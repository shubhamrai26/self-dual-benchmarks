module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 , y256 , y257 , y258 , y259 , y260 , y261 , y262 , y263 , y264 , y265 , y266 , y267 , y268 , y269 , y270 , y271 , y272 , y273 , y274 , y275 , y276 , y277 , y278 , y279 , y280 , y281 , y282 , y283 , y284 , y285 , y286 , y287 , y288 , y289 , y290 , y291 , y292 , y293 , y294 , y295 , y296 , y297 , y298 , y299 , y300 , y301 , y302 , y303 , y304 , y305 , y306 , y307 , y308 , y309 , y310 , y311 , y312 , y313 , y314 , y315 , y316 , y317 , y318 , y319 , y320 , y321 , y322 , y323 , y324 , y325 , y326 , y327 , y328 , y329 , y330 , y331 , y332 , y333 , y334 , y335 , y336 , y337 , y338 , y339 , y340 , y341 , y342 , y343 , y344 , y345 , y346 , y347 , y348 , y349 , y350 , y351 , y352 , y353 , y354 , y355 , y356 , y357 , y358 , y359 , y360 , y361 , y362 , y363 , y364 , y365 , y366 , y367 , y368 , y369 , y370 , y371 , y372 , y373 , y374 , y375 , y376 , y377 , y378 , y379 , y380 , y381 , y382 , y383 , y384 , y385 , y386 , y387 , y388 , y389 , y390 , y391 , y392 , y393 , y394 , y395 , y396 , y397 , y398 , y399 , y400 , y401 , y402 , y403 , y404 , y405 , y406 , y407 , y408 , y409 , y410 , y411 , y412 , y413 , y414 , y415 , y416 , y417 , y418 , y419 , y420 , y421 , y422 , y423 , y424 , y425 , y426 , y427 , y428 , y429 , y430 , y431 , y432 , y433 , y434 , y435 , y436 , y437 , y438 , y439 , y440 , y441 , y442 , y443 , y444 , y445 , y446 , y447 , y448 , y449 , y450 , y451 , y452 , y453 , y454 , y455 , y456 , y457 , y458 , y459 , y460 , y461 , y462 , y463 , y464 , y465 , y466 , y467 , y468 , y469 , y470 , y471 , y472 , y473 , y474 , y475 , y476 , y477 , y478 , y479 , y480 , y481 , y482 , y483 , y484 , y485 , y486 , y487 , y488 , y489 , y490 , y491 , y492 , y493 , y494 , y495 , y496 , y497 , y498 , y499 , y500 , y501 , y502 , y503 , y504 , y505 , y506 , y507 , y508 , y509 , y510 , y511 , y512 , y513 , y514 , y515 , y516 , y517 , y518 , y519 , y520 , y521 , y522 , y523 , y524 , y525 , y526 , y527 , y528 , y529 , y530 , y531 , y532 , y533 , y534 , y535 , y536 , y537 , y538 , y539 , y540 , y541 , y542 , y543 , y544 , y545 , y546 , y547 , y548 , y549 , y550 , y551 , y552 , y553 , y554 , y555 , y556 , y557 , y558 , y559 , y560 , y561 , y562 , y563 , y564 , y565 , y566 , y567 , y568 , y569 , y570 , y571 , y572 , y573 , y574 , y575 , y576 , y577 , y578 , y579 , y580 , y581 , y582 , y583 , y584 , y585 , y586 , y587 , y588 , y589 , y590 , y591 , y592 , y593 , y594 , y595 , y596 , y597 , y598 , y599 , y600 , y601 , y602 , y603 , y604 , y605 , y606 , y607 , y608 , y609 , y610 , y611 , y612 , y613 , y614 , y615 , y616 , y617 , y618 , y619 , y620 , y621 , y622 , y623 , y624 , y625 , y626 , y627 , y628 , y629 , y630 , y631 , y632 , y633 , y634 , y635 , y636 , y637 , y638 , y639 , y640 , y641 , y642 , y643 , y644 , y645 , y646 , y647 , y648 , y649 , y650 , y651 , y652 , y653 , y654 , y655 , y656 , y657 , y658 , y659 , y660 , y661 , y662 , y663 , y664 , y665 , y666 , y667 , y668 , y669 , y670 , y671 , y672 , y673 , y674 , y675 , y676 , y677 , y678 , y679 , y680 , y681 , y682 , y683 , y684 , y685 , y686 , y687 , y688 , y689 , y690 , y691 , y692 , y693 , y694 , y695 , y696 , y697 , y698 , y699 , y700 , y701 , y702 , y703 , y704 , y705 , y706 , y707 , y708 , y709 , y710 , y711 , y712 , y713 , y714 , y715 , y716 , y717 , y718 , y719 , y720 , y721 , y722 , y723 , y724 , y725 , y726 , y727 , y728 , y729 , y730 , y731 , y732 , y733 , y734 , y735 , y736 , y737 , y738 , y739 , y740 , y741 , y742 , y743 , y744 , y745 , y746 , y747 , y748 , y749 , y750 , y751 , y752 , y753 , y754 , y755 , y756 , y757 , y758 , y759 , y760 , y761 , y762 , y763 , y764 , y765 , y766 , y767 , y768 , y769 , y770 , y771 , y772 , y773 , y774 , y775 , y776 , y777 , y778 , y779 , y780 , y781 , y782 , y783 , y784 , y785 , y786 , y787 , y788 , y789 , y790 , y791 , y792 , y793 , y794 , y795 , y796 , y797 , y798 , y799 , y800 , y801 , y802 , y803 , y804 , y805 , y806 , y807 , y808 , y809 , y810 , y811 , y812 , y813 , y814 , y815 , y816 , y817 , y818 , y819 , y820 , y821 , y822 , y823 , y824 , y825 , y826 , y827 , y828 , y829 , y830 , y831 , y832 , y833 , y834 , y835 , y836 , y837 , y838 , y839 , y840 , y841 , y842 , y843 , y844 , y845 , y846 , y847 , y848 , y849 , y850 , y851 , y852 , y853 , y854 , y855 , y856 , y857 , y858 , y859 , y860 , y861 , y862 , y863 , y864 , y865 , y866 , y867 , y868 , y869 , y870 , y871 , y872 , y873 , y874 , y875 , y876 , y877 , y878 , y879 , y880 , y881 , y882 , y883 , y884 , y885 , y886 , y887 , y888 , y889 , y890 , y891 , y892 , y893 , y894 , y895 , y896 , y897 , y898 , y899 , y900 , y901 , y902 , y903 , y904 , y905 , y906 , y907 , y908 , y909 , y910 , y911 , y912 , y913 , y914 , y915 , y916 , y917 , y918 , y919 , y920 , y921 , y922 , y923 , y924 , y925 , y926 , y927 , y928 , y929 , y930 , y931 , y932 , y933 , y934 , y935 , y936 , y937 , y938 , y939 , y940 , y941 , y942 , y943 , y944 , y945 , y946 , y947 , y948 , y949 , y950 , y951 , y952 , y953 , y954 , y955 , y956 , y957 , y958 , y959 , y960 , y961 , y962 , y963 , y964 , y965 , y966 , y967 , y968 , y969 , y970 , y971 , y972 , y973 , y974 , y975 , y976 , y977 , y978 , y979 , y980 , y981 , y982 , y983 , y984 , y985 , y986 , y987 , y988 , y989 , y990 , y991 , y992 , y993 , y994 , y995 , y996 , y997 , y998 , y999 , y1000 , y1001 , y1002 , y1003 , y1004 , y1005 , y1006 , y1007 , y1008 , y1009 , y1010 , y1011 , y1012 , y1013 , y1014 , y1015 , y1016 , y1017 , y1018 , y1019 , y1020 , y1021 , y1022 , y1023 , y1024 , y1025 , y1026 , y1027 , y1028 , y1029 , y1030 , y1031 , y1032 , y1033 , y1034 , y1035 , y1036 , y1037 , y1038 , y1039 , y1040 , y1041 , y1042 , y1043 , y1044 , y1045 , y1046 , y1047 , y1048 , y1049 , y1050 , y1051 , y1052 , y1053 , y1054 , y1055 , y1056 , y1057 , y1058 , y1059 , y1060 , y1061 , y1062 , y1063 , y1064 , y1065 , y1066 , y1067 , y1068 , y1069 , y1070 , y1071 , y1072 , y1073 , y1074 , y1075 , y1076 , y1077 , y1078 , y1079 , y1080 , y1081 , y1082 , y1083 , y1084 , y1085 , y1086 , y1087 , y1088 , y1089 , y1090 , y1091 , y1092 , y1093 , y1094 , y1095 , y1096 , y1097 , y1098 , y1099 , y1100 , y1101 , y1102 , y1103 , y1104 , y1105 , y1106 , y1107 , y1108 , y1109 , y1110 , y1111 , y1112 , y1113 , y1114 , y1115 , y1116 , y1117 , y1118 , y1119 , y1120 , y1121 , y1122 , y1123 , y1124 , y1125 , y1126 , y1127 , y1128 , y1129 , y1130 , y1131 , y1132 , y1133 , y1134 , y1135 , y1136 , y1137 , y1138 , y1139 , y1140 , y1141 , y1142 , y1143 , y1144 , y1145 , y1146 , y1147 , y1148 , y1149 , y1150 , y1151 , y1152 , y1153 , y1154 , y1155 , y1156 , y1157 , y1158 , y1159 , y1160 , y1161 , y1162 , y1163 , y1164 , y1165 , y1166 , y1167 , y1168 , y1169 , y1170 , y1171 , y1172 , y1173 , y1174 , y1175 , y1176 , y1177 , y1178 , y1179 , y1180 , y1181 , y1182 , y1183 , y1184 , y1185 , y1186 , y1187 , y1188 , y1189 , y1190 , y1191 , y1192 , y1193 , y1194 , y1195 , y1196 , y1197 , y1198 , y1199 , y1200 , y1201 , y1202 , y1203 , y1204 , y1205 , y1206 , y1207 , y1208 , y1209 , y1210 , y1211 , y1212 , y1213 , y1214 , y1215 , y1216 , y1217 , y1218 , y1219 , y1220 , y1221 , y1222 , y1223 , y1224 , y1225 , y1226 , y1227 , y1228 , y1229 , y1230 , y1231 , y1232 , y1233 , y1234 , y1235 , y1236 , y1237 , y1238 , y1239 , y1240 , y1241 , y1242 , y1243 , y1244 , y1245 , y1246 , y1247 , y1248 , y1249 , y1250 , y1251 , y1252 , y1253 , y1254 , y1255 , y1256 , y1257 , y1258 , y1259 , y1260 , y1261 , y1262 , y1263 , y1264 , y1265 , y1266 , y1267 , y1268 , y1269 , y1270 , y1271 , y1272 , y1273 , y1274 , y1275 , y1276 , y1277 , y1278 , y1279 , y1280 , y1281 , y1282 , y1283 , y1284 , y1285 , y1286 , y1287 , y1288 , y1289 , y1290 , y1291 , y1292 , y1293 , y1294 , y1295 , y1296 , y1297 , y1298 , y1299 , y1300 , y1301 , y1302 , y1303 , y1304 , y1305 , y1306 , y1307 , y1308 , y1309 , y1310 , y1311 , y1312 , y1313 , y1314 , y1315 , y1316 , y1317 , y1318 , y1319 , y1320 , y1321 , y1322 , y1323 , y1324 , y1325 , y1326 , y1327 , y1328 , y1329 , y1330 , y1331 , y1332 , y1333 , y1334 , y1335 , y1336 , y1337 , y1338 , y1339 , y1340 , y1341 , y1342 , y1343 , y1344 , y1345 , y1346 , y1347 , y1348 , y1349 , y1350 , y1351 , y1352 , y1353 , y1354 , y1355 , y1356 , y1357 , y1358 , y1359 , y1360 , y1361 , y1362 , y1363 , y1364 , y1365 , y1366 , y1367 , y1368 , y1369 , y1370 , y1371 , y1372 , y1373 , y1374 , y1375 , y1376 , y1377 , y1378 , y1379 , y1380 , y1381 , y1382 , y1383 , y1384 , y1385 , y1386 , y1387 , y1388 , y1389 , y1390 , y1391 , y1392 , y1393 , y1394 , y1395 , y1396 , y1397 , y1398 , y1399 , y1400 , y1401 , y1402 , y1403 , y1404 , y1405 , y1406 , y1407 , y1408 , y1409 , y1410 , y1411 , y1412 , y1413 , y1414 , y1415 , y1416 , y1417 , y1418 , y1419 , y1420 , y1421 , y1422 , y1423 , y1424 , y1425 , y1426 , y1427 , y1428 , y1429 , y1430 , y1431 , y1432 , y1433 , y1434 , y1435 , y1436 , y1437 , y1438 , y1439 , y1440 , y1441 , y1442 , y1443 , y1444 , y1445 , y1446 , y1447 , y1448 , y1449 , y1450 , y1451 , y1452 , y1453 , y1454 , y1455 , y1456 , y1457 , y1458 , y1459 , y1460 , y1461 , y1462 , y1463 , y1464 , y1465 , y1466 , y1467 , y1468 , y1469 , y1470 , y1471 , y1472 , y1473 , y1474 , y1475 , y1476 , y1477 , y1478 , y1479 , y1480 , y1481 , y1482 , y1483 , y1484 , y1485 , y1486 , y1487 , y1488 , y1489 , y1490 , y1491 , y1492 , y1493 , y1494 , y1495 , y1496 , y1497 , y1498 , y1499 , y1500 , y1501 , y1502 , y1503 , y1504 , y1505 , y1506 , y1507 , y1508 , y1509 , y1510 , y1511 , y1512 , y1513 , y1514 , y1515 , y1516 , y1517 , y1518 , y1519 , y1520 , y1521 , y1522 , y1523 , y1524 , y1525 , y1526 , y1527 , y1528 , y1529 , y1530 , y1531 , y1532 , y1533 , y1534 , y1535 , y1536 , y1537 , y1538 , y1539 , y1540 , y1541 , y1542 , y1543 , y1544 , y1545 , y1546 , y1547 , y1548 , y1549 , y1550 , y1551 , y1552 , y1553 , y1554 , y1555 , y1556 , y1557 , y1558 , y1559 , y1560 , y1561 , y1562 , y1563 , y1564 , y1565 , y1566 , y1567 , y1568 , y1569 , y1570 , y1571 , y1572 , y1573 , y1574 , y1575 , y1576 , y1577 , y1578 , y1579 , y1580 , y1581 , y1582 , y1583 , y1584 , y1585 , y1586 , y1587 , y1588 , y1589 , y1590 , y1591 , y1592 , y1593 , y1594 , y1595 , y1596 , y1597 , y1598 , y1599 , y1600 , y1601 , y1602 , y1603 , y1604 , y1605 , y1606 , y1607 , y1608 , y1609 , y1610 , y1611 , y1612 , y1613 , y1614 , y1615 , y1616 , y1617 , y1618 , y1619 , y1620 , y1621 , y1622 , y1623 , y1624 , y1625 , y1626 , y1627 , y1628 , y1629 , y1630 , y1631 , y1632 , y1633 , y1634 , y1635 , y1636 , y1637 , y1638 , y1639 , y1640 , y1641 , y1642 , y1643 , y1644 , y1645 , y1646 , y1647 , y1648 , y1649 , y1650 , y1651 , y1652 , y1653 , y1654 , y1655 , y1656 , y1657 , y1658 , y1659 , y1660 , y1661 , y1662 , y1663 , y1664 , y1665 , y1666 , y1667 , y1668 , y1669 , y1670 , y1671 , y1672 , y1673 , y1674 , y1675 , y1676 , y1677 , y1678 , y1679 , y1680 , y1681 , y1682 , y1683 , y1684 , y1685 , y1686 , y1687 , y1688 , y1689 , y1690 , y1691 , y1692 , y1693 , y1694 , y1695 , y1696 , y1697 , y1698 , y1699 , y1700 , y1701 , y1702 , y1703 , y1704 , y1705 , y1706 , y1707 , y1708 , y1709 , y1710 , y1711 , y1712 , y1713 , y1714 , y1715 , y1716 , y1717 , y1718 , y1719 , y1720 , y1721 , y1722 , y1723 , y1724 , y1725 , y1726 , y1727 , y1728 , y1729 , y1730 , y1731 , y1732 , y1733 , y1734 , y1735 , y1736 , y1737 , y1738 , y1739 , y1740 , y1741 , y1742 , y1743 , y1744 , y1745 , y1746 , y1747 , y1748 , y1749 , y1750 , y1751 , y1752 , y1753 , y1754 , y1755 , y1756 , y1757 , y1758 , y1759 , y1760 , y1761 , y1762 , y1763 , y1764 , y1765 , y1766 , y1767 , y1768 , y1769 , y1770 , y1771 , y1772 , y1773 , y1774 , y1775 , y1776 , y1777 , y1778 , y1779 , y1780 , y1781 , y1782 , y1783 , y1784 , y1785 , y1786 , y1787 , y1788 , y1789 , y1790 , y1791 , y1792 , y1793 , y1794 , y1795 , y1796 , y1797 , y1798 , y1799 , y1800 , y1801 , y1802 , y1803 , y1804 , y1805 , y1806 , y1807 , y1808 , y1809 , y1810 , y1811 , y1812 , y1813 , y1814 , y1815 , y1816 , y1817 , y1818 , y1819 , y1820 , y1821 , y1822 , y1823 , y1824 , y1825 , y1826 , y1827 , y1828 , y1829 , y1830 , y1831 , y1832 , y1833 , y1834 , y1835 , y1836 , y1837 , y1838 , y1839 , y1840 , y1841 , y1842 , y1843 , y1844 , y1845 , y1846 , y1847 , y1848 , y1849 , y1850 , y1851 , y1852 , y1853 , y1854 , y1855 , y1856 , y1857 , y1858 , y1859 , y1860 , y1861 , y1862 , y1863 , y1864 , y1865 , y1866 , y1867 , y1868 , y1869 , y1870 , y1871 , y1872 , y1873 , y1874 , y1875 , y1876 , y1877 , y1878 , y1879 , y1880 , y1881 , y1882 , y1883 , y1884 , y1885 , y1886 , y1887 , y1888 , y1889 , y1890 , y1891 , y1892 , y1893 , y1894 , y1895 , y1896 , y1897 , y1898 , y1899 , y1900 , y1901 , y1902 , y1903 , y1904 , y1905 , y1906 , y1907 , y1908 , y1909 , y1910 , y1911 , y1912 , y1913 , y1914 , y1915 , y1916 , y1917 , y1918 , y1919 , y1920 , y1921 , y1922 , y1923 , y1924 , y1925 , y1926 , y1927 , y1928 , y1929 , y1930 , y1931 , y1932 , y1933 , y1934 , y1935 , y1936 , y1937 , y1938 , y1939 , y1940 , y1941 , y1942 , y1943 , y1944 , y1945 , y1946 , y1947 , y1948 , y1949 , y1950 , y1951 , y1952 , y1953 , y1954 , y1955 , y1956 , y1957 , y1958 , y1959 , y1960 , y1961 , y1962 , y1963 , y1964 , y1965 , y1966 , y1967 , y1968 , y1969 , y1970 , y1971 , y1972 , y1973 , y1974 , y1975 , y1976 , y1977 , y1978 , y1979 , y1980 , y1981 , y1982 , y1983 , y1984 , y1985 , y1986 , y1987 , y1988 , y1989 , y1990 , y1991 , y1992 , y1993 , y1994 , y1995 , y1996 , y1997 , y1998 , y1999 , y2000 , y2001 , y2002 , y2003 , y2004 , y2005 , y2006 , y2007 , y2008 , y2009 , y2010 , y2011 , y2012 , y2013 , y2014 , y2015 , y2016 , y2017 , y2018 , y2019 , y2020 , y2021 , y2022 , y2023 , y2024 , y2025 , y2026 , y2027 , y2028 , y2029 , y2030 , y2031 , y2032 , y2033 , y2034 , y2035 , y2036 , y2037 , y2038 , y2039 , y2040 , y2041 , y2042 , y2043 , y2044 , y2045 , y2046 , y2047 , y2048 , y2049 , y2050 , y2051 , y2052 , y2053 , y2054 , y2055 , y2056 , y2057 , y2058 , y2059 , y2060 , y2061 , y2062 , y2063 , y2064 , y2065 , y2066 , y2067 , y2068 , y2069 , y2070 , y2071 , y2072 , y2073 , y2074 , y2075 , y2076 , y2077 , y2078 , y2079 , y2080 , y2081 , y2082 , y2083 , y2084 , y2085 , y2086 , y2087 , y2088 , y2089 , y2090 , y2091 , y2092 , y2093 , y2094 , y2095 , y2096 , y2097 , y2098 , y2099 , y2100 , y2101 , y2102 , y2103 , y2104 , y2105 , y2106 , y2107 , y2108 , y2109 , y2110 , y2111 , y2112 , y2113 , y2114 , y2115 , y2116 , y2117 , y2118 , y2119 , y2120 , y2121 , y2122 , y2123 , y2124 , y2125 , y2126 , y2127 , y2128 , y2129 , y2130 , y2131 , y2132 , y2133 , y2134 , y2135 , y2136 , y2137 , y2138 , y2139 , y2140 , y2141 , y2142 , y2143 , y2144 , y2145 , y2146 , y2147 , y2148 , y2149 , y2150 , y2151 , y2152 , y2153 , y2154 , y2155 , y2156 , y2157 , y2158 , y2159 , y2160 , y2161 , y2162 , y2163 , y2164 , y2165 , y2166 , y2167 , y2168 , y2169 , y2170 , y2171 , y2172 , y2173 , y2174 , y2175 , y2176 , y2177 , y2178 , y2179 , y2180 , y2181 , y2182 , y2183 , y2184 , y2185 , y2186 , y2187 , y2188 , y2189 , y2190 , y2191 , y2192 , y2193 , y2194 , y2195 , y2196 , y2197 , y2198 , y2199 , y2200 , y2201 , y2202 , y2203 , y2204 , y2205 , y2206 , y2207 , y2208 , y2209 , y2210 , y2211 , y2212 , y2213 , y2214 , y2215 , y2216 , y2217 , y2218 , y2219 , y2220 , y2221 , y2222 , y2223 , y2224 , y2225 , y2226 , y2227 , y2228 , y2229 , y2230 , y2231 , y2232 , y2233 , y2234 , y2235 , y2236 , y2237 , y2238 , y2239 , y2240 , y2241 , y2242 , y2243 , y2244 , y2245 , y2246 , y2247 , y2248 , y2249 , y2250 , y2251 , y2252 , y2253 , y2254 , y2255 , y2256 , y2257 , y2258 , y2259 , y2260 , y2261 , y2262 , y2263 , y2264 , y2265 , y2266 , y2267 , y2268 , y2269 , y2270 , y2271 , y2272 , y2273 , y2274 , y2275 , y2276 , y2277 , y2278 , y2279 , y2280 , y2281 , y2282 , y2283 , y2284 , y2285 , y2286 , y2287 , y2288 , y2289 , y2290 , y2291 , y2292 , y2293 , y2294 , y2295 , y2296 , y2297 , y2298 , y2299 , y2300 , y2301 , y2302 , y2303 , y2304 , y2305 , y2306 , y2307 , y2308 , y2309 , y2310 , y2311 , y2312 , y2313 , y2314 , y2315 , y2316 , y2317 , y2318 , y2319 , y2320 , y2321 , y2322 , y2323 , y2324 , y2325 , y2326 , y2327 , y2328 , y2329 , y2330 , y2331 , y2332 , y2333 , y2334 , y2335 , y2336 , y2337 , y2338 , y2339 , y2340 , y2341 , y2342 , y2343 , y2344 , y2345 , y2346 , y2347 , y2348 , y2349 , y2350 , y2351 , y2352 , y2353 , y2354 , y2355 , y2356 , y2357 , y2358 , y2359 , y2360 , y2361 , y2362 , y2363 , y2364 , y2365 , y2366 , y2367 , y2368 , y2369 , y2370 , y2371 , y2372 , y2373 , y2374 , y2375 , y2376 , y2377 , y2378 , y2379 , y2380 , y2381 , y2382 , y2383 , y2384 , y2385 , y2386 , y2387 , y2388 , y2389 , y2390 , y2391 , y2392 , y2393 , y2394 , y2395 , y2396 , y2397 , y2398 , y2399 , y2400 , y2401 , y2402 , y2403 , y2404 , y2405 , y2406 , y2407 , y2408 , y2409 , y2410 , y2411 , y2412 , y2413 , y2414 , y2415 , y2416 , y2417 , y2418 , y2419 , y2420 , y2421 , y2422 , y2423 , y2424 , y2425 , y2426 , y2427 , y2428 , y2429 , y2430 , y2431 , y2432 , y2433 , y2434 , y2435 , y2436 , y2437 , y2438 , y2439 , y2440 , y2441 , y2442 , y2443 , y2444 , y2445 , y2446 , y2447 , y2448 , y2449 , y2450 , y2451 , y2452 , y2453 , y2454 , y2455 , y2456 , y2457 , y2458 , y2459 , y2460 , y2461 , y2462 , y2463 , y2464 , y2465 , y2466 , y2467 , y2468 , y2469 , y2470 , y2471 , y2472 , y2473 , y2474 , y2475 , y2476 , y2477 , y2478 , y2479 , y2480 , y2481 , y2482 , y2483 , y2484 , y2485 , y2486 , y2487 , y2488 , y2489 , y2490 , y2491 , y2492 , y2493 , y2494 , y2495 , y2496 , y2497 , y2498 , y2499 , y2500 , y2501 , y2502 , y2503 , y2504 , y2505 , y2506 , y2507 , y2508 , y2509 , y2510 , y2511 , y2512 , y2513 , y2514 , y2515 , y2516 , y2517 , y2518 , y2519 , y2520 , y2521 , y2522 , y2523 , y2524 , y2525 , y2526 , y2527 , y2528 , y2529 , y2530 , y2531 , y2532 , y2533 , y2534 , y2535 , y2536 , y2537 , y2538 , y2539 , y2540 , y2541 , y2542 , y2543 , y2544 , y2545 , y2546 , y2547 , y2548 , y2549 , y2550 , y2551 , y2552 , y2553 , y2554 , y2555 , y2556 , y2557 , y2558 , y2559 , y2560 , y2561 , y2562 , y2563 , y2564 , y2565 , y2566 , y2567 , y2568 , y2569 , y2570 , y2571 , y2572 , y2573 , y2574 , y2575 , y2576 , y2577 , y2578 , y2579 , y2580 , y2581 , y2582 , y2583 , y2584 , y2585 , y2586 , y2587 , y2588 , y2589 , y2590 , y2591 , y2592 , y2593 , y2594 , y2595 , y2596 , y2597 , y2598 , y2599 , y2600 , y2601 , y2602 , y2603 , y2604 , y2605 , y2606 , y2607 , y2608 , y2609 , y2610 , y2611 , y2612 , y2613 , y2614 , y2615 , y2616 , y2617 , y2618 , y2619 , y2620 , y2621 , y2622 , y2623 , y2624 , y2625 , y2626 , y2627 , y2628 , y2629 , y2630 , y2631 , y2632 , y2633 , y2634 , y2635 , y2636 , y2637 , y2638 , y2639 , y2640 , y2641 , y2642 , y2643 , y2644 , y2645 , y2646 , y2647 , y2648 , y2649 , y2650 , y2651 , y2652 , y2653 , y2654 , y2655 , y2656 , y2657 , y2658 , y2659 , y2660 , y2661 , y2662 , y2663 , y2664 , y2665 , y2666 , y2667 , y2668 , y2669 , y2670 , y2671 , y2672 , y2673 , y2674 , y2675 , y2676 , y2677 , y2678 , y2679 , y2680 , y2681 , y2682 , y2683 , y2684 , y2685 , y2686 , y2687 , y2688 , y2689 , y2690 , y2691 , y2692 , y2693 , y2694 , y2695 , y2696 , y2697 , y2698 , y2699 , y2700 , y2701 , y2702 , y2703 , y2704 , y2705 , y2706 , y2707 , y2708 , y2709 , y2710 , y2711 , y2712 , y2713 , y2714 , y2715 , y2716 , y2717 , y2718 , y2719 , y2720 , y2721 , y2722 , y2723 , y2724 , y2725 , y2726 , y2727 , y2728 , y2729 , y2730 , y2731 , y2732 , y2733 , y2734 , y2735 , y2736 , y2737 , y2738 , y2739 , y2740 , y2741 , y2742 , y2743 , y2744 , y2745 , y2746 , y2747 , y2748 , y2749 , y2750 , y2751 , y2752 , y2753 , y2754 , y2755 , y2756 , y2757 , y2758 , y2759 , y2760 , y2761 , y2762 , y2763 , y2764 , y2765 , y2766 , y2767 , y2768 , y2769 , y2770 , y2771 , y2772 , y2773 , y2774 , y2775 , y2776 , y2777 , y2778 , y2779 , y2780 , y2781 , y2782 , y2783 , y2784 , y2785 , y2786 , y2787 , y2788 , y2789 , y2790 , y2791 , y2792 , y2793 , y2794 , y2795 , y2796 , y2797 , y2798 , y2799 , y2800 , y2801 , y2802 , y2803 , y2804 , y2805 , y2806 , y2807 , y2808 , y2809 , y2810 , y2811 , y2812 , y2813 , y2814 , y2815 , y2816 , y2817 , y2818 , y2819 , y2820 , y2821 , y2822 , y2823 , y2824 , y2825 , y2826 , y2827 , y2828 , y2829 , y2830 , y2831 , y2832 , y2833 , y2834 , y2835 , y2836 , y2837 , y2838 , y2839 , y2840 , y2841 , y2842 , y2843 , y2844 , y2845 , y2846 , y2847 , y2848 , y2849 , y2850 , y2851 , y2852 , y2853 , y2854 , y2855 , y2856 , y2857 , y2858 , y2859 , y2860 , y2861 , y2862 , y2863 , y2864 , y2865 , y2866 , y2867 , y2868 , y2869 , y2870 , y2871 , y2872 , y2873 , y2874 , y2875 , y2876 , y2877 , y2878 , y2879 , y2880 , y2881 , y2882 , y2883 , y2884 , y2885 , y2886 , y2887 , y2888 , y2889 , y2890 , y2891 , y2892 , y2893 , y2894 , y2895 , y2896 , y2897 , y2898 , y2899 , y2900 , y2901 , y2902 , y2903 , y2904 , y2905 , y2906 , y2907 , y2908 , y2909 , y2910 , y2911 , y2912 , y2913 , y2914 , y2915 , y2916 , y2917 , y2918 , y2919 , y2920 , y2921 , y2922 , y2923 , y2924 , y2925 , y2926 , y2927 , y2928 , y2929 , y2930 , y2931 , y2932 , y2933 , y2934 , y2935 , y2936 , y2937 , y2938 , y2939 , y2940 , y2941 , y2942 , y2943 , y2944 , y2945 , y2946 , y2947 , y2948 , y2949 , y2950 , y2951 , y2952 , y2953 , y2954 , y2955 , y2956 , y2957 , y2958 , y2959 , y2960 , y2961 , y2962 , y2963 , y2964 , y2965 , y2966 , y2967 , y2968 , y2969 , y2970 , y2971 , y2972 , y2973 , y2974 , y2975 , y2976 , y2977 , y2978 , y2979 , y2980 , y2981 , y2982 , y2983 , y2984 , y2985 , y2986 , y2987 , y2988 , y2989 , y2990 , y2991 , y2992 , y2993 , y2994 , y2995 , y2996 , y2997 , y2998 , y2999 , y3000 , y3001 , y3002 , y3003 , y3004 , y3005 , y3006 , y3007 , y3008 , y3009 , y3010 , y3011 , y3012 , y3013 , y3014 , y3015 , y3016 , y3017 , y3018 , y3019 , y3020 , y3021 , y3022 , y3023 , y3024 , y3025 , y3026 , y3027 , y3028 , y3029 , y3030 , y3031 , y3032 , y3033 , y3034 , y3035 , y3036 , y3037 , y3038 , y3039 , y3040 , y3041 , y3042 , y3043 , y3044 , y3045 , y3046 , y3047 , y3048 , y3049 , y3050 , y3051 , y3052 , y3053 , y3054 , y3055 , y3056 , y3057 , y3058 , y3059 , y3060 , y3061 , y3062 , y3063 , y3064 , y3065 , y3066 , y3067 , y3068 , y3069 , y3070 , y3071 , y3072 , y3073 , y3074 , y3075 , y3076 , y3077 , y3078 , y3079 , y3080 , y3081 , y3082 , y3083 , y3084 , y3085 , y3086 , y3087 , y3088 , y3089 , y3090 , y3091 , y3092 , y3093 , y3094 , y3095 , y3096 , y3097 , y3098 , y3099 , y3100 , y3101 , y3102 , y3103 , y3104 , y3105 , y3106 , y3107 , y3108 , y3109 , y3110 , y3111 , y3112 , y3113 , y3114 , y3115 , y3116 , y3117 , y3118 , y3119 , y3120 , y3121 , y3122 , y3123 , y3124 , y3125 , y3126 , y3127 , y3128 , y3129 , y3130 , y3131 , y3132 , y3133 , y3134 , y3135 , y3136 , y3137 , y3138 , y3139 , y3140 , y3141 , y3142 , y3143 , y3144 , y3145 , y3146 , y3147 , y3148 , y3149 , y3150 , y3151 , y3152 , y3153 , y3154 , y3155 , y3156 , y3157 , y3158 , y3159 , y3160 , y3161 , y3162 , y3163 , y3164 , y3165 , y3166 , y3167 , y3168 , y3169 , y3170 , y3171 , y3172 , y3173 , y3174 , y3175 , y3176 , y3177 , y3178 , y3179 , y3180 , y3181 , y3182 , y3183 , y3184 , y3185 , y3186 , y3187 , y3188 , y3189 , y3190 , y3191 , y3192 , y3193 , y3194 , y3195 , y3196 , y3197 , y3198 , y3199 , y3200 , y3201 , y3202 , y3203 , y3204 , y3205 , y3206 , y3207 , y3208 , y3209 , y3210 , y3211 , y3212 , y3213 , y3214 , y3215 , y3216 , y3217 , y3218 , y3219 , y3220 , y3221 , y3222 , y3223 , y3224 , y3225 , y3226 , y3227 , y3228 , y3229 , y3230 , y3231 , y3232 , y3233 , y3234 , y3235 , y3236 , y3237 , y3238 , y3239 , y3240 , y3241 , y3242 , y3243 , y3244 , y3245 , y3246 , y3247 , y3248 , y3249 , y3250 , y3251 , y3252 , y3253 , y3254 , y3255 , y3256 , y3257 , y3258 , y3259 , y3260 , y3261 , y3262 , y3263 , y3264 , y3265 , y3266 , y3267 , y3268 , y3269 , y3270 , y3271 , y3272 , y3273 , y3274 , y3275 , y3276 , y3277 , y3278 , y3279 , y3280 , y3281 , y3282 , y3283 , y3284 , y3285 , y3286 , y3287 , y3288 , y3289 , y3290 , y3291 , y3292 , y3293 , y3294 , y3295 , y3296 , y3297 , y3298 , y3299 , y3300 , y3301 , y3302 , y3303 , y3304 , y3305 , y3306 , y3307 , y3308 , y3309 , y3310 , y3311 , y3312 , y3313 , y3314 , y3315 , y3316 , y3317 , y3318 , y3319 , y3320 , y3321 , y3322 , y3323 , y3324 , y3325 , y3326 , y3327 , y3328 , y3329 , y3330 , y3331 , y3332 , y3333 , y3334 , y3335 , y3336 , y3337 , y3338 , y3339 , y3340 , y3341 , y3342 , y3343 , y3344 , y3345 , y3346 , y3347 , y3348 , y3349 , y3350 , y3351 , y3352 , y3353 , y3354 , y3355 , y3356 , y3357 , y3358 , y3359 , y3360 , y3361 , y3362 , y3363 , y3364 , y3365 , y3366 , y3367 , y3368 , y3369 , y3370 , y3371 , y3372 , y3373 , y3374 , y3375 , y3376 , y3377 , y3378 , y3379 , y3380 , y3381 , y3382 , y3383 , y3384 , y3385 , y3386 , y3387 , y3388 , y3389 , y3390 , y3391 , y3392 , y3393 , y3394 , y3395 , y3396 , y3397 , y3398 , y3399 , y3400 , y3401 , y3402 , y3403 , y3404 , y3405 , y3406 , y3407 , y3408 , y3409 , y3410 , y3411 , y3412 , y3413 , y3414 , y3415 , y3416 , y3417 , y3418 , y3419 , y3420 , y3421 , y3422 , y3423 , y3424 , y3425 , y3426 , y3427 , y3428 , y3429 , y3430 , y3431 , y3432 , y3433 , y3434 , y3435 , y3436 , y3437 , y3438 , y3439 , y3440 , y3441 , y3442 , y3443 , y3444 , y3445 , y3446 , y3447 , y3448 , y3449 , y3450 , y3451 , y3452 , y3453 , y3454 , y3455 , y3456 , y3457 , y3458 , y3459 , y3460 , y3461 , y3462 , y3463 , y3464 , y3465 , y3466 , y3467 , y3468 , y3469 , y3470 , y3471 , y3472 , y3473 , y3474 , y3475 , y3476 , y3477 , y3478 , y3479 , y3480 , y3481 , y3482 , y3483 , y3484 , y3485 , y3486 , y3487 , y3488 , y3489 , y3490 , y3491 , y3492 , y3493 , y3494 , y3495 , y3496 , y3497 , y3498 , y3499 , y3500 , y3501 , y3502 , y3503 , y3504 , y3505 , y3506 , y3507 , y3508 , y3509 , y3510 , y3511 , y3512 , y3513 , y3514 , y3515 , y3516 , y3517 , y3518 , y3519 , y3520 , y3521 , y3522 , y3523 , y3524 , y3525 , y3526 , y3527 , y3528 , y3529 , y3530 , y3531 , y3532 , y3533 , y3534 , y3535 , y3536 , y3537 , y3538 , y3539 , y3540 , y3541 , y3542 , y3543 , y3544 , y3545 , y3546 , y3547 , y3548 , y3549 , y3550 , y3551 , y3552 , y3553 , y3554 , y3555 , y3556 , y3557 , y3558 , y3559 , y3560 , y3561 , y3562 , y3563 , y3564 , y3565 , y3566 , y3567 , y3568 , y3569 , y3570 , y3571 , y3572 , y3573 , y3574 , y3575 , y3576 , y3577 , y3578 , y3579 , y3580 , y3581 , y3582 , y3583 , y3584 , y3585 , y3586 , y3587 , y3588 , y3589 , y3590 , y3591 , y3592 , y3593 , y3594 , y3595 , y3596 , y3597 , y3598 , y3599 , y3600 , y3601 , y3602 , y3603 , y3604 , y3605 , y3606 , y3607 , y3608 , y3609 , y3610 , y3611 , y3612 , y3613 , y3614 , y3615 , y3616 , y3617 , y3618 , y3619 , y3620 , y3621 , y3622 , y3623 , y3624 , y3625 , y3626 , y3627 , y3628 , y3629 , y3630 , y3631 , y3632 , y3633 , y3634 , y3635 , y3636 , y3637 , y3638 , y3639 , y3640 , y3641 , y3642 , y3643 , y3644 , y3645 , y3646 , y3647 , y3648 , y3649 , y3650 , y3651 , y3652 , y3653 , y3654 , y3655 , y3656 , y3657 , y3658 , y3659 , y3660 , y3661 , y3662 , y3663 , y3664 , y3665 , y3666 , y3667 , y3668 , y3669 , y3670 , y3671 , y3672 , y3673 , y3674 , y3675 , y3676 , y3677 , y3678 , y3679 , y3680 , y3681 , y3682 , y3683 , y3684 , y3685 , y3686 , y3687 , y3688 , y3689 , y3690 , y3691 , y3692 , y3693 , y3694 , y3695 , y3696 , y3697 , y3698 , y3699 , y3700 , y3701 , y3702 , y3703 , y3704 , y3705 , y3706 , y3707 , y3708 , y3709 , y3710 , y3711 , y3712 , y3713 , y3714 , y3715 , y3716 , y3717 , y3718 , y3719 , y3720 , y3721 , y3722 , y3723 , y3724 , y3725 , y3726 , y3727 , y3728 , y3729 , y3730 , y3731 , y3732 , y3733 , y3734 , y3735 , y3736 , y3737 , y3738 , y3739 , y3740 , y3741 , y3742 , y3743 , y3744 , y3745 , y3746 , y3747 , y3748 , y3749 , y3750 , y3751 , y3752 , y3753 , y3754 , y3755 , y3756 , y3757 , y3758 , y3759 , y3760 , y3761 , y3762 , y3763 , y3764 , y3765 , y3766 , y3767 , y3768 , y3769 , y3770 , y3771 , y3772 , y3773 , y3774 , y3775 , y3776 , y3777 , y3778 , y3779 , y3780 , y3781 , y3782 , y3783 , y3784 , y3785 , y3786 , y3787 , y3788 , y3789 , y3790 , y3791 , y3792 , y3793 , y3794 , y3795 , y3796 , y3797 , y3798 , y3799 , y3800 , y3801 , y3802 , y3803 , y3804 , y3805 , y3806 , y3807 , y3808 , y3809 , y3810 , y3811 , y3812 , y3813 , y3814 , y3815 , y3816 , y3817 , y3818 , y3819 , y3820 , y3821 , y3822 , y3823 , y3824 , y3825 , y3826 , y3827 , y3828 , y3829 , y3830 , y3831 , y3832 , y3833 , y3834 , y3835 , y3836 , y3837 , y3838 , y3839 , y3840 , y3841 , y3842 , y3843 , y3844 , y3845 , y3846 , y3847 , y3848 , y3849 , y3850 , y3851 , y3852 , y3853 , y3854 , y3855 , y3856 , y3857 , y3858 , y3859 , y3860 , y3861 , y3862 , y3863 , y3864 , y3865 , y3866 , y3867 , y3868 , y3869 , y3870 , y3871 , y3872 , y3873 , y3874 , y3875 , y3876 , y3877 , y3878 , y3879 , y3880 , y3881 , y3882 , y3883 , y3884 , y3885 , y3886 , y3887 , y3888 , y3889 , y3890 , y3891 , y3892 , y3893 , y3894 , y3895 , y3896 , y3897 , y3898 , y3899 , y3900 , y3901 , y3902 , y3903 , y3904 , y3905 , y3906 , y3907 , y3908 , y3909 , y3910 , y3911 , y3912 , y3913 , y3914 , y3915 , y3916 , y3917 , y3918 , y3919 , y3920 , y3921 , y3922 , y3923 , y3924 , y3925 , y3926 , y3927 , y3928 , y3929 , y3930 , y3931 , y3932 , y3933 , y3934 , y3935 , y3936 , y3937 , y3938 , y3939 , y3940 , y3941 , y3942 , y3943 , y3944 , y3945 , y3946 , y3947 , y3948 , y3949 , y3950 , y3951 , y3952 , y3953 , y3954 , y3955 , y3956 , y3957 , y3958 , y3959 , y3960 , y3961 , y3962 , y3963 , y3964 , y3965 , y3966 , y3967 , y3968 , y3969 , y3970 , y3971 , y3972 , y3973 , y3974 , y3975 , y3976 , y3977 , y3978 , y3979 , y3980 , y3981 , y3982 , y3983 , y3984 , y3985 , y3986 , y3987 , y3988 , y3989 , y3990 , y3991 , y3992 , y3993 , y3994 , y3995 , y3996 , y3997 , y3998 , y3999 , y4000 , y4001 , y4002 , y4003 , y4004 , y4005 , y4006 , y4007 , y4008 , y4009 , y4010 , y4011 , y4012 , y4013 , y4014 , y4015 , y4016 , y4017 , y4018 , y4019 , y4020 , y4021 , y4022 , y4023 , y4024 , y4025 , y4026 , y4027 , y4028 , y4029 , y4030 , y4031 , y4032 , y4033 , y4034 , y4035 , y4036 , y4037 , y4038 , y4039 , y4040 , y4041 , y4042 , y4043 , y4044 , y4045 , y4046 , y4047 , y4048 , y4049 , y4050 , y4051 , y4052 , y4053 , y4054 , y4055 , y4056 , y4057 , y4058 , y4059 , y4060 , y4061 , y4062 , y4063 , y4064 , y4065 , y4066 , y4067 , y4068 , y4069 , y4070 , y4071 , y4072 , y4073 , y4074 , y4075 , y4076 , y4077 , y4078 , y4079 , y4080 , y4081 , y4082 , y4083 , y4084 , y4085 , y4086 , y4087 , y4088 , y4089 , y4090 , y4091 , y4092 , y4093 , y4094 , y4095 , y4096 , y4097 , y4098 , y4099 , y4100 , y4101 , y4102 , y4103 , y4104 , y4105 , y4106 , y4107 , y4108 , y4109 , y4110 , y4111 , y4112 , y4113 , y4114 , y4115 , y4116 , y4117 , y4118 , y4119 , y4120 , y4121 , y4122 , y4123 , y4124 , y4125 , y4126 , y4127 , y4128 , y4129 , y4130 , y4131 , y4132 , y4133 , y4134 , y4135 , y4136 , y4137 , y4138 , y4139 , y4140 , y4141 , y4142 , y4143 , y4144 , y4145 , y4146 , y4147 , y4148 , y4149 , y4150 , y4151 , y4152 , y4153 , y4154 , y4155 , y4156 , y4157 , y4158 , y4159 , y4160 , y4161 , y4162 , y4163 , y4164 , y4165 , y4166 , y4167 , y4168 , y4169 , y4170 , y4171 , y4172 , y4173 , y4174 , y4175 , y4176 , y4177 , y4178 , y4179 , y4180 , y4181 , y4182 , y4183 , y4184 , y4185 , y4186 , y4187 , y4188 , y4189 , y4190 , y4191 , y4192 , y4193 , y4194 , y4195 , y4196 , y4197 , y4198 , y4199 , y4200 , y4201 , y4202 , y4203 , y4204 , y4205 , y4206 , y4207 , y4208 , y4209 , y4210 , y4211 , y4212 , y4213 , y4214 , y4215 , y4216 , y4217 , y4218 , y4219 , y4220 , y4221 , y4222 , y4223 , y4224 , y4225 , y4226 , y4227 , y4228 , y4229 , y4230 , y4231 , y4232 , y4233 , y4234 , y4235 , y4236 , y4237 , y4238 , y4239 , y4240 , y4241 , y4242 , y4243 , y4244 , y4245 , y4246 , y4247 , y4248 , y4249 , y4250 , y4251 , y4252 , y4253 , y4254 , y4255 , y4256 , y4257 , y4258 , y4259 , y4260 , y4261 , y4262 , y4263 , y4264 , y4265 , y4266 , y4267 , y4268 , y4269 , y4270 , y4271 , y4272 , y4273 , y4274 , y4275 , y4276 , y4277 , y4278 , y4279 , y4280 , y4281 , y4282 , y4283 , y4284 , y4285 , y4286 , y4287 , y4288 , y4289 , y4290 , y4291 , y4292 , y4293 , y4294 , y4295 , y4296 , y4297 , y4298 , y4299 , y4300 , y4301 , y4302 , y4303 , y4304 , y4305 , y4306 , y4307 , y4308 , y4309 , y4310 , y4311 , y4312 , y4313 , y4314 , y4315 , y4316 , y4317 , y4318 , y4319 , y4320 , y4321 , y4322 , y4323 , y4324 , y4325 , y4326 , y4327 , y4328 , y4329 , y4330 , y4331 , y4332 , y4333 , y4334 , y4335 , y4336 , y4337 , y4338 , y4339 , y4340 , y4341 , y4342 , y4343 , y4344 , y4345 , y4346 , y4347 , y4348 , y4349 , y4350 , y4351 , y4352 , y4353 , y4354 , y4355 , y4356 , y4357 , y4358 , y4359 , y4360 , y4361 , y4362 , y4363 , y4364 , y4365 , y4366 , y4367 , y4368 , y4369 , y4370 , y4371 , y4372 , y4373 , y4374 , y4375 , y4376 , y4377 , y4378 , y4379 , y4380 , y4381 , y4382 , y4383 , y4384 , y4385 , y4386 , y4387 , y4388 , y4389 , y4390 , y4391 , y4392 , y4393 , y4394 , y4395 , y4396 , y4397 , y4398 , y4399 , y4400 , y4401 , y4402 , y4403 , y4404 , y4405 , y4406 , y4407 , y4408 , y4409 , y4410 , y4411 , y4412 , y4413 , y4414 , y4415 , y4416 , y4417 , y4418 , y4419 , y4420 , y4421 , y4422 , y4423 , y4424 , y4425 , y4426 , y4427 , y4428 , y4429 , y4430 , y4431 , y4432 , y4433 , y4434 , y4435 , y4436 , y4437 , y4438 , y4439 , y4440 , y4441 , y4442 , y4443 , y4444 , y4445 , y4446 , y4447 , y4448 , y4449 , y4450 , y4451 , y4452 , y4453 , y4454 , y4455 , y4456 , y4457 , y4458 , y4459 , y4460 , y4461 , y4462 , y4463 , y4464 , y4465 , y4466 , y4467 , y4468 , y4469 , y4470 , y4471 , y4472 , y4473 , y4474 , y4475 , y4476 , y4477 , y4478 , y4479 , y4480 , y4481 , y4482 , y4483 , y4484 , y4485 , y4486 , y4487 , y4488 , y4489 , y4490 , y4491 , y4492 , y4493 , y4494 , y4495 , y4496 , y4497 , y4498 , y4499 , y4500 , y4501 , y4502 , y4503 , y4504 , y4505 , y4506 , y4507 , y4508 , y4509 , y4510 , y4511 , y4512 , y4513 , y4514 , y4515 , y4516 , y4517 , y4518 , y4519 , y4520 , y4521 , y4522 , y4523 , y4524 , y4525 , y4526 , y4527 , y4528 , y4529 , y4530 , y4531 , y4532 , y4533 , y4534 , y4535 , y4536 , y4537 , y4538 , y4539 , y4540 , y4541 , y4542 , y4543 , y4544 , y4545 , y4546 , y4547 , y4548 , y4549 , y4550 , y4551 , y4552 , y4553 , y4554 , y4555 , y4556 , y4557 , y4558 , y4559 , y4560 , y4561 , y4562 , y4563 , y4564 , y4565 , y4566 , y4567 , y4568 , y4569 , y4570 , y4571 , y4572 , y4573 , y4574 , y4575 , y4576 , y4577 , y4578 , y4579 , y4580 , y4581 , y4582 , y4583 , y4584 , y4585 , y4586 , y4587 , y4588 , y4589 , y4590 , y4591 , y4592 , y4593 , y4594 , y4595 , y4596 , y4597 , y4598 , y4599 , y4600 , y4601 , y4602 , y4603 , y4604 , y4605 , y4606 , y4607 , y4608 , y4609 , y4610 , y4611 , y4612 , y4613 , y4614 , y4615 , y4616 , y4617 , y4618 , y4619 , y4620 , y4621 , y4622 , y4623 , y4624 , y4625 , y4626 , y4627 , y4628 , y4629 , y4630 , y4631 , y4632 , y4633 , y4634 , y4635 , y4636 , y4637 , y4638 , y4639 , y4640 , y4641 , y4642 , y4643 , y4644 , y4645 , y4646 , y4647 , y4648 , y4649 , y4650 , y4651 , y4652 , y4653 , y4654 , y4655 , y4656 , y4657 , y4658 , y4659 , y4660 , y4661 , y4662 , y4663 , y4664 , y4665 , y4666 , y4667 , y4668 , y4669 , y4670 , y4671 , y4672 , y4673 , y4674 , y4675 , y4676 , y4677 , y4678 , y4679 , y4680 , y4681 , y4682 , y4683 , y4684 , y4685 , y4686 , y4687 , y4688 , y4689 , y4690 , y4691 , y4692 , y4693 , y4694 , y4695 , y4696 , y4697 , y4698 , y4699 , y4700 , y4701 , y4702 , y4703 , y4704 , y4705 , y4706 , y4707 , y4708 , y4709 , y4710 , y4711 , y4712 , y4713 , y4714 , y4715 , y4716 , y4717 , y4718 , y4719 , y4720 , y4721 , y4722 , y4723 , y4724 , y4725 , y4726 , y4727 , y4728 , y4729 , y4730 , y4731 , y4732 , y4733 , y4734 , y4735 , y4736 , y4737 , y4738 , y4739 , y4740 , y4741 , y4742 , y4743 , y4744 , y4745 , y4746 , y4747 , y4748 , y4749 , y4750 , y4751 , y4752 , y4753 , y4754 , y4755 , y4756 , y4757 , y4758 , y4759 , y4760 , y4761 , y4762 , y4763 , y4764 , y4765 , y4766 , y4767 , y4768 , y4769 , y4770 , y4771 , y4772 , y4773 , y4774 , y4775 , y4776 , y4777 , y4778 , y4779 , y4780 , y4781 , y4782 , y4783 , y4784 , y4785 , y4786 , y4787 , y4788 , y4789 , y4790 , y4791 , y4792 , y4793 , y4794 , y4795 , y4796 , y4797 , y4798 , y4799 , y4800 , y4801 , y4802 , y4803 , y4804 , y4805 , y4806 , y4807 , y4808 , y4809 , y4810 , y4811 , y4812 , y4813 , y4814 , y4815 , y4816 , y4817 , y4818 , y4819 , y4820 , y4821 , y4822 , y4823 , y4824 , y4825 , y4826 , y4827 , y4828 , y4829 , y4830 , y4831 , y4832 , y4833 , y4834 , y4835 , y4836 , y4837 , y4838 , y4839 , y4840 , y4841 , y4842 , y4843 , y4844 , y4845 , y4846 , y4847 , y4848 , y4849 , y4850 , y4851 , y4852 , y4853 , y4854 , y4855 , y4856 , y4857 , y4858 , y4859 , y4860 , y4861 , y4862 , y4863 , y4864 , y4865 , y4866 , y4867 , y4868 , y4869 , y4870 , y4871 , y4872 , y4873 , y4874 , y4875 , y4876 , y4877 , y4878 , y4879 , y4880 , y4881 , y4882 , y4883 , y4884 , y4885 , y4886 , y4887 , y4888 , y4889 , y4890 , y4891 , y4892 , y4893 , y4894 , y4895 , y4896 , y4897 , y4898 , y4899 , y4900 , y4901 , y4902 , y4903 , y4904 , y4905 , y4906 , y4907 , y4908 , y4909 , y4910 , y4911 , y4912 , y4913 , y4914 , y4915 , y4916 , y4917 , y4918 , y4919 , y4920 , y4921 , y4922 , y4923 , y4924 , y4925 , y4926 , y4927 , y4928 , y4929 , y4930 , y4931 , y4932 , y4933 , y4934 , y4935 , y4936 , y4937 , y4938 , y4939 , y4940 , y4941 , y4942 , y4943 , y4944 , y4945 , y4946 , y4947 , y4948 , y4949 , y4950 , y4951 , y4952 , y4953 , y4954 , y4955 , y4956 , y4957 , y4958 , y4959 , y4960 , y4961 , y4962 , y4963 , y4964 , y4965 , y4966 , y4967 , y4968 , y4969 , y4970 , y4971 , y4972 , y4973 , y4974 , y4975 , y4976 , y4977 , y4978 , y4979 , y4980 , y4981 , y4982 , y4983 , y4984 , y4985 , y4986 , y4987 , y4988 , y4989 , y4990 , y4991 , y4992 , y4993 , y4994 , y4995 , y4996 , y4997 , y4998 , y4999 , y5000 , y5001 , y5002 , y5003 , y5004 , y5005 , y5006 , y5007 , y5008 , y5009 , y5010 , y5011 , y5012 , y5013 , y5014 , y5015 , y5016 , y5017 , y5018 , y5019 , y5020 , y5021 , y5022 , y5023 , y5024 , y5025 , y5026 , y5027 , y5028 , y5029 , y5030 , y5031 , y5032 , y5033 , y5034 , y5035 , y5036 , y5037 , y5038 , y5039 , y5040 , y5041 , y5042 , y5043 , y5044 , y5045 , y5046 , y5047 , y5048 , y5049 , y5050 , y5051 , y5052 , y5053 , y5054 , y5055 , y5056 , y5057 , y5058 , y5059 , y5060 , y5061 , y5062 , y5063 , y5064 , y5065 , y5066 , y5067 , y5068 , y5069 , y5070 , y5071 , y5072 , y5073 , y5074 , y5075 , y5076 , y5077 , y5078 , y5079 , y5080 , y5081 , y5082 , y5083 , y5084 , y5085 , y5086 , y5087 , y5088 , y5089 , y5090 , y5091 , y5092 , y5093 , y5094 , y5095 , y5096 , y5097 , y5098 , y5099 , y5100 , y5101 , y5102 , y5103 , y5104 , y5105 , y5106 , y5107 , y5108 , y5109 , y5110 , y5111 , y5112 , y5113 , y5114 , y5115 , y5116 , y5117 , y5118 , y5119 , y5120 , y5121 , y5122 , y5123 , y5124 , y5125 , y5126 , y5127 , y5128 , y5129 , y5130 , y5131 , y5132 , y5133 , y5134 , y5135 , y5136 , y5137 , y5138 , y5139 , y5140 , y5141 , y5142 , y5143 , y5144 , y5145 , y5146 , y5147 , y5148 , y5149 , y5150 , y5151 , y5152 , y5153 , y5154 , y5155 , y5156 , y5157 , y5158 , y5159 , y5160 , y5161 , y5162 , y5163 , y5164 , y5165 , y5166 , y5167 , y5168 , y5169 , y5170 , y5171 , y5172 , y5173 , y5174 , y5175 , y5176 , y5177 , y5178 , y5179 , y5180 , y5181 , y5182 , y5183 , y5184 , y5185 , y5186 , y5187 , y5188 , y5189 , y5190 , y5191 , y5192 , y5193 , y5194 , y5195 , y5196 , y5197 , y5198 , y5199 , y5200 , y5201 , y5202 , y5203 , y5204 , y5205 , y5206 , y5207 , y5208 , y5209 , y5210 , y5211 , y5212 , y5213 , y5214 , y5215 , y5216 , y5217 , y5218 , y5219 , y5220 , y5221 , y5222 , y5223 , y5224 , y5225 , y5226 , y5227 , y5228 , y5229 , y5230 , y5231 , y5232 , y5233 , y5234 , y5235 , y5236 , y5237 , y5238 , y5239 , y5240 , y5241 , y5242 , y5243 , y5244 , y5245 , y5246 , y5247 , y5248 , y5249 , y5250 , y5251 , y5252 , y5253 , y5254 , y5255 , y5256 , y5257 , y5258 , y5259 , y5260 , y5261 , y5262 , y5263 , y5264 , y5265 , y5266 , y5267 , y5268 , y5269 , y5270 , y5271 , y5272 , y5273 , y5274 , y5275 , y5276 , y5277 , y5278 , y5279 , y5280 , y5281 , y5282 , y5283 , y5284 , y5285 , y5286 , y5287 , y5288 , y5289 , y5290 , y5291 , y5292 , y5293 , y5294 , y5295 , y5296 , y5297 , y5298 , y5299 , y5300 , y5301 , y5302 , y5303 , y5304 , y5305 , y5306 , y5307 , y5308 , y5309 , y5310 , y5311 , y5312 , y5313 , y5314 , y5315 , y5316 , y5317 , y5318 , y5319 , y5320 , y5321 , y5322 , y5323 , y5324 , y5325 , y5326 , y5327 , y5328 , y5329 , y5330 , y5331 , y5332 , y5333 , y5334 , y5335 , y5336 , y5337 , y5338 , y5339 , y5340 , y5341 , y5342 , y5343 , y5344 , y5345 , y5346 , y5347 , y5348 , y5349 , y5350 , y5351 , y5352 , y5353 , y5354 , y5355 , y5356 , y5357 , y5358 , y5359 , y5360 , y5361 , y5362 , y5363 , y5364 , y5365 , y5366 , y5367 , y5368 , y5369 , y5370 , y5371 , y5372 , y5373 , y5374 , y5375 , y5376 , y5377 , y5378 , y5379 , y5380 , y5381 , y5382 , y5383 , y5384 , y5385 , y5386 , y5387 , y5388 , y5389 , y5390 , y5391 , y5392 , y5393 , y5394 , y5395 , y5396 , y5397 , y5398 , y5399 , y5400 , y5401 , y5402 , y5403 , y5404 , y5405 , y5406 , y5407 , y5408 , y5409 , y5410 , y5411 , y5412 , y5413 , y5414 , y5415 , y5416 , y5417 , y5418 , y5419 , y5420 , y5421 , y5422 , y5423 , y5424 , y5425 , y5426 , y5427 , y5428 , y5429 , y5430 , y5431 , y5432 , y5433 , y5434 , y5435 , y5436 , y5437 , y5438 , y5439 , y5440 , y5441 , y5442 , y5443 , y5444 , y5445 , y5446 , y5447 , y5448 , y5449 , y5450 , y5451 , y5452 , y5453 , y5454 , y5455 , y5456 , y5457 , y5458 , y5459 , y5460 , y5461 , y5462 , y5463 , y5464 , y5465 , y5466 , y5467 , y5468 , y5469 , y5470 , y5471 , y5472 , y5473 , y5474 , y5475 , y5476 , y5477 , y5478 , y5479 , y5480 , y5481 , y5482 , y5483 , y5484 , y5485 , y5486 , y5487 , y5488 , y5489 , y5490 , y5491 , y5492 , y5493 , y5494 , y5495 , y5496 , y5497 , y5498 , y5499 , y5500 , y5501 , y5502 , y5503 , y5504 , y5505 , y5506 , y5507 , y5508 , y5509 , y5510 , y5511 , y5512 , y5513 , y5514 , y5515 , y5516 , y5517 , y5518 , y5519 , y5520 , y5521 , y5522 , y5523 , y5524 , y5525 , y5526 , y5527 , y5528 , y5529 , y5530 , y5531 , y5532 , y5533 , y5534 , y5535 , y5536 , y5537 , y5538 , y5539 , y5540 , y5541 , y5542 , y5543 , y5544 , y5545 , y5546 , y5547 , y5548 , y5549 , y5550 , y5551 , y5552 , y5553 , y5554 , y5555 , y5556 , y5557 , y5558 , y5559 , y5560 , y5561 , y5562 , y5563 , y5564 , y5565 , y5566 , y5567 , y5568 , y5569 , y5570 , y5571 , y5572 , y5573 , y5574 , y5575 , y5576 , y5577 , y5578 , y5579 , y5580 , y5581 , y5582 , y5583 , y5584 , y5585 , y5586 , y5587 , y5588 , y5589 , y5590 , y5591 , y5592 , y5593 , y5594 , y5595 , y5596 , y5597 , y5598 , y5599 , y5600 , y5601 , y5602 , y5603 , y5604 , y5605 , y5606 , y5607 , y5608 , y5609 , y5610 , y5611 , y5612 , y5613 , y5614 , y5615 , y5616 , y5617 , y5618 , y5619 , y5620 , y5621 , y5622 , y5623 , y5624 , y5625 , y5626 , y5627 , y5628 , y5629 , y5630 , y5631 , y5632 , y5633 , y5634 , y5635 , y5636 , y5637 , y5638 , y5639 , y5640 , y5641 , y5642 , y5643 , y5644 , y5645 , y5646 , y5647 , y5648 , y5649 , y5650 , y5651 , y5652 , y5653 , y5654 , y5655 , y5656 , y5657 , y5658 , y5659 , y5660 , y5661 , y5662 , y5663 , y5664 , y5665 , y5666 , y5667 , y5668 , y5669 , y5670 , y5671 , y5672 , y5673 , y5674 , y5675 , y5676 , y5677 , y5678 , y5679 , y5680 , y5681 , y5682 , y5683 , y5684 , y5685 , y5686 , y5687 , y5688 , y5689 , y5690 , y5691 , y5692 , y5693 , y5694 , y5695 , y5696 , y5697 , y5698 , y5699 , y5700 , y5701 , y5702 , y5703 , y5704 , y5705 , y5706 , y5707 , y5708 , y5709 , y5710 , y5711 , y5712 , y5713 , y5714 , y5715 , y5716 , y5717 , y5718 , y5719 , y5720 , y5721 , y5722 , y5723 , y5724 , y5725 , y5726 , y5727 , y5728 , y5729 , y5730 , y5731 , y5732 , y5733 , y5734 , y5735 , y5736 , y5737 , y5738 , y5739 , y5740 , y5741 , y5742 , y5743 , y5744 , y5745 , y5746 , y5747 , y5748 , y5749 , y5750 , y5751 , y5752 , y5753 , y5754 , y5755 , y5756 , y5757 , y5758 , y5759 , y5760 , y5761 , y5762 , y5763 , y5764 , y5765 , y5766 , y5767 , y5768 , y5769 , y5770 , y5771 , y5772 , y5773 , y5774 , y5775 , y5776 , y5777 , y5778 , y5779 , y5780 , y5781 , y5782 , y5783 , y5784 , y5785 , y5786 , y5787 , y5788 , y5789 , y5790 , y5791 , y5792 , y5793 , y5794 , y5795 , y5796 , y5797 , y5798 , y5799 , y5800 , y5801 , y5802 , y5803 , y5804 , y5805 , y5806 , y5807 , y5808 , y5809 , y5810 , y5811 , y5812 , y5813 , y5814 , y5815 , y5816 , y5817 , y5818 , y5819 , y5820 , y5821 , y5822 , y5823 , y5824 , y5825 , y5826 , y5827 , y5828 , y5829 , y5830 , y5831 , y5832 , y5833 , y5834 , y5835 , y5836 , y5837 , y5838 , y5839 , y5840 , y5841 , y5842 , y5843 , y5844 , y5845 , y5846 , y5847 , y5848 , y5849 , y5850 , y5851 , y5852 , y5853 , y5854 , y5855 , y5856 , y5857 , y5858 , y5859 , y5860 , y5861 , y5862 , y5863 , y5864 , y5865 , y5866 , y5867 , y5868 , y5869 , y5870 , y5871 , y5872 , y5873 , y5874 , y5875 , y5876 , y5877 , y5878 , y5879 , y5880 , y5881 , y5882 , y5883 , y5884 , y5885 , y5886 , y5887 , y5888 , y5889 , y5890 , y5891 , y5892 , y5893 , y5894 , y5895 , y5896 , y5897 , y5898 , y5899 , y5900 , y5901 , y5902 , y5903 , y5904 , y5905 , y5906 , y5907 , y5908 , y5909 , y5910 , y5911 , y5912 , y5913 , y5914 , y5915 , y5916 , y5917 , y5918 , y5919 , y5920 , y5921 , y5922 , y5923 , y5924 , y5925 , y5926 , y5927 , y5928 , y5929 , y5930 , y5931 , y5932 , y5933 , y5934 , y5935 , y5936 , y5937 , y5938 , y5939 , y5940 , y5941 , y5942 , y5943 , y5944 , y5945 , y5946 , y5947 , y5948 , y5949 , y5950 , y5951 , y5952 , y5953 , y5954 , y5955 , y5956 , y5957 , y5958 , y5959 , y5960 , y5961 , y5962 , y5963 , y5964 , y5965 , y5966 , y5967 , y5968 , y5969 , y5970 , y5971 , y5972 , y5973 , y5974 , y5975 , y5976 , y5977 , y5978 , y5979 , y5980 , y5981 , y5982 , y5983 , y5984 , y5985 , y5986 , y5987 , y5988 , y5989 , y5990 , y5991 , y5992 , y5993 , y5994 , y5995 , y5996 , y5997 , y5998 , y5999 , y6000 , y6001 , y6002 , y6003 , y6004 , y6005 , y6006 , y6007 , y6008 , y6009 , y6010 , y6011 , y6012 , y6013 , y6014 , y6015 , y6016 , y6017 , y6018 , y6019 , y6020 , y6021 , y6022 , y6023 , y6024 , y6025 , y6026 , y6027 , y6028 , y6029 , y6030 , y6031 , y6032 , y6033 , y6034 , y6035 , y6036 , y6037 , y6038 , y6039 , y6040 , y6041 , y6042 , y6043 , y6044 , y6045 , y6046 , y6047 , y6048 , y6049 , y6050 , y6051 , y6052 , y6053 , y6054 , y6055 , y6056 , y6057 , y6058 , y6059 , y6060 , y6061 , y6062 , y6063 , y6064 , y6065 , y6066 , y6067 , y6068 , y6069 , y6070 , y6071 , y6072 , y6073 , y6074 , y6075 , y6076 , y6077 , y6078 , y6079 , y6080 , y6081 , y6082 , y6083 , y6084 , y6085 , y6086 , y6087 , y6088 , y6089 , y6090 , y6091 , y6092 , y6093 , y6094 , y6095 , y6096 , y6097 , y6098 , y6099 , y6100 , y6101 , y6102 , y6103 , y6104 , y6105 , y6106 , y6107 , y6108 , y6109 , y6110 , y6111 , y6112 , y6113 , y6114 , y6115 , y6116 , y6117 , y6118 , y6119 , y6120 , y6121 , y6122 , y6123 , y6124 , y6125 , y6126 , y6127 , y6128 , y6129 , y6130 , y6131 , y6132 , y6133 , y6134 , y6135 , y6136 , y6137 , y6138 , y6139 , y6140 , y6141 , y6142 , y6143 , y6144 , y6145 , y6146 , y6147 , y6148 , y6149 , y6150 , y6151 , y6152 , y6153 , y6154 , y6155 , y6156 , y6157 , y6158 , y6159 , y6160 , y6161 , y6162 , y6163 , y6164 , y6165 , y6166 , y6167 , y6168 , y6169 , y6170 , y6171 , y6172 , y6173 , y6174 , y6175 , y6176 , y6177 , y6178 , y6179 , y6180 , y6181 , y6182 , y6183 , y6184 , y6185 , y6186 , y6187 , y6188 , y6189 , y6190 , y6191 , y6192 , y6193 , y6194 , y6195 , y6196 , y6197 , y6198 , y6199 , y6200 , y6201 , y6202 , y6203 , y6204 , y6205 , y6206 , y6207 , y6208 , y6209 , y6210 , y6211 , y6212 , y6213 , y6214 , y6215 , y6216 , y6217 , y6218 , y6219 , y6220 , y6221 , y6222 , y6223 , y6224 , y6225 , y6226 , y6227 , y6228 , y6229 , y6230 , y6231 , y6232 , y6233 , y6234 , y6235 , y6236 , y6237 , y6238 , y6239 , y6240 , y6241 , y6242 , y6243 , y6244 , y6245 , y6246 , y6247 , y6248 , y6249 , y6250 , y6251 , y6252 , y6253 , y6254 , y6255 , y6256 , y6257 , y6258 , y6259 , y6260 , y6261 , y6262 , y6263 , y6264 , y6265 , y6266 , y6267 , y6268 , y6269 , y6270 , y6271 , y6272 , y6273 , y6274 , y6275 , y6276 , y6277 , y6278 , y6279 , y6280 , y6281 , y6282 , y6283 , y6284 , y6285 , y6286 , y6287 , y6288 , y6289 , y6290 , y6291 , y6292 , y6293 , y6294 , y6295 , y6296 , y6297 , y6298 , y6299 , y6300 , y6301 , y6302 , y6303 , y6304 , y6305 , y6306 , y6307 , y6308 , y6309 , y6310 , y6311 , y6312 , y6313 , y6314 , y6315 , y6316 , y6317 , y6318 , y6319 , y6320 , y6321 , y6322 , y6323 , y6324 , y6325 , y6326 , y6327 , y6328 , y6329 , y6330 , y6331 , y6332 , y6333 , y6334 , y6335 , y6336 , y6337 , y6338 , y6339 , y6340 , y6341 , y6342 , y6343 , y6344 , y6345 , y6346 , y6347 , y6348 , y6349 , y6350 , y6351 , y6352 , y6353 , y6354 , y6355 , y6356 , y6357 , y6358 , y6359 , y6360 , y6361 , y6362 , y6363 , y6364 , y6365 , y6366 , y6367 , y6368 , y6369 , y6370 , y6371 , y6372 , y6373 , y6374 , y6375 , y6376 , y6377 , y6378 , y6379 , y6380 , y6381 , y6382 , y6383 , y6384 , y6385 , y6386 , y6387 , y6388 , y6389 , y6390 , y6391 , y6392 , y6393 , y6394 , y6395 , y6396 , y6397 , y6398 , y6399 , y6400 , y6401 , y6402 , y6403 , y6404 , y6405 , y6406 , y6407 , y6408 , y6409 , y6410 , y6411 , y6412 , y6413 , y6414 , y6415 , y6416 , y6417 , y6418 , y6419 , y6420 , y6421 , y6422 , y6423 , y6424 , y6425 , y6426 , y6427 , y6428 , y6429 , y6430 , y6431 , y6432 , y6433 , y6434 , y6435 , y6436 , y6437 , y6438 , y6439 , y6440 , y6441 , y6442 , y6443 , y6444 , y6445 , y6446 , y6447 , y6448 , y6449 , y6450 , y6451 , y6452 , y6453 , y6454 , y6455 , y6456 , y6457 , y6458 , y6459 , y6460 , y6461 , y6462 , y6463 , y6464 , y6465 , y6466 , y6467 , y6468 , y6469 , y6470 , y6471 , y6472 , y6473 , y6474 , y6475 , y6476 , y6477 , y6478 , y6479 , y6480 , y6481 , y6482 , y6483 , y6484 , y6485 , y6486 , y6487 , y6488 , y6489 , y6490 , y6491 , y6492 , y6493 , y6494 , y6495 , y6496 , y6497 , y6498 , y6499 , y6500 , y6501 , y6502 , y6503 , y6504 , y6505 , y6506 , y6507 , y6508 , y6509 , y6510 , y6511 , y6512 , y6513 , y6514 , y6515 , y6516 , y6517 , y6518 , y6519 , y6520 , y6521 , y6522 , y6523 , y6524 , y6525 , y6526 , y6527 , y6528 , y6529 , y6530 , y6531 , y6532 , y6533 , y6534 , y6535 , y6536 , y6537 , y6538 , y6539 , y6540 , y6541 , y6542 , y6543 , y6544 , y6545 , y6546 , y6547 , y6548 , y6549 , y6550 , y6551 , y6552 , y6553 , y6554 , y6555 , y6556 , y6557 , y6558 , y6559 , y6560 , y6561 , y6562 , y6563 , y6564 , y6565 , y6566 , y6567 , y6568 , y6569 , y6570 , y6571 , y6572 , y6573 , y6574 , y6575 , y6576 , y6577 , y6578 , y6579 , y6580 , y6581 , y6582 , y6583 , y6584 , y6585 , y6586 , y6587 , y6588 , y6589 , y6590 , y6591 , y6592 , y6593 , y6594 , y6595 , y6596 , y6597 , y6598 , y6599 , y6600 , y6601 , y6602 , y6603 , y6604 , y6605 , y6606 , y6607 , y6608 , y6609 , y6610 , y6611 , y6612 , y6613 , y6614 , y6615 , y6616 , y6617 , y6618 , y6619 , y6620 , y6621 , y6622 , y6623 , y6624 , y6625 , y6626 , y6627 , y6628 , y6629 , y6630 , y6631 , y6632 , y6633 , y6634 , y6635 , y6636 , y6637 , y6638 , y6639 , y6640 , y6641 , y6642 , y6643 , y6644 , y6645 , y6646 , y6647 , y6648 , y6649 , y6650 , y6651 , y6652 , y6653 , y6654 , y6655 , y6656 , y6657 , y6658 , y6659 , y6660 , y6661 , y6662 , y6663 , y6664 , y6665 , y6666 , y6667 , y6668 , y6669 , y6670 , y6671 , y6672 , y6673 , y6674 , y6675 , y6676 , y6677 , y6678 , y6679 , y6680 , y6681 , y6682 , y6683 , y6684 , y6685 , y6686 , y6687 , y6688 , y6689 , y6690 , y6691 , y6692 , y6693 , y6694 , y6695 , y6696 , y6697 , y6698 , y6699 , y6700 , y6701 , y6702 , y6703 , y6704 , y6705 , y6706 , y6707 , y6708 , y6709 , y6710 , y6711 , y6712 , y6713 , y6714 , y6715 , y6716 , y6717 , y6718 , y6719 , y6720 , y6721 , y6722 , y6723 , y6724 , y6725 , y6726 , y6727 , y6728 , y6729 , y6730 , y6731 , y6732 , y6733 , y6734 , y6735 , y6736 , y6737 , y6738 , y6739 , y6740 , y6741 , y6742 , y6743 , y6744 , y6745 , y6746 , y6747 , y6748 , y6749 , y6750 , y6751 , y6752 , y6753 , y6754 , y6755 , y6756 , y6757 , y6758 , y6759 , y6760 , y6761 , y6762 , y6763 , y6764 , y6765 , y6766 , y6767 , y6768 , y6769 , y6770 , y6771 , y6772 , y6773 , y6774 , y6775 , y6776 , y6777 , y6778 , y6779 , y6780 , y6781 , y6782 , y6783 , y6784 , y6785 , y6786 , y6787 , y6788 , y6789 , y6790 , y6791 , y6792 , y6793 , y6794 , y6795 , y6796 , y6797 , y6798 , y6799 , y6800 , y6801 , y6802 , y6803 , y6804 , y6805 , y6806 , y6807 , y6808 , y6809 , y6810 , y6811 , y6812 , y6813 , y6814 , y6815 , y6816 , y6817 , y6818 , y6819 , y6820 , y6821 , y6822 , y6823 , y6824 , y6825 , y6826 , y6827 , y6828 , y6829 , y6830 , y6831 , y6832 , y6833 , y6834 , y6835 , y6836 , y6837 , y6838 , y6839 , y6840 , y6841 , y6842 , y6843 , y6844 , y6845 , y6846 , y6847 , y6848 , y6849 , y6850 , y6851 , y6852 , y6853 , y6854 , y6855 , y6856 , y6857 , y6858 , y6859 , y6860 , y6861 , y6862 , y6863 , y6864 , y6865 , y6866 , y6867 , y6868 , y6869 , y6870 , y6871 , y6872 , y6873 , y6874 , y6875 , y6876 , y6877 , y6878 , y6879 , y6880 , y6881 , y6882 , y6883 , y6884 , y6885 , y6886 , y6887 , y6888 , y6889 , y6890 , y6891 , y6892 , y6893 , y6894 , y6895 , y6896 , y6897 , y6898 , y6899 , y6900 , y6901 , y6902 , y6903 , y6904 , y6905 , y6906 , y6907 , y6908 , y6909 , y6910 , y6911 , y6912 , y6913 , y6914 , y6915 , y6916 , y6917 , y6918 , y6919 , y6920 , y6921 , y6922 , y6923 , y6924 , y6925 , y6926 , y6927 , y6928 , y6929 , y6930 , y6931 , y6932 , y6933 , y6934 , y6935 , y6936 , y6937 , y6938 , y6939 , y6940 , y6941 , y6942 , y6943 , y6944 , y6945 , y6946 , y6947 , y6948 , y6949 , y6950 , y6951 , y6952 , y6953 , y6954 , y6955 , y6956 , y6957 , y6958 , y6959 , y6960 , y6961 , y6962 , y6963 , y6964 , y6965 , y6966 , y6967 , y6968 , y6969 , y6970 , y6971 , y6972 , y6973 , y6974 , y6975 , y6976 , y6977 , y6978 , y6979 , y6980 , y6981 , y6982 , y6983 , y6984 , y6985 , y6986 , y6987 , y6988 , y6989 , y6990 , y6991 , y6992 , y6993 , y6994 , y6995 , y6996 , y6997 , y6998 , y6999 , y7000 , y7001 , y7002 , y7003 , y7004 , y7005 , y7006 , y7007 , y7008 , y7009 , y7010 , y7011 , y7012 , y7013 , y7014 , y7015 , y7016 , y7017 , y7018 , y7019 , y7020 , y7021 , y7022 , y7023 , y7024 , y7025 , y7026 , y7027 , y7028 , y7029 , y7030 , y7031 , y7032 , y7033 , y7034 , y7035 , y7036 , y7037 , y7038 , y7039 , y7040 , y7041 , y7042 , y7043 , y7044 , y7045 , y7046 , y7047 , y7048 , y7049 , y7050 , y7051 , y7052 , y7053 , y7054 , y7055 , y7056 , y7057 , y7058 , y7059 , y7060 , y7061 , y7062 , y7063 , y7064 , y7065 , y7066 , y7067 , y7068 , y7069 , y7070 , y7071 , y7072 , y7073 , y7074 , y7075 , y7076 , y7077 , y7078 , y7079 , y7080 , y7081 , y7082 , y7083 , y7084 , y7085 , y7086 , y7087 , y7088 , y7089 , y7090 , y7091 , y7092 , y7093 , y7094 , y7095 , y7096 , y7097 , y7098 , y7099 , y7100 , y7101 , y7102 , y7103 , y7104 , y7105 , y7106 , y7107 , y7108 , y7109 , y7110 , y7111 , y7112 , y7113 , y7114 , y7115 , y7116 , y7117 , y7118 , y7119 , y7120 , y7121 , y7122 , y7123 , y7124 , y7125 , y7126 , y7127 , y7128 , y7129 , y7130 , y7131 , y7132 , y7133 , y7134 , y7135 , y7136 , y7137 , y7138 , y7139 , y7140 , y7141 , y7142 , y7143 , y7144 , y7145 , y7146 , y7147 , y7148 , y7149 , y7150 , y7151 , y7152 , y7153 , y7154 , y7155 , y7156 , y7157 , y7158 , y7159 , y7160 , y7161 , y7162 , y7163 , y7164 , y7165 , y7166 , y7167 , y7168 , y7169 , y7170 , y7171 , y7172 , y7173 , y7174 , y7175 , y7176 , y7177 , y7178 , y7179 , y7180 , y7181 , y7182 , y7183 , y7184 , y7185 , y7186 , y7187 , y7188 , y7189 , y7190 , y7191 , y7192 , y7193 , y7194 , y7195 , y7196 , y7197 , y7198 , y7199 , y7200 , y7201 , y7202 , y7203 , y7204 , y7205 , y7206 , y7207 , y7208 , y7209 , y7210 , y7211 , y7212 , y7213 , y7214 , y7215 , y7216 , y7217 , y7218 , y7219 , y7220 , y7221 , y7222 , y7223 , y7224 , y7225 , y7226 , y7227 , y7228 , y7229 , y7230 , y7231 , y7232 , y7233 , y7234 , y7235 , y7236 , y7237 , y7238 , y7239 , y7240 , y7241 , y7242 , y7243 , y7244 , y7245 , y7246 , y7247 , y7248 , y7249 , y7250 , y7251 , y7252 , y7253 , y7254 , y7255 , y7256 , y7257 , y7258 , y7259 , y7260 , y7261 , y7262 , y7263 , y7264 , y7265 , y7266 , y7267 , y7268 , y7269 , y7270 , y7271 , y7272 , y7273 , y7274 , y7275 , y7276 , y7277 , y7278 , y7279 , y7280 , y7281 , y7282 , y7283 , y7284 , y7285 , y7286 , y7287 , y7288 , y7289 , y7290 , y7291 , y7292 , y7293 , y7294 , y7295 , y7296 , y7297 , y7298 , y7299 , y7300 , y7301 , y7302 , y7303 , y7304 , y7305 , y7306 , y7307 , y7308 , y7309 , y7310 , y7311 , y7312 , y7313 , y7314 , y7315 , y7316 , y7317 , y7318 , y7319 , y7320 , y7321 , y7322 , y7323 , y7324 , y7325 , y7326 , y7327 , y7328 , y7329 , y7330 , y7331 , y7332 , y7333 , y7334 , y7335 , y7336 , y7337 , y7338 , y7339 , y7340 , y7341 , y7342 , y7343 , y7344 , y7345 , y7346 , y7347 , y7348 , y7349 , y7350 , y7351 , y7352 , y7353 , y7354 , y7355 , y7356 , y7357 , y7358 , y7359 , y7360 , y7361 , y7362 , y7363 , y7364 , y7365 , y7366 , y7367 , y7368 , y7369 , y7370 , y7371 , y7372 , y7373 , y7374 , y7375 , y7376 , y7377 , y7378 , y7379 , y7380 , y7381 , y7382 , y7383 , y7384 , y7385 , y7386 , y7387 , y7388 , y7389 , y7390 , y7391 , y7392 , y7393 , y7394 , y7395 , y7396 , y7397 , y7398 , y7399 , y7400 , y7401 , y7402 , y7403 , y7404 , y7405 , y7406 , y7407 , y7408 , y7409 , y7410 , y7411 , y7412 , y7413 , y7414 , y7415 , y7416 , y7417 , y7418 , y7419 , y7420 , y7421 , y7422 , y7423 , y7424 , y7425 , y7426 , y7427 , y7428 , y7429 , y7430 , y7431 , y7432 , y7433 , y7434 , y7435 , y7436 , y7437 , y7438 , y7439 , y7440 , y7441 , y7442 , y7443 , y7444 , y7445 , y7446 , y7447 , y7448 , y7449 , y7450 , y7451 , y7452 , y7453 , y7454 , y7455 , y7456 , y7457 , y7458 , y7459 , y7460 , y7461 , y7462 , y7463 , y7464 , y7465 , y7466 , y7467 , y7468 , y7469 , y7470 , y7471 , y7472 , y7473 , y7474 , y7475 , y7476 , y7477 , y7478 , y7479 , y7480 , y7481 , y7482 , y7483 , y7484 , y7485 , y7486 , y7487 , y7488 , y7489 , y7490 , y7491 , y7492 , y7493 , y7494 , y7495 , y7496 , y7497 , y7498 , y7499 , y7500 , y7501 , y7502 , y7503 , y7504 , y7505 , y7506 , y7507 , y7508 , y7509 , y7510 , y7511 , y7512 , y7513 , y7514 , y7515 , y7516 , y7517 , y7518 , y7519 , y7520 , y7521 , y7522 , y7523 , y7524 , y7525 , y7526 , y7527 , y7528 , y7529 , y7530 , y7531 , y7532 , y7533 , y7534 , y7535 , y7536 , y7537 , y7538 , y7539 , y7540 , y7541 , y7542 , y7543 , y7544 , y7545 , y7546 , y7547 , y7548 , y7549 , y7550 , y7551 , y7552 , y7553 , y7554 , y7555 , y7556 , y7557 , y7558 , y7559 , y7560 , y7561 , y7562 , y7563 , y7564 , y7565 , y7566 , y7567 , y7568 , y7569 , y7570 , y7571 , y7572 , y7573 , y7574 , y7575 , y7576 , y7577 , y7578 , y7579 , y7580 , y7581 , y7582 , y7583 , y7584 , y7585 , y7586 , y7587 , y7588 , y7589 , y7590 , y7591 , y7592 , y7593 , y7594 , y7595 , y7596 , y7597 , y7598 , y7599 , y7600 , y7601 , y7602 , y7603 , y7604 , y7605 , y7606 , y7607 , y7608 , y7609 , y7610 , y7611 , y7612 , y7613 , y7614 , y7615 , y7616 , y7617 , y7618 , y7619 , y7620 , y7621 , y7622 , y7623 , y7624 , y7625 , y7626 , y7627 , y7628 , y7629 , y7630 , y7631 , y7632 , y7633 , y7634 , y7635 , y7636 , y7637 , y7638 , y7639 , y7640 , y7641 , y7642 , y7643 , y7644 , y7645 , y7646 , y7647 , y7648 , y7649 , y7650 , y7651 , y7652 , y7653 , y7654 , y7655 , y7656 , y7657 , y7658 , y7659 , y7660 , y7661 , y7662 , y7663 , y7664 , y7665 , y7666 , y7667 , y7668 , y7669 , y7670 , y7671 , y7672 , y7673 , y7674 , y7675 , y7676 , y7677 , y7678 , y7679 , y7680 , y7681 , y7682 , y7683 , y7684 , y7685 , y7686 , y7687 , y7688 , y7689 , y7690 , y7691 , y7692 , y7693 , y7694 , y7695 , y7696 , y7697 , y7698 , y7699 , y7700 , y7701 , y7702 , y7703 , y7704 , y7705 , y7706 , y7707 , y7708 , y7709 , y7710 , y7711 , y7712 , y7713 , y7714 , y7715 , y7716 , y7717 , y7718 , y7719 , y7720 , y7721 , y7722 , y7723 , y7724 , y7725 , y7726 , y7727 , y7728 , y7729 , y7730 , y7731 , y7732 , y7733 , y7734 , y7735 , y7736 , y7737 , y7738 , y7739 , y7740 , y7741 , y7742 , y7743 , y7744 , y7745 , y7746 , y7747 , y7748 , y7749 , y7750 , y7751 , y7752 , y7753 , y7754 , y7755 , y7756 , y7757 , y7758 , y7759 , y7760 , y7761 , y7762 , y7763 , y7764 , y7765 , y7766 , y7767 , y7768 , y7769 , y7770 , y7771 , y7772 , y7773 , y7774 , y7775 , y7776 , y7777 , y7778 , y7779 , y7780 , y7781 , y7782 , y7783 , y7784 , y7785 , y7786 , y7787 , y7788 , y7789 , y7790 , y7791 , y7792 , y7793 , y7794 , y7795 , y7796 , y7797 , y7798 , y7799 , y7800 , y7801 , y7802 , y7803 , y7804 , y7805 , y7806 , y7807 , y7808 , y7809 , y7810 , y7811 , y7812 , y7813 , y7814 , y7815 , y7816 , y7817 , y7818 , y7819 , y7820 , y7821 , y7822 , y7823 , y7824 , y7825 , y7826 , y7827 , y7828 , y7829 , y7830 , y7831 , y7832 , y7833 , y7834 , y7835 , y7836 , y7837 , y7838 , y7839 , y7840 , y7841 , y7842 , y7843 , y7844 , y7845 , y7846 , y7847 , y7848 , y7849 , y7850 , y7851 , y7852 , y7853 , y7854 , y7855 , y7856 , y7857 , y7858 , y7859 , y7860 , y7861 , y7862 , y7863 , y7864 , y7865 , y7866 , y7867 , y7868 , y7869 , y7870 , y7871 , y7872 , y7873 , y7874 , y7875 , y7876 , y7877 , y7878 , y7879 , y7880 , y7881 , y7882 , y7883 , y7884 , y7885 , y7886 , y7887 , y7888 , y7889 , y7890 , y7891 , y7892 , y7893 , y7894 , y7895 , y7896 , y7897 , y7898 , y7899 , y7900 , y7901 , y7902 , y7903 , y7904 , y7905 , y7906 , y7907 , y7908 , y7909 , y7910 , y7911 , y7912 , y7913 , y7914 , y7915 , y7916 , y7917 , y7918 , y7919 , y7920 , y7921 , y7922 , y7923 , y7924 , y7925 , y7926 , y7927 , y7928 , y7929 , y7930 , y7931 , y7932 , y7933 , y7934 , y7935 , y7936 , y7937 , y7938 , y7939 , y7940 , y7941 , y7942 , y7943 , y7944 , y7945 , y7946 , y7947 , y7948 , y7949 , y7950 , y7951 , y7952 , y7953 , y7954 , y7955 , y7956 , y7957 , y7958 , y7959 , y7960 , y7961 , y7962 , y7963 , y7964 , y7965 , y7966 , y7967 , y7968 , y7969 , y7970 , y7971 , y7972 , y7973 , y7974 , y7975 , y7976 , y7977 , y7978 , y7979 , y7980 , y7981 , y7982 , y7983 , y7984 , y7985 , y7986 , y7987 , y7988 , y7989 , y7990 , y7991 , y7992 , y7993 , y7994 , y7995 , y7996 , y7997 , y7998 , y7999 , y8000 , y8001 , y8002 , y8003 , y8004 , y8005 , y8006 , y8007 , y8008 , y8009 , y8010 , y8011 , y8012 , y8013 , y8014 , y8015 , y8016 , y8017 , y8018 , y8019 , y8020 , y8021 , y8022 , y8023 , y8024 , y8025 , y8026 , y8027 , y8028 , y8029 , y8030 , y8031 , y8032 , y8033 , y8034 , y8035 , y8036 , y8037 , y8038 , y8039 , y8040 , y8041 , y8042 , y8043 , y8044 , y8045 , y8046 , y8047 , y8048 , y8049 , y8050 , y8051 , y8052 , y8053 , y8054 , y8055 , y8056 , y8057 , y8058 , y8059 , y8060 , y8061 , y8062 , y8063 , y8064 , y8065 , y8066 , y8067 , y8068 , y8069 , y8070 , y8071 , y8072 , y8073 , y8074 , y8075 , y8076 , y8077 , y8078 , y8079 , y8080 , y8081 , y8082 , y8083 , y8084 , y8085 , y8086 , y8087 , y8088 , y8089 , y8090 , y8091 , y8092 , y8093 , y8094 , y8095 , y8096 , y8097 , y8098 , y8099 , y8100 , y8101 , y8102 , y8103 , y8104 , y8105 , y8106 , y8107 , y8108 , y8109 , y8110 , y8111 , y8112 , y8113 , y8114 , y8115 , y8116 , y8117 , y8118 , y8119 , y8120 , y8121 , y8122 , y8123 , y8124 , y8125 , y8126 , y8127 , y8128 , y8129 , y8130 , y8131 , y8132 , y8133 , y8134 , y8135 , y8136 , y8137 , y8138 , y8139 , y8140 , y8141 , y8142 , y8143 , y8144 , y8145 , y8146 , y8147 , y8148 , y8149 , y8150 , y8151 , y8152 , y8153 , y8154 , y8155 , y8156 , y8157 , y8158 , y8159 , y8160 , y8161 , y8162 , y8163 , y8164 , y8165 , y8166 , y8167 , y8168 , y8169 , y8170 , y8171 , y8172 , y8173 , y8174 , y8175 , y8176 , y8177 , y8178 , y8179 , y8180 , y8181 , y8182 , y8183 , y8184 , y8185 , y8186 , y8187 , y8188 , y8189 , y8190 , y8191 , y8192 , y8193 , y8194 , y8195 , y8196 , y8197 , y8198 , y8199 , y8200 , y8201 , y8202 , y8203 , y8204 , y8205 , y8206 , y8207 , y8208 , y8209 , y8210 , y8211 , y8212 , y8213 , y8214 , y8215 , y8216 , y8217 , y8218 , y8219 , y8220 , y8221 , y8222 , y8223 , y8224 , y8225 , y8226 , y8227 , y8228 , y8229 , y8230 , y8231 , y8232 , y8233 , y8234 , y8235 , y8236 , y8237 , y8238 , y8239 , y8240 , y8241 , y8242 , y8243 , y8244 , y8245 , y8246 , y8247 , y8248 , y8249 , y8250 , y8251 , y8252 , y8253 , y8254 , y8255 , y8256 , y8257 , y8258 , y8259 , y8260 , y8261 , y8262 , y8263 , y8264 , y8265 , y8266 , y8267 , y8268 , y8269 , y8270 , y8271 , y8272 , y8273 , y8274 , y8275 , y8276 , y8277 , y8278 , y8279 , y8280 , y8281 , y8282 , y8283 , y8284 , y8285 , y8286 , y8287 , y8288 , y8289 , y8290 , y8291 , y8292 , y8293 , y8294 , y8295 , y8296 , y8297 , y8298 , y8299 , y8300 , y8301 , y8302 , y8303 , y8304 , y8305 , y8306 , y8307 , y8308 , y8309 , y8310 , y8311 , y8312 , y8313 , y8314 , y8315 , y8316 , y8317 , y8318 , y8319 , y8320 , y8321 , y8322 , y8323 , y8324 , y8325 , y8326 , y8327 , y8328 , y8329 , y8330 , y8331 , y8332 , y8333 , y8334 , y8335 , y8336 , y8337 , y8338 , y8339 , y8340 , y8341 , y8342 , y8343 , y8344 , y8345 , y8346 , y8347 , y8348 , y8349 , y8350 , y8351 , y8352 , y8353 , y8354 , y8355 , y8356 , y8357 , y8358 , y8359 , y8360 , y8361 , y8362 , y8363 , y8364 , y8365 , y8366 , y8367 , y8368 , y8369 , y8370 , y8371 , y8372 , y8373 , y8374 , y8375 , y8376 , y8377 , y8378 , y8379 , y8380 , y8381 , y8382 , y8383 , y8384 , y8385 , y8386 , y8387 , y8388 , y8389 , y8390 , y8391 , y8392 , y8393 , y8394 , y8395 , y8396 , y8397 , y8398 , y8399 , y8400 , y8401 , y8402 , y8403 , y8404 , y8405 , y8406 , y8407 , y8408 , y8409 , y8410 , y8411 , y8412 , y8413 , y8414 , y8415 , y8416 , y8417 , y8418 , y8419 , y8420 , y8421 , y8422 , y8423 , y8424 , y8425 , y8426 , y8427 , y8428 , y8429 , y8430 , y8431 , y8432 , y8433 , y8434 , y8435 , y8436 , y8437 , y8438 , y8439 , y8440 , y8441 , y8442 , y8443 , y8444 , y8445 , y8446 , y8447 , y8448 , y8449 , y8450 , y8451 , y8452 , y8453 , y8454 , y8455 , y8456 , y8457 , y8458 , y8459 , y8460 , y8461 , y8462 , y8463 , y8464 , y8465 , y8466 , y8467 , y8468 , y8469 , y8470 , y8471 , y8472 , y8473 , y8474 , y8475 , y8476 , y8477 , y8478 , y8479 , y8480 , y8481 , y8482 , y8483 , y8484 , y8485 , y8486 , y8487 , y8488 , y8489 , y8490 , y8491 , y8492 , y8493 , y8494 , y8495 , y8496 , y8497 , y8498 , y8499 , y8500 , y8501 , y8502 , y8503 , y8504 , y8505 , y8506 , y8507 , y8508 , y8509 , y8510 , y8511 , y8512 , y8513 , y8514 , y8515 , y8516 , y8517 , y8518 , y8519 , y8520 , y8521 , y8522 , y8523 , y8524 , y8525 , y8526 , y8527 , y8528 , y8529 , y8530 , y8531 , y8532 , y8533 , y8534 , y8535 , y8536 , y8537 , y8538 , y8539 , y8540 , y8541 , y8542 , y8543 , y8544 , y8545 , y8546 , y8547 , y8548 , y8549 , y8550 , y8551 , y8552 , y8553 , y8554 , y8555 , y8556 , y8557 , y8558 , y8559 , y8560 , y8561 , y8562 , y8563 , y8564 , y8565 , y8566 , y8567 , y8568 , y8569 , y8570 , y8571 , y8572 , y8573 , y8574 , y8575 , y8576 , y8577 , y8578 , y8579 , y8580 , y8581 , y8582 , y8583 , y8584 , y8585 , y8586 , y8587 , y8588 , y8589 , y8590 , y8591 , y8592 , y8593 , y8594 , y8595 , y8596 , y8597 , y8598 , y8599 , y8600 , y8601 , y8602 , y8603 , y8604 , y8605 , y8606 , y8607 , y8608 , y8609 , y8610 , y8611 , y8612 , y8613 , y8614 , y8615 , y8616 , y8617 , y8618 , y8619 , y8620 , y8621 , y8622 , y8623 , y8624 , y8625 , y8626 , y8627 , y8628 , y8629 , y8630 , y8631 , y8632 , y8633 , y8634 , y8635 , y8636 , y8637 , y8638 , y8639 , y8640 , y8641 , y8642 , y8643 , y8644 , y8645 , y8646 , y8647 , y8648 , y8649 , y8650 , y8651 , y8652 , y8653 , y8654 , y8655 , y8656 , y8657 , y8658 , y8659 , y8660 , y8661 , y8662 , y8663 , y8664 , y8665 , y8666 , y8667 , y8668 , y8669 , y8670 , y8671 , y8672 , y8673 , y8674 , y8675 , y8676 , y8677 , y8678 , y8679 , y8680 , y8681 , y8682 , y8683 , y8684 , y8685 , y8686 , y8687 , y8688 , y8689 , y8690 , y8691 , y8692 , y8693 , y8694 , y8695 , y8696 , y8697 , y8698 , y8699 , y8700 , y8701 , y8702 , y8703 , y8704 , y8705 , y8706 , y8707 , y8708 , y8709 , y8710 , y8711 , y8712 , y8713 , y8714 , y8715 , y8716 , y8717 , y8718 , y8719 , y8720 , y8721 , y8722 , y8723 , y8724 , y8725 , y8726 , y8727 , y8728 , y8729 , y8730 , y8731 , y8732 , y8733 , y8734 , y8735 , y8736 , y8737 , y8738 , y8739 , y8740 , y8741 , y8742 , y8743 , y8744 , y8745 , y8746 , y8747 , y8748 , y8749 , y8750 , y8751 , y8752 , y8753 , y8754 , y8755 , y8756 , y8757 , y8758 , y8759 , y8760 , y8761 , y8762 , y8763 , y8764 , y8765 , y8766 , y8767 , y8768 , y8769 , y8770 , y8771 , y8772 , y8773 , y8774 , y8775 , y8776 , y8777 , y8778 , y8779 , y8780 , y8781 , y8782 , y8783 , y8784 , y8785 , y8786 , y8787 , y8788 , y8789 , y8790 , y8791 , y8792 , y8793 , y8794 , y8795 , y8796 , y8797 , y8798 , y8799 , y8800 , y8801 , y8802 , y8803 , y8804 , y8805 , y8806 , y8807 , y8808 , y8809 , y8810 , y8811 , y8812 , y8813 , y8814 , y8815 , y8816 , y8817 , y8818 , y8819 , y8820 , y8821 , y8822 , y8823 , y8824 , y8825 , y8826 , y8827 , y8828 , y8829 , y8830 , y8831 , y8832 , y8833 , y8834 , y8835 , y8836 , y8837 , y8838 , y8839 , y8840 , y8841 , y8842 , y8843 , y8844 , y8845 , y8846 , y8847 , y8848 , y8849 , y8850 , y8851 , y8852 , y8853 , y8854 , y8855 , y8856 , y8857 , y8858 , y8859 , y8860 , y8861 , y8862 , y8863 , y8864 , y8865 , y8866 , y8867 , y8868 , y8869 , y8870 , y8871 , y8872 , y8873 , y8874 , y8875 , y8876 , y8877 , y8878 , y8879 , y8880 , y8881 , y8882 , y8883 , y8884 , y8885 , y8886 , y8887 , y8888 , y8889 , y8890 , y8891 , y8892 , y8893 , y8894 , y8895 , y8896 , y8897 , y8898 , y8899 , y8900 , y8901 , y8902 , y8903 , y8904 , y8905 , y8906 , y8907 , y8908 , y8909 , y8910 , y8911 , y8912 , y8913 , y8914 , y8915 , y8916 , y8917 , y8918 , y8919 , y8920 , y8921 , y8922 , y8923 , y8924 , y8925 , y8926 , y8927 , y8928 , y8929 , y8930 , y8931 , y8932 , y8933 , y8934 , y8935 , y8936 , y8937 , y8938 , y8939 , y8940 , y8941 , y8942 , y8943 , y8944 , y8945 , y8946 , y8947 , y8948 , y8949 , y8950 , y8951 , y8952 , y8953 , y8954 , y8955 , y8956 , y8957 , y8958 , y8959 , y8960 , y8961 , y8962 , y8963 , y8964 , y8965 , y8966 , y8967 , y8968 , y8969 , y8970 , y8971 , y8972 , y8973 , y8974 , y8975 , y8976 , y8977 , y8978 , y8979 , y8980 , y8981 , y8982 , y8983 , y8984 , y8985 , y8986 , y8987 , y8988 , y8989 , y8990 , y8991 , y8992 , y8993 , y8994 , y8995 , y8996 , y8997 , y8998 , y8999 , y9000 , y9001 , y9002 , y9003 , y9004 , y9005 , y9006 , y9007 , y9008 , y9009 , y9010 , y9011 , y9012 , y9013 , y9014 , y9015 , y9016 , y9017 , y9018 , y9019 , y9020 , y9021 , y9022 , y9023 , y9024 , y9025 , y9026 , y9027 , y9028 , y9029 , y9030 , y9031 , y9032 , y9033 , y9034 , y9035 , y9036 , y9037 , y9038 , y9039 , y9040 , y9041 , y9042 , y9043 , y9044 , y9045 , y9046 , y9047 , y9048 , y9049 , y9050 , y9051 , y9052 , y9053 , y9054 , y9055 , y9056 , y9057 , y9058 , y9059 , y9060 , y9061 , y9062 , y9063 , y9064 , y9065 , y9066 , y9067 , y9068 , y9069 , y9070 , y9071 , y9072 , y9073 , y9074 , y9075 , y9076 , y9077 , y9078 , y9079 , y9080 , y9081 , y9082 , y9083 , y9084 , y9085 , y9086 , y9087 , y9088 , y9089 , y9090 , y9091 , y9092 , y9093 , y9094 , y9095 , y9096 , y9097 , y9098 , y9099 , y9100 , y9101 , y9102 , y9103 , y9104 , y9105 , y9106 , y9107 , y9108 , y9109 , y9110 , y9111 , y9112 , y9113 , y9114 , y9115 , y9116 , y9117 , y9118 , y9119 , y9120 , y9121 , y9122 , y9123 , y9124 , y9125 , y9126 , y9127 , y9128 , y9129 , y9130 , y9131 , y9132 , y9133 , y9134 , y9135 , y9136 , y9137 , y9138 , y9139 , y9140 , y9141 , y9142 , y9143 , y9144 , y9145 , y9146 , y9147 , y9148 , y9149 , y9150 , y9151 , y9152 , y9153 , y9154 , y9155 , y9156 , y9157 , y9158 , y9159 , y9160 , y9161 , y9162 , y9163 , y9164 , y9165 , y9166 , y9167 , y9168 , y9169 , y9170 , y9171 , y9172 , y9173 , y9174 , y9175 , y9176 , y9177 , y9178 , y9179 , y9180 , y9181 , y9182 , y9183 , y9184 , y9185 , y9186 , y9187 , y9188 , y9189 , y9190 , y9191 , y9192 , y9193 , y9194 , y9195 , y9196 , y9197 , y9198 , y9199 , y9200 , y9201 , y9202 , y9203 , y9204 , y9205 , y9206 , y9207 , y9208 , y9209 , y9210 , y9211 , y9212 , y9213 , y9214 , y9215 , y9216 , y9217 , y9218 , y9219 , y9220 , y9221 , y9222 , y9223 , y9224 , y9225 , y9226 , y9227 , y9228 , y9229 , y9230 , y9231 , y9232 , y9233 , y9234 , y9235 , y9236 , y9237 , y9238 , y9239 , y9240 , y9241 , y9242 , y9243 , y9244 , y9245 , y9246 , y9247 , y9248 , y9249 , y9250 , y9251 , y9252 , y9253 , y9254 , y9255 , y9256 , y9257 , y9258 , y9259 , y9260 , y9261 , y9262 , y9263 , y9264 , y9265 , y9266 , y9267 , y9268 , y9269 , y9270 , y9271 , y9272 , y9273 , y9274 , y9275 , y9276 , y9277 , y9278 , y9279 , y9280 , y9281 , y9282 , y9283 , y9284 , y9285 , y9286 , y9287 , y9288 , y9289 , y9290 , y9291 , y9292 , y9293 , y9294 , y9295 , y9296 , y9297 , y9298 , y9299 , y9300 , y9301 , y9302 , y9303 , y9304 , y9305 , y9306 , y9307 , y9308 , y9309 , y9310 , y9311 , y9312 , y9313 , y9314 , y9315 , y9316 , y9317 , y9318 , y9319 , y9320 , y9321 , y9322 , y9323 , y9324 , y9325 , y9326 , y9327 , y9328 , y9329 , y9330 , y9331 , y9332 , y9333 , y9334 , y9335 , y9336 , y9337 , y9338 , y9339 , y9340 , y9341 , y9342 , y9343 , y9344 , y9345 , y9346 , y9347 , y9348 , y9349 , y9350 , y9351 , y9352 , y9353 , y9354 , y9355 , y9356 , y9357 , y9358 , y9359 , y9360 , y9361 , y9362 , y9363 , y9364 , y9365 , y9366 , y9367 , y9368 , y9369 , y9370 , y9371 , y9372 , y9373 , y9374 , y9375 , y9376 , y9377 , y9378 , y9379 , y9380 , y9381 , y9382 , y9383 , y9384 , y9385 , y9386 , y9387 , y9388 , y9389 , y9390 , y9391 , y9392 , y9393 , y9394 , y9395 , y9396 , y9397 , y9398 , y9399 , y9400 , y9401 , y9402 , y9403 , y9404 , y9405 , y9406 , y9407 , y9408 , y9409 , y9410 , y9411 , y9412 , y9413 , y9414 , y9415 , y9416 , y9417 , y9418 , y9419 , y9420 , y9421 , y9422 , y9423 , y9424 , y9425 , y9426 , y9427 , y9428 , y9429 , y9430 , y9431 , y9432 , y9433 , y9434 , y9435 , y9436 , y9437 , y9438 , y9439 , y9440 , y9441 , y9442 , y9443 , y9444 , y9445 , y9446 , y9447 , y9448 , y9449 , y9450 , y9451 , y9452 , y9453 , y9454 , y9455 , y9456 , y9457 , y9458 , y9459 , y9460 , y9461 , y9462 , y9463 , y9464 , y9465 , y9466 , y9467 , y9468 , y9469 , y9470 , y9471 , y9472 , y9473 , y9474 , y9475 , y9476 , y9477 , y9478 , y9479 , y9480 , y9481 , y9482 , y9483 , y9484 , y9485 , y9486 , y9487 , y9488 , y9489 , y9490 , y9491 , y9492 , y9493 , y9494 , y9495 , y9496 , y9497 , y9498 , y9499 , y9500 , y9501 , y9502 , y9503 , y9504 , y9505 , y9506 , y9507 , y9508 , y9509 , y9510 , y9511 , y9512 , y9513 , y9514 , y9515 , y9516 , y9517 , y9518 , y9519 , y9520 , y9521 , y9522 , y9523 , y9524 , y9525 , y9526 , y9527 , y9528 , y9529 , y9530 , y9531 , y9532 , y9533 , y9534 , y9535 , y9536 , y9537 , y9538 , y9539 , y9540 , y9541 , y9542 , y9543 , y9544 , y9545 , y9546 , y9547 , y9548 , y9549 , y9550 , y9551 , y9552 , y9553 , y9554 , y9555 , y9556 , y9557 , y9558 , y9559 , y9560 , y9561 , y9562 , y9563 , y9564 , y9565 , y9566 , y9567 , y9568 , y9569 , y9570 , y9571 , y9572 , y9573 , y9574 , y9575 , y9576 , y9577 , y9578 , y9579 , y9580 , y9581 , y9582 , y9583 , y9584 , y9585 , y9586 , y9587 , y9588 , y9589 , y9590 , y9591 , y9592 , y9593 , y9594 , y9595 , y9596 , y9597 , y9598 , y9599 , y9600 , y9601 , y9602 , y9603 , y9604 , y9605 , y9606 , y9607 , y9608 , y9609 , y9610 , y9611 , y9612 , y9613 , y9614 , y9615 , y9616 , y9617 , y9618 , y9619 , y9620 , y9621 , y9622 , y9623 , y9624 , y9625 , y9626 , y9627 , y9628 , y9629 , y9630 , y9631 , y9632 , y9633 , y9634 , y9635 , y9636 , y9637 , y9638 , y9639 , y9640 , y9641 , y9642 , y9643 , y9644 , y9645 , y9646 , y9647 , y9648 , y9649 , y9650 , y9651 , y9652 , y9653 , y9654 , y9655 , y9656 , y9657 , y9658 , y9659 , y9660 , y9661 , y9662 , y9663 , y9664 , y9665 , y9666 , y9667 , y9668 , y9669 , y9670 , y9671 , y9672 , y9673 , y9674 , y9675 , y9676 , y9677 , y9678 , y9679 , y9680 , y9681 , y9682 , y9683 , y9684 , y9685 , y9686 , y9687 , y9688 , y9689 , y9690 , y9691 , y9692 , y9693 , y9694 , y9695 , y9696 , y9697 , y9698 , y9699 , y9700 , y9701 , y9702 , y9703 , y9704 , y9705 , y9706 , y9707 , y9708 , y9709 , y9710 , y9711 , y9712 , y9713 , y9714 , y9715 , y9716 , y9717 , y9718 , y9719 , y9720 , y9721 , y9722 , y9723 , y9724 , y9725 , y9726 , y9727 , y9728 , y9729 , y9730 , y9731 , y9732 , y9733 , y9734 , y9735 , y9736 , y9737 , y9738 , y9739 , y9740 , y9741 , y9742 , y9743 , y9744 , y9745 , y9746 , y9747 , y9748 , y9749 , y9750 , y9751 , y9752 , y9753 , y9754 , y9755 , y9756 , y9757 , y9758 , y9759 , y9760 , y9761 , y9762 , y9763 , y9764 , y9765 , y9766 , y9767 , y9768 , y9769 , y9770 , y9771 , y9772 , y9773 , y9774 , y9775 , y9776 , y9777 , y9778 , y9779 , y9780 , y9781 , y9782 , y9783 , y9784 , y9785 , y9786 , y9787 , y9788 , y9789 , y9790 , y9791 , y9792 , y9793 , y9794 , y9795 , y9796 , y9797 , y9798 , y9799 , y9800 , y9801 , y9802 , y9803 , y9804 , y9805 , y9806 , y9807 , y9808 , y9809 , y9810 , y9811 , y9812 , y9813 , y9814 , y9815 , y9816 , y9817 , y9818 , y9819 , y9820 , y9821 , y9822 , y9823 , y9824 , y9825 , y9826 , y9827 , y9828 , y9829 , y9830 , y9831 , y9832 , y9833 , y9834 , y9835 , y9836 , y9837 , y9838 , y9839 , y9840 , y9841 , y9842 , y9843 , y9844 , y9845 , y9846 , y9847 , y9848 , y9849 , y9850 , y9851 , y9852 , y9853 , y9854 , y9855 , y9856 , y9857 , y9858 , y9859 , y9860 , y9861 , y9862 , y9863 , y9864 , y9865 , y9866 , y9867 , y9868 , y9869 , y9870 , y9871 , y9872 , y9873 , y9874 , y9875 , y9876 , y9877 , y9878 , y9879 , y9880 , y9881 , y9882 , y9883 , y9884 , y9885 , y9886 , y9887 , y9888 , y9889 , y9890 , y9891 , y9892 , y9893 , y9894 , y9895 , y9896 , y9897 , y9898 , y9899 , y9900 , y9901 , y9902 , y9903 , y9904 , y9905 , y9906 , y9907 , y9908 , y9909 , y9910 , y9911 , y9912 , y9913 , y9914 , y9915 , y9916 , y9917 , y9918 , y9919 , y9920 , y9921 , y9922 , y9923 , y9924 , y9925 , y9926 , y9927 , y9928 , y9929 , y9930 , y9931 , y9932 , y9933 , y9934 , y9935 , y9936 , y9937 , y9938 , y9939 , y9940 , y9941 , y9942 , y9943 , y9944 , y9945 , y9946 , y9947 , y9948 , y9949 , y9950 , y9951 , y9952 , y9953 , y9954 , y9955 , y9956 , y9957 , y9958 , y9959 , y9960 , y9961 , y9962 , y9963 , y9964 , y9965 , y9966 , y9967 , y9968 , y9969 , y9970 , y9971 , y9972 , y9973 , y9974 , y9975 , y9976 , y9977 , y9978 , y9979 , y9980 , y9981 , y9982 , y9983 , y9984 , y9985 , y9986 , y9987 , y9988 , y9989 , y9990 , y9991 , y9992 , y9993 , y9994 , y9995 , y9996 , y9997 , y9998 , y9999 , y10000 , y10001 , y10002 , y10003 , y10004 , y10005 , y10006 , y10007 , y10008 , y10009 , y10010 , y10011 , y10012 , y10013 , y10014 , y10015 , y10016 , y10017 , y10018 , y10019 , y10020 , y10021 , y10022 , y10023 , y10024 , y10025 , y10026 , y10027 , y10028 , y10029 , y10030 , y10031 , y10032 , y10033 , y10034 , y10035 , y10036 , y10037 , y10038 , y10039 , y10040 , y10041 , y10042 , y10043 , y10044 , y10045 , y10046 , y10047 , y10048 , y10049 , y10050 , y10051 , y10052 , y10053 , y10054 , y10055 , y10056 , y10057 , y10058 , y10059 , y10060 , y10061 , y10062 , y10063 , y10064 , y10065 , y10066 , y10067 , y10068 , y10069 , y10070 , y10071 , y10072 , y10073 , y10074 , y10075 , y10076 , y10077 , y10078 , y10079 , y10080 , y10081 , y10082 , y10083 , y10084 , y10085 , y10086 , y10087 , y10088 , y10089 , y10090 , y10091 , y10092 , y10093 , y10094 , y10095 , y10096 , y10097 , y10098 , y10099 , y10100 , y10101 , y10102 , y10103 , y10104 , y10105 , y10106 , y10107 , y10108 , y10109 , y10110 , y10111 , y10112 , y10113 , y10114 , y10115 , y10116 , y10117 , y10118 , y10119 , y10120 , y10121 , y10122 , y10123 , y10124 , y10125 , y10126 , y10127 , y10128 , y10129 , y10130 , y10131 , y10132 , y10133 , y10134 , y10135 , y10136 , y10137 , y10138 , y10139 , y10140 , y10141 , y10142 , y10143 , y10144 , y10145 , y10146 , y10147 , y10148 , y10149 , y10150 , y10151 , y10152 , y10153 , y10154 , y10155 , y10156 , y10157 , y10158 , y10159 , y10160 , y10161 , y10162 , y10163 , y10164 , y10165 , y10166 , y10167 , y10168 , y10169 , y10170 , y10171 , y10172 , y10173 , y10174 , y10175 , y10176 , y10177 , y10178 , y10179 , y10180 , y10181 , y10182 , y10183 , y10184 , y10185 , y10186 , y10187 , y10188 , y10189 , y10190 , y10191 , y10192 , y10193 , y10194 , y10195 , y10196 , y10197 , y10198 , y10199 , y10200 , y10201 , y10202 , y10203 , y10204 , y10205 , y10206 , y10207 , y10208 , y10209 , y10210 , y10211 , y10212 , y10213 , y10214 , y10215 , y10216 , y10217 , y10218 , y10219 , y10220 , y10221 , y10222 , y10223 , y10224 , y10225 , y10226 , y10227 , y10228 , y10229 , y10230 , y10231 , y10232 , y10233 , y10234 , y10235 , y10236 , y10237 , y10238 , y10239 , y10240 , y10241 , y10242 , y10243 , y10244 , y10245 , y10246 , y10247 , y10248 , y10249 , y10250 , y10251 , y10252 , y10253 , y10254 , y10255 , y10256 , y10257 , y10258 , y10259 , y10260 , y10261 , y10262 , y10263 , y10264 , y10265 , y10266 , y10267 , y10268 , y10269 , y10270 , y10271 , y10272 , y10273 , y10274 , y10275 , y10276 , y10277 , y10278 , y10279 , y10280 , y10281 , y10282 , y10283 , y10284 , y10285 , y10286 , y10287 , y10288 , y10289 , y10290 , y10291 , y10292 , y10293 , y10294 , y10295 , y10296 , y10297 , y10298 , y10299 , y10300 , y10301 , y10302 , y10303 , y10304 , y10305 , y10306 , y10307 , y10308 , y10309 , y10310 , y10311 , y10312 , y10313 , y10314 , y10315 , y10316 , y10317 , y10318 , y10319 , y10320 , y10321 , y10322 , y10323 , y10324 , y10325 , y10326 , y10327 , y10328 , y10329 , y10330 , y10331 , y10332 , y10333 , y10334 , y10335 , y10336 , y10337 , y10338 , y10339 , y10340 , y10341 , y10342 , y10343 , y10344 , y10345 , y10346 , y10347 , y10348 , y10349 , y10350 , y10351 , y10352 , y10353 , y10354 , y10355 , y10356 , y10357 , y10358 , y10359 , y10360 , y10361 , y10362 , y10363 , y10364 , y10365 , y10366 , y10367 , y10368 , y10369 , y10370 , y10371 , y10372 , y10373 , y10374 , y10375 , y10376 , y10377 , y10378 , y10379 , y10380 , y10381 , y10382 , y10383 , y10384 , y10385 , y10386 , y10387 , y10388 , y10389 , y10390 , y10391 , y10392 , y10393 , y10394 , y10395 , y10396 , y10397 , y10398 , y10399 , y10400 , y10401 , y10402 , y10403 , y10404 , y10405 , y10406 , y10407 , y10408 , y10409 , y10410 , y10411 , y10412 , y10413 , y10414 , y10415 , y10416 , y10417 , y10418 , y10419 , y10420 , y10421 , y10422 , y10423 , y10424 , y10425 , y10426 , y10427 , y10428 , y10429 , y10430 , y10431 , y10432 , y10433 , y10434 , y10435 , y10436 , y10437 , y10438 , y10439 , y10440 , y10441 , y10442 , y10443 , y10444 , y10445 , y10446 , y10447 , y10448 , y10449 , y10450 , y10451 , y10452 , y10453 , y10454 , y10455 , y10456 , y10457 , y10458 , y10459 , y10460 , y10461 , y10462 , y10463 , y10464 , y10465 , y10466 , y10467 , y10468 , y10469 , y10470 , y10471 , y10472 , y10473 , y10474 , y10475 , y10476 , y10477 , y10478 , y10479 , y10480 , y10481 , y10482 , y10483 , y10484 , y10485 , y10486 , y10487 , y10488 , y10489 , y10490 , y10491 , y10492 , y10493 , y10494 , y10495 , y10496 , y10497 , y10498 , y10499 , y10500 , y10501 , y10502 , y10503 , y10504 , y10505 , y10506 , y10507 , y10508 , y10509 , y10510 , y10511 , y10512 , y10513 , y10514 , y10515 , y10516 , y10517 , y10518 , y10519 , y10520 , y10521 , y10522 , y10523 , y10524 , y10525 , y10526 , y10527 , y10528 , y10529 , y10530 , y10531 , y10532 , y10533 , y10534 , y10535 , y10536 , y10537 , y10538 , y10539 , y10540 , y10541 , y10542 , y10543 , y10544 , y10545 , y10546 , y10547 , y10548 , y10549 , y10550 , y10551 , y10552 , y10553 , y10554 , y10555 , y10556 , y10557 , y10558 , y10559 , y10560 , y10561 , y10562 , y10563 , y10564 , y10565 , y10566 , y10567 , y10568 , y10569 , y10570 , y10571 , y10572 , y10573 , y10574 , y10575 , y10576 , y10577 , y10578 , y10579 , y10580 , y10581 , y10582 , y10583 , y10584 , y10585 , y10586 , y10587 , y10588 , y10589 , y10590 , y10591 , y10592 , y10593 , y10594 , y10595 , y10596 , y10597 , y10598 , y10599 , y10600 , y10601 , y10602 , y10603 , y10604 , y10605 , y10606 , y10607 , y10608 , y10609 , y10610 , y10611 , y10612 , y10613 , y10614 , y10615 , y10616 , y10617 , y10618 , y10619 , y10620 , y10621 , y10622 , y10623 , y10624 , y10625 , y10626 , y10627 , y10628 , y10629 , y10630 , y10631 , y10632 , y10633 , y10634 , y10635 , y10636 , y10637 , y10638 , y10639 , y10640 , y10641 , y10642 , y10643 , y10644 , y10645 , y10646 , y10647 , y10648 , y10649 , y10650 , y10651 , y10652 , y10653 , y10654 , y10655 , y10656 , y10657 , y10658 , y10659 , y10660 , y10661 , y10662 , y10663 , y10664 , y10665 , y10666 , y10667 , y10668 , y10669 , y10670 , y10671 , y10672 , y10673 , y10674 , y10675 , y10676 , y10677 , y10678 , y10679 , y10680 , y10681 , y10682 , y10683 , y10684 , y10685 , y10686 , y10687 , y10688 , y10689 , y10690 , y10691 , y10692 , y10693 , y10694 , y10695 , y10696 , y10697 , y10698 , y10699 , y10700 , y10701 , y10702 , y10703 , y10704 , y10705 , y10706 , y10707 , y10708 , y10709 , y10710 , y10711 , y10712 , y10713 , y10714 , y10715 , y10716 , y10717 , y10718 , y10719 , y10720 , y10721 , y10722 , y10723 , y10724 , y10725 , y10726 , y10727 , y10728 , y10729 , y10730 , y10731 , y10732 , y10733 , y10734 , y10735 , y10736 , y10737 , y10738 , y10739 , y10740 , y10741 , y10742 , y10743 , y10744 , y10745 , y10746 , y10747 , y10748 , y10749 , y10750 , y10751 , y10752 , y10753 , y10754 , y10755 , y10756 , y10757 , y10758 , y10759 , y10760 , y10761 , y10762 , y10763 , y10764 , y10765 , y10766 , y10767 , y10768 , y10769 , y10770 , y10771 , y10772 , y10773 , y10774 , y10775 , y10776 , y10777 , y10778 , y10779 , y10780 , y10781 , y10782 , y10783 , y10784 , y10785 , y10786 , y10787 , y10788 , y10789 , y10790 , y10791 , y10792 , y10793 , y10794 , y10795 , y10796 , y10797 , y10798 , y10799 , y10800 , y10801 , y10802 , y10803 , y10804 , y10805 , y10806 , y10807 , y10808 , y10809 , y10810 , y10811 , y10812 , y10813 , y10814 , y10815 , y10816 , y10817 , y10818 , y10819 , y10820 , y10821 , y10822 , y10823 , y10824 , y10825 , y10826 , y10827 , y10828 , y10829 , y10830 , y10831 , y10832 , y10833 , y10834 , y10835 , y10836 , y10837 , y10838 , y10839 , y10840 , y10841 , y10842 , y10843 , y10844 , y10845 , y10846 , y10847 , y10848 , y10849 , y10850 , y10851 , y10852 , y10853 , y10854 , y10855 , y10856 , y10857 , y10858 , y10859 , y10860 , y10861 , y10862 , y10863 , y10864 , y10865 , y10866 , y10867 , y10868 , y10869 , y10870 , y10871 , y10872 , y10873 , y10874 , y10875 , y10876 , y10877 , y10878 , y10879 , y10880 , y10881 , y10882 , y10883 , y10884 , y10885 , y10886 , y10887 , y10888 , y10889 , y10890 , y10891 , y10892 , y10893 , y10894 , y10895 , y10896 , y10897 , y10898 , y10899 , y10900 , y10901 , y10902 , y10903 , y10904 , y10905 , y10906 , y10907 , y10908 , y10909 , y10910 , y10911 , y10912 , y10913 , y10914 , y10915 , y10916 , y10917 , y10918 , y10919 , y10920 , y10921 , y10922 , y10923 , y10924 , y10925 , y10926 , y10927 , y10928 , y10929 , y10930 , y10931 , y10932 , y10933 , y10934 , y10935 , y10936 , y10937 , y10938 , y10939 , y10940 , y10941 , y10942 , y10943 , y10944 , y10945 , y10946 , y10947 , y10948 , y10949 , y10950 , y10951 , y10952 , y10953 , y10954 , y10955 , y10956 , y10957 , y10958 , y10959 , y10960 , y10961 , y10962 , y10963 , y10964 , y10965 , y10966 , y10967 , y10968 , y10969 , y10970 , y10971 , y10972 , y10973 , y10974 , y10975 , y10976 , y10977 , y10978 , y10979 , y10980 , y10981 , y10982 , y10983 , y10984 , y10985 , y10986 , y10987 , y10988 , y10989 , y10990 , y10991 , y10992 , y10993 , y10994 , y10995 , y10996 , y10997 , y10998 , y10999 , y11000 , y11001 , y11002 , y11003 , y11004 , y11005 , y11006 , y11007 , y11008 , y11009 , y11010 , y11011 , y11012 , y11013 , y11014 , y11015 , y11016 , y11017 , y11018 , y11019 , y11020 , y11021 , y11022 , y11023 , y11024 , y11025 , y11026 , y11027 , y11028 , y11029 , y11030 , y11031 , y11032 , y11033 , y11034 , y11035 , y11036 , y11037 , y11038 , y11039 , y11040 , y11041 , y11042 , y11043 , y11044 , y11045 , y11046 , y11047 , y11048 , y11049 , y11050 , y11051 , y11052 , y11053 , y11054 , y11055 , y11056 , y11057 , y11058 , y11059 , y11060 , y11061 , y11062 , y11063 , y11064 , y11065 , y11066 , y11067 , y11068 , y11069 , y11070 , y11071 , y11072 , y11073 , y11074 , y11075 , y11076 , y11077 , y11078 , y11079 , y11080 , y11081 , y11082 , y11083 , y11084 , y11085 , y11086 , y11087 , y11088 , y11089 , y11090 , y11091 , y11092 , y11093 , y11094 , y11095 , y11096 , y11097 , y11098 , y11099 , y11100 , y11101 , y11102 , y11103 , y11104 , y11105 , y11106 , y11107 , y11108 , y11109 , y11110 , y11111 , y11112 , y11113 , y11114 , y11115 , y11116 , y11117 , y11118 , y11119 , y11120 , y11121 , y11122 , y11123 , y11124 , y11125 , y11126 , y11127 , y11128 , y11129 , y11130 , y11131 , y11132 , y11133 , y11134 , y11135 , y11136 , y11137 , y11138 , y11139 , y11140 , y11141 , y11142 , y11143 , y11144 , y11145 , y11146 , y11147 , y11148 , y11149 , y11150 , y11151 , y11152 , y11153 , y11154 , y11155 , y11156 , y11157 , y11158 , y11159 , y11160 , y11161 , y11162 , y11163 , y11164 , y11165 , y11166 , y11167 , y11168 , y11169 , y11170 , y11171 , y11172 , y11173 , y11174 , y11175 , y11176 , y11177 , y11178 , y11179 , y11180 , y11181 , y11182 , y11183 , y11184 , y11185 , y11186 , y11187 , y11188 , y11189 , y11190 , y11191 , y11192 , y11193 , y11194 , y11195 , y11196 , y11197 , y11198 , y11199 , y11200 , y11201 , y11202 , y11203 , y11204 , y11205 , y11206 , y11207 , y11208 , y11209 , y11210 , y11211 , y11212 , y11213 , y11214 , y11215 , y11216 , y11217 , y11218 , y11219 , y11220 , y11221 , y11222 , y11223 , y11224 , y11225 , y11226 , y11227 , y11228 , y11229 , y11230 , y11231 , y11232 , y11233 , y11234 , y11235 , y11236 , y11237 , y11238 , y11239 , y11240 , y11241 , y11242 , y11243 , y11244 , y11245 , y11246 , y11247 , y11248 , y11249 , y11250 , y11251 , y11252 , y11253 , y11254 , y11255 , y11256 , y11257 , y11258 , y11259 , y11260 , y11261 , y11262 , y11263 , y11264 , y11265 , y11266 , y11267 , y11268 , y11269 , y11270 , y11271 , y11272 , y11273 , y11274 , y11275 , y11276 , y11277 , y11278 , y11279 , y11280 , y11281 , y11282 , y11283 , y11284 , y11285 , y11286 , y11287 , y11288 , y11289 , y11290 , y11291 , y11292 , y11293 , y11294 , y11295 , y11296 , y11297 , y11298 , y11299 , y11300 , y11301 , y11302 , y11303 , y11304 , y11305 , y11306 , y11307 , y11308 , y11309 , y11310 , y11311 , y11312 , y11313 , y11314 , y11315 , y11316 , y11317 , y11318 , y11319 , y11320 , y11321 , y11322 , y11323 , y11324 , y11325 , y11326 , y11327 , y11328 , y11329 , y11330 , y11331 , y11332 , y11333 , y11334 , y11335 , y11336 , y11337 , y11338 , y11339 , y11340 , y11341 , y11342 , y11343 , y11344 , y11345 , y11346 , y11347 , y11348 , y11349 , y11350 , y11351 , y11352 , y11353 , y11354 , y11355 , y11356 , y11357 , y11358 , y11359 , y11360 , y11361 , y11362 , y11363 , y11364 , y11365 , y11366 , y11367 , y11368 , y11369 , y11370 , y11371 , y11372 , y11373 , y11374 , y11375 , y11376 , y11377 , y11378 , y11379 , y11380 , y11381 , y11382 , y11383 , y11384 , y11385 , y11386 , y11387 , y11388 , y11389 , y11390 , y11391 , y11392 , y11393 , y11394 , y11395 , y11396 , y11397 , y11398 , y11399 , y11400 , y11401 , y11402 , y11403 , y11404 , y11405 , y11406 , y11407 , y11408 , y11409 , y11410 , y11411 , y11412 , y11413 , y11414 , y11415 , y11416 , y11417 , y11418 , y11419 , y11420 , y11421 , y11422 , y11423 , y11424 , y11425 , y11426 , y11427 , y11428 , y11429 , y11430 , y11431 , y11432 , y11433 , y11434 , y11435 , y11436 , y11437 , y11438 , y11439 , y11440 , y11441 , y11442 , y11443 , y11444 , y11445 , y11446 , y11447 , y11448 , y11449 , y11450 , y11451 , y11452 , y11453 , y11454 , y11455 , y11456 , y11457 , y11458 , y11459 , y11460 , y11461 , y11462 , y11463 , y11464 , y11465 , y11466 , y11467 , y11468 , y11469 , y11470 , y11471 , y11472 , y11473 , y11474 , y11475 , y11476 , y11477 , y11478 , y11479 , y11480 , y11481 , y11482 , y11483 , y11484 , y11485 , y11486 , y11487 , y11488 , y11489 , y11490 , y11491 , y11492 , y11493 , y11494 , y11495 , y11496 , y11497 , y11498 , y11499 , y11500 , y11501 , y11502 , y11503 , y11504 , y11505 , y11506 , y11507 , y11508 , y11509 , y11510 , y11511 , y11512 , y11513 , y11514 , y11515 , y11516 , y11517 , y11518 , y11519 , y11520 , y11521 , y11522 , y11523 , y11524 , y11525 , y11526 , y11527 , y11528 , y11529 , y11530 , y11531 , y11532 , y11533 , y11534 , y11535 , y11536 , y11537 , y11538 , y11539 , y11540 , y11541 , y11542 , y11543 , y11544 , y11545 , y11546 , y11547 , y11548 , y11549 , y11550 , y11551 , y11552 , y11553 , y11554 , y11555 , y11556 , y11557 , y11558 , y11559 , y11560 , y11561 , y11562 , y11563 , y11564 , y11565 , y11566 , y11567 , y11568 , y11569 , y11570 , y11571 , y11572 , y11573 , y11574 , y11575 , y11576 , y11577 , y11578 , y11579 , y11580 , y11581 , y11582 , y11583 , y11584 , y11585 , y11586 , y11587 , y11588 , y11589 , y11590 , y11591 , y11592 , y11593 , y11594 , y11595 , y11596 , y11597 , y11598 , y11599 , y11600 , y11601 , y11602 , y11603 , y11604 , y11605 , y11606 , y11607 , y11608 , y11609 , y11610 , y11611 , y11612 , y11613 , y11614 , y11615 , y11616 , y11617 , y11618 , y11619 , y11620 , y11621 , y11622 , y11623 , y11624 , y11625 , y11626 , y11627 , y11628 , y11629 , y11630 , y11631 , y11632 , y11633 , y11634 , y11635 , y11636 , y11637 , y11638 , y11639 , y11640 , y11641 , y11642 , y11643 , y11644 , y11645 , y11646 , y11647 , y11648 , y11649 , y11650 , y11651 , y11652 , y11653 , y11654 , y11655 , y11656 , y11657 , y11658 , y11659 , y11660 , y11661 , y11662 , y11663 , y11664 , y11665 , y11666 , y11667 , y11668 , y11669 , y11670 , y11671 , y11672 , y11673 , y11674 , y11675 , y11676 , y11677 , y11678 , y11679 , y11680 , y11681 , y11682 , y11683 , y11684 , y11685 , y11686 , y11687 , y11688 , y11689 , y11690 , y11691 , y11692 , y11693 , y11694 , y11695 , y11696 , y11697 , y11698 , y11699 , y11700 , y11701 , y11702 , y11703 , y11704 , y11705 , y11706 , y11707 , y11708 , y11709 , y11710 , y11711 , y11712 , y11713 , y11714 , y11715 , y11716 , y11717 , y11718 , y11719 , y11720 , y11721 , y11722 , y11723 , y11724 , y11725 , y11726 , y11727 , y11728 , y11729 , y11730 , y11731 , y11732 , y11733 , y11734 , y11735 , y11736 , y11737 , y11738 , y11739 , y11740 , y11741 , y11742 , y11743 , y11744 , y11745 , y11746 , y11747 , y11748 , y11749 , y11750 , y11751 , y11752 , y11753 , y11754 , y11755 , y11756 , y11757 , y11758 , y11759 , y11760 , y11761 , y11762 , y11763 , y11764 , y11765 , y11766 , y11767 , y11768 , y11769 , y11770 , y11771 , y11772 , y11773 , y11774 , y11775 , y11776 , y11777 , y11778 , y11779 , y11780 , y11781 , y11782 , y11783 , y11784 , y11785 , y11786 , y11787 , y11788 , y11789 , y11790 , y11791 , y11792 , y11793 , y11794 , y11795 , y11796 , y11797 , y11798 , y11799 , y11800 , y11801 , y11802 , y11803 , y11804 , y11805 , y11806 , y11807 , y11808 , y11809 , y11810 , y11811 , y11812 , y11813 , y11814 , y11815 , y11816 , y11817 , y11818 , y11819 , y11820 , y11821 , y11822 , y11823 , y11824 , y11825 , y11826 , y11827 , y11828 , y11829 , y11830 , y11831 , y11832 , y11833 , y11834 , y11835 , y11836 , y11837 , y11838 , y11839 , y11840 , y11841 , y11842 , y11843 , y11844 , y11845 , y11846 , y11847 , y11848 , y11849 , y11850 , y11851 , y11852 , y11853 , y11854 , y11855 , y11856 , y11857 , y11858 , y11859 , y11860 , y11861 , y11862 , y11863 , y11864 , y11865 , y11866 , y11867 , y11868 , y11869 , y11870 , y11871 , y11872 , y11873 , y11874 , y11875 , y11876 , y11877 , y11878 , y11879 , y11880 , y11881 , y11882 , y11883 , y11884 , y11885 , y11886 , y11887 , y11888 , y11889 , y11890 , y11891 , y11892 , y11893 , y11894 , y11895 , y11896 , y11897 , y11898 , y11899 , y11900 , y11901 , y11902 , y11903 , y11904 , y11905 , y11906 , y11907 , y11908 , y11909 , y11910 , y11911 , y11912 , y11913 , y11914 , y11915 , y11916 , y11917 , y11918 , y11919 , y11920 , y11921 , y11922 , y11923 , y11924 , y11925 , y11926 , y11927 , y11928 , y11929 , y11930 , y11931 , y11932 , y11933 , y11934 , y11935 , y11936 , y11937 , y11938 , y11939 , y11940 , y11941 , y11942 , y11943 , y11944 , y11945 , y11946 , y11947 , y11948 , y11949 , y11950 , y11951 , y11952 , y11953 , y11954 , y11955 , y11956 , y11957 , y11958 , y11959 , y11960 , y11961 , y11962 , y11963 , y11964 , y11965 , y11966 , y11967 , y11968 , y11969 , y11970 , y11971 , y11972 , y11973 , y11974 , y11975 , y11976 , y11977 , y11978 , y11979 , y11980 , y11981 , y11982 , y11983 , y11984 , y11985 , y11986 , y11987 , y11988 , y11989 , y11990 , y11991 , y11992 , y11993 , y11994 , y11995 , y11996 , y11997 , y11998 , y11999 , y12000 , y12001 , y12002 , y12003 , y12004 , y12005 , y12006 , y12007 , y12008 , y12009 , y12010 , y12011 , y12012 , y12013 , y12014 , y12015 , y12016 , y12017 , y12018 , y12019 , y12020 , y12021 , y12022 , y12023 , y12024 , y12025 , y12026 , y12027 , y12028 , y12029 , y12030 , y12031 , y12032 , y12033 , y12034 , y12035 , y12036 , y12037 , y12038 , y12039 , y12040 , y12041 , y12042 , y12043 , y12044 , y12045 , y12046 , y12047 , y12048 , y12049 , y12050 , y12051 , y12052 , y12053 , y12054 , y12055 , y12056 , y12057 , y12058 , y12059 , y12060 , y12061 , y12062 , y12063 , y12064 , y12065 , y12066 , y12067 , y12068 , y12069 , y12070 , y12071 , y12072 , y12073 , y12074 , y12075 , y12076 , y12077 , y12078 , y12079 , y12080 , y12081 , y12082 , y12083 , y12084 , y12085 , y12086 , y12087 , y12088 , y12089 , y12090 , y12091 , y12092 , y12093 , y12094 , y12095 , y12096 , y12097 , y12098 , y12099 , y12100 , y12101 , y12102 , y12103 , y12104 , y12105 , y12106 , y12107 , y12108 , y12109 , y12110 , y12111 , y12112 , y12113 , y12114 , y12115 , y12116 , y12117 , y12118 , y12119 , y12120 , y12121 , y12122 , y12123 , y12124 , y12125 , y12126 , y12127 , y12128 , y12129 , y12130 , y12131 , y12132 , y12133 , y12134 , y12135 , y12136 , y12137 , y12138 , y12139 , y12140 , y12141 , y12142 , y12143 , y12144 , y12145 , y12146 , y12147 , y12148 , y12149 , y12150 , y12151 , y12152 , y12153 , y12154 , y12155 , y12156 , y12157 , y12158 , y12159 , y12160 , y12161 , y12162 , y12163 , y12164 , y12165 , y12166 , y12167 , y12168 , y12169 , y12170 , y12171 , y12172 , y12173 , y12174 , y12175 , y12176 , y12177 , y12178 , y12179 , y12180 , y12181 , y12182 , y12183 , y12184 , y12185 , y12186 , y12187 , y12188 , y12189 , y12190 , y12191 , y12192 , y12193 , y12194 , y12195 , y12196 , y12197 , y12198 , y12199 , y12200 , y12201 , y12202 , y12203 , y12204 , y12205 , y12206 , y12207 , y12208 , y12209 , y12210 , y12211 , y12212 , y12213 , y12214 , y12215 , y12216 , y12217 , y12218 , y12219 , y12220 , y12221 , y12222 , y12223 , y12224 , y12225 , y12226 , y12227 , y12228 , y12229 , y12230 , y12231 , y12232 , y12233 , y12234 , y12235 , y12236 , y12237 , y12238 , y12239 , y12240 , y12241 , y12242 , y12243 , y12244 , y12245 , y12246 , y12247 , y12248 , y12249 , y12250 , y12251 , y12252 , y12253 , y12254 , y12255 , y12256 , y12257 , y12258 , y12259 , y12260 , y12261 , y12262 , y12263 , y12264 , y12265 , y12266 , y12267 , y12268 , y12269 , y12270 , y12271 , y12272 , y12273 , y12274 , y12275 , y12276 , y12277 , y12278 , y12279 , y12280 , y12281 , y12282 , y12283 , y12284 , y12285 , y12286 , y12287 , y12288 , y12289 , y12290 , y12291 , y12292 , y12293 , y12294 , y12295 , y12296 , y12297 , y12298 , y12299 , y12300 , y12301 , y12302 , y12303 , y12304 , y12305 , y12306 , y12307 , y12308 , y12309 , y12310 , y12311 , y12312 , y12313 , y12314 , y12315 , y12316 , y12317 , y12318 , y12319 , y12320 , y12321 , y12322 , y12323 , y12324 , y12325 , y12326 , y12327 , y12328 , y12329 , y12330 , y12331 , y12332 , y12333 , y12334 , y12335 , y12336 , y12337 , y12338 , y12339 , y12340 , y12341 , y12342 , y12343 , y12344 , y12345 , y12346 , y12347 , y12348 , y12349 , y12350 , y12351 , y12352 , y12353 , y12354 , y12355 , y12356 , y12357 , y12358 , y12359 , y12360 , y12361 , y12362 , y12363 , y12364 , y12365 , y12366 , y12367 , y12368 , y12369 , y12370 , y12371 , y12372 , y12373 , y12374 , y12375 , y12376 , y12377 , y12378 , y12379 , y12380 , y12381 , y12382 , y12383 , y12384 , y12385 , y12386 , y12387 , y12388 , y12389 , y12390 , y12391 , y12392 , y12393 , y12394 , y12395 , y12396 , y12397 , y12398 , y12399 , y12400 , y12401 , y12402 , y12403 , y12404 , y12405 , y12406 , y12407 , y12408 , y12409 , y12410 , y12411 , y12412 , y12413 , y12414 , y12415 , y12416 , y12417 , y12418 , y12419 , y12420 , y12421 , y12422 , y12423 , y12424 , y12425 , y12426 , y12427 , y12428 , y12429 , y12430 , y12431 , y12432 , y12433 , y12434 , y12435 , y12436 , y12437 , y12438 , y12439 , y12440 , y12441 , y12442 , y12443 , y12444 , y12445 , y12446 , y12447 , y12448 , y12449 , y12450 , y12451 , y12452 , y12453 , y12454 , y12455 , y12456 , y12457 , y12458 , y12459 , y12460 , y12461 , y12462 , y12463 , y12464 , y12465 , y12466 , y12467 , y12468 , y12469 , y12470 , y12471 , y12472 , y12473 , y12474 , y12475 , y12476 , y12477 , y12478 , y12479 , y12480 , y12481 , y12482 , y12483 , y12484 , y12485 , y12486 , y12487 , y12488 , y12489 , y12490 , y12491 , y12492 , y12493 , y12494 , y12495 , y12496 , y12497 , y12498 , y12499 , y12500 , y12501 , y12502 , y12503 , y12504 , y12505 , y12506 , y12507 , y12508 , y12509 , y12510 , y12511 , y12512 , y12513 , y12514 , y12515 , y12516 , y12517 , y12518 , y12519 , y12520 , y12521 , y12522 , y12523 , y12524 , y12525 , y12526 , y12527 , y12528 , y12529 , y12530 , y12531 , y12532 , y12533 , y12534 , y12535 , y12536 , y12537 , y12538 , y12539 , y12540 , y12541 , y12542 , y12543 , y12544 , y12545 , y12546 , y12547 , y12548 , y12549 , y12550 , y12551 , y12552 , y12553 , y12554 , y12555 , y12556 , y12557 , y12558 , y12559 , y12560 , y12561 , y12562 , y12563 , y12564 , y12565 , y12566 , y12567 , y12568 , y12569 , y12570 , y12571 , y12572 , y12573 , y12574 , y12575 , y12576 , y12577 , y12578 , y12579 , y12580 , y12581 , y12582 , y12583 , y12584 , y12585 , y12586 , y12587 , y12588 , y12589 , y12590 , y12591 , y12592 , y12593 , y12594 , y12595 , y12596 , y12597 , y12598 , y12599 , y12600 , y12601 , y12602 , y12603 , y12604 , y12605 , y12606 , y12607 , y12608 , y12609 , y12610 , y12611 , y12612 , y12613 , y12614 , y12615 , y12616 , y12617 , y12618 , y12619 , y12620 , y12621 , y12622 , y12623 , y12624 , y12625 , y12626 , y12627 , y12628 , y12629 , y12630 , y12631 , y12632 , y12633 , y12634 , y12635 , y12636 , y12637 , y12638 , y12639 , y12640 , y12641 , y12642 , y12643 , y12644 , y12645 , y12646 , y12647 , y12648 , y12649 , y12650 , y12651 , y12652 , y12653 , y12654 , y12655 , y12656 , y12657 , y12658 , y12659 , y12660 , y12661 , y12662 , y12663 , y12664 , y12665 , y12666 , y12667 , y12668 , y12669 , y12670 , y12671 , y12672 , y12673 , y12674 , y12675 , y12676 , y12677 , y12678 , y12679 , y12680 , y12681 , y12682 , y12683 , y12684 , y12685 , y12686 , y12687 , y12688 , y12689 , y12690 , y12691 , y12692 , y12693 , y12694 , y12695 , y12696 , y12697 , y12698 , y12699 , y12700 , y12701 , y12702 , y12703 , y12704 , y12705 , y12706 , y12707 , y12708 , y12709 , y12710 , y12711 , y12712 , y12713 , y12714 , y12715 , y12716 , y12717 , y12718 , y12719 , y12720 , y12721 , y12722 , y12723 , y12724 , y12725 , y12726 , y12727 , y12728 , y12729 , y12730 , y12731 , y12732 , y12733 , y12734 , y12735 , y12736 , y12737 , y12738 , y12739 , y12740 , y12741 , y12742 , y12743 , y12744 , y12745 , y12746 , y12747 , y12748 , y12749 , y12750 , y12751 , y12752 , y12753 , y12754 , y12755 , y12756 , y12757 , y12758 , y12759 , y12760 , y12761 , y12762 , y12763 , y12764 , y12765 , y12766 , y12767 , y12768 , y12769 , y12770 , y12771 , y12772 , y12773 , y12774 , y12775 , y12776 , y12777 , y12778 , y12779 , y12780 , y12781 , y12782 , y12783 , y12784 , y12785 , y12786 , y12787 , y12788 , y12789 , y12790 , y12791 , y12792 , y12793 , y12794 , y12795 , y12796 , y12797 , y12798 , y12799 , y12800 , y12801 , y12802 , y12803 , y12804 , y12805 , y12806 , y12807 , y12808 , y12809 , y12810 , y12811 , y12812 , y12813 , y12814 , y12815 , y12816 , y12817 , y12818 , y12819 , y12820 , y12821 , y12822 , y12823 , y12824 , y12825 , y12826 , y12827 , y12828 , y12829 , y12830 , y12831 , y12832 , y12833 , y12834 , y12835 , y12836 , y12837 , y12838 , y12839 , y12840 , y12841 , y12842 , y12843 , y12844 , y12845 , y12846 , y12847 , y12848 , y12849 , y12850 , y12851 , y12852 , y12853 , y12854 , y12855 , y12856 , y12857 , y12858 , y12859 , y12860 , y12861 , y12862 , y12863 , y12864 , y12865 , y12866 , y12867 , y12868 , y12869 , y12870 , y12871 , y12872 , y12873 , y12874 , y12875 , y12876 , y12877 , y12878 , y12879 , y12880 , y12881 , y12882 , y12883 , y12884 , y12885 , y12886 , y12887 , y12888 , y12889 , y12890 , y12891 , y12892 , y12893 , y12894 , y12895 , y12896 , y12897 , y12898 , y12899 , y12900 , y12901 , y12902 , y12903 , y12904 , y12905 , y12906 , y12907 , y12908 , y12909 , y12910 , y12911 , y12912 , y12913 , y12914 , y12915 , y12916 , y12917 , y12918 , y12919 , y12920 , y12921 , y12922 , y12923 , y12924 , y12925 , y12926 , y12927 , y12928 , y12929 , y12930 , y12931 , y12932 , y12933 , y12934 , y12935 , y12936 , y12937 , y12938 , y12939 , y12940 , y12941 , y12942 , y12943 , y12944 , y12945 , y12946 , y12947 , y12948 , y12949 , y12950 , y12951 , y12952 , y12953 , y12954 , y12955 , y12956 , y12957 , y12958 , y12959 , y12960 , y12961 , y12962 , y12963 , y12964 , y12965 , y12966 , y12967 , y12968 , y12969 , y12970 , y12971 , y12972 , y12973 , y12974 , y12975 , y12976 , y12977 , y12978 , y12979 , y12980 , y12981 , y12982 , y12983 , y12984 , y12985 , y12986 , y12987 , y12988 , y12989 , y12990 , y12991 , y12992 , y12993 , y12994 , y12995 , y12996 , y12997 , y12998 , y12999 , y13000 , y13001 , y13002 , y13003 , y13004 , y13005 , y13006 , y13007 , y13008 , y13009 , y13010 , y13011 , y13012 , y13013 , y13014 , y13015 , y13016 , y13017 , y13018 , y13019 , y13020 , y13021 , y13022 , y13023 , y13024 , y13025 , y13026 , y13027 , y13028 , y13029 , y13030 , y13031 , y13032 , y13033 , y13034 , y13035 , y13036 , y13037 , y13038 , y13039 , y13040 , y13041 , y13042 , y13043 , y13044 , y13045 , y13046 , y13047 , y13048 , y13049 , y13050 , y13051 , y13052 , y13053 , y13054 , y13055 , y13056 , y13057 , y13058 , y13059 , y13060 , y13061 , y13062 , y13063 , y13064 , y13065 , y13066 , y13067 , y13068 , y13069 , y13070 , y13071 , y13072 , y13073 , y13074 , y13075 , y13076 , y13077 , y13078 , y13079 , y13080 , y13081 , y13082 , y13083 , y13084 , y13085 , y13086 , y13087 , y13088 , y13089 , y13090 , y13091 , y13092 , y13093 , y13094 , y13095 , y13096 , y13097 , y13098 , y13099 , y13100 , y13101 , y13102 , y13103 , y13104 , y13105 , y13106 , y13107 , y13108 , y13109 , y13110 , y13111 , y13112 , y13113 , y13114 , y13115 , y13116 , y13117 , y13118 , y13119 , y13120 , y13121 , y13122 , y13123 , y13124 , y13125 , y13126 , y13127 , y13128 , y13129 , y13130 , y13131 , y13132 , y13133 , y13134 , y13135 , y13136 , y13137 , y13138 , y13139 , y13140 , y13141 , y13142 , y13143 , y13144 , y13145 , y13146 , y13147 , y13148 , y13149 , y13150 , y13151 , y13152 , y13153 , y13154 , y13155 , y13156 , y13157 , y13158 , y13159 , y13160 , y13161 , y13162 , y13163 , y13164 , y13165 , y13166 , y13167 , y13168 , y13169 , y13170 , y13171 , y13172 , y13173 , y13174 , y13175 , y13176 , y13177 , y13178 , y13179 , y13180 , y13181 , y13182 , y13183 , y13184 , y13185 , y13186 , y13187 , y13188 , y13189 , y13190 , y13191 , y13192 , y13193 , y13194 , y13195 , y13196 , y13197 , y13198 , y13199 , y13200 , y13201 , y13202 , y13203 , y13204 , y13205 , y13206 , y13207 , y13208 , y13209 , y13210 , y13211 , y13212 , y13213 , y13214 , y13215 , y13216 , y13217 , y13218 , y13219 , y13220 , y13221 , y13222 , y13223 , y13224 , y13225 , y13226 , y13227 , y13228 , y13229 , y13230 , y13231 , y13232 , y13233 , y13234 , y13235 , y13236 , y13237 , y13238 , y13239 , y13240 , y13241 , y13242 , y13243 , y13244 , y13245 , y13246 , y13247 , y13248 , y13249 , y13250 , y13251 , y13252 , y13253 , y13254 , y13255 , y13256 , y13257 , y13258 , y13259 , y13260 , y13261 , y13262 , y13263 , y13264 , y13265 , y13266 , y13267 , y13268 , y13269 , y13270 , y13271 , y13272 , y13273 , y13274 , y13275 , y13276 , y13277 , y13278 , y13279 , y13280 , y13281 , y13282 , y13283 , y13284 , y13285 , y13286 , y13287 , y13288 , y13289 , y13290 , y13291 , y13292 , y13293 , y13294 , y13295 , y13296 , y13297 , y13298 , y13299 , y13300 , y13301 , y13302 , y13303 , y13304 , y13305 , y13306 , y13307 , y13308 , y13309 , y13310 , y13311 , y13312 , y13313 , y13314 , y13315 , y13316 , y13317 , y13318 , y13319 , y13320 , y13321 , y13322 , y13323 , y13324 , y13325 , y13326 , y13327 , y13328 , y13329 , y13330 , y13331 , y13332 , y13333 , y13334 , y13335 , y13336 , y13337 , y13338 , y13339 , y13340 , y13341 , y13342 , y13343 , y13344 , y13345 , y13346 , y13347 , y13348 , y13349 , y13350 , y13351 , y13352 , y13353 , y13354 , y13355 , y13356 , y13357 , y13358 , y13359 , y13360 , y13361 , y13362 , y13363 , y13364 , y13365 , y13366 , y13367 , y13368 , y13369 , y13370 , y13371 , y13372 , y13373 , y13374 , y13375 , y13376 , y13377 , y13378 , y13379 , y13380 , y13381 , y13382 , y13383 , y13384 , y13385 , y13386 , y13387 , y13388 , y13389 , y13390 , y13391 , y13392 , y13393 , y13394 , y13395 , y13396 , y13397 , y13398 , y13399 , y13400 , y13401 , y13402 , y13403 , y13404 , y13405 , y13406 , y13407 , y13408 , y13409 , y13410 , y13411 , y13412 , y13413 , y13414 , y13415 , y13416 , y13417 , y13418 , y13419 , y13420 , y13421 , y13422 , y13423 , y13424 , y13425 , y13426 , y13427 , y13428 , y13429 , y13430 , y13431 , y13432 , y13433 , y13434 , y13435 , y13436 , y13437 , y13438 , y13439 , y13440 , y13441 , y13442 , y13443 , y13444 , y13445 , y13446 , y13447 , y13448 , y13449 , y13450 , y13451 , y13452 , y13453 , y13454 , y13455 , y13456 , y13457 , y13458 , y13459 , y13460 , y13461 , y13462 , y13463 , y13464 , y13465 , y13466 , y13467 , y13468 , y13469 , y13470 , y13471 , y13472 , y13473 , y13474 , y13475 , y13476 , y13477 , y13478 , y13479 , y13480 , y13481 , y13482 , y13483 , y13484 , y13485 , y13486 , y13487 , y13488 , y13489 , y13490 , y13491 , y13492 , y13493 , y13494 , y13495 , y13496 , y13497 , y13498 , y13499 , y13500 , y13501 , y13502 , y13503 , y13504 , y13505 , y13506 , y13507 , y13508 , y13509 , y13510 , y13511 , y13512 , y13513 , y13514 , y13515 , y13516 , y13517 , y13518 , y13519 , y13520 , y13521 , y13522 , y13523 , y13524 , y13525 , y13526 , y13527 , y13528 , y13529 , y13530 , y13531 , y13532 , y13533 , y13534 , y13535 , y13536 , y13537 , y13538 , y13539 , y13540 , y13541 , y13542 , y13543 , y13544 , y13545 , y13546 , y13547 , y13548 , y13549 , y13550 , y13551 , y13552 , y13553 , y13554 , y13555 , y13556 , y13557 , y13558 , y13559 , y13560 , y13561 , y13562 , y13563 , y13564 , y13565 , y13566 , y13567 , y13568 , y13569 , y13570 , y13571 , y13572 , y13573 , y13574 , y13575 , y13576 , y13577 , y13578 , y13579 , y13580 , y13581 , y13582 , y13583 , y13584 , y13585 , y13586 , y13587 , y13588 , y13589 , y13590 , y13591 , y13592 , y13593 , y13594 , y13595 , y13596 , y13597 , y13598 , y13599 , y13600 , y13601 , y13602 , y13603 , y13604 , y13605 , y13606 , y13607 , y13608 , y13609 , y13610 , y13611 , y13612 , y13613 , y13614 , y13615 , y13616 , y13617 , y13618 , y13619 , y13620 , y13621 , y13622 , y13623 , y13624 , y13625 , y13626 , y13627 , y13628 , y13629 , y13630 , y13631 , y13632 , y13633 , y13634 , y13635 , y13636 , y13637 , y13638 , y13639 , y13640 , y13641 , y13642 , y13643 , y13644 , y13645 , y13646 , y13647 , y13648 , y13649 , y13650 , y13651 , y13652 , y13653 , y13654 , y13655 , y13656 , y13657 , y13658 , y13659 , y13660 , y13661 , y13662 , y13663 , y13664 , y13665 , y13666 , y13667 , y13668 , y13669 , y13670 , y13671 , y13672 , y13673 , y13674 , y13675 , y13676 , y13677 , y13678 , y13679 , y13680 , y13681 , y13682 , y13683 , y13684 , y13685 , y13686 , y13687 , y13688 , y13689 , y13690 , y13691 , y13692 , y13693 , y13694 , y13695 , y13696 , y13697 , y13698 , y13699 , y13700 , y13701 , y13702 , y13703 , y13704 , y13705 , y13706 , y13707 , y13708 , y13709 , y13710 , y13711 , y13712 , y13713 , y13714 , y13715 , y13716 , y13717 , y13718 , y13719 , y13720 , y13721 , y13722 , y13723 , y13724 , y13725 , y13726 , y13727 , y13728 , y13729 , y13730 , y13731 , y13732 , y13733 , y13734 , y13735 , y13736 , y13737 , y13738 , y13739 , y13740 , y13741 , y13742 , y13743 , y13744 , y13745 , y13746 , y13747 , y13748 , y13749 , y13750 , y13751 , y13752 , y13753 , y13754 , y13755 , y13756 , y13757 , y13758 , y13759 , y13760 , y13761 , y13762 , y13763 , y13764 , y13765 , y13766 , y13767 , y13768 , y13769 , y13770 , y13771 , y13772 , y13773 , y13774 , y13775 , y13776 , y13777 , y13778 , y13779 , y13780 , y13781 , y13782 , y13783 , y13784 , y13785 , y13786 , y13787 , y13788 , y13789 , y13790 , y13791 , y13792 , y13793 , y13794 , y13795 , y13796 , y13797 , y13798 , y13799 , y13800 , y13801 , y13802 , y13803 , y13804 , y13805 , y13806 , y13807 , y13808 , y13809 , y13810 , y13811 , y13812 , y13813 , y13814 , y13815 , y13816 , y13817 , y13818 , y13819 , y13820 , y13821 , y13822 , y13823 , y13824 , y13825 , y13826 , y13827 , y13828 , y13829 , y13830 , y13831 , y13832 , y13833 , y13834 , y13835 , y13836 , y13837 , y13838 , y13839 , y13840 , y13841 , y13842 , y13843 , y13844 , y13845 , y13846 , y13847 , y13848 , y13849 , y13850 , y13851 , y13852 , y13853 , y13854 , y13855 , y13856 , y13857 , y13858 , y13859 , y13860 , y13861 , y13862 , y13863 , y13864 , y13865 , y13866 , y13867 , y13868 , y13869 , y13870 , y13871 , y13872 , y13873 , y13874 , y13875 , y13876 , y13877 , y13878 , y13879 , y13880 , y13881 , y13882 , y13883 , y13884 , y13885 , y13886 , y13887 , y13888 , y13889 , y13890 , y13891 , y13892 , y13893 , y13894 , y13895 , y13896 , y13897 , y13898 , y13899 , y13900 , y13901 , y13902 , y13903 , y13904 , y13905 , y13906 , y13907 , y13908 , y13909 , y13910 , y13911 , y13912 , y13913 , y13914 , y13915 , y13916 , y13917 , y13918 , y13919 , y13920 , y13921 , y13922 , y13923 , y13924 , y13925 , y13926 , y13927 , y13928 , y13929 , y13930 , y13931 , y13932 , y13933 , y13934 , y13935 , y13936 , y13937 , y13938 , y13939 , y13940 , y13941 , y13942 , y13943 , y13944 , y13945 , y13946 , y13947 , y13948 , y13949 , y13950 , y13951 , y13952 , y13953 , y13954 , y13955 , y13956 , y13957 , y13958 , y13959 , y13960 , y13961 , y13962 , y13963 , y13964 , y13965 , y13966 , y13967 , y13968 , y13969 , y13970 , y13971 , y13972 , y13973 , y13974 , y13975 , y13976 , y13977 , y13978 , y13979 , y13980 , y13981 , y13982 , y13983 , y13984 , y13985 , y13986 , y13987 , y13988 , y13989 , y13990 , y13991 , y13992 , y13993 , y13994 , y13995 , y13996 , y13997 , y13998 , y13999 , y14000 , y14001 , y14002 , y14003 , y14004 , y14005 , y14006 , y14007 , y14008 , y14009 , y14010 , y14011 , y14012 , y14013 , y14014 , y14015 , y14016 , y14017 , y14018 , y14019 , y14020 , y14021 , y14022 , y14023 , y14024 , y14025 , y14026 , y14027 , y14028 , y14029 , y14030 , y14031 , y14032 , y14033 , y14034 , y14035 , y14036 , y14037 , y14038 , y14039 , y14040 , y14041 , y14042 , y14043 , y14044 , y14045 , y14046 , y14047 , y14048 , y14049 , y14050 , y14051 , y14052 , y14053 , y14054 , y14055 , y14056 , y14057 , y14058 , y14059 , y14060 , y14061 , y14062 , y14063 , y14064 , y14065 , y14066 , y14067 , y14068 , y14069 , y14070 , y14071 , y14072 , y14073 , y14074 , y14075 , y14076 , y14077 , y14078 , y14079 , y14080 , y14081 , y14082 , y14083 , y14084 , y14085 , y14086 , y14087 , y14088 , y14089 , y14090 , y14091 , y14092 , y14093 , y14094 , y14095 , y14096 , y14097 , y14098 , y14099 , y14100 , y14101 , y14102 , y14103 , y14104 , y14105 , y14106 , y14107 , y14108 , y14109 , y14110 , y14111 , y14112 , y14113 , y14114 , y14115 , y14116 , y14117 , y14118 , y14119 , y14120 , y14121 , y14122 , y14123 , y14124 , y14125 , y14126 , y14127 , y14128 , y14129 , y14130 , y14131 , y14132 , y14133 , y14134 , y14135 , y14136 , y14137 , y14138 , y14139 , y14140 , y14141 , y14142 , y14143 , y14144 , y14145 , y14146 , y14147 , y14148 , y14149 , y14150 , y14151 , y14152 , y14153 , y14154 , y14155 , y14156 , y14157 , y14158 , y14159 , y14160 , y14161 , y14162 , y14163 , y14164 , y14165 , y14166 , y14167 , y14168 , y14169 , y14170 , y14171 , y14172 , y14173 , y14174 , y14175 , y14176 , y14177 , y14178 , y14179 , y14180 , y14181 , y14182 , y14183 , y14184 , y14185 , y14186 , y14187 , y14188 , y14189 , y14190 , y14191 , y14192 , y14193 , y14194 , y14195 , y14196 , y14197 , y14198 , y14199 , y14200 , y14201 , y14202 , y14203 , y14204 , y14205 , y14206 , y14207 , y14208 , y14209 , y14210 , y14211 , y14212 , y14213 , y14214 , y14215 , y14216 , y14217 , y14218 , y14219 , y14220 , y14221 , y14222 , y14223 , y14224 , y14225 , y14226 , y14227 , y14228 , y14229 , y14230 , y14231 , y14232 , y14233 , y14234 , y14235 , y14236 , y14237 , y14238 , y14239 , y14240 , y14241 , y14242 , y14243 , y14244 , y14245 , y14246 , y14247 , y14248 , y14249 , y14250 , y14251 , y14252 , y14253 , y14254 , y14255 , y14256 , y14257 , y14258 , y14259 , y14260 , y14261 , y14262 , y14263 , y14264 , y14265 , y14266 , y14267 , y14268 , y14269 , y14270 , y14271 , y14272 , y14273 , y14274 , y14275 , y14276 , y14277 , y14278 , y14279 , y14280 , y14281 , y14282 , y14283 , y14284 , y14285 , y14286 , y14287 , y14288 , y14289 , y14290 , y14291 , y14292 , y14293 , y14294 , y14295 , y14296 , y14297 , y14298 , y14299 , y14300 , y14301 , y14302 , y14303 , y14304 , y14305 , y14306 , y14307 , y14308 , y14309 , y14310 , y14311 , y14312 , y14313 , y14314 , y14315 , y14316 , y14317 , y14318 , y14319 , y14320 , y14321 , y14322 , y14323 , y14324 , y14325 , y14326 , y14327 , y14328 , y14329 , y14330 , y14331 , y14332 , y14333 , y14334 , y14335 , y14336 , y14337 , y14338 , y14339 , y14340 , y14341 , y14342 , y14343 , y14344 , y14345 , y14346 , y14347 , y14348 , y14349 , y14350 , y14351 , y14352 , y14353 , y14354 , y14355 , y14356 , y14357 , y14358 , y14359 , y14360 , y14361 , y14362 , y14363 , y14364 , y14365 , y14366 , y14367 , y14368 , y14369 , y14370 , y14371 , y14372 , y14373 , y14374 , y14375 , y14376 , y14377 , y14378 , y14379 , y14380 , y14381 , y14382 , y14383 , y14384 , y14385 , y14386 , y14387 , y14388 , y14389 , y14390 , y14391 , y14392 , y14393 , y14394 , y14395 , y14396 , y14397 , y14398 , y14399 , y14400 , y14401 , y14402 , y14403 , y14404 , y14405 , y14406 , y14407 , y14408 , y14409 , y14410 , y14411 , y14412 , y14413 , y14414 , y14415 , y14416 , y14417 , y14418 , y14419 , y14420 , y14421 , y14422 , y14423 , y14424 , y14425 , y14426 , y14427 , y14428 , y14429 , y14430 , y14431 , y14432 , y14433 , y14434 , y14435 , y14436 , y14437 , y14438 , y14439 , y14440 , y14441 , y14442 , y14443 , y14444 , y14445 , y14446 , y14447 , y14448 , y14449 , y14450 , y14451 , y14452 , y14453 , y14454 , y14455 , y14456 , y14457 , y14458 , y14459 , y14460 , y14461 , y14462 , y14463 , y14464 , y14465 , y14466 , y14467 , y14468 , y14469 , y14470 , y14471 , y14472 , y14473 , y14474 , y14475 , y14476 , y14477 , y14478 , y14479 , y14480 , y14481 , y14482 , y14483 , y14484 , y14485 , y14486 , y14487 , y14488 , y14489 , y14490 , y14491 , y14492 , y14493 , y14494 , y14495 , y14496 , y14497 , y14498 , y14499 , y14500 , y14501 , y14502 , y14503 , y14504 , y14505 , y14506 , y14507 , y14508 , y14509 , y14510 , y14511 , y14512 , y14513 , y14514 , y14515 , y14516 , y14517 , y14518 , y14519 , y14520 , y14521 , y14522 , y14523 , y14524 , y14525 , y14526 , y14527 , y14528 , y14529 , y14530 , y14531 , y14532 , y14533 , y14534 , y14535 , y14536 , y14537 , y14538 , y14539 , y14540 , y14541 , y14542 , y14543 , y14544 , y14545 , y14546 , y14547 , y14548 , y14549 , y14550 , y14551 , y14552 , y14553 , y14554 , y14555 , y14556 , y14557 , y14558 , y14559 , y14560 , y14561 , y14562 , y14563 , y14564 , y14565 , y14566 , y14567 , y14568 , y14569 , y14570 , y14571 , y14572 , y14573 , y14574 , y14575 , y14576 , y14577 , y14578 , y14579 , y14580 , y14581 , y14582 , y14583 , y14584 , y14585 , y14586 , y14587 , y14588 , y14589 , y14590 , y14591 , y14592 , y14593 , y14594 , y14595 , y14596 , y14597 , y14598 , y14599 , y14600 , y14601 , y14602 , y14603 , y14604 , y14605 , y14606 , y14607 , y14608 , y14609 , y14610 , y14611 , y14612 , y14613 , y14614 , y14615 , y14616 , y14617 , y14618 , y14619 , y14620 , y14621 , y14622 , y14623 , y14624 , y14625 , y14626 , y14627 , y14628 , y14629 , y14630 , y14631 , y14632 , y14633 , y14634 , y14635 , y14636 , y14637 , y14638 , y14639 , y14640 , y14641 , y14642 , y14643 , y14644 , y14645 , y14646 , y14647 , y14648 , y14649 , y14650 , y14651 , y14652 , y14653 , y14654 , y14655 , y14656 , y14657 , y14658 , y14659 , y14660 , y14661 , y14662 , y14663 , y14664 , y14665 , y14666 , y14667 , y14668 , y14669 , y14670 , y14671 , y14672 , y14673 , y14674 , y14675 , y14676 , y14677 , y14678 , y14679 , y14680 , y14681 , y14682 , y14683 , y14684 , y14685 , y14686 , y14687 , y14688 , y14689 , y14690 , y14691 , y14692 , y14693 , y14694 , y14695 , y14696 , y14697 , y14698 , y14699 , y14700 , y14701 , y14702 , y14703 , y14704 , y14705 , y14706 , y14707 , y14708 , y14709 , y14710 , y14711 , y14712 , y14713 , y14714 , y14715 , y14716 , y14717 , y14718 , y14719 , y14720 , y14721 , y14722 , y14723 , y14724 , y14725 , y14726 , y14727 , y14728 , y14729 , y14730 , y14731 , y14732 , y14733 , y14734 , y14735 , y14736 , y14737 , y14738 , y14739 , y14740 , y14741 , y14742 , y14743 , y14744 , y14745 , y14746 , y14747 , y14748 , y14749 , y14750 , y14751 , y14752 , y14753 , y14754 , y14755 , y14756 , y14757 , y14758 , y14759 , y14760 , y14761 , y14762 , y14763 , y14764 , y14765 , y14766 , y14767 , y14768 , y14769 , y14770 , y14771 , y14772 , y14773 , y14774 , y14775 , y14776 , y14777 , y14778 , y14779 , y14780 , y14781 , y14782 , y14783 , y14784 , y14785 , y14786 , y14787 , y14788 , y14789 , y14790 , y14791 , y14792 , y14793 , y14794 , y14795 , y14796 , y14797 , y14798 , y14799 , y14800 , y14801 , y14802 , y14803 , y14804 , y14805 , y14806 , y14807 , y14808 , y14809 , y14810 , y14811 , y14812 , y14813 , y14814 , y14815 , y14816 , y14817 , y14818 , y14819 , y14820 , y14821 , y14822 , y14823 , y14824 , y14825 , y14826 , y14827 , y14828 , y14829 , y14830 , y14831 , y14832 , y14833 , y14834 , y14835 , y14836 , y14837 , y14838 , y14839 , y14840 , y14841 , y14842 , y14843 , y14844 , y14845 , y14846 , y14847 , y14848 , y14849 , y14850 , y14851 , y14852 , y14853 , y14854 , y14855 , y14856 , y14857 , y14858 , y14859 , y14860 , y14861 , y14862 , y14863 , y14864 , y14865 , y14866 , y14867 , y14868 , y14869 , y14870 , y14871 , y14872 , y14873 , y14874 , y14875 , y14876 , y14877 , y14878 , y14879 , y14880 , y14881 , y14882 , y14883 , y14884 , y14885 , y14886 , y14887 , y14888 , y14889 , y14890 , y14891 , y14892 , y14893 , y14894 , y14895 , y14896 , y14897 , y14898 , y14899 , y14900 , y14901 , y14902 , y14903 , y14904 , y14905 , y14906 , y14907 , y14908 , y14909 , y14910 , y14911 , y14912 , y14913 , y14914 , y14915 , y14916 , y14917 , y14918 , y14919 , y14920 , y14921 , y14922 , y14923 , y14924 , y14925 , y14926 , y14927 , y14928 , y14929 , y14930 , y14931 , y14932 , y14933 , y14934 , y14935 , y14936 , y14937 , y14938 , y14939 , y14940 , y14941 , y14942 , y14943 , y14944 , y14945 , y14946 , y14947 , y14948 , y14949 , y14950 , y14951 , y14952 , y14953 , y14954 , y14955 , y14956 , y14957 , y14958 , y14959 , y14960 , y14961 , y14962 , y14963 , y14964 , y14965 , y14966 , y14967 , y14968 , y14969 , y14970 , y14971 , y14972 , y14973 , y14974 , y14975 , y14976 , y14977 , y14978 , y14979 , y14980 , y14981 , y14982 , y14983 , y14984 , y14985 , y14986 , y14987 , y14988 , y14989 , y14990 , y14991 , y14992 , y14993 , y14994 , y14995 , y14996 , y14997 , y14998 , y14999 , y15000 , y15001 , y15002 , y15003 , y15004 , y15005 , y15006 , y15007 , y15008 , y15009 , y15010 , y15011 , y15012 , y15013 , y15014 , y15015 , y15016 , y15017 , y15018 , y15019 , y15020 , y15021 , y15022 , y15023 , y15024 , y15025 , y15026 , y15027 , y15028 , y15029 , y15030 , y15031 , y15032 , y15033 , y15034 , y15035 , y15036 , y15037 , y15038 , y15039 , y15040 , y15041 , y15042 , y15043 , y15044 , y15045 , y15046 , y15047 , y15048 , y15049 , y15050 , y15051 , y15052 , y15053 , y15054 , y15055 , y15056 , y15057 , y15058 , y15059 , y15060 , y15061 , y15062 , y15063 , y15064 , y15065 , y15066 , y15067 , y15068 , y15069 , y15070 , y15071 , y15072 , y15073 , y15074 , y15075 , y15076 , y15077 , y15078 , y15079 , y15080 , y15081 , y15082 , y15083 , y15084 , y15085 , y15086 , y15087 , y15088 , y15089 , y15090 , y15091 , y15092 , y15093 , y15094 , y15095 , y15096 , y15097 , y15098 , y15099 , y15100 , y15101 , y15102 , y15103 , y15104 , y15105 , y15106 , y15107 , y15108 , y15109 , y15110 , y15111 , y15112 , y15113 , y15114 , y15115 , y15116 , y15117 , y15118 , y15119 , y15120 , y15121 , y15122 , y15123 , y15124 , y15125 , y15126 , y15127 , y15128 , y15129 , y15130 , y15131 , y15132 , y15133 , y15134 , y15135 , y15136 , y15137 , y15138 , y15139 , y15140 , y15141 , y15142 , y15143 , y15144 , y15145 , y15146 , y15147 , y15148 , y15149 , y15150 , y15151 , y15152 , y15153 , y15154 , y15155 , y15156 , y15157 , y15158 , y15159 , y15160 , y15161 , y15162 , y15163 , y15164 , y15165 , y15166 , y15167 , y15168 , y15169 , y15170 , y15171 , y15172 , y15173 , y15174 , y15175 , y15176 , y15177 , y15178 , y15179 , y15180 , y15181 , y15182 , y15183 , y15184 , y15185 , y15186 , y15187 , y15188 , y15189 , y15190 , y15191 , y15192 , y15193 , y15194 , y15195 , y15196 , y15197 , y15198 , y15199 , y15200 , y15201 , y15202 , y15203 , y15204 , y15205 , y15206 , y15207 , y15208 , y15209 , y15210 , y15211 , y15212 , y15213 , y15214 , y15215 , y15216 , y15217 , y15218 , y15219 , y15220 , y15221 , y15222 , y15223 , y15224 , y15225 , y15226 , y15227 , y15228 , y15229 , y15230 , y15231 , y15232 , y15233 , y15234 , y15235 , y15236 , y15237 , y15238 , y15239 , y15240 , y15241 , y15242 , y15243 , y15244 , y15245 , y15246 , y15247 , y15248 , y15249 , y15250 , y15251 , y15252 , y15253 , y15254 , y15255 , y15256 , y15257 , y15258 , y15259 , y15260 , y15261 , y15262 , y15263 , y15264 , y15265 , y15266 , y15267 , y15268 , y15269 , y15270 , y15271 , y15272 , y15273 , y15274 , y15275 , y15276 , y15277 , y15278 , y15279 , y15280 , y15281 , y15282 , y15283 , y15284 , y15285 , y15286 , y15287 , y15288 , y15289 , y15290 , y15291 , y15292 , y15293 , y15294 , y15295 , y15296 , y15297 , y15298 , y15299 , y15300 , y15301 , y15302 , y15303 , y15304 , y15305 , y15306 , y15307 , y15308 , y15309 , y15310 , y15311 , y15312 , y15313 , y15314 , y15315 , y15316 , y15317 , y15318 , y15319 , y15320 , y15321 , y15322 , y15323 , y15324 , y15325 , y15326 , y15327 , y15328 , y15329 , y15330 , y15331 , y15332 , y15333 , y15334 , y15335 , y15336 , y15337 , y15338 , y15339 , y15340 , y15341 , y15342 , y15343 , y15344 , y15345 , y15346 , y15347 , y15348 , y15349 , y15350 , y15351 , y15352 , y15353 , y15354 , y15355 , y15356 , y15357 , y15358 , y15359 , y15360 , y15361 , y15362 , y15363 , y15364 , y15365 , y15366 , y15367 , y15368 , y15369 , y15370 , y15371 , y15372 , y15373 , y15374 , y15375 , y15376 , y15377 , y15378 , y15379 , y15380 , y15381 , y15382 , y15383 , y15384 , y15385 , y15386 , y15387 , y15388 , y15389 , y15390 , y15391 , y15392 , y15393 , y15394 , y15395 , y15396 , y15397 , y15398 , y15399 , y15400 , y15401 , y15402 , y15403 , y15404 , y15405 , y15406 , y15407 , y15408 , y15409 , y15410 , y15411 , y15412 , y15413 , y15414 , y15415 , y15416 , y15417 , y15418 , y15419 , y15420 , y15421 , y15422 , y15423 , y15424 , y15425 , y15426 , y15427 , y15428 , y15429 , y15430 , y15431 , y15432 , y15433 , y15434 , y15435 , y15436 , y15437 , y15438 , y15439 , y15440 , y15441 , y15442 , y15443 , y15444 , y15445 , y15446 , y15447 , y15448 , y15449 , y15450 , y15451 , y15452 , y15453 , y15454 , y15455 , y15456 , y15457 , y15458 , y15459 , y15460 , y15461 , y15462 , y15463 , y15464 , y15465 , y15466 , y15467 , y15468 , y15469 , y15470 , y15471 , y15472 , y15473 , y15474 , y15475 , y15476 , y15477 , y15478 , y15479 , y15480 , y15481 , y15482 , y15483 , y15484 , y15485 , y15486 , y15487 , y15488 , y15489 , y15490 , y15491 , y15492 , y15493 , y15494 , y15495 , y15496 , y15497 , y15498 , y15499 , y15500 , y15501 , y15502 , y15503 , y15504 , y15505 , y15506 , y15507 , y15508 , y15509 , y15510 , y15511 , y15512 , y15513 , y15514 , y15515 , y15516 , y15517 , y15518 , y15519 , y15520 , y15521 , y15522 , y15523 , y15524 , y15525 , y15526 , y15527 , y15528 , y15529 , y15530 , y15531 , y15532 , y15533 , y15534 , y15535 , y15536 , y15537 , y15538 , y15539 , y15540 , y15541 , y15542 , y15543 , y15544 , y15545 , y15546 , y15547 , y15548 , y15549 , y15550 , y15551 , y15552 , y15553 , y15554 , y15555 , y15556 , y15557 , y15558 , y15559 , y15560 , y15561 , y15562 , y15563 , y15564 , y15565 , y15566 , y15567 , y15568 , y15569 , y15570 , y15571 , y15572 , y15573 , y15574 , y15575 , y15576 , y15577 , y15578 , y15579 , y15580 , y15581 , y15582 , y15583 , y15584 , y15585 , y15586 , y15587 , y15588 , y15589 , y15590 , y15591 , y15592 , y15593 , y15594 , y15595 , y15596 , y15597 , y15598 , y15599 , y15600 , y15601 , y15602 , y15603 , y15604 , y15605 , y15606 , y15607 , y15608 , y15609 , y15610 , y15611 , y15612 , y15613 , y15614 , y15615 , y15616 , y15617 , y15618 , y15619 , y15620 , y15621 , y15622 , y15623 , y15624 , y15625 , y15626 , y15627 , y15628 , y15629 , y15630 , y15631 , y15632 , y15633 , y15634 , y15635 , y15636 , y15637 , y15638 , y15639 , y15640 , y15641 , y15642 , y15643 , y15644 , y15645 , y15646 , y15647 , y15648 , y15649 , y15650 , y15651 , y15652 , y15653 , y15654 , y15655 , y15656 , y15657 , y15658 , y15659 , y15660 , y15661 , y15662 , y15663 , y15664 , y15665 , y15666 , y15667 , y15668 , y15669 , y15670 , y15671 , y15672 , y15673 , y15674 , y15675 , y15676 , y15677 , y15678 , y15679 , y15680 , y15681 , y15682 , y15683 , y15684 , y15685 , y15686 , y15687 , y15688 , y15689 , y15690 , y15691 , y15692 , y15693 , y15694 , y15695 , y15696 , y15697 , y15698 , y15699 , y15700 , y15701 , y15702 , y15703 , y15704 , y15705 , y15706 , y15707 , y15708 , y15709 , y15710 , y15711 , y15712 , y15713 , y15714 , y15715 , y15716 , y15717 , y15718 , y15719 , y15720 , y15721 , y15722 , y15723 , y15724 , y15725 , y15726 , y15727 , y15728 , y15729 , y15730 , y15731 , y15732 , y15733 , y15734 , y15735 , y15736 , y15737 , y15738 , y15739 , y15740 , y15741 , y15742 , y15743 , y15744 , y15745 , y15746 , y15747 , y15748 , y15749 , y15750 , y15751 , y15752 , y15753 , y15754 , y15755 , y15756 , y15757 , y15758 , y15759 , y15760 , y15761 , y15762 , y15763 , y15764 , y15765 , y15766 , y15767 , y15768 , y15769 , y15770 , y15771 , y15772 , y15773 , y15774 , y15775 , y15776 , y15777 , y15778 , y15779 , y15780 , y15781 , y15782 , y15783 , y15784 , y15785 , y15786 , y15787 , y15788 , y15789 , y15790 , y15791 , y15792 , y15793 , y15794 , y15795 , y15796 , y15797 , y15798 , y15799 , y15800 , y15801 , y15802 , y15803 , y15804 , y15805 , y15806 , y15807 , y15808 , y15809 , y15810 , y15811 , y15812 , y15813 , y15814 , y15815 , y15816 , y15817 , y15818 , y15819 , y15820 , y15821 , y15822 , y15823 , y15824 , y15825 , y15826 , y15827 , y15828 , y15829 , y15830 , y15831 , y15832 , y15833 , y15834 , y15835 , y15836 , y15837 , y15838 , y15839 , y15840 , y15841 , y15842 , y15843 , y15844 , y15845 , y15846 , y15847 , y15848 , y15849 , y15850 , y15851 , y15852 , y15853 , y15854 , y15855 , y15856 , y15857 , y15858 , y15859 , y15860 , y15861 , y15862 , y15863 , y15864 , y15865 , y15866 , y15867 , y15868 , y15869 , y15870 , y15871 , y15872 , y15873 , y15874 , y15875 , y15876 , y15877 , y15878 , y15879 , y15880 , y15881 , y15882 , y15883 , y15884 , y15885 , y15886 , y15887 , y15888 , y15889 , y15890 , y15891 , y15892 , y15893 , y15894 , y15895 , y15896 , y15897 , y15898 , y15899 , y15900 , y15901 , y15902 , y15903 , y15904 , y15905 , y15906 , y15907 , y15908 , y15909 , y15910 , y15911 , y15912 , y15913 , y15914 , y15915 , y15916 , y15917 , y15918 , y15919 , y15920 , y15921 , y15922 , y15923 , y15924 , y15925 , y15926 , y15927 , y15928 , y15929 , y15930 , y15931 , y15932 , y15933 , y15934 , y15935 , y15936 , y15937 , y15938 , y15939 , y15940 , y15941 , y15942 , y15943 , y15944 , y15945 , y15946 , y15947 , y15948 , y15949 , y15950 , y15951 , y15952 , y15953 , y15954 , y15955 , y15956 , y15957 , y15958 , y15959 , y15960 , y15961 , y15962 , y15963 , y15964 , y15965 , y15966 , y15967 , y15968 , y15969 , y15970 , y15971 , y15972 , y15973 , y15974 , y15975 , y15976 , y15977 , y15978 , y15979 , y15980 , y15981 , y15982 , y15983 , y15984 , y15985 , y15986 , y15987 , y15988 , y15989 , y15990 , y15991 , y15992 , y15993 , y15994 , y15995 , y15996 , y15997 , y15998 , y15999 , y16000 , y16001 , y16002 , y16003 , y16004 , y16005 , y16006 , y16007 , y16008 , y16009 , y16010 , y16011 , y16012 , y16013 , y16014 , y16015 , y16016 , y16017 , y16018 , y16019 , y16020 , y16021 , y16022 , y16023 , y16024 , y16025 , y16026 , y16027 , y16028 , y16029 , y16030 , y16031 , y16032 , y16033 , y16034 , y16035 , y16036 , y16037 , y16038 , y16039 , y16040 , y16041 , y16042 , y16043 , y16044 , y16045 , y16046 , y16047 , y16048 , y16049 , y16050 , y16051 , y16052 , y16053 , y16054 , y16055 , y16056 , y16057 , y16058 , y16059 , y16060 , y16061 , y16062 , y16063 , y16064 , y16065 , y16066 , y16067 , y16068 , y16069 , y16070 , y16071 , y16072 , y16073 , y16074 , y16075 , y16076 , y16077 , y16078 , y16079 , y16080 , y16081 , y16082 , y16083 , y16084 , y16085 , y16086 , y16087 , y16088 , y16089 , y16090 , y16091 , y16092 , y16093 , y16094 , y16095 , y16096 , y16097 , y16098 , y16099 , y16100 , y16101 , y16102 , y16103 , y16104 , y16105 , y16106 , y16107 , y16108 , y16109 , y16110 , y16111 , y16112 , y16113 , y16114 , y16115 , y16116 , y16117 , y16118 , y16119 , y16120 , y16121 , y16122 , y16123 , y16124 , y16125 , y16126 , y16127 , y16128 , y16129 , y16130 , y16131 , y16132 , y16133 , y16134 , y16135 , y16136 , y16137 , y16138 , y16139 , y16140 , y16141 , y16142 , y16143 , y16144 , y16145 , y16146 , y16147 , y16148 , y16149 , y16150 , y16151 , y16152 , y16153 , y16154 , y16155 , y16156 , y16157 , y16158 , y16159 , y16160 , y16161 , y16162 , y16163 , y16164 , y16165 , y16166 , y16167 , y16168 , y16169 , y16170 , y16171 , y16172 , y16173 , y16174 , y16175 , y16176 , y16177 , y16178 , y16179 , y16180 , y16181 , y16182 , y16183 , y16184 , y16185 , y16186 , y16187 , y16188 , y16189 , y16190 , y16191 , y16192 , y16193 , y16194 , y16195 , y16196 , y16197 , y16198 , y16199 , y16200 , y16201 , y16202 , y16203 , y16204 , y16205 , y16206 , y16207 , y16208 , y16209 , y16210 , y16211 , y16212 , y16213 , y16214 , y16215 , y16216 , y16217 , y16218 , y16219 , y16220 , y16221 , y16222 , y16223 , y16224 , y16225 , y16226 , y16227 , y16228 , y16229 , y16230 , y16231 , y16232 , y16233 , y16234 , y16235 , y16236 , y16237 , y16238 , y16239 , y16240 , y16241 , y16242 , y16243 , y16244 , y16245 , y16246 , y16247 , y16248 , y16249 , y16250 , y16251 , y16252 , y16253 , y16254 , y16255 , y16256 , y16257 , y16258 , y16259 , y16260 , y16261 , y16262 , y16263 , y16264 , y16265 , y16266 , y16267 , y16268 , y16269 , y16270 , y16271 , y16272 , y16273 , y16274 , y16275 , y16276 , y16277 , y16278 , y16279 , y16280 , y16281 , y16282 , y16283 , y16284 , y16285 , y16286 , y16287 , y16288 , y16289 , y16290 , y16291 , y16292 , y16293 , y16294 , y16295 , y16296 , y16297 , y16298 , y16299 , y16300 , y16301 , y16302 , y16303 , y16304 , y16305 , y16306 , y16307 , y16308 , y16309 , y16310 , y16311 , y16312 , y16313 , y16314 , y16315 , y16316 , y16317 , y16318 , y16319 , y16320 , y16321 , y16322 , y16323 , y16324 , y16325 , y16326 , y16327 , y16328 , y16329 , y16330 , y16331 , y16332 , y16333 , y16334 , y16335 , y16336 , y16337 , y16338 , y16339 , y16340 , y16341 , y16342 , y16343 , y16344 , y16345 , y16346 , y16347 , y16348 , y16349 , y16350 , y16351 , y16352 , y16353 , y16354 , y16355 , y16356 , y16357 , y16358 , y16359 , y16360 , y16361 , y16362 , y16363 , y16364 , y16365 , y16366 , y16367 , y16368 , y16369 , y16370 , y16371 , y16372 , y16373 , y16374 , y16375 , y16376 , y16377 , y16378 , y16379 , y16380 , y16381 , y16382 , y16383 , y16384 , y16385 , y16386 , y16387 , y16388 , y16389 , y16390 , y16391 , y16392 , y16393 , y16394 , y16395 , y16396 , y16397 , y16398 , y16399 , y16400 , y16401 , y16402 , y16403 , y16404 , y16405 , y16406 , y16407 , y16408 , y16409 , y16410 , y16411 , y16412 , y16413 , y16414 , y16415 , y16416 , y16417 , y16418 , y16419 , y16420 , y16421 , y16422 , y16423 , y16424 , y16425 , y16426 , y16427 , y16428 , y16429 , y16430 , y16431 , y16432 , y16433 , y16434 , y16435 , y16436 , y16437 , y16438 , y16439 , y16440 , y16441 , y16442 , y16443 , y16444 , y16445 , y16446 , y16447 , y16448 , y16449 , y16450 , y16451 , y16452 , y16453 , y16454 , y16455 , y16456 , y16457 , y16458 , y16459 , y16460 , y16461 , y16462 , y16463 , y16464 , y16465 , y16466 , y16467 , y16468 , y16469 , y16470 , y16471 , y16472 , y16473 , y16474 , y16475 , y16476 , y16477 , y16478 , y16479 , y16480 , y16481 , y16482 , y16483 , y16484 , y16485 , y16486 , y16487 , y16488 , y16489 , y16490 , y16491 , y16492 , y16493 , y16494 , y16495 , y16496 , y16497 , y16498 , y16499 , y16500 , y16501 , y16502 , y16503 , y16504 , y16505 , y16506 , y16507 , y16508 , y16509 , y16510 , y16511 , y16512 , y16513 , y16514 , y16515 , y16516 , y16517 , y16518 , y16519 , y16520 , y16521 , y16522 , y16523 , y16524 , y16525 , y16526 , y16527 , y16528 , y16529 , y16530 , y16531 , y16532 , y16533 , y16534 , y16535 , y16536 , y16537 , y16538 , y16539 , y16540 , y16541 , y16542 , y16543 , y16544 , y16545 , y16546 , y16547 , y16548 , y16549 , y16550 , y16551 , y16552 , y16553 , y16554 , y16555 , y16556 , y16557 , y16558 , y16559 , y16560 , y16561 , y16562 , y16563 , y16564 , y16565 , y16566 , y16567 , y16568 , y16569 , y16570 , y16571 , y16572 , y16573 , y16574 , y16575 , y16576 , y16577 , y16578 , y16579 , y16580 , y16581 , y16582 , y16583 , y16584 , y16585 , y16586 , y16587 , y16588 , y16589 , y16590 , y16591 , y16592 , y16593 , y16594 , y16595 , y16596 , y16597 , y16598 , y16599 , y16600 , y16601 , y16602 , y16603 , y16604 , y16605 , y16606 , y16607 , y16608 , y16609 , y16610 , y16611 , y16612 , y16613 , y16614 , y16615 , y16616 , y16617 , y16618 , y16619 , y16620 , y16621 , y16622 , y16623 , y16624 , y16625 , y16626 , y16627 , y16628 , y16629 , y16630 , y16631 , y16632 , y16633 , y16634 , y16635 , y16636 , y16637 , y16638 , y16639 , y16640 , y16641 , y16642 , y16643 , y16644 , y16645 , y16646 , y16647 , y16648 , y16649 , y16650 , y16651 , y16652 , y16653 , y16654 , y16655 , y16656 , y16657 , y16658 , y16659 , y16660 , y16661 , y16662 , y16663 , y16664 , y16665 , y16666 , y16667 , y16668 , y16669 , y16670 , y16671 , y16672 , y16673 , y16674 , y16675 , y16676 , y16677 , y16678 , y16679 , y16680 , y16681 , y16682 , y16683 , y16684 , y16685 , y16686 , y16687 , y16688 , y16689 , y16690 , y16691 , y16692 , y16693 , y16694 , y16695 , y16696 , y16697 , y16698 , y16699 , y16700 , y16701 , y16702 , y16703 , y16704 , y16705 , y16706 , y16707 , y16708 , y16709 , y16710 , y16711 , y16712 , y16713 , y16714 , y16715 , y16716 , y16717 , y16718 , y16719 , y16720 , y16721 , y16722 , y16723 , y16724 , y16725 , y16726 , y16727 , y16728 , y16729 , y16730 , y16731 , y16732 , y16733 , y16734 , y16735 , y16736 , y16737 , y16738 , y16739 , y16740 , y16741 , y16742 , y16743 , y16744 , y16745 , y16746 , y16747 , y16748 , y16749 , y16750 , y16751 , y16752 , y16753 , y16754 , y16755 , y16756 , y16757 , y16758 , y16759 , y16760 , y16761 , y16762 , y16763 , y16764 , y16765 , y16766 , y16767 , y16768 , y16769 , y16770 , y16771 , y16772 , y16773 , y16774 , y16775 , y16776 , y16777 , y16778 , y16779 , y16780 , y16781 , y16782 , y16783 , y16784 , y16785 , y16786 , y16787 , y16788 , y16789 , y16790 , y16791 , y16792 , y16793 , y16794 , y16795 , y16796 , y16797 , y16798 , y16799 , y16800 , y16801 , y16802 , y16803 , y16804 , y16805 , y16806 , y16807 , y16808 , y16809 , y16810 , y16811 , y16812 , y16813 , y16814 , y16815 , y16816 , y16817 , y16818 , y16819 , y16820 , y16821 , y16822 , y16823 , y16824 , y16825 , y16826 , y16827 , y16828 , y16829 , y16830 , y16831 , y16832 , y16833 , y16834 , y16835 , y16836 , y16837 , y16838 , y16839 , y16840 , y16841 , y16842 , y16843 , y16844 , y16845 , y16846 , y16847 , y16848 , y16849 , y16850 , y16851 , y16852 , y16853 , y16854 , y16855 , y16856 , y16857 , y16858 , y16859 , y16860 , y16861 , y16862 , y16863 , y16864 , y16865 , y16866 , y16867 , y16868 , y16869 , y16870 , y16871 , y16872 , y16873 , y16874 , y16875 , y16876 , y16877 , y16878 , y16879 , y16880 , y16881 , y16882 , y16883 , y16884 , y16885 , y16886 , y16887 , y16888 , y16889 , y16890 , y16891 , y16892 , y16893 , y16894 , y16895 , y16896 , y16897 , y16898 , y16899 , y16900 , y16901 , y16902 , y16903 , y16904 , y16905 , y16906 , y16907 , y16908 , y16909 , y16910 , y16911 , y16912 , y16913 , y16914 , y16915 , y16916 , y16917 , y16918 , y16919 , y16920 , y16921 , y16922 , y16923 , y16924 , y16925 , y16926 , y16927 , y16928 , y16929 , y16930 , y16931 , y16932 , y16933 , y16934 , y16935 , y16936 , y16937 , y16938 , y16939 , y16940 , y16941 , y16942 , y16943 , y16944 , y16945 , y16946 , y16947 , y16948 , y16949 , y16950 , y16951 , y16952 , y16953 , y16954 , y16955 , y16956 , y16957 , y16958 , y16959 , y16960 , y16961 , y16962 , y16963 , y16964 , y16965 , y16966 , y16967 , y16968 , y16969 , y16970 , y16971 , y16972 , y16973 , y16974 , y16975 , y16976 , y16977 , y16978 , y16979 , y16980 , y16981 , y16982 , y16983 , y16984 , y16985 , y16986 , y16987 , y16988 , y16989 , y16990 , y16991 , y16992 , y16993 , y16994 , y16995 , y16996 , y16997 , y16998 , y16999 , y17000 , y17001 , y17002 , y17003 , y17004 , y17005 , y17006 , y17007 , y17008 , y17009 , y17010 , y17011 , y17012 , y17013 , y17014 , y17015 , y17016 , y17017 , y17018 , y17019 , y17020 , y17021 , y17022 , y17023 , y17024 , y17025 , y17026 , y17027 , y17028 , y17029 , y17030 , y17031 , y17032 , y17033 , y17034 , y17035 , y17036 , y17037 , y17038 , y17039 , y17040 , y17041 , y17042 , y17043 , y17044 , y17045 , y17046 , y17047 , y17048 , y17049 , y17050 , y17051 , y17052 , y17053 , y17054 , y17055 , y17056 , y17057 , y17058 , y17059 , y17060 , y17061 , y17062 , y17063 , y17064 , y17065 , y17066 , y17067 , y17068 , y17069 , y17070 , y17071 , y17072 , y17073 , y17074 , y17075 , y17076 , y17077 , y17078 , y17079 , y17080 , y17081 , y17082 , y17083 , y17084 , y17085 , y17086 , y17087 , y17088 , y17089 , y17090 , y17091 , y17092 , y17093 , y17094 , y17095 , y17096 , y17097 , y17098 , y17099 , y17100 , y17101 , y17102 , y17103 , y17104 , y17105 , y17106 , y17107 , y17108 , y17109 , y17110 , y17111 , y17112 , y17113 , y17114 , y17115 , y17116 , y17117 , y17118 , y17119 , y17120 , y17121 , y17122 , y17123 , y17124 , y17125 , y17126 , y17127 , y17128 , y17129 , y17130 , y17131 , y17132 , y17133 , y17134 , y17135 , y17136 , y17137 , y17138 , y17139 , y17140 , y17141 , y17142 , y17143 , y17144 , y17145 , y17146 , y17147 , y17148 , y17149 , y17150 , y17151 , y17152 , y17153 , y17154 , y17155 , y17156 , y17157 , y17158 , y17159 , y17160 , y17161 , y17162 , y17163 , y17164 , y17165 , y17166 , y17167 , y17168 , y17169 , y17170 , y17171 , y17172 , y17173 , y17174 , y17175 , y17176 , y17177 , y17178 , y17179 , y17180 , y17181 , y17182 , y17183 , y17184 , y17185 , y17186 , y17187 , y17188 , y17189 , y17190 , y17191 , y17192 , y17193 , y17194 , y17195 , y17196 , y17197 , y17198 , y17199 , y17200 , y17201 , y17202 , y17203 , y17204 , y17205 , y17206 , y17207 , y17208 , y17209 , y17210 , y17211 , y17212 , y17213 , y17214 , y17215 , y17216 , y17217 , y17218 , y17219 , y17220 , y17221 , y17222 , y17223 , y17224 , y17225 , y17226 , y17227 , y17228 , y17229 , y17230 , y17231 , y17232 , y17233 , y17234 , y17235 , y17236 , y17237 , y17238 , y17239 , y17240 , y17241 , y17242 , y17243 , y17244 , y17245 , y17246 , y17247 , y17248 , y17249 , y17250 , y17251 , y17252 , y17253 , y17254 , y17255 , y17256 , y17257 , y17258 , y17259 , y17260 , y17261 , y17262 , y17263 , y17264 , y17265 , y17266 , y17267 , y17268 , y17269 , y17270 , y17271 , y17272 , y17273 , y17274 , y17275 , y17276 , y17277 , y17278 , y17279 , y17280 , y17281 , y17282 , y17283 , y17284 , y17285 , y17286 , y17287 , y17288 , y17289 , y17290 , y17291 , y17292 , y17293 , y17294 , y17295 , y17296 , y17297 , y17298 , y17299 , y17300 , y17301 , y17302 , y17303 , y17304 , y17305 , y17306 , y17307 , y17308 , y17309 , y17310 , y17311 , y17312 , y17313 , y17314 , y17315 , y17316 , y17317 , y17318 , y17319 , y17320 , y17321 , y17322 , y17323 , y17324 , y17325 , y17326 , y17327 , y17328 , y17329 , y17330 , y17331 , y17332 , y17333 , y17334 , y17335 , y17336 , y17337 , y17338 , y17339 , y17340 , y17341 , y17342 , y17343 , y17344 , y17345 , y17346 , y17347 , y17348 , y17349 , y17350 , y17351 , y17352 , y17353 , y17354 , y17355 , y17356 , y17357 , y17358 , y17359 , y17360 , y17361 , y17362 , y17363 , y17364 , y17365 , y17366 , y17367 , y17368 , y17369 , y17370 , y17371 , y17372 , y17373 , y17374 , y17375 , y17376 , y17377 , y17378 , y17379 , y17380 , y17381 , y17382 , y17383 , y17384 , y17385 , y17386 , y17387 , y17388 , y17389 , y17390 , y17391 , y17392 , y17393 , y17394 , y17395 , y17396 , y17397 , y17398 , y17399 , y17400 , y17401 , y17402 , y17403 , y17404 , y17405 , y17406 , y17407 , y17408 , y17409 , y17410 , y17411 , y17412 , y17413 , y17414 , y17415 , y17416 , y17417 , y17418 , y17419 , y17420 , y17421 , y17422 , y17423 , y17424 , y17425 , y17426 , y17427 , y17428 , y17429 , y17430 , y17431 , y17432 , y17433 , y17434 , y17435 , y17436 , y17437 , y17438 , y17439 , y17440 , y17441 , y17442 , y17443 , y17444 , y17445 , y17446 , y17447 , y17448 , y17449 , y17450 , y17451 , y17452 , y17453 , y17454 , y17455 , y17456 , y17457 , y17458 , y17459 , y17460 , y17461 , y17462 , y17463 , y17464 , y17465 , y17466 , y17467 , y17468 , y17469 , y17470 , y17471 , y17472 , y17473 , y17474 , y17475 , y17476 , y17477 , y17478 , y17479 , y17480 , y17481 , y17482 , y17483 , y17484 , y17485 , y17486 , y17487 , y17488 , y17489 , y17490 , y17491 , y17492 , y17493 , y17494 , y17495 , y17496 , y17497 , y17498 , y17499 , y17500 , y17501 , y17502 , y17503 , y17504 , y17505 , y17506 , y17507 , y17508 , y17509 , y17510 , y17511 , y17512 , y17513 , y17514 , y17515 , y17516 , y17517 , y17518 , y17519 , y17520 , y17521 , y17522 , y17523 , y17524 , y17525 , y17526 , y17527 , y17528 , y17529 , y17530 , y17531 , y17532 , y17533 , y17534 , y17535 , y17536 , y17537 , y17538 , y17539 , y17540 , y17541 , y17542 , y17543 , y17544 , y17545 , y17546 , y17547 , y17548 , y17549 , y17550 , y17551 , y17552 , y17553 , y17554 , y17555 , y17556 , y17557 , y17558 , y17559 , y17560 , y17561 , y17562 , y17563 , y17564 , y17565 , y17566 , y17567 , y17568 , y17569 , y17570 , y17571 , y17572 , y17573 , y17574 , y17575 , y17576 , y17577 , y17578 , y17579 , y17580 , y17581 , y17582 , y17583 , y17584 , y17585 , y17586 , y17587 , y17588 , y17589 , y17590 , y17591 , y17592 , y17593 , y17594 , y17595 , y17596 , y17597 , y17598 , y17599 , y17600 , y17601 , y17602 , y17603 , y17604 , y17605 , y17606 , y17607 , y17608 , y17609 , y17610 , y17611 , y17612 , y17613 , y17614 , y17615 , y17616 , y17617 , y17618 , y17619 , y17620 , y17621 , y17622 , y17623 , y17624 , y17625 , y17626 , y17627 , y17628 , y17629 , y17630 , y17631 , y17632 , y17633 , y17634 , y17635 , y17636 , y17637 , y17638 , y17639 , y17640 , y17641 , y17642 , y17643 , y17644 , y17645 , y17646 , y17647 , y17648 , y17649 , y17650 , y17651 , y17652 , y17653 , y17654 , y17655 , y17656 , y17657 , y17658 , y17659 , y17660 , y17661 , y17662 , y17663 , y17664 , y17665 , y17666 , y17667 , y17668 , y17669 , y17670 , y17671 , y17672 , y17673 , y17674 , y17675 , y17676 , y17677 , y17678 , y17679 , y17680 , y17681 , y17682 , y17683 , y17684 , y17685 , y17686 , y17687 , y17688 , y17689 , y17690 , y17691 , y17692 , y17693 , y17694 , y17695 , y17696 , y17697 , y17698 , y17699 , y17700 , y17701 , y17702 , y17703 , y17704 , y17705 , y17706 , y17707 , y17708 , y17709 , y17710 , y17711 , y17712 , y17713 , y17714 , y17715 , y17716 , y17717 , y17718 , y17719 , y17720 , y17721 , y17722 , y17723 , y17724 , y17725 , y17726 , y17727 , y17728 , y17729 , y17730 , y17731 , y17732 , y17733 , y17734 , y17735 , y17736 , y17737 , y17738 , y17739 , y17740 , y17741 , y17742 , y17743 , y17744 , y17745 , y17746 , y17747 , y17748 , y17749 , y17750 , y17751 , y17752 , y17753 , y17754 , y17755 , y17756 , y17757 , y17758 , y17759 , y17760 , y17761 , y17762 , y17763 , y17764 , y17765 , y17766 , y17767 , y17768 , y17769 , y17770 , y17771 , y17772 , y17773 , y17774 , y17775 , y17776 , y17777 , y17778 , y17779 , y17780 , y17781 , y17782 , y17783 , y17784 , y17785 , y17786 , y17787 , y17788 , y17789 , y17790 , y17791 , y17792 , y17793 , y17794 , y17795 , y17796 , y17797 , y17798 , y17799 , y17800 , y17801 , y17802 , y17803 , y17804 , y17805 , y17806 , y17807 , y17808 , y17809 , y17810 , y17811 , y17812 , y17813 , y17814 , y17815 , y17816 , y17817 , y17818 , y17819 , y17820 , y17821 , y17822 , y17823 , y17824 , y17825 , y17826 , y17827 , y17828 , y17829 , y17830 , y17831 , y17832 , y17833 , y17834 , y17835 , y17836 , y17837 , y17838 , y17839 , y17840 , y17841 , y17842 , y17843 , y17844 , y17845 , y17846 , y17847 , y17848 , y17849 , y17850 , y17851 , y17852 , y17853 , y17854 , y17855 , y17856 , y17857 , y17858 , y17859 , y17860 , y17861 , y17862 , y17863 , y17864 , y17865 , y17866 , y17867 , y17868 , y17869 , y17870 , y17871 , y17872 , y17873 , y17874 , y17875 , y17876 , y17877 , y17878 , y17879 , y17880 , y17881 , y17882 , y17883 , y17884 , y17885 , y17886 , y17887 , y17888 , y17889 , y17890 , y17891 , y17892 , y17893 , y17894 , y17895 , y17896 , y17897 , y17898 , y17899 , y17900 , y17901 , y17902 , y17903 , y17904 , y17905 , y17906 , y17907 , y17908 , y17909 , y17910 , y17911 , y17912 , y17913 , y17914 , y17915 , y17916 , y17917 , y17918 , y17919 , y17920 , y17921 , y17922 , y17923 , y17924 , y17925 , y17926 , y17927 , y17928 , y17929 , y17930 , y17931 , y17932 , y17933 , y17934 , y17935 , y17936 , y17937 , y17938 , y17939 , y17940 , y17941 , y17942 , y17943 , y17944 , y17945 , y17946 , y17947 , y17948 , y17949 , y17950 , y17951 , y17952 , y17953 , y17954 , y17955 , y17956 , y17957 , y17958 , y17959 , y17960 , y17961 , y17962 , y17963 , y17964 , y17965 , y17966 , y17967 , y17968 , y17969 , y17970 , y17971 , y17972 , y17973 , y17974 , y17975 , y17976 , y17977 , y17978 , y17979 , y17980 , y17981 , y17982 , y17983 , y17984 , y17985 , y17986 , y17987 , y17988 , y17989 , y17990 , y17991 , y17992 , y17993 , y17994 , y17995 , y17996 , y17997 , y17998 , y17999 , y18000 , y18001 , y18002 , y18003 , y18004 , y18005 , y18006 , y18007 , y18008 , y18009 , y18010 , y18011 , y18012 , y18013 , y18014 , y18015 , y18016 , y18017 , y18018 , y18019 , y18020 , y18021 , y18022 , y18023 , y18024 , y18025 , y18026 , y18027 , y18028 , y18029 , y18030 , y18031 , y18032 , y18033 , y18034 , y18035 , y18036 , y18037 , y18038 , y18039 , y18040 , y18041 , y18042 , y18043 , y18044 , y18045 , y18046 , y18047 , y18048 , y18049 , y18050 , y18051 , y18052 , y18053 , y18054 , y18055 , y18056 , y18057 , y18058 , y18059 , y18060 , y18061 , y18062 , y18063 , y18064 , y18065 , y18066 , y18067 , y18068 , y18069 , y18070 , y18071 , y18072 , y18073 , y18074 , y18075 , y18076 , y18077 , y18078 , y18079 , y18080 , y18081 , y18082 , y18083 , y18084 , y18085 , y18086 , y18087 , y18088 , y18089 , y18090 , y18091 , y18092 , y18093 , y18094 , y18095 , y18096 , y18097 , y18098 , y18099 , y18100 , y18101 , y18102 , y18103 , y18104 , y18105 , y18106 , y18107 , y18108 , y18109 , y18110 , y18111 , y18112 , y18113 , y18114 , y18115 , y18116 , y18117 , y18118 , y18119 , y18120 , y18121 , y18122 , y18123 , y18124 , y18125 , y18126 , y18127 , y18128 , y18129 , y18130 , y18131 , y18132 , y18133 , y18134 , y18135 , y18136 , y18137 , y18138 , y18139 , y18140 , y18141 , y18142 , y18143 , y18144 , y18145 , y18146 , y18147 , y18148 , y18149 , y18150 , y18151 , y18152 , y18153 , y18154 , y18155 , y18156 , y18157 , y18158 , y18159 , y18160 , y18161 , y18162 , y18163 , y18164 , y18165 , y18166 , y18167 , y18168 , y18169 , y18170 , y18171 , y18172 , y18173 , y18174 , y18175 , y18176 , y18177 , y18178 , y18179 , y18180 , y18181 , y18182 , y18183 , y18184 , y18185 , y18186 , y18187 , y18188 , y18189 , y18190 , y18191 , y18192 , y18193 , y18194 , y18195 , y18196 , y18197 , y18198 , y18199 , y18200 , y18201 , y18202 , y18203 , y18204 , y18205 , y18206 , y18207 , y18208 , y18209 , y18210 , y18211 , y18212 , y18213 , y18214 , y18215 , y18216 , y18217 , y18218 , y18219 , y18220 , y18221 , y18222 , y18223 , y18224 , y18225 , y18226 , y18227 , y18228 , y18229 , y18230 , y18231 , y18232 , y18233 , y18234 , y18235 , y18236 , y18237 , y18238 , y18239 , y18240 , y18241 , y18242 , y18243 , y18244 , y18245 , y18246 , y18247 , y18248 , y18249 , y18250 , y18251 , y18252 , y18253 , y18254 , y18255 , y18256 , y18257 , y18258 , y18259 , y18260 , y18261 , y18262 , y18263 , y18264 , y18265 , y18266 , y18267 , y18268 , y18269 , y18270 , y18271 , y18272 , y18273 , y18274 , y18275 , y18276 , y18277 , y18278 , y18279 , y18280 , y18281 , y18282 , y18283 , y18284 , y18285 , y18286 , y18287 , y18288 , y18289 , y18290 , y18291 , y18292 , y18293 , y18294 , y18295 , y18296 , y18297 , y18298 , y18299 , y18300 , y18301 , y18302 , y18303 , y18304 , y18305 , y18306 , y18307 , y18308 , y18309 , y18310 , y18311 , y18312 , y18313 , y18314 , y18315 , y18316 , y18317 , y18318 , y18319 , y18320 , y18321 , y18322 , y18323 , y18324 , y18325 , y18326 , y18327 , y18328 , y18329 , y18330 , y18331 , y18332 , y18333 , y18334 , y18335 , y18336 , y18337 , y18338 , y18339 , y18340 , y18341 , y18342 , y18343 , y18344 , y18345 , y18346 , y18347 , y18348 , y18349 , y18350 , y18351 , y18352 , y18353 , y18354 , y18355 , y18356 , y18357 , y18358 , y18359 , y18360 , y18361 , y18362 , y18363 , y18364 , y18365 , y18366 , y18367 , y18368 , y18369 , y18370 , y18371 , y18372 , y18373 , y18374 , y18375 , y18376 , y18377 , y18378 , y18379 , y18380 , y18381 , y18382 , y18383 , y18384 , y18385 , y18386 , y18387 , y18388 , y18389 , y18390 , y18391 , y18392 , y18393 , y18394 , y18395 , y18396 , y18397 , y18398 , y18399 , y18400 , y18401 , y18402 , y18403 , y18404 , y18405 , y18406 , y18407 , y18408 , y18409 , y18410 , y18411 , y18412 , y18413 , y18414 , y18415 , y18416 , y18417 , y18418 , y18419 , y18420 , y18421 , y18422 , y18423 , y18424 , y18425 , y18426 , y18427 , y18428 , y18429 , y18430 , y18431 , y18432 , y18433 , y18434 , y18435 , y18436 , y18437 , y18438 , y18439 , y18440 , y18441 , y18442 , y18443 , y18444 , y18445 , y18446 , y18447 , y18448 , y18449 , y18450 , y18451 , y18452 , y18453 , y18454 , y18455 , y18456 , y18457 , y18458 , y18459 , y18460 , y18461 , y18462 , y18463 , y18464 , y18465 , y18466 , y18467 , y18468 , y18469 , y18470 , y18471 , y18472 , y18473 , y18474 , y18475 , y18476 , y18477 , y18478 , y18479 , y18480 , y18481 , y18482 , y18483 , y18484 , y18485 , y18486 , y18487 , y18488 , y18489 , y18490 , y18491 , y18492 , y18493 , y18494 , y18495 , y18496 , y18497 , y18498 , y18499 , y18500 , y18501 , y18502 , y18503 , y18504 , y18505 , y18506 , y18507 , y18508 , y18509 , y18510 , y18511 , y18512 , y18513 , y18514 , y18515 , y18516 , y18517 , y18518 , y18519 , y18520 , y18521 , y18522 , y18523 , y18524 , y18525 , y18526 , y18527 , y18528 , y18529 , y18530 , y18531 , y18532 , y18533 , y18534 , y18535 , y18536 , y18537 , y18538 , y18539 , y18540 , y18541 , y18542 , y18543 , y18544 , y18545 , y18546 , y18547 , y18548 , y18549 , y18550 , y18551 , y18552 , y18553 , y18554 , y18555 , y18556 , y18557 , y18558 , y18559 , y18560 , y18561 , y18562 , y18563 , y18564 , y18565 , y18566 , y18567 , y18568 , y18569 , y18570 , y18571 , y18572 , y18573 , y18574 , y18575 , y18576 , y18577 , y18578 , y18579 , y18580 , y18581 , y18582 , y18583 , y18584 , y18585 , y18586 , y18587 , y18588 , y18589 , y18590 , y18591 , y18592 , y18593 , y18594 , y18595 , y18596 , y18597 , y18598 , y18599 , y18600 , y18601 , y18602 , y18603 , y18604 , y18605 , y18606 , y18607 , y18608 , y18609 , y18610 , y18611 , y18612 , y18613 , y18614 , y18615 , y18616 , y18617 , y18618 , y18619 , y18620 , y18621 , y18622 , y18623 , y18624 , y18625 , y18626 , y18627 , y18628 , y18629 , y18630 , y18631 , y18632 , y18633 , y18634 , y18635 , y18636 , y18637 , y18638 , y18639 , y18640 , y18641 , y18642 , y18643 , y18644 , y18645 , y18646 , y18647 , y18648 , y18649 , y18650 , y18651 , y18652 , y18653 , y18654 , y18655 , y18656 , y18657 , y18658 , y18659 , y18660 , y18661 , y18662 , y18663 , y18664 , y18665 , y18666 , y18667 , y18668 , y18669 , y18670 , y18671 , y18672 , y18673 , y18674 , y18675 , y18676 , y18677 , y18678 , y18679 , y18680 , y18681 , y18682 , y18683 , y18684 , y18685 , y18686 , y18687 , y18688 , y18689 , y18690 , y18691 , y18692 , y18693 , y18694 , y18695 , y18696 , y18697 , y18698 , y18699 , y18700 , y18701 , y18702 , y18703 , y18704 , y18705 , y18706 , y18707 , y18708 , y18709 , y18710 , y18711 , y18712 , y18713 , y18714 , y18715 , y18716 , y18717 , y18718 , y18719 , y18720 , y18721 , y18722 , y18723 , y18724 , y18725 , y18726 , y18727 , y18728 , y18729 , y18730 , y18731 , y18732 , y18733 , y18734 , y18735 , y18736 , y18737 , y18738 , y18739 , y18740 , y18741 , y18742 , y18743 , y18744 , y18745 , y18746 , y18747 , y18748 , y18749 , y18750 , y18751 , y18752 , y18753 , y18754 , y18755 , y18756 , y18757 , y18758 , y18759 , y18760 , y18761 , y18762 , y18763 , y18764 , y18765 , y18766 , y18767 , y18768 , y18769 , y18770 , y18771 , y18772 , y18773 , y18774 , y18775 , y18776 , y18777 , y18778 , y18779 , y18780 , y18781 , y18782 , y18783 , y18784 , y18785 , y18786 , y18787 , y18788 , y18789 , y18790 , y18791 , y18792 , y18793 , y18794 , y18795 , y18796 , y18797 , y18798 , y18799 , y18800 , y18801 , y18802 , y18803 , y18804 , y18805 , y18806 , y18807 , y18808 , y18809 , y18810 , y18811 , y18812 , y18813 , y18814 , y18815 , y18816 , y18817 , y18818 , y18819 , y18820 , y18821 , y18822 , y18823 , y18824 , y18825 , y18826 , y18827 , y18828 , y18829 , y18830 , y18831 , y18832 , y18833 , y18834 , y18835 , y18836 , y18837 , y18838 , y18839 , y18840 , y18841 , y18842 , y18843 , y18844 , y18845 , y18846 , y18847 , y18848 , y18849 , y18850 , y18851 , y18852 , y18853 , y18854 , y18855 , y18856 , y18857 , y18858 , y18859 , y18860 , y18861 , y18862 , y18863 , y18864 , y18865 , y18866 , y18867 , y18868 , y18869 , y18870 , y18871 , y18872 , y18873 , y18874 , y18875 , y18876 , y18877 , y18878 , y18879 , y18880 , y18881 , y18882 , y18883 , y18884 , y18885 , y18886 , y18887 , y18888 , y18889 , y18890 , y18891 , y18892 , y18893 , y18894 , y18895 , y18896 , y18897 , y18898 , y18899 , y18900 , y18901 , y18902 , y18903 , y18904 , y18905 , y18906 , y18907 , y18908 , y18909 , y18910 , y18911 , y18912 , y18913 , y18914 , y18915 , y18916 , y18917 , y18918 , y18919 , y18920 , y18921 , y18922 , y18923 , y18924 , y18925 , y18926 , y18927 , y18928 , y18929 , y18930 , y18931 , y18932 , y18933 , y18934 , y18935 , y18936 , y18937 , y18938 , y18939 , y18940 , y18941 , y18942 , y18943 , y18944 , y18945 , y18946 , y18947 , y18948 , y18949 , y18950 , y18951 , y18952 , y18953 , y18954 , y18955 , y18956 , y18957 , y18958 , y18959 , y18960 , y18961 , y18962 , y18963 , y18964 , y18965 , y18966 , y18967 , y18968 , y18969 , y18970 , y18971 , y18972 , y18973 , y18974 , y18975 , y18976 , y18977 , y18978 , y18979 , y18980 , y18981 , y18982 , y18983 , y18984 , y18985 , y18986 , y18987 , y18988 , y18989 , y18990 , y18991 , y18992 , y18993 , y18994 , y18995 , y18996 , y18997 , y18998 , y18999 , y19000 , y19001 , y19002 , y19003 , y19004 , y19005 , y19006 , y19007 , y19008 , y19009 , y19010 , y19011 , y19012 , y19013 , y19014 , y19015 , y19016 , y19017 , y19018 , y19019 , y19020 , y19021 , y19022 , y19023 , y19024 , y19025 , y19026 , y19027 , y19028 , y19029 , y19030 , y19031 , y19032 , y19033 , y19034 , y19035 , y19036 , y19037 , y19038 , y19039 , y19040 , y19041 , y19042 , y19043 , y19044 , y19045 , y19046 , y19047 , y19048 , y19049 , y19050 , y19051 , y19052 , y19053 , y19054 , y19055 , y19056 , y19057 , y19058 , y19059 , y19060 , y19061 , y19062 , y19063 , y19064 , y19065 , y19066 , y19067 , y19068 , y19069 , y19070 , y19071 , y19072 , y19073 , y19074 , y19075 , y19076 , y19077 , y19078 , y19079 , y19080 , y19081 , y19082 , y19083 , y19084 , y19085 , y19086 , y19087 , y19088 , y19089 , y19090 , y19091 , y19092 , y19093 , y19094 , y19095 , y19096 , y19097 , y19098 , y19099 , y19100 , y19101 , y19102 , y19103 , y19104 , y19105 , y19106 , y19107 , y19108 , y19109 , y19110 , y19111 , y19112 , y19113 , y19114 , y19115 , y19116 , y19117 , y19118 , y19119 , y19120 , y19121 , y19122 , y19123 , y19124 , y19125 , y19126 , y19127 , y19128 , y19129 , y19130 , y19131 , y19132 , y19133 , y19134 , y19135 , y19136 , y19137 , y19138 , y19139 , y19140 , y19141 , y19142 , y19143 , y19144 , y19145 , y19146 , y19147 , y19148 , y19149 , y19150 , y19151 , y19152 , y19153 , y19154 , y19155 , y19156 , y19157 , y19158 , y19159 , y19160 , y19161 , y19162 , y19163 , y19164 , y19165 , y19166 , y19167 , y19168 , y19169 , y19170 , y19171 , y19172 , y19173 , y19174 , y19175 , y19176 , y19177 , y19178 , y19179 , y19180 , y19181 , y19182 , y19183 , y19184 , y19185 , y19186 , y19187 , y19188 , y19189 , y19190 , y19191 , y19192 , y19193 , y19194 , y19195 , y19196 , y19197 , y19198 , y19199 , y19200 , y19201 , y19202 , y19203 , y19204 , y19205 , y19206 , y19207 , y19208 , y19209 , y19210 , y19211 , y19212 , y19213 , y19214 , y19215 , y19216 , y19217 , y19218 , y19219 , y19220 , y19221 , y19222 , y19223 , y19224 , y19225 , y19226 , y19227 , y19228 , y19229 , y19230 , y19231 , y19232 , y19233 , y19234 , y19235 , y19236 , y19237 , y19238 , y19239 , y19240 , y19241 , y19242 , y19243 , y19244 , y19245 , y19246 , y19247 , y19248 , y19249 , y19250 , y19251 , y19252 , y19253 , y19254 , y19255 , y19256 , y19257 , y19258 , y19259 , y19260 , y19261 , y19262 , y19263 , y19264 , y19265 , y19266 , y19267 , y19268 , y19269 , y19270 , y19271 , y19272 , y19273 , y19274 , y19275 , y19276 , y19277 , y19278 , y19279 , y19280 , y19281 , y19282 , y19283 , y19284 , y19285 , y19286 , y19287 , y19288 , y19289 , y19290 , y19291 , y19292 , y19293 , y19294 , y19295 , y19296 , y19297 , y19298 , y19299 , y19300 , y19301 , y19302 , y19303 , y19304 , y19305 , y19306 , y19307 , y19308 , y19309 , y19310 , y19311 , y19312 , y19313 , y19314 , y19315 , y19316 , y19317 , y19318 , y19319 , y19320 , y19321 , y19322 , y19323 , y19324 , y19325 , y19326 , y19327 , y19328 , y19329 , y19330 , y19331 , y19332 , y19333 , y19334 , y19335 , y19336 , y19337 , y19338 , y19339 , y19340 , y19341 , y19342 , y19343 , y19344 , y19345 , y19346 , y19347 , y19348 , y19349 , y19350 , y19351 , y19352 , y19353 , y19354 , y19355 , y19356 , y19357 , y19358 , y19359 , y19360 , y19361 , y19362 , y19363 , y19364 , y19365 , y19366 , y19367 , y19368 , y19369 , y19370 , y19371 , y19372 , y19373 , y19374 , y19375 , y19376 , y19377 , y19378 , y19379 , y19380 , y19381 , y19382 , y19383 , y19384 , y19385 , y19386 , y19387 , y19388 , y19389 , y19390 , y19391 , y19392 , y19393 , y19394 , y19395 , y19396 , y19397 , y19398 , y19399 , y19400 , y19401 , y19402 , y19403 , y19404 , y19405 , y19406 , y19407 , y19408 , y19409 , y19410 , y19411 , y19412 , y19413 , y19414 , y19415 , y19416 , y19417 , y19418 , y19419 , y19420 , y19421 , y19422 , y19423 , y19424 , y19425 , y19426 , y19427 , y19428 , y19429 , y19430 , y19431 , y19432 , y19433 , y19434 , y19435 , y19436 , y19437 , y19438 , y19439 , y19440 , y19441 , y19442 , y19443 , y19444 , y19445 , y19446 , y19447 , y19448 , y19449 , y19450 , y19451 , y19452 , y19453 , y19454 , y19455 , y19456 , y19457 , y19458 , y19459 , y19460 , y19461 , y19462 , y19463 , y19464 , y19465 , y19466 , y19467 , y19468 , y19469 , y19470 , y19471 , y19472 , y19473 , y19474 , y19475 , y19476 , y19477 , y19478 , y19479 , y19480 , y19481 , y19482 , y19483 , y19484 , y19485 , y19486 , y19487 , y19488 , y19489 , y19490 , y19491 , y19492 , y19493 , y19494 , y19495 , y19496 , y19497 , y19498 , y19499 , y19500 , y19501 , y19502 , y19503 , y19504 , y19505 , y19506 , y19507 , y19508 , y19509 , y19510 , y19511 , y19512 , y19513 , y19514 , y19515 , y19516 , y19517 , y19518 , y19519 , y19520 , y19521 , y19522 , y19523 , y19524 , y19525 , y19526 , y19527 , y19528 , y19529 , y19530 , y19531 , y19532 , y19533 , y19534 , y19535 , y19536 , y19537 , y19538 , y19539 , y19540 , y19541 , y19542 , y19543 , y19544 , y19545 , y19546 , y19547 , y19548 , y19549 , y19550 , y19551 , y19552 , y19553 , y19554 , y19555 , y19556 , y19557 , y19558 , y19559 , y19560 , y19561 , y19562 , y19563 , y19564 , y19565 , y19566 , y19567 , y19568 , y19569 , y19570 , y19571 , y19572 , y19573 , y19574 , y19575 , y19576 , y19577 , y19578 , y19579 , y19580 , y19581 , y19582 , y19583 , y19584 , y19585 , y19586 , y19587 , y19588 , y19589 , y19590 , y19591 , y19592 , y19593 , y19594 , y19595 , y19596 , y19597 , y19598 , y19599 , y19600 , y19601 , y19602 , y19603 , y19604 , y19605 , y19606 , y19607 , y19608 , y19609 , y19610 , y19611 , y19612 , y19613 , y19614 , y19615 , y19616 , y19617 , y19618 , y19619 , y19620 , y19621 , y19622 , y19623 , y19624 , y19625 , y19626 , y19627 , y19628 , y19629 , y19630 , y19631 , y19632 , y19633 , y19634 , y19635 , y19636 , y19637 , y19638 , y19639 , y19640 , y19641 , y19642 , y19643 , y19644 , y19645 , y19646 , y19647 , y19648 , y19649 , y19650 , y19651 , y19652 , y19653 , y19654 , y19655 , y19656 , y19657 , y19658 , y19659 , y19660 , y19661 , y19662 , y19663 , y19664 , y19665 , y19666 , y19667 , y19668 , y19669 , y19670 , y19671 , y19672 , y19673 , y19674 , y19675 , y19676 , y19677 , y19678 , y19679 , y19680 , y19681 , y19682 , y19683 , y19684 , y19685 , y19686 , y19687 , y19688 , y19689 , y19690 , y19691 , y19692 , y19693 , y19694 , y19695 , y19696 , y19697 , y19698 , y19699 , y19700 , y19701 , y19702 , y19703 , y19704 , y19705 , y19706 , y19707 , y19708 , y19709 , y19710 , y19711 , y19712 , y19713 , y19714 , y19715 , y19716 , y19717 , y19718 , y19719 , y19720 , y19721 , y19722 , y19723 , y19724 , y19725 , y19726 , y19727 , y19728 , y19729 , y19730 , y19731 , y19732 , y19733 , y19734 , y19735 , y19736 , y19737 , y19738 , y19739 , y19740 , y19741 , y19742 , y19743 , y19744 , y19745 , y19746 , y19747 , y19748 , y19749 , y19750 , y19751 , y19752 , y19753 , y19754 , y19755 , y19756 , y19757 , y19758 , y19759 , y19760 , y19761 , y19762 , y19763 , y19764 , y19765 , y19766 , y19767 , y19768 , y19769 , y19770 , y19771 , y19772 , y19773 , y19774 , y19775 , y19776 , y19777 , y19778 , y19779 , y19780 , y19781 , y19782 , y19783 , y19784 , y19785 , y19786 , y19787 , y19788 , y19789 , y19790 , y19791 , y19792 , y19793 , y19794 , y19795 , y19796 , y19797 , y19798 , y19799 , y19800 , y19801 , y19802 , y19803 , y19804 , y19805 , y19806 , y19807 , y19808 , y19809 , y19810 , y19811 , y19812 , y19813 , y19814 , y19815 , y19816 , y19817 , y19818 , y19819 , y19820 , y19821 , y19822 , y19823 , y19824 , y19825 , y19826 , y19827 , y19828 , y19829 , y19830 , y19831 , y19832 , y19833 , y19834 , y19835 , y19836 , y19837 , y19838 , y19839 , y19840 , y19841 , y19842 , y19843 , y19844 , y19845 , y19846 , y19847 , y19848 , y19849 , y19850 , y19851 , y19852 , y19853 , y19854 , y19855 , y19856 , y19857 , y19858 , y19859 , y19860 , y19861 , y19862 , y19863 , y19864 , y19865 , y19866 , y19867 , y19868 , y19869 , y19870 , y19871 , y19872 , y19873 , y19874 , y19875 , y19876 , y19877 , y19878 , y19879 , y19880 , y19881 , y19882 , y19883 , y19884 , y19885 , y19886 , y19887 , y19888 , y19889 , y19890 , y19891 , y19892 , y19893 , y19894 , y19895 , y19896 , y19897 , y19898 , y19899 , y19900 , y19901 , y19902 , y19903 , y19904 , y19905 , y19906 , y19907 , y19908 , y19909 , y19910 , y19911 , y19912 , y19913 , y19914 , y19915 , y19916 , y19917 , y19918 , y19919 , y19920 , y19921 , y19922 , y19923 , y19924 , y19925 , y19926 , y19927 , y19928 , y19929 , y19930 , y19931 , y19932 , y19933 , y19934 , y19935 , y19936 , y19937 , y19938 , y19939 , y19940 , y19941 , y19942 , y19943 , y19944 , y19945 , y19946 , y19947 , y19948 , y19949 , y19950 , y19951 , y19952 , y19953 , y19954 , y19955 , y19956 , y19957 , y19958 , y19959 , y19960 , y19961 , y19962 , y19963 , y19964 , y19965 , y19966 , y19967 , y19968 , y19969 , y19970 , y19971 , y19972 , y19973 , y19974 , y19975 , y19976 , y19977 , y19978 , y19979 , y19980 , y19981 , y19982 , y19983 , y19984 , y19985 , y19986 , y19987 , y19988 , y19989 , y19990 , y19991 , y19992 , y19993 , y19994 , y19995 , y19996 , y19997 , y19998 , y19999 , y20000 , y20001 , y20002 , y20003 , y20004 , y20005 , y20006 , y20007 , y20008 , y20009 , y20010 , y20011 , y20012 , y20013 , y20014 , y20015 , y20016 , y20017 , y20018 , y20019 , y20020 , y20021 , y20022 , y20023 , y20024 , y20025 , y20026 , y20027 , y20028 , y20029 , y20030 , y20031 , y20032 , y20033 , y20034 , y20035 , y20036 , y20037 , y20038 , y20039 , y20040 , y20041 , y20042 , y20043 , y20044 , y20045 , y20046 , y20047 , y20048 , y20049 , y20050 , y20051 , y20052 , y20053 , y20054 , y20055 , y20056 , y20057 , y20058 , y20059 , y20060 , y20061 , y20062 , y20063 , y20064 , y20065 , y20066 , y20067 , y20068 , y20069 , y20070 , y20071 , y20072 , y20073 , y20074 , y20075 , y20076 , y20077 , y20078 , y20079 , y20080 , y20081 , y20082 , y20083 , y20084 , y20085 , y20086 , y20087 , y20088 , y20089 , y20090 , y20091 , y20092 , y20093 , y20094 , y20095 , y20096 , y20097 , y20098 , y20099 , y20100 , y20101 , y20102 , y20103 , y20104 , y20105 , y20106 , y20107 , y20108 , y20109 , y20110 , y20111 , y20112 , y20113 , y20114 , y20115 , y20116 , y20117 , y20118 , y20119 , y20120 , y20121 , y20122 , y20123 , y20124 , y20125 , y20126 , y20127 , y20128 , y20129 , y20130 , y20131 , y20132 , y20133 , y20134 , y20135 , y20136 , y20137 , y20138 , y20139 , y20140 , y20141 , y20142 , y20143 , y20144 , y20145 , y20146 , y20147 , y20148 , y20149 , y20150 , y20151 , y20152 , y20153 , y20154 , y20155 , y20156 , y20157 , y20158 , y20159 , y20160 , y20161 , y20162 , y20163 , y20164 , y20165 , y20166 , y20167 , y20168 , y20169 , y20170 , y20171 , y20172 , y20173 , y20174 , y20175 , y20176 , y20177 , y20178 , y20179 , y20180 , y20181 , y20182 , y20183 , y20184 , y20185 , y20186 , y20187 , y20188 , y20189 , y20190 , y20191 , y20192 , y20193 , y20194 , y20195 , y20196 , y20197 , y20198 , y20199 , y20200 , y20201 , y20202 , y20203 , y20204 , y20205 , y20206 , y20207 , y20208 , y20209 , y20210 , y20211 , y20212 , y20213 , y20214 , y20215 , y20216 , y20217 , y20218 , y20219 , y20220 , y20221 , y20222 , y20223 , y20224 , y20225 , y20226 , y20227 , y20228 , y20229 , y20230 , y20231 , y20232 , y20233 , y20234 , y20235 , y20236 , y20237 , y20238 , y20239 , y20240 , y20241 , y20242 , y20243 , y20244 , y20245 , y20246 , y20247 , y20248 , y20249 , y20250 , y20251 , y20252 , y20253 , y20254 , y20255 , y20256 , y20257 , y20258 , y20259 , y20260 , y20261 , y20262 , y20263 , y20264 , y20265 , y20266 , y20267 , y20268 , y20269 , y20270 , y20271 , y20272 , y20273 , y20274 , y20275 , y20276 , y20277 , y20278 , y20279 , y20280 , y20281 , y20282 , y20283 , y20284 , y20285 , y20286 , y20287 , y20288 , y20289 , y20290 , y20291 , y20292 , y20293 , y20294 , y20295 , y20296 , y20297 , y20298 , y20299 , y20300 , y20301 , y20302 , y20303 , y20304 , y20305 , y20306 , y20307 , y20308 , y20309 , y20310 , y20311 , y20312 , y20313 , y20314 , y20315 , y20316 , y20317 , y20318 , y20319 , y20320 , y20321 , y20322 , y20323 , y20324 , y20325 , y20326 , y20327 , y20328 , y20329 , y20330 , y20331 , y20332 , y20333 , y20334 , y20335 , y20336 , y20337 , y20338 , y20339 , y20340 , y20341 , y20342 , y20343 , y20344 , y20345 , y20346 , y20347 , y20348 , y20349 , y20350 , y20351 , y20352 , y20353 , y20354 , y20355 , y20356 , y20357 , y20358 , y20359 , y20360 , y20361 , y20362 , y20363 , y20364 , y20365 , y20366 , y20367 , y20368 , y20369 , y20370 , y20371 , y20372 , y20373 , y20374 , y20375 , y20376 , y20377 , y20378 , y20379 , y20380 , y20381 , y20382 , y20383 , y20384 , y20385 , y20386 , y20387 , y20388 , y20389 , y20390 , y20391 , y20392 , y20393 , y20394 , y20395 , y20396 , y20397 , y20398 , y20399 , y20400 , y20401 , y20402 , y20403 , y20404 , y20405 , y20406 , y20407 , y20408 , y20409 , y20410 , y20411 , y20412 , y20413 , y20414 , y20415 , y20416 , y20417 , y20418 , y20419 , y20420 , y20421 , y20422 , y20423 , y20424 , y20425 , y20426 , y20427 , y20428 , y20429 , y20430 , y20431 , y20432 , y20433 , y20434 , y20435 , y20436 , y20437 , y20438 , y20439 , y20440 , y20441 , y20442 , y20443 , y20444 , y20445 , y20446 , y20447 , y20448 , y20449 , y20450 , y20451 , y20452 , y20453 , y20454 , y20455 , y20456 , y20457 , y20458 , y20459 , y20460 , y20461 , y20462 , y20463 , y20464 , y20465 , y20466 , y20467 , y20468 , y20469 , y20470 , y20471 , y20472 , y20473 , y20474 , y20475 , y20476 , y20477 , y20478 , y20479 , y20480 , y20481 , y20482 , y20483 , y20484 , y20485 , y20486 , y20487 , y20488 , y20489 , y20490 , y20491 , y20492 , y20493 , y20494 , y20495 , y20496 , y20497 , y20498 , y20499 , y20500 , y20501 , y20502 , y20503 , y20504 , y20505 , y20506 , y20507 , y20508 , y20509 , y20510 , y20511 , y20512 , y20513 , y20514 , y20515 , y20516 , y20517 , y20518 , y20519 , y20520 , y20521 , y20522 , y20523 , y20524 , y20525 , y20526 , y20527 , y20528 , y20529 , y20530 , y20531 , y20532 , y20533 , y20534 , y20535 , y20536 , y20537 , y20538 , y20539 , y20540 , y20541 , y20542 , y20543 , y20544 , y20545 , y20546 , y20547 , y20548 , y20549 , y20550 , y20551 , y20552 , y20553 , y20554 , y20555 , y20556 , y20557 , y20558 , y20559 , y20560 , y20561 , y20562 , y20563 , y20564 , y20565 , y20566 , y20567 , y20568 , y20569 , y20570 , y20571 , y20572 , y20573 , y20574 , y20575 , y20576 , y20577 , y20578 , y20579 , y20580 , y20581 , y20582 , y20583 , y20584 , y20585 , y20586 , y20587 , y20588 , y20589 , y20590 , y20591 , y20592 , y20593 , y20594 , y20595 , y20596 , y20597 , y20598 , y20599 , y20600 , y20601 , y20602 , y20603 , y20604 , y20605 , y20606 , y20607 , y20608 , y20609 , y20610 , y20611 , y20612 , y20613 , y20614 , y20615 , y20616 , y20617 , y20618 , y20619 , y20620 , y20621 , y20622 , y20623 , y20624 , y20625 , y20626 , y20627 , y20628 , y20629 , y20630 , y20631 , y20632 , y20633 , y20634 , y20635 , y20636 , y20637 , y20638 , y20639 , y20640 , y20641 , y20642 , y20643 , y20644 , y20645 , y20646 , y20647 , y20648 , y20649 , y20650 , y20651 , y20652 , y20653 , y20654 , y20655 , y20656 , y20657 , y20658 , y20659 , y20660 , y20661 , y20662 , y20663 , y20664 , y20665 , y20666 , y20667 , y20668 , y20669 , y20670 , y20671 , y20672 , y20673 , y20674 , y20675 , y20676 , y20677 , y20678 , y20679 , y20680 , y20681 , y20682 , y20683 , y20684 , y20685 , y20686 , y20687 , y20688 , y20689 , y20690 , y20691 , y20692 , y20693 , y20694 , y20695 , y20696 , y20697 , y20698 , y20699 , y20700 , y20701 , y20702 , y20703 , y20704 , y20705 , y20706 , y20707 , y20708 , y20709 , y20710 , y20711 , y20712 , y20713 , y20714 , y20715 , y20716 , y20717 , y20718 , y20719 , y20720 , y20721 , y20722 , y20723 , y20724 , y20725 , y20726 , y20727 , y20728 , y20729 , y20730 , y20731 , y20732 , y20733 , y20734 , y20735 , y20736 , y20737 , y20738 , y20739 , y20740 , y20741 , y20742 , y20743 , y20744 , y20745 , y20746 , y20747 , y20748 , y20749 , y20750 , y20751 , y20752 , y20753 , y20754 , y20755 , y20756 , y20757 , y20758 , y20759 , y20760 , y20761 , y20762 , y20763 , y20764 , y20765 , y20766 , y20767 , y20768 , y20769 , y20770 , y20771 , y20772 , y20773 , y20774 , y20775 , y20776 , y20777 , y20778 , y20779 , y20780 , y20781 , y20782 , y20783 , y20784 , y20785 , y20786 , y20787 , y20788 , y20789 , y20790 , y20791 , y20792 , y20793 , y20794 , y20795 , y20796 , y20797 , y20798 , y20799 , y20800 , y20801 , y20802 , y20803 , y20804 , y20805 , y20806 , y20807 , y20808 , y20809 , y20810 , y20811 , y20812 , y20813 , y20814 , y20815 , y20816 , y20817 , y20818 , y20819 , y20820 , y20821 , y20822 , y20823 , y20824 , y20825 , y20826 , y20827 , y20828 , y20829 , y20830 , y20831 , y20832 , y20833 , y20834 , y20835 , y20836 , y20837 , y20838 , y20839 , y20840 , y20841 , y20842 , y20843 , y20844 , y20845 , y20846 , y20847 , y20848 , y20849 , y20850 , y20851 , y20852 , y20853 , y20854 , y20855 , y20856 , y20857 , y20858 , y20859 , y20860 , y20861 , y20862 , y20863 , y20864 , y20865 , y20866 , y20867 , y20868 , y20869 , y20870 , y20871 , y20872 , y20873 , y20874 , y20875 , y20876 , y20877 , y20878 , y20879 , y20880 , y20881 , y20882 , y20883 , y20884 , y20885 , y20886 , y20887 , y20888 , y20889 , y20890 , y20891 , y20892 , y20893 , y20894 , y20895 , y20896 , y20897 , y20898 , y20899 , y20900 , y20901 , y20902 , y20903 , y20904 , y20905 , y20906 , y20907 , y20908 , y20909 , y20910 , y20911 , y20912 , y20913 , y20914 , y20915 , y20916 , y20917 , y20918 , y20919 , y20920 , y20921 , y20922 , y20923 , y20924 , y20925 , y20926 , y20927 , y20928 , y20929 , y20930 , y20931 , y20932 , y20933 , y20934 , y20935 , y20936 , y20937 , y20938 , y20939 , y20940 , y20941 , y20942 , y20943 , y20944 , y20945 , y20946 , y20947 , y20948 , y20949 , y20950 , y20951 , y20952 , y20953 , y20954 , y20955 , y20956 , y20957 , y20958 , y20959 , y20960 , y20961 , y20962 , y20963 , y20964 , y20965 , y20966 , y20967 , y20968 , y20969 , y20970 , y20971 , y20972 , y20973 , y20974 , y20975 , y20976 , y20977 , y20978 , y20979 , y20980 , y20981 , y20982 , y20983 , y20984 , y20985 , y20986 , y20987 , y20988 , y20989 , y20990 , y20991 , y20992 , y20993 , y20994 , y20995 , y20996 , y20997 , y20998 , y20999 , y21000 , y21001 , y21002 , y21003 , y21004 , y21005 , y21006 , y21007 , y21008 , y21009 , y21010 , y21011 , y21012 , y21013 , y21014 , y21015 , y21016 , y21017 , y21018 , y21019 , y21020 , y21021 , y21022 , y21023 , y21024 , y21025 , y21026 , y21027 , y21028 , y21029 , y21030 , y21031 , y21032 , y21033 , y21034 , y21035 , y21036 , y21037 , y21038 , y21039 , y21040 , y21041 , y21042 , y21043 , y21044 , y21045 , y21046 , y21047 , y21048 , y21049 , y21050 , y21051 , y21052 , y21053 , y21054 , y21055 , y21056 , y21057 , y21058 , y21059 , y21060 , y21061 , y21062 , y21063 , y21064 , y21065 , y21066 , y21067 , y21068 , y21069 , y21070 , y21071 , y21072 , y21073 , y21074 , y21075 , y21076 , y21077 , y21078 , y21079 , y21080 , y21081 , y21082 , y21083 , y21084 , y21085 , y21086 , y21087 , y21088 , y21089 , y21090 , y21091 , y21092 , y21093 , y21094 , y21095 , y21096 , y21097 , y21098 , y21099 , y21100 , y21101 , y21102 , y21103 , y21104 , y21105 , y21106 , y21107 , y21108 , y21109 , y21110 , y21111 , y21112 , y21113 , y21114 , y21115 , y21116 , y21117 , y21118 , y21119 , y21120 , y21121 , y21122 , y21123 , y21124 , y21125 , y21126 , y21127 , y21128 , y21129 , y21130 , y21131 , y21132 , y21133 , y21134 , y21135 , y21136 , y21137 , y21138 , y21139 , y21140 , y21141 , y21142 , y21143 , y21144 , y21145 , y21146 , y21147 , y21148 , y21149 , y21150 , y21151 , y21152 , y21153 , y21154 , y21155 , y21156 , y21157 , y21158 , y21159 , y21160 , y21161 , y21162 , y21163 , y21164 , y21165 , y21166 , y21167 , y21168 , y21169 , y21170 , y21171 , y21172 , y21173 , y21174 , y21175 , y21176 , y21177 , y21178 , y21179 , y21180 , y21181 , y21182 , y21183 , y21184 , y21185 , y21186 , y21187 , y21188 , y21189 , y21190 , y21191 , y21192 , y21193 , y21194 , y21195 , y21196 , y21197 , y21198 , y21199 , y21200 , y21201 , y21202 , y21203 , y21204 , y21205 , y21206 , y21207 , y21208 , y21209 , y21210 , y21211 , y21212 , y21213 , y21214 , y21215 , y21216 , y21217 , y21218 , y21219 , y21220 , y21221 , y21222 , y21223 , y21224 , y21225 , y21226 , y21227 , y21228 , y21229 , y21230 , y21231 , y21232 , y21233 , y21234 , y21235 , y21236 , y21237 , y21238 , y21239 , y21240 , y21241 , y21242 , y21243 , y21244 , y21245 , y21246 , y21247 , y21248 , y21249 , y21250 , y21251 , y21252 , y21253 , y21254 , y21255 , y21256 , y21257 , y21258 , y21259 , y21260 , y21261 , y21262 , y21263 , y21264 , y21265 , y21266 , y21267 , y21268 , y21269 , y21270 , y21271 , y21272 , y21273 , y21274 , y21275 , y21276 , y21277 , y21278 , y21279 , y21280 , y21281 , y21282 , y21283 , y21284 , y21285 , y21286 , y21287 , y21288 , y21289 , y21290 , y21291 , y21292 , y21293 , y21294 , y21295 , y21296 , y21297 , y21298 , y21299 , y21300 , y21301 , y21302 , y21303 , y21304 , y21305 , y21306 , y21307 , y21308 , y21309 , y21310 , y21311 , y21312 , y21313 , y21314 , y21315 , y21316 , y21317 , y21318 , y21319 , y21320 , y21321 , y21322 , y21323 , y21324 , y21325 , y21326 , y21327 , y21328 , y21329 , y21330 , y21331 , y21332 , y21333 , y21334 , y21335 , y21336 , y21337 , y21338 , y21339 , y21340 , y21341 , y21342 , y21343 , y21344 , y21345 , y21346 , y21347 , y21348 , y21349 , y21350 , y21351 , y21352 , y21353 , y21354 , y21355 , y21356 , y21357 , y21358 , y21359 , y21360 , y21361 , y21362 , y21363 , y21364 , y21365 , y21366 , y21367 , y21368 , y21369 , y21370 , y21371 , y21372 , y21373 , y21374 , y21375 , y21376 , y21377 , y21378 , y21379 , y21380 , y21381 , y21382 , y21383 , y21384 , y21385 , y21386 , y21387 , y21388 , y21389 , y21390 , y21391 , y21392 , y21393 , y21394 , y21395 , y21396 , y21397 , y21398 , y21399 , y21400 , y21401 , y21402 , y21403 , y21404 , y21405 , y21406 , y21407 , y21408 , y21409 , y21410 , y21411 , y21412 , y21413 , y21414 , y21415 , y21416 , y21417 , y21418 , y21419 , y21420 , y21421 , y21422 , y21423 , y21424 , y21425 , y21426 , y21427 , y21428 , y21429 , y21430 , y21431 , y21432 , y21433 , y21434 , y21435 , y21436 , y21437 , y21438 , y21439 , y21440 , y21441 , y21442 , y21443 , y21444 , y21445 , y21446 , y21447 , y21448 , y21449 , y21450 , y21451 , y21452 , y21453 , y21454 , y21455 , y21456 , y21457 , y21458 , y21459 , y21460 , y21461 , y21462 , y21463 , y21464 , y21465 , y21466 , y21467 , y21468 , y21469 , y21470 , y21471 , y21472 , y21473 , y21474 , y21475 , y21476 , y21477 , y21478 , y21479 , y21480 , y21481 , y21482 , y21483 , y21484 , y21485 , y21486 , y21487 , y21488 , y21489 , y21490 , y21491 , y21492 , y21493 , y21494 , y21495 , y21496 , y21497 , y21498 , y21499 , y21500 , y21501 , y21502 , y21503 , y21504 , y21505 , y21506 , y21507 , y21508 , y21509 , y21510 , y21511 , y21512 , y21513 , y21514 , y21515 , y21516 , y21517 , y21518 , y21519 , y21520 , y21521 , y21522 , y21523 , y21524 , y21525 , y21526 , y21527 , y21528 , y21529 , y21530 , y21531 , y21532 , y21533 , y21534 , y21535 , y21536 , y21537 , y21538 , y21539 , y21540 , y21541 , y21542 , y21543 , y21544 , y21545 , y21546 , y21547 , y21548 , y21549 , y21550 , y21551 , y21552 , y21553 , y21554 , y21555 , y21556 , y21557 , y21558 , y21559 , y21560 , y21561 , y21562 , y21563 , y21564 , y21565 , y21566 , y21567 , y21568 , y21569 , y21570 , y21571 , y21572 , y21573 , y21574 , y21575 , y21576 , y21577 , y21578 , y21579 , y21580 , y21581 , y21582 , y21583 , y21584 , y21585 , y21586 , y21587 , y21588 , y21589 , y21590 , y21591 , y21592 , y21593 , y21594 , y21595 , y21596 , y21597 , y21598 , y21599 , y21600 , y21601 , y21602 , y21603 , y21604 , y21605 , y21606 , y21607 , y21608 , y21609 , y21610 , y21611 , y21612 , y21613 , y21614 , y21615 , y21616 , y21617 , y21618 , y21619 , y21620 , y21621 , y21622 , y21623 , y21624 , y21625 , y21626 , y21627 , y21628 , y21629 , y21630 , y21631 , y21632 , y21633 , y21634 , y21635 , y21636 , y21637 , y21638 , y21639 , y21640 , y21641 , y21642 , y21643 , y21644 , y21645 , y21646 , y21647 , y21648 , y21649 , y21650 , y21651 , y21652 , y21653 , y21654 , y21655 , y21656 , y21657 , y21658 , y21659 , y21660 , y21661 , y21662 , y21663 , y21664 , y21665 , y21666 , y21667 , y21668 , y21669 , y21670 , y21671 , y21672 , y21673 , y21674 , y21675 , y21676 , y21677 , y21678 , y21679 , y21680 , y21681 , y21682 , y21683 , y21684 , y21685 , y21686 , y21687 , y21688 , y21689 , y21690 , y21691 , y21692 , y21693 , y21694 , y21695 , y21696 , y21697 , y21698 , y21699 , y21700 , y21701 , y21702 , y21703 , y21704 , y21705 , y21706 , y21707 , y21708 , y21709 , y21710 , y21711 , y21712 , y21713 , y21714 , y21715 , y21716 , y21717 , y21718 , y21719 , y21720 , y21721 , y21722 , y21723 , y21724 , y21725 , y21726 , y21727 , y21728 , y21729 , y21730 , y21731 , y21732 , y21733 , y21734 , y21735 , y21736 , y21737 , y21738 , y21739 , y21740 , y21741 , y21742 , y21743 , y21744 , y21745 , y21746 , y21747 , y21748 , y21749 , y21750 , y21751 , y21752 , y21753 , y21754 , y21755 , y21756 , y21757 , y21758 , y21759 , y21760 , y21761 , y21762 , y21763 , y21764 , y21765 , y21766 , y21767 , y21768 , y21769 , y21770 , y21771 , y21772 , y21773 , y21774 , y21775 , y21776 , y21777 , y21778 , y21779 , y21780 , y21781 , y21782 , y21783 , y21784 , y21785 , y21786 , y21787 , y21788 , y21789 , y21790 , y21791 , y21792 , y21793 , y21794 , y21795 , y21796 , y21797 , y21798 , y21799 , y21800 , y21801 , y21802 , y21803 , y21804 , y21805 , y21806 , y21807 , y21808 , y21809 , y21810 , y21811 , y21812 , y21813 , y21814 , y21815 , y21816 , y21817 , y21818 , y21819 , y21820 , y21821 , y21822 , y21823 , y21824 , y21825 , y21826 , y21827 , y21828 , y21829 , y21830 , y21831 , y21832 , y21833 , y21834 , y21835 , y21836 , y21837 , y21838 , y21839 , y21840 , y21841 , y21842 , y21843 , y21844 , y21845 , y21846 , y21847 , y21848 , y21849 , y21850 , y21851 , y21852 , y21853 , y21854 , y21855 , y21856 , y21857 , y21858 , y21859 , y21860 , y21861 , y21862 , y21863 , y21864 , y21865 , y21866 , y21867 , y21868 , y21869 , y21870 , y21871 , y21872 , y21873 , y21874 , y21875 , y21876 , y21877 , y21878 , y21879 , y21880 , y21881 , y21882 , y21883 , y21884 , y21885 , y21886 , y21887 , y21888 , y21889 , y21890 , y21891 , y21892 , y21893 , y21894 , y21895 , y21896 , y21897 , y21898 , y21899 , y21900 , y21901 , y21902 , y21903 , y21904 , y21905 , y21906 , y21907 , y21908 , y21909 , y21910 , y21911 , y21912 , y21913 , y21914 , y21915 , y21916 , y21917 , y21918 , y21919 , y21920 , y21921 , y21922 , y21923 , y21924 , y21925 , y21926 , y21927 , y21928 , y21929 , y21930 , y21931 , y21932 , y21933 , y21934 , y21935 , y21936 , y21937 , y21938 , y21939 , y21940 , y21941 , y21942 , y21943 , y21944 , y21945 , y21946 , y21947 , y21948 , y21949 , y21950 , y21951 , y21952 , y21953 , y21954 , y21955 , y21956 , y21957 , y21958 , y21959 , y21960 , y21961 , y21962 , y21963 , y21964 , y21965 , y21966 , y21967 , y21968 , y21969 , y21970 , y21971 , y21972 , y21973 , y21974 , y21975 , y21976 , y21977 , y21978 , y21979 , y21980 , y21981 , y21982 , y21983 , y21984 , y21985 , y21986 , y21987 , y21988 , y21989 , y21990 , y21991 , y21992 , y21993 , y21994 , y21995 , y21996 , y21997 , y21998 , y21999 , y22000 , y22001 , y22002 , y22003 , y22004 , y22005 , y22006 , y22007 , y22008 , y22009 , y22010 , y22011 , y22012 , y22013 , y22014 , y22015 , y22016 , y22017 , y22018 , y22019 , y22020 , y22021 , y22022 , y22023 , y22024 , y22025 , y22026 , y22027 , y22028 , y22029 , y22030 , y22031 , y22032 , y22033 , y22034 , y22035 , y22036 , y22037 , y22038 , y22039 , y22040 , y22041 , y22042 , y22043 , y22044 , y22045 , y22046 , y22047 , y22048 , y22049 , y22050 , y22051 , y22052 , y22053 , y22054 , y22055 , y22056 , y22057 , y22058 , y22059 , y22060 , y22061 , y22062 , y22063 , y22064 , y22065 , y22066 , y22067 , y22068 , y22069 , y22070 , y22071 , y22072 , y22073 , y22074 , y22075 , y22076 , y22077 , y22078 , y22079 , y22080 , y22081 , y22082 , y22083 , y22084 , y22085 , y22086 , y22087 , y22088 , y22089 , y22090 , y22091 , y22092 , y22093 , y22094 , y22095 , y22096 , y22097 , y22098 , y22099 , y22100 , y22101 , y22102 , y22103 , y22104 , y22105 , y22106 , y22107 , y22108 , y22109 , y22110 , y22111 , y22112 , y22113 , y22114 , y22115 , y22116 , y22117 , y22118 , y22119 , y22120 , y22121 , y22122 , y22123 , y22124 , y22125 , y22126 , y22127 , y22128 , y22129 , y22130 , y22131 , y22132 , y22133 , y22134 , y22135 , y22136 , y22137 , y22138 , y22139 , y22140 , y22141 , y22142 , y22143 , y22144 , y22145 , y22146 , y22147 , y22148 , y22149 , y22150 , y22151 , y22152 , y22153 , y22154 , y22155 , y22156 , y22157 , y22158 , y22159 , y22160 , y22161 , y22162 , y22163 , y22164 , y22165 , y22166 , y22167 , y22168 , y22169 , y22170 , y22171 , y22172 , y22173 , y22174 , y22175 , y22176 , y22177 , y22178 , y22179 , y22180 , y22181 , y22182 , y22183 , y22184 , y22185 , y22186 , y22187 , y22188 , y22189 , y22190 , y22191 , y22192 , y22193 , y22194 , y22195 , y22196 , y22197 , y22198 , y22199 , y22200 , y22201 , y22202 , y22203 , y22204 , y22205 , y22206 , y22207 , y22208 , y22209 , y22210 , y22211 , y22212 , y22213 , y22214 , y22215 , y22216 , y22217 , y22218 , y22219 , y22220 , y22221 , y22222 , y22223 , y22224 , y22225 , y22226 , y22227 , y22228 , y22229 , y22230 , y22231 , y22232 , y22233 , y22234 , y22235 , y22236 , y22237 , y22238 , y22239 , y22240 , y22241 , y22242 , y22243 , y22244 , y22245 , y22246 , y22247 , y22248 , y22249 , y22250 , y22251 , y22252 , y22253 , y22254 , y22255 , y22256 , y22257 , y22258 , y22259 , y22260 , y22261 , y22262 , y22263 , y22264 , y22265 , y22266 , y22267 , y22268 , y22269 , y22270 , y22271 , y22272 , y22273 , y22274 , y22275 , y22276 , y22277 , y22278 , y22279 , y22280 , y22281 , y22282 , y22283 , y22284 , y22285 , y22286 , y22287 , y22288 , y22289 , y22290 , y22291 , y22292 , y22293 , y22294 , y22295 , y22296 , y22297 , y22298 , y22299 , y22300 , y22301 , y22302 , y22303 , y22304 , y22305 , y22306 , y22307 , y22308 , y22309 , y22310 , y22311 , y22312 , y22313 , y22314 , y22315 , y22316 , y22317 , y22318 , y22319 , y22320 , y22321 , y22322 , y22323 , y22324 , y22325 , y22326 , y22327 , y22328 , y22329 , y22330 , y22331 , y22332 , y22333 , y22334 , y22335 , y22336 , y22337 , y22338 , y22339 , y22340 , y22341 , y22342 , y22343 , y22344 , y22345 , y22346 , y22347 , y22348 , y22349 , y22350 , y22351 , y22352 , y22353 , y22354 , y22355 , y22356 , y22357 , y22358 , y22359 , y22360 , y22361 , y22362 , y22363 , y22364 , y22365 , y22366 , y22367 , y22368 , y22369 , y22370 , y22371 , y22372 , y22373 , y22374 , y22375 , y22376 , y22377 , y22378 , y22379 , y22380 , y22381 , y22382 , y22383 , y22384 , y22385 , y22386 , y22387 , y22388 , y22389 , y22390 , y22391 , y22392 , y22393 , y22394 , y22395 , y22396 , y22397 , y22398 , y22399 , y22400 , y22401 , y22402 , y22403 , y22404 , y22405 , y22406 , y22407 , y22408 , y22409 , y22410 , y22411 , y22412 , y22413 , y22414 , y22415 , y22416 , y22417 , y22418 , y22419 , y22420 , y22421 , y22422 , y22423 , y22424 , y22425 , y22426 , y22427 , y22428 , y22429 , y22430 , y22431 , y22432 , y22433 , y22434 , y22435 , y22436 , y22437 , y22438 , y22439 , y22440 , y22441 , y22442 , y22443 , y22444 , y22445 , y22446 , y22447 , y22448 , y22449 , y22450 , y22451 , y22452 , y22453 , y22454 , y22455 , y22456 , y22457 , y22458 , y22459 , y22460 , y22461 , y22462 , y22463 , y22464 , y22465 , y22466 , y22467 , y22468 , y22469 , y22470 , y22471 , y22472 , y22473 , y22474 , y22475 , y22476 , y22477 , y22478 , y22479 , y22480 , y22481 , y22482 , y22483 , y22484 , y22485 , y22486 , y22487 , y22488 , y22489 , y22490 , y22491 , y22492 , y22493 , y22494 , y22495 , y22496 , y22497 , y22498 , y22499 , y22500 , y22501 , y22502 , y22503 , y22504 , y22505 , y22506 , y22507 , y22508 , y22509 , y22510 , y22511 , y22512 , y22513 , y22514 , y22515 , y22516 , y22517 , y22518 , y22519 , y22520 , y22521 , y22522 , y22523 , y22524 , y22525 , y22526 , y22527 , y22528 , y22529 , y22530 , y22531 , y22532 , y22533 , y22534 , y22535 , y22536 , y22537 , y22538 , y22539 , y22540 , y22541 , y22542 , y22543 , y22544 , y22545 , y22546 , y22547 , y22548 , y22549 , y22550 , y22551 , y22552 , y22553 , y22554 , y22555 , y22556 , y22557 , y22558 , y22559 , y22560 , y22561 , y22562 , y22563 , y22564 , y22565 , y22566 , y22567 , y22568 , y22569 , y22570 , y22571 , y22572 , y22573 , y22574 , y22575 , y22576 , y22577 , y22578 , y22579 , y22580 , y22581 , y22582 , y22583 , y22584 , y22585 , y22586 , y22587 , y22588 , y22589 , y22590 , y22591 , y22592 , y22593 , y22594 , y22595 , y22596 , y22597 , y22598 , y22599 , y22600 , y22601 , y22602 , y22603 , y22604 , y22605 , y22606 , y22607 , y22608 , y22609 , y22610 , y22611 , y22612 , y22613 , y22614 , y22615 , y22616 , y22617 , y22618 , y22619 , y22620 , y22621 , y22622 , y22623 , y22624 , y22625 , y22626 , y22627 , y22628 , y22629 , y22630 , y22631 , y22632 , y22633 , y22634 , y22635 , y22636 , y22637 , y22638 , y22639 , y22640 , y22641 , y22642 , y22643 , y22644 , y22645 , y22646 , y22647 , y22648 , y22649 , y22650 , y22651 , y22652 , y22653 , y22654 , y22655 , y22656 , y22657 , y22658 , y22659 , y22660 , y22661 , y22662 , y22663 , y22664 , y22665 , y22666 , y22667 , y22668 , y22669 , y22670 , y22671 , y22672 , y22673 , y22674 , y22675 , y22676 , y22677 , y22678 , y22679 , y22680 , y22681 , y22682 , y22683 , y22684 , y22685 , y22686 , y22687 , y22688 , y22689 , y22690 , y22691 , y22692 , y22693 , y22694 , y22695 , y22696 , y22697 , y22698 , y22699 , y22700 , y22701 , y22702 , y22703 , y22704 , y22705 , y22706 , y22707 , y22708 , y22709 , y22710 , y22711 , y22712 , y22713 , y22714 , y22715 , y22716 , y22717 , y22718 , y22719 , y22720 , y22721 , y22722 , y22723 , y22724 , y22725 , y22726 , y22727 , y22728 , y22729 , y22730 , y22731 , y22732 , y22733 , y22734 , y22735 , y22736 , y22737 , y22738 , y22739 , y22740 , y22741 , y22742 , y22743 , y22744 , y22745 , y22746 , y22747 , y22748 , y22749 , y22750 , y22751 , y22752 , y22753 , y22754 , y22755 , y22756 , y22757 , y22758 , y22759 , y22760 , y22761 , y22762 , y22763 , y22764 , y22765 , y22766 , y22767 , y22768 , y22769 , y22770 , y22771 , y22772 , y22773 , y22774 , y22775 , y22776 , y22777 , y22778 , y22779 , y22780 , y22781 , y22782 , y22783 , y22784 , y22785 , y22786 , y22787 , y22788 , y22789 , y22790 , y22791 , y22792 , y22793 , y22794 , y22795 , y22796 , y22797 , y22798 , y22799 , y22800 , y22801 , y22802 , y22803 , y22804 , y22805 , y22806 , y22807 , y22808 , y22809 , y22810 , y22811 , y22812 , y22813 , y22814 , y22815 , y22816 , y22817 , y22818 , y22819 , y22820 , y22821 , y22822 , y22823 , y22824 , y22825 , y22826 , y22827 , y22828 , y22829 , y22830 , y22831 , y22832 , y22833 , y22834 , y22835 , y22836 , y22837 , y22838 , y22839 , y22840 , y22841 , y22842 , y22843 , y22844 , y22845 , y22846 , y22847 , y22848 , y22849 , y22850 , y22851 , y22852 , y22853 , y22854 , y22855 , y22856 , y22857 , y22858 , y22859 , y22860 , y22861 , y22862 , y22863 , y22864 , y22865 , y22866 , y22867 , y22868 , y22869 , y22870 , y22871 , y22872 , y22873 , y22874 , y22875 , y22876 , y22877 , y22878 , y22879 , y22880 , y22881 , y22882 , y22883 , y22884 , y22885 , y22886 , y22887 , y22888 , y22889 , y22890 , y22891 , y22892 , y22893 , y22894 , y22895 , y22896 , y22897 , y22898 , y22899 , y22900 , y22901 , y22902 , y22903 , y22904 , y22905 , y22906 , y22907 , y22908 , y22909 , y22910 , y22911 , y22912 , y22913 , y22914 , y22915 , y22916 , y22917 , y22918 , y22919 , y22920 , y22921 , y22922 , y22923 , y22924 , y22925 , y22926 , y22927 , y22928 , y22929 , y22930 , y22931 , y22932 , y22933 , y22934 , y22935 , y22936 , y22937 , y22938 , y22939 , y22940 , y22941 , y22942 , y22943 , y22944 , y22945 , y22946 , y22947 , y22948 , y22949 , y22950 , y22951 , y22952 , y22953 , y22954 , y22955 , y22956 , y22957 , y22958 , y22959 , y22960 , y22961 , y22962 , y22963 , y22964 , y22965 , y22966 , y22967 , y22968 , y22969 , y22970 , y22971 , y22972 , y22973 , y22974 , y22975 , y22976 , y22977 , y22978 , y22979 , y22980 , y22981 , y22982 , y22983 , y22984 , y22985 , y22986 , y22987 , y22988 , y22989 , y22990 , y22991 , y22992 , y22993 , y22994 , y22995 , y22996 , y22997 , y22998 , y22999 , y23000 , y23001 , y23002 , y23003 , y23004 , y23005 , y23006 , y23007 , y23008 , y23009 , y23010 , y23011 , y23012 , y23013 , y23014 , y23015 , y23016 , y23017 , y23018 , y23019 , y23020 , y23021 , y23022 , y23023 , y23024 , y23025 , y23026 , y23027 , y23028 , y23029 , y23030 , y23031 , y23032 , y23033 , y23034 , y23035 , y23036 , y23037 , y23038 , y23039 , y23040 , y23041 , y23042 , y23043 , y23044 , y23045 , y23046 , y23047 , y23048 , y23049 , y23050 , y23051 , y23052 , y23053 , y23054 , y23055 , y23056 , y23057 , y23058 , y23059 , y23060 , y23061 , y23062 , y23063 , y23064 , y23065 , y23066 , y23067 , y23068 , y23069 , y23070 , y23071 , y23072 , y23073 , y23074 , y23075 , y23076 , y23077 , y23078 , y23079 , y23080 , y23081 , y23082 , y23083 , y23084 , y23085 , y23086 , y23087 , y23088 , y23089 , y23090 , y23091 , y23092 , y23093 , y23094 , y23095 , y23096 , y23097 , y23098 , y23099 , y23100 , y23101 , y23102 , y23103 , y23104 , y23105 , y23106 , y23107 , y23108 , y23109 , y23110 , y23111 , y23112 , y23113 , y23114 , y23115 , y23116 , y23117 , y23118 , y23119 , y23120 , y23121 , y23122 , y23123 , y23124 , y23125 , y23126 , y23127 , y23128 , y23129 , y23130 , y23131 , y23132 , y23133 , y23134 , y23135 , y23136 , y23137 , y23138 , y23139 , y23140 , y23141 , y23142 , y23143 , y23144 , y23145 , y23146 , y23147 , y23148 , y23149 , y23150 , y23151 , y23152 , y23153 , y23154 , y23155 , y23156 , y23157 , y23158 , y23159 , y23160 , y23161 , y23162 , y23163 , y23164 , y23165 , y23166 , y23167 , y23168 , y23169 , y23170 , y23171 , y23172 , y23173 , y23174 , y23175 , y23176 , y23177 , y23178 , y23179 , y23180 , y23181 , y23182 , y23183 , y23184 , y23185 , y23186 , y23187 , y23188 , y23189 , y23190 , y23191 , y23192 , y23193 , y23194 , y23195 , y23196 , y23197 , y23198 , y23199 , y23200 , y23201 , y23202 , y23203 , y23204 , y23205 , y23206 , y23207 , y23208 , y23209 , y23210 , y23211 , y23212 , y23213 , y23214 , y23215 , y23216 , y23217 , y23218 , y23219 , y23220 , y23221 , y23222 , y23223 , y23224 , y23225 , y23226 , y23227 , y23228 , y23229 , y23230 , y23231 , y23232 , y23233 , y23234 , y23235 , y23236 , y23237 , y23238 , y23239 , y23240 , y23241 , y23242 , y23243 , y23244 , y23245 , y23246 , y23247 , y23248 , y23249 , y23250 , y23251 , y23252 , y23253 , y23254 , y23255 , y23256 , y23257 , y23258 , y23259 , y23260 , y23261 , y23262 , y23263 , y23264 , y23265 , y23266 , y23267 , y23268 , y23269 , y23270 , y23271 , y23272 , y23273 , y23274 , y23275 , y23276 , y23277 , y23278 , y23279 , y23280 , y23281 , y23282 , y23283 , y23284 , y23285 , y23286 , y23287 , y23288 , y23289 , y23290 , y23291 , y23292 , y23293 , y23294 , y23295 , y23296 , y23297 , y23298 , y23299 , y23300 , y23301 , y23302 , y23303 , y23304 , y23305 , y23306 , y23307 , y23308 , y23309 , y23310 , y23311 , y23312 , y23313 , y23314 , y23315 , y23316 , y23317 , y23318 , y23319 , y23320 , y23321 , y23322 , y23323 , y23324 , y23325 , y23326 , y23327 , y23328 , y23329 , y23330 , y23331 , y23332 , y23333 , y23334 , y23335 , y23336 , y23337 , y23338 , y23339 , y23340 , y23341 , y23342 , y23343 , y23344 , y23345 , y23346 , y23347 , y23348 , y23349 , y23350 , y23351 , y23352 , y23353 , y23354 , y23355 , y23356 , y23357 , y23358 , y23359 , y23360 , y23361 , y23362 , y23363 , y23364 , y23365 , y23366 , y23367 , y23368 , y23369 , y23370 , y23371 , y23372 , y23373 , y23374 , y23375 , y23376 , y23377 , y23378 , y23379 , y23380 , y23381 , y23382 , y23383 , y23384 , y23385 , y23386 , y23387 , y23388 , y23389 , y23390 , y23391 , y23392 , y23393 , y23394 , y23395 , y23396 , y23397 , y23398 , y23399 , y23400 , y23401 , y23402 , y23403 , y23404 , y23405 , y23406 , y23407 , y23408 , y23409 , y23410 , y23411 , y23412 , y23413 , y23414 , y23415 , y23416 , y23417 , y23418 , y23419 , y23420 , y23421 , y23422 , y23423 , y23424 , y23425 , y23426 , y23427 , y23428 , y23429 , y23430 , y23431 , y23432 , y23433 , y23434 , y23435 , y23436 , y23437 , y23438 , y23439 , y23440 , y23441 , y23442 , y23443 , y23444 , y23445 , y23446 , y23447 , y23448 , y23449 , y23450 , y23451 , y23452 , y23453 , y23454 , y23455 , y23456 , y23457 , y23458 , y23459 , y23460 , y23461 , y23462 , y23463 , y23464 , y23465 , y23466 , y23467 , y23468 , y23469 , y23470 , y23471 , y23472 , y23473 , y23474 , y23475 , y23476 , y23477 , y23478 , y23479 , y23480 , y23481 , y23482 , y23483 , y23484 , y23485 , y23486 , y23487 , y23488 , y23489 , y23490 , y23491 , y23492 , y23493 , y23494 , y23495 , y23496 , y23497 , y23498 , y23499 , y23500 , y23501 , y23502 , y23503 , y23504 , y23505 , y23506 , y23507 , y23508 , y23509 , y23510 , y23511 , y23512 , y23513 , y23514 , y23515 , y23516 , y23517 , y23518 , y23519 , y23520 , y23521 , y23522 , y23523 , y23524 , y23525 , y23526 , y23527 , y23528 , y23529 , y23530 , y23531 , y23532 , y23533 , y23534 , y23535 , y23536 , y23537 , y23538 , y23539 , y23540 , y23541 , y23542 , y23543 , y23544 , y23545 , y23546 , y23547 , y23548 , y23549 , y23550 , y23551 , y23552 , y23553 , y23554 , y23555 , y23556 , y23557 , y23558 , y23559 , y23560 , y23561 , y23562 , y23563 , y23564 , y23565 , y23566 , y23567 , y23568 , y23569 , y23570 , y23571 , y23572 , y23573 , y23574 , y23575 , y23576 , y23577 , y23578 , y23579 , y23580 , y23581 , y23582 , y23583 , y23584 , y23585 , y23586 , y23587 , y23588 , y23589 , y23590 , y23591 , y23592 , y23593 , y23594 , y23595 , y23596 , y23597 , y23598 , y23599 , y23600 , y23601 , y23602 , y23603 , y23604 , y23605 , y23606 , y23607 , y23608 , y23609 , y23610 , y23611 , y23612 , y23613 , y23614 , y23615 , y23616 , y23617 , y23618 , y23619 , y23620 , y23621 , y23622 , y23623 , y23624 , y23625 , y23626 , y23627 , y23628 , y23629 , y23630 , y23631 , y23632 , y23633 , y23634 , y23635 , y23636 , y23637 , y23638 , y23639 , y23640 , y23641 , y23642 , y23643 , y23644 , y23645 , y23646 , y23647 , y23648 , y23649 , y23650 , y23651 , y23652 , y23653 , y23654 , y23655 , y23656 , y23657 , y23658 , y23659 , y23660 , y23661 , y23662 , y23663 , y23664 , y23665 , y23666 , y23667 , y23668 , y23669 , y23670 , y23671 , y23672 , y23673 , y23674 , y23675 , y23676 , y23677 , y23678 , y23679 , y23680 , y23681 , y23682 , y23683 , y23684 , y23685 , y23686 , y23687 , y23688 , y23689 , y23690 , y23691 , y23692 , y23693 , y23694 , y23695 , y23696 , y23697 , y23698 , y23699 , y23700 , y23701 , y23702 , y23703 , y23704 , y23705 , y23706 , y23707 , y23708 , y23709 , y23710 , y23711 , y23712 , y23713 , y23714 , y23715 , y23716 , y23717 , y23718 , y23719 , y23720 , y23721 , y23722 , y23723 , y23724 , y23725 , y23726 , y23727 , y23728 , y23729 , y23730 , y23731 , y23732 , y23733 , y23734 , y23735 , y23736 , y23737 , y23738 , y23739 , y23740 , y23741 , y23742 , y23743 , y23744 , y23745 , y23746 , y23747 , y23748 , y23749 , y23750 , y23751 , y23752 , y23753 , y23754 , y23755 , y23756 , y23757 , y23758 , y23759 , y23760 , y23761 , y23762 , y23763 , y23764 , y23765 , y23766 , y23767 , y23768 , y23769 , y23770 , y23771 , y23772 , y23773 , y23774 , y23775 , y23776 , y23777 , y23778 , y23779 , y23780 , y23781 , y23782 , y23783 , y23784 , y23785 , y23786 , y23787 , y23788 , y23789 , y23790 , y23791 , y23792 , y23793 , y23794 , y23795 , y23796 , y23797 , y23798 , y23799 , y23800 , y23801 , y23802 , y23803 , y23804 , y23805 , y23806 , y23807 , y23808 , y23809 , y23810 , y23811 , y23812 , y23813 , y23814 , y23815 , y23816 , y23817 , y23818 , y23819 , y23820 , y23821 , y23822 , y23823 , y23824 , y23825 , y23826 , y23827 , y23828 , y23829 , y23830 , y23831 , y23832 , y23833 , y23834 , y23835 , y23836 , y23837 , y23838 , y23839 , y23840 , y23841 , y23842 , y23843 , y23844 , y23845 , y23846 , y23847 , y23848 , y23849 , y23850 , y23851 , y23852 , y23853 , y23854 , y23855 , y23856 , y23857 , y23858 , y23859 , y23860 , y23861 , y23862 , y23863 , y23864 , y23865 , y23866 , y23867 , y23868 , y23869 , y23870 , y23871 , y23872 , y23873 , y23874 , y23875 , y23876 , y23877 , y23878 , y23879 , y23880 , y23881 , y23882 , y23883 , y23884 , y23885 , y23886 , y23887 , y23888 , y23889 , y23890 , y23891 , y23892 , y23893 , y23894 , y23895 , y23896 , y23897 , y23898 , y23899 , y23900 , y23901 , y23902 , y23903 , y23904 , y23905 , y23906 , y23907 , y23908 , y23909 , y23910 , y23911 , y23912 , y23913 , y23914 , y23915 , y23916 , y23917 , y23918 , y23919 , y23920 , y23921 , y23922 , y23923 , y23924 , y23925 , y23926 , y23927 , y23928 , y23929 , y23930 , y23931 , y23932 , y23933 , y23934 , y23935 , y23936 , y23937 , y23938 , y23939 , y23940 , y23941 , y23942 , y23943 , y23944 , y23945 , y23946 , y23947 , y23948 , y23949 , y23950 , y23951 , y23952 , y23953 , y23954 , y23955 , y23956 , y23957 , y23958 , y23959 , y23960 , y23961 , y23962 , y23963 , y23964 , y23965 , y23966 , y23967 , y23968 , y23969 , y23970 , y23971 , y23972 , y23973 , y23974 , y23975 , y23976 , y23977 , y23978 , y23979 , y23980 , y23981 , y23982 , y23983 , y23984 , y23985 , y23986 , y23987 , y23988 , y23989 , y23990 , y23991 , y23992 , y23993 , y23994 , y23995 , y23996 , y23997 , y23998 , y23999 , y24000 , y24001 , y24002 , y24003 , y24004 , y24005 , y24006 , y24007 , y24008 , y24009 , y24010 , y24011 , y24012 , y24013 , y24014 , y24015 , y24016 , y24017 , y24018 , y24019 , y24020 , y24021 , y24022 , y24023 , y24024 , y24025 , y24026 , y24027 , y24028 , y24029 , y24030 , y24031 , y24032 , y24033 , y24034 , y24035 , y24036 , y24037 , y24038 , y24039 , y24040 , y24041 , y24042 , y24043 , y24044 , y24045 , y24046 , y24047 , y24048 , y24049 , y24050 , y24051 , y24052 , y24053 , y24054 , y24055 , y24056 , y24057 , y24058 , y24059 , y24060 , y24061 , y24062 , y24063 , y24064 , y24065 , y24066 , y24067 , y24068 , y24069 , y24070 , y24071 , y24072 , y24073 , y24074 , y24075 , y24076 , y24077 , y24078 , y24079 , y24080 , y24081 , y24082 , y24083 , y24084 , y24085 , y24086 , y24087 , y24088 , y24089 , y24090 , y24091 , y24092 , y24093 , y24094 , y24095 , y24096 , y24097 , y24098 , y24099 , y24100 , y24101 , y24102 , y24103 , y24104 , y24105 , y24106 , y24107 , y24108 , y24109 , y24110 , y24111 , y24112 , y24113 , y24114 , y24115 , y24116 , y24117 , y24118 , y24119 , y24120 , y24121 , y24122 , y24123 , y24124 , y24125 , y24126 , y24127 , y24128 , y24129 , y24130 , y24131 , y24132 , y24133 , y24134 , y24135 , y24136 , y24137 , y24138 , y24139 , y24140 , y24141 , y24142 , y24143 , y24144 , y24145 , y24146 , y24147 , y24148 , y24149 , y24150 , y24151 , y24152 , y24153 , y24154 , y24155 , y24156 , y24157 , y24158 , y24159 , y24160 , y24161 , y24162 , y24163 , y24164 , y24165 , y24166 , y24167 , y24168 , y24169 , y24170 , y24171 , y24172 , y24173 , y24174 , y24175 , y24176 , y24177 , y24178 , y24179 , y24180 , y24181 , y24182 , y24183 , y24184 , y24185 , y24186 , y24187 , y24188 , y24189 , y24190 , y24191 , y24192 , y24193 , y24194 , y24195 , y24196 , y24197 , y24198 , y24199 , y24200 , y24201 , y24202 , y24203 , y24204 , y24205 , y24206 , y24207 , y24208 , y24209 , y24210 , y24211 , y24212 , y24213 , y24214 , y24215 , y24216 , y24217 , y24218 , y24219 , y24220 , y24221 , y24222 , y24223 , y24224 , y24225 , y24226 , y24227 , y24228 , y24229 , y24230 , y24231 , y24232 , y24233 , y24234 , y24235 , y24236 , y24237 , y24238 , y24239 , y24240 , y24241 , y24242 , y24243 , y24244 , y24245 , y24246 , y24247 , y24248 , y24249 , y24250 , y24251 , y24252 , y24253 , y24254 , y24255 , y24256 , y24257 , y24258 , y24259 , y24260 , y24261 , y24262 , y24263 , y24264 , y24265 , y24266 , y24267 , y24268 , y24269 , y24270 , y24271 , y24272 , y24273 , y24274 , y24275 , y24276 , y24277 , y24278 , y24279 , y24280 , y24281 , y24282 , y24283 , y24284 , y24285 , y24286 , y24287 , y24288 , y24289 , y24290 , y24291 , y24292 , y24293 , y24294 , y24295 , y24296 , y24297 , y24298 , y24299 , y24300 , y24301 , y24302 , y24303 , y24304 , y24305 , y24306 , y24307 , y24308 , y24309 , y24310 , y24311 , y24312 , y24313 , y24314 , y24315 , y24316 , y24317 , y24318 , y24319 , y24320 , y24321 , y24322 , y24323 , y24324 , y24325 , y24326 , y24327 , y24328 , y24329 , y24330 , y24331 , y24332 , y24333 , y24334 , y24335 , y24336 , y24337 , y24338 , y24339 , y24340 , y24341 , y24342 , y24343 , y24344 , y24345 , y24346 , y24347 , y24348 , y24349 , y24350 , y24351 , y24352 , y24353 , y24354 , y24355 , y24356 , y24357 , y24358 , y24359 , y24360 , y24361 , y24362 , y24363 , y24364 , y24365 , y24366 , y24367 , y24368 , y24369 , y24370 , y24371 , y24372 , y24373 , y24374 , y24375 , y24376 , y24377 , y24378 , y24379 , y24380 , y24381 , y24382 , y24383 , y24384 , y24385 , y24386 , y24387 , y24388 , y24389 , y24390 , y24391 , y24392 , y24393 , y24394 , y24395 , y24396 , y24397 , y24398 , y24399 , y24400 , y24401 , y24402 , y24403 , y24404 , y24405 , y24406 , y24407 , y24408 , y24409 , y24410 , y24411 , y24412 , y24413 , y24414 , y24415 , y24416 , y24417 , y24418 , y24419 , y24420 , y24421 , y24422 , y24423 , y24424 , y24425 , y24426 , y24427 , y24428 , y24429 , y24430 , y24431 , y24432 , y24433 , y24434 , y24435 , y24436 , y24437 , y24438 , y24439 , y24440 , y24441 , y24442 , y24443 , y24444 , y24445 , y24446 , y24447 , y24448 , y24449 , y24450 , y24451 , y24452 , y24453 , y24454 , y24455 , y24456 , y24457 , y24458 , y24459 , y24460 , y24461 , y24462 , y24463 , y24464 , y24465 , y24466 , y24467 , y24468 , y24469 , y24470 , y24471 , y24472 , y24473 , y24474 , y24475 , y24476 , y24477 , y24478 , y24479 , y24480 , y24481 , y24482 , y24483 , y24484 , y24485 , y24486 , y24487 , y24488 , y24489 , y24490 , y24491 , y24492 , y24493 , y24494 , y24495 , y24496 , y24497 , y24498 , y24499 , y24500 , y24501 , y24502 , y24503 , y24504 , y24505 , y24506 , y24507 , y24508 , y24509 , y24510 , y24511 , y24512 , y24513 , y24514 , y24515 , y24516 , y24517 , y24518 , y24519 , y24520 , y24521 , y24522 , y24523 , y24524 , y24525 , y24526 , y24527 , y24528 , y24529 , y24530 , y24531 , y24532 , y24533 , y24534 , y24535 , y24536 , y24537 , y24538 , y24539 , y24540 , y24541 , y24542 , y24543 , y24544 , y24545 , y24546 , y24547 , y24548 , y24549 , y24550 , y24551 , y24552 , y24553 , y24554 , y24555 , y24556 , y24557 , y24558 , y24559 , y24560 , y24561 , y24562 , y24563 , y24564 , y24565 , y24566 , y24567 , y24568 , y24569 , y24570 , y24571 , y24572 , y24573 , y24574 , y24575 , y24576 , y24577 , y24578 , y24579 , y24580 , y24581 , y24582 , y24583 , y24584 , y24585 , y24586 , y24587 , y24588 , y24589 , y24590 , y24591 , y24592 , y24593 , y24594 , y24595 , y24596 , y24597 , y24598 , y24599 , y24600 , y24601 , y24602 , y24603 , y24604 , y24605 , y24606 , y24607 , y24608 , y24609 , y24610 , y24611 , y24612 , y24613 , y24614 , y24615 , y24616 , y24617 , y24618 , y24619 , y24620 , y24621 , y24622 , y24623 , y24624 , y24625 , y24626 , y24627 , y24628 , y24629 , y24630 , y24631 , y24632 , y24633 , y24634 , y24635 , y24636 , y24637 , y24638 , y24639 , y24640 , y24641 , y24642 , y24643 , y24644 , y24645 , y24646 , y24647 , y24648 , y24649 , y24650 , y24651 , y24652 , y24653 , y24654 , y24655 , y24656 , y24657 , y24658 , y24659 , y24660 , y24661 , y24662 , y24663 , y24664 , y24665 , y24666 , y24667 , y24668 , y24669 , y24670 , y24671 , y24672 , y24673 , y24674 , y24675 , y24676 , y24677 , y24678 , y24679 , y24680 , y24681 , y24682 , y24683 , y24684 , y24685 , y24686 , y24687 , y24688 , y24689 , y24690 , y24691 , y24692 , y24693 , y24694 , y24695 , y24696 , y24697 , y24698 , y24699 , y24700 , y24701 , y24702 , y24703 , y24704 , y24705 , y24706 , y24707 , y24708 , y24709 , y24710 , y24711 , y24712 , y24713 , y24714 , y24715 , y24716 , y24717 , y24718 , y24719 , y24720 , y24721 , y24722 , y24723 , y24724 , y24725 , y24726 , y24727 , y24728 , y24729 , y24730 , y24731 , y24732 , y24733 , y24734 , y24735 , y24736 , y24737 , y24738 , y24739 , y24740 , y24741 , y24742 , y24743 , y24744 , y24745 , y24746 , y24747 , y24748 , y24749 , y24750 , y24751 , y24752 , y24753 , y24754 , y24755 , y24756 , y24757 , y24758 , y24759 , y24760 , y24761 , y24762 , y24763 , y24764 , y24765 , y24766 , y24767 , y24768 , y24769 , y24770 , y24771 , y24772 , y24773 , y24774 , y24775 , y24776 , y24777 , y24778 , y24779 , y24780 , y24781 , y24782 , y24783 , y24784 , y24785 , y24786 , y24787 , y24788 , y24789 , y24790 , y24791 , y24792 , y24793 , y24794 , y24795 , y24796 , y24797 , y24798 , y24799 , y24800 , y24801 , y24802 , y24803 , y24804 , y24805 , y24806 , y24807 , y24808 , y24809 , y24810 , y24811 , y24812 , y24813 , y24814 , y24815 , y24816 , y24817 , y24818 , y24819 , y24820 , y24821 , y24822 , y24823 , y24824 , y24825 , y24826 , y24827 , y24828 , y24829 , y24830 , y24831 , y24832 , y24833 , y24834 , y24835 , y24836 , y24837 , y24838 , y24839 , y24840 , y24841 , y24842 , y24843 , y24844 , y24845 , y24846 , y24847 , y24848 , y24849 , y24850 , y24851 , y24852 , y24853 , y24854 , y24855 , y24856 , y24857 , y24858 , y24859 , y24860 , y24861 , y24862 , y24863 , y24864 , y24865 , y24866 , y24867 , y24868 , y24869 , y24870 , y24871 , y24872 , y24873 , y24874 , y24875 , y24876 , y24877 , y24878 , y24879 , y24880 , y24881 , y24882 , y24883 , y24884 , y24885 , y24886 , y24887 , y24888 , y24889 , y24890 , y24891 , y24892 , y24893 , y24894 , y24895 , y24896 , y24897 , y24898 , y24899 , y24900 , y24901 , y24902 , y24903 , y24904 , y24905 , y24906 , y24907 , y24908 , y24909 , y24910 , y24911 , y24912 , y24913 , y24914 , y24915 , y24916 , y24917 , y24918 , y24919 , y24920 , y24921 , y24922 , y24923 , y24924 , y24925 , y24926 , y24927 , y24928 , y24929 , y24930 , y24931 , y24932 , y24933 , y24934 , y24935 , y24936 , y24937 , y24938 , y24939 , y24940 , y24941 , y24942 , y24943 , y24944 , y24945 , y24946 , y24947 , y24948 , y24949 , y24950 , y24951 , y24952 , y24953 , y24954 , y24955 , y24956 , y24957 , y24958 , y24959 , y24960 , y24961 , y24962 , y24963 , y24964 , y24965 , y24966 , y24967 , y24968 , y24969 , y24970 , y24971 , y24972 , y24973 , y24974 , y24975 , y24976 , y24977 , y24978 , y24979 , y24980 , y24981 , y24982 , y24983 , y24984 , y24985 , y24986 , y24987 , y24988 , y24989 , y24990 , y24991 , y24992 , y24993 , y24994 , y24995 , y24996 , y24997 , y24998 , y24999 , y25000 , y25001 , y25002 , y25003 , y25004 , y25005 , y25006 , y25007 , y25008 , y25009 , y25010 , y25011 , y25012 , y25013 , y25014 , y25015 , y25016 , y25017 , y25018 , y25019 , y25020 , y25021 , y25022 , y25023 , y25024 , y25025 , y25026 , y25027 , y25028 , y25029 , y25030 , y25031 , y25032 , y25033 , y25034 , y25035 , y25036 , y25037 , y25038 , y25039 , y25040 , y25041 , y25042 , y25043 , y25044 , y25045 , y25046 , y25047 , y25048 , y25049 , y25050 , y25051 , y25052 , y25053 , y25054 , y25055 , y25056 , y25057 , y25058 , y25059 , y25060 , y25061 , y25062 , y25063 , y25064 , y25065 , y25066 , y25067 , y25068 , y25069 , y25070 , y25071 , y25072 , y25073 , y25074 , y25075 , y25076 , y25077 , y25078 , y25079 , y25080 , y25081 , y25082 , y25083 , y25084 , y25085 , y25086 , y25087 , y25088 , y25089 , y25090 , y25091 , y25092 , y25093 , y25094 , y25095 , y25096 , y25097 , y25098 , y25099 , y25100 , y25101 , y25102 , y25103 , y25104 , y25105 , y25106 , y25107 , y25108 , y25109 , y25110 , y25111 , y25112 , y25113 , y25114 , y25115 , y25116 , y25117 , y25118 , y25119 , y25120 , y25121 , y25122 , y25123 , y25124 , y25125 , y25126 , y25127 , y25128 , y25129 , y25130 , y25131 , y25132 , y25133 , y25134 , y25135 , y25136 , y25137 , y25138 , y25139 , y25140 , y25141 , y25142 , y25143 , y25144 , y25145 , y25146 , y25147 , y25148 , y25149 , y25150 , y25151 , y25152 , y25153 , y25154 , y25155 , y25156 , y25157 , y25158 , y25159 , y25160 , y25161 , y25162 , y25163 , y25164 , y25165 , y25166 , y25167 , y25168 , y25169 , y25170 , y25171 , y25172 , y25173 , y25174 , y25175 , y25176 , y25177 , y25178 , y25179 , y25180 , y25181 , y25182 , y25183 , y25184 , y25185 , y25186 , y25187 , y25188 , y25189 , y25190 , y25191 , y25192 , y25193 , y25194 , y25195 , y25196 , y25197 , y25198 , y25199 , y25200 , y25201 , y25202 , y25203 , y25204 , y25205 , y25206 , y25207 , y25208 , y25209 , y25210 , y25211 , y25212 , y25213 , y25214 , y25215 , y25216 , y25217 , y25218 , y25219 , y25220 , y25221 , y25222 , y25223 , y25224 , y25225 , y25226 , y25227 , y25228 , y25229 , y25230 , y25231 , y25232 , y25233 , y25234 , y25235 , y25236 , y25237 , y25238 , y25239 , y25240 , y25241 , y25242 , y25243 , y25244 , y25245 , y25246 , y25247 , y25248 , y25249 , y25250 , y25251 , y25252 , y25253 , y25254 , y25255 , y25256 , y25257 , y25258 , y25259 , y25260 , y25261 , y25262 , y25263 , y25264 , y25265 , y25266 , y25267 , y25268 , y25269 , y25270 , y25271 , y25272 , y25273 , y25274 , y25275 , y25276 , y25277 , y25278 , y25279 , y25280 , y25281 , y25282 , y25283 , y25284 , y25285 , y25286 , y25287 , y25288 , y25289 , y25290 , y25291 , y25292 , y25293 , y25294 , y25295 , y25296 , y25297 , y25298 , y25299 , y25300 , y25301 , y25302 , y25303 , y25304 , y25305 , y25306 , y25307 , y25308 , y25309 , y25310 , y25311 , y25312 , y25313 , y25314 , y25315 , y25316 , y25317 , y25318 , y25319 , y25320 , y25321 , y25322 , y25323 , y25324 , y25325 , y25326 , y25327 , y25328 , y25329 , y25330 , y25331 , y25332 , y25333 , y25334 , y25335 , y25336 , y25337 , y25338 , y25339 , y25340 , y25341 , y25342 , y25343 , y25344 , y25345 , y25346 , y25347 , y25348 , y25349 , y25350 , y25351 , y25352 , y25353 , y25354 , y25355 , y25356 , y25357 , y25358 , y25359 , y25360 , y25361 , y25362 , y25363 , y25364 , y25365 , y25366 , y25367 , y25368 , y25369 , y25370 , y25371 , y25372 , y25373 , y25374 , y25375 , y25376 , y25377 , y25378 , y25379 , y25380 , y25381 , y25382 , y25383 , y25384 , y25385 , y25386 , y25387 , y25388 , y25389 , y25390 , y25391 , y25392 , y25393 , y25394 , y25395 , y25396 , y25397 , y25398 , y25399 , y25400 , y25401 , y25402 , y25403 , y25404 , y25405 , y25406 , y25407 , y25408 , y25409 , y25410 , y25411 , y25412 , y25413 , y25414 , y25415 , y25416 , y25417 , y25418 , y25419 , y25420 , y25421 , y25422 , y25423 , y25424 , y25425 , y25426 , y25427 , y25428 , y25429 , y25430 , y25431 , y25432 , y25433 , y25434 , y25435 , y25436 , y25437 , y25438 , y25439 , y25440 , y25441 , y25442 , y25443 , y25444 , y25445 , y25446 , y25447 , y25448 , y25449 , y25450 , y25451 , y25452 , y25453 , y25454 , y25455 , y25456 , y25457 , y25458 , y25459 , y25460 , y25461 , y25462 , y25463 , y25464 , y25465 , y25466 , y25467 , y25468 , y25469 , y25470 , y25471 , y25472 , y25473 , y25474 , y25475 , y25476 , y25477 , y25478 , y25479 , y25480 , y25481 , y25482 , y25483 , y25484 , y25485 , y25486 , y25487 , y25488 , y25489 , y25490 , y25491 , y25492 , y25493 , y25494 , y25495 , y25496 , y25497 , y25498 , y25499 , y25500 , y25501 , y25502 , y25503 , y25504 , y25505 , y25506 , y25507 , y25508 , y25509 , y25510 , y25511 , y25512 , y25513 , y25514 , y25515 , y25516 , y25517 , y25518 , y25519 , y25520 , y25521 , y25522 , y25523 , y25524 , y25525 , y25526 , y25527 , y25528 , y25529 , y25530 , y25531 , y25532 , y25533 , y25534 , y25535 , y25536 , y25537 , y25538 , y25539 , y25540 , y25541 , y25542 , y25543 , y25544 , y25545 , y25546 , y25547 , y25548 , y25549 , y25550 , y25551 , y25552 , y25553 , y25554 , y25555 , y25556 , y25557 , y25558 , y25559 , y25560 , y25561 , y25562 , y25563 , y25564 , y25565 , y25566 , y25567 , y25568 , y25569 , y25570 , y25571 , y25572 , y25573 , y25574 , y25575 , y25576 , y25577 , y25578 , y25579 , y25580 , y25581 , y25582 , y25583 , y25584 , y25585 , y25586 , y25587 , y25588 , y25589 , y25590 , y25591 , y25592 , y25593 , y25594 , y25595 , y25596 , y25597 , y25598 , y25599 , y25600 , y25601 , y25602 , y25603 , y25604 , y25605 , y25606 , y25607 , y25608 , y25609 , y25610 , y25611 , y25612 , y25613 , y25614 , y25615 , y25616 , y25617 , y25618 , y25619 , y25620 , y25621 , y25622 , y25623 , y25624 , y25625 , y25626 , y25627 , y25628 , y25629 , y25630 , y25631 , y25632 , y25633 , y25634 , y25635 , y25636 , y25637 , y25638 , y25639 , y25640 , y25641 , y25642 , y25643 , y25644 , y25645 , y25646 , y25647 , y25648 , y25649 , y25650 , y25651 , y25652 , y25653 , y25654 , y25655 , y25656 , y25657 , y25658 , y25659 , y25660 , y25661 , y25662 , y25663 , y25664 , y25665 , y25666 , y25667 , y25668 , y25669 , y25670 , y25671 , y25672 , y25673 , y25674 , y25675 , y25676 , y25677 , y25678 , y25679 , y25680 , y25681 , y25682 , y25683 , y25684 , y25685 , y25686 , y25687 , y25688 , y25689 , y25690 , y25691 , y25692 , y25693 , y25694 , y25695 , y25696 , y25697 , y25698 , y25699 , y25700 , y25701 , y25702 , y25703 , y25704 , y25705 , y25706 , y25707 , y25708 , y25709 , y25710 , y25711 , y25712 , y25713 , y25714 , y25715 , y25716 , y25717 , y25718 , y25719 , y25720 , y25721 , y25722 , y25723 , y25724 , y25725 , y25726 , y25727 , y25728 , y25729 , y25730 , y25731 , y25732 , y25733 , y25734 , y25735 , y25736 , y25737 , y25738 , y25739 , y25740 , y25741 , y25742 , y25743 , y25744 , y25745 , y25746 , y25747 , y25748 , y25749 , y25750 , y25751 , y25752 , y25753 , y25754 , y25755 , y25756 , y25757 , y25758 , y25759 , y25760 , y25761 , y25762 , y25763 , y25764 , y25765 , y25766 , y25767 , y25768 , y25769 , y25770 , y25771 , y25772 , y25773 , y25774 , y25775 , y25776 , y25777 , y25778 , y25779 , y25780 , y25781 , y25782 , y25783 , y25784 , y25785 , y25786 , y25787 , y25788 , y25789 , y25790 , y25791 , y25792 , y25793 , y25794 , y25795 , y25796 , y25797 , y25798 , y25799 , y25800 , y25801 , y25802 , y25803 , y25804 , y25805 , y25806 , y25807 , y25808 , y25809 , y25810 , y25811 , y25812 , y25813 , y25814 , y25815 , y25816 , y25817 , y25818 , y25819 , y25820 , y25821 , y25822 , y25823 , y25824 , y25825 , y25826 , y25827 , y25828 , y25829 , y25830 , y25831 , y25832 , y25833 , y25834 , y25835 , y25836 , y25837 , y25838 , y25839 , y25840 , y25841 , y25842 , y25843 , y25844 , y25845 , y25846 , y25847 , y25848 , y25849 , y25850 , y25851 , y25852 , y25853 , y25854 , y25855 , y25856 , y25857 , y25858 , y25859 , y25860 , y25861 , y25862 , y25863 , y25864 , y25865 , y25866 , y25867 , y25868 , y25869 , y25870 , y25871 , y25872 , y25873 , y25874 , y25875 , y25876 , y25877 , y25878 , y25879 , y25880 , y25881 , y25882 , y25883 , y25884 , y25885 , y25886 , y25887 , y25888 , y25889 , y25890 , y25891 , y25892 , y25893 , y25894 , y25895 , y25896 , y25897 , y25898 , y25899 , y25900 , y25901 , y25902 , y25903 , y25904 , y25905 , y25906 , y25907 , y25908 , y25909 , y25910 , y25911 , y25912 , y25913 , y25914 , y25915 , y25916 , y25917 , y25918 , y25919 , y25920 , y25921 , y25922 , y25923 , y25924 , y25925 , y25926 , y25927 , y25928 , y25929 , y25930 , y25931 , y25932 , y25933 , y25934 , y25935 , y25936 , y25937 , y25938 , y25939 , y25940 , y25941 , y25942 , y25943 , y25944 , y25945 , y25946 , y25947 , y25948 , y25949 , y25950 , y25951 , y25952 , y25953 , y25954 , y25955 , y25956 , y25957 , y25958 , y25959 , y25960 , y25961 , y25962 , y25963 , y25964 , y25965 , y25966 , y25967 , y25968 , y25969 , y25970 , y25971 , y25972 , y25973 , y25974 , y25975 , y25976 , y25977 , y25978 , y25979 , y25980 , y25981 , y25982 , y25983 , y25984 , y25985 , y25986 , y25987 , y25988 , y25989 , y25990 , y25991 , y25992 , y25993 , y25994 , y25995 , y25996 , y25997 , y25998 , y25999 , y26000 , y26001 , y26002 , y26003 , y26004 , y26005 , y26006 , y26007 , y26008 , y26009 , y26010 , y26011 , y26012 , y26013 , y26014 , y26015 , y26016 , y26017 , y26018 , y26019 , y26020 , y26021 , y26022 , y26023 , y26024 , y26025 , y26026 , y26027 , y26028 , y26029 , y26030 , y26031 , y26032 , y26033 , y26034 , y26035 , y26036 , y26037 , y26038 , y26039 , y26040 , y26041 , y26042 , y26043 , y26044 , y26045 , y26046 , y26047 , y26048 , y26049 , y26050 , y26051 , y26052 , y26053 , y26054 , y26055 , y26056 , y26057 , y26058 , y26059 , y26060 , y26061 , y26062 , y26063 , y26064 , y26065 , y26066 , y26067 , y26068 , y26069 , y26070 , y26071 , y26072 , y26073 , y26074 , y26075 , y26076 , y26077 , y26078 , y26079 , y26080 , y26081 , y26082 , y26083 , y26084 , y26085 , y26086 , y26087 , y26088 , y26089 , y26090 , y26091 , y26092 , y26093 , y26094 , y26095 , y26096 , y26097 , y26098 , y26099 , y26100 , y26101 , y26102 , y26103 , y26104 , y26105 , y26106 , y26107 , y26108 , y26109 , y26110 , y26111 , y26112 , y26113 , y26114 , y26115 , y26116 , y26117 , y26118 , y26119 , y26120 , y26121 , y26122 , y26123 , y26124 , y26125 , y26126 , y26127 , y26128 , y26129 , y26130 , y26131 , y26132 , y26133 , y26134 , y26135 , y26136 , y26137 , y26138 , y26139 , y26140 , y26141 , y26142 , y26143 , y26144 , y26145 , y26146 , y26147 , y26148 , y26149 , y26150 , y26151 , y26152 , y26153 , y26154 , y26155 , y26156 , y26157 , y26158 , y26159 , y26160 , y26161 , y26162 , y26163 , y26164 , y26165 , y26166 , y26167 , y26168 , y26169 , y26170 , y26171 , y26172 , y26173 , y26174 , y26175 , y26176 , y26177 , y26178 , y26179 , y26180 , y26181 , y26182 , y26183 , y26184 , y26185 , y26186 , y26187 , y26188 , y26189 , y26190 , y26191 , y26192 , y26193 , y26194 , y26195 , y26196 , y26197 , y26198 , y26199 , y26200 , y26201 , y26202 , y26203 , y26204 , y26205 , y26206 , y26207 , y26208 , y26209 , y26210 , y26211 , y26212 , y26213 , y26214 , y26215 , y26216 , y26217 , y26218 , y26219 , y26220 , y26221 , y26222 , y26223 , y26224 , y26225 , y26226 , y26227 , y26228 , y26229 , y26230 , y26231 , y26232 , y26233 , y26234 , y26235 , y26236 , y26237 , y26238 , y26239 , y26240 , y26241 , y26242 , y26243 , y26244 , y26245 , y26246 , y26247 , y26248 , y26249 , y26250 , y26251 , y26252 , y26253 , y26254 , y26255 , y26256 , y26257 , y26258 , y26259 , y26260 , y26261 , y26262 , y26263 , y26264 , y26265 , y26266 , y26267 , y26268 , y26269 , y26270 , y26271 , y26272 , y26273 , y26274 , y26275 , y26276 , y26277 , y26278 , y26279 , y26280 , y26281 , y26282 , y26283 , y26284 , y26285 , y26286 , y26287 , y26288 , y26289 , y26290 , y26291 , y26292 , y26293 , y26294 , y26295 , y26296 , y26297 , y26298 , y26299 , y26300 , y26301 , y26302 , y26303 , y26304 , y26305 , y26306 , y26307 , y26308 , y26309 , y26310 , y26311 , y26312 , y26313 , y26314 , y26315 , y26316 , y26317 , y26318 , y26319 , y26320 , y26321 , y26322 , y26323 , y26324 , y26325 , y26326 , y26327 , y26328 , y26329 , y26330 , y26331 , y26332 , y26333 , y26334 , y26335 , y26336 , y26337 , y26338 , y26339 , y26340 , y26341 , y26342 , y26343 , y26344 , y26345 , y26346 , y26347 , y26348 , y26349 , y26350 , y26351 , y26352 , y26353 , y26354 , y26355 , y26356 , y26357 , y26358 , y26359 , y26360 , y26361 , y26362 , y26363 , y26364 , y26365 , y26366 , y26367 , y26368 , y26369 , y26370 , y26371 , y26372 , y26373 , y26374 , y26375 , y26376 , y26377 , y26378 , y26379 , y26380 , y26381 , y26382 , y26383 , y26384 , y26385 , y26386 , y26387 , y26388 , y26389 , y26390 , y26391 , y26392 , y26393 , y26394 , y26395 , y26396 , y26397 , y26398 , y26399 , y26400 , y26401 , y26402 , y26403 , y26404 , y26405 , y26406 , y26407 , y26408 , y26409 , y26410 , y26411 , y26412 , y26413 , y26414 , y26415 , y26416 , y26417 , y26418 , y26419 , y26420 , y26421 , y26422 , y26423 , y26424 , y26425 , y26426 , y26427 , y26428 , y26429 , y26430 , y26431 , y26432 , y26433 , y26434 , y26435 , y26436 , y26437 , y26438 , y26439 , y26440 , y26441 , y26442 , y26443 , y26444 , y26445 , y26446 , y26447 , y26448 , y26449 , y26450 , y26451 , y26452 , y26453 , y26454 , y26455 , y26456 , y26457 , y26458 , y26459 , y26460 , y26461 , y26462 , y26463 , y26464 , y26465 , y26466 , y26467 , y26468 , y26469 , y26470 , y26471 , y26472 , y26473 , y26474 , y26475 , y26476 , y26477 , y26478 , y26479 , y26480 , y26481 , y26482 , y26483 , y26484 , y26485 , y26486 , y26487 , y26488 , y26489 , y26490 , y26491 , y26492 , y26493 , y26494 , y26495 , y26496 , y26497 , y26498 , y26499 , y26500 , y26501 , y26502 , y26503 , y26504 , y26505 , y26506 , y26507 , y26508 , y26509 , y26510 , y26511 , y26512 , y26513 , y26514 , y26515 , y26516 , y26517 , y26518 , y26519 , y26520 , y26521 , y26522 , y26523 , y26524 , y26525 , y26526 , y26527 , y26528 , y26529 , y26530 , y26531 , y26532 , y26533 , y26534 , y26535 , y26536 , y26537 , y26538 , y26539 , y26540 , y26541 , y26542 , y26543 , y26544 , y26545 , y26546 , y26547 , y26548 , y26549 , y26550 , y26551 , y26552 , y26553 , y26554 , y26555 , y26556 , y26557 , y26558 , y26559 , y26560 , y26561 , y26562 , y26563 , y26564 , y26565 , y26566 , y26567 , y26568 , y26569 , y26570 , y26571 , y26572 , y26573 , y26574 , y26575 , y26576 , y26577 , y26578 , y26579 , y26580 , y26581 , y26582 , y26583 , y26584 , y26585 , y26586 , y26587 , y26588 , y26589 , y26590 , y26591 , y26592 , y26593 , y26594 , y26595 , y26596 , y26597 , y26598 , y26599 , y26600 , y26601 , y26602 , y26603 , y26604 , y26605 , y26606 , y26607 , y26608 , y26609 , y26610 , y26611 , y26612 , y26613 , y26614 , y26615 , y26616 , y26617 , y26618 , y26619 , y26620 , y26621 , y26622 , y26623 , y26624 , y26625 , y26626 , y26627 , y26628 , y26629 , y26630 , y26631 , y26632 , y26633 , y26634 , y26635 , y26636 , y26637 , y26638 , y26639 , y26640 , y26641 , y26642 , y26643 , y26644 , y26645 , y26646 , y26647 , y26648 , y26649 , y26650 , y26651 , y26652 , y26653 , y26654 , y26655 , y26656 , y26657 , y26658 , y26659 , y26660 , y26661 , y26662 , y26663 , y26664 , y26665 , y26666 , y26667 , y26668 , y26669 , y26670 , y26671 , y26672 , y26673 , y26674 , y26675 , y26676 , y26677 , y26678 , y26679 , y26680 , y26681 , y26682 , y26683 , y26684 , y26685 , y26686 , y26687 , y26688 , y26689 , y26690 , y26691 , y26692 , y26693 , y26694 , y26695 , y26696 , y26697 , y26698 , y26699 , y26700 , y26701 , y26702 , y26703 , y26704 , y26705 , y26706 , y26707 , y26708 , y26709 , y26710 , y26711 , y26712 , y26713 , y26714 , y26715 , y26716 , y26717 , y26718 , y26719 , y26720 , y26721 , y26722 , y26723 , y26724 , y26725 , y26726 , y26727 , y26728 , y26729 , y26730 , y26731 , y26732 , y26733 , y26734 , y26735 , y26736 , y26737 , y26738 , y26739 , y26740 , y26741 , y26742 , y26743 , y26744 , y26745 , y26746 , y26747 , y26748 , y26749 , y26750 , y26751 , y26752 , y26753 , y26754 , y26755 , y26756 , y26757 , y26758 , y26759 , y26760 , y26761 , y26762 , y26763 , y26764 , y26765 , y26766 , y26767 , y26768 , y26769 , y26770 , y26771 , y26772 , y26773 , y26774 , y26775 , y26776 , y26777 , y26778 , y26779 , y26780 , y26781 , y26782 , y26783 , y26784 , y26785 , y26786 , y26787 , y26788 , y26789 , y26790 , y26791 , y26792 , y26793 , y26794 , y26795 , y26796 , y26797 , y26798 , y26799 , y26800 , y26801 , y26802 , y26803 , y26804 , y26805 , y26806 , y26807 , y26808 , y26809 , y26810 , y26811 , y26812 , y26813 , y26814 , y26815 , y26816 , y26817 , y26818 , y26819 , y26820 , y26821 , y26822 , y26823 , y26824 , y26825 , y26826 , y26827 , y26828 , y26829 , y26830 , y26831 , y26832 , y26833 , y26834 , y26835 , y26836 , y26837 , y26838 , y26839 , y26840 , y26841 , y26842 , y26843 , y26844 , y26845 , y26846 , y26847 , y26848 , y26849 , y26850 , y26851 , y26852 , y26853 , y26854 , y26855 , y26856 , y26857 , y26858 , y26859 , y26860 , y26861 , y26862 , y26863 , y26864 , y26865 , y26866 , y26867 , y26868 , y26869 , y26870 , y26871 , y26872 , y26873 , y26874 , y26875 , y26876 , y26877 , y26878 , y26879 , y26880 , y26881 , y26882 , y26883 , y26884 , y26885 , y26886 , y26887 , y26888 , y26889 , y26890 , y26891 , y26892 , y26893 , y26894 , y26895 , y26896 , y26897 , y26898 , y26899 , y26900 , y26901 , y26902 , y26903 , y26904 , y26905 , y26906 , y26907 , y26908 , y26909 , y26910 , y26911 , y26912 , y26913 , y26914 , y26915 , y26916 , y26917 , y26918 , y26919 , y26920 , y26921 , y26922 , y26923 , y26924 , y26925 , y26926 , y26927 , y26928 , y26929 , y26930 , y26931 , y26932 , y26933 , y26934 , y26935 , y26936 , y26937 , y26938 , y26939 , y26940 , y26941 , y26942 , y26943 , y26944 , y26945 , y26946 , y26947 , y26948 , y26949 , y26950 , y26951 , y26952 , y26953 , y26954 , y26955 , y26956 , y26957 , y26958 , y26959 , y26960 , y26961 , y26962 , y26963 , y26964 , y26965 , y26966 , y26967 , y26968 , y26969 , y26970 , y26971 , y26972 , y26973 , y26974 , y26975 , y26976 , y26977 , y26978 , y26979 , y26980 , y26981 , y26982 , y26983 , y26984 , y26985 , y26986 , y26987 , y26988 , y26989 , y26990 , y26991 , y26992 , y26993 , y26994 , y26995 , y26996 , y26997 , y26998 , y26999 , y27000 , y27001 , y27002 , y27003 , y27004 , y27005 , y27006 , y27007 , y27008 , y27009 , y27010 , y27011 , y27012 , y27013 , y27014 , y27015 , y27016 , y27017 , y27018 , y27019 , y27020 , y27021 , y27022 , y27023 , y27024 , y27025 , y27026 , y27027 , y27028 , y27029 , y27030 , y27031 , y27032 , y27033 , y27034 , y27035 , y27036 , y27037 , y27038 , y27039 , y27040 , y27041 , y27042 , y27043 , y27044 , y27045 , y27046 , y27047 , y27048 , y27049 , y27050 , y27051 , y27052 , y27053 , y27054 , y27055 , y27056 , y27057 , y27058 , y27059 , y27060 , y27061 , y27062 , y27063 , y27064 , y27065 , y27066 , y27067 , y27068 , y27069 , y27070 , y27071 , y27072 , y27073 , y27074 , y27075 , y27076 , y27077 , y27078 , y27079 , y27080 , y27081 , y27082 , y27083 , y27084 , y27085 , y27086 , y27087 , y27088 , y27089 , y27090 , y27091 , y27092 , y27093 , y27094 , y27095 , y27096 , y27097 , y27098 , y27099 , y27100 , y27101 , y27102 , y27103 , y27104 , y27105 , y27106 , y27107 , y27108 , y27109 , y27110 , y27111 , y27112 , y27113 , y27114 , y27115 , y27116 , y27117 , y27118 , y27119 , y27120 , y27121 , y27122 , y27123 , y27124 , y27125 , y27126 , y27127 , y27128 , y27129 , y27130 , y27131 , y27132 , y27133 , y27134 , y27135 , y27136 , y27137 , y27138 , y27139 , y27140 , y27141 , y27142 , y27143 , y27144 , y27145 , y27146 , y27147 , y27148 , y27149 , y27150 , y27151 , y27152 , y27153 , y27154 , y27155 , y27156 , y27157 , y27158 , y27159 , y27160 , y27161 , y27162 , y27163 , y27164 , y27165 , y27166 , y27167 , y27168 , y27169 , y27170 , y27171 , y27172 , y27173 , y27174 , y27175 , y27176 , y27177 , y27178 , y27179 , y27180 , y27181 , y27182 , y27183 , y27184 , y27185 , y27186 , y27187 , y27188 , y27189 , y27190 , y27191 , y27192 , y27193 , y27194 , y27195 , y27196 , y27197 , y27198 , y27199 , y27200 , y27201 , y27202 , y27203 , y27204 , y27205 , y27206 , y27207 , y27208 , y27209 , y27210 , y27211 , y27212 , y27213 , y27214 , y27215 , y27216 , y27217 , y27218 , y27219 , y27220 , y27221 , y27222 , y27223 , y27224 , y27225 , y27226 , y27227 , y27228 , y27229 , y27230 , y27231 , y27232 , y27233 , y27234 , y27235 , y27236 , y27237 , y27238 , y27239 , y27240 , y27241 , y27242 , y27243 , y27244 , y27245 , y27246 , y27247 , y27248 , y27249 , y27250 , y27251 , y27252 , y27253 , y27254 , y27255 , y27256 , y27257 , y27258 , y27259 , y27260 , y27261 , y27262 , y27263 , y27264 , y27265 , y27266 , y27267 , y27268 , y27269 , y27270 , y27271 , y27272 , y27273 , y27274 , y27275 , y27276 , y27277 , y27278 , y27279 , y27280 , y27281 , y27282 , y27283 , y27284 , y27285 , y27286 , y27287 , y27288 , y27289 , y27290 , y27291 , y27292 , y27293 , y27294 , y27295 , y27296 , y27297 , y27298 , y27299 , y27300 , y27301 , y27302 , y27303 , y27304 , y27305 , y27306 , y27307 , y27308 , y27309 , y27310 , y27311 , y27312 , y27313 , y27314 , y27315 , y27316 , y27317 , y27318 , y27319 , y27320 , y27321 , y27322 , y27323 , y27324 , y27325 , y27326 , y27327 , y27328 , y27329 , y27330 , y27331 , y27332 , y27333 , y27334 , y27335 , y27336 , y27337 , y27338 , y27339 , y27340 , y27341 , y27342 , y27343 , y27344 , y27345 , y27346 , y27347 , y27348 , y27349 , y27350 , y27351 , y27352 , y27353 , y27354 , y27355 , y27356 , y27357 , y27358 , y27359 , y27360 , y27361 , y27362 , y27363 , y27364 , y27365 , y27366 , y27367 , y27368 , y27369 , y27370 , y27371 , y27372 , y27373 , y27374 , y27375 , y27376 , y27377 , y27378 , y27379 , y27380 , y27381 , y27382 , y27383 , y27384 , y27385 , y27386 , y27387 , y27388 , y27389 , y27390 , y27391 , y27392 , y27393 , y27394 , y27395 , y27396 , y27397 , y27398 , y27399 , y27400 , y27401 , y27402 , y27403 , y27404 , y27405 , y27406 , y27407 , y27408 , y27409 , y27410 , y27411 , y27412 , y27413 , y27414 , y27415 , y27416 , y27417 , y27418 , y27419 , y27420 , y27421 , y27422 , y27423 , y27424 , y27425 , y27426 , y27427 , y27428 , y27429 , y27430 , y27431 , y27432 , y27433 , y27434 , y27435 , y27436 , y27437 , y27438 , y27439 , y27440 , y27441 , y27442 , y27443 , y27444 , y27445 , y27446 , y27447 , y27448 , y27449 , y27450 , y27451 , y27452 , y27453 , y27454 , y27455 , y27456 , y27457 , y27458 , y27459 , y27460 , y27461 , y27462 , y27463 , y27464 , y27465 , y27466 , y27467 , y27468 , y27469 , y27470 , y27471 , y27472 , y27473 , y27474 , y27475 , y27476 , y27477 , y27478 , y27479 , y27480 , y27481 , y27482 , y27483 , y27484 , y27485 , y27486 , y27487 , y27488 , y27489 , y27490 , y27491 , y27492 , y27493 , y27494 , y27495 , y27496 , y27497 , y27498 , y27499 , y27500 , y27501 , y27502 , y27503 , y27504 , y27505 , y27506 , y27507 , y27508 , y27509 , y27510 , y27511 , y27512 , y27513 , y27514 , y27515 , y27516 , y27517 , y27518 , y27519 , y27520 , y27521 , y27522 , y27523 , y27524 , y27525 , y27526 , y27527 , y27528 , y27529 , y27530 , y27531 , y27532 , y27533 , y27534 , y27535 , y27536 , y27537 , y27538 , y27539 , y27540 , y27541 , y27542 , y27543 , y27544 , y27545 , y27546 , y27547 , y27548 , y27549 , y27550 , y27551 , y27552 , y27553 , y27554 , y27555 , y27556 , y27557 , y27558 , y27559 , y27560 , y27561 , y27562 , y27563 , y27564 , y27565 , y27566 , y27567 , y27568 , y27569 , y27570 , y27571 , y27572 , y27573 , y27574 , y27575 , y27576 , y27577 , y27578 , y27579 , y27580 , y27581 , y27582 , y27583 , y27584 , y27585 , y27586 , y27587 , y27588 , y27589 , y27590 , y27591 , y27592 , y27593 , y27594 , y27595 , y27596 , y27597 , y27598 , y27599 , y27600 , y27601 , y27602 , y27603 , y27604 , y27605 , y27606 , y27607 , y27608 , y27609 , y27610 , y27611 , y27612 , y27613 , y27614 , y27615 , y27616 , y27617 , y27618 , y27619 , y27620 , y27621 , y27622 , y27623 , y27624 , y27625 , y27626 , y27627 , y27628 , y27629 , y27630 , y27631 , y27632 , y27633 , y27634 , y27635 , y27636 , y27637 , y27638 , y27639 , y27640 , y27641 , y27642 , y27643 , y27644 , y27645 , y27646 , y27647 , y27648 , y27649 , y27650 , y27651 , y27652 , y27653 , y27654 , y27655 , y27656 , y27657 , y27658 , y27659 , y27660 , y27661 , y27662 , y27663 , y27664 , y27665 , y27666 , y27667 , y27668 , y27669 , y27670 , y27671 , y27672 , y27673 , y27674 , y27675 , y27676 , y27677 , y27678 , y27679 , y27680 , y27681 , y27682 , y27683 , y27684 , y27685 , y27686 , y27687 , y27688 , y27689 , y27690 , y27691 , y27692 , y27693 , y27694 , y27695 , y27696 , y27697 , y27698 , y27699 , y27700 , y27701 , y27702 , y27703 , y27704 , y27705 , y27706 , y27707 , y27708 , y27709 , y27710 , y27711 , y27712 , y27713 , y27714 , y27715 , y27716 , y27717 , y27718 , y27719 , y27720 , y27721 , y27722 , y27723 , y27724 , y27725 , y27726 , y27727 , y27728 , y27729 , y27730 , y27731 , y27732 , y27733 , y27734 , y27735 , y27736 , y27737 , y27738 , y27739 , y27740 , y27741 , y27742 , y27743 , y27744 , y27745 , y27746 , y27747 , y27748 , y27749 , y27750 , y27751 , y27752 , y27753 , y27754 , y27755 , y27756 , y27757 , y27758 , y27759 , y27760 , y27761 , y27762 , y27763 , y27764 , y27765 , y27766 , y27767 , y27768 , y27769 , y27770 , y27771 , y27772 , y27773 , y27774 , y27775 , y27776 , y27777 , y27778 , y27779 , y27780 , y27781 , y27782 , y27783 , y27784 , y27785 , y27786 , y27787 , y27788 , y27789 , y27790 , y27791 , y27792 , y27793 , y27794 , y27795 , y27796 , y27797 , y27798 , y27799 , y27800 , y27801 , y27802 , y27803 , y27804 , y27805 , y27806 , y27807 , y27808 , y27809 , y27810 , y27811 , y27812 , y27813 , y27814 , y27815 , y27816 , y27817 , y27818 , y27819 , y27820 , y27821 , y27822 , y27823 , y27824 , y27825 , y27826 , y27827 , y27828 , y27829 , y27830 , y27831 , y27832 , y27833 , y27834 , y27835 , y27836 , y27837 , y27838 , y27839 , y27840 , y27841 , y27842 , y27843 , y27844 , y27845 , y27846 , y27847 , y27848 , y27849 , y27850 , y27851 , y27852 , y27853 , y27854 , y27855 , y27856 , y27857 , y27858 , y27859 , y27860 , y27861 , y27862 , y27863 , y27864 , y27865 , y27866 , y27867 , y27868 , y27869 , y27870 , y27871 , y27872 , y27873 , y27874 , y27875 , y27876 , y27877 , y27878 , y27879 , y27880 , y27881 , y27882 , y27883 , y27884 , y27885 , y27886 , y27887 , y27888 , y27889 , y27890 , y27891 , y27892 , y27893 , y27894 , y27895 , y27896 , y27897 , y27898 , y27899 , y27900 , y27901 , y27902 , y27903 , y27904 , y27905 , y27906 , y27907 , y27908 , y27909 , y27910 , y27911 , y27912 , y27913 , y27914 , y27915 , y27916 , y27917 , y27918 , y27919 , y27920 , y27921 , y27922 , y27923 , y27924 , y27925 , y27926 , y27927 , y27928 , y27929 , y27930 , y27931 , y27932 , y27933 , y27934 , y27935 , y27936 , y27937 , y27938 , y27939 , y27940 , y27941 , y27942 , y27943 , y27944 , y27945 , y27946 , y27947 , y27948 , y27949 , y27950 , y27951 , y27952 , y27953 , y27954 , y27955 , y27956 , y27957 , y27958 , y27959 , y27960 , y27961 , y27962 , y27963 , y27964 , y27965 , y27966 , y27967 , y27968 , y27969 , y27970 , y27971 , y27972 , y27973 , y27974 , y27975 , y27976 , y27977 , y27978 , y27979 , y27980 , y27981 , y27982 , y27983 , y27984 , y27985 , y27986 , y27987 , y27988 , y27989 , y27990 , y27991 , y27992 , y27993 , y27994 , y27995 , y27996 , y27997 , y27998 , y27999 , y28000 , y28001 , y28002 , y28003 , y28004 , y28005 , y28006 , y28007 , y28008 , y28009 , y28010 , y28011 , y28012 , y28013 , y28014 , y28015 , y28016 , y28017 , y28018 , y28019 , y28020 , y28021 , y28022 , y28023 , y28024 , y28025 , y28026 , y28027 , y28028 , y28029 , y28030 , y28031 , y28032 , y28033 , y28034 , y28035 , y28036 , y28037 , y28038 , y28039 , y28040 , y28041 , y28042 , y28043 , y28044 , y28045 , y28046 , y28047 , y28048 , y28049 , y28050 , y28051 , y28052 , y28053 , y28054 , y28055 , y28056 , y28057 , y28058 , y28059 , y28060 , y28061 , y28062 , y28063 , y28064 , y28065 , y28066 , y28067 , y28068 , y28069 , y28070 , y28071 , y28072 , y28073 , y28074 , y28075 , y28076 , y28077 , y28078 , y28079 , y28080 , y28081 , y28082 , y28083 , y28084 , y28085 , y28086 , y28087 , y28088 , y28089 , y28090 , y28091 , y28092 , y28093 , y28094 , y28095 , y28096 , y28097 , y28098 , y28099 , y28100 , y28101 , y28102 , y28103 , y28104 , y28105 , y28106 , y28107 , y28108 , y28109 , y28110 , y28111 , y28112 , y28113 , y28114 , y28115 , y28116 , y28117 , y28118 , y28119 , y28120 , y28121 , y28122 , y28123 , y28124 , y28125 , y28126 , y28127 , y28128 , y28129 , y28130 , y28131 , y28132 , y28133 , y28134 , y28135 , y28136 , y28137 , y28138 , y28139 , y28140 , y28141 , y28142 , y28143 , y28144 , y28145 , y28146 , y28147 , y28148 , y28149 , y28150 , y28151 , y28152 , y28153 , y28154 , y28155 , y28156 , y28157 , y28158 , y28159 , y28160 , y28161 , y28162 , y28163 , y28164 , y28165 , y28166 , y28167 , y28168 , y28169 , y28170 , y28171 , y28172 , y28173 , y28174 , y28175 , y28176 , y28177 , y28178 , y28179 , y28180 , y28181 , y28182 , y28183 , y28184 , y28185 , y28186 , y28187 , y28188 , y28189 , y28190 , y28191 , y28192 , y28193 , y28194 , y28195 , y28196 , y28197 , y28198 , y28199 , y28200 , y28201 , y28202 , y28203 , y28204 , y28205 , y28206 , y28207 , y28208 , y28209 , y28210 , y28211 , y28212 , y28213 , y28214 , y28215 , y28216 , y28217 , y28218 , y28219 , y28220 , y28221 , y28222 , y28223 , y28224 , y28225 , y28226 , y28227 , y28228 , y28229 , y28230 , y28231 , y28232 , y28233 , y28234 , y28235 , y28236 , y28237 , y28238 , y28239 , y28240 , y28241 , y28242 , y28243 , y28244 , y28245 , y28246 , y28247 , y28248 , y28249 , y28250 , y28251 , y28252 , y28253 , y28254 , y28255 , y28256 , y28257 , y28258 , y28259 , y28260 , y28261 , y28262 , y28263 , y28264 , y28265 , y28266 , y28267 , y28268 , y28269 , y28270 , y28271 , y28272 , y28273 , y28274 , y28275 , y28276 , y28277 , y28278 , y28279 , y28280 , y28281 , y28282 , y28283 , y28284 , y28285 , y28286 , y28287 , y28288 , y28289 , y28290 , y28291 , y28292 , y28293 , y28294 , y28295 , y28296 , y28297 , y28298 , y28299 , y28300 , y28301 , y28302 , y28303 , y28304 , y28305 , y28306 , y28307 , y28308 , y28309 , y28310 , y28311 , y28312 , y28313 , y28314 , y28315 , y28316 , y28317 , y28318 , y28319 , y28320 , y28321 , y28322 , y28323 , y28324 , y28325 , y28326 , y28327 , y28328 , y28329 , y28330 , y28331 , y28332 , y28333 , y28334 , y28335 , y28336 , y28337 , y28338 , y28339 , y28340 , y28341 , y28342 , y28343 , y28344 , y28345 , y28346 , y28347 , y28348 , y28349 , y28350 , y28351 , y28352 , y28353 , y28354 , y28355 , y28356 , y28357 , y28358 , y28359 , y28360 , y28361 , y28362 , y28363 , y28364 , y28365 , y28366 , y28367 , y28368 , y28369 , y28370 , y28371 , y28372 , y28373 , y28374 , y28375 , y28376 , y28377 , y28378 , y28379 , y28380 , y28381 , y28382 , y28383 , y28384 , y28385 , y28386 , y28387 , y28388 , y28389 , y28390 , y28391 , y28392 , y28393 , y28394 , y28395 , y28396 , y28397 , y28398 , y28399 , y28400 , y28401 , y28402 , y28403 , y28404 , y28405 , y28406 , y28407 , y28408 , y28409 , y28410 , y28411 , y28412 , y28413 , y28414 , y28415 , y28416 , y28417 , y28418 , y28419 , y28420 , y28421 , y28422 , y28423 , y28424 , y28425 , y28426 , y28427 , y28428 , y28429 , y28430 , y28431 , y28432 , y28433 , y28434 , y28435 , y28436 , y28437 , y28438 , y28439 , y28440 , y28441 , y28442 , y28443 , y28444 , y28445 , y28446 , y28447 , y28448 , y28449 , y28450 , y28451 , y28452 , y28453 , y28454 , y28455 , y28456 , y28457 , y28458 , y28459 , y28460 , y28461 , y28462 , y28463 , y28464 , y28465 , y28466 , y28467 , y28468 , y28469 , y28470 , y28471 , y28472 , y28473 , y28474 , y28475 , y28476 , y28477 , y28478 , y28479 , y28480 , y28481 , y28482 , y28483 , y28484 , y28485 , y28486 , y28487 , y28488 , y28489 , y28490 , y28491 , y28492 , y28493 , y28494 , y28495 , y28496 , y28497 , y28498 , y28499 , y28500 , y28501 , y28502 , y28503 , y28504 , y28505 , y28506 , y28507 , y28508 , y28509 , y28510 , y28511 , y28512 , y28513 , y28514 , y28515 , y28516 , y28517 , y28518 , y28519 , y28520 , y28521 , y28522 , y28523 , y28524 , y28525 , y28526 , y28527 , y28528 , y28529 , y28530 , y28531 , y28532 , y28533 , y28534 , y28535 , y28536 , y28537 , y28538 , y28539 , y28540 , y28541 , y28542 , y28543 , y28544 , y28545 , y28546 , y28547 , y28548 , y28549 , y28550 , y28551 , y28552 , y28553 , y28554 , y28555 , y28556 , y28557 , y28558 , y28559 , y28560 , y28561 , y28562 , y28563 , y28564 , y28565 , y28566 , y28567 , y28568 , y28569 , y28570 , y28571 , y28572 , y28573 , y28574 , y28575 , y28576 , y28577 , y28578 , y28579 , y28580 , y28581 , y28582 , y28583 , y28584 , y28585 , y28586 , y28587 , y28588 , y28589 , y28590 , y28591 , y28592 , y28593 , y28594 , y28595 , y28596 , y28597 , y28598 , y28599 , y28600 , y28601 , y28602 , y28603 , y28604 , y28605 , y28606 , y28607 , y28608 , y28609 , y28610 , y28611 , y28612 , y28613 , y28614 , y28615 , y28616 , y28617 , y28618 , y28619 , y28620 , y28621 , y28622 , y28623 , y28624 , y28625 , y28626 , y28627 , y28628 , y28629 , y28630 , y28631 , y28632 , y28633 , y28634 , y28635 , y28636 , y28637 , y28638 , y28639 , y28640 , y28641 , y28642 , y28643 , y28644 , y28645 , y28646 , y28647 , y28648 , y28649 , y28650 , y28651 , y28652 , y28653 , y28654 , y28655 , y28656 , y28657 , y28658 , y28659 , y28660 , y28661 , y28662 , y28663 , y28664 , y28665 , y28666 , y28667 , y28668 , y28669 , y28670 , y28671 , y28672 , y28673 , y28674 , y28675 , y28676 , y28677 , y28678 , y28679 , y28680 , y28681 , y28682 , y28683 , y28684 , y28685 , y28686 , y28687 , y28688 , y28689 , y28690 , y28691 , y28692 , y28693 , y28694 , y28695 , y28696 , y28697 , y28698 , y28699 , y28700 , y28701 , y28702 , y28703 , y28704 , y28705 , y28706 , y28707 , y28708 , y28709 , y28710 , y28711 , y28712 , y28713 , y28714 , y28715 , y28716 , y28717 , y28718 , y28719 , y28720 , y28721 , y28722 , y28723 , y28724 , y28725 , y28726 , y28727 , y28728 , y28729 , y28730 , y28731 , y28732 , y28733 , y28734 , y28735 , y28736 , y28737 , y28738 , y28739 , y28740 , y28741 , y28742 , y28743 , y28744 , y28745 , y28746 , y28747 , y28748 , y28749 , y28750 , y28751 , y28752 , y28753 , y28754 , y28755 , y28756 , y28757 , y28758 , y28759 , y28760 , y28761 , y28762 , y28763 , y28764 , y28765 , y28766 , y28767 , y28768 , y28769 , y28770 , y28771 , y28772 , y28773 , y28774 , y28775 , y28776 , y28777 , y28778 , y28779 , y28780 , y28781 , y28782 , y28783 , y28784 , y28785 , y28786 , y28787 , y28788 , y28789 , y28790 , y28791 , y28792 , y28793 , y28794 , y28795 , y28796 , y28797 , y28798 , y28799 , y28800 , y28801 , y28802 , y28803 , y28804 , y28805 , y28806 , y28807 , y28808 , y28809 , y28810 , y28811 , y28812 , y28813 , y28814 , y28815 , y28816 , y28817 , y28818 , y28819 , y28820 , y28821 , y28822 , y28823 , y28824 , y28825 , y28826 , y28827 , y28828 , y28829 , y28830 , y28831 , y28832 , y28833 , y28834 , y28835 , y28836 , y28837 , y28838 , y28839 , y28840 , y28841 , y28842 , y28843 , y28844 , y28845 , y28846 , y28847 , y28848 , y28849 , y28850 , y28851 , y28852 , y28853 , y28854 , y28855 , y28856 , y28857 , y28858 , y28859 , y28860 , y28861 , y28862 , y28863 , y28864 , y28865 , y28866 , y28867 , y28868 , y28869 , y28870 , y28871 , y28872 , y28873 , y28874 , y28875 , y28876 , y28877 , y28878 , y28879 , y28880 , y28881 , y28882 , y28883 , y28884 , y28885 , y28886 , y28887 , y28888 , y28889 , y28890 , y28891 , y28892 , y28893 , y28894 , y28895 , y28896 , y28897 , y28898 , y28899 , y28900 , y28901 , y28902 , y28903 , y28904 , y28905 , y28906 , y28907 , y28908 , y28909 , y28910 , y28911 , y28912 , y28913 , y28914 , y28915 , y28916 , y28917 , y28918 , y28919 , y28920 , y28921 , y28922 , y28923 , y28924 , y28925 , y28926 , y28927 , y28928 , y28929 , y28930 , y28931 , y28932 , y28933 , y28934 , y28935 , y28936 , y28937 , y28938 , y28939 , y28940 , y28941 , y28942 , y28943 , y28944 , y28945 , y28946 , y28947 , y28948 , y28949 , y28950 , y28951 , y28952 , y28953 , y28954 , y28955 , y28956 , y28957 , y28958 , y28959 , y28960 , y28961 , y28962 , y28963 , y28964 , y28965 , y28966 , y28967 , y28968 , y28969 , y28970 , y28971 , y28972 , y28973 , y28974 , y28975 , y28976 , y28977 , y28978 , y28979 , y28980 , y28981 , y28982 , y28983 , y28984 , y28985 , y28986 , y28987 , y28988 , y28989 , y28990 , y28991 , y28992 , y28993 , y28994 , y28995 , y28996 , y28997 , y28998 , y28999 , y29000 , y29001 , y29002 , y29003 , y29004 , y29005 , y29006 , y29007 , y29008 , y29009 , y29010 , y29011 , y29012 , y29013 , y29014 , y29015 , y29016 , y29017 , y29018 , y29019 , y29020 , y29021 , y29022 , y29023 , y29024 , y29025 , y29026 , y29027 , y29028 , y29029 , y29030 , y29031 , y29032 , y29033 , y29034 , y29035 , y29036 , y29037 , y29038 , y29039 , y29040 , y29041 , y29042 , y29043 , y29044 , y29045 , y29046 , y29047 , y29048 , y29049 , y29050 , y29051 , y29052 , y29053 , y29054 , y29055 , y29056 , y29057 , y29058 , y29059 , y29060 , y29061 , y29062 , y29063 , y29064 , y29065 , y29066 , y29067 , y29068 , y29069 , y29070 , y29071 , y29072 , y29073 , y29074 , y29075 , y29076 , y29077 , y29078 , y29079 , y29080 , y29081 , y29082 , y29083 , y29084 , y29085 , y29086 , y29087 , y29088 , y29089 , y29090 , y29091 , y29092 , y29093 , y29094 , y29095 , y29096 , y29097 , y29098 , y29099 , y29100 , y29101 , y29102 , y29103 , y29104 , y29105 , y29106 , y29107 , y29108 , y29109 , y29110 , y29111 , y29112 , y29113 , y29114 , y29115 , y29116 , y29117 , y29118 , y29119 , y29120 , y29121 , y29122 , y29123 , y29124 , y29125 , y29126 , y29127 , y29128 , y29129 , y29130 , y29131 , y29132 , y29133 , y29134 , y29135 , y29136 , y29137 , y29138 , y29139 , y29140 , y29141 , y29142 , y29143 , y29144 , y29145 , y29146 , y29147 , y29148 , y29149 , y29150 , y29151 , y29152 , y29153 , y29154 , y29155 , y29156 , y29157 , y29158 , y29159 , y29160 , y29161 , y29162 , y29163 , y29164 , y29165 , y29166 , y29167 , y29168 , y29169 , y29170 , y29171 , y29172 , y29173 , y29174 , y29175 , y29176 , y29177 , y29178 , y29179 , y29180 , y29181 , y29182 , y29183 , y29184 , y29185 , y29186 , y29187 , y29188 , y29189 , y29190 , y29191 , y29192 , y29193 , y29194 , y29195 , y29196 , y29197 , y29198 , y29199 , y29200 , y29201 , y29202 , y29203 , y29204 , y29205 , y29206 , y29207 , y29208 , y29209 , y29210 , y29211 , y29212 , y29213 , y29214 , y29215 , y29216 , y29217 , y29218 , y29219 , y29220 , y29221 , y29222 , y29223 , y29224 , y29225 , y29226 , y29227 , y29228 , y29229 , y29230 , y29231 , y29232 , y29233 , y29234 , y29235 , y29236 , y29237 , y29238 , y29239 , y29240 , y29241 , y29242 , y29243 , y29244 , y29245 , y29246 , y29247 , y29248 , y29249 , y29250 , y29251 , y29252 , y29253 , y29254 , y29255 , y29256 , y29257 , y29258 , y29259 , y29260 , y29261 , y29262 , y29263 , y29264 , y29265 , y29266 , y29267 , y29268 , y29269 , y29270 , y29271 , y29272 , y29273 , y29274 , y29275 , y29276 , y29277 , y29278 , y29279 , y29280 , y29281 , y29282 , y29283 , y29284 , y29285 , y29286 , y29287 , y29288 , y29289 , y29290 , y29291 , y29292 , y29293 , y29294 , y29295 , y29296 , y29297 , y29298 , y29299 , y29300 , y29301 , y29302 , y29303 , y29304 , y29305 , y29306 , y29307 , y29308 , y29309 , y29310 , y29311 , y29312 , y29313 , y29314 , y29315 , y29316 , y29317 , y29318 , y29319 , y29320 , y29321 , y29322 , y29323 , y29324 , y29325 , y29326 , y29327 , y29328 , y29329 , y29330 , y29331 , y29332 , y29333 , y29334 , y29335 , y29336 , y29337 , y29338 , y29339 , y29340 , y29341 , y29342 , y29343 , y29344 , y29345 , y29346 , y29347 , y29348 , y29349 , y29350 , y29351 , y29352 , y29353 , y29354 , y29355 , y29356 , y29357 , y29358 , y29359 , y29360 , y29361 , y29362 , y29363 , y29364 , y29365 , y29366 , y29367 , y29368 , y29369 , y29370 , y29371 , y29372 , y29373 , y29374 , y29375 , y29376 , y29377 , y29378 , y29379 , y29380 , y29381 , y29382 , y29383 , y29384 , y29385 , y29386 , y29387 , y29388 , y29389 , y29390 , y29391 , y29392 , y29393 , y29394 , y29395 , y29396 , y29397 , y29398 , y29399 , y29400 , y29401 , y29402 , y29403 , y29404 , y29405 , y29406 , y29407 , y29408 , y29409 , y29410 , y29411 , y29412 , y29413 , y29414 , y29415 , y29416 , y29417 , y29418 , y29419 , y29420 , y29421 , y29422 , y29423 , y29424 , y29425 , y29426 , y29427 , y29428 , y29429 , y29430 , y29431 , y29432 , y29433 , y29434 , y29435 , y29436 , y29437 , y29438 , y29439 , y29440 , y29441 , y29442 , y29443 , y29444 , y29445 , y29446 , y29447 , y29448 , y29449 , y29450 , y29451 , y29452 , y29453 , y29454 , y29455 , y29456 , y29457 , y29458 , y29459 , y29460 , y29461 , y29462 , y29463 , y29464 , y29465 , y29466 , y29467 , y29468 , y29469 , y29470 , y29471 , y29472 , y29473 , y29474 , y29475 , y29476 , y29477 , y29478 , y29479 , y29480 , y29481 , y29482 , y29483 , y29484 , y29485 , y29486 , y29487 , y29488 , y29489 , y29490 , y29491 , y29492 , y29493 , y29494 , y29495 , y29496 , y29497 , y29498 , y29499 , y29500 , y29501 , y29502 , y29503 , y29504 , y29505 , y29506 , y29507 , y29508 , y29509 , y29510 , y29511 , y29512 , y29513 , y29514 , y29515 , y29516 , y29517 , y29518 , y29519 , y29520 , y29521 , y29522 , y29523 , y29524 , y29525 , y29526 , y29527 , y29528 , y29529 , y29530 , y29531 , y29532 , y29533 , y29534 , y29535 , y29536 , y29537 , y29538 , y29539 , y29540 , y29541 , y29542 , y29543 , y29544 , y29545 , y29546 , y29547 , y29548 , y29549 , y29550 , y29551 , y29552 , y29553 , y29554 , y29555 , y29556 , y29557 , y29558 , y29559 , y29560 , y29561 , y29562 , y29563 , y29564 , y29565 , y29566 , y29567 , y29568 , y29569 , y29570 , y29571 , y29572 , y29573 , y29574 , y29575 , y29576 , y29577 , y29578 , y29579 , y29580 , y29581 , y29582 , y29583 , y29584 , y29585 , y29586 , y29587 , y29588 , y29589 , y29590 , y29591 , y29592 , y29593 , y29594 , y29595 , y29596 , y29597 , y29598 , y29599 , y29600 , y29601 , y29602 , y29603 , y29604 , y29605 , y29606 , y29607 , y29608 , y29609 , y29610 , y29611 , y29612 , y29613 , y29614 , y29615 , y29616 , y29617 , y29618 , y29619 , y29620 , y29621 , y29622 , y29623 , y29624 , y29625 , y29626 , y29627 , y29628 , y29629 , y29630 , y29631 , y29632 , y29633 , y29634 , y29635 , y29636 , y29637 , y29638 , y29639 , y29640 , y29641 , y29642 , y29643 , y29644 , y29645 , y29646 , y29647 , y29648 , y29649 , y29650 , y29651 , y29652 , y29653 , y29654 , y29655 , y29656 , y29657 , y29658 , y29659 , y29660 , y29661 , y29662 , y29663 , y29664 , y29665 , y29666 , y29667 , y29668 , y29669 , y29670 , y29671 , y29672 , y29673 , y29674 , y29675 , y29676 , y29677 , y29678 , y29679 , y29680 , y29681 , y29682 , y29683 , y29684 , y29685 , y29686 , y29687 , y29688 , y29689 , y29690 , y29691 , y29692 , y29693 , y29694 , y29695 , y29696 , y29697 , y29698 , y29699 , y29700 , y29701 , y29702 , y29703 , y29704 , y29705 , y29706 , y29707 , y29708 , y29709 , y29710 , y29711 , y29712 , y29713 , y29714 , y29715 , y29716 , y29717 , y29718 , y29719 , y29720 , y29721 , y29722 , y29723 , y29724 , y29725 , y29726 , y29727 , y29728 , y29729 , y29730 , y29731 , y29732 , y29733 , y29734 , y29735 , y29736 , y29737 , y29738 , y29739 , y29740 , y29741 , y29742 , y29743 , y29744 , y29745 , y29746 , y29747 , y29748 , y29749 , y29750 , y29751 , y29752 , y29753 , y29754 , y29755 , y29756 , y29757 , y29758 , y29759 , y29760 , y29761 , y29762 , y29763 , y29764 , y29765 , y29766 , y29767 , y29768 , y29769 , y29770 , y29771 , y29772 , y29773 , y29774 , y29775 , y29776 , y29777 , y29778 , y29779 , y29780 , y29781 , y29782 , y29783 , y29784 , y29785 , y29786 , y29787 , y29788 , y29789 , y29790 , y29791 , y29792 , y29793 , y29794 , y29795 , y29796 , y29797 , y29798 , y29799 , y29800 , y29801 , y29802 , y29803 , y29804 , y29805 , y29806 , y29807 , y29808 , y29809 , y29810 , y29811 , y29812 , y29813 , y29814 , y29815 , y29816 , y29817 , y29818 , y29819 , y29820 , y29821 , y29822 , y29823 , y29824 , y29825 , y29826 , y29827 , y29828 , y29829 , y29830 , y29831 , y29832 , y29833 , y29834 , y29835 , y29836 , y29837 , y29838 , y29839 , y29840 , y29841 , y29842 , y29843 , y29844 , y29845 , y29846 , y29847 , y29848 , y29849 , y29850 , y29851 , y29852 , y29853 , y29854 , y29855 , y29856 , y29857 , y29858 , y29859 , y29860 , y29861 , y29862 , y29863 , y29864 , y29865 , y29866 , y29867 , y29868 , y29869 , y29870 , y29871 , y29872 , y29873 , y29874 , y29875 , y29876 , y29877 , y29878 , y29879 , y29880 , y29881 , y29882 , y29883 , y29884 , y29885 , y29886 , y29887 , y29888 , y29889 , y29890 , y29891 , y29892 , y29893 , y29894 , y29895 , y29896 , y29897 , y29898 , y29899 , y29900 , y29901 , y29902 , y29903 , y29904 , y29905 , y29906 , y29907 , y29908 , y29909 , y29910 , y29911 , y29912 , y29913 , y29914 , y29915 , y29916 , y29917 , y29918 , y29919 , y29920 , y29921 , y29922 , y29923 , y29924 , y29925 , y29926 , y29927 , y29928 , y29929 , y29930 , y29931 , y29932 , y29933 , y29934 , y29935 , y29936 , y29937 , y29938 , y29939 , y29940 , y29941 , y29942 , y29943 , y29944 , y29945 , y29946 , y29947 , y29948 , y29949 , y29950 , y29951 , y29952 , y29953 , y29954 , y29955 , y29956 , y29957 , y29958 , y29959 , y29960 , y29961 , y29962 , y29963 , y29964 , y29965 , y29966 , y29967 , y29968 , y29969 , y29970 , y29971 , y29972 , y29973 , y29974 , y29975 , y29976 , y29977 , y29978 , y29979 , y29980 , y29981 , y29982 , y29983 , y29984 , y29985 , y29986 , y29987 , y29988 , y29989 , y29990 , y29991 , y29992 , y29993 , y29994 , y29995 , y29996 , y29997 , y29998 , y29999 , y30000 , y30001 , y30002 , y30003 , y30004 , y30005 , y30006 , y30007 , y30008 , y30009 , y30010 , y30011 , y30012 , y30013 , y30014 , y30015 , y30016 , y30017 , y30018 , y30019 , y30020 , y30021 , y30022 , y30023 , y30024 , y30025 , y30026 , y30027 , y30028 , y30029 , y30030 , y30031 , y30032 , y30033 , y30034 , y30035 , y30036 , y30037 , y30038 , y30039 , y30040 , y30041 , y30042 , y30043 , y30044 , y30045 , y30046 , y30047 , y30048 , y30049 , y30050 , y30051 , y30052 , y30053 , y30054 , y30055 , y30056 , y30057 , y30058 , y30059 , y30060 , y30061 , y30062 , y30063 , y30064 , y30065 , y30066 , y30067 , y30068 , y30069 , y30070 , y30071 , y30072 , y30073 , y30074 , y30075 , y30076 , y30077 , y30078 , y30079 , y30080 , y30081 , y30082 , y30083 , y30084 , y30085 , y30086 , y30087 , y30088 , y30089 , y30090 , y30091 , y30092 , y30093 , y30094 , y30095 , y30096 , y30097 , y30098 , y30099 , y30100 , y30101 , y30102 , y30103 , y30104 , y30105 , y30106 , y30107 , y30108 , y30109 , y30110 , y30111 , y30112 , y30113 , y30114 , y30115 , y30116 , y30117 , y30118 , y30119 , y30120 , y30121 , y30122 , y30123 , y30124 , y30125 , y30126 , y30127 , y30128 , y30129 , y30130 , y30131 , y30132 , y30133 , y30134 , y30135 , y30136 , y30137 , y30138 , y30139 , y30140 , y30141 , y30142 , y30143 , y30144 , y30145 , y30146 , y30147 , y30148 , y30149 , y30150 , y30151 , y30152 , y30153 , y30154 , y30155 , y30156 , y30157 , y30158 , y30159 , y30160 , y30161 , y30162 , y30163 , y30164 , y30165 , y30166 , y30167 , y30168 , y30169 , y30170 , y30171 , y30172 , y30173 , y30174 , y30175 , y30176 , y30177 , y30178 , y30179 , y30180 , y30181 , y30182 , y30183 , y30184 , y30185 , y30186 , y30187 , y30188 , y30189 , y30190 , y30191 , y30192 , y30193 , y30194 , y30195 , y30196 , y30197 , y30198 , y30199 , y30200 , y30201 , y30202 , y30203 , y30204 , y30205 , y30206 , y30207 , y30208 , y30209 , y30210 , y30211 , y30212 , y30213 , y30214 , y30215 , y30216 , y30217 , y30218 , y30219 , y30220 , y30221 , y30222 , y30223 , y30224 , y30225 , y30226 , y30227 , y30228 , y30229 , y30230 , y30231 , y30232 , y30233 , y30234 , y30235 , y30236 , y30237 , y30238 , y30239 , y30240 , y30241 , y30242 , y30243 , y30244 , y30245 , y30246 , y30247 , y30248 , y30249 , y30250 , y30251 , y30252 , y30253 , y30254 , y30255 , y30256 , y30257 , y30258 , y30259 , y30260 , y30261 , y30262 , y30263 , y30264 , y30265 , y30266 , y30267 , y30268 , y30269 , y30270 , y30271 , y30272 , y30273 , y30274 , y30275 , y30276 , y30277 , y30278 , y30279 , y30280 , y30281 , y30282 , y30283 , y30284 , y30285 , y30286 , y30287 , y30288 , y30289 , y30290 , y30291 , y30292 , y30293 , y30294 , y30295 , y30296 , y30297 , y30298 , y30299 , y30300 , y30301 , y30302 , y30303 , y30304 , y30305 , y30306 , y30307 , y30308 , y30309 , y30310 , y30311 , y30312 , y30313 , y30314 , y30315 , y30316 , y30317 , y30318 , y30319 , y30320 , y30321 , y30322 , y30323 , y30324 , y30325 , y30326 , y30327 , y30328 , y30329 , y30330 , y30331 , y30332 , y30333 , y30334 , y30335 , y30336 , y30337 , y30338 , y30339 , y30340 , y30341 , y30342 , y30343 , y30344 , y30345 , y30346 , y30347 , y30348 , y30349 , y30350 , y30351 , y30352 , y30353 , y30354 , y30355 , y30356 , y30357 , y30358 , y30359 , y30360 , y30361 , y30362 , y30363 , y30364 , y30365 , y30366 , y30367 , y30368 , y30369 , y30370 , y30371 , y30372 , y30373 , y30374 , y30375 , y30376 , y30377 , y30378 , y30379 , y30380 , y30381 , y30382 , y30383 , y30384 , y30385 , y30386 , y30387 , y30388 , y30389 , y30390 , y30391 , y30392 , y30393 , y30394 , y30395 , y30396 , y30397 , y30398 , y30399 , y30400 , y30401 , y30402 , y30403 , y30404 , y30405 , y30406 , y30407 , y30408 , y30409 , y30410 , y30411 , y30412 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 , y256 , y257 , y258 , y259 , y260 , y261 , y262 , y263 , y264 , y265 , y266 , y267 , y268 , y269 , y270 , y271 , y272 , y273 , y274 , y275 , y276 , y277 , y278 , y279 , y280 , y281 , y282 , y283 , y284 , y285 , y286 , y287 , y288 , y289 , y290 , y291 , y292 , y293 , y294 , y295 , y296 , y297 , y298 , y299 , y300 , y301 , y302 , y303 , y304 , y305 , y306 , y307 , y308 , y309 , y310 , y311 , y312 , y313 , y314 , y315 , y316 , y317 , y318 , y319 , y320 , y321 , y322 , y323 , y324 , y325 , y326 , y327 , y328 , y329 , y330 , y331 , y332 , y333 , y334 , y335 , y336 , y337 , y338 , y339 , y340 , y341 , y342 , y343 , y344 , y345 , y346 , y347 , y348 , y349 , y350 , y351 , y352 , y353 , y354 , y355 , y356 , y357 , y358 , y359 , y360 , y361 , y362 , y363 , y364 , y365 , y366 , y367 , y368 , y369 , y370 , y371 , y372 , y373 , y374 , y375 , y376 , y377 , y378 , y379 , y380 , y381 , y382 , y383 , y384 , y385 , y386 , y387 , y388 , y389 , y390 , y391 , y392 , y393 , y394 , y395 , y396 , y397 , y398 , y399 , y400 , y401 , y402 , y403 , y404 , y405 , y406 , y407 , y408 , y409 , y410 , y411 , y412 , y413 , y414 , y415 , y416 , y417 , y418 , y419 , y420 , y421 , y422 , y423 , y424 , y425 , y426 , y427 , y428 , y429 , y430 , y431 , y432 , y433 , y434 , y435 , y436 , y437 , y438 , y439 , y440 , y441 , y442 , y443 , y444 , y445 , y446 , y447 , y448 , y449 , y450 , y451 , y452 , y453 , y454 , y455 , y456 , y457 , y458 , y459 , y460 , y461 , y462 , y463 , y464 , y465 , y466 , y467 , y468 , y469 , y470 , y471 , y472 , y473 , y474 , y475 , y476 , y477 , y478 , y479 , y480 , y481 , y482 , y483 , y484 , y485 , y486 , y487 , y488 , y489 , y490 , y491 , y492 , y493 , y494 , y495 , y496 , y497 , y498 , y499 , y500 , y501 , y502 , y503 , y504 , y505 , y506 , y507 , y508 , y509 , y510 , y511 , y512 , y513 , y514 , y515 , y516 , y517 , y518 , y519 , y520 , y521 , y522 , y523 , y524 , y525 , y526 , y527 , y528 , y529 , y530 , y531 , y532 , y533 , y534 , y535 , y536 , y537 , y538 , y539 , y540 , y541 , y542 , y543 , y544 , y545 , y546 , y547 , y548 , y549 , y550 , y551 , y552 , y553 , y554 , y555 , y556 , y557 , y558 , y559 , y560 , y561 , y562 , y563 , y564 , y565 , y566 , y567 , y568 , y569 , y570 , y571 , y572 , y573 , y574 , y575 , y576 , y577 , y578 , y579 , y580 , y581 , y582 , y583 , y584 , y585 , y586 , y587 , y588 , y589 , y590 , y591 , y592 , y593 , y594 , y595 , y596 , y597 , y598 , y599 , y600 , y601 , y602 , y603 , y604 , y605 , y606 , y607 , y608 , y609 , y610 , y611 , y612 , y613 , y614 , y615 , y616 , y617 , y618 , y619 , y620 , y621 , y622 , y623 , y624 , y625 , y626 , y627 , y628 , y629 , y630 , y631 , y632 , y633 , y634 , y635 , y636 , y637 , y638 , y639 , y640 , y641 , y642 , y643 , y644 , y645 , y646 , y647 , y648 , y649 , y650 , y651 , y652 , y653 , y654 , y655 , y656 , y657 , y658 , y659 , y660 , y661 , y662 , y663 , y664 , y665 , y666 , y667 , y668 , y669 , y670 , y671 , y672 , y673 , y674 , y675 , y676 , y677 , y678 , y679 , y680 , y681 , y682 , y683 , y684 , y685 , y686 , y687 , y688 , y689 , y690 , y691 , y692 , y693 , y694 , y695 , y696 , y697 , y698 , y699 , y700 , y701 , y702 , y703 , y704 , y705 , y706 , y707 , y708 , y709 , y710 , y711 , y712 , y713 , y714 , y715 , y716 , y717 , y718 , y719 , y720 , y721 , y722 , y723 , y724 , y725 , y726 , y727 , y728 , y729 , y730 , y731 , y732 , y733 , y734 , y735 , y736 , y737 , y738 , y739 , y740 , y741 , y742 , y743 , y744 , y745 , y746 , y747 , y748 , y749 , y750 , y751 , y752 , y753 , y754 , y755 , y756 , y757 , y758 , y759 , y760 , y761 , y762 , y763 , y764 , y765 , y766 , y767 , y768 , y769 , y770 , y771 , y772 , y773 , y774 , y775 , y776 , y777 , y778 , y779 , y780 , y781 , y782 , y783 , y784 , y785 , y786 , y787 , y788 , y789 , y790 , y791 , y792 , y793 , y794 , y795 , y796 , y797 , y798 , y799 , y800 , y801 , y802 , y803 , y804 , y805 , y806 , y807 , y808 , y809 , y810 , y811 , y812 , y813 , y814 , y815 , y816 , y817 , y818 , y819 , y820 , y821 , y822 , y823 , y824 , y825 , y826 , y827 , y828 , y829 , y830 , y831 , y832 , y833 , y834 , y835 , y836 , y837 , y838 , y839 , y840 , y841 , y842 , y843 , y844 , y845 , y846 , y847 , y848 , y849 , y850 , y851 , y852 , y853 , y854 , y855 , y856 , y857 , y858 , y859 , y860 , y861 , y862 , y863 , y864 , y865 , y866 , y867 , y868 , y869 , y870 , y871 , y872 , y873 , y874 , y875 , y876 , y877 , y878 , y879 , y880 , y881 , y882 , y883 , y884 , y885 , y886 , y887 , y888 , y889 , y890 , y891 , y892 , y893 , y894 , y895 , y896 , y897 , y898 , y899 , y900 , y901 , y902 , y903 , y904 , y905 , y906 , y907 , y908 , y909 , y910 , y911 , y912 , y913 , y914 , y915 , y916 , y917 , y918 , y919 , y920 , y921 , y922 , y923 , y924 , y925 , y926 , y927 , y928 , y929 , y930 , y931 , y932 , y933 , y934 , y935 , y936 , y937 , y938 , y939 , y940 , y941 , y942 , y943 , y944 , y945 , y946 , y947 , y948 , y949 , y950 , y951 , y952 , y953 , y954 , y955 , y956 , y957 , y958 , y959 , y960 , y961 , y962 , y963 , y964 , y965 , y966 , y967 , y968 , y969 , y970 , y971 , y972 , y973 , y974 , y975 , y976 , y977 , y978 , y979 , y980 , y981 , y982 , y983 , y984 , y985 , y986 , y987 , y988 , y989 , y990 , y991 , y992 , y993 , y994 , y995 , y996 , y997 , y998 , y999 , y1000 , y1001 , y1002 , y1003 , y1004 , y1005 , y1006 , y1007 , y1008 , y1009 , y1010 , y1011 , y1012 , y1013 , y1014 , y1015 , y1016 , y1017 , y1018 , y1019 , y1020 , y1021 , y1022 , y1023 , y1024 , y1025 , y1026 , y1027 , y1028 , y1029 , y1030 , y1031 , y1032 , y1033 , y1034 , y1035 , y1036 , y1037 , y1038 , y1039 , y1040 , y1041 , y1042 , y1043 , y1044 , y1045 , y1046 , y1047 , y1048 , y1049 , y1050 , y1051 , y1052 , y1053 , y1054 , y1055 , y1056 , y1057 , y1058 , y1059 , y1060 , y1061 , y1062 , y1063 , y1064 , y1065 , y1066 , y1067 , y1068 , y1069 , y1070 , y1071 , y1072 , y1073 , y1074 , y1075 , y1076 , y1077 , y1078 , y1079 , y1080 , y1081 , y1082 , y1083 , y1084 , y1085 , y1086 , y1087 , y1088 , y1089 , y1090 , y1091 , y1092 , y1093 , y1094 , y1095 , y1096 , y1097 , y1098 , y1099 , y1100 , y1101 , y1102 , y1103 , y1104 , y1105 , y1106 , y1107 , y1108 , y1109 , y1110 , y1111 , y1112 , y1113 , y1114 , y1115 , y1116 , y1117 , y1118 , y1119 , y1120 , y1121 , y1122 , y1123 , y1124 , y1125 , y1126 , y1127 , y1128 , y1129 , y1130 , y1131 , y1132 , y1133 , y1134 , y1135 , y1136 , y1137 , y1138 , y1139 , y1140 , y1141 , y1142 , y1143 , y1144 , y1145 , y1146 , y1147 , y1148 , y1149 , y1150 , y1151 , y1152 , y1153 , y1154 , y1155 , y1156 , y1157 , y1158 , y1159 , y1160 , y1161 , y1162 , y1163 , y1164 , y1165 , y1166 , y1167 , y1168 , y1169 , y1170 , y1171 , y1172 , y1173 , y1174 , y1175 , y1176 , y1177 , y1178 , y1179 , y1180 , y1181 , y1182 , y1183 , y1184 , y1185 , y1186 , y1187 , y1188 , y1189 , y1190 , y1191 , y1192 , y1193 , y1194 , y1195 , y1196 , y1197 , y1198 , y1199 , y1200 , y1201 , y1202 , y1203 , y1204 , y1205 , y1206 , y1207 , y1208 , y1209 , y1210 , y1211 , y1212 , y1213 , y1214 , y1215 , y1216 , y1217 , y1218 , y1219 , y1220 , y1221 , y1222 , y1223 , y1224 , y1225 , y1226 , y1227 , y1228 , y1229 , y1230 , y1231 , y1232 , y1233 , y1234 , y1235 , y1236 , y1237 , y1238 , y1239 , y1240 , y1241 , y1242 , y1243 , y1244 , y1245 , y1246 , y1247 , y1248 , y1249 , y1250 , y1251 , y1252 , y1253 , y1254 , y1255 , y1256 , y1257 , y1258 , y1259 , y1260 , y1261 , y1262 , y1263 , y1264 , y1265 , y1266 , y1267 , y1268 , y1269 , y1270 , y1271 , y1272 , y1273 , y1274 , y1275 , y1276 , y1277 , y1278 , y1279 , y1280 , y1281 , y1282 , y1283 , y1284 , y1285 , y1286 , y1287 , y1288 , y1289 , y1290 , y1291 , y1292 , y1293 , y1294 , y1295 , y1296 , y1297 , y1298 , y1299 , y1300 , y1301 , y1302 , y1303 , y1304 , y1305 , y1306 , y1307 , y1308 , y1309 , y1310 , y1311 , y1312 , y1313 , y1314 , y1315 , y1316 , y1317 , y1318 , y1319 , y1320 , y1321 , y1322 , y1323 , y1324 , y1325 , y1326 , y1327 , y1328 , y1329 , y1330 , y1331 , y1332 , y1333 , y1334 , y1335 , y1336 , y1337 , y1338 , y1339 , y1340 , y1341 , y1342 , y1343 , y1344 , y1345 , y1346 , y1347 , y1348 , y1349 , y1350 , y1351 , y1352 , y1353 , y1354 , y1355 , y1356 , y1357 , y1358 , y1359 , y1360 , y1361 , y1362 , y1363 , y1364 , y1365 , y1366 , y1367 , y1368 , y1369 , y1370 , y1371 , y1372 , y1373 , y1374 , y1375 , y1376 , y1377 , y1378 , y1379 , y1380 , y1381 , y1382 , y1383 , y1384 , y1385 , y1386 , y1387 , y1388 , y1389 , y1390 , y1391 , y1392 , y1393 , y1394 , y1395 , y1396 , y1397 , y1398 , y1399 , y1400 , y1401 , y1402 , y1403 , y1404 , y1405 , y1406 , y1407 , y1408 , y1409 , y1410 , y1411 , y1412 , y1413 , y1414 , y1415 , y1416 , y1417 , y1418 , y1419 , y1420 , y1421 , y1422 , y1423 , y1424 , y1425 , y1426 , y1427 , y1428 , y1429 , y1430 , y1431 , y1432 , y1433 , y1434 , y1435 , y1436 , y1437 , y1438 , y1439 , y1440 , y1441 , y1442 , y1443 , y1444 , y1445 , y1446 , y1447 , y1448 , y1449 , y1450 , y1451 , y1452 , y1453 , y1454 , y1455 , y1456 , y1457 , y1458 , y1459 , y1460 , y1461 , y1462 , y1463 , y1464 , y1465 , y1466 , y1467 , y1468 , y1469 , y1470 , y1471 , y1472 , y1473 , y1474 , y1475 , y1476 , y1477 , y1478 , y1479 , y1480 , y1481 , y1482 , y1483 , y1484 , y1485 , y1486 , y1487 , y1488 , y1489 , y1490 , y1491 , y1492 , y1493 , y1494 , y1495 , y1496 , y1497 , y1498 , y1499 , y1500 , y1501 , y1502 , y1503 , y1504 , y1505 , y1506 , y1507 , y1508 , y1509 , y1510 , y1511 , y1512 , y1513 , y1514 , y1515 , y1516 , y1517 , y1518 , y1519 , y1520 , y1521 , y1522 , y1523 , y1524 , y1525 , y1526 , y1527 , y1528 , y1529 , y1530 , y1531 , y1532 , y1533 , y1534 , y1535 , y1536 , y1537 , y1538 , y1539 , y1540 , y1541 , y1542 , y1543 , y1544 , y1545 , y1546 , y1547 , y1548 , y1549 , y1550 , y1551 , y1552 , y1553 , y1554 , y1555 , y1556 , y1557 , y1558 , y1559 , y1560 , y1561 , y1562 , y1563 , y1564 , y1565 , y1566 , y1567 , y1568 , y1569 , y1570 , y1571 , y1572 , y1573 , y1574 , y1575 , y1576 , y1577 , y1578 , y1579 , y1580 , y1581 , y1582 , y1583 , y1584 , y1585 , y1586 , y1587 , y1588 , y1589 , y1590 , y1591 , y1592 , y1593 , y1594 , y1595 , y1596 , y1597 , y1598 , y1599 , y1600 , y1601 , y1602 , y1603 , y1604 , y1605 , y1606 , y1607 , y1608 , y1609 , y1610 , y1611 , y1612 , y1613 , y1614 , y1615 , y1616 , y1617 , y1618 , y1619 , y1620 , y1621 , y1622 , y1623 , y1624 , y1625 , y1626 , y1627 , y1628 , y1629 , y1630 , y1631 , y1632 , y1633 , y1634 , y1635 , y1636 , y1637 , y1638 , y1639 , y1640 , y1641 , y1642 , y1643 , y1644 , y1645 , y1646 , y1647 , y1648 , y1649 , y1650 , y1651 , y1652 , y1653 , y1654 , y1655 , y1656 , y1657 , y1658 , y1659 , y1660 , y1661 , y1662 , y1663 , y1664 , y1665 , y1666 , y1667 , y1668 , y1669 , y1670 , y1671 , y1672 , y1673 , y1674 , y1675 , y1676 , y1677 , y1678 , y1679 , y1680 , y1681 , y1682 , y1683 , y1684 , y1685 , y1686 , y1687 , y1688 , y1689 , y1690 , y1691 , y1692 , y1693 , y1694 , y1695 , y1696 , y1697 , y1698 , y1699 , y1700 , y1701 , y1702 , y1703 , y1704 , y1705 , y1706 , y1707 , y1708 , y1709 , y1710 , y1711 , y1712 , y1713 , y1714 , y1715 , y1716 , y1717 , y1718 , y1719 , y1720 , y1721 , y1722 , y1723 , y1724 , y1725 , y1726 , y1727 , y1728 , y1729 , y1730 , y1731 , y1732 , y1733 , y1734 , y1735 , y1736 , y1737 , y1738 , y1739 , y1740 , y1741 , y1742 , y1743 , y1744 , y1745 , y1746 , y1747 , y1748 , y1749 , y1750 , y1751 , y1752 , y1753 , y1754 , y1755 , y1756 , y1757 , y1758 , y1759 , y1760 , y1761 , y1762 , y1763 , y1764 , y1765 , y1766 , y1767 , y1768 , y1769 , y1770 , y1771 , y1772 , y1773 , y1774 , y1775 , y1776 , y1777 , y1778 , y1779 , y1780 , y1781 , y1782 , y1783 , y1784 , y1785 , y1786 , y1787 , y1788 , y1789 , y1790 , y1791 , y1792 , y1793 , y1794 , y1795 , y1796 , y1797 , y1798 , y1799 , y1800 , y1801 , y1802 , y1803 , y1804 , y1805 , y1806 , y1807 , y1808 , y1809 , y1810 , y1811 , y1812 , y1813 , y1814 , y1815 , y1816 , y1817 , y1818 , y1819 , y1820 , y1821 , y1822 , y1823 , y1824 , y1825 , y1826 , y1827 , y1828 , y1829 , y1830 , y1831 , y1832 , y1833 , y1834 , y1835 , y1836 , y1837 , y1838 , y1839 , y1840 , y1841 , y1842 , y1843 , y1844 , y1845 , y1846 , y1847 , y1848 , y1849 , y1850 , y1851 , y1852 , y1853 , y1854 , y1855 , y1856 , y1857 , y1858 , y1859 , y1860 , y1861 , y1862 , y1863 , y1864 , y1865 , y1866 , y1867 , y1868 , y1869 , y1870 , y1871 , y1872 , y1873 , y1874 , y1875 , y1876 , y1877 , y1878 , y1879 , y1880 , y1881 , y1882 , y1883 , y1884 , y1885 , y1886 , y1887 , y1888 , y1889 , y1890 , y1891 , y1892 , y1893 , y1894 , y1895 , y1896 , y1897 , y1898 , y1899 , y1900 , y1901 , y1902 , y1903 , y1904 , y1905 , y1906 , y1907 , y1908 , y1909 , y1910 , y1911 , y1912 , y1913 , y1914 , y1915 , y1916 , y1917 , y1918 , y1919 , y1920 , y1921 , y1922 , y1923 , y1924 , y1925 , y1926 , y1927 , y1928 , y1929 , y1930 , y1931 , y1932 , y1933 , y1934 , y1935 , y1936 , y1937 , y1938 , y1939 , y1940 , y1941 , y1942 , y1943 , y1944 , y1945 , y1946 , y1947 , y1948 , y1949 , y1950 , y1951 , y1952 , y1953 , y1954 , y1955 , y1956 , y1957 , y1958 , y1959 , y1960 , y1961 , y1962 , y1963 , y1964 , y1965 , y1966 , y1967 , y1968 , y1969 , y1970 , y1971 , y1972 , y1973 , y1974 , y1975 , y1976 , y1977 , y1978 , y1979 , y1980 , y1981 , y1982 , y1983 , y1984 , y1985 , y1986 , y1987 , y1988 , y1989 , y1990 , y1991 , y1992 , y1993 , y1994 , y1995 , y1996 , y1997 , y1998 , y1999 , y2000 , y2001 , y2002 , y2003 , y2004 , y2005 , y2006 , y2007 , y2008 , y2009 , y2010 , y2011 , y2012 , y2013 , y2014 , y2015 , y2016 , y2017 , y2018 , y2019 , y2020 , y2021 , y2022 , y2023 , y2024 , y2025 , y2026 , y2027 , y2028 , y2029 , y2030 , y2031 , y2032 , y2033 , y2034 , y2035 , y2036 , y2037 , y2038 , y2039 , y2040 , y2041 , y2042 , y2043 , y2044 , y2045 , y2046 , y2047 , y2048 , y2049 , y2050 , y2051 , y2052 , y2053 , y2054 , y2055 , y2056 , y2057 , y2058 , y2059 , y2060 , y2061 , y2062 , y2063 , y2064 , y2065 , y2066 , y2067 , y2068 , y2069 , y2070 , y2071 , y2072 , y2073 , y2074 , y2075 , y2076 , y2077 , y2078 , y2079 , y2080 , y2081 , y2082 , y2083 , y2084 , y2085 , y2086 , y2087 , y2088 , y2089 , y2090 , y2091 , y2092 , y2093 , y2094 , y2095 , y2096 , y2097 , y2098 , y2099 , y2100 , y2101 , y2102 , y2103 , y2104 , y2105 , y2106 , y2107 , y2108 , y2109 , y2110 , y2111 , y2112 , y2113 , y2114 , y2115 , y2116 , y2117 , y2118 , y2119 , y2120 , y2121 , y2122 , y2123 , y2124 , y2125 , y2126 , y2127 , y2128 , y2129 , y2130 , y2131 , y2132 , y2133 , y2134 , y2135 , y2136 , y2137 , y2138 , y2139 , y2140 , y2141 , y2142 , y2143 , y2144 , y2145 , y2146 , y2147 , y2148 , y2149 , y2150 , y2151 , y2152 , y2153 , y2154 , y2155 , y2156 , y2157 , y2158 , y2159 , y2160 , y2161 , y2162 , y2163 , y2164 , y2165 , y2166 , y2167 , y2168 , y2169 , y2170 , y2171 , y2172 , y2173 , y2174 , y2175 , y2176 , y2177 , y2178 , y2179 , y2180 , y2181 , y2182 , y2183 , y2184 , y2185 , y2186 , y2187 , y2188 , y2189 , y2190 , y2191 , y2192 , y2193 , y2194 , y2195 , y2196 , y2197 , y2198 , y2199 , y2200 , y2201 , y2202 , y2203 , y2204 , y2205 , y2206 , y2207 , y2208 , y2209 , y2210 , y2211 , y2212 , y2213 , y2214 , y2215 , y2216 , y2217 , y2218 , y2219 , y2220 , y2221 , y2222 , y2223 , y2224 , y2225 , y2226 , y2227 , y2228 , y2229 , y2230 , y2231 , y2232 , y2233 , y2234 , y2235 , y2236 , y2237 , y2238 , y2239 , y2240 , y2241 , y2242 , y2243 , y2244 , y2245 , y2246 , y2247 , y2248 , y2249 , y2250 , y2251 , y2252 , y2253 , y2254 , y2255 , y2256 , y2257 , y2258 , y2259 , y2260 , y2261 , y2262 , y2263 , y2264 , y2265 , y2266 , y2267 , y2268 , y2269 , y2270 , y2271 , y2272 , y2273 , y2274 , y2275 , y2276 , y2277 , y2278 , y2279 , y2280 , y2281 , y2282 , y2283 , y2284 , y2285 , y2286 , y2287 , y2288 , y2289 , y2290 , y2291 , y2292 , y2293 , y2294 , y2295 , y2296 , y2297 , y2298 , y2299 , y2300 , y2301 , y2302 , y2303 , y2304 , y2305 , y2306 , y2307 , y2308 , y2309 , y2310 , y2311 , y2312 , y2313 , y2314 , y2315 , y2316 , y2317 , y2318 , y2319 , y2320 , y2321 , y2322 , y2323 , y2324 , y2325 , y2326 , y2327 , y2328 , y2329 , y2330 , y2331 , y2332 , y2333 , y2334 , y2335 , y2336 , y2337 , y2338 , y2339 , y2340 , y2341 , y2342 , y2343 , y2344 , y2345 , y2346 , y2347 , y2348 , y2349 , y2350 , y2351 , y2352 , y2353 , y2354 , y2355 , y2356 , y2357 , y2358 , y2359 , y2360 , y2361 , y2362 , y2363 , y2364 , y2365 , y2366 , y2367 , y2368 , y2369 , y2370 , y2371 , y2372 , y2373 , y2374 , y2375 , y2376 , y2377 , y2378 , y2379 , y2380 , y2381 , y2382 , y2383 , y2384 , y2385 , y2386 , y2387 , y2388 , y2389 , y2390 , y2391 , y2392 , y2393 , y2394 , y2395 , y2396 , y2397 , y2398 , y2399 , y2400 , y2401 , y2402 , y2403 , y2404 , y2405 , y2406 , y2407 , y2408 , y2409 , y2410 , y2411 , y2412 , y2413 , y2414 , y2415 , y2416 , y2417 , y2418 , y2419 , y2420 , y2421 , y2422 , y2423 , y2424 , y2425 , y2426 , y2427 , y2428 , y2429 , y2430 , y2431 , y2432 , y2433 , y2434 , y2435 , y2436 , y2437 , y2438 , y2439 , y2440 , y2441 , y2442 , y2443 , y2444 , y2445 , y2446 , y2447 , y2448 , y2449 , y2450 , y2451 , y2452 , y2453 , y2454 , y2455 , y2456 , y2457 , y2458 , y2459 , y2460 , y2461 , y2462 , y2463 , y2464 , y2465 , y2466 , y2467 , y2468 , y2469 , y2470 , y2471 , y2472 , y2473 , y2474 , y2475 , y2476 , y2477 , y2478 , y2479 , y2480 , y2481 , y2482 , y2483 , y2484 , y2485 , y2486 , y2487 , y2488 , y2489 , y2490 , y2491 , y2492 , y2493 , y2494 , y2495 , y2496 , y2497 , y2498 , y2499 , y2500 , y2501 , y2502 , y2503 , y2504 , y2505 , y2506 , y2507 , y2508 , y2509 , y2510 , y2511 , y2512 , y2513 , y2514 , y2515 , y2516 , y2517 , y2518 , y2519 , y2520 , y2521 , y2522 , y2523 , y2524 , y2525 , y2526 , y2527 , y2528 , y2529 , y2530 , y2531 , y2532 , y2533 , y2534 , y2535 , y2536 , y2537 , y2538 , y2539 , y2540 , y2541 , y2542 , y2543 , y2544 , y2545 , y2546 , y2547 , y2548 , y2549 , y2550 , y2551 , y2552 , y2553 , y2554 , y2555 , y2556 , y2557 , y2558 , y2559 , y2560 , y2561 , y2562 , y2563 , y2564 , y2565 , y2566 , y2567 , y2568 , y2569 , y2570 , y2571 , y2572 , y2573 , y2574 , y2575 , y2576 , y2577 , y2578 , y2579 , y2580 , y2581 , y2582 , y2583 , y2584 , y2585 , y2586 , y2587 , y2588 , y2589 , y2590 , y2591 , y2592 , y2593 , y2594 , y2595 , y2596 , y2597 , y2598 , y2599 , y2600 , y2601 , y2602 , y2603 , y2604 , y2605 , y2606 , y2607 , y2608 , y2609 , y2610 , y2611 , y2612 , y2613 , y2614 , y2615 , y2616 , y2617 , y2618 , y2619 , y2620 , y2621 , y2622 , y2623 , y2624 , y2625 , y2626 , y2627 , y2628 , y2629 , y2630 , y2631 , y2632 , y2633 , y2634 , y2635 , y2636 , y2637 , y2638 , y2639 , y2640 , y2641 , y2642 , y2643 , y2644 , y2645 , y2646 , y2647 , y2648 , y2649 , y2650 , y2651 , y2652 , y2653 , y2654 , y2655 , y2656 , y2657 , y2658 , y2659 , y2660 , y2661 , y2662 , y2663 , y2664 , y2665 , y2666 , y2667 , y2668 , y2669 , y2670 , y2671 , y2672 , y2673 , y2674 , y2675 , y2676 , y2677 , y2678 , y2679 , y2680 , y2681 , y2682 , y2683 , y2684 , y2685 , y2686 , y2687 , y2688 , y2689 , y2690 , y2691 , y2692 , y2693 , y2694 , y2695 , y2696 , y2697 , y2698 , y2699 , y2700 , y2701 , y2702 , y2703 , y2704 , y2705 , y2706 , y2707 , y2708 , y2709 , y2710 , y2711 , y2712 , y2713 , y2714 , y2715 , y2716 , y2717 , y2718 , y2719 , y2720 , y2721 , y2722 , y2723 , y2724 , y2725 , y2726 , y2727 , y2728 , y2729 , y2730 , y2731 , y2732 , y2733 , y2734 , y2735 , y2736 , y2737 , y2738 , y2739 , y2740 , y2741 , y2742 , y2743 , y2744 , y2745 , y2746 , y2747 , y2748 , y2749 , y2750 , y2751 , y2752 , y2753 , y2754 , y2755 , y2756 , y2757 , y2758 , y2759 , y2760 , y2761 , y2762 , y2763 , y2764 , y2765 , y2766 , y2767 , y2768 , y2769 , y2770 , y2771 , y2772 , y2773 , y2774 , y2775 , y2776 , y2777 , y2778 , y2779 , y2780 , y2781 , y2782 , y2783 , y2784 , y2785 , y2786 , y2787 , y2788 , y2789 , y2790 , y2791 , y2792 , y2793 , y2794 , y2795 , y2796 , y2797 , y2798 , y2799 , y2800 , y2801 , y2802 , y2803 , y2804 , y2805 , y2806 , y2807 , y2808 , y2809 , y2810 , y2811 , y2812 , y2813 , y2814 , y2815 , y2816 , y2817 , y2818 , y2819 , y2820 , y2821 , y2822 , y2823 , y2824 , y2825 , y2826 , y2827 , y2828 , y2829 , y2830 , y2831 , y2832 , y2833 , y2834 , y2835 , y2836 , y2837 , y2838 , y2839 , y2840 , y2841 , y2842 , y2843 , y2844 , y2845 , y2846 , y2847 , y2848 , y2849 , y2850 , y2851 , y2852 , y2853 , y2854 , y2855 , y2856 , y2857 , y2858 , y2859 , y2860 , y2861 , y2862 , y2863 , y2864 , y2865 , y2866 , y2867 , y2868 , y2869 , y2870 , y2871 , y2872 , y2873 , y2874 , y2875 , y2876 , y2877 , y2878 , y2879 , y2880 , y2881 , y2882 , y2883 , y2884 , y2885 , y2886 , y2887 , y2888 , y2889 , y2890 , y2891 , y2892 , y2893 , y2894 , y2895 , y2896 , y2897 , y2898 , y2899 , y2900 , y2901 , y2902 , y2903 , y2904 , y2905 , y2906 , y2907 , y2908 , y2909 , y2910 , y2911 , y2912 , y2913 , y2914 , y2915 , y2916 , y2917 , y2918 , y2919 , y2920 , y2921 , y2922 , y2923 , y2924 , y2925 , y2926 , y2927 , y2928 , y2929 , y2930 , y2931 , y2932 , y2933 , y2934 , y2935 , y2936 , y2937 , y2938 , y2939 , y2940 , y2941 , y2942 , y2943 , y2944 , y2945 , y2946 , y2947 , y2948 , y2949 , y2950 , y2951 , y2952 , y2953 , y2954 , y2955 , y2956 , y2957 , y2958 , y2959 , y2960 , y2961 , y2962 , y2963 , y2964 , y2965 , y2966 , y2967 , y2968 , y2969 , y2970 , y2971 , y2972 , y2973 , y2974 , y2975 , y2976 , y2977 , y2978 , y2979 , y2980 , y2981 , y2982 , y2983 , y2984 , y2985 , y2986 , y2987 , y2988 , y2989 , y2990 , y2991 , y2992 , y2993 , y2994 , y2995 , y2996 , y2997 , y2998 , y2999 , y3000 , y3001 , y3002 , y3003 , y3004 , y3005 , y3006 , y3007 , y3008 , y3009 , y3010 , y3011 , y3012 , y3013 , y3014 , y3015 , y3016 , y3017 , y3018 , y3019 , y3020 , y3021 , y3022 , y3023 , y3024 , y3025 , y3026 , y3027 , y3028 , y3029 , y3030 , y3031 , y3032 , y3033 , y3034 , y3035 , y3036 , y3037 , y3038 , y3039 , y3040 , y3041 , y3042 , y3043 , y3044 , y3045 , y3046 , y3047 , y3048 , y3049 , y3050 , y3051 , y3052 , y3053 , y3054 , y3055 , y3056 , y3057 , y3058 , y3059 , y3060 , y3061 , y3062 , y3063 , y3064 , y3065 , y3066 , y3067 , y3068 , y3069 , y3070 , y3071 , y3072 , y3073 , y3074 , y3075 , y3076 , y3077 , y3078 , y3079 , y3080 , y3081 , y3082 , y3083 , y3084 , y3085 , y3086 , y3087 , y3088 , y3089 , y3090 , y3091 , y3092 , y3093 , y3094 , y3095 , y3096 , y3097 , y3098 , y3099 , y3100 , y3101 , y3102 , y3103 , y3104 , y3105 , y3106 , y3107 , y3108 , y3109 , y3110 , y3111 , y3112 , y3113 , y3114 , y3115 , y3116 , y3117 , y3118 , y3119 , y3120 , y3121 , y3122 , y3123 , y3124 , y3125 , y3126 , y3127 , y3128 , y3129 , y3130 , y3131 , y3132 , y3133 , y3134 , y3135 , y3136 , y3137 , y3138 , y3139 , y3140 , y3141 , y3142 , y3143 , y3144 , y3145 , y3146 , y3147 , y3148 , y3149 , y3150 , y3151 , y3152 , y3153 , y3154 , y3155 , y3156 , y3157 , y3158 , y3159 , y3160 , y3161 , y3162 , y3163 , y3164 , y3165 , y3166 , y3167 , y3168 , y3169 , y3170 , y3171 , y3172 , y3173 , y3174 , y3175 , y3176 , y3177 , y3178 , y3179 , y3180 , y3181 , y3182 , y3183 , y3184 , y3185 , y3186 , y3187 , y3188 , y3189 , y3190 , y3191 , y3192 , y3193 , y3194 , y3195 , y3196 , y3197 , y3198 , y3199 , y3200 , y3201 , y3202 , y3203 , y3204 , y3205 , y3206 , y3207 , y3208 , y3209 , y3210 , y3211 , y3212 , y3213 , y3214 , y3215 , y3216 , y3217 , y3218 , y3219 , y3220 , y3221 , y3222 , y3223 , y3224 , y3225 , y3226 , y3227 , y3228 , y3229 , y3230 , y3231 , y3232 , y3233 , y3234 , y3235 , y3236 , y3237 , y3238 , y3239 , y3240 , y3241 , y3242 , y3243 , y3244 , y3245 , y3246 , y3247 , y3248 , y3249 , y3250 , y3251 , y3252 , y3253 , y3254 , y3255 , y3256 , y3257 , y3258 , y3259 , y3260 , y3261 , y3262 , y3263 , y3264 , y3265 , y3266 , y3267 , y3268 , y3269 , y3270 , y3271 , y3272 , y3273 , y3274 , y3275 , y3276 , y3277 , y3278 , y3279 , y3280 , y3281 , y3282 , y3283 , y3284 , y3285 , y3286 , y3287 , y3288 , y3289 , y3290 , y3291 , y3292 , y3293 , y3294 , y3295 , y3296 , y3297 , y3298 , y3299 , y3300 , y3301 , y3302 , y3303 , y3304 , y3305 , y3306 , y3307 , y3308 , y3309 , y3310 , y3311 , y3312 , y3313 , y3314 , y3315 , y3316 , y3317 , y3318 , y3319 , y3320 , y3321 , y3322 , y3323 , y3324 , y3325 , y3326 , y3327 , y3328 , y3329 , y3330 , y3331 , y3332 , y3333 , y3334 , y3335 , y3336 , y3337 , y3338 , y3339 , y3340 , y3341 , y3342 , y3343 , y3344 , y3345 , y3346 , y3347 , y3348 , y3349 , y3350 , y3351 , y3352 , y3353 , y3354 , y3355 , y3356 , y3357 , y3358 , y3359 , y3360 , y3361 , y3362 , y3363 , y3364 , y3365 , y3366 , y3367 , y3368 , y3369 , y3370 , y3371 , y3372 , y3373 , y3374 , y3375 , y3376 , y3377 , y3378 , y3379 , y3380 , y3381 , y3382 , y3383 , y3384 , y3385 , y3386 , y3387 , y3388 , y3389 , y3390 , y3391 , y3392 , y3393 , y3394 , y3395 , y3396 , y3397 , y3398 , y3399 , y3400 , y3401 , y3402 , y3403 , y3404 , y3405 , y3406 , y3407 , y3408 , y3409 , y3410 , y3411 , y3412 , y3413 , y3414 , y3415 , y3416 , y3417 , y3418 , y3419 , y3420 , y3421 , y3422 , y3423 , y3424 , y3425 , y3426 , y3427 , y3428 , y3429 , y3430 , y3431 , y3432 , y3433 , y3434 , y3435 , y3436 , y3437 , y3438 , y3439 , y3440 , y3441 , y3442 , y3443 , y3444 , y3445 , y3446 , y3447 , y3448 , y3449 , y3450 , y3451 , y3452 , y3453 , y3454 , y3455 , y3456 , y3457 , y3458 , y3459 , y3460 , y3461 , y3462 , y3463 , y3464 , y3465 , y3466 , y3467 , y3468 , y3469 , y3470 , y3471 , y3472 , y3473 , y3474 , y3475 , y3476 , y3477 , y3478 , y3479 , y3480 , y3481 , y3482 , y3483 , y3484 , y3485 , y3486 , y3487 , y3488 , y3489 , y3490 , y3491 , y3492 , y3493 , y3494 , y3495 , y3496 , y3497 , y3498 , y3499 , y3500 , y3501 , y3502 , y3503 , y3504 , y3505 , y3506 , y3507 , y3508 , y3509 , y3510 , y3511 , y3512 , y3513 , y3514 , y3515 , y3516 , y3517 , y3518 , y3519 , y3520 , y3521 , y3522 , y3523 , y3524 , y3525 , y3526 , y3527 , y3528 , y3529 , y3530 , y3531 , y3532 , y3533 , y3534 , y3535 , y3536 , y3537 , y3538 , y3539 , y3540 , y3541 , y3542 , y3543 , y3544 , y3545 , y3546 , y3547 , y3548 , y3549 , y3550 , y3551 , y3552 , y3553 , y3554 , y3555 , y3556 , y3557 , y3558 , y3559 , y3560 , y3561 , y3562 , y3563 , y3564 , y3565 , y3566 , y3567 , y3568 , y3569 , y3570 , y3571 , y3572 , y3573 , y3574 , y3575 , y3576 , y3577 , y3578 , y3579 , y3580 , y3581 , y3582 , y3583 , y3584 , y3585 , y3586 , y3587 , y3588 , y3589 , y3590 , y3591 , y3592 , y3593 , y3594 , y3595 , y3596 , y3597 , y3598 , y3599 , y3600 , y3601 , y3602 , y3603 , y3604 , y3605 , y3606 , y3607 , y3608 , y3609 , y3610 , y3611 , y3612 , y3613 , y3614 , y3615 , y3616 , y3617 , y3618 , y3619 , y3620 , y3621 , y3622 , y3623 , y3624 , y3625 , y3626 , y3627 , y3628 , y3629 , y3630 , y3631 , y3632 , y3633 , y3634 , y3635 , y3636 , y3637 , y3638 , y3639 , y3640 , y3641 , y3642 , y3643 , y3644 , y3645 , y3646 , y3647 , y3648 , y3649 , y3650 , y3651 , y3652 , y3653 , y3654 , y3655 , y3656 , y3657 , y3658 , y3659 , y3660 , y3661 , y3662 , y3663 , y3664 , y3665 , y3666 , y3667 , y3668 , y3669 , y3670 , y3671 , y3672 , y3673 , y3674 , y3675 , y3676 , y3677 , y3678 , y3679 , y3680 , y3681 , y3682 , y3683 , y3684 , y3685 , y3686 , y3687 , y3688 , y3689 , y3690 , y3691 , y3692 , y3693 , y3694 , y3695 , y3696 , y3697 , y3698 , y3699 , y3700 , y3701 , y3702 , y3703 , y3704 , y3705 , y3706 , y3707 , y3708 , y3709 , y3710 , y3711 , y3712 , y3713 , y3714 , y3715 , y3716 , y3717 , y3718 , y3719 , y3720 , y3721 , y3722 , y3723 , y3724 , y3725 , y3726 , y3727 , y3728 , y3729 , y3730 , y3731 , y3732 , y3733 , y3734 , y3735 , y3736 , y3737 , y3738 , y3739 , y3740 , y3741 , y3742 , y3743 , y3744 , y3745 , y3746 , y3747 , y3748 , y3749 , y3750 , y3751 , y3752 , y3753 , y3754 , y3755 , y3756 , y3757 , y3758 , y3759 , y3760 , y3761 , y3762 , y3763 , y3764 , y3765 , y3766 , y3767 , y3768 , y3769 , y3770 , y3771 , y3772 , y3773 , y3774 , y3775 , y3776 , y3777 , y3778 , y3779 , y3780 , y3781 , y3782 , y3783 , y3784 , y3785 , y3786 , y3787 , y3788 , y3789 , y3790 , y3791 , y3792 , y3793 , y3794 , y3795 , y3796 , y3797 , y3798 , y3799 , y3800 , y3801 , y3802 , y3803 , y3804 , y3805 , y3806 , y3807 , y3808 , y3809 , y3810 , y3811 , y3812 , y3813 , y3814 , y3815 , y3816 , y3817 , y3818 , y3819 , y3820 , y3821 , y3822 , y3823 , y3824 , y3825 , y3826 , y3827 , y3828 , y3829 , y3830 , y3831 , y3832 , y3833 , y3834 , y3835 , y3836 , y3837 , y3838 , y3839 , y3840 , y3841 , y3842 , y3843 , y3844 , y3845 , y3846 , y3847 , y3848 , y3849 , y3850 , y3851 , y3852 , y3853 , y3854 , y3855 , y3856 , y3857 , y3858 , y3859 , y3860 , y3861 , y3862 , y3863 , y3864 , y3865 , y3866 , y3867 , y3868 , y3869 , y3870 , y3871 , y3872 , y3873 , y3874 , y3875 , y3876 , y3877 , y3878 , y3879 , y3880 , y3881 , y3882 , y3883 , y3884 , y3885 , y3886 , y3887 , y3888 , y3889 , y3890 , y3891 , y3892 , y3893 , y3894 , y3895 , y3896 , y3897 , y3898 , y3899 , y3900 , y3901 , y3902 , y3903 , y3904 , y3905 , y3906 , y3907 , y3908 , y3909 , y3910 , y3911 , y3912 , y3913 , y3914 , y3915 , y3916 , y3917 , y3918 , y3919 , y3920 , y3921 , y3922 , y3923 , y3924 , y3925 , y3926 , y3927 , y3928 , y3929 , y3930 , y3931 , y3932 , y3933 , y3934 , y3935 , y3936 , y3937 , y3938 , y3939 , y3940 , y3941 , y3942 , y3943 , y3944 , y3945 , y3946 , y3947 , y3948 , y3949 , y3950 , y3951 , y3952 , y3953 , y3954 , y3955 , y3956 , y3957 , y3958 , y3959 , y3960 , y3961 , y3962 , y3963 , y3964 , y3965 , y3966 , y3967 , y3968 , y3969 , y3970 , y3971 , y3972 , y3973 , y3974 , y3975 , y3976 , y3977 , y3978 , y3979 , y3980 , y3981 , y3982 , y3983 , y3984 , y3985 , y3986 , y3987 , y3988 , y3989 , y3990 , y3991 , y3992 , y3993 , y3994 , y3995 , y3996 , y3997 , y3998 , y3999 , y4000 , y4001 , y4002 , y4003 , y4004 , y4005 , y4006 , y4007 , y4008 , y4009 , y4010 , y4011 , y4012 , y4013 , y4014 , y4015 , y4016 , y4017 , y4018 , y4019 , y4020 , y4021 , y4022 , y4023 , y4024 , y4025 , y4026 , y4027 , y4028 , y4029 , y4030 , y4031 , y4032 , y4033 , y4034 , y4035 , y4036 , y4037 , y4038 , y4039 , y4040 , y4041 , y4042 , y4043 , y4044 , y4045 , y4046 , y4047 , y4048 , y4049 , y4050 , y4051 , y4052 , y4053 , y4054 , y4055 , y4056 , y4057 , y4058 , y4059 , y4060 , y4061 , y4062 , y4063 , y4064 , y4065 , y4066 , y4067 , y4068 , y4069 , y4070 , y4071 , y4072 , y4073 , y4074 , y4075 , y4076 , y4077 , y4078 , y4079 , y4080 , y4081 , y4082 , y4083 , y4084 , y4085 , y4086 , y4087 , y4088 , y4089 , y4090 , y4091 , y4092 , y4093 , y4094 , y4095 , y4096 , y4097 , y4098 , y4099 , y4100 , y4101 , y4102 , y4103 , y4104 , y4105 , y4106 , y4107 , y4108 , y4109 , y4110 , y4111 , y4112 , y4113 , y4114 , y4115 , y4116 , y4117 , y4118 , y4119 , y4120 , y4121 , y4122 , y4123 , y4124 , y4125 , y4126 , y4127 , y4128 , y4129 , y4130 , y4131 , y4132 , y4133 , y4134 , y4135 , y4136 , y4137 , y4138 , y4139 , y4140 , y4141 , y4142 , y4143 , y4144 , y4145 , y4146 , y4147 , y4148 , y4149 , y4150 , y4151 , y4152 , y4153 , y4154 , y4155 , y4156 , y4157 , y4158 , y4159 , y4160 , y4161 , y4162 , y4163 , y4164 , y4165 , y4166 , y4167 , y4168 , y4169 , y4170 , y4171 , y4172 , y4173 , y4174 , y4175 , y4176 , y4177 , y4178 , y4179 , y4180 , y4181 , y4182 , y4183 , y4184 , y4185 , y4186 , y4187 , y4188 , y4189 , y4190 , y4191 , y4192 , y4193 , y4194 , y4195 , y4196 , y4197 , y4198 , y4199 , y4200 , y4201 , y4202 , y4203 , y4204 , y4205 , y4206 , y4207 , y4208 , y4209 , y4210 , y4211 , y4212 , y4213 , y4214 , y4215 , y4216 , y4217 , y4218 , y4219 , y4220 , y4221 , y4222 , y4223 , y4224 , y4225 , y4226 , y4227 , y4228 , y4229 , y4230 , y4231 , y4232 , y4233 , y4234 , y4235 , y4236 , y4237 , y4238 , y4239 , y4240 , y4241 , y4242 , y4243 , y4244 , y4245 , y4246 , y4247 , y4248 , y4249 , y4250 , y4251 , y4252 , y4253 , y4254 , y4255 , y4256 , y4257 , y4258 , y4259 , y4260 , y4261 , y4262 , y4263 , y4264 , y4265 , y4266 , y4267 , y4268 , y4269 , y4270 , y4271 , y4272 , y4273 , y4274 , y4275 , y4276 , y4277 , y4278 , y4279 , y4280 , y4281 , y4282 , y4283 , y4284 , y4285 , y4286 , y4287 , y4288 , y4289 , y4290 , y4291 , y4292 , y4293 , y4294 , y4295 , y4296 , y4297 , y4298 , y4299 , y4300 , y4301 , y4302 , y4303 , y4304 , y4305 , y4306 , y4307 , y4308 , y4309 , y4310 , y4311 , y4312 , y4313 , y4314 , y4315 , y4316 , y4317 , y4318 , y4319 , y4320 , y4321 , y4322 , y4323 , y4324 , y4325 , y4326 , y4327 , y4328 , y4329 , y4330 , y4331 , y4332 , y4333 , y4334 , y4335 , y4336 , y4337 , y4338 , y4339 , y4340 , y4341 , y4342 , y4343 , y4344 , y4345 , y4346 , y4347 , y4348 , y4349 , y4350 , y4351 , y4352 , y4353 , y4354 , y4355 , y4356 , y4357 , y4358 , y4359 , y4360 , y4361 , y4362 , y4363 , y4364 , y4365 , y4366 , y4367 , y4368 , y4369 , y4370 , y4371 , y4372 , y4373 , y4374 , y4375 , y4376 , y4377 , y4378 , y4379 , y4380 , y4381 , y4382 , y4383 , y4384 , y4385 , y4386 , y4387 , y4388 , y4389 , y4390 , y4391 , y4392 , y4393 , y4394 , y4395 , y4396 , y4397 , y4398 , y4399 , y4400 , y4401 , y4402 , y4403 , y4404 , y4405 , y4406 , y4407 , y4408 , y4409 , y4410 , y4411 , y4412 , y4413 , y4414 , y4415 , y4416 , y4417 , y4418 , y4419 , y4420 , y4421 , y4422 , y4423 , y4424 , y4425 , y4426 , y4427 , y4428 , y4429 , y4430 , y4431 , y4432 , y4433 , y4434 , y4435 , y4436 , y4437 , y4438 , y4439 , y4440 , y4441 , y4442 , y4443 , y4444 , y4445 , y4446 , y4447 , y4448 , y4449 , y4450 , y4451 , y4452 , y4453 , y4454 , y4455 , y4456 , y4457 , y4458 , y4459 , y4460 , y4461 , y4462 , y4463 , y4464 , y4465 , y4466 , y4467 , y4468 , y4469 , y4470 , y4471 , y4472 , y4473 , y4474 , y4475 , y4476 , y4477 , y4478 , y4479 , y4480 , y4481 , y4482 , y4483 , y4484 , y4485 , y4486 , y4487 , y4488 , y4489 , y4490 , y4491 , y4492 , y4493 , y4494 , y4495 , y4496 , y4497 , y4498 , y4499 , y4500 , y4501 , y4502 , y4503 , y4504 , y4505 , y4506 , y4507 , y4508 , y4509 , y4510 , y4511 , y4512 , y4513 , y4514 , y4515 , y4516 , y4517 , y4518 , y4519 , y4520 , y4521 , y4522 , y4523 , y4524 , y4525 , y4526 , y4527 , y4528 , y4529 , y4530 , y4531 , y4532 , y4533 , y4534 , y4535 , y4536 , y4537 , y4538 , y4539 , y4540 , y4541 , y4542 , y4543 , y4544 , y4545 , y4546 , y4547 , y4548 , y4549 , y4550 , y4551 , y4552 , y4553 , y4554 , y4555 , y4556 , y4557 , y4558 , y4559 , y4560 , y4561 , y4562 , y4563 , y4564 , y4565 , y4566 , y4567 , y4568 , y4569 , y4570 , y4571 , y4572 , y4573 , y4574 , y4575 , y4576 , y4577 , y4578 , y4579 , y4580 , y4581 , y4582 , y4583 , y4584 , y4585 , y4586 , y4587 , y4588 , y4589 , y4590 , y4591 , y4592 , y4593 , y4594 , y4595 , y4596 , y4597 , y4598 , y4599 , y4600 , y4601 , y4602 , y4603 , y4604 , y4605 , y4606 , y4607 , y4608 , y4609 , y4610 , y4611 , y4612 , y4613 , y4614 , y4615 , y4616 , y4617 , y4618 , y4619 , y4620 , y4621 , y4622 , y4623 , y4624 , y4625 , y4626 , y4627 , y4628 , y4629 , y4630 , y4631 , y4632 , y4633 , y4634 , y4635 , y4636 , y4637 , y4638 , y4639 , y4640 , y4641 , y4642 , y4643 , y4644 , y4645 , y4646 , y4647 , y4648 , y4649 , y4650 , y4651 , y4652 , y4653 , y4654 , y4655 , y4656 , y4657 , y4658 , y4659 , y4660 , y4661 , y4662 , y4663 , y4664 , y4665 , y4666 , y4667 , y4668 , y4669 , y4670 , y4671 , y4672 , y4673 , y4674 , y4675 , y4676 , y4677 , y4678 , y4679 , y4680 , y4681 , y4682 , y4683 , y4684 , y4685 , y4686 , y4687 , y4688 , y4689 , y4690 , y4691 , y4692 , y4693 , y4694 , y4695 , y4696 , y4697 , y4698 , y4699 , y4700 , y4701 , y4702 , y4703 , y4704 , y4705 , y4706 , y4707 , y4708 , y4709 , y4710 , y4711 , y4712 , y4713 , y4714 , y4715 , y4716 , y4717 , y4718 , y4719 , y4720 , y4721 , y4722 , y4723 , y4724 , y4725 , y4726 , y4727 , y4728 , y4729 , y4730 , y4731 , y4732 , y4733 , y4734 , y4735 , y4736 , y4737 , y4738 , y4739 , y4740 , y4741 , y4742 , y4743 , y4744 , y4745 , y4746 , y4747 , y4748 , y4749 , y4750 , y4751 , y4752 , y4753 , y4754 , y4755 , y4756 , y4757 , y4758 , y4759 , y4760 , y4761 , y4762 , y4763 , y4764 , y4765 , y4766 , y4767 , y4768 , y4769 , y4770 , y4771 , y4772 , y4773 , y4774 , y4775 , y4776 , y4777 , y4778 , y4779 , y4780 , y4781 , y4782 , y4783 , y4784 , y4785 , y4786 , y4787 , y4788 , y4789 , y4790 , y4791 , y4792 , y4793 , y4794 , y4795 , y4796 , y4797 , y4798 , y4799 , y4800 , y4801 , y4802 , y4803 , y4804 , y4805 , y4806 , y4807 , y4808 , y4809 , y4810 , y4811 , y4812 , y4813 , y4814 , y4815 , y4816 , y4817 , y4818 , y4819 , y4820 , y4821 , y4822 , y4823 , y4824 , y4825 , y4826 , y4827 , y4828 , y4829 , y4830 , y4831 , y4832 , y4833 , y4834 , y4835 , y4836 , y4837 , y4838 , y4839 , y4840 , y4841 , y4842 , y4843 , y4844 , y4845 , y4846 , y4847 , y4848 , y4849 , y4850 , y4851 , y4852 , y4853 , y4854 , y4855 , y4856 , y4857 , y4858 , y4859 , y4860 , y4861 , y4862 , y4863 , y4864 , y4865 , y4866 , y4867 , y4868 , y4869 , y4870 , y4871 , y4872 , y4873 , y4874 , y4875 , y4876 , y4877 , y4878 , y4879 , y4880 , y4881 , y4882 , y4883 , y4884 , y4885 , y4886 , y4887 , y4888 , y4889 , y4890 , y4891 , y4892 , y4893 , y4894 , y4895 , y4896 , y4897 , y4898 , y4899 , y4900 , y4901 , y4902 , y4903 , y4904 , y4905 , y4906 , y4907 , y4908 , y4909 , y4910 , y4911 , y4912 , y4913 , y4914 , y4915 , y4916 , y4917 , y4918 , y4919 , y4920 , y4921 , y4922 , y4923 , y4924 , y4925 , y4926 , y4927 , y4928 , y4929 , y4930 , y4931 , y4932 , y4933 , y4934 , y4935 , y4936 , y4937 , y4938 , y4939 , y4940 , y4941 , y4942 , y4943 , y4944 , y4945 , y4946 , y4947 , y4948 , y4949 , y4950 , y4951 , y4952 , y4953 , y4954 , y4955 , y4956 , y4957 , y4958 , y4959 , y4960 , y4961 , y4962 , y4963 , y4964 , y4965 , y4966 , y4967 , y4968 , y4969 , y4970 , y4971 , y4972 , y4973 , y4974 , y4975 , y4976 , y4977 , y4978 , y4979 , y4980 , y4981 , y4982 , y4983 , y4984 , y4985 , y4986 , y4987 , y4988 , y4989 , y4990 , y4991 , y4992 , y4993 , y4994 , y4995 , y4996 , y4997 , y4998 , y4999 , y5000 , y5001 , y5002 , y5003 , y5004 , y5005 , y5006 , y5007 , y5008 , y5009 , y5010 , y5011 , y5012 , y5013 , y5014 , y5015 , y5016 , y5017 , y5018 , y5019 , y5020 , y5021 , y5022 , y5023 , y5024 , y5025 , y5026 , y5027 , y5028 , y5029 , y5030 , y5031 , y5032 , y5033 , y5034 , y5035 , y5036 , y5037 , y5038 , y5039 , y5040 , y5041 , y5042 , y5043 , y5044 , y5045 , y5046 , y5047 , y5048 , y5049 , y5050 , y5051 , y5052 , y5053 , y5054 , y5055 , y5056 , y5057 , y5058 , y5059 , y5060 , y5061 , y5062 , y5063 , y5064 , y5065 , y5066 , y5067 , y5068 , y5069 , y5070 , y5071 , y5072 , y5073 , y5074 , y5075 , y5076 , y5077 , y5078 , y5079 , y5080 , y5081 , y5082 , y5083 , y5084 , y5085 , y5086 , y5087 , y5088 , y5089 , y5090 , y5091 , y5092 , y5093 , y5094 , y5095 , y5096 , y5097 , y5098 , y5099 , y5100 , y5101 , y5102 , y5103 , y5104 , y5105 , y5106 , y5107 , y5108 , y5109 , y5110 , y5111 , y5112 , y5113 , y5114 , y5115 , y5116 , y5117 , y5118 , y5119 , y5120 , y5121 , y5122 , y5123 , y5124 , y5125 , y5126 , y5127 , y5128 , y5129 , y5130 , y5131 , y5132 , y5133 , y5134 , y5135 , y5136 , y5137 , y5138 , y5139 , y5140 , y5141 , y5142 , y5143 , y5144 , y5145 , y5146 , y5147 , y5148 , y5149 , y5150 , y5151 , y5152 , y5153 , y5154 , y5155 , y5156 , y5157 , y5158 , y5159 , y5160 , y5161 , y5162 , y5163 , y5164 , y5165 , y5166 , y5167 , y5168 , y5169 , y5170 , y5171 , y5172 , y5173 , y5174 , y5175 , y5176 , y5177 , y5178 , y5179 , y5180 , y5181 , y5182 , y5183 , y5184 , y5185 , y5186 , y5187 , y5188 , y5189 , y5190 , y5191 , y5192 , y5193 , y5194 , y5195 , y5196 , y5197 , y5198 , y5199 , y5200 , y5201 , y5202 , y5203 , y5204 , y5205 , y5206 , y5207 , y5208 , y5209 , y5210 , y5211 , y5212 , y5213 , y5214 , y5215 , y5216 , y5217 , y5218 , y5219 , y5220 , y5221 , y5222 , y5223 , y5224 , y5225 , y5226 , y5227 , y5228 , y5229 , y5230 , y5231 , y5232 , y5233 , y5234 , y5235 , y5236 , y5237 , y5238 , y5239 , y5240 , y5241 , y5242 , y5243 , y5244 , y5245 , y5246 , y5247 , y5248 , y5249 , y5250 , y5251 , y5252 , y5253 , y5254 , y5255 , y5256 , y5257 , y5258 , y5259 , y5260 , y5261 , y5262 , y5263 , y5264 , y5265 , y5266 , y5267 , y5268 , y5269 , y5270 , y5271 , y5272 , y5273 , y5274 , y5275 , y5276 , y5277 , y5278 , y5279 , y5280 , y5281 , y5282 , y5283 , y5284 , y5285 , y5286 , y5287 , y5288 , y5289 , y5290 , y5291 , y5292 , y5293 , y5294 , y5295 , y5296 , y5297 , y5298 , y5299 , y5300 , y5301 , y5302 , y5303 , y5304 , y5305 , y5306 , y5307 , y5308 , y5309 , y5310 , y5311 , y5312 , y5313 , y5314 , y5315 , y5316 , y5317 , y5318 , y5319 , y5320 , y5321 , y5322 , y5323 , y5324 , y5325 , y5326 , y5327 , y5328 , y5329 , y5330 , y5331 , y5332 , y5333 , y5334 , y5335 , y5336 , y5337 , y5338 , y5339 , y5340 , y5341 , y5342 , y5343 , y5344 , y5345 , y5346 , y5347 , y5348 , y5349 , y5350 , y5351 , y5352 , y5353 , y5354 , y5355 , y5356 , y5357 , y5358 , y5359 , y5360 , y5361 , y5362 , y5363 , y5364 , y5365 , y5366 , y5367 , y5368 , y5369 , y5370 , y5371 , y5372 , y5373 , y5374 , y5375 , y5376 , y5377 , y5378 , y5379 , y5380 , y5381 , y5382 , y5383 , y5384 , y5385 , y5386 , y5387 , y5388 , y5389 , y5390 , y5391 , y5392 , y5393 , y5394 , y5395 , y5396 , y5397 , y5398 , y5399 , y5400 , y5401 , y5402 , y5403 , y5404 , y5405 , y5406 , y5407 , y5408 , y5409 , y5410 , y5411 , y5412 , y5413 , y5414 , y5415 , y5416 , y5417 , y5418 , y5419 , y5420 , y5421 , y5422 , y5423 , y5424 , y5425 , y5426 , y5427 , y5428 , y5429 , y5430 , y5431 , y5432 , y5433 , y5434 , y5435 , y5436 , y5437 , y5438 , y5439 , y5440 , y5441 , y5442 , y5443 , y5444 , y5445 , y5446 , y5447 , y5448 , y5449 , y5450 , y5451 , y5452 , y5453 , y5454 , y5455 , y5456 , y5457 , y5458 , y5459 , y5460 , y5461 , y5462 , y5463 , y5464 , y5465 , y5466 , y5467 , y5468 , y5469 , y5470 , y5471 , y5472 , y5473 , y5474 , y5475 , y5476 , y5477 , y5478 , y5479 , y5480 , y5481 , y5482 , y5483 , y5484 , y5485 , y5486 , y5487 , y5488 , y5489 , y5490 , y5491 , y5492 , y5493 , y5494 , y5495 , y5496 , y5497 , y5498 , y5499 , y5500 , y5501 , y5502 , y5503 , y5504 , y5505 , y5506 , y5507 , y5508 , y5509 , y5510 , y5511 , y5512 , y5513 , y5514 , y5515 , y5516 , y5517 , y5518 , y5519 , y5520 , y5521 , y5522 , y5523 , y5524 , y5525 , y5526 , y5527 , y5528 , y5529 , y5530 , y5531 , y5532 , y5533 , y5534 , y5535 , y5536 , y5537 , y5538 , y5539 , y5540 , y5541 , y5542 , y5543 , y5544 , y5545 , y5546 , y5547 , y5548 , y5549 , y5550 , y5551 , y5552 , y5553 , y5554 , y5555 , y5556 , y5557 , y5558 , y5559 , y5560 , y5561 , y5562 , y5563 , y5564 , y5565 , y5566 , y5567 , y5568 , y5569 , y5570 , y5571 , y5572 , y5573 , y5574 , y5575 , y5576 , y5577 , y5578 , y5579 , y5580 , y5581 , y5582 , y5583 , y5584 , y5585 , y5586 , y5587 , y5588 , y5589 , y5590 , y5591 , y5592 , y5593 , y5594 , y5595 , y5596 , y5597 , y5598 , y5599 , y5600 , y5601 , y5602 , y5603 , y5604 , y5605 , y5606 , y5607 , y5608 , y5609 , y5610 , y5611 , y5612 , y5613 , y5614 , y5615 , y5616 , y5617 , y5618 , y5619 , y5620 , y5621 , y5622 , y5623 , y5624 , y5625 , y5626 , y5627 , y5628 , y5629 , y5630 , y5631 , y5632 , y5633 , y5634 , y5635 , y5636 , y5637 , y5638 , y5639 , y5640 , y5641 , y5642 , y5643 , y5644 , y5645 , y5646 , y5647 , y5648 , y5649 , y5650 , y5651 , y5652 , y5653 , y5654 , y5655 , y5656 , y5657 , y5658 , y5659 , y5660 , y5661 , y5662 , y5663 , y5664 , y5665 , y5666 , y5667 , y5668 , y5669 , y5670 , y5671 , y5672 , y5673 , y5674 , y5675 , y5676 , y5677 , y5678 , y5679 , y5680 , y5681 , y5682 , y5683 , y5684 , y5685 , y5686 , y5687 , y5688 , y5689 , y5690 , y5691 , y5692 , y5693 , y5694 , y5695 , y5696 , y5697 , y5698 , y5699 , y5700 , y5701 , y5702 , y5703 , y5704 , y5705 , y5706 , y5707 , y5708 , y5709 , y5710 , y5711 , y5712 , y5713 , y5714 , y5715 , y5716 , y5717 , y5718 , y5719 , y5720 , y5721 , y5722 , y5723 , y5724 , y5725 , y5726 , y5727 , y5728 , y5729 , y5730 , y5731 , y5732 , y5733 , y5734 , y5735 , y5736 , y5737 , y5738 , y5739 , y5740 , y5741 , y5742 , y5743 , y5744 , y5745 , y5746 , y5747 , y5748 , y5749 , y5750 , y5751 , y5752 , y5753 , y5754 , y5755 , y5756 , y5757 , y5758 , y5759 , y5760 , y5761 , y5762 , y5763 , y5764 , y5765 , y5766 , y5767 , y5768 , y5769 , y5770 , y5771 , y5772 , y5773 , y5774 , y5775 , y5776 , y5777 , y5778 , y5779 , y5780 , y5781 , y5782 , y5783 , y5784 , y5785 , y5786 , y5787 , y5788 , y5789 , y5790 , y5791 , y5792 , y5793 , y5794 , y5795 , y5796 , y5797 , y5798 , y5799 , y5800 , y5801 , y5802 , y5803 , y5804 , y5805 , y5806 , y5807 , y5808 , y5809 , y5810 , y5811 , y5812 , y5813 , y5814 , y5815 , y5816 , y5817 , y5818 , y5819 , y5820 , y5821 , y5822 , y5823 , y5824 , y5825 , y5826 , y5827 , y5828 , y5829 , y5830 , y5831 , y5832 , y5833 , y5834 , y5835 , y5836 , y5837 , y5838 , y5839 , y5840 , y5841 , y5842 , y5843 , y5844 , y5845 , y5846 , y5847 , y5848 , y5849 , y5850 , y5851 , y5852 , y5853 , y5854 , y5855 , y5856 , y5857 , y5858 , y5859 , y5860 , y5861 , y5862 , y5863 , y5864 , y5865 , y5866 , y5867 , y5868 , y5869 , y5870 , y5871 , y5872 , y5873 , y5874 , y5875 , y5876 , y5877 , y5878 , y5879 , y5880 , y5881 , y5882 , y5883 , y5884 , y5885 , y5886 , y5887 , y5888 , y5889 , y5890 , y5891 , y5892 , y5893 , y5894 , y5895 , y5896 , y5897 , y5898 , y5899 , y5900 , y5901 , y5902 , y5903 , y5904 , y5905 , y5906 , y5907 , y5908 , y5909 , y5910 , y5911 , y5912 , y5913 , y5914 , y5915 , y5916 , y5917 , y5918 , y5919 , y5920 , y5921 , y5922 , y5923 , y5924 , y5925 , y5926 , y5927 , y5928 , y5929 , y5930 , y5931 , y5932 , y5933 , y5934 , y5935 , y5936 , y5937 , y5938 , y5939 , y5940 , y5941 , y5942 , y5943 , y5944 , y5945 , y5946 , y5947 , y5948 , y5949 , y5950 , y5951 , y5952 , y5953 , y5954 , y5955 , y5956 , y5957 , y5958 , y5959 , y5960 , y5961 , y5962 , y5963 , y5964 , y5965 , y5966 , y5967 , y5968 , y5969 , y5970 , y5971 , y5972 , y5973 , y5974 , y5975 , y5976 , y5977 , y5978 , y5979 , y5980 , y5981 , y5982 , y5983 , y5984 , y5985 , y5986 , y5987 , y5988 , y5989 , y5990 , y5991 , y5992 , y5993 , y5994 , y5995 , y5996 , y5997 , y5998 , y5999 , y6000 , y6001 , y6002 , y6003 , y6004 , y6005 , y6006 , y6007 , y6008 , y6009 , y6010 , y6011 , y6012 , y6013 , y6014 , y6015 , y6016 , y6017 , y6018 , y6019 , y6020 , y6021 , y6022 , y6023 , y6024 , y6025 , y6026 , y6027 , y6028 , y6029 , y6030 , y6031 , y6032 , y6033 , y6034 , y6035 , y6036 , y6037 , y6038 , y6039 , y6040 , y6041 , y6042 , y6043 , y6044 , y6045 , y6046 , y6047 , y6048 , y6049 , y6050 , y6051 , y6052 , y6053 , y6054 , y6055 , y6056 , y6057 , y6058 , y6059 , y6060 , y6061 , y6062 , y6063 , y6064 , y6065 , y6066 , y6067 , y6068 , y6069 , y6070 , y6071 , y6072 , y6073 , y6074 , y6075 , y6076 , y6077 , y6078 , y6079 , y6080 , y6081 , y6082 , y6083 , y6084 , y6085 , y6086 , y6087 , y6088 , y6089 , y6090 , y6091 , y6092 , y6093 , y6094 , y6095 , y6096 , y6097 , y6098 , y6099 , y6100 , y6101 , y6102 , y6103 , y6104 , y6105 , y6106 , y6107 , y6108 , y6109 , y6110 , y6111 , y6112 , y6113 , y6114 , y6115 , y6116 , y6117 , y6118 , y6119 , y6120 , y6121 , y6122 , y6123 , y6124 , y6125 , y6126 , y6127 , y6128 , y6129 , y6130 , y6131 , y6132 , y6133 , y6134 , y6135 , y6136 , y6137 , y6138 , y6139 , y6140 , y6141 , y6142 , y6143 , y6144 , y6145 , y6146 , y6147 , y6148 , y6149 , y6150 , y6151 , y6152 , y6153 , y6154 , y6155 , y6156 , y6157 , y6158 , y6159 , y6160 , y6161 , y6162 , y6163 , y6164 , y6165 , y6166 , y6167 , y6168 , y6169 , y6170 , y6171 , y6172 , y6173 , y6174 , y6175 , y6176 , y6177 , y6178 , y6179 , y6180 , y6181 , y6182 , y6183 , y6184 , y6185 , y6186 , y6187 , y6188 , y6189 , y6190 , y6191 , y6192 , y6193 , y6194 , y6195 , y6196 , y6197 , y6198 , y6199 , y6200 , y6201 , y6202 , y6203 , y6204 , y6205 , y6206 , y6207 , y6208 , y6209 , y6210 , y6211 , y6212 , y6213 , y6214 , y6215 , y6216 , y6217 , y6218 , y6219 , y6220 , y6221 , y6222 , y6223 , y6224 , y6225 , y6226 , y6227 , y6228 , y6229 , y6230 , y6231 , y6232 , y6233 , y6234 , y6235 , y6236 , y6237 , y6238 , y6239 , y6240 , y6241 , y6242 , y6243 , y6244 , y6245 , y6246 , y6247 , y6248 , y6249 , y6250 , y6251 , y6252 , y6253 , y6254 , y6255 , y6256 , y6257 , y6258 , y6259 , y6260 , y6261 , y6262 , y6263 , y6264 , y6265 , y6266 , y6267 , y6268 , y6269 , y6270 , y6271 , y6272 , y6273 , y6274 , y6275 , y6276 , y6277 , y6278 , y6279 , y6280 , y6281 , y6282 , y6283 , y6284 , y6285 , y6286 , y6287 , y6288 , y6289 , y6290 , y6291 , y6292 , y6293 , y6294 , y6295 , y6296 , y6297 , y6298 , y6299 , y6300 , y6301 , y6302 , y6303 , y6304 , y6305 , y6306 , y6307 , y6308 , y6309 , y6310 , y6311 , y6312 , y6313 , y6314 , y6315 , y6316 , y6317 , y6318 , y6319 , y6320 , y6321 , y6322 , y6323 , y6324 , y6325 , y6326 , y6327 , y6328 , y6329 , y6330 , y6331 , y6332 , y6333 , y6334 , y6335 , y6336 , y6337 , y6338 , y6339 , y6340 , y6341 , y6342 , y6343 , y6344 , y6345 , y6346 , y6347 , y6348 , y6349 , y6350 , y6351 , y6352 , y6353 , y6354 , y6355 , y6356 , y6357 , y6358 , y6359 , y6360 , y6361 , y6362 , y6363 , y6364 , y6365 , y6366 , y6367 , y6368 , y6369 , y6370 , y6371 , y6372 , y6373 , y6374 , y6375 , y6376 , y6377 , y6378 , y6379 , y6380 , y6381 , y6382 , y6383 , y6384 , y6385 , y6386 , y6387 , y6388 , y6389 , y6390 , y6391 , y6392 , y6393 , y6394 , y6395 , y6396 , y6397 , y6398 , y6399 , y6400 , y6401 , y6402 , y6403 , y6404 , y6405 , y6406 , y6407 , y6408 , y6409 , y6410 , y6411 , y6412 , y6413 , y6414 , y6415 , y6416 , y6417 , y6418 , y6419 , y6420 , y6421 , y6422 , y6423 , y6424 , y6425 , y6426 , y6427 , y6428 , y6429 , y6430 , y6431 , y6432 , y6433 , y6434 , y6435 , y6436 , y6437 , y6438 , y6439 , y6440 , y6441 , y6442 , y6443 , y6444 , y6445 , y6446 , y6447 , y6448 , y6449 , y6450 , y6451 , y6452 , y6453 , y6454 , y6455 , y6456 , y6457 , y6458 , y6459 , y6460 , y6461 , y6462 , y6463 , y6464 , y6465 , y6466 , y6467 , y6468 , y6469 , y6470 , y6471 , y6472 , y6473 , y6474 , y6475 , y6476 , y6477 , y6478 , y6479 , y6480 , y6481 , y6482 , y6483 , y6484 , y6485 , y6486 , y6487 , y6488 , y6489 , y6490 , y6491 , y6492 , y6493 , y6494 , y6495 , y6496 , y6497 , y6498 , y6499 , y6500 , y6501 , y6502 , y6503 , y6504 , y6505 , y6506 , y6507 , y6508 , y6509 , y6510 , y6511 , y6512 , y6513 , y6514 , y6515 , y6516 , y6517 , y6518 , y6519 , y6520 , y6521 , y6522 , y6523 , y6524 , y6525 , y6526 , y6527 , y6528 , y6529 , y6530 , y6531 , y6532 , y6533 , y6534 , y6535 , y6536 , y6537 , y6538 , y6539 , y6540 , y6541 , y6542 , y6543 , y6544 , y6545 , y6546 , y6547 , y6548 , y6549 , y6550 , y6551 , y6552 , y6553 , y6554 , y6555 , y6556 , y6557 , y6558 , y6559 , y6560 , y6561 , y6562 , y6563 , y6564 , y6565 , y6566 , y6567 , y6568 , y6569 , y6570 , y6571 , y6572 , y6573 , y6574 , y6575 , y6576 , y6577 , y6578 , y6579 , y6580 , y6581 , y6582 , y6583 , y6584 , y6585 , y6586 , y6587 , y6588 , y6589 , y6590 , y6591 , y6592 , y6593 , y6594 , y6595 , y6596 , y6597 , y6598 , y6599 , y6600 , y6601 , y6602 , y6603 , y6604 , y6605 , y6606 , y6607 , y6608 , y6609 , y6610 , y6611 , y6612 , y6613 , y6614 , y6615 , y6616 , y6617 , y6618 , y6619 , y6620 , y6621 , y6622 , y6623 , y6624 , y6625 , y6626 , y6627 , y6628 , y6629 , y6630 , y6631 , y6632 , y6633 , y6634 , y6635 , y6636 , y6637 , y6638 , y6639 , y6640 , y6641 , y6642 , y6643 , y6644 , y6645 , y6646 , y6647 , y6648 , y6649 , y6650 , y6651 , y6652 , y6653 , y6654 , y6655 , y6656 , y6657 , y6658 , y6659 , y6660 , y6661 , y6662 , y6663 , y6664 , y6665 , y6666 , y6667 , y6668 , y6669 , y6670 , y6671 , y6672 , y6673 , y6674 , y6675 , y6676 , y6677 , y6678 , y6679 , y6680 , y6681 , y6682 , y6683 , y6684 , y6685 , y6686 , y6687 , y6688 , y6689 , y6690 , y6691 , y6692 , y6693 , y6694 , y6695 , y6696 , y6697 , y6698 , y6699 , y6700 , y6701 , y6702 , y6703 , y6704 , y6705 , y6706 , y6707 , y6708 , y6709 , y6710 , y6711 , y6712 , y6713 , y6714 , y6715 , y6716 , y6717 , y6718 , y6719 , y6720 , y6721 , y6722 , y6723 , y6724 , y6725 , y6726 , y6727 , y6728 , y6729 , y6730 , y6731 , y6732 , y6733 , y6734 , y6735 , y6736 , y6737 , y6738 , y6739 , y6740 , y6741 , y6742 , y6743 , y6744 , y6745 , y6746 , y6747 , y6748 , y6749 , y6750 , y6751 , y6752 , y6753 , y6754 , y6755 , y6756 , y6757 , y6758 , y6759 , y6760 , y6761 , y6762 , y6763 , y6764 , y6765 , y6766 , y6767 , y6768 , y6769 , y6770 , y6771 , y6772 , y6773 , y6774 , y6775 , y6776 , y6777 , y6778 , y6779 , y6780 , y6781 , y6782 , y6783 , y6784 , y6785 , y6786 , y6787 , y6788 , y6789 , y6790 , y6791 , y6792 , y6793 , y6794 , y6795 , y6796 , y6797 , y6798 , y6799 , y6800 , y6801 , y6802 , y6803 , y6804 , y6805 , y6806 , y6807 , y6808 , y6809 , y6810 , y6811 , y6812 , y6813 , y6814 , y6815 , y6816 , y6817 , y6818 , y6819 , y6820 , y6821 , y6822 , y6823 , y6824 , y6825 , y6826 , y6827 , y6828 , y6829 , y6830 , y6831 , y6832 , y6833 , y6834 , y6835 , y6836 , y6837 , y6838 , y6839 , y6840 , y6841 , y6842 , y6843 , y6844 , y6845 , y6846 , y6847 , y6848 , y6849 , y6850 , y6851 , y6852 , y6853 , y6854 , y6855 , y6856 , y6857 , y6858 , y6859 , y6860 , y6861 , y6862 , y6863 , y6864 , y6865 , y6866 , y6867 , y6868 , y6869 , y6870 , y6871 , y6872 , y6873 , y6874 , y6875 , y6876 , y6877 , y6878 , y6879 , y6880 , y6881 , y6882 , y6883 , y6884 , y6885 , y6886 , y6887 , y6888 , y6889 , y6890 , y6891 , y6892 , y6893 , y6894 , y6895 , y6896 , y6897 , y6898 , y6899 , y6900 , y6901 , y6902 , y6903 , y6904 , y6905 , y6906 , y6907 , y6908 , y6909 , y6910 , y6911 , y6912 , y6913 , y6914 , y6915 , y6916 , y6917 , y6918 , y6919 , y6920 , y6921 , y6922 , y6923 , y6924 , y6925 , y6926 , y6927 , y6928 , y6929 , y6930 , y6931 , y6932 , y6933 , y6934 , y6935 , y6936 , y6937 , y6938 , y6939 , y6940 , y6941 , y6942 , y6943 , y6944 , y6945 , y6946 , y6947 , y6948 , y6949 , y6950 , y6951 , y6952 , y6953 , y6954 , y6955 , y6956 , y6957 , y6958 , y6959 , y6960 , y6961 , y6962 , y6963 , y6964 , y6965 , y6966 , y6967 , y6968 , y6969 , y6970 , y6971 , y6972 , y6973 , y6974 , y6975 , y6976 , y6977 , y6978 , y6979 , y6980 , y6981 , y6982 , y6983 , y6984 , y6985 , y6986 , y6987 , y6988 , y6989 , y6990 , y6991 , y6992 , y6993 , y6994 , y6995 , y6996 , y6997 , y6998 , y6999 , y7000 , y7001 , y7002 , y7003 , y7004 , y7005 , y7006 , y7007 , y7008 , y7009 , y7010 , y7011 , y7012 , y7013 , y7014 , y7015 , y7016 , y7017 , y7018 , y7019 , y7020 , y7021 , y7022 , y7023 , y7024 , y7025 , y7026 , y7027 , y7028 , y7029 , y7030 , y7031 , y7032 , y7033 , y7034 , y7035 , y7036 , y7037 , y7038 , y7039 , y7040 , y7041 , y7042 , y7043 , y7044 , y7045 , y7046 , y7047 , y7048 , y7049 , y7050 , y7051 , y7052 , y7053 , y7054 , y7055 , y7056 , y7057 , y7058 , y7059 , y7060 , y7061 , y7062 , y7063 , y7064 , y7065 , y7066 , y7067 , y7068 , y7069 , y7070 , y7071 , y7072 , y7073 , y7074 , y7075 , y7076 , y7077 , y7078 , y7079 , y7080 , y7081 , y7082 , y7083 , y7084 , y7085 , y7086 , y7087 , y7088 , y7089 , y7090 , y7091 , y7092 , y7093 , y7094 , y7095 , y7096 , y7097 , y7098 , y7099 , y7100 , y7101 , y7102 , y7103 , y7104 , y7105 , y7106 , y7107 , y7108 , y7109 , y7110 , y7111 , y7112 , y7113 , y7114 , y7115 , y7116 , y7117 , y7118 , y7119 , y7120 , y7121 , y7122 , y7123 , y7124 , y7125 , y7126 , y7127 , y7128 , y7129 , y7130 , y7131 , y7132 , y7133 , y7134 , y7135 , y7136 , y7137 , y7138 , y7139 , y7140 , y7141 , y7142 , y7143 , y7144 , y7145 , y7146 , y7147 , y7148 , y7149 , y7150 , y7151 , y7152 , y7153 , y7154 , y7155 , y7156 , y7157 , y7158 , y7159 , y7160 , y7161 , y7162 , y7163 , y7164 , y7165 , y7166 , y7167 , y7168 , y7169 , y7170 , y7171 , y7172 , y7173 , y7174 , y7175 , y7176 , y7177 , y7178 , y7179 , y7180 , y7181 , y7182 , y7183 , y7184 , y7185 , y7186 , y7187 , y7188 , y7189 , y7190 , y7191 , y7192 , y7193 , y7194 , y7195 , y7196 , y7197 , y7198 , y7199 , y7200 , y7201 , y7202 , y7203 , y7204 , y7205 , y7206 , y7207 , y7208 , y7209 , y7210 , y7211 , y7212 , y7213 , y7214 , y7215 , y7216 , y7217 , y7218 , y7219 , y7220 , y7221 , y7222 , y7223 , y7224 , y7225 , y7226 , y7227 , y7228 , y7229 , y7230 , y7231 , y7232 , y7233 , y7234 , y7235 , y7236 , y7237 , y7238 , y7239 , y7240 , y7241 , y7242 , y7243 , y7244 , y7245 , y7246 , y7247 , y7248 , y7249 , y7250 , y7251 , y7252 , y7253 , y7254 , y7255 , y7256 , y7257 , y7258 , y7259 , y7260 , y7261 , y7262 , y7263 , y7264 , y7265 , y7266 , y7267 , y7268 , y7269 , y7270 , y7271 , y7272 , y7273 , y7274 , y7275 , y7276 , y7277 , y7278 , y7279 , y7280 , y7281 , y7282 , y7283 , y7284 , y7285 , y7286 , y7287 , y7288 , y7289 , y7290 , y7291 , y7292 , y7293 , y7294 , y7295 , y7296 , y7297 , y7298 , y7299 , y7300 , y7301 , y7302 , y7303 , y7304 , y7305 , y7306 , y7307 , y7308 , y7309 , y7310 , y7311 , y7312 , y7313 , y7314 , y7315 , y7316 , y7317 , y7318 , y7319 , y7320 , y7321 , y7322 , y7323 , y7324 , y7325 , y7326 , y7327 , y7328 , y7329 , y7330 , y7331 , y7332 , y7333 , y7334 , y7335 , y7336 , y7337 , y7338 , y7339 , y7340 , y7341 , y7342 , y7343 , y7344 , y7345 , y7346 , y7347 , y7348 , y7349 , y7350 , y7351 , y7352 , y7353 , y7354 , y7355 , y7356 , y7357 , y7358 , y7359 , y7360 , y7361 , y7362 , y7363 , y7364 , y7365 , y7366 , y7367 , y7368 , y7369 , y7370 , y7371 , y7372 , y7373 , y7374 , y7375 , y7376 , y7377 , y7378 , y7379 , y7380 , y7381 , y7382 , y7383 , y7384 , y7385 , y7386 , y7387 , y7388 , y7389 , y7390 , y7391 , y7392 , y7393 , y7394 , y7395 , y7396 , y7397 , y7398 , y7399 , y7400 , y7401 , y7402 , y7403 , y7404 , y7405 , y7406 , y7407 , y7408 , y7409 , y7410 , y7411 , y7412 , y7413 , y7414 , y7415 , y7416 , y7417 , y7418 , y7419 , y7420 , y7421 , y7422 , y7423 , y7424 , y7425 , y7426 , y7427 , y7428 , y7429 , y7430 , y7431 , y7432 , y7433 , y7434 , y7435 , y7436 , y7437 , y7438 , y7439 , y7440 , y7441 , y7442 , y7443 , y7444 , y7445 , y7446 , y7447 , y7448 , y7449 , y7450 , y7451 , y7452 , y7453 , y7454 , y7455 , y7456 , y7457 , y7458 , y7459 , y7460 , y7461 , y7462 , y7463 , y7464 , y7465 , y7466 , y7467 , y7468 , y7469 , y7470 , y7471 , y7472 , y7473 , y7474 , y7475 , y7476 , y7477 , y7478 , y7479 , y7480 , y7481 , y7482 , y7483 , y7484 , y7485 , y7486 , y7487 , y7488 , y7489 , y7490 , y7491 , y7492 , y7493 , y7494 , y7495 , y7496 , y7497 , y7498 , y7499 , y7500 , y7501 , y7502 , y7503 , y7504 , y7505 , y7506 , y7507 , y7508 , y7509 , y7510 , y7511 , y7512 , y7513 , y7514 , y7515 , y7516 , y7517 , y7518 , y7519 , y7520 , y7521 , y7522 , y7523 , y7524 , y7525 , y7526 , y7527 , y7528 , y7529 , y7530 , y7531 , y7532 , y7533 , y7534 , y7535 , y7536 , y7537 , y7538 , y7539 , y7540 , y7541 , y7542 , y7543 , y7544 , y7545 , y7546 , y7547 , y7548 , y7549 , y7550 , y7551 , y7552 , y7553 , y7554 , y7555 , y7556 , y7557 , y7558 , y7559 , y7560 , y7561 , y7562 , y7563 , y7564 , y7565 , y7566 , y7567 , y7568 , y7569 , y7570 , y7571 , y7572 , y7573 , y7574 , y7575 , y7576 , y7577 , y7578 , y7579 , y7580 , y7581 , y7582 , y7583 , y7584 , y7585 , y7586 , y7587 , y7588 , y7589 , y7590 , y7591 , y7592 , y7593 , y7594 , y7595 , y7596 , y7597 , y7598 , y7599 , y7600 , y7601 , y7602 , y7603 , y7604 , y7605 , y7606 , y7607 , y7608 , y7609 , y7610 , y7611 , y7612 , y7613 , y7614 , y7615 , y7616 , y7617 , y7618 , y7619 , y7620 , y7621 , y7622 , y7623 , y7624 , y7625 , y7626 , y7627 , y7628 , y7629 , y7630 , y7631 , y7632 , y7633 , y7634 , y7635 , y7636 , y7637 , y7638 , y7639 , y7640 , y7641 , y7642 , y7643 , y7644 , y7645 , y7646 , y7647 , y7648 , y7649 , y7650 , y7651 , y7652 , y7653 , y7654 , y7655 , y7656 , y7657 , y7658 , y7659 , y7660 , y7661 , y7662 , y7663 , y7664 , y7665 , y7666 , y7667 , y7668 , y7669 , y7670 , y7671 , y7672 , y7673 , y7674 , y7675 , y7676 , y7677 , y7678 , y7679 , y7680 , y7681 , y7682 , y7683 , y7684 , y7685 , y7686 , y7687 , y7688 , y7689 , y7690 , y7691 , y7692 , y7693 , y7694 , y7695 , y7696 , y7697 , y7698 , y7699 , y7700 , y7701 , y7702 , y7703 , y7704 , y7705 , y7706 , y7707 , y7708 , y7709 , y7710 , y7711 , y7712 , y7713 , y7714 , y7715 , y7716 , y7717 , y7718 , y7719 , y7720 , y7721 , y7722 , y7723 , y7724 , y7725 , y7726 , y7727 , y7728 , y7729 , y7730 , y7731 , y7732 , y7733 , y7734 , y7735 , y7736 , y7737 , y7738 , y7739 , y7740 , y7741 , y7742 , y7743 , y7744 , y7745 , y7746 , y7747 , y7748 , y7749 , y7750 , y7751 , y7752 , y7753 , y7754 , y7755 , y7756 , y7757 , y7758 , y7759 , y7760 , y7761 , y7762 , y7763 , y7764 , y7765 , y7766 , y7767 , y7768 , y7769 , y7770 , y7771 , y7772 , y7773 , y7774 , y7775 , y7776 , y7777 , y7778 , y7779 , y7780 , y7781 , y7782 , y7783 , y7784 , y7785 , y7786 , y7787 , y7788 , y7789 , y7790 , y7791 , y7792 , y7793 , y7794 , y7795 , y7796 , y7797 , y7798 , y7799 , y7800 , y7801 , y7802 , y7803 , y7804 , y7805 , y7806 , y7807 , y7808 , y7809 , y7810 , y7811 , y7812 , y7813 , y7814 , y7815 , y7816 , y7817 , y7818 , y7819 , y7820 , y7821 , y7822 , y7823 , y7824 , y7825 , y7826 , y7827 , y7828 , y7829 , y7830 , y7831 , y7832 , y7833 , y7834 , y7835 , y7836 , y7837 , y7838 , y7839 , y7840 , y7841 , y7842 , y7843 , y7844 , y7845 , y7846 , y7847 , y7848 , y7849 , y7850 , y7851 , y7852 , y7853 , y7854 , y7855 , y7856 , y7857 , y7858 , y7859 , y7860 , y7861 , y7862 , y7863 , y7864 , y7865 , y7866 , y7867 , y7868 , y7869 , y7870 , y7871 , y7872 , y7873 , y7874 , y7875 , y7876 , y7877 , y7878 , y7879 , y7880 , y7881 , y7882 , y7883 , y7884 , y7885 , y7886 , y7887 , y7888 , y7889 , y7890 , y7891 , y7892 , y7893 , y7894 , y7895 , y7896 , y7897 , y7898 , y7899 , y7900 , y7901 , y7902 , y7903 , y7904 , y7905 , y7906 , y7907 , y7908 , y7909 , y7910 , y7911 , y7912 , y7913 , y7914 , y7915 , y7916 , y7917 , y7918 , y7919 , y7920 , y7921 , y7922 , y7923 , y7924 , y7925 , y7926 , y7927 , y7928 , y7929 , y7930 , y7931 , y7932 , y7933 , y7934 , y7935 , y7936 , y7937 , y7938 , y7939 , y7940 , y7941 , y7942 , y7943 , y7944 , y7945 , y7946 , y7947 , y7948 , y7949 , y7950 , y7951 , y7952 , y7953 , y7954 , y7955 , y7956 , y7957 , y7958 , y7959 , y7960 , y7961 , y7962 , y7963 , y7964 , y7965 , y7966 , y7967 , y7968 , y7969 , y7970 , y7971 , y7972 , y7973 , y7974 , y7975 , y7976 , y7977 , y7978 , y7979 , y7980 , y7981 , y7982 , y7983 , y7984 , y7985 , y7986 , y7987 , y7988 , y7989 , y7990 , y7991 , y7992 , y7993 , y7994 , y7995 , y7996 , y7997 , y7998 , y7999 , y8000 , y8001 , y8002 , y8003 , y8004 , y8005 , y8006 , y8007 , y8008 , y8009 , y8010 , y8011 , y8012 , y8013 , y8014 , y8015 , y8016 , y8017 , y8018 , y8019 , y8020 , y8021 , y8022 , y8023 , y8024 , y8025 , y8026 , y8027 , y8028 , y8029 , y8030 , y8031 , y8032 , y8033 , y8034 , y8035 , y8036 , y8037 , y8038 , y8039 , y8040 , y8041 , y8042 , y8043 , y8044 , y8045 , y8046 , y8047 , y8048 , y8049 , y8050 , y8051 , y8052 , y8053 , y8054 , y8055 , y8056 , y8057 , y8058 , y8059 , y8060 , y8061 , y8062 , y8063 , y8064 , y8065 , y8066 , y8067 , y8068 , y8069 , y8070 , y8071 , y8072 , y8073 , y8074 , y8075 , y8076 , y8077 , y8078 , y8079 , y8080 , y8081 , y8082 , y8083 , y8084 , y8085 , y8086 , y8087 , y8088 , y8089 , y8090 , y8091 , y8092 , y8093 , y8094 , y8095 , y8096 , y8097 , y8098 , y8099 , y8100 , y8101 , y8102 , y8103 , y8104 , y8105 , y8106 , y8107 , y8108 , y8109 , y8110 , y8111 , y8112 , y8113 , y8114 , y8115 , y8116 , y8117 , y8118 , y8119 , y8120 , y8121 , y8122 , y8123 , y8124 , y8125 , y8126 , y8127 , y8128 , y8129 , y8130 , y8131 , y8132 , y8133 , y8134 , y8135 , y8136 , y8137 , y8138 , y8139 , y8140 , y8141 , y8142 , y8143 , y8144 , y8145 , y8146 , y8147 , y8148 , y8149 , y8150 , y8151 , y8152 , y8153 , y8154 , y8155 , y8156 , y8157 , y8158 , y8159 , y8160 , y8161 , y8162 , y8163 , y8164 , y8165 , y8166 , y8167 , y8168 , y8169 , y8170 , y8171 , y8172 , y8173 , y8174 , y8175 , y8176 , y8177 , y8178 , y8179 , y8180 , y8181 , y8182 , y8183 , y8184 , y8185 , y8186 , y8187 , y8188 , y8189 , y8190 , y8191 , y8192 , y8193 , y8194 , y8195 , y8196 , y8197 , y8198 , y8199 , y8200 , y8201 , y8202 , y8203 , y8204 , y8205 , y8206 , y8207 , y8208 , y8209 , y8210 , y8211 , y8212 , y8213 , y8214 , y8215 , y8216 , y8217 , y8218 , y8219 , y8220 , y8221 , y8222 , y8223 , y8224 , y8225 , y8226 , y8227 , y8228 , y8229 , y8230 , y8231 , y8232 , y8233 , y8234 , y8235 , y8236 , y8237 , y8238 , y8239 , y8240 , y8241 , y8242 , y8243 , y8244 , y8245 , y8246 , y8247 , y8248 , y8249 , y8250 , y8251 , y8252 , y8253 , y8254 , y8255 , y8256 , y8257 , y8258 , y8259 , y8260 , y8261 , y8262 , y8263 , y8264 , y8265 , y8266 , y8267 , y8268 , y8269 , y8270 , y8271 , y8272 , y8273 , y8274 , y8275 , y8276 , y8277 , y8278 , y8279 , y8280 , y8281 , y8282 , y8283 , y8284 , y8285 , y8286 , y8287 , y8288 , y8289 , y8290 , y8291 , y8292 , y8293 , y8294 , y8295 , y8296 , y8297 , y8298 , y8299 , y8300 , y8301 , y8302 , y8303 , y8304 , y8305 , y8306 , y8307 , y8308 , y8309 , y8310 , y8311 , y8312 , y8313 , y8314 , y8315 , y8316 , y8317 , y8318 , y8319 , y8320 , y8321 , y8322 , y8323 , y8324 , y8325 , y8326 , y8327 , y8328 , y8329 , y8330 , y8331 , y8332 , y8333 , y8334 , y8335 , y8336 , y8337 , y8338 , y8339 , y8340 , y8341 , y8342 , y8343 , y8344 , y8345 , y8346 , y8347 , y8348 , y8349 , y8350 , y8351 , y8352 , y8353 , y8354 , y8355 , y8356 , y8357 , y8358 , y8359 , y8360 , y8361 , y8362 , y8363 , y8364 , y8365 , y8366 , y8367 , y8368 , y8369 , y8370 , y8371 , y8372 , y8373 , y8374 , y8375 , y8376 , y8377 , y8378 , y8379 , y8380 , y8381 , y8382 , y8383 , y8384 , y8385 , y8386 , y8387 , y8388 , y8389 , y8390 , y8391 , y8392 , y8393 , y8394 , y8395 , y8396 , y8397 , y8398 , y8399 , y8400 , y8401 , y8402 , y8403 , y8404 , y8405 , y8406 , y8407 , y8408 , y8409 , y8410 , y8411 , y8412 , y8413 , y8414 , y8415 , y8416 , y8417 , y8418 , y8419 , y8420 , y8421 , y8422 , y8423 , y8424 , y8425 , y8426 , y8427 , y8428 , y8429 , y8430 , y8431 , y8432 , y8433 , y8434 , y8435 , y8436 , y8437 , y8438 , y8439 , y8440 , y8441 , y8442 , y8443 , y8444 , y8445 , y8446 , y8447 , y8448 , y8449 , y8450 , y8451 , y8452 , y8453 , y8454 , y8455 , y8456 , y8457 , y8458 , y8459 , y8460 , y8461 , y8462 , y8463 , y8464 , y8465 , y8466 , y8467 , y8468 , y8469 , y8470 , y8471 , y8472 , y8473 , y8474 , y8475 , y8476 , y8477 , y8478 , y8479 , y8480 , y8481 , y8482 , y8483 , y8484 , y8485 , y8486 , y8487 , y8488 , y8489 , y8490 , y8491 , y8492 , y8493 , y8494 , y8495 , y8496 , y8497 , y8498 , y8499 , y8500 , y8501 , y8502 , y8503 , y8504 , y8505 , y8506 , y8507 , y8508 , y8509 , y8510 , y8511 , y8512 , y8513 , y8514 , y8515 , y8516 , y8517 , y8518 , y8519 , y8520 , y8521 , y8522 , y8523 , y8524 , y8525 , y8526 , y8527 , y8528 , y8529 , y8530 , y8531 , y8532 , y8533 , y8534 , y8535 , y8536 , y8537 , y8538 , y8539 , y8540 , y8541 , y8542 , y8543 , y8544 , y8545 , y8546 , y8547 , y8548 , y8549 , y8550 , y8551 , y8552 , y8553 , y8554 , y8555 , y8556 , y8557 , y8558 , y8559 , y8560 , y8561 , y8562 , y8563 , y8564 , y8565 , y8566 , y8567 , y8568 , y8569 , y8570 , y8571 , y8572 , y8573 , y8574 , y8575 , y8576 , y8577 , y8578 , y8579 , y8580 , y8581 , y8582 , y8583 , y8584 , y8585 , y8586 , y8587 , y8588 , y8589 , y8590 , y8591 , y8592 , y8593 , y8594 , y8595 , y8596 , y8597 , y8598 , y8599 , y8600 , y8601 , y8602 , y8603 , y8604 , y8605 , y8606 , y8607 , y8608 , y8609 , y8610 , y8611 , y8612 , y8613 , y8614 , y8615 , y8616 , y8617 , y8618 , y8619 , y8620 , y8621 , y8622 , y8623 , y8624 , y8625 , y8626 , y8627 , y8628 , y8629 , y8630 , y8631 , y8632 , y8633 , y8634 , y8635 , y8636 , y8637 , y8638 , y8639 , y8640 , y8641 , y8642 , y8643 , y8644 , y8645 , y8646 , y8647 , y8648 , y8649 , y8650 , y8651 , y8652 , y8653 , y8654 , y8655 , y8656 , y8657 , y8658 , y8659 , y8660 , y8661 , y8662 , y8663 , y8664 , y8665 , y8666 , y8667 , y8668 , y8669 , y8670 , y8671 , y8672 , y8673 , y8674 , y8675 , y8676 , y8677 , y8678 , y8679 , y8680 , y8681 , y8682 , y8683 , y8684 , y8685 , y8686 , y8687 , y8688 , y8689 , y8690 , y8691 , y8692 , y8693 , y8694 , y8695 , y8696 , y8697 , y8698 , y8699 , y8700 , y8701 , y8702 , y8703 , y8704 , y8705 , y8706 , y8707 , y8708 , y8709 , y8710 , y8711 , y8712 , y8713 , y8714 , y8715 , y8716 , y8717 , y8718 , y8719 , y8720 , y8721 , y8722 , y8723 , y8724 , y8725 , y8726 , y8727 , y8728 , y8729 , y8730 , y8731 , y8732 , y8733 , y8734 , y8735 , y8736 , y8737 , y8738 , y8739 , y8740 , y8741 , y8742 , y8743 , y8744 , y8745 , y8746 , y8747 , y8748 , y8749 , y8750 , y8751 , y8752 , y8753 , y8754 , y8755 , y8756 , y8757 , y8758 , y8759 , y8760 , y8761 , y8762 , y8763 , y8764 , y8765 , y8766 , y8767 , y8768 , y8769 , y8770 , y8771 , y8772 , y8773 , y8774 , y8775 , y8776 , y8777 , y8778 , y8779 , y8780 , y8781 , y8782 , y8783 , y8784 , y8785 , y8786 , y8787 , y8788 , y8789 , y8790 , y8791 , y8792 , y8793 , y8794 , y8795 , y8796 , y8797 , y8798 , y8799 , y8800 , y8801 , y8802 , y8803 , y8804 , y8805 , y8806 , y8807 , y8808 , y8809 , y8810 , y8811 , y8812 , y8813 , y8814 , y8815 , y8816 , y8817 , y8818 , y8819 , y8820 , y8821 , y8822 , y8823 , y8824 , y8825 , y8826 , y8827 , y8828 , y8829 , y8830 , y8831 , y8832 , y8833 , y8834 , y8835 , y8836 , y8837 , y8838 , y8839 , y8840 , y8841 , y8842 , y8843 , y8844 , y8845 , y8846 , y8847 , y8848 , y8849 , y8850 , y8851 , y8852 , y8853 , y8854 , y8855 , y8856 , y8857 , y8858 , y8859 , y8860 , y8861 , y8862 , y8863 , y8864 , y8865 , y8866 , y8867 , y8868 , y8869 , y8870 , y8871 , y8872 , y8873 , y8874 , y8875 , y8876 , y8877 , y8878 , y8879 , y8880 , y8881 , y8882 , y8883 , y8884 , y8885 , y8886 , y8887 , y8888 , y8889 , y8890 , y8891 , y8892 , y8893 , y8894 , y8895 , y8896 , y8897 , y8898 , y8899 , y8900 , y8901 , y8902 , y8903 , y8904 , y8905 , y8906 , y8907 , y8908 , y8909 , y8910 , y8911 , y8912 , y8913 , y8914 , y8915 , y8916 , y8917 , y8918 , y8919 , y8920 , y8921 , y8922 , y8923 , y8924 , y8925 , y8926 , y8927 , y8928 , y8929 , y8930 , y8931 , y8932 , y8933 , y8934 , y8935 , y8936 , y8937 , y8938 , y8939 , y8940 , y8941 , y8942 , y8943 , y8944 , y8945 , y8946 , y8947 , y8948 , y8949 , y8950 , y8951 , y8952 , y8953 , y8954 , y8955 , y8956 , y8957 , y8958 , y8959 , y8960 , y8961 , y8962 , y8963 , y8964 , y8965 , y8966 , y8967 , y8968 , y8969 , y8970 , y8971 , y8972 , y8973 , y8974 , y8975 , y8976 , y8977 , y8978 , y8979 , y8980 , y8981 , y8982 , y8983 , y8984 , y8985 , y8986 , y8987 , y8988 , y8989 , y8990 , y8991 , y8992 , y8993 , y8994 , y8995 , y8996 , y8997 , y8998 , y8999 , y9000 , y9001 , y9002 , y9003 , y9004 , y9005 , y9006 , y9007 , y9008 , y9009 , y9010 , y9011 , y9012 , y9013 , y9014 , y9015 , y9016 , y9017 , y9018 , y9019 , y9020 , y9021 , y9022 , y9023 , y9024 , y9025 , y9026 , y9027 , y9028 , y9029 , y9030 , y9031 , y9032 , y9033 , y9034 , y9035 , y9036 , y9037 , y9038 , y9039 , y9040 , y9041 , y9042 , y9043 , y9044 , y9045 , y9046 , y9047 , y9048 , y9049 , y9050 , y9051 , y9052 , y9053 , y9054 , y9055 , y9056 , y9057 , y9058 , y9059 , y9060 , y9061 , y9062 , y9063 , y9064 , y9065 , y9066 , y9067 , y9068 , y9069 , y9070 , y9071 , y9072 , y9073 , y9074 , y9075 , y9076 , y9077 , y9078 , y9079 , y9080 , y9081 , y9082 , y9083 , y9084 , y9085 , y9086 , y9087 , y9088 , y9089 , y9090 , y9091 , y9092 , y9093 , y9094 , y9095 , y9096 , y9097 , y9098 , y9099 , y9100 , y9101 , y9102 , y9103 , y9104 , y9105 , y9106 , y9107 , y9108 , y9109 , y9110 , y9111 , y9112 , y9113 , y9114 , y9115 , y9116 , y9117 , y9118 , y9119 , y9120 , y9121 , y9122 , y9123 , y9124 , y9125 , y9126 , y9127 , y9128 , y9129 , y9130 , y9131 , y9132 , y9133 , y9134 , y9135 , y9136 , y9137 , y9138 , y9139 , y9140 , y9141 , y9142 , y9143 , y9144 , y9145 , y9146 , y9147 , y9148 , y9149 , y9150 , y9151 , y9152 , y9153 , y9154 , y9155 , y9156 , y9157 , y9158 , y9159 , y9160 , y9161 , y9162 , y9163 , y9164 , y9165 , y9166 , y9167 , y9168 , y9169 , y9170 , y9171 , y9172 , y9173 , y9174 , y9175 , y9176 , y9177 , y9178 , y9179 , y9180 , y9181 , y9182 , y9183 , y9184 , y9185 , y9186 , y9187 , y9188 , y9189 , y9190 , y9191 , y9192 , y9193 , y9194 , y9195 , y9196 , y9197 , y9198 , y9199 , y9200 , y9201 , y9202 , y9203 , y9204 , y9205 , y9206 , y9207 , y9208 , y9209 , y9210 , y9211 , y9212 , y9213 , y9214 , y9215 , y9216 , y9217 , y9218 , y9219 , y9220 , y9221 , y9222 , y9223 , y9224 , y9225 , y9226 , y9227 , y9228 , y9229 , y9230 , y9231 , y9232 , y9233 , y9234 , y9235 , y9236 , y9237 , y9238 , y9239 , y9240 , y9241 , y9242 , y9243 , y9244 , y9245 , y9246 , y9247 , y9248 , y9249 , y9250 , y9251 , y9252 , y9253 , y9254 , y9255 , y9256 , y9257 , y9258 , y9259 , y9260 , y9261 , y9262 , y9263 , y9264 , y9265 , y9266 , y9267 , y9268 , y9269 , y9270 , y9271 , y9272 , y9273 , y9274 , y9275 , y9276 , y9277 , y9278 , y9279 , y9280 , y9281 , y9282 , y9283 , y9284 , y9285 , y9286 , y9287 , y9288 , y9289 , y9290 , y9291 , y9292 , y9293 , y9294 , y9295 , y9296 , y9297 , y9298 , y9299 , y9300 , y9301 , y9302 , y9303 , y9304 , y9305 , y9306 , y9307 , y9308 , y9309 , y9310 , y9311 , y9312 , y9313 , y9314 , y9315 , y9316 , y9317 , y9318 , y9319 , y9320 , y9321 , y9322 , y9323 , y9324 , y9325 , y9326 , y9327 , y9328 , y9329 , y9330 , y9331 , y9332 , y9333 , y9334 , y9335 , y9336 , y9337 , y9338 , y9339 , y9340 , y9341 , y9342 , y9343 , y9344 , y9345 , y9346 , y9347 , y9348 , y9349 , y9350 , y9351 , y9352 , y9353 , y9354 , y9355 , y9356 , y9357 , y9358 , y9359 , y9360 , y9361 , y9362 , y9363 , y9364 , y9365 , y9366 , y9367 , y9368 , y9369 , y9370 , y9371 , y9372 , y9373 , y9374 , y9375 , y9376 , y9377 , y9378 , y9379 , y9380 , y9381 , y9382 , y9383 , y9384 , y9385 , y9386 , y9387 , y9388 , y9389 , y9390 , y9391 , y9392 , y9393 , y9394 , y9395 , y9396 , y9397 , y9398 , y9399 , y9400 , y9401 , y9402 , y9403 , y9404 , y9405 , y9406 , y9407 , y9408 , y9409 , y9410 , y9411 , y9412 , y9413 , y9414 , y9415 , y9416 , y9417 , y9418 , y9419 , y9420 , y9421 , y9422 , y9423 , y9424 , y9425 , y9426 , y9427 , y9428 , y9429 , y9430 , y9431 , y9432 , y9433 , y9434 , y9435 , y9436 , y9437 , y9438 , y9439 , y9440 , y9441 , y9442 , y9443 , y9444 , y9445 , y9446 , y9447 , y9448 , y9449 , y9450 , y9451 , y9452 , y9453 , y9454 , y9455 , y9456 , y9457 , y9458 , y9459 , y9460 , y9461 , y9462 , y9463 , y9464 , y9465 , y9466 , y9467 , y9468 , y9469 , y9470 , y9471 , y9472 , y9473 , y9474 , y9475 , y9476 , y9477 , y9478 , y9479 , y9480 , y9481 , y9482 , y9483 , y9484 , y9485 , y9486 , y9487 , y9488 , y9489 , y9490 , y9491 , y9492 , y9493 , y9494 , y9495 , y9496 , y9497 , y9498 , y9499 , y9500 , y9501 , y9502 , y9503 , y9504 , y9505 , y9506 , y9507 , y9508 , y9509 , y9510 , y9511 , y9512 , y9513 , y9514 , y9515 , y9516 , y9517 , y9518 , y9519 , y9520 , y9521 , y9522 , y9523 , y9524 , y9525 , y9526 , y9527 , y9528 , y9529 , y9530 , y9531 , y9532 , y9533 , y9534 , y9535 , y9536 , y9537 , y9538 , y9539 , y9540 , y9541 , y9542 , y9543 , y9544 , y9545 , y9546 , y9547 , y9548 , y9549 , y9550 , y9551 , y9552 , y9553 , y9554 , y9555 , y9556 , y9557 , y9558 , y9559 , y9560 , y9561 , y9562 , y9563 , y9564 , y9565 , y9566 , y9567 , y9568 , y9569 , y9570 , y9571 , y9572 , y9573 , y9574 , y9575 , y9576 , y9577 , y9578 , y9579 , y9580 , y9581 , y9582 , y9583 , y9584 , y9585 , y9586 , y9587 , y9588 , y9589 , y9590 , y9591 , y9592 , y9593 , y9594 , y9595 , y9596 , y9597 , y9598 , y9599 , y9600 , y9601 , y9602 , y9603 , y9604 , y9605 , y9606 , y9607 , y9608 , y9609 , y9610 , y9611 , y9612 , y9613 , y9614 , y9615 , y9616 , y9617 , y9618 , y9619 , y9620 , y9621 , y9622 , y9623 , y9624 , y9625 , y9626 , y9627 , y9628 , y9629 , y9630 , y9631 , y9632 , y9633 , y9634 , y9635 , y9636 , y9637 , y9638 , y9639 , y9640 , y9641 , y9642 , y9643 , y9644 , y9645 , y9646 , y9647 , y9648 , y9649 , y9650 , y9651 , y9652 , y9653 , y9654 , y9655 , y9656 , y9657 , y9658 , y9659 , y9660 , y9661 , y9662 , y9663 , y9664 , y9665 , y9666 , y9667 , y9668 , y9669 , y9670 , y9671 , y9672 , y9673 , y9674 , y9675 , y9676 , y9677 , y9678 , y9679 , y9680 , y9681 , y9682 , y9683 , y9684 , y9685 , y9686 , y9687 , y9688 , y9689 , y9690 , y9691 , y9692 , y9693 , y9694 , y9695 , y9696 , y9697 , y9698 , y9699 , y9700 , y9701 , y9702 , y9703 , y9704 , y9705 , y9706 , y9707 , y9708 , y9709 , y9710 , y9711 , y9712 , y9713 , y9714 , y9715 , y9716 , y9717 , y9718 , y9719 , y9720 , y9721 , y9722 , y9723 , y9724 , y9725 , y9726 , y9727 , y9728 , y9729 , y9730 , y9731 , y9732 , y9733 , y9734 , y9735 , y9736 , y9737 , y9738 , y9739 , y9740 , y9741 , y9742 , y9743 , y9744 , y9745 , y9746 , y9747 , y9748 , y9749 , y9750 , y9751 , y9752 , y9753 , y9754 , y9755 , y9756 , y9757 , y9758 , y9759 , y9760 , y9761 , y9762 , y9763 , y9764 , y9765 , y9766 , y9767 , y9768 , y9769 , y9770 , y9771 , y9772 , y9773 , y9774 , y9775 , y9776 , y9777 , y9778 , y9779 , y9780 , y9781 , y9782 , y9783 , y9784 , y9785 , y9786 , y9787 , y9788 , y9789 , y9790 , y9791 , y9792 , y9793 , y9794 , y9795 , y9796 , y9797 , y9798 , y9799 , y9800 , y9801 , y9802 , y9803 , y9804 , y9805 , y9806 , y9807 , y9808 , y9809 , y9810 , y9811 , y9812 , y9813 , y9814 , y9815 , y9816 , y9817 , y9818 , y9819 , y9820 , y9821 , y9822 , y9823 , y9824 , y9825 , y9826 , y9827 , y9828 , y9829 , y9830 , y9831 , y9832 , y9833 , y9834 , y9835 , y9836 , y9837 , y9838 , y9839 , y9840 , y9841 , y9842 , y9843 , y9844 , y9845 , y9846 , y9847 , y9848 , y9849 , y9850 , y9851 , y9852 , y9853 , y9854 , y9855 , y9856 , y9857 , y9858 , y9859 , y9860 , y9861 , y9862 , y9863 , y9864 , y9865 , y9866 , y9867 , y9868 , y9869 , y9870 , y9871 , y9872 , y9873 , y9874 , y9875 , y9876 , y9877 , y9878 , y9879 , y9880 , y9881 , y9882 , y9883 , y9884 , y9885 , y9886 , y9887 , y9888 , y9889 , y9890 , y9891 , y9892 , y9893 , y9894 , y9895 , y9896 , y9897 , y9898 , y9899 , y9900 , y9901 , y9902 , y9903 , y9904 , y9905 , y9906 , y9907 , y9908 , y9909 , y9910 , y9911 , y9912 , y9913 , y9914 , y9915 , y9916 , y9917 , y9918 , y9919 , y9920 , y9921 , y9922 , y9923 , y9924 , y9925 , y9926 , y9927 , y9928 , y9929 , y9930 , y9931 , y9932 , y9933 , y9934 , y9935 , y9936 , y9937 , y9938 , y9939 , y9940 , y9941 , y9942 , y9943 , y9944 , y9945 , y9946 , y9947 , y9948 , y9949 , y9950 , y9951 , y9952 , y9953 , y9954 , y9955 , y9956 , y9957 , y9958 , y9959 , y9960 , y9961 , y9962 , y9963 , y9964 , y9965 , y9966 , y9967 , y9968 , y9969 , y9970 , y9971 , y9972 , y9973 , y9974 , y9975 , y9976 , y9977 , y9978 , y9979 , y9980 , y9981 , y9982 , y9983 , y9984 , y9985 , y9986 , y9987 , y9988 , y9989 , y9990 , y9991 , y9992 , y9993 , y9994 , y9995 , y9996 , y9997 , y9998 , y9999 , y10000 , y10001 , y10002 , y10003 , y10004 , y10005 , y10006 , y10007 , y10008 , y10009 , y10010 , y10011 , y10012 , y10013 , y10014 , y10015 , y10016 , y10017 , y10018 , y10019 , y10020 , y10021 , y10022 , y10023 , y10024 , y10025 , y10026 , y10027 , y10028 , y10029 , y10030 , y10031 , y10032 , y10033 , y10034 , y10035 , y10036 , y10037 , y10038 , y10039 , y10040 , y10041 , y10042 , y10043 , y10044 , y10045 , y10046 , y10047 , y10048 , y10049 , y10050 , y10051 , y10052 , y10053 , y10054 , y10055 , y10056 , y10057 , y10058 , y10059 , y10060 , y10061 , y10062 , y10063 , y10064 , y10065 , y10066 , y10067 , y10068 , y10069 , y10070 , y10071 , y10072 , y10073 , y10074 , y10075 , y10076 , y10077 , y10078 , y10079 , y10080 , y10081 , y10082 , y10083 , y10084 , y10085 , y10086 , y10087 , y10088 , y10089 , y10090 , y10091 , y10092 , y10093 , y10094 , y10095 , y10096 , y10097 , y10098 , y10099 , y10100 , y10101 , y10102 , y10103 , y10104 , y10105 , y10106 , y10107 , y10108 , y10109 , y10110 , y10111 , y10112 , y10113 , y10114 , y10115 , y10116 , y10117 , y10118 , y10119 , y10120 , y10121 , y10122 , y10123 , y10124 , y10125 , y10126 , y10127 , y10128 , y10129 , y10130 , y10131 , y10132 , y10133 , y10134 , y10135 , y10136 , y10137 , y10138 , y10139 , y10140 , y10141 , y10142 , y10143 , y10144 , y10145 , y10146 , y10147 , y10148 , y10149 , y10150 , y10151 , y10152 , y10153 , y10154 , y10155 , y10156 , y10157 , y10158 , y10159 , y10160 , y10161 , y10162 , y10163 , y10164 , y10165 , y10166 , y10167 , y10168 , y10169 , y10170 , y10171 , y10172 , y10173 , y10174 , y10175 , y10176 , y10177 , y10178 , y10179 , y10180 , y10181 , y10182 , y10183 , y10184 , y10185 , y10186 , y10187 , y10188 , y10189 , y10190 , y10191 , y10192 , y10193 , y10194 , y10195 , y10196 , y10197 , y10198 , y10199 , y10200 , y10201 , y10202 , y10203 , y10204 , y10205 , y10206 , y10207 , y10208 , y10209 , y10210 , y10211 , y10212 , y10213 , y10214 , y10215 , y10216 , y10217 , y10218 , y10219 , y10220 , y10221 , y10222 , y10223 , y10224 , y10225 , y10226 , y10227 , y10228 , y10229 , y10230 , y10231 , y10232 , y10233 , y10234 , y10235 , y10236 , y10237 , y10238 , y10239 , y10240 , y10241 , y10242 , y10243 , y10244 , y10245 , y10246 , y10247 , y10248 , y10249 , y10250 , y10251 , y10252 , y10253 , y10254 , y10255 , y10256 , y10257 , y10258 , y10259 , y10260 , y10261 , y10262 , y10263 , y10264 , y10265 , y10266 , y10267 , y10268 , y10269 , y10270 , y10271 , y10272 , y10273 , y10274 , y10275 , y10276 , y10277 , y10278 , y10279 , y10280 , y10281 , y10282 , y10283 , y10284 , y10285 , y10286 , y10287 , y10288 , y10289 , y10290 , y10291 , y10292 , y10293 , y10294 , y10295 , y10296 , y10297 , y10298 , y10299 , y10300 , y10301 , y10302 , y10303 , y10304 , y10305 , y10306 , y10307 , y10308 , y10309 , y10310 , y10311 , y10312 , y10313 , y10314 , y10315 , y10316 , y10317 , y10318 , y10319 , y10320 , y10321 , y10322 , y10323 , y10324 , y10325 , y10326 , y10327 , y10328 , y10329 , y10330 , y10331 , y10332 , y10333 , y10334 , y10335 , y10336 , y10337 , y10338 , y10339 , y10340 , y10341 , y10342 , y10343 , y10344 , y10345 , y10346 , y10347 , y10348 , y10349 , y10350 , y10351 , y10352 , y10353 , y10354 , y10355 , y10356 , y10357 , y10358 , y10359 , y10360 , y10361 , y10362 , y10363 , y10364 , y10365 , y10366 , y10367 , y10368 , y10369 , y10370 , y10371 , y10372 , y10373 , y10374 , y10375 , y10376 , y10377 , y10378 , y10379 , y10380 , y10381 , y10382 , y10383 , y10384 , y10385 , y10386 , y10387 , y10388 , y10389 , y10390 , y10391 , y10392 , y10393 , y10394 , y10395 , y10396 , y10397 , y10398 , y10399 , y10400 , y10401 , y10402 , y10403 , y10404 , y10405 , y10406 , y10407 , y10408 , y10409 , y10410 , y10411 , y10412 , y10413 , y10414 , y10415 , y10416 , y10417 , y10418 , y10419 , y10420 , y10421 , y10422 , y10423 , y10424 , y10425 , y10426 , y10427 , y10428 , y10429 , y10430 , y10431 , y10432 , y10433 , y10434 , y10435 , y10436 , y10437 , y10438 , y10439 , y10440 , y10441 , y10442 , y10443 , y10444 , y10445 , y10446 , y10447 , y10448 , y10449 , y10450 , y10451 , y10452 , y10453 , y10454 , y10455 , y10456 , y10457 , y10458 , y10459 , y10460 , y10461 , y10462 , y10463 , y10464 , y10465 , y10466 , y10467 , y10468 , y10469 , y10470 , y10471 , y10472 , y10473 , y10474 , y10475 , y10476 , y10477 , y10478 , y10479 , y10480 , y10481 , y10482 , y10483 , y10484 , y10485 , y10486 , y10487 , y10488 , y10489 , y10490 , y10491 , y10492 , y10493 , y10494 , y10495 , y10496 , y10497 , y10498 , y10499 , y10500 , y10501 , y10502 , y10503 , y10504 , y10505 , y10506 , y10507 , y10508 , y10509 , y10510 , y10511 , y10512 , y10513 , y10514 , y10515 , y10516 , y10517 , y10518 , y10519 , y10520 , y10521 , y10522 , y10523 , y10524 , y10525 , y10526 , y10527 , y10528 , y10529 , y10530 , y10531 , y10532 , y10533 , y10534 , y10535 , y10536 , y10537 , y10538 , y10539 , y10540 , y10541 , y10542 , y10543 , y10544 , y10545 , y10546 , y10547 , y10548 , y10549 , y10550 , y10551 , y10552 , y10553 , y10554 , y10555 , y10556 , y10557 , y10558 , y10559 , y10560 , y10561 , y10562 , y10563 , y10564 , y10565 , y10566 , y10567 , y10568 , y10569 , y10570 , y10571 , y10572 , y10573 , y10574 , y10575 , y10576 , y10577 , y10578 , y10579 , y10580 , y10581 , y10582 , y10583 , y10584 , y10585 , y10586 , y10587 , y10588 , y10589 , y10590 , y10591 , y10592 , y10593 , y10594 , y10595 , y10596 , y10597 , y10598 , y10599 , y10600 , y10601 , y10602 , y10603 , y10604 , y10605 , y10606 , y10607 , y10608 , y10609 , y10610 , y10611 , y10612 , y10613 , y10614 , y10615 , y10616 , y10617 , y10618 , y10619 , y10620 , y10621 , y10622 , y10623 , y10624 , y10625 , y10626 , y10627 , y10628 , y10629 , y10630 , y10631 , y10632 , y10633 , y10634 , y10635 , y10636 , y10637 , y10638 , y10639 , y10640 , y10641 , y10642 , y10643 , y10644 , y10645 , y10646 , y10647 , y10648 , y10649 , y10650 , y10651 , y10652 , y10653 , y10654 , y10655 , y10656 , y10657 , y10658 , y10659 , y10660 , y10661 , y10662 , y10663 , y10664 , y10665 , y10666 , y10667 , y10668 , y10669 , y10670 , y10671 , y10672 , y10673 , y10674 , y10675 , y10676 , y10677 , y10678 , y10679 , y10680 , y10681 , y10682 , y10683 , y10684 , y10685 , y10686 , y10687 , y10688 , y10689 , y10690 , y10691 , y10692 , y10693 , y10694 , y10695 , y10696 , y10697 , y10698 , y10699 , y10700 , y10701 , y10702 , y10703 , y10704 , y10705 , y10706 , y10707 , y10708 , y10709 , y10710 , y10711 , y10712 , y10713 , y10714 , y10715 , y10716 , y10717 , y10718 , y10719 , y10720 , y10721 , y10722 , y10723 , y10724 , y10725 , y10726 , y10727 , y10728 , y10729 , y10730 , y10731 , y10732 , y10733 , y10734 , y10735 , y10736 , y10737 , y10738 , y10739 , y10740 , y10741 , y10742 , y10743 , y10744 , y10745 , y10746 , y10747 , y10748 , y10749 , y10750 , y10751 , y10752 , y10753 , y10754 , y10755 , y10756 , y10757 , y10758 , y10759 , y10760 , y10761 , y10762 , y10763 , y10764 , y10765 , y10766 , y10767 , y10768 , y10769 , y10770 , y10771 , y10772 , y10773 , y10774 , y10775 , y10776 , y10777 , y10778 , y10779 , y10780 , y10781 , y10782 , y10783 , y10784 , y10785 , y10786 , y10787 , y10788 , y10789 , y10790 , y10791 , y10792 , y10793 , y10794 , y10795 , y10796 , y10797 , y10798 , y10799 , y10800 , y10801 , y10802 , y10803 , y10804 , y10805 , y10806 , y10807 , y10808 , y10809 , y10810 , y10811 , y10812 , y10813 , y10814 , y10815 , y10816 , y10817 , y10818 , y10819 , y10820 , y10821 , y10822 , y10823 , y10824 , y10825 , y10826 , y10827 , y10828 , y10829 , y10830 , y10831 , y10832 , y10833 , y10834 , y10835 , y10836 , y10837 , y10838 , y10839 , y10840 , y10841 , y10842 , y10843 , y10844 , y10845 , y10846 , y10847 , y10848 , y10849 , y10850 , y10851 , y10852 , y10853 , y10854 , y10855 , y10856 , y10857 , y10858 , y10859 , y10860 , y10861 , y10862 , y10863 , y10864 , y10865 , y10866 , y10867 , y10868 , y10869 , y10870 , y10871 , y10872 , y10873 , y10874 , y10875 , y10876 , y10877 , y10878 , y10879 , y10880 , y10881 , y10882 , y10883 , y10884 , y10885 , y10886 , y10887 , y10888 , y10889 , y10890 , y10891 , y10892 , y10893 , y10894 , y10895 , y10896 , y10897 , y10898 , y10899 , y10900 , y10901 , y10902 , y10903 , y10904 , y10905 , y10906 , y10907 , y10908 , y10909 , y10910 , y10911 , y10912 , y10913 , y10914 , y10915 , y10916 , y10917 , y10918 , y10919 , y10920 , y10921 , y10922 , y10923 , y10924 , y10925 , y10926 , y10927 , y10928 , y10929 , y10930 , y10931 , y10932 , y10933 , y10934 , y10935 , y10936 , y10937 , y10938 , y10939 , y10940 , y10941 , y10942 , y10943 , y10944 , y10945 , y10946 , y10947 , y10948 , y10949 , y10950 , y10951 , y10952 , y10953 , y10954 , y10955 , y10956 , y10957 , y10958 , y10959 , y10960 , y10961 , y10962 , y10963 , y10964 , y10965 , y10966 , y10967 , y10968 , y10969 , y10970 , y10971 , y10972 , y10973 , y10974 , y10975 , y10976 , y10977 , y10978 , y10979 , y10980 , y10981 , y10982 , y10983 , y10984 , y10985 , y10986 , y10987 , y10988 , y10989 , y10990 , y10991 , y10992 , y10993 , y10994 , y10995 , y10996 , y10997 , y10998 , y10999 , y11000 , y11001 , y11002 , y11003 , y11004 , y11005 , y11006 , y11007 , y11008 , y11009 , y11010 , y11011 , y11012 , y11013 , y11014 , y11015 , y11016 , y11017 , y11018 , y11019 , y11020 , y11021 , y11022 , y11023 , y11024 , y11025 , y11026 , y11027 , y11028 , y11029 , y11030 , y11031 , y11032 , y11033 , y11034 , y11035 , y11036 , y11037 , y11038 , y11039 , y11040 , y11041 , y11042 , y11043 , y11044 , y11045 , y11046 , y11047 , y11048 , y11049 , y11050 , y11051 , y11052 , y11053 , y11054 , y11055 , y11056 , y11057 , y11058 , y11059 , y11060 , y11061 , y11062 , y11063 , y11064 , y11065 , y11066 , y11067 , y11068 , y11069 , y11070 , y11071 , y11072 , y11073 , y11074 , y11075 , y11076 , y11077 , y11078 , y11079 , y11080 , y11081 , y11082 , y11083 , y11084 , y11085 , y11086 , y11087 , y11088 , y11089 , y11090 , y11091 , y11092 , y11093 , y11094 , y11095 , y11096 , y11097 , y11098 , y11099 , y11100 , y11101 , y11102 , y11103 , y11104 , y11105 , y11106 , y11107 , y11108 , y11109 , y11110 , y11111 , y11112 , y11113 , y11114 , y11115 , y11116 , y11117 , y11118 , y11119 , y11120 , y11121 , y11122 , y11123 , y11124 , y11125 , y11126 , y11127 , y11128 , y11129 , y11130 , y11131 , y11132 , y11133 , y11134 , y11135 , y11136 , y11137 , y11138 , y11139 , y11140 , y11141 , y11142 , y11143 , y11144 , y11145 , y11146 , y11147 , y11148 , y11149 , y11150 , y11151 , y11152 , y11153 , y11154 , y11155 , y11156 , y11157 , y11158 , y11159 , y11160 , y11161 , y11162 , y11163 , y11164 , y11165 , y11166 , y11167 , y11168 , y11169 , y11170 , y11171 , y11172 , y11173 , y11174 , y11175 , y11176 , y11177 , y11178 , y11179 , y11180 , y11181 , y11182 , y11183 , y11184 , y11185 , y11186 , y11187 , y11188 , y11189 , y11190 , y11191 , y11192 , y11193 , y11194 , y11195 , y11196 , y11197 , y11198 , y11199 , y11200 , y11201 , y11202 , y11203 , y11204 , y11205 , y11206 , y11207 , y11208 , y11209 , y11210 , y11211 , y11212 , y11213 , y11214 , y11215 , y11216 , y11217 , y11218 , y11219 , y11220 , y11221 , y11222 , y11223 , y11224 , y11225 , y11226 , y11227 , y11228 , y11229 , y11230 , y11231 , y11232 , y11233 , y11234 , y11235 , y11236 , y11237 , y11238 , y11239 , y11240 , y11241 , y11242 , y11243 , y11244 , y11245 , y11246 , y11247 , y11248 , y11249 , y11250 , y11251 , y11252 , y11253 , y11254 , y11255 , y11256 , y11257 , y11258 , y11259 , y11260 , y11261 , y11262 , y11263 , y11264 , y11265 , y11266 , y11267 , y11268 , y11269 , y11270 , y11271 , y11272 , y11273 , y11274 , y11275 , y11276 , y11277 , y11278 , y11279 , y11280 , y11281 , y11282 , y11283 , y11284 , y11285 , y11286 , y11287 , y11288 , y11289 , y11290 , y11291 , y11292 , y11293 , y11294 , y11295 , y11296 , y11297 , y11298 , y11299 , y11300 , y11301 , y11302 , y11303 , y11304 , y11305 , y11306 , y11307 , y11308 , y11309 , y11310 , y11311 , y11312 , y11313 , y11314 , y11315 , y11316 , y11317 , y11318 , y11319 , y11320 , y11321 , y11322 , y11323 , y11324 , y11325 , y11326 , y11327 , y11328 , y11329 , y11330 , y11331 , y11332 , y11333 , y11334 , y11335 , y11336 , y11337 , y11338 , y11339 , y11340 , y11341 , y11342 , y11343 , y11344 , y11345 , y11346 , y11347 , y11348 , y11349 , y11350 , y11351 , y11352 , y11353 , y11354 , y11355 , y11356 , y11357 , y11358 , y11359 , y11360 , y11361 , y11362 , y11363 , y11364 , y11365 , y11366 , y11367 , y11368 , y11369 , y11370 , y11371 , y11372 , y11373 , y11374 , y11375 , y11376 , y11377 , y11378 , y11379 , y11380 , y11381 , y11382 , y11383 , y11384 , y11385 , y11386 , y11387 , y11388 , y11389 , y11390 , y11391 , y11392 , y11393 , y11394 , y11395 , y11396 , y11397 , y11398 , y11399 , y11400 , y11401 , y11402 , y11403 , y11404 , y11405 , y11406 , y11407 , y11408 , y11409 , y11410 , y11411 , y11412 , y11413 , y11414 , y11415 , y11416 , y11417 , y11418 , y11419 , y11420 , y11421 , y11422 , y11423 , y11424 , y11425 , y11426 , y11427 , y11428 , y11429 , y11430 , y11431 , y11432 , y11433 , y11434 , y11435 , y11436 , y11437 , y11438 , y11439 , y11440 , y11441 , y11442 , y11443 , y11444 , y11445 , y11446 , y11447 , y11448 , y11449 , y11450 , y11451 , y11452 , y11453 , y11454 , y11455 , y11456 , y11457 , y11458 , y11459 , y11460 , y11461 , y11462 , y11463 , y11464 , y11465 , y11466 , y11467 , y11468 , y11469 , y11470 , y11471 , y11472 , y11473 , y11474 , y11475 , y11476 , y11477 , y11478 , y11479 , y11480 , y11481 , y11482 , y11483 , y11484 , y11485 , y11486 , y11487 , y11488 , y11489 , y11490 , y11491 , y11492 , y11493 , y11494 , y11495 , y11496 , y11497 , y11498 , y11499 , y11500 , y11501 , y11502 , y11503 , y11504 , y11505 , y11506 , y11507 , y11508 , y11509 , y11510 , y11511 , y11512 , y11513 , y11514 , y11515 , y11516 , y11517 , y11518 , y11519 , y11520 , y11521 , y11522 , y11523 , y11524 , y11525 , y11526 , y11527 , y11528 , y11529 , y11530 , y11531 , y11532 , y11533 , y11534 , y11535 , y11536 , y11537 , y11538 , y11539 , y11540 , y11541 , y11542 , y11543 , y11544 , y11545 , y11546 , y11547 , y11548 , y11549 , y11550 , y11551 , y11552 , y11553 , y11554 , y11555 , y11556 , y11557 , y11558 , y11559 , y11560 , y11561 , y11562 , y11563 , y11564 , y11565 , y11566 , y11567 , y11568 , y11569 , y11570 , y11571 , y11572 , y11573 , y11574 , y11575 , y11576 , y11577 , y11578 , y11579 , y11580 , y11581 , y11582 , y11583 , y11584 , y11585 , y11586 , y11587 , y11588 , y11589 , y11590 , y11591 , y11592 , y11593 , y11594 , y11595 , y11596 , y11597 , y11598 , y11599 , y11600 , y11601 , y11602 , y11603 , y11604 , y11605 , y11606 , y11607 , y11608 , y11609 , y11610 , y11611 , y11612 , y11613 , y11614 , y11615 , y11616 , y11617 , y11618 , y11619 , y11620 , y11621 , y11622 , y11623 , y11624 , y11625 , y11626 , y11627 , y11628 , y11629 , y11630 , y11631 , y11632 , y11633 , y11634 , y11635 , y11636 , y11637 , y11638 , y11639 , y11640 , y11641 , y11642 , y11643 , y11644 , y11645 , y11646 , y11647 , y11648 , y11649 , y11650 , y11651 , y11652 , y11653 , y11654 , y11655 , y11656 , y11657 , y11658 , y11659 , y11660 , y11661 , y11662 , y11663 , y11664 , y11665 , y11666 , y11667 , y11668 , y11669 , y11670 , y11671 , y11672 , y11673 , y11674 , y11675 , y11676 , y11677 , y11678 , y11679 , y11680 , y11681 , y11682 , y11683 , y11684 , y11685 , y11686 , y11687 , y11688 , y11689 , y11690 , y11691 , y11692 , y11693 , y11694 , y11695 , y11696 , y11697 , y11698 , y11699 , y11700 , y11701 , y11702 , y11703 , y11704 , y11705 , y11706 , y11707 , y11708 , y11709 , y11710 , y11711 , y11712 , y11713 , y11714 , y11715 , y11716 , y11717 , y11718 , y11719 , y11720 , y11721 , y11722 , y11723 , y11724 , y11725 , y11726 , y11727 , y11728 , y11729 , y11730 , y11731 , y11732 , y11733 , y11734 , y11735 , y11736 , y11737 , y11738 , y11739 , y11740 , y11741 , y11742 , y11743 , y11744 , y11745 , y11746 , y11747 , y11748 , y11749 , y11750 , y11751 , y11752 , y11753 , y11754 , y11755 , y11756 , y11757 , y11758 , y11759 , y11760 , y11761 , y11762 , y11763 , y11764 , y11765 , y11766 , y11767 , y11768 , y11769 , y11770 , y11771 , y11772 , y11773 , y11774 , y11775 , y11776 , y11777 , y11778 , y11779 , y11780 , y11781 , y11782 , y11783 , y11784 , y11785 , y11786 , y11787 , y11788 , y11789 , y11790 , y11791 , y11792 , y11793 , y11794 , y11795 , y11796 , y11797 , y11798 , y11799 , y11800 , y11801 , y11802 , y11803 , y11804 , y11805 , y11806 , y11807 , y11808 , y11809 , y11810 , y11811 , y11812 , y11813 , y11814 , y11815 , y11816 , y11817 , y11818 , y11819 , y11820 , y11821 , y11822 , y11823 , y11824 , y11825 , y11826 , y11827 , y11828 , y11829 , y11830 , y11831 , y11832 , y11833 , y11834 , y11835 , y11836 , y11837 , y11838 , y11839 , y11840 , y11841 , y11842 , y11843 , y11844 , y11845 , y11846 , y11847 , y11848 , y11849 , y11850 , y11851 , y11852 , y11853 , y11854 , y11855 , y11856 , y11857 , y11858 , y11859 , y11860 , y11861 , y11862 , y11863 , y11864 , y11865 , y11866 , y11867 , y11868 , y11869 , y11870 , y11871 , y11872 , y11873 , y11874 , y11875 , y11876 , y11877 , y11878 , y11879 , y11880 , y11881 , y11882 , y11883 , y11884 , y11885 , y11886 , y11887 , y11888 , y11889 , y11890 , y11891 , y11892 , y11893 , y11894 , y11895 , y11896 , y11897 , y11898 , y11899 , y11900 , y11901 , y11902 , y11903 , y11904 , y11905 , y11906 , y11907 , y11908 , y11909 , y11910 , y11911 , y11912 , y11913 , y11914 , y11915 , y11916 , y11917 , y11918 , y11919 , y11920 , y11921 , y11922 , y11923 , y11924 , y11925 , y11926 , y11927 , y11928 , y11929 , y11930 , y11931 , y11932 , y11933 , y11934 , y11935 , y11936 , y11937 , y11938 , y11939 , y11940 , y11941 , y11942 , y11943 , y11944 , y11945 , y11946 , y11947 , y11948 , y11949 , y11950 , y11951 , y11952 , y11953 , y11954 , y11955 , y11956 , y11957 , y11958 , y11959 , y11960 , y11961 , y11962 , y11963 , y11964 , y11965 , y11966 , y11967 , y11968 , y11969 , y11970 , y11971 , y11972 , y11973 , y11974 , y11975 , y11976 , y11977 , y11978 , y11979 , y11980 , y11981 , y11982 , y11983 , y11984 , y11985 , y11986 , y11987 , y11988 , y11989 , y11990 , y11991 , y11992 , y11993 , y11994 , y11995 , y11996 , y11997 , y11998 , y11999 , y12000 , y12001 , y12002 , y12003 , y12004 , y12005 , y12006 , y12007 , y12008 , y12009 , y12010 , y12011 , y12012 , y12013 , y12014 , y12015 , y12016 , y12017 , y12018 , y12019 , y12020 , y12021 , y12022 , y12023 , y12024 , y12025 , y12026 , y12027 , y12028 , y12029 , y12030 , y12031 , y12032 , y12033 , y12034 , y12035 , y12036 , y12037 , y12038 , y12039 , y12040 , y12041 , y12042 , y12043 , y12044 , y12045 , y12046 , y12047 , y12048 , y12049 , y12050 , y12051 , y12052 , y12053 , y12054 , y12055 , y12056 , y12057 , y12058 , y12059 , y12060 , y12061 , y12062 , y12063 , y12064 , y12065 , y12066 , y12067 , y12068 , y12069 , y12070 , y12071 , y12072 , y12073 , y12074 , y12075 , y12076 , y12077 , y12078 , y12079 , y12080 , y12081 , y12082 , y12083 , y12084 , y12085 , y12086 , y12087 , y12088 , y12089 , y12090 , y12091 , y12092 , y12093 , y12094 , y12095 , y12096 , y12097 , y12098 , y12099 , y12100 , y12101 , y12102 , y12103 , y12104 , y12105 , y12106 , y12107 , y12108 , y12109 , y12110 , y12111 , y12112 , y12113 , y12114 , y12115 , y12116 , y12117 , y12118 , y12119 , y12120 , y12121 , y12122 , y12123 , y12124 , y12125 , y12126 , y12127 , y12128 , y12129 , y12130 , y12131 , y12132 , y12133 , y12134 , y12135 , y12136 , y12137 , y12138 , y12139 , y12140 , y12141 , y12142 , y12143 , y12144 , y12145 , y12146 , y12147 , y12148 , y12149 , y12150 , y12151 , y12152 , y12153 , y12154 , y12155 , y12156 , y12157 , y12158 , y12159 , y12160 , y12161 , y12162 , y12163 , y12164 , y12165 , y12166 , y12167 , y12168 , y12169 , y12170 , y12171 , y12172 , y12173 , y12174 , y12175 , y12176 , y12177 , y12178 , y12179 , y12180 , y12181 , y12182 , y12183 , y12184 , y12185 , y12186 , y12187 , y12188 , y12189 , y12190 , y12191 , y12192 , y12193 , y12194 , y12195 , y12196 , y12197 , y12198 , y12199 , y12200 , y12201 , y12202 , y12203 , y12204 , y12205 , y12206 , y12207 , y12208 , y12209 , y12210 , y12211 , y12212 , y12213 , y12214 , y12215 , y12216 , y12217 , y12218 , y12219 , y12220 , y12221 , y12222 , y12223 , y12224 , y12225 , y12226 , y12227 , y12228 , y12229 , y12230 , y12231 , y12232 , y12233 , y12234 , y12235 , y12236 , y12237 , y12238 , y12239 , y12240 , y12241 , y12242 , y12243 , y12244 , y12245 , y12246 , y12247 , y12248 , y12249 , y12250 , y12251 , y12252 , y12253 , y12254 , y12255 , y12256 , y12257 , y12258 , y12259 , y12260 , y12261 , y12262 , y12263 , y12264 , y12265 , y12266 , y12267 , y12268 , y12269 , y12270 , y12271 , y12272 , y12273 , y12274 , y12275 , y12276 , y12277 , y12278 , y12279 , y12280 , y12281 , y12282 , y12283 , y12284 , y12285 , y12286 , y12287 , y12288 , y12289 , y12290 , y12291 , y12292 , y12293 , y12294 , y12295 , y12296 , y12297 , y12298 , y12299 , y12300 , y12301 , y12302 , y12303 , y12304 , y12305 , y12306 , y12307 , y12308 , y12309 , y12310 , y12311 , y12312 , y12313 , y12314 , y12315 , y12316 , y12317 , y12318 , y12319 , y12320 , y12321 , y12322 , y12323 , y12324 , y12325 , y12326 , y12327 , y12328 , y12329 , y12330 , y12331 , y12332 , y12333 , y12334 , y12335 , y12336 , y12337 , y12338 , y12339 , y12340 , y12341 , y12342 , y12343 , y12344 , y12345 , y12346 , y12347 , y12348 , y12349 , y12350 , y12351 , y12352 , y12353 , y12354 , y12355 , y12356 , y12357 , y12358 , y12359 , y12360 , y12361 , y12362 , y12363 , y12364 , y12365 , y12366 , y12367 , y12368 , y12369 , y12370 , y12371 , y12372 , y12373 , y12374 , y12375 , y12376 , y12377 , y12378 , y12379 , y12380 , y12381 , y12382 , y12383 , y12384 , y12385 , y12386 , y12387 , y12388 , y12389 , y12390 , y12391 , y12392 , y12393 , y12394 , y12395 , y12396 , y12397 , y12398 , y12399 , y12400 , y12401 , y12402 , y12403 , y12404 , y12405 , y12406 , y12407 , y12408 , y12409 , y12410 , y12411 , y12412 , y12413 , y12414 , y12415 , y12416 , y12417 , y12418 , y12419 , y12420 , y12421 , y12422 , y12423 , y12424 , y12425 , y12426 , y12427 , y12428 , y12429 , y12430 , y12431 , y12432 , y12433 , y12434 , y12435 , y12436 , y12437 , y12438 , y12439 , y12440 , y12441 , y12442 , y12443 , y12444 , y12445 , y12446 , y12447 , y12448 , y12449 , y12450 , y12451 , y12452 , y12453 , y12454 , y12455 , y12456 , y12457 , y12458 , y12459 , y12460 , y12461 , y12462 , y12463 , y12464 , y12465 , y12466 , y12467 , y12468 , y12469 , y12470 , y12471 , y12472 , y12473 , y12474 , y12475 , y12476 , y12477 , y12478 , y12479 , y12480 , y12481 , y12482 , y12483 , y12484 , y12485 , y12486 , y12487 , y12488 , y12489 , y12490 , y12491 , y12492 , y12493 , y12494 , y12495 , y12496 , y12497 , y12498 , y12499 , y12500 , y12501 , y12502 , y12503 , y12504 , y12505 , y12506 , y12507 , y12508 , y12509 , y12510 , y12511 , y12512 , y12513 , y12514 , y12515 , y12516 , y12517 , y12518 , y12519 , y12520 , y12521 , y12522 , y12523 , y12524 , y12525 , y12526 , y12527 , y12528 , y12529 , y12530 , y12531 , y12532 , y12533 , y12534 , y12535 , y12536 , y12537 , y12538 , y12539 , y12540 , y12541 , y12542 , y12543 , y12544 , y12545 , y12546 , y12547 , y12548 , y12549 , y12550 , y12551 , y12552 , y12553 , y12554 , y12555 , y12556 , y12557 , y12558 , y12559 , y12560 , y12561 , y12562 , y12563 , y12564 , y12565 , y12566 , y12567 , y12568 , y12569 , y12570 , y12571 , y12572 , y12573 , y12574 , y12575 , y12576 , y12577 , y12578 , y12579 , y12580 , y12581 , y12582 , y12583 , y12584 , y12585 , y12586 , y12587 , y12588 , y12589 , y12590 , y12591 , y12592 , y12593 , y12594 , y12595 , y12596 , y12597 , y12598 , y12599 , y12600 , y12601 , y12602 , y12603 , y12604 , y12605 , y12606 , y12607 , y12608 , y12609 , y12610 , y12611 , y12612 , y12613 , y12614 , y12615 , y12616 , y12617 , y12618 , y12619 , y12620 , y12621 , y12622 , y12623 , y12624 , y12625 , y12626 , y12627 , y12628 , y12629 , y12630 , y12631 , y12632 , y12633 , y12634 , y12635 , y12636 , y12637 , y12638 , y12639 , y12640 , y12641 , y12642 , y12643 , y12644 , y12645 , y12646 , y12647 , y12648 , y12649 , y12650 , y12651 , y12652 , y12653 , y12654 , y12655 , y12656 , y12657 , y12658 , y12659 , y12660 , y12661 , y12662 , y12663 , y12664 , y12665 , y12666 , y12667 , y12668 , y12669 , y12670 , y12671 , y12672 , y12673 , y12674 , y12675 , y12676 , y12677 , y12678 , y12679 , y12680 , y12681 , y12682 , y12683 , y12684 , y12685 , y12686 , y12687 , y12688 , y12689 , y12690 , y12691 , y12692 , y12693 , y12694 , y12695 , y12696 , y12697 , y12698 , y12699 , y12700 , y12701 , y12702 , y12703 , y12704 , y12705 , y12706 , y12707 , y12708 , y12709 , y12710 , y12711 , y12712 , y12713 , y12714 , y12715 , y12716 , y12717 , y12718 , y12719 , y12720 , y12721 , y12722 , y12723 , y12724 , y12725 , y12726 , y12727 , y12728 , y12729 , y12730 , y12731 , y12732 , y12733 , y12734 , y12735 , y12736 , y12737 , y12738 , y12739 , y12740 , y12741 , y12742 , y12743 , y12744 , y12745 , y12746 , y12747 , y12748 , y12749 , y12750 , y12751 , y12752 , y12753 , y12754 , y12755 , y12756 , y12757 , y12758 , y12759 , y12760 , y12761 , y12762 , y12763 , y12764 , y12765 , y12766 , y12767 , y12768 , y12769 , y12770 , y12771 , y12772 , y12773 , y12774 , y12775 , y12776 , y12777 , y12778 , y12779 , y12780 , y12781 , y12782 , y12783 , y12784 , y12785 , y12786 , y12787 , y12788 , y12789 , y12790 , y12791 , y12792 , y12793 , y12794 , y12795 , y12796 , y12797 , y12798 , y12799 , y12800 , y12801 , y12802 , y12803 , y12804 , y12805 , y12806 , y12807 , y12808 , y12809 , y12810 , y12811 , y12812 , y12813 , y12814 , y12815 , y12816 , y12817 , y12818 , y12819 , y12820 , y12821 , y12822 , y12823 , y12824 , y12825 , y12826 , y12827 , y12828 , y12829 , y12830 , y12831 , y12832 , y12833 , y12834 , y12835 , y12836 , y12837 , y12838 , y12839 , y12840 , y12841 , y12842 , y12843 , y12844 , y12845 , y12846 , y12847 , y12848 , y12849 , y12850 , y12851 , y12852 , y12853 , y12854 , y12855 , y12856 , y12857 , y12858 , y12859 , y12860 , y12861 , y12862 , y12863 , y12864 , y12865 , y12866 , y12867 , y12868 , y12869 , y12870 , y12871 , y12872 , y12873 , y12874 , y12875 , y12876 , y12877 , y12878 , y12879 , y12880 , y12881 , y12882 , y12883 , y12884 , y12885 , y12886 , y12887 , y12888 , y12889 , y12890 , y12891 , y12892 , y12893 , y12894 , y12895 , y12896 , y12897 , y12898 , y12899 , y12900 , y12901 , y12902 , y12903 , y12904 , y12905 , y12906 , y12907 , y12908 , y12909 , y12910 , y12911 , y12912 , y12913 , y12914 , y12915 , y12916 , y12917 , y12918 , y12919 , y12920 , y12921 , y12922 , y12923 , y12924 , y12925 , y12926 , y12927 , y12928 , y12929 , y12930 , y12931 , y12932 , y12933 , y12934 , y12935 , y12936 , y12937 , y12938 , y12939 , y12940 , y12941 , y12942 , y12943 , y12944 , y12945 , y12946 , y12947 , y12948 , y12949 , y12950 , y12951 , y12952 , y12953 , y12954 , y12955 , y12956 , y12957 , y12958 , y12959 , y12960 , y12961 , y12962 , y12963 , y12964 , y12965 , y12966 , y12967 , y12968 , y12969 , y12970 , y12971 , y12972 , y12973 , y12974 , y12975 , y12976 , y12977 , y12978 , y12979 , y12980 , y12981 , y12982 , y12983 , y12984 , y12985 , y12986 , y12987 , y12988 , y12989 , y12990 , y12991 , y12992 , y12993 , y12994 , y12995 , y12996 , y12997 , y12998 , y12999 , y13000 , y13001 , y13002 , y13003 , y13004 , y13005 , y13006 , y13007 , y13008 , y13009 , y13010 , y13011 , y13012 , y13013 , y13014 , y13015 , y13016 , y13017 , y13018 , y13019 , y13020 , y13021 , y13022 , y13023 , y13024 , y13025 , y13026 , y13027 , y13028 , y13029 , y13030 , y13031 , y13032 , y13033 , y13034 , y13035 , y13036 , y13037 , y13038 , y13039 , y13040 , y13041 , y13042 , y13043 , y13044 , y13045 , y13046 , y13047 , y13048 , y13049 , y13050 , y13051 , y13052 , y13053 , y13054 , y13055 , y13056 , y13057 , y13058 , y13059 , y13060 , y13061 , y13062 , y13063 , y13064 , y13065 , y13066 , y13067 , y13068 , y13069 , y13070 , y13071 , y13072 , y13073 , y13074 , y13075 , y13076 , y13077 , y13078 , y13079 , y13080 , y13081 , y13082 , y13083 , y13084 , y13085 , y13086 , y13087 , y13088 , y13089 , y13090 , y13091 , y13092 , y13093 , y13094 , y13095 , y13096 , y13097 , y13098 , y13099 , y13100 , y13101 , y13102 , y13103 , y13104 , y13105 , y13106 , y13107 , y13108 , y13109 , y13110 , y13111 , y13112 , y13113 , y13114 , y13115 , y13116 , y13117 , y13118 , y13119 , y13120 , y13121 , y13122 , y13123 , y13124 , y13125 , y13126 , y13127 , y13128 , y13129 , y13130 , y13131 , y13132 , y13133 , y13134 , y13135 , y13136 , y13137 , y13138 , y13139 , y13140 , y13141 , y13142 , y13143 , y13144 , y13145 , y13146 , y13147 , y13148 , y13149 , y13150 , y13151 , y13152 , y13153 , y13154 , y13155 , y13156 , y13157 , y13158 , y13159 , y13160 , y13161 , y13162 , y13163 , y13164 , y13165 , y13166 , y13167 , y13168 , y13169 , y13170 , y13171 , y13172 , y13173 , y13174 , y13175 , y13176 , y13177 , y13178 , y13179 , y13180 , y13181 , y13182 , y13183 , y13184 , y13185 , y13186 , y13187 , y13188 , y13189 , y13190 , y13191 , y13192 , y13193 , y13194 , y13195 , y13196 , y13197 , y13198 , y13199 , y13200 , y13201 , y13202 , y13203 , y13204 , y13205 , y13206 , y13207 , y13208 , y13209 , y13210 , y13211 , y13212 , y13213 , y13214 , y13215 , y13216 , y13217 , y13218 , y13219 , y13220 , y13221 , y13222 , y13223 , y13224 , y13225 , y13226 , y13227 , y13228 , y13229 , y13230 , y13231 , y13232 , y13233 , y13234 , y13235 , y13236 , y13237 , y13238 , y13239 , y13240 , y13241 , y13242 , y13243 , y13244 , y13245 , y13246 , y13247 , y13248 , y13249 , y13250 , y13251 , y13252 , y13253 , y13254 , y13255 , y13256 , y13257 , y13258 , y13259 , y13260 , y13261 , y13262 , y13263 , y13264 , y13265 , y13266 , y13267 , y13268 , y13269 , y13270 , y13271 , y13272 , y13273 , y13274 , y13275 , y13276 , y13277 , y13278 , y13279 , y13280 , y13281 , y13282 , y13283 , y13284 , y13285 , y13286 , y13287 , y13288 , y13289 , y13290 , y13291 , y13292 , y13293 , y13294 , y13295 , y13296 , y13297 , y13298 , y13299 , y13300 , y13301 , y13302 , y13303 , y13304 , y13305 , y13306 , y13307 , y13308 , y13309 , y13310 , y13311 , y13312 , y13313 , y13314 , y13315 , y13316 , y13317 , y13318 , y13319 , y13320 , y13321 , y13322 , y13323 , y13324 , y13325 , y13326 , y13327 , y13328 , y13329 , y13330 , y13331 , y13332 , y13333 , y13334 , y13335 , y13336 , y13337 , y13338 , y13339 , y13340 , y13341 , y13342 , y13343 , y13344 , y13345 , y13346 , y13347 , y13348 , y13349 , y13350 , y13351 , y13352 , y13353 , y13354 , y13355 , y13356 , y13357 , y13358 , y13359 , y13360 , y13361 , y13362 , y13363 , y13364 , y13365 , y13366 , y13367 , y13368 , y13369 , y13370 , y13371 , y13372 , y13373 , y13374 , y13375 , y13376 , y13377 , y13378 , y13379 , y13380 , y13381 , y13382 , y13383 , y13384 , y13385 , y13386 , y13387 , y13388 , y13389 , y13390 , y13391 , y13392 , y13393 , y13394 , y13395 , y13396 , y13397 , y13398 , y13399 , y13400 , y13401 , y13402 , y13403 , y13404 , y13405 , y13406 , y13407 , y13408 , y13409 , y13410 , y13411 , y13412 , y13413 , y13414 , y13415 , y13416 , y13417 , y13418 , y13419 , y13420 , y13421 , y13422 , y13423 , y13424 , y13425 , y13426 , y13427 , y13428 , y13429 , y13430 , y13431 , y13432 , y13433 , y13434 , y13435 , y13436 , y13437 , y13438 , y13439 , y13440 , y13441 , y13442 , y13443 , y13444 , y13445 , y13446 , y13447 , y13448 , y13449 , y13450 , y13451 , y13452 , y13453 , y13454 , y13455 , y13456 , y13457 , y13458 , y13459 , y13460 , y13461 , y13462 , y13463 , y13464 , y13465 , y13466 , y13467 , y13468 , y13469 , y13470 , y13471 , y13472 , y13473 , y13474 , y13475 , y13476 , y13477 , y13478 , y13479 , y13480 , y13481 , y13482 , y13483 , y13484 , y13485 , y13486 , y13487 , y13488 , y13489 , y13490 , y13491 , y13492 , y13493 , y13494 , y13495 , y13496 , y13497 , y13498 , y13499 , y13500 , y13501 , y13502 , y13503 , y13504 , y13505 , y13506 , y13507 , y13508 , y13509 , y13510 , y13511 , y13512 , y13513 , y13514 , y13515 , y13516 , y13517 , y13518 , y13519 , y13520 , y13521 , y13522 , y13523 , y13524 , y13525 , y13526 , y13527 , y13528 , y13529 , y13530 , y13531 , y13532 , y13533 , y13534 , y13535 , y13536 , y13537 , y13538 , y13539 , y13540 , y13541 , y13542 , y13543 , y13544 , y13545 , y13546 , y13547 , y13548 , y13549 , y13550 , y13551 , y13552 , y13553 , y13554 , y13555 , y13556 , y13557 , y13558 , y13559 , y13560 , y13561 , y13562 , y13563 , y13564 , y13565 , y13566 , y13567 , y13568 , y13569 , y13570 , y13571 , y13572 , y13573 , y13574 , y13575 , y13576 , y13577 , y13578 , y13579 , y13580 , y13581 , y13582 , y13583 , y13584 , y13585 , y13586 , y13587 , y13588 , y13589 , y13590 , y13591 , y13592 , y13593 , y13594 , y13595 , y13596 , y13597 , y13598 , y13599 , y13600 , y13601 , y13602 , y13603 , y13604 , y13605 , y13606 , y13607 , y13608 , y13609 , y13610 , y13611 , y13612 , y13613 , y13614 , y13615 , y13616 , y13617 , y13618 , y13619 , y13620 , y13621 , y13622 , y13623 , y13624 , y13625 , y13626 , y13627 , y13628 , y13629 , y13630 , y13631 , y13632 , y13633 , y13634 , y13635 , y13636 , y13637 , y13638 , y13639 , y13640 , y13641 , y13642 , y13643 , y13644 , y13645 , y13646 , y13647 , y13648 , y13649 , y13650 , y13651 , y13652 , y13653 , y13654 , y13655 , y13656 , y13657 , y13658 , y13659 , y13660 , y13661 , y13662 , y13663 , y13664 , y13665 , y13666 , y13667 , y13668 , y13669 , y13670 , y13671 , y13672 , y13673 , y13674 , y13675 , y13676 , y13677 , y13678 , y13679 , y13680 , y13681 , y13682 , y13683 , y13684 , y13685 , y13686 , y13687 , y13688 , y13689 , y13690 , y13691 , y13692 , y13693 , y13694 , y13695 , y13696 , y13697 , y13698 , y13699 , y13700 , y13701 , y13702 , y13703 , y13704 , y13705 , y13706 , y13707 , y13708 , y13709 , y13710 , y13711 , y13712 , y13713 , y13714 , y13715 , y13716 , y13717 , y13718 , y13719 , y13720 , y13721 , y13722 , y13723 , y13724 , y13725 , y13726 , y13727 , y13728 , y13729 , y13730 , y13731 , y13732 , y13733 , y13734 , y13735 , y13736 , y13737 , y13738 , y13739 , y13740 , y13741 , y13742 , y13743 , y13744 , y13745 , y13746 , y13747 , y13748 , y13749 , y13750 , y13751 , y13752 , y13753 , y13754 , y13755 , y13756 , y13757 , y13758 , y13759 , y13760 , y13761 , y13762 , y13763 , y13764 , y13765 , y13766 , y13767 , y13768 , y13769 , y13770 , y13771 , y13772 , y13773 , y13774 , y13775 , y13776 , y13777 , y13778 , y13779 , y13780 , y13781 , y13782 , y13783 , y13784 , y13785 , y13786 , y13787 , y13788 , y13789 , y13790 , y13791 , y13792 , y13793 , y13794 , y13795 , y13796 , y13797 , y13798 , y13799 , y13800 , y13801 , y13802 , y13803 , y13804 , y13805 , y13806 , y13807 , y13808 , y13809 , y13810 , y13811 , y13812 , y13813 , y13814 , y13815 , y13816 , y13817 , y13818 , y13819 , y13820 , y13821 , y13822 , y13823 , y13824 , y13825 , y13826 , y13827 , y13828 , y13829 , y13830 , y13831 , y13832 , y13833 , y13834 , y13835 , y13836 , y13837 , y13838 , y13839 , y13840 , y13841 , y13842 , y13843 , y13844 , y13845 , y13846 , y13847 , y13848 , y13849 , y13850 , y13851 , y13852 , y13853 , y13854 , y13855 , y13856 , y13857 , y13858 , y13859 , y13860 , y13861 , y13862 , y13863 , y13864 , y13865 , y13866 , y13867 , y13868 , y13869 , y13870 , y13871 , y13872 , y13873 , y13874 , y13875 , y13876 , y13877 , y13878 , y13879 , y13880 , y13881 , y13882 , y13883 , y13884 , y13885 , y13886 , y13887 , y13888 , y13889 , y13890 , y13891 , y13892 , y13893 , y13894 , y13895 , y13896 , y13897 , y13898 , y13899 , y13900 , y13901 , y13902 , y13903 , y13904 , y13905 , y13906 , y13907 , y13908 , y13909 , y13910 , y13911 , y13912 , y13913 , y13914 , y13915 , y13916 , y13917 , y13918 , y13919 , y13920 , y13921 , y13922 , y13923 , y13924 , y13925 , y13926 , y13927 , y13928 , y13929 , y13930 , y13931 , y13932 , y13933 , y13934 , y13935 , y13936 , y13937 , y13938 , y13939 , y13940 , y13941 , y13942 , y13943 , y13944 , y13945 , y13946 , y13947 , y13948 , y13949 , y13950 , y13951 , y13952 , y13953 , y13954 , y13955 , y13956 , y13957 , y13958 , y13959 , y13960 , y13961 , y13962 , y13963 , y13964 , y13965 , y13966 , y13967 , y13968 , y13969 , y13970 , y13971 , y13972 , y13973 , y13974 , y13975 , y13976 , y13977 , y13978 , y13979 , y13980 , y13981 , y13982 , y13983 , y13984 , y13985 , y13986 , y13987 , y13988 , y13989 , y13990 , y13991 , y13992 , y13993 , y13994 , y13995 , y13996 , y13997 , y13998 , y13999 , y14000 , y14001 , y14002 , y14003 , y14004 , y14005 , y14006 , y14007 , y14008 , y14009 , y14010 , y14011 , y14012 , y14013 , y14014 , y14015 , y14016 , y14017 , y14018 , y14019 , y14020 , y14021 , y14022 , y14023 , y14024 , y14025 , y14026 , y14027 , y14028 , y14029 , y14030 , y14031 , y14032 , y14033 , y14034 , y14035 , y14036 , y14037 , y14038 , y14039 , y14040 , y14041 , y14042 , y14043 , y14044 , y14045 , y14046 , y14047 , y14048 , y14049 , y14050 , y14051 , y14052 , y14053 , y14054 , y14055 , y14056 , y14057 , y14058 , y14059 , y14060 , y14061 , y14062 , y14063 , y14064 , y14065 , y14066 , y14067 , y14068 , y14069 , y14070 , y14071 , y14072 , y14073 , y14074 , y14075 , y14076 , y14077 , y14078 , y14079 , y14080 , y14081 , y14082 , y14083 , y14084 , y14085 , y14086 , y14087 , y14088 , y14089 , y14090 , y14091 , y14092 , y14093 , y14094 , y14095 , y14096 , y14097 , y14098 , y14099 , y14100 , y14101 , y14102 , y14103 , y14104 , y14105 , y14106 , y14107 , y14108 , y14109 , y14110 , y14111 , y14112 , y14113 , y14114 , y14115 , y14116 , y14117 , y14118 , y14119 , y14120 , y14121 , y14122 , y14123 , y14124 , y14125 , y14126 , y14127 , y14128 , y14129 , y14130 , y14131 , y14132 , y14133 , y14134 , y14135 , y14136 , y14137 , y14138 , y14139 , y14140 , y14141 , y14142 , y14143 , y14144 , y14145 , y14146 , y14147 , y14148 , y14149 , y14150 , y14151 , y14152 , y14153 , y14154 , y14155 , y14156 , y14157 , y14158 , y14159 , y14160 , y14161 , y14162 , y14163 , y14164 , y14165 , y14166 , y14167 , y14168 , y14169 , y14170 , y14171 , y14172 , y14173 , y14174 , y14175 , y14176 , y14177 , y14178 , y14179 , y14180 , y14181 , y14182 , y14183 , y14184 , y14185 , y14186 , y14187 , y14188 , y14189 , y14190 , y14191 , y14192 , y14193 , y14194 , y14195 , y14196 , y14197 , y14198 , y14199 , y14200 , y14201 , y14202 , y14203 , y14204 , y14205 , y14206 , y14207 , y14208 , y14209 , y14210 , y14211 , y14212 , y14213 , y14214 , y14215 , y14216 , y14217 , y14218 , y14219 , y14220 , y14221 , y14222 , y14223 , y14224 , y14225 , y14226 , y14227 , y14228 , y14229 , y14230 , y14231 , y14232 , y14233 , y14234 , y14235 , y14236 , y14237 , y14238 , y14239 , y14240 , y14241 , y14242 , y14243 , y14244 , y14245 , y14246 , y14247 , y14248 , y14249 , y14250 , y14251 , y14252 , y14253 , y14254 , y14255 , y14256 , y14257 , y14258 , y14259 , y14260 , y14261 , y14262 , y14263 , y14264 , y14265 , y14266 , y14267 , y14268 , y14269 , y14270 , y14271 , y14272 , y14273 , y14274 , y14275 , y14276 , y14277 , y14278 , y14279 , y14280 , y14281 , y14282 , y14283 , y14284 , y14285 , y14286 , y14287 , y14288 , y14289 , y14290 , y14291 , y14292 , y14293 , y14294 , y14295 , y14296 , y14297 , y14298 , y14299 , y14300 , y14301 , y14302 , y14303 , y14304 , y14305 , y14306 , y14307 , y14308 , y14309 , y14310 , y14311 , y14312 , y14313 , y14314 , y14315 , y14316 , y14317 , y14318 , y14319 , y14320 , y14321 , y14322 , y14323 , y14324 , y14325 , y14326 , y14327 , y14328 , y14329 , y14330 , y14331 , y14332 , y14333 , y14334 , y14335 , y14336 , y14337 , y14338 , y14339 , y14340 , y14341 , y14342 , y14343 , y14344 , y14345 , y14346 , y14347 , y14348 , y14349 , y14350 , y14351 , y14352 , y14353 , y14354 , y14355 , y14356 , y14357 , y14358 , y14359 , y14360 , y14361 , y14362 , y14363 , y14364 , y14365 , y14366 , y14367 , y14368 , y14369 , y14370 , y14371 , y14372 , y14373 , y14374 , y14375 , y14376 , y14377 , y14378 , y14379 , y14380 , y14381 , y14382 , y14383 , y14384 , y14385 , y14386 , y14387 , y14388 , y14389 , y14390 , y14391 , y14392 , y14393 , y14394 , y14395 , y14396 , y14397 , y14398 , y14399 , y14400 , y14401 , y14402 , y14403 , y14404 , y14405 , y14406 , y14407 , y14408 , y14409 , y14410 , y14411 , y14412 , y14413 , y14414 , y14415 , y14416 , y14417 , y14418 , y14419 , y14420 , y14421 , y14422 , y14423 , y14424 , y14425 , y14426 , y14427 , y14428 , y14429 , y14430 , y14431 , y14432 , y14433 , y14434 , y14435 , y14436 , y14437 , y14438 , y14439 , y14440 , y14441 , y14442 , y14443 , y14444 , y14445 , y14446 , y14447 , y14448 , y14449 , y14450 , y14451 , y14452 , y14453 , y14454 , y14455 , y14456 , y14457 , y14458 , y14459 , y14460 , y14461 , y14462 , y14463 , y14464 , y14465 , y14466 , y14467 , y14468 , y14469 , y14470 , y14471 , y14472 , y14473 , y14474 , y14475 , y14476 , y14477 , y14478 , y14479 , y14480 , y14481 , y14482 , y14483 , y14484 , y14485 , y14486 , y14487 , y14488 , y14489 , y14490 , y14491 , y14492 , y14493 , y14494 , y14495 , y14496 , y14497 , y14498 , y14499 , y14500 , y14501 , y14502 , y14503 , y14504 , y14505 , y14506 , y14507 , y14508 , y14509 , y14510 , y14511 , y14512 , y14513 , y14514 , y14515 , y14516 , y14517 , y14518 , y14519 , y14520 , y14521 , y14522 , y14523 , y14524 , y14525 , y14526 , y14527 , y14528 , y14529 , y14530 , y14531 , y14532 , y14533 , y14534 , y14535 , y14536 , y14537 , y14538 , y14539 , y14540 , y14541 , y14542 , y14543 , y14544 , y14545 , y14546 , y14547 , y14548 , y14549 , y14550 , y14551 , y14552 , y14553 , y14554 , y14555 , y14556 , y14557 , y14558 , y14559 , y14560 , y14561 , y14562 , y14563 , y14564 , y14565 , y14566 , y14567 , y14568 , y14569 , y14570 , y14571 , y14572 , y14573 , y14574 , y14575 , y14576 , y14577 , y14578 , y14579 , y14580 , y14581 , y14582 , y14583 , y14584 , y14585 , y14586 , y14587 , y14588 , y14589 , y14590 , y14591 , y14592 , y14593 , y14594 , y14595 , y14596 , y14597 , y14598 , y14599 , y14600 , y14601 , y14602 , y14603 , y14604 , y14605 , y14606 , y14607 , y14608 , y14609 , y14610 , y14611 , y14612 , y14613 , y14614 , y14615 , y14616 , y14617 , y14618 , y14619 , y14620 , y14621 , y14622 , y14623 , y14624 , y14625 , y14626 , y14627 , y14628 , y14629 , y14630 , y14631 , y14632 , y14633 , y14634 , y14635 , y14636 , y14637 , y14638 , y14639 , y14640 , y14641 , y14642 , y14643 , y14644 , y14645 , y14646 , y14647 , y14648 , y14649 , y14650 , y14651 , y14652 , y14653 , y14654 , y14655 , y14656 , y14657 , y14658 , y14659 , y14660 , y14661 , y14662 , y14663 , y14664 , y14665 , y14666 , y14667 , y14668 , y14669 , y14670 , y14671 , y14672 , y14673 , y14674 , y14675 , y14676 , y14677 , y14678 , y14679 , y14680 , y14681 , y14682 , y14683 , y14684 , y14685 , y14686 , y14687 , y14688 , y14689 , y14690 , y14691 , y14692 , y14693 , y14694 , y14695 , y14696 , y14697 , y14698 , y14699 , y14700 , y14701 , y14702 , y14703 , y14704 , y14705 , y14706 , y14707 , y14708 , y14709 , y14710 , y14711 , y14712 , y14713 , y14714 , y14715 , y14716 , y14717 , y14718 , y14719 , y14720 , y14721 , y14722 , y14723 , y14724 , y14725 , y14726 , y14727 , y14728 , y14729 , y14730 , y14731 , y14732 , y14733 , y14734 , y14735 , y14736 , y14737 , y14738 , y14739 , y14740 , y14741 , y14742 , y14743 , y14744 , y14745 , y14746 , y14747 , y14748 , y14749 , y14750 , y14751 , y14752 , y14753 , y14754 , y14755 , y14756 , y14757 , y14758 , y14759 , y14760 , y14761 , y14762 , y14763 , y14764 , y14765 , y14766 , y14767 , y14768 , y14769 , y14770 , y14771 , y14772 , y14773 , y14774 , y14775 , y14776 , y14777 , y14778 , y14779 , y14780 , y14781 , y14782 , y14783 , y14784 , y14785 , y14786 , y14787 , y14788 , y14789 , y14790 , y14791 , y14792 , y14793 , y14794 , y14795 , y14796 , y14797 , y14798 , y14799 , y14800 , y14801 , y14802 , y14803 , y14804 , y14805 , y14806 , y14807 , y14808 , y14809 , y14810 , y14811 , y14812 , y14813 , y14814 , y14815 , y14816 , y14817 , y14818 , y14819 , y14820 , y14821 , y14822 , y14823 , y14824 , y14825 , y14826 , y14827 , y14828 , y14829 , y14830 , y14831 , y14832 , y14833 , y14834 , y14835 , y14836 , y14837 , y14838 , y14839 , y14840 , y14841 , y14842 , y14843 , y14844 , y14845 , y14846 , y14847 , y14848 , y14849 , y14850 , y14851 , y14852 , y14853 , y14854 , y14855 , y14856 , y14857 , y14858 , y14859 , y14860 , y14861 , y14862 , y14863 , y14864 , y14865 , y14866 , y14867 , y14868 , y14869 , y14870 , y14871 , y14872 , y14873 , y14874 , y14875 , y14876 , y14877 , y14878 , y14879 , y14880 , y14881 , y14882 , y14883 , y14884 , y14885 , y14886 , y14887 , y14888 , y14889 , y14890 , y14891 , y14892 , y14893 , y14894 , y14895 , y14896 , y14897 , y14898 , y14899 , y14900 , y14901 , y14902 , y14903 , y14904 , y14905 , y14906 , y14907 , y14908 , y14909 , y14910 , y14911 , y14912 , y14913 , y14914 , y14915 , y14916 , y14917 , y14918 , y14919 , y14920 , y14921 , y14922 , y14923 , y14924 , y14925 , y14926 , y14927 , y14928 , y14929 , y14930 , y14931 , y14932 , y14933 , y14934 , y14935 , y14936 , y14937 , y14938 , y14939 , y14940 , y14941 , y14942 , y14943 , y14944 , y14945 , y14946 , y14947 , y14948 , y14949 , y14950 , y14951 , y14952 , y14953 , y14954 , y14955 , y14956 , y14957 , y14958 , y14959 , y14960 , y14961 , y14962 , y14963 , y14964 , y14965 , y14966 , y14967 , y14968 , y14969 , y14970 , y14971 , y14972 , y14973 , y14974 , y14975 , y14976 , y14977 , y14978 , y14979 , y14980 , y14981 , y14982 , y14983 , y14984 , y14985 , y14986 , y14987 , y14988 , y14989 , y14990 , y14991 , y14992 , y14993 , y14994 , y14995 , y14996 , y14997 , y14998 , y14999 , y15000 , y15001 , y15002 , y15003 , y15004 , y15005 , y15006 , y15007 , y15008 , y15009 , y15010 , y15011 , y15012 , y15013 , y15014 , y15015 , y15016 , y15017 , y15018 , y15019 , y15020 , y15021 , y15022 , y15023 , y15024 , y15025 , y15026 , y15027 , y15028 , y15029 , y15030 , y15031 , y15032 , y15033 , y15034 , y15035 , y15036 , y15037 , y15038 , y15039 , y15040 , y15041 , y15042 , y15043 , y15044 , y15045 , y15046 , y15047 , y15048 , y15049 , y15050 , y15051 , y15052 , y15053 , y15054 , y15055 , y15056 , y15057 , y15058 , y15059 , y15060 , y15061 , y15062 , y15063 , y15064 , y15065 , y15066 , y15067 , y15068 , y15069 , y15070 , y15071 , y15072 , y15073 , y15074 , y15075 , y15076 , y15077 , y15078 , y15079 , y15080 , y15081 , y15082 , y15083 , y15084 , y15085 , y15086 , y15087 , y15088 , y15089 , y15090 , y15091 , y15092 , y15093 , y15094 , y15095 , y15096 , y15097 , y15098 , y15099 , y15100 , y15101 , y15102 , y15103 , y15104 , y15105 , y15106 , y15107 , y15108 , y15109 , y15110 , y15111 , y15112 , y15113 , y15114 , y15115 , y15116 , y15117 , y15118 , y15119 , y15120 , y15121 , y15122 , y15123 , y15124 , y15125 , y15126 , y15127 , y15128 , y15129 , y15130 , y15131 , y15132 , y15133 , y15134 , y15135 , y15136 , y15137 , y15138 , y15139 , y15140 , y15141 , y15142 , y15143 , y15144 , y15145 , y15146 , y15147 , y15148 , y15149 , y15150 , y15151 , y15152 , y15153 , y15154 , y15155 , y15156 , y15157 , y15158 , y15159 , y15160 , y15161 , y15162 , y15163 , y15164 , y15165 , y15166 , y15167 , y15168 , y15169 , y15170 , y15171 , y15172 , y15173 , y15174 , y15175 , y15176 , y15177 , y15178 , y15179 , y15180 , y15181 , y15182 , y15183 , y15184 , y15185 , y15186 , y15187 , y15188 , y15189 , y15190 , y15191 , y15192 , y15193 , y15194 , y15195 , y15196 , y15197 , y15198 , y15199 , y15200 , y15201 , y15202 , y15203 , y15204 , y15205 , y15206 , y15207 , y15208 , y15209 , y15210 , y15211 , y15212 , y15213 , y15214 , y15215 , y15216 , y15217 , y15218 , y15219 , y15220 , y15221 , y15222 , y15223 , y15224 , y15225 , y15226 , y15227 , y15228 , y15229 , y15230 , y15231 , y15232 , y15233 , y15234 , y15235 , y15236 , y15237 , y15238 , y15239 , y15240 , y15241 , y15242 , y15243 , y15244 , y15245 , y15246 , y15247 , y15248 , y15249 , y15250 , y15251 , y15252 , y15253 , y15254 , y15255 , y15256 , y15257 , y15258 , y15259 , y15260 , y15261 , y15262 , y15263 , y15264 , y15265 , y15266 , y15267 , y15268 , y15269 , y15270 , y15271 , y15272 , y15273 , y15274 , y15275 , y15276 , y15277 , y15278 , y15279 , y15280 , y15281 , y15282 , y15283 , y15284 , y15285 , y15286 , y15287 , y15288 , y15289 , y15290 , y15291 , y15292 , y15293 , y15294 , y15295 , y15296 , y15297 , y15298 , y15299 , y15300 , y15301 , y15302 , y15303 , y15304 , y15305 , y15306 , y15307 , y15308 , y15309 , y15310 , y15311 , y15312 , y15313 , y15314 , y15315 , y15316 , y15317 , y15318 , y15319 , y15320 , y15321 , y15322 , y15323 , y15324 , y15325 , y15326 , y15327 , y15328 , y15329 , y15330 , y15331 , y15332 , y15333 , y15334 , y15335 , y15336 , y15337 , y15338 , y15339 , y15340 , y15341 , y15342 , y15343 , y15344 , y15345 , y15346 , y15347 , y15348 , y15349 , y15350 , y15351 , y15352 , y15353 , y15354 , y15355 , y15356 , y15357 , y15358 , y15359 , y15360 , y15361 , y15362 , y15363 , y15364 , y15365 , y15366 , y15367 , y15368 , y15369 , y15370 , y15371 , y15372 , y15373 , y15374 , y15375 , y15376 , y15377 , y15378 , y15379 , y15380 , y15381 , y15382 , y15383 , y15384 , y15385 , y15386 , y15387 , y15388 , y15389 , y15390 , y15391 , y15392 , y15393 , y15394 , y15395 , y15396 , y15397 , y15398 , y15399 , y15400 , y15401 , y15402 , y15403 , y15404 , y15405 , y15406 , y15407 , y15408 , y15409 , y15410 , y15411 , y15412 , y15413 , y15414 , y15415 , y15416 , y15417 , y15418 , y15419 , y15420 , y15421 , y15422 , y15423 , y15424 , y15425 , y15426 , y15427 , y15428 , y15429 , y15430 , y15431 , y15432 , y15433 , y15434 , y15435 , y15436 , y15437 , y15438 , y15439 , y15440 , y15441 , y15442 , y15443 , y15444 , y15445 , y15446 , y15447 , y15448 , y15449 , y15450 , y15451 , y15452 , y15453 , y15454 , y15455 , y15456 , y15457 , y15458 , y15459 , y15460 , y15461 , y15462 , y15463 , y15464 , y15465 , y15466 , y15467 , y15468 , y15469 , y15470 , y15471 , y15472 , y15473 , y15474 , y15475 , y15476 , y15477 , y15478 , y15479 , y15480 , y15481 , y15482 , y15483 , y15484 , y15485 , y15486 , y15487 , y15488 , y15489 , y15490 , y15491 , y15492 , y15493 , y15494 , y15495 , y15496 , y15497 , y15498 , y15499 , y15500 , y15501 , y15502 , y15503 , y15504 , y15505 , y15506 , y15507 , y15508 , y15509 , y15510 , y15511 , y15512 , y15513 , y15514 , y15515 , y15516 , y15517 , y15518 , y15519 , y15520 , y15521 , y15522 , y15523 , y15524 , y15525 , y15526 , y15527 , y15528 , y15529 , y15530 , y15531 , y15532 , y15533 , y15534 , y15535 , y15536 , y15537 , y15538 , y15539 , y15540 , y15541 , y15542 , y15543 , y15544 , y15545 , y15546 , y15547 , y15548 , y15549 , y15550 , y15551 , y15552 , y15553 , y15554 , y15555 , y15556 , y15557 , y15558 , y15559 , y15560 , y15561 , y15562 , y15563 , y15564 , y15565 , y15566 , y15567 , y15568 , y15569 , y15570 , y15571 , y15572 , y15573 , y15574 , y15575 , y15576 , y15577 , y15578 , y15579 , y15580 , y15581 , y15582 , y15583 , y15584 , y15585 , y15586 , y15587 , y15588 , y15589 , y15590 , y15591 , y15592 , y15593 , y15594 , y15595 , y15596 , y15597 , y15598 , y15599 , y15600 , y15601 , y15602 , y15603 , y15604 , y15605 , y15606 , y15607 , y15608 , y15609 , y15610 , y15611 , y15612 , y15613 , y15614 , y15615 , y15616 , y15617 , y15618 , y15619 , y15620 , y15621 , y15622 , y15623 , y15624 , y15625 , y15626 , y15627 , y15628 , y15629 , y15630 , y15631 , y15632 , y15633 , y15634 , y15635 , y15636 , y15637 , y15638 , y15639 , y15640 , y15641 , y15642 , y15643 , y15644 , y15645 , y15646 , y15647 , y15648 , y15649 , y15650 , y15651 , y15652 , y15653 , y15654 , y15655 , y15656 , y15657 , y15658 , y15659 , y15660 , y15661 , y15662 , y15663 , y15664 , y15665 , y15666 , y15667 , y15668 , y15669 , y15670 , y15671 , y15672 , y15673 , y15674 , y15675 , y15676 , y15677 , y15678 , y15679 , y15680 , y15681 , y15682 , y15683 , y15684 , y15685 , y15686 , y15687 , y15688 , y15689 , y15690 , y15691 , y15692 , y15693 , y15694 , y15695 , y15696 , y15697 , y15698 , y15699 , y15700 , y15701 , y15702 , y15703 , y15704 , y15705 , y15706 , y15707 , y15708 , y15709 , y15710 , y15711 , y15712 , y15713 , y15714 , y15715 , y15716 , y15717 , y15718 , y15719 , y15720 , y15721 , y15722 , y15723 , y15724 , y15725 , y15726 , y15727 , y15728 , y15729 , y15730 , y15731 , y15732 , y15733 , y15734 , y15735 , y15736 , y15737 , y15738 , y15739 , y15740 , y15741 , y15742 , y15743 , y15744 , y15745 , y15746 , y15747 , y15748 , y15749 , y15750 , y15751 , y15752 , y15753 , y15754 , y15755 , y15756 , y15757 , y15758 , y15759 , y15760 , y15761 , y15762 , y15763 , y15764 , y15765 , y15766 , y15767 , y15768 , y15769 , y15770 , y15771 , y15772 , y15773 , y15774 , y15775 , y15776 , y15777 , y15778 , y15779 , y15780 , y15781 , y15782 , y15783 , y15784 , y15785 , y15786 , y15787 , y15788 , y15789 , y15790 , y15791 , y15792 , y15793 , y15794 , y15795 , y15796 , y15797 , y15798 , y15799 , y15800 , y15801 , y15802 , y15803 , y15804 , y15805 , y15806 , y15807 , y15808 , y15809 , y15810 , y15811 , y15812 , y15813 , y15814 , y15815 , y15816 , y15817 , y15818 , y15819 , y15820 , y15821 , y15822 , y15823 , y15824 , y15825 , y15826 , y15827 , y15828 , y15829 , y15830 , y15831 , y15832 , y15833 , y15834 , y15835 , y15836 , y15837 , y15838 , y15839 , y15840 , y15841 , y15842 , y15843 , y15844 , y15845 , y15846 , y15847 , y15848 , y15849 , y15850 , y15851 , y15852 , y15853 , y15854 , y15855 , y15856 , y15857 , y15858 , y15859 , y15860 , y15861 , y15862 , y15863 , y15864 , y15865 , y15866 , y15867 , y15868 , y15869 , y15870 , y15871 , y15872 , y15873 , y15874 , y15875 , y15876 , y15877 , y15878 , y15879 , y15880 , y15881 , y15882 , y15883 , y15884 , y15885 , y15886 , y15887 , y15888 , y15889 , y15890 , y15891 , y15892 , y15893 , y15894 , y15895 , y15896 , y15897 , y15898 , y15899 , y15900 , y15901 , y15902 , y15903 , y15904 , y15905 , y15906 , y15907 , y15908 , y15909 , y15910 , y15911 , y15912 , y15913 , y15914 , y15915 , y15916 , y15917 , y15918 , y15919 , y15920 , y15921 , y15922 , y15923 , y15924 , y15925 , y15926 , y15927 , y15928 , y15929 , y15930 , y15931 , y15932 , y15933 , y15934 , y15935 , y15936 , y15937 , y15938 , y15939 , y15940 , y15941 , y15942 , y15943 , y15944 , y15945 , y15946 , y15947 , y15948 , y15949 , y15950 , y15951 , y15952 , y15953 , y15954 , y15955 , y15956 , y15957 , y15958 , y15959 , y15960 , y15961 , y15962 , y15963 , y15964 , y15965 , y15966 , y15967 , y15968 , y15969 , y15970 , y15971 , y15972 , y15973 , y15974 , y15975 , y15976 , y15977 , y15978 , y15979 , y15980 , y15981 , y15982 , y15983 , y15984 , y15985 , y15986 , y15987 , y15988 , y15989 , y15990 , y15991 , y15992 , y15993 , y15994 , y15995 , y15996 , y15997 , y15998 , y15999 , y16000 , y16001 , y16002 , y16003 , y16004 , y16005 , y16006 , y16007 , y16008 , y16009 , y16010 , y16011 , y16012 , y16013 , y16014 , y16015 , y16016 , y16017 , y16018 , y16019 , y16020 , y16021 , y16022 , y16023 , y16024 , y16025 , y16026 , y16027 , y16028 , y16029 , y16030 , y16031 , y16032 , y16033 , y16034 , y16035 , y16036 , y16037 , y16038 , y16039 , y16040 , y16041 , y16042 , y16043 , y16044 , y16045 , y16046 , y16047 , y16048 , y16049 , y16050 , y16051 , y16052 , y16053 , y16054 , y16055 , y16056 , y16057 , y16058 , y16059 , y16060 , y16061 , y16062 , y16063 , y16064 , y16065 , y16066 , y16067 , y16068 , y16069 , y16070 , y16071 , y16072 , y16073 , y16074 , y16075 , y16076 , y16077 , y16078 , y16079 , y16080 , y16081 , y16082 , y16083 , y16084 , y16085 , y16086 , y16087 , y16088 , y16089 , y16090 , y16091 , y16092 , y16093 , y16094 , y16095 , y16096 , y16097 , y16098 , y16099 , y16100 , y16101 , y16102 , y16103 , y16104 , y16105 , y16106 , y16107 , y16108 , y16109 , y16110 , y16111 , y16112 , y16113 , y16114 , y16115 , y16116 , y16117 , y16118 , y16119 , y16120 , y16121 , y16122 , y16123 , y16124 , y16125 , y16126 , y16127 , y16128 , y16129 , y16130 , y16131 , y16132 , y16133 , y16134 , y16135 , y16136 , y16137 , y16138 , y16139 , y16140 , y16141 , y16142 , y16143 , y16144 , y16145 , y16146 , y16147 , y16148 , y16149 , y16150 , y16151 , y16152 , y16153 , y16154 , y16155 , y16156 , y16157 , y16158 , y16159 , y16160 , y16161 , y16162 , y16163 , y16164 , y16165 , y16166 , y16167 , y16168 , y16169 , y16170 , y16171 , y16172 , y16173 , y16174 , y16175 , y16176 , y16177 , y16178 , y16179 , y16180 , y16181 , y16182 , y16183 , y16184 , y16185 , y16186 , y16187 , y16188 , y16189 , y16190 , y16191 , y16192 , y16193 , y16194 , y16195 , y16196 , y16197 , y16198 , y16199 , y16200 , y16201 , y16202 , y16203 , y16204 , y16205 , y16206 , y16207 , y16208 , y16209 , y16210 , y16211 , y16212 , y16213 , y16214 , y16215 , y16216 , y16217 , y16218 , y16219 , y16220 , y16221 , y16222 , y16223 , y16224 , y16225 , y16226 , y16227 , y16228 , y16229 , y16230 , y16231 , y16232 , y16233 , y16234 , y16235 , y16236 , y16237 , y16238 , y16239 , y16240 , y16241 , y16242 , y16243 , y16244 , y16245 , y16246 , y16247 , y16248 , y16249 , y16250 , y16251 , y16252 , y16253 , y16254 , y16255 , y16256 , y16257 , y16258 , y16259 , y16260 , y16261 , y16262 , y16263 , y16264 , y16265 , y16266 , y16267 , y16268 , y16269 , y16270 , y16271 , y16272 , y16273 , y16274 , y16275 , y16276 , y16277 , y16278 , y16279 , y16280 , y16281 , y16282 , y16283 , y16284 , y16285 , y16286 , y16287 , y16288 , y16289 , y16290 , y16291 , y16292 , y16293 , y16294 , y16295 , y16296 , y16297 , y16298 , y16299 , y16300 , y16301 , y16302 , y16303 , y16304 , y16305 , y16306 , y16307 , y16308 , y16309 , y16310 , y16311 , y16312 , y16313 , y16314 , y16315 , y16316 , y16317 , y16318 , y16319 , y16320 , y16321 , y16322 , y16323 , y16324 , y16325 , y16326 , y16327 , y16328 , y16329 , y16330 , y16331 , y16332 , y16333 , y16334 , y16335 , y16336 , y16337 , y16338 , y16339 , y16340 , y16341 , y16342 , y16343 , y16344 , y16345 , y16346 , y16347 , y16348 , y16349 , y16350 , y16351 , y16352 , y16353 , y16354 , y16355 , y16356 , y16357 , y16358 , y16359 , y16360 , y16361 , y16362 , y16363 , y16364 , y16365 , y16366 , y16367 , y16368 , y16369 , y16370 , y16371 , y16372 , y16373 , y16374 , y16375 , y16376 , y16377 , y16378 , y16379 , y16380 , y16381 , y16382 , y16383 , y16384 , y16385 , y16386 , y16387 , y16388 , y16389 , y16390 , y16391 , y16392 , y16393 , y16394 , y16395 , y16396 , y16397 , y16398 , y16399 , y16400 , y16401 , y16402 , y16403 , y16404 , y16405 , y16406 , y16407 , y16408 , y16409 , y16410 , y16411 , y16412 , y16413 , y16414 , y16415 , y16416 , y16417 , y16418 , y16419 , y16420 , y16421 , y16422 , y16423 , y16424 , y16425 , y16426 , y16427 , y16428 , y16429 , y16430 , y16431 , y16432 , y16433 , y16434 , y16435 , y16436 , y16437 , y16438 , y16439 , y16440 , y16441 , y16442 , y16443 , y16444 , y16445 , y16446 , y16447 , y16448 , y16449 , y16450 , y16451 , y16452 , y16453 , y16454 , y16455 , y16456 , y16457 , y16458 , y16459 , y16460 , y16461 , y16462 , y16463 , y16464 , y16465 , y16466 , y16467 , y16468 , y16469 , y16470 , y16471 , y16472 , y16473 , y16474 , y16475 , y16476 , y16477 , y16478 , y16479 , y16480 , y16481 , y16482 , y16483 , y16484 , y16485 , y16486 , y16487 , y16488 , y16489 , y16490 , y16491 , y16492 , y16493 , y16494 , y16495 , y16496 , y16497 , y16498 , y16499 , y16500 , y16501 , y16502 , y16503 , y16504 , y16505 , y16506 , y16507 , y16508 , y16509 , y16510 , y16511 , y16512 , y16513 , y16514 , y16515 , y16516 , y16517 , y16518 , y16519 , y16520 , y16521 , y16522 , y16523 , y16524 , y16525 , y16526 , y16527 , y16528 , y16529 , y16530 , y16531 , y16532 , y16533 , y16534 , y16535 , y16536 , y16537 , y16538 , y16539 , y16540 , y16541 , y16542 , y16543 , y16544 , y16545 , y16546 , y16547 , y16548 , y16549 , y16550 , y16551 , y16552 , y16553 , y16554 , y16555 , y16556 , y16557 , y16558 , y16559 , y16560 , y16561 , y16562 , y16563 , y16564 , y16565 , y16566 , y16567 , y16568 , y16569 , y16570 , y16571 , y16572 , y16573 , y16574 , y16575 , y16576 , y16577 , y16578 , y16579 , y16580 , y16581 , y16582 , y16583 , y16584 , y16585 , y16586 , y16587 , y16588 , y16589 , y16590 , y16591 , y16592 , y16593 , y16594 , y16595 , y16596 , y16597 , y16598 , y16599 , y16600 , y16601 , y16602 , y16603 , y16604 , y16605 , y16606 , y16607 , y16608 , y16609 , y16610 , y16611 , y16612 , y16613 , y16614 , y16615 , y16616 , y16617 , y16618 , y16619 , y16620 , y16621 , y16622 , y16623 , y16624 , y16625 , y16626 , y16627 , y16628 , y16629 , y16630 , y16631 , y16632 , y16633 , y16634 , y16635 , y16636 , y16637 , y16638 , y16639 , y16640 , y16641 , y16642 , y16643 , y16644 , y16645 , y16646 , y16647 , y16648 , y16649 , y16650 , y16651 , y16652 , y16653 , y16654 , y16655 , y16656 , y16657 , y16658 , y16659 , y16660 , y16661 , y16662 , y16663 , y16664 , y16665 , y16666 , y16667 , y16668 , y16669 , y16670 , y16671 , y16672 , y16673 , y16674 , y16675 , y16676 , y16677 , y16678 , y16679 , y16680 , y16681 , y16682 , y16683 , y16684 , y16685 , y16686 , y16687 , y16688 , y16689 , y16690 , y16691 , y16692 , y16693 , y16694 , y16695 , y16696 , y16697 , y16698 , y16699 , y16700 , y16701 , y16702 , y16703 , y16704 , y16705 , y16706 , y16707 , y16708 , y16709 , y16710 , y16711 , y16712 , y16713 , y16714 , y16715 , y16716 , y16717 , y16718 , y16719 , y16720 , y16721 , y16722 , y16723 , y16724 , y16725 , y16726 , y16727 , y16728 , y16729 , y16730 , y16731 , y16732 , y16733 , y16734 , y16735 , y16736 , y16737 , y16738 , y16739 , y16740 , y16741 , y16742 , y16743 , y16744 , y16745 , y16746 , y16747 , y16748 , y16749 , y16750 , y16751 , y16752 , y16753 , y16754 , y16755 , y16756 , y16757 , y16758 , y16759 , y16760 , y16761 , y16762 , y16763 , y16764 , y16765 , y16766 , y16767 , y16768 , y16769 , y16770 , y16771 , y16772 , y16773 , y16774 , y16775 , y16776 , y16777 , y16778 , y16779 , y16780 , y16781 , y16782 , y16783 , y16784 , y16785 , y16786 , y16787 , y16788 , y16789 , y16790 , y16791 , y16792 , y16793 , y16794 , y16795 , y16796 , y16797 , y16798 , y16799 , y16800 , y16801 , y16802 , y16803 , y16804 , y16805 , y16806 , y16807 , y16808 , y16809 , y16810 , y16811 , y16812 , y16813 , y16814 , y16815 , y16816 , y16817 , y16818 , y16819 , y16820 , y16821 , y16822 , y16823 , y16824 , y16825 , y16826 , y16827 , y16828 , y16829 , y16830 , y16831 , y16832 , y16833 , y16834 , y16835 , y16836 , y16837 , y16838 , y16839 , y16840 , y16841 , y16842 , y16843 , y16844 , y16845 , y16846 , y16847 , y16848 , y16849 , y16850 , y16851 , y16852 , y16853 , y16854 , y16855 , y16856 , y16857 , y16858 , y16859 , y16860 , y16861 , y16862 , y16863 , y16864 , y16865 , y16866 , y16867 , y16868 , y16869 , y16870 , y16871 , y16872 , y16873 , y16874 , y16875 , y16876 , y16877 , y16878 , y16879 , y16880 , y16881 , y16882 , y16883 , y16884 , y16885 , y16886 , y16887 , y16888 , y16889 , y16890 , y16891 , y16892 , y16893 , y16894 , y16895 , y16896 , y16897 , y16898 , y16899 , y16900 , y16901 , y16902 , y16903 , y16904 , y16905 , y16906 , y16907 , y16908 , y16909 , y16910 , y16911 , y16912 , y16913 , y16914 , y16915 , y16916 , y16917 , y16918 , y16919 , y16920 , y16921 , y16922 , y16923 , y16924 , y16925 , y16926 , y16927 , y16928 , y16929 , y16930 , y16931 , y16932 , y16933 , y16934 , y16935 , y16936 , y16937 , y16938 , y16939 , y16940 , y16941 , y16942 , y16943 , y16944 , y16945 , y16946 , y16947 , y16948 , y16949 , y16950 , y16951 , y16952 , y16953 , y16954 , y16955 , y16956 , y16957 , y16958 , y16959 , y16960 , y16961 , y16962 , y16963 , y16964 , y16965 , y16966 , y16967 , y16968 , y16969 , y16970 , y16971 , y16972 , y16973 , y16974 , y16975 , y16976 , y16977 , y16978 , y16979 , y16980 , y16981 , y16982 , y16983 , y16984 , y16985 , y16986 , y16987 , y16988 , y16989 , y16990 , y16991 , y16992 , y16993 , y16994 , y16995 , y16996 , y16997 , y16998 , y16999 , y17000 , y17001 , y17002 , y17003 , y17004 , y17005 , y17006 , y17007 , y17008 , y17009 , y17010 , y17011 , y17012 , y17013 , y17014 , y17015 , y17016 , y17017 , y17018 , y17019 , y17020 , y17021 , y17022 , y17023 , y17024 , y17025 , y17026 , y17027 , y17028 , y17029 , y17030 , y17031 , y17032 , y17033 , y17034 , y17035 , y17036 , y17037 , y17038 , y17039 , y17040 , y17041 , y17042 , y17043 , y17044 , y17045 , y17046 , y17047 , y17048 , y17049 , y17050 , y17051 , y17052 , y17053 , y17054 , y17055 , y17056 , y17057 , y17058 , y17059 , y17060 , y17061 , y17062 , y17063 , y17064 , y17065 , y17066 , y17067 , y17068 , y17069 , y17070 , y17071 , y17072 , y17073 , y17074 , y17075 , y17076 , y17077 , y17078 , y17079 , y17080 , y17081 , y17082 , y17083 , y17084 , y17085 , y17086 , y17087 , y17088 , y17089 , y17090 , y17091 , y17092 , y17093 , y17094 , y17095 , y17096 , y17097 , y17098 , y17099 , y17100 , y17101 , y17102 , y17103 , y17104 , y17105 , y17106 , y17107 , y17108 , y17109 , y17110 , y17111 , y17112 , y17113 , y17114 , y17115 , y17116 , y17117 , y17118 , y17119 , y17120 , y17121 , y17122 , y17123 , y17124 , y17125 , y17126 , y17127 , y17128 , y17129 , y17130 , y17131 , y17132 , y17133 , y17134 , y17135 , y17136 , y17137 , y17138 , y17139 , y17140 , y17141 , y17142 , y17143 , y17144 , y17145 , y17146 , y17147 , y17148 , y17149 , y17150 , y17151 , y17152 , y17153 , y17154 , y17155 , y17156 , y17157 , y17158 , y17159 , y17160 , y17161 , y17162 , y17163 , y17164 , y17165 , y17166 , y17167 , y17168 , y17169 , y17170 , y17171 , y17172 , y17173 , y17174 , y17175 , y17176 , y17177 , y17178 , y17179 , y17180 , y17181 , y17182 , y17183 , y17184 , y17185 , y17186 , y17187 , y17188 , y17189 , y17190 , y17191 , y17192 , y17193 , y17194 , y17195 , y17196 , y17197 , y17198 , y17199 , y17200 , y17201 , y17202 , y17203 , y17204 , y17205 , y17206 , y17207 , y17208 , y17209 , y17210 , y17211 , y17212 , y17213 , y17214 , y17215 , y17216 , y17217 , y17218 , y17219 , y17220 , y17221 , y17222 , y17223 , y17224 , y17225 , y17226 , y17227 , y17228 , y17229 , y17230 , y17231 , y17232 , y17233 , y17234 , y17235 , y17236 , y17237 , y17238 , y17239 , y17240 , y17241 , y17242 , y17243 , y17244 , y17245 , y17246 , y17247 , y17248 , y17249 , y17250 , y17251 , y17252 , y17253 , y17254 , y17255 , y17256 , y17257 , y17258 , y17259 , y17260 , y17261 , y17262 , y17263 , y17264 , y17265 , y17266 , y17267 , y17268 , y17269 , y17270 , y17271 , y17272 , y17273 , y17274 , y17275 , y17276 , y17277 , y17278 , y17279 , y17280 , y17281 , y17282 , y17283 , y17284 , y17285 , y17286 , y17287 , y17288 , y17289 , y17290 , y17291 , y17292 , y17293 , y17294 , y17295 , y17296 , y17297 , y17298 , y17299 , y17300 , y17301 , y17302 , y17303 , y17304 , y17305 , y17306 , y17307 , y17308 , y17309 , y17310 , y17311 , y17312 , y17313 , y17314 , y17315 , y17316 , y17317 , y17318 , y17319 , y17320 , y17321 , y17322 , y17323 , y17324 , y17325 , y17326 , y17327 , y17328 , y17329 , y17330 , y17331 , y17332 , y17333 , y17334 , y17335 , y17336 , y17337 , y17338 , y17339 , y17340 , y17341 , y17342 , y17343 , y17344 , y17345 , y17346 , y17347 , y17348 , y17349 , y17350 , y17351 , y17352 , y17353 , y17354 , y17355 , y17356 , y17357 , y17358 , y17359 , y17360 , y17361 , y17362 , y17363 , y17364 , y17365 , y17366 , y17367 , y17368 , y17369 , y17370 , y17371 , y17372 , y17373 , y17374 , y17375 , y17376 , y17377 , y17378 , y17379 , y17380 , y17381 , y17382 , y17383 , y17384 , y17385 , y17386 , y17387 , y17388 , y17389 , y17390 , y17391 , y17392 , y17393 , y17394 , y17395 , y17396 , y17397 , y17398 , y17399 , y17400 , y17401 , y17402 , y17403 , y17404 , y17405 , y17406 , y17407 , y17408 , y17409 , y17410 , y17411 , y17412 , y17413 , y17414 , y17415 , y17416 , y17417 , y17418 , y17419 , y17420 , y17421 , y17422 , y17423 , y17424 , y17425 , y17426 , y17427 , y17428 , y17429 , y17430 , y17431 , y17432 , y17433 , y17434 , y17435 , y17436 , y17437 , y17438 , y17439 , y17440 , y17441 , y17442 , y17443 , y17444 , y17445 , y17446 , y17447 , y17448 , y17449 , y17450 , y17451 , y17452 , y17453 , y17454 , y17455 , y17456 , y17457 , y17458 , y17459 , y17460 , y17461 , y17462 , y17463 , y17464 , y17465 , y17466 , y17467 , y17468 , y17469 , y17470 , y17471 , y17472 , y17473 , y17474 , y17475 , y17476 , y17477 , y17478 , y17479 , y17480 , y17481 , y17482 , y17483 , y17484 , y17485 , y17486 , y17487 , y17488 , y17489 , y17490 , y17491 , y17492 , y17493 , y17494 , y17495 , y17496 , y17497 , y17498 , y17499 , y17500 , y17501 , y17502 , y17503 , y17504 , y17505 , y17506 , y17507 , y17508 , y17509 , y17510 , y17511 , y17512 , y17513 , y17514 , y17515 , y17516 , y17517 , y17518 , y17519 , y17520 , y17521 , y17522 , y17523 , y17524 , y17525 , y17526 , y17527 , y17528 , y17529 , y17530 , y17531 , y17532 , y17533 , y17534 , y17535 , y17536 , y17537 , y17538 , y17539 , y17540 , y17541 , y17542 , y17543 , y17544 , y17545 , y17546 , y17547 , y17548 , y17549 , y17550 , y17551 , y17552 , y17553 , y17554 , y17555 , y17556 , y17557 , y17558 , y17559 , y17560 , y17561 , y17562 , y17563 , y17564 , y17565 , y17566 , y17567 , y17568 , y17569 , y17570 , y17571 , y17572 , y17573 , y17574 , y17575 , y17576 , y17577 , y17578 , y17579 , y17580 , y17581 , y17582 , y17583 , y17584 , y17585 , y17586 , y17587 , y17588 , y17589 , y17590 , y17591 , y17592 , y17593 , y17594 , y17595 , y17596 , y17597 , y17598 , y17599 , y17600 , y17601 , y17602 , y17603 , y17604 , y17605 , y17606 , y17607 , y17608 , y17609 , y17610 , y17611 , y17612 , y17613 , y17614 , y17615 , y17616 , y17617 , y17618 , y17619 , y17620 , y17621 , y17622 , y17623 , y17624 , y17625 , y17626 , y17627 , y17628 , y17629 , y17630 , y17631 , y17632 , y17633 , y17634 , y17635 , y17636 , y17637 , y17638 , y17639 , y17640 , y17641 , y17642 , y17643 , y17644 , y17645 , y17646 , y17647 , y17648 , y17649 , y17650 , y17651 , y17652 , y17653 , y17654 , y17655 , y17656 , y17657 , y17658 , y17659 , y17660 , y17661 , y17662 , y17663 , y17664 , y17665 , y17666 , y17667 , y17668 , y17669 , y17670 , y17671 , y17672 , y17673 , y17674 , y17675 , y17676 , y17677 , y17678 , y17679 , y17680 , y17681 , y17682 , y17683 , y17684 , y17685 , y17686 , y17687 , y17688 , y17689 , y17690 , y17691 , y17692 , y17693 , y17694 , y17695 , y17696 , y17697 , y17698 , y17699 , y17700 , y17701 , y17702 , y17703 , y17704 , y17705 , y17706 , y17707 , y17708 , y17709 , y17710 , y17711 , y17712 , y17713 , y17714 , y17715 , y17716 , y17717 , y17718 , y17719 , y17720 , y17721 , y17722 , y17723 , y17724 , y17725 , y17726 , y17727 , y17728 , y17729 , y17730 , y17731 , y17732 , y17733 , y17734 , y17735 , y17736 , y17737 , y17738 , y17739 , y17740 , y17741 , y17742 , y17743 , y17744 , y17745 , y17746 , y17747 , y17748 , y17749 , y17750 , y17751 , y17752 , y17753 , y17754 , y17755 , y17756 , y17757 , y17758 , y17759 , y17760 , y17761 , y17762 , y17763 , y17764 , y17765 , y17766 , y17767 , y17768 , y17769 , y17770 , y17771 , y17772 , y17773 , y17774 , y17775 , y17776 , y17777 , y17778 , y17779 , y17780 , y17781 , y17782 , y17783 , y17784 , y17785 , y17786 , y17787 , y17788 , y17789 , y17790 , y17791 , y17792 , y17793 , y17794 , y17795 , y17796 , y17797 , y17798 , y17799 , y17800 , y17801 , y17802 , y17803 , y17804 , y17805 , y17806 , y17807 , y17808 , y17809 , y17810 , y17811 , y17812 , y17813 , y17814 , y17815 , y17816 , y17817 , y17818 , y17819 , y17820 , y17821 , y17822 , y17823 , y17824 , y17825 , y17826 , y17827 , y17828 , y17829 , y17830 , y17831 , y17832 , y17833 , y17834 , y17835 , y17836 , y17837 , y17838 , y17839 , y17840 , y17841 , y17842 , y17843 , y17844 , y17845 , y17846 , y17847 , y17848 , y17849 , y17850 , y17851 , y17852 , y17853 , y17854 , y17855 , y17856 , y17857 , y17858 , y17859 , y17860 , y17861 , y17862 , y17863 , y17864 , y17865 , y17866 , y17867 , y17868 , y17869 , y17870 , y17871 , y17872 , y17873 , y17874 , y17875 , y17876 , y17877 , y17878 , y17879 , y17880 , y17881 , y17882 , y17883 , y17884 , y17885 , y17886 , y17887 , y17888 , y17889 , y17890 , y17891 , y17892 , y17893 , y17894 , y17895 , y17896 , y17897 , y17898 , y17899 , y17900 , y17901 , y17902 , y17903 , y17904 , y17905 , y17906 , y17907 , y17908 , y17909 , y17910 , y17911 , y17912 , y17913 , y17914 , y17915 , y17916 , y17917 , y17918 , y17919 , y17920 , y17921 , y17922 , y17923 , y17924 , y17925 , y17926 , y17927 , y17928 , y17929 , y17930 , y17931 , y17932 , y17933 , y17934 , y17935 , y17936 , y17937 , y17938 , y17939 , y17940 , y17941 , y17942 , y17943 , y17944 , y17945 , y17946 , y17947 , y17948 , y17949 , y17950 , y17951 , y17952 , y17953 , y17954 , y17955 , y17956 , y17957 , y17958 , y17959 , y17960 , y17961 , y17962 , y17963 , y17964 , y17965 , y17966 , y17967 , y17968 , y17969 , y17970 , y17971 , y17972 , y17973 , y17974 , y17975 , y17976 , y17977 , y17978 , y17979 , y17980 , y17981 , y17982 , y17983 , y17984 , y17985 , y17986 , y17987 , y17988 , y17989 , y17990 , y17991 , y17992 , y17993 , y17994 , y17995 , y17996 , y17997 , y17998 , y17999 , y18000 , y18001 , y18002 , y18003 , y18004 , y18005 , y18006 , y18007 , y18008 , y18009 , y18010 , y18011 , y18012 , y18013 , y18014 , y18015 , y18016 , y18017 , y18018 , y18019 , y18020 , y18021 , y18022 , y18023 , y18024 , y18025 , y18026 , y18027 , y18028 , y18029 , y18030 , y18031 , y18032 , y18033 , y18034 , y18035 , y18036 , y18037 , y18038 , y18039 , y18040 , y18041 , y18042 , y18043 , y18044 , y18045 , y18046 , y18047 , y18048 , y18049 , y18050 , y18051 , y18052 , y18053 , y18054 , y18055 , y18056 , y18057 , y18058 , y18059 , y18060 , y18061 , y18062 , y18063 , y18064 , y18065 , y18066 , y18067 , y18068 , y18069 , y18070 , y18071 , y18072 , y18073 , y18074 , y18075 , y18076 , y18077 , y18078 , y18079 , y18080 , y18081 , y18082 , y18083 , y18084 , y18085 , y18086 , y18087 , y18088 , y18089 , y18090 , y18091 , y18092 , y18093 , y18094 , y18095 , y18096 , y18097 , y18098 , y18099 , y18100 , y18101 , y18102 , y18103 , y18104 , y18105 , y18106 , y18107 , y18108 , y18109 , y18110 , y18111 , y18112 , y18113 , y18114 , y18115 , y18116 , y18117 , y18118 , y18119 , y18120 , y18121 , y18122 , y18123 , y18124 , y18125 , y18126 , y18127 , y18128 , y18129 , y18130 , y18131 , y18132 , y18133 , y18134 , y18135 , y18136 , y18137 , y18138 , y18139 , y18140 , y18141 , y18142 , y18143 , y18144 , y18145 , y18146 , y18147 , y18148 , y18149 , y18150 , y18151 , y18152 , y18153 , y18154 , y18155 , y18156 , y18157 , y18158 , y18159 , y18160 , y18161 , y18162 , y18163 , y18164 , y18165 , y18166 , y18167 , y18168 , y18169 , y18170 , y18171 , y18172 , y18173 , y18174 , y18175 , y18176 , y18177 , y18178 , y18179 , y18180 , y18181 , y18182 , y18183 , y18184 , y18185 , y18186 , y18187 , y18188 , y18189 , y18190 , y18191 , y18192 , y18193 , y18194 , y18195 , y18196 , y18197 , y18198 , y18199 , y18200 , y18201 , y18202 , y18203 , y18204 , y18205 , y18206 , y18207 , y18208 , y18209 , y18210 , y18211 , y18212 , y18213 , y18214 , y18215 , y18216 , y18217 , y18218 , y18219 , y18220 , y18221 , y18222 , y18223 , y18224 , y18225 , y18226 , y18227 , y18228 , y18229 , y18230 , y18231 , y18232 , y18233 , y18234 , y18235 , y18236 , y18237 , y18238 , y18239 , y18240 , y18241 , y18242 , y18243 , y18244 , y18245 , y18246 , y18247 , y18248 , y18249 , y18250 , y18251 , y18252 , y18253 , y18254 , y18255 , y18256 , y18257 , y18258 , y18259 , y18260 , y18261 , y18262 , y18263 , y18264 , y18265 , y18266 , y18267 , y18268 , y18269 , y18270 , y18271 , y18272 , y18273 , y18274 , y18275 , y18276 , y18277 , y18278 , y18279 , y18280 , y18281 , y18282 , y18283 , y18284 , y18285 , y18286 , y18287 , y18288 , y18289 , y18290 , y18291 , y18292 , y18293 , y18294 , y18295 , y18296 , y18297 , y18298 , y18299 , y18300 , y18301 , y18302 , y18303 , y18304 , y18305 , y18306 , y18307 , y18308 , y18309 , y18310 , y18311 , y18312 , y18313 , y18314 , y18315 , y18316 , y18317 , y18318 , y18319 , y18320 , y18321 , y18322 , y18323 , y18324 , y18325 , y18326 , y18327 , y18328 , y18329 , y18330 , y18331 , y18332 , y18333 , y18334 , y18335 , y18336 , y18337 , y18338 , y18339 , y18340 , y18341 , y18342 , y18343 , y18344 , y18345 , y18346 , y18347 , y18348 , y18349 , y18350 , y18351 , y18352 , y18353 , y18354 , y18355 , y18356 , y18357 , y18358 , y18359 , y18360 , y18361 , y18362 , y18363 , y18364 , y18365 , y18366 , y18367 , y18368 , y18369 , y18370 , y18371 , y18372 , y18373 , y18374 , y18375 , y18376 , y18377 , y18378 , y18379 , y18380 , y18381 , y18382 , y18383 , y18384 , y18385 , y18386 , y18387 , y18388 , y18389 , y18390 , y18391 , y18392 , y18393 , y18394 , y18395 , y18396 , y18397 , y18398 , y18399 , y18400 , y18401 , y18402 , y18403 , y18404 , y18405 , y18406 , y18407 , y18408 , y18409 , y18410 , y18411 , y18412 , y18413 , y18414 , y18415 , y18416 , y18417 , y18418 , y18419 , y18420 , y18421 , y18422 , y18423 , y18424 , y18425 , y18426 , y18427 , y18428 , y18429 , y18430 , y18431 , y18432 , y18433 , y18434 , y18435 , y18436 , y18437 , y18438 , y18439 , y18440 , y18441 , y18442 , y18443 , y18444 , y18445 , y18446 , y18447 , y18448 , y18449 , y18450 , y18451 , y18452 , y18453 , y18454 , y18455 , y18456 , y18457 , y18458 , y18459 , y18460 , y18461 , y18462 , y18463 , y18464 , y18465 , y18466 , y18467 , y18468 , y18469 , y18470 , y18471 , y18472 , y18473 , y18474 , y18475 , y18476 , y18477 , y18478 , y18479 , y18480 , y18481 , y18482 , y18483 , y18484 , y18485 , y18486 , y18487 , y18488 , y18489 , y18490 , y18491 , y18492 , y18493 , y18494 , y18495 , y18496 , y18497 , y18498 , y18499 , y18500 , y18501 , y18502 , y18503 , y18504 , y18505 , y18506 , y18507 , y18508 , y18509 , y18510 , y18511 , y18512 , y18513 , y18514 , y18515 , y18516 , y18517 , y18518 , y18519 , y18520 , y18521 , y18522 , y18523 , y18524 , y18525 , y18526 , y18527 , y18528 , y18529 , y18530 , y18531 , y18532 , y18533 , y18534 , y18535 , y18536 , y18537 , y18538 , y18539 , y18540 , y18541 , y18542 , y18543 , y18544 , y18545 , y18546 , y18547 , y18548 , y18549 , y18550 , y18551 , y18552 , y18553 , y18554 , y18555 , y18556 , y18557 , y18558 , y18559 , y18560 , y18561 , y18562 , y18563 , y18564 , y18565 , y18566 , y18567 , y18568 , y18569 , y18570 , y18571 , y18572 , y18573 , y18574 , y18575 , y18576 , y18577 , y18578 , y18579 , y18580 , y18581 , y18582 , y18583 , y18584 , y18585 , y18586 , y18587 , y18588 , y18589 , y18590 , y18591 , y18592 , y18593 , y18594 , y18595 , y18596 , y18597 , y18598 , y18599 , y18600 , y18601 , y18602 , y18603 , y18604 , y18605 , y18606 , y18607 , y18608 , y18609 , y18610 , y18611 , y18612 , y18613 , y18614 , y18615 , y18616 , y18617 , y18618 , y18619 , y18620 , y18621 , y18622 , y18623 , y18624 , y18625 , y18626 , y18627 , y18628 , y18629 , y18630 , y18631 , y18632 , y18633 , y18634 , y18635 , y18636 , y18637 , y18638 , y18639 , y18640 , y18641 , y18642 , y18643 , y18644 , y18645 , y18646 , y18647 , y18648 , y18649 , y18650 , y18651 , y18652 , y18653 , y18654 , y18655 , y18656 , y18657 , y18658 , y18659 , y18660 , y18661 , y18662 , y18663 , y18664 , y18665 , y18666 , y18667 , y18668 , y18669 , y18670 , y18671 , y18672 , y18673 , y18674 , y18675 , y18676 , y18677 , y18678 , y18679 , y18680 , y18681 , y18682 , y18683 , y18684 , y18685 , y18686 , y18687 , y18688 , y18689 , y18690 , y18691 , y18692 , y18693 , y18694 , y18695 , y18696 , y18697 , y18698 , y18699 , y18700 , y18701 , y18702 , y18703 , y18704 , y18705 , y18706 , y18707 , y18708 , y18709 , y18710 , y18711 , y18712 , y18713 , y18714 , y18715 , y18716 , y18717 , y18718 , y18719 , y18720 , y18721 , y18722 , y18723 , y18724 , y18725 , y18726 , y18727 , y18728 , y18729 , y18730 , y18731 , y18732 , y18733 , y18734 , y18735 , y18736 , y18737 , y18738 , y18739 , y18740 , y18741 , y18742 , y18743 , y18744 , y18745 , y18746 , y18747 , y18748 , y18749 , y18750 , y18751 , y18752 , y18753 , y18754 , y18755 , y18756 , y18757 , y18758 , y18759 , y18760 , y18761 , y18762 , y18763 , y18764 , y18765 , y18766 , y18767 , y18768 , y18769 , y18770 , y18771 , y18772 , y18773 , y18774 , y18775 , y18776 , y18777 , y18778 , y18779 , y18780 , y18781 , y18782 , y18783 , y18784 , y18785 , y18786 , y18787 , y18788 , y18789 , y18790 , y18791 , y18792 , y18793 , y18794 , y18795 , y18796 , y18797 , y18798 , y18799 , y18800 , y18801 , y18802 , y18803 , y18804 , y18805 , y18806 , y18807 , y18808 , y18809 , y18810 , y18811 , y18812 , y18813 , y18814 , y18815 , y18816 , y18817 , y18818 , y18819 , y18820 , y18821 , y18822 , y18823 , y18824 , y18825 , y18826 , y18827 , y18828 , y18829 , y18830 , y18831 , y18832 , y18833 , y18834 , y18835 , y18836 , y18837 , y18838 , y18839 , y18840 , y18841 , y18842 , y18843 , y18844 , y18845 , y18846 , y18847 , y18848 , y18849 , y18850 , y18851 , y18852 , y18853 , y18854 , y18855 , y18856 , y18857 , y18858 , y18859 , y18860 , y18861 , y18862 , y18863 , y18864 , y18865 , y18866 , y18867 , y18868 , y18869 , y18870 , y18871 , y18872 , y18873 , y18874 , y18875 , y18876 , y18877 , y18878 , y18879 , y18880 , y18881 , y18882 , y18883 , y18884 , y18885 , y18886 , y18887 , y18888 , y18889 , y18890 , y18891 , y18892 , y18893 , y18894 , y18895 , y18896 , y18897 , y18898 , y18899 , y18900 , y18901 , y18902 , y18903 , y18904 , y18905 , y18906 , y18907 , y18908 , y18909 , y18910 , y18911 , y18912 , y18913 , y18914 , y18915 , y18916 , y18917 , y18918 , y18919 , y18920 , y18921 , y18922 , y18923 , y18924 , y18925 , y18926 , y18927 , y18928 , y18929 , y18930 , y18931 , y18932 , y18933 , y18934 , y18935 , y18936 , y18937 , y18938 , y18939 , y18940 , y18941 , y18942 , y18943 , y18944 , y18945 , y18946 , y18947 , y18948 , y18949 , y18950 , y18951 , y18952 , y18953 , y18954 , y18955 , y18956 , y18957 , y18958 , y18959 , y18960 , y18961 , y18962 , y18963 , y18964 , y18965 , y18966 , y18967 , y18968 , y18969 , y18970 , y18971 , y18972 , y18973 , y18974 , y18975 , y18976 , y18977 , y18978 , y18979 , y18980 , y18981 , y18982 , y18983 , y18984 , y18985 , y18986 , y18987 , y18988 , y18989 , y18990 , y18991 , y18992 , y18993 , y18994 , y18995 , y18996 , y18997 , y18998 , y18999 , y19000 , y19001 , y19002 , y19003 , y19004 , y19005 , y19006 , y19007 , y19008 , y19009 , y19010 , y19011 , y19012 , y19013 , y19014 , y19015 , y19016 , y19017 , y19018 , y19019 , y19020 , y19021 , y19022 , y19023 , y19024 , y19025 , y19026 , y19027 , y19028 , y19029 , y19030 , y19031 , y19032 , y19033 , y19034 , y19035 , y19036 , y19037 , y19038 , y19039 , y19040 , y19041 , y19042 , y19043 , y19044 , y19045 , y19046 , y19047 , y19048 , y19049 , y19050 , y19051 , y19052 , y19053 , y19054 , y19055 , y19056 , y19057 , y19058 , y19059 , y19060 , y19061 , y19062 , y19063 , y19064 , y19065 , y19066 , y19067 , y19068 , y19069 , y19070 , y19071 , y19072 , y19073 , y19074 , y19075 , y19076 , y19077 , y19078 , y19079 , y19080 , y19081 , y19082 , y19083 , y19084 , y19085 , y19086 , y19087 , y19088 , y19089 , y19090 , y19091 , y19092 , y19093 , y19094 , y19095 , y19096 , y19097 , y19098 , y19099 , y19100 , y19101 , y19102 , y19103 , y19104 , y19105 , y19106 , y19107 , y19108 , y19109 , y19110 , y19111 , y19112 , y19113 , y19114 , y19115 , y19116 , y19117 , y19118 , y19119 , y19120 , y19121 , y19122 , y19123 , y19124 , y19125 , y19126 , y19127 , y19128 , y19129 , y19130 , y19131 , y19132 , y19133 , y19134 , y19135 , y19136 , y19137 , y19138 , y19139 , y19140 , y19141 , y19142 , y19143 , y19144 , y19145 , y19146 , y19147 , y19148 , y19149 , y19150 , y19151 , y19152 , y19153 , y19154 , y19155 , y19156 , y19157 , y19158 , y19159 , y19160 , y19161 , y19162 , y19163 , y19164 , y19165 , y19166 , y19167 , y19168 , y19169 , y19170 , y19171 , y19172 , y19173 , y19174 , y19175 , y19176 , y19177 , y19178 , y19179 , y19180 , y19181 , y19182 , y19183 , y19184 , y19185 , y19186 , y19187 , y19188 , y19189 , y19190 , y19191 , y19192 , y19193 , y19194 , y19195 , y19196 , y19197 , y19198 , y19199 , y19200 , y19201 , y19202 , y19203 , y19204 , y19205 , y19206 , y19207 , y19208 , y19209 , y19210 , y19211 , y19212 , y19213 , y19214 , y19215 , y19216 , y19217 , y19218 , y19219 , y19220 , y19221 , y19222 , y19223 , y19224 , y19225 , y19226 , y19227 , y19228 , y19229 , y19230 , y19231 , y19232 , y19233 , y19234 , y19235 , y19236 , y19237 , y19238 , y19239 , y19240 , y19241 , y19242 , y19243 , y19244 , y19245 , y19246 , y19247 , y19248 , y19249 , y19250 , y19251 , y19252 , y19253 , y19254 , y19255 , y19256 , y19257 , y19258 , y19259 , y19260 , y19261 , y19262 , y19263 , y19264 , y19265 , y19266 , y19267 , y19268 , y19269 , y19270 , y19271 , y19272 , y19273 , y19274 , y19275 , y19276 , y19277 , y19278 , y19279 , y19280 , y19281 , y19282 , y19283 , y19284 , y19285 , y19286 , y19287 , y19288 , y19289 , y19290 , y19291 , y19292 , y19293 , y19294 , y19295 , y19296 , y19297 , y19298 , y19299 , y19300 , y19301 , y19302 , y19303 , y19304 , y19305 , y19306 , y19307 , y19308 , y19309 , y19310 , y19311 , y19312 , y19313 , y19314 , y19315 , y19316 , y19317 , y19318 , y19319 , y19320 , y19321 , y19322 , y19323 , y19324 , y19325 , y19326 , y19327 , y19328 , y19329 , y19330 , y19331 , y19332 , y19333 , y19334 , y19335 , y19336 , y19337 , y19338 , y19339 , y19340 , y19341 , y19342 , y19343 , y19344 , y19345 , y19346 , y19347 , y19348 , y19349 , y19350 , y19351 , y19352 , y19353 , y19354 , y19355 , y19356 , y19357 , y19358 , y19359 , y19360 , y19361 , y19362 , y19363 , y19364 , y19365 , y19366 , y19367 , y19368 , y19369 , y19370 , y19371 , y19372 , y19373 , y19374 , y19375 , y19376 , y19377 , y19378 , y19379 , y19380 , y19381 , y19382 , y19383 , y19384 , y19385 , y19386 , y19387 , y19388 , y19389 , y19390 , y19391 , y19392 , y19393 , y19394 , y19395 , y19396 , y19397 , y19398 , y19399 , y19400 , y19401 , y19402 , y19403 , y19404 , y19405 , y19406 , y19407 , y19408 , y19409 , y19410 , y19411 , y19412 , y19413 , y19414 , y19415 , y19416 , y19417 , y19418 , y19419 , y19420 , y19421 , y19422 , y19423 , y19424 , y19425 , y19426 , y19427 , y19428 , y19429 , y19430 , y19431 , y19432 , y19433 , y19434 , y19435 , y19436 , y19437 , y19438 , y19439 , y19440 , y19441 , y19442 , y19443 , y19444 , y19445 , y19446 , y19447 , y19448 , y19449 , y19450 , y19451 , y19452 , y19453 , y19454 , y19455 , y19456 , y19457 , y19458 , y19459 , y19460 , y19461 , y19462 , y19463 , y19464 , y19465 , y19466 , y19467 , y19468 , y19469 , y19470 , y19471 , y19472 , y19473 , y19474 , y19475 , y19476 , y19477 , y19478 , y19479 , y19480 , y19481 , y19482 , y19483 , y19484 , y19485 , y19486 , y19487 , y19488 , y19489 , y19490 , y19491 , y19492 , y19493 , y19494 , y19495 , y19496 , y19497 , y19498 , y19499 , y19500 , y19501 , y19502 , y19503 , y19504 , y19505 , y19506 , y19507 , y19508 , y19509 , y19510 , y19511 , y19512 , y19513 , y19514 , y19515 , y19516 , y19517 , y19518 , y19519 , y19520 , y19521 , y19522 , y19523 , y19524 , y19525 , y19526 , y19527 , y19528 , y19529 , y19530 , y19531 , y19532 , y19533 , y19534 , y19535 , y19536 , y19537 , y19538 , y19539 , y19540 , y19541 , y19542 , y19543 , y19544 , y19545 , y19546 , y19547 , y19548 , y19549 , y19550 , y19551 , y19552 , y19553 , y19554 , y19555 , y19556 , y19557 , y19558 , y19559 , y19560 , y19561 , y19562 , y19563 , y19564 , y19565 , y19566 , y19567 , y19568 , y19569 , y19570 , y19571 , y19572 , y19573 , y19574 , y19575 , y19576 , y19577 , y19578 , y19579 , y19580 , y19581 , y19582 , y19583 , y19584 , y19585 , y19586 , y19587 , y19588 , y19589 , y19590 , y19591 , y19592 , y19593 , y19594 , y19595 , y19596 , y19597 , y19598 , y19599 , y19600 , y19601 , y19602 , y19603 , y19604 , y19605 , y19606 , y19607 , y19608 , y19609 , y19610 , y19611 , y19612 , y19613 , y19614 , y19615 , y19616 , y19617 , y19618 , y19619 , y19620 , y19621 , y19622 , y19623 , y19624 , y19625 , y19626 , y19627 , y19628 , y19629 , y19630 , y19631 , y19632 , y19633 , y19634 , y19635 , y19636 , y19637 , y19638 , y19639 , y19640 , y19641 , y19642 , y19643 , y19644 , y19645 , y19646 , y19647 , y19648 , y19649 , y19650 , y19651 , y19652 , y19653 , y19654 , y19655 , y19656 , y19657 , y19658 , y19659 , y19660 , y19661 , y19662 , y19663 , y19664 , y19665 , y19666 , y19667 , y19668 , y19669 , y19670 , y19671 , y19672 , y19673 , y19674 , y19675 , y19676 , y19677 , y19678 , y19679 , y19680 , y19681 , y19682 , y19683 , y19684 , y19685 , y19686 , y19687 , y19688 , y19689 , y19690 , y19691 , y19692 , y19693 , y19694 , y19695 , y19696 , y19697 , y19698 , y19699 , y19700 , y19701 , y19702 , y19703 , y19704 , y19705 , y19706 , y19707 , y19708 , y19709 , y19710 , y19711 , y19712 , y19713 , y19714 , y19715 , y19716 , y19717 , y19718 , y19719 , y19720 , y19721 , y19722 , y19723 , y19724 , y19725 , y19726 , y19727 , y19728 , y19729 , y19730 , y19731 , y19732 , y19733 , y19734 , y19735 , y19736 , y19737 , y19738 , y19739 , y19740 , y19741 , y19742 , y19743 , y19744 , y19745 , y19746 , y19747 , y19748 , y19749 , y19750 , y19751 , y19752 , y19753 , y19754 , y19755 , y19756 , y19757 , y19758 , y19759 , y19760 , y19761 , y19762 , y19763 , y19764 , y19765 , y19766 , y19767 , y19768 , y19769 , y19770 , y19771 , y19772 , y19773 , y19774 , y19775 , y19776 , y19777 , y19778 , y19779 , y19780 , y19781 , y19782 , y19783 , y19784 , y19785 , y19786 , y19787 , y19788 , y19789 , y19790 , y19791 , y19792 , y19793 , y19794 , y19795 , y19796 , y19797 , y19798 , y19799 , y19800 , y19801 , y19802 , y19803 , y19804 , y19805 , y19806 , y19807 , y19808 , y19809 , y19810 , y19811 , y19812 , y19813 , y19814 , y19815 , y19816 , y19817 , y19818 , y19819 , y19820 , y19821 , y19822 , y19823 , y19824 , y19825 , y19826 , y19827 , y19828 , y19829 , y19830 , y19831 , y19832 , y19833 , y19834 , y19835 , y19836 , y19837 , y19838 , y19839 , y19840 , y19841 , y19842 , y19843 , y19844 , y19845 , y19846 , y19847 , y19848 , y19849 , y19850 , y19851 , y19852 , y19853 , y19854 , y19855 , y19856 , y19857 , y19858 , y19859 , y19860 , y19861 , y19862 , y19863 , y19864 , y19865 , y19866 , y19867 , y19868 , y19869 , y19870 , y19871 , y19872 , y19873 , y19874 , y19875 , y19876 , y19877 , y19878 , y19879 , y19880 , y19881 , y19882 , y19883 , y19884 , y19885 , y19886 , y19887 , y19888 , y19889 , y19890 , y19891 , y19892 , y19893 , y19894 , y19895 , y19896 , y19897 , y19898 , y19899 , y19900 , y19901 , y19902 , y19903 , y19904 , y19905 , y19906 , y19907 , y19908 , y19909 , y19910 , y19911 , y19912 , y19913 , y19914 , y19915 , y19916 , y19917 , y19918 , y19919 , y19920 , y19921 , y19922 , y19923 , y19924 , y19925 , y19926 , y19927 , y19928 , y19929 , y19930 , y19931 , y19932 , y19933 , y19934 , y19935 , y19936 , y19937 , y19938 , y19939 , y19940 , y19941 , y19942 , y19943 , y19944 , y19945 , y19946 , y19947 , y19948 , y19949 , y19950 , y19951 , y19952 , y19953 , y19954 , y19955 , y19956 , y19957 , y19958 , y19959 , y19960 , y19961 , y19962 , y19963 , y19964 , y19965 , y19966 , y19967 , y19968 , y19969 , y19970 , y19971 , y19972 , y19973 , y19974 , y19975 , y19976 , y19977 , y19978 , y19979 , y19980 , y19981 , y19982 , y19983 , y19984 , y19985 , y19986 , y19987 , y19988 , y19989 , y19990 , y19991 , y19992 , y19993 , y19994 , y19995 , y19996 , y19997 , y19998 , y19999 , y20000 , y20001 , y20002 , y20003 , y20004 , y20005 , y20006 , y20007 , y20008 , y20009 , y20010 , y20011 , y20012 , y20013 , y20014 , y20015 , y20016 , y20017 , y20018 , y20019 , y20020 , y20021 , y20022 , y20023 , y20024 , y20025 , y20026 , y20027 , y20028 , y20029 , y20030 , y20031 , y20032 , y20033 , y20034 , y20035 , y20036 , y20037 , y20038 , y20039 , y20040 , y20041 , y20042 , y20043 , y20044 , y20045 , y20046 , y20047 , y20048 , y20049 , y20050 , y20051 , y20052 , y20053 , y20054 , y20055 , y20056 , y20057 , y20058 , y20059 , y20060 , y20061 , y20062 , y20063 , y20064 , y20065 , y20066 , y20067 , y20068 , y20069 , y20070 , y20071 , y20072 , y20073 , y20074 , y20075 , y20076 , y20077 , y20078 , y20079 , y20080 , y20081 , y20082 , y20083 , y20084 , y20085 , y20086 , y20087 , y20088 , y20089 , y20090 , y20091 , y20092 , y20093 , y20094 , y20095 , y20096 , y20097 , y20098 , y20099 , y20100 , y20101 , y20102 , y20103 , y20104 , y20105 , y20106 , y20107 , y20108 , y20109 , y20110 , y20111 , y20112 , y20113 , y20114 , y20115 , y20116 , y20117 , y20118 , y20119 , y20120 , y20121 , y20122 , y20123 , y20124 , y20125 , y20126 , y20127 , y20128 , y20129 , y20130 , y20131 , y20132 , y20133 , y20134 , y20135 , y20136 , y20137 , y20138 , y20139 , y20140 , y20141 , y20142 , y20143 , y20144 , y20145 , y20146 , y20147 , y20148 , y20149 , y20150 , y20151 , y20152 , y20153 , y20154 , y20155 , y20156 , y20157 , y20158 , y20159 , y20160 , y20161 , y20162 , y20163 , y20164 , y20165 , y20166 , y20167 , y20168 , y20169 , y20170 , y20171 , y20172 , y20173 , y20174 , y20175 , y20176 , y20177 , y20178 , y20179 , y20180 , y20181 , y20182 , y20183 , y20184 , y20185 , y20186 , y20187 , y20188 , y20189 , y20190 , y20191 , y20192 , y20193 , y20194 , y20195 , y20196 , y20197 , y20198 , y20199 , y20200 , y20201 , y20202 , y20203 , y20204 , y20205 , y20206 , y20207 , y20208 , y20209 , y20210 , y20211 , y20212 , y20213 , y20214 , y20215 , y20216 , y20217 , y20218 , y20219 , y20220 , y20221 , y20222 , y20223 , y20224 , y20225 , y20226 , y20227 , y20228 , y20229 , y20230 , y20231 , y20232 , y20233 , y20234 , y20235 , y20236 , y20237 , y20238 , y20239 , y20240 , y20241 , y20242 , y20243 , y20244 , y20245 , y20246 , y20247 , y20248 , y20249 , y20250 , y20251 , y20252 , y20253 , y20254 , y20255 , y20256 , y20257 , y20258 , y20259 , y20260 , y20261 , y20262 , y20263 , y20264 , y20265 , y20266 , y20267 , y20268 , y20269 , y20270 , y20271 , y20272 , y20273 , y20274 , y20275 , y20276 , y20277 , y20278 , y20279 , y20280 , y20281 , y20282 , y20283 , y20284 , y20285 , y20286 , y20287 , y20288 , y20289 , y20290 , y20291 , y20292 , y20293 , y20294 , y20295 , y20296 , y20297 , y20298 , y20299 , y20300 , y20301 , y20302 , y20303 , y20304 , y20305 , y20306 , y20307 , y20308 , y20309 , y20310 , y20311 , y20312 , y20313 , y20314 , y20315 , y20316 , y20317 , y20318 , y20319 , y20320 , y20321 , y20322 , y20323 , y20324 , y20325 , y20326 , y20327 , y20328 , y20329 , y20330 , y20331 , y20332 , y20333 , y20334 , y20335 , y20336 , y20337 , y20338 , y20339 , y20340 , y20341 , y20342 , y20343 , y20344 , y20345 , y20346 , y20347 , y20348 , y20349 , y20350 , y20351 , y20352 , y20353 , y20354 , y20355 , y20356 , y20357 , y20358 , y20359 , y20360 , y20361 , y20362 , y20363 , y20364 , y20365 , y20366 , y20367 , y20368 , y20369 , y20370 , y20371 , y20372 , y20373 , y20374 , y20375 , y20376 , y20377 , y20378 , y20379 , y20380 , y20381 , y20382 , y20383 , y20384 , y20385 , y20386 , y20387 , y20388 , y20389 , y20390 , y20391 , y20392 , y20393 , y20394 , y20395 , y20396 , y20397 , y20398 , y20399 , y20400 , y20401 , y20402 , y20403 , y20404 , y20405 , y20406 , y20407 , y20408 , y20409 , y20410 , y20411 , y20412 , y20413 , y20414 , y20415 , y20416 , y20417 , y20418 , y20419 , y20420 , y20421 , y20422 , y20423 , y20424 , y20425 , y20426 , y20427 , y20428 , y20429 , y20430 , y20431 , y20432 , y20433 , y20434 , y20435 , y20436 , y20437 , y20438 , y20439 , y20440 , y20441 , y20442 , y20443 , y20444 , y20445 , y20446 , y20447 , y20448 , y20449 , y20450 , y20451 , y20452 , y20453 , y20454 , y20455 , y20456 , y20457 , y20458 , y20459 , y20460 , y20461 , y20462 , y20463 , y20464 , y20465 , y20466 , y20467 , y20468 , y20469 , y20470 , y20471 , y20472 , y20473 , y20474 , y20475 , y20476 , y20477 , y20478 , y20479 , y20480 , y20481 , y20482 , y20483 , y20484 , y20485 , y20486 , y20487 , y20488 , y20489 , y20490 , y20491 , y20492 , y20493 , y20494 , y20495 , y20496 , y20497 , y20498 , y20499 , y20500 , y20501 , y20502 , y20503 , y20504 , y20505 , y20506 , y20507 , y20508 , y20509 , y20510 , y20511 , y20512 , y20513 , y20514 , y20515 , y20516 , y20517 , y20518 , y20519 , y20520 , y20521 , y20522 , y20523 , y20524 , y20525 , y20526 , y20527 , y20528 , y20529 , y20530 , y20531 , y20532 , y20533 , y20534 , y20535 , y20536 , y20537 , y20538 , y20539 , y20540 , y20541 , y20542 , y20543 , y20544 , y20545 , y20546 , y20547 , y20548 , y20549 , y20550 , y20551 , y20552 , y20553 , y20554 , y20555 , y20556 , y20557 , y20558 , y20559 , y20560 , y20561 , y20562 , y20563 , y20564 , y20565 , y20566 , y20567 , y20568 , y20569 , y20570 , y20571 , y20572 , y20573 , y20574 , y20575 , y20576 , y20577 , y20578 , y20579 , y20580 , y20581 , y20582 , y20583 , y20584 , y20585 , y20586 , y20587 , y20588 , y20589 , y20590 , y20591 , y20592 , y20593 , y20594 , y20595 , y20596 , y20597 , y20598 , y20599 , y20600 , y20601 , y20602 , y20603 , y20604 , y20605 , y20606 , y20607 , y20608 , y20609 , y20610 , y20611 , y20612 , y20613 , y20614 , y20615 , y20616 , y20617 , y20618 , y20619 , y20620 , y20621 , y20622 , y20623 , y20624 , y20625 , y20626 , y20627 , y20628 , y20629 , y20630 , y20631 , y20632 , y20633 , y20634 , y20635 , y20636 , y20637 , y20638 , y20639 , y20640 , y20641 , y20642 , y20643 , y20644 , y20645 , y20646 , y20647 , y20648 , y20649 , y20650 , y20651 , y20652 , y20653 , y20654 , y20655 , y20656 , y20657 , y20658 , y20659 , y20660 , y20661 , y20662 , y20663 , y20664 , y20665 , y20666 , y20667 , y20668 , y20669 , y20670 , y20671 , y20672 , y20673 , y20674 , y20675 , y20676 , y20677 , y20678 , y20679 , y20680 , y20681 , y20682 , y20683 , y20684 , y20685 , y20686 , y20687 , y20688 , y20689 , y20690 , y20691 , y20692 , y20693 , y20694 , y20695 , y20696 , y20697 , y20698 , y20699 , y20700 , y20701 , y20702 , y20703 , y20704 , y20705 , y20706 , y20707 , y20708 , y20709 , y20710 , y20711 , y20712 , y20713 , y20714 , y20715 , y20716 , y20717 , y20718 , y20719 , y20720 , y20721 , y20722 , y20723 , y20724 , y20725 , y20726 , y20727 , y20728 , y20729 , y20730 , y20731 , y20732 , y20733 , y20734 , y20735 , y20736 , y20737 , y20738 , y20739 , y20740 , y20741 , y20742 , y20743 , y20744 , y20745 , y20746 , y20747 , y20748 , y20749 , y20750 , y20751 , y20752 , y20753 , y20754 , y20755 , y20756 , y20757 , y20758 , y20759 , y20760 , y20761 , y20762 , y20763 , y20764 , y20765 , y20766 , y20767 , y20768 , y20769 , y20770 , y20771 , y20772 , y20773 , y20774 , y20775 , y20776 , y20777 , y20778 , y20779 , y20780 , y20781 , y20782 , y20783 , y20784 , y20785 , y20786 , y20787 , y20788 , y20789 , y20790 , y20791 , y20792 , y20793 , y20794 , y20795 , y20796 , y20797 , y20798 , y20799 , y20800 , y20801 , y20802 , y20803 , y20804 , y20805 , y20806 , y20807 , y20808 , y20809 , y20810 , y20811 , y20812 , y20813 , y20814 , y20815 , y20816 , y20817 , y20818 , y20819 , y20820 , y20821 , y20822 , y20823 , y20824 , y20825 , y20826 , y20827 , y20828 , y20829 , y20830 , y20831 , y20832 , y20833 , y20834 , y20835 , y20836 , y20837 , y20838 , y20839 , y20840 , y20841 , y20842 , y20843 , y20844 , y20845 , y20846 , y20847 , y20848 , y20849 , y20850 , y20851 , y20852 , y20853 , y20854 , y20855 , y20856 , y20857 , y20858 , y20859 , y20860 , y20861 , y20862 , y20863 , y20864 , y20865 , y20866 , y20867 , y20868 , y20869 , y20870 , y20871 , y20872 , y20873 , y20874 , y20875 , y20876 , y20877 , y20878 , y20879 , y20880 , y20881 , y20882 , y20883 , y20884 , y20885 , y20886 , y20887 , y20888 , y20889 , y20890 , y20891 , y20892 , y20893 , y20894 , y20895 , y20896 , y20897 , y20898 , y20899 , y20900 , y20901 , y20902 , y20903 , y20904 , y20905 , y20906 , y20907 , y20908 , y20909 , y20910 , y20911 , y20912 , y20913 , y20914 , y20915 , y20916 , y20917 , y20918 , y20919 , y20920 , y20921 , y20922 , y20923 , y20924 , y20925 , y20926 , y20927 , y20928 , y20929 , y20930 , y20931 , y20932 , y20933 , y20934 , y20935 , y20936 , y20937 , y20938 , y20939 , y20940 , y20941 , y20942 , y20943 , y20944 , y20945 , y20946 , y20947 , y20948 , y20949 , y20950 , y20951 , y20952 , y20953 , y20954 , y20955 , y20956 , y20957 , y20958 , y20959 , y20960 , y20961 , y20962 , y20963 , y20964 , y20965 , y20966 , y20967 , y20968 , y20969 , y20970 , y20971 , y20972 , y20973 , y20974 , y20975 , y20976 , y20977 , y20978 , y20979 , y20980 , y20981 , y20982 , y20983 , y20984 , y20985 , y20986 , y20987 , y20988 , y20989 , y20990 , y20991 , y20992 , y20993 , y20994 , y20995 , y20996 , y20997 , y20998 , y20999 , y21000 , y21001 , y21002 , y21003 , y21004 , y21005 , y21006 , y21007 , y21008 , y21009 , y21010 , y21011 , y21012 , y21013 , y21014 , y21015 , y21016 , y21017 , y21018 , y21019 , y21020 , y21021 , y21022 , y21023 , y21024 , y21025 , y21026 , y21027 , y21028 , y21029 , y21030 , y21031 , y21032 , y21033 , y21034 , y21035 , y21036 , y21037 , y21038 , y21039 , y21040 , y21041 , y21042 , y21043 , y21044 , y21045 , y21046 , y21047 , y21048 , y21049 , y21050 , y21051 , y21052 , y21053 , y21054 , y21055 , y21056 , y21057 , y21058 , y21059 , y21060 , y21061 , y21062 , y21063 , y21064 , y21065 , y21066 , y21067 , y21068 , y21069 , y21070 , y21071 , y21072 , y21073 , y21074 , y21075 , y21076 , y21077 , y21078 , y21079 , y21080 , y21081 , y21082 , y21083 , y21084 , y21085 , y21086 , y21087 , y21088 , y21089 , y21090 , y21091 , y21092 , y21093 , y21094 , y21095 , y21096 , y21097 , y21098 , y21099 , y21100 , y21101 , y21102 , y21103 , y21104 , y21105 , y21106 , y21107 , y21108 , y21109 , y21110 , y21111 , y21112 , y21113 , y21114 , y21115 , y21116 , y21117 , y21118 , y21119 , y21120 , y21121 , y21122 , y21123 , y21124 , y21125 , y21126 , y21127 , y21128 , y21129 , y21130 , y21131 , y21132 , y21133 , y21134 , y21135 , y21136 , y21137 , y21138 , y21139 , y21140 , y21141 , y21142 , y21143 , y21144 , y21145 , y21146 , y21147 , y21148 , y21149 , y21150 , y21151 , y21152 , y21153 , y21154 , y21155 , y21156 , y21157 , y21158 , y21159 , y21160 , y21161 , y21162 , y21163 , y21164 , y21165 , y21166 , y21167 , y21168 , y21169 , y21170 , y21171 , y21172 , y21173 , y21174 , y21175 , y21176 , y21177 , y21178 , y21179 , y21180 , y21181 , y21182 , y21183 , y21184 , y21185 , y21186 , y21187 , y21188 , y21189 , y21190 , y21191 , y21192 , y21193 , y21194 , y21195 , y21196 , y21197 , y21198 , y21199 , y21200 , y21201 , y21202 , y21203 , y21204 , y21205 , y21206 , y21207 , y21208 , y21209 , y21210 , y21211 , y21212 , y21213 , y21214 , y21215 , y21216 , y21217 , y21218 , y21219 , y21220 , y21221 , y21222 , y21223 , y21224 , y21225 , y21226 , y21227 , y21228 , y21229 , y21230 , y21231 , y21232 , y21233 , y21234 , y21235 , y21236 , y21237 , y21238 , y21239 , y21240 , y21241 , y21242 , y21243 , y21244 , y21245 , y21246 , y21247 , y21248 , y21249 , y21250 , y21251 , y21252 , y21253 , y21254 , y21255 , y21256 , y21257 , y21258 , y21259 , y21260 , y21261 , y21262 , y21263 , y21264 , y21265 , y21266 , y21267 , y21268 , y21269 , y21270 , y21271 , y21272 , y21273 , y21274 , y21275 , y21276 , y21277 , y21278 , y21279 , y21280 , y21281 , y21282 , y21283 , y21284 , y21285 , y21286 , y21287 , y21288 , y21289 , y21290 , y21291 , y21292 , y21293 , y21294 , y21295 , y21296 , y21297 , y21298 , y21299 , y21300 , y21301 , y21302 , y21303 , y21304 , y21305 , y21306 , y21307 , y21308 , y21309 , y21310 , y21311 , y21312 , y21313 , y21314 , y21315 , y21316 , y21317 , y21318 , y21319 , y21320 , y21321 , y21322 , y21323 , y21324 , y21325 , y21326 , y21327 , y21328 , y21329 , y21330 , y21331 , y21332 , y21333 , y21334 , y21335 , y21336 , y21337 , y21338 , y21339 , y21340 , y21341 , y21342 , y21343 , y21344 , y21345 , y21346 , y21347 , y21348 , y21349 , y21350 , y21351 , y21352 , y21353 , y21354 , y21355 , y21356 , y21357 , y21358 , y21359 , y21360 , y21361 , y21362 , y21363 , y21364 , y21365 , y21366 , y21367 , y21368 , y21369 , y21370 , y21371 , y21372 , y21373 , y21374 , y21375 , y21376 , y21377 , y21378 , y21379 , y21380 , y21381 , y21382 , y21383 , y21384 , y21385 , y21386 , y21387 , y21388 , y21389 , y21390 , y21391 , y21392 , y21393 , y21394 , y21395 , y21396 , y21397 , y21398 , y21399 , y21400 , y21401 , y21402 , y21403 , y21404 , y21405 , y21406 , y21407 , y21408 , y21409 , y21410 , y21411 , y21412 , y21413 , y21414 , y21415 , y21416 , y21417 , y21418 , y21419 , y21420 , y21421 , y21422 , y21423 , y21424 , y21425 , y21426 , y21427 , y21428 , y21429 , y21430 , y21431 , y21432 , y21433 , y21434 , y21435 , y21436 , y21437 , y21438 , y21439 , y21440 , y21441 , y21442 , y21443 , y21444 , y21445 , y21446 , y21447 , y21448 , y21449 , y21450 , y21451 , y21452 , y21453 , y21454 , y21455 , y21456 , y21457 , y21458 , y21459 , y21460 , y21461 , y21462 , y21463 , y21464 , y21465 , y21466 , y21467 , y21468 , y21469 , y21470 , y21471 , y21472 , y21473 , y21474 , y21475 , y21476 , y21477 , y21478 , y21479 , y21480 , y21481 , y21482 , y21483 , y21484 , y21485 , y21486 , y21487 , y21488 , y21489 , y21490 , y21491 , y21492 , y21493 , y21494 , y21495 , y21496 , y21497 , y21498 , y21499 , y21500 , y21501 , y21502 , y21503 , y21504 , y21505 , y21506 , y21507 , y21508 , y21509 , y21510 , y21511 , y21512 , y21513 , y21514 , y21515 , y21516 , y21517 , y21518 , y21519 , y21520 , y21521 , y21522 , y21523 , y21524 , y21525 , y21526 , y21527 , y21528 , y21529 , y21530 , y21531 , y21532 , y21533 , y21534 , y21535 , y21536 , y21537 , y21538 , y21539 , y21540 , y21541 , y21542 , y21543 , y21544 , y21545 , y21546 , y21547 , y21548 , y21549 , y21550 , y21551 , y21552 , y21553 , y21554 , y21555 , y21556 , y21557 , y21558 , y21559 , y21560 , y21561 , y21562 , y21563 , y21564 , y21565 , y21566 , y21567 , y21568 , y21569 , y21570 , y21571 , y21572 , y21573 , y21574 , y21575 , y21576 , y21577 , y21578 , y21579 , y21580 , y21581 , y21582 , y21583 , y21584 , y21585 , y21586 , y21587 , y21588 , y21589 , y21590 , y21591 , y21592 , y21593 , y21594 , y21595 , y21596 , y21597 , y21598 , y21599 , y21600 , y21601 , y21602 , y21603 , y21604 , y21605 , y21606 , y21607 , y21608 , y21609 , y21610 , y21611 , y21612 , y21613 , y21614 , y21615 , y21616 , y21617 , y21618 , y21619 , y21620 , y21621 , y21622 , y21623 , y21624 , y21625 , y21626 , y21627 , y21628 , y21629 , y21630 , y21631 , y21632 , y21633 , y21634 , y21635 , y21636 , y21637 , y21638 , y21639 , y21640 , y21641 , y21642 , y21643 , y21644 , y21645 , y21646 , y21647 , y21648 , y21649 , y21650 , y21651 , y21652 , y21653 , y21654 , y21655 , y21656 , y21657 , y21658 , y21659 , y21660 , y21661 , y21662 , y21663 , y21664 , y21665 , y21666 , y21667 , y21668 , y21669 , y21670 , y21671 , y21672 , y21673 , y21674 , y21675 , y21676 , y21677 , y21678 , y21679 , y21680 , y21681 , y21682 , y21683 , y21684 , y21685 , y21686 , y21687 , y21688 , y21689 , y21690 , y21691 , y21692 , y21693 , y21694 , y21695 , y21696 , y21697 , y21698 , y21699 , y21700 , y21701 , y21702 , y21703 , y21704 , y21705 , y21706 , y21707 , y21708 , y21709 , y21710 , y21711 , y21712 , y21713 , y21714 , y21715 , y21716 , y21717 , y21718 , y21719 , y21720 , y21721 , y21722 , y21723 , y21724 , y21725 , y21726 , y21727 , y21728 , y21729 , y21730 , y21731 , y21732 , y21733 , y21734 , y21735 , y21736 , y21737 , y21738 , y21739 , y21740 , y21741 , y21742 , y21743 , y21744 , y21745 , y21746 , y21747 , y21748 , y21749 , y21750 , y21751 , y21752 , y21753 , y21754 , y21755 , y21756 , y21757 , y21758 , y21759 , y21760 , y21761 , y21762 , y21763 , y21764 , y21765 , y21766 , y21767 , y21768 , y21769 , y21770 , y21771 , y21772 , y21773 , y21774 , y21775 , y21776 , y21777 , y21778 , y21779 , y21780 , y21781 , y21782 , y21783 , y21784 , y21785 , y21786 , y21787 , y21788 , y21789 , y21790 , y21791 , y21792 , y21793 , y21794 , y21795 , y21796 , y21797 , y21798 , y21799 , y21800 , y21801 , y21802 , y21803 , y21804 , y21805 , y21806 , y21807 , y21808 , y21809 , y21810 , y21811 , y21812 , y21813 , y21814 , y21815 , y21816 , y21817 , y21818 , y21819 , y21820 , y21821 , y21822 , y21823 , y21824 , y21825 , y21826 , y21827 , y21828 , y21829 , y21830 , y21831 , y21832 , y21833 , y21834 , y21835 , y21836 , y21837 , y21838 , y21839 , y21840 , y21841 , y21842 , y21843 , y21844 , y21845 , y21846 , y21847 , y21848 , y21849 , y21850 , y21851 , y21852 , y21853 , y21854 , y21855 , y21856 , y21857 , y21858 , y21859 , y21860 , y21861 , y21862 , y21863 , y21864 , y21865 , y21866 , y21867 , y21868 , y21869 , y21870 , y21871 , y21872 , y21873 , y21874 , y21875 , y21876 , y21877 , y21878 , y21879 , y21880 , y21881 , y21882 , y21883 , y21884 , y21885 , y21886 , y21887 , y21888 , y21889 , y21890 , y21891 , y21892 , y21893 , y21894 , y21895 , y21896 , y21897 , y21898 , y21899 , y21900 , y21901 , y21902 , y21903 , y21904 , y21905 , y21906 , y21907 , y21908 , y21909 , y21910 , y21911 , y21912 , y21913 , y21914 , y21915 , y21916 , y21917 , y21918 , y21919 , y21920 , y21921 , y21922 , y21923 , y21924 , y21925 , y21926 , y21927 , y21928 , y21929 , y21930 , y21931 , y21932 , y21933 , y21934 , y21935 , y21936 , y21937 , y21938 , y21939 , y21940 , y21941 , y21942 , y21943 , y21944 , y21945 , y21946 , y21947 , y21948 , y21949 , y21950 , y21951 , y21952 , y21953 , y21954 , y21955 , y21956 , y21957 , y21958 , y21959 , y21960 , y21961 , y21962 , y21963 , y21964 , y21965 , y21966 , y21967 , y21968 , y21969 , y21970 , y21971 , y21972 , y21973 , y21974 , y21975 , y21976 , y21977 , y21978 , y21979 , y21980 , y21981 , y21982 , y21983 , y21984 , y21985 , y21986 , y21987 , y21988 , y21989 , y21990 , y21991 , y21992 , y21993 , y21994 , y21995 , y21996 , y21997 , y21998 , y21999 , y22000 , y22001 , y22002 , y22003 , y22004 , y22005 , y22006 , y22007 , y22008 , y22009 , y22010 , y22011 , y22012 , y22013 , y22014 , y22015 , y22016 , y22017 , y22018 , y22019 , y22020 , y22021 , y22022 , y22023 , y22024 , y22025 , y22026 , y22027 , y22028 , y22029 , y22030 , y22031 , y22032 , y22033 , y22034 , y22035 , y22036 , y22037 , y22038 , y22039 , y22040 , y22041 , y22042 , y22043 , y22044 , y22045 , y22046 , y22047 , y22048 , y22049 , y22050 , y22051 , y22052 , y22053 , y22054 , y22055 , y22056 , y22057 , y22058 , y22059 , y22060 , y22061 , y22062 , y22063 , y22064 , y22065 , y22066 , y22067 , y22068 , y22069 , y22070 , y22071 , y22072 , y22073 , y22074 , y22075 , y22076 , y22077 , y22078 , y22079 , y22080 , y22081 , y22082 , y22083 , y22084 , y22085 , y22086 , y22087 , y22088 , y22089 , y22090 , y22091 , y22092 , y22093 , y22094 , y22095 , y22096 , y22097 , y22098 , y22099 , y22100 , y22101 , y22102 , y22103 , y22104 , y22105 , y22106 , y22107 , y22108 , y22109 , y22110 , y22111 , y22112 , y22113 , y22114 , y22115 , y22116 , y22117 , y22118 , y22119 , y22120 , y22121 , y22122 , y22123 , y22124 , y22125 , y22126 , y22127 , y22128 , y22129 , y22130 , y22131 , y22132 , y22133 , y22134 , y22135 , y22136 , y22137 , y22138 , y22139 , y22140 , y22141 , y22142 , y22143 , y22144 , y22145 , y22146 , y22147 , y22148 , y22149 , y22150 , y22151 , y22152 , y22153 , y22154 , y22155 , y22156 , y22157 , y22158 , y22159 , y22160 , y22161 , y22162 , y22163 , y22164 , y22165 , y22166 , y22167 , y22168 , y22169 , y22170 , y22171 , y22172 , y22173 , y22174 , y22175 , y22176 , y22177 , y22178 , y22179 , y22180 , y22181 , y22182 , y22183 , y22184 , y22185 , y22186 , y22187 , y22188 , y22189 , y22190 , y22191 , y22192 , y22193 , y22194 , y22195 , y22196 , y22197 , y22198 , y22199 , y22200 , y22201 , y22202 , y22203 , y22204 , y22205 , y22206 , y22207 , y22208 , y22209 , y22210 , y22211 , y22212 , y22213 , y22214 , y22215 , y22216 , y22217 , y22218 , y22219 , y22220 , y22221 , y22222 , y22223 , y22224 , y22225 , y22226 , y22227 , y22228 , y22229 , y22230 , y22231 , y22232 , y22233 , y22234 , y22235 , y22236 , y22237 , y22238 , y22239 , y22240 , y22241 , y22242 , y22243 , y22244 , y22245 , y22246 , y22247 , y22248 , y22249 , y22250 , y22251 , y22252 , y22253 , y22254 , y22255 , y22256 , y22257 , y22258 , y22259 , y22260 , y22261 , y22262 , y22263 , y22264 , y22265 , y22266 , y22267 , y22268 , y22269 , y22270 , y22271 , y22272 , y22273 , y22274 , y22275 , y22276 , y22277 , y22278 , y22279 , y22280 , y22281 , y22282 , y22283 , y22284 , y22285 , y22286 , y22287 , y22288 , y22289 , y22290 , y22291 , y22292 , y22293 , y22294 , y22295 , y22296 , y22297 , y22298 , y22299 , y22300 , y22301 , y22302 , y22303 , y22304 , y22305 , y22306 , y22307 , y22308 , y22309 , y22310 , y22311 , y22312 , y22313 , y22314 , y22315 , y22316 , y22317 , y22318 , y22319 , y22320 , y22321 , y22322 , y22323 , y22324 , y22325 , y22326 , y22327 , y22328 , y22329 , y22330 , y22331 , y22332 , y22333 , y22334 , y22335 , y22336 , y22337 , y22338 , y22339 , y22340 , y22341 , y22342 , y22343 , y22344 , y22345 , y22346 , y22347 , y22348 , y22349 , y22350 , y22351 , y22352 , y22353 , y22354 , y22355 , y22356 , y22357 , y22358 , y22359 , y22360 , y22361 , y22362 , y22363 , y22364 , y22365 , y22366 , y22367 , y22368 , y22369 , y22370 , y22371 , y22372 , y22373 , y22374 , y22375 , y22376 , y22377 , y22378 , y22379 , y22380 , y22381 , y22382 , y22383 , y22384 , y22385 , y22386 , y22387 , y22388 , y22389 , y22390 , y22391 , y22392 , y22393 , y22394 , y22395 , y22396 , y22397 , y22398 , y22399 , y22400 , y22401 , y22402 , y22403 , y22404 , y22405 , y22406 , y22407 , y22408 , y22409 , y22410 , y22411 , y22412 , y22413 , y22414 , y22415 , y22416 , y22417 , y22418 , y22419 , y22420 , y22421 , y22422 , y22423 , y22424 , y22425 , y22426 , y22427 , y22428 , y22429 , y22430 , y22431 , y22432 , y22433 , y22434 , y22435 , y22436 , y22437 , y22438 , y22439 , y22440 , y22441 , y22442 , y22443 , y22444 , y22445 , y22446 , y22447 , y22448 , y22449 , y22450 , y22451 , y22452 , y22453 , y22454 , y22455 , y22456 , y22457 , y22458 , y22459 , y22460 , y22461 , y22462 , y22463 , y22464 , y22465 , y22466 , y22467 , y22468 , y22469 , y22470 , y22471 , y22472 , y22473 , y22474 , y22475 , y22476 , y22477 , y22478 , y22479 , y22480 , y22481 , y22482 , y22483 , y22484 , y22485 , y22486 , y22487 , y22488 , y22489 , y22490 , y22491 , y22492 , y22493 , y22494 , y22495 , y22496 , y22497 , y22498 , y22499 , y22500 , y22501 , y22502 , y22503 , y22504 , y22505 , y22506 , y22507 , y22508 , y22509 , y22510 , y22511 , y22512 , y22513 , y22514 , y22515 , y22516 , y22517 , y22518 , y22519 , y22520 , y22521 , y22522 , y22523 , y22524 , y22525 , y22526 , y22527 , y22528 , y22529 , y22530 , y22531 , y22532 , y22533 , y22534 , y22535 , y22536 , y22537 , y22538 , y22539 , y22540 , y22541 , y22542 , y22543 , y22544 , y22545 , y22546 , y22547 , y22548 , y22549 , y22550 , y22551 , y22552 , y22553 , y22554 , y22555 , y22556 , y22557 , y22558 , y22559 , y22560 , y22561 , y22562 , y22563 , y22564 , y22565 , y22566 , y22567 , y22568 , y22569 , y22570 , y22571 , y22572 , y22573 , y22574 , y22575 , y22576 , y22577 , y22578 , y22579 , y22580 , y22581 , y22582 , y22583 , y22584 , y22585 , y22586 , y22587 , y22588 , y22589 , y22590 , y22591 , y22592 , y22593 , y22594 , y22595 , y22596 , y22597 , y22598 , y22599 , y22600 , y22601 , y22602 , y22603 , y22604 , y22605 , y22606 , y22607 , y22608 , y22609 , y22610 , y22611 , y22612 , y22613 , y22614 , y22615 , y22616 , y22617 , y22618 , y22619 , y22620 , y22621 , y22622 , y22623 , y22624 , y22625 , y22626 , y22627 , y22628 , y22629 , y22630 , y22631 , y22632 , y22633 , y22634 , y22635 , y22636 , y22637 , y22638 , y22639 , y22640 , y22641 , y22642 , y22643 , y22644 , y22645 , y22646 , y22647 , y22648 , y22649 , y22650 , y22651 , y22652 , y22653 , y22654 , y22655 , y22656 , y22657 , y22658 , y22659 , y22660 , y22661 , y22662 , y22663 , y22664 , y22665 , y22666 , y22667 , y22668 , y22669 , y22670 , y22671 , y22672 , y22673 , y22674 , y22675 , y22676 , y22677 , y22678 , y22679 , y22680 , y22681 , y22682 , y22683 , y22684 , y22685 , y22686 , y22687 , y22688 , y22689 , y22690 , y22691 , y22692 , y22693 , y22694 , y22695 , y22696 , y22697 , y22698 , y22699 , y22700 , y22701 , y22702 , y22703 , y22704 , y22705 , y22706 , y22707 , y22708 , y22709 , y22710 , y22711 , y22712 , y22713 , y22714 , y22715 , y22716 , y22717 , y22718 , y22719 , y22720 , y22721 , y22722 , y22723 , y22724 , y22725 , y22726 , y22727 , y22728 , y22729 , y22730 , y22731 , y22732 , y22733 , y22734 , y22735 , y22736 , y22737 , y22738 , y22739 , y22740 , y22741 , y22742 , y22743 , y22744 , y22745 , y22746 , y22747 , y22748 , y22749 , y22750 , y22751 , y22752 , y22753 , y22754 , y22755 , y22756 , y22757 , y22758 , y22759 , y22760 , y22761 , y22762 , y22763 , y22764 , y22765 , y22766 , y22767 , y22768 , y22769 , y22770 , y22771 , y22772 , y22773 , y22774 , y22775 , y22776 , y22777 , y22778 , y22779 , y22780 , y22781 , y22782 , y22783 , y22784 , y22785 , y22786 , y22787 , y22788 , y22789 , y22790 , y22791 , y22792 , y22793 , y22794 , y22795 , y22796 , y22797 , y22798 , y22799 , y22800 , y22801 , y22802 , y22803 , y22804 , y22805 , y22806 , y22807 , y22808 , y22809 , y22810 , y22811 , y22812 , y22813 , y22814 , y22815 , y22816 , y22817 , y22818 , y22819 , y22820 , y22821 , y22822 , y22823 , y22824 , y22825 , y22826 , y22827 , y22828 , y22829 , y22830 , y22831 , y22832 , y22833 , y22834 , y22835 , y22836 , y22837 , y22838 , y22839 , y22840 , y22841 , y22842 , y22843 , y22844 , y22845 , y22846 , y22847 , y22848 , y22849 , y22850 , y22851 , y22852 , y22853 , y22854 , y22855 , y22856 , y22857 , y22858 , y22859 , y22860 , y22861 , y22862 , y22863 , y22864 , y22865 , y22866 , y22867 , y22868 , y22869 , y22870 , y22871 , y22872 , y22873 , y22874 , y22875 , y22876 , y22877 , y22878 , y22879 , y22880 , y22881 , y22882 , y22883 , y22884 , y22885 , y22886 , y22887 , y22888 , y22889 , y22890 , y22891 , y22892 , y22893 , y22894 , y22895 , y22896 , y22897 , y22898 , y22899 , y22900 , y22901 , y22902 , y22903 , y22904 , y22905 , y22906 , y22907 , y22908 , y22909 , y22910 , y22911 , y22912 , y22913 , y22914 , y22915 , y22916 , y22917 , y22918 , y22919 , y22920 , y22921 , y22922 , y22923 , y22924 , y22925 , y22926 , y22927 , y22928 , y22929 , y22930 , y22931 , y22932 , y22933 , y22934 , y22935 , y22936 , y22937 , y22938 , y22939 , y22940 , y22941 , y22942 , y22943 , y22944 , y22945 , y22946 , y22947 , y22948 , y22949 , y22950 , y22951 , y22952 , y22953 , y22954 , y22955 , y22956 , y22957 , y22958 , y22959 , y22960 , y22961 , y22962 , y22963 , y22964 , y22965 , y22966 , y22967 , y22968 , y22969 , y22970 , y22971 , y22972 , y22973 , y22974 , y22975 , y22976 , y22977 , y22978 , y22979 , y22980 , y22981 , y22982 , y22983 , y22984 , y22985 , y22986 , y22987 , y22988 , y22989 , y22990 , y22991 , y22992 , y22993 , y22994 , y22995 , y22996 , y22997 , y22998 , y22999 , y23000 , y23001 , y23002 , y23003 , y23004 , y23005 , y23006 , y23007 , y23008 , y23009 , y23010 , y23011 , y23012 , y23013 , y23014 , y23015 , y23016 , y23017 , y23018 , y23019 , y23020 , y23021 , y23022 , y23023 , y23024 , y23025 , y23026 , y23027 , y23028 , y23029 , y23030 , y23031 , y23032 , y23033 , y23034 , y23035 , y23036 , y23037 , y23038 , y23039 , y23040 , y23041 , y23042 , y23043 , y23044 , y23045 , y23046 , y23047 , y23048 , y23049 , y23050 , y23051 , y23052 , y23053 , y23054 , y23055 , y23056 , y23057 , y23058 , y23059 , y23060 , y23061 , y23062 , y23063 , y23064 , y23065 , y23066 , y23067 , y23068 , y23069 , y23070 , y23071 , y23072 , y23073 , y23074 , y23075 , y23076 , y23077 , y23078 , y23079 , y23080 , y23081 , y23082 , y23083 , y23084 , y23085 , y23086 , y23087 , y23088 , y23089 , y23090 , y23091 , y23092 , y23093 , y23094 , y23095 , y23096 , y23097 , y23098 , y23099 , y23100 , y23101 , y23102 , y23103 , y23104 , y23105 , y23106 , y23107 , y23108 , y23109 , y23110 , y23111 , y23112 , y23113 , y23114 , y23115 , y23116 , y23117 , y23118 , y23119 , y23120 , y23121 , y23122 , y23123 , y23124 , y23125 , y23126 , y23127 , y23128 , y23129 , y23130 , y23131 , y23132 , y23133 , y23134 , y23135 , y23136 , y23137 , y23138 , y23139 , y23140 , y23141 , y23142 , y23143 , y23144 , y23145 , y23146 , y23147 , y23148 , y23149 , y23150 , y23151 , y23152 , y23153 , y23154 , y23155 , y23156 , y23157 , y23158 , y23159 , y23160 , y23161 , y23162 , y23163 , y23164 , y23165 , y23166 , y23167 , y23168 , y23169 , y23170 , y23171 , y23172 , y23173 , y23174 , y23175 , y23176 , y23177 , y23178 , y23179 , y23180 , y23181 , y23182 , y23183 , y23184 , y23185 , y23186 , y23187 , y23188 , y23189 , y23190 , y23191 , y23192 , y23193 , y23194 , y23195 , y23196 , y23197 , y23198 , y23199 , y23200 , y23201 , y23202 , y23203 , y23204 , y23205 , y23206 , y23207 , y23208 , y23209 , y23210 , y23211 , y23212 , y23213 , y23214 , y23215 , y23216 , y23217 , y23218 , y23219 , y23220 , y23221 , y23222 , y23223 , y23224 , y23225 , y23226 , y23227 , y23228 , y23229 , y23230 , y23231 , y23232 , y23233 , y23234 , y23235 , y23236 , y23237 , y23238 , y23239 , y23240 , y23241 , y23242 , y23243 , y23244 , y23245 , y23246 , y23247 , y23248 , y23249 , y23250 , y23251 , y23252 , y23253 , y23254 , y23255 , y23256 , y23257 , y23258 , y23259 , y23260 , y23261 , y23262 , y23263 , y23264 , y23265 , y23266 , y23267 , y23268 , y23269 , y23270 , y23271 , y23272 , y23273 , y23274 , y23275 , y23276 , y23277 , y23278 , y23279 , y23280 , y23281 , y23282 , y23283 , y23284 , y23285 , y23286 , y23287 , y23288 , y23289 , y23290 , y23291 , y23292 , y23293 , y23294 , y23295 , y23296 , y23297 , y23298 , y23299 , y23300 , y23301 , y23302 , y23303 , y23304 , y23305 , y23306 , y23307 , y23308 , y23309 , y23310 , y23311 , y23312 , y23313 , y23314 , y23315 , y23316 , y23317 , y23318 , y23319 , y23320 , y23321 , y23322 , y23323 , y23324 , y23325 , y23326 , y23327 , y23328 , y23329 , y23330 , y23331 , y23332 , y23333 , y23334 , y23335 , y23336 , y23337 , y23338 , y23339 , y23340 , y23341 , y23342 , y23343 , y23344 , y23345 , y23346 , y23347 , y23348 , y23349 , y23350 , y23351 , y23352 , y23353 , y23354 , y23355 , y23356 , y23357 , y23358 , y23359 , y23360 , y23361 , y23362 , y23363 , y23364 , y23365 , y23366 , y23367 , y23368 , y23369 , y23370 , y23371 , y23372 , y23373 , y23374 , y23375 , y23376 , y23377 , y23378 , y23379 , y23380 , y23381 , y23382 , y23383 , y23384 , y23385 , y23386 , y23387 , y23388 , y23389 , y23390 , y23391 , y23392 , y23393 , y23394 , y23395 , y23396 , y23397 , y23398 , y23399 , y23400 , y23401 , y23402 , y23403 , y23404 , y23405 , y23406 , y23407 , y23408 , y23409 , y23410 , y23411 , y23412 , y23413 , y23414 , y23415 , y23416 , y23417 , y23418 , y23419 , y23420 , y23421 , y23422 , y23423 , y23424 , y23425 , y23426 , y23427 , y23428 , y23429 , y23430 , y23431 , y23432 , y23433 , y23434 , y23435 , y23436 , y23437 , y23438 , y23439 , y23440 , y23441 , y23442 , y23443 , y23444 , y23445 , y23446 , y23447 , y23448 , y23449 , y23450 , y23451 , y23452 , y23453 , y23454 , y23455 , y23456 , y23457 , y23458 , y23459 , y23460 , y23461 , y23462 , y23463 , y23464 , y23465 , y23466 , y23467 , y23468 , y23469 , y23470 , y23471 , y23472 , y23473 , y23474 , y23475 , y23476 , y23477 , y23478 , y23479 , y23480 , y23481 , y23482 , y23483 , y23484 , y23485 , y23486 , y23487 , y23488 , y23489 , y23490 , y23491 , y23492 , y23493 , y23494 , y23495 , y23496 , y23497 , y23498 , y23499 , y23500 , y23501 , y23502 , y23503 , y23504 , y23505 , y23506 , y23507 , y23508 , y23509 , y23510 , y23511 , y23512 , y23513 , y23514 , y23515 , y23516 , y23517 , y23518 , y23519 , y23520 , y23521 , y23522 , y23523 , y23524 , y23525 , y23526 , y23527 , y23528 , y23529 , y23530 , y23531 , y23532 , y23533 , y23534 , y23535 , y23536 , y23537 , y23538 , y23539 , y23540 , y23541 , y23542 , y23543 , y23544 , y23545 , y23546 , y23547 , y23548 , y23549 , y23550 , y23551 , y23552 , y23553 , y23554 , y23555 , y23556 , y23557 , y23558 , y23559 , y23560 , y23561 , y23562 , y23563 , y23564 , y23565 , y23566 , y23567 , y23568 , y23569 , y23570 , y23571 , y23572 , y23573 , y23574 , y23575 , y23576 , y23577 , y23578 , y23579 , y23580 , y23581 , y23582 , y23583 , y23584 , y23585 , y23586 , y23587 , y23588 , y23589 , y23590 , y23591 , y23592 , y23593 , y23594 , y23595 , y23596 , y23597 , y23598 , y23599 , y23600 , y23601 , y23602 , y23603 , y23604 , y23605 , y23606 , y23607 , y23608 , y23609 , y23610 , y23611 , y23612 , y23613 , y23614 , y23615 , y23616 , y23617 , y23618 , y23619 , y23620 , y23621 , y23622 , y23623 , y23624 , y23625 , y23626 , y23627 , y23628 , y23629 , y23630 , y23631 , y23632 , y23633 , y23634 , y23635 , y23636 , y23637 , y23638 , y23639 , y23640 , y23641 , y23642 , y23643 , y23644 , y23645 , y23646 , y23647 , y23648 , y23649 , y23650 , y23651 , y23652 , y23653 , y23654 , y23655 , y23656 , y23657 , y23658 , y23659 , y23660 , y23661 , y23662 , y23663 , y23664 , y23665 , y23666 , y23667 , y23668 , y23669 , y23670 , y23671 , y23672 , y23673 , y23674 , y23675 , y23676 , y23677 , y23678 , y23679 , y23680 , y23681 , y23682 , y23683 , y23684 , y23685 , y23686 , y23687 , y23688 , y23689 , y23690 , y23691 , y23692 , y23693 , y23694 , y23695 , y23696 , y23697 , y23698 , y23699 , y23700 , y23701 , y23702 , y23703 , y23704 , y23705 , y23706 , y23707 , y23708 , y23709 , y23710 , y23711 , y23712 , y23713 , y23714 , y23715 , y23716 , y23717 , y23718 , y23719 , y23720 , y23721 , y23722 , y23723 , y23724 , y23725 , y23726 , y23727 , y23728 , y23729 , y23730 , y23731 , y23732 , y23733 , y23734 , y23735 , y23736 , y23737 , y23738 , y23739 , y23740 , y23741 , y23742 , y23743 , y23744 , y23745 , y23746 , y23747 , y23748 , y23749 , y23750 , y23751 , y23752 , y23753 , y23754 , y23755 , y23756 , y23757 , y23758 , y23759 , y23760 , y23761 , y23762 , y23763 , y23764 , y23765 , y23766 , y23767 , y23768 , y23769 , y23770 , y23771 , y23772 , y23773 , y23774 , y23775 , y23776 , y23777 , y23778 , y23779 , y23780 , y23781 , y23782 , y23783 , y23784 , y23785 , y23786 , y23787 , y23788 , y23789 , y23790 , y23791 , y23792 , y23793 , y23794 , y23795 , y23796 , y23797 , y23798 , y23799 , y23800 , y23801 , y23802 , y23803 , y23804 , y23805 , y23806 , y23807 , y23808 , y23809 , y23810 , y23811 , y23812 , y23813 , y23814 , y23815 , y23816 , y23817 , y23818 , y23819 , y23820 , y23821 , y23822 , y23823 , y23824 , y23825 , y23826 , y23827 , y23828 , y23829 , y23830 , y23831 , y23832 , y23833 , y23834 , y23835 , y23836 , y23837 , y23838 , y23839 , y23840 , y23841 , y23842 , y23843 , y23844 , y23845 , y23846 , y23847 , y23848 , y23849 , y23850 , y23851 , y23852 , y23853 , y23854 , y23855 , y23856 , y23857 , y23858 , y23859 , y23860 , y23861 , y23862 , y23863 , y23864 , y23865 , y23866 , y23867 , y23868 , y23869 , y23870 , y23871 , y23872 , y23873 , y23874 , y23875 , y23876 , y23877 , y23878 , y23879 , y23880 , y23881 , y23882 , y23883 , y23884 , y23885 , y23886 , y23887 , y23888 , y23889 , y23890 , y23891 , y23892 , y23893 , y23894 , y23895 , y23896 , y23897 , y23898 , y23899 , y23900 , y23901 , y23902 , y23903 , y23904 , y23905 , y23906 , y23907 , y23908 , y23909 , y23910 , y23911 , y23912 , y23913 , y23914 , y23915 , y23916 , y23917 , y23918 , y23919 , y23920 , y23921 , y23922 , y23923 , y23924 , y23925 , y23926 , y23927 , y23928 , y23929 , y23930 , y23931 , y23932 , y23933 , y23934 , y23935 , y23936 , y23937 , y23938 , y23939 , y23940 , y23941 , y23942 , y23943 , y23944 , y23945 , y23946 , y23947 , y23948 , y23949 , y23950 , y23951 , y23952 , y23953 , y23954 , y23955 , y23956 , y23957 , y23958 , y23959 , y23960 , y23961 , y23962 , y23963 , y23964 , y23965 , y23966 , y23967 , y23968 , y23969 , y23970 , y23971 , y23972 , y23973 , y23974 , y23975 , y23976 , y23977 , y23978 , y23979 , y23980 , y23981 , y23982 , y23983 , y23984 , y23985 , y23986 , y23987 , y23988 , y23989 , y23990 , y23991 , y23992 , y23993 , y23994 , y23995 , y23996 , y23997 , y23998 , y23999 , y24000 , y24001 , y24002 , y24003 , y24004 , y24005 , y24006 , y24007 , y24008 , y24009 , y24010 , y24011 , y24012 , y24013 , y24014 , y24015 , y24016 , y24017 , y24018 , y24019 , y24020 , y24021 , y24022 , y24023 , y24024 , y24025 , y24026 , y24027 , y24028 , y24029 , y24030 , y24031 , y24032 , y24033 , y24034 , y24035 , y24036 , y24037 , y24038 , y24039 , y24040 , y24041 , y24042 , y24043 , y24044 , y24045 , y24046 , y24047 , y24048 , y24049 , y24050 , y24051 , y24052 , y24053 , y24054 , y24055 , y24056 , y24057 , y24058 , y24059 , y24060 , y24061 , y24062 , y24063 , y24064 , y24065 , y24066 , y24067 , y24068 , y24069 , y24070 , y24071 , y24072 , y24073 , y24074 , y24075 , y24076 , y24077 , y24078 , y24079 , y24080 , y24081 , y24082 , y24083 , y24084 , y24085 , y24086 , y24087 , y24088 , y24089 , y24090 , y24091 , y24092 , y24093 , y24094 , y24095 , y24096 , y24097 , y24098 , y24099 , y24100 , y24101 , y24102 , y24103 , y24104 , y24105 , y24106 , y24107 , y24108 , y24109 , y24110 , y24111 , y24112 , y24113 , y24114 , y24115 , y24116 , y24117 , y24118 , y24119 , y24120 , y24121 , y24122 , y24123 , y24124 , y24125 , y24126 , y24127 , y24128 , y24129 , y24130 , y24131 , y24132 , y24133 , y24134 , y24135 , y24136 , y24137 , y24138 , y24139 , y24140 , y24141 , y24142 , y24143 , y24144 , y24145 , y24146 , y24147 , y24148 , y24149 , y24150 , y24151 , y24152 , y24153 , y24154 , y24155 , y24156 , y24157 , y24158 , y24159 , y24160 , y24161 , y24162 , y24163 , y24164 , y24165 , y24166 , y24167 , y24168 , y24169 , y24170 , y24171 , y24172 , y24173 , y24174 , y24175 , y24176 , y24177 , y24178 , y24179 , y24180 , y24181 , y24182 , y24183 , y24184 , y24185 , y24186 , y24187 , y24188 , y24189 , y24190 , y24191 , y24192 , y24193 , y24194 , y24195 , y24196 , y24197 , y24198 , y24199 , y24200 , y24201 , y24202 , y24203 , y24204 , y24205 , y24206 , y24207 , y24208 , y24209 , y24210 , y24211 , y24212 , y24213 , y24214 , y24215 , y24216 , y24217 , y24218 , y24219 , y24220 , y24221 , y24222 , y24223 , y24224 , y24225 , y24226 , y24227 , y24228 , y24229 , y24230 , y24231 , y24232 , y24233 , y24234 , y24235 , y24236 , y24237 , y24238 , y24239 , y24240 , y24241 , y24242 , y24243 , y24244 , y24245 , y24246 , y24247 , y24248 , y24249 , y24250 , y24251 , y24252 , y24253 , y24254 , y24255 , y24256 , y24257 , y24258 , y24259 , y24260 , y24261 , y24262 , y24263 , y24264 , y24265 , y24266 , y24267 , y24268 , y24269 , y24270 , y24271 , y24272 , y24273 , y24274 , y24275 , y24276 , y24277 , y24278 , y24279 , y24280 , y24281 , y24282 , y24283 , y24284 , y24285 , y24286 , y24287 , y24288 , y24289 , y24290 , y24291 , y24292 , y24293 , y24294 , y24295 , y24296 , y24297 , y24298 , y24299 , y24300 , y24301 , y24302 , y24303 , y24304 , y24305 , y24306 , y24307 , y24308 , y24309 , y24310 , y24311 , y24312 , y24313 , y24314 , y24315 , y24316 , y24317 , y24318 , y24319 , y24320 , y24321 , y24322 , y24323 , y24324 , y24325 , y24326 , y24327 , y24328 , y24329 , y24330 , y24331 , y24332 , y24333 , y24334 , y24335 , y24336 , y24337 , y24338 , y24339 , y24340 , y24341 , y24342 , y24343 , y24344 , y24345 , y24346 , y24347 , y24348 , y24349 , y24350 , y24351 , y24352 , y24353 , y24354 , y24355 , y24356 , y24357 , y24358 , y24359 , y24360 , y24361 , y24362 , y24363 , y24364 , y24365 , y24366 , y24367 , y24368 , y24369 , y24370 , y24371 , y24372 , y24373 , y24374 , y24375 , y24376 , y24377 , y24378 , y24379 , y24380 , y24381 , y24382 , y24383 , y24384 , y24385 , y24386 , y24387 , y24388 , y24389 , y24390 , y24391 , y24392 , y24393 , y24394 , y24395 , y24396 , y24397 , y24398 , y24399 , y24400 , y24401 , y24402 , y24403 , y24404 , y24405 , y24406 , y24407 , y24408 , y24409 , y24410 , y24411 , y24412 , y24413 , y24414 , y24415 , y24416 , y24417 , y24418 , y24419 , y24420 , y24421 , y24422 , y24423 , y24424 , y24425 , y24426 , y24427 , y24428 , y24429 , y24430 , y24431 , y24432 , y24433 , y24434 , y24435 , y24436 , y24437 , y24438 , y24439 , y24440 , y24441 , y24442 , y24443 , y24444 , y24445 , y24446 , y24447 , y24448 , y24449 , y24450 , y24451 , y24452 , y24453 , y24454 , y24455 , y24456 , y24457 , y24458 , y24459 , y24460 , y24461 , y24462 , y24463 , y24464 , y24465 , y24466 , y24467 , y24468 , y24469 , y24470 , y24471 , y24472 , y24473 , y24474 , y24475 , y24476 , y24477 , y24478 , y24479 , y24480 , y24481 , y24482 , y24483 , y24484 , y24485 , y24486 , y24487 , y24488 , y24489 , y24490 , y24491 , y24492 , y24493 , y24494 , y24495 , y24496 , y24497 , y24498 , y24499 , y24500 , y24501 , y24502 , y24503 , y24504 , y24505 , y24506 , y24507 , y24508 , y24509 , y24510 , y24511 , y24512 , y24513 , y24514 , y24515 , y24516 , y24517 , y24518 , y24519 , y24520 , y24521 , y24522 , y24523 , y24524 , y24525 , y24526 , y24527 , y24528 , y24529 , y24530 , y24531 , y24532 , y24533 , y24534 , y24535 , y24536 , y24537 , y24538 , y24539 , y24540 , y24541 , y24542 , y24543 , y24544 , y24545 , y24546 , y24547 , y24548 , y24549 , y24550 , y24551 , y24552 , y24553 , y24554 , y24555 , y24556 , y24557 , y24558 , y24559 , y24560 , y24561 , y24562 , y24563 , y24564 , y24565 , y24566 , y24567 , y24568 , y24569 , y24570 , y24571 , y24572 , y24573 , y24574 , y24575 , y24576 , y24577 , y24578 , y24579 , y24580 , y24581 , y24582 , y24583 , y24584 , y24585 , y24586 , y24587 , y24588 , y24589 , y24590 , y24591 , y24592 , y24593 , y24594 , y24595 , y24596 , y24597 , y24598 , y24599 , y24600 , y24601 , y24602 , y24603 , y24604 , y24605 , y24606 , y24607 , y24608 , y24609 , y24610 , y24611 , y24612 , y24613 , y24614 , y24615 , y24616 , y24617 , y24618 , y24619 , y24620 , y24621 , y24622 , y24623 , y24624 , y24625 , y24626 , y24627 , y24628 , y24629 , y24630 , y24631 , y24632 , y24633 , y24634 , y24635 , y24636 , y24637 , y24638 , y24639 , y24640 , y24641 , y24642 , y24643 , y24644 , y24645 , y24646 , y24647 , y24648 , y24649 , y24650 , y24651 , y24652 , y24653 , y24654 , y24655 , y24656 , y24657 , y24658 , y24659 , y24660 , y24661 , y24662 , y24663 , y24664 , y24665 , y24666 , y24667 , y24668 , y24669 , y24670 , y24671 , y24672 , y24673 , y24674 , y24675 , y24676 , y24677 , y24678 , y24679 , y24680 , y24681 , y24682 , y24683 , y24684 , y24685 , y24686 , y24687 , y24688 , y24689 , y24690 , y24691 , y24692 , y24693 , y24694 , y24695 , y24696 , y24697 , y24698 , y24699 , y24700 , y24701 , y24702 , y24703 , y24704 , y24705 , y24706 , y24707 , y24708 , y24709 , y24710 , y24711 , y24712 , y24713 , y24714 , y24715 , y24716 , y24717 , y24718 , y24719 , y24720 , y24721 , y24722 , y24723 , y24724 , y24725 , y24726 , y24727 , y24728 , y24729 , y24730 , y24731 , y24732 , y24733 , y24734 , y24735 , y24736 , y24737 , y24738 , y24739 , y24740 , y24741 , y24742 , y24743 , y24744 , y24745 , y24746 , y24747 , y24748 , y24749 , y24750 , y24751 , y24752 , y24753 , y24754 , y24755 , y24756 , y24757 , y24758 , y24759 , y24760 , y24761 , y24762 , y24763 , y24764 , y24765 , y24766 , y24767 , y24768 , y24769 , y24770 , y24771 , y24772 , y24773 , y24774 , y24775 , y24776 , y24777 , y24778 , y24779 , y24780 , y24781 , y24782 , y24783 , y24784 , y24785 , y24786 , y24787 , y24788 , y24789 , y24790 , y24791 , y24792 , y24793 , y24794 , y24795 , y24796 , y24797 , y24798 , y24799 , y24800 , y24801 , y24802 , y24803 , y24804 , y24805 , y24806 , y24807 , y24808 , y24809 , y24810 , y24811 , y24812 , y24813 , y24814 , y24815 , y24816 , y24817 , y24818 , y24819 , y24820 , y24821 , y24822 , y24823 , y24824 , y24825 , y24826 , y24827 , y24828 , y24829 , y24830 , y24831 , y24832 , y24833 , y24834 , y24835 , y24836 , y24837 , y24838 , y24839 , y24840 , y24841 , y24842 , y24843 , y24844 , y24845 , y24846 , y24847 , y24848 , y24849 , y24850 , y24851 , y24852 , y24853 , y24854 , y24855 , y24856 , y24857 , y24858 , y24859 , y24860 , y24861 , y24862 , y24863 , y24864 , y24865 , y24866 , y24867 , y24868 , y24869 , y24870 , y24871 , y24872 , y24873 , y24874 , y24875 , y24876 , y24877 , y24878 , y24879 , y24880 , y24881 , y24882 , y24883 , y24884 , y24885 , y24886 , y24887 , y24888 , y24889 , y24890 , y24891 , y24892 , y24893 , y24894 , y24895 , y24896 , y24897 , y24898 , y24899 , y24900 , y24901 , y24902 , y24903 , y24904 , y24905 , y24906 , y24907 , y24908 , y24909 , y24910 , y24911 , y24912 , y24913 , y24914 , y24915 , y24916 , y24917 , y24918 , y24919 , y24920 , y24921 , y24922 , y24923 , y24924 , y24925 , y24926 , y24927 , y24928 , y24929 , y24930 , y24931 , y24932 , y24933 , y24934 , y24935 , y24936 , y24937 , y24938 , y24939 , y24940 , y24941 , y24942 , y24943 , y24944 , y24945 , y24946 , y24947 , y24948 , y24949 , y24950 , y24951 , y24952 , y24953 , y24954 , y24955 , y24956 , y24957 , y24958 , y24959 , y24960 , y24961 , y24962 , y24963 , y24964 , y24965 , y24966 , y24967 , y24968 , y24969 , y24970 , y24971 , y24972 , y24973 , y24974 , y24975 , y24976 , y24977 , y24978 , y24979 , y24980 , y24981 , y24982 , y24983 , y24984 , y24985 , y24986 , y24987 , y24988 , y24989 , y24990 , y24991 , y24992 , y24993 , y24994 , y24995 , y24996 , y24997 , y24998 , y24999 , y25000 , y25001 , y25002 , y25003 , y25004 , y25005 , y25006 , y25007 , y25008 , y25009 , y25010 , y25011 , y25012 , y25013 , y25014 , y25015 , y25016 , y25017 , y25018 , y25019 , y25020 , y25021 , y25022 , y25023 , y25024 , y25025 , y25026 , y25027 , y25028 , y25029 , y25030 , y25031 , y25032 , y25033 , y25034 , y25035 , y25036 , y25037 , y25038 , y25039 , y25040 , y25041 , y25042 , y25043 , y25044 , y25045 , y25046 , y25047 , y25048 , y25049 , y25050 , y25051 , y25052 , y25053 , y25054 , y25055 , y25056 , y25057 , y25058 , y25059 , y25060 , y25061 , y25062 , y25063 , y25064 , y25065 , y25066 , y25067 , y25068 , y25069 , y25070 , y25071 , y25072 , y25073 , y25074 , y25075 , y25076 , y25077 , y25078 , y25079 , y25080 , y25081 , y25082 , y25083 , y25084 , y25085 , y25086 , y25087 , y25088 , y25089 , y25090 , y25091 , y25092 , y25093 , y25094 , y25095 , y25096 , y25097 , y25098 , y25099 , y25100 , y25101 , y25102 , y25103 , y25104 , y25105 , y25106 , y25107 , y25108 , y25109 , y25110 , y25111 , y25112 , y25113 , y25114 , y25115 , y25116 , y25117 , y25118 , y25119 , y25120 , y25121 , y25122 , y25123 , y25124 , y25125 , y25126 , y25127 , y25128 , y25129 , y25130 , y25131 , y25132 , y25133 , y25134 , y25135 , y25136 , y25137 , y25138 , y25139 , y25140 , y25141 , y25142 , y25143 , y25144 , y25145 , y25146 , y25147 , y25148 , y25149 , y25150 , y25151 , y25152 , y25153 , y25154 , y25155 , y25156 , y25157 , y25158 , y25159 , y25160 , y25161 , y25162 , y25163 , y25164 , y25165 , y25166 , y25167 , y25168 , y25169 , y25170 , y25171 , y25172 , y25173 , y25174 , y25175 , y25176 , y25177 , y25178 , y25179 , y25180 , y25181 , y25182 , y25183 , y25184 , y25185 , y25186 , y25187 , y25188 , y25189 , y25190 , y25191 , y25192 , y25193 , y25194 , y25195 , y25196 , y25197 , y25198 , y25199 , y25200 , y25201 , y25202 , y25203 , y25204 , y25205 , y25206 , y25207 , y25208 , y25209 , y25210 , y25211 , y25212 , y25213 , y25214 , y25215 , y25216 , y25217 , y25218 , y25219 , y25220 , y25221 , y25222 , y25223 , y25224 , y25225 , y25226 , y25227 , y25228 , y25229 , y25230 , y25231 , y25232 , y25233 , y25234 , y25235 , y25236 , y25237 , y25238 , y25239 , y25240 , y25241 , y25242 , y25243 , y25244 , y25245 , y25246 , y25247 , y25248 , y25249 , y25250 , y25251 , y25252 , y25253 , y25254 , y25255 , y25256 , y25257 , y25258 , y25259 , y25260 , y25261 , y25262 , y25263 , y25264 , y25265 , y25266 , y25267 , y25268 , y25269 , y25270 , y25271 , y25272 , y25273 , y25274 , y25275 , y25276 , y25277 , y25278 , y25279 , y25280 , y25281 , y25282 , y25283 , y25284 , y25285 , y25286 , y25287 , y25288 , y25289 , y25290 , y25291 , y25292 , y25293 , y25294 , y25295 , y25296 , y25297 , y25298 , y25299 , y25300 , y25301 , y25302 , y25303 , y25304 , y25305 , y25306 , y25307 , y25308 , y25309 , y25310 , y25311 , y25312 , y25313 , y25314 , y25315 , y25316 , y25317 , y25318 , y25319 , y25320 , y25321 , y25322 , y25323 , y25324 , y25325 , y25326 , y25327 , y25328 , y25329 , y25330 , y25331 , y25332 , y25333 , y25334 , y25335 , y25336 , y25337 , y25338 , y25339 , y25340 , y25341 , y25342 , y25343 , y25344 , y25345 , y25346 , y25347 , y25348 , y25349 , y25350 , y25351 , y25352 , y25353 , y25354 , y25355 , y25356 , y25357 , y25358 , y25359 , y25360 , y25361 , y25362 , y25363 , y25364 , y25365 , y25366 , y25367 , y25368 , y25369 , y25370 , y25371 , y25372 , y25373 , y25374 , y25375 , y25376 , y25377 , y25378 , y25379 , y25380 , y25381 , y25382 , y25383 , y25384 , y25385 , y25386 , y25387 , y25388 , y25389 , y25390 , y25391 , y25392 , y25393 , y25394 , y25395 , y25396 , y25397 , y25398 , y25399 , y25400 , y25401 , y25402 , y25403 , y25404 , y25405 , y25406 , y25407 , y25408 , y25409 , y25410 , y25411 , y25412 , y25413 , y25414 , y25415 , y25416 , y25417 , y25418 , y25419 , y25420 , y25421 , y25422 , y25423 , y25424 , y25425 , y25426 , y25427 , y25428 , y25429 , y25430 , y25431 , y25432 , y25433 , y25434 , y25435 , y25436 , y25437 , y25438 , y25439 , y25440 , y25441 , y25442 , y25443 , y25444 , y25445 , y25446 , y25447 , y25448 , y25449 , y25450 , y25451 , y25452 , y25453 , y25454 , y25455 , y25456 , y25457 , y25458 , y25459 , y25460 , y25461 , y25462 , y25463 , y25464 , y25465 , y25466 , y25467 , y25468 , y25469 , y25470 , y25471 , y25472 , y25473 , y25474 , y25475 , y25476 , y25477 , y25478 , y25479 , y25480 , y25481 , y25482 , y25483 , y25484 , y25485 , y25486 , y25487 , y25488 , y25489 , y25490 , y25491 , y25492 , y25493 , y25494 , y25495 , y25496 , y25497 , y25498 , y25499 , y25500 , y25501 , y25502 , y25503 , y25504 , y25505 , y25506 , y25507 , y25508 , y25509 , y25510 , y25511 , y25512 , y25513 , y25514 , y25515 , y25516 , y25517 , y25518 , y25519 , y25520 , y25521 , y25522 , y25523 , y25524 , y25525 , y25526 , y25527 , y25528 , y25529 , y25530 , y25531 , y25532 , y25533 , y25534 , y25535 , y25536 , y25537 , y25538 , y25539 , y25540 , y25541 , y25542 , y25543 , y25544 , y25545 , y25546 , y25547 , y25548 , y25549 , y25550 , y25551 , y25552 , y25553 , y25554 , y25555 , y25556 , y25557 , y25558 , y25559 , y25560 , y25561 , y25562 , y25563 , y25564 , y25565 , y25566 , y25567 , y25568 , y25569 , y25570 , y25571 , y25572 , y25573 , y25574 , y25575 , y25576 , y25577 , y25578 , y25579 , y25580 , y25581 , y25582 , y25583 , y25584 , y25585 , y25586 , y25587 , y25588 , y25589 , y25590 , y25591 , y25592 , y25593 , y25594 , y25595 , y25596 , y25597 , y25598 , y25599 , y25600 , y25601 , y25602 , y25603 , y25604 , y25605 , y25606 , y25607 , y25608 , y25609 , y25610 , y25611 , y25612 , y25613 , y25614 , y25615 , y25616 , y25617 , y25618 , y25619 , y25620 , y25621 , y25622 , y25623 , y25624 , y25625 , y25626 , y25627 , y25628 , y25629 , y25630 , y25631 , y25632 , y25633 , y25634 , y25635 , y25636 , y25637 , y25638 , y25639 , y25640 , y25641 , y25642 , y25643 , y25644 , y25645 , y25646 , y25647 , y25648 , y25649 , y25650 , y25651 , y25652 , y25653 , y25654 , y25655 , y25656 , y25657 , y25658 , y25659 , y25660 , y25661 , y25662 , y25663 , y25664 , y25665 , y25666 , y25667 , y25668 , y25669 , y25670 , y25671 , y25672 , y25673 , y25674 , y25675 , y25676 , y25677 , y25678 , y25679 , y25680 , y25681 , y25682 , y25683 , y25684 , y25685 , y25686 , y25687 , y25688 , y25689 , y25690 , y25691 , y25692 , y25693 , y25694 , y25695 , y25696 , y25697 , y25698 , y25699 , y25700 , y25701 , y25702 , y25703 , y25704 , y25705 , y25706 , y25707 , y25708 , y25709 , y25710 , y25711 , y25712 , y25713 , y25714 , y25715 , y25716 , y25717 , y25718 , y25719 , y25720 , y25721 , y25722 , y25723 , y25724 , y25725 , y25726 , y25727 , y25728 , y25729 , y25730 , y25731 , y25732 , y25733 , y25734 , y25735 , y25736 , y25737 , y25738 , y25739 , y25740 , y25741 , y25742 , y25743 , y25744 , y25745 , y25746 , y25747 , y25748 , y25749 , y25750 , y25751 , y25752 , y25753 , y25754 , y25755 , y25756 , y25757 , y25758 , y25759 , y25760 , y25761 , y25762 , y25763 , y25764 , y25765 , y25766 , y25767 , y25768 , y25769 , y25770 , y25771 , y25772 , y25773 , y25774 , y25775 , y25776 , y25777 , y25778 , y25779 , y25780 , y25781 , y25782 , y25783 , y25784 , y25785 , y25786 , y25787 , y25788 , y25789 , y25790 , y25791 , y25792 , y25793 , y25794 , y25795 , y25796 , y25797 , y25798 , y25799 , y25800 , y25801 , y25802 , y25803 , y25804 , y25805 , y25806 , y25807 , y25808 , y25809 , y25810 , y25811 , y25812 , y25813 , y25814 , y25815 , y25816 , y25817 , y25818 , y25819 , y25820 , y25821 , y25822 , y25823 , y25824 , y25825 , y25826 , y25827 , y25828 , y25829 , y25830 , y25831 , y25832 , y25833 , y25834 , y25835 , y25836 , y25837 , y25838 , y25839 , y25840 , y25841 , y25842 , y25843 , y25844 , y25845 , y25846 , y25847 , y25848 , y25849 , y25850 , y25851 , y25852 , y25853 , y25854 , y25855 , y25856 , y25857 , y25858 , y25859 , y25860 , y25861 , y25862 , y25863 , y25864 , y25865 , y25866 , y25867 , y25868 , y25869 , y25870 , y25871 , y25872 , y25873 , y25874 , y25875 , y25876 , y25877 , y25878 , y25879 , y25880 , y25881 , y25882 , y25883 , y25884 , y25885 , y25886 , y25887 , y25888 , y25889 , y25890 , y25891 , y25892 , y25893 , y25894 , y25895 , y25896 , y25897 , y25898 , y25899 , y25900 , y25901 , y25902 , y25903 , y25904 , y25905 , y25906 , y25907 , y25908 , y25909 , y25910 , y25911 , y25912 , y25913 , y25914 , y25915 , y25916 , y25917 , y25918 , y25919 , y25920 , y25921 , y25922 , y25923 , y25924 , y25925 , y25926 , y25927 , y25928 , y25929 , y25930 , y25931 , y25932 , y25933 , y25934 , y25935 , y25936 , y25937 , y25938 , y25939 , y25940 , y25941 , y25942 , y25943 , y25944 , y25945 , y25946 , y25947 , y25948 , y25949 , y25950 , y25951 , y25952 , y25953 , y25954 , y25955 , y25956 , y25957 , y25958 , y25959 , y25960 , y25961 , y25962 , y25963 , y25964 , y25965 , y25966 , y25967 , y25968 , y25969 , y25970 , y25971 , y25972 , y25973 , y25974 , y25975 , y25976 , y25977 , y25978 , y25979 , y25980 , y25981 , y25982 , y25983 , y25984 , y25985 , y25986 , y25987 , y25988 , y25989 , y25990 , y25991 , y25992 , y25993 , y25994 , y25995 , y25996 , y25997 , y25998 , y25999 , y26000 , y26001 , y26002 , y26003 , y26004 , y26005 , y26006 , y26007 , y26008 , y26009 , y26010 , y26011 , y26012 , y26013 , y26014 , y26015 , y26016 , y26017 , y26018 , y26019 , y26020 , y26021 , y26022 , y26023 , y26024 , y26025 , y26026 , y26027 , y26028 , y26029 , y26030 , y26031 , y26032 , y26033 , y26034 , y26035 , y26036 , y26037 , y26038 , y26039 , y26040 , y26041 , y26042 , y26043 , y26044 , y26045 , y26046 , y26047 , y26048 , y26049 , y26050 , y26051 , y26052 , y26053 , y26054 , y26055 , y26056 , y26057 , y26058 , y26059 , y26060 , y26061 , y26062 , y26063 , y26064 , y26065 , y26066 , y26067 , y26068 , y26069 , y26070 , y26071 , y26072 , y26073 , y26074 , y26075 , y26076 , y26077 , y26078 , y26079 , y26080 , y26081 , y26082 , y26083 , y26084 , y26085 , y26086 , y26087 , y26088 , y26089 , y26090 , y26091 , y26092 , y26093 , y26094 , y26095 , y26096 , y26097 , y26098 , y26099 , y26100 , y26101 , y26102 , y26103 , y26104 , y26105 , y26106 , y26107 , y26108 , y26109 , y26110 , y26111 , y26112 , y26113 , y26114 , y26115 , y26116 , y26117 , y26118 , y26119 , y26120 , y26121 , y26122 , y26123 , y26124 , y26125 , y26126 , y26127 , y26128 , y26129 , y26130 , y26131 , y26132 , y26133 , y26134 , y26135 , y26136 , y26137 , y26138 , y26139 , y26140 , y26141 , y26142 , y26143 , y26144 , y26145 , y26146 , y26147 , y26148 , y26149 , y26150 , y26151 , y26152 , y26153 , y26154 , y26155 , y26156 , y26157 , y26158 , y26159 , y26160 , y26161 , y26162 , y26163 , y26164 , y26165 , y26166 , y26167 , y26168 , y26169 , y26170 , y26171 , y26172 , y26173 , y26174 , y26175 , y26176 , y26177 , y26178 , y26179 , y26180 , y26181 , y26182 , y26183 , y26184 , y26185 , y26186 , y26187 , y26188 , y26189 , y26190 , y26191 , y26192 , y26193 , y26194 , y26195 , y26196 , y26197 , y26198 , y26199 , y26200 , y26201 , y26202 , y26203 , y26204 , y26205 , y26206 , y26207 , y26208 , y26209 , y26210 , y26211 , y26212 , y26213 , y26214 , y26215 , y26216 , y26217 , y26218 , y26219 , y26220 , y26221 , y26222 , y26223 , y26224 , y26225 , y26226 , y26227 , y26228 , y26229 , y26230 , y26231 , y26232 , y26233 , y26234 , y26235 , y26236 , y26237 , y26238 , y26239 , y26240 , y26241 , y26242 , y26243 , y26244 , y26245 , y26246 , y26247 , y26248 , y26249 , y26250 , y26251 , y26252 , y26253 , y26254 , y26255 , y26256 , y26257 , y26258 , y26259 , y26260 , y26261 , y26262 , y26263 , y26264 , y26265 , y26266 , y26267 , y26268 , y26269 , y26270 , y26271 , y26272 , y26273 , y26274 , y26275 , y26276 , y26277 , y26278 , y26279 , y26280 , y26281 , y26282 , y26283 , y26284 , y26285 , y26286 , y26287 , y26288 , y26289 , y26290 , y26291 , y26292 , y26293 , y26294 , y26295 , y26296 , y26297 , y26298 , y26299 , y26300 , y26301 , y26302 , y26303 , y26304 , y26305 , y26306 , y26307 , y26308 , y26309 , y26310 , y26311 , y26312 , y26313 , y26314 , y26315 , y26316 , y26317 , y26318 , y26319 , y26320 , y26321 , y26322 , y26323 , y26324 , y26325 , y26326 , y26327 , y26328 , y26329 , y26330 , y26331 , y26332 , y26333 , y26334 , y26335 , y26336 , y26337 , y26338 , y26339 , y26340 , y26341 , y26342 , y26343 , y26344 , y26345 , y26346 , y26347 , y26348 , y26349 , y26350 , y26351 , y26352 , y26353 , y26354 , y26355 , y26356 , y26357 , y26358 , y26359 , y26360 , y26361 , y26362 , y26363 , y26364 , y26365 , y26366 , y26367 , y26368 , y26369 , y26370 , y26371 , y26372 , y26373 , y26374 , y26375 , y26376 , y26377 , y26378 , y26379 , y26380 , y26381 , y26382 , y26383 , y26384 , y26385 , y26386 , y26387 , y26388 , y26389 , y26390 , y26391 , y26392 , y26393 , y26394 , y26395 , y26396 , y26397 , y26398 , y26399 , y26400 , y26401 , y26402 , y26403 , y26404 , y26405 , y26406 , y26407 , y26408 , y26409 , y26410 , y26411 , y26412 , y26413 , y26414 , y26415 , y26416 , y26417 , y26418 , y26419 , y26420 , y26421 , y26422 , y26423 , y26424 , y26425 , y26426 , y26427 , y26428 , y26429 , y26430 , y26431 , y26432 , y26433 , y26434 , y26435 , y26436 , y26437 , y26438 , y26439 , y26440 , y26441 , y26442 , y26443 , y26444 , y26445 , y26446 , y26447 , y26448 , y26449 , y26450 , y26451 , y26452 , y26453 , y26454 , y26455 , y26456 , y26457 , y26458 , y26459 , y26460 , y26461 , y26462 , y26463 , y26464 , y26465 , y26466 , y26467 , y26468 , y26469 , y26470 , y26471 , y26472 , y26473 , y26474 , y26475 , y26476 , y26477 , y26478 , y26479 , y26480 , y26481 , y26482 , y26483 , y26484 , y26485 , y26486 , y26487 , y26488 , y26489 , y26490 , y26491 , y26492 , y26493 , y26494 , y26495 , y26496 , y26497 , y26498 , y26499 , y26500 , y26501 , y26502 , y26503 , y26504 , y26505 , y26506 , y26507 , y26508 , y26509 , y26510 , y26511 , y26512 , y26513 , y26514 , y26515 , y26516 , y26517 , y26518 , y26519 , y26520 , y26521 , y26522 , y26523 , y26524 , y26525 , y26526 , y26527 , y26528 , y26529 , y26530 , y26531 , y26532 , y26533 , y26534 , y26535 , y26536 , y26537 , y26538 , y26539 , y26540 , y26541 , y26542 , y26543 , y26544 , y26545 , y26546 , y26547 , y26548 , y26549 , y26550 , y26551 , y26552 , y26553 , y26554 , y26555 , y26556 , y26557 , y26558 , y26559 , y26560 , y26561 , y26562 , y26563 , y26564 , y26565 , y26566 , y26567 , y26568 , y26569 , y26570 , y26571 , y26572 , y26573 , y26574 , y26575 , y26576 , y26577 , y26578 , y26579 , y26580 , y26581 , y26582 , y26583 , y26584 , y26585 , y26586 , y26587 , y26588 , y26589 , y26590 , y26591 , y26592 , y26593 , y26594 , y26595 , y26596 , y26597 , y26598 , y26599 , y26600 , y26601 , y26602 , y26603 , y26604 , y26605 , y26606 , y26607 , y26608 , y26609 , y26610 , y26611 , y26612 , y26613 , y26614 , y26615 , y26616 , y26617 , y26618 , y26619 , y26620 , y26621 , y26622 , y26623 , y26624 , y26625 , y26626 , y26627 , y26628 , y26629 , y26630 , y26631 , y26632 , y26633 , y26634 , y26635 , y26636 , y26637 , y26638 , y26639 , y26640 , y26641 , y26642 , y26643 , y26644 , y26645 , y26646 , y26647 , y26648 , y26649 , y26650 , y26651 , y26652 , y26653 , y26654 , y26655 , y26656 , y26657 , y26658 , y26659 , y26660 , y26661 , y26662 , y26663 , y26664 , y26665 , y26666 , y26667 , y26668 , y26669 , y26670 , y26671 , y26672 , y26673 , y26674 , y26675 , y26676 , y26677 , y26678 , y26679 , y26680 , y26681 , y26682 , y26683 , y26684 , y26685 , y26686 , y26687 , y26688 , y26689 , y26690 , y26691 , y26692 , y26693 , y26694 , y26695 , y26696 , y26697 , y26698 , y26699 , y26700 , y26701 , y26702 , y26703 , y26704 , y26705 , y26706 , y26707 , y26708 , y26709 , y26710 , y26711 , y26712 , y26713 , y26714 , y26715 , y26716 , y26717 , y26718 , y26719 , y26720 , y26721 , y26722 , y26723 , y26724 , y26725 , y26726 , y26727 , y26728 , y26729 , y26730 , y26731 , y26732 , y26733 , y26734 , y26735 , y26736 , y26737 , y26738 , y26739 , y26740 , y26741 , y26742 , y26743 , y26744 , y26745 , y26746 , y26747 , y26748 , y26749 , y26750 , y26751 , y26752 , y26753 , y26754 , y26755 , y26756 , y26757 , y26758 , y26759 , y26760 , y26761 , y26762 , y26763 , y26764 , y26765 , y26766 , y26767 , y26768 , y26769 , y26770 , y26771 , y26772 , y26773 , y26774 , y26775 , y26776 , y26777 , y26778 , y26779 , y26780 , y26781 , y26782 , y26783 , y26784 , y26785 , y26786 , y26787 , y26788 , y26789 , y26790 , y26791 , y26792 , y26793 , y26794 , y26795 , y26796 , y26797 , y26798 , y26799 , y26800 , y26801 , y26802 , y26803 , y26804 , y26805 , y26806 , y26807 , y26808 , y26809 , y26810 , y26811 , y26812 , y26813 , y26814 , y26815 , y26816 , y26817 , y26818 , y26819 , y26820 , y26821 , y26822 , y26823 , y26824 , y26825 , y26826 , y26827 , y26828 , y26829 , y26830 , y26831 , y26832 , y26833 , y26834 , y26835 , y26836 , y26837 , y26838 , y26839 , y26840 , y26841 , y26842 , y26843 , y26844 , y26845 , y26846 , y26847 , y26848 , y26849 , y26850 , y26851 , y26852 , y26853 , y26854 , y26855 , y26856 , y26857 , y26858 , y26859 , y26860 , y26861 , y26862 , y26863 , y26864 , y26865 , y26866 , y26867 , y26868 , y26869 , y26870 , y26871 , y26872 , y26873 , y26874 , y26875 , y26876 , y26877 , y26878 , y26879 , y26880 , y26881 , y26882 , y26883 , y26884 , y26885 , y26886 , y26887 , y26888 , y26889 , y26890 , y26891 , y26892 , y26893 , y26894 , y26895 , y26896 , y26897 , y26898 , y26899 , y26900 , y26901 , y26902 , y26903 , y26904 , y26905 , y26906 , y26907 , y26908 , y26909 , y26910 , y26911 , y26912 , y26913 , y26914 , y26915 , y26916 , y26917 , y26918 , y26919 , y26920 , y26921 , y26922 , y26923 , y26924 , y26925 , y26926 , y26927 , y26928 , y26929 , y26930 , y26931 , y26932 , y26933 , y26934 , y26935 , y26936 , y26937 , y26938 , y26939 , y26940 , y26941 , y26942 , y26943 , y26944 , y26945 , y26946 , y26947 , y26948 , y26949 , y26950 , y26951 , y26952 , y26953 , y26954 , y26955 , y26956 , y26957 , y26958 , y26959 , y26960 , y26961 , y26962 , y26963 , y26964 , y26965 , y26966 , y26967 , y26968 , y26969 , y26970 , y26971 , y26972 , y26973 , y26974 , y26975 , y26976 , y26977 , y26978 , y26979 , y26980 , y26981 , y26982 , y26983 , y26984 , y26985 , y26986 , y26987 , y26988 , y26989 , y26990 , y26991 , y26992 , y26993 , y26994 , y26995 , y26996 , y26997 , y26998 , y26999 , y27000 , y27001 , y27002 , y27003 , y27004 , y27005 , y27006 , y27007 , y27008 , y27009 , y27010 , y27011 , y27012 , y27013 , y27014 , y27015 , y27016 , y27017 , y27018 , y27019 , y27020 , y27021 , y27022 , y27023 , y27024 , y27025 , y27026 , y27027 , y27028 , y27029 , y27030 , y27031 , y27032 , y27033 , y27034 , y27035 , y27036 , y27037 , y27038 , y27039 , y27040 , y27041 , y27042 , y27043 , y27044 , y27045 , y27046 , y27047 , y27048 , y27049 , y27050 , y27051 , y27052 , y27053 , y27054 , y27055 , y27056 , y27057 , y27058 , y27059 , y27060 , y27061 , y27062 , y27063 , y27064 , y27065 , y27066 , y27067 , y27068 , y27069 , y27070 , y27071 , y27072 , y27073 , y27074 , y27075 , y27076 , y27077 , y27078 , y27079 , y27080 , y27081 , y27082 , y27083 , y27084 , y27085 , y27086 , y27087 , y27088 , y27089 , y27090 , y27091 , y27092 , y27093 , y27094 , y27095 , y27096 , y27097 , y27098 , y27099 , y27100 , y27101 , y27102 , y27103 , y27104 , y27105 , y27106 , y27107 , y27108 , y27109 , y27110 , y27111 , y27112 , y27113 , y27114 , y27115 , y27116 , y27117 , y27118 , y27119 , y27120 , y27121 , y27122 , y27123 , y27124 , y27125 , y27126 , y27127 , y27128 , y27129 , y27130 , y27131 , y27132 , y27133 , y27134 , y27135 , y27136 , y27137 , y27138 , y27139 , y27140 , y27141 , y27142 , y27143 , y27144 , y27145 , y27146 , y27147 , y27148 , y27149 , y27150 , y27151 , y27152 , y27153 , y27154 , y27155 , y27156 , y27157 , y27158 , y27159 , y27160 , y27161 , y27162 , y27163 , y27164 , y27165 , y27166 , y27167 , y27168 , y27169 , y27170 , y27171 , y27172 , y27173 , y27174 , y27175 , y27176 , y27177 , y27178 , y27179 , y27180 , y27181 , y27182 , y27183 , y27184 , y27185 , y27186 , y27187 , y27188 , y27189 , y27190 , y27191 , y27192 , y27193 , y27194 , y27195 , y27196 , y27197 , y27198 , y27199 , y27200 , y27201 , y27202 , y27203 , y27204 , y27205 , y27206 , y27207 , y27208 , y27209 , y27210 , y27211 , y27212 , y27213 , y27214 , y27215 , y27216 , y27217 , y27218 , y27219 , y27220 , y27221 , y27222 , y27223 , y27224 , y27225 , y27226 , y27227 , y27228 , y27229 , y27230 , y27231 , y27232 , y27233 , y27234 , y27235 , y27236 , y27237 , y27238 , y27239 , y27240 , y27241 , y27242 , y27243 , y27244 , y27245 , y27246 , y27247 , y27248 , y27249 , y27250 , y27251 , y27252 , y27253 , y27254 , y27255 , y27256 , y27257 , y27258 , y27259 , y27260 , y27261 , y27262 , y27263 , y27264 , y27265 , y27266 , y27267 , y27268 , y27269 , y27270 , y27271 , y27272 , y27273 , y27274 , y27275 , y27276 , y27277 , y27278 , y27279 , y27280 , y27281 , y27282 , y27283 , y27284 , y27285 , y27286 , y27287 , y27288 , y27289 , y27290 , y27291 , y27292 , y27293 , y27294 , y27295 , y27296 , y27297 , y27298 , y27299 , y27300 , y27301 , y27302 , y27303 , y27304 , y27305 , y27306 , y27307 , y27308 , y27309 , y27310 , y27311 , y27312 , y27313 , y27314 , y27315 , y27316 , y27317 , y27318 , y27319 , y27320 , y27321 , y27322 , y27323 , y27324 , y27325 , y27326 , y27327 , y27328 , y27329 , y27330 , y27331 , y27332 , y27333 , y27334 , y27335 , y27336 , y27337 , y27338 , y27339 , y27340 , y27341 , y27342 , y27343 , y27344 , y27345 , y27346 , y27347 , y27348 , y27349 , y27350 , y27351 , y27352 , y27353 , y27354 , y27355 , y27356 , y27357 , y27358 , y27359 , y27360 , y27361 , y27362 , y27363 , y27364 , y27365 , y27366 , y27367 , y27368 , y27369 , y27370 , y27371 , y27372 , y27373 , y27374 , y27375 , y27376 , y27377 , y27378 , y27379 , y27380 , y27381 , y27382 , y27383 , y27384 , y27385 , y27386 , y27387 , y27388 , y27389 , y27390 , y27391 , y27392 , y27393 , y27394 , y27395 , y27396 , y27397 , y27398 , y27399 , y27400 , y27401 , y27402 , y27403 , y27404 , y27405 , y27406 , y27407 , y27408 , y27409 , y27410 , y27411 , y27412 , y27413 , y27414 , y27415 , y27416 , y27417 , y27418 , y27419 , y27420 , y27421 , y27422 , y27423 , y27424 , y27425 , y27426 , y27427 , y27428 , y27429 , y27430 , y27431 , y27432 , y27433 , y27434 , y27435 , y27436 , y27437 , y27438 , y27439 , y27440 , y27441 , y27442 , y27443 , y27444 , y27445 , y27446 , y27447 , y27448 , y27449 , y27450 , y27451 , y27452 , y27453 , y27454 , y27455 , y27456 , y27457 , y27458 , y27459 , y27460 , y27461 , y27462 , y27463 , y27464 , y27465 , y27466 , y27467 , y27468 , y27469 , y27470 , y27471 , y27472 , y27473 , y27474 , y27475 , y27476 , y27477 , y27478 , y27479 , y27480 , y27481 , y27482 , y27483 , y27484 , y27485 , y27486 , y27487 , y27488 , y27489 , y27490 , y27491 , y27492 , y27493 , y27494 , y27495 , y27496 , y27497 , y27498 , y27499 , y27500 , y27501 , y27502 , y27503 , y27504 , y27505 , y27506 , y27507 , y27508 , y27509 , y27510 , y27511 , y27512 , y27513 , y27514 , y27515 , y27516 , y27517 , y27518 , y27519 , y27520 , y27521 , y27522 , y27523 , y27524 , y27525 , y27526 , y27527 , y27528 , y27529 , y27530 , y27531 , y27532 , y27533 , y27534 , y27535 , y27536 , y27537 , y27538 , y27539 , y27540 , y27541 , y27542 , y27543 , y27544 , y27545 , y27546 , y27547 , y27548 , y27549 , y27550 , y27551 , y27552 , y27553 , y27554 , y27555 , y27556 , y27557 , y27558 , y27559 , y27560 , y27561 , y27562 , y27563 , y27564 , y27565 , y27566 , y27567 , y27568 , y27569 , y27570 , y27571 , y27572 , y27573 , y27574 , y27575 , y27576 , y27577 , y27578 , y27579 , y27580 , y27581 , y27582 , y27583 , y27584 , y27585 , y27586 , y27587 , y27588 , y27589 , y27590 , y27591 , y27592 , y27593 , y27594 , y27595 , y27596 , y27597 , y27598 , y27599 , y27600 , y27601 , y27602 , y27603 , y27604 , y27605 , y27606 , y27607 , y27608 , y27609 , y27610 , y27611 , y27612 , y27613 , y27614 , y27615 , y27616 , y27617 , y27618 , y27619 , y27620 , y27621 , y27622 , y27623 , y27624 , y27625 , y27626 , y27627 , y27628 , y27629 , y27630 , y27631 , y27632 , y27633 , y27634 , y27635 , y27636 , y27637 , y27638 , y27639 , y27640 , y27641 , y27642 , y27643 , y27644 , y27645 , y27646 , y27647 , y27648 , y27649 , y27650 , y27651 , y27652 , y27653 , y27654 , y27655 , y27656 , y27657 , y27658 , y27659 , y27660 , y27661 , y27662 , y27663 , y27664 , y27665 , y27666 , y27667 , y27668 , y27669 , y27670 , y27671 , y27672 , y27673 , y27674 , y27675 , y27676 , y27677 , y27678 , y27679 , y27680 , y27681 , y27682 , y27683 , y27684 , y27685 , y27686 , y27687 , y27688 , y27689 , y27690 , y27691 , y27692 , y27693 , y27694 , y27695 , y27696 , y27697 , y27698 , y27699 , y27700 , y27701 , y27702 , y27703 , y27704 , y27705 , y27706 , y27707 , y27708 , y27709 , y27710 , y27711 , y27712 , y27713 , y27714 , y27715 , y27716 , y27717 , y27718 , y27719 , y27720 , y27721 , y27722 , y27723 , y27724 , y27725 , y27726 , y27727 , y27728 , y27729 , y27730 , y27731 , y27732 , y27733 , y27734 , y27735 , y27736 , y27737 , y27738 , y27739 , y27740 , y27741 , y27742 , y27743 , y27744 , y27745 , y27746 , y27747 , y27748 , y27749 , y27750 , y27751 , y27752 , y27753 , y27754 , y27755 , y27756 , y27757 , y27758 , y27759 , y27760 , y27761 , y27762 , y27763 , y27764 , y27765 , y27766 , y27767 , y27768 , y27769 , y27770 , y27771 , y27772 , y27773 , y27774 , y27775 , y27776 , y27777 , y27778 , y27779 , y27780 , y27781 , y27782 , y27783 , y27784 , y27785 , y27786 , y27787 , y27788 , y27789 , y27790 , y27791 , y27792 , y27793 , y27794 , y27795 , y27796 , y27797 , y27798 , y27799 , y27800 , y27801 , y27802 , y27803 , y27804 , y27805 , y27806 , y27807 , y27808 , y27809 , y27810 , y27811 , y27812 , y27813 , y27814 , y27815 , y27816 , y27817 , y27818 , y27819 , y27820 , y27821 , y27822 , y27823 , y27824 , y27825 , y27826 , y27827 , y27828 , y27829 , y27830 , y27831 , y27832 , y27833 , y27834 , y27835 , y27836 , y27837 , y27838 , y27839 , y27840 , y27841 , y27842 , y27843 , y27844 , y27845 , y27846 , y27847 , y27848 , y27849 , y27850 , y27851 , y27852 , y27853 , y27854 , y27855 , y27856 , y27857 , y27858 , y27859 , y27860 , y27861 , y27862 , y27863 , y27864 , y27865 , y27866 , y27867 , y27868 , y27869 , y27870 , y27871 , y27872 , y27873 , y27874 , y27875 , y27876 , y27877 , y27878 , y27879 , y27880 , y27881 , y27882 , y27883 , y27884 , y27885 , y27886 , y27887 , y27888 , y27889 , y27890 , y27891 , y27892 , y27893 , y27894 , y27895 , y27896 , y27897 , y27898 , y27899 , y27900 , y27901 , y27902 , y27903 , y27904 , y27905 , y27906 , y27907 , y27908 , y27909 , y27910 , y27911 , y27912 , y27913 , y27914 , y27915 , y27916 , y27917 , y27918 , y27919 , y27920 , y27921 , y27922 , y27923 , y27924 , y27925 , y27926 , y27927 , y27928 , y27929 , y27930 , y27931 , y27932 , y27933 , y27934 , y27935 , y27936 , y27937 , y27938 , y27939 , y27940 , y27941 , y27942 , y27943 , y27944 , y27945 , y27946 , y27947 , y27948 , y27949 , y27950 , y27951 , y27952 , y27953 , y27954 , y27955 , y27956 , y27957 , y27958 , y27959 , y27960 , y27961 , y27962 , y27963 , y27964 , y27965 , y27966 , y27967 , y27968 , y27969 , y27970 , y27971 , y27972 , y27973 , y27974 , y27975 , y27976 , y27977 , y27978 , y27979 , y27980 , y27981 , y27982 , y27983 , y27984 , y27985 , y27986 , y27987 , y27988 , y27989 , y27990 , y27991 , y27992 , y27993 , y27994 , y27995 , y27996 , y27997 , y27998 , y27999 , y28000 , y28001 , y28002 , y28003 , y28004 , y28005 , y28006 , y28007 , y28008 , y28009 , y28010 , y28011 , y28012 , y28013 , y28014 , y28015 , y28016 , y28017 , y28018 , y28019 , y28020 , y28021 , y28022 , y28023 , y28024 , y28025 , y28026 , y28027 , y28028 , y28029 , y28030 , y28031 , y28032 , y28033 , y28034 , y28035 , y28036 , y28037 , y28038 , y28039 , y28040 , y28041 , y28042 , y28043 , y28044 , y28045 , y28046 , y28047 , y28048 , y28049 , y28050 , y28051 , y28052 , y28053 , y28054 , y28055 , y28056 , y28057 , y28058 , y28059 , y28060 , y28061 , y28062 , y28063 , y28064 , y28065 , y28066 , y28067 , y28068 , y28069 , y28070 , y28071 , y28072 , y28073 , y28074 , y28075 , y28076 , y28077 , y28078 , y28079 , y28080 , y28081 , y28082 , y28083 , y28084 , y28085 , y28086 , y28087 , y28088 , y28089 , y28090 , y28091 , y28092 , y28093 , y28094 , y28095 , y28096 , y28097 , y28098 , y28099 , y28100 , y28101 , y28102 , y28103 , y28104 , y28105 , y28106 , y28107 , y28108 , y28109 , y28110 , y28111 , y28112 , y28113 , y28114 , y28115 , y28116 , y28117 , y28118 , y28119 , y28120 , y28121 , y28122 , y28123 , y28124 , y28125 , y28126 , y28127 , y28128 , y28129 , y28130 , y28131 , y28132 , y28133 , y28134 , y28135 , y28136 , y28137 , y28138 , y28139 , y28140 , y28141 , y28142 , y28143 , y28144 , y28145 , y28146 , y28147 , y28148 , y28149 , y28150 , y28151 , y28152 , y28153 , y28154 , y28155 , y28156 , y28157 , y28158 , y28159 , y28160 , y28161 , y28162 , y28163 , y28164 , y28165 , y28166 , y28167 , y28168 , y28169 , y28170 , y28171 , y28172 , y28173 , y28174 , y28175 , y28176 , y28177 , y28178 , y28179 , y28180 , y28181 , y28182 , y28183 , y28184 , y28185 , y28186 , y28187 , y28188 , y28189 , y28190 , y28191 , y28192 , y28193 , y28194 , y28195 , y28196 , y28197 , y28198 , y28199 , y28200 , y28201 , y28202 , y28203 , y28204 , y28205 , y28206 , y28207 , y28208 , y28209 , y28210 , y28211 , y28212 , y28213 , y28214 , y28215 , y28216 , y28217 , y28218 , y28219 , y28220 , y28221 , y28222 , y28223 , y28224 , y28225 , y28226 , y28227 , y28228 , y28229 , y28230 , y28231 , y28232 , y28233 , y28234 , y28235 , y28236 , y28237 , y28238 , y28239 , y28240 , y28241 , y28242 , y28243 , y28244 , y28245 , y28246 , y28247 , y28248 , y28249 , y28250 , y28251 , y28252 , y28253 , y28254 , y28255 , y28256 , y28257 , y28258 , y28259 , y28260 , y28261 , y28262 , y28263 , y28264 , y28265 , y28266 , y28267 , y28268 , y28269 , y28270 , y28271 , y28272 , y28273 , y28274 , y28275 , y28276 , y28277 , y28278 , y28279 , y28280 , y28281 , y28282 , y28283 , y28284 , y28285 , y28286 , y28287 , y28288 , y28289 , y28290 , y28291 , y28292 , y28293 , y28294 , y28295 , y28296 , y28297 , y28298 , y28299 , y28300 , y28301 , y28302 , y28303 , y28304 , y28305 , y28306 , y28307 , y28308 , y28309 , y28310 , y28311 , y28312 , y28313 , y28314 , y28315 , y28316 , y28317 , y28318 , y28319 , y28320 , y28321 , y28322 , y28323 , y28324 , y28325 , y28326 , y28327 , y28328 , y28329 , y28330 , y28331 , y28332 , y28333 , y28334 , y28335 , y28336 , y28337 , y28338 , y28339 , y28340 , y28341 , y28342 , y28343 , y28344 , y28345 , y28346 , y28347 , y28348 , y28349 , y28350 , y28351 , y28352 , y28353 , y28354 , y28355 , y28356 , y28357 , y28358 , y28359 , y28360 , y28361 , y28362 , y28363 , y28364 , y28365 , y28366 , y28367 , y28368 , y28369 , y28370 , y28371 , y28372 , y28373 , y28374 , y28375 , y28376 , y28377 , y28378 , y28379 , y28380 , y28381 , y28382 , y28383 , y28384 , y28385 , y28386 , y28387 , y28388 , y28389 , y28390 , y28391 , y28392 , y28393 , y28394 , y28395 , y28396 , y28397 , y28398 , y28399 , y28400 , y28401 , y28402 , y28403 , y28404 , y28405 , y28406 , y28407 , y28408 , y28409 , y28410 , y28411 , y28412 , y28413 , y28414 , y28415 , y28416 , y28417 , y28418 , y28419 , y28420 , y28421 , y28422 , y28423 , y28424 , y28425 , y28426 , y28427 , y28428 , y28429 , y28430 , y28431 , y28432 , y28433 , y28434 , y28435 , y28436 , y28437 , y28438 , y28439 , y28440 , y28441 , y28442 , y28443 , y28444 , y28445 , y28446 , y28447 , y28448 , y28449 , y28450 , y28451 , y28452 , y28453 , y28454 , y28455 , y28456 , y28457 , y28458 , y28459 , y28460 , y28461 , y28462 , y28463 , y28464 , y28465 , y28466 , y28467 , y28468 , y28469 , y28470 , y28471 , y28472 , y28473 , y28474 , y28475 , y28476 , y28477 , y28478 , y28479 , y28480 , y28481 , y28482 , y28483 , y28484 , y28485 , y28486 , y28487 , y28488 , y28489 , y28490 , y28491 , y28492 , y28493 , y28494 , y28495 , y28496 , y28497 , y28498 , y28499 , y28500 , y28501 , y28502 , y28503 , y28504 , y28505 , y28506 , y28507 , y28508 , y28509 , y28510 , y28511 , y28512 , y28513 , y28514 , y28515 , y28516 , y28517 , y28518 , y28519 , y28520 , y28521 , y28522 , y28523 , y28524 , y28525 , y28526 , y28527 , y28528 , y28529 , y28530 , y28531 , y28532 , y28533 , y28534 , y28535 , y28536 , y28537 , y28538 , y28539 , y28540 , y28541 , y28542 , y28543 , y28544 , y28545 , y28546 , y28547 , y28548 , y28549 , y28550 , y28551 , y28552 , y28553 , y28554 , y28555 , y28556 , y28557 , y28558 , y28559 , y28560 , y28561 , y28562 , y28563 , y28564 , y28565 , y28566 , y28567 , y28568 , y28569 , y28570 , y28571 , y28572 , y28573 , y28574 , y28575 , y28576 , y28577 , y28578 , y28579 , y28580 , y28581 , y28582 , y28583 , y28584 , y28585 , y28586 , y28587 , y28588 , y28589 , y28590 , y28591 , y28592 , y28593 , y28594 , y28595 , y28596 , y28597 , y28598 , y28599 , y28600 , y28601 , y28602 , y28603 , y28604 , y28605 , y28606 , y28607 , y28608 , y28609 , y28610 , y28611 , y28612 , y28613 , y28614 , y28615 , y28616 , y28617 , y28618 , y28619 , y28620 , y28621 , y28622 , y28623 , y28624 , y28625 , y28626 , y28627 , y28628 , y28629 , y28630 , y28631 , y28632 , y28633 , y28634 , y28635 , y28636 , y28637 , y28638 , y28639 , y28640 , y28641 , y28642 , y28643 , y28644 , y28645 , y28646 , y28647 , y28648 , y28649 , y28650 , y28651 , y28652 , y28653 , y28654 , y28655 , y28656 , y28657 , y28658 , y28659 , y28660 , y28661 , y28662 , y28663 , y28664 , y28665 , y28666 , y28667 , y28668 , y28669 , y28670 , y28671 , y28672 , y28673 , y28674 , y28675 , y28676 , y28677 , y28678 , y28679 , y28680 , y28681 , y28682 , y28683 , y28684 , y28685 , y28686 , y28687 , y28688 , y28689 , y28690 , y28691 , y28692 , y28693 , y28694 , y28695 , y28696 , y28697 , y28698 , y28699 , y28700 , y28701 , y28702 , y28703 , y28704 , y28705 , y28706 , y28707 , y28708 , y28709 , y28710 , y28711 , y28712 , y28713 , y28714 , y28715 , y28716 , y28717 , y28718 , y28719 , y28720 , y28721 , y28722 , y28723 , y28724 , y28725 , y28726 , y28727 , y28728 , y28729 , y28730 , y28731 , y28732 , y28733 , y28734 , y28735 , y28736 , y28737 , y28738 , y28739 , y28740 , y28741 , y28742 , y28743 , y28744 , y28745 , y28746 , y28747 , y28748 , y28749 , y28750 , y28751 , y28752 , y28753 , y28754 , y28755 , y28756 , y28757 , y28758 , y28759 , y28760 , y28761 , y28762 , y28763 , y28764 , y28765 , y28766 , y28767 , y28768 , y28769 , y28770 , y28771 , y28772 , y28773 , y28774 , y28775 , y28776 , y28777 , y28778 , y28779 , y28780 , y28781 , y28782 , y28783 , y28784 , y28785 , y28786 , y28787 , y28788 , y28789 , y28790 , y28791 , y28792 , y28793 , y28794 , y28795 , y28796 , y28797 , y28798 , y28799 , y28800 , y28801 , y28802 , y28803 , y28804 , y28805 , y28806 , y28807 , y28808 , y28809 , y28810 , y28811 , y28812 , y28813 , y28814 , y28815 , y28816 , y28817 , y28818 , y28819 , y28820 , y28821 , y28822 , y28823 , y28824 , y28825 , y28826 , y28827 , y28828 , y28829 , y28830 , y28831 , y28832 , y28833 , y28834 , y28835 , y28836 , y28837 , y28838 , y28839 , y28840 , y28841 , y28842 , y28843 , y28844 , y28845 , y28846 , y28847 , y28848 , y28849 , y28850 , y28851 , y28852 , y28853 , y28854 , y28855 , y28856 , y28857 , y28858 , y28859 , y28860 , y28861 , y28862 , y28863 , y28864 , y28865 , y28866 , y28867 , y28868 , y28869 , y28870 , y28871 , y28872 , y28873 , y28874 , y28875 , y28876 , y28877 , y28878 , y28879 , y28880 , y28881 , y28882 , y28883 , y28884 , y28885 , y28886 , y28887 , y28888 , y28889 , y28890 , y28891 , y28892 , y28893 , y28894 , y28895 , y28896 , y28897 , y28898 , y28899 , y28900 , y28901 , y28902 , y28903 , y28904 , y28905 , y28906 , y28907 , y28908 , y28909 , y28910 , y28911 , y28912 , y28913 , y28914 , y28915 , y28916 , y28917 , y28918 , y28919 , y28920 , y28921 , y28922 , y28923 , y28924 , y28925 , y28926 , y28927 , y28928 , y28929 , y28930 , y28931 , y28932 , y28933 , y28934 , y28935 , y28936 , y28937 , y28938 , y28939 , y28940 , y28941 , y28942 , y28943 , y28944 , y28945 , y28946 , y28947 , y28948 , y28949 , y28950 , y28951 , y28952 , y28953 , y28954 , y28955 , y28956 , y28957 , y28958 , y28959 , y28960 , y28961 , y28962 , y28963 , y28964 , y28965 , y28966 , y28967 , y28968 , y28969 , y28970 , y28971 , y28972 , y28973 , y28974 , y28975 , y28976 , y28977 , y28978 , y28979 , y28980 , y28981 , y28982 , y28983 , y28984 , y28985 , y28986 , y28987 , y28988 , y28989 , y28990 , y28991 , y28992 , y28993 , y28994 , y28995 , y28996 , y28997 , y28998 , y28999 , y29000 , y29001 , y29002 , y29003 , y29004 , y29005 , y29006 , y29007 , y29008 , y29009 , y29010 , y29011 , y29012 , y29013 , y29014 , y29015 , y29016 , y29017 , y29018 , y29019 , y29020 , y29021 , y29022 , y29023 , y29024 , y29025 , y29026 , y29027 , y29028 , y29029 , y29030 , y29031 , y29032 , y29033 , y29034 , y29035 , y29036 , y29037 , y29038 , y29039 , y29040 , y29041 , y29042 , y29043 , y29044 , y29045 , y29046 , y29047 , y29048 , y29049 , y29050 , y29051 , y29052 , y29053 , y29054 , y29055 , y29056 , y29057 , y29058 , y29059 , y29060 , y29061 , y29062 , y29063 , y29064 , y29065 , y29066 , y29067 , y29068 , y29069 , y29070 , y29071 , y29072 , y29073 , y29074 , y29075 , y29076 , y29077 , y29078 , y29079 , y29080 , y29081 , y29082 , y29083 , y29084 , y29085 , y29086 , y29087 , y29088 , y29089 , y29090 , y29091 , y29092 , y29093 , y29094 , y29095 , y29096 , y29097 , y29098 , y29099 , y29100 , y29101 , y29102 , y29103 , y29104 , y29105 , y29106 , y29107 , y29108 , y29109 , y29110 , y29111 , y29112 , y29113 , y29114 , y29115 , y29116 , y29117 , y29118 , y29119 , y29120 , y29121 , y29122 , y29123 , y29124 , y29125 , y29126 , y29127 , y29128 , y29129 , y29130 , y29131 , y29132 , y29133 , y29134 , y29135 , y29136 , y29137 , y29138 , y29139 , y29140 , y29141 , y29142 , y29143 , y29144 , y29145 , y29146 , y29147 , y29148 , y29149 , y29150 , y29151 , y29152 , y29153 , y29154 , y29155 , y29156 , y29157 , y29158 , y29159 , y29160 , y29161 , y29162 , y29163 , y29164 , y29165 , y29166 , y29167 , y29168 , y29169 , y29170 , y29171 , y29172 , y29173 , y29174 , y29175 , y29176 , y29177 , y29178 , y29179 , y29180 , y29181 , y29182 , y29183 , y29184 , y29185 , y29186 , y29187 , y29188 , y29189 , y29190 , y29191 , y29192 , y29193 , y29194 , y29195 , y29196 , y29197 , y29198 , y29199 , y29200 , y29201 , y29202 , y29203 , y29204 , y29205 , y29206 , y29207 , y29208 , y29209 , y29210 , y29211 , y29212 , y29213 , y29214 , y29215 , y29216 , y29217 , y29218 , y29219 , y29220 , y29221 , y29222 , y29223 , y29224 , y29225 , y29226 , y29227 , y29228 , y29229 , y29230 , y29231 , y29232 , y29233 , y29234 , y29235 , y29236 , y29237 , y29238 , y29239 , y29240 , y29241 , y29242 , y29243 , y29244 , y29245 , y29246 , y29247 , y29248 , y29249 , y29250 , y29251 , y29252 , y29253 , y29254 , y29255 , y29256 , y29257 , y29258 , y29259 , y29260 , y29261 , y29262 , y29263 , y29264 , y29265 , y29266 , y29267 , y29268 , y29269 , y29270 , y29271 , y29272 , y29273 , y29274 , y29275 , y29276 , y29277 , y29278 , y29279 , y29280 , y29281 , y29282 , y29283 , y29284 , y29285 , y29286 , y29287 , y29288 , y29289 , y29290 , y29291 , y29292 , y29293 , y29294 , y29295 , y29296 , y29297 , y29298 , y29299 , y29300 , y29301 , y29302 , y29303 , y29304 , y29305 , y29306 , y29307 , y29308 , y29309 , y29310 , y29311 , y29312 , y29313 , y29314 , y29315 , y29316 , y29317 , y29318 , y29319 , y29320 , y29321 , y29322 , y29323 , y29324 , y29325 , y29326 , y29327 , y29328 , y29329 , y29330 , y29331 , y29332 , y29333 , y29334 , y29335 , y29336 , y29337 , y29338 , y29339 , y29340 , y29341 , y29342 , y29343 , y29344 , y29345 , y29346 , y29347 , y29348 , y29349 , y29350 , y29351 , y29352 , y29353 , y29354 , y29355 , y29356 , y29357 , y29358 , y29359 , y29360 , y29361 , y29362 , y29363 , y29364 , y29365 , y29366 , y29367 , y29368 , y29369 , y29370 , y29371 , y29372 , y29373 , y29374 , y29375 , y29376 , y29377 , y29378 , y29379 , y29380 , y29381 , y29382 , y29383 , y29384 , y29385 , y29386 , y29387 , y29388 , y29389 , y29390 , y29391 , y29392 , y29393 , y29394 , y29395 , y29396 , y29397 , y29398 , y29399 , y29400 , y29401 , y29402 , y29403 , y29404 , y29405 , y29406 , y29407 , y29408 , y29409 , y29410 , y29411 , y29412 , y29413 , y29414 , y29415 , y29416 , y29417 , y29418 , y29419 , y29420 , y29421 , y29422 , y29423 , y29424 , y29425 , y29426 , y29427 , y29428 , y29429 , y29430 , y29431 , y29432 , y29433 , y29434 , y29435 , y29436 , y29437 , y29438 , y29439 , y29440 , y29441 , y29442 , y29443 , y29444 , y29445 , y29446 , y29447 , y29448 , y29449 , y29450 , y29451 , y29452 , y29453 , y29454 , y29455 , y29456 , y29457 , y29458 , y29459 , y29460 , y29461 , y29462 , y29463 , y29464 , y29465 , y29466 , y29467 , y29468 , y29469 , y29470 , y29471 , y29472 , y29473 , y29474 , y29475 , y29476 , y29477 , y29478 , y29479 , y29480 , y29481 , y29482 , y29483 , y29484 , y29485 , y29486 , y29487 , y29488 , y29489 , y29490 , y29491 , y29492 , y29493 , y29494 , y29495 , y29496 , y29497 , y29498 , y29499 , y29500 , y29501 , y29502 , y29503 , y29504 , y29505 , y29506 , y29507 , y29508 , y29509 , y29510 , y29511 , y29512 , y29513 , y29514 , y29515 , y29516 , y29517 , y29518 , y29519 , y29520 , y29521 , y29522 , y29523 , y29524 , y29525 , y29526 , y29527 , y29528 , y29529 , y29530 , y29531 , y29532 , y29533 , y29534 , y29535 , y29536 , y29537 , y29538 , y29539 , y29540 , y29541 , y29542 , y29543 , y29544 , y29545 , y29546 , y29547 , y29548 , y29549 , y29550 , y29551 , y29552 , y29553 , y29554 , y29555 , y29556 , y29557 , y29558 , y29559 , y29560 , y29561 , y29562 , y29563 , y29564 , y29565 , y29566 , y29567 , y29568 , y29569 , y29570 , y29571 , y29572 , y29573 , y29574 , y29575 , y29576 , y29577 , y29578 , y29579 , y29580 , y29581 , y29582 , y29583 , y29584 , y29585 , y29586 , y29587 , y29588 , y29589 , y29590 , y29591 , y29592 , y29593 , y29594 , y29595 , y29596 , y29597 , y29598 , y29599 , y29600 , y29601 , y29602 , y29603 , y29604 , y29605 , y29606 , y29607 , y29608 , y29609 , y29610 , y29611 , y29612 , y29613 , y29614 , y29615 , y29616 , y29617 , y29618 , y29619 , y29620 , y29621 , y29622 , y29623 , y29624 , y29625 , y29626 , y29627 , y29628 , y29629 , y29630 , y29631 , y29632 , y29633 , y29634 , y29635 , y29636 , y29637 , y29638 , y29639 , y29640 , y29641 , y29642 , y29643 , y29644 , y29645 , y29646 , y29647 , y29648 , y29649 , y29650 , y29651 , y29652 , y29653 , y29654 , y29655 , y29656 , y29657 , y29658 , y29659 , y29660 , y29661 , y29662 , y29663 , y29664 , y29665 , y29666 , y29667 , y29668 , y29669 , y29670 , y29671 , y29672 , y29673 , y29674 , y29675 , y29676 , y29677 , y29678 , y29679 , y29680 , y29681 , y29682 , y29683 , y29684 , y29685 , y29686 , y29687 , y29688 , y29689 , y29690 , y29691 , y29692 , y29693 , y29694 , y29695 , y29696 , y29697 , y29698 , y29699 , y29700 , y29701 , y29702 , y29703 , y29704 , y29705 , y29706 , y29707 , y29708 , y29709 , y29710 , y29711 , y29712 , y29713 , y29714 , y29715 , y29716 , y29717 , y29718 , y29719 , y29720 , y29721 , y29722 , y29723 , y29724 , y29725 , y29726 , y29727 , y29728 , y29729 , y29730 , y29731 , y29732 , y29733 , y29734 , y29735 , y29736 , y29737 , y29738 , y29739 , y29740 , y29741 , y29742 , y29743 , y29744 , y29745 , y29746 , y29747 , y29748 , y29749 , y29750 , y29751 , y29752 , y29753 , y29754 , y29755 , y29756 , y29757 , y29758 , y29759 , y29760 , y29761 , y29762 , y29763 , y29764 , y29765 , y29766 , y29767 , y29768 , y29769 , y29770 , y29771 , y29772 , y29773 , y29774 , y29775 , y29776 , y29777 , y29778 , y29779 , y29780 , y29781 , y29782 , y29783 , y29784 , y29785 , y29786 , y29787 , y29788 , y29789 , y29790 , y29791 , y29792 , y29793 , y29794 , y29795 , y29796 , y29797 , y29798 , y29799 , y29800 , y29801 , y29802 , y29803 , y29804 , y29805 , y29806 , y29807 , y29808 , y29809 , y29810 , y29811 , y29812 , y29813 , y29814 , y29815 , y29816 , y29817 , y29818 , y29819 , y29820 , y29821 , y29822 , y29823 , y29824 , y29825 , y29826 , y29827 , y29828 , y29829 , y29830 , y29831 , y29832 , y29833 , y29834 , y29835 , y29836 , y29837 , y29838 , y29839 , y29840 , y29841 , y29842 , y29843 , y29844 , y29845 , y29846 , y29847 , y29848 , y29849 , y29850 , y29851 , y29852 , y29853 , y29854 , y29855 , y29856 , y29857 , y29858 , y29859 , y29860 , y29861 , y29862 , y29863 , y29864 , y29865 , y29866 , y29867 , y29868 , y29869 , y29870 , y29871 , y29872 , y29873 , y29874 , y29875 , y29876 , y29877 , y29878 , y29879 , y29880 , y29881 , y29882 , y29883 , y29884 , y29885 , y29886 , y29887 , y29888 , y29889 , y29890 , y29891 , y29892 , y29893 , y29894 , y29895 , y29896 , y29897 , y29898 , y29899 , y29900 , y29901 , y29902 , y29903 , y29904 , y29905 , y29906 , y29907 , y29908 , y29909 , y29910 , y29911 , y29912 , y29913 , y29914 , y29915 , y29916 , y29917 , y29918 , y29919 , y29920 , y29921 , y29922 , y29923 , y29924 , y29925 , y29926 , y29927 , y29928 , y29929 , y29930 , y29931 , y29932 , y29933 , y29934 , y29935 , y29936 , y29937 , y29938 , y29939 , y29940 , y29941 , y29942 , y29943 , y29944 , y29945 , y29946 , y29947 , y29948 , y29949 , y29950 , y29951 , y29952 , y29953 , y29954 , y29955 , y29956 , y29957 , y29958 , y29959 , y29960 , y29961 , y29962 , y29963 , y29964 , y29965 , y29966 , y29967 , y29968 , y29969 , y29970 , y29971 , y29972 , y29973 , y29974 , y29975 , y29976 , y29977 , y29978 , y29979 , y29980 , y29981 , y29982 , y29983 , y29984 , y29985 , y29986 , y29987 , y29988 , y29989 , y29990 , y29991 , y29992 , y29993 , y29994 , y29995 , y29996 , y29997 , y29998 , y29999 , y30000 , y30001 , y30002 , y30003 , y30004 , y30005 , y30006 , y30007 , y30008 , y30009 , y30010 , y30011 , y30012 , y30013 , y30014 , y30015 , y30016 , y30017 , y30018 , y30019 , y30020 , y30021 , y30022 , y30023 , y30024 , y30025 , y30026 , y30027 , y30028 , y30029 , y30030 , y30031 , y30032 , y30033 , y30034 , y30035 , y30036 , y30037 , y30038 , y30039 , y30040 , y30041 , y30042 , y30043 , y30044 , y30045 , y30046 , y30047 , y30048 , y30049 , y30050 , y30051 , y30052 , y30053 , y30054 , y30055 , y30056 , y30057 , y30058 , y30059 , y30060 , y30061 , y30062 , y30063 , y30064 , y30065 , y30066 , y30067 , y30068 , y30069 , y30070 , y30071 , y30072 , y30073 , y30074 , y30075 , y30076 , y30077 , y30078 , y30079 , y30080 , y30081 , y30082 , y30083 , y30084 , y30085 , y30086 , y30087 , y30088 , y30089 , y30090 , y30091 , y30092 , y30093 , y30094 , y30095 , y30096 , y30097 , y30098 , y30099 , y30100 , y30101 , y30102 , y30103 , y30104 , y30105 , y30106 , y30107 , y30108 , y30109 , y30110 , y30111 , y30112 , y30113 , y30114 , y30115 , y30116 , y30117 , y30118 , y30119 , y30120 , y30121 , y30122 , y30123 , y30124 , y30125 , y30126 , y30127 , y30128 , y30129 , y30130 , y30131 , y30132 , y30133 , y30134 , y30135 , y30136 , y30137 , y30138 , y30139 , y30140 , y30141 , y30142 , y30143 , y30144 , y30145 , y30146 , y30147 , y30148 , y30149 , y30150 , y30151 , y30152 , y30153 , y30154 , y30155 , y30156 , y30157 , y30158 , y30159 , y30160 , y30161 , y30162 , y30163 , y30164 , y30165 , y30166 , y30167 , y30168 , y30169 , y30170 , y30171 , y30172 , y30173 , y30174 , y30175 , y30176 , y30177 , y30178 , y30179 , y30180 , y30181 , y30182 , y30183 , y30184 , y30185 , y30186 , y30187 , y30188 , y30189 , y30190 , y30191 , y30192 , y30193 , y30194 , y30195 , y30196 , y30197 , y30198 , y30199 , y30200 , y30201 , y30202 , y30203 , y30204 , y30205 , y30206 , y30207 , y30208 , y30209 , y30210 , y30211 , y30212 , y30213 , y30214 , y30215 , y30216 , y30217 , y30218 , y30219 , y30220 , y30221 , y30222 , y30223 , y30224 , y30225 , y30226 , y30227 , y30228 , y30229 , y30230 , y30231 , y30232 , y30233 , y30234 , y30235 , y30236 , y30237 , y30238 , y30239 , y30240 , y30241 , y30242 , y30243 , y30244 , y30245 , y30246 , y30247 , y30248 , y30249 , y30250 , y30251 , y30252 , y30253 , y30254 , y30255 , y30256 , y30257 , y30258 , y30259 , y30260 , y30261 , y30262 , y30263 , y30264 , y30265 , y30266 , y30267 , y30268 , y30269 , y30270 , y30271 , y30272 , y30273 , y30274 , y30275 , y30276 , y30277 , y30278 , y30279 , y30280 , y30281 , y30282 , y30283 , y30284 , y30285 , y30286 , y30287 , y30288 , y30289 , y30290 , y30291 , y30292 , y30293 , y30294 , y30295 , y30296 , y30297 , y30298 , y30299 , y30300 , y30301 , y30302 , y30303 , y30304 , y30305 , y30306 , y30307 , y30308 , y30309 , y30310 , y30311 , y30312 , y30313 , y30314 , y30315 , y30316 , y30317 , y30318 , y30319 , y30320 , y30321 , y30322 , y30323 , y30324 , y30325 , y30326 , y30327 , y30328 , y30329 , y30330 , y30331 , y30332 , y30333 , y30334 , y30335 , y30336 , y30337 , y30338 , y30339 , y30340 , y30341 , y30342 , y30343 , y30344 , y30345 , y30346 , y30347 , y30348 , y30349 , y30350 , y30351 , y30352 , y30353 , y30354 , y30355 , y30356 , y30357 , y30358 , y30359 , y30360 , y30361 , y30362 , y30363 , y30364 , y30365 , y30366 , y30367 , y30368 , y30369 , y30370 , y30371 , y30372 , y30373 , y30374 , y30375 , y30376 , y30377 , y30378 , y30379 , y30380 , y30381 , y30382 , y30383 , y30384 , y30385 , y30386 , y30387 , y30388 , y30389 , y30390 , y30391 , y30392 , y30393 , y30394 , y30395 , y30396 , y30397 , y30398 , y30399 , y30400 , y30401 , y30402 , y30403 , y30404 , y30405 , y30406 , y30407 , y30408 , y30409 , y30410 , y30411 , y30412 ;
  wire n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , n18511 , n18512 , n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , n18679 , n18680 , n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , n18709 , n18710 , n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , n18841 , n18842 , n18843 , n18844 , n18845 , n18846 , n18847 , n18848 , n18849 , n18850 , n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , n18870 , n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , n18891 , n18892 , n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , n18910 , n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , n18921 , n18922 , n18923 , n18924 , n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , n18969 , n18970 , n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , n18977 , n18978 , n18979 , n18980 , n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , n18989 , n18990 , n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , n18999 , n19000 , n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , n19017 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , n19029 , n19030 , n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , n19037 , n19038 , n19039 , n19040 , n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , n19049 , n19050 , n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , n19060 , n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , n19067 , n19068 , n19069 , n19070 , n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , n19079 , n19080 , n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , n19089 , n19090 , n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , n19099 , n19100 , n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , n19137 , n19138 , n19139 , n19140 , n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , n19157 , n19158 , n19159 , n19160 , n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , n19167 , n19168 , n19169 , n19170 , n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , n19179 , n19180 , n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , n19189 , n19190 , n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , n19198 , n19199 , n19200 , n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , n19210 , n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , n19217 , n19218 , n19219 , n19220 , n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , n19229 , n19230 , n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , n19239 , n19240 , n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , n19249 , n19250 , n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , n19259 , n19260 , n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , n19279 , n19280 , n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , n19287 , n19288 , n19289 , n19290 , n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , n19297 , n19298 , n19299 , n19300 , n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , n19309 , n19310 , n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , n19319 , n19320 , n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , n19329 , n19330 , n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , n19339 , n19340 , n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , n19359 , n19360 , n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , n19369 , n19370 , n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , n19379 , n19380 , n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19387 , n19388 , n19389 , n19390 , n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , n19400 , n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , n19410 , n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , n19417 , n19418 , n19419 , n19420 , n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , n19440 , n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , n19450 , n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , n19459 , n19460 , n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , n19470 , n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , n19529 , n19530 , n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , n19550 , n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , n19567 , n19568 , n19569 , n19570 , n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , n19587 , n19588 , n19589 , n19590 , n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , n19619 , n19620 , n19621 , n19622 , n19623 , n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , n19670 , n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , n19711 , n19712 , n19713 , n19714 , n19715 , n19716 , n19717 , n19718 , n19719 , n19720 , n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , n19737 , n19738 , n19739 , n19740 , n19741 , n19742 , n19743 , n19744 , n19745 , n19746 , n19747 , n19748 , n19749 , n19750 , n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , n19757 , n19758 , n19759 , n19760 , n19761 , n19762 , n19763 , n19764 , n19765 , n19766 , n19767 , n19768 , n19769 , n19770 , n19771 , n19772 , n19773 , n19774 , n19775 , n19776 , n19777 , n19778 , n19779 , n19780 , n19781 , n19782 , n19783 , n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , n19791 , n19792 , n19793 , n19794 , n19795 , n19796 , n19797 , n19798 , n19799 , n19800 , n19801 , n19802 , n19803 , n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , n19811 , n19812 , n19813 , n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , n19821 , n19822 , n19823 , n19824 , n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , n19831 , n19832 , n19833 , n19834 , n19835 , n19836 , n19837 , n19838 , n19839 , n19840 , n19841 , n19842 , n19843 , n19844 , n19845 , n19846 , n19847 , n19848 , n19849 , n19850 , n19851 , n19852 , n19853 , n19854 , n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , n19861 , n19862 , n19863 , n19864 , n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , n19871 , n19872 , n19873 , n19874 , n19875 , n19876 , n19877 , n19878 , n19879 , n19880 , n19881 , n19882 , n19883 , n19884 , n19885 , n19886 , n19887 , n19888 , n19889 , n19890 , n19891 , n19892 , n19893 , n19894 , n19895 , n19896 , n19897 , n19898 , n19899 , n19900 , n19901 , n19902 , n19903 , n19904 , n19905 , n19906 , n19907 , n19908 , n19909 , n19910 , n19911 , n19912 , n19913 , n19914 , n19915 , n19916 , n19917 , n19918 , n19919 , n19920 , n19921 , n19922 , n19923 , n19924 , n19925 , n19926 , n19927 , n19928 , n19929 , n19930 , n19931 , n19932 , n19933 , n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , n19940 , n19941 , n19942 , n19943 , n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , n19951 , n19952 , n19953 , n19954 , n19955 , n19956 , n19957 , n19958 , n19959 , n19960 , n19961 , n19962 , n19963 , n19964 , n19965 , n19966 , n19967 , n19968 , n19969 , n19970 , n19971 , n19972 , n19973 , n19974 , n19975 , n19976 , n19977 , n19978 , n19979 , n19980 , n19981 , n19982 , n19983 , n19984 , n19985 , n19986 , n19987 , n19988 , n19989 , n19990 , n19991 , n19992 , n19993 , n19994 , n19995 , n19996 , n19997 , n19998 , n19999 , n20000 , n20001 , n20002 , n20003 , n20004 , n20005 , n20006 , n20007 , n20008 , n20009 , n20010 , n20011 , n20012 , n20013 , n20014 , n20015 , n20016 , n20017 , n20018 , n20019 , n20020 , n20021 , n20022 , n20023 , n20024 , n20025 , n20026 , n20027 , n20028 , n20029 , n20030 , n20031 , n20032 , n20033 , n20034 , n20035 , n20036 , n20037 , n20038 , n20039 , n20040 , n20041 , n20042 , n20043 , n20044 , n20045 , n20046 , n20047 , n20048 , n20049 , n20050 , n20051 , n20052 , n20053 , n20054 , n20055 , n20056 , n20057 , n20058 , n20059 , n20060 , n20061 , n20062 , n20063 , n20064 , n20065 , n20066 , n20067 , n20068 , n20069 , n20070 , n20071 , n20072 , n20073 , n20074 , n20075 , n20076 , n20077 , n20078 , n20079 , n20080 , n20081 , n20082 , n20083 , n20084 , n20085 , n20086 , n20087 , n20088 , n20089 , n20090 , n20091 , n20092 , n20093 , n20094 , n20095 , n20096 , n20097 , n20098 , n20099 , n20100 , n20101 , n20102 , n20103 , n20104 , n20105 , n20106 , n20107 , n20108 , n20109 , n20110 , n20111 , n20112 , n20113 , n20114 , n20115 , n20116 , n20117 , n20118 , n20119 , n20120 , n20121 , n20122 , n20123 , n20124 , n20125 , n20126 , n20127 , n20128 , n20129 , n20130 , n20131 , n20132 , n20133 , n20134 , n20135 , n20136 , n20137 , n20138 , n20139 , n20140 , n20141 , n20142 , n20143 , n20144 , n20145 , n20146 , n20147 , n20148 , n20149 , n20150 , n20151 , n20152 , n20153 , n20154 , n20155 , n20156 , n20157 , n20158 , n20159 , n20160 , n20161 , n20162 , n20163 , n20164 , n20165 , n20166 , n20167 , n20168 , n20169 , n20170 , n20171 , n20172 , n20173 , n20174 , n20175 , n20176 , n20177 , n20178 , n20179 , n20180 , n20181 , n20182 , n20183 , n20184 , n20185 , n20186 , n20187 , n20188 , n20189 , n20190 , n20191 , n20192 , n20193 , n20194 , n20195 , n20196 , n20197 , n20198 , n20199 , n20200 , n20201 , n20202 , n20203 , n20204 , n20205 , n20206 , n20207 , n20208 , n20209 , n20210 , n20211 , n20212 , n20213 , n20214 , n20215 , n20216 , n20217 , n20218 , n20219 , n20220 , n20221 , n20222 , n20223 , n20224 , n20225 , n20226 , n20227 , n20228 , n20229 , n20230 , n20231 , n20232 , n20233 , n20234 , n20235 , n20236 , n20237 , n20238 , n20239 , n20240 , n20241 , n20242 , n20243 , n20244 , n20245 , n20246 , n20247 , n20248 , n20249 , n20250 , n20251 , n20252 , n20253 , n20254 , n20255 , n20256 , n20257 , n20258 , n20259 , n20260 , n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , n20267 , n20268 , n20269 , n20270 , n20271 , n20272 , n20273 , n20274 , n20275 , n20276 , n20277 , n20278 , n20279 , n20280 , n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , n20287 , n20288 , n20289 , n20290 , n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , n20297 , n20298 , n20299 , n20300 , n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , n20307 , n20308 , n20309 , n20310 , n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , n20317 , n20318 , n20319 , n20320 , n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , n20327 , n20328 , n20329 , n20330 , n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , n20337 , n20338 , n20339 , n20340 , n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , n20347 , n20348 , n20349 , n20350 , n20351 , n20352 , n20353 , n20354 , n20355 , n20356 , n20357 , n20358 , n20359 , n20360 , n20361 , n20362 , n20363 , n20364 , n20365 , n20366 , n20367 , n20368 , n20369 , n20370 , n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , n20377 , n20378 , n20379 , n20380 , n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , n20389 , n20390 , n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , n20397 , n20398 , n20399 , n20400 , n20401 , n20402 , n20403 , n20404 , n20405 , n20406 , n20407 , n20408 , n20409 , n20410 , n20411 , n20412 , n20413 , n20414 , n20415 , n20416 , n20417 , n20418 , n20419 , n20420 , n20421 , n20422 , n20423 , n20424 , n20425 , n20426 , n20427 , n20428 , n20429 , n20430 , n20431 , n20432 , n20433 , n20434 , n20435 , n20436 , n20437 , n20438 , n20439 , n20440 , n20441 , n20442 , n20443 , n20444 , n20445 , n20446 , n20447 , n20448 , n20449 , n20450 , n20451 , n20452 , n20453 , n20454 , n20455 , n20456 , n20457 , n20458 , n20459 , n20460 , n20461 , n20462 , n20463 , n20464 , n20465 , n20466 , n20467 , n20468 , n20469 , n20470 , n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , n20477 , n20478 , n20479 , n20480 , n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , n20487 , n20488 , n20489 , n20490 , n20491 , n20492 , n20493 , n20494 , n20495 , n20496 , n20497 , n20498 , n20499 , n20500 , n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , n20507 , n20508 , n20509 , n20510 , n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , n20519 , n20520 , n20521 , n20522 , n20523 , n20524 , n20525 , n20526 , n20527 , n20528 , n20529 , n20530 , n20531 , n20532 , n20533 , n20534 , n20535 , n20536 , n20537 , n20538 , n20539 , n20540 , n20541 , n20542 , n20543 , n20544 , n20545 , n20546 , n20547 , n20548 , n20549 , n20550 , n20551 , n20552 , n20553 , n20554 , n20555 , n20556 , n20557 , n20558 , n20559 , n20560 , n20561 , n20562 , n20563 , n20564 , n20565 , n20566 , n20567 , n20568 , n20569 , n20570 , n20571 , n20572 , n20573 , n20574 , n20575 , n20576 , n20577 , n20578 , n20579 , n20580 , n20581 , n20582 , n20583 , n20584 , n20585 , n20586 , n20587 , n20588 , n20589 , n20590 , n20591 , n20592 , n20593 , n20594 , n20595 , n20596 , n20597 , n20598 , n20599 , n20600 , n20601 , n20602 , n20603 , n20604 , n20605 , n20606 , n20607 , n20608 , n20609 , n20610 , n20611 , n20612 , n20613 , n20614 , n20615 , n20616 , n20617 , n20618 , n20619 , n20620 , n20621 , n20622 , n20623 , n20624 , n20625 , n20626 , n20627 , n20628 , n20629 , n20630 , n20631 , n20632 , n20633 , n20634 , n20635 , n20636 , n20637 , n20638 , n20639 , n20640 , n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , n20647 , n20648 , n20649 , n20650 , n20651 , n20652 , n20653 , n20654 , n20655 , n20656 , n20657 , n20658 , n20659 , n20660 , n20661 , n20662 , n20663 , n20664 , n20665 , n20666 , n20667 , n20668 , n20669 , n20670 , n20671 , n20672 , n20673 , n20674 , n20675 , n20676 , n20677 , n20678 , n20679 , n20680 , n20681 , n20682 , n20683 , n20684 , n20685 , n20686 , n20687 , n20688 , n20689 , n20690 , n20691 , n20692 , n20693 , n20694 , n20695 , n20696 , n20697 , n20698 , n20699 , n20700 , n20701 , n20702 , n20703 , n20704 , n20705 , n20706 , n20707 , n20708 , n20709 , n20710 , n20711 , n20712 , n20713 , n20714 , n20715 , n20716 , n20717 , n20718 , n20719 , n20720 , n20721 , n20722 , n20723 , n20724 , n20725 , n20726 , n20727 , n20728 , n20729 , n20730 , n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , n20737 , n20738 , n20739 , n20740 , n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , n20747 , n20748 , n20749 , n20750 , n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , n20757 , n20758 , n20759 , n20760 , n20761 , n20762 , n20763 , n20764 , n20765 , n20766 , n20767 , n20768 , n20769 , n20770 , n20771 , n20772 , n20773 , n20774 , n20775 , n20776 , n20777 , n20778 , n20779 , n20780 , n20781 , n20782 , n20783 , n20784 , n20785 , n20786 , n20787 , n20788 , n20789 , n20790 , n20791 , n20792 , n20793 , n20794 , n20795 , n20796 , n20797 , n20798 , n20799 , n20800 , n20801 , n20802 , n20803 , n20804 , n20805 , n20806 , n20807 , n20808 , n20809 , n20810 , n20811 , n20812 , n20813 , n20814 , n20815 , n20816 , n20817 , n20818 , n20819 , n20820 , n20821 , n20822 , n20823 , n20824 , n20825 , n20826 , n20827 , n20828 , n20829 , n20830 , n20831 , n20832 , n20833 , n20834 , n20835 , n20836 , n20837 , n20838 , n20839 , n20840 , n20841 , n20842 , n20843 , n20844 , n20845 , n20846 , n20847 , n20848 , n20849 , n20850 , n20851 , n20852 , n20853 , n20854 , n20855 , n20856 , n20857 , n20858 , n20859 , n20860 , n20861 , n20862 , n20863 , n20864 , n20865 , n20866 , n20867 , n20868 , n20869 , n20870 , n20871 , n20872 , n20873 , n20874 , n20875 , n20876 , n20877 , n20878 , n20879 , n20880 , n20881 , n20882 , n20883 , n20884 , n20885 , n20886 , n20887 , n20888 , n20889 , n20890 , n20891 , n20892 , n20893 , n20894 , n20895 , n20896 , n20897 , n20898 , n20899 , n20900 , n20901 , n20902 , n20903 , n20904 , n20905 , n20906 , n20907 , n20908 , n20909 , n20910 , n20911 , n20912 , n20913 , n20914 , n20915 , n20916 , n20917 , n20918 , n20919 , n20920 , n20921 , n20922 , n20923 , n20924 , n20925 , n20926 , n20927 , n20928 , n20929 , n20930 , n20931 , n20932 , n20933 , n20934 , n20935 , n20936 , n20937 , n20938 , n20939 , n20940 , n20941 , n20942 , n20943 , n20944 , n20945 , n20946 , n20947 , n20948 , n20949 , n20950 , n20951 , n20952 , n20953 , n20954 , n20955 , n20956 , n20957 , n20958 , n20959 , n20960 , n20961 , n20962 , n20963 , n20964 , n20965 , n20966 , n20967 , n20968 , n20969 , n20970 , n20971 , n20972 , n20973 , n20974 , n20975 , n20976 , n20977 , n20978 , n20979 , n20980 , n20981 , n20982 , n20983 , n20984 , n20985 , n20986 , n20987 , n20988 , n20989 , n20990 , n20991 , n20992 , n20993 , n20994 , n20995 , n20996 , n20997 , n20998 , n20999 , n21000 , n21001 , n21002 , n21003 , n21004 , n21005 , n21006 , n21007 , n21008 , n21009 , n21010 , n21011 , n21012 , n21013 , n21014 , n21015 , n21016 , n21017 , n21018 , n21019 , n21020 , n21021 , n21022 , n21023 , n21024 , n21025 , n21026 , n21027 , n21028 , n21029 , n21030 , n21031 , n21032 , n21033 , n21034 , n21035 , n21036 , n21037 , n21038 , n21039 , n21040 , n21041 , n21042 , n21043 , n21044 , n21045 , n21046 , n21047 , n21048 , n21049 , n21050 , n21051 , n21052 , n21053 , n21054 , n21055 , n21056 , n21057 , n21058 , n21059 , n21060 , n21061 , n21062 , n21063 , n21064 , n21065 , n21066 , n21067 , n21068 , n21069 , n21070 , n21071 , n21072 , n21073 , n21074 , n21075 , n21076 , n21077 , n21078 , n21079 , n21080 , n21081 , n21082 , n21083 , n21084 , n21085 , n21086 , n21087 , n21088 , n21089 , n21090 , n21091 , n21092 , n21093 , n21094 , n21095 , n21096 , n21097 , n21098 , n21099 , n21100 , n21101 , n21102 , n21103 , n21104 , n21105 , n21106 , n21107 , n21108 , n21109 , n21110 , n21111 , n21112 , n21113 , n21114 , n21115 , n21116 , n21117 , n21118 , n21119 , n21120 , n21121 , n21122 , n21123 , n21124 , n21125 , n21126 , n21127 , n21128 , n21129 , n21130 , n21131 , n21132 , n21133 , n21134 , n21135 , n21136 , n21137 , n21138 , n21139 , n21140 , n21141 , n21142 , n21143 , n21144 , n21145 , n21146 , n21147 , n21148 , n21149 , n21150 , n21151 , n21152 , n21153 , n21154 , n21155 , n21156 , n21157 , n21158 , n21159 , n21160 , n21161 , n21162 , n21163 , n21164 , n21165 , n21166 , n21167 , n21168 , n21169 , n21170 , n21171 , n21172 , n21173 , n21174 , n21175 , n21176 , n21177 , n21178 , n21179 , n21180 , n21181 , n21182 , n21183 , n21184 , n21185 , n21186 , n21187 , n21188 , n21189 , n21190 , n21191 , n21192 , n21193 , n21194 , n21195 , n21196 , n21197 , n21198 , n21199 , n21200 , n21201 , n21202 , n21203 , n21204 , n21205 , n21206 , n21207 , n21208 , n21209 , n21210 , n21211 , n21212 , n21213 , n21214 , n21215 , n21216 , n21217 , n21218 , n21219 , n21220 , n21221 , n21222 , n21223 , n21224 , n21225 , n21226 , n21227 , n21228 , n21229 , n21230 , n21231 , n21232 , n21233 , n21234 , n21235 , n21236 , n21237 , n21238 , n21239 , n21240 , n21241 , n21242 , n21243 , n21244 , n21245 , n21246 , n21247 , n21248 , n21249 , n21250 , n21251 , n21252 , n21253 , n21254 , n21255 , n21256 , n21257 , n21258 , n21259 , n21260 , n21261 , n21262 , n21263 , n21264 , n21265 , n21266 , n21267 , n21268 , n21269 , n21270 , n21271 , n21272 , n21273 , n21274 , n21275 , n21276 , n21277 , n21278 , n21279 , n21280 , n21281 , n21282 , n21283 , n21284 , n21285 , n21286 , n21287 , n21288 , n21289 , n21290 , n21291 , n21292 , n21293 , n21294 , n21295 , n21296 , n21297 , n21298 , n21299 , n21300 , n21301 , n21302 , n21303 , n21304 , n21305 , n21306 , n21307 , n21308 , n21309 , n21310 , n21311 , n21312 , n21313 , n21314 , n21315 , n21316 , n21317 , n21318 , n21319 , n21320 , n21321 , n21322 , n21323 , n21324 , n21325 , n21326 , n21327 , n21328 , n21329 , n21330 , n21331 , n21332 , n21333 , n21334 , n21335 , n21336 , n21337 , n21338 , n21339 , n21340 , n21341 , n21342 , n21343 , n21344 , n21345 , n21346 , n21347 , n21348 , n21349 , n21350 , n21351 , n21352 , n21353 , n21354 , n21355 , n21356 , n21357 , n21358 , n21359 , n21360 , n21361 , n21362 , n21363 , n21364 , n21365 , n21366 , n21367 , n21368 , n21369 , n21370 , n21371 , n21372 , n21373 , n21374 , n21375 , n21376 , n21377 , n21378 , n21379 , n21380 , n21381 , n21382 , n21383 , n21384 , n21385 , n21386 , n21387 , n21388 , n21389 , n21390 , n21391 , n21392 , n21393 , n21394 , n21395 , n21396 , n21397 , n21398 , n21399 , n21400 , n21401 , n21402 , n21403 , n21404 , n21405 , n21406 , n21407 , n21408 , n21409 , n21410 , n21411 , n21412 , n21413 , n21414 , n21415 , n21416 , n21417 , n21418 , n21419 , n21420 , n21421 , n21422 , n21423 , n21424 , n21425 , n21426 , n21427 , n21428 , n21429 , n21430 , n21431 , n21432 , n21433 , n21434 , n21435 , n21436 , n21437 , n21438 , n21439 , n21440 , n21441 , n21442 , n21443 , n21444 , n21445 , n21446 , n21447 , n21448 , n21449 , n21450 , n21451 , n21452 , n21453 , n21454 , n21455 , n21456 , n21457 , n21458 , n21459 , n21460 , n21461 , n21462 , n21463 , n21464 , n21465 , n21466 , n21467 , n21468 , n21469 , n21470 , n21471 , n21472 , n21473 , n21474 , n21475 , n21476 , n21477 , n21478 , n21479 , n21480 , n21481 , n21482 , n21483 , n21484 , n21485 , n21486 , n21487 , n21488 , n21489 , n21490 , n21491 , n21492 , n21493 , n21494 , n21495 , n21496 , n21497 , n21498 , n21499 , n21500 , n21501 , n21502 , n21503 , n21504 , n21505 , n21506 , n21507 , n21508 , n21509 , n21510 , n21511 , n21512 , n21513 , n21514 , n21515 , n21516 , n21517 , n21518 , n21519 , n21520 , n21521 , n21522 , n21523 , n21524 , n21525 , n21526 , n21527 , n21528 , n21529 , n21530 , n21531 , n21532 , n21533 , n21534 , n21535 , n21536 , n21537 , n21538 , n21539 , n21540 , n21541 , n21542 , n21543 , n21544 , n21545 , n21546 , n21547 , n21548 , n21549 , n21550 , n21551 , n21552 , n21553 , n21554 , n21555 , n21556 , n21557 , n21558 , n21559 , n21560 , n21561 , n21562 , n21563 , n21564 , n21565 , n21566 , n21567 , n21568 , n21569 , n21570 , n21571 , n21572 , n21573 , n21574 , n21575 , n21576 , n21577 , n21578 , n21579 , n21580 , n21581 , n21582 , n21583 , n21584 , n21585 , n21586 , n21587 , n21588 , n21589 , n21590 , n21591 , n21592 , n21593 , n21594 , n21595 , n21596 , n21597 , n21598 , n21599 , n21600 , n21601 , n21602 , n21603 , n21604 , n21605 , n21606 , n21607 , n21608 , n21609 , n21610 , n21611 , n21612 , n21613 , n21614 , n21615 , n21616 , n21617 , n21618 , n21619 , n21620 , n21621 , n21622 , n21623 , n21624 , n21625 , n21626 , n21627 , n21628 , n21629 , n21630 , n21631 , n21632 , n21633 , n21634 , n21635 , n21636 , n21637 , n21638 , n21639 , n21640 , n21641 , n21642 , n21643 , n21644 , n21645 , n21646 , n21647 , n21648 , n21649 , n21650 , n21651 , n21652 , n21653 , n21654 , n21655 , n21656 , n21657 , n21658 , n21659 , n21660 , n21661 , n21662 , n21663 , n21664 , n21665 , n21666 , n21667 , n21668 , n21669 , n21670 , n21671 , n21672 , n21673 , n21674 , n21675 , n21676 , n21677 , n21678 , n21679 , n21680 , n21681 , n21682 , n21683 , n21684 , n21685 , n21686 , n21687 , n21688 , n21689 , n21690 , n21691 , n21692 , n21693 , n21694 , n21695 , n21696 , n21697 , n21698 , n21699 , n21700 , n21701 , n21702 , n21703 , n21704 , n21705 , n21706 , n21707 , n21708 , n21709 , n21710 , n21711 , n21712 , n21713 , n21714 , n21715 , n21716 , n21717 , n21718 , n21719 , n21720 , n21721 , n21722 , n21723 , n21724 , n21725 , n21726 , n21727 , n21728 , n21729 , n21730 , n21731 , n21732 , n21733 , n21734 , n21735 , n21736 , n21737 , n21738 , n21739 , n21740 , n21741 , n21742 , n21743 , n21744 , n21745 , n21746 , n21747 , n21748 , n21749 , n21750 , n21751 , n21752 , n21753 , n21754 , n21755 , n21756 , n21757 , n21758 , n21759 , n21760 , n21761 , n21762 , n21763 , n21764 , n21765 , n21766 , n21767 , n21768 , n21769 , n21770 , n21771 , n21772 , n21773 , n21774 , n21775 , n21776 , n21777 , n21778 , n21779 , n21780 , n21781 , n21782 , n21783 , n21784 , n21785 , n21786 , n21787 , n21788 , n21789 , n21790 , n21791 , n21792 , n21793 , n21794 , n21795 , n21796 , n21797 , n21798 , n21799 , n21800 , n21801 , n21802 , n21803 , n21804 , n21805 , n21806 , n21807 , n21808 , n21809 , n21810 , n21811 , n21812 , n21813 , n21814 , n21815 , n21816 , n21817 , n21818 , n21819 , n21820 , n21821 , n21822 , n21823 , n21824 , n21825 , n21826 , n21827 , n21828 , n21829 , n21830 , n21831 , n21832 , n21833 , n21834 , n21835 , n21836 , n21837 , n21838 , n21839 , n21840 , n21841 , n21842 , n21843 , n21844 , n21845 , n21846 , n21847 , n21848 , n21849 , n21850 , n21851 , n21852 , n21853 , n21854 , n21855 , n21856 , n21857 , n21858 , n21859 , n21860 , n21861 , n21862 , n21863 , n21864 , n21865 , n21866 , n21867 , n21868 , n21869 , n21870 , n21871 , n21872 , n21873 , n21874 , n21875 , n21876 , n21877 , n21878 , n21879 , n21880 , n21881 , n21882 , n21883 , n21884 , n21885 , n21886 , n21887 , n21888 , n21889 , n21890 , n21891 , n21892 , n21893 , n21894 , n21895 , n21896 , n21897 , n21898 , n21899 , n21900 , n21901 , n21902 , n21903 , n21904 , n21905 , n21906 , n21907 , n21908 , n21909 , n21910 , n21911 , n21912 , n21913 , n21914 , n21915 , n21916 , n21917 , n21918 , n21919 , n21920 , n21921 , n21922 , n21923 , n21924 , n21925 , n21926 , n21927 , n21928 , n21929 , n21930 , n21931 , n21932 , n21933 , n21934 , n21935 , n21936 , n21937 , n21938 , n21939 , n21940 , n21941 , n21942 , n21943 , n21944 , n21945 , n21946 , n21947 , n21948 , n21949 , n21950 , n21951 , n21952 , n21953 , n21954 , n21955 , n21956 , n21957 , n21958 , n21959 , n21960 , n21961 , n21962 , n21963 , n21964 , n21965 , n21966 , n21967 , n21968 , n21969 , n21970 , n21971 , n21972 , n21973 , n21974 , n21975 , n21976 , n21977 , n21978 , n21979 , n21980 , n21981 , n21982 , n21983 , n21984 , n21985 , n21986 , n21987 , n21988 , n21989 , n21990 , n21991 , n21992 , n21993 , n21994 , n21995 , n21996 , n21997 , n21998 , n21999 , n22000 , n22001 , n22002 , n22003 , n22004 , n22005 , n22006 , n22007 , n22008 , n22009 , n22010 , n22011 , n22012 , n22013 , n22014 , n22015 , n22016 , n22017 , n22018 , n22019 , n22020 , n22021 , n22022 , n22023 , n22024 , n22025 , n22026 , n22027 , n22028 , n22029 , n22030 , n22031 , n22032 , n22033 , n22034 , n22035 , n22036 , n22037 , n22038 , n22039 , n22040 , n22041 , n22042 , n22043 , n22044 , n22045 , n22046 , n22047 , n22048 , n22049 , n22050 , n22051 , n22052 , n22053 , n22054 , n22055 , n22056 , n22057 , n22058 , n22059 , n22060 , n22061 , n22062 , n22063 , n22064 , n22065 , n22066 , n22067 , n22068 , n22069 , n22070 , n22071 , n22072 , n22073 , n22074 , n22075 , n22076 , n22077 , n22078 , n22079 , n22080 , n22081 , n22082 , n22083 , n22084 , n22085 , n22086 , n22087 , n22088 , n22089 , n22090 , n22091 , n22092 , n22093 , n22094 , n22095 , n22096 , n22097 , n22098 , n22099 , n22100 , n22101 , n22102 , n22103 , n22104 , n22105 , n22106 , n22107 , n22108 , n22109 , n22110 , n22111 , n22112 , n22113 , n22114 , n22115 , n22116 , n22117 , n22118 , n22119 , n22120 , n22121 , n22122 , n22123 , n22124 , n22125 , n22126 , n22127 , n22128 , n22129 , n22130 , n22131 , n22132 , n22133 , n22134 , n22135 , n22136 , n22137 , n22138 , n22139 , n22140 , n22141 , n22142 , n22143 , n22144 , n22145 , n22146 , n22147 , n22148 , n22149 , n22150 , n22151 , n22152 , n22153 , n22154 , n22155 , n22156 , n22157 , n22158 , n22159 , n22160 , n22161 , n22162 , n22163 , n22164 , n22165 , n22166 , n22167 , n22168 , n22169 , n22170 , n22171 , n22172 , n22173 , n22174 , n22175 , n22176 , n22177 , n22178 , n22179 , n22180 , n22181 , n22182 , n22183 , n22184 , n22185 , n22186 , n22187 , n22188 , n22189 , n22190 , n22191 , n22192 , n22193 , n22194 , n22195 , n22196 , n22197 , n22198 , n22199 , n22200 , n22201 , n22202 , n22203 , n22204 , n22205 , n22206 , n22207 , n22208 , n22209 , n22210 , n22211 , n22212 , n22213 , n22214 , n22215 , n22216 , n22217 , n22218 , n22219 , n22220 , n22221 , n22222 , n22223 , n22224 , n22225 , n22226 , n22227 , n22228 , n22229 , n22230 , n22231 , n22232 , n22233 , n22234 , n22235 , n22236 , n22237 , n22238 , n22239 , n22240 , n22241 , n22242 , n22243 , n22244 , n22245 , n22246 , n22247 , n22248 , n22249 , n22250 , n22251 , n22252 , n22253 , n22254 , n22255 , n22256 , n22257 , n22258 , n22259 , n22260 , n22261 , n22262 , n22263 , n22264 , n22265 , n22266 , n22267 , n22268 , n22269 , n22270 , n22271 , n22272 , n22273 , n22274 , n22275 , n22276 , n22277 , n22278 , n22279 , n22280 , n22281 , n22282 , n22283 , n22284 , n22285 , n22286 , n22287 , n22288 , n22289 , n22290 , n22291 , n22292 , n22293 , n22294 , n22295 , n22296 , n22297 , n22298 , n22299 , n22300 , n22301 , n22302 , n22303 , n22304 , n22305 , n22306 , n22307 , n22308 , n22309 , n22310 , n22311 , n22312 , n22313 , n22314 , n22315 , n22316 , n22317 , n22318 , n22319 , n22320 , n22321 , n22322 , n22323 , n22324 , n22325 , n22326 , n22327 , n22328 , n22329 , n22330 , n22331 , n22332 , n22333 , n22334 , n22335 , n22336 , n22337 , n22338 , n22339 , n22340 , n22341 , n22342 , n22343 , n22344 , n22345 , n22346 , n22347 , n22348 , n22349 , n22350 , n22351 , n22352 , n22353 , n22354 , n22355 , n22356 , n22357 , n22358 , n22359 , n22360 , n22361 , n22362 , n22363 , n22364 , n22365 , n22366 , n22367 , n22368 , n22369 , n22370 , n22371 , n22372 , n22373 , n22374 , n22375 , n22376 , n22377 , n22378 , n22379 , n22380 , n22381 , n22382 , n22383 , n22384 , n22385 , n22386 , n22387 , n22388 , n22389 , n22390 , n22391 , n22392 , n22393 , n22394 , n22395 , n22396 , n22397 , n22398 , n22399 , n22400 , n22401 , n22402 , n22403 , n22404 , n22405 , n22406 , n22407 , n22408 , n22409 , n22410 , n22411 , n22412 , n22413 , n22414 , n22415 , n22416 , n22417 , n22418 , n22419 , n22420 , n22421 , n22422 , n22423 , n22424 , n22425 , n22426 , n22427 , n22428 , n22429 , n22430 , n22431 , n22432 , n22433 , n22434 , n22435 , n22436 , n22437 , n22438 , n22439 , n22440 , n22441 , n22442 , n22443 , n22444 , n22445 , n22446 , n22447 , n22448 , n22449 , n22450 , n22451 , n22452 , n22453 , n22454 , n22455 , n22456 , n22457 , n22458 , n22459 , n22460 , n22461 , n22462 , n22463 , n22464 , n22465 , n22466 , n22467 , n22468 , n22469 , n22470 , n22471 , n22472 , n22473 , n22474 , n22475 , n22476 , n22477 , n22478 , n22479 , n22480 , n22481 , n22482 , n22483 , n22484 , n22485 , n22486 , n22487 , n22488 , n22489 , n22490 , n22491 , n22492 , n22493 , n22494 , n22495 , n22496 , n22497 , n22498 , n22499 , n22500 , n22501 , n22502 , n22503 , n22504 , n22505 , n22506 , n22507 , n22508 , n22509 , n22510 , n22511 , n22512 , n22513 , n22514 , n22515 , n22516 , n22517 , n22518 , n22519 , n22520 , n22521 , n22522 , n22523 , n22524 , n22525 , n22526 , n22527 , n22528 , n22529 , n22530 , n22531 , n22532 , n22533 , n22534 , n22535 , n22536 , n22537 , n22538 , n22539 , n22540 , n22541 , n22542 , n22543 , n22544 , n22545 , n22546 , n22547 , n22548 , n22549 , n22550 , n22551 , n22552 , n22553 , n22554 , n22555 , n22556 , n22557 , n22558 , n22559 , n22560 , n22561 , n22562 , n22563 , n22564 , n22565 , n22566 , n22567 , n22568 , n22569 , n22570 , n22571 , n22572 , n22573 , n22574 , n22575 , n22576 , n22577 , n22578 , n22579 , n22580 , n22581 , n22582 , n22583 , n22584 , n22585 , n22586 , n22587 , n22588 , n22589 , n22590 , n22591 , n22592 , n22593 , n22594 , n22595 , n22596 , n22597 , n22598 , n22599 , n22600 , n22601 , n22602 , n22603 , n22604 , n22605 , n22606 , n22607 , n22608 , n22609 , n22610 , n22611 , n22612 , n22613 , n22614 , n22615 , n22616 , n22617 , n22618 , n22619 , n22620 , n22621 , n22622 , n22623 , n22624 , n22625 , n22626 , n22627 , n22628 , n22629 , n22630 , n22631 , n22632 , n22633 , n22634 , n22635 , n22636 , n22637 , n22638 , n22639 , n22640 , n22641 , n22642 , n22643 , n22644 , n22645 , n22646 , n22647 , n22648 , n22649 , n22650 , n22651 , n22652 , n22653 , n22654 , n22655 , n22656 , n22657 , n22658 , n22659 , n22660 , n22661 , n22662 , n22663 , n22664 , n22665 , n22666 , n22667 , n22668 , n22669 , n22670 , n22671 , n22672 , n22673 , n22674 , n22675 , n22676 , n22677 , n22678 , n22679 , n22680 , n22681 , n22682 , n22683 , n22684 , n22685 , n22686 , n22687 , n22688 , n22689 , n22690 , n22691 , n22692 , n22693 , n22694 , n22695 , n22696 , n22697 , n22698 , n22699 , n22700 , n22701 , n22702 , n22703 , n22704 , n22705 , n22706 , n22707 , n22708 , n22709 , n22710 , n22711 , n22712 , n22713 , n22714 , n22715 , n22716 , n22717 , n22718 , n22719 , n22720 , n22721 , n22722 , n22723 , n22724 , n22725 , n22726 , n22727 , n22728 , n22729 , n22730 , n22731 , n22732 , n22733 , n22734 , n22735 , n22736 , n22737 , n22738 , n22739 , n22740 , n22741 , n22742 , n22743 , n22744 , n22745 , n22746 , n22747 , n22748 , n22749 , n22750 , n22751 , n22752 , n22753 , n22754 , n22755 , n22756 , n22757 , n22758 , n22759 , n22760 , n22761 , n22762 , n22763 , n22764 , n22765 , n22766 , n22767 , n22768 , n22769 , n22770 , n22771 , n22772 , n22773 , n22774 , n22775 , n22776 , n22777 , n22778 , n22779 , n22780 , n22781 , n22782 , n22783 , n22784 , n22785 , n22786 , n22787 , n22788 , n22789 , n22790 , n22791 , n22792 , n22793 , n22794 , n22795 , n22796 , n22797 , n22798 , n22799 , n22800 , n22801 , n22802 , n22803 , n22804 , n22805 , n22806 , n22807 , n22808 , n22809 , n22810 , n22811 , n22812 , n22813 , n22814 , n22815 , n22816 , n22817 , n22818 , n22819 , n22820 , n22821 , n22822 , n22823 , n22824 , n22825 , n22826 , n22827 , n22828 , n22829 , n22830 , n22831 , n22832 , n22833 , n22834 , n22835 , n22836 , n22837 , n22838 , n22839 , n22840 , n22841 , n22842 , n22843 , n22844 , n22845 , n22846 , n22847 , n22848 , n22849 , n22850 , n22851 , n22852 , n22853 , n22854 , n22855 , n22856 , n22857 , n22858 , n22859 , n22860 , n22861 , n22862 , n22863 , n22864 , n22865 , n22866 , n22867 , n22868 , n22869 , n22870 , n22871 , n22872 , n22873 , n22874 , n22875 , n22876 , n22877 , n22878 , n22879 , n22880 , n22881 , n22882 , n22883 , n22884 , n22885 , n22886 , n22887 , n22888 , n22889 , n22890 , n22891 , n22892 , n22893 , n22894 , n22895 , n22896 , n22897 , n22898 , n22899 , n22900 , n22901 , n22902 , n22903 , n22904 , n22905 , n22906 , n22907 , n22908 , n22909 , n22910 , n22911 , n22912 , n22913 , n22914 , n22915 , n22916 , n22917 , n22918 , n22919 , n22920 , n22921 , n22922 , n22923 , n22924 , n22925 , n22926 , n22927 , n22928 , n22929 , n22930 , n22931 , n22932 , n22933 , n22934 , n22935 , n22936 , n22937 , n22938 , n22939 , n22940 , n22941 , n22942 , n22943 , n22944 , n22945 , n22946 , n22947 , n22948 , n22949 , n22950 , n22951 , n22952 , n22953 , n22954 , n22955 , n22956 , n22957 , n22958 , n22959 , n22960 , n22961 , n22962 , n22963 , n22964 , n22965 , n22966 , n22967 , n22968 , n22969 , n22970 , n22971 , n22972 , n22973 , n22974 , n22975 , n22976 , n22977 , n22978 , n22979 , n22980 , n22981 , n22982 , n22983 , n22984 , n22985 , n22986 , n22987 , n22988 , n22989 , n22990 , n22991 , n22992 , n22993 , n22994 , n22995 , n22996 , n22997 , n22998 , n22999 , n23000 , n23001 , n23002 , n23003 , n23004 , n23005 , n23006 , n23007 , n23008 , n23009 , n23010 , n23011 , n23012 , n23013 , n23014 , n23015 , n23016 , n23017 , n23018 , n23019 , n23020 , n23021 , n23022 , n23023 , n23024 , n23025 , n23026 , n23027 , n23028 , n23029 , n23030 , n23031 , n23032 , n23033 , n23034 , n23035 , n23036 , n23037 , n23038 , n23039 , n23040 , n23041 , n23042 , n23043 , n23044 , n23045 , n23046 , n23047 , n23048 , n23049 , n23050 , n23051 , n23052 , n23053 , n23054 , n23055 , n23056 , n23057 , n23058 , n23059 , n23060 , n23061 , n23062 , n23063 , n23064 , n23065 , n23066 , n23067 , n23068 , n23069 , n23070 , n23071 , n23072 , n23073 , n23074 , n23075 , n23076 , n23077 , n23078 , n23079 , n23080 , n23081 , n23082 , n23083 , n23084 , n23085 , n23086 , n23087 , n23088 , n23089 , n23090 , n23091 , n23092 , n23093 , n23094 , n23095 , n23096 , n23097 , n23098 , n23099 , n23100 , n23101 , n23102 , n23103 , n23104 , n23105 , n23106 , n23107 , n23108 , n23109 , n23110 , n23111 , n23112 , n23113 , n23114 , n23115 , n23116 , n23117 , n23118 , n23119 , n23120 , n23121 , n23122 , n23123 , n23124 , n23125 , n23126 , n23127 , n23128 , n23129 , n23130 , n23131 , n23132 , n23133 , n23134 , n23135 , n23136 , n23137 , n23138 , n23139 , n23140 , n23141 , n23142 , n23143 , n23144 , n23145 , n23146 , n23147 , n23148 , n23149 , n23150 , n23151 , n23152 , n23153 , n23154 , n23155 , n23156 , n23157 , n23158 , n23159 , n23160 , n23161 , n23162 , n23163 , n23164 , n23165 , n23166 , n23167 , n23168 , n23169 , n23170 , n23171 , n23172 , n23173 , n23174 , n23175 , n23176 , n23177 , n23178 , n23179 , n23180 , n23181 , n23182 , n23183 , n23184 , n23185 , n23186 , n23187 , n23188 , n23189 , n23190 , n23191 , n23192 , n23193 , n23194 , n23195 , n23196 , n23197 , n23198 , n23199 , n23200 , n23201 , n23202 , n23203 , n23204 , n23205 , n23206 , n23207 , n23208 , n23209 , n23210 , n23211 , n23212 , n23213 , n23214 , n23215 , n23216 , n23217 , n23218 , n23219 , n23220 , n23221 , n23222 , n23223 , n23224 , n23225 , n23226 , n23227 , n23228 , n23229 , n23230 , n23231 , n23232 , n23233 , n23234 , n23235 , n23236 , n23237 , n23238 , n23239 , n23240 , n23241 , n23242 , n23243 , n23244 , n23245 , n23246 , n23247 , n23248 , n23249 , n23250 , n23251 , n23252 , n23253 , n23254 , n23255 , n23256 , n23257 , n23258 , n23259 , n23260 , n23261 , n23262 , n23263 , n23264 , n23265 , n23266 , n23267 , n23268 , n23269 , n23270 , n23271 , n23272 , n23273 , n23274 , n23275 , n23276 , n23277 , n23278 , n23279 , n23280 , n23281 , n23282 , n23283 , n23284 , n23285 , n23286 , n23287 , n23288 , n23289 , n23290 , n23291 , n23292 , n23293 , n23294 , n23295 , n23296 , n23297 , n23298 , n23299 , n23300 , n23301 , n23302 , n23303 , n23304 , n23305 , n23306 , n23307 , n23308 , n23309 , n23310 , n23311 , n23312 , n23313 , n23314 , n23315 , n23316 , n23317 , n23318 , n23319 , n23320 , n23321 , n23322 , n23323 , n23324 , n23325 , n23326 , n23327 , n23328 , n23329 , n23330 , n23331 , n23332 , n23333 , n23334 , n23335 , n23336 , n23337 , n23338 , n23339 , n23340 , n23341 , n23342 , n23343 , n23344 , n23345 , n23346 , n23347 , n23348 , n23349 , n23350 , n23351 , n23352 , n23353 , n23354 , n23355 , n23356 , n23357 , n23358 , n23359 , n23360 , n23361 , n23362 , n23363 , n23364 , n23365 , n23366 , n23367 , n23368 , n23369 , n23370 , n23371 , n23372 , n23373 , n23374 , n23375 , n23376 , n23377 , n23378 , n23379 , n23380 , n23381 , n23382 , n23383 , n23384 , n23385 , n23386 , n23387 , n23388 , n23389 , n23390 , n23391 , n23392 , n23393 , n23394 , n23395 , n23396 , n23397 , n23398 , n23399 , n23400 , n23401 , n23402 , n23403 , n23404 , n23405 , n23406 , n23407 , n23408 , n23409 , n23410 , n23411 , n23412 , n23413 , n23414 , n23415 , n23416 , n23417 , n23418 , n23419 , n23420 , n23421 , n23422 , n23423 , n23424 , n23425 , n23426 , n23427 , n23428 , n23429 , n23430 , n23431 , n23432 , n23433 , n23434 , n23435 , n23436 , n23437 , n23438 , n23439 , n23440 , n23441 , n23442 , n23443 , n23444 , n23445 , n23446 , n23447 , n23448 , n23449 , n23450 , n23451 , n23452 , n23453 , n23454 , n23455 , n23456 , n23457 , n23458 , n23459 , n23460 , n23461 , n23462 , n23463 , n23464 , n23465 , n23466 , n23467 , n23468 , n23469 , n23470 , n23471 , n23472 , n23473 , n23474 , n23475 , n23476 , n23477 , n23478 , n23479 , n23480 , n23481 , n23482 , n23483 , n23484 , n23485 , n23486 , n23487 , n23488 , n23489 , n23490 , n23491 , n23492 , n23493 , n23494 , n23495 , n23496 , n23497 , n23498 , n23499 , n23500 , n23501 , n23502 , n23503 , n23504 , n23505 , n23506 , n23507 , n23508 , n23509 , n23510 , n23511 , n23512 , n23513 , n23514 , n23515 , n23516 , n23517 , n23518 , n23519 , n23520 , n23521 , n23522 , n23523 , n23524 , n23525 , n23526 , n23527 , n23528 , n23529 , n23530 , n23531 , n23532 , n23533 , n23534 , n23535 , n23536 , n23537 , n23538 , n23539 , n23540 , n23541 , n23542 , n23543 , n23544 , n23545 , n23546 , n23547 , n23548 , n23549 , n23550 , n23551 , n23552 , n23553 , n23554 , n23555 , n23556 , n23557 , n23558 , n23559 , n23560 , n23561 , n23562 , n23563 , n23564 , n23565 , n23566 , n23567 , n23568 , n23569 , n23570 , n23571 , n23572 , n23573 , n23574 , n23575 , n23576 , n23577 , n23578 , n23579 , n23580 , n23581 , n23582 , n23583 , n23584 , n23585 , n23586 , n23587 , n23588 , n23589 , n23590 , n23591 , n23592 , n23593 , n23594 , n23595 , n23596 , n23597 , n23598 , n23599 , n23600 , n23601 , n23602 , n23603 , n23604 , n23605 , n23606 , n23607 , n23608 , n23609 , n23610 , n23611 , n23612 , n23613 , n23614 , n23615 , n23616 , n23617 , n23618 , n23619 , n23620 , n23621 , n23622 , n23623 , n23624 , n23625 , n23626 , n23627 , n23628 , n23629 , n23630 , n23631 , n23632 , n23633 , n23634 , n23635 , n23636 , n23637 , n23638 , n23639 , n23640 , n23641 , n23642 , n23643 , n23644 , n23645 , n23646 , n23647 , n23648 , n23649 , n23650 , n23651 , n23652 , n23653 , n23654 , n23655 , n23656 , n23657 , n23658 , n23659 , n23660 , n23661 , n23662 , n23663 , n23664 , n23665 , n23666 , n23667 , n23668 , n23669 , n23670 , n23671 , n23672 , n23673 , n23674 , n23675 , n23676 , n23677 , n23678 , n23679 , n23680 , n23681 , n23682 , n23683 , n23684 , n23685 , n23686 , n23687 , n23688 , n23689 , n23690 , n23691 , n23692 , n23693 , n23694 , n23695 , n23696 , n23697 , n23698 , n23699 , n23700 , n23701 , n23702 , n23703 , n23704 , n23705 , n23706 , n23707 , n23708 , n23709 , n23710 , n23711 , n23712 , n23713 , n23714 , n23715 , n23716 , n23717 , n23718 , n23719 , n23720 , n23721 , n23722 , n23723 , n23724 , n23725 , n23726 , n23727 , n23728 , n23729 , n23730 , n23731 , n23732 , n23733 , n23734 , n23735 , n23736 , n23737 , n23738 , n23739 , n23740 , n23741 , n23742 , n23743 , n23744 , n23745 , n23746 , n23747 , n23748 , n23749 , n23750 , n23751 , n23752 , n23753 , n23754 , n23755 , n23756 , n23757 , n23758 , n23759 , n23760 , n23761 , n23762 , n23763 , n23764 , n23765 , n23766 , n23767 , n23768 , n23769 , n23770 , n23771 , n23772 , n23773 , n23774 , n23775 , n23776 , n23777 , n23778 , n23779 , n23780 , n23781 , n23782 , n23783 , n23784 , n23785 , n23786 , n23787 , n23788 , n23789 , n23790 , n23791 , n23792 , n23793 , n23794 , n23795 , n23796 , n23797 , n23798 , n23799 , n23800 , n23801 , n23802 , n23803 , n23804 , n23805 , n23806 , n23807 , n23808 , n23809 , n23810 , n23811 , n23812 , n23813 , n23814 , n23815 , n23816 , n23817 , n23818 , n23819 , n23820 , n23821 , n23822 , n23823 , n23824 , n23825 , n23826 , n23827 , n23828 , n23829 , n23830 , n23831 , n23832 , n23833 , n23834 , n23835 , n23836 , n23837 , n23838 , n23839 , n23840 , n23841 , n23842 , n23843 , n23844 , n23845 , n23846 , n23847 , n23848 , n23849 , n23850 , n23851 , n23852 , n23853 , n23854 , n23855 , n23856 , n23857 , n23858 , n23859 , n23860 , n23861 , n23862 , n23863 , n23864 , n23865 , n23866 , n23867 , n23868 , n23869 , n23870 , n23871 , n23872 , n23873 , n23874 , n23875 , n23876 , n23877 , n23878 , n23879 , n23880 , n23881 , n23882 , n23883 , n23884 , n23885 , n23886 , n23887 , n23888 , n23889 , n23890 , n23891 , n23892 , n23893 , n23894 , n23895 , n23896 , n23897 , n23898 , n23899 , n23900 , n23901 , n23902 , n23903 , n23904 , n23905 , n23906 , n23907 , n23908 , n23909 , n23910 , n23911 , n23912 , n23913 , n23914 , n23915 , n23916 , n23917 , n23918 , n23919 , n23920 , n23921 , n23922 , n23923 , n23924 , n23925 , n23926 , n23927 , n23928 , n23929 , n23930 , n23931 , n23932 , n23933 , n23934 , n23935 , n23936 , n23937 , n23938 , n23939 , n23940 , n23941 , n23942 , n23943 , n23944 , n23945 , n23946 , n23947 , n23948 , n23949 , n23950 , n23951 , n23952 , n23953 , n23954 , n23955 , n23956 , n23957 , n23958 , n23959 , n23960 , n23961 , n23962 , n23963 , n23964 , n23965 , n23966 , n23967 , n23968 , n23969 , n23970 , n23971 , n23972 , n23973 , n23974 , n23975 , n23976 , n23977 , n23978 , n23979 , n23980 , n23981 , n23982 , n23983 , n23984 , n23985 , n23986 , n23987 , n23988 , n23989 , n23990 , n23991 , n23992 , n23993 , n23994 , n23995 , n23996 , n23997 , n23998 , n23999 , n24000 , n24001 , n24002 , n24003 , n24004 , n24005 , n24006 , n24007 , n24008 , n24009 , n24010 , n24011 , n24012 , n24013 , n24014 , n24015 , n24016 , n24017 , n24018 , n24019 , n24020 , n24021 , n24022 , n24023 , n24024 , n24025 , n24026 , n24027 , n24028 , n24029 , n24030 , n24031 , n24032 , n24033 , n24034 , n24035 , n24036 , n24037 , n24038 , n24039 , n24040 , n24041 , n24042 , n24043 , n24044 , n24045 , n24046 , n24047 , n24048 , n24049 , n24050 , n24051 , n24052 , n24053 , n24054 , n24055 , n24056 , n24057 , n24058 , n24059 , n24060 , n24061 , n24062 , n24063 , n24064 , n24065 , n24066 , n24067 , n24068 , n24069 , n24070 , n24071 , n24072 , n24073 , n24074 , n24075 , n24076 , n24077 , n24078 , n24079 , n24080 , n24081 , n24082 , n24083 , n24084 , n24085 , n24086 , n24087 , n24088 , n24089 , n24090 , n24091 , n24092 , n24093 , n24094 , n24095 , n24096 , n24097 , n24098 , n24099 , n24100 , n24101 , n24102 , n24103 , n24104 , n24105 , n24106 , n24107 , n24108 , n24109 , n24110 , n24111 , n24112 , n24113 , n24114 , n24115 , n24116 , n24117 , n24118 , n24119 , n24120 , n24121 , n24122 , n24123 , n24124 , n24125 , n24126 , n24127 , n24128 , n24129 , n24130 , n24131 , n24132 , n24133 , n24134 , n24135 , n24136 , n24137 , n24138 , n24139 , n24140 , n24141 , n24142 , n24143 , n24144 , n24145 , n24146 , n24147 , n24148 , n24149 , n24150 , n24151 , n24152 , n24153 , n24154 , n24155 , n24156 , n24157 , n24158 , n24159 , n24160 , n24161 , n24162 , n24163 , n24164 , n24165 , n24166 , n24167 , n24168 , n24169 , n24170 , n24171 , n24172 , n24173 , n24174 , n24175 , n24176 , n24177 , n24178 , n24179 , n24180 , n24181 , n24182 , n24183 , n24184 , n24185 , n24186 , n24187 , n24188 , n24189 , n24190 , n24191 , n24192 , n24193 , n24194 , n24195 , n24196 , n24197 , n24198 , n24199 , n24200 , n24201 , n24202 , n24203 , n24204 , n24205 , n24206 , n24207 , n24208 , n24209 , n24210 , n24211 , n24212 , n24213 , n24214 , n24215 , n24216 , n24217 , n24218 , n24219 , n24220 , n24221 , n24222 , n24223 , n24224 , n24225 , n24226 , n24227 , n24228 , n24229 , n24230 , n24231 , n24232 , n24233 , n24234 , n24235 , n24236 , n24237 , n24238 , n24239 , n24240 , n24241 , n24242 , n24243 , n24244 , n24245 , n24246 , n24247 , n24248 , n24249 , n24250 , n24251 , n24252 , n24253 , n24254 , n24255 , n24256 , n24257 , n24258 , n24259 , n24260 , n24261 , n24262 , n24263 , n24264 , n24265 , n24266 , n24267 , n24268 , n24269 , n24270 , n24271 , n24272 , n24273 , n24274 , n24275 , n24276 , n24277 , n24278 , n24279 , n24280 , n24281 , n24282 , n24283 , n24284 , n24285 , n24286 , n24287 , n24288 , n24289 , n24290 , n24291 , n24292 , n24293 , n24294 , n24295 , n24296 , n24297 , n24298 , n24299 , n24300 , n24301 , n24302 , n24303 , n24304 , n24305 , n24306 , n24307 , n24308 , n24309 , n24310 , n24311 , n24312 , n24313 , n24314 , n24315 , n24316 , n24317 , n24318 , n24319 , n24320 , n24321 , n24322 , n24323 , n24324 , n24325 , n24326 , n24327 , n24328 , n24329 , n24330 , n24331 , n24332 , n24333 , n24334 , n24335 , n24336 , n24337 , n24338 , n24339 , n24340 , n24341 , n24342 , n24343 , n24344 , n24345 , n24346 , n24347 , n24348 , n24349 , n24350 , n24351 , n24352 , n24353 , n24354 , n24355 , n24356 , n24357 , n24358 , n24359 , n24360 , n24361 , n24362 , n24363 , n24364 , n24365 , n24366 , n24367 , n24368 , n24369 , n24370 , n24371 , n24372 , n24373 , n24374 , n24375 , n24376 , n24377 , n24378 , n24379 , n24380 , n24381 , n24382 , n24383 , n24384 , n24385 , n24386 , n24387 , n24388 , n24389 , n24390 , n24391 , n24392 , n24393 , n24394 , n24395 , n24396 , n24397 , n24398 , n24399 , n24400 , n24401 , n24402 , n24403 , n24404 , n24405 , n24406 , n24407 , n24408 , n24409 , n24410 , n24411 , n24412 , n24413 , n24414 , n24415 , n24416 , n24417 , n24418 , n24419 , n24420 , n24421 , n24422 , n24423 , n24424 , n24425 , n24426 , n24427 , n24428 , n24429 , n24430 , n24431 , n24432 , n24433 , n24434 , n24435 , n24436 , n24437 , n24438 , n24439 , n24440 , n24441 , n24442 , n24443 , n24444 , n24445 , n24446 , n24447 , n24448 , n24449 , n24450 , n24451 , n24452 , n24453 , n24454 , n24455 , n24456 , n24457 , n24458 , n24459 , n24460 , n24461 , n24462 , n24463 , n24464 , n24465 , n24466 , n24467 , n24468 , n24469 , n24470 , n24471 , n24472 , n24473 , n24474 , n24475 , n24476 , n24477 , n24478 , n24479 , n24480 , n24481 , n24482 , n24483 , n24484 , n24485 , n24486 , n24487 , n24488 , n24489 , n24490 , n24491 , n24492 , n24493 , n24494 , n24495 , n24496 , n24497 , n24498 , n24499 , n24500 , n24501 , n24502 , n24503 , n24504 , n24505 , n24506 , n24507 , n24508 , n24509 , n24510 , n24511 , n24512 , n24513 , n24514 , n24515 , n24516 , n24517 , n24518 , n24519 , n24520 , n24521 , n24522 , n24523 , n24524 , n24525 , n24526 , n24527 , n24528 , n24529 , n24530 , n24531 , n24532 , n24533 , n24534 , n24535 , n24536 , n24537 , n24538 , n24539 , n24540 , n24541 , n24542 , n24543 , n24544 , n24545 , n24546 , n24547 , n24548 , n24549 , n24550 , n24551 , n24552 , n24553 , n24554 , n24555 , n24556 , n24557 , n24558 , n24559 , n24560 , n24561 , n24562 , n24563 , n24564 , n24565 , n24566 , n24567 , n24568 , n24569 , n24570 , n24571 , n24572 , n24573 , n24574 , n24575 , n24576 , n24577 , n24578 , n24579 , n24580 , n24581 , n24582 , n24583 , n24584 , n24585 , n24586 , n24587 , n24588 , n24589 , n24590 , n24591 , n24592 , n24593 , n24594 , n24595 , n24596 , n24597 , n24598 , n24599 , n24600 , n24601 , n24602 , n24603 , n24604 , n24605 , n24606 , n24607 , n24608 , n24609 , n24610 , n24611 , n24612 , n24613 , n24614 , n24615 , n24616 , n24617 , n24618 , n24619 , n24620 , n24621 , n24622 , n24623 , n24624 , n24625 , n24626 , n24627 , n24628 , n24629 , n24630 , n24631 , n24632 , n24633 , n24634 , n24635 , n24636 , n24637 , n24638 , n24639 , n24640 , n24641 , n24642 , n24643 , n24644 , n24645 , n24646 , n24647 , n24648 , n24649 , n24650 , n24651 , n24652 , n24653 , n24654 , n24655 , n24656 , n24657 , n24658 , n24659 , n24660 , n24661 , n24662 , n24663 , n24664 , n24665 , n24666 , n24667 , n24668 , n24669 , n24670 , n24671 , n24672 , n24673 , n24674 , n24675 , n24676 , n24677 , n24678 , n24679 , n24680 , n24681 , n24682 , n24683 , n24684 , n24685 , n24686 , n24687 , n24688 , n24689 , n24690 , n24691 , n24692 , n24693 , n24694 , n24695 , n24696 , n24697 , n24698 , n24699 , n24700 , n24701 , n24702 , n24703 , n24704 , n24705 , n24706 , n24707 , n24708 , n24709 , n24710 , n24711 , n24712 , n24713 , n24714 , n24715 , n24716 , n24717 , n24718 , n24719 , n24720 , n24721 , n24722 , n24723 , n24724 , n24725 , n24726 , n24727 , n24728 , n24729 , n24730 , n24731 , n24732 , n24733 , n24734 , n24735 , n24736 , n24737 , n24738 , n24739 , n24740 , n24741 , n24742 , n24743 , n24744 , n24745 , n24746 , n24747 , n24748 , n24749 , n24750 , n24751 , n24752 , n24753 , n24754 , n24755 , n24756 , n24757 , n24758 , n24759 , n24760 , n24761 , n24762 , n24763 , n24764 , n24765 , n24766 , n24767 , n24768 , n24769 , n24770 , n24771 , n24772 , n24773 , n24774 , n24775 , n24776 , n24777 , n24778 , n24779 , n24780 , n24781 , n24782 , n24783 , n24784 , n24785 , n24786 , n24787 , n24788 , n24789 , n24790 , n24791 , n24792 , n24793 , n24794 , n24795 , n24796 , n24797 , n24798 , n24799 , n24800 , n24801 , n24802 , n24803 , n24804 , n24805 , n24806 , n24807 , n24808 , n24809 , n24810 , n24811 , n24812 , n24813 , n24814 , n24815 , n24816 , n24817 , n24818 , n24819 , n24820 , n24821 , n24822 , n24823 , n24824 , n24825 , n24826 , n24827 , n24828 , n24829 , n24830 , n24831 , n24832 , n24833 , n24834 , n24835 , n24836 , n24837 , n24838 , n24839 , n24840 , n24841 , n24842 , n24843 , n24844 , n24845 , n24846 , n24847 , n24848 , n24849 , n24850 , n24851 , n24852 , n24853 , n24854 , n24855 , n24856 , n24857 , n24858 , n24859 , n24860 , n24861 , n24862 , n24863 , n24864 , n24865 , n24866 , n24867 , n24868 , n24869 , n24870 , n24871 , n24872 , n24873 , n24874 , n24875 , n24876 , n24877 , n24878 , n24879 , n24880 , n24881 , n24882 , n24883 , n24884 , n24885 , n24886 , n24887 , n24888 , n24889 , n24890 , n24891 , n24892 , n24893 , n24894 , n24895 , n24896 , n24897 , n24898 , n24899 , n24900 , n24901 , n24902 , n24903 , n24904 , n24905 , n24906 , n24907 , n24908 , n24909 , n24910 , n24911 , n24912 , n24913 , n24914 , n24915 , n24916 , n24917 , n24918 , n24919 , n24920 , n24921 , n24922 , n24923 , n24924 , n24925 , n24926 , n24927 , n24928 , n24929 , n24930 , n24931 , n24932 , n24933 , n24934 , n24935 , n24936 , n24937 , n24938 , n24939 , n24940 , n24941 , n24942 , n24943 , n24944 , n24945 , n24946 , n24947 , n24948 , n24949 , n24950 , n24951 , n24952 , n24953 , n24954 , n24955 , n24956 , n24957 , n24958 , n24959 , n24960 , n24961 , n24962 , n24963 , n24964 , n24965 , n24966 , n24967 , n24968 , n24969 , n24970 , n24971 , n24972 , n24973 , n24974 , n24975 , n24976 , n24977 , n24978 , n24979 , n24980 , n24981 , n24982 , n24983 , n24984 , n24985 , n24986 , n24987 , n24988 , n24989 , n24990 , n24991 , n24992 , n24993 , n24994 , n24995 , n24996 , n24997 , n24998 , n24999 , n25000 , n25001 , n25002 , n25003 , n25004 , n25005 , n25006 , n25007 , n25008 , n25009 , n25010 , n25011 , n25012 , n25013 , n25014 , n25015 , n25016 , n25017 , n25018 , n25019 , n25020 , n25021 , n25022 , n25023 , n25024 , n25025 , n25026 , n25027 , n25028 , n25029 , n25030 , n25031 , n25032 , n25033 , n25034 , n25035 , n25036 , n25037 , n25038 , n25039 , n25040 , n25041 , n25042 , n25043 , n25044 , n25045 , n25046 , n25047 , n25048 , n25049 , n25050 , n25051 , n25052 , n25053 , n25054 , n25055 , n25056 , n25057 , n25058 , n25059 , n25060 , n25061 , n25062 , n25063 , n25064 , n25065 , n25066 , n25067 , n25068 , n25069 , n25070 , n25071 , n25072 , n25073 , n25074 , n25075 , n25076 , n25077 , n25078 , n25079 , n25080 , n25081 , n25082 , n25083 , n25084 , n25085 , n25086 , n25087 , n25088 , n25089 , n25090 , n25091 , n25092 , n25093 , n25094 , n25095 , n25096 , n25097 , n25098 , n25099 , n25100 , n25101 , n25102 , n25103 , n25104 , n25105 , n25106 , n25107 , n25108 , n25109 , n25110 , n25111 , n25112 , n25113 , n25114 , n25115 , n25116 , n25117 , n25118 , n25119 , n25120 , n25121 , n25122 , n25123 , n25124 , n25125 , n25126 , n25127 , n25128 , n25129 , n25130 , n25131 , n25132 , n25133 , n25134 , n25135 , n25136 , n25137 , n25138 , n25139 , n25140 , n25141 , n25142 , n25143 , n25144 , n25145 , n25146 , n25147 , n25148 , n25149 , n25150 , n25151 , n25152 , n25153 , n25154 , n25155 , n25156 , n25157 , n25158 , n25159 , n25160 , n25161 , n25162 , n25163 , n25164 , n25165 , n25166 , n25167 , n25168 , n25169 , n25170 , n25171 , n25172 , n25173 , n25174 , n25175 , n25176 , n25177 , n25178 , n25179 , n25180 , n25181 , n25182 , n25183 , n25184 , n25185 , n25186 , n25187 , n25188 , n25189 , n25190 , n25191 , n25192 , n25193 , n25194 , n25195 , n25196 , n25197 , n25198 , n25199 , n25200 , n25201 , n25202 , n25203 , n25204 , n25205 , n25206 , n25207 , n25208 , n25209 , n25210 , n25211 , n25212 , n25213 , n25214 , n25215 , n25216 , n25217 , n25218 , n25219 , n25220 , n25221 , n25222 , n25223 , n25224 , n25225 , n25226 , n25227 , n25228 , n25229 , n25230 , n25231 , n25232 , n25233 , n25234 , n25235 , n25236 , n25237 , n25238 , n25239 , n25240 , n25241 , n25242 , n25243 , n25244 , n25245 , n25246 , n25247 , n25248 , n25249 , n25250 , n25251 , n25252 , n25253 , n25254 , n25255 , n25256 , n25257 , n25258 , n25259 , n25260 , n25261 , n25262 , n25263 , n25264 , n25265 , n25266 , n25267 , n25268 , n25269 , n25270 , n25271 , n25272 , n25273 , n25274 , n25275 , n25276 , n25277 , n25278 , n25279 , n25280 , n25281 , n25282 , n25283 , n25284 , n25285 , n25286 , n25287 , n25288 , n25289 , n25290 , n25291 , n25292 , n25293 , n25294 , n25295 , n25296 , n25297 , n25298 , n25299 , n25300 , n25301 , n25302 , n25303 , n25304 , n25305 , n25306 , n25307 , n25308 , n25309 , n25310 , n25311 , n25312 , n25313 , n25314 , n25315 , n25316 , n25317 , n25318 , n25319 , n25320 , n25321 , n25322 , n25323 , n25324 , n25325 , n25326 , n25327 , n25328 , n25329 , n25330 , n25331 , n25332 , n25333 , n25334 , n25335 , n25336 , n25337 , n25338 , n25339 , n25340 , n25341 , n25342 , n25343 , n25344 , n25345 , n25346 , n25347 , n25348 , n25349 , n25350 , n25351 , n25352 , n25353 , n25354 , n25355 , n25356 , n25357 , n25358 , n25359 , n25360 , n25361 , n25362 , n25363 , n25364 , n25365 , n25366 , n25367 , n25368 , n25369 , n25370 , n25371 , n25372 , n25373 , n25374 , n25375 , n25376 , n25377 , n25378 , n25379 , n25380 , n25381 , n25382 , n25383 , n25384 , n25385 , n25386 , n25387 , n25388 , n25389 , n25390 , n25391 , n25392 , n25393 , n25394 , n25395 , n25396 , n25397 , n25398 , n25399 , n25400 , n25401 , n25402 , n25403 , n25404 , n25405 , n25406 , n25407 , n25408 , n25409 , n25410 , n25411 , n25412 , n25413 , n25414 , n25415 , n25416 , n25417 , n25418 , n25419 , n25420 , n25421 , n25422 , n25423 , n25424 , n25425 , n25426 , n25427 , n25428 , n25429 , n25430 , n25431 , n25432 , n25433 , n25434 , n25435 , n25436 , n25437 , n25438 , n25439 , n25440 , n25441 , n25442 , n25443 , n25444 , n25445 , n25446 , n25447 , n25448 , n25449 , n25450 , n25451 , n25452 , n25453 , n25454 , n25455 , n25456 , n25457 , n25458 , n25459 , n25460 , n25461 , n25462 , n25463 , n25464 , n25465 , n25466 , n25467 , n25468 , n25469 , n25470 , n25471 , n25472 , n25473 , n25474 , n25475 , n25476 , n25477 , n25478 , n25479 , n25480 , n25481 , n25482 , n25483 , n25484 , n25485 , n25486 , n25487 , n25488 , n25489 , n25490 , n25491 , n25492 , n25493 , n25494 , n25495 , n25496 , n25497 , n25498 , n25499 , n25500 , n25501 , n25502 , n25503 , n25504 , n25505 , n25506 , n25507 , n25508 , n25509 , n25510 , n25511 , n25512 , n25513 , n25514 , n25515 , n25516 , n25517 , n25518 , n25519 , n25520 , n25521 , n25522 , n25523 , n25524 , n25525 , n25526 , n25527 , n25528 , n25529 , n25530 , n25531 , n25532 , n25533 , n25534 , n25535 , n25536 , n25537 , n25538 , n25539 , n25540 , n25541 , n25542 , n25543 , n25544 , n25545 , n25546 , n25547 , n25548 , n25549 , n25550 , n25551 , n25552 , n25553 , n25554 , n25555 , n25556 , n25557 , n25558 , n25559 , n25560 , n25561 , n25562 , n25563 , n25564 , n25565 , n25566 , n25567 , n25568 , n25569 , n25570 , n25571 , n25572 , n25573 , n25574 , n25575 , n25576 , n25577 , n25578 , n25579 , n25580 , n25581 , n25582 , n25583 , n25584 , n25585 , n25586 , n25587 , n25588 , n25589 , n25590 , n25591 , n25592 , n25593 , n25594 , n25595 , n25596 , n25597 , n25598 , n25599 , n25600 , n25601 , n25602 , n25603 , n25604 , n25605 , n25606 , n25607 , n25608 , n25609 , n25610 , n25611 , n25612 , n25613 , n25614 , n25615 , n25616 , n25617 , n25618 , n25619 , n25620 , n25621 , n25622 , n25623 , n25624 , n25625 , n25626 , n25627 , n25628 , n25629 , n25630 , n25631 , n25632 , n25633 , n25634 , n25635 , n25636 , n25637 , n25638 , n25639 , n25640 , n25641 , n25642 , n25643 , n25644 , n25645 , n25646 , n25647 , n25648 , n25649 , n25650 , n25651 , n25652 , n25653 , n25654 , n25655 , n25656 , n25657 , n25658 , n25659 , n25660 , n25661 , n25662 , n25663 , n25664 , n25665 , n25666 , n25667 , n25668 , n25669 , n25670 , n25671 , n25672 , n25673 , n25674 , n25675 , n25676 , n25677 , n25678 , n25679 , n25680 , n25681 , n25682 , n25683 , n25684 , n25685 , n25686 , n25687 , n25688 , n25689 , n25690 , n25691 , n25692 , n25693 , n25694 , n25695 , n25696 , n25697 , n25698 , n25699 , n25700 , n25701 , n25702 , n25703 , n25704 , n25705 , n25706 , n25707 , n25708 , n25709 , n25710 , n25711 , n25712 , n25713 , n25714 , n25715 , n25716 , n25717 , n25718 , n25719 , n25720 , n25721 , n25722 , n25723 , n25724 , n25725 , n25726 , n25727 , n25728 , n25729 , n25730 , n25731 , n25732 , n25733 , n25734 , n25735 , n25736 , n25737 , n25738 , n25739 , n25740 , n25741 , n25742 , n25743 , n25744 , n25745 , n25746 , n25747 , n25748 , n25749 , n25750 , n25751 , n25752 , n25753 , n25754 , n25755 , n25756 , n25757 , n25758 , n25759 , n25760 , n25761 , n25762 , n25763 , n25764 , n25765 , n25766 , n25767 , n25768 , n25769 , n25770 , n25771 , n25772 , n25773 , n25774 , n25775 , n25776 , n25777 , n25778 , n25779 , n25780 , n25781 , n25782 , n25783 , n25784 , n25785 , n25786 , n25787 , n25788 , n25789 , n25790 , n25791 , n25792 , n25793 , n25794 , n25795 , n25796 , n25797 , n25798 , n25799 , n25800 , n25801 , n25802 , n25803 , n25804 , n25805 , n25806 , n25807 , n25808 , n25809 , n25810 , n25811 , n25812 , n25813 , n25814 , n25815 , n25816 , n25817 , n25818 , n25819 , n25820 , n25821 , n25822 , n25823 , n25824 , n25825 , n25826 , n25827 , n25828 , n25829 , n25830 , n25831 , n25832 , n25833 , n25834 , n25835 , n25836 , n25837 , n25838 , n25839 , n25840 , n25841 , n25842 , n25843 , n25844 , n25845 , n25846 , n25847 , n25848 , n25849 , n25850 , n25851 , n25852 , n25853 , n25854 , n25855 , n25856 , n25857 , n25858 , n25859 , n25860 , n25861 , n25862 , n25863 , n25864 , n25865 , n25866 , n25867 , n25868 , n25869 , n25870 , n25871 , n25872 , n25873 , n25874 , n25875 , n25876 , n25877 , n25878 , n25879 , n25880 , n25881 , n25882 , n25883 , n25884 , n25885 , n25886 , n25887 , n25888 , n25889 , n25890 , n25891 , n25892 , n25893 , n25894 , n25895 , n25896 , n25897 , n25898 , n25899 , n25900 , n25901 , n25902 , n25903 , n25904 , n25905 , n25906 , n25907 , n25908 , n25909 , n25910 , n25911 , n25912 , n25913 , n25914 , n25915 , n25916 , n25917 , n25918 , n25919 , n25920 , n25921 , n25922 , n25923 , n25924 , n25925 , n25926 , n25927 , n25928 , n25929 , n25930 , n25931 , n25932 , n25933 , n25934 , n25935 , n25936 , n25937 , n25938 , n25939 , n25940 , n25941 , n25942 , n25943 , n25944 , n25945 , n25946 , n25947 , n25948 , n25949 , n25950 , n25951 , n25952 , n25953 , n25954 , n25955 , n25956 , n25957 , n25958 , n25959 , n25960 , n25961 , n25962 , n25963 , n25964 , n25965 , n25966 , n25967 , n25968 , n25969 , n25970 , n25971 , n25972 , n25973 , n25974 , n25975 , n25976 , n25977 , n25978 , n25979 , n25980 , n25981 , n25982 , n25983 , n25984 , n25985 , n25986 , n25987 , n25988 , n25989 , n25990 , n25991 , n25992 , n25993 , n25994 , n25995 , n25996 , n25997 , n25998 , n25999 , n26000 , n26001 , n26002 , n26003 , n26004 , n26005 , n26006 , n26007 , n26008 , n26009 , n26010 , n26011 , n26012 , n26013 , n26014 , n26015 , n26016 , n26017 , n26018 , n26019 , n26020 , n26021 , n26022 , n26023 , n26024 , n26025 , n26026 , n26027 , n26028 , n26029 , n26030 , n26031 , n26032 , n26033 , n26034 , n26035 , n26036 , n26037 , n26038 , n26039 , n26040 , n26041 , n26042 , n26043 , n26044 , n26045 , n26046 , n26047 , n26048 , n26049 , n26050 , n26051 , n26052 , n26053 , n26054 , n26055 , n26056 , n26057 , n26058 , n26059 , n26060 , n26061 , n26062 , n26063 , n26064 , n26065 , n26066 , n26067 , n26068 , n26069 , n26070 , n26071 , n26072 , n26073 , n26074 , n26075 , n26076 , n26077 , n26078 , n26079 , n26080 , n26081 , n26082 , n26083 , n26084 , n26085 , n26086 , n26087 , n26088 , n26089 , n26090 , n26091 , n26092 , n26093 , n26094 , n26095 , n26096 , n26097 , n26098 , n26099 , n26100 , n26101 , n26102 , n26103 , n26104 , n26105 , n26106 , n26107 , n26108 , n26109 , n26110 , n26111 , n26112 , n26113 , n26114 , n26115 , n26116 , n26117 , n26118 , n26119 , n26120 , n26121 , n26122 , n26123 , n26124 , n26125 , n26126 , n26127 , n26128 , n26129 , n26130 , n26131 , n26132 , n26133 , n26134 , n26135 , n26136 , n26137 , n26138 , n26139 , n26140 , n26141 , n26142 , n26143 , n26144 , n26145 , n26146 , n26147 , n26148 , n26149 , n26150 , n26151 , n26152 , n26153 , n26154 , n26155 , n26156 , n26157 , n26158 , n26159 , n26160 , n26161 , n26162 , n26163 , n26164 , n26165 , n26166 , n26167 , n26168 , n26169 , n26170 , n26171 , n26172 , n26173 , n26174 , n26175 , n26176 , n26177 , n26178 , n26179 , n26180 , n26181 , n26182 , n26183 , n26184 , n26185 , n26186 , n26187 , n26188 , n26189 , n26190 , n26191 , n26192 , n26193 , n26194 , n26195 , n26196 , n26197 , n26198 , n26199 , n26200 , n26201 , n26202 , n26203 , n26204 , n26205 , n26206 , n26207 , n26208 , n26209 , n26210 , n26211 , n26212 , n26213 , n26214 , n26215 , n26216 , n26217 , n26218 , n26219 , n26220 , n26221 , n26222 , n26223 , n26224 , n26225 , n26226 , n26227 , n26228 , n26229 , n26230 , n26231 , n26232 , n26233 , n26234 , n26235 , n26236 , n26237 , n26238 , n26239 , n26240 , n26241 , n26242 , n26243 , n26244 , n26245 , n26246 , n26247 , n26248 , n26249 , n26250 , n26251 , n26252 , n26253 , n26254 , n26255 , n26256 , n26257 , n26258 , n26259 , n26260 , n26261 , n26262 , n26263 , n26264 , n26265 , n26266 , n26267 , n26268 , n26269 , n26270 , n26271 , n26272 , n26273 , n26274 , n26275 , n26276 , n26277 , n26278 , n26279 , n26280 , n26281 , n26282 , n26283 , n26284 , n26285 , n26286 , n26287 , n26288 , n26289 , n26290 , n26291 , n26292 , n26293 , n26294 , n26295 , n26296 , n26297 , n26298 , n26299 , n26300 , n26301 , n26302 , n26303 , n26304 , n26305 , n26306 , n26307 , n26308 , n26309 , n26310 , n26311 , n26312 , n26313 , n26314 , n26315 , n26316 , n26317 , n26318 , n26319 , n26320 , n26321 , n26322 , n26323 , n26324 , n26325 , n26326 , n26327 , n26328 , n26329 , n26330 , n26331 , n26332 , n26333 , n26334 , n26335 , n26336 , n26337 , n26338 , n26339 , n26340 , n26341 , n26342 , n26343 , n26344 , n26345 , n26346 , n26347 , n26348 , n26349 , n26350 , n26351 , n26352 , n26353 , n26354 , n26355 , n26356 , n26357 , n26358 , n26359 , n26360 , n26361 , n26362 , n26363 , n26364 , n26365 , n26366 , n26367 , n26368 , n26369 , n26370 , n26371 , n26372 , n26373 , n26374 , n26375 , n26376 , n26377 , n26378 , n26379 , n26380 , n26381 , n26382 , n26383 , n26384 , n26385 , n26386 , n26387 , n26388 , n26389 , n26390 , n26391 , n26392 , n26393 , n26394 , n26395 , n26396 , n26397 , n26398 , n26399 , n26400 , n26401 , n26402 , n26403 , n26404 , n26405 , n26406 , n26407 , n26408 , n26409 , n26410 , n26411 , n26412 , n26413 , n26414 , n26415 , n26416 , n26417 , n26418 , n26419 , n26420 , n26421 , n26422 , n26423 , n26424 , n26425 , n26426 , n26427 , n26428 , n26429 , n26430 , n26431 , n26432 , n26433 , n26434 , n26435 , n26436 , n26437 , n26438 , n26439 , n26440 , n26441 , n26442 , n26443 , n26444 , n26445 , n26446 , n26447 , n26448 , n26449 , n26450 , n26451 , n26452 , n26453 , n26454 , n26455 , n26456 , n26457 , n26458 , n26459 , n26460 , n26461 , n26462 , n26463 , n26464 , n26465 , n26466 , n26467 , n26468 , n26469 , n26470 , n26471 , n26472 , n26473 , n26474 , n26475 , n26476 , n26477 , n26478 , n26479 , n26480 , n26481 , n26482 , n26483 , n26484 , n26485 , n26486 , n26487 , n26488 , n26489 , n26490 , n26491 , n26492 , n26493 , n26494 , n26495 , n26496 , n26497 , n26498 , n26499 , n26500 , n26501 , n26502 , n26503 , n26504 , n26505 , n26506 , n26507 , n26508 , n26509 , n26510 , n26511 , n26512 , n26513 , n26514 , n26515 , n26516 , n26517 , n26518 , n26519 , n26520 , n26521 , n26522 , n26523 , n26524 , n26525 , n26526 , n26527 , n26528 , n26529 , n26530 , n26531 , n26532 , n26533 , n26534 , n26535 , n26536 , n26537 , n26538 , n26539 , n26540 , n26541 , n26542 , n26543 , n26544 , n26545 , n26546 , n26547 , n26548 , n26549 , n26550 , n26551 , n26552 , n26553 , n26554 , n26555 , n26556 , n26557 , n26558 , n26559 , n26560 , n26561 , n26562 , n26563 , n26564 , n26565 , n26566 , n26567 , n26568 , n26569 , n26570 , n26571 , n26572 , n26573 , n26574 , n26575 , n26576 , n26577 , n26578 , n26579 , n26580 , n26581 , n26582 , n26583 , n26584 , n26585 , n26586 , n26587 , n26588 , n26589 , n26590 , n26591 , n26592 , n26593 , n26594 , n26595 , n26596 , n26597 , n26598 , n26599 , n26600 , n26601 , n26602 , n26603 , n26604 , n26605 , n26606 , n26607 , n26608 , n26609 , n26610 , n26611 , n26612 , n26613 , n26614 , n26615 , n26616 , n26617 , n26618 , n26619 , n26620 , n26621 , n26622 , n26623 , n26624 , n26625 , n26626 , n26627 , n26628 , n26629 , n26630 , n26631 , n26632 , n26633 , n26634 , n26635 , n26636 , n26637 , n26638 , n26639 , n26640 , n26641 , n26642 , n26643 , n26644 , n26645 , n26646 , n26647 , n26648 , n26649 , n26650 , n26651 , n26652 , n26653 , n26654 , n26655 , n26656 , n26657 , n26658 , n26659 , n26660 , n26661 , n26662 , n26663 , n26664 , n26665 , n26666 , n26667 , n26668 , n26669 , n26670 , n26671 , n26672 , n26673 , n26674 , n26675 , n26676 , n26677 , n26678 , n26679 , n26680 , n26681 , n26682 , n26683 , n26684 , n26685 , n26686 , n26687 , n26688 , n26689 , n26690 , n26691 , n26692 , n26693 , n26694 , n26695 , n26696 , n26697 , n26698 , n26699 , n26700 , n26701 , n26702 , n26703 , n26704 , n26705 , n26706 , n26707 , n26708 , n26709 , n26710 , n26711 , n26712 , n26713 , n26714 , n26715 , n26716 , n26717 , n26718 , n26719 , n26720 , n26721 , n26722 , n26723 , n26724 , n26725 , n26726 , n26727 , n26728 , n26729 , n26730 , n26731 , n26732 , n26733 , n26734 , n26735 , n26736 , n26737 , n26738 , n26739 , n26740 , n26741 , n26742 , n26743 , n26744 , n26745 , n26746 , n26747 , n26748 , n26749 , n26750 , n26751 , n26752 , n26753 , n26754 , n26755 , n26756 , n26757 , n26758 , n26759 , n26760 , n26761 , n26762 , n26763 , n26764 , n26765 , n26766 , n26767 , n26768 , n26769 , n26770 , n26771 , n26772 , n26773 , n26774 , n26775 , n26776 , n26777 , n26778 , n26779 , n26780 , n26781 , n26782 , n26783 , n26784 , n26785 , n26786 , n26787 , n26788 , n26789 , n26790 , n26791 , n26792 , n26793 , n26794 , n26795 , n26796 , n26797 , n26798 , n26799 , n26800 , n26801 , n26802 , n26803 , n26804 , n26805 , n26806 , n26807 , n26808 , n26809 , n26810 , n26811 , n26812 , n26813 , n26814 , n26815 , n26816 , n26817 , n26818 , n26819 , n26820 , n26821 , n26822 , n26823 , n26824 , n26825 , n26826 , n26827 , n26828 , n26829 , n26830 , n26831 , n26832 , n26833 , n26834 , n26835 , n26836 , n26837 , n26838 , n26839 , n26840 , n26841 , n26842 , n26843 , n26844 , n26845 , n26846 , n26847 , n26848 , n26849 , n26850 , n26851 , n26852 , n26853 , n26854 , n26855 , n26856 , n26857 , n26858 , n26859 , n26860 , n26861 , n26862 , n26863 , n26864 , n26865 , n26866 , n26867 , n26868 , n26869 , n26870 , n26871 , n26872 , n26873 , n26874 , n26875 , n26876 , n26877 , n26878 , n26879 , n26880 , n26881 , n26882 , n26883 , n26884 , n26885 , n26886 , n26887 , n26888 , n26889 , n26890 , n26891 , n26892 , n26893 , n26894 , n26895 , n26896 , n26897 , n26898 , n26899 , n26900 , n26901 , n26902 , n26903 , n26904 , n26905 , n26906 , n26907 , n26908 , n26909 , n26910 , n26911 , n26912 , n26913 , n26914 , n26915 , n26916 , n26917 , n26918 , n26919 , n26920 , n26921 , n26922 , n26923 , n26924 , n26925 , n26926 , n26927 , n26928 , n26929 , n26930 , n26931 , n26932 , n26933 , n26934 , n26935 , n26936 , n26937 , n26938 , n26939 , n26940 , n26941 , n26942 , n26943 , n26944 , n26945 , n26946 , n26947 , n26948 , n26949 , n26950 , n26951 , n26952 , n26953 , n26954 , n26955 , n26956 , n26957 , n26958 , n26959 , n26960 , n26961 , n26962 , n26963 , n26964 , n26965 , n26966 , n26967 , n26968 , n26969 , n26970 , n26971 , n26972 , n26973 , n26974 , n26975 , n26976 , n26977 , n26978 , n26979 , n26980 , n26981 , n26982 , n26983 , n26984 , n26985 , n26986 , n26987 , n26988 , n26989 , n26990 , n26991 , n26992 , n26993 , n26994 , n26995 , n26996 , n26997 , n26998 , n26999 , n27000 , n27001 , n27002 , n27003 , n27004 , n27005 , n27006 , n27007 , n27008 , n27009 , n27010 , n27011 , n27012 , n27013 , n27014 , n27015 , n27016 , n27017 , n27018 , n27019 , n27020 , n27021 , n27022 , n27023 , n27024 , n27025 , n27026 , n27027 , n27028 , n27029 , n27030 , n27031 , n27032 , n27033 , n27034 , n27035 , n27036 , n27037 , n27038 , n27039 , n27040 , n27041 , n27042 , n27043 , n27044 , n27045 , n27046 , n27047 , n27048 , n27049 , n27050 , n27051 , n27052 , n27053 , n27054 , n27055 , n27056 , n27057 , n27058 , n27059 , n27060 , n27061 , n27062 , n27063 , n27064 , n27065 , n27066 , n27067 , n27068 , n27069 , n27070 , n27071 , n27072 , n27073 , n27074 , n27075 , n27076 , n27077 , n27078 , n27079 , n27080 , n27081 , n27082 , n27083 , n27084 , n27085 , n27086 , n27087 , n27088 , n27089 , n27090 , n27091 , n27092 , n27093 , n27094 , n27095 , n27096 , n27097 , n27098 , n27099 , n27100 , n27101 , n27102 , n27103 , n27104 , n27105 , n27106 , n27107 , n27108 , n27109 , n27110 , n27111 , n27112 , n27113 , n27114 , n27115 , n27116 , n27117 , n27118 , n27119 , n27120 , n27121 , n27122 , n27123 , n27124 , n27125 , n27126 , n27127 , n27128 , n27129 , n27130 , n27131 , n27132 , n27133 , n27134 , n27135 , n27136 , n27137 , n27138 , n27139 , n27140 , n27141 , n27142 , n27143 , n27144 , n27145 , n27146 , n27147 , n27148 , n27149 , n27150 , n27151 , n27152 , n27153 , n27154 , n27155 , n27156 , n27157 , n27158 , n27159 , n27160 , n27161 , n27162 , n27163 , n27164 , n27165 , n27166 , n27167 , n27168 , n27169 , n27170 , n27171 , n27172 , n27173 , n27174 , n27175 , n27176 , n27177 , n27178 , n27179 , n27180 , n27181 , n27182 , n27183 , n27184 , n27185 , n27186 , n27187 , n27188 , n27189 , n27190 , n27191 , n27192 , n27193 , n27194 , n27195 , n27196 , n27197 , n27198 , n27199 , n27200 , n27201 , n27202 , n27203 , n27204 , n27205 , n27206 , n27207 , n27208 , n27209 , n27210 , n27211 , n27212 , n27213 , n27214 , n27215 , n27216 , n27217 , n27218 , n27219 , n27220 , n27221 , n27222 , n27223 , n27224 , n27225 , n27226 , n27227 , n27228 , n27229 , n27230 , n27231 , n27232 , n27233 , n27234 , n27235 , n27236 , n27237 , n27238 , n27239 , n27240 , n27241 , n27242 , n27243 , n27244 , n27245 , n27246 , n27247 , n27248 , n27249 , n27250 , n27251 , n27252 , n27253 , n27254 , n27255 , n27256 , n27257 , n27258 , n27259 , n27260 , n27261 , n27262 , n27263 , n27264 , n27265 , n27266 , n27267 , n27268 , n27269 , n27270 , n27271 , n27272 , n27273 , n27274 , n27275 , n27276 , n27277 , n27278 , n27279 , n27280 , n27281 , n27282 , n27283 , n27284 , n27285 , n27286 , n27287 , n27288 , n27289 , n27290 , n27291 , n27292 , n27293 , n27294 , n27295 , n27296 , n27297 , n27298 , n27299 , n27300 , n27301 , n27302 , n27303 , n27304 , n27305 , n27306 , n27307 , n27308 , n27309 , n27310 , n27311 , n27312 , n27313 , n27314 , n27315 , n27316 , n27317 , n27318 , n27319 , n27320 , n27321 , n27322 , n27323 , n27324 , n27325 , n27326 , n27327 , n27328 , n27329 , n27330 , n27331 , n27332 , n27333 , n27334 , n27335 , n27336 , n27337 , n27338 , n27339 , n27340 , n27341 , n27342 , n27343 , n27344 , n27345 , n27346 , n27347 , n27348 , n27349 , n27350 , n27351 , n27352 , n27353 , n27354 , n27355 , n27356 , n27357 , n27358 , n27359 , n27360 , n27361 , n27362 , n27363 , n27364 , n27365 , n27366 , n27367 , n27368 , n27369 , n27370 , n27371 , n27372 , n27373 , n27374 , n27375 , n27376 , n27377 , n27378 , n27379 , n27380 , n27381 , n27382 , n27383 , n27384 , n27385 , n27386 , n27387 , n27388 , n27389 , n27390 , n27391 , n27392 , n27393 , n27394 , n27395 , n27396 , n27397 , n27398 , n27399 , n27400 , n27401 , n27402 , n27403 , n27404 , n27405 , n27406 , n27407 , n27408 , n27409 , n27410 , n27411 , n27412 , n27413 , n27414 , n27415 , n27416 , n27417 , n27418 , n27419 , n27420 , n27421 , n27422 , n27423 , n27424 , n27425 , n27426 , n27427 , n27428 , n27429 , n27430 , n27431 , n27432 , n27433 , n27434 , n27435 , n27436 , n27437 , n27438 , n27439 , n27440 , n27441 , n27442 , n27443 , n27444 , n27445 , n27446 , n27447 , n27448 , n27449 , n27450 , n27451 , n27452 , n27453 , n27454 , n27455 , n27456 , n27457 , n27458 , n27459 , n27460 , n27461 , n27462 , n27463 , n27464 , n27465 , n27466 , n27467 , n27468 , n27469 , n27470 , n27471 , n27472 , n27473 , n27474 , n27475 , n27476 , n27477 , n27478 , n27479 , n27480 , n27481 , n27482 , n27483 , n27484 , n27485 , n27486 , n27487 , n27488 , n27489 , n27490 , n27491 , n27492 , n27493 , n27494 , n27495 , n27496 , n27497 , n27498 , n27499 , n27500 , n27501 , n27502 , n27503 , n27504 , n27505 , n27506 , n27507 , n27508 , n27509 , n27510 , n27511 , n27512 , n27513 , n27514 , n27515 , n27516 , n27517 , n27518 , n27519 , n27520 , n27521 , n27522 , n27523 , n27524 , n27525 , n27526 , n27527 , n27528 , n27529 , n27530 , n27531 , n27532 , n27533 , n27534 , n27535 , n27536 , n27537 , n27538 , n27539 , n27540 , n27541 , n27542 , n27543 , n27544 , n27545 , n27546 , n27547 , n27548 , n27549 , n27550 , n27551 , n27552 , n27553 , n27554 , n27555 , n27556 , n27557 , n27558 , n27559 , n27560 , n27561 , n27562 , n27563 , n27564 , n27565 , n27566 , n27567 , n27568 , n27569 , n27570 , n27571 , n27572 , n27573 , n27574 , n27575 , n27576 , n27577 , n27578 , n27579 , n27580 , n27581 , n27582 , n27583 , n27584 , n27585 , n27586 , n27587 , n27588 , n27589 , n27590 , n27591 , n27592 , n27593 , n27594 , n27595 , n27596 , n27597 , n27598 , n27599 , n27600 , n27601 , n27602 , n27603 , n27604 , n27605 , n27606 , n27607 , n27608 , n27609 , n27610 , n27611 , n27612 , n27613 , n27614 , n27615 , n27616 , n27617 , n27618 , n27619 , n27620 , n27621 , n27622 , n27623 , n27624 , n27625 , n27626 , n27627 , n27628 , n27629 , n27630 , n27631 , n27632 , n27633 , n27634 , n27635 , n27636 , n27637 , n27638 , n27639 , n27640 , n27641 , n27642 , n27643 , n27644 , n27645 , n27646 , n27647 , n27648 , n27649 , n27650 , n27651 , n27652 , n27653 , n27654 , n27655 , n27656 , n27657 , n27658 , n27659 , n27660 , n27661 , n27662 , n27663 , n27664 , n27665 , n27666 , n27667 , n27668 , n27669 , n27670 , n27671 , n27672 , n27673 , n27674 , n27675 , n27676 , n27677 , n27678 , n27679 , n27680 , n27681 , n27682 , n27683 , n27684 , n27685 , n27686 , n27687 , n27688 , n27689 , n27690 , n27691 , n27692 , n27693 , n27694 , n27695 , n27696 , n27697 , n27698 , n27699 , n27700 , n27701 , n27702 , n27703 , n27704 , n27705 , n27706 , n27707 , n27708 , n27709 , n27710 , n27711 , n27712 , n27713 , n27714 , n27715 , n27716 , n27717 , n27718 , n27719 , n27720 , n27721 , n27722 , n27723 , n27724 , n27725 , n27726 , n27727 , n27728 , n27729 , n27730 , n27731 , n27732 , n27733 , n27734 , n27735 , n27736 , n27737 , n27738 , n27739 , n27740 , n27741 , n27742 , n27743 , n27744 , n27745 , n27746 , n27747 , n27748 , n27749 , n27750 , n27751 , n27752 , n27753 , n27754 , n27755 , n27756 , n27757 , n27758 , n27759 , n27760 , n27761 , n27762 , n27763 , n27764 , n27765 , n27766 , n27767 , n27768 , n27769 , n27770 , n27771 , n27772 , n27773 , n27774 , n27775 , n27776 , n27777 , n27778 , n27779 , n27780 , n27781 , n27782 , n27783 , n27784 , n27785 , n27786 , n27787 , n27788 , n27789 , n27790 , n27791 , n27792 , n27793 , n27794 , n27795 , n27796 , n27797 , n27798 , n27799 , n27800 , n27801 , n27802 , n27803 , n27804 , n27805 , n27806 , n27807 , n27808 , n27809 , n27810 , n27811 , n27812 , n27813 , n27814 , n27815 , n27816 , n27817 , n27818 , n27819 , n27820 , n27821 , n27822 , n27823 , n27824 , n27825 , n27826 , n27827 , n27828 , n27829 , n27830 , n27831 , n27832 , n27833 , n27834 , n27835 , n27836 , n27837 , n27838 , n27839 , n27840 , n27841 , n27842 , n27843 , n27844 , n27845 , n27846 , n27847 , n27848 , n27849 , n27850 , n27851 , n27852 , n27853 , n27854 , n27855 , n27856 , n27857 , n27858 , n27859 , n27860 , n27861 , n27862 , n27863 , n27864 , n27865 , n27866 , n27867 , n27868 , n27869 , n27870 , n27871 , n27872 , n27873 , n27874 , n27875 , n27876 , n27877 , n27878 , n27879 , n27880 , n27881 , n27882 , n27883 , n27884 , n27885 , n27886 , n27887 , n27888 , n27889 , n27890 , n27891 , n27892 , n27893 , n27894 , n27895 , n27896 , n27897 , n27898 , n27899 , n27900 , n27901 , n27902 , n27903 , n27904 , n27905 , n27906 , n27907 , n27908 , n27909 , n27910 , n27911 , n27912 , n27913 , n27914 , n27915 , n27916 , n27917 , n27918 , n27919 , n27920 , n27921 , n27922 , n27923 , n27924 , n27925 , n27926 , n27927 , n27928 , n27929 , n27930 , n27931 , n27932 , n27933 , n27934 , n27935 , n27936 , n27937 , n27938 , n27939 , n27940 , n27941 , n27942 , n27943 , n27944 , n27945 , n27946 , n27947 , n27948 , n27949 , n27950 , n27951 , n27952 , n27953 , n27954 , n27955 , n27956 , n27957 , n27958 , n27959 , n27960 , n27961 , n27962 , n27963 , n27964 , n27965 , n27966 , n27967 , n27968 , n27969 , n27970 , n27971 , n27972 , n27973 , n27974 , n27975 , n27976 , n27977 , n27978 , n27979 , n27980 , n27981 , n27982 , n27983 , n27984 , n27985 , n27986 , n27987 , n27988 , n27989 , n27990 , n27991 , n27992 , n27993 , n27994 , n27995 , n27996 , n27997 , n27998 , n27999 , n28000 , n28001 , n28002 , n28003 , n28004 , n28005 , n28006 , n28007 , n28008 , n28009 , n28010 , n28011 , n28012 , n28013 , n28014 , n28015 , n28016 , n28017 , n28018 , n28019 , n28020 , n28021 , n28022 , n28023 , n28024 , n28025 , n28026 , n28027 , n28028 , n28029 , n28030 , n28031 , n28032 , n28033 , n28034 , n28035 , n28036 , n28037 , n28038 , n28039 , n28040 , n28041 , n28042 , n28043 , n28044 , n28045 , n28046 , n28047 , n28048 , n28049 , n28050 , n28051 , n28052 , n28053 , n28054 , n28055 , n28056 , n28057 , n28058 , n28059 , n28060 , n28061 , n28062 , n28063 , n28064 , n28065 , n28066 , n28067 , n28068 , n28069 , n28070 , n28071 , n28072 , n28073 , n28074 , n28075 , n28076 , n28077 , n28078 , n28079 , n28080 , n28081 , n28082 , n28083 , n28084 , n28085 , n28086 , n28087 , n28088 , n28089 , n28090 , n28091 , n28092 , n28093 , n28094 , n28095 , n28096 , n28097 , n28098 , n28099 , n28100 , n28101 , n28102 , n28103 , n28104 , n28105 , n28106 , n28107 , n28108 , n28109 , n28110 , n28111 , n28112 , n28113 , n28114 , n28115 , n28116 , n28117 , n28118 , n28119 , n28120 , n28121 , n28122 , n28123 , n28124 , n28125 , n28126 , n28127 , n28128 , n28129 , n28130 , n28131 , n28132 , n28133 , n28134 , n28135 , n28136 , n28137 , n28138 , n28139 , n28140 , n28141 , n28142 , n28143 , n28144 , n28145 , n28146 , n28147 , n28148 , n28149 , n28150 , n28151 , n28152 , n28153 , n28154 , n28155 , n28156 , n28157 , n28158 , n28159 , n28160 , n28161 , n28162 , n28163 , n28164 , n28165 , n28166 , n28167 , n28168 , n28169 , n28170 , n28171 , n28172 , n28173 , n28174 , n28175 , n28176 , n28177 , n28178 , n28179 , n28180 , n28181 , n28182 , n28183 , n28184 , n28185 , n28186 , n28187 , n28188 , n28189 , n28190 , n28191 , n28192 , n28193 , n28194 , n28195 , n28196 , n28197 , n28198 , n28199 , n28200 , n28201 , n28202 , n28203 , n28204 , n28205 , n28206 , n28207 , n28208 , n28209 , n28210 , n28211 , n28212 , n28213 , n28214 , n28215 , n28216 , n28217 , n28218 , n28219 , n28220 , n28221 , n28222 , n28223 , n28224 , n28225 , n28226 , n28227 , n28228 , n28229 , n28230 , n28231 , n28232 , n28233 , n28234 , n28235 , n28236 , n28237 , n28238 , n28239 , n28240 , n28241 , n28242 , n28243 , n28244 , n28245 , n28246 , n28247 , n28248 , n28249 , n28250 , n28251 , n28252 , n28253 , n28254 , n28255 , n28256 , n28257 , n28258 , n28259 , n28260 , n28261 , n28262 , n28263 , n28264 , n28265 , n28266 , n28267 , n28268 , n28269 , n28270 , n28271 , n28272 , n28273 , n28274 , n28275 , n28276 , n28277 , n28278 , n28279 , n28280 , n28281 , n28282 , n28283 , n28284 , n28285 , n28286 , n28287 , n28288 , n28289 , n28290 , n28291 , n28292 , n28293 , n28294 , n28295 , n28296 , n28297 , n28298 , n28299 , n28300 , n28301 , n28302 , n28303 , n28304 , n28305 , n28306 , n28307 , n28308 , n28309 , n28310 , n28311 , n28312 , n28313 , n28314 , n28315 , n28316 , n28317 , n28318 , n28319 , n28320 , n28321 , n28322 , n28323 , n28324 , n28325 , n28326 , n28327 , n28328 , n28329 , n28330 , n28331 , n28332 , n28333 , n28334 , n28335 , n28336 , n28337 , n28338 , n28339 , n28340 , n28341 , n28342 , n28343 , n28344 , n28345 , n28346 , n28347 , n28348 , n28349 , n28350 , n28351 , n28352 , n28353 , n28354 , n28355 , n28356 , n28357 , n28358 , n28359 , n28360 , n28361 , n28362 , n28363 , n28364 , n28365 , n28366 , n28367 , n28368 , n28369 , n28370 , n28371 , n28372 , n28373 , n28374 , n28375 , n28376 , n28377 , n28378 , n28379 , n28380 , n28381 , n28382 , n28383 , n28384 , n28385 , n28386 , n28387 , n28388 , n28389 , n28390 , n28391 , n28392 , n28393 , n28394 , n28395 , n28396 , n28397 , n28398 , n28399 , n28400 , n28401 , n28402 , n28403 , n28404 , n28405 , n28406 , n28407 , n28408 , n28409 , n28410 , n28411 , n28412 , n28413 , n28414 , n28415 , n28416 , n28417 , n28418 , n28419 , n28420 , n28421 , n28422 , n28423 , n28424 , n28425 , n28426 , n28427 , n28428 , n28429 , n28430 , n28431 , n28432 , n28433 , n28434 , n28435 , n28436 , n28437 , n28438 , n28439 , n28440 , n28441 , n28442 , n28443 , n28444 , n28445 , n28446 , n28447 , n28448 , n28449 , n28450 , n28451 , n28452 , n28453 , n28454 , n28455 , n28456 , n28457 , n28458 , n28459 , n28460 , n28461 , n28462 , n28463 , n28464 , n28465 , n28466 , n28467 , n28468 , n28469 , n28470 , n28471 , n28472 , n28473 , n28474 , n28475 , n28476 , n28477 , n28478 , n28479 , n28480 , n28481 , n28482 , n28483 , n28484 , n28485 , n28486 , n28487 , n28488 , n28489 , n28490 , n28491 , n28492 , n28493 , n28494 , n28495 , n28496 , n28497 , n28498 , n28499 , n28500 , n28501 , n28502 , n28503 , n28504 , n28505 , n28506 , n28507 , n28508 , n28509 , n28510 , n28511 , n28512 , n28513 , n28514 , n28515 , n28516 , n28517 , n28518 , n28519 , n28520 , n28521 , n28522 , n28523 , n28524 , n28525 , n28526 , n28527 , n28528 , n28529 , n28530 , n28531 , n28532 , n28533 , n28534 , n28535 , n28536 , n28537 , n28538 , n28539 , n28540 , n28541 , n28542 , n28543 , n28544 , n28545 , n28546 , n28547 , n28548 , n28549 , n28550 , n28551 , n28552 , n28553 , n28554 , n28555 , n28556 , n28557 , n28558 , n28559 , n28560 , n28561 , n28562 , n28563 , n28564 , n28565 , n28566 , n28567 , n28568 , n28569 , n28570 , n28571 , n28572 , n28573 , n28574 , n28575 , n28576 , n28577 , n28578 , n28579 , n28580 , n28581 , n28582 , n28583 , n28584 , n28585 , n28586 , n28587 , n28588 , n28589 , n28590 , n28591 , n28592 , n28593 , n28594 , n28595 , n28596 , n28597 , n28598 , n28599 , n28600 , n28601 , n28602 , n28603 , n28604 , n28605 , n28606 , n28607 , n28608 , n28609 , n28610 , n28611 , n28612 , n28613 , n28614 , n28615 , n28616 , n28617 , n28618 , n28619 , n28620 , n28621 , n28622 , n28623 , n28624 , n28625 , n28626 , n28627 , n28628 , n28629 , n28630 , n28631 , n28632 , n28633 , n28634 , n28635 , n28636 , n28637 , n28638 , n28639 , n28640 , n28641 , n28642 , n28643 , n28644 , n28645 , n28646 , n28647 , n28648 , n28649 , n28650 , n28651 , n28652 , n28653 , n28654 , n28655 , n28656 , n28657 , n28658 , n28659 , n28660 , n28661 , n28662 , n28663 , n28664 , n28665 , n28666 , n28667 , n28668 , n28669 , n28670 , n28671 , n28672 , n28673 , n28674 , n28675 , n28676 , n28677 , n28678 , n28679 , n28680 , n28681 , n28682 , n28683 , n28684 , n28685 , n28686 , n28687 , n28688 , n28689 , n28690 , n28691 , n28692 , n28693 , n28694 , n28695 , n28696 , n28697 , n28698 , n28699 , n28700 , n28701 , n28702 , n28703 , n28704 , n28705 , n28706 , n28707 , n28708 , n28709 , n28710 , n28711 , n28712 , n28713 , n28714 , n28715 , n28716 , n28717 , n28718 , n28719 , n28720 , n28721 , n28722 , n28723 , n28724 , n28725 , n28726 , n28727 , n28728 , n28729 , n28730 , n28731 , n28732 , n28733 , n28734 , n28735 , n28736 , n28737 , n28738 , n28739 , n28740 , n28741 , n28742 , n28743 , n28744 , n28745 , n28746 , n28747 , n28748 , n28749 , n28750 , n28751 , n28752 , n28753 , n28754 , n28755 , n28756 , n28757 , n28758 , n28759 , n28760 , n28761 , n28762 , n28763 , n28764 , n28765 , n28766 , n28767 , n28768 , n28769 , n28770 , n28771 , n28772 , n28773 , n28774 , n28775 , n28776 , n28777 , n28778 , n28779 , n28780 , n28781 , n28782 , n28783 , n28784 , n28785 , n28786 , n28787 , n28788 , n28789 , n28790 , n28791 , n28792 , n28793 , n28794 , n28795 , n28796 , n28797 , n28798 , n28799 , n28800 , n28801 , n28802 , n28803 , n28804 , n28805 , n28806 , n28807 , n28808 , n28809 , n28810 , n28811 , n28812 , n28813 , n28814 , n28815 , n28816 , n28817 , n28818 , n28819 , n28820 , n28821 , n28822 , n28823 , n28824 , n28825 , n28826 , n28827 , n28828 , n28829 , n28830 , n28831 , n28832 , n28833 , n28834 , n28835 , n28836 , n28837 , n28838 , n28839 , n28840 , n28841 , n28842 , n28843 , n28844 , n28845 , n28846 , n28847 , n28848 , n28849 , n28850 , n28851 , n28852 , n28853 , n28854 , n28855 , n28856 , n28857 , n28858 , n28859 , n28860 , n28861 , n28862 , n28863 , n28864 , n28865 , n28866 , n28867 , n28868 , n28869 , n28870 , n28871 , n28872 , n28873 , n28874 , n28875 , n28876 , n28877 , n28878 , n28879 , n28880 , n28881 , n28882 , n28883 , n28884 , n28885 , n28886 , n28887 , n28888 , n28889 , n28890 , n28891 , n28892 , n28893 , n28894 , n28895 , n28896 , n28897 , n28898 , n28899 , n28900 , n28901 , n28902 , n28903 , n28904 , n28905 , n28906 , n28907 , n28908 , n28909 , n28910 , n28911 , n28912 , n28913 , n28914 , n28915 , n28916 , n28917 , n28918 , n28919 , n28920 , n28921 , n28922 , n28923 , n28924 , n28925 , n28926 , n28927 , n28928 , n28929 , n28930 , n28931 , n28932 , n28933 , n28934 , n28935 , n28936 , n28937 , n28938 , n28939 , n28940 , n28941 , n28942 , n28943 , n28944 , n28945 , n28946 , n28947 , n28948 , n28949 , n28950 , n28951 , n28952 , n28953 , n28954 , n28955 , n28956 , n28957 , n28958 , n28959 , n28960 , n28961 , n28962 , n28963 , n28964 , n28965 , n28966 , n28967 , n28968 , n28969 , n28970 , n28971 , n28972 , n28973 , n28974 , n28975 , n28976 , n28977 , n28978 , n28979 , n28980 , n28981 , n28982 , n28983 , n28984 , n28985 , n28986 , n28987 , n28988 , n28989 , n28990 , n28991 , n28992 , n28993 , n28994 , n28995 , n28996 , n28997 , n28998 , n28999 , n29000 , n29001 , n29002 , n29003 , n29004 , n29005 , n29006 , n29007 , n29008 , n29009 , n29010 , n29011 , n29012 , n29013 , n29014 , n29015 , n29016 , n29017 , n29018 , n29019 , n29020 , n29021 , n29022 , n29023 , n29024 , n29025 , n29026 , n29027 , n29028 , n29029 , n29030 , n29031 , n29032 , n29033 , n29034 , n29035 , n29036 , n29037 , n29038 , n29039 , n29040 , n29041 , n29042 , n29043 , n29044 , n29045 , n29046 , n29047 , n29048 , n29049 , n29050 , n29051 , n29052 , n29053 , n29054 , n29055 , n29056 , n29057 , n29058 , n29059 , n29060 , n29061 , n29062 , n29063 , n29064 , n29065 , n29066 , n29067 , n29068 , n29069 , n29070 , n29071 , n29072 , n29073 , n29074 , n29075 , n29076 , n29077 , n29078 , n29079 , n29080 , n29081 , n29082 , n29083 , n29084 , n29085 , n29086 , n29087 , n29088 , n29089 , n29090 , n29091 , n29092 , n29093 , n29094 , n29095 , n29096 , n29097 , n29098 , n29099 , n29100 , n29101 , n29102 , n29103 , n29104 , n29105 , n29106 , n29107 , n29108 , n29109 , n29110 , n29111 , n29112 , n29113 , n29114 , n29115 , n29116 , n29117 , n29118 , n29119 , n29120 , n29121 , n29122 , n29123 , n29124 , n29125 , n29126 , n29127 , n29128 , n29129 , n29130 , n29131 , n29132 , n29133 , n29134 , n29135 , n29136 , n29137 , n29138 , n29139 , n29140 , n29141 , n29142 , n29143 , n29144 , n29145 , n29146 , n29147 , n29148 , n29149 , n29150 , n29151 , n29152 , n29153 , n29154 , n29155 , n29156 , n29157 , n29158 , n29159 , n29160 , n29161 , n29162 , n29163 , n29164 , n29165 , n29166 , n29167 , n29168 , n29169 , n29170 , n29171 , n29172 , n29173 , n29174 , n29175 , n29176 , n29177 , n29178 , n29179 , n29180 , n29181 , n29182 , n29183 , n29184 , n29185 , n29186 , n29187 , n29188 , n29189 , n29190 , n29191 , n29192 , n29193 , n29194 , n29195 , n29196 , n29197 , n29198 , n29199 , n29200 , n29201 , n29202 , n29203 , n29204 , n29205 , n29206 , n29207 , n29208 , n29209 , n29210 , n29211 , n29212 , n29213 , n29214 , n29215 , n29216 , n29217 , n29218 , n29219 , n29220 , n29221 , n29222 , n29223 , n29224 , n29225 , n29226 , n29227 , n29228 , n29229 , n29230 , n29231 , n29232 , n29233 , n29234 , n29235 , n29236 , n29237 , n29238 , n29239 , n29240 , n29241 , n29242 , n29243 , n29244 , n29245 , n29246 , n29247 , n29248 , n29249 , n29250 , n29251 , n29252 , n29253 , n29254 , n29255 , n29256 , n29257 , n29258 , n29259 , n29260 , n29261 , n29262 , n29263 , n29264 , n29265 , n29266 , n29267 , n29268 , n29269 , n29270 , n29271 , n29272 , n29273 , n29274 , n29275 , n29276 , n29277 , n29278 , n29279 , n29280 , n29281 , n29282 , n29283 , n29284 , n29285 , n29286 , n29287 , n29288 , n29289 , n29290 , n29291 , n29292 , n29293 , n29294 , n29295 , n29296 , n29297 , n29298 , n29299 , n29300 , n29301 , n29302 , n29303 , n29304 , n29305 , n29306 , n29307 , n29308 , n29309 , n29310 , n29311 , n29312 , n29313 , n29314 , n29315 , n29316 , n29317 , n29318 , n29319 , n29320 , n29321 , n29322 , n29323 , n29324 , n29325 , n29326 , n29327 , n29328 , n29329 , n29330 , n29331 , n29332 , n29333 , n29334 , n29335 , n29336 , n29337 , n29338 , n29339 , n29340 , n29341 , n29342 , n29343 , n29344 , n29345 , n29346 , n29347 , n29348 , n29349 , n29350 , n29351 , n29352 , n29353 , n29354 , n29355 , n29356 , n29357 , n29358 , n29359 , n29360 , n29361 , n29362 , n29363 , n29364 , n29365 , n29366 , n29367 , n29368 , n29369 , n29370 , n29371 , n29372 , n29373 , n29374 , n29375 , n29376 , n29377 , n29378 , n29379 , n29380 , n29381 , n29382 , n29383 , n29384 , n29385 , n29386 , n29387 , n29388 , n29389 , n29390 , n29391 , n29392 , n29393 , n29394 , n29395 , n29396 , n29397 , n29398 , n29399 , n29400 , n29401 , n29402 , n29403 , n29404 , n29405 , n29406 , n29407 , n29408 , n29409 , n29410 , n29411 , n29412 , n29413 , n29414 , n29415 , n29416 , n29417 , n29418 , n29419 , n29420 , n29421 , n29422 , n29423 , n29424 , n29425 , n29426 , n29427 , n29428 , n29429 , n29430 , n29431 , n29432 , n29433 , n29434 , n29435 , n29436 , n29437 , n29438 , n29439 , n29440 , n29441 , n29442 , n29443 , n29444 , n29445 , n29446 , n29447 , n29448 , n29449 , n29450 , n29451 , n29452 , n29453 , n29454 , n29455 , n29456 , n29457 , n29458 , n29459 , n29460 , n29461 , n29462 , n29463 , n29464 , n29465 , n29466 , n29467 , n29468 , n29469 , n29470 , n29471 , n29472 , n29473 , n29474 , n29475 , n29476 , n29477 , n29478 , n29479 , n29480 , n29481 , n29482 , n29483 , n29484 , n29485 , n29486 , n29487 , n29488 , n29489 , n29490 , n29491 , n29492 , n29493 , n29494 , n29495 , n29496 , n29497 , n29498 , n29499 , n29500 , n29501 , n29502 , n29503 , n29504 , n29505 , n29506 , n29507 , n29508 , n29509 , n29510 , n29511 , n29512 , n29513 , n29514 , n29515 , n29516 , n29517 , n29518 , n29519 , n29520 , n29521 , n29522 , n29523 , n29524 , n29525 , n29526 , n29527 , n29528 , n29529 , n29530 , n29531 , n29532 , n29533 , n29534 , n29535 , n29536 , n29537 , n29538 , n29539 , n29540 , n29541 , n29542 , n29543 , n29544 , n29545 , n29546 , n29547 , n29548 , n29549 , n29550 , n29551 , n29552 , n29553 , n29554 , n29555 , n29556 , n29557 , n29558 , n29559 , n29560 , n29561 , n29562 , n29563 , n29564 , n29565 , n29566 , n29567 , n29568 , n29569 , n29570 , n29571 , n29572 , n29573 , n29574 , n29575 , n29576 , n29577 , n29578 , n29579 , n29580 , n29581 , n29582 , n29583 , n29584 , n29585 , n29586 , n29587 , n29588 , n29589 , n29590 , n29591 , n29592 , n29593 , n29594 , n29595 , n29596 , n29597 , n29598 , n29599 , n29600 , n29601 , n29602 , n29603 , n29604 , n29605 , n29606 , n29607 , n29608 , n29609 , n29610 , n29611 , n29612 , n29613 , n29614 , n29615 , n29616 , n29617 , n29618 , n29619 , n29620 , n29621 , n29622 , n29623 , n29624 , n29625 , n29626 , n29627 , n29628 , n29629 , n29630 , n29631 , n29632 , n29633 , n29634 , n29635 , n29636 , n29637 , n29638 , n29639 , n29640 , n29641 , n29642 , n29643 , n29644 , n29645 , n29646 , n29647 , n29648 , n29649 , n29650 , n29651 , n29652 , n29653 , n29654 , n29655 , n29656 , n29657 , n29658 , n29659 , n29660 , n29661 , n29662 , n29663 , n29664 , n29665 , n29666 , n29667 , n29668 , n29669 , n29670 , n29671 , n29672 , n29673 , n29674 , n29675 , n29676 , n29677 , n29678 , n29679 , n29680 , n29681 , n29682 , n29683 , n29684 , n29685 , n29686 , n29687 , n29688 , n29689 , n29690 , n29691 , n29692 , n29693 , n29694 , n29695 , n29696 , n29697 , n29698 , n29699 , n29700 , n29701 , n29702 , n29703 , n29704 , n29705 , n29706 , n29707 , n29708 , n29709 , n29710 , n29711 , n29712 , n29713 , n29714 , n29715 , n29716 , n29717 , n29718 , n29719 , n29720 , n29721 , n29722 , n29723 , n29724 , n29725 , n29726 , n29727 , n29728 , n29729 , n29730 , n29731 , n29732 , n29733 , n29734 , n29735 , n29736 , n29737 , n29738 , n29739 , n29740 , n29741 , n29742 , n29743 , n29744 , n29745 , n29746 , n29747 , n29748 , n29749 , n29750 , n29751 , n29752 , n29753 , n29754 , n29755 , n29756 , n29757 , n29758 , n29759 , n29760 , n29761 , n29762 , n29763 , n29764 , n29765 , n29766 , n29767 , n29768 , n29769 , n29770 , n29771 , n29772 , n29773 , n29774 , n29775 , n29776 , n29777 , n29778 , n29779 , n29780 , n29781 , n29782 , n29783 , n29784 , n29785 , n29786 , n29787 , n29788 , n29789 , n29790 , n29791 , n29792 , n29793 , n29794 , n29795 , n29796 , n29797 , n29798 , n29799 , n29800 , n29801 , n29802 , n29803 , n29804 , n29805 , n29806 , n29807 , n29808 , n29809 , n29810 , n29811 , n29812 , n29813 , n29814 , n29815 , n29816 , n29817 , n29818 , n29819 , n29820 , n29821 , n29822 , n29823 , n29824 , n29825 , n29826 , n29827 , n29828 , n29829 , n29830 , n29831 , n29832 , n29833 , n29834 , n29835 , n29836 , n29837 , n29838 , n29839 , n29840 , n29841 , n29842 , n29843 , n29844 , n29845 , n29846 , n29847 , n29848 , n29849 , n29850 , n29851 , n29852 , n29853 , n29854 , n29855 , n29856 , n29857 , n29858 , n29859 , n29860 , n29861 , n29862 , n29863 , n29864 , n29865 , n29866 , n29867 , n29868 , n29869 , n29870 , n29871 , n29872 , n29873 , n29874 , n29875 , n29876 , n29877 , n29878 , n29879 , n29880 , n29881 , n29882 , n29883 , n29884 , n29885 , n29886 , n29887 , n29888 , n29889 , n29890 , n29891 , n29892 , n29893 , n29894 , n29895 , n29896 , n29897 , n29898 , n29899 , n29900 , n29901 , n29902 , n29903 , n29904 , n29905 , n29906 , n29907 , n29908 , n29909 , n29910 , n29911 , n29912 , n29913 , n29914 , n29915 , n29916 , n29917 , n29918 , n29919 , n29920 , n29921 , n29922 , n29923 , n29924 , n29925 , n29926 , n29927 , n29928 , n29929 , n29930 , n29931 , n29932 , n29933 , n29934 , n29935 , n29936 , n29937 , n29938 , n29939 , n29940 , n29941 , n29942 , n29943 , n29944 , n29945 , n29946 , n29947 , n29948 , n29949 , n29950 , n29951 , n29952 , n29953 , n29954 , n29955 , n29956 , n29957 , n29958 , n29959 , n29960 , n29961 , n29962 , n29963 , n29964 , n29965 , n29966 , n29967 , n29968 , n29969 , n29970 , n29971 , n29972 , n29973 , n29974 , n29975 , n29976 , n29977 , n29978 , n29979 , n29980 , n29981 , n29982 , n29983 , n29984 , n29985 , n29986 , n29987 , n29988 , n29989 , n29990 , n29991 , n29992 , n29993 , n29994 , n29995 , n29996 , n29997 , n29998 , n29999 , n30000 , n30001 , n30002 , n30003 , n30004 , n30005 , n30006 , n30007 , n30008 , n30009 , n30010 , n30011 , n30012 , n30013 , n30014 , n30015 , n30016 , n30017 , n30018 , n30019 , n30020 , n30021 , n30022 , n30023 , n30024 , n30025 , n30026 , n30027 , n30028 , n30029 , n30030 , n30031 , n30032 , n30033 , n30034 , n30035 , n30036 , n30037 , n30038 , n30039 , n30040 , n30041 , n30042 , n30043 , n30044 , n30045 , n30046 , n30047 , n30048 , n30049 , n30050 , n30051 , n30052 , n30053 , n30054 , n30055 , n30056 , n30057 , n30058 , n30059 , n30060 , n30061 , n30062 , n30063 , n30064 , n30065 , n30066 , n30067 , n30068 , n30069 , n30070 , n30071 , n30072 , n30073 , n30074 , n30075 , n30076 , n30077 , n30078 , n30079 , n30080 , n30081 , n30082 , n30083 , n30084 , n30085 , n30086 , n30087 , n30088 , n30089 , n30090 , n30091 , n30092 , n30093 , n30094 , n30095 , n30096 , n30097 , n30098 , n30099 , n30100 , n30101 , n30102 , n30103 , n30104 , n30105 , n30106 , n30107 , n30108 , n30109 , n30110 , n30111 , n30112 , n30113 , n30114 , n30115 , n30116 , n30117 , n30118 , n30119 , n30120 , n30121 , n30122 , n30123 , n30124 , n30125 , n30126 , n30127 , n30128 , n30129 , n30130 , n30131 , n30132 , n30133 , n30134 , n30135 , n30136 , n30137 , n30138 , n30139 , n30140 , n30141 , n30142 , n30143 , n30144 , n30145 , n30146 , n30147 , n30148 , n30149 , n30150 , n30151 , n30152 , n30153 , n30154 , n30155 , n30156 , n30157 , n30158 , n30159 , n30160 , n30161 , n30162 , n30163 , n30164 , n30165 , n30166 , n30167 , n30168 , n30169 , n30170 , n30171 , n30172 , n30173 , n30174 , n30175 , n30176 , n30177 , n30178 , n30179 , n30180 , n30181 , n30182 , n30183 , n30184 , n30185 , n30186 , n30187 , n30188 , n30189 , n30190 , n30191 , n30192 , n30193 , n30194 , n30195 , n30196 , n30197 , n30198 , n30199 , n30200 , n30201 , n30202 , n30203 , n30204 , n30205 , n30206 , n30207 , n30208 , n30209 , n30210 , n30211 , n30212 , n30213 , n30214 , n30215 , n30216 , n30217 , n30218 , n30219 , n30220 , n30221 , n30222 , n30223 , n30224 , n30225 , n30226 , n30227 , n30228 , n30229 , n30230 , n30231 , n30232 , n30233 , n30234 , n30235 , n30236 , n30237 , n30238 , n30239 , n30240 , n30241 , n30242 , n30243 , n30244 , n30245 , n30246 , n30247 , n30248 , n30249 , n30250 , n30251 , n30252 , n30253 , n30254 , n30255 , n30256 , n30257 , n30258 , n30259 , n30260 , n30261 , n30262 , n30263 , n30264 , n30265 , n30266 , n30267 , n30268 , n30269 , n30270 , n30271 , n30272 , n30273 , n30274 , n30275 , n30276 , n30277 , n30278 , n30279 , n30280 , n30281 , n30282 , n30283 , n30284 , n30285 , n30286 , n30287 , n30288 , n30289 , n30290 , n30291 , n30292 , n30293 , n30294 , n30295 , n30296 , n30297 , n30298 , n30299 , n30300 , n30301 , n30302 , n30303 , n30304 , n30305 , n30306 , n30307 , n30308 , n30309 , n30310 , n30311 , n30312 , n30313 , n30314 , n30315 , n30316 , n30317 , n30318 , n30319 , n30320 , n30321 , n30322 , n30323 , n30324 , n30325 , n30326 , n30327 , n30328 , n30329 , n30330 , n30331 , n30332 , n30333 , n30334 , n30335 , n30336 , n30337 , n30338 , n30339 , n30340 , n30341 , n30342 , n30343 , n30344 , n30345 , n30346 , n30347 , n30348 , n30349 , n30350 , n30351 , n30352 , n30353 , n30354 , n30355 , n30356 , n30357 , n30358 , n30359 , n30360 , n30361 , n30362 , n30363 , n30364 , n30365 , n30366 , n30367 , n30368 , n30369 , n30370 , n30371 , n30372 , n30373 , n30374 , n30375 , n30376 , n30377 , n30378 , n30379 , n30380 , n30381 , n30382 , n30383 , n30384 , n30385 , n30386 , n30387 , n30388 , n30389 , n30390 , n30391 , n30392 , n30393 , n30394 , n30395 , n30396 , n30397 , n30398 , n30399 , n30400 , n30401 , n30402 , n30403 , n30404 , n30405 , n30406 , n30407 , n30408 , n30409 , n30410 , n30411 , n30412 , n30413 , n30414 , n30415 , n30416 , n30417 , n30418 , n30419 , n30420 , n30421 , n30422 , n30423 , n30424 , n30425 , n30426 , n30427 , n30428 , n30429 , n30430 , n30431 , n30432 , n30433 , n30434 , n30435 , n30436 , n30437 , n30438 , n30439 , n30440 , n30441 , n30442 , n30443 , n30444 , n30445 , n30446 , n30447 , n30448 , n30449 , n30450 , n30451 , n30452 , n30453 , n30454 , n30455 , n30456 , n30457 , n30458 , n30459 , n30460 , n30461 , n30462 , n30463 , n30464 , n30465 , n30466 , n30467 , n30468 , n30469 , n30470 , n30471 , n30472 , n30473 , n30474 , n30475 , n30476 , n30477 , n30478 , n30479 , n30480 , n30481 , n30482 , n30483 , n30484 , n30485 , n30486 , n30487 , n30488 , n30489 , n30490 , n30491 , n30492 , n30493 , n30494 , n30495 , n30496 , n30497 , n30498 , n30499 , n30500 , n30501 , n30502 , n30503 , n30504 , n30505 , n30506 , n30507 , n30508 , n30509 , n30510 , n30511 , n30512 , n30513 , n30514 , n30515 , n30516 , n30517 , n30518 , n30519 , n30520 , n30521 , n30522 , n30523 , n30524 , n30525 , n30526 , n30527 , n30528 , n30529 , n30530 , n30531 , n30532 , n30533 , n30534 , n30535 , n30536 , n30537 , n30538 , n30539 , n30540 , n30541 , n30542 , n30543 , n30544 , n30545 , n30546 , n30547 , n30548 , n30549 , n30550 , n30551 , n30552 , n30553 , n30554 , n30555 , n30556 , n30557 , n30558 , n30559 , n30560 , n30561 , n30562 , n30563 , n30564 , n30565 , n30566 , n30567 , n30568 , n30569 , n30570 , n30571 , n30572 , n30573 , n30574 , n30575 , n30576 , n30577 , n30578 , n30579 , n30580 , n30581 , n30582 , n30583 , n30584 , n30585 , n30586 , n30587 , n30588 , n30589 , n30590 , n30591 , n30592 , n30593 , n30594 , n30595 , n30596 , n30597 , n30598 , n30599 , n30600 , n30601 , n30602 , n30603 , n30604 , n30605 , n30606 , n30607 , n30608 , n30609 , n30610 , n30611 , n30612 , n30613 , n30614 , n30615 , n30616 , n30617 , n30618 , n30619 , n30620 , n30621 , n30622 , n30623 , n30624 , n30625 , n30626 , n30627 , n30628 , n30629 , n30630 , n30631 , n30632 , n30633 , n30634 , n30635 , n30636 , n30637 , n30638 , n30639 , n30640 , n30641 , n30642 , n30643 , n30644 , n30645 , n30646 , n30647 , n30648 , n30649 , n30650 , n30651 , n30652 , n30653 , n30654 , n30655 , n30656 , n30657 , n30658 , n30659 , n30660 , n30661 , n30662 , n30663 , n30664 , n30665 , n30666 , n30667 , n30668 , n30669 , n30670 , n30671 , n30672 , n30673 , n30674 , n30675 , n30676 , n30677 , n30678 , n30679 , n30680 , n30681 , n30682 , n30683 , n30684 , n30685 , n30686 , n30687 , n30688 , n30689 , n30690 , n30691 , n30692 , n30693 , n30694 , n30695 , n30696 , n30697 , n30698 , n30699 , n30700 , n30701 , n30702 , n30703 , n30704 , n30705 , n30706 , n30707 , n30708 , n30709 , n30710 , n30711 , n30712 , n30713 , n30714 , n30715 , n30716 , n30717 , n30718 , n30719 , n30720 , n30721 , n30722 , n30723 , n30724 , n30725 , n30726 , n30727 , n30728 , n30729 , n30730 , n30731 , n30732 , n30733 , n30734 , n30735 , n30736 , n30737 , n30738 , n30739 , n30740 , n30741 , n30742 , n30743 , n30744 , n30745 , n30746 , n30747 , n30748 , n30749 , n30750 , n30751 , n30752 , n30753 , n30754 , n30755 , n30756 , n30757 , n30758 , n30759 , n30760 , n30761 , n30762 , n30763 , n30764 , n30765 , n30766 , n30767 , n30768 , n30769 , n30770 , n30771 , n30772 , n30773 , n30774 , n30775 , n30776 , n30777 , n30778 , n30779 , n30780 , n30781 , n30782 , n30783 , n30784 , n30785 , n30786 , n30787 , n30788 , n30789 , n30790 , n30791 , n30792 , n30793 , n30794 , n30795 , n30796 , n30797 , n30798 , n30799 , n30800 , n30801 , n30802 , n30803 , n30804 , n30805 , n30806 , n30807 , n30808 , n30809 , n30810 , n30811 , n30812 , n30813 , n30814 , n30815 , n30816 , n30817 , n30818 , n30819 , n30820 , n30821 , n30822 , n30823 , n30824 , n30825 , n30826 , n30827 , n30828 , n30829 , n30830 , n30831 , n30832 , n30833 , n30834 , n30835 , n30836 , n30837 , n30838 , n30839 , n30840 , n30841 , n30842 , n30843 , n30844 , n30845 , n30846 , n30847 , n30848 , n30849 , n30850 , n30851 , n30852 , n30853 , n30854 , n30855 , n30856 , n30857 , n30858 , n30859 , n30860 , n30861 , n30862 , n30863 , n30864 , n30865 , n30866 , n30867 , n30868 , n30869 , n30870 , n30871 , n30872 , n30873 , n30874 , n30875 , n30876 , n30877 , n30878 , n30879 , n30880 , n30881 , n30882 , n30883 , n30884 , n30885 , n30886 , n30887 , n30888 , n30889 , n30890 , n30891 , n30892 , n30893 , n30894 , n30895 , n30896 , n30897 , n30898 , n30899 , n30900 , n30901 , n30902 , n30903 , n30904 , n30905 , n30906 , n30907 , n30908 , n30909 , n30910 , n30911 , n30912 , n30913 , n30914 , n30915 , n30916 , n30917 , n30918 , n30919 , n30920 , n30921 , n30922 , n30923 , n30924 , n30925 , n30926 , n30927 , n30928 , n30929 , n30930 , n30931 , n30932 , n30933 , n30934 , n30935 , n30936 , n30937 , n30938 , n30939 , n30940 , n30941 , n30942 , n30943 , n30944 , n30945 , n30946 , n30947 , n30948 , n30949 , n30950 , n30951 , n30952 , n30953 , n30954 , n30955 , n30956 , n30957 , n30958 , n30959 , n30960 , n30961 , n30962 , n30963 , n30964 , n30965 , n30966 , n30967 , n30968 , n30969 , n30970 , n30971 , n30972 , n30973 , n30974 , n30975 , n30976 , n30977 , n30978 , n30979 , n30980 , n30981 , n30982 , n30983 , n30984 , n30985 , n30986 , n30987 , n30988 , n30989 , n30990 , n30991 , n30992 , n30993 , n30994 , n30995 , n30996 , n30997 , n30998 , n30999 , n31000 , n31001 , n31002 , n31003 , n31004 , n31005 , n31006 , n31007 , n31008 , n31009 , n31010 , n31011 , n31012 , n31013 , n31014 , n31015 , n31016 , n31017 , n31018 , n31019 , n31020 , n31021 , n31022 , n31023 , n31024 , n31025 , n31026 , n31027 , n31028 , n31029 , n31030 , n31031 , n31032 , n31033 , n31034 , n31035 , n31036 , n31037 , n31038 , n31039 , n31040 , n31041 , n31042 , n31043 , n31044 , n31045 , n31046 , n31047 , n31048 , n31049 , n31050 , n31051 , n31052 , n31053 , n31054 , n31055 , n31056 , n31057 , n31058 , n31059 , n31060 , n31061 , n31062 , n31063 , n31064 , n31065 , n31066 , n31067 , n31068 , n31069 , n31070 , n31071 , n31072 , n31073 , n31074 , n31075 , n31076 , n31077 , n31078 , n31079 , n31080 , n31081 , n31082 , n31083 , n31084 , n31085 , n31086 , n31087 , n31088 , n31089 , n31090 , n31091 , n31092 , n31093 , n31094 , n31095 , n31096 , n31097 , n31098 , n31099 , n31100 , n31101 , n31102 , n31103 , n31104 , n31105 , n31106 , n31107 , n31108 , n31109 , n31110 , n31111 , n31112 , n31113 , n31114 , n31115 , n31116 , n31117 , n31118 , n31119 , n31120 , n31121 , n31122 , n31123 , n31124 , n31125 , n31126 , n31127 , n31128 , n31129 , n31130 , n31131 , n31132 , n31133 , n31134 , n31135 , n31136 , n31137 , n31138 , n31139 , n31140 , n31141 , n31142 , n31143 , n31144 , n31145 , n31146 , n31147 , n31148 , n31149 , n31150 , n31151 , n31152 , n31153 , n31154 , n31155 , n31156 , n31157 , n31158 , n31159 , n31160 , n31161 , n31162 , n31163 , n31164 , n31165 , n31166 , n31167 , n31168 , n31169 , n31170 , n31171 , n31172 , n31173 , n31174 , n31175 , n31176 , n31177 , n31178 , n31179 , n31180 , n31181 , n31182 , n31183 , n31184 , n31185 , n31186 , n31187 , n31188 , n31189 , n31190 , n31191 , n31192 , n31193 , n31194 , n31195 , n31196 , n31197 , n31198 , n31199 , n31200 , n31201 , n31202 , n31203 , n31204 , n31205 , n31206 , n31207 , n31208 , n31209 , n31210 , n31211 , n31212 , n31213 , n31214 , n31215 , n31216 , n31217 , n31218 , n31219 , n31220 , n31221 , n31222 , n31223 , n31224 , n31225 , n31226 , n31227 , n31228 , n31229 , n31230 , n31231 , n31232 , n31233 , n31234 , n31235 , n31236 , n31237 , n31238 , n31239 , n31240 , n31241 , n31242 , n31243 , n31244 , n31245 , n31246 , n31247 , n31248 , n31249 , n31250 , n31251 , n31252 , n31253 , n31254 , n31255 , n31256 , n31257 , n31258 , n31259 , n31260 , n31261 , n31262 , n31263 , n31264 , n31265 , n31266 , n31267 , n31268 , n31269 , n31270 , n31271 , n31272 , n31273 , n31274 , n31275 , n31276 , n31277 , n31278 , n31279 , n31280 , n31281 , n31282 , n31283 , n31284 , n31285 , n31286 , n31287 , n31288 , n31289 , n31290 , n31291 , n31292 , n31293 , n31294 , n31295 , n31296 , n31297 , n31298 , n31299 , n31300 , n31301 , n31302 , n31303 , n31304 , n31305 , n31306 , n31307 , n31308 , n31309 , n31310 , n31311 , n31312 , n31313 , n31314 , n31315 , n31316 , n31317 , n31318 , n31319 , n31320 , n31321 , n31322 , n31323 , n31324 , n31325 , n31326 , n31327 , n31328 , n31329 , n31330 , n31331 , n31332 , n31333 , n31334 , n31335 , n31336 , n31337 , n31338 , n31339 , n31340 , n31341 , n31342 , n31343 , n31344 , n31345 , n31346 , n31347 , n31348 , n31349 , n31350 , n31351 , n31352 , n31353 , n31354 , n31355 , n31356 , n31357 , n31358 , n31359 , n31360 , n31361 , n31362 , n31363 , n31364 , n31365 , n31366 , n31367 , n31368 , n31369 , n31370 , n31371 , n31372 , n31373 , n31374 , n31375 , n31376 , n31377 , n31378 , n31379 , n31380 , n31381 , n31382 , n31383 , n31384 , n31385 , n31386 , n31387 , n31388 , n31389 , n31390 , n31391 , n31392 , n31393 , n31394 , n31395 , n31396 , n31397 , n31398 , n31399 , n31400 , n31401 , n31402 , n31403 , n31404 , n31405 , n31406 , n31407 , n31408 , n31409 , n31410 , n31411 , n31412 , n31413 , n31414 , n31415 , n31416 , n31417 , n31418 , n31419 , n31420 , n31421 , n31422 , n31423 , n31424 , n31425 , n31426 , n31427 , n31428 , n31429 , n31430 , n31431 , n31432 , n31433 , n31434 , n31435 , n31436 , n31437 , n31438 , n31439 , n31440 , n31441 , n31442 , n31443 , n31444 , n31445 , n31446 , n31447 , n31448 , n31449 , n31450 , n31451 , n31452 , n31453 , n31454 , n31455 , n31456 , n31457 , n31458 , n31459 , n31460 , n31461 , n31462 , n31463 , n31464 , n31465 , n31466 , n31467 , n31468 , n31469 , n31470 , n31471 , n31472 , n31473 , n31474 , n31475 , n31476 , n31477 , n31478 , n31479 , n31480 , n31481 , n31482 , n31483 , n31484 , n31485 , n31486 , n31487 , n31488 , n31489 , n31490 , n31491 , n31492 , n31493 , n31494 , n31495 , n31496 , n31497 , n31498 , n31499 , n31500 , n31501 , n31502 , n31503 , n31504 , n31505 , n31506 , n31507 , n31508 , n31509 , n31510 , n31511 , n31512 , n31513 , n31514 , n31515 , n31516 , n31517 , n31518 , n31519 , n31520 , n31521 , n31522 , n31523 , n31524 , n31525 , n31526 , n31527 , n31528 , n31529 , n31530 , n31531 , n31532 , n31533 , n31534 , n31535 , n31536 , n31537 , n31538 , n31539 , n31540 , n31541 , n31542 , n31543 , n31544 , n31545 , n31546 , n31547 , n31548 , n31549 , n31550 , n31551 , n31552 , n31553 , n31554 , n31555 , n31556 , n31557 , n31558 , n31559 , n31560 , n31561 , n31562 , n31563 , n31564 , n31565 , n31566 , n31567 , n31568 , n31569 , n31570 , n31571 , n31572 , n31573 , n31574 , n31575 , n31576 , n31577 , n31578 , n31579 , n31580 , n31581 , n31582 , n31583 , n31584 , n31585 , n31586 , n31587 , n31588 , n31589 , n31590 , n31591 , n31592 , n31593 , n31594 , n31595 , n31596 , n31597 , n31598 , n31599 , n31600 , n31601 , n31602 , n31603 , n31604 , n31605 , n31606 , n31607 , n31608 , n31609 , n31610 , n31611 , n31612 , n31613 , n31614 , n31615 , n31616 , n31617 , n31618 , n31619 , n31620 , n31621 , n31622 , n31623 , n31624 , n31625 , n31626 , n31627 , n31628 , n31629 , n31630 , n31631 , n31632 , n31633 , n31634 , n31635 , n31636 , n31637 , n31638 , n31639 , n31640 , n31641 , n31642 , n31643 , n31644 , n31645 , n31646 , n31647 , n31648 , n31649 , n31650 , n31651 , n31652 , n31653 , n31654 , n31655 , n31656 , n31657 , n31658 , n31659 , n31660 , n31661 , n31662 , n31663 , n31664 , n31665 , n31666 , n31667 , n31668 , n31669 , n31670 , n31671 , n31672 , n31673 , n31674 , n31675 , n31676 , n31677 , n31678 , n31679 , n31680 , n31681 , n31682 , n31683 , n31684 , n31685 , n31686 , n31687 , n31688 , n31689 , n31690 , n31691 , n31692 , n31693 , n31694 , n31695 , n31696 , n31697 , n31698 , n31699 , n31700 , n31701 , n31702 , n31703 , n31704 , n31705 , n31706 , n31707 , n31708 , n31709 , n31710 , n31711 , n31712 , n31713 , n31714 , n31715 , n31716 , n31717 , n31718 , n31719 , n31720 , n31721 , n31722 , n31723 , n31724 , n31725 , n31726 , n31727 , n31728 , n31729 , n31730 , n31731 , n31732 , n31733 , n31734 , n31735 , n31736 , n31737 , n31738 , n31739 , n31740 , n31741 , n31742 , n31743 , n31744 , n31745 , n31746 , n31747 , n31748 , n31749 , n31750 , n31751 , n31752 , n31753 , n31754 , n31755 , n31756 , n31757 , n31758 , n31759 , n31760 , n31761 , n31762 , n31763 , n31764 , n31765 , n31766 , n31767 , n31768 , n31769 , n31770 , n31771 , n31772 , n31773 , n31774 , n31775 , n31776 , n31777 , n31778 , n31779 , n31780 , n31781 , n31782 , n31783 , n31784 , n31785 , n31786 , n31787 , n31788 , n31789 , n31790 , n31791 , n31792 , n31793 , n31794 , n31795 , n31796 , n31797 , n31798 , n31799 , n31800 , n31801 , n31802 , n31803 , n31804 , n31805 , n31806 , n31807 , n31808 , n31809 , n31810 , n31811 , n31812 , n31813 , n31814 , n31815 , n31816 , n31817 , n31818 , n31819 , n31820 , n31821 , n31822 , n31823 , n31824 , n31825 , n31826 , n31827 , n31828 , n31829 , n31830 , n31831 , n31832 , n31833 , n31834 , n31835 , n31836 , n31837 , n31838 , n31839 , n31840 , n31841 , n31842 , n31843 , n31844 , n31845 , n31846 , n31847 , n31848 , n31849 , n31850 , n31851 , n31852 , n31853 , n31854 , n31855 , n31856 , n31857 , n31858 , n31859 , n31860 , n31861 , n31862 , n31863 , n31864 , n31865 , n31866 , n31867 , n31868 , n31869 , n31870 , n31871 , n31872 , n31873 , n31874 , n31875 , n31876 , n31877 , n31878 , n31879 , n31880 , n31881 , n31882 , n31883 , n31884 , n31885 , n31886 , n31887 , n31888 , n31889 , n31890 , n31891 , n31892 , n31893 , n31894 , n31895 , n31896 , n31897 , n31898 , n31899 , n31900 , n31901 , n31902 , n31903 , n31904 , n31905 , n31906 , n31907 , n31908 , n31909 , n31910 , n31911 , n31912 , n31913 , n31914 , n31915 , n31916 , n31917 , n31918 , n31919 , n31920 , n31921 , n31922 , n31923 , n31924 , n31925 , n31926 , n31927 , n31928 , n31929 , n31930 , n31931 , n31932 , n31933 , n31934 , n31935 , n31936 , n31937 , n31938 , n31939 , n31940 , n31941 , n31942 , n31943 , n31944 , n31945 , n31946 , n31947 , n31948 , n31949 , n31950 , n31951 , n31952 , n31953 , n31954 , n31955 , n31956 , n31957 , n31958 , n31959 , n31960 , n31961 , n31962 , n31963 , n31964 , n31965 , n31966 , n31967 , n31968 , n31969 , n31970 , n31971 , n31972 , n31973 , n31974 , n31975 , n31976 , n31977 , n31978 , n31979 , n31980 , n31981 , n31982 , n31983 , n31984 , n31985 , n31986 , n31987 , n31988 , n31989 , n31990 , n31991 , n31992 , n31993 , n31994 , n31995 , n31996 , n31997 , n31998 , n31999 , n32000 , n32001 , n32002 , n32003 , n32004 , n32005 , n32006 , n32007 , n32008 , n32009 , n32010 , n32011 , n32012 , n32013 , n32014 , n32015 , n32016 , n32017 , n32018 , n32019 , n32020 , n32021 , n32022 , n32023 , n32024 , n32025 , n32026 , n32027 , n32028 , n32029 , n32030 , n32031 , n32032 , n32033 , n32034 , n32035 , n32036 , n32037 , n32038 , n32039 , n32040 , n32041 , n32042 , n32043 , n32044 , n32045 , n32046 , n32047 , n32048 , n32049 , n32050 , n32051 , n32052 , n32053 , n32054 , n32055 , n32056 , n32057 , n32058 , n32059 , n32060 , n32061 , n32062 , n32063 , n32064 , n32065 , n32066 , n32067 , n32068 , n32069 , n32070 , n32071 , n32072 , n32073 , n32074 , n32075 , n32076 , n32077 , n32078 , n32079 , n32080 , n32081 , n32082 , n32083 , n32084 , n32085 , n32086 , n32087 , n32088 , n32089 , n32090 , n32091 , n32092 , n32093 , n32094 , n32095 , n32096 , n32097 , n32098 , n32099 , n32100 , n32101 , n32102 , n32103 , n32104 , n32105 , n32106 , n32107 , n32108 , n32109 , n32110 , n32111 , n32112 , n32113 , n32114 , n32115 , n32116 , n32117 , n32118 , n32119 , n32120 , n32121 , n32122 , n32123 , n32124 , n32125 , n32126 , n32127 , n32128 , n32129 , n32130 , n32131 , n32132 , n32133 , n32134 , n32135 , n32136 , n32137 , n32138 , n32139 , n32140 , n32141 , n32142 , n32143 , n32144 , n32145 , n32146 , n32147 , n32148 , n32149 , n32150 , n32151 , n32152 , n32153 , n32154 , n32155 , n32156 , n32157 , n32158 , n32159 , n32160 , n32161 , n32162 , n32163 , n32164 , n32165 , n32166 , n32167 , n32168 , n32169 , n32170 , n32171 , n32172 , n32173 , n32174 , n32175 , n32176 , n32177 , n32178 , n32179 , n32180 , n32181 , n32182 , n32183 , n32184 , n32185 , n32186 , n32187 , n32188 , n32189 , n32190 , n32191 , n32192 , n32193 , n32194 , n32195 , n32196 , n32197 , n32198 , n32199 , n32200 , n32201 , n32202 , n32203 , n32204 , n32205 , n32206 , n32207 , n32208 , n32209 , n32210 , n32211 , n32212 , n32213 , n32214 , n32215 , n32216 , n32217 , n32218 , n32219 , n32220 , n32221 , n32222 , n32223 , n32224 , n32225 , n32226 , n32227 , n32228 , n32229 , n32230 , n32231 , n32232 , n32233 , n32234 , n32235 , n32236 , n32237 , n32238 , n32239 , n32240 , n32241 , n32242 , n32243 , n32244 , n32245 , n32246 , n32247 , n32248 , n32249 , n32250 , n32251 , n32252 , n32253 , n32254 , n32255 , n32256 , n32257 , n32258 , n32259 , n32260 , n32261 , n32262 , n32263 , n32264 , n32265 , n32266 , n32267 , n32268 , n32269 , n32270 , n32271 , n32272 , n32273 , n32274 , n32275 , n32276 , n32277 , n32278 , n32279 , n32280 , n32281 , n32282 , n32283 , n32284 , n32285 , n32286 , n32287 , n32288 , n32289 , n32290 , n32291 , n32292 , n32293 , n32294 , n32295 , n32296 , n32297 , n32298 , n32299 , n32300 , n32301 , n32302 , n32303 , n32304 , n32305 , n32306 , n32307 , n32308 , n32309 , n32310 , n32311 , n32312 , n32313 , n32314 , n32315 , n32316 , n32317 , n32318 , n32319 , n32320 , n32321 , n32322 , n32323 , n32324 , n32325 , n32326 , n32327 , n32328 , n32329 , n32330 , n32331 , n32332 , n32333 , n32334 , n32335 , n32336 , n32337 , n32338 , n32339 , n32340 , n32341 , n32342 , n32343 , n32344 , n32345 , n32346 , n32347 , n32348 , n32349 , n32350 , n32351 , n32352 , n32353 , n32354 , n32355 , n32356 , n32357 , n32358 , n32359 , n32360 , n32361 , n32362 , n32363 , n32364 , n32365 , n32366 , n32367 , n32368 , n32369 , n32370 , n32371 , n32372 , n32373 , n32374 , n32375 , n32376 , n32377 , n32378 , n32379 , n32380 , n32381 , n32382 , n32383 , n32384 , n32385 , n32386 , n32387 , n32388 , n32389 , n32390 , n32391 , n32392 , n32393 , n32394 , n32395 , n32396 , n32397 , n32398 , n32399 , n32400 , n32401 , n32402 , n32403 , n32404 , n32405 , n32406 , n32407 , n32408 , n32409 , n32410 , n32411 , n32412 , n32413 , n32414 , n32415 , n32416 , n32417 , n32418 , n32419 , n32420 , n32421 , n32422 , n32423 , n32424 , n32425 , n32426 , n32427 , n32428 , n32429 , n32430 , n32431 , n32432 , n32433 , n32434 , n32435 , n32436 , n32437 , n32438 , n32439 , n32440 , n32441 , n32442 , n32443 , n32444 , n32445 , n32446 , n32447 , n32448 , n32449 , n32450 , n32451 , n32452 , n32453 , n32454 , n32455 , n32456 , n32457 , n32458 , n32459 , n32460 , n32461 , n32462 , n32463 , n32464 , n32465 , n32466 , n32467 , n32468 , n32469 , n32470 , n32471 , n32472 , n32473 , n32474 , n32475 , n32476 , n32477 , n32478 , n32479 , n32480 , n32481 , n32482 , n32483 , n32484 , n32485 , n32486 , n32487 , n32488 , n32489 , n32490 , n32491 , n32492 , n32493 , n32494 , n32495 , n32496 , n32497 , n32498 , n32499 , n32500 , n32501 , n32502 , n32503 , n32504 , n32505 , n32506 , n32507 , n32508 , n32509 , n32510 , n32511 , n32512 , n32513 , n32514 , n32515 , n32516 , n32517 , n32518 , n32519 , n32520 , n32521 , n32522 , n32523 , n32524 , n32525 , n32526 , n32527 , n32528 , n32529 , n32530 , n32531 , n32532 , n32533 , n32534 , n32535 , n32536 , n32537 , n32538 , n32539 , n32540 , n32541 , n32542 , n32543 , n32544 , n32545 , n32546 , n32547 , n32548 , n32549 , n32550 , n32551 , n32552 , n32553 , n32554 , n32555 , n32556 , n32557 , n32558 , n32559 , n32560 , n32561 , n32562 , n32563 , n32564 , n32565 , n32566 , n32567 , n32568 , n32569 , n32570 , n32571 , n32572 , n32573 , n32574 , n32575 , n32576 , n32577 , n32578 , n32579 , n32580 , n32581 , n32582 , n32583 , n32584 , n32585 , n32586 , n32587 , n32588 , n32589 , n32590 , n32591 , n32592 , n32593 , n32594 , n32595 , n32596 , n32597 , n32598 , n32599 , n32600 , n32601 , n32602 , n32603 , n32604 , n32605 , n32606 , n32607 , n32608 , n32609 , n32610 , n32611 , n32612 , n32613 , n32614 , n32615 , n32616 , n32617 , n32618 , n32619 , n32620 , n32621 , n32622 , n32623 , n32624 , n32625 , n32626 , n32627 , n32628 , n32629 , n32630 , n32631 , n32632 , n32633 , n32634 , n32635 , n32636 , n32637 , n32638 , n32639 , n32640 , n32641 , n32642 , n32643 , n32644 , n32645 , n32646 , n32647 , n32648 , n32649 , n32650 , n32651 , n32652 , n32653 , n32654 , n32655 , n32656 , n32657 , n32658 , n32659 , n32660 , n32661 , n32662 , n32663 , n32664 , n32665 , n32666 , n32667 , n32668 , n32669 , n32670 , n32671 , n32672 , n32673 , n32674 , n32675 , n32676 , n32677 , n32678 , n32679 , n32680 , n32681 , n32682 , n32683 , n32684 , n32685 , n32686 , n32687 , n32688 , n32689 , n32690 , n32691 , n32692 , n32693 , n32694 , n32695 , n32696 , n32697 , n32698 , n32699 , n32700 , n32701 , n32702 , n32703 , n32704 , n32705 , n32706 , n32707 , n32708 , n32709 , n32710 , n32711 , n32712 , n32713 , n32714 , n32715 , n32716 , n32717 , n32718 , n32719 , n32720 , n32721 , n32722 , n32723 , n32724 , n32725 , n32726 , n32727 , n32728 , n32729 , n32730 , n32731 , n32732 , n32733 , n32734 , n32735 , n32736 , n32737 , n32738 , n32739 , n32740 , n32741 , n32742 , n32743 , n32744 , n32745 , n32746 , n32747 , n32748 , n32749 , n32750 , n32751 , n32752 , n32753 , n32754 , n32755 , n32756 , n32757 , n32758 , n32759 , n32760 , n32761 , n32762 , n32763 , n32764 , n32765 , n32766 , n32767 , n32768 , n32769 , n32770 , n32771 , n32772 , n32773 , n32774 , n32775 , n32776 , n32777 , n32778 , n32779 , n32780 , n32781 , n32782 , n32783 , n32784 , n32785 , n32786 , n32787 , n32788 , n32789 , n32790 , n32791 , n32792 , n32793 , n32794 , n32795 , n32796 , n32797 , n32798 , n32799 , n32800 , n32801 , n32802 , n32803 , n32804 , n32805 , n32806 , n32807 , n32808 , n32809 , n32810 , n32811 , n32812 , n32813 , n32814 , n32815 , n32816 , n32817 , n32818 , n32819 , n32820 , n32821 , n32822 , n32823 , n32824 , n32825 , n32826 , n32827 , n32828 , n32829 , n32830 , n32831 , n32832 , n32833 , n32834 , n32835 , n32836 , n32837 , n32838 , n32839 , n32840 , n32841 , n32842 , n32843 , n32844 , n32845 , n32846 , n32847 , n32848 , n32849 , n32850 , n32851 , n32852 , n32853 , n32854 , n32855 , n32856 , n32857 , n32858 , n32859 , n32860 , n32861 , n32862 , n32863 , n32864 , n32865 , n32866 , n32867 , n32868 , n32869 , n32870 , n32871 , n32872 , n32873 , n32874 , n32875 , n32876 , n32877 , n32878 , n32879 , n32880 , n32881 , n32882 , n32883 , n32884 , n32885 , n32886 , n32887 , n32888 , n32889 , n32890 , n32891 , n32892 , n32893 , n32894 , n32895 , n32896 , n32897 , n32898 , n32899 , n32900 , n32901 , n32902 , n32903 , n32904 , n32905 , n32906 , n32907 , n32908 , n32909 , n32910 , n32911 , n32912 , n32913 , n32914 , n32915 , n32916 , n32917 , n32918 , n32919 , n32920 , n32921 , n32922 , n32923 , n32924 , n32925 , n32926 , n32927 , n32928 , n32929 , n32930 , n32931 , n32932 , n32933 , n32934 , n32935 , n32936 , n32937 , n32938 , n32939 , n32940 , n32941 , n32942 , n32943 , n32944 , n32945 , n32946 , n32947 , n32948 , n32949 , n32950 , n32951 , n32952 , n32953 , n32954 , n32955 , n32956 , n32957 , n32958 , n32959 , n32960 , n32961 , n32962 , n32963 , n32964 , n32965 , n32966 , n32967 , n32968 , n32969 , n32970 , n32971 , n32972 , n32973 , n32974 , n32975 , n32976 , n32977 , n32978 , n32979 , n32980 , n32981 , n32982 , n32983 , n32984 , n32985 , n32986 , n32987 , n32988 , n32989 , n32990 , n32991 , n32992 , n32993 , n32994 , n32995 , n32996 , n32997 , n32998 , n32999 , n33000 , n33001 , n33002 , n33003 , n33004 , n33005 , n33006 , n33007 , n33008 , n33009 , n33010 , n33011 , n33012 , n33013 , n33014 , n33015 , n33016 , n33017 , n33018 , n33019 , n33020 , n33021 , n33022 , n33023 , n33024 , n33025 , n33026 , n33027 , n33028 , n33029 , n33030 , n33031 , n33032 , n33033 , n33034 , n33035 , n33036 , n33037 , n33038 , n33039 , n33040 , n33041 , n33042 , n33043 , n33044 , n33045 , n33046 , n33047 , n33048 , n33049 , n33050 , n33051 , n33052 , n33053 , n33054 , n33055 , n33056 , n33057 , n33058 , n33059 , n33060 , n33061 , n33062 , n33063 , n33064 , n33065 , n33066 , n33067 , n33068 , n33069 , n33070 , n33071 , n33072 , n33073 , n33074 , n33075 , n33076 , n33077 , n33078 , n33079 , n33080 , n33081 , n33082 , n33083 , n33084 , n33085 , n33086 , n33087 , n33088 , n33089 , n33090 , n33091 , n33092 , n33093 , n33094 , n33095 , n33096 , n33097 , n33098 , n33099 , n33100 , n33101 , n33102 , n33103 , n33104 , n33105 , n33106 , n33107 , n33108 , n33109 , n33110 , n33111 , n33112 , n33113 , n33114 , n33115 , n33116 , n33117 , n33118 , n33119 , n33120 , n33121 , n33122 , n33123 , n33124 , n33125 , n33126 , n33127 , n33128 , n33129 , n33130 , n33131 , n33132 , n33133 , n33134 , n33135 , n33136 , n33137 , n33138 , n33139 , n33140 , n33141 , n33142 , n33143 , n33144 , n33145 , n33146 , n33147 , n33148 , n33149 , n33150 , n33151 , n33152 , n33153 , n33154 , n33155 , n33156 , n33157 , n33158 , n33159 , n33160 , n33161 , n33162 , n33163 , n33164 , n33165 , n33166 , n33167 , n33168 , n33169 , n33170 , n33171 , n33172 , n33173 , n33174 , n33175 , n33176 , n33177 , n33178 , n33179 , n33180 , n33181 , n33182 , n33183 , n33184 , n33185 , n33186 , n33187 , n33188 , n33189 , n33190 , n33191 , n33192 , n33193 , n33194 , n33195 , n33196 , n33197 , n33198 , n33199 , n33200 , n33201 , n33202 , n33203 , n33204 , n33205 , n33206 , n33207 , n33208 , n33209 , n33210 , n33211 , n33212 , n33213 , n33214 , n33215 , n33216 , n33217 , n33218 , n33219 , n33220 , n33221 , n33222 , n33223 , n33224 , n33225 , n33226 , n33227 , n33228 , n33229 , n33230 , n33231 , n33232 , n33233 , n33234 , n33235 , n33236 , n33237 , n33238 , n33239 , n33240 , n33241 , n33242 , n33243 , n33244 , n33245 , n33246 , n33247 , n33248 , n33249 , n33250 , n33251 , n33252 , n33253 , n33254 , n33255 , n33256 , n33257 , n33258 , n33259 , n33260 , n33261 , n33262 , n33263 , n33264 , n33265 , n33266 , n33267 , n33268 , n33269 , n33270 , n33271 , n33272 , n33273 , n33274 , n33275 , n33276 , n33277 , n33278 , n33279 , n33280 , n33281 , n33282 , n33283 , n33284 , n33285 , n33286 , n33287 , n33288 , n33289 , n33290 , n33291 , n33292 , n33293 , n33294 , n33295 , n33296 , n33297 , n33298 , n33299 , n33300 , n33301 , n33302 , n33303 , n33304 , n33305 , n33306 , n33307 , n33308 , n33309 , n33310 , n33311 , n33312 , n33313 , n33314 , n33315 , n33316 , n33317 , n33318 , n33319 , n33320 , n33321 , n33322 , n33323 , n33324 , n33325 , n33326 , n33327 , n33328 , n33329 , n33330 , n33331 , n33332 , n33333 , n33334 , n33335 , n33336 , n33337 , n33338 , n33339 , n33340 , n33341 , n33342 , n33343 , n33344 , n33345 , n33346 , n33347 , n33348 , n33349 , n33350 , n33351 , n33352 , n33353 , n33354 , n33355 , n33356 , n33357 , n33358 , n33359 , n33360 , n33361 , n33362 , n33363 , n33364 , n33365 , n33366 , n33367 , n33368 , n33369 , n33370 , n33371 , n33372 , n33373 , n33374 , n33375 , n33376 , n33377 , n33378 , n33379 , n33380 , n33381 , n33382 , n33383 , n33384 , n33385 , n33386 , n33387 , n33388 , n33389 , n33390 , n33391 , n33392 , n33393 , n33394 , n33395 , n33396 , n33397 , n33398 , n33399 , n33400 , n33401 , n33402 , n33403 , n33404 , n33405 , n33406 , n33407 , n33408 , n33409 , n33410 , n33411 , n33412 , n33413 , n33414 , n33415 , n33416 , n33417 , n33418 , n33419 , n33420 , n33421 , n33422 , n33423 , n33424 , n33425 , n33426 , n33427 , n33428 , n33429 , n33430 , n33431 , n33432 , n33433 , n33434 , n33435 , n33436 , n33437 , n33438 , n33439 , n33440 , n33441 , n33442 , n33443 , n33444 , n33445 , n33446 , n33447 , n33448 , n33449 , n33450 , n33451 , n33452 , n33453 , n33454 , n33455 , n33456 , n33457 , n33458 , n33459 , n33460 , n33461 , n33462 , n33463 , n33464 , n33465 , n33466 , n33467 , n33468 , n33469 , n33470 , n33471 , n33472 , n33473 , n33474 , n33475 , n33476 , n33477 , n33478 , n33479 , n33480 , n33481 , n33482 , n33483 , n33484 , n33485 , n33486 , n33487 , n33488 , n33489 , n33490 , n33491 , n33492 , n33493 , n33494 , n33495 , n33496 , n33497 , n33498 , n33499 , n33500 , n33501 , n33502 , n33503 , n33504 , n33505 , n33506 , n33507 , n33508 , n33509 , n33510 , n33511 , n33512 , n33513 , n33514 , n33515 , n33516 , n33517 , n33518 , n33519 , n33520 , n33521 , n33522 , n33523 , n33524 , n33525 , n33526 , n33527 , n33528 , n33529 , n33530 , n33531 , n33532 , n33533 , n33534 , n33535 , n33536 , n33537 , n33538 , n33539 , n33540 , n33541 , n33542 , n33543 , n33544 , n33545 , n33546 , n33547 , n33548 , n33549 , n33550 , n33551 , n33552 , n33553 , n33554 , n33555 , n33556 , n33557 , n33558 , n33559 , n33560 , n33561 , n33562 , n33563 , n33564 , n33565 , n33566 , n33567 , n33568 , n33569 , n33570 , n33571 , n33572 , n33573 , n33574 , n33575 , n33576 , n33577 , n33578 , n33579 , n33580 , n33581 , n33582 , n33583 , n33584 , n33585 , n33586 , n33587 , n33588 , n33589 , n33590 , n33591 , n33592 , n33593 , n33594 , n33595 , n33596 , n33597 , n33598 , n33599 , n33600 , n33601 , n33602 , n33603 , n33604 , n33605 , n33606 , n33607 , n33608 , n33609 , n33610 , n33611 , n33612 , n33613 , n33614 , n33615 , n33616 , n33617 , n33618 , n33619 , n33620 , n33621 , n33622 , n33623 , n33624 , n33625 , n33626 , n33627 , n33628 , n33629 , n33630 , n33631 , n33632 , n33633 , n33634 , n33635 , n33636 , n33637 , n33638 , n33639 , n33640 , n33641 , n33642 , n33643 , n33644 , n33645 , n33646 , n33647 , n33648 , n33649 , n33650 , n33651 , n33652 , n33653 , n33654 , n33655 , n33656 , n33657 , n33658 , n33659 , n33660 , n33661 , n33662 , n33663 , n33664 , n33665 , n33666 , n33667 , n33668 , n33669 , n33670 , n33671 , n33672 , n33673 , n33674 , n33675 , n33676 , n33677 , n33678 , n33679 , n33680 , n33681 , n33682 , n33683 , n33684 , n33685 , n33686 , n33687 , n33688 , n33689 , n33690 , n33691 , n33692 , n33693 , n33694 , n33695 , n33696 , n33697 , n33698 , n33699 , n33700 , n33701 , n33702 , n33703 , n33704 , n33705 , n33706 , n33707 , n33708 , n33709 , n33710 , n33711 , n33712 , n33713 , n33714 , n33715 , n33716 , n33717 , n33718 , n33719 , n33720 , n33721 , n33722 , n33723 , n33724 , n33725 , n33726 , n33727 , n33728 , n33729 , n33730 , n33731 , n33732 , n33733 , n33734 , n33735 , n33736 , n33737 , n33738 , n33739 , n33740 , n33741 , n33742 , n33743 , n33744 , n33745 , n33746 , n33747 , n33748 , n33749 , n33750 , n33751 , n33752 , n33753 , n33754 , n33755 , n33756 , n33757 , n33758 , n33759 , n33760 , n33761 , n33762 , n33763 , n33764 , n33765 , n33766 , n33767 , n33768 , n33769 , n33770 , n33771 , n33772 , n33773 , n33774 , n33775 , n33776 , n33777 , n33778 , n33779 , n33780 , n33781 , n33782 , n33783 , n33784 , n33785 , n33786 , n33787 , n33788 , n33789 , n33790 , n33791 , n33792 , n33793 , n33794 , n33795 , n33796 , n33797 , n33798 , n33799 , n33800 , n33801 , n33802 , n33803 , n33804 , n33805 , n33806 , n33807 , n33808 , n33809 , n33810 , n33811 , n33812 , n33813 , n33814 , n33815 , n33816 , n33817 , n33818 , n33819 , n33820 , n33821 , n33822 , n33823 , n33824 , n33825 , n33826 , n33827 , n33828 , n33829 , n33830 , n33831 , n33832 , n33833 , n33834 , n33835 , n33836 , n33837 , n33838 , n33839 , n33840 , n33841 , n33842 , n33843 , n33844 , n33845 , n33846 , n33847 , n33848 , n33849 , n33850 , n33851 , n33852 , n33853 , n33854 , n33855 , n33856 , n33857 , n33858 , n33859 , n33860 , n33861 , n33862 , n33863 , n33864 , n33865 , n33866 , n33867 , n33868 , n33869 , n33870 , n33871 , n33872 , n33873 , n33874 , n33875 , n33876 , n33877 , n33878 , n33879 , n33880 , n33881 , n33882 , n33883 , n33884 , n33885 , n33886 , n33887 , n33888 , n33889 , n33890 , n33891 , n33892 , n33893 , n33894 , n33895 , n33896 , n33897 , n33898 , n33899 , n33900 , n33901 , n33902 , n33903 , n33904 , n33905 , n33906 , n33907 , n33908 , n33909 , n33910 , n33911 , n33912 , n33913 , n33914 , n33915 , n33916 , n33917 , n33918 , n33919 , n33920 , n33921 , n33922 , n33923 , n33924 , n33925 , n33926 , n33927 , n33928 , n33929 , n33930 , n33931 , n33932 , n33933 , n33934 , n33935 , n33936 , n33937 , n33938 , n33939 , n33940 , n33941 , n33942 , n33943 , n33944 , n33945 , n33946 , n33947 , n33948 , n33949 , n33950 , n33951 , n33952 , n33953 , n33954 , n33955 , n33956 , n33957 , n33958 , n33959 , n33960 , n33961 , n33962 , n33963 , n33964 , n33965 , n33966 , n33967 , n33968 , n33969 , n33970 , n33971 , n33972 , n33973 , n33974 , n33975 , n33976 , n33977 , n33978 , n33979 , n33980 , n33981 , n33982 , n33983 , n33984 , n33985 , n33986 , n33987 , n33988 , n33989 , n33990 , n33991 , n33992 , n33993 , n33994 , n33995 , n33996 , n33997 , n33998 , n33999 , n34000 , n34001 , n34002 , n34003 , n34004 , n34005 , n34006 , n34007 , n34008 , n34009 , n34010 , n34011 , n34012 , n34013 , n34014 , n34015 , n34016 , n34017 , n34018 , n34019 , n34020 , n34021 , n34022 , n34023 , n34024 , n34025 , n34026 , n34027 , n34028 , n34029 , n34030 , n34031 , n34032 , n34033 , n34034 , n34035 , n34036 , n34037 , n34038 , n34039 , n34040 , n34041 , n34042 , n34043 , n34044 , n34045 , n34046 , n34047 , n34048 , n34049 , n34050 , n34051 , n34052 , n34053 , n34054 , n34055 , n34056 , n34057 , n34058 , n34059 , n34060 , n34061 , n34062 , n34063 , n34064 , n34065 , n34066 , n34067 , n34068 , n34069 , n34070 , n34071 , n34072 , n34073 , n34074 , n34075 , n34076 , n34077 , n34078 , n34079 , n34080 , n34081 , n34082 , n34083 , n34084 , n34085 , n34086 , n34087 , n34088 , n34089 , n34090 , n34091 , n34092 , n34093 , n34094 , n34095 , n34096 , n34097 , n34098 , n34099 , n34100 , n34101 , n34102 , n34103 , n34104 , n34105 , n34106 , n34107 , n34108 , n34109 , n34110 , n34111 , n34112 , n34113 , n34114 , n34115 , n34116 , n34117 , n34118 , n34119 , n34120 , n34121 , n34122 , n34123 , n34124 , n34125 , n34126 , n34127 , n34128 , n34129 , n34130 , n34131 , n34132 , n34133 , n34134 , n34135 , n34136 , n34137 , n34138 , n34139 , n34140 , n34141 , n34142 , n34143 , n34144 , n34145 , n34146 , n34147 , n34148 , n34149 , n34150 , n34151 , n34152 , n34153 , n34154 , n34155 , n34156 , n34157 , n34158 , n34159 , n34160 , n34161 , n34162 , n34163 , n34164 , n34165 , n34166 , n34167 , n34168 , n34169 , n34170 , n34171 , n34172 , n34173 , n34174 , n34175 , n34176 , n34177 , n34178 , n34179 , n34180 , n34181 , n34182 , n34183 , n34184 , n34185 , n34186 , n34187 , n34188 , n34189 , n34190 , n34191 , n34192 , n34193 , n34194 , n34195 , n34196 , n34197 , n34198 , n34199 , n34200 , n34201 , n34202 , n34203 , n34204 , n34205 , n34206 , n34207 , n34208 , n34209 , n34210 , n34211 , n34212 , n34213 , n34214 , n34215 , n34216 , n34217 , n34218 , n34219 , n34220 , n34221 , n34222 , n34223 , n34224 , n34225 , n34226 , n34227 , n34228 , n34229 , n34230 , n34231 , n34232 , n34233 , n34234 , n34235 , n34236 , n34237 , n34238 , n34239 , n34240 , n34241 , n34242 , n34243 , n34244 , n34245 , n34246 , n34247 , n34248 , n34249 , n34250 , n34251 , n34252 , n34253 , n34254 , n34255 , n34256 , n34257 , n34258 , n34259 , n34260 , n34261 , n34262 , n34263 , n34264 , n34265 , n34266 , n34267 , n34268 , n34269 , n34270 , n34271 , n34272 , n34273 , n34274 , n34275 , n34276 , n34277 , n34278 , n34279 , n34280 , n34281 , n34282 , n34283 , n34284 , n34285 , n34286 , n34287 , n34288 , n34289 , n34290 , n34291 , n34292 , n34293 , n34294 , n34295 , n34296 , n34297 , n34298 , n34299 , n34300 , n34301 , n34302 , n34303 , n34304 , n34305 , n34306 , n34307 , n34308 , n34309 , n34310 , n34311 , n34312 , n34313 , n34314 , n34315 , n34316 , n34317 , n34318 , n34319 , n34320 , n34321 , n34322 , n34323 , n34324 , n34325 , n34326 , n34327 , n34328 , n34329 , n34330 , n34331 , n34332 , n34333 , n34334 , n34335 , n34336 , n34337 , n34338 , n34339 , n34340 , n34341 , n34342 , n34343 , n34344 , n34345 , n34346 , n34347 , n34348 , n34349 , n34350 , n34351 , n34352 , n34353 , n34354 , n34355 , n34356 , n34357 , n34358 , n34359 , n34360 , n34361 , n34362 , n34363 , n34364 , n34365 , n34366 , n34367 , n34368 , n34369 , n34370 , n34371 , n34372 , n34373 , n34374 , n34375 , n34376 , n34377 , n34378 , n34379 , n34380 , n34381 , n34382 , n34383 , n34384 , n34385 , n34386 , n34387 , n34388 , n34389 , n34390 , n34391 , n34392 , n34393 , n34394 , n34395 , n34396 , n34397 , n34398 , n34399 , n34400 , n34401 , n34402 , n34403 , n34404 , n34405 , n34406 , n34407 , n34408 , n34409 , n34410 , n34411 , n34412 , n34413 , n34414 , n34415 , n34416 , n34417 , n34418 , n34419 , n34420 , n34421 , n34422 , n34423 , n34424 , n34425 , n34426 , n34427 , n34428 , n34429 , n34430 , n34431 , n34432 , n34433 , n34434 , n34435 , n34436 , n34437 , n34438 , n34439 , n34440 , n34441 , n34442 , n34443 , n34444 , n34445 , n34446 , n34447 , n34448 , n34449 , n34450 , n34451 , n34452 , n34453 , n34454 , n34455 , n34456 , n34457 , n34458 , n34459 , n34460 , n34461 , n34462 , n34463 , n34464 , n34465 , n34466 , n34467 , n34468 , n34469 , n34470 , n34471 , n34472 , n34473 , n34474 , n34475 , n34476 , n34477 , n34478 , n34479 , n34480 , n34481 , n34482 , n34483 , n34484 , n34485 , n34486 , n34487 , n34488 , n34489 , n34490 , n34491 , n34492 , n34493 , n34494 , n34495 , n34496 , n34497 , n34498 , n34499 , n34500 , n34501 , n34502 , n34503 , n34504 , n34505 , n34506 , n34507 , n34508 , n34509 , n34510 , n34511 , n34512 , n34513 , n34514 , n34515 , n34516 , n34517 , n34518 , n34519 , n34520 , n34521 , n34522 , n34523 , n34524 , n34525 , n34526 , n34527 , n34528 , n34529 , n34530 , n34531 , n34532 , n34533 , n34534 , n34535 , n34536 , n34537 , n34538 , n34539 , n34540 , n34541 , n34542 , n34543 , n34544 , n34545 , n34546 , n34547 , n34548 , n34549 , n34550 , n34551 , n34552 , n34553 , n34554 , n34555 , n34556 , n34557 , n34558 , n34559 , n34560 , n34561 , n34562 , n34563 , n34564 , n34565 , n34566 , n34567 , n34568 , n34569 , n34570 , n34571 , n34572 , n34573 , n34574 , n34575 , n34576 , n34577 , n34578 , n34579 , n34580 , n34581 , n34582 , n34583 , n34584 , n34585 , n34586 , n34587 , n34588 , n34589 , n34590 , n34591 , n34592 , n34593 , n34594 , n34595 , n34596 , n34597 , n34598 , n34599 , n34600 , n34601 , n34602 , n34603 , n34604 , n34605 , n34606 , n34607 , n34608 , n34609 , n34610 , n34611 , n34612 , n34613 , n34614 , n34615 , n34616 , n34617 , n34618 , n34619 , n34620 , n34621 , n34622 , n34623 , n34624 , n34625 , n34626 , n34627 , n34628 , n34629 , n34630 , n34631 , n34632 , n34633 , n34634 , n34635 , n34636 , n34637 , n34638 , n34639 , n34640 , n34641 , n34642 , n34643 , n34644 , n34645 , n34646 , n34647 , n34648 , n34649 , n34650 , n34651 , n34652 , n34653 , n34654 , n34655 , n34656 , n34657 , n34658 , n34659 , n34660 , n34661 , n34662 , n34663 , n34664 , n34665 , n34666 , n34667 , n34668 , n34669 , n34670 , n34671 , n34672 , n34673 , n34674 , n34675 , n34676 , n34677 , n34678 , n34679 , n34680 , n34681 , n34682 , n34683 , n34684 , n34685 , n34686 , n34687 , n34688 , n34689 , n34690 , n34691 , n34692 , n34693 , n34694 , n34695 , n34696 , n34697 , n34698 , n34699 , n34700 , n34701 , n34702 , n34703 , n34704 , n34705 , n34706 , n34707 , n34708 , n34709 , n34710 , n34711 , n34712 , n34713 , n34714 , n34715 , n34716 , n34717 , n34718 , n34719 , n34720 , n34721 , n34722 , n34723 , n34724 , n34725 , n34726 , n34727 , n34728 , n34729 , n34730 , n34731 , n34732 , n34733 , n34734 , n34735 , n34736 , n34737 , n34738 , n34739 , n34740 , n34741 , n34742 , n34743 , n34744 , n34745 , n34746 , n34747 , n34748 , n34749 , n34750 , n34751 , n34752 , n34753 , n34754 , n34755 , n34756 , n34757 , n34758 , n34759 , n34760 , n34761 , n34762 , n34763 , n34764 , n34765 , n34766 , n34767 , n34768 , n34769 , n34770 , n34771 , n34772 , n34773 , n34774 , n34775 , n34776 , n34777 , n34778 , n34779 , n34780 , n34781 , n34782 , n34783 , n34784 , n34785 , n34786 , n34787 , n34788 , n34789 , n34790 , n34791 , n34792 , n34793 , n34794 , n34795 , n34796 , n34797 , n34798 , n34799 , n34800 , n34801 , n34802 , n34803 , n34804 , n34805 , n34806 , n34807 , n34808 , n34809 , n34810 , n34811 , n34812 , n34813 , n34814 , n34815 , n34816 , n34817 , n34818 , n34819 , n34820 , n34821 , n34822 , n34823 , n34824 , n34825 , n34826 , n34827 , n34828 , n34829 , n34830 , n34831 , n34832 , n34833 , n34834 , n34835 , n34836 , n34837 , n34838 , n34839 , n34840 , n34841 , n34842 , n34843 , n34844 , n34845 , n34846 , n34847 , n34848 , n34849 , n34850 , n34851 , n34852 , n34853 , n34854 , n34855 , n34856 , n34857 , n34858 , n34859 , n34860 , n34861 , n34862 , n34863 , n34864 , n34865 , n34866 , n34867 , n34868 , n34869 , n34870 , n34871 , n34872 , n34873 , n34874 , n34875 , n34876 , n34877 , n34878 , n34879 , n34880 , n34881 , n34882 , n34883 , n34884 , n34885 , n34886 , n34887 , n34888 , n34889 , n34890 , n34891 , n34892 , n34893 , n34894 , n34895 , n34896 , n34897 , n34898 , n34899 , n34900 , n34901 , n34902 , n34903 , n34904 , n34905 , n34906 , n34907 , n34908 , n34909 , n34910 , n34911 , n34912 , n34913 , n34914 , n34915 , n34916 , n34917 , n34918 , n34919 , n34920 , n34921 , n34922 , n34923 , n34924 , n34925 , n34926 , n34927 , n34928 , n34929 , n34930 , n34931 , n34932 , n34933 , n34934 , n34935 , n34936 , n34937 , n34938 , n34939 , n34940 , n34941 , n34942 , n34943 , n34944 , n34945 , n34946 , n34947 , n34948 , n34949 , n34950 , n34951 , n34952 , n34953 , n34954 , n34955 , n34956 , n34957 , n34958 , n34959 , n34960 , n34961 , n34962 , n34963 , n34964 , n34965 , n34966 , n34967 , n34968 , n34969 , n34970 , n34971 , n34972 , n34973 , n34974 , n34975 , n34976 , n34977 , n34978 , n34979 , n34980 , n34981 , n34982 , n34983 , n34984 , n34985 , n34986 , n34987 , n34988 , n34989 , n34990 , n34991 , n34992 , n34993 , n34994 , n34995 , n34996 , n34997 , n34998 , n34999 , n35000 , n35001 , n35002 , n35003 , n35004 , n35005 , n35006 , n35007 , n35008 , n35009 , n35010 , n35011 , n35012 , n35013 , n35014 , n35015 , n35016 , n35017 , n35018 , n35019 , n35020 , n35021 , n35022 , n35023 , n35024 , n35025 , n35026 , n35027 , n35028 , n35029 , n35030 , n35031 , n35032 , n35033 , n35034 , n35035 , n35036 , n35037 , n35038 , n35039 , n35040 , n35041 , n35042 , n35043 , n35044 , n35045 , n35046 , n35047 , n35048 , n35049 , n35050 , n35051 , n35052 , n35053 , n35054 , n35055 , n35056 , n35057 , n35058 , n35059 , n35060 , n35061 , n35062 , n35063 , n35064 , n35065 , n35066 , n35067 , n35068 , n35069 , n35070 , n35071 , n35072 , n35073 , n35074 , n35075 , n35076 , n35077 , n35078 , n35079 , n35080 , n35081 , n35082 , n35083 , n35084 , n35085 , n35086 , n35087 , n35088 , n35089 , n35090 , n35091 , n35092 , n35093 , n35094 , n35095 , n35096 , n35097 , n35098 , n35099 , n35100 , n35101 , n35102 , n35103 , n35104 , n35105 , n35106 , n35107 , n35108 , n35109 , n35110 , n35111 , n35112 , n35113 , n35114 , n35115 , n35116 , n35117 , n35118 , n35119 , n35120 , n35121 , n35122 , n35123 , n35124 , n35125 , n35126 , n35127 , n35128 , n35129 , n35130 , n35131 , n35132 , n35133 , n35134 , n35135 , n35136 , n35137 , n35138 , n35139 , n35140 , n35141 , n35142 , n35143 , n35144 , n35145 , n35146 , n35147 , n35148 , n35149 , n35150 , n35151 , n35152 , n35153 , n35154 , n35155 , n35156 , n35157 , n35158 , n35159 , n35160 , n35161 , n35162 , n35163 , n35164 , n35165 , n35166 , n35167 , n35168 , n35169 , n35170 , n35171 , n35172 , n35173 , n35174 , n35175 , n35176 , n35177 , n35178 , n35179 , n35180 , n35181 , n35182 , n35183 , n35184 , n35185 , n35186 , n35187 , n35188 , n35189 , n35190 , n35191 , n35192 , n35193 , n35194 , n35195 , n35196 , n35197 , n35198 , n35199 , n35200 , n35201 , n35202 , n35203 , n35204 , n35205 , n35206 , n35207 , n35208 , n35209 , n35210 , n35211 , n35212 , n35213 , n35214 , n35215 , n35216 , n35217 , n35218 , n35219 , n35220 , n35221 , n35222 , n35223 , n35224 , n35225 , n35226 , n35227 , n35228 , n35229 , n35230 , n35231 , n35232 , n35233 , n35234 , n35235 , n35236 , n35237 , n35238 , n35239 , n35240 , n35241 , n35242 , n35243 , n35244 , n35245 , n35246 , n35247 , n35248 , n35249 , n35250 , n35251 , n35252 , n35253 , n35254 , n35255 , n35256 , n35257 , n35258 , n35259 , n35260 , n35261 , n35262 , n35263 , n35264 , n35265 , n35266 , n35267 , n35268 , n35269 , n35270 , n35271 , n35272 , n35273 , n35274 , n35275 , n35276 , n35277 , n35278 , n35279 , n35280 , n35281 , n35282 , n35283 , n35284 , n35285 , n35286 , n35287 , n35288 , n35289 , n35290 , n35291 , n35292 , n35293 , n35294 , n35295 , n35296 , n35297 , n35298 , n35299 , n35300 , n35301 , n35302 , n35303 , n35304 , n35305 , n35306 , n35307 , n35308 , n35309 , n35310 , n35311 , n35312 , n35313 , n35314 , n35315 , n35316 , n35317 , n35318 , n35319 , n35320 , n35321 , n35322 , n35323 , n35324 , n35325 , n35326 , n35327 , n35328 , n35329 , n35330 , n35331 , n35332 , n35333 , n35334 , n35335 , n35336 , n35337 , n35338 , n35339 , n35340 , n35341 , n35342 , n35343 , n35344 , n35345 , n35346 , n35347 , n35348 , n35349 , n35350 , n35351 , n35352 , n35353 , n35354 , n35355 , n35356 , n35357 , n35358 , n35359 , n35360 , n35361 , n35362 , n35363 , n35364 , n35365 , n35366 , n35367 , n35368 , n35369 , n35370 , n35371 , n35372 , n35373 , n35374 , n35375 , n35376 , n35377 , n35378 , n35379 , n35380 , n35381 , n35382 , n35383 , n35384 , n35385 , n35386 , n35387 , n35388 , n35389 , n35390 , n35391 , n35392 , n35393 , n35394 , n35395 , n35396 , n35397 , n35398 , n35399 , n35400 , n35401 , n35402 , n35403 , n35404 , n35405 , n35406 , n35407 , n35408 , n35409 , n35410 , n35411 , n35412 , n35413 , n35414 , n35415 , n35416 , n35417 , n35418 , n35419 , n35420 , n35421 , n35422 , n35423 , n35424 , n35425 , n35426 , n35427 , n35428 , n35429 , n35430 , n35431 , n35432 , n35433 , n35434 , n35435 , n35436 , n35437 , n35438 , n35439 , n35440 , n35441 , n35442 , n35443 , n35444 , n35445 , n35446 , n35447 , n35448 , n35449 , n35450 , n35451 , n35452 , n35453 , n35454 , n35455 , n35456 , n35457 , n35458 , n35459 , n35460 , n35461 , n35462 , n35463 , n35464 , n35465 , n35466 , n35467 , n35468 , n35469 , n35470 , n35471 , n35472 , n35473 , n35474 , n35475 , n35476 , n35477 , n35478 , n35479 , n35480 , n35481 , n35482 , n35483 , n35484 , n35485 , n35486 , n35487 , n35488 , n35489 , n35490 , n35491 , n35492 , n35493 , n35494 , n35495 , n35496 , n35497 , n35498 , n35499 , n35500 , n35501 , n35502 , n35503 , n35504 , n35505 , n35506 , n35507 , n35508 , n35509 , n35510 , n35511 , n35512 , n35513 , n35514 , n35515 , n35516 , n35517 , n35518 , n35519 , n35520 , n35521 , n35522 , n35523 , n35524 , n35525 , n35526 , n35527 , n35528 , n35529 , n35530 , n35531 , n35532 , n35533 , n35534 , n35535 , n35536 , n35537 , n35538 , n35539 , n35540 , n35541 , n35542 , n35543 , n35544 , n35545 , n35546 , n35547 , n35548 , n35549 , n35550 , n35551 , n35552 , n35553 , n35554 , n35555 , n35556 , n35557 , n35558 , n35559 , n35560 , n35561 , n35562 , n35563 , n35564 , n35565 , n35566 , n35567 , n35568 , n35569 , n35570 , n35571 , n35572 , n35573 , n35574 , n35575 , n35576 , n35577 , n35578 , n35579 , n35580 , n35581 , n35582 , n35583 , n35584 , n35585 , n35586 , n35587 , n35588 , n35589 , n35590 , n35591 , n35592 , n35593 , n35594 , n35595 , n35596 , n35597 , n35598 , n35599 , n35600 , n35601 , n35602 , n35603 , n35604 , n35605 , n35606 , n35607 , n35608 , n35609 , n35610 , n35611 , n35612 , n35613 , n35614 , n35615 , n35616 , n35617 , n35618 , n35619 , n35620 , n35621 , n35622 , n35623 , n35624 , n35625 , n35626 , n35627 , n35628 , n35629 , n35630 , n35631 , n35632 , n35633 , n35634 , n35635 , n35636 , n35637 , n35638 , n35639 , n35640 , n35641 , n35642 , n35643 , n35644 , n35645 , n35646 , n35647 , n35648 , n35649 , n35650 , n35651 , n35652 , n35653 , n35654 , n35655 , n35656 , n35657 , n35658 , n35659 , n35660 , n35661 , n35662 , n35663 , n35664 , n35665 , n35666 , n35667 , n35668 , n35669 , n35670 , n35671 , n35672 , n35673 , n35674 , n35675 , n35676 , n35677 , n35678 , n35679 , n35680 , n35681 , n35682 , n35683 , n35684 , n35685 , n35686 , n35687 , n35688 , n35689 , n35690 , n35691 , n35692 , n35693 , n35694 , n35695 , n35696 , n35697 , n35698 , n35699 , n35700 , n35701 , n35702 , n35703 , n35704 , n35705 , n35706 , n35707 , n35708 , n35709 , n35710 , n35711 , n35712 , n35713 , n35714 , n35715 , n35716 , n35717 , n35718 , n35719 , n35720 , n35721 , n35722 , n35723 , n35724 , n35725 , n35726 , n35727 , n35728 , n35729 , n35730 , n35731 , n35732 , n35733 , n35734 , n35735 , n35736 , n35737 , n35738 , n35739 , n35740 , n35741 , n35742 , n35743 , n35744 , n35745 , n35746 , n35747 , n35748 , n35749 , n35750 , n35751 , n35752 , n35753 , n35754 , n35755 , n35756 , n35757 , n35758 , n35759 , n35760 , n35761 , n35762 , n35763 , n35764 , n35765 , n35766 , n35767 , n35768 , n35769 , n35770 , n35771 , n35772 , n35773 , n35774 , n35775 , n35776 , n35777 , n35778 , n35779 , n35780 , n35781 , n35782 , n35783 , n35784 , n35785 , n35786 , n35787 , n35788 , n35789 , n35790 , n35791 , n35792 , n35793 , n35794 , n35795 , n35796 , n35797 , n35798 , n35799 , n35800 , n35801 , n35802 , n35803 , n35804 , n35805 , n35806 , n35807 , n35808 , n35809 , n35810 , n35811 , n35812 , n35813 , n35814 , n35815 , n35816 , n35817 , n35818 , n35819 , n35820 , n35821 , n35822 , n35823 , n35824 , n35825 , n35826 , n35827 , n35828 , n35829 , n35830 , n35831 , n35832 , n35833 , n35834 , n35835 , n35836 , n35837 , n35838 , n35839 , n35840 , n35841 , n35842 , n35843 , n35844 , n35845 , n35846 , n35847 , n35848 , n35849 , n35850 , n35851 , n35852 , n35853 , n35854 , n35855 , n35856 , n35857 , n35858 , n35859 , n35860 , n35861 , n35862 , n35863 , n35864 , n35865 , n35866 , n35867 , n35868 , n35869 , n35870 , n35871 , n35872 , n35873 , n35874 , n35875 , n35876 , n35877 , n35878 , n35879 , n35880 , n35881 , n35882 , n35883 , n35884 , n35885 , n35886 , n35887 , n35888 , n35889 , n35890 , n35891 , n35892 , n35893 , n35894 , n35895 , n35896 , n35897 , n35898 , n35899 , n35900 , n35901 , n35902 , n35903 , n35904 , n35905 , n35906 , n35907 , n35908 , n35909 , n35910 , n35911 , n35912 , n35913 , n35914 , n35915 , n35916 , n35917 , n35918 , n35919 , n35920 , n35921 , n35922 , n35923 , n35924 , n35925 , n35926 , n35927 , n35928 , n35929 , n35930 , n35931 , n35932 , n35933 , n35934 , n35935 , n35936 , n35937 , n35938 , n35939 , n35940 , n35941 , n35942 , n35943 , n35944 , n35945 , n35946 , n35947 , n35948 , n35949 , n35950 , n35951 , n35952 , n35953 , n35954 , n35955 , n35956 , n35957 , n35958 , n35959 , n35960 , n35961 , n35962 , n35963 , n35964 , n35965 , n35966 , n35967 , n35968 , n35969 , n35970 , n35971 , n35972 , n35973 , n35974 , n35975 , n35976 , n35977 , n35978 , n35979 , n35980 , n35981 , n35982 , n35983 , n35984 , n35985 , n35986 , n35987 , n35988 , n35989 , n35990 , n35991 , n35992 , n35993 , n35994 , n35995 , n35996 , n35997 , n35998 , n35999 , n36000 , n36001 , n36002 , n36003 , n36004 , n36005 , n36006 , n36007 , n36008 , n36009 , n36010 , n36011 , n36012 , n36013 , n36014 , n36015 , n36016 , n36017 , n36018 , n36019 , n36020 , n36021 , n36022 , n36023 , n36024 , n36025 , n36026 , n36027 , n36028 , n36029 , n36030 , n36031 , n36032 , n36033 , n36034 , n36035 , n36036 , n36037 , n36038 , n36039 , n36040 , n36041 , n36042 , n36043 , n36044 , n36045 , n36046 , n36047 , n36048 , n36049 , n36050 , n36051 , n36052 , n36053 , n36054 , n36055 , n36056 , n36057 , n36058 , n36059 , n36060 , n36061 , n36062 , n36063 , n36064 , n36065 , n36066 , n36067 , n36068 , n36069 , n36070 , n36071 , n36072 , n36073 , n36074 , n36075 , n36076 , n36077 , n36078 , n36079 , n36080 , n36081 , n36082 , n36083 , n36084 , n36085 , n36086 , n36087 , n36088 , n36089 , n36090 , n36091 , n36092 , n36093 , n36094 , n36095 , n36096 , n36097 , n36098 , n36099 , n36100 , n36101 , n36102 , n36103 , n36104 , n36105 , n36106 , n36107 , n36108 , n36109 , n36110 , n36111 , n36112 , n36113 , n36114 , n36115 , n36116 , n36117 , n36118 , n36119 , n36120 , n36121 , n36122 , n36123 , n36124 , n36125 , n36126 , n36127 , n36128 , n36129 , n36130 , n36131 , n36132 , n36133 , n36134 , n36135 , n36136 , n36137 , n36138 , n36139 , n36140 , n36141 , n36142 , n36143 , n36144 , n36145 , n36146 , n36147 , n36148 , n36149 , n36150 , n36151 , n36152 , n36153 , n36154 , n36155 , n36156 , n36157 , n36158 , n36159 , n36160 , n36161 , n36162 , n36163 , n36164 , n36165 , n36166 , n36167 , n36168 , n36169 , n36170 , n36171 , n36172 , n36173 , n36174 , n36175 , n36176 , n36177 , n36178 , n36179 , n36180 , n36181 , n36182 , n36183 , n36184 , n36185 , n36186 , n36187 , n36188 , n36189 , n36190 , n36191 , n36192 , n36193 , n36194 , n36195 , n36196 , n36197 , n36198 , n36199 , n36200 , n36201 , n36202 , n36203 , n36204 , n36205 , n36206 , n36207 , n36208 , n36209 , n36210 , n36211 , n36212 , n36213 , n36214 , n36215 , n36216 , n36217 , n36218 , n36219 , n36220 , n36221 , n36222 , n36223 , n36224 , n36225 , n36226 , n36227 , n36228 , n36229 , n36230 , n36231 , n36232 , n36233 , n36234 , n36235 , n36236 , n36237 , n36238 , n36239 , n36240 , n36241 , n36242 , n36243 , n36244 , n36245 , n36246 , n36247 , n36248 , n36249 , n36250 , n36251 , n36252 , n36253 , n36254 , n36255 , n36256 , n36257 , n36258 , n36259 , n36260 , n36261 , n36262 , n36263 , n36264 , n36265 , n36266 , n36267 , n36268 , n36269 , n36270 , n36271 , n36272 , n36273 , n36274 , n36275 , n36276 , n36277 , n36278 , n36279 , n36280 , n36281 , n36282 , n36283 , n36284 , n36285 , n36286 , n36287 , n36288 , n36289 , n36290 , n36291 , n36292 , n36293 , n36294 , n36295 , n36296 , n36297 , n36298 , n36299 , n36300 , n36301 , n36302 , n36303 , n36304 , n36305 , n36306 , n36307 , n36308 , n36309 , n36310 , n36311 , n36312 , n36313 , n36314 , n36315 , n36316 , n36317 , n36318 , n36319 , n36320 , n36321 , n36322 , n36323 , n36324 , n36325 , n36326 , n36327 , n36328 , n36329 , n36330 , n36331 , n36332 , n36333 , n36334 , n36335 , n36336 , n36337 , n36338 , n36339 , n36340 , n36341 , n36342 , n36343 , n36344 , n36345 , n36346 , n36347 , n36348 , n36349 , n36350 , n36351 , n36352 , n36353 , n36354 , n36355 , n36356 , n36357 , n36358 , n36359 , n36360 , n36361 , n36362 , n36363 , n36364 , n36365 , n36366 , n36367 , n36368 , n36369 , n36370 , n36371 , n36372 , n36373 , n36374 , n36375 , n36376 , n36377 , n36378 , n36379 , n36380 , n36381 , n36382 , n36383 , n36384 , n36385 , n36386 , n36387 , n36388 , n36389 , n36390 , n36391 , n36392 , n36393 , n36394 , n36395 , n36396 , n36397 , n36398 , n36399 , n36400 , n36401 , n36402 , n36403 , n36404 , n36405 , n36406 , n36407 , n36408 , n36409 , n36410 , n36411 , n36412 , n36413 , n36414 , n36415 , n36416 , n36417 , n36418 , n36419 , n36420 , n36421 , n36422 , n36423 , n36424 , n36425 , n36426 , n36427 , n36428 , n36429 , n36430 , n36431 , n36432 , n36433 , n36434 , n36435 , n36436 , n36437 , n36438 , n36439 , n36440 , n36441 , n36442 , n36443 , n36444 , n36445 , n36446 , n36447 , n36448 , n36449 , n36450 , n36451 , n36452 , n36453 , n36454 , n36455 , n36456 , n36457 , n36458 , n36459 , n36460 , n36461 , n36462 , n36463 , n36464 , n36465 , n36466 , n36467 , n36468 , n36469 , n36470 , n36471 , n36472 , n36473 , n36474 , n36475 , n36476 , n36477 , n36478 , n36479 , n36480 , n36481 , n36482 , n36483 , n36484 , n36485 , n36486 , n36487 , n36488 , n36489 , n36490 , n36491 , n36492 , n36493 , n36494 , n36495 , n36496 , n36497 , n36498 , n36499 , n36500 , n36501 , n36502 , n36503 , n36504 , n36505 , n36506 , n36507 , n36508 , n36509 , n36510 , n36511 , n36512 , n36513 , n36514 , n36515 , n36516 , n36517 , n36518 , n36519 , n36520 , n36521 , n36522 , n36523 , n36524 , n36525 , n36526 , n36527 , n36528 , n36529 , n36530 , n36531 , n36532 , n36533 , n36534 , n36535 , n36536 , n36537 , n36538 , n36539 , n36540 , n36541 , n36542 , n36543 , n36544 , n36545 , n36546 , n36547 , n36548 , n36549 , n36550 , n36551 , n36552 , n36553 , n36554 , n36555 , n36556 , n36557 , n36558 , n36559 , n36560 , n36561 , n36562 , n36563 , n36564 , n36565 , n36566 , n36567 , n36568 , n36569 , n36570 , n36571 , n36572 , n36573 , n36574 , n36575 , n36576 , n36577 , n36578 , n36579 , n36580 , n36581 , n36582 , n36583 , n36584 , n36585 , n36586 , n36587 , n36588 , n36589 , n36590 , n36591 , n36592 , n36593 , n36594 , n36595 , n36596 , n36597 , n36598 , n36599 , n36600 , n36601 , n36602 , n36603 , n36604 , n36605 , n36606 , n36607 , n36608 , n36609 , n36610 , n36611 , n36612 , n36613 , n36614 , n36615 , n36616 , n36617 , n36618 , n36619 , n36620 , n36621 , n36622 , n36623 , n36624 , n36625 , n36626 , n36627 , n36628 , n36629 , n36630 , n36631 , n36632 , n36633 , n36634 , n36635 , n36636 , n36637 , n36638 , n36639 , n36640 , n36641 , n36642 , n36643 , n36644 , n36645 , n36646 , n36647 , n36648 , n36649 , n36650 , n36651 , n36652 , n36653 , n36654 , n36655 , n36656 , n36657 , n36658 , n36659 , n36660 , n36661 , n36662 , n36663 , n36664 , n36665 , n36666 , n36667 , n36668 , n36669 , n36670 , n36671 , n36672 , n36673 , n36674 , n36675 , n36676 , n36677 , n36678 , n36679 , n36680 , n36681 , n36682 , n36683 , n36684 , n36685 , n36686 , n36687 , n36688 , n36689 , n36690 , n36691 , n36692 , n36693 , n36694 , n36695 , n36696 , n36697 , n36698 , n36699 , n36700 , n36701 , n36702 , n36703 , n36704 , n36705 , n36706 , n36707 , n36708 , n36709 , n36710 , n36711 , n36712 , n36713 , n36714 , n36715 , n36716 , n36717 , n36718 , n36719 , n36720 , n36721 , n36722 , n36723 , n36724 , n36725 , n36726 , n36727 , n36728 , n36729 , n36730 , n36731 , n36732 , n36733 , n36734 , n36735 , n36736 , n36737 , n36738 , n36739 , n36740 , n36741 , n36742 , n36743 , n36744 , n36745 , n36746 , n36747 , n36748 , n36749 , n36750 , n36751 , n36752 , n36753 , n36754 , n36755 , n36756 , n36757 , n36758 , n36759 , n36760 , n36761 , n36762 , n36763 , n36764 , n36765 , n36766 , n36767 , n36768 , n36769 , n36770 , n36771 , n36772 , n36773 , n36774 , n36775 , n36776 , n36777 , n36778 , n36779 , n36780 , n36781 , n36782 , n36783 , n36784 , n36785 , n36786 , n36787 , n36788 , n36789 , n36790 , n36791 , n36792 , n36793 , n36794 , n36795 , n36796 , n36797 , n36798 , n36799 , n36800 , n36801 , n36802 , n36803 , n36804 , n36805 , n36806 , n36807 , n36808 , n36809 , n36810 , n36811 , n36812 , n36813 , n36814 , n36815 , n36816 , n36817 , n36818 , n36819 , n36820 , n36821 , n36822 , n36823 , n36824 , n36825 , n36826 , n36827 , n36828 , n36829 , n36830 , n36831 , n36832 , n36833 , n36834 , n36835 , n36836 , n36837 , n36838 , n36839 , n36840 , n36841 , n36842 , n36843 , n36844 , n36845 , n36846 , n36847 , n36848 , n36849 , n36850 , n36851 , n36852 , n36853 , n36854 , n36855 , n36856 , n36857 , n36858 , n36859 , n36860 , n36861 , n36862 , n36863 , n36864 , n36865 , n36866 , n36867 , n36868 , n36869 , n36870 , n36871 , n36872 , n36873 , n36874 , n36875 , n36876 , n36877 , n36878 , n36879 , n36880 , n36881 , n36882 , n36883 , n36884 , n36885 , n36886 , n36887 , n36888 , n36889 , n36890 , n36891 , n36892 , n36893 , n36894 , n36895 , n36896 , n36897 , n36898 , n36899 , n36900 , n36901 , n36902 , n36903 , n36904 , n36905 , n36906 , n36907 , n36908 , n36909 , n36910 , n36911 , n36912 , n36913 , n36914 , n36915 , n36916 , n36917 , n36918 , n36919 , n36920 , n36921 , n36922 , n36923 , n36924 , n36925 , n36926 , n36927 , n36928 , n36929 , n36930 , n36931 , n36932 , n36933 , n36934 , n36935 , n36936 , n36937 , n36938 , n36939 , n36940 , n36941 , n36942 , n36943 , n36944 , n36945 , n36946 , n36947 , n36948 , n36949 , n36950 , n36951 , n36952 , n36953 , n36954 , n36955 , n36956 , n36957 , n36958 , n36959 , n36960 , n36961 , n36962 , n36963 , n36964 , n36965 , n36966 , n36967 , n36968 , n36969 , n36970 , n36971 , n36972 , n36973 , n36974 , n36975 , n36976 , n36977 , n36978 , n36979 , n36980 , n36981 , n36982 , n36983 , n36984 , n36985 , n36986 , n36987 , n36988 , n36989 , n36990 , n36991 , n36992 , n36993 , n36994 , n36995 , n36996 , n36997 , n36998 , n36999 , n37000 , n37001 , n37002 , n37003 , n37004 , n37005 , n37006 , n37007 , n37008 , n37009 , n37010 , n37011 , n37012 , n37013 , n37014 , n37015 , n37016 , n37017 , n37018 , n37019 , n37020 , n37021 , n37022 , n37023 , n37024 , n37025 , n37026 , n37027 , n37028 , n37029 , n37030 , n37031 , n37032 , n37033 , n37034 , n37035 , n37036 , n37037 , n37038 , n37039 , n37040 , n37041 , n37042 , n37043 , n37044 , n37045 , n37046 , n37047 , n37048 , n37049 , n37050 , n37051 , n37052 , n37053 , n37054 , n37055 , n37056 , n37057 , n37058 , n37059 , n37060 , n37061 , n37062 , n37063 , n37064 , n37065 , n37066 , n37067 , n37068 , n37069 , n37070 , n37071 , n37072 , n37073 , n37074 , n37075 , n37076 , n37077 , n37078 , n37079 , n37080 , n37081 , n37082 , n37083 , n37084 , n37085 , n37086 , n37087 , n37088 , n37089 , n37090 , n37091 , n37092 , n37093 , n37094 , n37095 , n37096 , n37097 , n37098 , n37099 , n37100 , n37101 , n37102 , n37103 , n37104 , n37105 , n37106 , n37107 , n37108 , n37109 , n37110 , n37111 , n37112 , n37113 , n37114 , n37115 , n37116 , n37117 , n37118 , n37119 , n37120 , n37121 , n37122 , n37123 , n37124 , n37125 , n37126 , n37127 , n37128 , n37129 , n37130 , n37131 , n37132 , n37133 , n37134 , n37135 , n37136 , n37137 , n37138 , n37139 , n37140 , n37141 , n37142 , n37143 , n37144 , n37145 , n37146 , n37147 , n37148 , n37149 , n37150 , n37151 , n37152 , n37153 , n37154 , n37155 , n37156 , n37157 , n37158 , n37159 , n37160 , n37161 , n37162 , n37163 , n37164 , n37165 , n37166 , n37167 , n37168 , n37169 , n37170 , n37171 , n37172 , n37173 , n37174 , n37175 , n37176 , n37177 , n37178 , n37179 , n37180 , n37181 , n37182 , n37183 , n37184 , n37185 , n37186 , n37187 , n37188 , n37189 , n37190 , n37191 , n37192 , n37193 , n37194 , n37195 , n37196 , n37197 , n37198 , n37199 , n37200 , n37201 , n37202 , n37203 , n37204 , n37205 , n37206 , n37207 , n37208 , n37209 , n37210 , n37211 , n37212 , n37213 , n37214 , n37215 , n37216 , n37217 , n37218 , n37219 , n37220 , n37221 , n37222 , n37223 , n37224 , n37225 , n37226 , n37227 , n37228 , n37229 , n37230 , n37231 , n37232 , n37233 , n37234 , n37235 , n37236 , n37237 , n37238 , n37239 , n37240 , n37241 , n37242 , n37243 , n37244 , n37245 , n37246 , n37247 , n37248 , n37249 , n37250 , n37251 , n37252 , n37253 , n37254 , n37255 , n37256 , n37257 , n37258 , n37259 , n37260 , n37261 , n37262 , n37263 , n37264 , n37265 , n37266 , n37267 , n37268 , n37269 , n37270 , n37271 , n37272 , n37273 , n37274 , n37275 , n37276 , n37277 , n37278 , n37279 , n37280 , n37281 , n37282 , n37283 , n37284 , n37285 , n37286 , n37287 , n37288 , n37289 , n37290 , n37291 , n37292 , n37293 , n37294 , n37295 , n37296 , n37297 , n37298 , n37299 , n37300 , n37301 , n37302 , n37303 , n37304 , n37305 , n37306 , n37307 , n37308 , n37309 , n37310 , n37311 , n37312 , n37313 , n37314 , n37315 , n37316 , n37317 , n37318 , n37319 , n37320 , n37321 , n37322 , n37323 , n37324 , n37325 , n37326 , n37327 , n37328 , n37329 , n37330 , n37331 , n37332 , n37333 , n37334 , n37335 , n37336 , n37337 , n37338 , n37339 , n37340 , n37341 , n37342 , n37343 , n37344 , n37345 , n37346 , n37347 , n37348 , n37349 , n37350 , n37351 , n37352 , n37353 , n37354 , n37355 , n37356 , n37357 , n37358 , n37359 , n37360 , n37361 , n37362 , n37363 , n37364 , n37365 , n37366 , n37367 , n37368 , n37369 , n37370 , n37371 , n37372 , n37373 , n37374 , n37375 , n37376 , n37377 , n37378 , n37379 , n37380 , n37381 , n37382 , n37383 , n37384 , n37385 , n37386 , n37387 , n37388 , n37389 , n37390 , n37391 , n37392 , n37393 , n37394 , n37395 , n37396 , n37397 , n37398 , n37399 , n37400 , n37401 , n37402 , n37403 , n37404 , n37405 , n37406 , n37407 , n37408 , n37409 , n37410 , n37411 , n37412 , n37413 , n37414 , n37415 , n37416 , n37417 , n37418 , n37419 , n37420 , n37421 , n37422 , n37423 , n37424 , n37425 , n37426 , n37427 , n37428 , n37429 , n37430 , n37431 , n37432 , n37433 , n37434 , n37435 , n37436 , n37437 , n37438 , n37439 , n37440 , n37441 , n37442 , n37443 , n37444 , n37445 , n37446 , n37447 , n37448 , n37449 , n37450 , n37451 , n37452 , n37453 , n37454 , n37455 , n37456 , n37457 , n37458 , n37459 , n37460 , n37461 , n37462 , n37463 , n37464 , n37465 , n37466 , n37467 , n37468 , n37469 , n37470 , n37471 , n37472 , n37473 , n37474 , n37475 , n37476 , n37477 , n37478 , n37479 , n37480 , n37481 , n37482 , n37483 , n37484 , n37485 , n37486 , n37487 , n37488 , n37489 , n37490 , n37491 , n37492 , n37493 , n37494 , n37495 , n37496 , n37497 , n37498 , n37499 , n37500 , n37501 , n37502 , n37503 , n37504 , n37505 , n37506 , n37507 , n37508 , n37509 , n37510 , n37511 , n37512 , n37513 , n37514 , n37515 , n37516 , n37517 , n37518 , n37519 , n37520 , n37521 , n37522 , n37523 , n37524 , n37525 , n37526 , n37527 , n37528 , n37529 , n37530 , n37531 , n37532 , n37533 , n37534 , n37535 , n37536 , n37537 , n37538 , n37539 , n37540 , n37541 , n37542 , n37543 , n37544 , n37545 , n37546 , n37547 , n37548 , n37549 , n37550 , n37551 , n37552 , n37553 , n37554 , n37555 , n37556 , n37557 , n37558 , n37559 , n37560 , n37561 , n37562 , n37563 , n37564 , n37565 , n37566 , n37567 , n37568 , n37569 , n37570 , n37571 , n37572 , n37573 , n37574 , n37575 , n37576 , n37577 , n37578 , n37579 , n37580 , n37581 , n37582 , n37583 , n37584 , n37585 , n37586 , n37587 , n37588 , n37589 , n37590 , n37591 , n37592 , n37593 , n37594 , n37595 , n37596 , n37597 , n37598 , n37599 , n37600 , n37601 , n37602 , n37603 , n37604 , n37605 , n37606 , n37607 , n37608 , n37609 , n37610 , n37611 , n37612 , n37613 , n37614 , n37615 , n37616 , n37617 , n37618 , n37619 , n37620 , n37621 , n37622 , n37623 , n37624 , n37625 , n37626 , n37627 , n37628 , n37629 , n37630 , n37631 , n37632 , n37633 , n37634 , n37635 , n37636 , n37637 , n37638 , n37639 , n37640 , n37641 , n37642 , n37643 , n37644 , n37645 , n37646 , n37647 , n37648 , n37649 , n37650 , n37651 , n37652 , n37653 , n37654 , n37655 , n37656 , n37657 , n37658 , n37659 , n37660 , n37661 , n37662 , n37663 , n37664 , n37665 , n37666 , n37667 , n37668 , n37669 , n37670 , n37671 , n37672 , n37673 , n37674 , n37675 , n37676 , n37677 , n37678 , n37679 , n37680 , n37681 , n37682 , n37683 , n37684 , n37685 , n37686 , n37687 , n37688 , n37689 , n37690 , n37691 , n37692 , n37693 , n37694 , n37695 , n37696 , n37697 , n37698 , n37699 , n37700 , n37701 , n37702 , n37703 , n37704 , n37705 , n37706 , n37707 , n37708 , n37709 , n37710 , n37711 , n37712 , n37713 , n37714 , n37715 , n37716 , n37717 , n37718 , n37719 , n37720 , n37721 , n37722 , n37723 , n37724 , n37725 , n37726 , n37727 , n37728 , n37729 , n37730 , n37731 , n37732 , n37733 , n37734 , n37735 , n37736 , n37737 , n37738 , n37739 , n37740 , n37741 , n37742 , n37743 , n37744 , n37745 , n37746 , n37747 , n37748 , n37749 , n37750 , n37751 , n37752 , n37753 , n37754 , n37755 , n37756 , n37757 , n37758 , n37759 , n37760 , n37761 , n37762 , n37763 , n37764 , n37765 , n37766 , n37767 , n37768 , n37769 , n37770 , n37771 , n37772 , n37773 , n37774 , n37775 , n37776 , n37777 , n37778 , n37779 , n37780 , n37781 , n37782 , n37783 , n37784 , n37785 , n37786 , n37787 , n37788 , n37789 , n37790 , n37791 , n37792 , n37793 , n37794 , n37795 , n37796 , n37797 , n37798 , n37799 , n37800 , n37801 , n37802 , n37803 , n37804 , n37805 , n37806 , n37807 , n37808 , n37809 , n37810 , n37811 , n37812 , n37813 , n37814 , n37815 , n37816 , n37817 , n37818 , n37819 , n37820 , n37821 , n37822 , n37823 , n37824 , n37825 , n37826 , n37827 , n37828 , n37829 , n37830 , n37831 , n37832 , n37833 , n37834 , n37835 , n37836 , n37837 , n37838 , n37839 , n37840 , n37841 , n37842 , n37843 , n37844 , n37845 , n37846 , n37847 , n37848 , n37849 , n37850 , n37851 , n37852 , n37853 , n37854 , n37855 , n37856 , n37857 , n37858 , n37859 , n37860 , n37861 , n37862 , n37863 , n37864 , n37865 , n37866 , n37867 , n37868 , n37869 , n37870 , n37871 , n37872 , n37873 , n37874 , n37875 , n37876 , n37877 , n37878 , n37879 , n37880 , n37881 , n37882 , n37883 , n37884 , n37885 , n37886 , n37887 , n37888 , n37889 , n37890 , n37891 , n37892 , n37893 , n37894 , n37895 , n37896 , n37897 , n37898 , n37899 , n37900 , n37901 , n37902 , n37903 , n37904 , n37905 , n37906 , n37907 , n37908 , n37909 , n37910 , n37911 , n37912 , n37913 , n37914 , n37915 , n37916 , n37917 , n37918 , n37919 , n37920 , n37921 , n37922 , n37923 , n37924 , n37925 , n37926 , n37927 , n37928 , n37929 , n37930 , n37931 , n37932 , n37933 , n37934 , n37935 , n37936 , n37937 , n37938 , n37939 , n37940 , n37941 , n37942 , n37943 , n37944 , n37945 , n37946 , n37947 , n37948 , n37949 , n37950 , n37951 , n37952 , n37953 , n37954 , n37955 , n37956 , n37957 , n37958 , n37959 , n37960 , n37961 , n37962 , n37963 , n37964 , n37965 , n37966 , n37967 , n37968 , n37969 , n37970 , n37971 , n37972 , n37973 , n37974 , n37975 , n37976 , n37977 , n37978 , n37979 , n37980 , n37981 , n37982 , n37983 , n37984 , n37985 , n37986 , n37987 , n37988 , n37989 , n37990 , n37991 , n37992 , n37993 , n37994 , n37995 , n37996 , n37997 , n37998 , n37999 , n38000 , n38001 , n38002 , n38003 , n38004 , n38005 , n38006 , n38007 , n38008 , n38009 , n38010 , n38011 , n38012 , n38013 , n38014 , n38015 , n38016 , n38017 , n38018 , n38019 , n38020 , n38021 , n38022 , n38023 , n38024 , n38025 , n38026 , n38027 , n38028 , n38029 , n38030 , n38031 , n38032 , n38033 , n38034 , n38035 , n38036 , n38037 , n38038 , n38039 , n38040 , n38041 , n38042 , n38043 , n38044 , n38045 , n38046 , n38047 , n38048 , n38049 , n38050 , n38051 , n38052 , n38053 , n38054 , n38055 , n38056 , n38057 , n38058 , n38059 , n38060 , n38061 , n38062 , n38063 , n38064 , n38065 , n38066 , n38067 , n38068 , n38069 , n38070 , n38071 , n38072 , n38073 , n38074 , n38075 , n38076 , n38077 , n38078 , n38079 , n38080 , n38081 , n38082 , n38083 , n38084 , n38085 , n38086 , n38087 , n38088 , n38089 , n38090 , n38091 , n38092 , n38093 , n38094 , n38095 , n38096 , n38097 , n38098 , n38099 , n38100 , n38101 , n38102 , n38103 , n38104 , n38105 , n38106 , n38107 , n38108 , n38109 , n38110 , n38111 , n38112 , n38113 , n38114 , n38115 , n38116 , n38117 , n38118 , n38119 , n38120 , n38121 , n38122 , n38123 , n38124 , n38125 , n38126 , n38127 , n38128 , n38129 , n38130 , n38131 , n38132 , n38133 , n38134 , n38135 , n38136 , n38137 , n38138 , n38139 , n38140 , n38141 , n38142 , n38143 , n38144 , n38145 , n38146 , n38147 , n38148 , n38149 , n38150 , n38151 , n38152 , n38153 , n38154 , n38155 , n38156 , n38157 , n38158 , n38159 , n38160 , n38161 , n38162 , n38163 , n38164 , n38165 , n38166 , n38167 , n38168 , n38169 , n38170 , n38171 , n38172 , n38173 , n38174 , n38175 , n38176 , n38177 , n38178 , n38179 , n38180 , n38181 , n38182 , n38183 , n38184 , n38185 , n38186 , n38187 , n38188 , n38189 , n38190 , n38191 , n38192 , n38193 , n38194 , n38195 , n38196 , n38197 , n38198 , n38199 , n38200 , n38201 , n38202 , n38203 , n38204 , n38205 , n38206 , n38207 , n38208 , n38209 , n38210 , n38211 , n38212 , n38213 , n38214 , n38215 , n38216 , n38217 , n38218 , n38219 , n38220 , n38221 , n38222 , n38223 , n38224 , n38225 , n38226 , n38227 , n38228 , n38229 , n38230 , n38231 , n38232 , n38233 , n38234 , n38235 , n38236 , n38237 , n38238 , n38239 , n38240 , n38241 , n38242 , n38243 , n38244 , n38245 , n38246 , n38247 , n38248 , n38249 , n38250 , n38251 , n38252 , n38253 , n38254 , n38255 , n38256 , n38257 , n38258 , n38259 , n38260 , n38261 , n38262 , n38263 , n38264 , n38265 , n38266 , n38267 , n38268 , n38269 , n38270 , n38271 , n38272 , n38273 , n38274 , n38275 , n38276 , n38277 , n38278 , n38279 , n38280 , n38281 , n38282 , n38283 , n38284 , n38285 , n38286 , n38287 , n38288 , n38289 , n38290 , n38291 , n38292 , n38293 , n38294 , n38295 , n38296 , n38297 , n38298 , n38299 , n38300 , n38301 , n38302 , n38303 , n38304 , n38305 , n38306 , n38307 , n38308 , n38309 , n38310 , n38311 , n38312 , n38313 , n38314 , n38315 , n38316 , n38317 , n38318 , n38319 , n38320 , n38321 , n38322 , n38323 , n38324 , n38325 , n38326 , n38327 , n38328 , n38329 , n38330 , n38331 , n38332 , n38333 , n38334 , n38335 , n38336 , n38337 , n38338 , n38339 , n38340 , n38341 , n38342 , n38343 , n38344 , n38345 , n38346 , n38347 , n38348 , n38349 , n38350 , n38351 , n38352 , n38353 , n38354 , n38355 , n38356 , n38357 , n38358 , n38359 , n38360 , n38361 , n38362 , n38363 , n38364 , n38365 , n38366 , n38367 , n38368 , n38369 , n38370 , n38371 , n38372 , n38373 , n38374 , n38375 , n38376 , n38377 , n38378 , n38379 , n38380 , n38381 , n38382 , n38383 , n38384 , n38385 , n38386 , n38387 , n38388 , n38389 , n38390 , n38391 , n38392 , n38393 , n38394 , n38395 , n38396 , n38397 , n38398 , n38399 , n38400 , n38401 , n38402 , n38403 , n38404 , n38405 , n38406 , n38407 , n38408 , n38409 , n38410 , n38411 , n38412 , n38413 , n38414 , n38415 , n38416 , n38417 , n38418 , n38419 , n38420 , n38421 , n38422 , n38423 , n38424 , n38425 , n38426 , n38427 , n38428 , n38429 , n38430 , n38431 , n38432 , n38433 , n38434 , n38435 , n38436 , n38437 , n38438 , n38439 , n38440 , n38441 , n38442 , n38443 , n38444 , n38445 , n38446 , n38447 , n38448 , n38449 , n38450 , n38451 , n38452 , n38453 , n38454 , n38455 , n38456 , n38457 , n38458 , n38459 , n38460 , n38461 , n38462 , n38463 , n38464 , n38465 , n38466 , n38467 , n38468 , n38469 , n38470 , n38471 , n38472 , n38473 , n38474 , n38475 , n38476 , n38477 , n38478 , n38479 , n38480 , n38481 , n38482 , n38483 , n38484 , n38485 , n38486 , n38487 , n38488 , n38489 , n38490 , n38491 , n38492 , n38493 , n38494 , n38495 , n38496 , n38497 , n38498 , n38499 , n38500 , n38501 , n38502 , n38503 , n38504 , n38505 , n38506 , n38507 , n38508 , n38509 , n38510 , n38511 , n38512 , n38513 , n38514 , n38515 , n38516 , n38517 , n38518 , n38519 , n38520 , n38521 , n38522 , n38523 , n38524 , n38525 , n38526 , n38527 , n38528 , n38529 , n38530 , n38531 , n38532 , n38533 , n38534 , n38535 , n38536 , n38537 , n38538 , n38539 , n38540 , n38541 , n38542 , n38543 , n38544 , n38545 , n38546 , n38547 , n38548 , n38549 , n38550 , n38551 , n38552 , n38553 , n38554 , n38555 , n38556 , n38557 , n38558 , n38559 , n38560 , n38561 , n38562 , n38563 , n38564 , n38565 , n38566 , n38567 , n38568 , n38569 , n38570 , n38571 , n38572 , n38573 , n38574 , n38575 , n38576 , n38577 , n38578 , n38579 , n38580 , n38581 , n38582 , n38583 , n38584 , n38585 , n38586 , n38587 , n38588 , n38589 , n38590 , n38591 , n38592 , n38593 , n38594 , n38595 , n38596 , n38597 , n38598 , n38599 , n38600 , n38601 , n38602 , n38603 , n38604 , n38605 , n38606 , n38607 , n38608 , n38609 , n38610 , n38611 , n38612 , n38613 , n38614 , n38615 , n38616 , n38617 , n38618 , n38619 , n38620 , n38621 , n38622 , n38623 , n38624 , n38625 , n38626 , n38627 , n38628 , n38629 , n38630 , n38631 , n38632 , n38633 , n38634 , n38635 , n38636 , n38637 , n38638 , n38639 , n38640 , n38641 , n38642 , n38643 , n38644 , n38645 , n38646 , n38647 , n38648 , n38649 , n38650 , n38651 , n38652 , n38653 , n38654 , n38655 , n38656 , n38657 , n38658 , n38659 , n38660 , n38661 , n38662 , n38663 , n38664 , n38665 , n38666 , n38667 , n38668 , n38669 , n38670 , n38671 , n38672 , n38673 , n38674 , n38675 , n38676 , n38677 , n38678 , n38679 , n38680 , n38681 , n38682 , n38683 , n38684 , n38685 , n38686 , n38687 , n38688 , n38689 , n38690 , n38691 , n38692 , n38693 , n38694 , n38695 , n38696 , n38697 , n38698 , n38699 , n38700 , n38701 , n38702 , n38703 , n38704 , n38705 , n38706 , n38707 , n38708 , n38709 , n38710 , n38711 , n38712 , n38713 , n38714 , n38715 , n38716 , n38717 , n38718 , n38719 , n38720 , n38721 , n38722 , n38723 , n38724 , n38725 , n38726 , n38727 , n38728 , n38729 , n38730 , n38731 , n38732 , n38733 , n38734 , n38735 , n38736 , n38737 , n38738 , n38739 , n38740 , n38741 , n38742 , n38743 , n38744 , n38745 , n38746 , n38747 , n38748 , n38749 , n38750 , n38751 , n38752 , n38753 , n38754 , n38755 , n38756 , n38757 , n38758 , n38759 , n38760 , n38761 , n38762 , n38763 , n38764 , n38765 , n38766 , n38767 , n38768 , n38769 , n38770 , n38771 , n38772 , n38773 , n38774 , n38775 , n38776 , n38777 , n38778 , n38779 , n38780 , n38781 , n38782 , n38783 , n38784 , n38785 , n38786 , n38787 , n38788 , n38789 , n38790 , n38791 , n38792 , n38793 , n38794 , n38795 , n38796 , n38797 , n38798 , n38799 , n38800 , n38801 , n38802 , n38803 , n38804 , n38805 , n38806 , n38807 , n38808 , n38809 , n38810 , n38811 , n38812 , n38813 , n38814 , n38815 , n38816 , n38817 , n38818 , n38819 , n38820 , n38821 , n38822 , n38823 , n38824 , n38825 , n38826 , n38827 , n38828 , n38829 , n38830 , n38831 , n38832 , n38833 , n38834 , n38835 , n38836 , n38837 , n38838 , n38839 , n38840 , n38841 , n38842 , n38843 , n38844 , n38845 , n38846 , n38847 , n38848 , n38849 , n38850 , n38851 , n38852 , n38853 , n38854 , n38855 , n38856 , n38857 , n38858 , n38859 , n38860 , n38861 , n38862 , n38863 , n38864 , n38865 , n38866 , n38867 , n38868 , n38869 , n38870 , n38871 , n38872 , n38873 , n38874 , n38875 , n38876 , n38877 , n38878 , n38879 , n38880 , n38881 , n38882 , n38883 , n38884 , n38885 , n38886 , n38887 , n38888 , n38889 , n38890 , n38891 , n38892 , n38893 , n38894 , n38895 , n38896 , n38897 , n38898 , n38899 , n38900 , n38901 , n38902 , n38903 , n38904 , n38905 , n38906 , n38907 , n38908 , n38909 , n38910 , n38911 , n38912 , n38913 , n38914 , n38915 , n38916 , n38917 , n38918 , n38919 , n38920 , n38921 , n38922 , n38923 , n38924 , n38925 , n38926 , n38927 , n38928 , n38929 , n38930 , n38931 , n38932 , n38933 , n38934 , n38935 , n38936 , n38937 , n38938 , n38939 , n38940 , n38941 , n38942 , n38943 , n38944 , n38945 , n38946 , n38947 , n38948 , n38949 , n38950 , n38951 , n38952 , n38953 , n38954 , n38955 , n38956 , n38957 , n38958 , n38959 , n38960 , n38961 , n38962 , n38963 , n38964 , n38965 , n38966 , n38967 , n38968 , n38969 , n38970 , n38971 , n38972 , n38973 , n38974 , n38975 , n38976 , n38977 , n38978 , n38979 , n38980 , n38981 , n38982 , n38983 , n38984 , n38985 , n38986 , n38987 , n38988 , n38989 , n38990 , n38991 , n38992 , n38993 , n38994 , n38995 , n38996 , n38997 , n38998 , n38999 , n39000 , n39001 , n39002 , n39003 , n39004 , n39005 , n39006 , n39007 , n39008 , n39009 , n39010 , n39011 , n39012 , n39013 , n39014 , n39015 , n39016 , n39017 , n39018 , n39019 , n39020 , n39021 , n39022 , n39023 , n39024 , n39025 , n39026 , n39027 , n39028 , n39029 , n39030 , n39031 , n39032 , n39033 , n39034 , n39035 , n39036 , n39037 , n39038 , n39039 , n39040 , n39041 , n39042 , n39043 , n39044 , n39045 , n39046 , n39047 , n39048 , n39049 , n39050 , n39051 , n39052 , n39053 , n39054 , n39055 , n39056 , n39057 , n39058 , n39059 , n39060 , n39061 , n39062 , n39063 , n39064 , n39065 , n39066 , n39067 , n39068 , n39069 , n39070 , n39071 , n39072 , n39073 , n39074 , n39075 , n39076 , n39077 , n39078 , n39079 , n39080 , n39081 , n39082 , n39083 , n39084 , n39085 , n39086 , n39087 , n39088 , n39089 , n39090 , n39091 , n39092 , n39093 , n39094 , n39095 , n39096 , n39097 , n39098 , n39099 , n39100 , n39101 , n39102 , n39103 , n39104 , n39105 , n39106 , n39107 , n39108 , n39109 , n39110 , n39111 , n39112 , n39113 , n39114 , n39115 , n39116 , n39117 , n39118 , n39119 , n39120 , n39121 , n39122 , n39123 , n39124 , n39125 , n39126 , n39127 , n39128 , n39129 , n39130 , n39131 , n39132 , n39133 , n39134 , n39135 , n39136 , n39137 , n39138 , n39139 , n39140 , n39141 , n39142 , n39143 , n39144 , n39145 , n39146 , n39147 , n39148 , n39149 , n39150 , n39151 , n39152 , n39153 , n39154 , n39155 , n39156 , n39157 , n39158 , n39159 , n39160 , n39161 , n39162 , n39163 , n39164 , n39165 , n39166 , n39167 , n39168 , n39169 , n39170 , n39171 , n39172 , n39173 , n39174 , n39175 , n39176 , n39177 , n39178 , n39179 , n39180 , n39181 , n39182 , n39183 , n39184 , n39185 , n39186 , n39187 , n39188 , n39189 , n39190 , n39191 , n39192 , n39193 , n39194 , n39195 , n39196 , n39197 , n39198 , n39199 , n39200 , n39201 , n39202 , n39203 , n39204 , n39205 , n39206 , n39207 , n39208 , n39209 , n39210 , n39211 , n39212 , n39213 , n39214 , n39215 , n39216 , n39217 , n39218 , n39219 , n39220 , n39221 , n39222 , n39223 , n39224 , n39225 , n39226 , n39227 , n39228 , n39229 , n39230 , n39231 , n39232 , n39233 , n39234 , n39235 , n39236 , n39237 , n39238 , n39239 , n39240 , n39241 , n39242 , n39243 , n39244 , n39245 , n39246 , n39247 , n39248 , n39249 , n39250 , n39251 , n39252 , n39253 , n39254 , n39255 , n39256 , n39257 , n39258 , n39259 , n39260 , n39261 , n39262 , n39263 , n39264 , n39265 , n39266 , n39267 , n39268 , n39269 , n39270 , n39271 , n39272 , n39273 , n39274 , n39275 , n39276 , n39277 , n39278 , n39279 , n39280 , n39281 , n39282 , n39283 , n39284 , n39285 , n39286 , n39287 , n39288 , n39289 , n39290 , n39291 , n39292 , n39293 , n39294 , n39295 , n39296 , n39297 , n39298 , n39299 , n39300 , n39301 , n39302 , n39303 , n39304 , n39305 , n39306 , n39307 , n39308 , n39309 , n39310 , n39311 , n39312 , n39313 , n39314 , n39315 , n39316 , n39317 , n39318 , n39319 , n39320 , n39321 , n39322 , n39323 , n39324 , n39325 , n39326 , n39327 , n39328 , n39329 , n39330 , n39331 , n39332 , n39333 , n39334 , n39335 , n39336 , n39337 , n39338 , n39339 , n39340 , n39341 , n39342 , n39343 , n39344 , n39345 , n39346 , n39347 , n39348 , n39349 , n39350 , n39351 , n39352 , n39353 , n39354 , n39355 , n39356 , n39357 , n39358 , n39359 , n39360 , n39361 , n39362 , n39363 , n39364 , n39365 , n39366 , n39367 , n39368 , n39369 , n39370 , n39371 , n39372 , n39373 , n39374 , n39375 , n39376 , n39377 , n39378 , n39379 , n39380 , n39381 , n39382 , n39383 , n39384 , n39385 , n39386 , n39387 , n39388 , n39389 , n39390 , n39391 , n39392 , n39393 , n39394 , n39395 , n39396 , n39397 , n39398 , n39399 , n39400 , n39401 , n39402 , n39403 , n39404 , n39405 , n39406 , n39407 , n39408 , n39409 , n39410 , n39411 , n39412 , n39413 , n39414 , n39415 , n39416 , n39417 , n39418 , n39419 , n39420 , n39421 , n39422 , n39423 , n39424 , n39425 , n39426 , n39427 , n39428 , n39429 , n39430 , n39431 , n39432 , n39433 , n39434 , n39435 , n39436 , n39437 , n39438 , n39439 , n39440 , n39441 , n39442 , n39443 , n39444 , n39445 , n39446 , n39447 , n39448 , n39449 , n39450 , n39451 , n39452 , n39453 , n39454 , n39455 , n39456 , n39457 , n39458 , n39459 , n39460 , n39461 , n39462 , n39463 , n39464 , n39465 , n39466 , n39467 , n39468 , n39469 , n39470 , n39471 , n39472 , n39473 , n39474 , n39475 , n39476 , n39477 , n39478 , n39479 , n39480 , n39481 , n39482 , n39483 , n39484 , n39485 , n39486 , n39487 , n39488 , n39489 , n39490 , n39491 , n39492 , n39493 , n39494 , n39495 , n39496 , n39497 , n39498 , n39499 , n39500 , n39501 , n39502 , n39503 , n39504 , n39505 , n39506 , n39507 , n39508 , n39509 , n39510 , n39511 , n39512 , n39513 , n39514 , n39515 , n39516 , n39517 , n39518 , n39519 , n39520 , n39521 , n39522 , n39523 , n39524 , n39525 , n39526 , n39527 , n39528 , n39529 , n39530 , n39531 , n39532 , n39533 , n39534 , n39535 , n39536 , n39537 , n39538 , n39539 , n39540 , n39541 , n39542 , n39543 , n39544 , n39545 , n39546 , n39547 , n39548 , n39549 , n39550 , n39551 , n39552 , n39553 , n39554 , n39555 , n39556 , n39557 , n39558 , n39559 , n39560 , n39561 , n39562 , n39563 , n39564 , n39565 , n39566 , n39567 , n39568 , n39569 , n39570 , n39571 , n39572 , n39573 , n39574 , n39575 , n39576 , n39577 , n39578 , n39579 , n39580 , n39581 , n39582 , n39583 , n39584 , n39585 , n39586 , n39587 , n39588 , n39589 , n39590 , n39591 , n39592 , n39593 , n39594 , n39595 , n39596 , n39597 , n39598 , n39599 , n39600 , n39601 , n39602 , n39603 , n39604 , n39605 , n39606 , n39607 , n39608 , n39609 , n39610 , n39611 , n39612 , n39613 , n39614 , n39615 , n39616 , n39617 , n39618 , n39619 , n39620 , n39621 , n39622 , n39623 , n39624 , n39625 , n39626 , n39627 , n39628 , n39629 , n39630 , n39631 , n39632 , n39633 , n39634 , n39635 , n39636 , n39637 , n39638 , n39639 , n39640 , n39641 , n39642 , n39643 , n39644 , n39645 , n39646 , n39647 , n39648 , n39649 , n39650 , n39651 , n39652 , n39653 , n39654 , n39655 , n39656 , n39657 , n39658 , n39659 , n39660 , n39661 , n39662 , n39663 , n39664 , n39665 , n39666 , n39667 , n39668 , n39669 , n39670 , n39671 , n39672 , n39673 , n39674 , n39675 , n39676 , n39677 , n39678 , n39679 , n39680 , n39681 , n39682 , n39683 , n39684 , n39685 , n39686 , n39687 , n39688 , n39689 , n39690 , n39691 , n39692 , n39693 , n39694 , n39695 , n39696 , n39697 , n39698 , n39699 , n39700 , n39701 , n39702 , n39703 , n39704 , n39705 , n39706 , n39707 , n39708 , n39709 , n39710 , n39711 , n39712 , n39713 , n39714 , n39715 , n39716 , n39717 , n39718 , n39719 , n39720 , n39721 , n39722 , n39723 , n39724 , n39725 , n39726 , n39727 , n39728 , n39729 , n39730 , n39731 , n39732 , n39733 , n39734 , n39735 , n39736 , n39737 , n39738 , n39739 , n39740 , n39741 , n39742 , n39743 , n39744 , n39745 , n39746 , n39747 , n39748 , n39749 , n39750 , n39751 , n39752 , n39753 , n39754 , n39755 , n39756 , n39757 , n39758 , n39759 , n39760 , n39761 , n39762 , n39763 , n39764 , n39765 , n39766 , n39767 , n39768 , n39769 , n39770 , n39771 , n39772 , n39773 , n39774 , n39775 , n39776 , n39777 , n39778 , n39779 , n39780 , n39781 , n39782 , n39783 , n39784 , n39785 , n39786 , n39787 , n39788 , n39789 , n39790 , n39791 , n39792 , n39793 , n39794 , n39795 , n39796 , n39797 , n39798 , n39799 , n39800 , n39801 , n39802 , n39803 , n39804 , n39805 , n39806 , n39807 , n39808 , n39809 , n39810 , n39811 , n39812 , n39813 , n39814 , n39815 , n39816 , n39817 , n39818 , n39819 , n39820 , n39821 , n39822 , n39823 , n39824 , n39825 , n39826 , n39827 , n39828 , n39829 , n39830 , n39831 , n39832 , n39833 , n39834 , n39835 , n39836 , n39837 , n39838 , n39839 , n39840 , n39841 , n39842 , n39843 , n39844 , n39845 , n39846 , n39847 , n39848 , n39849 , n39850 , n39851 , n39852 , n39853 , n39854 , n39855 , n39856 , n39857 , n39858 , n39859 , n39860 , n39861 , n39862 , n39863 , n39864 , n39865 , n39866 , n39867 , n39868 , n39869 , n39870 , n39871 , n39872 , n39873 , n39874 , n39875 , n39876 , n39877 , n39878 , n39879 , n39880 , n39881 , n39882 , n39883 , n39884 , n39885 , n39886 , n39887 , n39888 , n39889 , n39890 , n39891 , n39892 , n39893 , n39894 , n39895 , n39896 , n39897 , n39898 , n39899 , n39900 , n39901 , n39902 , n39903 , n39904 , n39905 , n39906 , n39907 , n39908 , n39909 , n39910 , n39911 , n39912 , n39913 , n39914 , n39915 , n39916 , n39917 , n39918 , n39919 , n39920 , n39921 , n39922 , n39923 , n39924 , n39925 , n39926 , n39927 , n39928 , n39929 , n39930 , n39931 , n39932 , n39933 , n39934 , n39935 , n39936 , n39937 , n39938 , n39939 , n39940 , n39941 , n39942 , n39943 , n39944 , n39945 , n39946 , n39947 , n39948 , n39949 , n39950 , n39951 , n39952 , n39953 , n39954 , n39955 , n39956 , n39957 , n39958 , n39959 , n39960 , n39961 , n39962 , n39963 , n39964 , n39965 , n39966 , n39967 , n39968 , n39969 , n39970 , n39971 , n39972 , n39973 , n39974 , n39975 , n39976 , n39977 , n39978 , n39979 , n39980 , n39981 , n39982 , n39983 , n39984 , n39985 , n39986 , n39987 , n39988 , n39989 , n39990 , n39991 , n39992 , n39993 , n39994 , n39995 , n39996 , n39997 , n39998 , n39999 , n40000 , n40001 , n40002 , n40003 , n40004 , n40005 , n40006 , n40007 , n40008 , n40009 , n40010 , n40011 , n40012 , n40013 , n40014 , n40015 , n40016 , n40017 , n40018 , n40019 , n40020 , n40021 , n40022 , n40023 , n40024 , n40025 , n40026 , n40027 , n40028 , n40029 , n40030 , n40031 , n40032 , n40033 , n40034 , n40035 , n40036 , n40037 , n40038 , n40039 , n40040 , n40041 , n40042 , n40043 , n40044 , n40045 , n40046 , n40047 , n40048 , n40049 , n40050 , n40051 , n40052 , n40053 , n40054 , n40055 , n40056 , n40057 , n40058 , n40059 , n40060 , n40061 , n40062 , n40063 , n40064 , n40065 , n40066 , n40067 , n40068 , n40069 , n40070 , n40071 , n40072 , n40073 , n40074 , n40075 , n40076 , n40077 , n40078 , n40079 , n40080 , n40081 , n40082 , n40083 , n40084 , n40085 , n40086 , n40087 , n40088 , n40089 , n40090 , n40091 , n40092 , n40093 , n40094 , n40095 , n40096 , n40097 , n40098 , n40099 , n40100 , n40101 , n40102 , n40103 , n40104 , n40105 , n40106 , n40107 , n40108 , n40109 , n40110 , n40111 , n40112 , n40113 , n40114 , n40115 , n40116 , n40117 , n40118 , n40119 , n40120 , n40121 , n40122 , n40123 , n40124 , n40125 , n40126 , n40127 , n40128 , n40129 , n40130 , n40131 , n40132 , n40133 , n40134 , n40135 , n40136 , n40137 , n40138 , n40139 , n40140 , n40141 , n40142 , n40143 , n40144 , n40145 , n40146 , n40147 , n40148 , n40149 , n40150 , n40151 , n40152 , n40153 , n40154 , n40155 , n40156 , n40157 , n40158 , n40159 , n40160 , n40161 , n40162 , n40163 , n40164 , n40165 , n40166 , n40167 , n40168 , n40169 , n40170 , n40171 , n40172 , n40173 , n40174 , n40175 , n40176 , n40177 , n40178 , n40179 , n40180 , n40181 , n40182 , n40183 , n40184 , n40185 , n40186 , n40187 , n40188 , n40189 , n40190 , n40191 , n40192 , n40193 , n40194 , n40195 , n40196 , n40197 , n40198 , n40199 , n40200 , n40201 , n40202 , n40203 , n40204 , n40205 , n40206 , n40207 , n40208 , n40209 , n40210 , n40211 , n40212 , n40213 , n40214 , n40215 , n40216 , n40217 , n40218 , n40219 , n40220 , n40221 , n40222 , n40223 , n40224 , n40225 , n40226 , n40227 , n40228 , n40229 , n40230 , n40231 , n40232 , n40233 , n40234 , n40235 , n40236 , n40237 , n40238 , n40239 , n40240 , n40241 , n40242 , n40243 , n40244 , n40245 , n40246 , n40247 , n40248 , n40249 , n40250 , n40251 , n40252 , n40253 , n40254 , n40255 , n40256 , n40257 , n40258 , n40259 , n40260 , n40261 , n40262 , n40263 , n40264 , n40265 , n40266 , n40267 , n40268 , n40269 , n40270 , n40271 , n40272 , n40273 , n40274 , n40275 , n40276 , n40277 , n40278 , n40279 , n40280 , n40281 , n40282 , n40283 , n40284 , n40285 , n40286 , n40287 , n40288 , n40289 , n40290 , n40291 , n40292 , n40293 , n40294 , n40295 , n40296 , n40297 , n40298 , n40299 , n40300 , n40301 , n40302 , n40303 , n40304 , n40305 , n40306 , n40307 , n40308 , n40309 , n40310 , n40311 , n40312 , n40313 , n40314 , n40315 , n40316 , n40317 , n40318 , n40319 , n40320 , n40321 , n40322 , n40323 , n40324 , n40325 , n40326 , n40327 , n40328 , n40329 , n40330 , n40331 , n40332 , n40333 , n40334 , n40335 , n40336 , n40337 , n40338 , n40339 , n40340 , n40341 , n40342 , n40343 , n40344 , n40345 , n40346 , n40347 , n40348 , n40349 , n40350 , n40351 , n40352 , n40353 , n40354 , n40355 , n40356 , n40357 , n40358 , n40359 , n40360 , n40361 , n40362 , n40363 , n40364 , n40365 , n40366 , n40367 , n40368 , n40369 , n40370 , n40371 , n40372 , n40373 , n40374 , n40375 , n40376 , n40377 , n40378 , n40379 , n40380 , n40381 , n40382 , n40383 , n40384 , n40385 , n40386 , n40387 , n40388 , n40389 , n40390 , n40391 , n40392 , n40393 , n40394 , n40395 , n40396 , n40397 , n40398 , n40399 , n40400 , n40401 , n40402 , n40403 , n40404 , n40405 , n40406 , n40407 , n40408 , n40409 , n40410 , n40411 , n40412 , n40413 , n40414 , n40415 , n40416 , n40417 , n40418 , n40419 , n40420 , n40421 , n40422 , n40423 , n40424 , n40425 , n40426 , n40427 , n40428 , n40429 , n40430 , n40431 , n40432 , n40433 , n40434 , n40435 , n40436 , n40437 , n40438 , n40439 , n40440 , n40441 , n40442 , n40443 , n40444 , n40445 , n40446 , n40447 , n40448 , n40449 , n40450 , n40451 , n40452 , n40453 , n40454 , n40455 , n40456 , n40457 , n40458 , n40459 , n40460 , n40461 , n40462 , n40463 , n40464 , n40465 , n40466 , n40467 , n40468 , n40469 , n40470 , n40471 , n40472 , n40473 , n40474 , n40475 , n40476 , n40477 , n40478 , n40479 , n40480 , n40481 , n40482 , n40483 , n40484 , n40485 , n40486 , n40487 , n40488 , n40489 , n40490 , n40491 , n40492 , n40493 , n40494 , n40495 , n40496 , n40497 , n40498 , n40499 , n40500 , n40501 , n40502 , n40503 , n40504 , n40505 , n40506 , n40507 , n40508 , n40509 , n40510 , n40511 , n40512 , n40513 , n40514 , n40515 , n40516 , n40517 , n40518 , n40519 , n40520 , n40521 , n40522 , n40523 , n40524 , n40525 , n40526 , n40527 , n40528 , n40529 , n40530 , n40531 , n40532 , n40533 , n40534 , n40535 , n40536 , n40537 , n40538 , n40539 , n40540 , n40541 , n40542 , n40543 , n40544 , n40545 , n40546 , n40547 , n40548 , n40549 , n40550 , n40551 , n40552 , n40553 , n40554 , n40555 , n40556 , n40557 , n40558 , n40559 , n40560 , n40561 , n40562 , n40563 , n40564 , n40565 , n40566 , n40567 , n40568 , n40569 , n40570 , n40571 , n40572 , n40573 , n40574 , n40575 , n40576 , n40577 , n40578 , n40579 , n40580 , n40581 , n40582 , n40583 , n40584 , n40585 , n40586 , n40587 , n40588 , n40589 , n40590 , n40591 , n40592 , n40593 , n40594 , n40595 , n40596 , n40597 , n40598 , n40599 , n40600 , n40601 , n40602 , n40603 , n40604 , n40605 , n40606 , n40607 , n40608 , n40609 , n40610 , n40611 , n40612 , n40613 , n40614 , n40615 , n40616 , n40617 , n40618 , n40619 , n40620 , n40621 , n40622 , n40623 , n40624 , n40625 , n40626 , n40627 , n40628 , n40629 , n40630 , n40631 , n40632 , n40633 , n40634 , n40635 , n40636 , n40637 , n40638 , n40639 , n40640 , n40641 , n40642 , n40643 , n40644 , n40645 , n40646 , n40647 , n40648 , n40649 , n40650 , n40651 , n40652 , n40653 , n40654 , n40655 , n40656 , n40657 , n40658 , n40659 , n40660 , n40661 , n40662 , n40663 , n40664 , n40665 , n40666 , n40667 , n40668 , n40669 , n40670 , n40671 , n40672 , n40673 , n40674 , n40675 , n40676 , n40677 , n40678 , n40679 , n40680 , n40681 , n40682 , n40683 , n40684 , n40685 , n40686 , n40687 , n40688 , n40689 , n40690 , n40691 , n40692 , n40693 , n40694 , n40695 , n40696 , n40697 , n40698 , n40699 , n40700 , n40701 , n40702 , n40703 , n40704 , n40705 , n40706 , n40707 , n40708 , n40709 , n40710 , n40711 , n40712 , n40713 , n40714 , n40715 , n40716 , n40717 , n40718 , n40719 , n40720 , n40721 , n40722 , n40723 , n40724 , n40725 , n40726 , n40727 , n40728 , n40729 , n40730 , n40731 , n40732 , n40733 , n40734 , n40735 , n40736 , n40737 , n40738 , n40739 , n40740 , n40741 , n40742 , n40743 , n40744 , n40745 , n40746 , n40747 , n40748 , n40749 , n40750 , n40751 , n40752 , n40753 , n40754 , n40755 , n40756 , n40757 , n40758 , n40759 , n40760 , n40761 , n40762 , n40763 , n40764 , n40765 , n40766 , n40767 , n40768 , n40769 , n40770 , n40771 , n40772 , n40773 , n40774 , n40775 , n40776 , n40777 , n40778 , n40779 , n40780 , n40781 , n40782 , n40783 , n40784 , n40785 , n40786 , n40787 , n40788 , n40789 , n40790 , n40791 , n40792 , n40793 , n40794 , n40795 , n40796 , n40797 , n40798 , n40799 , n40800 , n40801 , n40802 , n40803 , n40804 , n40805 , n40806 , n40807 , n40808 , n40809 , n40810 , n40811 , n40812 , n40813 , n40814 , n40815 , n40816 , n40817 , n40818 , n40819 , n40820 , n40821 , n40822 , n40823 , n40824 , n40825 , n40826 , n40827 , n40828 , n40829 , n40830 , n40831 , n40832 , n40833 , n40834 , n40835 , n40836 , n40837 , n40838 , n40839 , n40840 , n40841 , n40842 , n40843 , n40844 , n40845 , n40846 , n40847 , n40848 , n40849 , n40850 , n40851 , n40852 , n40853 , n40854 , n40855 , n40856 , n40857 , n40858 , n40859 , n40860 , n40861 , n40862 , n40863 , n40864 , n40865 , n40866 , n40867 , n40868 , n40869 , n40870 , n40871 , n40872 , n40873 , n40874 , n40875 , n40876 , n40877 , n40878 , n40879 , n40880 , n40881 , n40882 , n40883 , n40884 , n40885 , n40886 , n40887 , n40888 , n40889 , n40890 , n40891 , n40892 , n40893 , n40894 , n40895 , n40896 , n40897 , n40898 , n40899 , n40900 , n40901 , n40902 , n40903 , n40904 , n40905 , n40906 , n40907 , n40908 , n40909 , n40910 , n40911 , n40912 , n40913 , n40914 , n40915 , n40916 , n40917 , n40918 , n40919 , n40920 , n40921 , n40922 , n40923 , n40924 , n40925 , n40926 , n40927 , n40928 , n40929 , n40930 , n40931 , n40932 , n40933 , n40934 , n40935 , n40936 , n40937 , n40938 , n40939 , n40940 , n40941 , n40942 , n40943 , n40944 , n40945 , n40946 , n40947 , n40948 , n40949 , n40950 , n40951 , n40952 , n40953 , n40954 , n40955 , n40956 , n40957 , n40958 , n40959 , n40960 , n40961 , n40962 , n40963 , n40964 , n40965 , n40966 , n40967 , n40968 , n40969 , n40970 , n40971 , n40972 , n40973 , n40974 , n40975 , n40976 , n40977 , n40978 , n40979 , n40980 , n40981 , n40982 , n40983 , n40984 , n40985 , n40986 , n40987 , n40988 , n40989 , n40990 , n40991 , n40992 , n40993 , n40994 , n40995 , n40996 , n40997 , n40998 , n40999 , n41000 , n41001 , n41002 , n41003 , n41004 , n41005 , n41006 , n41007 , n41008 , n41009 , n41010 , n41011 , n41012 , n41013 , n41014 , n41015 , n41016 , n41017 , n41018 , n41019 , n41020 , n41021 , n41022 , n41023 , n41024 , n41025 , n41026 , n41027 , n41028 , n41029 , n41030 , n41031 , n41032 , n41033 , n41034 , n41035 , n41036 , n41037 , n41038 , n41039 , n41040 , n41041 , n41042 , n41043 , n41044 , n41045 , n41046 , n41047 , n41048 , n41049 , n41050 , n41051 , n41052 , n41053 , n41054 , n41055 , n41056 , n41057 , n41058 , n41059 , n41060 , n41061 , n41062 , n41063 , n41064 , n41065 , n41066 , n41067 , n41068 , n41069 , n41070 , n41071 , n41072 , n41073 , n41074 , n41075 , n41076 , n41077 , n41078 , n41079 , n41080 , n41081 , n41082 , n41083 , n41084 , n41085 , n41086 , n41087 , n41088 , n41089 , n41090 , n41091 , n41092 , n41093 , n41094 , n41095 , n41096 , n41097 , n41098 , n41099 , n41100 , n41101 , n41102 , n41103 , n41104 , n41105 , n41106 , n41107 , n41108 , n41109 , n41110 , n41111 , n41112 , n41113 , n41114 , n41115 , n41116 , n41117 , n41118 , n41119 , n41120 , n41121 , n41122 , n41123 , n41124 , n41125 , n41126 , n41127 , n41128 , n41129 , n41130 , n41131 , n41132 , n41133 , n41134 , n41135 , n41136 , n41137 , n41138 , n41139 , n41140 , n41141 , n41142 , n41143 , n41144 , n41145 , n41146 , n41147 , n41148 , n41149 , n41150 , n41151 , n41152 , n41153 , n41154 , n41155 , n41156 , n41157 , n41158 , n41159 , n41160 , n41161 , n41162 , n41163 , n41164 , n41165 , n41166 , n41167 , n41168 , n41169 , n41170 , n41171 , n41172 , n41173 , n41174 , n41175 , n41176 , n41177 , n41178 , n41179 , n41180 , n41181 , n41182 , n41183 , n41184 , n41185 , n41186 , n41187 , n41188 , n41189 , n41190 , n41191 , n41192 , n41193 , n41194 , n41195 , n41196 , n41197 , n41198 , n41199 , n41200 , n41201 , n41202 , n41203 , n41204 , n41205 , n41206 , n41207 , n41208 , n41209 , n41210 , n41211 , n41212 , n41213 , n41214 , n41215 , n41216 , n41217 , n41218 , n41219 , n41220 , n41221 , n41222 , n41223 , n41224 , n41225 , n41226 , n41227 , n41228 , n41229 , n41230 , n41231 , n41232 , n41233 , n41234 , n41235 , n41236 , n41237 , n41238 , n41239 , n41240 , n41241 , n41242 , n41243 , n41244 , n41245 , n41246 , n41247 , n41248 , n41249 , n41250 , n41251 , n41252 , n41253 , n41254 , n41255 , n41256 , n41257 , n41258 , n41259 , n41260 , n41261 , n41262 , n41263 , n41264 , n41265 , n41266 , n41267 , n41268 , n41269 , n41270 , n41271 , n41272 , n41273 , n41274 , n41275 , n41276 , n41277 , n41278 , n41279 , n41280 , n41281 , n41282 , n41283 , n41284 , n41285 , n41286 , n41287 , n41288 , n41289 , n41290 , n41291 , n41292 , n41293 , n41294 , n41295 , n41296 , n41297 , n41298 , n41299 , n41300 , n41301 , n41302 , n41303 , n41304 , n41305 , n41306 , n41307 , n41308 , n41309 , n41310 , n41311 , n41312 , n41313 , n41314 , n41315 , n41316 , n41317 , n41318 , n41319 , n41320 , n41321 , n41322 , n41323 , n41324 , n41325 , n41326 , n41327 , n41328 , n41329 , n41330 , n41331 , n41332 , n41333 , n41334 , n41335 , n41336 , n41337 , n41338 , n41339 , n41340 , n41341 , n41342 , n41343 , n41344 , n41345 , n41346 , n41347 , n41348 , n41349 , n41350 , n41351 , n41352 , n41353 , n41354 , n41355 , n41356 , n41357 , n41358 , n41359 , n41360 , n41361 , n41362 , n41363 , n41364 , n41365 , n41366 , n41367 , n41368 , n41369 , n41370 , n41371 , n41372 , n41373 , n41374 , n41375 , n41376 , n41377 , n41378 , n41379 , n41380 , n41381 , n41382 , n41383 , n41384 , n41385 , n41386 , n41387 , n41388 , n41389 , n41390 , n41391 , n41392 , n41393 , n41394 , n41395 , n41396 , n41397 , n41398 , n41399 , n41400 , n41401 , n41402 , n41403 , n41404 , n41405 , n41406 , n41407 , n41408 , n41409 , n41410 , n41411 , n41412 , n41413 , n41414 , n41415 , n41416 , n41417 , n41418 , n41419 , n41420 , n41421 , n41422 , n41423 , n41424 , n41425 , n41426 , n41427 , n41428 , n41429 , n41430 , n41431 , n41432 , n41433 , n41434 , n41435 , n41436 , n41437 , n41438 , n41439 , n41440 , n41441 , n41442 , n41443 , n41444 , n41445 , n41446 , n41447 , n41448 , n41449 , n41450 , n41451 , n41452 , n41453 , n41454 , n41455 , n41456 , n41457 , n41458 , n41459 , n41460 , n41461 , n41462 , n41463 , n41464 , n41465 , n41466 , n41467 , n41468 , n41469 , n41470 , n41471 , n41472 , n41473 , n41474 , n41475 , n41476 , n41477 , n41478 , n41479 , n41480 , n41481 , n41482 , n41483 , n41484 , n41485 , n41486 , n41487 , n41488 , n41489 , n41490 , n41491 , n41492 , n41493 , n41494 , n41495 , n41496 , n41497 , n41498 , n41499 , n41500 , n41501 , n41502 , n41503 , n41504 , n41505 , n41506 , n41507 , n41508 , n41509 , n41510 , n41511 , n41512 , n41513 , n41514 , n41515 , n41516 , n41517 , n41518 , n41519 , n41520 , n41521 , n41522 , n41523 , n41524 , n41525 , n41526 , n41527 , n41528 , n41529 , n41530 , n41531 , n41532 , n41533 , n41534 , n41535 , n41536 , n41537 , n41538 , n41539 , n41540 , n41541 , n41542 , n41543 , n41544 , n41545 , n41546 , n41547 , n41548 , n41549 , n41550 , n41551 , n41552 , n41553 , n41554 , n41555 , n41556 , n41557 , n41558 , n41559 , n41560 , n41561 , n41562 , n41563 , n41564 , n41565 , n41566 , n41567 , n41568 , n41569 , n41570 , n41571 , n41572 , n41573 , n41574 , n41575 , n41576 , n41577 , n41578 , n41579 , n41580 , n41581 , n41582 , n41583 , n41584 , n41585 , n41586 , n41587 , n41588 , n41589 , n41590 , n41591 , n41592 , n41593 , n41594 , n41595 , n41596 , n41597 , n41598 , n41599 , n41600 , n41601 , n41602 , n41603 , n41604 , n41605 , n41606 , n41607 , n41608 , n41609 , n41610 , n41611 , n41612 , n41613 , n41614 , n41615 , n41616 , n41617 , n41618 , n41619 , n41620 , n41621 , n41622 , n41623 , n41624 , n41625 , n41626 , n41627 , n41628 , n41629 , n41630 , n41631 , n41632 , n41633 , n41634 , n41635 , n41636 , n41637 , n41638 , n41639 , n41640 , n41641 , n41642 , n41643 , n41644 , n41645 , n41646 , n41647 , n41648 , n41649 , n41650 , n41651 , n41652 , n41653 , n41654 , n41655 , n41656 , n41657 , n41658 , n41659 , n41660 , n41661 , n41662 , n41663 , n41664 , n41665 , n41666 , n41667 , n41668 , n41669 , n41670 , n41671 , n41672 , n41673 , n41674 , n41675 , n41676 , n41677 , n41678 , n41679 , n41680 , n41681 , n41682 , n41683 , n41684 , n41685 , n41686 , n41687 , n41688 , n41689 , n41690 , n41691 , n41692 , n41693 , n41694 , n41695 , n41696 , n41697 , n41698 , n41699 , n41700 , n41701 , n41702 , n41703 , n41704 , n41705 , n41706 , n41707 , n41708 , n41709 , n41710 , n41711 , n41712 , n41713 , n41714 , n41715 , n41716 , n41717 , n41718 , n41719 , n41720 , n41721 , n41722 , n41723 , n41724 , n41725 , n41726 , n41727 , n41728 , n41729 , n41730 , n41731 , n41732 , n41733 , n41734 , n41735 , n41736 , n41737 , n41738 , n41739 , n41740 , n41741 , n41742 , n41743 , n41744 , n41745 , n41746 , n41747 , n41748 , n41749 , n41750 , n41751 , n41752 , n41753 , n41754 , n41755 , n41756 , n41757 , n41758 , n41759 , n41760 , n41761 , n41762 , n41763 , n41764 , n41765 , n41766 , n41767 , n41768 , n41769 , n41770 , n41771 , n41772 , n41773 , n41774 , n41775 , n41776 , n41777 , n41778 , n41779 , n41780 , n41781 , n41782 , n41783 , n41784 , n41785 , n41786 , n41787 , n41788 , n41789 , n41790 , n41791 , n41792 , n41793 , n41794 , n41795 , n41796 , n41797 , n41798 , n41799 , n41800 , n41801 , n41802 , n41803 , n41804 , n41805 , n41806 , n41807 , n41808 , n41809 , n41810 , n41811 , n41812 , n41813 , n41814 , n41815 , n41816 , n41817 , n41818 , n41819 , n41820 , n41821 , n41822 , n41823 , n41824 , n41825 , n41826 , n41827 , n41828 , n41829 , n41830 , n41831 , n41832 , n41833 , n41834 , n41835 , n41836 , n41837 , n41838 , n41839 , n41840 , n41841 , n41842 , n41843 , n41844 , n41845 , n41846 , n41847 , n41848 , n41849 , n41850 , n41851 , n41852 , n41853 , n41854 , n41855 , n41856 , n41857 , n41858 , n41859 , n41860 , n41861 , n41862 , n41863 , n41864 , n41865 , n41866 , n41867 , n41868 , n41869 , n41870 , n41871 , n41872 , n41873 , n41874 , n41875 , n41876 , n41877 , n41878 , n41879 , n41880 , n41881 , n41882 , n41883 , n41884 , n41885 , n41886 , n41887 , n41888 , n41889 , n41890 , n41891 , n41892 , n41893 , n41894 , n41895 , n41896 , n41897 , n41898 , n41899 , n41900 , n41901 , n41902 , n41903 , n41904 , n41905 , n41906 , n41907 , n41908 , n41909 , n41910 , n41911 , n41912 , n41913 , n41914 , n41915 , n41916 , n41917 , n41918 , n41919 , n41920 , n41921 , n41922 , n41923 , n41924 , n41925 , n41926 , n41927 , n41928 , n41929 , n41930 , n41931 , n41932 , n41933 , n41934 , n41935 , n41936 , n41937 , n41938 , n41939 , n41940 , n41941 , n41942 , n41943 , n41944 , n41945 , n41946 , n41947 , n41948 , n41949 , n41950 , n41951 , n41952 , n41953 , n41954 , n41955 , n41956 , n41957 , n41958 , n41959 , n41960 , n41961 , n41962 , n41963 , n41964 , n41965 , n41966 , n41967 , n41968 , n41969 , n41970 , n41971 , n41972 , n41973 , n41974 , n41975 , n41976 , n41977 , n41978 , n41979 , n41980 , n41981 , n41982 , n41983 , n41984 , n41985 , n41986 , n41987 , n41988 , n41989 , n41990 , n41991 , n41992 , n41993 , n41994 , n41995 , n41996 , n41997 , n41998 , n41999 , n42000 , n42001 , n42002 , n42003 , n42004 , n42005 , n42006 , n42007 , n42008 , n42009 , n42010 , n42011 , n42012 , n42013 , n42014 , n42015 , n42016 , n42017 , n42018 , n42019 , n42020 , n42021 , n42022 , n42023 , n42024 , n42025 , n42026 , n42027 , n42028 , n42029 , n42030 , n42031 , n42032 , n42033 , n42034 , n42035 , n42036 , n42037 , n42038 , n42039 , n42040 , n42041 , n42042 , n42043 , n42044 , n42045 , n42046 , n42047 , n42048 , n42049 , n42050 , n42051 , n42052 , n42053 , n42054 , n42055 , n42056 , n42057 , n42058 , n42059 , n42060 , n42061 , n42062 , n42063 , n42064 , n42065 , n42066 , n42067 , n42068 , n42069 , n42070 , n42071 , n42072 , n42073 , n42074 , n42075 , n42076 , n42077 , n42078 , n42079 , n42080 , n42081 , n42082 , n42083 , n42084 , n42085 , n42086 , n42087 , n42088 , n42089 , n42090 , n42091 , n42092 , n42093 , n42094 , n42095 , n42096 , n42097 , n42098 , n42099 , n42100 , n42101 , n42102 , n42103 , n42104 , n42105 , n42106 , n42107 , n42108 , n42109 , n42110 , n42111 , n42112 , n42113 , n42114 , n42115 , n42116 , n42117 , n42118 , n42119 , n42120 , n42121 , n42122 , n42123 , n42124 , n42125 , n42126 , n42127 , n42128 , n42129 , n42130 , n42131 , n42132 , n42133 , n42134 , n42135 , n42136 , n42137 , n42138 , n42139 , n42140 , n42141 , n42142 , n42143 , n42144 , n42145 , n42146 , n42147 , n42148 , n42149 , n42150 , n42151 , n42152 , n42153 , n42154 , n42155 , n42156 , n42157 , n42158 , n42159 , n42160 , n42161 , n42162 , n42163 , n42164 , n42165 , n42166 , n42167 , n42168 , n42169 , n42170 , n42171 , n42172 , n42173 , n42174 , n42175 , n42176 , n42177 , n42178 , n42179 , n42180 , n42181 , n42182 , n42183 , n42184 , n42185 , n42186 , n42187 , n42188 , n42189 , n42190 , n42191 , n42192 , n42193 , n42194 , n42195 , n42196 , n42197 , n42198 , n42199 , n42200 , n42201 , n42202 , n42203 , n42204 , n42205 , n42206 , n42207 , n42208 , n42209 , n42210 , n42211 , n42212 , n42213 , n42214 , n42215 , n42216 , n42217 , n42218 , n42219 , n42220 , n42221 , n42222 , n42223 , n42224 , n42225 , n42226 , n42227 , n42228 , n42229 , n42230 , n42231 , n42232 , n42233 , n42234 , n42235 , n42236 , n42237 , n42238 , n42239 , n42240 , n42241 , n42242 , n42243 , n42244 , n42245 , n42246 , n42247 , n42248 , n42249 , n42250 , n42251 , n42252 , n42253 , n42254 , n42255 , n42256 , n42257 , n42258 , n42259 , n42260 , n42261 , n42262 , n42263 , n42264 , n42265 , n42266 , n42267 , n42268 , n42269 , n42270 , n42271 , n42272 , n42273 , n42274 , n42275 , n42276 , n42277 , n42278 , n42279 , n42280 , n42281 , n42282 , n42283 , n42284 , n42285 , n42286 , n42287 , n42288 , n42289 , n42290 , n42291 , n42292 , n42293 , n42294 , n42295 , n42296 , n42297 , n42298 , n42299 , n42300 , n42301 , n42302 , n42303 , n42304 , n42305 , n42306 , n42307 , n42308 , n42309 , n42310 , n42311 , n42312 , n42313 , n42314 , n42315 , n42316 , n42317 , n42318 , n42319 , n42320 , n42321 , n42322 , n42323 , n42324 , n42325 , n42326 , n42327 , n42328 , n42329 , n42330 , n42331 , n42332 , n42333 , n42334 , n42335 , n42336 , n42337 , n42338 , n42339 , n42340 , n42341 , n42342 , n42343 , n42344 , n42345 , n42346 , n42347 , n42348 , n42349 , n42350 , n42351 , n42352 , n42353 , n42354 , n42355 , n42356 , n42357 , n42358 , n42359 , n42360 , n42361 , n42362 , n42363 , n42364 , n42365 , n42366 , n42367 , n42368 , n42369 , n42370 , n42371 , n42372 , n42373 , n42374 , n42375 , n42376 , n42377 , n42378 , n42379 , n42380 , n42381 , n42382 , n42383 , n42384 , n42385 , n42386 , n42387 , n42388 , n42389 , n42390 , n42391 , n42392 , n42393 , n42394 , n42395 , n42396 , n42397 , n42398 , n42399 , n42400 , n42401 , n42402 , n42403 , n42404 , n42405 , n42406 , n42407 , n42408 , n42409 , n42410 , n42411 , n42412 , n42413 , n42414 , n42415 , n42416 , n42417 , n42418 , n42419 , n42420 , n42421 , n42422 , n42423 , n42424 , n42425 , n42426 , n42427 , n42428 , n42429 , n42430 , n42431 , n42432 , n42433 , n42434 , n42435 , n42436 , n42437 , n42438 , n42439 , n42440 , n42441 , n42442 , n42443 , n42444 , n42445 , n42446 , n42447 , n42448 , n42449 , n42450 , n42451 , n42452 , n42453 , n42454 , n42455 , n42456 , n42457 , n42458 , n42459 , n42460 , n42461 , n42462 , n42463 , n42464 , n42465 , n42466 , n42467 , n42468 , n42469 , n42470 , n42471 , n42472 , n42473 , n42474 , n42475 , n42476 , n42477 , n42478 , n42479 , n42480 , n42481 , n42482 , n42483 , n42484 , n42485 , n42486 , n42487 , n42488 , n42489 , n42490 , n42491 , n42492 , n42493 , n42494 , n42495 , n42496 , n42497 , n42498 , n42499 , n42500 , n42501 , n42502 , n42503 , n42504 , n42505 , n42506 , n42507 , n42508 , n42509 , n42510 , n42511 , n42512 , n42513 , n42514 , n42515 , n42516 , n42517 , n42518 , n42519 , n42520 , n42521 , n42522 , n42523 , n42524 , n42525 , n42526 , n42527 , n42528 , n42529 , n42530 , n42531 , n42532 , n42533 , n42534 , n42535 , n42536 , n42537 , n42538 , n42539 , n42540 , n42541 , n42542 , n42543 , n42544 , n42545 , n42546 , n42547 , n42548 , n42549 , n42550 , n42551 , n42552 , n42553 , n42554 , n42555 , n42556 , n42557 , n42558 , n42559 , n42560 , n42561 , n42562 , n42563 , n42564 , n42565 , n42566 , n42567 , n42568 , n42569 , n42570 , n42571 , n42572 , n42573 , n42574 , n42575 , n42576 , n42577 , n42578 , n42579 , n42580 , n42581 , n42582 , n42583 , n42584 , n42585 , n42586 , n42587 , n42588 , n42589 , n42590 , n42591 , n42592 , n42593 , n42594 , n42595 , n42596 , n42597 , n42598 , n42599 , n42600 , n42601 , n42602 , n42603 , n42604 , n42605 , n42606 , n42607 , n42608 , n42609 , n42610 , n42611 , n42612 , n42613 , n42614 , n42615 , n42616 , n42617 , n42618 , n42619 , n42620 , n42621 , n42622 , n42623 , n42624 , n42625 , n42626 , n42627 , n42628 , n42629 , n42630 , n42631 , n42632 , n42633 , n42634 , n42635 , n42636 , n42637 , n42638 , n42639 , n42640 , n42641 , n42642 , n42643 , n42644 , n42645 , n42646 , n42647 , n42648 , n42649 , n42650 , n42651 , n42652 , n42653 , n42654 , n42655 , n42656 , n42657 , n42658 , n42659 , n42660 , n42661 , n42662 , n42663 , n42664 , n42665 , n42666 , n42667 , n42668 , n42669 , n42670 , n42671 , n42672 , n42673 , n42674 , n42675 , n42676 , n42677 , n42678 , n42679 , n42680 , n42681 , n42682 , n42683 , n42684 , n42685 , n42686 , n42687 , n42688 , n42689 , n42690 , n42691 , n42692 , n42693 , n42694 , n42695 , n42696 , n42697 , n42698 , n42699 , n42700 , n42701 , n42702 , n42703 , n42704 , n42705 , n42706 , n42707 , n42708 , n42709 , n42710 , n42711 , n42712 , n42713 , n42714 , n42715 , n42716 , n42717 , n42718 , n42719 , n42720 , n42721 , n42722 , n42723 , n42724 , n42725 , n42726 , n42727 , n42728 , n42729 , n42730 , n42731 , n42732 , n42733 , n42734 , n42735 , n42736 , n42737 , n42738 , n42739 , n42740 , n42741 , n42742 , n42743 , n42744 , n42745 , n42746 , n42747 , n42748 , n42749 , n42750 , n42751 , n42752 , n42753 , n42754 , n42755 , n42756 , n42757 , n42758 , n42759 , n42760 , n42761 , n42762 , n42763 , n42764 , n42765 , n42766 , n42767 , n42768 , n42769 , n42770 , n42771 , n42772 , n42773 , n42774 , n42775 , n42776 , n42777 , n42778 , n42779 , n42780 , n42781 , n42782 , n42783 , n42784 , n42785 , n42786 , n42787 , n42788 , n42789 , n42790 , n42791 , n42792 , n42793 , n42794 , n42795 , n42796 , n42797 , n42798 , n42799 , n42800 , n42801 , n42802 , n42803 , n42804 , n42805 , n42806 , n42807 , n42808 , n42809 , n42810 , n42811 , n42812 , n42813 , n42814 , n42815 , n42816 , n42817 , n42818 , n42819 , n42820 , n42821 , n42822 , n42823 , n42824 , n42825 , n42826 , n42827 , n42828 , n42829 , n42830 , n42831 , n42832 , n42833 , n42834 , n42835 , n42836 , n42837 , n42838 , n42839 , n42840 , n42841 , n42842 , n42843 , n42844 , n42845 , n42846 , n42847 , n42848 , n42849 , n42850 , n42851 , n42852 , n42853 , n42854 , n42855 , n42856 , n42857 , n42858 , n42859 , n42860 , n42861 , n42862 , n42863 , n42864 , n42865 , n42866 , n42867 , n42868 , n42869 , n42870 , n42871 , n42872 , n42873 , n42874 , n42875 , n42876 , n42877 , n42878 , n42879 , n42880 , n42881 , n42882 , n42883 , n42884 , n42885 , n42886 , n42887 , n42888 , n42889 , n42890 , n42891 , n42892 , n42893 , n42894 , n42895 , n42896 , n42897 , n42898 , n42899 , n42900 , n42901 , n42902 , n42903 , n42904 , n42905 , n42906 , n42907 , n42908 , n42909 , n42910 , n42911 , n42912 , n42913 , n42914 , n42915 , n42916 , n42917 , n42918 , n42919 , n42920 , n42921 , n42922 , n42923 , n42924 , n42925 , n42926 , n42927 , n42928 , n42929 , n42930 , n42931 , n42932 , n42933 , n42934 , n42935 , n42936 , n42937 , n42938 , n42939 , n42940 , n42941 , n42942 , n42943 , n42944 , n42945 , n42946 , n42947 , n42948 , n42949 , n42950 , n42951 , n42952 , n42953 , n42954 , n42955 , n42956 , n42957 , n42958 , n42959 , n42960 , n42961 , n42962 , n42963 , n42964 , n42965 , n42966 , n42967 , n42968 , n42969 , n42970 , n42971 , n42972 , n42973 , n42974 , n42975 , n42976 , n42977 , n42978 , n42979 , n42980 , n42981 , n42982 , n42983 , n42984 , n42985 , n42986 , n42987 , n42988 , n42989 , n42990 , n42991 , n42992 , n42993 , n42994 , n42995 , n42996 , n42997 , n42998 , n42999 , n43000 , n43001 , n43002 , n43003 , n43004 , n43005 , n43006 , n43007 , n43008 , n43009 , n43010 , n43011 , n43012 , n43013 , n43014 , n43015 , n43016 , n43017 , n43018 , n43019 , n43020 , n43021 , n43022 , n43023 , n43024 , n43025 , n43026 , n43027 , n43028 , n43029 , n43030 , n43031 , n43032 , n43033 , n43034 , n43035 , n43036 , n43037 , n43038 , n43039 , n43040 , n43041 , n43042 , n43043 , n43044 , n43045 , n43046 , n43047 , n43048 , n43049 , n43050 , n43051 , n43052 , n43053 , n43054 , n43055 , n43056 , n43057 , n43058 , n43059 , n43060 , n43061 , n43062 , n43063 , n43064 , n43065 , n43066 , n43067 , n43068 , n43069 , n43070 , n43071 , n43072 , n43073 , n43074 , n43075 , n43076 , n43077 , n43078 , n43079 , n43080 , n43081 , n43082 , n43083 , n43084 , n43085 , n43086 , n43087 , n43088 , n43089 , n43090 , n43091 , n43092 , n43093 , n43094 , n43095 , n43096 , n43097 , n43098 , n43099 , n43100 , n43101 , n43102 , n43103 , n43104 , n43105 , n43106 , n43107 , n43108 , n43109 , n43110 , n43111 , n43112 , n43113 , n43114 , n43115 , n43116 , n43117 , n43118 , n43119 , n43120 , n43121 , n43122 , n43123 , n43124 , n43125 , n43126 , n43127 , n43128 , n43129 , n43130 , n43131 , n43132 , n43133 , n43134 , n43135 , n43136 , n43137 , n43138 , n43139 , n43140 , n43141 , n43142 , n43143 , n43144 , n43145 , n43146 , n43147 , n43148 , n43149 , n43150 , n43151 , n43152 , n43153 , n43154 , n43155 , n43156 , n43157 , n43158 , n43159 , n43160 , n43161 , n43162 , n43163 , n43164 , n43165 , n43166 , n43167 , n43168 , n43169 , n43170 , n43171 , n43172 , n43173 , n43174 , n43175 , n43176 , n43177 , n43178 , n43179 , n43180 , n43181 , n43182 , n43183 , n43184 , n43185 , n43186 , n43187 , n43188 , n43189 , n43190 , n43191 , n43192 , n43193 , n43194 , n43195 , n43196 , n43197 , n43198 , n43199 , n43200 , n43201 , n43202 , n43203 , n43204 , n43205 , n43206 , n43207 , n43208 , n43209 , n43210 , n43211 , n43212 , n43213 , n43214 , n43215 , n43216 , n43217 , n43218 , n43219 , n43220 , n43221 , n43222 , n43223 , n43224 , n43225 , n43226 , n43227 , n43228 , n43229 , n43230 , n43231 , n43232 , n43233 , n43234 , n43235 , n43236 , n43237 , n43238 , n43239 , n43240 , n43241 , n43242 , n43243 , n43244 , n43245 , n43246 , n43247 , n43248 , n43249 , n43250 , n43251 , n43252 , n43253 , n43254 , n43255 , n43256 , n43257 , n43258 , n43259 , n43260 , n43261 , n43262 , n43263 , n43264 , n43265 , n43266 , n43267 , n43268 , n43269 , n43270 , n43271 , n43272 , n43273 , n43274 , n43275 , n43276 , n43277 , n43278 , n43279 , n43280 , n43281 , n43282 , n43283 , n43284 , n43285 , n43286 , n43287 , n43288 , n43289 , n43290 , n43291 , n43292 , n43293 , n43294 , n43295 , n43296 , n43297 , n43298 , n43299 , n43300 , n43301 , n43302 , n43303 , n43304 , n43305 , n43306 , n43307 , n43308 , n43309 , n43310 , n43311 , n43312 , n43313 , n43314 , n43315 , n43316 , n43317 , n43318 , n43319 , n43320 , n43321 , n43322 , n43323 , n43324 , n43325 , n43326 , n43327 , n43328 , n43329 , n43330 , n43331 , n43332 , n43333 , n43334 , n43335 , n43336 , n43337 , n43338 , n43339 , n43340 , n43341 , n43342 , n43343 , n43344 , n43345 , n43346 , n43347 , n43348 , n43349 , n43350 , n43351 , n43352 , n43353 , n43354 , n43355 , n43356 , n43357 , n43358 , n43359 , n43360 , n43361 , n43362 , n43363 , n43364 , n43365 , n43366 , n43367 , n43368 , n43369 , n43370 , n43371 , n43372 , n43373 , n43374 , n43375 , n43376 , n43377 , n43378 , n43379 , n43380 , n43381 , n43382 , n43383 , n43384 , n43385 , n43386 , n43387 , n43388 , n43389 , n43390 , n43391 , n43392 , n43393 , n43394 , n43395 , n43396 , n43397 , n43398 , n43399 , n43400 , n43401 , n43402 , n43403 , n43404 , n43405 , n43406 , n43407 , n43408 , n43409 , n43410 , n43411 , n43412 , n43413 , n43414 , n43415 , n43416 , n43417 , n43418 , n43419 , n43420 , n43421 , n43422 , n43423 , n43424 , n43425 , n43426 , n43427 , n43428 , n43429 , n43430 , n43431 , n43432 , n43433 , n43434 , n43435 , n43436 , n43437 , n43438 , n43439 , n43440 , n43441 , n43442 , n43443 , n43444 , n43445 , n43446 , n43447 , n43448 , n43449 , n43450 , n43451 , n43452 , n43453 , n43454 , n43455 , n43456 , n43457 , n43458 , n43459 , n43460 , n43461 , n43462 , n43463 , n43464 , n43465 , n43466 , n43467 , n43468 , n43469 , n43470 , n43471 , n43472 , n43473 , n43474 , n43475 , n43476 , n43477 , n43478 , n43479 , n43480 , n43481 , n43482 , n43483 , n43484 , n43485 , n43486 , n43487 , n43488 , n43489 , n43490 , n43491 , n43492 , n43493 , n43494 , n43495 , n43496 , n43497 , n43498 , n43499 , n43500 , n43501 , n43502 , n43503 , n43504 , n43505 , n43506 , n43507 , n43508 , n43509 , n43510 , n43511 , n43512 , n43513 , n43514 , n43515 , n43516 , n43517 , n43518 , n43519 , n43520 , n43521 , n43522 , n43523 , n43524 , n43525 , n43526 , n43527 , n43528 , n43529 , n43530 , n43531 , n43532 , n43533 , n43534 , n43535 , n43536 , n43537 , n43538 , n43539 , n43540 , n43541 , n43542 , n43543 , n43544 , n43545 , n43546 , n43547 , n43548 , n43549 , n43550 , n43551 , n43552 , n43553 , n43554 , n43555 , n43556 , n43557 , n43558 , n43559 , n43560 , n43561 , n43562 , n43563 , n43564 , n43565 , n43566 , n43567 , n43568 , n43569 , n43570 , n43571 , n43572 , n43573 , n43574 , n43575 , n43576 , n43577 , n43578 , n43579 , n43580 , n43581 , n43582 , n43583 , n43584 , n43585 , n43586 , n43587 , n43588 , n43589 , n43590 , n43591 , n43592 , n43593 , n43594 , n43595 , n43596 , n43597 , n43598 , n43599 , n43600 , n43601 , n43602 , n43603 , n43604 , n43605 , n43606 , n43607 , n43608 , n43609 , n43610 , n43611 , n43612 , n43613 , n43614 , n43615 , n43616 , n43617 , n43618 , n43619 , n43620 , n43621 , n43622 , n43623 , n43624 , n43625 , n43626 , n43627 , n43628 , n43629 , n43630 , n43631 , n43632 , n43633 , n43634 , n43635 , n43636 , n43637 , n43638 , n43639 , n43640 , n43641 , n43642 , n43643 , n43644 , n43645 , n43646 , n43647 , n43648 , n43649 , n43650 , n43651 , n43652 , n43653 , n43654 , n43655 , n43656 , n43657 , n43658 , n43659 , n43660 , n43661 , n43662 , n43663 , n43664 , n43665 , n43666 , n43667 , n43668 , n43669 , n43670 , n43671 , n43672 , n43673 , n43674 , n43675 , n43676 , n43677 , n43678 , n43679 , n43680 , n43681 , n43682 , n43683 , n43684 , n43685 , n43686 , n43687 , n43688 , n43689 , n43690 , n43691 , n43692 , n43693 , n43694 , n43695 , n43696 , n43697 , n43698 , n43699 , n43700 , n43701 , n43702 , n43703 , n43704 , n43705 , n43706 , n43707 , n43708 , n43709 , n43710 , n43711 , n43712 , n43713 , n43714 , n43715 , n43716 , n43717 , n43718 , n43719 , n43720 , n43721 , n43722 , n43723 , n43724 , n43725 , n43726 , n43727 , n43728 , n43729 , n43730 , n43731 , n43732 , n43733 , n43734 , n43735 , n43736 , n43737 , n43738 , n43739 , n43740 , n43741 , n43742 , n43743 , n43744 , n43745 , n43746 , n43747 , n43748 , n43749 , n43750 , n43751 , n43752 , n43753 , n43754 , n43755 , n43756 , n43757 , n43758 , n43759 , n43760 , n43761 , n43762 , n43763 , n43764 , n43765 , n43766 , n43767 , n43768 , n43769 , n43770 , n43771 , n43772 , n43773 , n43774 , n43775 , n43776 , n43777 , n43778 , n43779 , n43780 , n43781 , n43782 , n43783 , n43784 , n43785 , n43786 , n43787 , n43788 , n43789 , n43790 , n43791 , n43792 , n43793 , n43794 , n43795 , n43796 , n43797 , n43798 , n43799 , n43800 , n43801 , n43802 , n43803 , n43804 , n43805 , n43806 , n43807 , n43808 , n43809 , n43810 , n43811 , n43812 , n43813 , n43814 , n43815 , n43816 , n43817 , n43818 , n43819 , n43820 , n43821 , n43822 , n43823 , n43824 , n43825 , n43826 , n43827 , n43828 , n43829 , n43830 , n43831 , n43832 , n43833 , n43834 , n43835 , n43836 , n43837 , n43838 , n43839 , n43840 , n43841 , n43842 , n43843 , n43844 , n43845 , n43846 , n43847 , n43848 , n43849 , n43850 , n43851 , n43852 , n43853 , n43854 , n43855 , n43856 , n43857 , n43858 , n43859 , n43860 , n43861 , n43862 , n43863 , n43864 , n43865 , n43866 , n43867 , n43868 , n43869 , n43870 , n43871 , n43872 , n43873 , n43874 , n43875 , n43876 , n43877 , n43878 , n43879 , n43880 , n43881 , n43882 , n43883 , n43884 , n43885 , n43886 , n43887 , n43888 , n43889 , n43890 , n43891 , n43892 , n43893 , n43894 , n43895 , n43896 , n43897 , n43898 , n43899 , n43900 , n43901 , n43902 , n43903 , n43904 , n43905 , n43906 , n43907 , n43908 , n43909 , n43910 , n43911 , n43912 , n43913 , n43914 , n43915 , n43916 , n43917 , n43918 , n43919 , n43920 , n43921 , n43922 , n43923 , n43924 , n43925 , n43926 , n43927 , n43928 , n43929 , n43930 , n43931 , n43932 , n43933 , n43934 , n43935 , n43936 , n43937 , n43938 , n43939 , n43940 , n43941 , n43942 , n43943 , n43944 , n43945 , n43946 , n43947 , n43948 , n43949 , n43950 , n43951 , n43952 , n43953 , n43954 , n43955 , n43956 , n43957 , n43958 , n43959 , n43960 , n43961 , n43962 , n43963 , n43964 , n43965 , n43966 , n43967 , n43968 , n43969 , n43970 , n43971 , n43972 , n43973 , n43974 , n43975 , n43976 , n43977 , n43978 , n43979 , n43980 , n43981 , n43982 , n43983 , n43984 , n43985 , n43986 , n43987 , n43988 , n43989 , n43990 , n43991 , n43992 , n43993 , n43994 , n43995 , n43996 , n43997 , n43998 , n43999 , n44000 , n44001 , n44002 , n44003 , n44004 , n44005 , n44006 , n44007 , n44008 , n44009 , n44010 , n44011 , n44012 , n44013 , n44014 , n44015 , n44016 , n44017 , n44018 , n44019 , n44020 , n44021 , n44022 , n44023 , n44024 , n44025 , n44026 , n44027 , n44028 , n44029 , n44030 , n44031 , n44032 , n44033 , n44034 , n44035 , n44036 , n44037 , n44038 , n44039 , n44040 , n44041 , n44042 , n44043 , n44044 , n44045 , n44046 , n44047 , n44048 , n44049 , n44050 , n44051 , n44052 , n44053 , n44054 , n44055 , n44056 , n44057 , n44058 , n44059 , n44060 , n44061 , n44062 , n44063 , n44064 , n44065 , n44066 , n44067 , n44068 , n44069 , n44070 , n44071 , n44072 , n44073 , n44074 , n44075 , n44076 , n44077 , n44078 , n44079 , n44080 , n44081 , n44082 , n44083 , n44084 , n44085 , n44086 , n44087 , n44088 , n44089 , n44090 , n44091 , n44092 , n44093 , n44094 , n44095 , n44096 , n44097 , n44098 , n44099 , n44100 , n44101 , n44102 , n44103 , n44104 , n44105 , n44106 , n44107 , n44108 , n44109 , n44110 , n44111 , n44112 , n44113 , n44114 , n44115 , n44116 , n44117 , n44118 , n44119 , n44120 , n44121 , n44122 , n44123 , n44124 , n44125 , n44126 , n44127 , n44128 , n44129 , n44130 , n44131 , n44132 , n44133 , n44134 , n44135 , n44136 , n44137 , n44138 , n44139 , n44140 , n44141 , n44142 , n44143 , n44144 , n44145 , n44146 , n44147 , n44148 , n44149 , n44150 , n44151 , n44152 , n44153 , n44154 , n44155 , n44156 , n44157 , n44158 , n44159 , n44160 , n44161 , n44162 , n44163 , n44164 , n44165 , n44166 , n44167 , n44168 , n44169 , n44170 , n44171 , n44172 , n44173 , n44174 , n44175 , n44176 , n44177 , n44178 , n44179 , n44180 , n44181 , n44182 , n44183 , n44184 , n44185 , n44186 , n44187 , n44188 , n44189 , n44190 , n44191 , n44192 , n44193 , n44194 , n44195 , n44196 , n44197 , n44198 , n44199 , n44200 , n44201 , n44202 , n44203 , n44204 , n44205 , n44206 , n44207 , n44208 , n44209 , n44210 , n44211 , n44212 , n44213 , n44214 , n44215 , n44216 , n44217 , n44218 , n44219 , n44220 , n44221 , n44222 , n44223 , n44224 , n44225 , n44226 , n44227 , n44228 , n44229 , n44230 , n44231 , n44232 , n44233 , n44234 , n44235 , n44236 , n44237 , n44238 , n44239 , n44240 , n44241 , n44242 , n44243 , n44244 , n44245 , n44246 , n44247 , n44248 , n44249 , n44250 , n44251 , n44252 , n44253 , n44254 , n44255 , n44256 , n44257 , n44258 , n44259 , n44260 , n44261 , n44262 , n44263 , n44264 , n44265 , n44266 , n44267 , n44268 , n44269 , n44270 , n44271 , n44272 , n44273 , n44274 , n44275 , n44276 , n44277 , n44278 , n44279 , n44280 , n44281 , n44282 , n44283 , n44284 , n44285 , n44286 , n44287 , n44288 , n44289 , n44290 , n44291 , n44292 , n44293 , n44294 , n44295 , n44296 , n44297 , n44298 , n44299 , n44300 , n44301 , n44302 , n44303 , n44304 , n44305 , n44306 , n44307 , n44308 , n44309 , n44310 , n44311 , n44312 , n44313 , n44314 , n44315 , n44316 , n44317 , n44318 , n44319 , n44320 , n44321 , n44322 , n44323 , n44324 , n44325 , n44326 , n44327 , n44328 , n44329 , n44330 , n44331 , n44332 , n44333 , n44334 , n44335 , n44336 , n44337 , n44338 , n44339 , n44340 , n44341 , n44342 , n44343 , n44344 , n44345 , n44346 , n44347 , n44348 , n44349 , n44350 , n44351 , n44352 , n44353 , n44354 , n44355 , n44356 , n44357 , n44358 , n44359 , n44360 , n44361 , n44362 , n44363 , n44364 , n44365 , n44366 , n44367 , n44368 , n44369 , n44370 , n44371 , n44372 , n44373 , n44374 , n44375 , n44376 , n44377 , n44378 , n44379 , n44380 , n44381 , n44382 , n44383 , n44384 , n44385 , n44386 , n44387 , n44388 , n44389 , n44390 , n44391 , n44392 , n44393 , n44394 , n44395 , n44396 , n44397 , n44398 , n44399 , n44400 , n44401 , n44402 , n44403 , n44404 , n44405 , n44406 , n44407 , n44408 , n44409 , n44410 , n44411 , n44412 , n44413 , n44414 , n44415 , n44416 , n44417 , n44418 , n44419 , n44420 , n44421 , n44422 , n44423 , n44424 , n44425 , n44426 , n44427 , n44428 , n44429 , n44430 , n44431 , n44432 , n44433 , n44434 , n44435 , n44436 , n44437 , n44438 , n44439 , n44440 , n44441 , n44442 , n44443 , n44444 , n44445 , n44446 , n44447 , n44448 , n44449 , n44450 , n44451 , n44452 , n44453 , n44454 , n44455 , n44456 , n44457 , n44458 , n44459 , n44460 , n44461 , n44462 , n44463 , n44464 , n44465 , n44466 , n44467 , n44468 , n44469 , n44470 , n44471 , n44472 , n44473 , n44474 , n44475 , n44476 , n44477 , n44478 , n44479 , n44480 , n44481 , n44482 , n44483 , n44484 , n44485 , n44486 , n44487 , n44488 , n44489 , n44490 , n44491 , n44492 , n44493 , n44494 , n44495 , n44496 , n44497 , n44498 , n44499 , n44500 , n44501 , n44502 , n44503 , n44504 , n44505 , n44506 , n44507 , n44508 , n44509 , n44510 , n44511 , n44512 , n44513 , n44514 , n44515 , n44516 , n44517 , n44518 , n44519 , n44520 , n44521 , n44522 , n44523 , n44524 , n44525 , n44526 , n44527 , n44528 , n44529 , n44530 , n44531 , n44532 , n44533 , n44534 , n44535 , n44536 , n44537 , n44538 , n44539 , n44540 , n44541 , n44542 , n44543 , n44544 , n44545 , n44546 , n44547 , n44548 , n44549 , n44550 , n44551 , n44552 , n44553 , n44554 , n44555 , n44556 , n44557 , n44558 , n44559 , n44560 , n44561 , n44562 , n44563 , n44564 , n44565 , n44566 , n44567 , n44568 , n44569 , n44570 , n44571 , n44572 , n44573 , n44574 , n44575 , n44576 , n44577 , n44578 , n44579 , n44580 , n44581 , n44582 , n44583 , n44584 , n44585 , n44586 , n44587 , n44588 , n44589 , n44590 , n44591 , n44592 , n44593 , n44594 , n44595 , n44596 , n44597 , n44598 , n44599 , n44600 , n44601 , n44602 , n44603 , n44604 , n44605 , n44606 , n44607 , n44608 , n44609 , n44610 , n44611 , n44612 , n44613 , n44614 , n44615 , n44616 , n44617 , n44618 , n44619 , n44620 , n44621 , n44622 , n44623 , n44624 , n44625 , n44626 , n44627 , n44628 , n44629 , n44630 , n44631 , n44632 , n44633 , n44634 , n44635 , n44636 , n44637 , n44638 , n44639 , n44640 , n44641 , n44642 , n44643 , n44644 , n44645 , n44646 , n44647 , n44648 , n44649 , n44650 , n44651 , n44652 , n44653 , n44654 , n44655 , n44656 , n44657 , n44658 , n44659 , n44660 , n44661 , n44662 , n44663 , n44664 , n44665 , n44666 , n44667 , n44668 , n44669 , n44670 , n44671 , n44672 , n44673 , n44674 , n44675 , n44676 , n44677 , n44678 , n44679 , n44680 , n44681 , n44682 , n44683 , n44684 , n44685 , n44686 , n44687 , n44688 , n44689 , n44690 , n44691 , n44692 , n44693 , n44694 , n44695 , n44696 , n44697 , n44698 , n44699 , n44700 , n44701 , n44702 , n44703 , n44704 , n44705 , n44706 , n44707 , n44708 , n44709 , n44710 , n44711 , n44712 , n44713 , n44714 , n44715 , n44716 , n44717 , n44718 , n44719 , n44720 , n44721 , n44722 , n44723 , n44724 , n44725 , n44726 , n44727 , n44728 , n44729 , n44730 , n44731 , n44732 , n44733 , n44734 , n44735 , n44736 , n44737 , n44738 , n44739 , n44740 , n44741 , n44742 , n44743 , n44744 , n44745 , n44746 , n44747 , n44748 , n44749 , n44750 , n44751 , n44752 , n44753 , n44754 , n44755 , n44756 , n44757 , n44758 , n44759 , n44760 , n44761 , n44762 , n44763 , n44764 , n44765 , n44766 , n44767 , n44768 , n44769 , n44770 , n44771 , n44772 , n44773 , n44774 , n44775 , n44776 , n44777 , n44778 , n44779 , n44780 , n44781 , n44782 , n44783 , n44784 , n44785 , n44786 , n44787 , n44788 , n44789 , n44790 , n44791 , n44792 , n44793 , n44794 , n44795 , n44796 , n44797 , n44798 , n44799 , n44800 , n44801 , n44802 , n44803 , n44804 , n44805 , n44806 , n44807 , n44808 , n44809 , n44810 , n44811 , n44812 , n44813 , n44814 , n44815 , n44816 , n44817 , n44818 , n44819 , n44820 , n44821 , n44822 , n44823 , n44824 , n44825 , n44826 , n44827 , n44828 , n44829 , n44830 , n44831 , n44832 , n44833 , n44834 , n44835 , n44836 , n44837 , n44838 , n44839 , n44840 , n44841 , n44842 , n44843 , n44844 , n44845 , n44846 , n44847 , n44848 , n44849 , n44850 , n44851 , n44852 , n44853 , n44854 , n44855 , n44856 , n44857 , n44858 , n44859 , n44860 , n44861 , n44862 , n44863 , n44864 , n44865 , n44866 , n44867 , n44868 , n44869 , n44870 , n44871 , n44872 , n44873 , n44874 , n44875 , n44876 , n44877 , n44878 , n44879 , n44880 , n44881 , n44882 , n44883 , n44884 , n44885 , n44886 , n44887 , n44888 , n44889 , n44890 , n44891 , n44892 , n44893 , n44894 , n44895 , n44896 , n44897 , n44898 , n44899 , n44900 , n44901 , n44902 , n44903 , n44904 , n44905 , n44906 , n44907 , n44908 , n44909 , n44910 , n44911 , n44912 , n44913 , n44914 , n44915 , n44916 , n44917 , n44918 , n44919 , n44920 , n44921 , n44922 , n44923 , n44924 , n44925 , n44926 , n44927 , n44928 , n44929 , n44930 , n44931 , n44932 , n44933 , n44934 , n44935 , n44936 , n44937 , n44938 , n44939 , n44940 , n44941 , n44942 , n44943 , n44944 , n44945 , n44946 , n44947 , n44948 , n44949 , n44950 , n44951 , n44952 , n44953 , n44954 , n44955 , n44956 , n44957 , n44958 , n44959 , n44960 , n44961 , n44962 , n44963 , n44964 , n44965 , n44966 , n44967 , n44968 , n44969 , n44970 , n44971 , n44972 , n44973 , n44974 , n44975 , n44976 , n44977 , n44978 , n44979 , n44980 , n44981 , n44982 , n44983 , n44984 , n44985 , n44986 , n44987 , n44988 , n44989 , n44990 , n44991 , n44992 , n44993 , n44994 , n44995 , n44996 , n44997 , n44998 , n44999 , n45000 , n45001 , n45002 , n45003 , n45004 , n45005 , n45006 , n45007 , n45008 , n45009 , n45010 , n45011 , n45012 , n45013 , n45014 , n45015 , n45016 , n45017 , n45018 , n45019 , n45020 , n45021 , n45022 , n45023 , n45024 , n45025 , n45026 , n45027 , n45028 , n45029 , n45030 , n45031 , n45032 , n45033 , n45034 , n45035 , n45036 , n45037 , n45038 , n45039 , n45040 , n45041 , n45042 , n45043 , n45044 , n45045 , n45046 , n45047 , n45048 , n45049 , n45050 , n45051 , n45052 , n45053 , n45054 , n45055 , n45056 , n45057 , n45058 , n45059 , n45060 , n45061 , n45062 , n45063 , n45064 , n45065 , n45066 , n45067 , n45068 , n45069 , n45070 , n45071 , n45072 , n45073 , n45074 , n45075 , n45076 , n45077 , n45078 , n45079 , n45080 , n45081 , n45082 , n45083 , n45084 , n45085 , n45086 , n45087 , n45088 , n45089 , n45090 , n45091 , n45092 , n45093 , n45094 , n45095 , n45096 , n45097 , n45098 , n45099 , n45100 , n45101 , n45102 , n45103 , n45104 , n45105 , n45106 , n45107 , n45108 , n45109 , n45110 , n45111 , n45112 , n45113 , n45114 , n45115 , n45116 , n45117 , n45118 , n45119 , n45120 , n45121 , n45122 , n45123 , n45124 , n45125 , n45126 , n45127 , n45128 , n45129 , n45130 , n45131 , n45132 , n45133 , n45134 , n45135 , n45136 , n45137 , n45138 , n45139 , n45140 , n45141 , n45142 , n45143 , n45144 , n45145 , n45146 , n45147 , n45148 , n45149 , n45150 , n45151 , n45152 , n45153 , n45154 , n45155 , n45156 , n45157 , n45158 , n45159 , n45160 , n45161 , n45162 , n45163 , n45164 , n45165 , n45166 , n45167 , n45168 , n45169 , n45170 , n45171 , n45172 , n45173 , n45174 , n45175 , n45176 , n45177 , n45178 , n45179 , n45180 , n45181 , n45182 , n45183 , n45184 , n45185 , n45186 , n45187 , n45188 , n45189 , n45190 , n45191 , n45192 , n45193 , n45194 , n45195 , n45196 , n45197 , n45198 , n45199 , n45200 , n45201 , n45202 , n45203 , n45204 , n45205 , n45206 , n45207 , n45208 , n45209 , n45210 , n45211 , n45212 , n45213 , n45214 , n45215 , n45216 , n45217 , n45218 , n45219 , n45220 , n45221 , n45222 , n45223 , n45224 , n45225 , n45226 , n45227 , n45228 , n45229 , n45230 , n45231 , n45232 , n45233 , n45234 , n45235 , n45236 , n45237 , n45238 , n45239 , n45240 , n45241 , n45242 , n45243 , n45244 , n45245 , n45246 , n45247 , n45248 , n45249 , n45250 , n45251 , n45252 , n45253 , n45254 , n45255 , n45256 , n45257 , n45258 , n45259 , n45260 , n45261 , n45262 , n45263 , n45264 , n45265 , n45266 , n45267 , n45268 , n45269 , n45270 , n45271 , n45272 , n45273 , n45274 , n45275 , n45276 , n45277 , n45278 , n45279 , n45280 , n45281 , n45282 , n45283 , n45284 , n45285 , n45286 , n45287 , n45288 , n45289 , n45290 , n45291 , n45292 , n45293 , n45294 , n45295 , n45296 , n45297 , n45298 , n45299 , n45300 , n45301 , n45302 , n45303 , n45304 , n45305 , n45306 , n45307 , n45308 , n45309 , n45310 , n45311 , n45312 , n45313 , n45314 , n45315 , n45316 , n45317 , n45318 , n45319 , n45320 , n45321 , n45322 , n45323 , n45324 , n45325 , n45326 , n45327 , n45328 , n45329 , n45330 , n45331 , n45332 , n45333 , n45334 , n45335 , n45336 , n45337 , n45338 , n45339 , n45340 , n45341 , n45342 , n45343 , n45344 , n45345 , n45346 , n45347 , n45348 , n45349 , n45350 , n45351 , n45352 , n45353 , n45354 , n45355 , n45356 , n45357 , n45358 , n45359 , n45360 , n45361 , n45362 , n45363 , n45364 , n45365 , n45366 , n45367 , n45368 , n45369 , n45370 , n45371 , n45372 , n45373 , n45374 , n45375 , n45376 , n45377 , n45378 , n45379 , n45380 , n45381 , n45382 , n45383 , n45384 , n45385 , n45386 , n45387 , n45388 , n45389 , n45390 , n45391 , n45392 , n45393 , n45394 , n45395 , n45396 , n45397 , n45398 , n45399 , n45400 , n45401 , n45402 , n45403 , n45404 , n45405 , n45406 , n45407 , n45408 , n45409 , n45410 , n45411 , n45412 , n45413 , n45414 , n45415 , n45416 , n45417 , n45418 , n45419 , n45420 , n45421 , n45422 , n45423 , n45424 , n45425 , n45426 , n45427 , n45428 , n45429 , n45430 , n45431 , n45432 , n45433 , n45434 , n45435 , n45436 , n45437 , n45438 , n45439 , n45440 , n45441 , n45442 , n45443 , n45444 , n45445 , n45446 , n45447 , n45448 , n45449 , n45450 , n45451 , n45452 , n45453 , n45454 , n45455 , n45456 , n45457 , n45458 , n45459 , n45460 , n45461 , n45462 , n45463 , n45464 , n45465 , n45466 , n45467 , n45468 , n45469 , n45470 , n45471 , n45472 , n45473 , n45474 , n45475 , n45476 , n45477 , n45478 , n45479 , n45480 , n45481 , n45482 , n45483 , n45484 , n45485 , n45486 , n45487 , n45488 , n45489 , n45490 , n45491 , n45492 , n45493 , n45494 , n45495 , n45496 , n45497 , n45498 , n45499 , n45500 , n45501 , n45502 , n45503 , n45504 , n45505 , n45506 , n45507 , n45508 , n45509 , n45510 , n45511 , n45512 , n45513 , n45514 , n45515 , n45516 , n45517 , n45518 , n45519 , n45520 , n45521 , n45522 , n45523 , n45524 , n45525 , n45526 , n45527 , n45528 , n45529 , n45530 , n45531 , n45532 , n45533 , n45534 , n45535 , n45536 , n45537 , n45538 , n45539 , n45540 , n45541 , n45542 , n45543 , n45544 , n45545 , n45546 , n45547 , n45548 , n45549 , n45550 , n45551 , n45552 , n45553 , n45554 , n45555 , n45556 , n45557 , n45558 , n45559 , n45560 , n45561 , n45562 , n45563 , n45564 , n45565 , n45566 , n45567 , n45568 , n45569 , n45570 , n45571 , n45572 , n45573 , n45574 , n45575 , n45576 , n45577 , n45578 , n45579 , n45580 , n45581 , n45582 , n45583 , n45584 , n45585 , n45586 , n45587 , n45588 , n45589 , n45590 , n45591 , n45592 , n45593 , n45594 , n45595 , n45596 , n45597 , n45598 , n45599 , n45600 , n45601 , n45602 , n45603 , n45604 , n45605 , n45606 , n45607 , n45608 , n45609 , n45610 , n45611 , n45612 , n45613 , n45614 , n45615 , n45616 , n45617 , n45618 , n45619 , n45620 , n45621 , n45622 , n45623 , n45624 , n45625 , n45626 , n45627 , n45628 , n45629 , n45630 , n45631 , n45632 , n45633 , n45634 , n45635 , n45636 , n45637 , n45638 , n45639 , n45640 , n45641 , n45642 , n45643 , n45644 , n45645 , n45646 , n45647 , n45648 , n45649 , n45650 , n45651 , n45652 , n45653 , n45654 , n45655 , n45656 , n45657 , n45658 , n45659 , n45660 , n45661 , n45662 , n45663 , n45664 , n45665 , n45666 , n45667 , n45668 , n45669 , n45670 , n45671 , n45672 , n45673 , n45674 , n45675 , n45676 , n45677 , n45678 , n45679 , n45680 , n45681 , n45682 , n45683 , n45684 , n45685 , n45686 , n45687 , n45688 , n45689 , n45690 , n45691 , n45692 , n45693 , n45694 , n45695 , n45696 , n45697 , n45698 , n45699 , n45700 , n45701 , n45702 , n45703 , n45704 , n45705 , n45706 , n45707 , n45708 , n45709 , n45710 , n45711 , n45712 , n45713 , n45714 , n45715 , n45716 , n45717 , n45718 , n45719 , n45720 , n45721 , n45722 , n45723 , n45724 , n45725 , n45726 , n45727 , n45728 , n45729 , n45730 , n45731 , n45732 , n45733 , n45734 , n45735 , n45736 , n45737 , n45738 , n45739 , n45740 , n45741 , n45742 , n45743 , n45744 , n45745 , n45746 , n45747 , n45748 , n45749 , n45750 , n45751 , n45752 , n45753 , n45754 , n45755 , n45756 , n45757 , n45758 , n45759 , n45760 , n45761 , n45762 , n45763 , n45764 , n45765 , n45766 , n45767 , n45768 , n45769 , n45770 , n45771 , n45772 , n45773 , n45774 , n45775 , n45776 , n45777 , n45778 , n45779 , n45780 , n45781 , n45782 , n45783 , n45784 , n45785 , n45786 , n45787 , n45788 , n45789 , n45790 , n45791 , n45792 , n45793 , n45794 , n45795 , n45796 , n45797 , n45798 , n45799 , n45800 , n45801 , n45802 , n45803 , n45804 , n45805 , n45806 , n45807 , n45808 , n45809 , n45810 , n45811 , n45812 , n45813 , n45814 , n45815 , n45816 , n45817 , n45818 , n45819 , n45820 , n45821 , n45822 , n45823 , n45824 , n45825 , n45826 , n45827 , n45828 , n45829 , n45830 , n45831 , n45832 , n45833 , n45834 , n45835 , n45836 , n45837 , n45838 , n45839 , n45840 , n45841 , n45842 , n45843 , n45844 , n45845 , n45846 , n45847 , n45848 , n45849 , n45850 , n45851 , n45852 , n45853 , n45854 , n45855 , n45856 , n45857 , n45858 , n45859 , n45860 , n45861 , n45862 , n45863 , n45864 , n45865 , n45866 , n45867 , n45868 , n45869 , n45870 , n45871 , n45872 , n45873 , n45874 , n45875 , n45876 , n45877 , n45878 , n45879 , n45880 , n45881 , n45882 , n45883 , n45884 , n45885 , n45886 , n45887 , n45888 , n45889 , n45890 , n45891 , n45892 , n45893 , n45894 , n45895 , n45896 , n45897 , n45898 , n45899 , n45900 , n45901 , n45902 , n45903 , n45904 , n45905 , n45906 , n45907 , n45908 , n45909 , n45910 , n45911 , n45912 , n45913 , n45914 , n45915 , n45916 , n45917 , n45918 , n45919 , n45920 , n45921 , n45922 , n45923 , n45924 , n45925 , n45926 , n45927 , n45928 , n45929 , n45930 , n45931 , n45932 , n45933 , n45934 , n45935 , n45936 , n45937 , n45938 , n45939 , n45940 , n45941 , n45942 , n45943 , n45944 , n45945 , n45946 , n45947 , n45948 , n45949 , n45950 , n45951 , n45952 , n45953 , n45954 , n45955 , n45956 , n45957 , n45958 , n45959 , n45960 , n45961 , n45962 , n45963 , n45964 , n45965 , n45966 , n45967 , n45968 , n45969 , n45970 , n45971 , n45972 , n45973 , n45974 , n45975 , n45976 , n45977 , n45978 , n45979 , n45980 , n45981 , n45982 , n45983 , n45984 , n45985 , n45986 , n45987 , n45988 , n45989 , n45990 , n45991 , n45992 , n45993 , n45994 , n45995 , n45996 , n45997 , n45998 , n45999 , n46000 , n46001 , n46002 , n46003 , n46004 , n46005 , n46006 , n46007 , n46008 , n46009 , n46010 , n46011 , n46012 , n46013 , n46014 , n46015 , n46016 , n46017 , n46018 , n46019 , n46020 , n46021 , n46022 , n46023 , n46024 , n46025 , n46026 , n46027 , n46028 , n46029 , n46030 , n46031 , n46032 , n46033 , n46034 , n46035 , n46036 , n46037 , n46038 , n46039 , n46040 , n46041 , n46042 , n46043 , n46044 , n46045 , n46046 , n46047 , n46048 , n46049 , n46050 , n46051 , n46052 , n46053 , n46054 , n46055 , n46056 , n46057 , n46058 , n46059 , n46060 , n46061 , n46062 , n46063 , n46064 , n46065 , n46066 , n46067 , n46068 , n46069 , n46070 , n46071 , n46072 , n46073 , n46074 , n46075 , n46076 , n46077 , n46078 , n46079 , n46080 , n46081 , n46082 , n46083 , n46084 , n46085 , n46086 , n46087 , n46088 , n46089 , n46090 , n46091 , n46092 , n46093 , n46094 , n46095 , n46096 , n46097 , n46098 , n46099 , n46100 , n46101 , n46102 , n46103 , n46104 , n46105 , n46106 , n46107 , n46108 , n46109 , n46110 , n46111 , n46112 , n46113 , n46114 , n46115 , n46116 , n46117 , n46118 , n46119 , n46120 , n46121 , n46122 , n46123 , n46124 , n46125 , n46126 , n46127 , n46128 , n46129 , n46130 , n46131 , n46132 , n46133 , n46134 , n46135 , n46136 , n46137 , n46138 , n46139 , n46140 , n46141 , n46142 , n46143 , n46144 , n46145 , n46146 , n46147 , n46148 , n46149 , n46150 , n46151 , n46152 , n46153 , n46154 , n46155 , n46156 , n46157 , n46158 , n46159 , n46160 , n46161 , n46162 , n46163 , n46164 , n46165 , n46166 , n46167 , n46168 , n46169 , n46170 , n46171 , n46172 , n46173 , n46174 , n46175 , n46176 , n46177 , n46178 , n46179 , n46180 , n46181 , n46182 , n46183 , n46184 , n46185 , n46186 , n46187 , n46188 , n46189 , n46190 , n46191 , n46192 , n46193 , n46194 , n46195 , n46196 , n46197 , n46198 , n46199 , n46200 , n46201 , n46202 , n46203 , n46204 , n46205 , n46206 , n46207 , n46208 , n46209 , n46210 , n46211 , n46212 , n46213 , n46214 , n46215 , n46216 , n46217 , n46218 , n46219 , n46220 , n46221 , n46222 , n46223 , n46224 , n46225 , n46226 , n46227 , n46228 , n46229 , n46230 , n46231 , n46232 , n46233 , n46234 , n46235 , n46236 , n46237 , n46238 , n46239 , n46240 , n46241 , n46242 , n46243 , n46244 , n46245 , n46246 , n46247 , n46248 , n46249 , n46250 , n46251 , n46252 , n46253 , n46254 , n46255 , n46256 , n46257 , n46258 , n46259 , n46260 , n46261 , n46262 , n46263 , n46264 , n46265 , n46266 , n46267 , n46268 , n46269 , n46270 , n46271 , n46272 , n46273 , n46274 , n46275 , n46276 , n46277 , n46278 , n46279 , n46280 , n46281 , n46282 , n46283 , n46284 , n46285 , n46286 , n46287 , n46288 , n46289 , n46290 , n46291 , n46292 , n46293 , n46294 , n46295 , n46296 , n46297 , n46298 , n46299 , n46300 , n46301 , n46302 , n46303 , n46304 , n46305 , n46306 , n46307 , n46308 , n46309 , n46310 , n46311 , n46312 , n46313 , n46314 , n46315 , n46316 , n46317 , n46318 , n46319 , n46320 , n46321 , n46322 , n46323 , n46324 , n46325 , n46326 , n46327 , n46328 , n46329 , n46330 , n46331 , n46332 , n46333 , n46334 , n46335 , n46336 , n46337 , n46338 , n46339 , n46340 , n46341 , n46342 , n46343 , n46344 , n46345 , n46346 , n46347 , n46348 , n46349 , n46350 , n46351 , n46352 , n46353 , n46354 , n46355 , n46356 , n46357 , n46358 , n46359 , n46360 , n46361 , n46362 , n46363 , n46364 , n46365 , n46366 , n46367 , n46368 , n46369 , n46370 , n46371 , n46372 , n46373 , n46374 , n46375 , n46376 , n46377 , n46378 , n46379 , n46380 , n46381 , n46382 , n46383 , n46384 , n46385 , n46386 , n46387 , n46388 , n46389 , n46390 , n46391 , n46392 , n46393 , n46394 , n46395 , n46396 , n46397 , n46398 , n46399 , n46400 , n46401 , n46402 , n46403 , n46404 , n46405 , n46406 , n46407 , n46408 , n46409 , n46410 , n46411 , n46412 , n46413 , n46414 , n46415 , n46416 , n46417 , n46418 , n46419 , n46420 , n46421 , n46422 , n46423 , n46424 , n46425 , n46426 , n46427 , n46428 , n46429 , n46430 , n46431 , n46432 , n46433 , n46434 , n46435 , n46436 , n46437 , n46438 , n46439 , n46440 , n46441 , n46442 , n46443 , n46444 , n46445 , n46446 , n46447 , n46448 , n46449 , n46450 , n46451 , n46452 , n46453 , n46454 , n46455 , n46456 , n46457 , n46458 , n46459 , n46460 , n46461 , n46462 , n46463 , n46464 , n46465 , n46466 , n46467 , n46468 , n46469 , n46470 , n46471 , n46472 , n46473 , n46474 , n46475 , n46476 , n46477 , n46478 , n46479 , n46480 , n46481 , n46482 , n46483 , n46484 , n46485 , n46486 , n46487 , n46488 , n46489 , n46490 , n46491 , n46492 , n46493 , n46494 , n46495 , n46496 , n46497 , n46498 , n46499 , n46500 , n46501 , n46502 , n46503 , n46504 , n46505 , n46506 , n46507 , n46508 , n46509 , n46510 , n46511 , n46512 , n46513 , n46514 , n46515 , n46516 , n46517 , n46518 , n46519 , n46520 , n46521 , n46522 , n46523 , n46524 , n46525 , n46526 , n46527 , n46528 , n46529 , n46530 , n46531 , n46532 , n46533 , n46534 , n46535 , n46536 , n46537 , n46538 , n46539 , n46540 , n46541 , n46542 , n46543 , n46544 , n46545 , n46546 , n46547 , n46548 , n46549 , n46550 , n46551 , n46552 , n46553 , n46554 , n46555 , n46556 , n46557 , n46558 , n46559 , n46560 , n46561 , n46562 , n46563 , n46564 , n46565 , n46566 , n46567 , n46568 , n46569 , n46570 , n46571 , n46572 , n46573 , n46574 , n46575 , n46576 , n46577 , n46578 , n46579 , n46580 , n46581 , n46582 , n46583 , n46584 , n46585 , n46586 , n46587 , n46588 , n46589 , n46590 , n46591 , n46592 , n46593 , n46594 , n46595 , n46596 , n46597 , n46598 , n46599 , n46600 , n46601 , n46602 , n46603 , n46604 , n46605 , n46606 , n46607 , n46608 , n46609 , n46610 , n46611 , n46612 , n46613 , n46614 , n46615 , n46616 , n46617 , n46618 , n46619 , n46620 , n46621 , n46622 , n46623 , n46624 , n46625 , n46626 , n46627 , n46628 , n46629 , n46630 , n46631 , n46632 , n46633 , n46634 , n46635 , n46636 , n46637 , n46638 , n46639 , n46640 , n46641 , n46642 , n46643 , n46644 , n46645 , n46646 , n46647 , n46648 , n46649 , n46650 , n46651 , n46652 , n46653 , n46654 , n46655 , n46656 , n46657 , n46658 , n46659 , n46660 , n46661 , n46662 , n46663 , n46664 , n46665 , n46666 , n46667 , n46668 , n46669 , n46670 , n46671 , n46672 , n46673 , n46674 , n46675 , n46676 , n46677 , n46678 , n46679 , n46680 , n46681 , n46682 , n46683 , n46684 , n46685 , n46686 , n46687 , n46688 , n46689 , n46690 , n46691 , n46692 , n46693 , n46694 , n46695 , n46696 , n46697 , n46698 , n46699 , n46700 , n46701 , n46702 , n46703 , n46704 , n46705 , n46706 , n46707 , n46708 , n46709 , n46710 , n46711 , n46712 , n46713 , n46714 , n46715 , n46716 , n46717 , n46718 , n46719 , n46720 , n46721 , n46722 , n46723 , n46724 , n46725 , n46726 , n46727 , n46728 , n46729 , n46730 , n46731 , n46732 , n46733 , n46734 , n46735 , n46736 , n46737 , n46738 , n46739 , n46740 , n46741 , n46742 , n46743 , n46744 , n46745 , n46746 , n46747 , n46748 , n46749 , n46750 , n46751 , n46752 , n46753 , n46754 , n46755 , n46756 , n46757 , n46758 , n46759 , n46760 , n46761 , n46762 , n46763 , n46764 , n46765 , n46766 , n46767 , n46768 , n46769 , n46770 , n46771 , n46772 , n46773 , n46774 , n46775 , n46776 , n46777 , n46778 , n46779 , n46780 , n46781 , n46782 , n46783 , n46784 , n46785 , n46786 , n46787 , n46788 , n46789 , n46790 , n46791 , n46792 , n46793 , n46794 , n46795 , n46796 , n46797 , n46798 , n46799 , n46800 , n46801 , n46802 , n46803 , n46804 , n46805 , n46806 , n46807 , n46808 , n46809 , n46810 , n46811 , n46812 , n46813 , n46814 , n46815 , n46816 , n46817 , n46818 , n46819 , n46820 , n46821 , n46822 , n46823 , n46824 , n46825 , n46826 , n46827 , n46828 , n46829 , n46830 , n46831 , n46832 , n46833 , n46834 , n46835 , n46836 , n46837 , n46838 , n46839 , n46840 , n46841 , n46842 , n46843 , n46844 , n46845 , n46846 , n46847 , n46848 , n46849 , n46850 , n46851 , n46852 , n46853 , n46854 , n46855 , n46856 , n46857 , n46858 , n46859 , n46860 , n46861 , n46862 , n46863 , n46864 , n46865 , n46866 , n46867 , n46868 , n46869 , n46870 , n46871 , n46872 , n46873 , n46874 , n46875 , n46876 , n46877 , n46878 , n46879 , n46880 , n46881 , n46882 , n46883 , n46884 , n46885 , n46886 , n46887 , n46888 , n46889 , n46890 , n46891 , n46892 , n46893 , n46894 , n46895 , n46896 , n46897 , n46898 , n46899 , n46900 , n46901 , n46902 , n46903 , n46904 , n46905 , n46906 , n46907 , n46908 , n46909 , n46910 , n46911 , n46912 , n46913 , n46914 , n46915 , n46916 , n46917 , n46918 , n46919 , n46920 , n46921 , n46922 , n46923 , n46924 , n46925 , n46926 , n46927 , n46928 , n46929 , n46930 , n46931 , n46932 , n46933 , n46934 , n46935 , n46936 , n46937 , n46938 , n46939 , n46940 , n46941 , n46942 , n46943 , n46944 , n46945 , n46946 , n46947 , n46948 , n46949 , n46950 , n46951 , n46952 , n46953 , n46954 , n46955 , n46956 , n46957 , n46958 , n46959 , n46960 , n46961 , n46962 , n46963 , n46964 , n46965 , n46966 , n46967 , n46968 , n46969 , n46970 , n46971 , n46972 , n46973 , n46974 , n46975 , n46976 , n46977 , n46978 , n46979 , n46980 , n46981 , n46982 , n46983 , n46984 , n46985 , n46986 , n46987 , n46988 , n46989 , n46990 , n46991 , n46992 , n46993 , n46994 , n46995 , n46996 , n46997 , n46998 , n46999 , n47000 , n47001 , n47002 , n47003 , n47004 , n47005 , n47006 , n47007 , n47008 , n47009 , n47010 , n47011 , n47012 , n47013 , n47014 , n47015 , n47016 , n47017 , n47018 , n47019 , n47020 , n47021 , n47022 , n47023 , n47024 , n47025 , n47026 , n47027 , n47028 , n47029 , n47030 , n47031 , n47032 , n47033 , n47034 , n47035 , n47036 , n47037 , n47038 , n47039 , n47040 , n47041 , n47042 , n47043 , n47044 , n47045 , n47046 , n47047 , n47048 , n47049 , n47050 , n47051 , n47052 , n47053 , n47054 , n47055 , n47056 , n47057 , n47058 , n47059 , n47060 , n47061 , n47062 , n47063 , n47064 , n47065 , n47066 , n47067 , n47068 , n47069 , n47070 , n47071 , n47072 , n47073 , n47074 , n47075 , n47076 , n47077 , n47078 , n47079 , n47080 , n47081 , n47082 , n47083 , n47084 , n47085 , n47086 , n47087 , n47088 , n47089 , n47090 , n47091 , n47092 , n47093 , n47094 , n47095 , n47096 , n47097 , n47098 , n47099 , n47100 , n47101 , n47102 , n47103 , n47104 , n47105 , n47106 , n47107 , n47108 , n47109 , n47110 , n47111 , n47112 , n47113 , n47114 , n47115 , n47116 , n47117 , n47118 , n47119 , n47120 , n47121 , n47122 , n47123 , n47124 , n47125 , n47126 , n47127 , n47128 , n47129 , n47130 , n47131 , n47132 , n47133 , n47134 , n47135 , n47136 , n47137 , n47138 , n47139 , n47140 , n47141 , n47142 , n47143 , n47144 , n47145 , n47146 , n47147 , n47148 , n47149 , n47150 , n47151 , n47152 , n47153 , n47154 , n47155 , n47156 , n47157 , n47158 , n47159 , n47160 , n47161 , n47162 , n47163 , n47164 , n47165 , n47166 , n47167 , n47168 , n47169 , n47170 , n47171 , n47172 , n47173 , n47174 , n47175 , n47176 , n47177 , n47178 , n47179 , n47180 , n47181 , n47182 , n47183 , n47184 , n47185 , n47186 , n47187 , n47188 , n47189 , n47190 , n47191 , n47192 , n47193 , n47194 , n47195 , n47196 , n47197 , n47198 , n47199 , n47200 , n47201 , n47202 , n47203 , n47204 , n47205 , n47206 , n47207 , n47208 , n47209 , n47210 , n47211 , n47212 , n47213 , n47214 , n47215 , n47216 , n47217 , n47218 , n47219 , n47220 , n47221 , n47222 , n47223 , n47224 , n47225 , n47226 , n47227 , n47228 , n47229 , n47230 , n47231 , n47232 , n47233 , n47234 , n47235 , n47236 , n47237 , n47238 , n47239 , n47240 , n47241 , n47242 , n47243 , n47244 , n47245 , n47246 , n47247 , n47248 , n47249 , n47250 , n47251 , n47252 , n47253 , n47254 , n47255 , n47256 , n47257 , n47258 , n47259 , n47260 , n47261 , n47262 , n47263 , n47264 , n47265 , n47266 , n47267 , n47268 , n47269 , n47270 , n47271 , n47272 , n47273 , n47274 , n47275 , n47276 , n47277 , n47278 , n47279 , n47280 , n47281 , n47282 , n47283 , n47284 , n47285 , n47286 , n47287 , n47288 , n47289 , n47290 , n47291 , n47292 , n47293 , n47294 , n47295 , n47296 , n47297 , n47298 , n47299 , n47300 , n47301 , n47302 , n47303 , n47304 , n47305 , n47306 , n47307 , n47308 , n47309 , n47310 , n47311 , n47312 , n47313 , n47314 , n47315 , n47316 , n47317 , n47318 , n47319 , n47320 , n47321 , n47322 , n47323 , n47324 , n47325 , n47326 , n47327 , n47328 , n47329 , n47330 , n47331 , n47332 , n47333 , n47334 , n47335 , n47336 , n47337 , n47338 , n47339 , n47340 , n47341 , n47342 , n47343 , n47344 , n47345 , n47346 , n47347 , n47348 , n47349 , n47350 , n47351 , n47352 , n47353 , n47354 , n47355 , n47356 , n47357 , n47358 , n47359 , n47360 , n47361 , n47362 , n47363 , n47364 , n47365 , n47366 , n47367 , n47368 , n47369 , n47370 , n47371 , n47372 , n47373 , n47374 , n47375 , n47376 , n47377 , n47378 , n47379 , n47380 , n47381 , n47382 , n47383 , n47384 , n47385 , n47386 , n47387 , n47388 , n47389 , n47390 , n47391 , n47392 , n47393 , n47394 , n47395 , n47396 , n47397 , n47398 , n47399 , n47400 , n47401 , n47402 , n47403 , n47404 , n47405 , n47406 , n47407 , n47408 , n47409 , n47410 , n47411 , n47412 , n47413 , n47414 , n47415 , n47416 , n47417 , n47418 , n47419 , n47420 , n47421 , n47422 , n47423 , n47424 , n47425 , n47426 , n47427 , n47428 , n47429 , n47430 , n47431 , n47432 , n47433 , n47434 , n47435 , n47436 , n47437 , n47438 , n47439 , n47440 , n47441 , n47442 , n47443 , n47444 , n47445 , n47446 , n47447 , n47448 , n47449 , n47450 , n47451 , n47452 , n47453 , n47454 , n47455 , n47456 , n47457 , n47458 , n47459 , n47460 , n47461 , n47462 , n47463 , n47464 , n47465 , n47466 , n47467 , n47468 , n47469 , n47470 , n47471 , n47472 , n47473 , n47474 , n47475 , n47476 , n47477 , n47478 , n47479 , n47480 , n47481 , n47482 , n47483 , n47484 , n47485 , n47486 , n47487 , n47488 , n47489 , n47490 , n47491 , n47492 , n47493 , n47494 , n47495 , n47496 , n47497 , n47498 , n47499 , n47500 , n47501 , n47502 , n47503 , n47504 , n47505 , n47506 , n47507 , n47508 , n47509 , n47510 , n47511 , n47512 , n47513 , n47514 , n47515 , n47516 , n47517 , n47518 , n47519 , n47520 , n47521 , n47522 , n47523 , n47524 , n47525 , n47526 , n47527 , n47528 , n47529 , n47530 , n47531 , n47532 , n47533 , n47534 , n47535 , n47536 , n47537 , n47538 , n47539 , n47540 , n47541 , n47542 , n47543 , n47544 , n47545 , n47546 , n47547 , n47548 , n47549 , n47550 , n47551 , n47552 , n47553 , n47554 , n47555 , n47556 , n47557 , n47558 , n47559 , n47560 , n47561 , n47562 , n47563 , n47564 , n47565 , n47566 , n47567 , n47568 , n47569 , n47570 , n47571 , n47572 , n47573 , n47574 , n47575 , n47576 , n47577 , n47578 , n47579 , n47580 , n47581 , n47582 , n47583 , n47584 , n47585 , n47586 , n47587 , n47588 , n47589 , n47590 , n47591 , n47592 , n47593 , n47594 , n47595 , n47596 , n47597 , n47598 , n47599 , n47600 , n47601 , n47602 , n47603 , n47604 , n47605 , n47606 , n47607 , n47608 , n47609 , n47610 , n47611 , n47612 , n47613 , n47614 , n47615 , n47616 , n47617 , n47618 , n47619 , n47620 , n47621 , n47622 , n47623 , n47624 , n47625 , n47626 , n47627 , n47628 , n47629 , n47630 , n47631 , n47632 , n47633 , n47634 , n47635 , n47636 , n47637 , n47638 , n47639 , n47640 , n47641 , n47642 , n47643 , n47644 , n47645 , n47646 , n47647 , n47648 , n47649 , n47650 , n47651 , n47652 , n47653 , n47654 , n47655 , n47656 , n47657 , n47658 , n47659 , n47660 , n47661 , n47662 , n47663 , n47664 , n47665 , n47666 , n47667 , n47668 , n47669 , n47670 , n47671 , n47672 , n47673 , n47674 , n47675 , n47676 , n47677 , n47678 , n47679 , n47680 , n47681 , n47682 , n47683 , n47684 , n47685 , n47686 , n47687 , n47688 , n47689 , n47690 , n47691 , n47692 , n47693 , n47694 , n47695 , n47696 , n47697 , n47698 , n47699 , n47700 , n47701 , n47702 , n47703 , n47704 , n47705 , n47706 , n47707 , n47708 , n47709 , n47710 , n47711 , n47712 , n47713 , n47714 , n47715 , n47716 , n47717 , n47718 , n47719 , n47720 , n47721 , n47722 , n47723 , n47724 , n47725 , n47726 , n47727 , n47728 , n47729 , n47730 , n47731 , n47732 , n47733 , n47734 , n47735 , n47736 , n47737 , n47738 , n47739 , n47740 , n47741 , n47742 , n47743 , n47744 , n47745 , n47746 , n47747 , n47748 , n47749 , n47750 , n47751 , n47752 , n47753 , n47754 , n47755 , n47756 , n47757 , n47758 , n47759 , n47760 , n47761 , n47762 , n47763 , n47764 , n47765 , n47766 , n47767 , n47768 , n47769 , n47770 , n47771 , n47772 , n47773 , n47774 , n47775 , n47776 , n47777 , n47778 , n47779 , n47780 , n47781 , n47782 , n47783 , n47784 , n47785 , n47786 , n47787 , n47788 , n47789 , n47790 , n47791 , n47792 , n47793 , n47794 , n47795 , n47796 , n47797 , n47798 , n47799 , n47800 , n47801 , n47802 , n47803 , n47804 , n47805 , n47806 , n47807 , n47808 , n47809 , n47810 , n47811 , n47812 , n47813 , n47814 , n47815 , n47816 , n47817 , n47818 , n47819 , n47820 , n47821 , n47822 , n47823 , n47824 , n47825 , n47826 , n47827 , n47828 , n47829 , n47830 , n47831 , n47832 , n47833 , n47834 , n47835 , n47836 , n47837 , n47838 , n47839 , n47840 , n47841 , n47842 , n47843 , n47844 , n47845 , n47846 , n47847 , n47848 , n47849 , n47850 , n47851 , n47852 , n47853 , n47854 , n47855 , n47856 , n47857 , n47858 , n47859 , n47860 , n47861 , n47862 , n47863 , n47864 , n47865 , n47866 , n47867 , n47868 , n47869 , n47870 , n47871 , n47872 , n47873 , n47874 , n47875 , n47876 , n47877 , n47878 , n47879 , n47880 , n47881 , n47882 , n47883 , n47884 , n47885 , n47886 , n47887 , n47888 , n47889 , n47890 , n47891 , n47892 , n47893 , n47894 , n47895 , n47896 , n47897 , n47898 , n47899 , n47900 , n47901 , n47902 , n47903 , n47904 , n47905 , n47906 , n47907 , n47908 , n47909 , n47910 , n47911 , n47912 , n47913 , n47914 , n47915 , n47916 , n47917 , n47918 , n47919 , n47920 , n47921 , n47922 , n47923 , n47924 , n47925 , n47926 , n47927 , n47928 , n47929 , n47930 , n47931 , n47932 , n47933 , n47934 , n47935 , n47936 , n47937 , n47938 , n47939 , n47940 , n47941 , n47942 , n47943 , n47944 , n47945 , n47946 , n47947 , n47948 , n47949 , n47950 , n47951 , n47952 , n47953 , n47954 , n47955 , n47956 , n47957 , n47958 , n47959 , n47960 , n47961 , n47962 , n47963 , n47964 , n47965 , n47966 , n47967 , n47968 , n47969 , n47970 , n47971 , n47972 , n47973 , n47974 , n47975 , n47976 , n47977 , n47978 , n47979 , n47980 , n47981 , n47982 , n47983 , n47984 , n47985 , n47986 , n47987 , n47988 , n47989 , n47990 , n47991 , n47992 , n47993 , n47994 , n47995 , n47996 , n47997 , n47998 , n47999 , n48000 , n48001 , n48002 , n48003 , n48004 , n48005 , n48006 , n48007 , n48008 , n48009 , n48010 , n48011 , n48012 , n48013 , n48014 , n48015 , n48016 , n48017 , n48018 , n48019 , n48020 , n48021 , n48022 , n48023 , n48024 , n48025 , n48026 , n48027 , n48028 , n48029 , n48030 , n48031 , n48032 , n48033 , n48034 , n48035 , n48036 , n48037 , n48038 , n48039 , n48040 , n48041 , n48042 , n48043 , n48044 , n48045 , n48046 , n48047 , n48048 , n48049 , n48050 , n48051 , n48052 , n48053 , n48054 , n48055 , n48056 , n48057 , n48058 , n48059 , n48060 , n48061 , n48062 , n48063 , n48064 , n48065 , n48066 , n48067 , n48068 , n48069 , n48070 , n48071 , n48072 , n48073 , n48074 , n48075 , n48076 , n48077 , n48078 , n48079 , n48080 , n48081 , n48082 , n48083 , n48084 , n48085 , n48086 , n48087 , n48088 , n48089 , n48090 , n48091 , n48092 , n48093 , n48094 , n48095 , n48096 , n48097 , n48098 , n48099 , n48100 , n48101 , n48102 , n48103 , n48104 , n48105 , n48106 , n48107 , n48108 , n48109 , n48110 , n48111 , n48112 , n48113 , n48114 , n48115 , n48116 , n48117 , n48118 , n48119 , n48120 , n48121 , n48122 , n48123 , n48124 , n48125 , n48126 , n48127 , n48128 , n48129 , n48130 , n48131 , n48132 , n48133 , n48134 , n48135 , n48136 , n48137 , n48138 , n48139 , n48140 , n48141 , n48142 , n48143 , n48144 , n48145 , n48146 , n48147 , n48148 , n48149 , n48150 , n48151 , n48152 , n48153 , n48154 , n48155 , n48156 , n48157 , n48158 , n48159 , n48160 , n48161 , n48162 , n48163 , n48164 , n48165 , n48166 , n48167 , n48168 , n48169 , n48170 , n48171 , n48172 , n48173 , n48174 , n48175 , n48176 , n48177 , n48178 , n48179 , n48180 , n48181 , n48182 , n48183 , n48184 , n48185 , n48186 , n48187 , n48188 , n48189 , n48190 , n48191 , n48192 , n48193 , n48194 , n48195 , n48196 , n48197 , n48198 , n48199 , n48200 , n48201 , n48202 , n48203 , n48204 , n48205 , n48206 , n48207 , n48208 , n48209 , n48210 , n48211 , n48212 , n48213 , n48214 , n48215 , n48216 , n48217 , n48218 , n48219 , n48220 , n48221 , n48222 , n48223 , n48224 , n48225 , n48226 , n48227 , n48228 , n48229 , n48230 , n48231 , n48232 , n48233 , n48234 , n48235 , n48236 , n48237 , n48238 , n48239 , n48240 , n48241 , n48242 , n48243 , n48244 , n48245 , n48246 , n48247 , n48248 , n48249 , n48250 , n48251 , n48252 , n48253 , n48254 , n48255 , n48256 , n48257 , n48258 , n48259 , n48260 , n48261 , n48262 , n48263 , n48264 , n48265 , n48266 , n48267 , n48268 , n48269 , n48270 , n48271 , n48272 , n48273 , n48274 , n48275 , n48276 , n48277 , n48278 , n48279 , n48280 , n48281 , n48282 , n48283 , n48284 , n48285 , n48286 , n48287 , n48288 , n48289 , n48290 , n48291 , n48292 , n48293 , n48294 , n48295 , n48296 , n48297 , n48298 , n48299 , n48300 , n48301 , n48302 , n48303 , n48304 , n48305 , n48306 , n48307 , n48308 , n48309 , n48310 , n48311 , n48312 , n48313 , n48314 , n48315 , n48316 , n48317 , n48318 , n48319 , n48320 , n48321 , n48322 , n48323 , n48324 , n48325 , n48326 , n48327 , n48328 , n48329 , n48330 , n48331 , n48332 , n48333 , n48334 , n48335 , n48336 , n48337 , n48338 , n48339 , n48340 , n48341 , n48342 , n48343 , n48344 , n48345 , n48346 , n48347 , n48348 , n48349 , n48350 , n48351 , n48352 , n48353 , n48354 , n48355 , n48356 , n48357 , n48358 , n48359 , n48360 , n48361 , n48362 , n48363 , n48364 , n48365 , n48366 , n48367 , n48368 , n48369 , n48370 , n48371 , n48372 , n48373 , n48374 , n48375 , n48376 , n48377 , n48378 , n48379 , n48380 , n48381 , n48382 , n48383 , n48384 , n48385 , n48386 , n48387 , n48388 , n48389 , n48390 , n48391 , n48392 , n48393 , n48394 , n48395 , n48396 , n48397 , n48398 , n48399 , n48400 , n48401 , n48402 , n48403 , n48404 , n48405 , n48406 , n48407 , n48408 , n48409 , n48410 , n48411 , n48412 , n48413 , n48414 , n48415 , n48416 , n48417 , n48418 , n48419 , n48420 , n48421 , n48422 , n48423 , n48424 , n48425 , n48426 , n48427 , n48428 , n48429 , n48430 , n48431 , n48432 , n48433 , n48434 , n48435 , n48436 , n48437 , n48438 , n48439 , n48440 , n48441 , n48442 , n48443 , n48444 , n48445 , n48446 , n48447 , n48448 , n48449 , n48450 , n48451 , n48452 , n48453 , n48454 , n48455 , n48456 , n48457 , n48458 , n48459 , n48460 , n48461 , n48462 , n48463 , n48464 , n48465 , n48466 , n48467 , n48468 , n48469 , n48470 , n48471 , n48472 , n48473 , n48474 , n48475 , n48476 , n48477 , n48478 , n48479 , n48480 , n48481 , n48482 , n48483 , n48484 , n48485 , n48486 , n48487 , n48488 , n48489 , n48490 , n48491 , n48492 , n48493 , n48494 , n48495 , n48496 , n48497 , n48498 , n48499 , n48500 , n48501 , n48502 , n48503 , n48504 , n48505 , n48506 , n48507 , n48508 , n48509 , n48510 , n48511 , n48512 , n48513 , n48514 , n48515 , n48516 , n48517 , n48518 , n48519 , n48520 , n48521 , n48522 , n48523 , n48524 , n48525 , n48526 , n48527 , n48528 , n48529 , n48530 , n48531 , n48532 , n48533 , n48534 , n48535 , n48536 , n48537 , n48538 , n48539 , n48540 , n48541 , n48542 , n48543 , n48544 , n48545 , n48546 , n48547 , n48548 , n48549 , n48550 , n48551 , n48552 , n48553 , n48554 , n48555 , n48556 , n48557 , n48558 , n48559 , n48560 , n48561 , n48562 , n48563 , n48564 , n48565 , n48566 , n48567 , n48568 , n48569 , n48570 , n48571 , n48572 , n48573 , n48574 , n48575 , n48576 , n48577 , n48578 , n48579 , n48580 , n48581 , n48582 , n48583 , n48584 , n48585 , n48586 , n48587 , n48588 , n48589 , n48590 , n48591 , n48592 , n48593 , n48594 , n48595 , n48596 , n48597 , n48598 , n48599 , n48600 , n48601 , n48602 , n48603 , n48604 , n48605 , n48606 , n48607 , n48608 , n48609 , n48610 , n48611 , n48612 , n48613 , n48614 , n48615 , n48616 , n48617 , n48618 , n48619 , n48620 , n48621 , n48622 , n48623 , n48624 , n48625 , n48626 , n48627 , n48628 , n48629 , n48630 , n48631 , n48632 , n48633 , n48634 , n48635 , n48636 , n48637 , n48638 , n48639 , n48640 , n48641 , n48642 , n48643 , n48644 , n48645 , n48646 , n48647 , n48648 , n48649 , n48650 , n48651 , n48652 , n48653 , n48654 , n48655 , n48656 , n48657 , n48658 , n48659 , n48660 , n48661 , n48662 , n48663 , n48664 , n48665 , n48666 , n48667 , n48668 , n48669 , n48670 , n48671 , n48672 , n48673 , n48674 , n48675 , n48676 , n48677 , n48678 , n48679 , n48680 , n48681 , n48682 , n48683 , n48684 , n48685 , n48686 , n48687 , n48688 , n48689 , n48690 , n48691 , n48692 , n48693 , n48694 , n48695 , n48696 , n48697 , n48698 , n48699 , n48700 , n48701 , n48702 , n48703 , n48704 , n48705 , n48706 , n48707 , n48708 , n48709 , n48710 , n48711 , n48712 , n48713 , n48714 , n48715 , n48716 , n48717 , n48718 , n48719 , n48720 , n48721 , n48722 , n48723 , n48724 , n48725 , n48726 , n48727 , n48728 , n48729 , n48730 , n48731 , n48732 , n48733 , n48734 , n48735 , n48736 , n48737 , n48738 , n48739 , n48740 , n48741 , n48742 , n48743 , n48744 , n48745 , n48746 , n48747 , n48748 , n48749 , n48750 , n48751 , n48752 , n48753 , n48754 , n48755 , n48756 , n48757 , n48758 , n48759 , n48760 , n48761 , n48762 , n48763 , n48764 , n48765 , n48766 , n48767 , n48768 , n48769 , n48770 , n48771 , n48772 , n48773 , n48774 , n48775 , n48776 , n48777 , n48778 , n48779 , n48780 , n48781 , n48782 , n48783 , n48784 , n48785 , n48786 , n48787 , n48788 , n48789 , n48790 , n48791 , n48792 , n48793 , n48794 , n48795 , n48796 , n48797 , n48798 , n48799 , n48800 , n48801 , n48802 , n48803 , n48804 , n48805 , n48806 , n48807 , n48808 , n48809 , n48810 , n48811 , n48812 , n48813 , n48814 , n48815 , n48816 , n48817 , n48818 , n48819 , n48820 , n48821 , n48822 , n48823 , n48824 , n48825 , n48826 , n48827 , n48828 , n48829 , n48830 , n48831 , n48832 , n48833 , n48834 , n48835 , n48836 , n48837 , n48838 , n48839 , n48840 , n48841 , n48842 , n48843 , n48844 , n48845 , n48846 , n48847 , n48848 , n48849 , n48850 , n48851 , n48852 , n48853 , n48854 , n48855 , n48856 , n48857 , n48858 , n48859 , n48860 , n48861 , n48862 , n48863 , n48864 , n48865 , n48866 , n48867 , n48868 , n48869 , n48870 , n48871 , n48872 , n48873 , n48874 , n48875 , n48876 , n48877 , n48878 , n48879 , n48880 , n48881 , n48882 , n48883 , n48884 , n48885 , n48886 , n48887 , n48888 , n48889 , n48890 , n48891 , n48892 , n48893 , n48894 , n48895 , n48896 , n48897 , n48898 , n48899 , n48900 , n48901 , n48902 , n48903 , n48904 , n48905 , n48906 , n48907 , n48908 , n48909 , n48910 , n48911 , n48912 , n48913 , n48914 , n48915 , n48916 , n48917 , n48918 , n48919 , n48920 , n48921 , n48922 , n48923 , n48924 , n48925 , n48926 , n48927 , n48928 , n48929 , n48930 , n48931 , n48932 , n48933 , n48934 , n48935 , n48936 , n48937 , n48938 , n48939 , n48940 , n48941 , n48942 , n48943 , n48944 , n48945 , n48946 , n48947 , n48948 , n48949 , n48950 , n48951 , n48952 , n48953 , n48954 , n48955 , n48956 , n48957 , n48958 , n48959 , n48960 , n48961 , n48962 , n48963 , n48964 , n48965 , n48966 , n48967 , n48968 , n48969 , n48970 , n48971 , n48972 , n48973 , n48974 , n48975 , n48976 , n48977 , n48978 , n48979 , n48980 , n48981 , n48982 , n48983 , n48984 , n48985 , n48986 , n48987 , n48988 , n48989 , n48990 , n48991 , n48992 , n48993 , n48994 , n48995 , n48996 , n48997 , n48998 , n48999 , n49000 , n49001 , n49002 , n49003 , n49004 , n49005 , n49006 , n49007 , n49008 , n49009 , n49010 , n49011 , n49012 , n49013 , n49014 , n49015 , n49016 , n49017 , n49018 , n49019 , n49020 , n49021 , n49022 , n49023 , n49024 , n49025 , n49026 , n49027 , n49028 , n49029 , n49030 , n49031 , n49032 , n49033 , n49034 , n49035 , n49036 , n49037 , n49038 , n49039 , n49040 , n49041 , n49042 , n49043 , n49044 , n49045 , n49046 , n49047 , n49048 , n49049 , n49050 , n49051 , n49052 , n49053 , n49054 , n49055 , n49056 , n49057 , n49058 , n49059 , n49060 , n49061 , n49062 , n49063 , n49064 , n49065 , n49066 , n49067 , n49068 , n49069 , n49070 , n49071 , n49072 , n49073 , n49074 , n49075 , n49076 , n49077 , n49078 , n49079 , n49080 , n49081 , n49082 , n49083 , n49084 , n49085 , n49086 , n49087 , n49088 , n49089 , n49090 , n49091 , n49092 , n49093 , n49094 , n49095 , n49096 , n49097 , n49098 , n49099 , n49100 , n49101 , n49102 , n49103 , n49104 , n49105 , n49106 , n49107 , n49108 , n49109 , n49110 , n49111 , n49112 , n49113 , n49114 , n49115 , n49116 , n49117 , n49118 , n49119 , n49120 , n49121 , n49122 , n49123 , n49124 , n49125 , n49126 , n49127 , n49128 , n49129 , n49130 , n49131 , n49132 , n49133 , n49134 , n49135 , n49136 , n49137 , n49138 , n49139 , n49140 , n49141 , n49142 , n49143 , n49144 , n49145 , n49146 , n49147 , n49148 , n49149 , n49150 , n49151 , n49152 , n49153 , n49154 , n49155 , n49156 , n49157 , n49158 , n49159 , n49160 , n49161 , n49162 , n49163 , n49164 , n49165 , n49166 , n49167 , n49168 , n49169 , n49170 , n49171 , n49172 , n49173 , n49174 , n49175 , n49176 , n49177 , n49178 , n49179 , n49180 , n49181 , n49182 , n49183 , n49184 , n49185 , n49186 , n49187 , n49188 , n49189 , n49190 , n49191 , n49192 , n49193 , n49194 , n49195 , n49196 , n49197 , n49198 , n49199 , n49200 , n49201 , n49202 , n49203 , n49204 , n49205 , n49206 , n49207 , n49208 , n49209 , n49210 , n49211 , n49212 , n49213 , n49214 , n49215 , n49216 , n49217 , n49218 , n49219 , n49220 , n49221 , n49222 , n49223 , n49224 , n49225 , n49226 , n49227 , n49228 , n49229 , n49230 , n49231 , n49232 , n49233 , n49234 , n49235 , n49236 , n49237 , n49238 , n49239 , n49240 , n49241 , n49242 , n49243 , n49244 , n49245 , n49246 , n49247 , n49248 , n49249 , n49250 , n49251 , n49252 , n49253 , n49254 , n49255 , n49256 , n49257 , n49258 , n49259 , n49260 , n49261 , n49262 , n49263 , n49264 , n49265 , n49266 , n49267 , n49268 , n49269 , n49270 , n49271 , n49272 , n49273 , n49274 , n49275 , n49276 , n49277 , n49278 , n49279 , n49280 , n49281 , n49282 , n49283 , n49284 , n49285 , n49286 , n49287 , n49288 , n49289 , n49290 , n49291 , n49292 , n49293 , n49294 , n49295 , n49296 , n49297 , n49298 , n49299 , n49300 , n49301 , n49302 , n49303 , n49304 , n49305 , n49306 , n49307 , n49308 , n49309 , n49310 , n49311 , n49312 , n49313 , n49314 , n49315 , n49316 , n49317 , n49318 , n49319 , n49320 , n49321 , n49322 , n49323 , n49324 , n49325 , n49326 , n49327 , n49328 , n49329 , n49330 , n49331 , n49332 , n49333 , n49334 , n49335 , n49336 , n49337 , n49338 , n49339 , n49340 , n49341 , n49342 , n49343 , n49344 , n49345 , n49346 , n49347 , n49348 , n49349 , n49350 , n49351 , n49352 , n49353 , n49354 , n49355 , n49356 , n49357 , n49358 , n49359 , n49360 , n49361 , n49362 , n49363 , n49364 , n49365 , n49366 , n49367 , n49368 , n49369 , n49370 , n49371 , n49372 , n49373 , n49374 , n49375 , n49376 , n49377 , n49378 , n49379 , n49380 , n49381 , n49382 , n49383 , n49384 , n49385 , n49386 , n49387 , n49388 , n49389 , n49390 , n49391 , n49392 , n49393 , n49394 , n49395 , n49396 , n49397 , n49398 , n49399 , n49400 , n49401 , n49402 , n49403 , n49404 , n49405 , n49406 , n49407 , n49408 , n49409 , n49410 , n49411 , n49412 , n49413 , n49414 , n49415 , n49416 , n49417 , n49418 , n49419 , n49420 , n49421 , n49422 , n49423 , n49424 , n49425 , n49426 , n49427 , n49428 , n49429 , n49430 , n49431 , n49432 , n49433 , n49434 , n49435 , n49436 , n49437 , n49438 , n49439 , n49440 , n49441 , n49442 , n49443 , n49444 , n49445 , n49446 , n49447 , n49448 , n49449 , n49450 , n49451 , n49452 , n49453 , n49454 , n49455 , n49456 , n49457 , n49458 , n49459 , n49460 , n49461 , n49462 , n49463 , n49464 , n49465 , n49466 , n49467 , n49468 , n49469 , n49470 , n49471 , n49472 , n49473 , n49474 , n49475 , n49476 , n49477 , n49478 , n49479 , n49480 , n49481 , n49482 , n49483 , n49484 , n49485 , n49486 , n49487 , n49488 , n49489 , n49490 , n49491 , n49492 , n49493 , n49494 , n49495 , n49496 , n49497 , n49498 , n49499 , n49500 , n49501 , n49502 , n49503 , n49504 , n49505 , n49506 , n49507 , n49508 , n49509 , n49510 , n49511 , n49512 , n49513 , n49514 , n49515 , n49516 , n49517 , n49518 , n49519 , n49520 , n49521 , n49522 , n49523 , n49524 , n49525 , n49526 , n49527 , n49528 , n49529 , n49530 , n49531 , n49532 , n49533 , n49534 , n49535 , n49536 , n49537 , n49538 , n49539 , n49540 , n49541 , n49542 , n49543 , n49544 , n49545 , n49546 , n49547 , n49548 , n49549 , n49550 , n49551 , n49552 , n49553 , n49554 , n49555 , n49556 , n49557 , n49558 , n49559 , n49560 , n49561 , n49562 , n49563 , n49564 , n49565 , n49566 , n49567 , n49568 , n49569 , n49570 , n49571 , n49572 , n49573 , n49574 , n49575 , n49576 , n49577 , n49578 , n49579 , n49580 , n49581 , n49582 , n49583 , n49584 , n49585 , n49586 , n49587 , n49588 , n49589 , n49590 , n49591 , n49592 , n49593 , n49594 , n49595 , n49596 , n49597 , n49598 , n49599 , n49600 , n49601 , n49602 , n49603 , n49604 , n49605 , n49606 , n49607 , n49608 , n49609 , n49610 , n49611 , n49612 , n49613 , n49614 , n49615 , n49616 , n49617 , n49618 , n49619 , n49620 , n49621 , n49622 , n49623 , n49624 , n49625 , n49626 , n49627 , n49628 , n49629 , n49630 , n49631 , n49632 , n49633 , n49634 , n49635 , n49636 , n49637 , n49638 , n49639 , n49640 , n49641 , n49642 , n49643 , n49644 , n49645 , n49646 , n49647 , n49648 , n49649 , n49650 , n49651 , n49652 , n49653 , n49654 , n49655 , n49656 , n49657 , n49658 , n49659 , n49660 , n49661 , n49662 , n49663 , n49664 , n49665 , n49666 , n49667 , n49668 , n49669 , n49670 , n49671 , n49672 , n49673 , n49674 , n49675 , n49676 , n49677 , n49678 , n49679 , n49680 , n49681 , n49682 , n49683 , n49684 , n49685 , n49686 , n49687 , n49688 , n49689 , n49690 , n49691 , n49692 , n49693 , n49694 , n49695 , n49696 , n49697 , n49698 , n49699 , n49700 , n49701 , n49702 , n49703 , n49704 , n49705 , n49706 , n49707 , n49708 , n49709 , n49710 , n49711 , n49712 , n49713 , n49714 , n49715 , n49716 , n49717 , n49718 , n49719 , n49720 , n49721 , n49722 , n49723 , n49724 , n49725 , n49726 , n49727 , n49728 , n49729 , n49730 , n49731 , n49732 , n49733 , n49734 , n49735 , n49736 , n49737 , n49738 , n49739 , n49740 , n49741 , n49742 , n49743 , n49744 , n49745 , n49746 , n49747 , n49748 , n49749 , n49750 , n49751 , n49752 , n49753 , n49754 , n49755 , n49756 , n49757 , n49758 , n49759 , n49760 , n49761 , n49762 , n49763 , n49764 , n49765 , n49766 , n49767 , n49768 , n49769 , n49770 , n49771 , n49772 , n49773 , n49774 , n49775 , n49776 , n49777 , n49778 , n49779 , n49780 , n49781 , n49782 , n49783 , n49784 , n49785 , n49786 , n49787 , n49788 , n49789 , n49790 , n49791 , n49792 , n49793 , n49794 , n49795 , n49796 , n49797 , n49798 , n49799 , n49800 , n49801 , n49802 , n49803 , n49804 , n49805 , n49806 , n49807 , n49808 , n49809 , n49810 , n49811 , n49812 , n49813 , n49814 , n49815 , n49816 , n49817 , n49818 , n49819 , n49820 , n49821 , n49822 , n49823 , n49824 , n49825 , n49826 , n49827 , n49828 , n49829 , n49830 , n49831 , n49832 , n49833 , n49834 , n49835 , n49836 , n49837 , n49838 , n49839 , n49840 , n49841 , n49842 , n49843 , n49844 , n49845 , n49846 , n49847 , n49848 , n49849 , n49850 , n49851 , n49852 , n49853 , n49854 , n49855 , n49856 , n49857 , n49858 , n49859 , n49860 , n49861 , n49862 , n49863 , n49864 , n49865 , n49866 , n49867 , n49868 , n49869 , n49870 , n49871 , n49872 , n49873 , n49874 , n49875 , n49876 , n49877 , n49878 , n49879 , n49880 , n49881 , n49882 , n49883 , n49884 , n49885 , n49886 , n49887 , n49888 , n49889 , n49890 , n49891 , n49892 , n49893 , n49894 , n49895 , n49896 , n49897 , n49898 , n49899 , n49900 , n49901 , n49902 , n49903 , n49904 , n49905 , n49906 , n49907 , n49908 , n49909 , n49910 , n49911 , n49912 , n49913 , n49914 , n49915 , n49916 , n49917 , n49918 , n49919 , n49920 , n49921 , n49922 , n49923 , n49924 , n49925 , n49926 , n49927 , n49928 , n49929 , n49930 , n49931 , n49932 , n49933 , n49934 , n49935 , n49936 , n49937 , n49938 , n49939 , n49940 , n49941 , n49942 , n49943 , n49944 , n49945 , n49946 , n49947 , n49948 , n49949 , n49950 , n49951 , n49952 , n49953 , n49954 , n49955 , n49956 , n49957 , n49958 , n49959 , n49960 , n49961 , n49962 , n49963 , n49964 , n49965 , n49966 , n49967 , n49968 , n49969 , n49970 , n49971 , n49972 , n49973 , n49974 , n49975 , n49976 , n49977 , n49978 , n49979 , n49980 , n49981 , n49982 , n49983 , n49984 , n49985 , n49986 , n49987 , n49988 , n49989 , n49990 , n49991 , n49992 , n49993 , n49994 , n49995 , n49996 , n49997 , n49998 , n49999 , n50000 , n50001 , n50002 , n50003 , n50004 , n50005 , n50006 , n50007 , n50008 , n50009 , n50010 , n50011 , n50012 , n50013 , n50014 , n50015 , n50016 , n50017 , n50018 , n50019 , n50020 , n50021 , n50022 , n50023 , n50024 , n50025 , n50026 , n50027 , n50028 , n50029 , n50030 , n50031 , n50032 , n50033 , n50034 , n50035 , n50036 , n50037 , n50038 , n50039 , n50040 , n50041 , n50042 , n50043 , n50044 , n50045 , n50046 , n50047 , n50048 , n50049 , n50050 , n50051 , n50052 , n50053 , n50054 , n50055 , n50056 , n50057 , n50058 , n50059 , n50060 , n50061 , n50062 , n50063 , n50064 , n50065 , n50066 , n50067 , n50068 , n50069 , n50070 , n50071 , n50072 , n50073 , n50074 , n50075 , n50076 , n50077 , n50078 , n50079 , n50080 , n50081 , n50082 , n50083 , n50084 , n50085 , n50086 , n50087 , n50088 , n50089 , n50090 , n50091 , n50092 , n50093 , n50094 , n50095 , n50096 , n50097 , n50098 , n50099 , n50100 , n50101 , n50102 , n50103 , n50104 , n50105 , n50106 , n50107 , n50108 , n50109 , n50110 , n50111 , n50112 , n50113 , n50114 , n50115 , n50116 , n50117 , n50118 , n50119 , n50120 , n50121 , n50122 , n50123 , n50124 , n50125 , n50126 , n50127 , n50128 , n50129 , n50130 , n50131 , n50132 , n50133 , n50134 , n50135 , n50136 , n50137 , n50138 , n50139 , n50140 , n50141 , n50142 , n50143 , n50144 , n50145 , n50146 , n50147 , n50148 , n50149 , n50150 , n50151 , n50152 , n50153 , n50154 , n50155 , n50156 , n50157 , n50158 , n50159 , n50160 , n50161 , n50162 , n50163 , n50164 , n50165 , n50166 , n50167 , n50168 , n50169 , n50170 , n50171 , n50172 , n50173 , n50174 , n50175 , n50176 , n50177 , n50178 , n50179 , n50180 , n50181 , n50182 , n50183 , n50184 , n50185 , n50186 , n50187 , n50188 , n50189 , n50190 , n50191 , n50192 , n50193 , n50194 , n50195 , n50196 , n50197 , n50198 , n50199 , n50200 , n50201 , n50202 , n50203 , n50204 , n50205 , n50206 , n50207 , n50208 , n50209 , n50210 , n50211 , n50212 , n50213 , n50214 , n50215 , n50216 , n50217 , n50218 , n50219 , n50220 , n50221 , n50222 , n50223 , n50224 , n50225 , n50226 , n50227 , n50228 , n50229 , n50230 , n50231 , n50232 , n50233 , n50234 , n50235 , n50236 , n50237 , n50238 , n50239 , n50240 , n50241 , n50242 , n50243 , n50244 , n50245 , n50246 , n50247 , n50248 , n50249 , n50250 , n50251 , n50252 , n50253 , n50254 , n50255 , n50256 , n50257 , n50258 , n50259 , n50260 , n50261 , n50262 , n50263 , n50264 , n50265 , n50266 , n50267 , n50268 , n50269 , n50270 , n50271 , n50272 , n50273 , n50274 , n50275 , n50276 , n50277 , n50278 , n50279 , n50280 , n50281 , n50282 , n50283 , n50284 , n50285 , n50286 , n50287 , n50288 , n50289 , n50290 , n50291 , n50292 , n50293 , n50294 , n50295 , n50296 , n50297 , n50298 , n50299 , n50300 , n50301 , n50302 , n50303 , n50304 , n50305 , n50306 , n50307 , n50308 , n50309 , n50310 , n50311 , n50312 , n50313 , n50314 , n50315 , n50316 , n50317 , n50318 , n50319 , n50320 , n50321 , n50322 , n50323 , n50324 , n50325 , n50326 , n50327 , n50328 , n50329 , n50330 , n50331 , n50332 , n50333 , n50334 , n50335 , n50336 , n50337 , n50338 , n50339 , n50340 , n50341 , n50342 , n50343 , n50344 , n50345 , n50346 , n50347 , n50348 , n50349 , n50350 , n50351 , n50352 , n50353 , n50354 , n50355 , n50356 , n50357 , n50358 , n50359 , n50360 , n50361 , n50362 , n50363 , n50364 , n50365 , n50366 , n50367 , n50368 , n50369 , n50370 , n50371 , n50372 , n50373 , n50374 , n50375 , n50376 , n50377 , n50378 , n50379 , n50380 , n50381 , n50382 , n50383 , n50384 , n50385 , n50386 , n50387 , n50388 , n50389 , n50390 , n50391 , n50392 , n50393 , n50394 , n50395 , n50396 , n50397 , n50398 , n50399 , n50400 , n50401 , n50402 , n50403 , n50404 , n50405 , n50406 , n50407 , n50408 , n50409 , n50410 , n50411 , n50412 , n50413 , n50414 , n50415 , n50416 , n50417 , n50418 , n50419 , n50420 , n50421 , n50422 , n50423 , n50424 , n50425 , n50426 , n50427 , n50428 , n50429 , n50430 , n50431 , n50432 , n50433 , n50434 , n50435 , n50436 , n50437 , n50438 , n50439 , n50440 , n50441 , n50442 , n50443 , n50444 , n50445 , n50446 , n50447 , n50448 , n50449 , n50450 , n50451 , n50452 , n50453 , n50454 , n50455 , n50456 , n50457 , n50458 , n50459 , n50460 , n50461 , n50462 , n50463 , n50464 , n50465 , n50466 , n50467 , n50468 , n50469 , n50470 , n50471 , n50472 , n50473 , n50474 , n50475 , n50476 , n50477 , n50478 , n50479 , n50480 , n50481 , n50482 , n50483 , n50484 , n50485 , n50486 , n50487 , n50488 , n50489 , n50490 , n50491 , n50492 , n50493 , n50494 , n50495 , n50496 , n50497 , n50498 , n50499 , n50500 , n50501 , n50502 , n50503 ;
  assign n13 = x11 ^ x7 ^ x4 ;
  assign n14 = x3 & ~n13 ;
  assign n15 = ~x7 & n14 ;
  assign n16 = x4 & x6 ;
  assign n17 = n16 ^ x0 ^ 1'b0 ;
  assign n18 = x3 & x4 ;
  assign n19 = ~x0 & n18 ;
  assign n20 = x0 & x11 ;
  assign n21 = n20 ^ x8 ^ 1'b0 ;
  assign n28 = ( ~x6 & x7 ) | ( ~x6 & x8 ) | ( x7 & x8 ) ;
  assign n22 = x2 ^ x0 ^ 1'b0 ;
  assign n23 = x5 & n22 ;
  assign n29 = n23 ^ x11 ^ 1'b0 ;
  assign n30 = n28 & n29 ;
  assign n26 = n20 ^ x0 ^ 1'b0 ;
  assign n24 = ~n13 & n23 ;
  assign n25 = n24 ^ n19 ^ 1'b0 ;
  assign n27 = n26 ^ n25 ^ x1 ;
  assign n31 = n30 ^ n27 ^ 1'b0 ;
  assign n32 = ~n26 & n27 ;
  assign n33 = n32 ^ n30 ^ 1'b0 ;
  assign n34 = x10 & ~n33 ;
  assign n35 = ~x5 & n34 ;
  assign n36 = n23 | n31 ;
  assign n37 = x0 & ~n33 ;
  assign n38 = n37 ^ n31 ^ 1'b0 ;
  assign n46 = n23 & ~n26 ;
  assign n47 = n21 & n46 ;
  assign n42 = n30 ^ n19 ^ 1'b0 ;
  assign n43 = n28 & ~n42 ;
  assign n44 = ( x9 & n28 ) | ( x9 & ~n43 ) | ( n28 & ~n43 ) ;
  assign n39 = x5 & x6 ;
  assign n40 = n26 & n39 ;
  assign n41 = x7 & ~n40 ;
  assign n45 = n44 ^ n41 ^ 1'b0 ;
  assign n48 = n47 ^ n45 ^ x3 ;
  assign n49 = n48 ^ n47 ^ n17 ;
  assign n50 = x9 ^ x6 ^ 1'b0 ;
  assign n51 = ~n19 & n50 ;
  assign n52 = n25 ^ x7 ^ x6 ;
  assign n53 = x8 ^ x2 ^ 1'b0 ;
  assign n54 = ~n15 & n53 ;
  assign n55 = ~n52 & n54 ;
  assign n56 = n31 & n55 ;
  assign n57 = n56 ^ x3 ^ x2 ;
  assign n58 = n57 ^ n56 ^ x11 ;
  assign n59 = ~n17 & n43 ;
  assign n60 = n59 ^ x10 ^ 1'b0 ;
  assign n61 = n30 & ~n60 ;
  assign n62 = n61 ^ x1 ^ 1'b0 ;
  assign n63 = ~n48 & n62 ;
  assign n64 = n31 | n52 ;
  assign n65 = n64 ^ n33 ^ 1'b0 ;
  assign n66 = n60 ^ x8 ^ 1'b0 ;
  assign n67 = n65 | n66 ;
  assign n68 = n54 & ~n67 ;
  assign n69 = ~n63 & n68 ;
  assign n70 = n30 & ~n65 ;
  assign n71 = n13 & n70 ;
  assign n72 = n23 ^ x6 ^ 1'b0 ;
  assign n73 = x1 & n72 ;
  assign n74 = n69 ^ n48 ^ n13 ;
  assign n75 = n74 ^ n27 ^ 1'b0 ;
  assign n76 = n44 & n75 ;
  assign n78 = x9 ^ x7 ^ 1'b0 ;
  assign n79 = x11 & n78 ;
  assign n77 = n23 & ~n27 ;
  assign n80 = n79 ^ n77 ^ 1'b0 ;
  assign n81 = x10 & ~n80 ;
  assign n82 = x2 & n81 ;
  assign n83 = n82 ^ n31 ^ 1'b0 ;
  assign n84 = n54 & ~n77 ;
  assign n85 = ~n51 & n84 ;
  assign n86 = ( x3 & ~x5 ) | ( x3 & n28 ) | ( ~x5 & n28 ) ;
  assign n87 = x3 & n86 ;
  assign n88 = n87 ^ n27 ^ 1'b0 ;
  assign n89 = n88 ^ n61 ^ 1'b0 ;
  assign n90 = n76 ^ n36 ^ 1'b0 ;
  assign n91 = n89 & n90 ;
  assign n92 = x5 & ~n47 ;
  assign n93 = ~x7 & n92 ;
  assign n94 = n79 & n88 ;
  assign n95 = n94 ^ n67 ^ 1'b0 ;
  assign n96 = n27 & n95 ;
  assign n97 = ~n56 & n96 ;
  assign n98 = n97 ^ n54 ^ 1'b0 ;
  assign n99 = x4 & ~n98 ;
  assign n100 = ~n91 & n99 ;
  assign n102 = n54 ^ n38 ^ 1'b0 ;
  assign n103 = x2 & n102 ;
  assign n101 = n49 & n63 ;
  assign n104 = n103 ^ n101 ^ 1'b0 ;
  assign n105 = n44 & n53 ;
  assign n106 = n105 ^ n56 ^ n31 ;
  assign n107 = n96 ^ n81 ^ n21 ;
  assign n108 = n107 ^ n17 ^ 1'b0 ;
  assign n109 = n20 | n108 ;
  assign n110 = n33 & ~n109 ;
  assign n111 = x6 & ~n110 ;
  assign n112 = n111 ^ n30 ^ 1'b0 ;
  assign n113 = n15 ^ x4 ^ 1'b0 ;
  assign n114 = n23 & n79 ;
  assign n115 = n13 & n114 ;
  assign n116 = n30 ^ x3 ^ 1'b0 ;
  assign n117 = ~n77 & n116 ;
  assign n118 = n115 | n117 ;
  assign n119 = n118 ^ n116 ^ 1'b0 ;
  assign n120 = ~n20 & n78 ;
  assign n121 = n120 ^ n17 ^ 1'b0 ;
  assign n122 = ( ~n57 & n112 ) | ( ~n57 & n121 ) | ( n112 & n121 ) ;
  assign n123 = n45 ^ n27 ^ 1'b0 ;
  assign n124 = n36 & ~n123 ;
  assign n125 = n45 ^ x9 ^ 1'b0 ;
  assign n126 = n81 & ~n125 ;
  assign n127 = ( n21 & ~n58 ) | ( n21 & n96 ) | ( ~n58 & n96 ) ;
  assign n128 = x9 & ~n20 ;
  assign n129 = n128 ^ n108 ^ 1'b0 ;
  assign n130 = n51 ^ n25 ^ 1'b0 ;
  assign n131 = ~n27 & n130 ;
  assign n132 = ( n35 & ~n48 ) | ( n35 & n61 ) | ( ~n48 & n61 ) ;
  assign n133 = n43 ^ n13 ^ 1'b0 ;
  assign n134 = n133 ^ n120 ^ 1'b0 ;
  assign n135 = n94 | n134 ;
  assign n136 = n61 | n135 ;
  assign n138 = x8 & n26 ;
  assign n137 = x2 & n23 ;
  assign n139 = n138 ^ n137 ^ 1'b0 ;
  assign n140 = x6 | n139 ;
  assign n141 = x11 & ~n119 ;
  assign n142 = ~x9 & n141 ;
  assign n143 = x9 & n96 ;
  assign n144 = ~n73 & n143 ;
  assign n145 = ~n40 & n81 ;
  assign n146 = n145 ^ n51 ^ 1'b0 ;
  assign n147 = n146 ^ n35 ^ x10 ;
  assign n148 = n103 & ~n147 ;
  assign n149 = x11 & n31 ;
  assign n150 = n27 & n149 ;
  assign n151 = x5 & n49 ;
  assign n152 = ~n57 & n151 ;
  assign n153 = n27 & ~n152 ;
  assign n154 = n153 ^ n25 ^ 1'b0 ;
  assign n157 = ~n56 & n81 ;
  assign n158 = n47 & n157 ;
  assign n159 = n108 & ~n158 ;
  assign n155 = n113 & n121 ;
  assign n156 = n71 | n155 ;
  assign n160 = n159 ^ n156 ^ 1'b0 ;
  assign n161 = n63 & ~n106 ;
  assign n162 = n144 & n161 ;
  assign n163 = n35 ^ n27 ^ 1'b0 ;
  assign n164 = ( ~x1 & x6 ) | ( ~x1 & n163 ) | ( x6 & n163 ) ;
  assign n169 = n81 ^ n77 ^ n33 ;
  assign n165 = n115 ^ n74 ^ n27 ;
  assign n166 = n165 ^ n107 ^ 1'b0 ;
  assign n167 = n27 & n166 ;
  assign n168 = n54 & n167 ;
  assign n170 = n169 ^ n168 ^ 1'b0 ;
  assign n171 = n27 & n170 ;
  assign n172 = n112 ^ n63 ^ 1'b0 ;
  assign n173 = n125 | n172 ;
  assign n174 = n27 & ~n173 ;
  assign n175 = ~n91 & n174 ;
  assign n176 = n44 & ~n175 ;
  assign n177 = ~n49 & n176 ;
  assign n178 = n26 | n60 ;
  assign n179 = n88 & ~n178 ;
  assign n180 = n83 & ~n133 ;
  assign n181 = n180 ^ n63 ^ 1'b0 ;
  assign n182 = n179 & ~n181 ;
  assign n183 = ( x8 & n52 ) | ( x8 & ~n121 ) | ( n52 & ~n121 ) ;
  assign n184 = ( n17 & n61 ) | ( n17 & ~n159 ) | ( n61 & ~n159 ) ;
  assign n185 = n44 ^ n21 ^ 1'b0 ;
  assign n186 = n93 | n185 ;
  assign n187 = n186 ^ n138 ^ 1'b0 ;
  assign n188 = n52 | n187 ;
  assign n189 = n188 ^ n186 ^ 1'b0 ;
  assign n190 = ~n93 & n138 ;
  assign n191 = n181 & n190 ;
  assign n194 = n35 ^ n21 ^ 1'b0 ;
  assign n192 = n56 & ~n85 ;
  assign n193 = n49 & ~n192 ;
  assign n195 = n194 ^ n193 ^ 1'b0 ;
  assign n198 = n165 ^ n43 ^ 1'b0 ;
  assign n199 = ~n71 & n198 ;
  assign n196 = n71 | n158 ;
  assign n197 = n196 ^ n74 ^ 1'b0 ;
  assign n200 = n199 ^ n197 ^ n100 ;
  assign n201 = n200 ^ n144 ^ 1'b0 ;
  assign n202 = n139 | n201 ;
  assign n203 = n67 ^ n51 ^ 1'b0 ;
  assign n204 = n13 | n203 ;
  assign n205 = n126 & n204 ;
  assign n206 = n135 | n205 ;
  assign n207 = n202 & ~n206 ;
  assign n208 = n36 & n63 ;
  assign n209 = n51 ^ n47 ^ 1'b0 ;
  assign n210 = ~n112 & n209 ;
  assign n211 = n210 ^ n63 ^ 1'b0 ;
  assign n212 = n208 & n211 ;
  assign n213 = n73 ^ n61 ^ n23 ;
  assign n214 = n179 ^ n49 ^ x3 ;
  assign n215 = n214 ^ n126 ^ 1'b0 ;
  assign n216 = ~n213 & n215 ;
  assign n217 = ~n47 & n103 ;
  assign n218 = n217 ^ n74 ^ 1'b0 ;
  assign n219 = ~n184 & n218 ;
  assign n220 = n107 & n120 ;
  assign n221 = n38 ^ x4 ^ 1'b0 ;
  assign n222 = ( n60 & ~n100 ) | ( n60 & n221 ) | ( ~n100 & n221 ) ;
  assign n223 = n56 & ~n222 ;
  assign n224 = n223 ^ n94 ^ n65 ;
  assign n225 = ( n103 & n131 ) | ( n103 & n224 ) | ( n131 & n224 ) ;
  assign n227 = n204 ^ n61 ^ 1'b0 ;
  assign n226 = n169 ^ n98 ^ n91 ;
  assign n228 = n227 ^ n226 ^ 1'b0 ;
  assign n229 = n60 | n147 ;
  assign n230 = n229 ^ n54 ^ 1'b0 ;
  assign n231 = ~n228 & n230 ;
  assign n232 = n182 ^ n147 ^ 1'b0 ;
  assign n233 = n167 & n232 ;
  assign n234 = n223 ^ n83 ^ x5 ;
  assign n235 = ~n88 & n150 ;
  assign n236 = n235 ^ x6 ^ 1'b0 ;
  assign n237 = ~n183 & n236 ;
  assign n238 = n163 ^ n125 ^ 1'b0 ;
  assign n239 = n163 & ~n238 ;
  assign n240 = x1 & n144 ;
  assign n241 = n240 ^ n21 ^ 1'b0 ;
  assign n242 = n148 ^ n124 ^ 1'b0 ;
  assign n243 = n56 | n242 ;
  assign n244 = ( n113 & ~n241 ) | ( n113 & n243 ) | ( ~n241 & n243 ) ;
  assign n245 = n139 ^ n77 ^ 1'b0 ;
  assign n246 = ~n189 & n245 ;
  assign n247 = n27 & ~n162 ;
  assign n248 = n116 & n247 ;
  assign n249 = n218 & ~n248 ;
  assign n250 = ~n204 & n244 ;
  assign n253 = x1 & n147 ;
  assign n251 = x2 & ~n43 ;
  assign n252 = n150 | n251 ;
  assign n254 = n253 ^ n252 ^ 1'b0 ;
  assign n255 = n93 ^ n73 ^ 1'b0 ;
  assign n256 = n149 | n205 ;
  assign n257 = n13 & ~n256 ;
  assign n258 = n255 | n257 ;
  assign n259 = n175 & ~n258 ;
  assign n260 = n244 ^ n183 ^ 1'b0 ;
  assign n262 = n100 | n142 ;
  assign n263 = n262 ^ n138 ^ 1'b0 ;
  assign n261 = n224 ^ n202 ^ n27 ;
  assign n264 = n263 ^ n261 ^ 1'b0 ;
  assign n265 = ~n56 & n132 ;
  assign n266 = x1 | n192 ;
  assign n267 = n266 ^ n227 ^ 1'b0 ;
  assign n268 = n124 | n140 ;
  assign n269 = n58 | n268 ;
  assign n270 = ( ~n149 & n159 ) | ( ~n149 & n173 ) | ( n159 & n173 ) ;
  assign n271 = n270 ^ n216 ^ n17 ;
  assign n272 = n56 ^ x2 ^ 1'b0 ;
  assign n273 = x9 & ~n272 ;
  assign n274 = n224 & n273 ;
  assign n275 = ~n54 & n274 ;
  assign n276 = ~n69 & n81 ;
  assign n277 = ~n107 & n276 ;
  assign n278 = n112 | n119 ;
  assign n279 = n61 | n278 ;
  assign n280 = ( n36 & n54 ) | ( n36 & n152 ) | ( n54 & n152 ) ;
  assign n281 = n280 ^ n126 ^ 1'b0 ;
  assign n282 = n56 & n281 ;
  assign n283 = n122 & ~n211 ;
  assign n284 = n283 ^ n105 ^ 1'b0 ;
  assign n285 = ~n67 & n284 ;
  assign n286 = ~n57 & n285 ;
  assign n288 = n107 ^ n105 ^ 1'b0 ;
  assign n289 = n288 ^ n67 ^ 1'b0 ;
  assign n290 = ~n112 & n289 ;
  assign n287 = n208 ^ n45 ^ 1'b0 ;
  assign n291 = n290 ^ n287 ^ 1'b0 ;
  assign n292 = n124 ^ x2 ^ 1'b0 ;
  assign n293 = n155 | n218 ;
  assign n294 = n293 ^ n33 ^ 1'b0 ;
  assign n295 = n266 | n294 ;
  assign n296 = n295 ^ n290 ^ n181 ;
  assign n297 = n57 & n265 ;
  assign n298 = n40 & ~n65 ;
  assign n299 = n165 & ~n298 ;
  assign n300 = n285 ^ n81 ^ 1'b0 ;
  assign n301 = ~n33 & n300 ;
  assign n304 = n273 ^ n235 ^ 1'b0 ;
  assign n305 = ~n179 & n304 ;
  assign n302 = n192 & ~n204 ;
  assign n303 = n61 & ~n302 ;
  assign n306 = n305 ^ n303 ^ 1'b0 ;
  assign n307 = n218 ^ n124 ^ 1'b0 ;
  assign n308 = n147 & ~n155 ;
  assign n309 = n307 & n308 ;
  assign n310 = n209 ^ n91 ^ 1'b0 ;
  assign n311 = ~n224 & n310 ;
  assign n312 = n311 ^ n65 ^ 1'b0 ;
  assign n313 = n25 & ~n47 ;
  assign n314 = ~n76 & n313 ;
  assign n315 = n295 & ~n314 ;
  assign n316 = ~n271 & n315 ;
  assign n317 = n115 ^ x0 ^ 1'b0 ;
  assign n318 = n317 ^ n69 ^ n52 ;
  assign n319 = n318 ^ n51 ^ 1'b0 ;
  assign n320 = n54 & n319 ;
  assign n321 = n320 ^ n148 ^ 1'b0 ;
  assign n322 = n35 | n321 ;
  assign n323 = n17 & ~n144 ;
  assign n324 = n323 ^ n57 ^ 1'b0 ;
  assign n325 = n322 | n324 ;
  assign n330 = n94 ^ n85 ^ 1'b0 ;
  assign n326 = ~n48 & n213 ;
  assign n327 = n326 ^ n139 ^ 1'b0 ;
  assign n328 = n304 | n327 ;
  assign n329 = ~n112 & n328 ;
  assign n331 = n330 ^ n329 ^ 1'b0 ;
  assign n332 = ~n213 & n223 ;
  assign n333 = ~n113 & n332 ;
  assign n334 = ~n150 & n333 ;
  assign n335 = n120 ^ x7 ^ 1'b0 ;
  assign n336 = ~x6 & n209 ;
  assign n337 = n261 ^ n229 ^ 1'b0 ;
  assign n338 = n249 & ~n337 ;
  assign n343 = n54 | n115 ;
  assign n339 = n54 ^ n27 ^ 1'b0 ;
  assign n340 = n339 ^ n63 ^ 1'b0 ;
  assign n341 = n318 & n340 ;
  assign n342 = ~x2 & n341 ;
  assign n344 = n343 ^ n342 ^ n89 ;
  assign n345 = n330 ^ n323 ^ 1'b0 ;
  assign n346 = n345 ^ n261 ^ 1'b0 ;
  assign n347 = n344 | n346 ;
  assign n348 = n249 ^ n208 ^ 1'b0 ;
  assign n349 = n147 & n348 ;
  assign n350 = n200 ^ n27 ^ 1'b0 ;
  assign n351 = n197 & n350 ;
  assign n352 = x2 & ~n351 ;
  assign n354 = n144 ^ x7 ^ 1'b0 ;
  assign n355 = x2 & n354 ;
  assign n356 = n355 ^ n253 ^ 1'b0 ;
  assign n357 = ( n69 & n116 ) | ( n69 & ~n356 ) | ( n116 & ~n356 ) ;
  assign n353 = ~n19 & n171 ;
  assign n358 = n357 ^ n353 ^ 1'b0 ;
  assign n359 = n192 ^ n121 ^ 1'b0 ;
  assign n360 = n213 | n359 ;
  assign n361 = n360 ^ n61 ^ 1'b0 ;
  assign n362 = n330 | n361 ;
  assign n365 = ( n130 & n155 ) | ( n130 & ~n179 ) | ( n155 & ~n179 ) ;
  assign n363 = n285 ^ n57 ^ 1'b0 ;
  assign n364 = n349 & n363 ;
  assign n366 = n365 ^ n364 ^ 1'b0 ;
  assign n367 = ~n79 & n212 ;
  assign n368 = n246 ^ n105 ^ 1'b0 ;
  assign n373 = n140 ^ n57 ^ 1'b0 ;
  assign n374 = n373 ^ n261 ^ n121 ;
  assign n369 = n213 | n223 ;
  assign n370 = n15 | n369 ;
  assign n371 = n93 & ~n370 ;
  assign n372 = ~n112 & n371 ;
  assign n375 = n374 ^ n372 ^ 1'b0 ;
  assign n376 = ~n323 & n375 ;
  assign n377 = n67 | n104 ;
  assign n378 = n117 & ~n377 ;
  assign n379 = n378 ^ x7 ^ 1'b0 ;
  assign n380 = n222 ^ n189 ^ 1'b0 ;
  assign n381 = n380 ^ n325 ^ 1'b0 ;
  assign n382 = n51 & ~n381 ;
  assign n386 = n177 ^ n125 ^ 1'b0 ;
  assign n383 = ~n112 & n130 ;
  assign n384 = n383 ^ n235 ^ 1'b0 ;
  assign n385 = n115 | n384 ;
  assign n387 = n386 ^ n385 ^ 1'b0 ;
  assign n388 = ( n21 & n254 ) | ( n21 & ~n387 ) | ( n254 & ~n387 ) ;
  assign n389 = x2 & ~n77 ;
  assign n390 = n48 & n389 ;
  assign n391 = n119 | n390 ;
  assign n392 = n17 & ~n391 ;
  assign n393 = n392 ^ n146 ^ n61 ;
  assign n394 = n76 & ~n88 ;
  assign n395 = ~n25 & n394 ;
  assign n396 = n23 & n395 ;
  assign n397 = n396 ^ n322 ^ n221 ;
  assign n398 = n227 ^ n56 ^ 1'b0 ;
  assign n399 = n398 ^ n98 ^ 1'b0 ;
  assign n400 = x6 & ~n399 ;
  assign n401 = n400 ^ n113 ^ 1'b0 ;
  assign n402 = n320 ^ n144 ^ 1'b0 ;
  assign n403 = ( n93 & n211 ) | ( n93 & n402 ) | ( n211 & n402 ) ;
  assign n404 = n20 | n40 ;
  assign n405 = n117 ^ n26 ^ 1'b0 ;
  assign n406 = ~n152 & n405 ;
  assign n407 = x4 & ~n85 ;
  assign n408 = ~n406 & n407 ;
  assign n409 = n408 ^ n177 ^ n146 ;
  assign n410 = n79 & n409 ;
  assign n411 = n410 ^ n320 ^ 1'b0 ;
  assign n412 = n147 ^ n51 ^ 1'b0 ;
  assign n413 = x5 & n113 ;
  assign n414 = n47 & n413 ;
  assign n415 = n202 ^ n116 ^ 1'b0 ;
  assign n416 = x8 & ~n288 ;
  assign n417 = n415 & n416 ;
  assign n418 = n417 ^ n380 ^ 1'b0 ;
  assign n419 = ~n414 & n418 ;
  assign n420 = ( x1 & n33 ) | ( x1 & n125 ) | ( n33 & n125 ) ;
  assign n421 = n420 ^ n221 ^ 1'b0 ;
  assign n422 = n27 & ~n421 ;
  assign n423 = ~n225 & n422 ;
  assign n424 = n305 ^ n255 ^ 1'b0 ;
  assign n425 = ~n414 & n424 ;
  assign n427 = n138 ^ n120 ^ 1'b0 ;
  assign n428 = ~n69 & n427 ;
  assign n429 = ~n35 & n221 ;
  assign n430 = n429 ^ n139 ^ 1'b0 ;
  assign n431 = n430 ^ n228 ^ 1'b0 ;
  assign n432 = n431 ^ x11 ^ 1'b0 ;
  assign n433 = ( n150 & ~n428 ) | ( n150 & n432 ) | ( ~n428 & n432 ) ;
  assign n426 = n121 & n124 ;
  assign n434 = n433 ^ n426 ^ 1'b0 ;
  assign n435 = n181 ^ n179 ^ 1'b0 ;
  assign n436 = ~n19 & n435 ;
  assign n437 = n105 ^ n94 ^ 1'b0 ;
  assign n438 = n436 & ~n437 ;
  assign n439 = n33 ^ n15 ^ 1'b0 ;
  assign n440 = n160 ^ n96 ^ 1'b0 ;
  assign n441 = n439 & n440 ;
  assign n442 = n163 ^ n52 ^ 1'b0 ;
  assign n443 = n384 & ~n442 ;
  assign n444 = ~n211 & n443 ;
  assign n445 = ~n441 & n444 ;
  assign n446 = n35 & n182 ;
  assign n447 = n446 ^ n182 ^ n148 ;
  assign n448 = n447 ^ n136 ^ 1'b0 ;
  assign n449 = n76 & n402 ;
  assign n450 = n205 & n449 ;
  assign n451 = n163 ^ n133 ^ 1'b0 ;
  assign n452 = ~n88 & n417 ;
  assign n453 = x8 & n61 ;
  assign n454 = n115 | n330 ;
  assign n455 = n121 & ~n417 ;
  assign n456 = ~n129 & n455 ;
  assign n457 = ~n112 & n113 ;
  assign n458 = ~n223 & n457 ;
  assign n459 = ( ~n261 & n267 ) | ( ~n261 & n458 ) | ( n267 & n458 ) ;
  assign n460 = n239 & n459 ;
  assign n461 = ~n320 & n460 ;
  assign n462 = ~n67 & n120 ;
  assign n463 = ~n363 & n462 ;
  assign n464 = n224 & ~n463 ;
  assign n465 = n464 ^ x6 ^ 1'b0 ;
  assign n466 = ~n275 & n465 ;
  assign n467 = n15 | n131 ;
  assign n468 = n467 ^ n175 ^ 1'b0 ;
  assign n469 = n458 ^ n67 ^ 1'b0 ;
  assign n470 = ~n15 & n469 ;
  assign n471 = ~n85 & n121 ;
  assign n472 = n471 ^ n147 ^ n115 ;
  assign n473 = n188 ^ n150 ^ 1'b0 ;
  assign n474 = ( n392 & n418 ) | ( n392 & n473 ) | ( n418 & n473 ) ;
  assign n475 = n36 & n61 ;
  assign n476 = n474 | n475 ;
  assign n477 = n476 ^ n216 ^ 1'b0 ;
  assign n478 = n273 ^ n177 ^ 1'b0 ;
  assign n479 = n125 & n478 ;
  assign n480 = n384 ^ n38 ^ 1'b0 ;
  assign n481 = n290 | n480 ;
  assign n482 = n366 & ~n481 ;
  assign n483 = n61 & ~n465 ;
  assign n484 = n483 ^ n397 ^ 1'b0 ;
  assign n485 = n221 ^ n119 ^ 1'b0 ;
  assign n486 = x6 & n432 ;
  assign n487 = n485 & n486 ;
  assign n488 = ( ~n98 & n315 ) | ( ~n98 & n487 ) | ( n315 & n487 ) ;
  assign n489 = n369 ^ n186 ^ 1'b0 ;
  assign n490 = n227 ^ n104 ^ x4 ;
  assign n491 = n104 | n490 ;
  assign n492 = n144 | n491 ;
  assign n493 = n325 | n492 ;
  assign n494 = n214 ^ n147 ^ n67 ;
  assign n495 = n494 ^ n384 ^ n317 ;
  assign n499 = n369 ^ n173 ^ 1'b0 ;
  assign n500 = n160 & n499 ;
  assign n496 = ~n251 & n286 ;
  assign n497 = ~n400 & n496 ;
  assign n498 = ( n170 & ~n411 ) | ( n170 & n497 ) | ( ~n411 & n497 ) ;
  assign n501 = n500 ^ n498 ^ 1'b0 ;
  assign n502 = ~n152 & n501 ;
  assign n503 = ~n207 & n280 ;
  assign n504 = n503 ^ n227 ^ 1'b0 ;
  assign n505 = n147 & n504 ;
  assign n506 = n285 ^ n205 ^ n188 ;
  assign n507 = n49 & ~n433 ;
  assign n508 = n378 & n507 ;
  assign n509 = n244 ^ n131 ^ n88 ;
  assign n510 = n509 ^ n323 ^ 1'b0 ;
  assign n511 = n28 & n115 ;
  assign n512 = n122 | n511 ;
  assign n513 = n512 ^ n73 ^ 1'b0 ;
  assign n514 = x6 & n513 ;
  assign n515 = n48 & n514 ;
  assign n516 = n515 ^ n110 ^ 1'b0 ;
  assign n517 = n290 & n516 ;
  assign n518 = n216 | n261 ;
  assign n519 = n422 ^ n296 ^ 1'b0 ;
  assign n520 = n519 ^ n371 ^ 1'b0 ;
  assign n521 = ~n518 & n520 ;
  assign n522 = n318 & n320 ;
  assign n523 = ~n83 & n522 ;
  assign n524 = n126 & ~n428 ;
  assign n525 = n524 ^ n183 ^ 1'b0 ;
  assign n526 = n437 ^ n338 ^ 1'b0 ;
  assign n527 = x11 & n526 ;
  assign n528 = ~n17 & n244 ;
  assign n529 = n170 & n222 ;
  assign n530 = n529 ^ n119 ^ 1'b0 ;
  assign n531 = n100 ^ n89 ^ 1'b0 ;
  assign n532 = n530 & ~n531 ;
  assign n533 = ~n411 & n532 ;
  assign n534 = n343 ^ n285 ^ 1'b0 ;
  assign n535 = n363 & ~n534 ;
  assign n538 = x2 & ~n302 ;
  assign n539 = ~n63 & n538 ;
  assign n540 = n539 ^ n194 ^ 1'b0 ;
  assign n541 = n540 ^ x1 ^ 1'b0 ;
  assign n536 = n73 & n222 ;
  assign n537 = ~n21 & n536 ;
  assign n542 = n541 ^ n537 ^ 1'b0 ;
  assign n543 = ~n445 & n472 ;
  assign n544 = n144 | n541 ;
  assign n545 = n544 ^ n25 ^ 1'b0 ;
  assign n546 = ~n67 & n392 ;
  assign n547 = n546 ^ n188 ^ 1'b0 ;
  assign n548 = n317 ^ n227 ^ 1'b0 ;
  assign n549 = n301 | n548 ;
  assign n550 = ~n150 & n241 ;
  assign n551 = ~n402 & n550 ;
  assign n552 = n209 & n551 ;
  assign n553 = n552 ^ n290 ^ 1'b0 ;
  assign n555 = ( n83 & n244 ) | ( n83 & n453 ) | ( n244 & n453 ) ;
  assign n556 = n36 ^ x1 ^ 1'b0 ;
  assign n557 = ~n356 & n556 ;
  assign n558 = n557 ^ n21 ^ 1'b0 ;
  assign n559 = n555 & ~n558 ;
  assign n554 = n243 | n523 ;
  assign n560 = n559 ^ n554 ^ 1'b0 ;
  assign n561 = ( ~n45 & n88 ) | ( ~n45 & n177 ) | ( n88 & n177 ) ;
  assign n562 = ~n56 & n561 ;
  assign n563 = n541 | n562 ;
  assign n567 = n83 & n314 ;
  assign n568 = n567 ^ n408 ^ 1'b0 ;
  assign n569 = n241 & n532 ;
  assign n570 = ~n568 & n569 ;
  assign n564 = n446 ^ n135 ^ n86 ;
  assign n565 = ~n49 & n564 ;
  assign n566 = n19 | n565 ;
  assign n571 = n570 ^ n566 ^ 1'b0 ;
  assign n572 = n89 & n152 ;
  assign n573 = n124 | n275 ;
  assign n574 = n572 | n573 ;
  assign n578 = ~n54 & n61 ;
  assign n577 = n98 | n216 ;
  assign n576 = n503 ^ n301 ^ 1'b0 ;
  assign n579 = n578 ^ n577 ^ n576 ;
  assign n580 = n365 & n579 ;
  assign n581 = n580 ^ n132 ^ 1'b0 ;
  assign n575 = n23 & n188 ;
  assign n582 = n581 ^ n575 ^ 1'b0 ;
  assign n583 = ~n124 & n283 ;
  assign n584 = n420 & n583 ;
  assign n585 = n211 ^ n159 ^ 1'b0 ;
  assign n586 = n135 | n585 ;
  assign n587 = n458 | n586 ;
  assign n588 = n251 & ~n587 ;
  assign n589 = x1 & ~n224 ;
  assign n590 = n589 ^ n120 ^ 1'b0 ;
  assign n591 = n590 ^ n560 ^ 1'b0 ;
  assign n592 = n417 ^ x1 ^ 1'b0 ;
  assign n593 = n110 & ~n592 ;
  assign n594 = n551 ^ n235 ^ 1'b0 ;
  assign n595 = ~n33 & n594 ;
  assign n596 = ~n188 & n498 ;
  assign n597 = n596 ^ n533 ^ 1'b0 ;
  assign n598 = n147 & n188 ;
  assign n599 = n234 ^ n183 ^ 1'b0 ;
  assign n600 = ~n52 & n599 ;
  assign n601 = n212 & n600 ;
  assign n602 = n452 ^ n388 ^ n85 ;
  assign n603 = n601 | n602 ;
  assign n604 = n224 | n603 ;
  assign n605 = n546 ^ n386 ^ 1'b0 ;
  assign n606 = ( n552 & ~n600 ) | ( n552 & n605 ) | ( ~n600 & n605 ) ;
  assign n607 = n287 | n606 ;
  assign n608 = n330 | n363 ;
  assign n609 = n593 ^ n264 ^ 1'b0 ;
  assign n610 = n27 ^ x4 ^ 1'b0 ;
  assign n611 = ~n296 & n610 ;
  assign n612 = ( ~n228 & n423 ) | ( ~n228 & n611 ) | ( n423 & n611 ) ;
  assign n613 = ~n219 & n345 ;
  assign n614 = ~n451 & n613 ;
  assign n615 = n414 ^ n191 ^ n36 ;
  assign n616 = n103 & n334 ;
  assign n617 = n602 & n616 ;
  assign n618 = ~n31 & n194 ;
  assign n619 = n618 ^ n150 ^ 1'b0 ;
  assign n620 = ( n316 & ~n358 ) | ( n316 & n619 ) | ( ~n358 & n619 ) ;
  assign n621 = n620 ^ n138 ^ 1'b0 ;
  assign n622 = n52 | n621 ;
  assign n623 = n445 ^ n251 ^ 1'b0 ;
  assign n624 = n160 ^ n76 ^ 1'b0 ;
  assign n625 = ~n623 & n624 ;
  assign n626 = x6 & n527 ;
  assign n627 = n626 ^ n525 ^ 1'b0 ;
  assign n629 = n63 & n96 ;
  assign n630 = n629 ^ n514 ^ 1'b0 ;
  assign n631 = n133 | n280 ;
  assign n632 = ~n630 & n631 ;
  assign n633 = n330 & n632 ;
  assign n628 = n335 | n540 ;
  assign n634 = n633 ^ n628 ^ 1'b0 ;
  assign n635 = n155 ^ n105 ^ 1'b0 ;
  assign n636 = n565 ^ n513 ^ 1'b0 ;
  assign n637 = n615 & ~n636 ;
  assign n638 = n184 & ~n395 ;
  assign n639 = n390 | n638 ;
  assign n640 = n639 ^ n125 ^ 1'b0 ;
  assign n641 = n468 & ~n640 ;
  assign n642 = n69 & n107 ;
  assign n643 = ~n162 & n306 ;
  assign n644 = n643 ^ n403 ^ 1'b0 ;
  assign n645 = n644 ^ n56 ^ 1'b0 ;
  assign n646 = n642 | n645 ;
  assign n647 = n119 | n646 ;
  assign n648 = n205 ^ n38 ^ 1'b0 ;
  assign n649 = n648 ^ n439 ^ 1'b0 ;
  assign n650 = ~n191 & n649 ;
  assign n651 = n650 ^ n561 ^ 1'b0 ;
  assign n652 = n651 ^ n641 ^ n339 ;
  assign n653 = x9 & ~n139 ;
  assign n654 = n653 ^ n170 ^ 1'b0 ;
  assign n655 = n342 ^ n226 ^ x3 ;
  assign n656 = n655 ^ n273 ^ 1'b0 ;
  assign n657 = ~n654 & n656 ;
  assign n658 = n398 & ~n620 ;
  assign n659 = ~n657 & n658 ;
  assign n660 = n439 ^ x7 ^ 1'b0 ;
  assign n661 = ~n640 & n660 ;
  assign n662 = n167 & ~n228 ;
  assign n663 = ~n233 & n662 ;
  assign n664 = ~n85 & n663 ;
  assign n665 = n406 & ~n664 ;
  assign n666 = n665 ^ n380 ^ 1'b0 ;
  assign n667 = ( ~n200 & n661 ) | ( ~n200 & n666 ) | ( n661 & n666 ) ;
  assign n668 = n334 & n484 ;
  assign n669 = ~n610 & n668 ;
  assign n670 = n669 ^ n309 ^ 1'b0 ;
  assign n671 = n645 | n670 ;
  assign n672 = n260 ^ n113 ^ 1'b0 ;
  assign n673 = n35 & n672 ;
  assign n674 = n380 & n673 ;
  assign n675 = n674 ^ n265 ^ 1'b0 ;
  assign n676 = n450 & n451 ;
  assign n677 = ( x0 & n296 ) | ( x0 & ~n676 ) | ( n296 & ~n676 ) ;
  assign n679 = n125 | n188 ;
  assign n680 = n173 & ~n679 ;
  assign n681 = n100 & ~n680 ;
  assign n678 = n214 & ~n610 ;
  assign n682 = n681 ^ n678 ^ 1'b0 ;
  assign n683 = n248 & ~n458 ;
  assign n684 = n492 ^ n160 ^ 1'b0 ;
  assign n685 = n572 ^ n297 ^ 1'b0 ;
  assign n686 = n685 ^ n362 ^ 1'b0 ;
  assign n687 = n684 & n686 ;
  assign n691 = n437 ^ n17 ^ 1'b0 ;
  assign n692 = n436 & ~n691 ;
  assign n688 = n286 & ~n371 ;
  assign n689 = n327 & n688 ;
  assign n690 = n411 & n689 ;
  assign n693 = n692 ^ n690 ^ 1'b0 ;
  assign n694 = n317 | n693 ;
  assign n695 = n568 ^ n452 ^ n110 ;
  assign n696 = n239 | n695 ;
  assign n697 = n642 ^ n81 ^ 1'b0 ;
  assign n698 = n291 & ~n697 ;
  assign n700 = n110 | n292 ;
  assign n699 = n200 ^ n31 ^ 1'b0 ;
  assign n701 = n700 ^ n699 ^ n481 ;
  assign n702 = n479 & n530 ;
  assign n703 = n702 ^ n191 ^ 1'b0 ;
  assign n704 = n265 | n342 ;
  assign n705 = n588 ^ n98 ^ 1'b0 ;
  assign n706 = n231 & n705 ;
  assign n707 = ~x1 & n280 ;
  assign n708 = n36 & ~n707 ;
  assign n709 = n249 ^ n131 ^ 1'b0 ;
  assign n710 = n709 ^ n666 ^ n305 ;
  assign n711 = n345 ^ n271 ^ 1'b0 ;
  assign n712 = n241 & n711 ;
  assign n713 = n27 & ~n317 ;
  assign n714 = n713 ^ n124 ^ 1'b0 ;
  assign n715 = n152 | n714 ;
  assign n716 = n712 | n715 ;
  assign n717 = n344 & ~n548 ;
  assign n719 = ~n417 & n432 ;
  assign n720 = ~n358 & n719 ;
  assign n718 = n318 & ~n607 ;
  assign n721 = n720 ^ n718 ^ 1'b0 ;
  assign n723 = n93 ^ n47 ^ 1'b0 ;
  assign n724 = ~n285 & n723 ;
  assign n722 = n409 & ~n420 ;
  assign n725 = n724 ^ n722 ^ 1'b0 ;
  assign n726 = n725 ^ n482 ^ 1'b0 ;
  assign n727 = n601 | n726 ;
  assign n728 = n417 ^ n368 ^ 1'b0 ;
  assign n729 = ~n139 & n728 ;
  assign n730 = n131 | n422 ;
  assign n731 = n730 ^ n264 ^ 1'b0 ;
  assign n732 = n255 & n731 ;
  assign n733 = n333 ^ n120 ^ 1'b0 ;
  assign n734 = n733 ^ n26 ^ 1'b0 ;
  assign n735 = n734 ^ n598 ^ 1'b0 ;
  assign n736 = ~n205 & n735 ;
  assign n737 = n162 & ~n397 ;
  assign n738 = n390 ^ n298 ^ 1'b0 ;
  assign n739 = ~n584 & n738 ;
  assign n740 = ~n737 & n739 ;
  assign n741 = n563 ^ n497 ^ n406 ;
  assign n742 = ~n685 & n724 ;
  assign n743 = ~n314 & n673 ;
  assign n744 = n743 ^ n724 ^ 1'b0 ;
  assign n745 = n244 & n744 ;
  assign n746 = ~n251 & n351 ;
  assign n747 = n746 ^ n266 ^ n23 ;
  assign n750 = n692 ^ n298 ^ 1'b0 ;
  assign n748 = n121 & n231 ;
  assign n749 = ~x10 & n748 ;
  assign n751 = n750 ^ n749 ^ 1'b0 ;
  assign n752 = n129 & ~n401 ;
  assign n753 = n282 ^ x9 ^ 1'b0 ;
  assign n755 = n200 & n244 ;
  assign n756 = n31 | n755 ;
  assign n757 = n581 & ~n756 ;
  assign n754 = n115 | n226 ;
  assign n758 = n757 ^ n754 ^ 1'b0 ;
  assign n759 = n254 ^ n44 ^ 1'b0 ;
  assign n760 = n436 & n759 ;
  assign n761 = n552 & n760 ;
  assign n762 = n761 ^ n503 ^ 1'b0 ;
  assign n763 = n762 ^ n146 ^ 1'b0 ;
  assign n764 = ~n606 & n763 ;
  assign n765 = n339 ^ n126 ^ 1'b0 ;
  assign n766 = n703 & ~n765 ;
  assign n767 = n248 & ~n373 ;
  assign n768 = ( n65 & n362 ) | ( n65 & ~n767 ) | ( n362 & ~n767 ) ;
  assign n769 = n597 ^ n282 ^ 1'b0 ;
  assign n770 = n588 | n769 ;
  assign n771 = ~n47 & n765 ;
  assign n772 = n771 ^ n339 ^ 1'b0 ;
  assign n773 = n772 ^ n581 ^ 1'b0 ;
  assign n774 = n246 ^ n57 ^ 1'b0 ;
  assign n775 = n774 ^ n119 ^ 1'b0 ;
  assign n776 = n661 & ~n775 ;
  assign n777 = n776 ^ n517 ^ 1'b0 ;
  assign n778 = n746 ^ x6 ^ 1'b0 ;
  assign n779 = ~n468 & n637 ;
  assign n780 = n779 ^ n710 ^ 1'b0 ;
  assign n781 = n681 ^ n61 ^ 1'b0 ;
  assign n782 = n194 | n204 ;
  assign n783 = n288 | n782 ;
  assign n784 = n576 ^ x11 ^ 1'b0 ;
  assign n785 = ~n783 & n784 ;
  assign n786 = n576 & n785 ;
  assign n787 = n259 | n575 ;
  assign n788 = n540 & ~n694 ;
  assign n789 = n489 & n788 ;
  assign n790 = n789 ^ n541 ^ 1'b0 ;
  assign n791 = n94 & ~n205 ;
  assign n792 = n130 & n791 ;
  assign n793 = n458 | n664 ;
  assign n794 = n500 & ~n627 ;
  assign n795 = n793 & n794 ;
  assign n796 = ~n645 & n795 ;
  assign n797 = n796 ^ n591 ^ 1'b0 ;
  assign n798 = n749 | n797 ;
  assign n800 = n540 ^ n322 ^ 1'b0 ;
  assign n799 = ~n307 & n373 ;
  assign n801 = n800 ^ n799 ^ 1'b0 ;
  assign n802 = n173 & n418 ;
  assign n803 = n802 ^ n266 ^ 1'b0 ;
  assign n804 = n546 | n803 ;
  assign n805 = ( n448 & n801 ) | ( n448 & ~n804 ) | ( n801 & ~n804 ) ;
  assign n806 = n620 ^ n262 ^ 1'b0 ;
  assign n807 = ~n150 & n382 ;
  assign n808 = n326 & n807 ;
  assign n809 = n322 ^ n106 ^ 1'b0 ;
  assign n810 = n809 ^ n309 ^ 1'b0 ;
  assign n811 = n221 & n810 ;
  assign n812 = n811 ^ n40 ^ 1'b0 ;
  assign n813 = n167 | n421 ;
  assign n814 = n376 & n813 ;
  assign n815 = ~n208 & n814 ;
  assign n816 = n283 & n400 ;
  assign n817 = n257 & n816 ;
  assign n818 = n815 | n817 ;
  assign n819 = n812 | n818 ;
  assign n820 = n105 | n450 ;
  assign n821 = n815 ^ n704 ^ 1'b0 ;
  assign n822 = n83 ^ n25 ^ n23 ;
  assign n823 = n651 | n822 ;
  assign n824 = ~n305 & n823 ;
  assign n825 = n824 ^ n527 ^ 1'b0 ;
  assign n826 = n334 & ~n572 ;
  assign n827 = n826 ^ n572 ^ 1'b0 ;
  assign n828 = n567 ^ n331 ^ n214 ;
  assign n829 = n673 ^ x7 ^ 1'b0 ;
  assign n830 = n150 | n179 ;
  assign n831 = n732 & ~n830 ;
  assign n832 = ~n392 & n792 ;
  assign n833 = x3 & ~n108 ;
  assign n839 = ( ~n23 & n273 ) | ( ~n23 & n298 ) | ( n273 & n298 ) ;
  assign n834 = n317 ^ x6 ^ 1'b0 ;
  assign n835 = n147 & ~n834 ;
  assign n836 = n489 ^ n422 ^ 1'b0 ;
  assign n837 = n835 & ~n836 ;
  assign n838 = ~n45 & n837 ;
  assign n840 = n839 ^ n838 ^ 1'b0 ;
  assign n841 = n216 & n415 ;
  assign n842 = n540 ^ n127 ^ 1'b0 ;
  assign n843 = n461 | n842 ;
  assign n844 = n219 & ~n843 ;
  assign n845 = n170 & n226 ;
  assign n846 = n845 ^ n610 ^ 1'b0 ;
  assign n849 = n333 ^ n248 ^ 1'b0 ;
  assign n847 = n122 | n326 ;
  assign n848 = n76 | n847 ;
  assign n850 = n849 ^ n848 ^ 1'b0 ;
  assign n851 = n433 ^ n183 ^ 1'b0 ;
  assign n852 = n126 ^ n63 ^ 1'b0 ;
  assign n853 = n73 & ~n852 ;
  assign n854 = ~x3 & n853 ;
  assign n855 = n333 ^ n221 ^ 1'b0 ;
  assign n856 = n855 ^ n615 ^ 1'b0 ;
  assign n857 = n644 ^ n110 ^ 1'b0 ;
  assign n858 = n857 ^ n720 ^ 1'b0 ;
  assign n859 = n858 ^ n282 ^ 1'b0 ;
  assign n860 = n856 | n859 ;
  assign n861 = ( ~n47 & n474 ) | ( ~n47 & n676 ) | ( n474 & n676 ) ;
  assign n862 = n625 ^ n340 ^ 1'b0 ;
  assign n863 = n664 ^ n395 ^ 1'b0 ;
  assign n864 = ~n222 & n863 ;
  assign n865 = n255 & n439 ;
  assign n866 = n865 ^ n614 ^ 1'b0 ;
  assign n867 = n67 | n866 ;
  assign n872 = n49 | n106 ;
  assign n873 = ~n127 & n314 ;
  assign n874 = ( n541 & n872 ) | ( n541 & n873 ) | ( n872 & n873 ) ;
  assign n868 = n638 ^ n390 ^ n228 ;
  assign n869 = n868 ^ n334 ^ 1'b0 ;
  assign n870 = ~n630 & n869 ;
  assign n871 = ~n582 & n870 ;
  assign n875 = n874 ^ n871 ^ 1'b0 ;
  assign n876 = n430 & ~n642 ;
  assign n877 = n876 ^ n373 ^ 1'b0 ;
  assign n878 = ( n135 & n226 ) | ( n135 & n582 ) | ( n226 & n582 ) ;
  assign n879 = x11 & ~n390 ;
  assign n880 = ~n478 & n879 ;
  assign n881 = n21 | n139 ;
  assign n882 = n480 ^ n225 ^ 1'b0 ;
  assign n883 = n881 | n882 ;
  assign n884 = n250 & ~n883 ;
  assign n885 = n254 & n382 ;
  assign n886 = n147 & ~n885 ;
  assign n887 = n169 | n390 ;
  assign n888 = n49 & ~n887 ;
  assign n889 = n888 ^ n220 ^ 1'b0 ;
  assign n890 = ( n490 & n543 ) | ( n490 & ~n889 ) | ( n543 & ~n889 ) ;
  assign n891 = n49 & n208 ;
  assign n892 = n81 & ~n357 ;
  assign n893 = n227 & n315 ;
  assign n894 = ~n892 & n893 ;
  assign n895 = n572 ^ n323 ^ 1'b0 ;
  assign n896 = n894 | n895 ;
  assign n897 = n369 ^ n135 ^ 1'b0 ;
  assign n898 = ~n304 & n897 ;
  assign n899 = n86 & ~n898 ;
  assign n900 = n899 ^ n233 ^ 1'b0 ;
  assign n901 = n57 & ~n900 ;
  assign n902 = n459 ^ n165 ^ 1'b0 ;
  assign n903 = n533 | n902 ;
  assign n904 = n903 ^ n697 ^ 1'b0 ;
  assign n905 = n291 ^ n104 ^ 1'b0 ;
  assign n906 = n690 | n905 ;
  assign n907 = n40 & ~n906 ;
  assign n908 = n631 ^ n188 ^ 1'b0 ;
  assign n909 = n600 & n908 ;
  assign n910 = n909 ^ n227 ^ 1'b0 ;
  assign n911 = n126 & n910 ;
  assign n913 = n390 ^ n26 ^ 1'b0 ;
  assign n914 = ~n173 & n913 ;
  assign n912 = ~n577 & n788 ;
  assign n915 = n914 ^ n912 ^ 1'b0 ;
  assign n916 = n307 & n595 ;
  assign n917 = n863 | n916 ;
  assign n919 = n835 & ~n899 ;
  assign n918 = n108 & ~n541 ;
  assign n920 = n919 ^ n918 ^ n85 ;
  assign n921 = n627 ^ n625 ^ 1'b0 ;
  assign n922 = n858 | n921 ;
  assign n924 = ~n77 & n211 ;
  assign n925 = ~n343 & n924 ;
  assign n926 = n392 & n925 ;
  assign n923 = n52 | n448 ;
  assign n927 = n926 ^ n923 ^ 1'b0 ;
  assign n928 = n367 & ~n922 ;
  assign n929 = n928 ^ n832 ^ 1'b0 ;
  assign n930 = n35 | n158 ;
  assign n931 = n930 ^ n76 ^ 1'b0 ;
  assign n932 = ~n772 & n931 ;
  assign n933 = n222 & n235 ;
  assign n934 = ~n849 & n933 ;
  assign n935 = n150 ^ n126 ^ 1'b0 ;
  assign n936 = n225 & ~n935 ;
  assign n937 = n936 ^ n234 ^ 1'b0 ;
  assign n938 = n934 | n937 ;
  assign n939 = n261 ^ n251 ^ 1'b0 ;
  assign n940 = n398 & n939 ;
  assign n941 = n822 ^ n28 ^ 1'b0 ;
  assign n942 = n181 | n941 ;
  assign n943 = n384 | n942 ;
  assign n944 = n873 & ~n943 ;
  assign n945 = n54 & ~n944 ;
  assign n946 = n452 & n945 ;
  assign n947 = n940 & ~n946 ;
  assign n948 = n698 & n947 ;
  assign n949 = n948 ^ n757 ^ 1'b0 ;
  assign n950 = n533 | n641 ;
  assign n951 = n45 | n65 ;
  assign n952 = n98 & ~n951 ;
  assign n953 = n952 ^ n856 ^ 1'b0 ;
  assign n954 = n208 & n953 ;
  assign n955 = ~n420 & n737 ;
  assign n956 = n955 ^ n498 ^ 1'b0 ;
  assign n957 = n956 ^ n645 ^ 1'b0 ;
  assign n958 = n279 & n545 ;
  assign n959 = ~n957 & n958 ;
  assign n960 = x6 & n848 ;
  assign n961 = n169 & n960 ;
  assign n962 = n458 ^ n76 ^ 1'b0 ;
  assign n963 = n138 & ~n962 ;
  assign n964 = n963 ^ n961 ^ 1'b0 ;
  assign n965 = n961 | n964 ;
  assign n966 = n737 | n961 ;
  assign n967 = ~n881 & n966 ;
  assign n968 = n404 | n890 ;
  assign n969 = x6 & n522 ;
  assign n970 = n154 & n969 ;
  assign n971 = ( ~n212 & n503 ) | ( ~n212 & n970 ) | ( n503 & n970 ) ;
  assign n972 = n890 & ~n971 ;
  assign n973 = n746 ^ n422 ^ 1'b0 ;
  assign n974 = n105 & n973 ;
  assign n975 = n525 & ~n796 ;
  assign n976 = n86 & ~n251 ;
  assign n977 = n454 ^ n340 ^ 1'b0 ;
  assign n978 = n418 & ~n977 ;
  assign n979 = ~n47 & n280 ;
  assign n980 = n979 ^ n113 ^ 1'b0 ;
  assign n981 = n980 ^ n809 ^ 1'b0 ;
  assign n982 = n978 & ~n981 ;
  assign n983 = ~n154 & n982 ;
  assign n984 = ~n631 & n983 ;
  assign n985 = n292 & ~n783 ;
  assign n986 = n243 | n690 ;
  assign n987 = n408 & ~n986 ;
  assign n988 = n638 | n987 ;
  assign n989 = ~n86 & n758 ;
  assign n990 = n23 & n872 ;
  assign n991 = ~n171 & n990 ;
  assign n992 = n733 ^ n133 ^ 1'b0 ;
  assign n993 = n991 | n992 ;
  assign n994 = n205 | n880 ;
  assign n995 = n994 ^ n17 ^ 1'b0 ;
  assign n996 = n942 | n995 ;
  assign n997 = n996 ^ n615 ^ n56 ;
  assign n998 = n147 | n997 ;
  assign n999 = ~n130 & n430 ;
  assign n1000 = ~n915 & n999 ;
  assign n1001 = n563 | n584 ;
  assign n1002 = n931 | n1001 ;
  assign n1003 = n1002 ^ n503 ^ 1'b0 ;
  assign n1004 = n441 | n911 ;
  assign n1005 = n227 ^ n222 ^ 1'b0 ;
  assign n1006 = ~n468 & n727 ;
  assign n1007 = n1005 & ~n1006 ;
  assign n1009 = n224 ^ n205 ^ 1'b0 ;
  assign n1008 = n233 & n522 ;
  assign n1010 = n1009 ^ n1008 ^ 1'b0 ;
  assign n1011 = n85 ^ n38 ^ 1'b0 ;
  assign n1012 = n54 & ~n1011 ;
  assign n1013 = ~n420 & n1012 ;
  assign n1014 = n1013 ^ n478 ^ 1'b0 ;
  assign n1015 = n1014 ^ n136 ^ 1'b0 ;
  assign n1016 = ~n873 & n1015 ;
  assign n1017 = ~n667 & n1016 ;
  assign n1018 = n508 & n1017 ;
  assign n1019 = n307 | n552 ;
  assign n1020 = n1018 & ~n1019 ;
  assign n1021 = n1020 ^ n560 ^ 1'b0 ;
  assign n1022 = n223 & n837 ;
  assign n1023 = ~n220 & n1022 ;
  assign n1024 = ( ~n188 & n852 ) | ( ~n188 & n1023 ) | ( n852 & n1023 ) ;
  assign n1025 = n438 & n902 ;
  assign n1026 = n418 ^ n376 ^ 1'b0 ;
  assign n1027 = ~n680 & n1026 ;
  assign n1028 = n388 & ~n395 ;
  assign n1029 = ~n1027 & n1028 ;
  assign n1030 = n40 | n999 ;
  assign n1031 = n1030 ^ n19 ^ 1'b0 ;
  assign n1032 = n474 | n1031 ;
  assign n1033 = n635 ^ n138 ^ 1'b0 ;
  assign n1034 = n309 ^ n154 ^ 1'b0 ;
  assign n1035 = ~n563 & n1034 ;
  assign n1036 = ~n365 & n1035 ;
  assign n1037 = n1036 ^ n808 ^ 1'b0 ;
  assign n1038 = n1033 & n1037 ;
  assign n1039 = ~n422 & n799 ;
  assign n1040 = n1039 ^ n600 ^ 1'b0 ;
  assign n1041 = n317 | n798 ;
  assign n1042 = n1041 ^ n586 ^ 1'b0 ;
  assign n1043 = n130 & ~n442 ;
  assign n1044 = ~n349 & n1043 ;
  assign n1045 = ( ~n641 & n862 ) | ( ~n641 & n1044 ) | ( n862 & n1044 ) ;
  assign n1046 = n200 & n259 ;
  assign n1047 = n1046 ^ n387 ^ 1'b0 ;
  assign n1048 = n432 & n1047 ;
  assign n1049 = n1048 ^ n398 ^ 1'b0 ;
  assign n1050 = ~n110 & n1049 ;
  assign n1051 = n1050 ^ n437 ^ 1'b0 ;
  assign n1052 = ~n468 & n1051 ;
  assign n1053 = x4 & ~n952 ;
  assign n1054 = ~n1052 & n1053 ;
  assign n1055 = n1045 & n1054 ;
  assign n1056 = n1055 ^ n577 ^ n489 ;
  assign n1057 = ~n412 & n877 ;
  assign n1059 = ~n124 & n799 ;
  assign n1060 = n991 & n1059 ;
  assign n1061 = n477 & ~n1060 ;
  assign n1062 = n1061 ^ x8 ^ 1'b0 ;
  assign n1058 = n229 ^ n28 ^ 1'b0 ;
  assign n1063 = n1062 ^ n1058 ^ 1'b0 ;
  assign n1064 = n27 & n465 ;
  assign n1065 = n1064 ^ n919 ^ n417 ;
  assign n1066 = ( n896 & n934 ) | ( n896 & ~n1044 ) | ( n934 & ~n1044 ) ;
  assign n1067 = n331 ^ n146 ^ 1'b0 ;
  assign n1068 = n260 & ~n1067 ;
  assign n1069 = ~n495 & n961 ;
  assign n1070 = n1069 ^ n194 ^ 1'b0 ;
  assign n1071 = n1068 & n1070 ;
  assign n1072 = n131 | n885 ;
  assign n1073 = n421 | n1072 ;
  assign n1074 = n331 & ~n411 ;
  assign n1075 = n1074 ^ n47 ^ 1'b0 ;
  assign n1076 = n1075 ^ n523 ^ 1'b0 ;
  assign n1077 = n260 | n1076 ;
  assign n1078 = n854 ^ n371 ^ n326 ;
  assign n1079 = n508 ^ n401 ^ n132 ;
  assign n1080 = n511 | n1079 ;
  assign n1081 = n1080 ^ n749 ^ 1'b0 ;
  assign n1082 = n305 | n1081 ;
  assign n1083 = n1082 ^ n490 ^ 1'b0 ;
  assign n1084 = n199 & ~n325 ;
  assign n1085 = ~n212 & n1084 ;
  assign n1086 = n631 & n737 ;
  assign n1087 = n454 & n1086 ;
  assign n1088 = n875 ^ n155 ^ 1'b0 ;
  assign n1089 = n390 | n1088 ;
  assign n1090 = ~n452 & n687 ;
  assign n1091 = n100 | n889 ;
  assign n1092 = n898 | n1091 ;
  assign n1093 = ~n328 & n1092 ;
  assign n1094 = ~n709 & n1093 ;
  assign n1095 = n1033 ^ n297 ^ 1'b0 ;
  assign n1101 = n124 & ~n431 ;
  assign n1102 = n1052 & ~n1101 ;
  assign n1103 = n1102 ^ n54 ^ 1'b0 ;
  assign n1098 = n539 ^ x0 ^ 1'b0 ;
  assign n1099 = n239 & ~n1098 ;
  assign n1096 = n360 & ~n767 ;
  assign n1097 = x0 & ~n1096 ;
  assign n1100 = n1099 ^ n1097 ^ 1'b0 ;
  assign n1104 = n1103 ^ n1100 ^ n271 ;
  assign n1105 = n451 & n1045 ;
  assign n1106 = n204 ^ n43 ^ 1'b0 ;
  assign n1107 = n30 & ~n1106 ;
  assign n1108 = ~n312 & n1107 ;
  assign n1109 = ~n61 & n1108 ;
  assign n1110 = n793 & ~n1054 ;
  assign n1111 = n1109 | n1110 ;
  assign n1112 = n56 & n765 ;
  assign n1113 = ~n1060 & n1112 ;
  assign n1114 = n1113 ^ n851 ^ 1'b0 ;
  assign n1115 = n942 ^ n659 ^ 1'b0 ;
  assign n1116 = ~n459 & n1115 ;
  assign n1117 = n1031 ^ n766 ^ n675 ;
  assign n1118 = n456 & n1117 ;
  assign n1119 = ~x5 & n167 ;
  assign n1120 = n1119 ^ n131 ^ 1'b0 ;
  assign n1121 = n212 & ~n1120 ;
  assign n1122 = ( n584 & ~n710 ) | ( n584 & n957 ) | ( ~n710 & n957 ) ;
  assign n1123 = n195 & ~n1122 ;
  assign n1124 = ~n23 & n327 ;
  assign n1125 = n619 ^ n606 ^ 1'b0 ;
  assign n1126 = n85 | n1125 ;
  assign n1127 = n1126 ^ n133 ^ 1'b0 ;
  assign n1128 = n25 & n1127 ;
  assign n1129 = n205 | n326 ;
  assign n1130 = n1033 | n1129 ;
  assign n1131 = n257 | n277 ;
  assign n1132 = n343 | n559 ;
  assign n1133 = n1132 ^ n363 ^ 1'b0 ;
  assign n1134 = n409 & n1133 ;
  assign n1135 = n673 ^ n582 ^ 1'b0 ;
  assign n1136 = n404 | n1135 ;
  assign n1139 = ~n251 & n600 ;
  assign n1140 = n1139 ^ n255 ^ 1'b0 ;
  assign n1137 = n270 & n380 ;
  assign n1138 = n1137 ^ n44 ^ 1'b0 ;
  assign n1141 = n1140 ^ n1138 ^ 1'b0 ;
  assign n1142 = n279 & n841 ;
  assign n1143 = n902 ^ n588 ^ 1'b0 ;
  assign n1144 = n1142 & n1143 ;
  assign n1145 = n423 ^ n86 ^ n56 ;
  assign n1146 = n852 ^ n437 ^ 1'b0 ;
  assign n1147 = n1146 ^ n360 ^ 1'b0 ;
  assign n1148 = n25 & n189 ;
  assign n1149 = n1148 ^ n695 ^ 1'b0 ;
  assign n1150 = ~n1147 & n1149 ;
  assign n1151 = ~n149 & n227 ;
  assign n1152 = n1151 ^ n228 ^ 1'b0 ;
  assign n1153 = n1152 ^ n579 ^ 1'b0 ;
  assign n1154 = n1150 & n1153 ;
  assign n1155 = n20 & n765 ;
  assign n1156 = n685 | n1155 ;
  assign n1157 = n1156 ^ n113 ^ 1'b0 ;
  assign n1158 = n129 & n406 ;
  assign n1159 = ~n320 & n1158 ;
  assign n1160 = n1159 ^ n851 ^ 1'b0 ;
  assign n1161 = n249 & n1160 ;
  assign n1162 = n226 ^ n115 ^ 1'b0 ;
  assign n1163 = n536 & ~n1162 ;
  assign n1164 = n661 ^ n623 ^ n47 ;
  assign n1165 = n1163 & ~n1164 ;
  assign n1166 = n91 & n1027 ;
  assign n1167 = n1096 & n1166 ;
  assign n1168 = n446 ^ n26 ^ 1'b0 ;
  assign n1169 = n27 & ~n1168 ;
  assign n1170 = ( n253 & n317 ) | ( n253 & ~n1169 ) | ( n317 & ~n1169 ) ;
  assign n1171 = n147 & ~n1170 ;
  assign n1172 = n1171 ^ n452 ^ 1'b0 ;
  assign n1173 = n447 & ~n1172 ;
  assign n1174 = n113 | n548 ;
  assign n1175 = n133 | n140 ;
  assign n1176 = n243 & ~n1175 ;
  assign n1177 = n1174 & ~n1176 ;
  assign n1178 = n301 & n1068 ;
  assign n1179 = n406 & n1178 ;
  assign n1180 = n181 ^ n27 ^ 1'b0 ;
  assign n1181 = n20 | n1180 ;
  assign n1182 = n23 & n94 ;
  assign n1183 = n1181 | n1182 ;
  assign n1184 = n1183 ^ n541 ^ 1'b0 ;
  assign n1185 = ~n533 & n1184 ;
  assign n1186 = n1138 & n1185 ;
  assign n1187 = n395 ^ n365 ^ 1'b0 ;
  assign n1188 = ~n539 & n712 ;
  assign n1189 = ~n73 & n1188 ;
  assign n1190 = n1187 & n1189 ;
  assign n1191 = ( n164 & n345 ) | ( n164 & n372 ) | ( n345 & n372 ) ;
  assign n1192 = n1191 ^ n716 ^ 1'b0 ;
  assign n1193 = ~n586 & n608 ;
  assign n1194 = n1193 ^ n275 ^ 1'b0 ;
  assign n1195 = ~n390 & n931 ;
  assign n1196 = ~n1194 & n1195 ;
  assign n1197 = x1 & n885 ;
  assign n1198 = n590 & n1197 ;
  assign n1199 = n132 | n1198 ;
  assign n1203 = n160 & n494 ;
  assign n1204 = n1203 ^ n224 ^ 1'b0 ;
  assign n1201 = n229 ^ n51 ^ 1'b0 ;
  assign n1202 = ( x0 & n47 ) | ( x0 & n1201 ) | ( n47 & n1201 ) ;
  assign n1205 = n1204 ^ n1202 ^ n318 ;
  assign n1206 = n1012 & ~n1205 ;
  assign n1207 = n393 & n1206 ;
  assign n1200 = n592 & n1092 ;
  assign n1208 = n1207 ^ n1200 ^ n392 ;
  assign n1209 = ~n13 & n76 ;
  assign n1210 = n1208 & n1209 ;
  assign n1211 = n110 & n315 ;
  assign n1212 = n695 & ~n889 ;
  assign n1213 = n1212 ^ n696 ^ n79 ;
  assign n1214 = ~n248 & n655 ;
  assign n1215 = ~n521 & n1214 ;
  assign n1216 = ( n325 & n354 ) | ( n325 & n598 ) | ( n354 & n598 ) ;
  assign n1222 = ~n420 & n868 ;
  assign n1223 = n85 & n1222 ;
  assign n1220 = n116 | n347 ;
  assign n1221 = n44 | n1220 ;
  assign n1224 = n1223 ^ n1221 ^ 1'b0 ;
  assign n1217 = n844 ^ n233 ^ 1'b0 ;
  assign n1218 = n1217 ^ n1020 ^ 1'b0 ;
  assign n1219 = n57 & ~n1218 ;
  assign n1225 = n1224 ^ n1219 ^ 1'b0 ;
  assign n1226 = n598 & ~n1225 ;
  assign n1227 = ~n286 & n868 ;
  assign n1228 = ~n497 & n983 ;
  assign n1229 = ~n43 & n1228 ;
  assign n1230 = n1229 ^ n733 ^ n492 ;
  assign n1231 = n694 | n1014 ;
  assign n1232 = n372 | n890 ;
  assign n1233 = n150 & ~n1232 ;
  assign n1234 = n1233 ^ n17 ^ 1'b0 ;
  assign n1235 = ~x9 & n898 ;
  assign n1236 = n1235 ^ n315 ^ 1'b0 ;
  assign n1237 = n452 | n1236 ;
  assign n1238 = n472 & n1199 ;
  assign n1239 = n845 & n1130 ;
  assign n1240 = n1239 ^ n208 ^ 1'b0 ;
  assign n1241 = ~n1231 & n1240 ;
  assign n1242 = n305 | n637 ;
  assign n1243 = n1242 ^ n439 ^ 1'b0 ;
  assign n1244 = n657 & ~n829 ;
  assign n1245 = n1148 | n1244 ;
  assign n1246 = ( ~n181 & n543 ) | ( ~n181 & n732 ) | ( n543 & n732 ) ;
  assign n1247 = n1246 ^ n160 ^ 1'b0 ;
  assign n1248 = ~n219 & n269 ;
  assign n1249 = n1248 ^ n855 ^ 1'b0 ;
  assign n1250 = n362 | n1249 ;
  assign n1251 = n387 & ~n1250 ;
  assign n1252 = ~n602 & n1217 ;
  assign n1253 = ~n260 & n1252 ;
  assign n1254 = n1253 ^ n1186 ^ 1'b0 ;
  assign n1257 = n19 | n497 ;
  assign n1255 = ~n307 & n707 ;
  assign n1256 = n1255 ^ n140 ^ 1'b0 ;
  assign n1258 = n1257 ^ n1256 ^ n167 ;
  assign n1259 = n49 & n527 ;
  assign n1260 = ~n1258 & n1259 ;
  assign n1261 = n1260 ^ n973 ^ 1'b0 ;
  assign n1262 = n738 & n961 ;
  assign n1263 = n746 ^ n452 ^ 1'b0 ;
  assign n1264 = ( ~n703 & n1262 ) | ( ~n703 & n1263 ) | ( n1262 & n1263 ) ;
  assign n1265 = n732 ^ n404 ^ 1'b0 ;
  assign n1266 = ~n49 & n1265 ;
  assign n1267 = n13 | n28 ;
  assign n1268 = n188 ^ x8 ^ 1'b0 ;
  assign n1269 = n1055 & ~n1268 ;
  assign n1270 = ~n727 & n924 ;
  assign n1271 = ~n36 & n1270 ;
  assign n1274 = n568 ^ n227 ^ 1'b0 ;
  assign n1275 = n339 & n1274 ;
  assign n1272 = n999 ^ n170 ^ 1'b0 ;
  assign n1273 = n749 | n1272 ;
  assign n1276 = n1275 ^ n1273 ^ 1'b0 ;
  assign n1277 = n564 ^ n269 ^ 1'b0 ;
  assign n1278 = n1033 & ~n1277 ;
  assign n1279 = n459 & ~n663 ;
  assign n1280 = n1279 ^ n826 ^ 1'b0 ;
  assign n1281 = n1278 & ~n1280 ;
  assign n1282 = n1281 ^ n825 ^ 1'b0 ;
  assign n1283 = n451 & n1282 ;
  assign n1284 = n132 | n1241 ;
  assign n1285 = n890 & ~n1191 ;
  assign n1286 = n475 & ~n582 ;
  assign n1287 = n1286 ^ n547 ^ 1'b0 ;
  assign n1288 = n223 & ~n1287 ;
  assign n1289 = n1285 & n1288 ;
  assign n1290 = n796 & n1289 ;
  assign n1291 = ~n503 & n1290 ;
  assign n1292 = n487 ^ n384 ^ 1'b0 ;
  assign n1293 = n673 & n1292 ;
  assign n1294 = n1293 ^ n229 ^ 1'b0 ;
  assign n1295 = n312 | n1294 ;
  assign n1296 = n220 & ~n1295 ;
  assign n1297 = n1296 ^ n304 ^ 1'b0 ;
  assign n1298 = n163 & n365 ;
  assign n1299 = n1298 ^ n983 ^ n568 ;
  assign n1300 = ~n226 & n257 ;
  assign n1301 = n310 & n625 ;
  assign n1303 = n619 ^ n35 ^ 1'b0 ;
  assign n1304 = ~n480 & n1303 ;
  assign n1302 = x6 & ~n993 ;
  assign n1305 = n1304 ^ n1302 ^ 1'b0 ;
  assign n1306 = n1235 ^ n316 ^ 1'b0 ;
  assign n1307 = n1306 ^ n73 ^ 1'b0 ;
  assign n1308 = n248 ^ n119 ^ 1'b0 ;
  assign n1309 = n205 | n1062 ;
  assign n1310 = x6 | n1309 ;
  assign n1311 = ~n250 & n489 ;
  assign n1312 = n1311 ^ n518 ^ 1'b0 ;
  assign n1313 = n1047 & ~n1312 ;
  assign n1314 = n220 & ~n1229 ;
  assign n1315 = n1314 ^ n254 ^ 1'b0 ;
  assign n1316 = ~n431 & n809 ;
  assign n1317 = n160 & ~n461 ;
  assign n1318 = n1317 ^ n195 ^ 1'b0 ;
  assign n1319 = ~n260 & n1318 ;
  assign n1320 = n1319 ^ n905 ^ 1'b0 ;
  assign n1321 = ( n288 & n530 ) | ( n288 & n855 ) | ( n530 & n855 ) ;
  assign n1322 = ~n135 & n508 ;
  assign n1323 = n494 ^ n67 ^ 1'b0 ;
  assign n1325 = ~n226 & n379 ;
  assign n1324 = ~n136 & n688 ;
  assign n1326 = n1325 ^ n1324 ^ 1'b0 ;
  assign n1327 = ~n27 & n339 ;
  assign n1328 = n1327 ^ n199 ^ 1'b0 ;
  assign n1329 = x2 & ~n1328 ;
  assign n1330 = ~n459 & n849 ;
  assign n1331 = n47 & n1330 ;
  assign n1333 = n25 & n222 ;
  assign n1334 = n1333 ^ n723 ^ 1'b0 ;
  assign n1332 = n54 & ~n135 ;
  assign n1335 = n1334 ^ n1332 ^ 1'b0 ;
  assign n1336 = n892 & n1014 ;
  assign n1337 = n1023 & n1336 ;
  assign n1338 = n983 ^ n214 ^ 1'b0 ;
  assign n1339 = ~n390 & n1338 ;
  assign n1340 = n1339 ^ n487 ^ 1'b0 ;
  assign n1341 = n441 & n873 ;
  assign n1342 = n783 & n1341 ;
  assign n1343 = n746 ^ n26 ^ 1'b0 ;
  assign n1344 = n1343 ^ n1107 ^ 1'b0 ;
  assign n1345 = n488 ^ n315 ^ 1'b0 ;
  assign n1346 = ~n107 & n1184 ;
  assign n1347 = n344 ^ n57 ^ 1'b0 ;
  assign n1348 = ~n468 & n1025 ;
  assign n1349 = ~n1347 & n1348 ;
  assign n1351 = n369 ^ n246 ^ n160 ;
  assign n1350 = ~n159 & n974 ;
  assign n1352 = n1351 ^ n1350 ^ 1'b0 ;
  assign n1353 = n649 ^ n103 ^ 1'b0 ;
  assign n1354 = n471 ^ n183 ^ 1'b0 ;
  assign n1355 = n40 & ~n1354 ;
  assign n1356 = n517 ^ n197 ^ 1'b0 ;
  assign n1357 = n707 ^ n448 ^ 1'b0 ;
  assign n1358 = n1356 | n1357 ;
  assign n1359 = n1358 ^ n905 ^ 1'b0 ;
  assign n1360 = n835 & n1359 ;
  assign n1361 = n988 ^ n511 ^ 1'b0 ;
  assign n1362 = x9 & ~n952 ;
  assign n1363 = n1362 ^ n322 ^ 1'b0 ;
  assign n1364 = ~n851 & n1363 ;
  assign n1365 = n1364 ^ n456 ^ 1'b0 ;
  assign n1366 = n765 ^ n392 ^ 1'b0 ;
  assign n1367 = n1366 ^ n49 ^ 1'b0 ;
  assign n1368 = n938 | n1367 ;
  assign n1369 = n1123 & ~n1368 ;
  assign n1370 = ( n582 & n745 ) | ( n582 & ~n1369 ) | ( n745 & ~n1369 ) ;
  assign n1371 = n825 ^ n712 ^ n58 ;
  assign n1372 = n685 & n1371 ;
  assign n1373 = n592 | n1031 ;
  assign n1374 = n1373 ^ n983 ^ 1'b0 ;
  assign n1375 = x3 & n1374 ;
  assign n1376 = n890 & n1375 ;
  assign n1377 = n1376 ^ n861 ^ 1'b0 ;
  assign n1378 = n931 ^ n173 ^ 1'b0 ;
  assign n1379 = ~n867 & n1378 ;
  assign n1380 = n720 | n1207 ;
  assign n1381 = n910 & ~n1380 ;
  assign n1382 = n270 & ~n617 ;
  assign n1383 = n1336 & ~n1382 ;
  assign n1384 = ~n1131 & n1383 ;
  assign n1385 = n1384 ^ n86 ^ 1'b0 ;
  assign n1386 = n1142 ^ n224 ^ 1'b0 ;
  assign n1387 = n286 | n880 ;
  assign n1388 = n1387 ^ n1194 ^ 1'b0 ;
  assign n1389 = n720 | n1388 ;
  assign n1390 = n453 & n1389 ;
  assign n1391 = n432 ^ n212 ^ n199 ;
  assign n1392 = n331 | n541 ;
  assign n1393 = n502 & ~n1392 ;
  assign n1394 = n1393 ^ n854 ^ 1'b0 ;
  assign n1395 = ( n100 & n1391 ) | ( n100 & n1394 ) | ( n1391 & n1394 ) ;
  assign n1396 = n1194 ^ n311 ^ 1'b0 ;
  assign n1397 = n1396 ^ n1012 ^ 1'b0 ;
  assign n1398 = n1271 | n1397 ;
  assign n1399 = n1251 | n1369 ;
  assign n1400 = x6 | n1399 ;
  assign n1401 = n861 ^ n825 ^ n356 ;
  assign n1402 = ~n851 & n1401 ;
  assign n1403 = n1402 ^ n376 ^ 1'b0 ;
  assign n1406 = ~n250 & n513 ;
  assign n1407 = n1406 ^ n466 ^ 1'b0 ;
  assign n1408 = n741 & ~n1407 ;
  assign n1404 = n527 & n936 ;
  assign n1405 = ~n820 & n1404 ;
  assign n1409 = n1408 ^ n1405 ^ 1'b0 ;
  assign n1410 = n989 ^ n796 ^ n339 ;
  assign n1411 = n328 & n1389 ;
  assign n1414 = n28 & ~n173 ;
  assign n1415 = n547 ^ n244 ^ 1'b0 ;
  assign n1416 = n1414 & ~n1415 ;
  assign n1412 = ~n149 & n434 ;
  assign n1413 = n360 & n1412 ;
  assign n1417 = n1416 ^ n1413 ^ 1'b0 ;
  assign n1418 = n65 | n1417 ;
  assign n1419 = n1109 ^ n311 ^ 1'b0 ;
  assign n1420 = n226 & ~n1161 ;
  assign n1421 = n608 & ~n663 ;
  assign n1422 = n1421 ^ n564 ^ 1'b0 ;
  assign n1423 = ~n344 & n1422 ;
  assign n1424 = n1420 & n1423 ;
  assign n1425 = n139 | n778 ;
  assign n1426 = n1425 ^ n1356 ^ n26 ;
  assign n1427 = n1267 ^ n241 ^ 1'b0 ;
  assign n1428 = n1038 & ~n1427 ;
  assign n1429 = n668 ^ n542 ^ 1'b0 ;
  assign n1430 = n1429 ^ n890 ^ 1'b0 ;
  assign n1434 = n533 ^ n239 ^ 1'b0 ;
  assign n1431 = n776 ^ n30 ^ 1'b0 ;
  assign n1432 = ( n323 & n956 ) | ( n323 & ~n993 ) | ( n956 & ~n993 ) ;
  assign n1433 = n1431 & ~n1432 ;
  assign n1435 = n1434 ^ n1433 ^ 1'b0 ;
  assign n1436 = n259 & n440 ;
  assign n1437 = n1436 ^ n967 ^ n251 ;
  assign n1438 = n1343 ^ n901 ^ n849 ;
  assign n1439 = n1438 ^ n67 ^ 1'b0 ;
  assign n1440 = n681 & n1152 ;
  assign n1441 = n1440 ^ n160 ^ 1'b0 ;
  assign n1442 = n508 | n1441 ;
  assign n1443 = n926 ^ n304 ^ 1'b0 ;
  assign n1444 = ~n1029 & n1443 ;
  assign n1445 = ~n517 & n1444 ;
  assign n1447 = n218 | n905 ;
  assign n1448 = n1447 ^ n261 ^ 1'b0 ;
  assign n1449 = ( ~n119 & n159 ) | ( ~n119 & n1448 ) | ( n159 & n1448 ) ;
  assign n1450 = n1449 ^ n1256 ^ 1'b0 ;
  assign n1446 = n1105 ^ n862 ^ 1'b0 ;
  assign n1451 = n1450 ^ n1446 ^ n199 ;
  assign n1452 = n1077 ^ n890 ^ 1'b0 ;
  assign n1453 = n600 & n1452 ;
  assign n1454 = n36 & ~n898 ;
  assign n1455 = ~n280 & n1033 ;
  assign n1456 = n358 & ~n661 ;
  assign n1457 = n1456 ^ n793 ^ 1'b0 ;
  assign n1458 = n402 & n1457 ;
  assign n1459 = ( n322 & n991 ) | ( n322 & n1458 ) | ( n991 & n1458 ) ;
  assign n1460 = n1198 & ~n1459 ;
  assign n1461 = n1455 | n1460 ;
  assign n1462 = n304 | n1152 ;
  assign n1463 = n889 ^ n766 ^ 1'b0 ;
  assign n1464 = n513 & ~n1463 ;
  assign n1467 = ~n357 & n645 ;
  assign n1465 = n296 & n1414 ;
  assign n1466 = ~n889 & n1465 ;
  assign n1468 = n1467 ^ n1466 ^ 1'b0 ;
  assign n1469 = n1464 & n1468 ;
  assign n1475 = n498 & ~n510 ;
  assign n1476 = n1475 ^ n189 ^ 1'b0 ;
  assign n1470 = n169 ^ x6 ^ 1'b0 ;
  assign n1471 = n265 | n1470 ;
  assign n1472 = n219 | n714 ;
  assign n1473 = n1472 ^ n880 ^ 1'b0 ;
  assign n1474 = n1471 | n1473 ;
  assign n1477 = n1476 ^ n1474 ^ 1'b0 ;
  assign n1478 = ~n330 & n1277 ;
  assign n1479 = n1478 ^ n667 ^ 1'b0 ;
  assign n1480 = n1479 ^ n1023 ^ n257 ;
  assign n1481 = ( ~n374 & n1477 ) | ( ~n374 & n1480 ) | ( n1477 & n1480 ) ;
  assign n1482 = n600 ^ n314 ^ 1'b0 ;
  assign n1483 = n417 | n1482 ;
  assign n1484 = n1483 ^ n785 ^ 1'b0 ;
  assign n1485 = ~n1202 & n1425 ;
  assign n1486 = n221 ^ n132 ^ 1'b0 ;
  assign n1487 = n126 & n1052 ;
  assign n1488 = ~n1005 & n1487 ;
  assign n1489 = n1486 & ~n1488 ;
  assign n1490 = n805 & n1489 ;
  assign n1491 = n1490 ^ n840 ^ 1'b0 ;
  assign n1492 = n857 ^ n231 ^ 1'b0 ;
  assign n1493 = n602 | n1492 ;
  assign n1494 = n588 | n667 ;
  assign n1495 = n1004 | n1494 ;
  assign n1496 = n1495 ^ n1409 ^ 1'b0 ;
  assign n1497 = ~n1493 & n1496 ;
  assign n1498 = n833 & n1322 ;
  assign n1499 = n1498 ^ n873 ^ 1'b0 ;
  assign n1500 = n1271 ^ n527 ^ 1'b0 ;
  assign n1501 = n28 | n1500 ;
  assign n1502 = n1080 & n1320 ;
  assign n1503 = ~n56 & n470 ;
  assign n1504 = n1503 ^ n286 ^ 1'b0 ;
  assign n1505 = n703 ^ n320 ^ 1'b0 ;
  assign n1506 = n1024 & ~n1173 ;
  assign n1507 = n382 & n1466 ;
  assign n1509 = n944 ^ n584 ^ 1'b0 ;
  assign n1510 = n1336 & n1509 ;
  assign n1508 = n312 ^ n304 ^ 1'b0 ;
  assign n1511 = n1510 ^ n1508 ^ n451 ;
  assign n1512 = n110 | n565 ;
  assign n1513 = n478 | n1512 ;
  assign n1514 = n637 ^ n209 ^ 1'b0 ;
  assign n1515 = n721 & ~n808 ;
  assign n1516 = n1515 ^ n1244 ^ 1'b0 ;
  assign n1517 = n262 | n1192 ;
  assign n1518 = ( ~n133 & n323 ) | ( ~n133 & n675 ) | ( n323 & n675 ) ;
  assign n1519 = ~n944 & n1518 ;
  assign n1520 = n1519 ^ n1338 ^ 1'b0 ;
  assign n1521 = ( n452 & ~n463 ) | ( n452 & n648 ) | ( ~n463 & n648 ) ;
  assign n1522 = n1521 ^ x6 ^ 1'b0 ;
  assign n1523 = n1414 ^ n1087 ^ n822 ;
  assign n1524 = n207 | n1523 ;
  assign n1525 = n821 | n1524 ;
  assign n1526 = n197 ^ n40 ^ 1'b0 ;
  assign n1527 = n1300 & n1526 ;
  assign n1528 = n1527 ^ n597 ^ 1'b0 ;
  assign n1529 = n792 | n880 ;
  assign n1530 = n231 | n1529 ;
  assign n1531 = n826 & ~n1530 ;
  assign n1533 = n931 ^ n468 ^ 1'b0 ;
  assign n1534 = n688 & ~n1533 ;
  assign n1532 = n1345 & n1460 ;
  assign n1535 = n1534 ^ n1532 ^ 1'b0 ;
  assign n1536 = n765 ^ n139 ^ 1'b0 ;
  assign n1537 = n541 | n1536 ;
  assign n1538 = n265 & ~n1537 ;
  assign n1539 = n96 & n806 ;
  assign n1543 = n105 & n430 ;
  assign n1544 = ( n165 & n630 ) | ( n165 & n1543 ) | ( n630 & n1543 ) ;
  assign n1545 = n1544 ^ n1334 ^ n138 ;
  assign n1540 = n456 & ~n564 ;
  assign n1541 = ~n459 & n1540 ;
  assign n1542 = n296 & n1541 ;
  assign n1546 = n1545 ^ n1542 ^ n851 ;
  assign n1547 = ~n750 & n1546 ;
  assign n1548 = n1547 ^ n1403 ^ 1'b0 ;
  assign n1551 = n152 & n331 ;
  assign n1549 = n727 | n1201 ;
  assign n1550 = n1549 ^ n488 ^ 1'b0 ;
  assign n1552 = n1551 ^ n1550 ^ 1'b0 ;
  assign n1553 = n136 & ~n970 ;
  assign n1554 = ( n592 & n908 ) | ( n592 & ~n1553 ) | ( n908 & ~n1553 ) ;
  assign n1555 = n1554 ^ n48 ^ 1'b0 ;
  assign n1556 = n403 | n1555 ;
  assign n1557 = n1554 ^ n121 ^ 1'b0 ;
  assign n1558 = ~n1556 & n1557 ;
  assign n1559 = n235 & n848 ;
  assign n1560 = ~n1558 & n1559 ;
  assign n1561 = n17 | n169 ;
  assign n1562 = n125 | n1035 ;
  assign n1563 = n896 | n1562 ;
  assign n1564 = ( n200 & n673 ) | ( n200 & n709 ) | ( n673 & n709 ) ;
  assign n1565 = ~n411 & n835 ;
  assign n1566 = ~n1564 & n1565 ;
  assign n1567 = n1566 ^ n996 ^ 1'b0 ;
  assign n1568 = n1387 ^ n717 ^ 1'b0 ;
  assign n1569 = n1568 ^ n1201 ^ 1'b0 ;
  assign n1570 = ~n344 & n1569 ;
  assign n1571 = n799 & ~n1570 ;
  assign n1572 = ~n1049 & n1134 ;
  assign n1573 = n1571 & n1572 ;
  assign n1574 = n164 & ~n423 ;
  assign n1575 = n1574 ^ n1301 ^ 1'b0 ;
  assign n1576 = ~n997 & n1575 ;
  assign n1577 = ~n1103 & n1335 ;
  assign n1578 = n1577 ^ n1170 ^ 1'b0 ;
  assign n1579 = n241 & ~n1040 ;
  assign n1580 = n1579 ^ n887 ^ 1'b0 ;
  assign n1581 = ~n1186 & n1580 ;
  assign n1582 = n1581 ^ n813 ^ 1'b0 ;
  assign n1583 = n25 & ~n356 ;
  assign n1584 = n1583 ^ n222 ^ 1'b0 ;
  assign n1585 = n27 & ~n551 ;
  assign n1586 = n1584 & n1585 ;
  assign n1587 = n865 ^ n600 ^ 1'b0 ;
  assign n1588 = ~n463 & n1587 ;
  assign n1589 = n690 & n1588 ;
  assign n1590 = ( n452 & ~n1586 ) | ( n452 & n1589 ) | ( ~n1586 & n1589 ) ;
  assign n1591 = ( n1123 & ~n1582 ) | ( n1123 & n1590 ) | ( ~n1582 & n1590 ) ;
  assign n1592 = x1 | n263 ;
  assign n1593 = n647 & n1592 ;
  assign n1594 = ~n1172 & n1593 ;
  assign n1595 = n1004 & n1550 ;
  assign n1596 = n1595 ^ n1329 ^ 1'b0 ;
  assign n1597 = n768 | n1596 ;
  assign n1598 = n1597 ^ n133 ^ 1'b0 ;
  assign n1599 = n1395 ^ n817 ^ 1'b0 ;
  assign n1600 = n360 | n892 ;
  assign n1601 = n1600 ^ n720 ^ 1'b0 ;
  assign n1602 = n557 & n1601 ;
  assign n1603 = n1602 ^ n131 ^ 1'b0 ;
  assign n1604 = n1420 ^ n318 ^ 1'b0 ;
  assign n1605 = n1163 & ~n1604 ;
  assign n1606 = n676 ^ n169 ^ 1'b0 ;
  assign n1607 = ~n1189 & n1606 ;
  assign n1608 = n1109 | n1607 ;
  assign n1609 = n619 ^ n344 ^ 1'b0 ;
  assign n1610 = n1024 | n1083 ;
  assign n1611 = n1610 ^ n856 ^ 1'b0 ;
  assign n1612 = ~n207 & n451 ;
  assign n1613 = n1612 ^ n290 ^ 1'b0 ;
  assign n1614 = n765 ^ n454 ^ 1'b0 ;
  assign n1615 = n1613 | n1614 ;
  assign n1616 = n1142 & ~n1615 ;
  assign n1617 = n1616 ^ n204 ^ 1'b0 ;
  assign n1618 = n1617 ^ n1196 ^ n266 ;
  assign n1619 = n517 ^ x9 ^ 1'b0 ;
  assign n1620 = ~n683 & n1619 ;
  assign n1621 = n535 ^ n277 ^ 1'b0 ;
  assign n1622 = n148 | n1621 ;
  assign n1623 = ( n15 & n1241 ) | ( n15 & ~n1622 ) | ( n1241 & ~n1622 ) ;
  assign n1624 = n1623 ^ n1004 ^ 1'b0 ;
  assign n1625 = n751 ^ n376 ^ 1'b0 ;
  assign n1626 = ~n234 & n1578 ;
  assign n1627 = n634 & n1626 ;
  assign n1628 = n106 & ~n1207 ;
  assign n1629 = n1628 ^ n418 ^ 1'b0 ;
  assign n1630 = ~n772 & n1469 ;
  assign n1631 = n1630 ^ n584 ^ 1'b0 ;
  assign n1632 = n1352 ^ n264 ^ 1'b0 ;
  assign n1633 = ~n1466 & n1632 ;
  assign n1634 = n1633 ^ x0 ^ 1'b0 ;
  assign n1635 = ~n19 & n1634 ;
  assign n1636 = ( n61 & n528 ) | ( n61 & ~n959 ) | ( n528 & ~n959 ) ;
  assign n1637 = n1205 ^ n815 ^ 1'b0 ;
  assign n1641 = n463 ^ n440 ^ 1'b0 ;
  assign n1642 = n1641 ^ n997 ^ 1'b0 ;
  assign n1643 = n475 | n1642 ;
  assign n1644 = n1262 & n1643 ;
  assign n1645 = n1542 ^ n870 ^ 1'b0 ;
  assign n1646 = n842 ^ n74 ^ 1'b0 ;
  assign n1647 = n1645 | n1646 ;
  assign n1648 = ( n611 & ~n1644 ) | ( n611 & n1647 ) | ( ~n1644 & n1647 ) ;
  assign n1638 = n605 & ~n1189 ;
  assign n1639 = ~n170 & n1638 ;
  assign n1640 = n1451 & ~n1639 ;
  assign n1649 = n1648 ^ n1640 ^ 1'b0 ;
  assign n1650 = n780 & n790 ;
  assign n1651 = n61 & n611 ;
  assign n1652 = ~n737 & n1651 ;
  assign n1653 = n511 & ~n1652 ;
  assign n1654 = n669 & ~n1087 ;
  assign n1655 = n26 & n744 ;
  assign n1656 = n302 & n727 ;
  assign n1657 = n380 ^ n188 ^ 1'b0 ;
  assign n1658 = n910 & ~n1289 ;
  assign n1659 = n901 ^ n450 ^ 1'b0 ;
  assign n1660 = n936 | n1615 ;
  assign n1661 = ~n700 & n1660 ;
  assign n1662 = n1553 & n1661 ;
  assign n1663 = n1659 | n1662 ;
  assign n1664 = n820 ^ n722 ^ 1'b0 ;
  assign n1665 = ~n183 & n279 ;
  assign n1666 = n1665 ^ n266 ^ 1'b0 ;
  assign n1667 = n514 | n1666 ;
  assign n1668 = n572 & ~n1110 ;
  assign n1669 = n1667 & ~n1668 ;
  assign n1670 = ~n850 & n1669 ;
  assign n1671 = ~n146 & n1670 ;
  assign n1672 = ~n138 & n1671 ;
  assign n1673 = n608 | n1411 ;
  assign n1674 = n1673 ^ n1563 ^ 1'b0 ;
  assign n1675 = n844 ^ n113 ^ 1'b0 ;
  assign n1676 = n978 & ~n1675 ;
  assign n1677 = ~n1078 & n1676 ;
  assign n1678 = ~n77 & n271 ;
  assign n1679 = n1678 ^ n227 ^ 1'b0 ;
  assign n1680 = n1679 ^ n515 ^ 1'b0 ;
  assign n1681 = n1295 | n1680 ;
  assign n1682 = n768 & ~n1681 ;
  assign n1683 = n1677 | n1682 ;
  assign n1684 = n173 & ~n1683 ;
  assign n1688 = n809 ^ n459 ^ x2 ;
  assign n1685 = n485 | n593 ;
  assign n1686 = n213 | n1685 ;
  assign n1687 = n724 | n1686 ;
  assign n1689 = n1688 ^ n1687 ^ 1'b0 ;
  assign n1690 = n1124 ^ n83 ^ 1'b0 ;
  assign n1691 = ~n567 & n1352 ;
  assign n1692 = n700 | n1584 ;
  assign n1693 = n982 | n1692 ;
  assign n1694 = n470 & ~n1693 ;
  assign n1695 = n1694 ^ n106 ^ 1'b0 ;
  assign n1696 = ~n968 & n1695 ;
  assign n1697 = n1696 ^ n15 ^ 1'b0 ;
  assign n1698 = ~n1315 & n1697 ;
  assign n1699 = n1698 ^ n1267 ^ 1'b0 ;
  assign n1700 = n1483 ^ n861 ^ 1'b0 ;
  assign n1701 = n926 ^ n481 ^ 1'b0 ;
  assign n1702 = n885 ^ n112 ^ 1'b0 ;
  assign n1703 = n802 | n1702 ;
  assign n1704 = n540 | n564 ;
  assign n1705 = n1551 | n1704 ;
  assign n1707 = ( n25 & n73 ) | ( n25 & ~n83 ) | ( n73 & ~n83 ) ;
  assign n1708 = ~n362 & n1707 ;
  assign n1709 = ~n282 & n1708 ;
  assign n1710 = n1709 ^ n509 ^ 1'b0 ;
  assign n1711 = n575 | n1710 ;
  assign n1706 = n492 & n625 ;
  assign n1712 = n1711 ^ n1706 ^ 1'b0 ;
  assign n1713 = n1712 ^ n423 ^ 1'b0 ;
  assign n1714 = n889 | n1713 ;
  assign n1715 = ( ~n976 & n1705 ) | ( ~n976 & n1714 ) | ( n1705 & n1714 ) ;
  assign n1716 = n996 & n1189 ;
  assign n1717 = n1031 ^ n251 ^ 1'b0 ;
  assign n1718 = ~n40 & n978 ;
  assign n1719 = ~n1198 & n1718 ;
  assign n1720 = n1717 & n1719 ;
  assign n1721 = n1460 ^ n1243 ^ 1'b0 ;
  assign n1722 = n875 & ~n971 ;
  assign n1723 = n1722 ^ n414 ^ 1'b0 ;
  assign n1724 = n1121 & ~n1723 ;
  assign n1725 = ~n881 & n1092 ;
  assign n1726 = n817 & n1725 ;
  assign n1727 = n1726 ^ n676 ^ 1'b0 ;
  assign n1728 = n1724 | n1727 ;
  assign n1729 = n1401 ^ n1056 ^ n454 ;
  assign n1730 = n956 ^ n163 ^ 1'b0 ;
  assign n1731 = ~n588 & n1730 ;
  assign n1732 = n163 & ~n384 ;
  assign n1733 = n1732 ^ n936 ^ 1'b0 ;
  assign n1734 = n673 & n1733 ;
  assign n1735 = n1347 & n1734 ;
  assign n1736 = n265 & n1735 ;
  assign n1737 = n1731 & ~n1736 ;
  assign n1738 = n1622 & n1737 ;
  assign n1739 = ( n1094 & n1627 ) | ( n1094 & ~n1738 ) | ( n1627 & ~n1738 ) ;
  assign n1740 = n1476 ^ n738 ^ n228 ;
  assign n1741 = ( n49 & n1627 ) | ( n49 & n1740 ) | ( n1627 & n1740 ) ;
  assign n1742 = n661 | n907 ;
  assign n1743 = n487 & n1742 ;
  assign n1744 = n340 & ~n600 ;
  assign n1745 = n527 ^ n49 ^ 1'b0 ;
  assign n1746 = ~n1744 & n1745 ;
  assign n1747 = n1746 ^ n683 ^ 1'b0 ;
  assign n1748 = ~n1586 & n1747 ;
  assign n1749 = ~n167 & n1748 ;
  assign n1750 = n1064 ^ n931 ^ 1'b0 ;
  assign n1751 = n1750 ^ n459 ^ 1'b0 ;
  assign n1752 = n439 & ~n1751 ;
  assign n1753 = n884 ^ n26 ^ 1'b0 ;
  assign n1754 = ~n541 & n823 ;
  assign n1755 = n1286 & n1754 ;
  assign n1756 = n1755 ^ n801 ^ n340 ;
  assign n1757 = n1753 | n1756 ;
  assign n1758 = n347 & ~n1757 ;
  assign n1759 = n251 | n439 ;
  assign n1760 = n839 & ~n1759 ;
  assign n1761 = n890 ^ n765 ^ 1'b0 ;
  assign n1762 = n1761 ^ n877 ^ 1'b0 ;
  assign n1763 = n515 | n1762 ;
  assign n1764 = n1392 | n1763 ;
  assign n1765 = ( n167 & n732 ) | ( n167 & ~n835 ) | ( n732 & ~n835 ) ;
  assign n1766 = n1707 ^ n96 ^ 1'b0 ;
  assign n1767 = n919 & n1766 ;
  assign n1768 = n1767 ^ n439 ^ 1'b0 ;
  assign n1769 = n1768 ^ n688 ^ 1'b0 ;
  assign n1770 = n1331 ^ n949 ^ 1'b0 ;
  assign n1771 = n968 & n1770 ;
  assign n1772 = ~n1182 & n1265 ;
  assign n1773 = ~n40 & n1052 ;
  assign n1774 = ~n950 & n1773 ;
  assign n1775 = ( n263 & n1772 ) | ( n263 & n1774 ) | ( n1772 & n1774 ) ;
  assign n1777 = n717 ^ n408 ^ 1'b0 ;
  assign n1778 = ~n1568 & n1777 ;
  assign n1776 = ~n297 & n760 ;
  assign n1779 = n1778 ^ n1776 ^ 1'b0 ;
  assign n1780 = n655 & ~n1411 ;
  assign n1781 = n1780 ^ n147 ^ 1'b0 ;
  assign n1782 = n146 ^ n132 ^ 1'b0 ;
  assign n1783 = n642 | n1782 ;
  assign n1785 = ( x9 & n279 ) | ( x9 & ~n635 ) | ( n279 & ~n635 ) ;
  assign n1784 = n625 & n733 ;
  assign n1786 = n1785 ^ n1784 ^ 1'b0 ;
  assign n1787 = n1286 | n1786 ;
  assign n1788 = n800 & ~n1787 ;
  assign n1790 = ~n1476 & n1539 ;
  assign n1789 = n40 & n734 ;
  assign n1791 = n1790 ^ n1789 ^ 1'b0 ;
  assign n1792 = ~n181 & n1111 ;
  assign n1793 = n28 & n351 ;
  assign n1794 = n1793 ^ n129 ^ 1'b0 ;
  assign n1795 = n152 | n1794 ;
  assign n1796 = n1795 ^ n205 ^ 1'b0 ;
  assign n1797 = n1796 ^ n1123 ^ 1'b0 ;
  assign n1798 = n827 & n1797 ;
  assign n1799 = n942 | n1159 ;
  assign n1800 = n1798 | n1799 ;
  assign n1801 = n1385 ^ n539 ^ 1'b0 ;
  assign n1802 = ~n1181 & n1801 ;
  assign n1803 = n855 ^ n546 ^ 1'b0 ;
  assign n1804 = n1803 ^ n703 ^ 1'b0 ;
  assign n1805 = n1551 ^ n365 ^ 1'b0 ;
  assign n1806 = ~n224 & n1805 ;
  assign n1807 = ~n1031 & n1806 ;
  assign n1808 = ~n502 & n1807 ;
  assign n1809 = n49 & ~n1361 ;
  assign n1810 = ~n402 & n765 ;
  assign n1811 = n1810 ^ n1789 ^ 1'b0 ;
  assign n1812 = n619 | n1750 ;
  assign n1813 = n754 | n1812 ;
  assign n1814 = x3 | n1813 ;
  assign n1815 = n1056 & n1394 ;
  assign n1816 = n1815 ^ n403 ^ 1'b0 ;
  assign n1817 = n1707 ^ n112 ^ 1'b0 ;
  assign n1818 = n675 & ~n1817 ;
  assign n1819 = ~n1605 & n1818 ;
  assign n1820 = n1432 ^ n575 ^ 1'b0 ;
  assign n1821 = n1767 & n1820 ;
  assign n1822 = n1821 ^ x6 ^ 1'b0 ;
  assign n1823 = n1409 & n1822 ;
  assign n1824 = n915 ^ n495 ^ 1'b0 ;
  assign n1825 = ~n420 & n1824 ;
  assign n1826 = ~n481 & n605 ;
  assign n1827 = n1826 ^ n1539 ^ 1'b0 ;
  assign n1828 = n1825 & n1827 ;
  assign n1829 = n591 | n1828 ;
  assign n1830 = n1331 ^ n1321 ^ 1'b0 ;
  assign n1831 = n28 | n1744 ;
  assign n1832 = n1831 ^ n93 ^ 1'b0 ;
  assign n1833 = n1655 ^ n1424 ^ 1'b0 ;
  assign n1834 = n239 & n1833 ;
  assign n1835 = n747 ^ n226 ^ 1'b0 ;
  assign n1836 = ~n956 & n1371 ;
  assign n1837 = n1836 ^ n560 ^ 1'b0 ;
  assign n1838 = n26 | n1648 ;
  assign n1839 = n503 ^ n388 ^ 1'b0 ;
  assign n1840 = n1839 ^ n1134 ^ 1'b0 ;
  assign n1841 = n1335 & n1840 ;
  assign n1842 = ~n177 & n1669 ;
  assign n1843 = n1064 ^ n360 ^ 1'b0 ;
  assign n1844 = n902 ^ n192 ^ 1'b0 ;
  assign n1845 = n1843 | n1844 ;
  assign n1846 = n465 ^ n28 ^ 1'b0 ;
  assign n1847 = ~n110 & n1846 ;
  assign n1848 = n1847 ^ n304 ^ 1'b0 ;
  assign n1849 = n150 | n1540 ;
  assign n1850 = n311 | n1173 ;
  assign n1851 = n244 & ~n1850 ;
  assign n1856 = n744 ^ n338 ^ 1'b0 ;
  assign n1857 = ~n1143 & n1856 ;
  assign n1852 = n74 | n563 ;
  assign n1853 = n952 ^ n808 ^ n750 ;
  assign n1854 = n1852 & n1853 ;
  assign n1855 = ~n481 & n1854 ;
  assign n1858 = n1857 ^ n1855 ^ 1'b0 ;
  assign n1860 = n351 & ~n1177 ;
  assign n1861 = ~n760 & n1860 ;
  assign n1859 = n21 & ~n1697 ;
  assign n1862 = n1861 ^ n1859 ^ 1'b0 ;
  assign n1863 = n1381 & n1862 ;
  assign n1867 = n1049 ^ n124 ^ 1'b0 ;
  assign n1868 = n1867 ^ n117 ^ 1'b0 ;
  assign n1869 = n366 | n1868 ;
  assign n1870 = n511 & ~n1869 ;
  assign n1864 = n957 & ~n1121 ;
  assign n1865 = n1138 ^ n541 ^ 1'b0 ;
  assign n1866 = n1864 | n1865 ;
  assign n1871 = n1870 ^ n1866 ^ 1'b0 ;
  assign n1872 = n1871 ^ n782 ^ 1'b0 ;
  assign n1873 = ( n295 & n619 ) | ( n295 & n1409 ) | ( n619 & n1409 ) ;
  assign n1874 = ~n1093 & n1818 ;
  assign n1875 = ~n1873 & n1874 ;
  assign n1876 = n952 ^ n798 ^ 1'b0 ;
  assign n1877 = n330 | n605 ;
  assign n1878 = n83 & n159 ;
  assign n1879 = n1877 & ~n1878 ;
  assign n1880 = n1879 ^ n1845 ^ 1'b0 ;
  assign n1881 = n1774 | n1880 ;
  assign n1882 = n661 | n1881 ;
  assign n1883 = n1439 ^ n88 ^ 1'b0 ;
  assign n1884 = n972 & n1691 ;
  assign n1885 = n852 ^ n124 ^ 1'b0 ;
  assign n1886 = n36 & n1885 ;
  assign n1887 = n1886 ^ n807 ^ 1'b0 ;
  assign n1888 = n1868 & n1887 ;
  assign n1889 = n1888 ^ n574 ^ 1'b0 ;
  assign n1890 = n297 | n1889 ;
  assign n1891 = n219 & ~n1890 ;
  assign n1892 = n931 | n1891 ;
  assign n1893 = ( n112 & n967 ) | ( n112 & ~n1561 ) | ( n967 & ~n1561 ) ;
  assign n1894 = n393 | n1006 ;
  assign n1895 = n1894 ^ n528 ^ 1'b0 ;
  assign n1896 = n1895 ^ n515 ^ 1'b0 ;
  assign n1897 = ~n398 & n441 ;
  assign n1898 = n344 | n1897 ;
  assign n1900 = n225 & ~n588 ;
  assign n1899 = n823 & n828 ;
  assign n1901 = n1900 ^ n1899 ^ 1'b0 ;
  assign n1902 = ~n1898 & n1901 ;
  assign n1903 = n545 ^ n494 ^ 1'b0 ;
  assign n1904 = n494 & n1903 ;
  assign n1905 = ( n221 & n1027 ) | ( n221 & ~n1904 ) | ( n1027 & ~n1904 ) ;
  assign n1906 = ~n205 & n1905 ;
  assign n1907 = n1906 ^ n1905 ^ 1'b0 ;
  assign n1908 = n1054 ^ n846 ^ 1'b0 ;
  assign n1909 = n1908 ^ n263 ^ 1'b0 ;
  assign n1910 = n488 & ~n1909 ;
  assign n1911 = n1443 ^ n798 ^ n280 ;
  assign n1914 = n642 ^ n263 ^ 1'b0 ;
  assign n1912 = ~n606 & n1456 ;
  assign n1913 = n605 & n1912 ;
  assign n1915 = n1914 ^ n1913 ^ 1'b0 ;
  assign n1917 = n712 ^ n234 ^ n133 ;
  assign n1916 = x10 & ~n371 ;
  assign n1918 = n1917 ^ n1916 ^ 1'b0 ;
  assign n1919 = n645 | n1073 ;
  assign n1920 = n1919 ^ n619 ^ 1'b0 ;
  assign n1921 = n1920 ^ n1346 ^ n1105 ;
  assign n1922 = n209 ^ n154 ^ 1'b0 ;
  assign n1923 = n1141 & ~n1922 ;
  assign n1924 = ~n354 & n1923 ;
  assign n1925 = n878 ^ n845 ^ 1'b0 ;
  assign n1926 = n874 ^ n481 ^ 1'b0 ;
  assign n1927 = ~n695 & n1926 ;
  assign n1928 = n1174 & ~n1413 ;
  assign n1929 = n1927 & n1928 ;
  assign n1930 = n1662 ^ n1002 ^ n140 ;
  assign n1931 = n86 & ~n1930 ;
  assign n1932 = ~x3 & n1931 ;
  assign n1933 = n588 ^ n150 ^ 1'b0 ;
  assign n1934 = n821 & ~n1933 ;
  assign n1935 = ~n103 & n1934 ;
  assign n1936 = n841 & n980 ;
  assign n1939 = n781 & ~n920 ;
  assign n1937 = n591 & ~n1677 ;
  assign n1938 = n1937 ^ n764 ^ n220 ;
  assign n1940 = n1939 ^ n1938 ^ 1'b0 ;
  assign n1941 = n1936 & n1940 ;
  assign n1942 = n266 & ~n468 ;
  assign n1943 = n1942 ^ n999 ^ 1'b0 ;
  assign n1944 = n563 & n1943 ;
  assign n1945 = n1574 & n1944 ;
  assign n1946 = ( n709 & ~n747 ) | ( n709 & n1570 ) | ( ~n747 & n1570 ) ;
  assign n1947 = n826 & n1946 ;
  assign n1948 = n173 | n1112 ;
  assign n1949 = n961 & ~n1948 ;
  assign n1950 = ~n588 & n723 ;
  assign n1951 = ~n1628 & n1950 ;
  assign n1954 = n301 & ~n1198 ;
  assign n1955 = n510 & n1954 ;
  assign n1952 = n301 & ~n1652 ;
  assign n1953 = ~n841 & n1952 ;
  assign n1956 = n1955 ^ n1953 ^ 1'b0 ;
  assign n1957 = n1956 ^ n1192 ^ 1'b0 ;
  assign n1958 = n1951 | n1957 ;
  assign n1959 = n386 | n1473 ;
  assign n1960 = n1639 & ~n1959 ;
  assign n1961 = n1960 ^ n717 ^ 1'b0 ;
  assign n1962 = n822 ^ n342 ^ 1'b0 ;
  assign n1963 = ~n533 & n742 ;
  assign n1964 = n1962 & n1963 ;
  assign n1965 = n1961 | n1964 ;
  assign n1966 = n454 & ~n1965 ;
  assign n1967 = n602 ^ n553 ^ 1'b0 ;
  assign n1968 = ( n447 & n877 ) | ( n447 & ~n1967 ) | ( n877 & ~n1967 ) ;
  assign n1969 = n746 ^ n89 ^ 1'b0 ;
  assign n1970 = ~n805 & n1969 ;
  assign n1971 = ~n929 & n1970 ;
  assign n1972 = n772 | n1971 ;
  assign n1973 = ( n1514 & n1654 ) | ( n1514 & n1972 ) | ( n1654 & n1972 ) ;
  assign n1974 = ~n127 & n254 ;
  assign n1975 = n205 & n1974 ;
  assign n1976 = n1653 & n1975 ;
  assign n1977 = n335 | n495 ;
  assign n1978 = n1977 ^ n351 ^ 1'b0 ;
  assign n1979 = n552 ^ n352 ^ 1'b0 ;
  assign n1980 = n1978 & ~n1979 ;
  assign n1981 = n808 | n1659 ;
  assign n1982 = n331 & n1347 ;
  assign n1983 = n1982 ^ n765 ^ 1'b0 ;
  assign n1984 = ( n766 & n1221 ) | ( n766 & n1983 ) | ( n1221 & n1983 ) ;
  assign n1985 = n1984 ^ n692 ^ 1'b0 ;
  assign n1986 = n1891 ^ n83 ^ 1'b0 ;
  assign n1987 = n408 | n697 ;
  assign n1988 = n592 ^ n139 ^ 1'b0 ;
  assign n1989 = n298 & ~n1111 ;
  assign n1990 = n546 ^ n448 ^ 1'b0 ;
  assign n1991 = n23 & n1990 ;
  assign n1992 = n1329 & n1991 ;
  assign n1993 = n1736 & n1992 ;
  assign n1994 = n896 ^ n880 ^ n668 ;
  assign n1995 = n294 & n338 ;
  assign n1996 = n1995 ^ n67 ^ 1'b0 ;
  assign n1997 = n150 | n1996 ;
  assign n1998 = n1994 | n1997 ;
  assign n1999 = n1998 ^ n1915 ^ 1'b0 ;
  assign n2000 = n553 ^ n372 ^ 1'b0 ;
  assign n2001 = n734 & ~n1023 ;
  assign n2002 = n2000 & n2001 ;
  assign n2006 = n582 ^ n43 ^ 1'b0 ;
  assign n2003 = n1075 & n1345 ;
  assign n2004 = n2003 ^ n588 ^ 1'b0 ;
  assign n2005 = n2004 ^ n1215 ^ 1'b0 ;
  assign n2007 = n2006 ^ n2005 ^ 1'b0 ;
  assign n2008 = n1845 ^ n241 ^ 1'b0 ;
  assign n2009 = n733 & ~n1224 ;
  assign n2010 = ~n810 & n2009 ;
  assign n2013 = n439 & n1050 ;
  assign n2014 = n2013 ^ n227 ^ 1'b0 ;
  assign n2015 = ~n762 & n2014 ;
  assign n2016 = n822 & n2015 ;
  assign n2011 = n976 | n1901 ;
  assign n2012 = n2011 ^ n28 ^ 1'b0 ;
  assign n2017 = n2016 ^ n2012 ^ n345 ;
  assign n2018 = n851 ^ n528 ^ 1'b0 ;
  assign n2019 = n1045 & n2018 ;
  assign n2020 = n1978 ^ n368 ^ 1'b0 ;
  assign n2021 = n983 | n2020 ;
  assign n2022 = n1201 & ~n2021 ;
  assign n2023 = n454 | n1691 ;
  assign n2024 = n1932 ^ n744 ^ 1'b0 ;
  assign n2027 = ~n732 & n983 ;
  assign n2028 = ~n1119 & n2027 ;
  assign n2026 = ~n393 & n552 ;
  assign n2029 = n2028 ^ n2026 ^ 1'b0 ;
  assign n2025 = n129 & ~n428 ;
  assign n2030 = n2029 ^ n2025 ^ 1'b0 ;
  assign n2031 = n965 ^ n105 ^ 1'b0 ;
  assign n2032 = n2031 ^ n749 ^ 1'b0 ;
  assign n2033 = ~n339 & n1707 ;
  assign n2034 = n1264 ^ n901 ^ 1'b0 ;
  assign n2035 = n179 | n1870 ;
  assign n2036 = n2035 ^ n1980 ^ 1'b0 ;
  assign n2037 = n1045 & n2036 ;
  assign n2038 = n2037 ^ n681 ^ 1'b0 ;
  assign n2039 = ~n422 & n2038 ;
  assign n2040 = n89 & ~n1191 ;
  assign n2041 = n2040 ^ n1816 ^ n873 ;
  assign n2042 = n195 & n216 ;
  assign n2043 = n1540 & n2042 ;
  assign n2044 = n2043 ^ n1267 ^ 1'b0 ;
  assign n2045 = n521 & ~n709 ;
  assign n2046 = n1234 ^ n248 ^ 1'b0 ;
  assign n2047 = ~n433 & n1588 ;
  assign n2048 = n840 & n2047 ;
  assign n2049 = n592 & n1189 ;
  assign n2050 = n2049 ^ n1576 ^ n1306 ;
  assign n2051 = n1633 ^ n837 ^ 1'b0 ;
  assign n2052 = n1726 ^ n488 ^ 1'b0 ;
  assign n2053 = ~n1186 & n2052 ;
  assign n2054 = ( ~n318 & n924 ) | ( ~n318 & n2053 ) | ( n924 & n2053 ) ;
  assign n2055 = n2051 & ~n2054 ;
  assign n2056 = n1770 ^ n680 ^ 1'b0 ;
  assign n2057 = ~n873 & n1068 ;
  assign n2058 = n2057 ^ n680 ^ 1'b0 ;
  assign n2059 = n2058 ^ n588 ^ 1'b0 ;
  assign n2060 = n2056 | n2059 ;
  assign n2061 = ~n347 & n408 ;
  assign n2062 = n398 | n1224 ;
  assign n2063 = n600 & ~n2062 ;
  assign n2064 = x3 & n1027 ;
  assign n2065 = n2064 ^ n593 ^ 1'b0 ;
  assign n2066 = n2065 ^ n188 ^ 1'b0 ;
  assign n2071 = n651 & ~n741 ;
  assign n2072 = n2071 ^ n565 ^ 1'b0 ;
  assign n2068 = ~n322 & n1093 ;
  assign n2069 = ~n226 & n1365 ;
  assign n2070 = n2068 & n2069 ;
  assign n2073 = n2072 ^ n2070 ^ 1'b0 ;
  assign n2074 = n2073 ^ n1886 ^ n255 ;
  assign n2075 = ~n259 & n920 ;
  assign n2076 = ~n2074 & n2075 ;
  assign n2067 = n1023 ^ n511 ^ 1'b0 ;
  assign n2077 = n2076 ^ n2067 ^ 1'b0 ;
  assign n2078 = n131 & n1289 ;
  assign n2079 = n2078 ^ n631 ^ n404 ;
  assign n2080 = n1546 & n2079 ;
  assign n2081 = n796 ^ n459 ^ n458 ;
  assign n2082 = n648 ^ n362 ^ 1'b0 ;
  assign n2083 = n2082 ^ n1912 ^ 1'b0 ;
  assign n2084 = n2083 ^ n1763 ^ 1'b0 ;
  assign n2085 = ~n2081 & n2084 ;
  assign n2086 = ( ~n634 & n808 ) | ( ~n634 & n1304 ) | ( n808 & n1304 ) ;
  assign n2087 = n1592 & n2086 ;
  assign n2089 = n1054 ^ n1047 ^ 1'b0 ;
  assign n2090 = n1414 & ~n2089 ;
  assign n2088 = n124 | n227 ;
  assign n2091 = n2090 ^ n2088 ^ 1'b0 ;
  assign n2092 = n1525 ^ n144 ^ 1'b0 ;
  assign n2093 = n828 & n2092 ;
  assign n2094 = n400 & ~n936 ;
  assign n2095 = n1312 ^ n842 ^ 1'b0 ;
  assign n2096 = n839 & n2095 ;
  assign n2097 = n2096 ^ n929 ^ 1'b0 ;
  assign n2098 = ( n396 & n1730 ) | ( n396 & ~n2097 ) | ( n1730 & ~n2097 ) ;
  assign n2099 = n545 ^ n47 ^ 1'b0 ;
  assign n2100 = n1522 | n2099 ;
  assign n2101 = n2100 ^ n571 ^ 1'b0 ;
  assign n2102 = n919 & n2101 ;
  assign n2103 = ~n572 & n1823 ;
  assign n2104 = n922 ^ n173 ^ 1'b0 ;
  assign n2105 = n2104 ^ n917 ^ 1'b0 ;
  assign n2106 = n1876 & ~n2105 ;
  assign n2107 = n1743 ^ n700 ^ 1'b0 ;
  assign n2108 = n331 & ~n2107 ;
  assign n2109 = n782 ^ n131 ^ 1'b0 ;
  assign n2110 = n1675 ^ n290 ^ 1'b0 ;
  assign n2111 = ~n1726 & n1857 ;
  assign n2112 = n2111 ^ n1653 ^ 1'b0 ;
  assign n2113 = n1042 | n1904 ;
  assign n2114 = ( n744 & ~n2065 ) | ( n744 & n2113 ) | ( ~n2065 & n2113 ) ;
  assign n2115 = n1832 | n2032 ;
  assign n2116 = n2114 | n2115 ;
  assign n2117 = ~x6 & n786 ;
  assign n2118 = n347 | n2117 ;
  assign n2119 = n2118 ^ n1744 ^ 1'b0 ;
  assign n2120 = n81 & n2119 ;
  assign n2121 = n112 | n782 ;
  assign n2122 = n985 & ~n1540 ;
  assign n2123 = n2121 & n2122 ;
  assign n2124 = n2018 & n2123 ;
  assign n2125 = n2124 ^ n1052 ^ 1'b0 ;
  assign n2126 = n417 | n2125 ;
  assign n2127 = n1336 | n2126 ;
  assign n2128 = n261 ^ n28 ^ 1'b0 ;
  assign n2129 = n423 ^ n305 ^ 1'b0 ;
  assign n2130 = n684 & ~n1543 ;
  assign n2131 = ~n1094 & n2130 ;
  assign n2132 = n1398 & n2131 ;
  assign n2133 = n414 & ~n1123 ;
  assign n2134 = ( n1955 & n2132 ) | ( n1955 & ~n2133 ) | ( n2132 & ~n2133 ) ;
  assign n2135 = ~n98 & n239 ;
  assign n2136 = n640 & n2135 ;
  assign n2137 = n335 | n415 ;
  assign n2138 = ( ~n1167 & n1516 ) | ( ~n1167 & n2137 ) | ( n1516 & n2137 ) ;
  assign n2139 = n244 ^ n194 ^ 1'b0 ;
  assign n2140 = n2139 ^ n839 ^ 1'b0 ;
  assign n2141 = n646 & n2140 ;
  assign n2142 = n582 ^ n17 ^ 1'b0 ;
  assign n2143 = n246 & n2142 ;
  assign n2144 = n1221 & n2143 ;
  assign n2145 = n2144 ^ n1803 ^ 1'b0 ;
  assign n2146 = n1337 | n1523 ;
  assign n2147 = ~n225 & n1884 ;
  assign n2148 = n2147 ^ n1441 ^ 1'b0 ;
  assign n2149 = n1483 ^ x11 ^ 1'b0 ;
  assign n2150 = ~n592 & n2149 ;
  assign n2151 = n1560 ^ n466 ^ 1'b0 ;
  assign n2152 = ~n1238 & n2151 ;
  assign n2153 = n2152 ^ n849 ^ 1'b0 ;
  assign n2154 = n2150 & ~n2153 ;
  assign n2155 = ~n13 & n433 ;
  assign n2156 = n1212 ^ n500 ^ 1'b0 ;
  assign n2157 = n1344 | n2156 ;
  assign n2158 = n1971 ^ n56 ^ 1'b0 ;
  assign n2159 = ( n652 & ~n1345 ) | ( n652 & n1707 ) | ( ~n1345 & n1707 ) ;
  assign n2164 = n33 | n453 ;
  assign n2165 = n506 | n2164 ;
  assign n2166 = n2165 ^ n645 ^ 1'b0 ;
  assign n2160 = n875 & n1329 ;
  assign n2161 = n2160 ^ n548 ^ 1'b0 ;
  assign n2162 = n2161 ^ x5 ^ 1'b0 ;
  assign n2163 = ~n1036 & n2162 ;
  assign n2167 = n2166 ^ n2163 ^ 1'b0 ;
  assign n2168 = n1835 | n2167 ;
  assign n2169 = n809 & ~n993 ;
  assign n2170 = n2169 ^ n1821 ^ 1'b0 ;
  assign n2171 = ~n485 & n1980 ;
  assign n2172 = n2171 ^ n1868 ^ 1'b0 ;
  assign n2173 = n195 & ~n757 ;
  assign n2174 = ~n2172 & n2173 ;
  assign n2175 = n1811 & n2174 ;
  assign n2176 = n1598 & n2091 ;
  assign n2177 = n683 ^ n536 ^ 1'b0 ;
  assign n2178 = ~n1212 & n2177 ;
  assign n2179 = n839 ^ n612 ^ 1'b0 ;
  assign n2180 = n2179 ^ n684 ^ 1'b0 ;
  assign n2181 = n1229 | n2180 ;
  assign n2182 = x8 & ~n2181 ;
  assign n2183 = n2182 ^ n1938 ^ 1'b0 ;
  assign n2184 = ~n2178 & n2183 ;
  assign n2185 = n793 ^ n338 ^ 1'b0 ;
  assign n2186 = n1320 & n2185 ;
  assign n2187 = ~n362 & n478 ;
  assign n2188 = n2187 ^ n815 ^ 1'b0 ;
  assign n2189 = n2188 ^ n395 ^ n35 ;
  assign n2190 = n470 & ~n1707 ;
  assign n2191 = n2190 ^ n744 ^ 1'b0 ;
  assign n2192 = ~n2189 & n2191 ;
  assign n2193 = ( n657 & ~n839 ) | ( n657 & n2192 ) | ( ~n839 & n2192 ) ;
  assign n2194 = ~n1843 & n2193 ;
  assign n2195 = ~n2188 & n2194 ;
  assign n2196 = n296 ^ n267 ^ 1'b0 ;
  assign n2197 = n19 | n2196 ;
  assign n2198 = n387 | n2197 ;
  assign n2199 = n74 | n2198 ;
  assign n2200 = ~n347 & n2199 ;
  assign n2201 = n2200 ^ n1058 ^ 1'b0 ;
  assign n2202 = n2201 ^ n186 ^ 1'b0 ;
  assign n2203 = n2177 | n2202 ;
  assign n2204 = n522 & n774 ;
  assign n2205 = n148 & ~n832 ;
  assign n2206 = ~n506 & n2205 ;
  assign n2207 = ( n205 & n239 ) | ( n205 & n2206 ) | ( n239 & n2206 ) ;
  assign n2208 = n1208 | n1365 ;
  assign n2209 = n677 & n2208 ;
  assign n2210 = ~n1685 & n2209 ;
  assign n2211 = x6 & n751 ;
  assign n2212 = ( ~n541 & n1284 ) | ( ~n541 & n1304 ) | ( n1284 & n1304 ) ;
  assign n2213 = n722 ^ n541 ^ 1'b0 ;
  assign n2214 = n2213 ^ n1016 ^ n52 ;
  assign n2215 = n980 ^ n340 ^ 1'b0 ;
  assign n2216 = n20 | n2215 ;
  assign n2217 = n1189 | n2216 ;
  assign n2221 = n961 ^ n533 ^ 1'b0 ;
  assign n2222 = ~n993 & n2221 ;
  assign n2218 = n1376 ^ n1124 ^ 1'b0 ;
  assign n2219 = ( n682 & n1995 ) | ( n682 & n2218 ) | ( n1995 & n2218 ) ;
  assign n2220 = n365 & n2219 ;
  assign n2223 = n2222 ^ n2220 ^ 1'b0 ;
  assign n2224 = n1235 ^ n148 ^ 1'b0 ;
  assign n2225 = n1119 & n2224 ;
  assign n2226 = n2225 ^ n676 ^ n582 ;
  assign n2227 = n965 & ~n2226 ;
  assign n2228 = n890 & ~n1278 ;
  assign n2229 = n1205 & ~n2228 ;
  assign n2230 = ~n374 & n1921 ;
  assign n2231 = ~n1750 & n2016 ;
  assign n2232 = n1418 ^ n418 ^ n286 ;
  assign n2233 = ( n162 & ~n1858 ) | ( n162 & n2232 ) | ( ~n1858 & n2232 ) ;
  assign n2234 = n530 & ~n1594 ;
  assign n2235 = n927 & n2234 ;
  assign n2236 = ( n208 & n326 ) | ( n208 & n970 ) | ( n326 & n970 ) ;
  assign n2237 = ~n395 & n1641 ;
  assign n2238 = n2236 & n2237 ;
  assign n2239 = n1476 ^ n970 ^ 1'b0 ;
  assign n2240 = n2238 & ~n2239 ;
  assign n2241 = n833 & n885 ;
  assign n2242 = n1867 & n2241 ;
  assign n2243 = ~n571 & n2242 ;
  assign n2244 = n2243 ^ n390 ^ 1'b0 ;
  assign n2245 = n493 & ~n709 ;
  assign n2246 = n2245 ^ x5 ^ 1'b0 ;
  assign n2247 = n1099 | n1347 ;
  assign n2248 = ( n363 & n1293 ) | ( n363 & n1677 ) | ( n1293 & n1677 ) ;
  assign n2249 = n688 & n1439 ;
  assign n2250 = ~n2248 & n2249 ;
  assign n2251 = n1040 | n1419 ;
  assign n2252 = n225 | n2251 ;
  assign n2253 = n13 & n2077 ;
  assign n2254 = n584 & n1518 ;
  assign n2255 = n995 ^ n149 ^ 1'b0 ;
  assign n2256 = ~n2254 & n2255 ;
  assign n2257 = ( n758 & ~n1277 ) | ( n758 & n2058 ) | ( ~n1277 & n2058 ) ;
  assign n2258 = n1216 | n1491 ;
  assign n2259 = n40 | n2258 ;
  assign n2260 = n752 & ~n2259 ;
  assign n2261 = ( ~n1664 & n2257 ) | ( ~n1664 & n2260 ) | ( n2257 & n2260 ) ;
  assign n2262 = n714 ^ n257 ^ n125 ;
  assign n2263 = n744 & ~n2100 ;
  assign n2264 = ~n2262 & n2263 ;
  assign n2265 = ( n684 & ~n737 ) | ( n684 & n2264 ) | ( ~n737 & n2264 ) ;
  assign n2267 = ~n69 & n1647 ;
  assign n2268 = ~n372 & n2267 ;
  assign n2266 = ~n1271 & n1943 ;
  assign n2269 = n2268 ^ n2266 ^ 1'b0 ;
  assign n2270 = n2155 & ~n2269 ;
  assign n2272 = n924 ^ n837 ^ 1'b0 ;
  assign n2271 = n555 & n2014 ;
  assign n2273 = n2272 ^ n2271 ^ 1'b0 ;
  assign n2274 = n781 ^ n586 ^ 1'b0 ;
  assign n2275 = n738 & ~n2274 ;
  assign n2276 = ~n2273 & n2275 ;
  assign n2277 = n2276 ^ n1933 ^ 1'b0 ;
  assign n2278 = n2277 ^ n1624 ^ 1'b0 ;
  assign n2279 = n864 | n2278 ;
  assign n2281 = n774 & ~n1430 ;
  assign n2282 = n159 & n2281 ;
  assign n2283 = n2282 ^ n801 ^ 1'b0 ;
  assign n2280 = n105 & ~n2228 ;
  assign n2284 = n2283 ^ n2280 ^ 1'b0 ;
  assign n2285 = n2284 ^ n932 ^ 1'b0 ;
  assign n2286 = n1425 & n2285 ;
  assign n2287 = ( n1367 & n1607 ) | ( n1367 & ~n1880 ) | ( n1607 & ~n1880 ) ;
  assign n2288 = ( n107 & n124 ) | ( n107 & n2287 ) | ( n124 & n2287 ) ;
  assign n2289 = n2236 ^ n1200 ^ 1'b0 ;
  assign n2290 = n729 & ~n2289 ;
  assign n2291 = n440 & ~n2290 ;
  assign n2292 = ( n130 & ~n861 ) | ( n130 & n2137 ) | ( ~n861 & n2137 ) ;
  assign n2293 = n720 ^ n304 ^ 1'b0 ;
  assign n2294 = n2292 & n2293 ;
  assign n2302 = n2022 ^ n223 ^ 1'b0 ;
  assign n2303 = n192 & ~n2302 ;
  assign n2295 = n320 & ~n325 ;
  assign n2296 = n2295 ^ n440 ^ 1'b0 ;
  assign n2297 = n2137 ^ n432 ^ 1'b0 ;
  assign n2298 = n714 | n2297 ;
  assign n2299 = n2296 | n2298 ;
  assign n2300 = n2299 ^ n1744 ^ 1'b0 ;
  assign n2301 = ~n1933 & n2300 ;
  assign n2304 = n2303 ^ n2301 ^ 1'b0 ;
  assign n2305 = n1627 | n2304 ;
  assign n2306 = n1729 | n2305 ;
  assign n2307 = n2306 ^ n1486 ^ 1'b0 ;
  assign n2308 = n2294 & n2307 ;
  assign n2309 = n94 & ~n1697 ;
  assign n2310 = n458 & ~n2062 ;
  assign n2311 = n1394 & n2310 ;
  assign n2312 = n2024 ^ n179 ^ 1'b0 ;
  assign n2313 = n113 & ~n2312 ;
  assign n2314 = n54 & n1697 ;
  assign n2315 = n61 & n2314 ;
  assign n2316 = n2315 ^ n2046 ^ n17 ;
  assign n2317 = n523 | n2262 ;
  assign n2318 = n2317 ^ n2283 ^ 1'b0 ;
  assign n2319 = n2318 ^ n1542 ^ 1'b0 ;
  assign n2320 = n1052 ^ n839 ^ n746 ;
  assign n2321 = n2166 ^ n867 ^ 1'b0 ;
  assign n2327 = n1223 | n1257 ;
  assign n2322 = n956 ^ n753 ^ 1'b0 ;
  assign n2323 = n235 & n2272 ;
  assign n2324 = n2323 ^ n1003 ^ 1'b0 ;
  assign n2325 = ~n2322 & n2324 ;
  assign n2326 = ~n1116 & n2325 ;
  assign n2328 = n2327 ^ n2326 ^ n344 ;
  assign n2329 = ~n347 & n1071 ;
  assign n2330 = n2329 ^ n218 ^ 1'b0 ;
  assign n2331 = ( n63 & n800 ) | ( n63 & ~n2330 ) | ( n800 & ~n2330 ) ;
  assign n2332 = n466 | n1109 ;
  assign n2333 = n360 | n2332 ;
  assign n2334 = n2318 & ~n2333 ;
  assign n2335 = n51 & ~n2143 ;
  assign n2336 = n542 | n2008 ;
  assign n2337 = n135 & n2014 ;
  assign n2338 = n967 | n2337 ;
  assign n2339 = n1668 & n2338 ;
  assign n2340 = ~n1721 & n2339 ;
  assign n2341 = n108 | n2098 ;
  assign n2346 = n673 ^ n419 ^ 1'b0 ;
  assign n2347 = ~n1027 & n2346 ;
  assign n2345 = n299 & ~n1745 ;
  assign n2348 = n2347 ^ n2345 ^ 1'b0 ;
  assign n2342 = n1534 & ~n1553 ;
  assign n2343 = n2342 ^ n791 ^ 1'b0 ;
  assign n2344 = ~n1609 & n2343 ;
  assign n2349 = n2348 ^ n2344 ^ 1'b0 ;
  assign n2350 = n1419 ^ n1134 ^ n983 ;
  assign n2351 = n2350 ^ n1284 ^ 1'b0 ;
  assign n2352 = n1534 ^ n707 ^ n481 ;
  assign n2353 = ( ~n475 & n2315 ) | ( ~n475 & n2352 ) | ( n2315 & n2352 ) ;
  assign n2354 = ~n305 & n1453 ;
  assign n2355 = n2354 ^ n1198 ^ 1'b0 ;
  assign n2356 = n1327 ^ n555 ^ 1'b0 ;
  assign n2357 = n714 | n2356 ;
  assign n2358 = n235 | n2357 ;
  assign n2359 = n546 & n1510 ;
  assign n2360 = n2358 & ~n2359 ;
  assign n2361 = ~n2355 & n2360 ;
  assign n2362 = ~n533 & n2361 ;
  assign n2363 = n170 | n1794 ;
  assign n2364 = n2363 ^ n270 ^ 1'b0 ;
  assign n2365 = n1298 & n2364 ;
  assign n2366 = n2365 ^ n2173 ^ 1'b0 ;
  assign n2367 = n2024 ^ n1464 ^ 1'b0 ;
  assign n2368 = ( n1081 & n2014 ) | ( n1081 & n2317 ) | ( n2014 & n2317 ) ;
  assign n2369 = n2368 ^ n749 ^ 1'b0 ;
  assign n2370 = n1246 & ~n2369 ;
  assign n2371 = n841 & n2370 ;
  assign n2372 = n43 & ~n802 ;
  assign n2373 = n1060 & n2372 ;
  assign n2374 = n165 & ~n2373 ;
  assign n2375 = n139 | n317 ;
  assign n2376 = n1953 & ~n2375 ;
  assign n2380 = ~n207 & n1306 ;
  assign n2377 = n2095 ^ n349 ^ 1'b0 ;
  assign n2378 = n2377 ^ n1392 ^ 1'b0 ;
  assign n2379 = n1792 | n2378 ;
  assign n2381 = n2380 ^ n2379 ^ 1'b0 ;
  assign n2382 = n1363 ^ n588 ^ 1'b0 ;
  assign n2383 = n333 ^ n191 ^ 1'b0 ;
  assign n2384 = ~n1181 & n2383 ;
  assign n2385 = ~n907 & n2384 ;
  assign n2386 = n2385 ^ n1117 ^ 1'b0 ;
  assign n2387 = n465 & ~n988 ;
  assign n2388 = ~n1207 & n1229 ;
  assign n2389 = n2388 ^ n968 ^ 1'b0 ;
  assign n2390 = n749 & n2389 ;
  assign n2391 = ~n1409 & n2158 ;
  assign n2392 = n2390 & ~n2391 ;
  assign n2393 = ~n706 & n2392 ;
  assign n2394 = ~n667 & n1340 ;
  assign n2395 = n275 | n542 ;
  assign n2396 = n373 | n2395 ;
  assign n2397 = n2396 ^ n177 ^ 1'b0 ;
  assign n2398 = n2397 ^ n777 ^ 1'b0 ;
  assign n2399 = ( ~n21 & n2394 ) | ( ~n21 & n2398 ) | ( n2394 & n2398 ) ;
  assign n2400 = ~n57 & n1667 ;
  assign n2401 = n2231 & n2400 ;
  assign n2402 = n237 & ~n255 ;
  assign n2403 = n186 & n2402 ;
  assign n2404 = n725 | n2403 ;
  assign n2405 = n2404 ^ n791 ^ n651 ;
  assign n2406 = ~n1038 & n2405 ;
  assign n2407 = n924 & n1720 ;
  assign n2408 = ~n395 & n2347 ;
  assign n2409 = ( n1882 & n2407 ) | ( n1882 & n2408 ) | ( n2407 & n2408 ) ;
  assign n2410 = ~n591 & n2409 ;
  assign n2411 = n2410 ^ n2391 ^ 1'b0 ;
  assign n2415 = n1049 | n1169 ;
  assign n2416 = n2415 ^ n20 ^ 1'b0 ;
  assign n2417 = n1336 & n2416 ;
  assign n2418 = n929 ^ n418 ^ 1'b0 ;
  assign n2419 = n1744 & n2418 ;
  assign n2420 = n2417 & n2419 ;
  assign n2412 = n1367 | n1694 ;
  assign n2413 = n1014 & ~n2412 ;
  assign n2414 = n2322 | n2413 ;
  assign n2421 = n2420 ^ n2414 ^ 1'b0 ;
  assign n2422 = ~n2401 & n2421 ;
  assign n2423 = ~n1554 & n2422 ;
  assign n2425 = n965 ^ n318 ^ n23 ;
  assign n2424 = ~n767 & n1340 ;
  assign n2426 = n2425 ^ n2424 ^ n1066 ;
  assign n2427 = ~n1246 & n1540 ;
  assign n2428 = ~n356 & n2427 ;
  assign n2429 = n79 | n1261 ;
  assign n2430 = n2072 ^ n98 ^ 1'b0 ;
  assign n2431 = n2429 | n2430 ;
  assign n2432 = ~n734 & n975 ;
  assign n2433 = ( ~n1740 & n2022 ) | ( ~n1740 & n2432 ) | ( n2022 & n2432 ) ;
  assign n2434 = n404 & n482 ;
  assign n2435 = ~n160 & n2434 ;
  assign n2436 = n1443 & ~n2435 ;
  assign n2437 = n2436 ^ n2377 ^ 1'b0 ;
  assign n2438 = n103 & ~n1014 ;
  assign n2439 = n2438 ^ n1363 ^ n510 ;
  assign n2440 = n219 | n870 ;
  assign n2441 = ~n2439 & n2440 ;
  assign n2442 = ~n392 & n2441 ;
  assign n2443 = n1428 ^ n807 ^ 1'b0 ;
  assign n2444 = n1064 ^ n820 ^ 1'b0 ;
  assign n2445 = n2444 ^ n1947 ^ n1243 ;
  assign n2446 = n1173 & n2445 ;
  assign n2447 = n1728 ^ n870 ^ 1'b0 ;
  assign n2448 = n1351 & n2447 ;
  assign n2449 = ~n680 & n1490 ;
  assign n2450 = ~n1460 & n2449 ;
  assign n2451 = ~n1723 & n2450 ;
  assign n2452 = n488 & ~n2155 ;
  assign n2453 = n919 & ~n1755 ;
  assign n2454 = n2453 ^ n765 ^ 1'b0 ;
  assign n2455 = ~n1586 & n2454 ;
  assign n2456 = n2455 ^ n1703 ^ n845 ;
  assign n2457 = n237 & n1163 ;
  assign n2458 = n2457 ^ n395 ^ 1'b0 ;
  assign n2459 = n131 | n1205 ;
  assign n2460 = n2459 ^ n294 ^ 1'b0 ;
  assign n2461 = n1071 | n2460 ;
  assign n2462 = n2461 ^ n2118 ^ 1'b0 ;
  assign n2463 = n2356 ^ n453 ^ 1'b0 ;
  assign n2464 = n2463 ^ n195 ^ 1'b0 ;
  assign n2465 = ~n749 & n2464 ;
  assign n2466 = n21 & ~n593 ;
  assign n2467 = n2466 ^ n2077 ^ 1'b0 ;
  assign n2468 = n1867 ^ n785 ^ 1'b0 ;
  assign n2469 = n2468 ^ n126 ^ 1'b0 ;
  assign n2470 = n1237 ^ n231 ^ 1'b0 ;
  assign n2471 = n642 & ~n2470 ;
  assign n2472 = ( ~n316 & n1932 ) | ( ~n316 & n2471 ) | ( n1932 & n2471 ) ;
  assign n2473 = n844 | n2273 ;
  assign n2474 = n2473 ^ n36 ^ 1'b0 ;
  assign n2475 = n2114 & n2150 ;
  assign n2476 = ~n239 & n2475 ;
  assign n2477 = n2437 ^ n1344 ^ 1'b0 ;
  assign n2478 = n793 | n2477 ;
  assign n2479 = n220 & ~n1756 ;
  assign n2480 = n2479 ^ n989 ^ 1'b0 ;
  assign n2481 = ~n1134 & n2453 ;
  assign n2482 = n1980 & ~n2481 ;
  assign n2483 = n1439 & ~n2482 ;
  assign n2484 = n344 | n961 ;
  assign n2485 = n1615 | n2484 ;
  assign n2486 = n2273 & ~n2485 ;
  assign n2487 = n1445 | n2486 ;
  assign n2488 = n774 | n2487 ;
  assign n2489 = n2100 ^ n1873 ^ 1'b0 ;
  assign n2490 = ~n620 & n1100 ;
  assign n2491 = n211 & n2490 ;
  assign n2492 = n2491 ^ n676 ^ 1'b0 ;
  assign n2493 = n1042 | n1372 ;
  assign n2494 = n2493 ^ n1740 ^ 1'b0 ;
  assign n2495 = n749 & n1469 ;
  assign n2496 = n2188 ^ n527 ^ 1'b0 ;
  assign n2497 = n2495 & n2496 ;
  assign n2498 = n1542 & n2497 ;
  assign n2499 = n2117 & ~n2483 ;
  assign n2500 = ~n1695 & n2499 ;
  assign n2501 = n968 ^ n458 ^ n302 ;
  assign n2502 = n1107 & ~n2501 ;
  assign n2503 = ~n586 & n1365 ;
  assign n2504 = n2503 ^ n2082 ^ 1'b0 ;
  assign n2505 = n1536 ^ n1241 ^ 1'b0 ;
  assign n2506 = ~n553 & n2505 ;
  assign n2507 = n2506 ^ n2087 ^ 1'b0 ;
  assign n2508 = n74 | n451 ;
  assign n2509 = n1760 & n2508 ;
  assign n2510 = n2509 ^ n1821 ^ 1'b0 ;
  assign n2511 = n1556 ^ n521 ^ 1'b0 ;
  assign n2512 = n1246 & ~n2511 ;
  assign n2513 = n1223 | n2446 ;
  assign n2517 = n1226 ^ n288 ^ 1'b0 ;
  assign n2514 = n2352 ^ n772 ^ 1'b0 ;
  assign n2515 = n600 & n2514 ;
  assign n2516 = n2102 & n2515 ;
  assign n2518 = n2517 ^ n2516 ^ 1'b0 ;
  assign n2519 = n1124 ^ n130 ^ 1'b0 ;
  assign n2520 = n1677 & n2519 ;
  assign n2521 = n2520 ^ n1443 ^ 1'b0 ;
  assign n2522 = n2213 ^ n461 ^ 1'b0 ;
  assign n2523 = n2522 ^ n2098 ^ 1'b0 ;
  assign n2524 = n1064 ^ n379 ^ 1'b0 ;
  assign n2525 = n181 ^ x10 ^ 1'b0 ;
  assign n2526 = n2524 & n2525 ;
  assign n2528 = n1458 ^ n508 ^ 1'b0 ;
  assign n2529 = n277 | n2528 ;
  assign n2527 = ( ~x8 & n1422 ) | ( ~x8 & n2068 ) | ( n1422 & n2068 ) ;
  assign n2530 = n2529 ^ n2527 ^ 1'b0 ;
  assign n2531 = n2526 & n2530 ;
  assign n2532 = n2177 ^ n2109 ^ 1'b0 ;
  assign n2533 = n710 & ~n1878 ;
  assign n2534 = n2533 ^ n1511 ^ 1'b0 ;
  assign n2535 = n664 | n2534 ;
  assign n2536 = ( ~n747 & n1622 ) | ( ~n747 & n1694 ) | ( n1622 & n1694 ) ;
  assign n2537 = ~n1513 & n1752 ;
  assign n2538 = n2537 ^ n1714 ^ 1'b0 ;
  assign n2539 = n2536 | n2538 ;
  assign n2540 = n938 ^ n645 ^ 1'b0 ;
  assign n2541 = n1832 ^ n1414 ^ 1'b0 ;
  assign n2542 = n2541 ^ n765 ^ 1'b0 ;
  assign n2543 = n2540 & ~n2542 ;
  assign n2544 = n1439 ^ n792 ^ 1'b0 ;
  assign n2545 = n2036 & ~n2544 ;
  assign n2546 = n625 & n2545 ;
  assign n2547 = n683 & n2546 ;
  assign n2548 = n751 ^ n694 ^ n363 ;
  assign n2549 = n2548 ^ n2110 ^ 1'b0 ;
  assign n2550 = n620 | n2042 ;
  assign n2551 = ( ~n315 & n518 ) | ( ~n315 & n2550 ) | ( n518 & n2550 ) ;
  assign n2552 = n1045 & n1592 ;
  assign n2553 = n2368 & n2552 ;
  assign n2554 = n2553 ^ n409 ^ 1'b0 ;
  assign n2555 = n493 & n1712 ;
  assign n2556 = n2260 ^ n259 ^ 1'b0 ;
  assign n2557 = ~n841 & n2143 ;
  assign n2558 = n2557 ^ n959 ^ 1'b0 ;
  assign n2559 = n2558 ^ n625 ^ 1'b0 ;
  assign n2560 = n2556 | n2559 ;
  assign n2561 = n45 | n371 ;
  assign n2562 = n1569 | n2561 ;
  assign n2563 = n2562 ^ n2222 ^ x5 ;
  assign n2564 = n1570 ^ n477 ^ 1'b0 ;
  assign n2565 = n1889 ^ n466 ^ 1'b0 ;
  assign n2566 = n1745 & ~n2565 ;
  assign n2567 = n2222 ^ n443 ^ 1'b0 ;
  assign n2568 = n2567 ^ n652 ^ 1'b0 ;
  assign n2569 = n162 & ~n1286 ;
  assign n2570 = n1010 & n1755 ;
  assign n2571 = n1980 & ~n2570 ;
  assign n2575 = n450 ^ n173 ^ 1'b0 ;
  assign n2576 = n221 & ~n231 ;
  assign n2577 = n2575 | n2576 ;
  assign n2572 = n1736 ^ n365 ^ 1'b0 ;
  assign n2573 = n2572 ^ n807 ^ 1'b0 ;
  assign n2574 = n1169 & n2573 ;
  assign n2578 = n2577 ^ n2574 ^ n67 ;
  assign n2580 = n229 ^ n115 ^ 1'b0 ;
  assign n2579 = ~n560 & n2452 ;
  assign n2581 = n2580 ^ n2579 ^ 1'b0 ;
  assign n2582 = n615 & ~n911 ;
  assign n2583 = n1212 & n2582 ;
  assign n2584 = n2583 ^ n631 ^ 1'b0 ;
  assign n2585 = n1672 | n2584 ;
  assign n2586 = n1650 & ~n2585 ;
  assign n2587 = n1114 & ~n2586 ;
  assign n2588 = n344 ^ n76 ^ 1'b0 ;
  assign n2589 = n2580 ^ n428 ^ 1'b0 ;
  assign n2590 = x6 & n61 ;
  assign n2591 = n2590 ^ n862 ^ 1'b0 ;
  assign n2592 = n2591 ^ n1016 ^ 1'b0 ;
  assign n2593 = n2589 & ~n2592 ;
  assign n2594 = n1624 & n2371 ;
  assign n2595 = n1664 ^ n144 ^ 1'b0 ;
  assign n2597 = n1337 & ~n1686 ;
  assign n2598 = n2597 ^ n1098 ^ 1'b0 ;
  assign n2599 = n1697 | n2598 ;
  assign n2600 = n2599 ^ n661 ^ 1'b0 ;
  assign n2596 = n1340 & n2331 ;
  assign n2601 = n2600 ^ n2596 ^ 1'b0 ;
  assign n2608 = n1806 ^ n445 ^ 1'b0 ;
  assign n2609 = n227 & ~n2608 ;
  assign n2602 = ~n316 & n398 ;
  assign n2603 = n568 ^ n521 ^ 1'b0 ;
  assign n2604 = n2197 ^ n765 ^ 1'b0 ;
  assign n2605 = ( n1694 & ~n2603 ) | ( n1694 & n2604 ) | ( ~n2603 & n2604 ) ;
  assign n2606 = n2605 ^ n2589 ^ 1'b0 ;
  assign n2607 = n2602 & ~n2606 ;
  assign n2610 = n2609 ^ n2607 ^ 1'b0 ;
  assign n2611 = n1645 | n2610 ;
  assign n2612 = n2611 ^ n1908 ^ 1'b0 ;
  assign n2614 = n372 ^ x4 ^ 1'b0 ;
  assign n2615 = ~n1790 & n2614 ;
  assign n2613 = n484 & n1660 ;
  assign n2616 = n2615 ^ n2613 ^ 1'b0 ;
  assign n2617 = n1562 | n2616 ;
  assign n2618 = n2617 ^ n659 ^ 1'b0 ;
  assign n2619 = n619 ^ n239 ^ n51 ;
  assign n2620 = ~n387 & n600 ;
  assign n2621 = n265 & n2620 ;
  assign n2622 = ~n144 & n1697 ;
  assign n2623 = n2621 & n2622 ;
  assign n2624 = n764 & n806 ;
  assign n2625 = ~n1395 & n2624 ;
  assign n2626 = n2625 ^ n1865 ^ 1'b0 ;
  assign n2627 = n202 & ~n1465 ;
  assign n2628 = n1116 & ~n2470 ;
  assign n2629 = n2628 ^ n982 ^ 1'b0 ;
  assign n2630 = n1010 & n2629 ;
  assign n2631 = n440 & n648 ;
  assign n2632 = ~n1152 & n2631 ;
  assign n2633 = n74 & ~n150 ;
  assign n2634 = ~n2632 & n2633 ;
  assign n2635 = n2266 & ~n2287 ;
  assign n2636 = n1865 | n2467 ;
  assign n2637 = n1504 | n2636 ;
  assign n2638 = n365 & ~n758 ;
  assign n2639 = n1984 & n2455 ;
  assign n2640 = n135 | n1749 ;
  assign n2641 = n2640 ^ n787 ^ n588 ;
  assign n2642 = n393 | n870 ;
  assign n2643 = n2642 ^ n1003 ^ 1'b0 ;
  assign n2644 = n2643 ^ n2472 ^ 1'b0 ;
  assign n2645 = n2130 ^ n1742 ^ 1'b0 ;
  assign n2646 = ~n1422 & n2645 ;
  assign n2647 = ~n737 & n2646 ;
  assign n2648 = n1517 ^ n1207 ^ 1'b0 ;
  assign n2649 = n2386 ^ n509 ^ n439 ;
  assign n2650 = n2347 ^ n1434 ^ 1'b0 ;
  assign n2651 = ~n110 & n318 ;
  assign n2652 = n2651 ^ n572 ^ 1'b0 ;
  assign n2653 = n1814 & n2652 ;
  assign n2654 = n721 ^ x11 ^ 1'b0 ;
  assign n2655 = n1847 & n2654 ;
  assign n2656 = n305 & n1318 ;
  assign n2657 = n2655 & ~n2656 ;
  assign n2658 = n2017 ^ n861 ^ n330 ;
  assign n2659 = ~n1714 & n2658 ;
  assign n2660 = n2659 ^ n287 ^ 1'b0 ;
  assign n2661 = n1365 ^ n331 ^ n61 ;
  assign n2662 = n2661 ^ n1307 ^ 1'b0 ;
  assign n2663 = ~n497 & n514 ;
  assign n2664 = n1796 | n2388 ;
  assign n2665 = n2664 ^ n465 ^ 1'b0 ;
  assign n2666 = n1600 & ~n1880 ;
  assign n2667 = n2666 ^ n2236 ^ 1'b0 ;
  assign n2668 = n661 & ~n2667 ;
  assign n2669 = n2668 ^ n1802 ^ 1'b0 ;
  assign n2670 = ~n1325 & n1591 ;
  assign n2671 = n949 & n2615 ;
  assign n2672 = n952 | n1845 ;
  assign n2673 = n1083 & ~n2672 ;
  assign n2674 = n1605 & n2673 ;
  assign n2676 = n2417 ^ n568 ^ 1'b0 ;
  assign n2677 = n1543 & n2676 ;
  assign n2675 = n508 & n1264 ;
  assign n2678 = n2677 ^ n2675 ^ n1336 ;
  assign n2679 = n1407 ^ n649 ^ 1'b0 ;
  assign n2680 = n2679 ^ n475 ^ n96 ;
  assign n2681 = n1033 & n1081 ;
  assign n2682 = ( ~n1177 & n1316 ) | ( ~n1177 & n2681 ) | ( n1316 & n2681 ) ;
  assign n2683 = n1176 ^ n93 ^ 1'b0 ;
  assign n2684 = ~n177 & n2683 ;
  assign n2685 = n2074 ^ n874 ^ 1'b0 ;
  assign n2686 = n2685 ^ n445 ^ 1'b0 ;
  assign n2688 = n682 & ~n965 ;
  assign n2687 = n998 & n1310 ;
  assign n2689 = n2688 ^ n2687 ^ 1'b0 ;
  assign n2690 = n1753 ^ n369 ^ 1'b0 ;
  assign n2691 = n54 & n2690 ;
  assign n2692 = n2691 ^ n1745 ^ 1'b0 ;
  assign n2693 = n667 & ~n2692 ;
  assign n2696 = n619 & n782 ;
  assign n2697 = ~n1092 & n2696 ;
  assign n2694 = n593 ^ n347 ^ 1'b0 ;
  assign n2695 = n2694 ^ n965 ^ 1'b0 ;
  assign n2698 = n2697 ^ n2695 ^ n226 ;
  assign n2703 = n2100 ^ n186 ^ 1'b0 ;
  assign n2704 = n2045 & ~n2703 ;
  assign n2705 = n1949 & n2704 ;
  assign n2699 = n74 | n1198 ;
  assign n2700 = n2699 ^ n322 ^ 1'b0 ;
  assign n2701 = n1469 & ~n2700 ;
  assign n2702 = n521 & ~n2701 ;
  assign n2706 = n2705 ^ n2702 ^ 1'b0 ;
  assign n2707 = ~n205 & n2462 ;
  assign n2708 = n2707 ^ n1548 ^ 1'b0 ;
  assign n2709 = n2708 ^ n1742 ^ 1'b0 ;
  assign n2710 = n695 | n891 ;
  assign n2711 = n1802 | n2710 ;
  assign n2712 = n43 & ~n255 ;
  assign n2713 = ~n2669 & n2712 ;
  assign n2714 = n31 | n140 ;
  assign n2715 = n1967 & ~n2714 ;
  assign n2716 = n2356 | n2715 ;
  assign n2717 = n1644 ^ n1111 ^ 1'b0 ;
  assign n2718 = n79 & ~n2717 ;
  assign n2719 = ~n86 & n2718 ;
  assign n2726 = n362 & n1695 ;
  assign n2720 = n837 & ~n1174 ;
  assign n2721 = n2720 ^ n19 ^ 1'b0 ;
  assign n2723 = n690 ^ n510 ^ n487 ;
  assign n2722 = n858 | n1419 ;
  assign n2724 = n2723 ^ n2722 ^ 1'b0 ;
  assign n2725 = n2721 & n2724 ;
  assign n2727 = n2726 ^ n2725 ^ 1'b0 ;
  assign n2728 = n781 ^ n720 ^ 1'b0 ;
  assign n2729 = n1542 ^ n868 ^ 1'b0 ;
  assign n2730 = n2697 | n2729 ;
  assign n2731 = n347 | n2730 ;
  assign n2732 = n2731 ^ n1229 ^ 1'b0 ;
  assign n2733 = n1955 & ~n2732 ;
  assign n2734 = n2492 ^ n2393 ^ 1'b0 ;
  assign n2735 = n2607 & n2734 ;
  assign n2736 = n189 | n1006 ;
  assign n2743 = n1020 ^ n208 ^ 1'b0 ;
  assign n2744 = ~n52 & n2743 ;
  assign n2745 = n1131 & n2744 ;
  assign n2737 = n376 & n1112 ;
  assign n2738 = n2737 ^ n1182 ^ 1'b0 ;
  assign n2739 = ~n1016 & n2738 ;
  assign n2740 = n475 ^ n169 ^ 1'b0 ;
  assign n2741 = ~n2739 & n2740 ;
  assign n2742 = n2145 & n2741 ;
  assign n2746 = n2745 ^ n2742 ^ 1'b0 ;
  assign n2747 = n1365 & n2373 ;
  assign n2748 = n758 ^ n515 ^ 1'b0 ;
  assign n2749 = n782 & ~n2748 ;
  assign n2750 = n1641 & n2252 ;
  assign n2751 = ~n1416 & n2750 ;
  assign n2752 = n2749 & ~n2751 ;
  assign n2753 = n2747 & n2752 ;
  assign n2754 = ~n475 & n1953 ;
  assign n2755 = n327 & ~n2754 ;
  assign n2756 = n1431 ^ n703 ^ 1'b0 ;
  assign n2757 = n2756 ^ n835 ^ 1'b0 ;
  assign n2758 = ~n1376 & n2757 ;
  assign n2759 = n2023 ^ n340 ^ 1'b0 ;
  assign n2760 = n2758 & n2759 ;
  assign n2761 = n795 | n1800 ;
  assign n2762 = ~n922 & n2761 ;
  assign n2763 = n2760 ^ x1 ^ 1'b0 ;
  assign n2764 = n1122 ^ n40 ^ 1'b0 ;
  assign n2765 = n983 ^ n296 ^ 1'b0 ;
  assign n2766 = ~n2016 & n2765 ;
  assign n2767 = ~n2764 & n2766 ;
  assign n2768 = ~n896 & n1172 ;
  assign n2769 = n2768 ^ n1849 ^ 1'b0 ;
  assign n2770 = n549 | n620 ;
  assign n2771 = ~n1422 & n2451 ;
  assign n2772 = x1 | n2039 ;
  assign n2773 = n1208 ^ n390 ^ n286 ;
  assign n2774 = n1000 | n2773 ;
  assign n2775 = n2774 ^ n1542 ^ 1'b0 ;
  assign n2776 = n1584 ^ n148 ^ 1'b0 ;
  assign n2777 = ~n116 & n2199 ;
  assign n2778 = ~n1179 & n2777 ;
  assign n2779 = ( ~n458 & n1939 ) | ( ~n458 & n2778 ) | ( n1939 & n2778 ) ;
  assign n2780 = n1221 & ~n1900 ;
  assign n2781 = n2780 ^ n1508 ^ 1'b0 ;
  assign n2784 = n453 & n518 ;
  assign n2782 = n1539 ^ n590 ^ 1'b0 ;
  assign n2783 = n89 & n2782 ;
  assign n2785 = n2784 ^ n2783 ^ 1'b0 ;
  assign n2786 = n929 & n2785 ;
  assign n2787 = n2781 & n2786 ;
  assign n2790 = n1219 ^ n224 ^ 1'b0 ;
  assign n2788 = ~n417 & n525 ;
  assign n2789 = n2788 ^ n732 ^ 1'b0 ;
  assign n2791 = n2790 ^ n2789 ^ n1072 ;
  assign n2792 = n1172 ^ n372 ^ 1'b0 ;
  assign n2793 = n438 & ~n2362 ;
  assign n2794 = ~n2792 & n2793 ;
  assign n2795 = n1914 ^ n911 ^ 1'b0 ;
  assign n2796 = n347 | n2795 ;
  assign n2797 = n2796 ^ n798 ^ 1'b0 ;
  assign n2798 = n229 | n2797 ;
  assign n2799 = n1327 & ~n2798 ;
  assign n2800 = n2589 & n2799 ;
  assign n2801 = ~n649 & n2800 ;
  assign n2802 = n2801 ^ n801 ^ 1'b0 ;
  assign n2803 = n641 ^ n349 ^ 1'b0 ;
  assign n2804 = n104 & ~n2803 ;
  assign n2805 = ~n746 & n2804 ;
  assign n2806 = n428 & n914 ;
  assign n2807 = n2806 ^ n387 ^ 1'b0 ;
  assign n2808 = ~n219 & n737 ;
  assign n2809 = ~n1615 & n2808 ;
  assign n2810 = n2809 ^ n445 ^ 1'b0 ;
  assign n2811 = ~n1578 & n2363 ;
  assign n2812 = n2810 & n2811 ;
  assign n2813 = ~n1356 & n2812 ;
  assign n2814 = ~n2697 & n2754 ;
  assign n2815 = ~n1422 & n2814 ;
  assign n2816 = n38 & n1812 ;
  assign n2817 = n2816 ^ n331 ^ 1'b0 ;
  assign n2818 = n1264 & n2817 ;
  assign n2819 = n1216 & ~n2380 ;
  assign n2820 = n2819 ^ n35 ^ 1'b0 ;
  assign n2821 = n2820 ^ n2017 ^ 1'b0 ;
  assign n2822 = ~n920 & n2247 ;
  assign n2823 = ~n1378 & n2045 ;
  assign n2824 = n1845 & n2823 ;
  assign n2825 = n443 & n765 ;
  assign n2826 = ~n126 & n2825 ;
  assign n2827 = n2826 ^ n229 ^ 1'b0 ;
  assign n2828 = n874 | n2827 ;
  assign n2829 = n2140 & ~n2828 ;
  assign n2830 = n2275 & n2829 ;
  assign n2831 = n2824 & n2830 ;
  assign n2834 = ~n1437 & n2095 ;
  assign n2835 = n295 & n2834 ;
  assign n2832 = n441 | n546 ;
  assign n2833 = n2832 ^ n806 ^ 1'b0 ;
  assign n2836 = n2835 ^ n2833 ^ 1'b0 ;
  assign n2837 = n1335 & ~n2836 ;
  assign n2838 = n1837 & ~n2837 ;
  assign n2839 = ~n586 & n2580 ;
  assign n2840 = n2839 ^ n248 ^ 1'b0 ;
  assign n2841 = n2840 ^ n2273 ^ 1'b0 ;
  assign n2842 = n1968 & n2841 ;
  assign n2843 = ~n1607 & n2842 ;
  assign n2844 = n2484 ^ n841 ^ 1'b0 ;
  assign n2845 = n733 & ~n2844 ;
  assign n2846 = n1454 & ~n2638 ;
  assign n2847 = n2778 & n2810 ;
  assign n2848 = n1838 | n2846 ;
  assign n2849 = n2349 ^ n1707 ^ 1'b0 ;
  assign n2850 = ~n619 & n914 ;
  assign n2851 = n2850 ^ n224 ^ 1'b0 ;
  assign n2852 = n2851 ^ n2108 ^ 1'b0 ;
  assign n2853 = n1068 ^ n139 ^ 1'b0 ;
  assign n2854 = n515 & ~n2853 ;
  assign n2855 = n105 & ~n998 ;
  assign n2856 = n1649 ^ n1574 ^ n1551 ;
  assign n2857 = n2856 ^ n45 ^ 1'b0 ;
  assign n2858 = n376 & ~n2361 ;
  assign n2859 = n2858 ^ n1269 ^ 1'b0 ;
  assign n2860 = n2175 & ~n2859 ;
  assign n2861 = n1327 & ~n2104 ;
  assign n2862 = n640 & n2861 ;
  assign n2863 = n1558 ^ n802 ^ 1'b0 ;
  assign n2864 = n736 & ~n2863 ;
  assign n2865 = n1054 & n2864 ;
  assign n2866 = ~n562 & n849 ;
  assign n2867 = n179 & n2866 ;
  assign n2868 = n315 & ~n770 ;
  assign n2869 = n2867 & n2868 ;
  assign n2870 = n433 ^ n43 ^ 1'b0 ;
  assign n2871 = n549 & ~n2870 ;
  assign n2872 = n1331 | n1739 ;
  assign n2873 = n2872 ^ n605 ^ n79 ;
  assign n2874 = n2871 & ~n2873 ;
  assign n2875 = ( n121 & n463 ) | ( n121 & ~n559 ) | ( n463 & ~n559 ) ;
  assign n2876 = ~n122 & n1566 ;
  assign n2886 = n2322 ^ n746 ^ 1'b0 ;
  assign n2887 = n2886 ^ n1191 ^ 1'b0 ;
  assign n2888 = ~n481 & n2887 ;
  assign n2889 = n2888 ^ n1453 ^ 1'b0 ;
  assign n2890 = n434 & n2889 ;
  assign n2882 = n592 | n1845 ;
  assign n2883 = n1818 | n2882 ;
  assign n2884 = ~n1569 & n2883 ;
  assign n2885 = ~n1105 & n2884 ;
  assign n2877 = n1796 ^ n1347 ^ 1'b0 ;
  assign n2878 = n181 | n2877 ;
  assign n2879 = n1284 & ~n2878 ;
  assign n2880 = n880 | n2376 ;
  assign n2881 = n2879 & ~n2880 ;
  assign n2891 = n2890 ^ n2885 ^ n2881 ;
  assign n2892 = n1050 & n1112 ;
  assign n2893 = n2892 ^ n1202 ^ 1'b0 ;
  assign n2895 = ( x3 & n451 ) | ( x3 & n2463 ) | ( n451 & n2463 ) ;
  assign n2894 = n1679 ^ n188 ^ 1'b0 ;
  assign n2896 = n2895 ^ n2894 ^ 1'b0 ;
  assign n2897 = n1260 | n2896 ;
  assign n2898 = n2857 | n2897 ;
  assign n2899 = n2122 | n2898 ;
  assign n2900 = n1765 ^ n991 ^ 1'b0 ;
  assign n2901 = ~n997 & n2865 ;
  assign n2902 = n1994 & n2208 ;
  assign n2903 = n1798 & n2902 ;
  assign n2904 = n854 & n2903 ;
  assign n2905 = n2838 ^ n1418 ^ 1'b0 ;
  assign n2906 = n1871 & ~n2778 ;
  assign n2907 = n1469 & n1540 ;
  assign n2908 = n716 ^ n402 ^ 1'b0 ;
  assign n2909 = ~n671 & n2908 ;
  assign n2910 = n2745 | n2909 ;
  assign n2911 = n489 & ~n896 ;
  assign n2912 = n2181 & n2911 ;
  assign n2913 = n2912 ^ n2252 ^ 1'b0 ;
  assign n2914 = n2910 & ~n2913 ;
  assign n2915 = ( ~n465 & n905 ) | ( ~n465 & n2388 ) | ( n905 & n2388 ) ;
  assign n2916 = n1853 & ~n2915 ;
  assign n2917 = ~n699 & n2238 ;
  assign n2918 = n249 | n798 ;
  assign n2919 = n2918 ^ n2356 ^ 1'b0 ;
  assign n2920 = ( n744 & n880 ) | ( n744 & n1467 ) | ( n880 & n1467 ) ;
  assign n2921 = n2920 ^ n612 ^ 1'b0 ;
  assign n2922 = n2921 ^ n2552 ^ n2100 ;
  assign n2923 = n2205 ^ n1966 ^ 1'b0 ;
  assign n2924 = n2679 ^ n212 ^ 1'b0 ;
  assign n2925 = n1338 & ~n2631 ;
  assign n2926 = n1574 ^ n182 ^ 1'b0 ;
  assign n2927 = n2926 ^ n360 ^ 1'b0 ;
  assign n2928 = n35 & ~n244 ;
  assign n2929 = n2927 & n2928 ;
  assign n2930 = n2351 ^ n2053 ^ n1338 ;
  assign n2931 = n1925 | n2859 ;
  assign n2932 = n810 | n2931 ;
  assign n2935 = n447 ^ n21 ^ 1'b0 ;
  assign n2936 = n459 & n1307 ;
  assign n2937 = n2935 & n2936 ;
  assign n2934 = n2541 ^ n362 ^ 1'b0 ;
  assign n2933 = n1215 | n2832 ;
  assign n2938 = n2937 ^ n2934 ^ n2933 ;
  assign n2939 = n306 ^ n290 ^ 1'b0 ;
  assign n2940 = ~n1584 & n2939 ;
  assign n2941 = ~n152 & n2940 ;
  assign n2942 = n806 & n1079 ;
  assign n2943 = ~n2941 & n2942 ;
  assign n2944 = n1657 ^ n1081 ^ 1'b0 ;
  assign n2945 = ~n922 & n2944 ;
  assign n2946 = n2945 ^ x6 ^ 1'b0 ;
  assign n2947 = n835 & ~n2946 ;
  assign n2948 = ~n290 & n2947 ;
  assign n2949 = ~n47 & n1551 ;
  assign n2950 = n878 & n2949 ;
  assign n2951 = n1167 | n2950 ;
  assign n2952 = ~n630 & n1099 ;
  assign n2953 = n829 & n934 ;
  assign n2954 = n1176 | n2953 ;
  assign n2955 = n2226 | n2730 ;
  assign n2956 = n1146 | n1249 ;
  assign n2957 = n1497 & ~n2956 ;
  assign n2958 = n1933 & n2957 ;
  assign n2959 = n2958 ^ n2199 ^ 1'b0 ;
  assign n2960 = n2104 & ~n2959 ;
  assign n2961 = n963 ^ n936 ^ n703 ;
  assign n2962 = n2961 ^ n867 ^ 1'b0 ;
  assign n2963 = n2872 ^ n839 ^ 1'b0 ;
  assign n2964 = n349 & ~n2963 ;
  assign n2965 = n2962 & n2964 ;
  assign n2966 = n2965 ^ n2480 ^ 1'b0 ;
  assign n2967 = ~n244 & n1493 ;
  assign n2972 = n608 & ~n1014 ;
  assign n2973 = ~x6 & n2972 ;
  assign n2968 = n1101 ^ n973 ^ 1'b0 ;
  assign n2969 = n2968 ^ n738 ^ 1'b0 ;
  assign n2970 = n567 & n2969 ;
  assign n2971 = n2045 & ~n2970 ;
  assign n2974 = n2973 ^ n2971 ^ 1'b0 ;
  assign n2975 = n1551 & ~n2974 ;
  assign n2976 = n1770 | n2975 ;
  assign n2977 = n219 | n2726 ;
  assign n2978 = n2446 & ~n2977 ;
  assign n2979 = n2833 ^ n2282 ^ 1'b0 ;
  assign n2980 = n2283 | n2979 ;
  assign n2981 = n459 & ~n2980 ;
  assign n2982 = n1045 ^ n944 ^ 1'b0 ;
  assign n2983 = n1395 | n2982 ;
  assign n2984 = n1804 ^ n619 ^ 1'b0 ;
  assign n2985 = n1379 & n2984 ;
  assign n2986 = n2985 ^ n152 ^ 1'b0 ;
  assign n2989 = n211 | n1411 ;
  assign n2990 = n237 & ~n1753 ;
  assign n2991 = n2990 ^ n1414 ^ 1'b0 ;
  assign n2992 = n2991 ^ n344 ^ 1'b0 ;
  assign n2993 = n2989 | n2992 ;
  assign n2994 = n2108 & ~n2993 ;
  assign n2987 = n250 & ~n2828 ;
  assign n2988 = n1907 | n2987 ;
  assign n2995 = n2994 ^ n2988 ^ 1'b0 ;
  assign n2996 = n400 ^ n267 ^ 1'b0 ;
  assign n2997 = n1845 | n2996 ;
  assign n2998 = n2995 | n2997 ;
  assign n2999 = n873 ^ n760 ^ n652 ;
  assign n3000 = ( n757 & n1295 ) | ( n757 & ~n1624 ) | ( n1295 & ~n1624 ) ;
  assign n3001 = ( n708 & n2999 ) | ( n708 & ~n3000 ) | ( n2999 & ~n3000 ) ;
  assign n3002 = n2127 ^ n477 ^ 1'b0 ;
  assign n3003 = n3001 & n3002 ;
  assign n3004 = n712 ^ x8 ^ 1'b0 ;
  assign n3005 = n3004 ^ n898 ^ 1'b0 ;
  assign n3006 = n144 & ~n3005 ;
  assign n3007 = n738 & n1863 ;
  assign n3008 = ~n3006 & n3007 ;
  assign n3009 = n619 | n1983 ;
  assign n3010 = n3009 ^ n1645 ^ 1'b0 ;
  assign n3011 = n2202 & n3010 ;
  assign n3012 = n3011 ^ n1289 ^ 1'b0 ;
  assign n3013 = ~n105 & n380 ;
  assign n3014 = n1811 ^ n724 ^ 1'b0 ;
  assign n3015 = n2371 & n3014 ;
  assign n3016 = ~n1286 & n3015 ;
  assign n3017 = n3016 ^ n1505 ^ 1'b0 ;
  assign n3018 = n3009 ^ n1418 ^ 1'b0 ;
  assign n3019 = ~n386 & n3018 ;
  assign n3020 = n3019 ^ n2442 ^ 1'b0 ;
  assign n3021 = ~n182 & n1479 ;
  assign n3022 = n1378 ^ n783 ^ 1'b0 ;
  assign n3023 = n105 & n3022 ;
  assign n3024 = n1130 & n3023 ;
  assign n3025 = ~n3021 & n3024 ;
  assign n3026 = n872 & ~n963 ;
  assign n3027 = n1027 & ~n1295 ;
  assign n3028 = ( ~n43 & n89 ) | ( ~n43 & n875 ) | ( n89 & n875 ) ;
  assign n3029 = ~n1405 & n3028 ;
  assign n3030 = n3029 ^ n924 ^ 1'b0 ;
  assign n3031 = n224 & ~n2130 ;
  assign n3032 = n105 & n3031 ;
  assign n3033 = n3032 ^ n2370 ^ 1'b0 ;
  assign n3034 = n1528 ^ n1335 ^ 1'b0 ;
  assign n3035 = n910 ^ n611 ^ n231 ;
  assign n3036 = n1391 & ~n3035 ;
  assign n3037 = n1065 & n1724 ;
  assign n3038 = n3037 ^ n2941 ^ 1'b0 ;
  assign n3039 = n3036 | n3038 ;
  assign n3040 = n144 & ~n2092 ;
  assign n3041 = ~n1566 & n3040 ;
  assign n3042 = n2395 ^ n1533 ^ x11 ;
  assign n3043 = n2826 | n3042 ;
  assign n3044 = n3043 ^ n277 ^ 1'b0 ;
  assign n3045 = n1588 & ~n1732 ;
  assign n3046 = n1261 | n3045 ;
  assign n3047 = n3046 ^ n415 ^ 1'b0 ;
  assign n3048 = n1420 ^ n474 ^ 1'b0 ;
  assign n3049 = ~n1531 & n3048 ;
  assign n3050 = n3049 ^ n418 ^ 1'b0 ;
  assign n3051 = n796 | n1029 ;
  assign n3052 = n3051 ^ n1044 ^ 1'b0 ;
  assign n3053 = n1271 | n3052 ;
  assign n3054 = n586 & ~n3053 ;
  assign n3055 = ~n777 & n908 ;
  assign n3056 = n633 & n3055 ;
  assign n3057 = n287 | n3056 ;
  assign n3058 = n3057 ^ n1200 ^ 1'b0 ;
  assign n3059 = n655 & ~n2664 ;
  assign n3060 = ~n3058 & n3059 ;
  assign n3061 = n1465 ^ n720 ^ 1'b0 ;
  assign n3062 = ~n3060 & n3061 ;
  assign n3063 = ( ~n2407 & n2791 ) | ( ~n2407 & n3062 ) | ( n2791 & n3062 ) ;
  assign n3064 = n44 & n472 ;
  assign n3065 = n3064 ^ n846 ^ 1'b0 ;
  assign n3066 = n451 & n3065 ;
  assign n3067 = n2571 ^ n598 ^ 1'b0 ;
  assign n3068 = n545 & n3067 ;
  assign n3069 = n560 & ~n1143 ;
  assign n3070 = n3069 ^ n1967 ^ 1'b0 ;
  assign n3077 = n488 & n1578 ;
  assign n3078 = ~n1530 & n3077 ;
  assign n3071 = n88 & n380 ;
  assign n3072 = n477 & ~n578 ;
  assign n3073 = n3072 ^ n1005 ^ n28 ;
  assign n3074 = n1785 & ~n3073 ;
  assign n3075 = ~n3071 & n3074 ;
  assign n3076 = n1136 | n3075 ;
  assign n3079 = n3078 ^ n3076 ^ 1'b0 ;
  assign n3080 = n924 & ~n3079 ;
  assign n3081 = n458 & n2045 ;
  assign n3082 = n3028 ^ n600 ^ 1'b0 ;
  assign n3083 = ( n651 & n3081 ) | ( n651 & n3082 ) | ( n3081 & n3082 ) ;
  assign n3084 = n901 & ~n1369 ;
  assign n3085 = ~n1322 & n3084 ;
  assign n3086 = n3085 ^ n2048 ^ 1'b0 ;
  assign n3087 = n1849 & n2482 ;
  assign n3088 = n3087 ^ n2444 ^ 1'b0 ;
  assign n3089 = n3088 ^ n751 ^ 1'b0 ;
  assign n3090 = n3086 & ~n3089 ;
  assign n3091 = n3011 ^ n1240 ^ 1'b0 ;
  assign n3092 = n372 ^ n229 ^ 1'b0 ;
  assign n3093 = n1337 | n3092 ;
  assign n3094 = n3093 ^ n1334 ^ n1003 ;
  assign n3095 = ~n575 & n800 ;
  assign n3096 = ( n1211 & ~n1306 ) | ( n1211 & n3095 ) | ( ~n1306 & n3095 ) ;
  assign n3097 = ~n688 & n2055 ;
  assign n3098 = n1247 ^ n567 ^ 1'b0 ;
  assign n3099 = n3098 ^ n669 ^ 1'b0 ;
  assign n3100 = n3099 ^ n1036 ^ 1'b0 ;
  assign n3101 = n3097 | n3100 ;
  assign n3107 = n1933 ^ n1186 ^ n340 ;
  assign n3104 = n1861 ^ n924 ^ 1'b0 ;
  assign n3105 = ~n887 & n3104 ;
  assign n3106 = n327 & ~n3105 ;
  assign n3108 = n3107 ^ n3106 ^ n858 ;
  assign n3109 = n3108 ^ n2232 ^ 1'b0 ;
  assign n3102 = n890 | n1650 ;
  assign n3103 = n2348 | n3102 ;
  assign n3110 = n3109 ^ n3103 ^ 1'b0 ;
  assign n3111 = ~n175 & n2583 ;
  assign n3112 = n1497 & n2600 ;
  assign n3113 = n1517 & ~n3008 ;
  assign n3114 = n2781 ^ n1629 ^ n38 ;
  assign n3115 = n896 | n3075 ;
  assign n3117 = n1479 ^ n179 ^ 1'b0 ;
  assign n3118 = n312 | n3117 ;
  assign n3116 = n209 & n1863 ;
  assign n3119 = n3118 ^ n3116 ^ n1691 ;
  assign n3120 = n541 ^ n425 ^ 1'b0 ;
  assign n3121 = n1159 | n3120 ;
  assign n3122 = n1340 & n3121 ;
  assign n3123 = ~n479 & n3099 ;
  assign n3124 = n738 | n1009 ;
  assign n3125 = ~x3 & n1742 ;
  assign n3126 = n1533 | n3125 ;
  assign n3127 = n3126 ^ n2614 ^ 1'b0 ;
  assign n3128 = n96 & n2531 ;
  assign n3129 = n3128 ^ n1504 ^ 1'b0 ;
  assign n3130 = n318 & ~n3129 ;
  assign n3131 = n3130 ^ n1143 ^ 1'b0 ;
  assign n3132 = n466 & ~n1164 ;
  assign n3133 = ~n1007 & n3132 ;
  assign n3138 = n2525 ^ n825 ^ 1'b0 ;
  assign n3139 = n27 & n3138 ;
  assign n3134 = n194 & ~n793 ;
  assign n3135 = ~n547 & n3134 ;
  assign n3136 = n3135 ^ n1291 ^ 1'b0 ;
  assign n3137 = n1891 | n3136 ;
  assign n3140 = n3139 ^ n3137 ^ 1'b0 ;
  assign n3141 = ~n2328 & n2807 ;
  assign n3142 = n567 & n1980 ;
  assign n3143 = ~n261 & n1853 ;
  assign n3144 = n44 ^ x6 ^ 1'b0 ;
  assign n3145 = n28 & n3144 ;
  assign n3146 = ( n159 & n422 ) | ( n159 & n3145 ) | ( n422 & n3145 ) ;
  assign n3147 = n852 | n3146 ;
  assign n3149 = n805 ^ n597 ^ 1'b0 ;
  assign n3150 = ~n445 & n3149 ;
  assign n3151 = n3150 ^ n2780 ^ 1'b0 ;
  assign n3152 = ~n1403 & n3151 ;
  assign n3148 = ~n796 & n1104 ;
  assign n3153 = n3152 ^ n3148 ^ 1'b0 ;
  assign n3154 = x1 & n1969 ;
  assign n3155 = ~n2086 & n3154 ;
  assign n3156 = n160 & ~n3155 ;
  assign n3157 = n3156 ^ n2727 ^ 1'b0 ;
  assign n3158 = n2034 ^ n1299 ^ 1'b0 ;
  assign n3160 = n398 ^ n133 ^ 1'b0 ;
  assign n3161 = n3160 ^ n540 ^ 1'b0 ;
  assign n3162 = n3161 ^ n1750 ^ 1'b0 ;
  assign n3159 = ~n839 & n2968 ;
  assign n3163 = n3162 ^ n3159 ^ 1'b0 ;
  assign n3164 = n706 & ~n780 ;
  assign n3165 = ~n635 & n3164 ;
  assign n3166 = n58 & n1176 ;
  assign n3167 = n1961 ^ n152 ^ 1'b0 ;
  assign n3169 = ~n592 & n668 ;
  assign n3170 = n633 | n3169 ;
  assign n3171 = n3170 ^ n306 ^ 1'b0 ;
  assign n3172 = n3171 ^ n863 ^ 1'b0 ;
  assign n3168 = n49 & ~n458 ;
  assign n3173 = n3172 ^ n3168 ^ 1'b0 ;
  assign n3174 = ( n3166 & ~n3167 ) | ( n3166 & n3173 ) | ( ~n3167 & n3173 ) ;
  assign n3175 = n3174 ^ n3169 ^ 1'b0 ;
  assign n3176 = n3165 | n3175 ;
  assign n3177 = n3176 ^ n1049 ^ 1'b0 ;
  assign n3178 = n2813 & n3177 ;
  assign n3179 = n1042 & n2543 ;
  assign n3181 = n2404 & n3045 ;
  assign n3180 = ~n179 & n2114 ;
  assign n3182 = n3181 ^ n3180 ^ 1'b0 ;
  assign n3183 = n1289 & n3182 ;
  assign n3184 = n197 & n3183 ;
  assign n3185 = n497 & n3184 ;
  assign n3186 = n828 & n3185 ;
  assign n3187 = n2594 ^ n1275 ^ 1'b0 ;
  assign n3188 = n409 ^ n344 ^ 1'b0 ;
  assign n3189 = n33 ^ x4 ^ 1'b0 ;
  assign n3190 = n560 | n3189 ;
  assign n3191 = n2030 & ~n3190 ;
  assign n3192 = ~n523 & n3191 ;
  assign n3193 = n1131 & n3192 ;
  assign n3194 = ~n3188 & n3193 ;
  assign n3195 = n362 | n1911 ;
  assign n3196 = n124 & ~n3195 ;
  assign n3197 = ~n3194 & n3196 ;
  assign n3198 = n2435 ^ n667 ^ 1'b0 ;
  assign n3199 = n246 & n3198 ;
  assign n3200 = ~n415 & n760 ;
  assign n3201 = n3200 ^ n2046 ^ 1'b0 ;
  assign n3202 = n3201 ^ n3194 ^ 1'b0 ;
  assign n3204 = n150 & ~n582 ;
  assign n3205 = ~n1340 & n3204 ;
  assign n3203 = n2067 & ~n3153 ;
  assign n3206 = n3205 ^ n3203 ^ 1'b0 ;
  assign n3207 = n1205 | n1340 ;
  assign n3208 = ~n133 & n1443 ;
  assign n3209 = ~n733 & n3208 ;
  assign n3210 = ( ~n450 & n954 ) | ( ~n450 & n3209 ) | ( n954 & n3209 ) ;
  assign n3211 = n2426 & ~n3210 ;
  assign n3212 = n1596 ^ n199 ^ 1'b0 ;
  assign n3213 = n3212 ^ n878 ^ 1'b0 ;
  assign n3214 = n647 & n2937 ;
  assign n3215 = n3214 ^ n57 ^ 1'b0 ;
  assign n3216 = n2808 & ~n3215 ;
  assign n3217 = n428 & n810 ;
  assign n3218 = n3217 ^ n582 ^ 1'b0 ;
  assign n3219 = n878 & n3218 ;
  assign n3224 = n1403 | n2028 ;
  assign n3222 = ~n423 & n2439 ;
  assign n3223 = n3222 ^ n727 ^ 1'b0 ;
  assign n3220 = n328 & n1788 ;
  assign n3221 = n3220 ^ n1753 ^ 1'b0 ;
  assign n3225 = n3224 ^ n3223 ^ n3221 ;
  assign n3226 = n1322 & n1837 ;
  assign n3227 = n2678 ^ n2349 ^ 1'b0 ;
  assign n3228 = n1823 & n2304 ;
  assign n3229 = n2850 ^ n73 ^ 1'b0 ;
  assign n3230 = ~n387 & n2222 ;
  assign n3231 = n3230 ^ n552 ^ 1'b0 ;
  assign n3233 = n1024 ^ n880 ^ 1'b0 ;
  assign n3232 = n2117 & n2139 ;
  assign n3234 = n3233 ^ n3232 ^ 1'b0 ;
  assign n3235 = ~n3231 & n3234 ;
  assign n3236 = n2773 ^ n390 ^ 1'b0 ;
  assign n3237 = ~n622 & n1505 ;
  assign n3238 = n3237 ^ n1536 ^ 1'b0 ;
  assign n3239 = n1146 & n3238 ;
  assign n3240 = n880 & ~n1490 ;
  assign n3241 = n571 | n614 ;
  assign n3242 = n1396 & ~n3241 ;
  assign n3243 = ~n2451 & n3242 ;
  assign n3244 = n1226 ^ n1016 ^ 1'b0 ;
  assign n3245 = n2580 & n3244 ;
  assign n3246 = n717 & ~n1714 ;
  assign n3247 = n1845 ^ n891 ^ 1'b0 ;
  assign n3248 = ~n3246 & n3247 ;
  assign n3249 = n3245 & n3248 ;
  assign n3250 = n588 & n3249 ;
  assign n3251 = ( n539 & n806 ) | ( n539 & ~n2240 ) | ( n806 & ~n2240 ) ;
  assign n3252 = n2014 ^ n619 ^ 1'b0 ;
  assign n3253 = n3252 ^ n1021 ^ 1'b0 ;
  assign n3254 = n57 & ~n3253 ;
  assign n3256 = n221 & ~n473 ;
  assign n3257 = n3256 ^ n1101 ^ 1'b0 ;
  assign n3255 = n2358 & ~n2472 ;
  assign n3258 = n3257 ^ n3255 ^ 1'b0 ;
  assign n3259 = ( ~n27 & n3254 ) | ( ~n27 & n3258 ) | ( n3254 & n3258 ) ;
  assign n3260 = n1179 & n1194 ;
  assign n3261 = n3260 ^ n2820 ^ 1'b0 ;
  assign n3262 = ( n1291 & ~n1347 ) | ( n1291 & n3261 ) | ( ~n1347 & n3261 ) ;
  assign n3263 = n579 & n877 ;
  assign n3264 = n3263 ^ n801 ^ 1'b0 ;
  assign n3265 = n360 ^ n104 ^ 1'b0 ;
  assign n3266 = n3265 ^ n2366 ^ 1'b0 ;
  assign n3267 = n3264 & n3266 ;
  assign n3268 = n3262 & n3267 ;
  assign n3269 = n45 | n1284 ;
  assign n3270 = n3269 ^ n944 ^ 1'b0 ;
  assign n3271 = n2656 ^ n1285 ^ 1'b0 ;
  assign n3272 = n3183 ^ n1915 ^ n1182 ;
  assign n3273 = n1904 ^ n1020 ^ 1'b0 ;
  assign n3274 = n3272 | n3273 ;
  assign n3275 = n186 | n694 ;
  assign n3276 = n3275 ^ n509 ^ 1'b0 ;
  assign n3277 = n1828 ^ n88 ^ 1'b0 ;
  assign n3278 = n1354 | n3277 ;
  assign n3279 = n205 & n1144 ;
  assign n3280 = ~n213 & n1242 ;
  assign n3281 = ~n3279 & n3280 ;
  assign n3282 = n3281 ^ n2205 ^ 1'b0 ;
  assign n3283 = n2206 & n3282 ;
  assign n3284 = ~n2208 & n3283 ;
  assign n3285 = n3278 | n3284 ;
  assign n3286 = ~n541 & n695 ;
  assign n3287 = ~n1016 & n3286 ;
  assign n3288 = n652 ^ x7 ^ 1'b0 ;
  assign n3289 = n911 & n3288 ;
  assign n3290 = ( n130 & n1182 ) | ( n130 & ~n3289 ) | ( n1182 & ~n3289 ) ;
  assign n3291 = n2065 ^ n1847 ^ 1'b0 ;
  assign n3292 = n311 & n3291 ;
  assign n3293 = ( n940 & ~n2420 ) | ( n940 & n3292 ) | ( ~n2420 & n3292 ) ;
  assign n3294 = n484 & n1312 ;
  assign n3295 = n192 & n3294 ;
  assign n3296 = n415 & ~n3295 ;
  assign n3297 = ~n2371 & n3296 ;
  assign n3298 = n795 | n2989 ;
  assign n3299 = ( n192 & ~n1304 ) | ( n192 & n3298 ) | ( ~n1304 & n3298 ) ;
  assign n3300 = n2139 ^ n1878 ^ n541 ;
  assign n3301 = n331 & ~n3300 ;
  assign n3302 = n3301 ^ n1775 ^ 1'b0 ;
  assign n3303 = n459 & n1912 ;
  assign n3304 = n1413 | n3303 ;
  assign n3305 = n3304 ^ n283 ^ 1'b0 ;
  assign n3306 = n3305 ^ n1845 ^ n415 ;
  assign n3307 = n3306 ^ n1863 ^ 1'b0 ;
  assign n3308 = n2851 ^ n1918 ^ 1'b0 ;
  assign n3309 = ~n342 & n1914 ;
  assign n3310 = n48 & n3309 ;
  assign n3311 = n625 ^ n622 ^ 1'b0 ;
  assign n3312 = n1477 & ~n3311 ;
  assign n3313 = n3310 | n3312 ;
  assign n3314 = n1582 ^ n1280 ^ 1'b0 ;
  assign n3315 = n1325 & ~n3314 ;
  assign n3316 = n1144 ^ n57 ^ 1'b0 ;
  assign n3317 = ~n3315 & n3316 ;
  assign n3318 = n3317 ^ n635 ^ 1'b0 ;
  assign n3319 = n402 ^ n152 ^ 1'b0 ;
  assign n3320 = n3319 ^ n3026 ^ 1'b0 ;
  assign n3322 = ~n352 & n1712 ;
  assign n3323 = ~n1069 & n3322 ;
  assign n3321 = n373 | n2429 ;
  assign n3324 = n3323 ^ n3321 ^ 1'b0 ;
  assign n3325 = ~n1672 & n3324 ;
  assign n3326 = n1164 | n3325 ;
  assign n3327 = n3326 ^ n2322 ^ 1'b0 ;
  assign n3328 = n2151 & ~n3327 ;
  assign n3329 = n2550 ^ n1080 ^ 1'b0 ;
  assign n3330 = ~n1985 & n3329 ;
  assign n3331 = n1004 & ~n2070 ;
  assign n3332 = n2515 & n3331 ;
  assign n3333 = n3332 ^ n255 ^ 1'b0 ;
  assign n3334 = ( n91 & n2473 ) | ( n91 & ~n3333 ) | ( n2473 & ~n3333 ) ;
  assign n3337 = n2460 | n3085 ;
  assign n3338 = n3337 ^ n3137 ^ 1'b0 ;
  assign n3335 = ~n447 & n2524 ;
  assign n3336 = n3265 & ~n3335 ;
  assign n3339 = n3338 ^ n3336 ^ 1'b0 ;
  assign n3340 = n323 | n1622 ;
  assign n3341 = n3340 ^ n1266 ^ 1'b0 ;
  assign n3342 = n2669 ^ n2082 ^ 1'b0 ;
  assign n3343 = ~n666 & n3342 ;
  assign n3344 = ~n1875 & n3343 ;
  assign n3345 = ~n1688 & n3344 ;
  assign n3346 = n2016 | n2019 ;
  assign n3347 = n3346 ^ n227 ^ 1'b0 ;
  assign n3348 = n454 ^ n356 ^ 1'b0 ;
  assign n3349 = n1829 & n3348 ;
  assign n3350 = ( ~n2216 & n2445 ) | ( ~n2216 & n2770 ) | ( n2445 & n2770 ) ;
  assign n3351 = n1526 & n3350 ;
  assign n3352 = n1004 ^ n105 ^ 1'b0 ;
  assign n3353 = n2806 ^ n1918 ^ 1'b0 ;
  assign n3356 = n122 | n362 ;
  assign n3357 = n3356 ^ n110 ^ 1'b0 ;
  assign n3354 = n2061 ^ n808 ^ 1'b0 ;
  assign n3355 = n571 | n3354 ;
  assign n3358 = n3357 ^ n3355 ^ 1'b0 ;
  assign n3360 = n154 | n540 ;
  assign n3361 = n3360 ^ n896 ^ 1'b0 ;
  assign n3359 = n228 | n1845 ;
  assign n3362 = n3361 ^ n3359 ^ 1'b0 ;
  assign n3363 = ~n1466 & n3362 ;
  assign n3364 = n3363 ^ n1454 ^ n1434 ;
  assign n3368 = ~n2131 & n2758 ;
  assign n3369 = n796 & n3368 ;
  assign n3370 = n918 | n3369 ;
  assign n3365 = n1278 & n1561 ;
  assign n3366 = n3365 ^ n2370 ^ 1'b0 ;
  assign n3367 = n3366 ^ n401 ^ 1'b0 ;
  assign n3371 = n3370 ^ n3367 ^ 1'b0 ;
  assign n3372 = ( n188 & n315 ) | ( n188 & ~n400 ) | ( n315 & ~n400 ) ;
  assign n3373 = n2157 ^ n2019 ^ 1'b0 ;
  assign n3374 = n3140 & n3373 ;
  assign n3375 = n1466 ^ n1092 ^ 1'b0 ;
  assign n3376 = n3211 ^ n1202 ^ 1'b0 ;
  assign n3377 = n3066 & n3376 ;
  assign n3378 = n870 & ~n2411 ;
  assign n3379 = n2332 | n2665 ;
  assign n3381 = n3246 ^ n431 ^ 1'b0 ;
  assign n3382 = n135 | n3381 ;
  assign n3380 = n758 & ~n2604 ;
  assign n3383 = n3382 ^ n3380 ^ 1'b0 ;
  assign n3384 = n861 ^ n785 ^ n327 ;
  assign n3385 = n382 & n3384 ;
  assign n3386 = ~n3383 & n3385 ;
  assign n3387 = n1306 | n2279 ;
  assign n3388 = n666 & ~n3387 ;
  assign n3389 = n3388 ^ n793 ^ n782 ;
  assign n3390 = n86 & ~n649 ;
  assign n3391 = ( n541 & n555 ) | ( n541 & n3390 ) | ( n555 & n3390 ) ;
  assign n3392 = n3391 ^ n2070 ^ n1933 ;
  assign n3393 = n1800 ^ n1329 ^ 1'b0 ;
  assign n3394 = n1811 | n1872 ;
  assign n3395 = n3393 | n3394 ;
  assign n3396 = n1264 & n3395 ;
  assign n3397 = n3392 & n3396 ;
  assign n3398 = n1534 | n3218 ;
  assign n3399 = n3398 ^ n915 ^ 1'b0 ;
  assign n3400 = n2644 & n3399 ;
  assign n3401 = n2440 ^ n1947 ^ 1'b0 ;
  assign n3402 = n3400 & n3401 ;
  assign n3403 = n1729 ^ n458 ^ 1'b0 ;
  assign n3404 = n401 & ~n3224 ;
  assign n3405 = n3404 ^ n2799 ^ 1'b0 ;
  assign n3406 = n961 & ~n2987 ;
  assign n3407 = n3406 ^ n1385 ^ 1'b0 ;
  assign n3408 = ~n3405 & n3407 ;
  assign n3409 = n1050 ^ n755 ^ 1'b0 ;
  assign n3410 = n539 & ~n3409 ;
  assign n3411 = ~n67 & n551 ;
  assign n3412 = n3411 ^ n2137 ^ n1411 ;
  assign n3413 = ( n1848 & n3167 ) | ( n1848 & ~n3412 ) | ( n3167 & ~n3412 ) ;
  assign n3414 = n1534 | n3091 ;
  assign n3415 = n1254 & ~n2205 ;
  assign n3416 = n3415 ^ n2042 ^ 1'b0 ;
  assign n3417 = n1313 & n3416 ;
  assign n3418 = n1917 ^ n536 ^ 1'b0 ;
  assign n3419 = n1821 & n2526 ;
  assign n3420 = n3419 ^ n1915 ^ 1'b0 ;
  assign n3421 = n2631 ^ n1967 ^ 1'b0 ;
  assign n3422 = n3420 & ~n3421 ;
  assign n3425 = x11 & n924 ;
  assign n3423 = n2631 ^ n2248 ^ n1745 ;
  assign n3424 = ~n754 & n3423 ;
  assign n3426 = n3425 ^ n3424 ^ n966 ;
  assign n3427 = n2683 & n3426 ;
  assign n3428 = n3427 ^ n3052 ^ 1'b0 ;
  assign n3429 = ( ~n13 & n152 ) | ( ~n13 & n393 ) | ( n152 & n393 ) ;
  assign n3430 = ~n1688 & n1997 ;
  assign n3431 = n3147 & ~n3430 ;
  assign n3432 = ~n401 & n3431 ;
  assign n3434 = ( ~n207 & n459 ) | ( ~n207 & n2356 ) | ( n459 & n2356 ) ;
  assign n3433 = n409 & n1114 ;
  assign n3435 = n3434 ^ n3433 ^ 1'b0 ;
  assign n3436 = n536 & ~n831 ;
  assign n3437 = ~n470 & n3436 ;
  assign n3438 = n3437 ^ n1143 ^ 1'b0 ;
  assign n3439 = n1217 & n3438 ;
  assign n3440 = n799 & ~n1094 ;
  assign n3441 = ~n119 & n3333 ;
  assign n3442 = n1915 ^ n737 ^ 1'b0 ;
  assign n3443 = n2851 & n3442 ;
  assign n3444 = n1945 & ~n2083 ;
  assign n3445 = n980 | n3444 ;
  assign n3446 = n911 & n1083 ;
  assign n3447 = n3446 ^ n1132 ^ 1'b0 ;
  assign n3448 = n3447 ^ n3319 ^ 1'b0 ;
  assign n3449 = n770 | n1432 ;
  assign n3450 = n3449 ^ n2502 ^ 1'b0 ;
  assign n3451 = n3450 ^ n3201 ^ n1962 ;
  assign n3452 = n2257 & ~n2381 ;
  assign n3453 = ~n1804 & n3452 ;
  assign n3454 = n254 & ~n652 ;
  assign n3455 = n3454 ^ n845 ^ 1'b0 ;
  assign n3456 = n2000 ^ n112 ^ 1'b0 ;
  assign n3457 = n1551 & n3456 ;
  assign n3458 = n3457 ^ n536 ^ 1'b0 ;
  assign n3459 = n3455 & n3458 ;
  assign n3464 = n2529 ^ n2381 ^ n525 ;
  assign n3460 = n1010 ^ x10 ^ 1'b0 ;
  assign n3461 = n657 & n3460 ;
  assign n3462 = n2327 & n3461 ;
  assign n3463 = n3040 | n3462 ;
  assign n3465 = n3464 ^ n3463 ^ 1'b0 ;
  assign n3466 = n3176 ^ n2643 ^ n2540 ;
  assign n3467 = ~n506 & n2874 ;
  assign n3468 = n3444 ^ n2403 ^ 1'b0 ;
  assign n3469 = ~n459 & n3468 ;
  assign n3470 = n1234 & n1476 ;
  assign n3471 = n3432 ^ n2821 ^ 1'b0 ;
  assign n3472 = n2023 ^ n239 ^ 1'b0 ;
  assign n3473 = n2155 & n3472 ;
  assign n3474 = n3473 ^ n2193 ^ n1608 ;
  assign n3475 = n255 & ~n1714 ;
  assign n3476 = ~n699 & n2770 ;
  assign n3477 = n3476 ^ n492 ^ 1'b0 ;
  assign n3480 = n1351 ^ n1056 ^ 1'b0 ;
  assign n3481 = n1381 ^ n867 ^ 1'b0 ;
  assign n3482 = ~n3480 & n3481 ;
  assign n3478 = n1546 ^ n197 ^ 1'b0 ;
  assign n3479 = n1546 & n3478 ;
  assign n3483 = n3482 ^ n3479 ^ n2603 ;
  assign n3484 = n2379 ^ n2233 ^ 1'b0 ;
  assign n3485 = n3484 ^ n2186 ^ 1'b0 ;
  assign n3486 = n3261 & ~n3485 ;
  assign n3487 = n327 & ~n1325 ;
  assign n3488 = n3487 ^ n83 ^ 1'b0 ;
  assign n3489 = ( n612 & n2856 ) | ( n612 & n3301 ) | ( n2856 & n3301 ) ;
  assign n3490 = n1582 & n1591 ;
  assign n3491 = n139 | n2619 ;
  assign n3492 = n2527 & ~n3491 ;
  assign n3493 = n3492 ^ n481 ^ 1'b0 ;
  assign n3494 = ~n891 & n3493 ;
  assign n3495 = n2393 ^ n2034 ^ 1'b0 ;
  assign n3496 = ~n1003 & n3495 ;
  assign n3499 = n1126 | n1629 ;
  assign n3500 = n3499 ^ n1984 ^ 1'b0 ;
  assign n3497 = ~n1972 & n2330 ;
  assign n3498 = n3497 ^ n2847 ^ 1'b0 ;
  assign n3501 = n3500 ^ n3498 ^ 1'b0 ;
  assign n3502 = ~n2150 & n2833 ;
  assign n3503 = n2349 ^ n202 ^ 1'b0 ;
  assign n3504 = n1800 & ~n3503 ;
  assign n3505 = n2647 | n3504 ;
  assign n3506 = ~n368 & n2420 ;
  assign n3507 = n108 & n3506 ;
  assign n3508 = ~n680 & n1521 ;
  assign n3509 = n3508 ^ n562 ^ 1'b0 ;
  assign n3510 = n3507 | n3509 ;
  assign n3511 = n1707 ^ n110 ^ 1'b0 ;
  assign n3512 = n2923 | n3511 ;
  assign n3517 = ( n764 & n970 ) | ( n764 & n1880 ) | ( n970 & n1880 ) ;
  assign n3513 = ~n488 & n2225 ;
  assign n3514 = n1173 & ~n2773 ;
  assign n3515 = n3513 | n3514 ;
  assign n3516 = n3515 ^ n2502 ^ 1'b0 ;
  assign n3518 = n3517 ^ n3516 ^ n2828 ;
  assign n3519 = n3518 ^ n57 ^ 1'b0 ;
  assign n3520 = ~n1800 & n3483 ;
  assign n3521 = n3049 ^ n2645 ^ 1'b0 ;
  assign n3522 = n1728 & n3521 ;
  assign n3523 = n2807 & ~n3167 ;
  assign n3524 = n3447 & n3523 ;
  assign n3526 = n1454 ^ n1346 ^ 1'b0 ;
  assign n3525 = n243 | n384 ;
  assign n3527 = n3526 ^ n3525 ^ 1'b0 ;
  assign n3528 = ~n1291 & n3527 ;
  assign n3529 = n3528 ^ n1161 ^ 1'b0 ;
  assign n3530 = n86 & n2885 ;
  assign n3531 = n3530 ^ n390 ^ 1'b0 ;
  assign n3532 = n3531 ^ n683 ^ 1'b0 ;
  assign n3533 = ~n1101 & n3532 ;
  assign n3534 = n2615 ^ n547 ^ 1'b0 ;
  assign n3535 = ~n808 & n3534 ;
  assign n3536 = n633 | n708 ;
  assign n3537 = n2155 ^ n1551 ^ 1'b0 ;
  assign n3538 = n3537 ^ n2413 ^ 1'b0 ;
  assign n3539 = n2998 & ~n3538 ;
  assign n3540 = n1783 ^ n1608 ^ 1'b0 ;
  assign n3541 = n1327 & ~n3540 ;
  assign n3542 = n3160 | n3541 ;
  assign n3543 = n3542 ^ n401 ^ 1'b0 ;
  assign n3544 = n959 & ~n1540 ;
  assign n3545 = ~n1511 & n3544 ;
  assign n3546 = n144 | n474 ;
  assign n3547 = n3546 ^ n1336 ^ 1'b0 ;
  assign n3548 = ( n815 & n914 ) | ( n815 & n3547 ) | ( n914 & n3547 ) ;
  assign n3549 = n3548 ^ n2758 ^ 1'b0 ;
  assign n3550 = n2492 ^ n1428 ^ n1369 ;
  assign n3554 = n2267 ^ n692 ^ 1'b0 ;
  assign n3551 = n1481 & n1943 ;
  assign n3552 = n3551 ^ n3264 ^ 1'b0 ;
  assign n3553 = n1685 | n3552 ;
  assign n3555 = n3554 ^ n3553 ^ 1'b0 ;
  assign n3556 = n3555 ^ n2473 ^ x11 ;
  assign n3557 = n105 & ~n1198 ;
  assign n3558 = n607 & n3557 ;
  assign n3559 = n877 & ~n1865 ;
  assign n3560 = n3559 ^ n2155 ^ 1'b0 ;
  assign n3561 = n3045 ^ n1107 ^ 1'b0 ;
  assign n3562 = n968 | n3561 ;
  assign n3563 = n351 & ~n752 ;
  assign n3564 = n3563 ^ n417 ^ 1'b0 ;
  assign n3565 = ( n220 & n942 ) | ( n220 & ~n1068 ) | ( n942 & ~n1068 ) ;
  assign n3566 = n3060 | n3565 ;
  assign n3567 = ( n3562 & n3564 ) | ( n3562 & n3566 ) | ( n3564 & n3566 ) ;
  assign n3568 = ( ~n854 & n2327 ) | ( ~n854 & n2861 ) | ( n2327 & n2861 ) ;
  assign n3569 = n1284 | n2324 ;
  assign n3570 = n414 ^ n314 ^ 1'b0 ;
  assign n3571 = ~n3569 & n3570 ;
  assign n3572 = ~n1083 & n3571 ;
  assign n3573 = ~n1170 & n2700 ;
  assign n3574 = n282 ^ n183 ^ 1'b0 ;
  assign n3575 = n1790 ^ n1685 ^ 1'b0 ;
  assign n3576 = n738 & ~n3575 ;
  assign n3577 = n1078 ^ n362 ^ 1'b0 ;
  assign n3578 = ~n561 & n1121 ;
  assign n3579 = n3578 ^ n2317 ^ n2128 ;
  assign n3580 = n1756 ^ n1414 ^ 1'b0 ;
  assign n3582 = n1901 | n2082 ;
  assign n3581 = n1838 | n2831 ;
  assign n3583 = n3582 ^ n3581 ^ 1'b0 ;
  assign n3584 = n144 & ~n1099 ;
  assign n3585 = n3584 ^ n2199 ^ 1'b0 ;
  assign n3586 = n1800 & n3585 ;
  assign n3587 = n2347 ^ n2208 ^ n1057 ;
  assign n3588 = n3586 & n3587 ;
  assign n3589 = n2334 ^ n1809 ^ 1'b0 ;
  assign n3590 = n2910 ^ n2762 ^ 1'b0 ;
  assign n3591 = n3589 & ~n3590 ;
  assign n3592 = ~n497 & n2118 ;
  assign n3593 = n612 & ~n1405 ;
  assign n3594 = n3593 ^ n2185 ^ 1'b0 ;
  assign n3595 = n1659 ^ n541 ^ n295 ;
  assign n3596 = n3595 ^ n968 ^ 1'b0 ;
  assign n3597 = ~n3594 & n3596 ;
  assign n3598 = n3592 & ~n3597 ;
  assign n3599 = n1701 & n2648 ;
  assign n3600 = n640 & n1843 ;
  assign n3602 = n2580 ^ n450 ^ 1'b0 ;
  assign n3601 = ~n1993 & n2141 ;
  assign n3603 = n3602 ^ n3601 ^ n3037 ;
  assign n3604 = n2621 ^ n439 ^ 1'b0 ;
  assign n3605 = n1336 & ~n3604 ;
  assign n3606 = n3605 ^ n802 ^ 1'b0 ;
  assign n3607 = n1918 & ~n3606 ;
  assign n3608 = n530 & n576 ;
  assign n3609 = n3608 ^ n2886 ^ 1'b0 ;
  assign n3610 = n43 & n3609 ;
  assign n3611 = n3607 & ~n3610 ;
  assign n3612 = ~n85 & n3477 ;
  assign n3613 = n1499 ^ n1005 ^ 1'b0 ;
  assign n3614 = n3613 ^ n311 ^ 1'b0 ;
  assign n3615 = n1988 ^ n1212 ^ 1'b0 ;
  assign n3616 = n283 & ~n3615 ;
  assign n3617 = ~n434 & n3616 ;
  assign n3618 = n539 | n1779 ;
  assign n3619 = n2275 ^ n1772 ^ n1016 ;
  assign n3620 = n1114 & n3619 ;
  assign n3621 = n135 | n3620 ;
  assign n3622 = n3621 ^ n1378 ^ 1'b0 ;
  assign n3623 = n171 & ~n2252 ;
  assign n3626 = n3265 & ~n3472 ;
  assign n3624 = n2168 | n2735 ;
  assign n3625 = n3624 ^ n559 ^ 1'b0 ;
  assign n3627 = n3626 ^ n3625 ^ 1'b0 ;
  assign n3628 = ~n1170 & n3627 ;
  assign n3629 = n918 & ~n2591 ;
  assign n3630 = n3629 ^ n783 ^ 1'b0 ;
  assign n3631 = n1845 & n3630 ;
  assign n3633 = n3111 ^ n173 ^ 1'b0 ;
  assign n3634 = ~n1189 & n3633 ;
  assign n3632 = n2031 ^ n1550 ^ 1'b0 ;
  assign n3635 = n3634 ^ n3632 ^ n280 ;
  assign n3636 = n3124 & ~n3224 ;
  assign n3637 = n3078 ^ n2070 ^ n976 ;
  assign n3638 = n2614 ^ n2014 ^ 1'b0 ;
  assign n3639 = n3638 ^ n480 ^ 1'b0 ;
  assign n3640 = ~n697 & n3613 ;
  assign n3641 = ~n220 & n3640 ;
  assign n3642 = n3641 ^ n3636 ^ 1'b0 ;
  assign n3643 = n3639 & n3642 ;
  assign n3644 = n439 | n3238 ;
  assign n3645 = ~n307 & n1608 ;
  assign n3646 = n3645 ^ n563 ^ 1'b0 ;
  assign n3647 = n2471 ^ n786 ^ 1'b0 ;
  assign n3648 = n3646 | n3647 ;
  assign n3649 = n3648 ^ n1093 ^ 1'b0 ;
  assign n3650 = n1615 | n3649 ;
  assign n3651 = n1652 & ~n3650 ;
  assign n3652 = ( n894 & ~n3644 ) | ( n894 & n3651 ) | ( ~n3644 & n3651 ) ;
  assign n3654 = n781 & ~n1327 ;
  assign n3655 = n1917 & n3654 ;
  assign n3656 = n2754 & ~n3655 ;
  assign n3657 = ~n829 & n3656 ;
  assign n3653 = n1411 | n3513 ;
  assign n3658 = n3657 ^ n3653 ^ 1'b0 ;
  assign n3659 = n1358 ^ n1099 ^ 1'b0 ;
  assign n3660 = n1004 & ~n3659 ;
  assign n3661 = n2439 ^ n1714 ^ 1'b0 ;
  assign n3662 = n3660 & ~n3661 ;
  assign n3663 = n975 & ~n1546 ;
  assign n3664 = n1560 ^ n625 ^ 1'b0 ;
  assign n3665 = n3664 ^ n412 ^ 1'b0 ;
  assign n3666 = n2417 & n3111 ;
  assign n3667 = n2318 & n3666 ;
  assign n3668 = n3486 | n3667 ;
  assign n3669 = n2233 & ~n2893 ;
  assign n3671 = n2053 ^ n257 ^ 1'b0 ;
  assign n3670 = n850 ^ n798 ^ 1'b0 ;
  assign n3672 = n3671 ^ n3670 ^ 1'b0 ;
  assign n3673 = n874 ^ n362 ^ 1'b0 ;
  assign n3674 = n1009 | n3673 ;
  assign n3675 = n3592 ^ n2784 ^ 1'b0 ;
  assign n3676 = n261 & n3675 ;
  assign n3677 = n1510 ^ n184 ^ 1'b0 ;
  assign n3678 = n2061 & ~n3677 ;
  assign n3679 = n1072 ^ n135 ^ 1'b0 ;
  assign n3680 = n129 & n3679 ;
  assign n3681 = n1464 & n3680 ;
  assign n3682 = ~n3678 & n3681 ;
  assign n3684 = n749 ^ n237 ^ 1'b0 ;
  assign n3685 = n28 | n3684 ;
  assign n3683 = n2570 ^ n227 ^ 1'b0 ;
  assign n3686 = n3685 ^ n3683 ^ 1'b0 ;
  assign n3687 = n3686 ^ n1852 ^ 1'b0 ;
  assign n3688 = n2562 ^ n1609 ^ n1502 ;
  assign n3689 = n3688 ^ n3647 ^ 1'b0 ;
  assign n3690 = n2481 | n3689 ;
  assign n3691 = n1109 ^ n83 ^ 1'b0 ;
  assign n3692 = n1600 & n3145 ;
  assign n3693 = n3692 ^ n1707 ^ 1'b0 ;
  assign n3694 = ~n229 & n3693 ;
  assign n3695 = n3694 ^ n1304 ^ 1'b0 ;
  assign n3696 = n3695 ^ n2922 ^ n94 ;
  assign n3697 = ~n1533 & n1770 ;
  assign n3698 = n3697 ^ n2632 ^ 1'b0 ;
  assign n3699 = n3698 ^ n2101 ^ 1'b0 ;
  assign n3700 = n2492 & ~n3699 ;
  assign n3701 = n745 & n3095 ;
  assign n3702 = n335 ^ n89 ^ 1'b0 ;
  assign n3703 = n3701 & ~n3702 ;
  assign n3706 = n886 | n2273 ;
  assign n3707 = n3706 ^ n579 ^ 1'b0 ;
  assign n3704 = n326 ^ n259 ^ 1'b0 ;
  assign n3705 = n3704 ^ n485 ^ 1'b0 ;
  assign n3708 = n3707 ^ n3705 ^ 1'b0 ;
  assign n3709 = n664 ^ n484 ^ 1'b0 ;
  assign n3710 = n982 | n3709 ;
  assign n3711 = n1745 & ~n3710 ;
  assign n3712 = n1378 & n3711 ;
  assign n3713 = n1267 ^ n725 ^ 1'b0 ;
  assign n3714 = n3712 | n3713 ;
  assign n3715 = n3714 ^ n3232 ^ 1'b0 ;
  assign n3716 = n3715 ^ n1372 ^ 1'b0 ;
  assign n3717 = n1956 ^ n740 ^ 1'b0 ;
  assign n3718 = ~n757 & n3717 ;
  assign n3719 = n342 | n1491 ;
  assign n3720 = n3719 ^ n100 ^ 1'b0 ;
  assign n3721 = n3658 | n3720 ;
  assign n3722 = n828 ^ n634 ^ 1'b0 ;
  assign n3723 = n3721 | n3722 ;
  assign n3724 = ~n2634 & n3135 ;
  assign n3725 = ~n1538 & n2394 ;
  assign n3726 = n61 | n98 ;
  assign n3727 = n472 & ~n1060 ;
  assign n3728 = ~n1152 & n3727 ;
  assign n3729 = ~n2036 & n3728 ;
  assign n3730 = n466 & n3729 ;
  assign n3731 = n2292 ^ n150 ^ 1'b0 ;
  assign n3732 = n254 & n737 ;
  assign n3733 = n2350 ^ n2292 ^ 1'b0 ;
  assign n3734 = n316 | n3733 ;
  assign n3735 = n3732 & n3734 ;
  assign n3736 = n998 & n1865 ;
  assign n3737 = n286 & ~n1724 ;
  assign n3738 = n3737 ^ n1863 ^ 1'b0 ;
  assign n3739 = n1905 & ~n3738 ;
  assign n3740 = ~x11 & n3739 ;
  assign n3741 = n354 | n356 ;
  assign n3742 = n1461 ^ n1394 ^ n373 ;
  assign n3743 = n3742 ^ n2202 ^ 1'b0 ;
  assign n3744 = n3254 & ~n3743 ;
  assign n3745 = n3744 ^ n1432 ^ 1'b0 ;
  assign n3746 = n354 | n2097 ;
  assign n3747 = n3361 | n3746 ;
  assign n3748 = ( n419 & ~n1146 ) | ( n419 & n1434 ) | ( ~n1146 & n1434 ) ;
  assign n3749 = ( n1174 & n1221 ) | ( n1174 & n3748 ) | ( n1221 & n3748 ) ;
  assign n3750 = n820 ^ n492 ^ 1'b0 ;
  assign n3751 = n3749 & n3750 ;
  assign n3752 = ~n3747 & n3751 ;
  assign n3753 = ~n3745 & n3752 ;
  assign n3754 = n1052 & ~n1471 ;
  assign n3755 = n3754 ^ n418 ^ 1'b0 ;
  assign n3756 = n299 | n1533 ;
  assign n3757 = n1420 | n3756 ;
  assign n3758 = n542 & n3693 ;
  assign n3759 = n158 ^ n35 ^ n30 ;
  assign n3760 = n3759 ^ n1535 ^ n447 ;
  assign n3761 = n3760 ^ n2873 ^ 1'b0 ;
  assign n3762 = n1000 ^ n901 ^ n47 ;
  assign n3763 = n3762 ^ n3121 ^ 1'b0 ;
  assign n3764 = n2655 ^ n58 ^ 1'b0 ;
  assign n3765 = n856 | n2776 ;
  assign n3766 = n3764 | n3765 ;
  assign n3767 = n3602 ^ n1742 ^ 1'b0 ;
  assign n3768 = n450 | n3767 ;
  assign n3769 = n3768 ^ n1867 ^ 1'b0 ;
  assign n3770 = n790 & n3769 ;
  assign n3771 = n819 & ~n889 ;
  assign n3772 = n1467 & n3771 ;
  assign n3773 = n3772 ^ n1101 ^ 1'b0 ;
  assign n3774 = ~n296 & n3773 ;
  assign n3775 = n1641 & n3774 ;
  assign n3777 = n1688 ^ n852 ^ 1'b0 ;
  assign n3776 = n1260 | n1682 ;
  assign n3778 = n3777 ^ n3776 ^ 1'b0 ;
  assign n3779 = ( n3770 & ~n3775 ) | ( n3770 & n3778 ) | ( ~n3775 & n3778 ) ;
  assign n3780 = n3766 ^ n582 ^ 1'b0 ;
  assign n3781 = ( n1267 & n1304 ) | ( n1267 & ~n1804 ) | ( n1304 & ~n1804 ) ;
  assign n3782 = n2336 & ~n3031 ;
  assign n3783 = n3781 & n3782 ;
  assign n3789 = n1211 ^ n488 ^ 1'b0 ;
  assign n3786 = ~n414 & n855 ;
  assign n3787 = ~n126 & n3786 ;
  assign n3788 = n1312 | n3787 ;
  assign n3790 = n3789 ^ n3788 ^ n2507 ;
  assign n3791 = n2270 & ~n3790 ;
  assign n3784 = n1656 | n2100 ;
  assign n3785 = n827 | n3784 ;
  assign n3792 = n3791 ^ n3785 ^ 1'b0 ;
  assign n3793 = n2486 ^ n911 ^ 1'b0 ;
  assign n3794 = ~n1329 & n3793 ;
  assign n3796 = n330 & n1242 ;
  assign n3797 = n3796 ^ n474 ^ 1'b0 ;
  assign n3795 = n2143 ^ n1075 ^ 1'b0 ;
  assign n3798 = n3797 ^ n3795 ^ 1'b0 ;
  assign n3799 = n3056 ^ n227 ^ 1'b0 ;
  assign n3800 = n147 & ~n3799 ;
  assign n3801 = n2100 ^ n588 ^ 1'b0 ;
  assign n3802 = n1252 & n3801 ;
  assign n3803 = n1510 & n2706 ;
  assign n3804 = n2816 & n3803 ;
  assign n3805 = ( ~n3800 & n3802 ) | ( ~n3800 & n3804 ) | ( n3802 & n3804 ) ;
  assign n3806 = n347 & ~n3268 ;
  assign n3807 = n3806 ^ n1315 ^ 1'b0 ;
  assign n3808 = ~n1851 & n2535 ;
  assign n3809 = n74 & n3808 ;
  assign n3810 = n3461 ^ n1217 ^ 1'b0 ;
  assign n3811 = n2895 & n3810 ;
  assign n3812 = ~n548 & n3811 ;
  assign n3813 = n445 & n3812 ;
  assign n3816 = n488 ^ n81 ^ 1'b0 ;
  assign n3817 = ~n31 & n3816 ;
  assign n3818 = n1800 & n3817 ;
  assign n3819 = n3818 ^ n508 ^ 1'b0 ;
  assign n3820 = n1186 | n3819 ;
  assign n3821 = n786 & ~n2028 ;
  assign n3822 = n3821 ^ n144 ^ 1'b0 ;
  assign n3823 = ( ~n318 & n3323 ) | ( ~n318 & n3822 ) | ( n3323 & n3822 ) ;
  assign n3824 = n2840 & ~n3823 ;
  assign n3825 = n1728 & n3824 ;
  assign n3826 = ~n3820 & n3825 ;
  assign n3814 = ( n669 & n832 ) | ( n669 & n1845 ) | ( n832 & n1845 ) ;
  assign n3815 = n3327 | n3814 ;
  assign n3827 = n3826 ^ n3815 ^ 1'b0 ;
  assign n3828 = n1563 ^ n1491 ^ n983 ;
  assign n3829 = n2816 ^ n1383 ^ 1'b0 ;
  assign n3830 = n2833 & ~n3829 ;
  assign n3831 = n1842 & n3830 ;
  assign n3832 = n2616 | n3831 ;
  assign n3833 = n3828 | n3832 ;
  assign n3834 = n484 & ~n2189 ;
  assign n3835 = n3834 ^ n1695 ^ 1'b0 ;
  assign n3836 = n563 ^ n159 ^ 1'b0 ;
  assign n3837 = n253 & ~n3836 ;
  assign n3838 = ( n443 & ~n1410 ) | ( n443 & n3837 ) | ( ~n1410 & n3837 ) ;
  assign n3839 = ( n47 & ~n305 ) | ( n47 & n331 ) | ( ~n305 & n331 ) ;
  assign n3840 = n273 & n3839 ;
  assign n3841 = n3838 & ~n3840 ;
  assign n3842 = n3835 & n3841 ;
  assign n3843 = n1159 ^ n800 ^ 1'b0 ;
  assign n3844 = n2256 & ~n3843 ;
  assign n3845 = n3844 ^ n2439 ^ 1'b0 ;
  assign n3846 = n1230 & ~n3845 ;
  assign n3847 = n3846 ^ n2663 ^ 1'b0 ;
  assign n3848 = n3847 ^ n3268 ^ 1'b0 ;
  assign n3850 = n98 | n1709 ;
  assign n3851 = n3850 ^ n2355 ^ 1'b0 ;
  assign n3849 = ~n740 & n1462 ;
  assign n3852 = n3851 ^ n3849 ^ 1'b0 ;
  assign n3853 = n1584 ^ n1344 ^ 1'b0 ;
  assign n3854 = ~n61 & n1295 ;
  assign n3855 = ~n2859 & n3854 ;
  assign n3856 = n3685 & n3855 ;
  assign n3857 = n3566 ^ n1083 ^ 1'b0 ;
  assign n3858 = n877 & n3857 ;
  assign n3859 = n1142 & ~n3111 ;
  assign n3860 = n3858 & n3859 ;
  assign n3861 = n3860 ^ n2132 ^ 1'b0 ;
  assign n3862 = n924 | n3772 ;
  assign n3863 = n3862 ^ n1649 ^ 1'b0 ;
  assign n3864 = n3863 ^ n3707 ^ 1'b0 ;
  assign n3865 = n225 & ~n815 ;
  assign n3866 = n188 & n3865 ;
  assign n3867 = ( n220 & ~n595 ) | ( n220 & n1318 ) | ( ~n595 & n1318 ) ;
  assign n3868 = n2478 ^ n140 ^ 1'b0 ;
  assign n3869 = n3867 & n3868 ;
  assign n3870 = n2838 ^ n2824 ^ 1'b0 ;
  assign n3871 = n3869 & n3870 ;
  assign n3872 = ~n3866 & n3871 ;
  assign n3873 = ~n290 & n3872 ;
  assign n3874 = ~n2054 & n3399 ;
  assign n3875 = ( n3113 & n3122 ) | ( n3113 & n3874 ) | ( n3122 & n3874 ) ;
  assign n3876 = n2201 ^ n1035 ^ 1'b0 ;
  assign n3879 = n609 | n1014 ;
  assign n3880 = n530 | n3879 ;
  assign n3881 = n1010 & n3880 ;
  assign n3877 = n2910 ^ n1398 ^ n347 ;
  assign n3878 = n2841 & ~n3877 ;
  assign n3882 = n3881 ^ n3878 ^ 1'b0 ;
  assign n3883 = n3446 ^ n1571 ^ 1'b0 ;
  assign n3884 = n1419 & n3883 ;
  assign n3885 = n1843 ^ n1690 ^ 1'b0 ;
  assign n3886 = ~n1947 & n1969 ;
  assign n3887 = ( n801 & ~n905 ) | ( n801 & n1363 ) | ( ~n905 & n1363 ) ;
  assign n3888 = n304 | n2238 ;
  assign n3889 = n420 & ~n3888 ;
  assign n3890 = n3887 & ~n3889 ;
  assign n3891 = ~n2087 & n3238 ;
  assign n3892 = ~n228 & n924 ;
  assign n3893 = n3892 ^ n1591 ^ 1'b0 ;
  assign n3894 = n1231 | n1808 ;
  assign n3895 = n2060 ^ n1670 ^ n56 ;
  assign n3896 = n835 & ~n3895 ;
  assign n3897 = n1016 & ~n3665 ;
  assign n3898 = ~n1522 & n2845 ;
  assign n3899 = n3898 ^ n352 ^ 1'b0 ;
  assign n3900 = n615 & ~n2987 ;
  assign n3901 = n3900 ^ n2932 ^ 1'b0 ;
  assign n3902 = ( n880 & ~n1370 ) | ( n880 & n2632 ) | ( ~n1370 & n2632 ) ;
  assign n3903 = n3902 ^ n825 ^ 1'b0 ;
  assign n3904 = ( n1635 & ~n1644 ) | ( n1635 & n2781 ) | ( ~n1644 & n2781 ) ;
  assign n3905 = n1435 ^ n804 ^ 1'b0 ;
  assign n3906 = n2005 & ~n3905 ;
  assign n3907 = n3612 & n3906 ;
  assign n3908 = n470 ^ n218 ^ 1'b0 ;
  assign n3909 = n197 & ~n3908 ;
  assign n3910 = n2917 & n3909 ;
  assign n3911 = ~n3907 & n3910 ;
  assign n3912 = n2638 ^ n1445 ^ n484 ;
  assign n3913 = n411 | n1204 ;
  assign n3914 = n1880 | n2391 ;
  assign n3915 = n1337 & ~n3914 ;
  assign n3916 = n3566 | n3915 ;
  assign n3917 = n1198 & ~n3916 ;
  assign n3919 = ~n271 & n765 ;
  assign n3918 = n3195 ^ n2429 ^ 1'b0 ;
  assign n3920 = n3919 ^ n3918 ^ n2066 ;
  assign n3921 = n1009 & ~n1240 ;
  assign n3922 = n950 & ~n2481 ;
  assign n3923 = ~n3592 & n3922 ;
  assign n3924 = n1918 & ~n3486 ;
  assign n3925 = n1927 ^ n1625 ^ 1'b0 ;
  assign n3926 = ~n366 & n3925 ;
  assign n3927 = ~n2066 & n3926 ;
  assign n3928 = ( n154 & n902 ) | ( n154 & ~n1092 ) | ( n902 & ~n1092 ) ;
  assign n3929 = n2600 ^ n667 ^ 1'b0 ;
  assign n3930 = n298 & ~n3929 ;
  assign n3931 = ~n1759 & n3930 ;
  assign n3932 = n3928 & n3931 ;
  assign n3933 = n1967 ^ n148 ^ 1'b0 ;
  assign n3934 = n3933 ^ n3264 ^ 1'b0 ;
  assign n3935 = ~n155 & n257 ;
  assign n3936 = n3935 ^ n277 ^ 1'b0 ;
  assign n3937 = n3936 ^ n2780 ^ 1'b0 ;
  assign n3942 = n1845 ^ n162 ^ 1'b0 ;
  assign n3943 = n3942 ^ n1351 ^ 1'b0 ;
  assign n3938 = n1237 ^ n126 ^ 1'b0 ;
  assign n3939 = n1320 & ~n3938 ;
  assign n3940 = n2423 & n3939 ;
  assign n3941 = n209 & ~n3940 ;
  assign n3944 = n3943 ^ n3941 ^ 1'b0 ;
  assign n3945 = n1922 | n2137 ;
  assign n3946 = n3945 ^ n751 ^ 1'b0 ;
  assign n3947 = ( n1365 & n2577 ) | ( n1365 & n3946 ) | ( n2577 & n3946 ) ;
  assign n3948 = n3947 ^ n500 ^ 1'b0 ;
  assign n3949 = ~n1987 & n3948 ;
  assign n3950 = n3949 ^ n1871 ^ 1'b0 ;
  assign n3951 = n2929 ^ n1570 ^ 1'b0 ;
  assign n3952 = n1002 & ~n1312 ;
  assign n3953 = n2888 ^ n2852 ^ 1'b0 ;
  assign n3954 = ( n701 & n2063 ) | ( n701 & n2739 ) | ( n2063 & n2739 ) ;
  assign n3955 = n2139 | n3954 ;
  assign n3956 = n1804 ^ n277 ^ 1'b0 ;
  assign n3957 = n340 & ~n3956 ;
  assign n3958 = n3957 ^ n3742 ^ n683 ;
  assign n3959 = n2735 & n3958 ;
  assign n3960 = n2136 ^ n1356 ^ 1'b0 ;
  assign n3961 = ~n2507 & n3960 ;
  assign n3962 = ( n588 & ~n3086 ) | ( n588 & n3961 ) | ( ~n3086 & n3961 ) ;
  assign n3963 = n1438 | n2486 ;
  assign n3964 = n3173 & ~n3963 ;
  assign n3965 = n3964 ^ n2628 ^ 1'b0 ;
  assign n3966 = n2114 | n3965 ;
  assign n3968 = ~x0 & n54 ;
  assign n3969 = n1845 ^ n432 ^ 1'b0 ;
  assign n3970 = n3968 | n3969 ;
  assign n3967 = ~n384 & n1181 ;
  assign n3971 = n3970 ^ n3967 ^ n2298 ;
  assign n3972 = n1469 & ~n2044 ;
  assign n3973 = ~n571 & n1513 ;
  assign n3974 = n3973 ^ n3378 ^ 1'b0 ;
  assign n3975 = n706 & n2000 ;
  assign n3976 = n3527 & ~n3975 ;
  assign n3977 = n600 & n3976 ;
  assign n3978 = n2092 ^ n253 ^ 1'b0 ;
  assign n3979 = n3977 | n3978 ;
  assign n3980 = n2630 & n2927 ;
  assign n3981 = n791 & n1601 ;
  assign n3982 = n398 & ~n3981 ;
  assign n3983 = n1639 & ~n3446 ;
  assign n3984 = ~n1305 & n2653 ;
  assign n3985 = n3984 ^ n3072 ^ 1'b0 ;
  assign n3986 = n1568 | n3453 ;
  assign n3987 = n998 | n3986 ;
  assign n3988 = ~n591 & n1591 ;
  assign n3989 = n3988 ^ n144 ^ 1'b0 ;
  assign n3990 = n3989 ^ n997 ^ 1'b0 ;
  assign n3991 = n3935 ^ n233 ^ 1'b0 ;
  assign n3992 = n3991 ^ n1152 ^ n47 ;
  assign n3993 = n3088 ^ n2556 ^ 1'b0 ;
  assign n3994 = n17 | n331 ;
  assign n3995 = n3994 ^ n1027 ^ 1'b0 ;
  assign n3996 = ( n1716 & n3991 ) | ( n1716 & n3995 ) | ( n3991 & n3995 ) ;
  assign n3997 = n1546 ^ n1449 ^ 1'b0 ;
  assign n3998 = ~n3443 & n3997 ;
  assign n3999 = ~n506 & n3998 ;
  assign n4000 = n3996 & n3999 ;
  assign n4001 = n948 ^ n387 ^ 1'b0 ;
  assign n4002 = n202 | n3851 ;
  assign n4003 = n4002 ^ n3118 ^ 1'b0 ;
  assign n4004 = n3646 | n4003 ;
  assign n4005 = ~n477 & n2113 ;
  assign n4006 = n3757 ^ n3459 ^ 1'b0 ;
  assign n4007 = n1580 ^ n363 ^ 1'b0 ;
  assign n4008 = n4007 ^ n764 ^ 1'b0 ;
  assign n4009 = n162 & ~n4008 ;
  assign n4010 = n3429 & ~n3909 ;
  assign n4011 = n335 | n1024 ;
  assign n4012 = n4011 ^ n533 ^ 1'b0 ;
  assign n4013 = n1832 ^ n120 ^ 1'b0 ;
  assign n4014 = n4013 ^ n2572 ^ 1'b0 ;
  assign n4015 = ( n1109 & n4012 ) | ( n1109 & ~n4014 ) | ( n4012 & ~n4014 ) ;
  assign n4016 = n283 & n946 ;
  assign n4017 = n4016 ^ n1263 ^ 1'b0 ;
  assign n4018 = n1542 ^ n310 ^ 1'b0 ;
  assign n4019 = n3430 & ~n4018 ;
  assign n4020 = n3746 ^ n436 ^ 1'b0 ;
  assign n4021 = n4020 ^ n2219 ^ 1'b0 ;
  assign n4022 = n3105 | n4021 ;
  assign n4023 = n1269 & n2650 ;
  assign n4024 = n3449 & n4023 ;
  assign n4025 = ~n2340 & n4024 ;
  assign n4026 = n1863 ^ n487 ^ 1'b0 ;
  assign n4028 = n3132 ^ n2701 ^ 1'b0 ;
  assign n4027 = n3270 ^ n2114 ^ n1306 ;
  assign n4029 = n4028 ^ n4027 ^ 1'b0 ;
  assign n4030 = ( n2374 & n3109 ) | ( n2374 & n4029 ) | ( n3109 & n4029 ) ;
  assign n4031 = n774 & n2837 ;
  assign n4032 = n4031 ^ n1829 ^ 1'b0 ;
  assign n4033 = n4032 ^ n3695 ^ 1'b0 ;
  assign n4034 = n1574 & n4033 ;
  assign n4035 = n4034 ^ n3245 ^ 1'b0 ;
  assign n4036 = n3258 & n4035 ;
  assign n4037 = ~n2317 & n3280 ;
  assign n4038 = ~n265 & n1668 ;
  assign n4039 = ~n4037 & n4038 ;
  assign n4040 = n1173 ^ n296 ^ 1'b0 ;
  assign n4042 = ~n192 & n798 ;
  assign n4043 = ~n561 & n1313 ;
  assign n4044 = ~n1450 & n4043 ;
  assign n4045 = n4044 ^ n3416 ^ 1'b0 ;
  assign n4046 = ~n4042 & n4045 ;
  assign n4047 = n4046 ^ n2155 ^ 1'b0 ;
  assign n4048 = n1090 & n4047 ;
  assign n4041 = ( n706 & ~n1943 ) | ( n706 & n3388 ) | ( ~n1943 & n3388 ) ;
  assign n4049 = n4048 ^ n4041 ^ 1'b0 ;
  assign n4050 = n4040 & n4049 ;
  assign n4051 = n2694 & ~n3562 ;
  assign n4052 = n1469 & n1548 ;
  assign n4053 = n88 & n4052 ;
  assign n4054 = n1761 & n4053 ;
  assign n4055 = n1946 & n3817 ;
  assign n4056 = n4055 ^ n220 ^ 1'b0 ;
  assign n4057 = n4056 ^ n2103 ^ 1'b0 ;
  assign n4058 = x5 & n4057 ;
  assign n4060 = n2090 ^ n342 ^ 1'b0 ;
  assign n4059 = ( n25 & n2045 ) | ( n25 & n3649 ) | ( n2045 & n3649 ) ;
  assign n4061 = n4060 ^ n4059 ^ n3556 ;
  assign n4062 = n1378 | n1448 ;
  assign n4063 = n1244 & ~n4062 ;
  assign n4064 = ~n106 & n1173 ;
  assign n4065 = n4064 ^ n2103 ^ 1'b0 ;
  assign n4066 = n3560 ^ n423 ^ 1'b0 ;
  assign n4067 = n2536 ^ n1336 ^ 1'b0 ;
  assign n4068 = n3748 & ~n4067 ;
  assign n4069 = n4068 ^ n2735 ^ 1'b0 ;
  assign n4070 = ~n3667 & n4069 ;
  assign n4071 = n543 & n3701 ;
  assign n4072 = ~n4070 & n4071 ;
  assign n4073 = n546 ^ n490 ^ 1'b0 ;
  assign n4074 = n598 & n4073 ;
  assign n4075 = n3384 & ~n4074 ;
  assign n4076 = n1050 ^ n448 ^ 1'b0 ;
  assign n4077 = n150 & n4076 ;
  assign n4078 = ~n2848 & n4077 ;
  assign n4079 = n4078 ^ n584 ^ 1'b0 ;
  assign n4080 = n2673 ^ n1161 ^ 1'b0 ;
  assign n4081 = ( ~n1558 & n1761 ) | ( ~n1558 & n3906 ) | ( n1761 & n3906 ) ;
  assign n4082 = n2621 | n4081 ;
  assign n4083 = n4082 ^ n767 ^ 1'b0 ;
  assign n4084 = ( ~n439 & n885 ) | ( ~n439 & n2852 ) | ( n885 & n2852 ) ;
  assign n4085 = n2533 ^ n1497 ^ n961 ;
  assign n4086 = n4085 ^ n3688 ^ n2374 ;
  assign n4087 = n3892 | n4086 ;
  assign n4088 = ~n1466 & n3224 ;
  assign n4089 = ~n2031 & n4088 ;
  assign n4090 = n3861 ^ n887 ^ 1'b0 ;
  assign n4091 = ~n316 & n3789 ;
  assign n4092 = n4091 ^ n2578 ^ 1'b0 ;
  assign n4093 = n2408 ^ n1033 ^ 1'b0 ;
  assign n4094 = n1729 ^ n858 ^ 1'b0 ;
  assign n4095 = n4094 ^ n1244 ^ 1'b0 ;
  assign n4096 = n4093 | n4095 ;
  assign n4097 = n4096 ^ n3052 ^ 1'b0 ;
  assign n4098 = n612 & ~n3639 ;
  assign n4099 = n2094 ^ n1738 ^ 1'b0 ;
  assign n4100 = ~n1686 & n4099 ;
  assign n4101 = ~n275 & n488 ;
  assign n4104 = ~n286 & n3072 ;
  assign n4102 = n1029 | n2000 ;
  assign n4103 = ~n1089 & n4102 ;
  assign n4105 = n4104 ^ n4103 ^ 1'b0 ;
  assign n4106 = n3384 ^ n2775 ^ n1469 ;
  assign n4107 = n4106 ^ n2641 ^ 1'b0 ;
  assign n4108 = n2661 | n4107 ;
  assign n4109 = n249 & n1987 ;
  assign n4110 = ~n94 & n2721 ;
  assign n4111 = n4109 & n4110 ;
  assign n4112 = n877 | n1911 ;
  assign n4113 = n4112 ^ n505 ^ 1'b0 ;
  assign n4114 = n2881 & ~n3437 ;
  assign n4116 = n502 & n1582 ;
  assign n4115 = n2958 | n3081 ;
  assign n4117 = n4116 ^ n4115 ^ 1'b0 ;
  assign n4118 = n1355 & ~n4117 ;
  assign n4119 = ~n3637 & n4118 ;
  assign n4120 = n2400 ^ n1442 ^ 1'b0 ;
  assign n4121 = n1552 & n4120 ;
  assign n4122 = n4121 ^ n1760 ^ n746 ;
  assign n4123 = n1242 & ~n3232 ;
  assign n4124 = n367 & n782 ;
  assign n4125 = n4124 ^ n179 ^ 1'b0 ;
  assign n4126 = n3962 ^ n3927 ^ 1'b0 ;
  assign n4130 = n318 & n3620 ;
  assign n4131 = n4130 ^ n1694 ^ 1'b0 ;
  assign n4127 = n1418 | n1650 ;
  assign n4128 = n1416 & ~n4127 ;
  assign n4129 = n1112 & n4128 ;
  assign n4132 = n4131 ^ n4129 ^ 1'b0 ;
  assign n4133 = ( n800 & ~n1096 ) | ( n800 & n1930 ) | ( ~n1096 & n1930 ) ;
  assign n4134 = n2765 & ~n4133 ;
  assign n4135 = n4134 ^ n1688 ^ 1'b0 ;
  assign n4137 = n1684 & ~n1928 ;
  assign n4136 = n2028 ^ n1426 ^ 1'b0 ;
  assign n4138 = n4137 ^ n4136 ^ 1'b0 ;
  assign n4139 = ~n754 & n1865 ;
  assign n4145 = n1920 ^ n1637 ^ 1'b0 ;
  assign n4146 = n1445 & ~n4145 ;
  assign n4140 = n582 ^ n105 ^ 1'b0 ;
  assign n4141 = n120 | n4140 ;
  assign n4142 = n967 & ~n4141 ;
  assign n4143 = n4142 ^ n432 ^ 1'b0 ;
  assign n4144 = n1226 & n4143 ;
  assign n4147 = n4146 ^ n4144 ^ 1'b0 ;
  assign n4150 = n1062 ^ n541 ^ 1'b0 ;
  assign n4151 = n781 & n4150 ;
  assign n4152 = n2888 & n4151 ;
  assign n4153 = ~n2754 & n4152 ;
  assign n4148 = n2190 ^ n288 ^ 1'b0 ;
  assign n4149 = n4148 ^ n2504 ^ n1343 ;
  assign n4154 = n4153 ^ n4149 ^ 1'b0 ;
  assign n4155 = n40 & n48 ;
  assign n4162 = n3023 ^ n506 ^ 1'b0 ;
  assign n4156 = ~n1260 & n3139 ;
  assign n4157 = n4156 ^ n451 ^ 1'b0 ;
  assign n4158 = n849 & ~n1143 ;
  assign n4159 = n4158 ^ n2347 ^ 1'b0 ;
  assign n4160 = n4159 ^ n3967 ^ 1'b0 ;
  assign n4161 = n4157 & ~n4160 ;
  assign n4163 = n4162 ^ n4161 ^ 1'b0 ;
  assign n4164 = n108 & ~n1305 ;
  assign n4165 = n2820 | n4164 ;
  assign n4166 = n484 | n4165 ;
  assign n4167 = ~n2510 & n4133 ;
  assign n4168 = ~n762 & n1469 ;
  assign n4169 = x7 & ~n4017 ;
  assign n4170 = n4168 & n4169 ;
  assign n4171 = n1083 ^ n390 ^ 1'b0 ;
  assign n4172 = n949 ^ n551 ^ 1'b0 ;
  assign n4173 = n694 & n4172 ;
  assign n4174 = n3223 & ~n4173 ;
  assign n4175 = n1569 & n2519 ;
  assign n4176 = ~n1289 & n4175 ;
  assign n4177 = n4176 ^ n374 ^ 1'b0 ;
  assign n4178 = n3118 | n4177 ;
  assign n4179 = ~n1245 & n4030 ;
  assign n4181 = n1558 & ~n3361 ;
  assign n4182 = n4181 ^ n737 ^ 1'b0 ;
  assign n4180 = ~n33 & n1403 ;
  assign n4183 = n4182 ^ n4180 ^ n2309 ;
  assign n4184 = n984 & ~n995 ;
  assign n4185 = ~n447 & n4184 ;
  assign n4186 = n3476 ^ n677 ^ 1'b0 ;
  assign n4187 = ~n1930 & n4186 ;
  assign n4189 = n2253 ^ n1852 ^ 1'b0 ;
  assign n4188 = n400 & n2016 ;
  assign n4190 = n4189 ^ n4188 ^ 1'b0 ;
  assign n4191 = n1716 | n4190 ;
  assign n4192 = n1353 | n3647 ;
  assign n4193 = n3949 | n4192 ;
  assign n4194 = ( n27 & ~n2131 ) | ( n27 & n3093 ) | ( ~n2131 & n3093 ) ;
  assign n4195 = n2520 ^ n1605 ^ 1'b0 ;
  assign n4196 = n120 & ~n140 ;
  assign n4197 = ~n4195 & n4196 ;
  assign n4198 = n3464 | n4197 ;
  assign n4199 = n1707 | n4198 ;
  assign n4200 = n1240 ^ n277 ^ 1'b0 ;
  assign n4201 = n582 & n4200 ;
  assign n4202 = n3298 ^ n3101 ^ 1'b0 ;
  assign n4203 = ~n1560 & n4202 ;
  assign n4204 = ~n3665 & n4203 ;
  assign n4205 = n4204 ^ n3141 ^ 1'b0 ;
  assign n4206 = n2321 ^ n1205 ^ n219 ;
  assign n4207 = n770 & n3147 ;
  assign n4208 = n732 & n1462 ;
  assign n4209 = n3818 ^ n707 ^ 1'b0 ;
  assign n4210 = n4208 & n4209 ;
  assign n4211 = ~n4207 & n4210 ;
  assign n4212 = n578 & ~n1655 ;
  assign n4213 = n4212 ^ n3805 ^ 1'b0 ;
  assign n4214 = n826 ^ n810 ^ 1'b0 ;
  assign n4215 = n2155 ^ n1182 ^ 1'b0 ;
  assign n4216 = n630 | n694 ;
  assign n4217 = ~n1280 & n4216 ;
  assign n4218 = ~n821 & n4217 ;
  assign n4219 = n344 | n4218 ;
  assign n4220 = n3414 & ~n4219 ;
  assign n4221 = n625 & n961 ;
  assign n4222 = n439 & ~n1252 ;
  assign n4223 = n1525 & n2656 ;
  assign n4224 = n4222 & n4223 ;
  assign n4225 = n2771 | n4224 ;
  assign n4226 = n2267 & ~n4225 ;
  assign n4227 = ~n973 & n2145 ;
  assign n4228 = ~n555 & n4227 ;
  assign n4229 = n4228 ^ n1809 ^ 1'b0 ;
  assign n4230 = n4229 ^ n2394 ^ 1'b0 ;
  assign n4231 = ~n445 & n4230 ;
  assign n4232 = n1035 & n1383 ;
  assign n4233 = n4232 ^ n130 ^ 1'b0 ;
  assign n4234 = n3484 & ~n4233 ;
  assign n4235 = ~n56 & n1849 ;
  assign n4236 = n649 & ~n2507 ;
  assign n4237 = n2363 & n3562 ;
  assign n4238 = ~n568 & n4237 ;
  assign n4239 = ~n1508 & n2571 ;
  assign n4240 = ~n1422 & n4239 ;
  assign n4241 = n1295 & ~n2502 ;
  assign n4242 = n1267 & n1283 ;
  assign n4243 = n661 & n4242 ;
  assign n4244 = n4243 ^ n4145 ^ 1'b0 ;
  assign n4245 = ( n162 & n1075 ) | ( n162 & ~n2046 ) | ( n1075 & ~n2046 ) ;
  assign n4246 = ( n572 & n1830 ) | ( n572 & ~n2326 ) | ( n1830 & ~n2326 ) ;
  assign n4247 = n4245 & n4246 ;
  assign n4248 = ~n4244 & n4247 ;
  assign n4249 = n2787 ^ n2077 ^ 1'b0 ;
  assign n4250 = n192 & ~n4249 ;
  assign n4251 = ~n758 & n1688 ;
  assign n4252 = n828 & n2871 ;
  assign n4254 = n249 & ~n2145 ;
  assign n4253 = ~n239 & n3502 ;
  assign n4255 = n4254 ^ n4253 ^ 1'b0 ;
  assign n4256 = n2994 & n4255 ;
  assign n4257 = ( ~n356 & n1078 ) | ( ~n356 & n1700 ) | ( n1078 & n1700 ) ;
  assign n4258 = n666 | n1023 ;
  assign n4259 = n2205 & ~n4258 ;
  assign n4260 = n362 & ~n4259 ;
  assign n4261 = n2184 | n2682 ;
  assign n4262 = n2732 ^ n1971 ^ 1'b0 ;
  assign n4263 = n839 & n4262 ;
  assign n4264 = n4263 ^ n2828 ^ n1675 ;
  assign n4266 = n2050 ^ n946 ^ 1'b0 ;
  assign n4267 = ~n2070 & n4266 ;
  assign n4265 = n690 | n1655 ;
  assign n4268 = n4267 ^ n4265 ^ 1'b0 ;
  assign n4269 = n3766 | n3852 ;
  assign n4270 = n3514 ^ n3124 ^ 1'b0 ;
  assign n4271 = n4050 ^ n2087 ^ n914 ;
  assign n4272 = n345 & n1516 ;
  assign n4273 = n4272 ^ n259 ^ 1'b0 ;
  assign n4274 = n4273 ^ n620 ^ 1'b0 ;
  assign n4275 = n768 & ~n1908 ;
  assign n4276 = ~n4214 & n4275 ;
  assign n4277 = n3482 ^ n1016 ^ 1'b0 ;
  assign n4278 = ~n1434 & n4277 ;
  assign n4279 = n3566 ^ n3045 ^ n2078 ;
  assign n4280 = ( ~n316 & n668 ) | ( ~n316 & n2219 ) | ( n668 & n2219 ) ;
  assign n4281 = n4280 ^ n4082 ^ 1'b0 ;
  assign n4282 = n1830 | n4281 ;
  assign n4283 = n149 | n4282 ;
  assign n4284 = n4283 ^ n3264 ^ 1'b0 ;
  assign n4285 = n1486 ^ n1189 ^ 1'b0 ;
  assign n4286 = ~n40 & n171 ;
  assign n4287 = ~n52 & n4286 ;
  assign n4288 = n1705 & ~n2236 ;
  assign n4289 = n4287 & n4288 ;
  assign n4290 = n3282 ^ n1798 ^ 1'b0 ;
  assign n4291 = ~n2815 & n3949 ;
  assign n4292 = n4291 ^ n2661 ^ 1'b0 ;
  assign n4293 = n4290 | n4292 ;
  assign n4294 = n4293 ^ n1625 ^ 1'b0 ;
  assign n4295 = n2104 ^ n1141 ^ 1'b0 ;
  assign n4296 = n498 ^ n362 ^ 1'b0 ;
  assign n4297 = n142 | n2130 ;
  assign n4298 = ( n1150 & n3539 ) | ( n1150 & n4297 ) | ( n3539 & n4297 ) ;
  assign n4299 = ~n2922 & n4298 ;
  assign n4300 = n846 ^ n754 ^ 1'b0 ;
  assign n4301 = n4300 ^ n1845 ^ 1'b0 ;
  assign n4302 = n4116 & ~n4301 ;
  assign n4303 = n2132 & ~n2247 ;
  assign n4304 = ~n4302 & n4303 ;
  assign n4305 = n3153 & n4304 ;
  assign n4306 = n4305 ^ n3961 ^ 1'b0 ;
  assign n4307 = n1460 | n4306 ;
  assign n4308 = n697 | n4307 ;
  assign n4309 = n4308 ^ n3280 ^ 1'b0 ;
  assign n4310 = n409 & n2368 ;
  assign n4311 = n4310 ^ n1023 ^ 1'b0 ;
  assign n4312 = n4311 ^ n3297 ^ 1'b0 ;
  assign n4313 = ( n625 & ~n911 ) | ( n625 & n2645 ) | ( ~n911 & n2645 ) ;
  assign n4314 = n2934 ^ n2000 ^ 1'b0 ;
  assign n4315 = ~n2604 & n4314 ;
  assign n4316 = n1121 & n2102 ;
  assign n4317 = n4316 ^ n349 ^ 1'b0 ;
  assign n4318 = n1178 ^ n1094 ^ 1'b0 ;
  assign n4319 = n1464 | n4318 ;
  assign n4320 = n1159 | n4319 ;
  assign n4321 = n106 & ~n4320 ;
  assign n4322 = n901 | n4321 ;
  assign n4323 = n447 & ~n880 ;
  assign n4324 = n4323 ^ x8 ^ 1'b0 ;
  assign n4325 = ( ~n3313 & n3496 ) | ( ~n3313 & n3774 ) | ( n3496 & n3774 ) ;
  assign n4326 = n997 ^ n578 ^ n318 ;
  assign n4327 = n1190 ^ n1090 ^ 1'b0 ;
  assign n4328 = ~n35 & n2166 ;
  assign n4329 = n4328 ^ n4284 ^ n2789 ;
  assign n4330 = n2505 ^ n1843 ^ 1'b0 ;
  assign n4331 = ~n117 & n4330 ;
  assign n4332 = n3355 & n4331 ;
  assign n4333 = n542 ^ n27 ^ 1'b0 ;
  assign n4334 = n1257 | n4333 ;
  assign n4335 = n3271 & ~n4334 ;
  assign n4336 = n3349 ^ n967 ^ 1'b0 ;
  assign n4337 = n459 | n4336 ;
  assign n4338 = n4337 ^ n2883 ^ 1'b0 ;
  assign n4339 = n3520 ^ n3179 ^ 1'b0 ;
  assign n4340 = n3006 & ~n4339 ;
  assign n4341 = n366 & ~n942 ;
  assign n4342 = n3909 & n4341 ;
  assign n4343 = ~n4340 & n4342 ;
  assign n4344 = n2796 ^ n1637 ^ 1'b0 ;
  assign n4345 = n4344 ^ n409 ^ 1'b0 ;
  assign n4346 = n2779 | n4345 ;
  assign n4347 = n673 & n2632 ;
  assign n4348 = n2313 ^ n1370 ^ n339 ;
  assign n4349 = n2589 ^ n2163 ^ 1'b0 ;
  assign n4350 = n2210 ^ n1198 ^ 1'b0 ;
  assign n4351 = n709 & n1620 ;
  assign n4352 = n1471 ^ x7 ^ 1'b0 ;
  assign n4353 = n4351 | n4352 ;
  assign n4354 = n2458 ^ n182 ^ 1'b0 ;
  assign n4355 = n2077 & ~n4354 ;
  assign n4356 = n793 | n1806 ;
  assign n4357 = n1123 & ~n4356 ;
  assign n4359 = n2816 ^ n298 ^ 1'b0 ;
  assign n4360 = n635 & n4359 ;
  assign n4358 = ~n1201 & n2472 ;
  assign n4361 = n4360 ^ n4358 ^ 1'b0 ;
  assign n4362 = ~n2403 & n4104 ;
  assign n4363 = ~n2141 & n4362 ;
  assign n4364 = n4363 ^ n3187 ^ n1065 ;
  assign n4365 = n2338 ^ n1857 ^ 1'b0 ;
  assign n4366 = n4365 ^ n3225 ^ 1'b0 ;
  assign n4367 = n754 | n1386 ;
  assign n4369 = n1810 & ~n2743 ;
  assign n4368 = n2635 ^ n2580 ^ 1'b0 ;
  assign n4370 = n4369 ^ n4368 ^ n3179 ;
  assign n4371 = n1625 & n2502 ;
  assign n4372 = n4371 ^ n3447 ^ 1'b0 ;
  assign n4373 = ~n1953 & n3006 ;
  assign n4374 = ~n2873 & n4373 ;
  assign n4375 = n4374 ^ n3582 ^ 1'b0 ;
  assign n4376 = n312 | n4375 ;
  assign n4377 = n3290 & n4376 ;
  assign n4378 = n3221 ^ n2691 ^ 1'b0 ;
  assign n4379 = n778 & ~n2094 ;
  assign n4380 = n2688 | n4379 ;
  assign n4381 = n521 | n755 ;
  assign n4382 = n2004 | n3977 ;
  assign n4383 = n4382 ^ n229 ^ 1'b0 ;
  assign n4384 = n1208 | n4383 ;
  assign n4385 = n488 & n2628 ;
  assign n4386 = n4385 ^ n1337 ^ 1'b0 ;
  assign n4387 = n489 & n1124 ;
  assign n4388 = n959 & n4387 ;
  assign n4389 = n1189 & ~n1853 ;
  assign n4390 = ~n1288 & n1313 ;
  assign n4391 = ~n840 & n4390 ;
  assign n4392 = ~n987 & n4185 ;
  assign n4393 = n4173 ^ n2806 ^ 1'b0 ;
  assign n4394 = n2811 | n4393 ;
  assign n4395 = ~n3254 & n4394 ;
  assign n4399 = n755 ^ n110 ^ 1'b0 ;
  assign n4400 = n4399 ^ n2082 ^ 1'b0 ;
  assign n4396 = n347 & n502 ;
  assign n4397 = n3049 & ~n4396 ;
  assign n4398 = ~n1761 & n4397 ;
  assign n4401 = n4400 ^ n4398 ^ 1'b0 ;
  assign n4402 = n3327 | n4401 ;
  assign n4403 = ( n1240 & ~n1743 ) | ( n1240 & n4070 ) | ( ~n1743 & n4070 ) ;
  assign n4404 = n241 & ~n822 ;
  assign n4405 = n4404 ^ n76 ^ 1'b0 ;
  assign n4406 = n4405 ^ n2765 ^ n2381 ;
  assign n4407 = n33 | n2694 ;
  assign n4408 = n3544 ^ n1361 ^ 1'b0 ;
  assign n4409 = ~n2218 & n4408 ;
  assign n4410 = n2810 ^ n223 ^ 1'b0 ;
  assign n4411 = n2607 ^ n823 ^ 1'b0 ;
  assign n4412 = ~n1331 & n3547 ;
  assign n4413 = n4412 ^ n568 ^ 1'b0 ;
  assign n4414 = n237 & ~n4413 ;
  assign n4415 = n4411 & n4414 ;
  assign n4416 = n1318 & ~n2638 ;
  assign n4417 = n129 & ~n4269 ;
  assign n4418 = ~n2148 & n4417 ;
  assign n4419 = n1395 ^ n552 ^ 1'b0 ;
  assign n4420 = ( n746 & n3734 ) | ( n746 & ~n4419 ) | ( n3734 & ~n4419 ) ;
  assign n4421 = n345 & ~n1170 ;
  assign n4422 = n4421 ^ n707 ^ 1'b0 ;
  assign n4423 = n2387 ^ n2108 ^ 1'b0 ;
  assign n4424 = n1278 & ~n1994 ;
  assign n4425 = ~n4423 & n4424 ;
  assign n4426 = n1914 ^ n1329 ^ 1'b0 ;
  assign n4427 = ~n474 & n4426 ;
  assign n4428 = n3061 | n4427 ;
  assign n4429 = n3840 ^ n3766 ^ n2566 ;
  assign n4430 = n4429 ^ n2108 ^ 1'b0 ;
  assign n4431 = n4430 ^ n472 ^ 1'b0 ;
  assign n4432 = n2098 & n4431 ;
  assign n4433 = n244 | n3082 ;
  assign n4434 = n76 & n169 ;
  assign n4435 = n4433 & ~n4434 ;
  assign n4436 = n2508 ^ n76 ^ 1'b0 ;
  assign n4437 = n3405 | n3913 ;
  assign n4438 = n3573 & ~n4437 ;
  assign n4439 = n2340 ^ n1534 ^ 1'b0 ;
  assign n4440 = n1165 & n4439 ;
  assign n4441 = n982 & n4440 ;
  assign n4442 = n4441 ^ n57 ^ 1'b0 ;
  assign n4443 = ~n1060 & n3851 ;
  assign n4444 = n4443 ^ n1911 ^ 1'b0 ;
  assign n4445 = ~n2824 & n4444 ;
  assign n4446 = n20 & n4445 ;
  assign n4447 = n2448 ^ n1922 ^ 1'b0 ;
  assign n4448 = ( n1090 & n1392 ) | ( n1090 & ~n1673 ) | ( n1392 & ~n1673 ) ;
  assign n4449 = n3533 ^ n214 ^ 1'b0 ;
  assign n4450 = n1641 & n2837 ;
  assign n4451 = n1956 & n4450 ;
  assign n4452 = n3805 ^ n3026 ^ n851 ;
  assign n4453 = n1939 | n2700 ;
  assign n4454 = n4452 | n4453 ;
  assign n4455 = n1956 | n4454 ;
  assign n4456 = n3088 & n3998 ;
  assign n4457 = n4456 ^ n465 ^ 1'b0 ;
  assign n4458 = ~n136 & n2682 ;
  assign n4459 = n4458 ^ n1460 ^ 1'b0 ;
  assign n4460 = n755 | n841 ;
  assign n4464 = ~n342 & n954 ;
  assign n4462 = ~n333 & n1912 ;
  assign n4463 = n4462 ^ n2413 ^ 1'b0 ;
  assign n4465 = n4464 ^ n4463 ^ 1'b0 ;
  assign n4466 = n243 | n4465 ;
  assign n4461 = ~n1036 & n1442 ;
  assign n4467 = n4466 ^ n4461 ^ 1'b0 ;
  assign n4468 = n1385 | n4467 ;
  assign n4469 = n4460 | n4468 ;
  assign n4470 = n2756 | n4469 ;
  assign n4475 = ~n518 & n1128 ;
  assign n4476 = n4475 ^ n218 ^ 1'b0 ;
  assign n4474 = ~n154 & n3021 ;
  assign n4477 = n4476 ^ n4474 ^ 1'b0 ;
  assign n4471 = n144 & n1121 ;
  assign n4472 = n4471 ^ n712 ^ 1'b0 ;
  assign n4473 = ~n347 & n4472 ;
  assign n4478 = n4477 ^ n4473 ^ n4419 ;
  assign n4479 = n2117 | n4478 ;
  assign n4480 = n3726 ^ n1069 ^ 1'b0 ;
  assign n4481 = n3902 ^ n1783 ^ n1398 ;
  assign n4482 = n2030 | n3789 ;
  assign n4483 = n950 | n4482 ;
  assign n4484 = ~n4476 & n4483 ;
  assign n4485 = ~n4138 & n4484 ;
  assign n4486 = n1455 & n2236 ;
  assign n4487 = n1925 ^ n1506 ^ n924 ;
  assign n4488 = n4016 ^ n373 ^ 1'b0 ;
  assign n4489 = n43 & ~n4488 ;
  assign n4490 = n4489 ^ n2794 ^ 1'b0 ;
  assign n4491 = n4487 | n4490 ;
  assign n4492 = ~n2912 & n4461 ;
  assign n4493 = ~n547 & n1887 ;
  assign n4494 = n312 | n4493 ;
  assign n4495 = n4494 ^ n753 ^ 1'b0 ;
  assign n4496 = n901 ^ n605 ^ 1'b0 ;
  assign n4497 = n88 | n481 ;
  assign n4498 = ~n1073 & n2833 ;
  assign n4499 = n4498 ^ n1007 ^ 1'b0 ;
  assign n4500 = n2317 & n3140 ;
  assign n4501 = n4500 ^ n1653 ^ 1'b0 ;
  assign n4502 = n1518 & ~n2859 ;
  assign n4503 = n4502 ^ n1825 ^ 1'b0 ;
  assign n4504 = n1695 | n4503 ;
  assign n4505 = n776 & n4504 ;
  assign n4506 = n3822 ^ n1441 ^ n406 ;
  assign n4510 = n3744 ^ n3657 ^ 1'b0 ;
  assign n4511 = n195 & n4510 ;
  assign n4507 = n2862 ^ n551 ^ 1'b0 ;
  assign n4508 = n4002 & n4507 ;
  assign n4509 = n2101 & n4508 ;
  assign n4512 = n4511 ^ n4509 ^ 1'b0 ;
  assign n4514 = ~n326 & n3126 ;
  assign n4515 = n4514 ^ n694 ^ 1'b0 ;
  assign n4516 = n3933 ^ n3006 ^ 1'b0 ;
  assign n4517 = ~n4515 & n4516 ;
  assign n4513 = n305 | n2097 ;
  assign n4518 = n4517 ^ n4513 ^ 1'b0 ;
  assign n4523 = n873 | n961 ;
  assign n4519 = n2730 ^ n808 ^ 1'b0 ;
  assign n4520 = n4519 ^ n3457 ^ 1'b0 ;
  assign n4521 = n2783 & ~n4520 ;
  assign n4522 = n2155 | n4521 ;
  assign n4524 = n4523 ^ n4522 ^ 1'b0 ;
  assign n4525 = ~n3858 & n4524 ;
  assign n4526 = n3580 | n3953 ;
  assign n4527 = n511 ^ n225 ^ 1'b0 ;
  assign n4528 = n1518 & ~n4527 ;
  assign n4529 = n4528 ^ n539 ^ 1'b0 ;
  assign n4530 = n842 | n4529 ;
  assign n4531 = n2924 & ~n4530 ;
  assign n4532 = ~n1596 & n4531 ;
  assign n4533 = n1438 & ~n2332 ;
  assign n4534 = ~n826 & n1090 ;
  assign n4535 = ~n4533 & n4534 ;
  assign n4536 = n183 & n3704 ;
  assign n4537 = n1510 | n4536 ;
  assign n4540 = n4351 ^ n1966 ^ 1'b0 ;
  assign n4541 = n4540 ^ n221 ^ 1'b0 ;
  assign n4542 = n974 & n4541 ;
  assign n4538 = n2612 & n2650 ;
  assign n4539 = n1207 | n4538 ;
  assign n4543 = n4542 ^ n4539 ^ 1'b0 ;
  assign n4544 = n4543 ^ n2486 ^ 1'b0 ;
  assign n4549 = n829 & ~n2468 ;
  assign n4550 = ~n1237 & n4549 ;
  assign n4545 = n1944 ^ n1428 ^ n946 ;
  assign n4546 = n1767 | n4545 ;
  assign n4547 = n3314 & n4546 ;
  assign n4548 = n3484 | n4547 ;
  assign n4551 = n4550 ^ n4548 ^ 1'b0 ;
  assign n4552 = n357 | n4551 ;
  assign n4553 = n4552 ^ n600 ^ 1'b0 ;
  assign n4554 = n2204 ^ n150 ^ 1'b0 ;
  assign n4555 = ~n1276 & n2063 ;
  assign n4556 = n4555 ^ n1798 ^ 1'b0 ;
  assign n4557 = n1688 | n2139 ;
  assign n4558 = n2596 | n4557 ;
  assign n4559 = ~n477 & n4558 ;
  assign n4560 = n3325 | n4048 ;
  assign n4561 = ( n1282 & n2859 ) | ( n1282 & ~n3600 ) | ( n2859 & ~n3600 ) ;
  assign n4562 = n1914 & n4197 ;
  assign n4563 = n699 ^ n21 ^ 1'b0 ;
  assign n4564 = n3364 ^ n1659 ^ 1'b0 ;
  assign n4565 = n1513 ^ n52 ^ 1'b0 ;
  assign n4566 = n292 & ~n4565 ;
  assign n4567 = n1072 | n4566 ;
  assign n4568 = ~n1387 & n4567 ;
  assign n4569 = n2233 | n4568 ;
  assign n4570 = n3858 ^ n1170 ^ 1'b0 ;
  assign n4571 = n2022 & ~n4570 ;
  assign n4572 = ( n20 & n1066 ) | ( n20 & n1256 ) | ( n1066 & n1256 ) ;
  assign n4573 = n4572 ^ n2810 ^ n644 ;
  assign n4574 = ~n1398 & n4573 ;
  assign n4575 = n4574 ^ n3738 ^ 1'b0 ;
  assign n4576 = n968 | n1372 ;
  assign n4577 = n4575 & n4576 ;
  assign n4578 = n4571 & n4577 ;
  assign n4579 = n821 ^ n184 ^ 1'b0 ;
  assign n4580 = n4579 ^ n296 ^ 1'b0 ;
  assign n4581 = n226 | n4580 ;
  assign n4582 = n1231 | n4581 ;
  assign n4583 = n441 | n4582 ;
  assign n4584 = n3736 | n4583 ;
  assign n4585 = n982 & ~n4584 ;
  assign n4586 = n1504 & n1573 ;
  assign n4587 = n212 & ~n1050 ;
  assign n4588 = n1767 ^ n1215 ^ 1'b0 ;
  assign n4589 = n3690 ^ n315 ^ 1'b0 ;
  assign n4590 = n884 & n4589 ;
  assign n4591 = n3724 & n4590 ;
  assign n4592 = n404 & n4591 ;
  assign n4593 = ~n4588 & n4592 ;
  assign n4594 = n490 ^ n489 ^ 1'b0 ;
  assign n4595 = n894 | n4594 ;
  assign n4596 = n2332 & ~n4595 ;
  assign n4597 = n4596 ^ n3009 ^ 1'b0 ;
  assign n4599 = n1301 & n2393 ;
  assign n4600 = n822 | n1685 ;
  assign n4601 = n4600 ^ n3746 ^ 1'b0 ;
  assign n4602 = ~n2929 & n4601 ;
  assign n4603 = n216 & n4602 ;
  assign n4604 = ~n4599 & n4603 ;
  assign n4598 = n806 & ~n1343 ;
  assign n4605 = n4604 ^ n4598 ^ 1'b0 ;
  assign n4606 = n564 | n654 ;
  assign n4607 = n162 & ~n4606 ;
  assign n4608 = n533 & ~n4607 ;
  assign n4609 = n1912 ^ n1700 ^ 1'b0 ;
  assign n4610 = n839 & n4609 ;
  assign n4611 = ~n3725 & n4610 ;
  assign n4612 = n883 & n4611 ;
  assign n4613 = n1796 ^ n271 ^ 1'b0 ;
  assign n4614 = n4613 ^ n766 ^ 1'b0 ;
  assign n4615 = n2640 | n4614 ;
  assign n4616 = n4615 ^ n3564 ^ 1'b0 ;
  assign n4617 = n4612 | n4616 ;
  assign n4618 = n4617 ^ n379 ^ 1'b0 ;
  assign n4619 = n4618 ^ n2308 ^ 1'b0 ;
  assign n4620 = n1395 | n3867 ;
  assign n4621 = n79 | n4620 ;
  assign n4622 = n495 | n1853 ;
  assign n4623 = n4622 ^ n1307 ^ 1'b0 ;
  assign n4624 = n298 & n4623 ;
  assign n4625 = n3685 ^ n1477 ^ 1'b0 ;
  assign n4626 = n1196 | n4625 ;
  assign n4627 = n617 | n4626 ;
  assign n4628 = n4624 & ~n4627 ;
  assign n4629 = ~n4621 & n4628 ;
  assign n4630 = n3833 ^ n2694 ^ 1'b0 ;
  assign n4631 = n1157 & ~n4630 ;
  assign n4632 = n3761 ^ n2481 ^ 1'b0 ;
  assign n4633 = n3306 & n4632 ;
  assign n4634 = n2217 & n4633 ;
  assign n4635 = n2045 & ~n2501 ;
  assign n4636 = n183 & ~n1966 ;
  assign n4637 = n1664 | n3239 ;
  assign n4638 = ~n1794 & n4637 ;
  assign n4639 = n4638 ^ n265 ^ 1'b0 ;
  assign n4640 = n1118 & ~n1448 ;
  assign n4641 = n4640 ^ n2303 ^ 1'b0 ;
  assign n4642 = n3232 & ~n4641 ;
  assign n4643 = ~n286 & n4642 ;
  assign n4644 = n1829 & n4528 ;
  assign n4645 = n1794 ^ n315 ^ 1'b0 ;
  assign n4646 = n4645 ^ n1079 ^ 1'b0 ;
  assign n4647 = n1083 ^ n846 ^ 1'b0 ;
  assign n4648 = n2747 | n4647 ;
  assign n4649 = ~n48 & n229 ;
  assign n4650 = n3951 & n4649 ;
  assign n4651 = n3166 ^ n1653 ^ 1'b0 ;
  assign n4652 = n4177 & n4651 ;
  assign n4653 = n4652 ^ n4037 ^ 1'b0 ;
  assign n4661 = n683 | n1014 ;
  assign n4662 = n4661 ^ n3584 ^ 1'b0 ;
  assign n4654 = n443 & n492 ;
  assign n4655 = n295 & n4654 ;
  assign n4656 = ~n1948 & n1991 ;
  assign n4657 = n4656 ^ n606 ^ 1'b0 ;
  assign n4658 = n2420 & ~n3449 ;
  assign n4659 = ~n4657 & n4658 ;
  assign n4660 = ~n4655 & n4659 ;
  assign n4663 = n4662 ^ n4660 ^ 1'b0 ;
  assign n4664 = n717 | n4663 ;
  assign n4665 = n539 & ~n2803 ;
  assign n4666 = n412 & n4665 ;
  assign n4667 = n2890 ^ n1995 ^ n795 ;
  assign n4670 = n395 & n479 ;
  assign n4668 = ( n2881 & n3231 ) | ( n2881 & n4200 ) | ( n3231 & n4200 ) ;
  assign n4669 = n219 | n4668 ;
  assign n4671 = n4670 ^ n4669 ^ 1'b0 ;
  assign n4672 = n4671 ^ n547 ^ 1'b0 ;
  assign n4675 = n1148 ^ n1077 ^ 1'b0 ;
  assign n4673 = n774 & n798 ;
  assign n4674 = n4673 ^ n620 ^ 1'b0 ;
  assign n4676 = n4675 ^ n4674 ^ n1276 ;
  assign n4677 = ~n315 & n2962 ;
  assign n4678 = n4677 ^ n767 ^ 1'b0 ;
  assign n4679 = n1077 | n4678 ;
  assign n4680 = n1291 | n1386 ;
  assign n4681 = n659 & ~n4680 ;
  assign n4682 = n873 & n1301 ;
  assign n4683 = n4682 ^ n2973 ^ 1'b0 ;
  assign n4684 = ~n110 & n903 ;
  assign n4685 = n4684 ^ n844 ^ 1'b0 ;
  assign n4686 = n4685 ^ n1753 ^ 1'b0 ;
  assign n4687 = n4683 & ~n4686 ;
  assign n4688 = n582 | n4687 ;
  assign n4689 = n96 & ~n4688 ;
  assign n4690 = n4689 ^ n3687 ^ 1'b0 ;
  assign n4691 = n541 | n4690 ;
  assign n4692 = n708 & ~n3746 ;
  assign n4693 = ~n2675 & n4692 ;
  assign n4694 = n940 | n1024 ;
  assign n4695 = n3789 ^ n766 ^ 1'b0 ;
  assign n4696 = n4694 | n4695 ;
  assign n4697 = n4693 | n4696 ;
  assign n4698 = n4697 ^ n3190 ^ 1'b0 ;
  assign n4699 = n2749 ^ n1670 ^ 1'b0 ;
  assign n4700 = ~n3918 & n4699 ;
  assign n4701 = n868 ^ n508 ^ 1'b0 ;
  assign n4702 = n283 ^ n277 ^ 1'b0 ;
  assign n4703 = n4702 ^ n3766 ^ 1'b0 ;
  assign n4704 = n4701 & n4703 ;
  assign n4707 = n625 & ~n4573 ;
  assign n4708 = ~n1072 & n4707 ;
  assign n4709 = n4708 ^ n1441 ^ 1'b0 ;
  assign n4710 = ( ~n539 & n3124 ) | ( ~n539 & n4709 ) | ( n3124 & n4709 ) ;
  assign n4705 = n959 ^ n287 ^ 1'b0 ;
  assign n4706 = ~n4380 & n4705 ;
  assign n4711 = n4710 ^ n4706 ^ 1'b0 ;
  assign n4712 = n2927 & ~n3742 ;
  assign n4713 = n1989 & ~n4712 ;
  assign n4714 = n4713 ^ n3693 ^ 1'b0 ;
  assign n4715 = ~n1095 & n2246 ;
  assign n4716 = n1845 & n4715 ;
  assign n4717 = n4714 & ~n4716 ;
  assign n4718 = ~n3307 & n4717 ;
  assign n4719 = n4718 ^ n2964 ^ n2377 ;
  assign n4720 = n3576 & ~n4719 ;
  assign n4721 = ~n1280 & n1545 ;
  assign n4722 = n4721 ^ n1623 ^ 1'b0 ;
  assign n4723 = n2077 & n3469 ;
  assign n4724 = n4723 ^ n1335 ^ 1'b0 ;
  assign n4731 = n545 & n1221 ;
  assign n4730 = ~n183 & n358 ;
  assign n4732 = n4731 ^ n4730 ^ 1'b0 ;
  assign n4725 = n1352 | n2708 ;
  assign n4726 = n211 | n2449 ;
  assign n4727 = n4726 ^ n1124 ^ 1'b0 ;
  assign n4728 = n4727 ^ n1096 ^ 1'b0 ;
  assign n4729 = n4725 & n4728 ;
  assign n4733 = n4732 ^ n4729 ^ n4705 ;
  assign n4734 = n1884 | n3145 ;
  assign n4735 = n218 & n2439 ;
  assign n4736 = n2072 & n4735 ;
  assign n4737 = n4736 ^ n1420 ^ 1'b0 ;
  assign n4738 = n4737 ^ n2524 ^ 1'b0 ;
  assign n4740 = ~n169 & n283 ;
  assign n4739 = n1105 & ~n3975 ;
  assign n4741 = n4740 ^ n4739 ^ 1'b0 ;
  assign n4742 = ~n40 & n3303 ;
  assign n4743 = n4742 ^ n1085 ^ 1'b0 ;
  assign n4744 = n3220 & ~n4743 ;
  assign n4745 = n4135 ^ n2294 ^ 1'b0 ;
  assign n4746 = n791 | n2472 ;
  assign n4747 = n4675 ^ n2605 ^ n2461 ;
  assign n4748 = ~n4746 & n4747 ;
  assign n4749 = n249 & n4748 ;
  assign n4750 = ~n2564 & n4749 ;
  assign n4751 = n3105 ^ n253 ^ 1'b0 ;
  assign n4752 = n3923 ^ n2876 ^ 1'b0 ;
  assign n4753 = n4751 & ~n4752 ;
  assign n4759 = ~n3565 & n3691 ;
  assign n4760 = n4759 ^ n3049 ^ 1'b0 ;
  assign n4754 = n481 | n1012 ;
  assign n4755 = ~n3552 & n4754 ;
  assign n4756 = n3699 ^ n372 ^ 1'b0 ;
  assign n4757 = ~n916 & n4756 ;
  assign n4758 = n4755 & n4757 ;
  assign n4761 = n4760 ^ n4758 ^ 1'b0 ;
  assign n4762 = n1631 & ~n3858 ;
  assign n4763 = ~n1419 & n1513 ;
  assign n4764 = ~n3487 & n4763 ;
  assign n4765 = n431 | n2406 ;
  assign n4766 = n2739 | n4765 ;
  assign n4767 = n4764 & ~n4766 ;
  assign n4768 = ~n4762 & n4767 ;
  assign n4769 = n1234 & ~n3366 ;
  assign n4770 = n4769 ^ n2993 ^ 1'b0 ;
  assign n4771 = n4770 ^ n3996 ^ 1'b0 ;
  assign n4772 = n3406 | n4771 ;
  assign n4773 = n4768 | n4772 ;
  assign n4774 = n4773 ^ n3757 ^ 1'b0 ;
  assign n4775 = n2347 ^ n448 ^ n277 ;
  assign n4776 = n3909 ^ n3837 ^ n49 ;
  assign n4777 = n2082 & ~n4776 ;
  assign n4778 = n4777 ^ n4010 ^ 1'b0 ;
  assign n4779 = n1720 ^ n1300 ^ 1'b0 ;
  assign n4780 = n1826 & ~n4779 ;
  assign n4781 = n2883 & ~n4780 ;
  assign n4782 = n600 & ~n4781 ;
  assign n4783 = n551 & ~n4782 ;
  assign n4784 = n4783 ^ n2063 ^ 1'b0 ;
  assign n4785 = n3744 ^ n1589 ^ 1'b0 ;
  assign n4786 = n1865 | n4785 ;
  assign n4787 = n1589 | n4786 ;
  assign n4788 = ~n2650 & n2764 ;
  assign n4789 = n136 & n4788 ;
  assign n4790 = n4789 ^ n1479 ^ 1'b0 ;
  assign n4794 = n1251 | n1361 ;
  assign n4795 = ~n3008 & n4794 ;
  assign n4791 = n374 | n2728 ;
  assign n4792 = n2083 & ~n4791 ;
  assign n4793 = n915 & ~n4792 ;
  assign n4796 = n4795 ^ n4793 ^ 1'b0 ;
  assign n4797 = n3473 ^ n27 ^ 1'b0 ;
  assign n4798 = n996 ^ n212 ^ 1'b0 ;
  assign n4799 = n2266 & n4798 ;
  assign n4800 = n4799 ^ n1069 ^ 1'b0 ;
  assign n4801 = n4609 ^ n1853 ^ 1'b0 ;
  assign n4802 = n4801 ^ n2649 ^ 1'b0 ;
  assign n4803 = n2398 & ~n3324 ;
  assign n4804 = n3080 & n4803 ;
  assign n4805 = n4422 ^ n2275 ^ 1'b0 ;
  assign n4806 = ~n2767 & n2816 ;
  assign n4807 = ~n4805 & n4806 ;
  assign n4808 = n3545 | n4807 ;
  assign n4809 = x1 & n1073 ;
  assign n4810 = n4809 ^ n2681 ^ 1'b0 ;
  assign n4811 = n2395 ^ n1308 ^ 1'b0 ;
  assign n4812 = n578 & ~n4811 ;
  assign n4813 = ( n3774 & n4810 ) | ( n3774 & ~n4812 ) | ( n4810 & ~n4812 ) ;
  assign n4814 = n4233 & n4423 ;
  assign n4815 = ~n104 & n4007 ;
  assign n4816 = n275 & n4815 ;
  assign n4817 = n4816 ^ n1507 ^ 1'b0 ;
  assign n4821 = ~n663 & n1625 ;
  assign n4822 = ~n367 & n4821 ;
  assign n4818 = n667 & ~n2483 ;
  assign n4819 = n4818 ^ n160 ^ 1'b0 ;
  assign n4820 = n2438 & ~n4819 ;
  assign n4823 = n4822 ^ n4820 ^ 1'b0 ;
  assign n4824 = ~n4194 & n4823 ;
  assign n4825 = ~n2244 & n4596 ;
  assign n4826 = n4825 ^ n430 ^ 1'b0 ;
  assign n4827 = n4826 ^ n1443 ^ 1'b0 ;
  assign n4828 = n2377 | n2397 ;
  assign n4829 = n1740 | n4828 ;
  assign n4830 = ~n1918 & n4829 ;
  assign n4831 = n4830 ^ n2607 ^ 1'b0 ;
  assign n4832 = n2045 & n4831 ;
  assign n4833 = n2930 | n3261 ;
  assign n4834 = ( n125 & n2067 ) | ( n125 & ~n4833 ) | ( n2067 & ~n4833 ) ;
  assign n4835 = n2081 ^ n848 ^ 1'b0 ;
  assign n4836 = n1391 | n2664 ;
  assign n4837 = n4835 | n4836 ;
  assign n4838 = n2881 | n4837 ;
  assign n4839 = ~n4834 & n4838 ;
  assign n4840 = n4718 & n4839 ;
  assign n4841 = ( n1816 & n4542 ) | ( n1816 & n4840 ) | ( n4542 & n4840 ) ;
  assign n4842 = n340 & n1165 ;
  assign n4843 = n4842 ^ n2435 ^ 1'b0 ;
  assign n4844 = n4064 ^ n1361 ^ 1'b0 ;
  assign n4845 = n387 & n4844 ;
  assign n4846 = ( n1211 & n2155 ) | ( n1211 & n4845 ) | ( n2155 & n4845 ) ;
  assign n4847 = ~n56 & n1712 ;
  assign n4848 = n4846 & n4847 ;
  assign n4854 = n800 ^ n465 ^ 1'b0 ;
  assign n4855 = n334 & n4854 ;
  assign n4856 = n2583 | n4855 ;
  assign n4849 = ~n1212 & n1312 ;
  assign n4850 = n277 | n2102 ;
  assign n4851 = n2824 | n4850 ;
  assign n4852 = n1448 & ~n4851 ;
  assign n4853 = n4849 & n4852 ;
  assign n4857 = n4856 ^ n4853 ^ 1'b0 ;
  assign n4858 = n2332 | n4448 ;
  assign n4859 = n1709 ^ n445 ^ 1'b0 ;
  assign n4860 = n4859 ^ n846 ^ 1'b0 ;
  assign n4861 = ~n392 & n402 ;
  assign n4862 = n3284 & n4861 ;
  assign n4863 = n3153 & ~n4147 ;
  assign n4864 = n1767 & ~n4472 ;
  assign n4865 = n2631 & ~n4864 ;
  assign n4866 = n2408 ^ n1705 ^ 1'b0 ;
  assign n4867 = n1208 | n1437 ;
  assign n4868 = n1823 | n4867 ;
  assign n4869 = n4203 & n4868 ;
  assign n4870 = n588 & n4869 ;
  assign n4871 = n1469 & ~n2267 ;
  assign n4872 = n4871 ^ n3977 ^ 1'b0 ;
  assign n4873 = n4701 & n4872 ;
  assign n4874 = n637 & n3206 ;
  assign n4875 = n4874 ^ n2062 ^ 1'b0 ;
  assign n4876 = n3757 & n4875 ;
  assign n4877 = n4876 ^ n1398 ^ 1'b0 ;
  assign n4878 = n1476 & ~n3297 ;
  assign n4879 = n792 & n4878 ;
  assign n4880 = n52 & ~n4879 ;
  assign n4881 = ~n3198 & n4880 ;
  assign n4882 = n4485 | n4881 ;
  assign n4883 = n857 & ~n4882 ;
  assign n4884 = n2397 & n4457 ;
  assign n4885 = n4483 ^ n3363 ^ 1'b0 ;
  assign n4886 = ( n590 & n991 ) | ( n590 & ~n4885 ) | ( n991 & ~n4885 ) ;
  assign n4887 = n1729 ^ n535 ^ 1'b0 ;
  assign n4888 = ~n607 & n4887 ;
  assign n4889 = n65 | n1794 ;
  assign n4890 = n1601 | n4889 ;
  assign n4891 = n4835 | n4890 ;
  assign n4892 = n1857 & n4891 ;
  assign n4893 = n4892 ^ n2915 ^ 1'b0 ;
  assign n4894 = ( n302 & n561 ) | ( n302 & ~n1147 ) | ( n561 & ~n1147 ) ;
  assign n4895 = x0 & n4894 ;
  assign n4896 = n4895 ^ n124 ^ 1'b0 ;
  assign n4897 = n802 | n4896 ;
  assign n4898 = n3471 & ~n4897 ;
  assign n4899 = n4898 ^ n4407 ^ 1'b0 ;
  assign n4900 = ~n177 & n796 ;
  assign n4901 = n374 & n4900 ;
  assign n4902 = n4901 ^ n2799 ^ 1'b0 ;
  assign n4903 = n220 & n3798 ;
  assign n4904 = n2914 & n4173 ;
  assign n4905 = n695 & n4904 ;
  assign n4906 = n4280 ^ n1009 ^ 1'b0 ;
  assign n4907 = n924 & ~n4906 ;
  assign n4908 = n3160 ^ n910 ^ 1'b0 ;
  assign n4909 = n4907 & n4908 ;
  assign n4912 = n285 | n717 ;
  assign n4913 = ~n541 & n4912 ;
  assign n4914 = n1383 & n4683 ;
  assign n4915 = ~n1803 & n4914 ;
  assign n4916 = ~n4913 & n4915 ;
  assign n4910 = n4754 ^ n269 ^ 1'b0 ;
  assign n4911 = n541 & ~n4910 ;
  assign n4917 = n4916 ^ n4911 ^ 1'b0 ;
  assign n4918 = ( n1379 & n1775 ) | ( n1379 & n2577 ) | ( n1775 & n2577 ) ;
  assign n4919 = n2225 & n4918 ;
  assign n4920 = n1943 ^ n528 ^ 1'b0 ;
  assign n4921 = ( n422 & ~n737 ) | ( n422 & n4920 ) | ( ~n737 & n4920 ) ;
  assign n4926 = ~n260 & n543 ;
  assign n4924 = ~n1534 & n3473 ;
  assign n4922 = ( ~n2813 & n3146 ) | ( ~n2813 & n3392 ) | ( n3146 & n3392 ) ;
  assign n4923 = n4157 & ~n4922 ;
  assign n4925 = n4924 ^ n4923 ^ 1'b0 ;
  assign n4927 = n4926 ^ n4925 ^ 1'b0 ;
  assign n4928 = n466 & ~n4927 ;
  assign n4929 = n2273 ^ n535 ^ 1'b0 ;
  assign n4930 = n957 & ~n4929 ;
  assign n4931 = n4930 ^ n439 ^ 1'b0 ;
  assign n4933 = n1988 ^ n1369 ^ 1'b0 ;
  assign n4932 = n1283 ^ n1154 ^ 1'b0 ;
  assign n4934 = n4933 ^ n4932 ^ 1'b0 ;
  assign n4935 = n4931 | n4934 ;
  assign n4937 = n1693 ^ n659 ^ 1'b0 ;
  assign n4936 = n437 & ~n3792 ;
  assign n4938 = n4937 ^ n4936 ^ 1'b0 ;
  assign n4939 = n417 & ~n3399 ;
  assign n4940 = n4939 ^ n2314 ^ n2061 ;
  assign n4941 = ~n466 & n4634 ;
  assign n4942 = n487 & ~n4007 ;
  assign n4946 = ~n192 & n4698 ;
  assign n4943 = n640 | n2179 ;
  assign n4944 = n4943 ^ n1960 ^ 1'b0 ;
  assign n4945 = n4944 ^ n1231 ^ 1'b0 ;
  assign n4947 = n4946 ^ n4945 ^ 1'b0 ;
  assign n4948 = n514 ^ n271 ^ 1'b0 ;
  assign n4949 = n3085 ^ n1352 ^ 1'b0 ;
  assign n4952 = n421 & n2428 ;
  assign n4950 = n3126 ^ n1744 ^ 1'b0 ;
  assign n4951 = n1118 & ~n4950 ;
  assign n4953 = n4952 ^ n4951 ^ 1'b0 ;
  assign n4954 = n4949 & n4953 ;
  assign n4955 = n4954 ^ n243 ^ 1'b0 ;
  assign n4964 = ~n1763 & n3367 ;
  assign n4965 = n4964 ^ n1989 ^ 1'b0 ;
  assign n4966 = n4965 ^ n2252 ^ 1'b0 ;
  assign n4967 = n2257 & n4966 ;
  assign n4968 = ~n1534 & n4967 ;
  assign n4956 = n150 | n1907 ;
  assign n4957 = n929 & ~n3409 ;
  assign n4958 = n4957 ^ n3513 ^ 1'b0 ;
  assign n4959 = n205 & n2065 ;
  assign n4960 = n4959 ^ n1136 ^ 1'b0 ;
  assign n4961 = ~n593 & n4960 ;
  assign n4962 = ~n4958 & n4961 ;
  assign n4963 = n4956 & ~n4962 ;
  assign n4969 = n4968 ^ n4963 ^ 1'b0 ;
  assign n4970 = n4403 ^ n1177 ^ 1'b0 ;
  assign n4971 = n4409 ^ n2593 ^ 1'b0 ;
  assign n4972 = n3179 & ~n4167 ;
  assign n4973 = n4972 ^ n3582 ^ 1'b0 ;
  assign n4974 = n1078 & n3667 ;
  assign n4975 = n4974 ^ n1488 ^ 1'b0 ;
  assign n4976 = ~n1289 & n3469 ;
  assign n4977 = n2671 ^ n214 ^ 1'b0 ;
  assign n4978 = n2826 ^ n2214 ^ 1'b0 ;
  assign n4979 = ~n2139 & n4978 ;
  assign n4980 = n3783 & ~n4451 ;
  assign n4981 = ( n1983 & ~n3924 ) | ( n1983 & n4195 ) | ( ~n3924 & n4195 ) ;
  assign n4982 = x6 & n2883 ;
  assign n4984 = n1761 ^ n562 ^ 1'b0 ;
  assign n4985 = n727 | n1598 ;
  assign n4986 = n4984 | n4985 ;
  assign n4987 = ~n1454 & n4986 ;
  assign n4988 = n4987 ^ n3248 ^ 1'b0 ;
  assign n4983 = ( n1654 & n2435 ) | ( n1654 & n3797 ) | ( n2435 & n3797 ) ;
  assign n4989 = n4988 ^ n4983 ^ 1'b0 ;
  assign n4990 = ~n224 & n1460 ;
  assign n4991 = n4990 ^ n1907 ^ 1'b0 ;
  assign n4992 = n3818 ^ n328 ^ 1'b0 ;
  assign n4993 = n4054 & n4992 ;
  assign n4994 = n2505 & n4993 ;
  assign n4995 = n4994 ^ n2626 ^ 1'b0 ;
  assign n4996 = ~n175 & n1312 ;
  assign n4997 = n4996 ^ n1811 ^ 1'b0 ;
  assign n4998 = n4997 ^ n4381 ^ 1'b0 ;
  assign n4999 = n3845 | n4998 ;
  assign n5000 = n2935 ^ n229 ^ 1'b0 ;
  assign n5001 = ~n2205 & n5000 ;
  assign n5002 = n920 & ~n5001 ;
  assign n5003 = ~n4999 & n5002 ;
  assign n5004 = n4675 ^ n959 ^ 1'b0 ;
  assign n5005 = n5004 ^ n1688 ^ 1'b0 ;
  assign n5006 = n725 & ~n2781 ;
  assign n5007 = n5006 ^ n3058 ^ 1'b0 ;
  assign n5008 = n2236 | n5007 ;
  assign n5009 = n3577 & ~n5008 ;
  assign n5010 = n5009 ^ n640 ^ 1'b0 ;
  assign n5011 = n5010 ^ n1326 ^ 1'b0 ;
  assign n5012 = ~n2310 & n5011 ;
  assign n5013 = n119 | n451 ;
  assign n5014 = n205 | n5013 ;
  assign n5015 = n5014 ^ n2764 ^ n1546 ;
  assign n5016 = n1927 & ~n2004 ;
  assign n5017 = n709 | n5016 ;
  assign n5018 = n1505 | n5017 ;
  assign n5019 = n1104 & ~n3867 ;
  assign n5020 = n188 & n5019 ;
  assign n5021 = n5020 ^ n2033 ^ 1'b0 ;
  assign n5022 = n5021 ^ n940 ^ 1'b0 ;
  assign n5023 = n2480 ^ n404 ^ 1'b0 ;
  assign n5024 = n3284 ^ n305 ^ 1'b0 ;
  assign n5025 = n2114 & n5024 ;
  assign n5026 = n2895 ^ n431 ^ 1'b0 ;
  assign n5027 = n5026 ^ n3787 ^ n2504 ;
  assign n5028 = n1207 ^ n1066 ^ 1'b0 ;
  assign n5029 = ~n910 & n3989 ;
  assign n5030 = n5029 ^ n3150 ^ 1'b0 ;
  assign n5032 = ( n487 & ~n813 ) | ( n487 & n1620 ) | ( ~n813 & n1620 ) ;
  assign n5031 = n2811 ^ n819 ^ n263 ;
  assign n5033 = n5032 ^ n5031 ^ n221 ;
  assign n5034 = n2492 | n5033 ;
  assign n5035 = n5034 ^ n422 ^ 1'b0 ;
  assign n5036 = n5030 | n5035 ;
  assign n5037 = n1546 | n3162 ;
  assign n5038 = n2114 & ~n2527 ;
  assign n5039 = n5038 ^ n2508 ^ 1'b0 ;
  assign n5040 = n5037 & ~n5039 ;
  assign n5041 = n1901 ^ n798 ^ 1'b0 ;
  assign n5042 = n4757 | n5041 ;
  assign n5043 = n1633 & n3751 ;
  assign n5044 = n2893 & n5043 ;
  assign n5045 = n5044 ^ n3382 ^ 1'b0 ;
  assign n5046 = ( n905 & ~n2761 ) | ( n905 & n4850 ) | ( ~n2761 & n4850 ) ;
  assign n5047 = n2388 | n5046 ;
  assign n5048 = ( n3861 & n4267 ) | ( n3861 & n5047 ) | ( n4267 & n5047 ) ;
  assign n5049 = n2569 & ~n4709 ;
  assign n5050 = n5049 ^ n4960 ^ 1'b0 ;
  assign n5051 = n774 & n5050 ;
  assign n5052 = n924 & n5051 ;
  assign n5053 = n1480 ^ n108 ^ 1'b0 ;
  assign n5054 = n1589 & n5053 ;
  assign n5055 = n3474 | n5054 ;
  assign n5056 = ~n3641 & n4671 ;
  assign n5057 = ~n565 & n5056 ;
  assign n5058 = n1528 ^ n543 ^ 1'b0 ;
  assign n5059 = ~n213 & n1660 ;
  assign n5063 = n698 & ~n1728 ;
  assign n5060 = n757 | n3009 ;
  assign n5061 = n5060 ^ n1659 ^ 1'b0 ;
  assign n5062 = ~n322 & n5061 ;
  assign n5064 = n5063 ^ n5062 ^ 1'b0 ;
  assign n5065 = n2600 ^ n489 ^ 1'b0 ;
  assign n5069 = ~n1164 & n3411 ;
  assign n5066 = n2894 ^ n2367 ^ 1'b0 ;
  assign n5067 = n1007 & n5066 ;
  assign n5068 = ~n368 & n5067 ;
  assign n5070 = n5069 ^ n5068 ^ 1'b0 ;
  assign n5071 = n395 & ~n3036 ;
  assign n5072 = n4080 & n5071 ;
  assign n5073 = n668 | n2835 ;
  assign n5074 = n1516 & ~n2250 ;
  assign n5075 = n5074 ^ n93 ^ 1'b0 ;
  assign n5076 = ~n5073 & n5075 ;
  assign n5077 = n5076 ^ n1816 ^ 1'b0 ;
  assign n5078 = n1811 ^ n1558 ^ 1'b0 ;
  assign n5079 = n4085 ^ n1654 ^ n1594 ;
  assign n5080 = n2998 ^ n2030 ^ 1'b0 ;
  assign n5081 = n1382 & n5080 ;
  assign n5082 = n2404 ^ n431 ^ 1'b0 ;
  assign n5083 = n2820 | n5082 ;
  assign n5084 = ( n721 & n3357 ) | ( n721 & ~n5083 ) | ( n3357 & ~n5083 ) ;
  assign n5085 = ( n423 & n1298 ) | ( n423 & ~n1338 ) | ( n1298 & ~n1338 ) ;
  assign n5086 = n5084 & ~n5085 ;
  assign n5087 = n5086 ^ n2756 ^ 1'b0 ;
  assign n5088 = n619 & ~n5087 ;
  assign n5089 = n2554 | n3464 ;
  assign n5090 = n5089 ^ n3778 ^ 1'b0 ;
  assign n5091 = n5088 & n5090 ;
  assign n5092 = n738 & n2455 ;
  assign n5093 = n227 & n5092 ;
  assign n5094 = n1385 | n4848 ;
  assign n5095 = n5094 ^ n3974 ^ 1'b0 ;
  assign n5097 = n401 & n510 ;
  assign n5098 = n5097 ^ n2703 ^ 1'b0 ;
  assign n5099 = ~n1081 & n5098 ;
  assign n5096 = ~n652 & n2101 ;
  assign n5100 = n5099 ^ n5096 ^ n3989 ;
  assign n5101 = n676 | n5100 ;
  assign n5102 = n1098 & n2201 ;
  assign n5103 = n5102 ^ n1192 ^ 1'b0 ;
  assign n5104 = ( n1530 & n1752 ) | ( n1530 & n3823 ) | ( n1752 & n3823 ) ;
  assign n5105 = n5104 ^ n438 ^ 1'b0 ;
  assign n5106 = n4079 & n5105 ;
  assign n5107 = n1545 ^ n1521 ^ 1'b0 ;
  assign n5108 = n5107 ^ n48 ^ 1'b0 ;
  assign n5109 = n2150 & ~n2267 ;
  assign n5110 = n567 & ~n1624 ;
  assign n5111 = n225 | n1664 ;
  assign n5112 = n5111 ^ n2848 ^ 1'b0 ;
  assign n5113 = n5110 | n5112 ;
  assign n5114 = n2380 ^ n212 ^ 1'b0 ;
  assign n5115 = n5114 ^ n2110 ^ 1'b0 ;
  assign n5116 = n5113 & ~n5115 ;
  assign n5117 = n150 & ~n5116 ;
  assign n5118 = n5109 & n5117 ;
  assign n5128 = n2440 | n3045 ;
  assign n5129 = n3802 & n5128 ;
  assign n5130 = n5129 ^ n2955 ^ 1'b0 ;
  assign n5119 = n1563 | n1655 ;
  assign n5120 = n5119 ^ n4141 ^ 1'b0 ;
  assign n5124 = ( ~n1141 & n1662 ) | ( ~n1141 & n2501 ) | ( n1662 & n2501 ) ;
  assign n5121 = n942 & n1981 ;
  assign n5122 = n5121 ^ n4600 ^ 1'b0 ;
  assign n5123 = n2801 & ~n5122 ;
  assign n5125 = n5124 ^ n5123 ^ 1'b0 ;
  assign n5126 = n3437 | n5125 ;
  assign n5127 = n5120 | n5126 ;
  assign n5131 = n5130 ^ n5127 ^ 1'b0 ;
  assign n5132 = ~n539 & n2335 ;
  assign n5134 = n3252 ^ n2185 ^ 1'b0 ;
  assign n5135 = n2547 | n5134 ;
  assign n5136 = n5135 ^ n3339 ^ 1'b0 ;
  assign n5133 = ~n263 & n4236 ;
  assign n5137 = n5136 ^ n5133 ^ 1'b0 ;
  assign n5138 = n5132 & ~n5137 ;
  assign n5139 = ~n294 & n347 ;
  assign n5140 = n492 ^ n414 ^ 1'b0 ;
  assign n5141 = n3450 & ~n5140 ;
  assign n5142 = n1275 & n4273 ;
  assign n5143 = n5142 ^ n4484 ^ 1'b0 ;
  assign n5144 = n67 & n2741 ;
  assign n5145 = n2580 ^ n1620 ^ n1300 ;
  assign n5146 = n5145 ^ n1845 ^ 1'b0 ;
  assign n5147 = n3490 & ~n5146 ;
  assign n5148 = n966 & n2314 ;
  assign n5149 = n2223 & n5148 ;
  assign n5150 = n45 | n286 ;
  assign n5151 = n5150 ^ n2040 ^ n831 ;
  assign n5152 = n5151 ^ n3772 ^ 1'b0 ;
  assign n5153 = n1705 & ~n5152 ;
  assign n5154 = n5149 & n5153 ;
  assign n5155 = n1657 ^ n1455 ^ 1'b0 ;
  assign n5156 = n4919 & n5155 ;
  assign n5157 = n5154 & n5156 ;
  assign n5158 = n1854 & n2273 ;
  assign n5159 = n5158 ^ n5078 ^ 1'b0 ;
  assign n5160 = n5097 | n5159 ;
  assign n5161 = n3536 ^ n255 ^ 1'b0 ;
  assign n5162 = n4645 ^ n2637 ^ 1'b0 ;
  assign n5163 = ~n1907 & n5162 ;
  assign n5164 = n398 & ~n1438 ;
  assign n5165 = n5164 ^ n1273 ^ 1'b0 ;
  assign n5166 = ~n2753 & n3594 ;
  assign n5167 = ~n2374 & n3748 ;
  assign n5168 = n861 & n1428 ;
  assign n5169 = n2428 & n5168 ;
  assign n5170 = n5169 ^ n1184 ^ 1'b0 ;
  assign n5171 = n4154 | n5170 ;
  assign n5172 = n5171 ^ n533 ^ 1'b0 ;
  assign n5173 = n1744 ^ n508 ^ 1'b0 ;
  assign n5174 = n1533 | n5173 ;
  assign n5175 = n5174 ^ n88 ^ 1'b0 ;
  assign n5176 = ( n21 & n167 ) | ( n21 & n615 ) | ( n167 & n615 ) ;
  assign n5177 = n5176 ^ n132 ^ 1'b0 ;
  assign n5178 = ~n528 & n5177 ;
  assign n5179 = n2173 ^ n1456 ^ 1'b0 ;
  assign n5180 = n5179 ^ n508 ^ 1'b0 ;
  assign n5181 = n3437 & n5180 ;
  assign n5182 = ~n2306 & n2495 ;
  assign n5183 = n4153 ^ n2113 ^ 1'b0 ;
  assign n5184 = ~n3035 & n5183 ;
  assign n5188 = n2403 ^ n1442 ^ 1'b0 ;
  assign n5189 = ~n3996 & n5188 ;
  assign n5190 = ~n1246 & n2202 ;
  assign n5191 = n5190 ^ n2628 ^ 1'b0 ;
  assign n5192 = n3306 & ~n5191 ;
  assign n5193 = n5192 ^ n2317 ^ 1'b0 ;
  assign n5194 = n5189 | n5193 ;
  assign n5185 = n4038 ^ n2683 ^ 1'b0 ;
  assign n5186 = n3804 & ~n4095 ;
  assign n5187 = ( ~n291 & n5185 ) | ( ~n291 & n5186 ) | ( n5185 & n5186 ) ;
  assign n5195 = n5194 ^ n5187 ^ 1'b0 ;
  assign n5196 = n2147 & n3535 ;
  assign n5197 = n5196 ^ n2796 ^ 1'b0 ;
  assign n5198 = ~n2103 & n5197 ;
  assign n5199 = n1875 & n5198 ;
  assign n5200 = ~n695 & n3826 ;
  assign n5201 = n1608 ^ n1562 ^ 1'b0 ;
  assign n5202 = n1988 ^ n165 ^ 1'b0 ;
  assign n5203 = n1308 & ~n5202 ;
  assign n5204 = n5203 ^ n3891 ^ 1'b0 ;
  assign n5205 = n5204 ^ n767 ^ 1'b0 ;
  assign n5206 = ~n4351 & n5205 ;
  assign n5207 = n2146 ^ n1410 ^ 1'b0 ;
  assign n5208 = ~n1865 & n5207 ;
  assign n5209 = ~n592 & n5208 ;
  assign n5211 = n2460 ^ n1566 ^ n306 ;
  assign n5210 = n1392 & ~n2460 ;
  assign n5212 = n5211 ^ n5210 ^ 1'b0 ;
  assign n5213 = n808 | n3939 ;
  assign n5214 = n5213 ^ n1615 ^ 1'b0 ;
  assign n5215 = n2904 ^ n1458 ^ 1'b0 ;
  assign n5216 = n5215 ^ n2956 ^ n2918 ;
  assign n5217 = n1233 ^ n105 ^ 1'b0 ;
  assign n5218 = n5217 ^ n1428 ^ 1'b0 ;
  assign n5219 = n4355 ^ n3444 ^ 1'b0 ;
  assign n5220 = n3442 & n5219 ;
  assign n5221 = n5220 ^ n1690 ^ 1'b0 ;
  assign n5222 = ( n863 & ~n3426 ) | ( n863 & n3835 ) | ( ~n3426 & n3835 ) ;
  assign n5223 = n4651 & n5222 ;
  assign n5224 = n5223 ^ n3867 ^ 1'b0 ;
  assign n5225 = n1379 ^ n465 ^ 1'b0 ;
  assign n5226 = n3188 | n5225 ;
  assign n5227 = n5226 ^ n2808 ^ n1685 ;
  assign n5228 = n2946 ^ n2588 ^ 1'b0 ;
  assign n5229 = n5228 ^ n4755 ^ n43 ;
  assign n5230 = n428 | n5229 ;
  assign n5231 = n5230 ^ n3517 ^ 1'b0 ;
  assign n5232 = ~n959 & n5231 ;
  assign n5233 = n2806 | n3646 ;
  assign n5234 = n5233 ^ n91 ^ 1'b0 ;
  assign n5235 = n3338 | n5234 ;
  assign n5239 = n2120 & n4596 ;
  assign n5240 = n5239 ^ n910 ^ 1'b0 ;
  assign n5241 = n5240 ^ n3587 ^ 1'b0 ;
  assign n5236 = n3125 ^ n1714 ^ n760 ;
  assign n5237 = n3928 | n5236 ;
  assign n5238 = n1079 & n5237 ;
  assign n5242 = n5241 ^ n5238 ^ 1'b0 ;
  assign n5243 = n910 ^ n179 ^ 1'b0 ;
  assign n5244 = n5242 & ~n5243 ;
  assign n5245 = n4322 ^ n867 ^ 1'b0 ;
  assign n5246 = n1803 ^ n687 ^ 1'b0 ;
  assign n5247 = n2046 & ~n5246 ;
  assign n5248 = n2170 | n5247 ;
  assign n5249 = n5248 ^ n2709 ^ 1'b0 ;
  assign n5250 = ~n1531 & n5249 ;
  assign n5251 = n86 & ~n148 ;
  assign n5252 = n2719 | n5073 ;
  assign n5253 = n5251 | n5252 ;
  assign n5254 = n133 & n5253 ;
  assign n5255 = n2097 ^ n1473 ^ 1'b0 ;
  assign n5256 = n555 & n5255 ;
  assign n5257 = n3531 ^ n1548 ^ 1'b0 ;
  assign n5258 = n3232 & n5057 ;
  assign n5259 = n2907 ^ n1811 ^ 1'b0 ;
  assign n5260 = n1477 & n2223 ;
  assign n5262 = ( n1141 & n3434 ) | ( n1141 & n3881 ) | ( n3434 & n3881 ) ;
  assign n5263 = ( n1847 & ~n2960 ) | ( n1847 & n5262 ) | ( ~n2960 & n5262 ) ;
  assign n5261 = n2783 & ~n2872 ;
  assign n5264 = n5263 ^ n5261 ^ 1'b0 ;
  assign n5265 = n699 | n772 ;
  assign n5266 = n5265 ^ n821 ^ 1'b0 ;
  assign n5267 = ( n104 & n1924 ) | ( n104 & n5266 ) | ( n1924 & n5266 ) ;
  assign n5268 = n5267 ^ n1306 ^ 1'b0 ;
  assign n5269 = n944 | n1271 ;
  assign n5270 = n1027 | n5269 ;
  assign n5272 = n785 & n885 ;
  assign n5273 = n5272 ^ n1299 ^ 1'b0 ;
  assign n5274 = n5273 ^ n4519 ^ 1'b0 ;
  assign n5275 = n5274 ^ n3867 ^ 1'b0 ;
  assign n5276 = n489 & n5275 ;
  assign n5271 = n4326 & ~n4698 ;
  assign n5277 = n5276 ^ n5271 ^ 1'b0 ;
  assign n5278 = n89 & n3490 ;
  assign n5279 = n3095 & n5278 ;
  assign n5280 = n291 | n4990 ;
  assign n5281 = n5280 ^ n1367 ^ 1'b0 ;
  assign n5282 = n310 & ~n5281 ;
  assign n5283 = n5282 ^ n3207 ^ 1'b0 ;
  assign n5284 = n423 | n5283 ;
  assign n5285 = n4025 ^ n2668 ^ 1'b0 ;
  assign n5286 = n2951 | n4341 ;
  assign n5287 = x8 & ~n1241 ;
  assign n5288 = n5287 ^ n1438 ^ 1'b0 ;
  assign n5289 = ( ~n1363 & n2049 ) | ( ~n1363 & n5288 ) | ( n2049 & n5288 ) ;
  assign n5290 = n5289 ^ n140 ^ 1'b0 ;
  assign n5291 = n3983 & ~n5065 ;
  assign n5292 = n5291 ^ n1984 ^ 1'b0 ;
  assign n5293 = n988 & ~n2458 ;
  assign n5294 = ( n83 & n2288 ) | ( n83 & n2758 ) | ( n2288 & n2758 ) ;
  assign n5295 = n5294 ^ n1988 ^ 1'b0 ;
  assign n5296 = ( n809 & ~n5293 ) | ( n809 & n5295 ) | ( ~n5293 & n5295 ) ;
  assign n5297 = n1922 ^ n290 ^ 1'b0 ;
  assign n5298 = n1999 ^ n1419 ^ 1'b0 ;
  assign n5299 = ~n508 & n3869 ;
  assign n5300 = ~n1601 & n5299 ;
  assign n5301 = n1551 & ~n2210 ;
  assign n5302 = ~n74 & n5301 ;
  assign n5303 = n1845 | n5302 ;
  assign n5304 = n5303 ^ n3378 ^ n1124 ;
  assign n5305 = n5304 ^ n1578 ^ 1'b0 ;
  assign n5306 = n5249 ^ n3430 ^ 1'b0 ;
  assign n5307 = n1769 & ~n3700 ;
  assign n5308 = n5306 & n5307 ;
  assign n5309 = n567 ^ n406 ^ 1'b0 ;
  assign n5310 = n5309 ^ n4140 ^ 1'b0 ;
  assign n5311 = n2787 ^ n43 ^ 1'b0 ;
  assign n5312 = n844 | n1432 ;
  assign n5313 = n2885 | n5312 ;
  assign n5314 = n4698 | n4853 ;
  assign n5315 = n253 & ~n2050 ;
  assign n5316 = n19 & n5315 ;
  assign n5317 = n478 & ~n4579 ;
  assign n5318 = n4132 | n5317 ;
  assign n5319 = n3802 | n5318 ;
  assign n5321 = n1118 & ~n2017 ;
  assign n5322 = n171 & ~n5321 ;
  assign n5323 = n5322 ^ n4539 ^ 1'b0 ;
  assign n5320 = ~n1631 & n2580 ;
  assign n5324 = n5323 ^ n5320 ^ 1'b0 ;
  assign n5325 = n56 & ~n2987 ;
  assign n5326 = n5325 ^ n1434 ^ 1'b0 ;
  assign n5327 = n56 & ~n5326 ;
  assign n5328 = n5327 ^ n770 ^ 1'b0 ;
  assign n5329 = n4285 & n5328 ;
  assign n5330 = ~n2614 & n4092 ;
  assign n5331 = n5330 ^ n1105 ^ 1'b0 ;
  assign n5332 = ( n1063 & n5329 ) | ( n1063 & n5331 ) | ( n5329 & n5331 ) ;
  assign n5333 = n707 & n1491 ;
  assign n5334 = n5247 ^ n1186 ^ 1'b0 ;
  assign n5335 = ~n5333 & n5334 ;
  assign n5336 = ~n4267 & n5335 ;
  assign n5337 = n1416 & ~n3160 ;
  assign n5338 = ~n412 & n5337 ;
  assign n5339 = n4738 & ~n5338 ;
  assign n5340 = n5336 & n5339 ;
  assign n5341 = n79 & ~n2806 ;
  assign n5342 = n234 & n5341 ;
  assign n5343 = n2351 & ~n5342 ;
  assign n5344 = n5343 ^ n1194 ^ 1'b0 ;
  assign n5345 = n1872 ^ n251 ^ 1'b0 ;
  assign n5346 = ~n5344 & n5345 ;
  assign n5347 = n740 | n2973 ;
  assign n5348 = n5347 ^ n2095 ^ 1'b0 ;
  assign n5349 = ~n21 & n5348 ;
  assign n5350 = n837 ^ n451 ^ 1'b0 ;
  assign n5357 = n1631 ^ n896 ^ 1'b0 ;
  assign n5351 = n1117 & ~n2388 ;
  assign n5352 = ~n2832 & n5351 ;
  assign n5353 = n974 | n5352 ;
  assign n5354 = n5353 ^ n2407 ^ 1'b0 ;
  assign n5355 = ( n311 & ~n776 ) | ( n311 & n5354 ) | ( ~n776 & n5354 ) ;
  assign n5356 = n3859 & ~n5355 ;
  assign n5358 = n5357 ^ n5356 ^ 1'b0 ;
  assign n5359 = ( n2787 & n3125 ) | ( n2787 & n5358 ) | ( n3125 & n5358 ) ;
  assign n5360 = n5350 & ~n5359 ;
  assign n5361 = ~n2401 & n5354 ;
  assign n5362 = ~n3418 & n5361 ;
  assign n5363 = n1760 ^ n1439 ^ n1400 ;
  assign n5364 = ( ~n47 & n2806 ) | ( ~n47 & n5363 ) | ( n2806 & n5363 ) ;
  assign n5365 = n5364 ^ n4030 ^ 1'b0 ;
  assign n5366 = n5365 ^ n1898 ^ 1'b0 ;
  assign n5367 = n439 & n2547 ;
  assign n5368 = n4252 ^ n2250 ^ 1'b0 ;
  assign n5369 = n4233 ^ n2532 ^ 1'b0 ;
  assign n5370 = n369 | n1471 ;
  assign n5371 = n1320 | n5370 ;
  assign n5372 = n1431 & n3325 ;
  assign n5373 = n5371 & ~n5372 ;
  assign n5374 = ~n5369 & n5373 ;
  assign n5375 = n2178 | n2219 ;
  assign n5376 = n4980 & n5375 ;
  assign n5377 = n5376 ^ n2900 ^ 1'b0 ;
  assign n5378 = n825 | n1326 ;
  assign n5379 = ( n600 & n2484 ) | ( n600 & ~n5378 ) | ( n2484 & ~n5378 ) ;
  assign n5380 = n598 & n5379 ;
  assign n5381 = n130 & ~n5380 ;
  assign n5382 = n2796 | n2799 ;
  assign n5383 = n1215 & ~n2137 ;
  assign n5384 = n5383 ^ n458 ^ 1'b0 ;
  assign n5385 = ~n4367 & n5384 ;
  assign n5386 = ~n934 & n2909 ;
  assign n5387 = ~n212 & n5386 ;
  assign n5388 = n3730 ^ n2451 ^ 1'b0 ;
  assign n5389 = ~n1349 & n1907 ;
  assign n5390 = n5388 & n5389 ;
  assign n5391 = ~n249 & n1321 ;
  assign n5392 = ~n1628 & n3909 ;
  assign n5393 = n3181 ^ n861 ^ 1'b0 ;
  assign n5394 = n5392 & ~n5393 ;
  assign n5399 = n1282 & ~n1887 ;
  assign n5400 = n5399 ^ n3179 ^ 1'b0 ;
  assign n5395 = n170 | n541 ;
  assign n5396 = n3887 | n5395 ;
  assign n5397 = n5396 ^ n3080 ^ n2068 ;
  assign n5398 = n1466 | n5397 ;
  assign n5401 = n5400 ^ n5398 ^ 1'b0 ;
  assign n5402 = ~n362 & n532 ;
  assign n5403 = ( n717 & ~n1896 ) | ( n717 & n2492 ) | ( ~n1896 & n2492 ) ;
  assign n5404 = n5403 ^ n2927 ^ 1'b0 ;
  assign n5405 = n2319 & ~n3687 ;
  assign n5406 = n1607 ^ n1217 ^ 1'b0 ;
  assign n5407 = ~n1471 & n3108 ;
  assign n5408 = n5407 ^ n225 ^ 1'b0 ;
  assign n5409 = n5406 | n5408 ;
  assign n5410 = n5405 | n5409 ;
  assign n5411 = ( n1057 & n1109 ) | ( n1057 & n5410 ) | ( n1109 & n5410 ) ;
  assign n5412 = n4013 ^ n959 ^ 1'b0 ;
  assign n5413 = ~n1246 & n5412 ;
  assign n5414 = n3990 ^ n1558 ^ 1'b0 ;
  assign n5417 = ( n1300 & ~n2086 ) | ( n1300 & n2675 ) | ( ~n2086 & n2675 ) ;
  assign n5415 = n2891 | n4394 ;
  assign n5416 = n4615 & ~n5415 ;
  assign n5418 = n5417 ^ n5416 ^ 1'b0 ;
  assign n5419 = n5204 & ~n5418 ;
  assign n5420 = n3964 ^ n73 ^ 1'b0 ;
  assign n5421 = n1689 ^ n15 ^ 1'b0 ;
  assign n5422 = n219 | n5421 ;
  assign n5423 = n5422 ^ n4624 ^ 1'b0 ;
  assign n5424 = n2229 & ~n5423 ;
  assign n5425 = n5420 & n5424 ;
  assign n5426 = ~n2139 & n3417 ;
  assign n5432 = n3946 ^ n1734 ^ 1'b0 ;
  assign n5433 = n999 & n5393 ;
  assign n5434 = n5433 ^ n2361 ^ 1'b0 ;
  assign n5435 = n5432 & ~n5434 ;
  assign n5427 = n1450 & n2020 ;
  assign n5428 = n5427 ^ n2310 ^ 1'b0 ;
  assign n5429 = n3680 & n5428 ;
  assign n5430 = ~n2758 & n5429 ;
  assign n5431 = n5430 ^ n5273 ^ n1237 ;
  assign n5436 = n5435 ^ n5431 ^ 1'b0 ;
  assign n5437 = ~n445 & n5436 ;
  assign n5438 = n5437 ^ n1865 ^ 1'b0 ;
  assign n5439 = n400 | n2605 ;
  assign n5440 = n3867 & ~n5030 ;
  assign n5441 = ~n5439 & n5440 ;
  assign n5442 = n765 & n2531 ;
  assign n5444 = n3017 & n3472 ;
  assign n5443 = n983 ^ n204 ^ 1'b0 ;
  assign n5445 = n5444 ^ n5443 ^ 1'b0 ;
  assign n5446 = n2050 ^ n1099 ^ 1'b0 ;
  assign n5447 = n3347 | n3982 ;
  assign n5448 = ~n4948 & n4954 ;
  assign n5449 = n1148 & n5448 ;
  assign n5450 = n586 & ~n1204 ;
  assign n5451 = n5450 ^ n3199 ^ 1'b0 ;
  assign n5452 = n4535 | n5146 ;
  assign n5453 = n1513 ^ n1280 ^ n1192 ;
  assign n5454 = n619 | n2216 ;
  assign n5455 = ~n4302 & n5454 ;
  assign n5456 = n408 & ~n1803 ;
  assign n5458 = n3299 ^ n1732 ^ 1'b0 ;
  assign n5457 = n880 | n3705 ;
  assign n5459 = n5458 ^ n5457 ^ 1'b0 ;
  assign n5460 = n1622 | n5459 ;
  assign n5461 = n2662 | n5460 ;
  assign n5463 = n1699 ^ n950 ^ 1'b0 ;
  assign n5462 = n737 | n5357 ;
  assign n5464 = n5463 ^ n5462 ^ 1'b0 ;
  assign n5465 = n4235 ^ n821 ^ n74 ;
  assign n5466 = n488 & ~n1471 ;
  assign n5467 = ~n1266 & n2637 ;
  assign n5468 = ~n1179 & n4158 ;
  assign n5469 = n340 | n1875 ;
  assign n5470 = n5468 & ~n5469 ;
  assign n5471 = n5470 ^ n3507 ^ 1'b0 ;
  assign n5472 = n1596 | n2976 ;
  assign n5473 = n1552 ^ n1544 ^ 1'b0 ;
  assign n5474 = n5473 ^ n4639 ^ 1'b0 ;
  assign n5475 = n694 | n2652 ;
  assign n5476 = n2346 ^ n1553 ^ 1'b0 ;
  assign n5477 = n2023 & ~n5476 ;
  assign n5478 = n5475 & n5477 ;
  assign n5479 = ( n1251 & n4119 ) | ( n1251 & n5478 ) | ( n4119 & n5478 ) ;
  assign n5480 = n997 ^ n987 ^ 1'b0 ;
  assign n5481 = n3601 | n5480 ;
  assign n5482 = n5481 ^ n4007 ^ 1'b0 ;
  assign n5483 = n418 | n2327 ;
  assign n5484 = ( n425 & n2178 ) | ( n425 & n5483 ) | ( n2178 & n5483 ) ;
  assign n5485 = n5484 ^ n246 ^ 1'b0 ;
  assign n5486 = n3418 & ~n5282 ;
  assign n5487 = n4229 & n5486 ;
  assign n5488 = n2470 ^ n48 ^ 1'b0 ;
  assign n5489 = ~n5030 & n5488 ;
  assign n5490 = ( n582 & n2588 ) | ( n582 & ~n4400 ) | ( n2588 & ~n4400 ) ;
  assign n5491 = n842 | n2236 ;
  assign n5492 = n946 | n5491 ;
  assign n5493 = ~n2771 & n5492 ;
  assign n5494 = n781 & n3848 ;
  assign n5495 = n519 & n5494 ;
  assign n5496 = ~n671 & n2440 ;
  assign n5497 = ~n966 & n5496 ;
  assign n5498 = n3176 | n4910 ;
  assign n5499 = n5497 | n5498 ;
  assign n5500 = n5499 ^ n1709 ^ 1'b0 ;
  assign n5501 = n5495 | n5500 ;
  assign n5502 = n96 & n290 ;
  assign n5503 = ~n722 & n5502 ;
  assign n5504 = n5503 ^ n682 ^ 1'b0 ;
  assign n5505 = n5504 ^ n2859 ^ n2095 ;
  assign n5506 = ~n622 & n5485 ;
  assign n5507 = ~n3191 & n5506 ;
  assign n5508 = ~n1020 & n3333 ;
  assign n5509 = ~n553 & n5197 ;
  assign n5510 = ~n1213 & n5509 ;
  assign n5511 = n2568 ^ n831 ^ 1'b0 ;
  assign n5512 = n2894 | n5511 ;
  assign n5513 = n5512 ^ n4065 ^ 1'b0 ;
  assign n5514 = n1897 & n5513 ;
  assign n5515 = n408 | n456 ;
  assign n5516 = n5515 ^ n1003 ^ 1'b0 ;
  assign n5517 = ( n1237 & n1275 ) | ( n1237 & ~n5516 ) | ( n1275 & ~n5516 ) ;
  assign n5518 = n2205 & n5517 ;
  assign n5519 = n5518 ^ n3240 ^ 1'b0 ;
  assign n5520 = n459 & n3989 ;
  assign n5521 = n5520 ^ n2888 ^ 1'b0 ;
  assign n5522 = n506 | n5521 ;
  assign n5523 = n5519 & n5522 ;
  assign n5524 = n2901 ^ n942 ^ 1'b0 ;
  assign n5525 = n3961 & ~n5524 ;
  assign n5526 = n737 | n2377 ;
  assign n5527 = n357 | n5526 ;
  assign n5528 = n2080 | n5527 ;
  assign n5529 = ~n5122 & n5124 ;
  assign n5530 = n79 & n4722 ;
  assign n5531 = ~n5529 & n5530 ;
  assign n5534 = n162 & ~n2272 ;
  assign n5532 = n1580 & ~n2132 ;
  assign n5533 = n3837 & n5532 ;
  assign n5535 = n5534 ^ n5533 ^ 1'b0 ;
  assign n5537 = n1826 ^ n641 ^ 1'b0 ;
  assign n5538 = n3964 | n5537 ;
  assign n5536 = n3517 | n3573 ;
  assign n5539 = n5538 ^ n5536 ^ 1'b0 ;
  assign n5540 = n5365 ^ n5155 ^ 1'b0 ;
  assign n5541 = n1109 ^ n519 ^ 1'b0 ;
  assign n5542 = ~n2894 & n3897 ;
  assign n5543 = ~n5541 & n5542 ;
  assign n5544 = n5492 ^ n283 ^ 1'b0 ;
  assign n5545 = n1877 ^ n1045 ^ 1'b0 ;
  assign n5546 = ~n2663 & n5545 ;
  assign n5547 = n4485 ^ n3240 ^ 1'b0 ;
  assign n5548 = n1886 ^ n765 ^ 1'b0 ;
  assign n5549 = n4954 & ~n5548 ;
  assign n5550 = ~n3566 & n4511 ;
  assign n5551 = n459 & n5550 ;
  assign n5552 = n4945 ^ n2019 ^ 1'b0 ;
  assign n5553 = n4434 ^ n1104 ^ 1'b0 ;
  assign n5554 = n5553 ^ n49 ^ 1'b0 ;
  assign n5555 = n5554 ^ n2855 ^ 1'b0 ;
  assign n5556 = n4694 ^ n488 ^ 1'b0 ;
  assign n5557 = n2706 & ~n5556 ;
  assign n5560 = n1068 & n4674 ;
  assign n5561 = n5560 ^ n1834 ^ 1'b0 ;
  assign n5558 = n103 & ~n3183 ;
  assign n5559 = n682 & n5558 ;
  assign n5562 = n5561 ^ n5559 ^ 1'b0 ;
  assign n5563 = n2894 ^ n1033 ^ 1'b0 ;
  assign n5564 = n5073 ^ n2541 ^ n1136 ;
  assign n5565 = n841 & ~n5564 ;
  assign n5566 = n5565 ^ n2628 ^ 1'b0 ;
  assign n5567 = ~n1825 & n2673 ;
  assign n5568 = n2053 & ~n5567 ;
  assign n5569 = n2205 & n5568 ;
  assign n5570 = n5569 ^ n3607 ^ 1'b0 ;
  assign n5571 = n4626 ^ n1912 ^ 1'b0 ;
  assign n5572 = n5380 ^ n2677 ^ 1'b0 ;
  assign n5573 = n5572 ^ n5552 ^ n3232 ;
  assign n5574 = n487 | n4030 ;
  assign n5575 = ~n602 & n1208 ;
  assign n5576 = n3112 ^ n2151 ^ n1732 ;
  assign n5577 = n2189 ^ n1755 ^ 1'b0 ;
  assign n5578 = ~n357 & n5577 ;
  assign n5579 = ( ~n1369 & n3301 ) | ( ~n1369 & n5578 ) | ( n3301 & n5578 ) ;
  assign n5580 = n3366 ^ n2445 ^ 1'b0 ;
  assign n5581 = n5580 ^ n4311 ^ 1'b0 ;
  assign n5582 = n1740 & n4006 ;
  assign n5583 = n831 & n5582 ;
  assign n5584 = n5583 ^ n1027 ^ n396 ;
  assign n5585 = n2508 ^ n107 ^ 1'b0 ;
  assign n5586 = n2953 & n5585 ;
  assign n5587 = n5181 & n5586 ;
  assign n5588 = n3121 ^ n2520 ^ 1'b0 ;
  assign n5589 = n3071 & n5588 ;
  assign n5590 = n5589 ^ n1914 ^ 1'b0 ;
  assign n5591 = n3379 & n5590 ;
  assign n5592 = n5226 ^ n3390 ^ n1271 ;
  assign n5593 = n1548 | n3392 ;
  assign n5594 = n2593 ^ n2326 ^ n886 ;
  assign n5598 = n736 ^ n515 ^ 1'b0 ;
  assign n5597 = n1349 | n4103 ;
  assign n5599 = n5598 ^ n5597 ^ 1'b0 ;
  assign n5595 = ( n551 & n4093 ) | ( n551 & ~n4464 ) | ( n4093 & ~n4464 ) ;
  assign n5596 = ~n2283 & n5595 ;
  assign n5600 = n5599 ^ n5596 ^ 1'b0 ;
  assign n5601 = n880 & ~n1656 ;
  assign n5602 = ~n995 & n5601 ;
  assign n5603 = n2995 ^ n1271 ^ 1'b0 ;
  assign n5604 = n3845 | n5603 ;
  assign n5605 = n5604 ^ n2080 ^ 1'b0 ;
  assign n5606 = ~n2288 & n5605 ;
  assign n5607 = n5602 & ~n5606 ;
  assign n5608 = n527 & ~n2859 ;
  assign n5609 = n5608 ^ n3972 ^ 1'b0 ;
  assign n5610 = n3209 & n5236 ;
  assign n5611 = n358 & n1266 ;
  assign n5612 = n5611 ^ n2915 ^ 1'b0 ;
  assign n5613 = ~n5610 & n5612 ;
  assign n5614 = n5613 ^ n434 ^ 1'b0 ;
  assign n5615 = n3441 & n5614 ;
  assign n5618 = n1548 & n2603 ;
  assign n5616 = n2794 ^ n2157 ^ n1611 ;
  assign n5617 = ~n2394 & n5616 ;
  assign n5619 = n5618 ^ n5617 ^ 1'b0 ;
  assign n5620 = n5355 ^ n3195 ^ 1'b0 ;
  assign n5621 = ~n4879 & n5620 ;
  assign n5622 = n1396 | n4529 ;
  assign n5623 = n61 & ~n5622 ;
  assign n5624 = n4579 & ~n4650 ;
  assign n5628 = ( n503 & ~n793 ) | ( n503 & n1420 ) | ( ~n793 & n1420 ) ;
  assign n5629 = n5628 ^ n2861 ^ 1'b0 ;
  assign n5625 = ~n3734 & n3947 ;
  assign n5626 = n155 & n5625 ;
  assign n5627 = n5454 & n5626 ;
  assign n5630 = n5629 ^ n5627 ^ 1'b0 ;
  assign n5631 = n4263 & ~n5286 ;
  assign n5632 = n5631 ^ n760 ^ 1'b0 ;
  assign n5633 = n1342 & ~n3932 ;
  assign n5634 = n188 | n1611 ;
  assign n5635 = n5634 ^ n5249 ^ 1'b0 ;
  assign n5636 = n5633 | n5635 ;
  assign n5637 = n1852 ^ n1567 ^ n302 ;
  assign n5638 = n1978 ^ n1501 ^ 1'b0 ;
  assign n5639 = ~n5637 & n5638 ;
  assign n5640 = n2663 & n3909 ;
  assign n5641 = n1295 & n5640 ;
  assign n5642 = n5641 ^ n3698 ^ 1'b0 ;
  assign n5643 = n2413 ^ n588 ^ 1'b0 ;
  assign n5644 = n1543 & n5643 ;
  assign n5645 = n3167 & n5644 ;
  assign n5646 = n810 | n1050 ;
  assign n5647 = n5646 ^ n3124 ^ n2587 ;
  assign n5648 = n4263 ^ n1016 ^ 1'b0 ;
  assign n5649 = ( n2875 & n4100 ) | ( n2875 & n5648 ) | ( n4100 & n5648 ) ;
  assign n5650 = n44 & ~n4668 ;
  assign n5651 = n2971 & n5650 ;
  assign n5652 = n307 ^ n288 ^ 1'b0 ;
  assign n5653 = n2985 & n3954 ;
  assign n5654 = ~n5652 & n5653 ;
  assign n5655 = n3818 | n5654 ;
  assign n5656 = n3482 ^ n1280 ^ 1'b0 ;
  assign n5657 = n910 ^ n406 ^ 1'b0 ;
  assign n5658 = n1184 & ~n5657 ;
  assign n5659 = n527 & n5658 ;
  assign n5660 = n2337 & n5659 ;
  assign n5661 = n1738 | n5660 ;
  assign n5662 = n5217 | n5661 ;
  assign n5663 = n5662 ^ n4997 ^ 1'b0 ;
  assign n5664 = ~n5656 & n5663 ;
  assign n5665 = n2058 ^ n522 ^ 1'b0 ;
  assign n5666 = ~n2852 & n5665 ;
  assign n5667 = ~n58 & n5666 ;
  assign n5668 = ~n968 & n5667 ;
  assign n5670 = n1814 & n1853 ;
  assign n5671 = n2474 & n5670 ;
  assign n5669 = n398 & n1670 ;
  assign n5672 = n5671 ^ n5669 ^ 1'b0 ;
  assign n5673 = n2092 ^ n755 ^ 1'b0 ;
  assign n5674 = n3537 ^ n477 ^ 1'b0 ;
  assign n5675 = n5167 & n5674 ;
  assign n5676 = n126 | n3932 ;
  assign n5677 = n3287 ^ n477 ^ 1'b0 ;
  assign n5678 = n2321 & ~n3064 ;
  assign n5679 = ~n5390 & n5678 ;
  assign n5680 = ~n3228 & n5679 ;
  assign n5681 = ~n1240 & n4074 ;
  assign n5682 = ( ~n1297 & n5328 ) | ( ~n1297 & n5681 ) | ( n5328 & n5681 ) ;
  assign n5683 = ~n508 & n5682 ;
  assign n5684 = ~n1371 & n5683 ;
  assign n5685 = n2753 ^ n652 ^ 1'b0 ;
  assign n5686 = n61 & ~n4849 ;
  assign n5687 = n5686 ^ n5079 ^ n601 ;
  assign n5688 = ~n983 & n1949 ;
  assign n5689 = ( n437 & n894 ) | ( n437 & n5688 ) | ( n894 & n5688 ) ;
  assign n5690 = n5689 ^ n4984 ^ 1'b0 ;
  assign n5691 = n3940 & n5690 ;
  assign n5692 = n1599 ^ n98 ^ 1'b0 ;
  assign n5693 = n5168 ^ n3137 ^ n2522 ;
  assign n5694 = n3731 & ~n5693 ;
  assign n5695 = ~n5692 & n5694 ;
  assign n5696 = ~n372 & n611 ;
  assign n5697 = n5696 ^ n2550 ^ 1'b0 ;
  assign n5698 = n4036 & ~n5697 ;
  assign n5699 = n5698 ^ n4622 ^ 1'b0 ;
  assign n5700 = n2790 | n4751 ;
  assign n5701 = n1749 ^ n1694 ^ 1'b0 ;
  assign n5702 = n539 | n5701 ;
  assign n5703 = n3086 & n5702 ;
  assign n5704 = ~n1697 & n5703 ;
  assign n5705 = n1182 & n3586 ;
  assign n5706 = n5705 ^ x6 ^ 1'b0 ;
  assign n5707 = n2935 ^ n1772 ^ 1'b0 ;
  assign n5708 = n5707 ^ n181 ^ 1'b0 ;
  assign n5709 = ~n694 & n5708 ;
  assign n5710 = n2901 & n5709 ;
  assign n5711 = n3544 ^ n1251 ^ 1'b0 ;
  assign n5714 = n360 | n1904 ;
  assign n5712 = n2065 ^ n205 ^ 1'b0 ;
  assign n5713 = ~n717 & n5712 ;
  assign n5715 = n5714 ^ n5713 ^ 1'b0 ;
  assign n5716 = n5711 | n5715 ;
  assign n5717 = n1202 & ~n5716 ;
  assign n5718 = ~n1997 & n4207 ;
  assign n5719 = n1573 & n5718 ;
  assign n5720 = n1550 & ~n5719 ;
  assign n5721 = ~n4546 & n5720 ;
  assign n5722 = n884 ^ n785 ^ 1'b0 ;
  assign n5723 = n5722 ^ n3947 ^ 1'b0 ;
  assign n5724 = n5721 | n5723 ;
  assign n5725 = n219 & n1546 ;
  assign n5726 = n5725 ^ n3428 ^ 1'b0 ;
  assign n5727 = n1291 ^ n539 ^ 1'b0 ;
  assign n5728 = n4838 ^ n4808 ^ 1'b0 ;
  assign n5729 = n191 | n5728 ;
  assign n5730 = n5727 & ~n5729 ;
  assign n5731 = n5429 | n5538 ;
  assign n5732 = n2045 ^ n967 ^ 1'b0 ;
  assign n5733 = ~n1396 & n5732 ;
  assign n5734 = n5733 ^ n3805 ^ 1'b0 ;
  assign n5736 = n130 & ~n2304 ;
  assign n5737 = n2104 ^ n421 ^ 1'b0 ;
  assign n5738 = n5736 & ~n5737 ;
  assign n5735 = n1216 & n1230 ;
  assign n5739 = n5738 ^ n5735 ^ 1'b0 ;
  assign n5740 = n3384 ^ n2850 ^ 1'b0 ;
  assign n5741 = n2048 ^ n390 ^ 1'b0 ;
  assign n5742 = n5741 ^ n1915 ^ 1'b0 ;
  assign n5743 = n5740 & ~n5742 ;
  assign n5744 = n27 | n1439 ;
  assign n5745 = ~n4843 & n5744 ;
  assign n5746 = ~n2927 & n5393 ;
  assign n5747 = n5746 ^ n263 ^ 1'b0 ;
  assign n5748 = n1305 & n1445 ;
  assign n5749 = ~n5747 & n5748 ;
  assign n5750 = ( n2431 & n3278 ) | ( n2431 & n4025 ) | ( n3278 & n4025 ) ;
  assign n5751 = ~n25 & n5702 ;
  assign n5752 = n108 | n2946 ;
  assign n5753 = n5437 | n5752 ;
  assign n5754 = n1283 & ~n1685 ;
  assign n5755 = n125 & n5754 ;
  assign n5756 = n646 & ~n1363 ;
  assign n5757 = ( n2432 & n2468 ) | ( n2432 & n5756 ) | ( n2468 & n5756 ) ;
  assign n5758 = n645 & ~n5757 ;
  assign n5759 = ( ~n1741 & n5755 ) | ( ~n1741 & n5758 ) | ( n5755 & n5758 ) ;
  assign n5760 = n826 & n5759 ;
  assign n5761 = n3738 ^ n2362 ^ 1'b0 ;
  assign n5762 = ~n2560 & n5761 ;
  assign n5763 = ( n3690 & ~n3990 ) | ( n3690 & n5573 ) | ( ~n3990 & n5573 ) ;
  assign n5764 = n2603 ^ n27 ^ 1'b0 ;
  assign n5765 = n1200 & ~n5764 ;
  assign n5766 = n4321 & n5765 ;
  assign n5767 = n5766 ^ n5546 ^ n2861 ;
  assign n5768 = n2637 ^ n2138 ^ 1'b0 ;
  assign n5769 = n1656 ^ n1576 ^ 1'b0 ;
  assign n5770 = n2529 | n5224 ;
  assign n5771 = n5769 | n5770 ;
  assign n5772 = n4331 ^ n2491 ^ 1'b0 ;
  assign n5773 = n2568 & ~n5772 ;
  assign n5780 = n2038 ^ n279 ^ 1'b0 ;
  assign n5781 = n1878 | n5780 ;
  assign n5777 = n255 & ~n2406 ;
  assign n5778 = n4143 & n5777 ;
  assign n5774 = n2670 ^ n354 ^ 1'b0 ;
  assign n5775 = ~n3696 & n5774 ;
  assign n5776 = ~n3700 & n5775 ;
  assign n5779 = n5778 ^ n5776 ^ 1'b0 ;
  assign n5782 = n5781 ^ n5779 ^ 1'b0 ;
  assign n5783 = ~n5042 & n5782 ;
  assign n5784 = n280 & n5027 ;
  assign n5785 = ~n4690 & n5784 ;
  assign n5786 = n1592 ^ n1543 ^ 1'b0 ;
  assign n5787 = n38 & n277 ;
  assign n5788 = n5787 ^ n1763 ^ 1'b0 ;
  assign n5789 = n5786 & n5788 ;
  assign n5790 = n1508 ^ n1269 ^ 1'b0 ;
  assign n5791 = n1377 | n5790 ;
  assign n5792 = n2473 | n5791 ;
  assign n5793 = n5792 ^ n2090 ^ 1'b0 ;
  assign n5794 = n1617 ^ n154 ^ 1'b0 ;
  assign n5795 = n1087 | n5794 ;
  assign n5796 = ~n1349 & n1366 ;
  assign n5797 = n5796 ^ n74 ^ 1'b0 ;
  assign n5798 = n2850 ^ n1753 ^ 1'b0 ;
  assign n5799 = ( n638 & ~n5571 ) | ( n638 & n5798 ) | ( ~n5571 & n5798 ) ;
  assign n5800 = n1685 & n4855 ;
  assign n5801 = n5800 ^ n4063 ^ 1'b0 ;
  assign n5802 = n2603 ^ n765 ^ n489 ;
  assign n5803 = n5802 ^ n3764 ^ 1'b0 ;
  assign n5804 = n3866 ^ n362 ^ 1'b0 ;
  assign n5805 = ~n3791 & n5804 ;
  assign n5806 = n5805 ^ n1182 ^ n142 ;
  assign n5807 = n140 | n5806 ;
  assign n5808 = n4341 ^ n725 ^ 1'b0 ;
  assign n5809 = n96 & n5808 ;
  assign n5810 = n5809 ^ n3153 ^ 1'b0 ;
  assign n5811 = n4525 & ~n5758 ;
  assign n5812 = n5532 & ~n5811 ;
  assign n5813 = n482 & ~n559 ;
  assign n5814 = ~n1142 & n5813 ;
  assign n5815 = n790 & n1395 ;
  assign n5816 = n2918 & ~n5815 ;
  assign n5817 = n5395 ^ n3114 ^ 1'b0 ;
  assign n5818 = ~n564 & n5817 ;
  assign n5819 = n2340 & ~n3977 ;
  assign n5823 = n584 & ~n1694 ;
  assign n5824 = n1157 & n5823 ;
  assign n5825 = n1590 & ~n5824 ;
  assign n5826 = n1374 ^ n999 ^ 1'b0 ;
  assign n5827 = n5825 | n5826 ;
  assign n5820 = n5417 ^ n2343 ^ 1'b0 ;
  assign n5821 = ~n840 & n5820 ;
  assign n5822 = n2358 & n5821 ;
  assign n5828 = n5827 ^ n5822 ^ 1'b0 ;
  assign n5829 = n1002 & ~n5828 ;
  assign n5830 = n5809 ^ n1821 ^ 1'b0 ;
  assign n5831 = ~n244 & n5830 ;
  assign n5832 = ~n1271 & n5831 ;
  assign n5833 = n1941 | n2435 ;
  assign n5834 = n530 & ~n4179 ;
  assign n5835 = n5833 & ~n5834 ;
  assign n5836 = n3658 ^ n27 ^ 1'b0 ;
  assign n5842 = n4545 ^ n1960 ^ 1'b0 ;
  assign n5843 = n5357 ^ n3667 ^ 1'b0 ;
  assign n5844 = ~n5842 & n5843 ;
  assign n5837 = ~n1845 & n2888 ;
  assign n5838 = ~n481 & n1504 ;
  assign n5839 = n894 & n5838 ;
  assign n5840 = n5839 ^ n2337 ^ n560 ;
  assign n5841 = n5837 & ~n5840 ;
  assign n5845 = n5844 ^ n5841 ^ 1'b0 ;
  assign n5846 = n3066 & ~n5779 ;
  assign n5847 = n5846 ^ n2391 ^ 1'b0 ;
  assign n5848 = n2723 ^ n2377 ^ 1'b0 ;
  assign n5849 = ~n997 & n5848 ;
  assign n5850 = ~n4105 & n5381 ;
  assign n5851 = ~n1915 & n3647 ;
  assign n5852 = n819 ^ n508 ^ 1'b0 ;
  assign n5853 = n3167 | n5852 ;
  assign n5854 = n5853 ^ n3037 ^ 1'b0 ;
  assign n5855 = n103 & n920 ;
  assign n5856 = ~n5854 & n5855 ;
  assign n5857 = n1077 & ~n5856 ;
  assign n5858 = n1491 | n2228 ;
  assign n5859 = n5858 ^ n4148 ^ 1'b0 ;
  assign n5860 = n5859 ^ n5037 ^ 1'b0 ;
  assign n5861 = n1969 & n5860 ;
  assign n5862 = n1466 | n5504 ;
  assign n5863 = n5862 ^ n438 ^ 1'b0 ;
  assign n5864 = n889 & n5553 ;
  assign n5865 = n205 | n1951 ;
  assign n5866 = n5865 ^ n2163 ^ n296 ;
  assign n5867 = n5866 ^ n508 ^ 1'b0 ;
  assign n5868 = ~n1918 & n5028 ;
  assign n5869 = n1936 ^ n67 ^ 1'b0 ;
  assign n5870 = n4208 & n5869 ;
  assign n5871 = n2216 & n5870 ;
  assign n5872 = ( ~n479 & n1110 ) | ( ~n479 & n1371 ) | ( n1110 & n1371 ) ;
  assign n5873 = n5360 & ~n5872 ;
  assign n5874 = n396 ^ n23 ^ 1'b0 ;
  assign n5875 = n1458 & n5874 ;
  assign n5876 = ~n2332 & n5875 ;
  assign n5877 = n874 & n5876 ;
  assign n5878 = n2925 ^ n2588 ^ 1'b0 ;
  assign n5879 = ~n2772 & n5878 ;
  assign n5880 = n3145 & ~n3759 ;
  assign n5881 = ~n917 & n2397 ;
  assign n5882 = n224 | n1908 ;
  assign n5883 = n160 | n5882 ;
  assign n5884 = n81 & n5883 ;
  assign n5885 = ~n5881 & n5884 ;
  assign n5886 = n222 & n2626 ;
  assign n5887 = n171 | n5886 ;
  assign n5888 = n5887 ^ n1717 ^ 1'b0 ;
  assign n5889 = n4720 & n5888 ;
  assign n5890 = n5885 & n5889 ;
  assign n5891 = n4312 ^ n3021 ^ 1'b0 ;
  assign n5892 = n4671 & ~n5891 ;
  assign n5893 = n5071 ^ n1570 ^ 1'b0 ;
  assign n5894 = n5893 ^ n3325 ^ 1'b0 ;
  assign n5895 = ~n4259 & n5894 ;
  assign n5896 = ~n5892 & n5895 ;
  assign n5897 = n1673 | n2955 ;
  assign n5906 = n4079 ^ n1062 ^ 1'b0 ;
  assign n5899 = n694 ^ n521 ^ 1'b0 ;
  assign n5900 = ~n368 & n5899 ;
  assign n5901 = n1322 & n5900 ;
  assign n5898 = n1569 ^ n563 ^ 1'b0 ;
  assign n5902 = n5901 ^ n5898 ^ n2796 ;
  assign n5903 = n5354 ^ n1636 ^ 1'b0 ;
  assign n5904 = n1732 & n5903 ;
  assign n5905 = n5902 & n5904 ;
  assign n5907 = n5906 ^ n5905 ^ 1'b0 ;
  assign n5908 = ~n5302 & n5907 ;
  assign n5909 = n4967 ^ n4539 ^ 1'b0 ;
  assign n5910 = ~n384 & n598 ;
  assign n5911 = n5910 ^ n2040 ^ 1'b0 ;
  assign n5912 = n5909 | n5911 ;
  assign n5913 = n339 & ~n1493 ;
  assign n5914 = ~n200 & n5913 ;
  assign n5915 = n503 | n5914 ;
  assign n5916 = n3774 ^ n968 ^ 1'b0 ;
  assign n5917 = n5916 ^ n4849 ^ 1'b0 ;
  assign n5918 = n362 & ~n439 ;
  assign n5919 = n3044 & n5918 ;
  assign n5920 = n5919 ^ n1742 ^ 1'b0 ;
  assign n5921 = ( n2943 & n3280 ) | ( n2943 & ~n5920 ) | ( n3280 & ~n5920 ) ;
  assign n5922 = n2377 | n2474 ;
  assign n5923 = n2474 & ~n5922 ;
  assign n5924 = n562 | n2291 ;
  assign n5925 = n5924 ^ n2727 ^ 1'b0 ;
  assign n5926 = ~n5923 & n5925 ;
  assign n5927 = n5923 & n5926 ;
  assign n5928 = ~n2184 & n4588 ;
  assign n5929 = n2635 & n5928 ;
  assign n5930 = ( n43 & ~n1237 ) | ( n43 & n5929 ) | ( ~n1237 & n5929 ) ;
  assign n5931 = n5927 | n5930 ;
  assign n5932 = n5931 ^ n5868 ^ 1'b0 ;
  assign n5933 = n551 | n3374 ;
  assign n5934 = n3450 & ~n3985 ;
  assign n5935 = ~n2425 & n5934 ;
  assign n5936 = n3756 & ~n5935 ;
  assign n5937 = n2930 & ~n2958 ;
  assign n5938 = n93 | n132 ;
  assign n5939 = n1387 & ~n1872 ;
  assign n5940 = n5938 & ~n5939 ;
  assign n5941 = n5940 ^ n3389 ^ 1'b0 ;
  assign n5942 = ~n2820 & n5941 ;
  assign n5943 = n5942 ^ n4233 ^ 1'b0 ;
  assign n5944 = n5937 & ~n5943 ;
  assign n5945 = n1701 & ~n5944 ;
  assign n5946 = n5629 ^ n2743 ^ n347 ;
  assign n5947 = n2072 & ~n4108 ;
  assign n5948 = ~n5012 & n5947 ;
  assign n5949 = n3475 & n4748 ;
  assign n5950 = n2283 & n5949 ;
  assign n5951 = ~n801 & n1821 ;
  assign n5952 = n5951 ^ n804 ^ 1'b0 ;
  assign n5953 = n5952 ^ n3052 ^ 1'b0 ;
  assign n5954 = n4117 ^ n2924 ^ n395 ;
  assign n5955 = n414 | n1392 ;
  assign n5956 = n5954 & ~n5955 ;
  assign n5957 = ( n402 & ~n2394 ) | ( n402 & n3315 ) | ( ~n2394 & n3315 ) ;
  assign n5958 = n5957 ^ n3537 ^ 1'b0 ;
  assign n5959 = n1140 & ~n1438 ;
  assign n5960 = n1383 & ~n2397 ;
  assign n5961 = n5960 ^ n1540 ^ 1'b0 ;
  assign n5962 = n1975 | n5961 ;
  assign n5963 = n5962 ^ n1263 ^ 1'b0 ;
  assign n5964 = n1591 ^ n267 ^ 1'b0 ;
  assign n5965 = n5963 & n5964 ;
  assign n5966 = n5959 & n5965 ;
  assign n5967 = n5966 ^ n817 ^ 1'b0 ;
  assign n5968 = n3856 | n4474 ;
  assign n5969 = n2408 | n5968 ;
  assign n5970 = n4913 ^ n2610 ^ 1'b0 ;
  assign n5971 = n2656 & n4142 ;
  assign n5972 = n1264 & ~n4390 ;
  assign n5973 = ~n2315 & n5972 ;
  assign n5974 = n5973 ^ n3449 ^ 1'b0 ;
  assign n5975 = n184 | n563 ;
  assign n5976 = n5975 ^ n539 ^ 1'b0 ;
  assign n5977 = n5976 ^ n2270 ^ 1'b0 ;
  assign n5978 = n4063 | n5977 ;
  assign n5979 = n880 & n1910 ;
  assign n5980 = ~n1104 & n5979 ;
  assign n5981 = ( n229 & n645 ) | ( n229 & ~n1459 ) | ( n645 & ~n1459 ) ;
  assign n5982 = n3257 & ~n5981 ;
  assign n5983 = n2833 & n5234 ;
  assign n5984 = n5983 ^ n362 ^ 1'b0 ;
  assign n5985 = ~n541 & n3580 ;
  assign n5986 = n5985 ^ n43 ^ 1'b0 ;
  assign n5988 = n3609 ^ n3052 ^ 1'b0 ;
  assign n5987 = ~n5293 & n5380 ;
  assign n5989 = n5988 ^ n5987 ^ 1'b0 ;
  assign n5990 = n782 & n3333 ;
  assign n5991 = n5990 ^ n3442 ^ 1'b0 ;
  assign n5992 = n5991 ^ n3800 ^ 1'b0 ;
  assign n5993 = ~n5641 & n5992 ;
  assign n5994 = ~n2290 & n5993 ;
  assign n5995 = n4685 ^ n3634 ^ 1'b0 ;
  assign n5996 = ~n2492 & n3961 ;
  assign n5997 = n5996 ^ n3257 ^ 1'b0 ;
  assign n5998 = n620 | n4039 ;
  assign n5999 = n5998 ^ n823 ^ 1'b0 ;
  assign n6000 = ( n911 & ~n5997 ) | ( n911 & n5999 ) | ( ~n5997 & n5999 ) ;
  assign n6001 = ~n4008 & n4778 ;
  assign n6002 = n5914 ^ n1349 ^ 1'b0 ;
  assign n6006 = n2226 | n2568 ;
  assign n6003 = n1999 ^ n349 ^ 1'b0 ;
  assign n6004 = n4809 ^ n2349 ^ 1'b0 ;
  assign n6005 = n6003 & ~n6004 ;
  assign n6007 = n6006 ^ n6005 ^ 1'b0 ;
  assign n6008 = ~n1054 & n2794 ;
  assign n6009 = n3837 & n6008 ;
  assign n6011 = n1546 ^ n1535 ^ 1'b0 ;
  assign n6010 = n1618 & ~n4169 ;
  assign n6012 = n6011 ^ n6010 ^ 1'b0 ;
  assign n6013 = n2532 | n2664 ;
  assign n6014 = n6013 ^ n1884 ^ 1'b0 ;
  assign n6015 = n6012 | n6014 ;
  assign n6016 = n5288 & ~n5628 ;
  assign n6017 = n3255 ^ n492 ^ 1'b0 ;
  assign n6018 = n4510 & ~n6017 ;
  assign n6019 = ~n140 & n3445 ;
  assign n6020 = ~n1104 & n5936 ;
  assign n6021 = n3542 ^ n2178 ^ 1'b0 ;
  assign n6022 = n546 | n2779 ;
  assign n6023 = n6021 & ~n6022 ;
  assign n6024 = n6020 | n6023 ;
  assign n6025 = ( n438 & n2548 ) | ( n438 & n3384 ) | ( n2548 & n3384 ) ;
  assign n6026 = n6025 ^ n1340 ^ 1'b0 ;
  assign n6027 = n1391 | n1655 ;
  assign n6028 = n6027 ^ n560 ^ 1'b0 ;
  assign n6029 = n96 & ~n6028 ;
  assign n6030 = n4962 ^ n4826 ^ 1'b0 ;
  assign n6031 = n6030 ^ n4364 ^ 1'b0 ;
  assign n6032 = n6029 & ~n6031 ;
  assign n6033 = n5821 ^ n1997 ^ 1'b0 ;
  assign n6034 = n1119 ^ n980 ^ 1'b0 ;
  assign n6035 = n517 & ~n6034 ;
  assign n6036 = n3840 & n5989 ;
  assign n6037 = n2593 & n3027 ;
  assign n6038 = n2201 & ~n6037 ;
  assign n6039 = n468 & n4704 ;
  assign n6041 = n1506 | n3826 ;
  assign n6040 = n3651 ^ n1152 ^ 1'b0 ;
  assign n6042 = n6041 ^ n6040 ^ n938 ;
  assign n6043 = n6042 ^ n5406 ^ 1'b0 ;
  assign n6044 = n1789 ^ n598 ^ 1'b0 ;
  assign n6045 = n306 & ~n6044 ;
  assign n6046 = n5174 ^ n363 ^ 1'b0 ;
  assign n6047 = n6045 & ~n6046 ;
  assign n6048 = ( ~n117 & n901 ) | ( ~n117 & n1556 ) | ( n901 & n1556 ) ;
  assign n6049 = n6047 & n6048 ;
  assign n6050 = n1083 & n6049 ;
  assign n6051 = ~n2829 & n6050 ;
  assign n6052 = n5470 ^ n4667 ^ 1'b0 ;
  assign n6053 = n2097 ^ n362 ^ 1'b0 ;
  assign n6054 = n5216 & ~n6053 ;
  assign n6057 = n3390 ^ n2166 ^ n21 ;
  assign n6055 = n2446 ^ n1172 ^ 1'b0 ;
  assign n6056 = n3884 & ~n6055 ;
  assign n6058 = n6057 ^ n6056 ^ 1'b0 ;
  assign n6059 = n488 & ~n631 ;
  assign n6060 = n6059 ^ n3864 ^ 1'b0 ;
  assign n6061 = n1800 & ~n5579 ;
  assign n6062 = n2973 & n6061 ;
  assign n6063 = n6062 ^ n2746 ^ 1'b0 ;
  assign n6064 = n2575 ^ n294 ^ 1'b0 ;
  assign n6065 = n2403 | n6064 ;
  assign n6066 = n2218 ^ n1047 ^ 1'b0 ;
  assign n6067 = ~n122 & n6066 ;
  assign n6068 = ~n6065 & n6067 ;
  assign n6069 = n4712 & n6068 ;
  assign n6070 = ~n535 & n2423 ;
  assign n6071 = n2960 ^ n1155 ^ 1'b0 ;
  assign n6072 = n365 & n5491 ;
  assign n6073 = n6072 ^ n1908 ^ 1'b0 ;
  assign n6074 = n6071 | n6073 ;
  assign n6075 = n2377 ^ n1590 ^ 1'b0 ;
  assign n6076 = n3312 & ~n4523 ;
  assign n6077 = ~n3691 & n6076 ;
  assign n6078 = n6077 ^ n312 ^ 1'b0 ;
  assign n6079 = n6075 & n6078 ;
  assign n6080 = n1586 ^ n582 ^ 1'b0 ;
  assign n6081 = ~n3866 & n6058 ;
  assign n6082 = ~n785 & n3502 ;
  assign n6083 = ~n1473 & n5547 ;
  assign n6087 = ~n831 & n5601 ;
  assign n6088 = n148 & n6087 ;
  assign n6089 = n6088 ^ n2749 ^ 1'b0 ;
  assign n6090 = n86 & ~n6089 ;
  assign n6091 = n982 & n6090 ;
  assign n6092 = n6091 ^ n3738 ^ 1'b0 ;
  assign n6093 = n3724 | n6092 ;
  assign n6084 = n2038 | n5107 ;
  assign n6085 = n4036 | n6084 ;
  assign n6086 = n833 & ~n6085 ;
  assign n6094 = n6093 ^ n6086 ^ 1'b0 ;
  assign n6095 = n707 & n2381 ;
  assign n6096 = n565 & ~n4657 ;
  assign n6097 = n6095 | n6096 ;
  assign n6098 = n6097 ^ n3098 ^ 1'b0 ;
  assign n6099 = n126 & ~n1119 ;
  assign n6100 = n506 & ~n6099 ;
  assign n6101 = ~n749 & n1953 ;
  assign n6102 = n1280 & ~n6101 ;
  assign n6103 = ( n3562 & n4341 ) | ( n3562 & ~n5357 ) | ( n4341 & ~n5357 ) ;
  assign n6104 = n3516 & n3621 ;
  assign n6105 = n3891 & n6104 ;
  assign n6106 = ~n6103 & n6105 ;
  assign n6107 = n192 | n887 ;
  assign n6108 = n1073 & ~n6107 ;
  assign n6109 = n357 | n6108 ;
  assign n6110 = n1744 | n6109 ;
  assign n6111 = n2189 & n6110 ;
  assign n6112 = n5549 ^ n372 ^ 1'b0 ;
  assign n6113 = ~n1594 & n2371 ;
  assign n6114 = ~n74 & n6113 ;
  assign n6115 = n2358 & ~n6114 ;
  assign n6116 = n6115 ^ n703 ^ 1'b0 ;
  assign n6117 = n6116 ^ n998 ^ n513 ;
  assign n6118 = n1941 & n6117 ;
  assign n6119 = ~n723 & n6118 ;
  assign n6120 = n6119 ^ n1845 ^ 1'b0 ;
  assign n6121 = n2675 & ~n6120 ;
  assign n6122 = n5641 ^ n4982 ^ 1'b0 ;
  assign n6123 = n6122 ^ n5898 ^ 1'b0 ;
  assign n6124 = n397 | n6123 ;
  assign n6125 = n509 & n2155 ;
  assign n6126 = n6125 ^ n808 ^ n423 ;
  assign n6127 = ~n2745 & n3599 ;
  assign n6128 = ~n808 & n985 ;
  assign n6129 = n929 & n5008 ;
  assign n6130 = n1217 & n6129 ;
  assign n6131 = n663 & n6130 ;
  assign n6132 = n5352 ^ n299 ^ 1'b0 ;
  assign n6133 = ( ~n854 & n2472 ) | ( ~n854 & n6132 ) | ( n2472 & n6132 ) ;
  assign n6134 = ~n48 & n6133 ;
  assign n6135 = ~n5151 & n6134 ;
  assign n6136 = n5010 ^ n4275 ^ n1794 ;
  assign n6137 = n1411 | n1711 ;
  assign n6138 = n1390 & ~n6137 ;
  assign n6139 = n6138 ^ n1544 ^ 1'b0 ;
  assign n6140 = n968 & ~n6139 ;
  assign n6141 = ~n205 & n1618 ;
  assign n6142 = n6141 ^ n1877 ^ 1'b0 ;
  assign n6143 = n260 & n1991 ;
  assign n6144 = ~n681 & n6143 ;
  assign n6145 = ~n1323 & n6144 ;
  assign n6146 = n2419 & ~n2736 ;
  assign n6147 = n6145 & n6146 ;
  assign n6148 = n4999 ^ n2319 ^ 1'b0 ;
  assign n6149 = n2317 & ~n6148 ;
  assign n6150 = n1327 & ~n3959 ;
  assign n6151 = ~n6149 & n6150 ;
  assign n6152 = n2650 & ~n6151 ;
  assign n6153 = n6152 ^ n3594 ^ 1'b0 ;
  assign n6154 = n6153 ^ n5139 ^ 1'b0 ;
  assign n6155 = n25 & ~n2094 ;
  assign n6156 = n6155 ^ n1308 ^ 1'b0 ;
  assign n6157 = n1477 ^ n521 ^ 1'b0 ;
  assign n6158 = n547 & ~n2560 ;
  assign n6159 = ~n6157 & n6158 ;
  assign n6160 = ~n1103 & n1208 ;
  assign n6161 = n6160 ^ n4360 ^ 1'b0 ;
  assign n6162 = ~n2885 & n6161 ;
  assign n6163 = n2138 ^ n1080 ^ 1'b0 ;
  assign n6164 = n1485 & n6163 ;
  assign n6165 = ~n4394 & n4605 ;
  assign n6166 = n5646 ^ n1865 ^ 1'b0 ;
  assign n6167 = ~n1908 & n3688 ;
  assign n6168 = n5566 & n6167 ;
  assign n6169 = n3245 & ~n4116 ;
  assign n6170 = n2507 & n6169 ;
  assign n6171 = n4291 & ~n6170 ;
  assign n6172 = ~n2641 & n6171 ;
  assign n6173 = n6172 ^ n86 ^ 1'b0 ;
  assign n6174 = ~n2267 & n6173 ;
  assign n6175 = ~n1223 & n6174 ;
  assign n6176 = n917 ^ n798 ^ 1'b0 ;
  assign n6177 = n4457 & ~n6176 ;
  assign n6178 = n3794 ^ n376 ^ 1'b0 ;
  assign n6179 = ~n3602 & n6178 ;
  assign n6180 = n3412 & ~n6179 ;
  assign n6181 = n1983 ^ n931 ^ 1'b0 ;
  assign n6182 = n2104 | n4539 ;
  assign n6183 = n3971 | n6182 ;
  assign n6184 = ~n162 & n4080 ;
  assign n6185 = n2460 ^ n318 ^ 1'b0 ;
  assign n6186 = n1405 | n2022 ;
  assign n6187 = n6186 ^ n1321 ^ 1'b0 ;
  assign n6188 = ~n6185 & n6187 ;
  assign n6189 = n1080 & n6188 ;
  assign n6190 = n1832 | n5861 ;
  assign n6191 = n1918 ^ n1003 ^ 1'b0 ;
  assign n6192 = n1921 & n6191 ;
  assign n6193 = n6192 ^ n3155 ^ 1'b0 ;
  assign n6194 = ~n3729 & n6193 ;
  assign n6195 = n2413 & n6194 ;
  assign n6201 = n936 & n3680 ;
  assign n6202 = ~n4102 & n6201 ;
  assign n6203 = ~n1920 & n6202 ;
  assign n6196 = n892 & n2034 ;
  assign n6197 = n854 | n6196 ;
  assign n6198 = x7 | n6197 ;
  assign n6199 = ~n184 & n6198 ;
  assign n6200 = n6199 ^ n3912 ^ 1'b0 ;
  assign n6204 = n6203 ^ n6200 ^ 1'b0 ;
  assign n6205 = n4169 | n6204 ;
  assign n6206 = n1045 & ~n2367 ;
  assign n6213 = n1691 ^ n360 ^ 1'b0 ;
  assign n6207 = n2403 ^ n2124 ^ 1'b0 ;
  assign n6208 = ~n2680 & n6207 ;
  assign n6209 = ~n959 & n2660 ;
  assign n6210 = ~n3333 & n6209 ;
  assign n6211 = n6208 & ~n6210 ;
  assign n6212 = n6211 ^ n5324 ^ 1'b0 ;
  assign n6214 = n6213 ^ n6212 ^ 1'b0 ;
  assign n6215 = ~n6206 & n6214 ;
  assign n6216 = ~n878 & n2618 ;
  assign n6217 = n3302 ^ n1377 ^ 1'b0 ;
  assign n6218 = n495 & n5971 ;
  assign n6219 = n194 | n1058 ;
  assign n6220 = n2971 | n6219 ;
  assign n6221 = n6220 ^ n1199 ^ 1'b0 ;
  assign n6222 = n56 & n910 ;
  assign n6223 = ~n220 & n6222 ;
  assign n6224 = n1320 | n6223 ;
  assign n6225 = ( n2811 & ~n5395 ) | ( n2811 & n6224 ) | ( ~n5395 & n6224 ) ;
  assign n6226 = n2700 ^ n854 ^ 1'b0 ;
  assign n6227 = n1933 & n6226 ;
  assign n6228 = ~n3127 & n3358 ;
  assign n6229 = n149 & ~n6228 ;
  assign n6230 = n1929 & ~n4988 ;
  assign n6231 = n1266 ^ n848 ^ 1'b0 ;
  assign n6232 = n6231 ^ n3894 ^ 1'b0 ;
  assign n6233 = n5564 ^ n3050 ^ n2821 ;
  assign n6234 = ( ~n3602 & n6232 ) | ( ~n3602 & n6233 ) | ( n6232 & n6233 ) ;
  assign n6235 = n1207 & ~n1726 ;
  assign n6236 = n4506 ^ n2253 ^ n327 ;
  assign n6237 = n1878 ^ n271 ^ 1'b0 ;
  assign n6238 = n2995 & ~n6237 ;
  assign n6239 = n1181 | n2855 ;
  assign n6240 = n2352 | n6239 ;
  assign n6241 = n6240 ^ n2283 ^ n1298 ;
  assign n6242 = n2277 & ~n3484 ;
  assign n6243 = n6242 ^ n2166 ^ 1'b0 ;
  assign n6246 = n249 & n2884 ;
  assign n6247 = ~n4859 & n6246 ;
  assign n6244 = n1536 ^ n428 ^ 1'b0 ;
  assign n6245 = n3449 | n6244 ;
  assign n6248 = n6247 ^ n6245 ^ n924 ;
  assign n6249 = n6248 ^ n91 ^ 1'b0 ;
  assign n6250 = n6243 & n6249 ;
  assign n6251 = n5345 ^ n228 ^ 1'b0 ;
  assign n6252 = n3569 | n6251 ;
  assign n6253 = n1497 & ~n4732 ;
  assign n6254 = n4653 & n6253 ;
  assign n6255 = n6254 ^ n4740 ^ 1'b0 ;
  assign n6256 = n2721 ^ n2691 ^ 1'b0 ;
  assign n6257 = n3849 ^ n2664 ^ 1'b0 ;
  assign n6258 = ( ~n971 & n3968 ) | ( ~n971 & n5682 ) | ( n3968 & n5682 ) ;
  assign n6259 = n4228 | n4740 ;
  assign n6260 = n44 & n6259 ;
  assign n6261 = ~n1032 & n6260 ;
  assign n6262 = n1087 ^ n625 ^ 1'b0 ;
  assign n6263 = n3989 & ~n4197 ;
  assign n6264 = n5135 & n6263 ;
  assign n6265 = n6264 ^ n2904 ^ 1'b0 ;
  assign n6266 = n3021 & n3213 ;
  assign n6267 = n6266 ^ n312 ^ 1'b0 ;
  assign n6268 = n1237 | n2028 ;
  assign n6269 = n6268 ^ n2739 ^ 1'b0 ;
  assign n6270 = n3211 | n6269 ;
  assign n6271 = n4446 & ~n6270 ;
  assign n6272 = ( ~n734 & n1477 ) | ( ~n734 & n1534 ) | ( n1477 & n1534 ) ;
  assign n6273 = n5449 ^ n835 ^ 1'b0 ;
  assign n6274 = n1796 ^ x11 ^ 1'b0 ;
  assign n6275 = n6274 ^ n186 ^ 1'b0 ;
  assign n6276 = n2051 & ~n4668 ;
  assign n6277 = n6276 ^ n3992 ^ 1'b0 ;
  assign n6278 = n379 & n1798 ;
  assign n6279 = n6278 ^ n3173 ^ 1'b0 ;
  assign n6280 = ( n1756 & n2300 ) | ( n1756 & n6193 ) | ( n2300 & n6193 ) ;
  assign n6281 = n107 | n3327 ;
  assign n6282 = n2922 & n6281 ;
  assign n6283 = ~n1344 & n6282 ;
  assign n6284 = n707 & ~n4519 ;
  assign n6285 = ~n2225 & n6284 ;
  assign n6286 = n6285 ^ n1816 ^ 1'b0 ;
  assign n6287 = ~n4885 & n6286 ;
  assign n6288 = n2862 ^ n2853 ^ 1'b0 ;
  assign n6289 = n6288 ^ n4849 ^ 1'b0 ;
  assign n6290 = n6289 ^ n987 ^ 1'b0 ;
  assign n6291 = n2902 & ~n2912 ;
  assign n6292 = n6291 ^ n2267 ^ 1'b0 ;
  assign n6293 = n2776 | n6292 ;
  assign n6294 = ~n753 & n887 ;
  assign n6295 = ~n1299 & n3306 ;
  assign n6296 = n6294 & n6295 ;
  assign n6297 = n3533 ^ n2267 ^ 1'b0 ;
  assign n6298 = n1422 | n6297 ;
  assign n6299 = ~n1083 & n6298 ;
  assign n6300 = ~n3157 & n6191 ;
  assign n6301 = n1582 ^ n833 ^ 1'b0 ;
  assign n6302 = n896 | n6301 ;
  assign n6303 = n3631 & ~n6302 ;
  assign n6304 = n768 & n6303 ;
  assign n6305 = ( n2197 & n2760 ) | ( n2197 & ~n6304 ) | ( n2760 & ~n6304 ) ;
  assign n6306 = n6305 ^ n2373 ^ 1'b0 ;
  assign n6307 = n4712 | n6306 ;
  assign n6308 = n1407 ^ n1040 ^ 1'b0 ;
  assign n6309 = ~n280 & n2537 ;
  assign n6310 = n1576 & ~n6309 ;
  assign n6311 = n2137 & ~n2872 ;
  assign n6312 = n135 & ~n1736 ;
  assign n6313 = n4183 | n6312 ;
  assign n6314 = n6311 & ~n6313 ;
  assign n6315 = n4100 & n5901 ;
  assign n6316 = ~n5854 & n6315 ;
  assign n6317 = n414 ^ n288 ^ 1'b0 ;
  assign n6318 = ~n3169 & n6317 ;
  assign n6319 = n2094 ^ n700 ^ 1'b0 ;
  assign n6320 = n6318 & n6319 ;
  assign n6321 = ~n1282 & n4088 ;
  assign n6322 = n1224 & ~n3155 ;
  assign n6323 = n481 | n3566 ;
  assign n6324 = n1770 & ~n6323 ;
  assign n6325 = ~n6322 & n6324 ;
  assign n6326 = ~n1724 & n4422 ;
  assign n6327 = n6326 ^ n6176 ^ 1'b0 ;
  assign n6328 = n6325 | n6327 ;
  assign n6329 = n3474 | n6328 ;
  assign n6330 = n6321 | n6329 ;
  assign n6331 = n4079 & ~n6330 ;
  assign n6332 = n6331 ^ n4515 ^ n1408 ;
  assign n6333 = n1198 | n3280 ;
  assign n6334 = n6333 ^ n421 ^ 1'b0 ;
  assign n6335 = n3776 | n6334 ;
  assign n6337 = n889 ^ n40 ^ 1'b0 ;
  assign n6336 = n774 & ~n2801 ;
  assign n6338 = n6337 ^ n6336 ^ 1'b0 ;
  assign n6339 = ~n2601 & n2929 ;
  assign n6340 = n6339 ^ n6042 ^ n21 ;
  assign n6341 = n850 | n2373 ;
  assign n6342 = n2891 & ~n6341 ;
  assign n6343 = n1407 & ~n6342 ;
  assign n6344 = n3417 | n3794 ;
  assign n6345 = ( n129 & n1691 ) | ( n129 & ~n1806 ) | ( n1691 & ~n1806 ) ;
  assign n6346 = n1843 ^ n1020 ^ 1'b0 ;
  assign n6347 = ~n6269 & n6346 ;
  assign n6348 = ( n1955 & n6345 ) | ( n1955 & n6347 ) | ( n6345 & n6347 ) ;
  assign n6349 = ~n1744 & n2365 ;
  assign n6350 = n6349 ^ n887 ^ 1'b0 ;
  assign n6353 = n2685 ^ n205 ^ 1'b0 ;
  assign n6351 = ~n3695 & n4781 ;
  assign n6352 = n6351 ^ n3634 ^ 1'b0 ;
  assign n6354 = n6353 ^ n6352 ^ n690 ;
  assign n6355 = n4231 & ~n6176 ;
  assign n6356 = n6355 ^ n5986 ^ n2600 ;
  assign n6359 = ~n767 & n2296 ;
  assign n6360 = ~n623 & n6359 ;
  assign n6361 = ~n682 & n6360 ;
  assign n6362 = n1461 & n6361 ;
  assign n6357 = ~n330 & n4912 ;
  assign n6358 = n582 & n6357 ;
  assign n6363 = n6362 ^ n6358 ^ n5586 ;
  assign n6364 = n6248 & ~n6363 ;
  assign n6365 = n5473 & n6364 ;
  assign n6366 = n615 & ~n1501 ;
  assign n6367 = n6366 ^ n4999 ^ 1'b0 ;
  assign n6368 = n5475 | n6367 ;
  assign n6369 = n5190 ^ n542 ^ 1'b0 ;
  assign n6370 = n433 | n6369 ;
  assign n6371 = ~n2789 & n6198 ;
  assign n6372 = n6371 ^ n378 ^ 1'b0 ;
  assign n6373 = n6342 ^ n6296 ^ n1184 ;
  assign n6374 = n1182 & ~n6373 ;
  assign n6375 = ~n1582 & n6374 ;
  assign n6376 = ( n3450 & ~n4741 ) | ( n3450 & n6375 ) | ( ~n4741 & n6375 ) ;
  assign n6377 = n2113 ^ n1439 ^ 1'b0 ;
  assign n6378 = ~n392 & n2967 ;
  assign n6379 = n5235 & n6378 ;
  assign n6380 = n6379 ^ n4179 ^ 1'b0 ;
  assign n6381 = n6380 ^ n4478 ^ n666 ;
  assign n6382 = n1981 ^ n191 ^ 1'b0 ;
  assign n6383 = n1582 | n6382 ;
  assign n6384 = n177 & ~n2189 ;
  assign n6385 = n6384 ^ n1385 ^ 1'b0 ;
  assign n6386 = n1929 & n6385 ;
  assign n6387 = n6386 ^ n3668 ^ 1'b0 ;
  assign n6388 = n6387 ^ n2999 ^ 1'b0 ;
  assign n6389 = n1066 & ~n6388 ;
  assign n6391 = n5246 ^ n1830 ^ 1'b0 ;
  assign n6392 = ~n1488 & n6391 ;
  assign n6390 = ~n5137 & n5768 ;
  assign n6393 = n6392 ^ n6390 ^ 1'b0 ;
  assign n6396 = n5032 ^ n1346 ^ 1'b0 ;
  assign n6394 = n1948 ^ n280 ^ 1'b0 ;
  assign n6395 = n1650 | n6394 ;
  assign n6397 = n6396 ^ n6395 ^ 1'b0 ;
  assign n6398 = n1020 & n4461 ;
  assign n6399 = n5342 ^ n1690 ^ n565 ;
  assign n6400 = n6399 ^ n2403 ^ 1'b0 ;
  assign n6401 = n4000 | n6400 ;
  assign n6402 = n6401 ^ n4866 ^ 1'b0 ;
  assign n6403 = n1262 & n6402 ;
  assign n6404 = ~n5478 & n6403 ;
  assign n6405 = ( n163 & n593 ) | ( n163 & n2040 ) | ( n593 & n2040 ) ;
  assign n6406 = n1420 | n2609 ;
  assign n6407 = n2512 ^ n2060 ^ 1'b0 ;
  assign n6408 = x7 & ~n6407 ;
  assign n6409 = n886 & ~n6408 ;
  assign n6410 = n578 & ~n6081 ;
  assign n6411 = ~n3959 & n4570 ;
  assign n6412 = n2905 & ~n6411 ;
  assign n6413 = n664 & n6412 ;
  assign n6414 = n1150 & n3105 ;
  assign n6415 = n4229 & n6414 ;
  assign n6416 = n5675 ^ n452 ^ 1'b0 ;
  assign n6417 = n6416 ^ n754 ^ 1'b0 ;
  assign n6418 = ~n694 & n3333 ;
  assign n6419 = n6418 ^ n2584 ^ 1'b0 ;
  assign n6420 = n6075 ^ n5940 ^ 1'b0 ;
  assign n6421 = n6419 & ~n6420 ;
  assign n6422 = n6421 ^ n3558 ^ 1'b0 ;
  assign n6423 = n1812 | n6422 ;
  assign n6424 = n5245 ^ n2197 ^ 1'b0 ;
  assign n6425 = n5397 ^ n2235 ^ 1'b0 ;
  assign n6426 = ~n849 & n6425 ;
  assign n6427 = n6138 ^ n620 ^ n584 ;
  assign n6428 = n6427 ^ n1558 ^ 1'b0 ;
  assign n6429 = n4228 & n6428 ;
  assign n6430 = n688 & ~n1526 ;
  assign n6431 = n5609 ^ n459 ^ 1'b0 ;
  assign n6432 = ~n4093 & n6112 ;
  assign n6433 = n6432 ^ n5760 ^ 1'b0 ;
  assign n6434 = ( ~n447 & n1832 ) | ( ~n447 & n4246 ) | ( n1832 & n4246 ) ;
  assign n6435 = n6059 ^ n2869 ^ 1'b0 ;
  assign n6436 = n3749 | n3958 ;
  assign n6437 = ( n1023 & ~n1429 ) | ( n1023 & n3181 ) | ( ~n1429 & n3181 ) ;
  assign n6438 = n6436 | n6437 ;
  assign n6439 = n6438 ^ n152 ^ 1'b0 ;
  assign n6440 = ~n31 & n3105 ;
  assign n6441 = n1571 & n6440 ;
  assign n6442 = n3429 ^ n356 ^ 1'b0 ;
  assign n6443 = n4228 ^ n1479 ^ 1'b0 ;
  assign n6444 = n3678 & ~n6443 ;
  assign n6445 = n5128 ^ n1539 ^ 1'b0 ;
  assign n6446 = n790 & n6445 ;
  assign n6447 = n6444 & n6446 ;
  assign n6448 = n1976 ^ n1408 ^ 1'b0 ;
  assign n6449 = n557 & ~n6448 ;
  assign n6450 = n6449 ^ n1798 ^ n481 ;
  assign n6451 = n1112 & ~n3209 ;
  assign n6452 = ~n6450 & n6451 ;
  assign n6453 = n2128 & n3454 ;
  assign n6454 = n6452 & n6453 ;
  assign n6455 = n4193 & ~n6181 ;
  assign n6456 = n6213 ^ n5991 ^ 1'b0 ;
  assign n6457 = n970 & n1336 ;
  assign n6458 = ( ~n1922 & n1984 ) | ( ~n1922 & n4495 ) | ( n1984 & n4495 ) ;
  assign n6459 = n575 | n1714 ;
  assign n6460 = n6459 ^ n3357 ^ 1'b0 ;
  assign n6461 = n6460 ^ n5420 ^ 1'b0 ;
  assign n6462 = n4537 & ~n6461 ;
  assign n6463 = n971 & n6462 ;
  assign n6464 = n2893 | n3236 ;
  assign n6465 = n6464 ^ n1764 ^ 1'b0 ;
  assign n6466 = n911 & n4034 ;
  assign n6467 = ~n6465 & n6466 ;
  assign n6468 = n5139 & n6467 ;
  assign n6471 = n243 | n466 ;
  assign n6472 = n108 & ~n6471 ;
  assign n6469 = n3544 ^ n2406 ^ 1'b0 ;
  assign n6470 = n81 & n6469 ;
  assign n6473 = n6472 ^ n6470 ^ 1'b0 ;
  assign n6478 = n2524 ^ n732 ^ 1'b0 ;
  assign n6479 = n1143 | n6478 ;
  assign n6480 = n1812 | n6479 ;
  assign n6481 = n6480 ^ n3123 ^ 1'b0 ;
  assign n6474 = n2442 ^ n1110 ^ 1'b0 ;
  assign n6475 = n3416 & ~n6474 ;
  assign n6476 = ~n808 & n6475 ;
  assign n6477 = n214 & ~n6476 ;
  assign n6482 = n6481 ^ n6477 ^ 1'b0 ;
  assign n6483 = n6048 ^ n265 ^ 1'b0 ;
  assign n6484 = n2583 | n4343 ;
  assign n6485 = n1803 & ~n6484 ;
  assign n6486 = n6485 ^ n2193 ^ 1'b0 ;
  assign n6487 = n2852 ^ n894 ^ 1'b0 ;
  assign n6488 = ~n1014 & n6487 ;
  assign n6489 = n3064 & ~n6488 ;
  assign n6490 = ~n1843 & n3003 ;
  assign n6491 = n1083 & n6490 ;
  assign n6492 = ~n6489 & n6491 ;
  assign n6493 = n1459 ^ n1288 ^ 1'b0 ;
  assign n6494 = n225 | n6493 ;
  assign n6495 = n4588 ^ n1933 ^ 1'b0 ;
  assign n6496 = n806 & ~n6495 ;
  assign n6497 = n425 ^ n417 ^ 1'b0 ;
  assign n6498 = n6496 & ~n6497 ;
  assign n6499 = n6498 ^ n3778 ^ 1'b0 ;
  assign n6500 = n1207 | n6499 ;
  assign n6501 = ~n6494 & n6500 ;
  assign n6502 = ~n1857 & n6501 ;
  assign n6503 = n2779 | n6502 ;
  assign n6504 = n4416 | n6503 ;
  assign n6505 = n3271 ^ n2770 ^ 1'b0 ;
  assign n6506 = n1497 & n6505 ;
  assign n6507 = n6506 ^ n4754 ^ 1'b0 ;
  assign n6508 = ~n1755 & n5063 ;
  assign n6509 = n6508 ^ n4155 ^ 1'b0 ;
  assign n6510 = n3285 & n5809 ;
  assign n6511 = n6510 ^ n2275 ^ 1'b0 ;
  assign n6517 = n5031 ^ n1072 ^ 1'b0 ;
  assign n6518 = n2217 | n6517 ;
  assign n6519 = n2539 ^ n368 ^ 1'b0 ;
  assign n6520 = n812 & n6519 ;
  assign n6521 = n6520 ^ n1063 ^ 1'b0 ;
  assign n6522 = ~n6518 & n6521 ;
  assign n6512 = n2443 ^ n508 ^ 1'b0 ;
  assign n6513 = ~n1655 & n2760 ;
  assign n6514 = n6513 ^ n21 ^ 1'b0 ;
  assign n6515 = n6512 & ~n6514 ;
  assign n6516 = ~n503 & n6515 ;
  assign n6523 = n6522 ^ n6516 ^ 1'b0 ;
  assign n6524 = n2541 | n5759 ;
  assign n6525 = ( n619 & ~n3435 ) | ( n619 & n6264 ) | ( ~n3435 & n6264 ) ;
  assign n6526 = ( n130 & n950 ) | ( n130 & n2481 ) | ( n950 & n2481 ) ;
  assign n6527 = ( n112 & n280 ) | ( n112 & n6526 ) | ( n280 & n6526 ) ;
  assign n6528 = n1049 | n6527 ;
  assign n6529 = ~n6525 & n6528 ;
  assign n6530 = n6529 ^ n1684 ^ 1'b0 ;
  assign n6532 = n237 & ~n2478 ;
  assign n6533 = ~n5096 & n6532 ;
  assign n6531 = n3367 & ~n4082 ;
  assign n6534 = n6533 ^ n6531 ^ 1'b0 ;
  assign n6535 = n5841 & ~n6534 ;
  assign n6536 = ~n3193 & n6359 ;
  assign n6537 = ~n6535 & n6536 ;
  assign n6538 = ~n4328 & n5417 ;
  assign n6539 = n48 & ~n5680 ;
  assign n6540 = ( n6262 & n6538 ) | ( n6262 & ~n6539 ) | ( n6538 & ~n6539 ) ;
  assign n6541 = n2226 | n5330 ;
  assign n6542 = n6541 ^ n1306 ^ 1'b0 ;
  assign n6543 = n6542 ^ n1743 ^ 1'b0 ;
  assign n6547 = ~n124 & n2508 ;
  assign n6548 = ~n1221 & n6547 ;
  assign n6549 = n6548 ^ n2112 ^ 1'b0 ;
  assign n6550 = ~n563 & n6549 ;
  assign n6545 = n752 & n2365 ;
  assign n6546 = ~n5551 & n6545 ;
  assign n6551 = n6550 ^ n6546 ^ 1'b0 ;
  assign n6544 = n1876 & n3261 ;
  assign n6552 = n6551 ^ n6544 ^ 1'b0 ;
  assign n6553 = n6543 & n6552 ;
  assign n6554 = n2904 | n4776 ;
  assign n6555 = n465 | n6554 ;
  assign n6556 = n6555 ^ n676 ^ 1'b0 ;
  assign n6557 = ( n2404 & n2891 ) | ( n2404 & n6556 ) | ( n2891 & n6556 ) ;
  assign n6558 = n4020 ^ n2066 ^ 1'b0 ;
  assign n6559 = n2807 & ~n6558 ;
  assign n6560 = x3 | n1562 ;
  assign n6561 = n698 | n1167 ;
  assign n6562 = n6560 | n6561 ;
  assign n6563 = ~n1488 & n6562 ;
  assign n6564 = n4267 & ~n6563 ;
  assign n6565 = n6559 & ~n6564 ;
  assign n6566 = ~n2550 & n6565 ;
  assign n6568 = n45 & ~n770 ;
  assign n6567 = ~n3609 & n4685 ;
  assign n6569 = n6568 ^ n6567 ^ 1'b0 ;
  assign n6570 = ( n277 & n4481 ) | ( n277 & n6569 ) | ( n4481 & n6569 ) ;
  assign n6571 = n4775 ^ n182 ^ 1'b0 ;
  assign n6572 = n1551 & n6571 ;
  assign n6573 = n6033 & ~n6217 ;
  assign n6574 = n3835 | n3927 ;
  assign n6575 = ~n1973 & n3867 ;
  assign n6576 = n6575 ^ n3788 ^ n1488 ;
  assign n6577 = ~n148 & n2236 ;
  assign n6578 = ~n1234 & n6577 ;
  assign n6579 = n4698 | n4824 ;
  assign n6580 = n6578 & ~n6579 ;
  assign n6581 = n1426 & n2033 ;
  assign n6582 = ~n1411 & n1811 ;
  assign n6583 = n6582 ^ n3539 ^ 1'b0 ;
  assign n6584 = n6583 ^ n4698 ^ 1'b0 ;
  assign n6585 = n6584 ^ n2927 ^ n1868 ;
  assign n6586 = n200 | n4429 ;
  assign n6587 = n3519 ^ n1588 ^ 1'b0 ;
  assign n6588 = n6586 | n6587 ;
  assign n6594 = n3556 ^ n1872 ^ 1'b0 ;
  assign n6589 = n5111 ^ n205 ^ 1'b0 ;
  assign n6590 = ~n2030 & n6589 ;
  assign n6591 = n6590 ^ n323 ^ 1'b0 ;
  assign n6592 = ~n3966 & n6591 ;
  assign n6593 = n4813 & n6592 ;
  assign n6595 = n6594 ^ n6593 ^ 1'b0 ;
  assign n6596 = n3723 & ~n4672 ;
  assign n6597 = n3646 & n4622 ;
  assign n6598 = n6597 ^ n2598 ^ 1'b0 ;
  assign n6599 = n6596 | n6598 ;
  assign n6600 = n3070 ^ n1298 ^ 1'b0 ;
  assign n6601 = n6600 ^ n2907 ^ 1'b0 ;
  assign n6602 = n1770 & n6228 ;
  assign n6603 = n2137 ^ n2080 ^ 1'b0 ;
  assign n6604 = n6602 & n6603 ;
  assign n6605 = ( n1657 & n3508 ) | ( n1657 & n4607 ) | ( n3508 & n4607 ) ;
  assign n6606 = n253 & n1298 ;
  assign n6607 = n6606 ^ n2078 ^ 1'b0 ;
  assign n6608 = n6607 ^ n2828 ^ n105 ;
  assign n6609 = n774 | n985 ;
  assign n6610 = n6609 ^ n2048 ^ 1'b0 ;
  assign n6611 = n488 & n2641 ;
  assign n6612 = n6611 ^ n2347 ^ 1'b0 ;
  assign n6613 = n2192 & n6612 ;
  assign n6614 = n2104 & n5392 ;
  assign n6615 = ~n549 & n6614 ;
  assign n6616 = n6615 ^ n1741 ^ 1'b0 ;
  assign n6617 = n1306 | n1745 ;
  assign n6618 = n4103 ^ n3162 ^ 1'b0 ;
  assign n6619 = n3418 & n6618 ;
  assign n6620 = n975 | n1152 ;
  assign n6621 = n3198 & n6620 ;
  assign n6624 = n914 & n1350 ;
  assign n6625 = ~n2614 & n6624 ;
  assign n6622 = n1212 ^ n652 ^ 1'b0 ;
  assign n6623 = n6622 ^ n5758 ^ 1'b0 ;
  assign n6626 = n6625 ^ n6623 ^ 1'b0 ;
  assign n6627 = n4710 ^ n362 ^ 1'b0 ;
  assign n6628 = n6626 & ~n6627 ;
  assign n6629 = ( n3466 & n5454 ) | ( n3466 & n6035 ) | ( n5454 & n6035 ) ;
  assign n6630 = n6629 ^ n6570 ^ 1'b0 ;
  assign n6631 = n4218 | n6409 ;
  assign n6632 = n5079 ^ n4109 ^ 1'b0 ;
  assign n6633 = n6385 ^ n6154 ^ 1'b0 ;
  assign n6634 = n2442 ^ n2086 ^ 1'b0 ;
  assign n6635 = n1543 & n6634 ;
  assign n6636 = n6201 & n6576 ;
  assign n6637 = ~n6635 & n6636 ;
  assign n6638 = n850 | n6637 ;
  assign n6639 = n4148 & n5562 ;
  assign n6640 = n1837 & n6639 ;
  assign n6641 = ( ~n2038 & n4653 ) | ( ~n2038 & n6640 ) | ( n4653 & n6640 ) ;
  assign n6642 = n5929 ^ n1533 ^ 1'b0 ;
  assign n6643 = ~n4814 & n6642 ;
  assign n6644 = n2851 & ~n3715 ;
  assign n6645 = n6644 ^ n6481 ^ 1'b0 ;
  assign n6646 = n1124 | n2769 ;
  assign n6647 = n1211 & ~n2258 ;
  assign n6648 = n3276 & ~n6647 ;
  assign n6649 = n6648 ^ n2481 ^ 1'b0 ;
  assign n6650 = n4328 & n6649 ;
  assign n6651 = ~n1461 & n5321 ;
  assign n6652 = n4224 | n6651 ;
  assign n6653 = n6652 ^ n1644 ^ 1'b0 ;
  assign n6654 = n1700 | n1896 ;
  assign n6655 = n6654 ^ n3165 ^ 1'b0 ;
  assign n6656 = n1732 & n6655 ;
  assign n6657 = n5967 ^ n5699 ^ n2068 ;
  assign n6658 = ~n1933 & n2212 ;
  assign n6659 = n1300 & n6658 ;
  assign n6660 = n6659 ^ n806 ^ 1'b0 ;
  assign n6661 = n130 & ~n6660 ;
  assign n6662 = n4515 & n6661 ;
  assign n6663 = n3633 ^ n1534 ^ 1'b0 ;
  assign n6664 = n6663 ^ n5219 ^ 1'b0 ;
  assign n6665 = n6664 ^ n915 ^ 1'b0 ;
  assign n6666 = n5599 ^ n1065 ^ 1'b0 ;
  assign n6667 = n3971 & ~n6666 ;
  assign n6668 = n20 & ~n4395 ;
  assign n6669 = n6668 ^ n2852 ^ 1'b0 ;
  assign n6670 = n5294 & n5624 ;
  assign n6671 = n828 & ~n2761 ;
  assign n6672 = n1244 ^ n668 ^ n219 ;
  assign n6673 = n5059 ^ n2661 ^ 1'b0 ;
  assign n6674 = n6672 | n6673 ;
  assign n6675 = ( ~n1338 & n6671 ) | ( ~n1338 & n6674 ) | ( n6671 & n6674 ) ;
  assign n6676 = n301 | n3783 ;
  assign n6677 = n6676 ^ n5610 ^ 1'b0 ;
  assign n6678 = n2771 | n6677 ;
  assign n6679 = ~n481 & n3621 ;
  assign n6680 = ~n3998 & n6679 ;
  assign n6681 = n3766 ^ n1488 ^ 1'b0 ;
  assign n6682 = n1098 & n3631 ;
  assign n6683 = ~n489 & n6682 ;
  assign n6684 = n831 | n1049 ;
  assign n6685 = n6684 ^ n4061 ^ 1'b0 ;
  assign n6686 = n446 & n1285 ;
  assign n6687 = n6686 ^ n1235 ^ 1'b0 ;
  assign n6688 = ~n1093 & n3946 ;
  assign n6689 = n104 | n6688 ;
  assign n6690 = n2065 | n6689 ;
  assign n6691 = n2669 & n5432 ;
  assign n6692 = ~n6690 & n6691 ;
  assign n6693 = n5809 ^ n1624 ^ 1'b0 ;
  assign n6694 = n2356 | n6693 ;
  assign n6695 = ~n6581 & n6694 ;
  assign n6696 = ~n574 & n800 ;
  assign n6697 = n5132 | n6696 ;
  assign n6698 = ~n1517 & n2288 ;
  assign n6699 = ~n6522 & n6698 ;
  assign n6700 = n4135 | n5179 ;
  assign n6701 = n5293 ^ n2881 ^ n877 ;
  assign n6702 = n207 | n6701 ;
  assign n6703 = n842 | n1031 ;
  assign n6704 = n6703 ^ n4459 ^ 1'b0 ;
  assign n6705 = n2933 ^ n1843 ^ 1'b0 ;
  assign n6706 = n6705 ^ n600 ^ 1'b0 ;
  assign n6707 = n1495 & n6706 ;
  assign n6708 = n813 & n3319 ;
  assign n6709 = n6708 ^ n533 ^ 1'b0 ;
  assign n6710 = n6709 ^ n5113 ^ 1'b0 ;
  assign n6711 = n521 & ~n6710 ;
  assign n6712 = n6711 ^ n533 ^ 1'b0 ;
  assign n6713 = n3886 ^ n2480 ^ n717 ;
  assign n6714 = n3484 ^ n1152 ^ 1'b0 ;
  assign n6715 = n6714 ^ n3095 ^ 1'b0 ;
  assign n6716 = n2813 & ~n6715 ;
  assign n6717 = n4762 ^ n1038 ^ 1'b0 ;
  assign n6718 = n6701 ^ n2773 ^ 1'b0 ;
  assign n6719 = ~n466 & n2915 ;
  assign n6720 = n6718 & ~n6719 ;
  assign n6721 = n635 & ~n988 ;
  assign n6722 = n2031 & n6721 ;
  assign n6723 = n6722 ^ n1313 ^ n927 ;
  assign n6724 = n2306 & ~n5190 ;
  assign n6725 = n6723 & n6724 ;
  assign n6726 = n4881 & ~n6725 ;
  assign n6728 = n368 | n442 ;
  assign n6729 = n2056 & ~n6728 ;
  assign n6727 = n5616 ^ n3854 ^ n1718 ;
  assign n6730 = n6729 ^ n6727 ^ n3488 ;
  assign n6731 = n5872 & ~n6730 ;
  assign n6732 = n1800 & n6255 ;
  assign n6733 = ~n773 & n5725 ;
  assign n6734 = n6733 ^ n2698 ^ 1'b0 ;
  assign n6735 = n5377 | n6734 ;
  assign n6736 = n755 & ~n6735 ;
  assign n6737 = n4091 ^ n3270 ^ 1'b0 ;
  assign n6738 = ~n3078 & n6737 ;
  assign n6741 = n1647 & ~n6245 ;
  assign n6739 = n4868 ^ n3734 ^ 1'b0 ;
  assign n6740 = n3876 & ~n6739 ;
  assign n6742 = n6741 ^ n6740 ^ 1'b0 ;
  assign n6743 = n3257 ^ n296 ^ 1'b0 ;
  assign n6744 = ( n4163 & n5250 ) | ( n4163 & ~n6743 ) | ( n5250 & ~n6743 ) ;
  assign n6745 = n2802 | n5954 ;
  assign n6746 = n700 | n6745 ;
  assign n6747 = n6744 & ~n6746 ;
  assign n6748 = n578 | n2635 ;
  assign n6749 = n6748 ^ n6352 ^ n4179 ;
  assign n6750 = n115 & n1327 ;
  assign n6751 = n3703 ^ n3399 ^ 1'b0 ;
  assign n6753 = n6743 ^ n6099 ^ 1'b0 ;
  assign n6752 = n1521 | n3993 ;
  assign n6754 = n6753 ^ n6752 ^ 1'b0 ;
  assign n6755 = n1654 ^ n1152 ^ 1'b0 ;
  assign n6756 = n340 & n6755 ;
  assign n6757 = n6756 ^ n3169 ^ n2328 ;
  assign n6758 = ~n1981 & n6757 ;
  assign n6759 = n6758 ^ n3514 ^ 1'b0 ;
  assign n6760 = n768 | n1159 ;
  assign n6761 = n13 | n3759 ;
  assign n6762 = n3564 ^ n3258 ^ 1'b0 ;
  assign n6763 = n200 & n6762 ;
  assign n6764 = ~n1159 & n5350 ;
  assign n6765 = n1771 & ~n3327 ;
  assign n6766 = n1251 ^ n1024 ^ n535 ;
  assign n6767 = n213 | n342 ;
  assign n6768 = n6767 ^ n1293 ^ 1'b0 ;
  assign n6769 = ~n5490 & n6768 ;
  assign n6770 = n3031 & n6057 ;
  assign n6773 = ( ~n2314 & n4063 ) | ( ~n2314 & n4505 ) | ( n4063 & n4505 ) ;
  assign n6771 = n1848 ^ n158 ^ 1'b0 ;
  assign n6772 = n2252 | n6771 ;
  assign n6774 = n6773 ^ n6772 ^ 1'b0 ;
  assign n6775 = n83 & n358 ;
  assign n6776 = n1789 | n5058 ;
  assign n6777 = ( n2989 & ~n3434 ) | ( n2989 & n6776 ) | ( ~n3434 & n6776 ) ;
  assign n6778 = n1469 | n1652 ;
  assign n6779 = n6778 ^ n2708 ^ 1'b0 ;
  assign n6780 = n378 & ~n654 ;
  assign n6781 = n320 & ~n5202 ;
  assign n6782 = ~n2367 & n6781 ;
  assign n6783 = n6782 ^ n1207 ^ 1'b0 ;
  assign n6784 = n5353 & n6783 ;
  assign n6785 = ( ~n477 & n731 ) | ( ~n477 & n6784 ) | ( n731 & n6784 ) ;
  assign n6786 = n279 & n2014 ;
  assign n6787 = n6786 ^ n1528 ^ 1'b0 ;
  assign n6788 = n2199 & ~n4381 ;
  assign n6789 = n5827 & n6788 ;
  assign n6793 = ~n667 & n4677 ;
  assign n6794 = n3760 & n6793 ;
  assign n6790 = n216 & ~n1962 ;
  assign n6791 = n6790 ^ n6048 ^ 1'b0 ;
  assign n6792 = ~n2236 & n6791 ;
  assign n6795 = n6794 ^ n6792 ^ 1'b0 ;
  assign n6796 = n6789 | n6795 ;
  assign n6797 = n6796 ^ n1765 ^ n162 ;
  assign n6798 = n406 & ~n2705 ;
  assign n6799 = ~n5464 & n6798 ;
  assign n6800 = n2417 ^ n1146 ^ 1'b0 ;
  assign n6801 = n1141 & n3588 ;
  assign n6802 = n4278 & n6801 ;
  assign n6803 = n6800 & ~n6802 ;
  assign n6804 = n6799 & n6803 ;
  assign n6805 = n3044 ^ n2778 ^ n56 ;
  assign n6806 = n6172 | n6805 ;
  assign n6807 = n5174 ^ n1528 ^ 1'b0 ;
  assign n6808 = n6806 | n6807 ;
  assign n6809 = n3345 & ~n6808 ;
  assign n6810 = n1657 | n3895 ;
  assign n6811 = n1994 & ~n6810 ;
  assign n6812 = n6811 ^ n5001 ^ 1'b0 ;
  assign n6813 = n952 | n6812 ;
  assign n6814 = n5042 | n6813 ;
  assign n6815 = ( n4591 & n5362 ) | ( n4591 & n5546 ) | ( n5362 & n5546 ) ;
  assign n6816 = n1165 & ~n6294 ;
  assign n6817 = ~n5497 & n6816 ;
  assign n6818 = n6817 ^ n2754 ^ n2619 ;
  assign n6819 = n2340 ^ n652 ^ 1'b0 ;
  assign n6820 = n4381 | n6819 ;
  assign n6821 = n2706 & ~n6554 ;
  assign n6822 = n6821 ^ n4289 ^ 1'b0 ;
  assign n6823 = n6820 | n6822 ;
  assign n6824 = n6823 ^ n2314 ^ n737 ;
  assign n6825 = n4248 ^ n189 ^ 1'b0 ;
  assign n6826 = n4473 ^ n620 ^ 1'b0 ;
  assign n6827 = n4702 & n6826 ;
  assign n6828 = ~n1922 & n2225 ;
  assign n6829 = ~n6827 & n6828 ;
  assign n6830 = n226 & n4182 ;
  assign n6831 = n1837 & n6830 ;
  assign n6832 = n6831 ^ n4127 ^ 1'b0 ;
  assign n6833 = n6729 ^ n4203 ^ 1'b0 ;
  assign n6834 = n352 | n1038 ;
  assign n6835 = n6834 ^ n192 ^ 1'b0 ;
  assign n6836 = n5632 | n6835 ;
  assign n6837 = n4422 ^ n484 ^ 1'b0 ;
  assign n6838 = n1843 | n6837 ;
  assign n6839 = n320 & n6838 ;
  assign n6840 = ~n5637 & n5807 ;
  assign n6841 = ~n6839 & n6840 ;
  assign n6842 = n1005 & n6318 ;
  assign n6843 = ~n3173 & n6842 ;
  assign n6844 = ~n1877 & n6843 ;
  assign n6845 = n3516 ^ n211 ^ 1'b0 ;
  assign n6846 = n4946 | n6845 ;
  assign n6847 = n6846 ^ n2282 ^ 1'b0 ;
  assign n6848 = n3680 & n5437 ;
  assign n6849 = ~n6667 & n6848 ;
  assign n6850 = n6092 & ~n6849 ;
  assign n6851 = n3477 ^ n3319 ^ 1'b0 ;
  assign n6852 = n5824 | n6632 ;
  assign n6854 = n363 | n1286 ;
  assign n6853 = n2098 & n6149 ;
  assign n6855 = n6854 ^ n6853 ^ 1'b0 ;
  assign n6856 = n124 & ~n2332 ;
  assign n6857 = n1893 ^ n226 ^ 1'b0 ;
  assign n6858 = n2675 ^ n2664 ^ n645 ;
  assign n6859 = n6857 | n6858 ;
  assign n6860 = n6856 | n6859 ;
  assign n6861 = n2051 & ~n4222 ;
  assign n6862 = ~n4005 & n6861 ;
  assign n6863 = ~n6860 & n6862 ;
  assign n6864 = ~n1578 & n1768 ;
  assign n6865 = n244 & n855 ;
  assign n6866 = n6865 ^ n2512 ^ 1'b0 ;
  assign n6867 = ~n5989 & n6866 ;
  assign n6868 = ( n2155 & n6864 ) | ( n2155 & n6867 ) | ( n6864 & n6867 ) ;
  assign n6869 = n335 & n6868 ;
  assign n6870 = n1731 ^ n1025 ^ 1'b0 ;
  assign n6871 = n6870 ^ n2146 ^ n334 ;
  assign n6872 = n1701 & ~n6871 ;
  assign n6873 = n698 | n6872 ;
  assign n6874 = n6873 ^ n770 ^ 1'b0 ;
  assign n6875 = n5909 ^ n1385 ^ 1'b0 ;
  assign n6876 = n1811 & ~n6875 ;
  assign n6877 = n688 & ~n2240 ;
  assign n6878 = n140 & n6877 ;
  assign n6879 = n4609 ^ n2724 ^ 1'b0 ;
  assign n6880 = ~n1774 & n6879 ;
  assign n6881 = ~n829 & n2614 ;
  assign n6882 = x11 & ~n6881 ;
  assign n6883 = ~n1130 & n6882 ;
  assign n6884 = n1469 & ~n6883 ;
  assign n6885 = ~n6880 & n6884 ;
  assign n6886 = n515 & ~n6885 ;
  assign n6887 = n4214 ^ n2726 ^ 1'b0 ;
  assign n6888 = n2673 | n6887 ;
  assign n6889 = ( n1861 & n4761 ) | ( n1861 & ~n6888 ) | ( n4761 & ~n6888 ) ;
  assign n6890 = n6889 ^ n6128 ^ 1'b0 ;
  assign n6891 = n1321 | n2604 ;
  assign n6892 = n4551 & n5977 ;
  assign n6893 = n4683 ^ n4662 ^ n3592 ;
  assign n6894 = ( ~n1648 & n2541 ) | ( ~n1648 & n6893 ) | ( n2541 & n6893 ) ;
  assign n6895 = n1063 & n6894 ;
  assign n6896 = n6892 | n6895 ;
  assign n6897 = n1636 & n1731 ;
  assign n6898 = n3185 & n6897 ;
  assign n6899 = n4850 & n6709 ;
  assign n6900 = ~n5507 & n6899 ;
  assign n6901 = n5693 & n6900 ;
  assign n6902 = n3524 ^ n2352 ^ 1'b0 ;
  assign n6904 = ( n1143 & ~n1398 ) | ( n1143 & n3437 ) | ( ~n1398 & n3437 ) ;
  assign n6903 = n1063 ^ n107 ^ 1'b0 ;
  assign n6905 = n6904 ^ n6903 ^ 1'b0 ;
  assign n6906 = n6016 & ~n6905 ;
  assign n6907 = n1173 ^ n224 ^ 1'b0 ;
  assign n6908 = n5839 ^ n4187 ^ 1'b0 ;
  assign n6909 = n6908 ^ n6695 ^ 1'b0 ;
  assign n6910 = n5052 & n6909 ;
  assign n6911 = n4813 & n6876 ;
  assign n6913 = n43 & n3098 ;
  assign n6914 = n6913 ^ n35 ^ 1'b0 ;
  assign n6912 = n3403 & ~n4026 ;
  assign n6915 = n6914 ^ n6912 ^ 1'b0 ;
  assign n6916 = ~n6758 & n6915 ;
  assign n6917 = n6916 ^ n2202 ^ 1'b0 ;
  assign n6918 = n6917 ^ n6274 ^ 1'b0 ;
  assign n6919 = n1109 | n6918 ;
  assign n6921 = n1497 & n3537 ;
  assign n6922 = ~n194 & n6921 ;
  assign n6923 = n4302 & ~n6922 ;
  assign n6920 = n1000 & ~n6302 ;
  assign n6924 = n6923 ^ n6920 ^ 1'b0 ;
  assign n6925 = n1946 & n4707 ;
  assign n6926 = n4698 | n6106 ;
  assign n6927 = n607 ^ n477 ^ 1'b0 ;
  assign n6928 = n6041 | n6927 ;
  assign n6929 = n3101 ^ n2925 ^ 1'b0 ;
  assign n6930 = n6043 | n6929 ;
  assign n6931 = n978 & ~n1347 ;
  assign n6932 = n4082 | n6931 ;
  assign n6933 = n6932 ^ n1308 ^ 1'b0 ;
  assign n6934 = n6933 ^ n5839 ^ 1'b0 ;
  assign n6935 = n6934 ^ n5791 ^ n3518 ;
  assign n6936 = ~n1267 & n2808 ;
  assign n6937 = n6936 ^ n1219 ^ 1'b0 ;
  assign n6938 = n3412 ^ n706 ^ 1'b0 ;
  assign n6939 = n6937 | n6938 ;
  assign n6940 = n2087 ^ n67 ^ 1'b0 ;
  assign n6941 = n2639 ^ n432 ^ 1'b0 ;
  assign n6942 = n4710 & n5022 ;
  assign n6943 = n3904 ^ n996 ^ 1'b0 ;
  assign n6944 = ( ~n2637 & n5266 ) | ( ~n2637 & n5629 ) | ( n5266 & n5629 ) ;
  assign n6945 = n5982 ^ n2460 ^ 1'b0 ;
  assign n6946 = n2588 ^ n1065 ^ 1'b0 ;
  assign n6947 = n3892 ^ n2521 ^ 1'b0 ;
  assign n6948 = n2679 | n6947 ;
  assign n6949 = n2978 ^ n2708 ^ 1'b0 ;
  assign n6950 = n194 & ~n3972 ;
  assign n6951 = n1964 ^ n83 ^ 1'b0 ;
  assign n6953 = n1693 & ~n4173 ;
  assign n6952 = n1215 & n2146 ;
  assign n6954 = n6953 ^ n6952 ^ 1'b0 ;
  assign n6955 = n456 | n6954 ;
  assign n6956 = n681 & ~n1224 ;
  assign n6957 = n110 & n6956 ;
  assign n6958 = n4066 & ~n6957 ;
  assign n6959 = n6256 & n6958 ;
  assign n6960 = n253 & ~n3095 ;
  assign n6961 = n6960 ^ n4535 ^ 1'b0 ;
  assign n6962 = n694 & n6961 ;
  assign n6963 = n6962 ^ n200 ^ 1'b0 ;
  assign n6964 = n5431 ^ n2697 ^ n582 ;
  assign n6965 = n963 & n6406 ;
  assign n6966 = n5093 & n6965 ;
  assign n6967 = n1374 & n6880 ;
  assign n6968 = n4321 & n6967 ;
  assign n6969 = n6968 ^ n428 ^ 1'b0 ;
  assign n6970 = n4543 | n6969 ;
  assign n6971 = n609 & ~n6970 ;
  assign n6972 = n6971 ^ n4300 ^ 1'b0 ;
  assign n6974 = ~n663 & n3700 ;
  assign n6975 = n6974 ^ n924 ^ 1'b0 ;
  assign n6973 = n3562 & n6344 ;
  assign n6976 = n6975 ^ n6973 ^ 1'b0 ;
  assign n6977 = n1563 | n3710 ;
  assign n6978 = n6976 | n6977 ;
  assign n6979 = n2223 | n2600 ;
  assign n6980 = n489 | n938 ;
  assign n6981 = ~n6979 & n6980 ;
  assign n6982 = n6198 ^ n1451 ^ 1'b0 ;
  assign n6983 = ~n453 & n3012 ;
  assign n6984 = n4795 & n6983 ;
  assign n6985 = n6984 ^ n6629 ^ 1'b0 ;
  assign n6986 = n5201 ^ n4980 ^ n3826 ;
  assign n6987 = n983 | n3358 ;
  assign n6988 = n6987 ^ n135 ^ 1'b0 ;
  assign n6989 = n6988 ^ n6878 ^ 1'b0 ;
  assign n6990 = n902 & n2273 ;
  assign n6991 = n1260 ^ n907 ^ 1'b0 ;
  assign n6992 = n2455 ^ n2291 ^ 1'b0 ;
  assign n6993 = n1601 & ~n6992 ;
  assign n6994 = n6993 ^ n4999 ^ 1'b0 ;
  assign n6995 = ( n3409 & n6991 ) | ( n3409 & n6994 ) | ( n6991 & n6994 ) ;
  assign n6996 = n4555 & n6995 ;
  assign n6997 = ~n459 & n541 ;
  assign n6998 = ~n297 & n867 ;
  assign n6999 = ~n6997 & n6998 ;
  assign n7000 = n2862 & n3586 ;
  assign n7001 = n2472 & ~n7000 ;
  assign n7002 = n2905 & ~n7001 ;
  assign n7003 = n6704 & n7002 ;
  assign n7008 = n840 ^ n179 ^ 1'b0 ;
  assign n7004 = n2303 ^ n314 ^ 1'b0 ;
  assign n7005 = ~n69 & n7004 ;
  assign n7006 = n1647 | n7005 ;
  assign n7007 = n1136 & ~n7006 ;
  assign n7009 = n7008 ^ n7007 ^ 1'b0 ;
  assign n7010 = n6871 & n7009 ;
  assign n7011 = n5130 ^ n1867 ^ n1422 ;
  assign n7012 = n1955 & ~n7011 ;
  assign n7019 = n1740 ^ n1473 ^ n182 ;
  assign n7016 = n3867 ^ n2363 ^ n325 ;
  assign n7013 = ~n1898 & n4986 ;
  assign n7014 = n458 & n7013 ;
  assign n7015 = n7014 ^ n3129 ^ 1'b0 ;
  assign n7017 = n7016 ^ n7015 ^ 1'b0 ;
  assign n7018 = n4504 & ~n7017 ;
  assign n7020 = n7019 ^ n7018 ^ 1'b0 ;
  assign n7021 = n5719 ^ n5107 ^ 1'b0 ;
  assign n7022 = ~n6796 & n7021 ;
  assign n7023 = n3372 & ~n5699 ;
  assign n7024 = n371 & ~n620 ;
  assign n7025 = n5976 & n7024 ;
  assign n7026 = n388 ^ n149 ^ 1'b0 ;
  assign n7027 = n7025 & ~n7026 ;
  assign n7028 = ~n4937 & n7027 ;
  assign n7029 = ~n344 & n7028 ;
  assign n7030 = n4555 ^ n1289 ^ 1'b0 ;
  assign n7031 = n4405 & ~n5612 ;
  assign n7032 = ~n3934 & n7031 ;
  assign n7033 = n1772 & n7032 ;
  assign n7034 = n1896 | n7033 ;
  assign n7035 = n1050 & n4416 ;
  assign n7036 = n7035 ^ n3758 ^ 1'b0 ;
  assign n7037 = n3080 | n4550 ;
  assign n7038 = n7037 ^ n5682 ^ 1'b0 ;
  assign n7039 = n3461 & n3639 ;
  assign n7040 = n7039 ^ n6870 ^ 1'b0 ;
  assign n7041 = ~n948 & n7040 ;
  assign n7044 = n3177 ^ n2262 ^ 1'b0 ;
  assign n7045 = ( ~n1576 & n2175 ) | ( ~n1576 & n7044 ) | ( n2175 & n7044 ) ;
  assign n7042 = n1243 ^ n56 ^ 1'b0 ;
  assign n7043 = n414 | n7042 ;
  assign n7046 = n7045 ^ n7043 ^ 1'b0 ;
  assign n7047 = ( ~n4814 & n5266 ) | ( ~n4814 & n7046 ) | ( n5266 & n7046 ) ;
  assign n7048 = n362 | n2150 ;
  assign n7049 = n2273 | n5317 ;
  assign n7050 = n7049 ^ n1235 ^ 1'b0 ;
  assign n7051 = n5594 ^ n3058 ^ n2883 ;
  assign n7052 = ( ~n2223 & n7050 ) | ( ~n2223 & n7051 ) | ( n7050 & n7051 ) ;
  assign n7053 = ( n1558 & n7048 ) | ( n1558 & n7052 ) | ( n7048 & n7052 ) ;
  assign n7054 = n1620 ^ n1618 ^ 1'b0 ;
  assign n7055 = n7054 ^ n1363 ^ 1'b0 ;
  assign n7056 = ~n1935 & n7055 ;
  assign n7057 = n112 & n7056 ;
  assign n7058 = n7057 ^ n1484 ^ 1'b0 ;
  assign n7059 = n83 & n3924 ;
  assign n7060 = n7059 ^ n4510 ^ n3633 ;
  assign n7061 = n7058 & n7060 ;
  assign n7062 = n1021 & n2387 ;
  assign n7063 = n2109 & ~n7062 ;
  assign n7065 = n2845 & ~n3695 ;
  assign n7066 = n1413 & n7065 ;
  assign n7064 = n1465 | n2576 ;
  assign n7067 = n7066 ^ n7064 ^ 1'b0 ;
  assign n7068 = n1336 & ~n2881 ;
  assign n7069 = n7068 ^ n378 ^ 1'b0 ;
  assign n7070 = ~n5660 & n7069 ;
  assign n7071 = n1865 & n7070 ;
  assign n7072 = n7071 ^ n4583 ^ 1'b0 ;
  assign n7073 = ~n7067 & n7072 ;
  assign n7074 = n2922 & ~n4088 ;
  assign n7075 = n1674 & n7074 ;
  assign n7076 = n5449 & n7075 ;
  assign n7077 = n316 & n3143 ;
  assign n7078 = ~n233 & n7077 ;
  assign n7079 = ~n1252 & n6667 ;
  assign n7080 = n5828 ^ n5023 ^ 1'b0 ;
  assign n7081 = n6827 & n7061 ;
  assign n7082 = n3415 & n3566 ;
  assign n7083 = ~n3779 & n7082 ;
  assign n7084 = ~n3992 & n7083 ;
  assign n7085 = n2377 ^ n2306 ^ 1'b0 ;
  assign n7086 = ~n7046 & n7085 ;
  assign n7087 = n2448 ^ n36 ^ 1'b0 ;
  assign n7088 = n7087 ^ n1143 ^ 1'b0 ;
  assign n7089 = n2865 | n3226 ;
  assign n7092 = n3980 ^ n2080 ^ 1'b0 ;
  assign n7090 = n2569 & ~n5667 ;
  assign n7091 = n7090 ^ n3940 ^ 1'b0 ;
  assign n7093 = n7092 ^ n7091 ^ 1'b0 ;
  assign n7094 = n5142 | n5504 ;
  assign n7095 = n7094 ^ n5949 ^ 1'b0 ;
  assign n7097 = n2000 ^ n311 ^ 1'b0 ;
  assign n7098 = n7097 ^ n4610 ^ 1'b0 ;
  assign n7099 = ~n654 & n7098 ;
  assign n7100 = n2079 & ~n7099 ;
  assign n7096 = n5433 ^ n3696 ^ n1525 ;
  assign n7101 = n7100 ^ n7096 ^ 1'b0 ;
  assign n7102 = n3017 | n7101 ;
  assign n7103 = n7102 ^ n5095 ^ 1'b0 ;
  assign n7104 = n6054 & n7103 ;
  assign n7105 = n205 | n3097 ;
  assign n7106 = n7105 ^ n835 ^ 1'b0 ;
  assign n7107 = ~n541 & n5968 ;
  assign n7108 = ~n560 & n1732 ;
  assign n7109 = n58 & n5787 ;
  assign n7110 = n4189 | n7109 ;
  assign n7111 = n1617 & n5004 ;
  assign n7112 = n1968 ^ n1826 ^ 1'b0 ;
  assign n7113 = n7112 ^ n6594 ^ 1'b0 ;
  assign n7114 = n1130 & ~n7113 ;
  assign n7115 = n7114 ^ n6026 ^ 1'b0 ;
  assign n7116 = ~n7111 & n7115 ;
  assign n7117 = ~n7110 & n7116 ;
  assign n7118 = n7117 ^ n1939 ^ 1'b0 ;
  assign n7119 = n428 | n5491 ;
  assign n7120 = n7119 ^ n5316 ^ 1'b0 ;
  assign n7121 = n4536 & n7120 ;
  assign n7122 = n638 | n874 ;
  assign n7123 = n2435 & ~n7122 ;
  assign n7124 = n3595 | n7123 ;
  assign n7125 = n5417 & ~n6012 ;
  assign n7126 = n340 & n1405 ;
  assign n7127 = ~n79 & n7126 ;
  assign n7128 = ~n402 & n4533 ;
  assign n7129 = n3348 ^ n146 ^ 1'b0 ;
  assign n7130 = ~n423 & n7129 ;
  assign n7131 = n5179 & n7130 ;
  assign n7132 = ~n259 & n7019 ;
  assign n7133 = n4451 & n5138 ;
  assign n7134 = n311 & n6182 ;
  assign n7135 = n7134 ^ n3218 ^ 1'b0 ;
  assign n7136 = n541 | n6886 ;
  assign n7137 = n1876 ^ n349 ^ 1'b0 ;
  assign n7138 = n7137 ^ n150 ^ 1'b0 ;
  assign n7139 = n4056 & ~n7138 ;
  assign n7140 = n6538 ^ n3383 ^ 1'b0 ;
  assign n7141 = n5242 ^ n4677 ^ 1'b0 ;
  assign n7142 = n2120 | n7141 ;
  assign n7143 = n7077 ^ n177 ^ 1'b0 ;
  assign n7145 = n129 | n4007 ;
  assign n7144 = n3554 | n6966 ;
  assign n7146 = n7145 ^ n7144 ^ 1'b0 ;
  assign n7148 = n6647 ^ n4407 ^ 1'b0 ;
  assign n7149 = n7148 ^ n3064 ^ 1'b0 ;
  assign n7147 = n2491 & ~n5803 ;
  assign n7150 = n7149 ^ n7147 ^ 1'b0 ;
  assign n7151 = ~n1455 & n4116 ;
  assign n7152 = ( ~n235 & n2980 ) | ( ~n235 & n3064 ) | ( n2980 & n3064 ) ;
  assign n7153 = n959 & n7152 ;
  assign n7154 = n179 | n3577 ;
  assign n7158 = n4268 & ~n4359 ;
  assign n7159 = n7158 ^ n2821 ^ 1'b0 ;
  assign n7155 = n2455 & n2853 ;
  assign n7156 = n7155 ^ n3402 ^ 1'b0 ;
  assign n7157 = n1347 & n7156 ;
  assign n7160 = n7159 ^ n7157 ^ 1'b0 ;
  assign n7161 = n250 | n1506 ;
  assign n7162 = n7161 ^ n604 ^ 1'b0 ;
  assign n7163 = n7162 ^ n15 ^ 1'b0 ;
  assign n7164 = n152 & ~n7163 ;
  assign n7165 = n5839 ^ n4540 ^ 1'b0 ;
  assign n7166 = n800 & ~n854 ;
  assign n7167 = n5316 & n7166 ;
  assign n7168 = n3928 | n7167 ;
  assign n7169 = n2767 & ~n7168 ;
  assign n7170 = n2040 ^ n208 ^ 1'b0 ;
  assign n7171 = n4274 & n7170 ;
  assign n7172 = n4372 & n7171 ;
  assign n7173 = n5150 ^ n3300 ^ 1'b0 ;
  assign n7174 = n1734 & n7173 ;
  assign n7175 = n6538 & ~n7174 ;
  assign n7176 = n3539 ^ n3066 ^ 1'b0 ;
  assign n7177 = n2186 ^ n1764 ^ n998 ;
  assign n7178 = n6080 & n7177 ;
  assign n7179 = n1251 & n7178 ;
  assign n7180 = n6980 & ~n7179 ;
  assign n7181 = n3805 | n7180 ;
  assign n7182 = n7176 | n7181 ;
  assign n7186 = n549 | n3250 ;
  assign n7187 = ( n1050 & n1943 ) | ( n1050 & ~n7186 ) | ( n1943 & ~n7186 ) ;
  assign n7183 = n262 | n1789 ;
  assign n7184 = n1405 & ~n7183 ;
  assign n7185 = n7184 ^ n3361 ^ 1'b0 ;
  assign n7188 = n7187 ^ n7185 ^ 1'b0 ;
  assign n7189 = n574 | n7188 ;
  assign n7192 = n1964 | n3979 ;
  assign n7193 = n2155 & ~n7192 ;
  assign n7190 = ~n959 & n2202 ;
  assign n7191 = ~n2014 & n7190 ;
  assign n7194 = n7193 ^ n7191 ^ 1'b0 ;
  assign n7195 = n1491 | n7194 ;
  assign n7196 = n2951 ^ n2409 ^ 1'b0 ;
  assign n7197 = n27 & ~n7196 ;
  assign n7198 = ~n2279 & n4632 ;
  assign n7199 = ( n1244 & n5181 ) | ( n1244 & n7198 ) | ( n5181 & n7198 ) ;
  assign n7200 = n2975 & n3178 ;
  assign n7204 = n2895 | n3839 ;
  assign n7205 = n3610 ^ n171 ^ 1'b0 ;
  assign n7206 = n7204 | n7205 ;
  assign n7201 = n2721 ^ n207 ^ 1'b0 ;
  assign n7202 = n1523 | n7201 ;
  assign n7203 = n5385 & ~n7202 ;
  assign n7207 = n7206 ^ n7203 ^ 1'b0 ;
  assign n7208 = n765 | n2282 ;
  assign n7209 = n7208 ^ n3577 ^ 1'b0 ;
  assign n7210 = ~n85 & n940 ;
  assign n7211 = ~n940 & n7210 ;
  assign n7212 = n1191 & ~n2619 ;
  assign n7213 = n2619 & n7212 ;
  assign n7214 = n901 & n7213 ;
  assign n7215 = ~n3710 & n7214 ;
  assign n7216 = n3710 & n7215 ;
  assign n7217 = n7211 | n7216 ;
  assign n7218 = n7211 & ~n7217 ;
  assign n7221 = n638 | n822 ;
  assign n7222 = n822 & ~n7221 ;
  assign n7223 = n140 | n395 ;
  assign n7224 = n7222 & ~n7223 ;
  assign n7225 = x0 & ~n7224 ;
  assign n7226 = ~x0 & n7225 ;
  assign n7227 = n108 | n7226 ;
  assign n7228 = n108 & ~n7227 ;
  assign n7229 = n4855 & ~n7228 ;
  assign n7230 = n7228 & n7229 ;
  assign n7219 = n4964 ^ n197 ^ 1'b0 ;
  assign n7220 = n7219 ^ n2336 ^ 1'b0 ;
  assign n7231 = n7230 ^ n7220 ^ 1'b0 ;
  assign n7232 = n7218 | n7231 ;
  assign n7233 = ( n1055 & n1454 ) | ( n1055 & n3266 ) | ( n1454 & n3266 ) ;
  assign n7234 = n6694 & n7233 ;
  assign n7235 = n2956 | n5320 ;
  assign n7236 = n7235 ^ n572 ^ 1'b0 ;
  assign n7237 = n2159 ^ n378 ^ 1'b0 ;
  assign n7238 = n3521 & n7237 ;
  assign n7239 = n1202 & n1370 ;
  assign n7240 = n6099 ^ n5390 ^ 1'b0 ;
  assign n7241 = n3112 & ~n4831 ;
  assign n7242 = n2452 & ~n7241 ;
  assign n7243 = n1546 & n5925 ;
  assign n7244 = n1306 | n3686 ;
  assign n7245 = n2753 & ~n7244 ;
  assign n7246 = ~n3121 & n4965 ;
  assign n7247 = n7246 ^ n3114 ^ n154 ;
  assign n7248 = ( n5756 & ~n7245 ) | ( n5756 & n7247 ) | ( ~n7245 & n7247 ) ;
  assign n7249 = ~n625 & n1336 ;
  assign n7250 = n7249 ^ n2309 ^ 1'b0 ;
  assign n7251 = n1526 & ~n7250 ;
  assign n7252 = n7251 ^ n695 ^ 1'b0 ;
  assign n7253 = n81 & n7252 ;
  assign n7254 = n7253 ^ n3856 ^ 1'b0 ;
  assign n7255 = n1063 & n1254 ;
  assign n7256 = n7255 ^ n1553 ^ 1'b0 ;
  assign n7257 = n7256 ^ n6486 ^ 1'b0 ;
  assign n7258 = n1948 | n4328 ;
  assign n7259 = n3487 | n7258 ;
  assign n7260 = n4517 & n7259 ;
  assign n7261 = n1488 & n7260 ;
  assign n7262 = n7261 ^ n6333 ^ 1'b0 ;
  assign n7263 = n302 & n3979 ;
  assign n7264 = n6128 | n6172 ;
  assign n7265 = n7263 & ~n7264 ;
  assign n7266 = n4295 | n4705 ;
  assign n7267 = n7266 ^ n3777 ^ n1961 ;
  assign n7268 = n5918 & n7267 ;
  assign n7269 = n1843 ^ n1666 ^ 1'b0 ;
  assign n7270 = n1199 & ~n1450 ;
  assign n7271 = n481 & ~n7270 ;
  assign n7272 = n7271 ^ n1576 ^ 1'b0 ;
  assign n7273 = n3896 ^ n1694 ^ 1'b0 ;
  assign n7274 = n7273 ^ n2869 ^ 1'b0 ;
  assign n7275 = n1863 & n7274 ;
  assign n7276 = n1967 | n4858 ;
  assign n7277 = n5099 ^ n2374 ^ 1'b0 ;
  assign n7278 = ~n4285 & n7277 ;
  assign n7280 = n5333 ^ n582 ^ 1'b0 ;
  assign n7281 = n868 & ~n7280 ;
  assign n7282 = n7281 ^ n415 ^ 1'b0 ;
  assign n7279 = n1918 & n2552 ;
  assign n7283 = n7282 ^ n7279 ^ 1'b0 ;
  assign n7284 = n2048 & n5130 ;
  assign n7285 = ( n523 & n4235 ) | ( n523 & n7284 ) | ( n4235 & n7284 ) ;
  assign n7286 = n387 & ~n7285 ;
  assign n7287 = ~n7283 & n7286 ;
  assign n7288 = n2860 | n5745 ;
  assign n7289 = n253 & ~n1912 ;
  assign n7290 = n1695 ^ n1511 ^ n1036 ;
  assign n7291 = ~n1299 & n7290 ;
  assign n7292 = n7291 ^ n5510 ^ 1'b0 ;
  assign n7293 = n5672 ^ n5667 ^ n1490 ;
  assign n7294 = n2090 & n3124 ;
  assign n7295 = n7290 ^ n1718 ^ 1'b0 ;
  assign n7296 = ~n5693 & n7295 ;
  assign n7297 = n7296 ^ n2833 ^ n2444 ;
  assign n7298 = n79 | n5701 ;
  assign n7299 = n535 & ~n7298 ;
  assign n7300 = ~x10 & n7299 ;
  assign n7301 = ~n4571 & n6073 ;
  assign n7302 = ~n6449 & n7301 ;
  assign n7303 = ~n606 & n2771 ;
  assign n7304 = n7303 ^ n466 ^ 1'b0 ;
  assign n7305 = n7304 ^ n1707 ^ n1251 ;
  assign n7306 = n1967 | n4796 ;
  assign n7307 = n1728 & ~n7306 ;
  assign n7308 = n4770 ^ n4254 ^ 1'b0 ;
  assign n7309 = n2082 & ~n3297 ;
  assign n7310 = n345 & n2495 ;
  assign n7311 = ~n365 & n7310 ;
  assign n7312 = ~n4776 & n7311 ;
  assign n7313 = ~n2961 & n7312 ;
  assign n7314 = n5179 ^ n2042 ^ 1'b0 ;
  assign n7315 = ~n1329 & n4280 ;
  assign n7316 = n7315 ^ n889 ^ 1'b0 ;
  assign n7317 = n7057 & n7316 ;
  assign n7318 = n292 & ~n1456 ;
  assign n7319 = n7318 ^ n287 ^ 1'b0 ;
  assign n7320 = ~n1208 & n7319 ;
  assign n7321 = n7320 ^ n2265 ^ 1'b0 ;
  assign n7322 = ( n1291 & ~n2184 ) | ( n1291 & n5147 ) | ( ~n2184 & n5147 ) ;
  assign n7323 = ~n1295 & n7322 ;
  assign n7324 = n7323 ^ n6927 ^ 1'b0 ;
  assign n7331 = n2077 & ~n2594 ;
  assign n7332 = ~n1464 & n7331 ;
  assign n7325 = ~n2343 & n5371 ;
  assign n7326 = n963 & ~n7325 ;
  assign n7327 = n220 & n3279 ;
  assign n7328 = n7326 | n7327 ;
  assign n7329 = n742 | n7328 ;
  assign n7330 = ~n6722 & n7329 ;
  assign n7333 = n7332 ^ n7330 ^ 1'b0 ;
  assign n7334 = n243 | n5001 ;
  assign n7335 = n7334 ^ n3671 ^ 1'b0 ;
  assign n7336 = n26 | n1434 ;
  assign n7337 = n1837 & ~n7336 ;
  assign n7338 = n21 & n3166 ;
  assign n7339 = ~n3633 & n4030 ;
  assign n7340 = ~n7338 & n7339 ;
  assign n7341 = n7337 | n7340 ;
  assign n7342 = n7335 | n7341 ;
  assign n7343 = ~n397 & n846 ;
  assign n7344 = n451 & n7343 ;
  assign n7345 = n4493 | n5084 ;
  assign n7346 = n7344 & ~n7345 ;
  assign n7347 = n7342 & ~n7346 ;
  assign n7348 = n6506 ^ n2024 ^ 1'b0 ;
  assign n7349 = n2060 & ~n3707 ;
  assign n7350 = n2010 & n6156 ;
  assign n7351 = n4088 & n5615 ;
  assign n7356 = n2038 ^ n1381 ^ n365 ;
  assign n7357 = n6436 | n7356 ;
  assign n7358 = n7357 ^ n282 ^ 1'b0 ;
  assign n7359 = ~n163 & n7358 ;
  assign n7352 = n4046 ^ n3957 ^ n1204 ;
  assign n7353 = n1726 & n7352 ;
  assign n7354 = ~n3428 & n7353 ;
  assign n7355 = n2133 | n7354 ;
  assign n7360 = n7359 ^ n7355 ^ 1'b0 ;
  assign n7361 = n2694 | n3649 ;
  assign n7362 = n1405 | n2993 ;
  assign n7363 = n6243 & ~n6745 ;
  assign n7364 = n322 & n7363 ;
  assign n7365 = n7362 | n7364 ;
  assign n7366 = n7361 & ~n7365 ;
  assign n7367 = ~n645 & n6761 ;
  assign n7368 = n6206 ^ n2140 ^ 1'b0 ;
  assign n7369 = n1560 & ~n4027 ;
  assign n7370 = n6447 & ~n7089 ;
  assign n7371 = n738 ^ n254 ^ 1'b0 ;
  assign n7372 = ~n3312 & n7371 ;
  assign n7373 = n7372 ^ n1005 ^ 1'b0 ;
  assign n7374 = n2394 | n7373 ;
  assign n7375 = n5781 ^ n1460 ^ 1'b0 ;
  assign n7376 = n1065 & ~n2848 ;
  assign n7377 = ~n856 & n4533 ;
  assign n7378 = n6820 | n7377 ;
  assign n7379 = n5748 | n7378 ;
  assign n7380 = n4561 ^ n3272 ^ n2785 ;
  assign n7381 = n910 & ~n7380 ;
  assign n7382 = ~n6092 & n7381 ;
  assign n7383 = n6937 ^ n1732 ^ 1'b0 ;
  assign n7384 = n1739 & ~n4809 ;
  assign n7385 = n1685 & ~n3214 ;
  assign n7386 = ~n7384 & n7385 ;
  assign n7387 = ~n4197 & n7386 ;
  assign n7388 = n7387 ^ n1261 ^ 1'b0 ;
  assign n7389 = n810 ^ n38 ^ 1'b0 ;
  assign n7390 = ( ~n325 & n343 ) | ( ~n325 & n3240 ) | ( n343 & n3240 ) ;
  assign n7391 = n6273 | n7390 ;
  assign n7392 = n3351 & n3833 ;
  assign n7393 = ~n4008 & n7392 ;
  assign n7394 = n3745 & ~n7393 ;
  assign n7395 = ~n296 & n7099 ;
  assign n7396 = n447 & n7395 ;
  assign n7397 = n1988 | n7396 ;
  assign n7398 = n2082 ^ n331 ^ 1'b0 ;
  assign n7399 = n7398 ^ n2713 ^ 1'b0 ;
  assign n7400 = n7399 ^ n6322 ^ 1'b0 ;
  assign n7401 = n360 & n2133 ;
  assign n7402 = n5469 & ~n7401 ;
  assign n7403 = n7084 | n7402 ;
  assign n7404 = n5317 | n7234 ;
  assign n7405 = n6771 ^ n6080 ^ 1'b0 ;
  assign n7406 = n3845 ^ n685 ^ 1'b0 ;
  assign n7407 = n4029 & n7406 ;
  assign n7408 = n4157 & ~n7407 ;
  assign n7409 = n2954 ^ n1522 ^ 1'b0 ;
  assign n7410 = n7408 & n7409 ;
  assign n7412 = ~n1275 & n3220 ;
  assign n7413 = n7412 ^ n3258 ^ 1'b0 ;
  assign n7411 = n2311 | n4858 ;
  assign n7414 = n7413 ^ n7411 ^ 1'b0 ;
  assign n7415 = n2562 ^ n430 ^ 1'b0 ;
  assign n7416 = n2871 & ~n7415 ;
  assign n7417 = n7416 ^ n5958 ^ 1'b0 ;
  assign n7418 = n6764 & ~n7417 ;
  assign n7419 = n3398 ^ n2877 ^ 1'b0 ;
  assign n7420 = n259 & ~n7419 ;
  assign n7421 = n7420 ^ n2495 ^ 1'b0 ;
  assign n7422 = ( n1845 & n4980 ) | ( n1845 & ~n7421 ) | ( n4980 & ~n7421 ) ;
  assign n7423 = ( n1267 & n1829 ) | ( n1267 & n6621 ) | ( n1829 & n6621 ) ;
  assign n7424 = n2529 | n3115 ;
  assign n7425 = n7424 ^ n1584 ^ 1'b0 ;
  assign n7426 = n7208 | n7425 ;
  assign n7427 = n7426 ^ n6681 ^ 1'b0 ;
  assign n7428 = n5886 & ~n6043 ;
  assign n7429 = ~n5642 & n7428 ;
  assign n7430 = n4019 & ~n7429 ;
  assign n7431 = n692 & n3536 ;
  assign n7432 = ~n3536 & n7431 ;
  assign n7433 = n567 | n2172 ;
  assign n7434 = n2172 & ~n7433 ;
  assign n7435 = n7432 | n7434 ;
  assign n7436 = n7432 & ~n7435 ;
  assign n7437 = ~n1204 & n3295 ;
  assign n7438 = ~n633 & n7437 ;
  assign n7439 = n633 & n7438 ;
  assign n7440 = n7439 ^ n6621 ^ 1'b0 ;
  assign n7441 = n7436 | n7440 ;
  assign n7442 = n4564 ^ n2724 ^ n1570 ;
  assign n7443 = n3195 ^ n335 ^ 1'b0 ;
  assign n7444 = n7443 ^ n3934 ^ n88 ;
  assign n7445 = n3090 & ~n4010 ;
  assign n7446 = ~n7444 & n7445 ;
  assign n7447 = ~n474 & n1644 ;
  assign n7448 = ( n358 & ~n1620 ) | ( n358 & n1889 ) | ( ~n1620 & n1889 ) ;
  assign n7449 = n7448 ^ n150 ^ 1'b0 ;
  assign n7450 = n5466 & n7449 ;
  assign n7451 = n7450 ^ n1973 ^ 1'b0 ;
  assign n7452 = n122 | n2655 ;
  assign n7453 = n395 | n7452 ;
  assign n7454 = n411 & ~n7453 ;
  assign n7455 = ( n892 & ~n4764 ) | ( n892 & n7354 ) | ( ~n4764 & n7354 ) ;
  assign n7456 = n3536 ^ n440 ^ n44 ;
  assign n7457 = ~n6722 & n7456 ;
  assign n7458 = n6861 ^ n579 ^ 1'b0 ;
  assign n7459 = n5070 ^ n2647 ^ 1'b0 ;
  assign n7460 = ~n3054 & n4602 ;
  assign n7461 = n592 | n7460 ;
  assign n7462 = n7461 ^ n819 ^ 1'b0 ;
  assign n7463 = n5340 | n7462 ;
  assign n7464 = n7463 ^ n1065 ^ n855 ;
  assign n7465 = n6871 ^ n968 ^ 1'b0 ;
  assign n7466 = n1786 | n7465 ;
  assign n7467 = n6323 ^ n4587 ^ 1'b0 ;
  assign n7468 = n2193 & ~n4287 ;
  assign n7469 = n7468 ^ n4536 ^ 1'b0 ;
  assign n7470 = n1201 | n4477 ;
  assign n7471 = n5860 & ~n7470 ;
  assign n7472 = n7471 ^ n6225 ^ 1'b0 ;
  assign n7473 = n7469 | n7472 ;
  assign n7474 = n5021 & ~n7473 ;
  assign n7475 = n6996 & ~n7474 ;
  assign n7476 = n4958 ^ n2036 ^ n1386 ;
  assign n7477 = n7476 ^ n1993 ^ 1'b0 ;
  assign n7478 = n286 & ~n682 ;
  assign n7479 = n7478 ^ n2309 ^ 1'b0 ;
  assign n7480 = n4296 | n5329 ;
  assign n7481 = ~n326 & n4200 ;
  assign n7482 = n7481 ^ n165 ^ 1'b0 ;
  assign n7483 = ~n954 & n1770 ;
  assign n7484 = n5788 | n7483 ;
  assign n7485 = n4329 & ~n4432 ;
  assign n7486 = n2389 & ~n3766 ;
  assign n7487 = n2833 | n7486 ;
  assign n7488 = n7487 ^ n3361 ^ 1'b0 ;
  assign n7489 = n51 & n675 ;
  assign n7490 = n7489 ^ n472 ^ 1'b0 ;
  assign n7491 = ( ~n4855 & n5733 ) | ( ~n4855 & n7490 ) | ( n5733 & n7490 ) ;
  assign n7492 = ( n514 & n2975 ) | ( n514 & ~n3314 ) | ( n2975 & ~n3314 ) ;
  assign n7493 = n188 & ~n1152 ;
  assign n7494 = n6237 & ~n7493 ;
  assign n7495 = n3361 ^ n796 ^ 1'b0 ;
  assign n7496 = n3818 & n5689 ;
  assign n7497 = ~n7495 & n7496 ;
  assign n7498 = ( n588 & ~n5061 ) | ( n588 & n5897 ) | ( ~n5061 & n5897 ) ;
  assign n7499 = ( ~n2172 & n4092 ) | ( ~n2172 & n6114 ) | ( n4092 & n6114 ) ;
  assign n7500 = n1945 & n6383 ;
  assign n7501 = n2619 ^ n1886 ^ n1469 ;
  assign n7502 = n581 ^ n362 ^ 1'b0 ;
  assign n7503 = ~n2062 & n3353 ;
  assign n7504 = n7503 ^ n3097 ^ 1'b0 ;
  assign n7505 = ~n2136 & n7504 ;
  assign n7506 = n2258 & n7505 ;
  assign n7507 = n7502 & n7506 ;
  assign n7508 = n288 | n1094 ;
  assign n7509 = n5405 | n7508 ;
  assign n7510 = ~n2304 & n7509 ;
  assign n7511 = n4050 ^ n1534 ^ 1'b0 ;
  assign n7512 = n4472 | n7511 ;
  assign n7513 = n4092 & ~n7512 ;
  assign n7514 = ( n695 & n7510 ) | ( n695 & n7513 ) | ( n7510 & n7513 ) ;
  assign n7515 = ( n1260 & n2041 ) | ( n1260 & ~n6006 ) | ( n2041 & ~n6006 ) ;
  assign n7516 = n7245 ^ n1327 ^ 1'b0 ;
  assign n7517 = ~n7515 & n7516 ;
  assign n7518 = ~n7514 & n7517 ;
  assign n7519 = n4583 & n6450 ;
  assign n7520 = n459 & n7519 ;
  assign n7521 = n340 & n7520 ;
  assign n7522 = n6613 ^ n466 ^ n425 ;
  assign n7523 = n7104 ^ n5128 ^ 1'b0 ;
  assign n7524 = n6267 ^ n3167 ^ 1'b0 ;
  assign n7525 = n673 & n1422 ;
  assign n7526 = n7525 ^ n3166 ^ 1'b0 ;
  assign n7527 = n7526 ^ n2468 ^ 1'b0 ;
  assign n7528 = n7524 & n7527 ;
  assign n7529 = n5052 & n5231 ;
  assign n7530 = n3293 & n3665 ;
  assign n7531 = n7530 ^ n1251 ^ 1'b0 ;
  assign n7532 = n3423 & ~n5154 ;
  assign n7533 = n150 | n5120 ;
  assign n7534 = n7533 ^ n2403 ^ 1'b0 ;
  assign n7535 = n3823 | n7534 ;
  assign n7536 = n3418 | n7535 ;
  assign n7537 = n7536 ^ n392 ^ 1'b0 ;
  assign n7538 = ( n105 & n192 ) | ( n105 & n2792 ) | ( n192 & n2792 ) ;
  assign n7539 = ( n188 & n1880 ) | ( n188 & ~n2826 ) | ( n1880 & ~n2826 ) ;
  assign n7540 = n7071 | n7539 ;
  assign n7541 = n3671 | n7540 ;
  assign n7542 = n7541 ^ n182 ^ 1'b0 ;
  assign n7543 = n2985 ^ n1649 ^ 1'b0 ;
  assign n7544 = ~n968 & n7543 ;
  assign n7545 = ~n1439 & n7544 ;
  assign n7546 = n6576 ^ n2921 ^ n1320 ;
  assign n7547 = n5938 ^ n2137 ^ n753 ;
  assign n7548 = n1771 ^ n790 ^ 1'b0 ;
  assign n7549 = ~n7547 & n7548 ;
  assign n7550 = n4343 & ~n5124 ;
  assign n7551 = n3861 ^ n582 ^ 1'b0 ;
  assign n7552 = n4954 & n7551 ;
  assign n7553 = n7552 ^ n1697 ^ 1'b0 ;
  assign n7554 = ~n7550 & n7553 ;
  assign n7555 = ~n2175 & n2471 ;
  assign n7556 = n2474 & n7555 ;
  assign n7557 = n4667 & ~n7556 ;
  assign n7558 = n997 & n7557 ;
  assign n7559 = n972 & n4735 ;
  assign n7560 = n7559 ^ n112 ^ 1'b0 ;
  assign n7561 = n1991 & n7560 ;
  assign n7562 = n7561 ^ n4722 ^ 1'b0 ;
  assign n7563 = n4201 | n7562 ;
  assign n7564 = n4331 | n7563 ;
  assign n7565 = n2533 | n5612 ;
  assign n7566 = n1852 & ~n2921 ;
  assign n7567 = n315 & n7566 ;
  assign n7568 = n7027 ^ n58 ^ 1'b0 ;
  assign n7569 = n160 & ~n1551 ;
  assign n7570 = ~n4570 & n7569 ;
  assign n7571 = n249 & n3646 ;
  assign n7572 = n7571 ^ n209 ^ 1'b0 ;
  assign n7573 = n2885 | n7572 ;
  assign n7574 = n7573 ^ n6856 ^ 1'b0 ;
  assign n7575 = n7574 ^ n5333 ^ 1'b0 ;
  assign n7576 = n3698 | n7575 ;
  assign n7577 = n4206 | n7576 ;
  assign n7578 = n7437 & ~n7577 ;
  assign n7579 = ~n124 & n1669 ;
  assign n7580 = n3082 & ~n7579 ;
  assign n7581 = n7580 ^ n2771 ^ 1'b0 ;
  assign n7582 = n2758 & n5652 ;
  assign n7583 = n3652 ^ n2489 ^ 1'b0 ;
  assign n7584 = n3892 ^ n3613 ^ 1'b0 ;
  assign n7585 = n1098 & n7584 ;
  assign n7586 = n7585 ^ n1462 ^ 1'b0 ;
  assign n7587 = n2883 ^ n975 ^ 1'b0 ;
  assign n7588 = ~n21 & n7587 ;
  assign n7589 = n625 & n7588 ;
  assign n7590 = ( n1459 & n2568 ) | ( n1459 & ~n5469 ) | ( n2568 & ~n5469 ) ;
  assign n7591 = n1664 & n3867 ;
  assign n7592 = n5458 | n7591 ;
  assign n7593 = n6176 & ~n7592 ;
  assign n7594 = n189 | n3641 ;
  assign n7595 = n2408 & ~n7594 ;
  assign n7596 = n7595 ^ n6294 ^ n3741 ;
  assign n7597 = n312 | n2417 ;
  assign n7598 = ( n6889 & ~n7596 ) | ( n6889 & n7597 ) | ( ~n7596 & n7597 ) ;
  assign n7599 = n6392 ^ n4819 ^ 1'b0 ;
  assign n7600 = n2311 | n7599 ;
  assign n7601 = n1883 | n7600 ;
  assign n7602 = ~n6914 & n7601 ;
  assign n7603 = n7602 ^ n5551 ^ 1'b0 ;
  assign n7604 = n4732 | n7603 ;
  assign n7605 = ~n5652 & n6021 ;
  assign n7606 = n7604 | n7605 ;
  assign n7607 = n6912 ^ n1700 ^ 1'b0 ;
  assign n7608 = n2548 ^ n1119 ^ 1'b0 ;
  assign n7609 = n3190 | n7608 ;
  assign n7610 = n7501 ^ n4213 ^ 1'b0 ;
  assign n7611 = n7609 | n7610 ;
  assign n7612 = n2152 ^ n98 ^ 1'b0 ;
  assign n7613 = n3909 & ~n7612 ;
  assign n7614 = n2355 & ~n6121 ;
  assign n7615 = ~n2374 & n4254 ;
  assign n7616 = n7614 & n7615 ;
  assign n7617 = n261 & ~n2935 ;
  assign n7618 = n7617 ^ n3574 ^ n2304 ;
  assign n7621 = n2614 ^ n292 ^ 1'b0 ;
  assign n7622 = n5725 & ~n7621 ;
  assign n7623 = ~n5765 & n7622 ;
  assign n7619 = ~n1656 & n2128 ;
  assign n7620 = n7619 ^ n1176 ^ 1'b0 ;
  assign n7624 = n7623 ^ n7620 ^ 1'b0 ;
  assign n7625 = ~n250 & n2810 ;
  assign n7626 = n3760 & n7625 ;
  assign n7627 = n7626 ^ n2960 ^ n2604 ;
  assign n7628 = ( n2228 & ~n3450 ) | ( n2228 & n4725 ) | ( ~n3450 & n4725 ) ;
  assign n7629 = n5988 ^ n1897 ^ 1'b0 ;
  assign n7630 = ~n7628 & n7629 ;
  assign n7631 = ~n7627 & n7630 ;
  assign n7632 = n3416 | n4914 ;
  assign n7633 = n6161 & ~n7299 ;
  assign n7634 = n311 & ~n541 ;
  assign n7635 = ( n564 & n4539 ) | ( n564 & n7634 ) | ( n4539 & n7634 ) ;
  assign n7636 = n2680 ^ n262 ^ 1'b0 ;
  assign n7637 = n3229 & n7636 ;
  assign n7638 = ~n3610 & n7637 ;
  assign n7639 = n7638 ^ n3001 ^ 1'b0 ;
  assign n7640 = ~n1312 & n4714 ;
  assign n7641 = n1202 & ~n7640 ;
  assign n7642 = n3172 & n7641 ;
  assign n7643 = ~n6504 & n7642 ;
  assign n7644 = n4211 ^ n637 ^ 1'b0 ;
  assign n7645 = n6934 & ~n7644 ;
  assign n7646 = n6842 ^ n1517 ^ 1'b0 ;
  assign n7647 = n4651 & ~n7646 ;
  assign n7649 = n3660 ^ n563 ^ 1'b0 ;
  assign n7650 = n7649 ^ n3245 ^ 1'b0 ;
  assign n7651 = ~n4570 & n7650 ;
  assign n7648 = n3113 ^ n1511 ^ 1'b0 ;
  assign n7652 = n7651 ^ n7648 ^ n1511 ;
  assign n7653 = n367 & ~n1276 ;
  assign n7654 = ~n870 & n3730 ;
  assign n7655 = n7653 & n7654 ;
  assign n7656 = n7655 ^ n7324 ^ 1'b0 ;
  assign n7657 = n4007 ^ n742 ^ n362 ;
  assign n7658 = n2802 | n7657 ;
  assign n7659 = ~n299 & n972 ;
  assign n7660 = ( n33 & n606 ) | ( n33 & ~n7659 ) | ( n606 & ~n7659 ) ;
  assign n7661 = ( n661 & n2569 ) | ( n661 & n7660 ) | ( n2569 & n7660 ) ;
  assign n7662 = n7661 ^ n1145 ^ 1'b0 ;
  assign n7663 = n1545 & ~n7662 ;
  assign n7664 = ~n4595 & n7663 ;
  assign n7665 = ( n1063 & n6423 ) | ( n1063 & n7664 ) | ( n6423 & n7664 ) ;
  assign n7666 = n6988 ^ n2901 ^ 1'b0 ;
  assign n7668 = ~n3438 & n4511 ;
  assign n7667 = ~n2647 & n5849 ;
  assign n7669 = n7668 ^ n7667 ^ 1'b0 ;
  assign n7670 = n7516 ^ n2541 ^ 1'b0 ;
  assign n7672 = ( ~n1109 & n3139 ) | ( ~n1109 & n4809 ) | ( n3139 & n4809 ) ;
  assign n7671 = n3611 & n3759 ;
  assign n7673 = n7672 ^ n7671 ^ 1'b0 ;
  assign n7674 = n4612 ^ n4525 ^ 1'b0 ;
  assign n7675 = n3285 ^ n2709 ^ n1182 ;
  assign n7676 = ( n1066 & n7674 ) | ( n1066 & ~n7675 ) | ( n7674 & ~n7675 ) ;
  assign n7677 = n170 | n1390 ;
  assign n7678 = ( ~n1031 & n2691 ) | ( ~n1031 & n5240 ) | ( n2691 & n5240 ) ;
  assign n7679 = n7678 ^ n3779 ^ 1'b0 ;
  assign n7680 = ~n1306 & n7679 ;
  assign n7681 = n7680 ^ n3146 ^ 1'b0 ;
  assign n7682 = ( n6082 & ~n7677 ) | ( n6082 & n7681 ) | ( ~n7677 & n7681 ) ;
  assign n7683 = ~n3535 & n3611 ;
  assign n7684 = n7277 & n7683 ;
  assign n7685 = n7684 ^ n7655 ^ 1'b0 ;
  assign n7686 = n7685 ^ n6526 ^ 1'b0 ;
  assign n7687 = n5514 ^ n1877 ^ 1'b0 ;
  assign n7688 = n746 & ~n1381 ;
  assign n7689 = n7687 & n7688 ;
  assign n7690 = n7689 ^ n1514 ^ 1'b0 ;
  assign n7691 = n3132 ^ n35 ^ 1'b0 ;
  assign n7692 = n3181 | n3567 ;
  assign n7693 = n7692 ^ n2317 ^ 1'b0 ;
  assign n7694 = n1845 & n5146 ;
  assign n7695 = ~n6226 & n7694 ;
  assign n7696 = ~n1378 & n5781 ;
  assign n7697 = n7696 ^ n5022 ^ 1'b0 ;
  assign n7698 = n7697 ^ n2073 ^ 1'b0 ;
  assign n7699 = n2456 & ~n7698 ;
  assign n7700 = ~n135 & n6172 ;
  assign n7701 = n1769 & n7700 ;
  assign n7702 = n5514 & n7701 ;
  assign n7703 = n2230 | n5503 ;
  assign n7704 = n7703 ^ n883 ^ 1'b0 ;
  assign n7705 = n741 | n3300 ;
  assign n7706 = n4359 | n7702 ;
  assign n7707 = n749 & ~n7706 ;
  assign n7708 = ( n2270 & ~n2460 ) | ( n2270 & n2572 ) | ( ~n2460 & n2572 ) ;
  assign n7709 = n712 & n7708 ;
  assign n7710 = n2558 & n7709 ;
  assign n7711 = n551 & ~n4394 ;
  assign n7712 = n7711 ^ n5111 ^ 1'b0 ;
  assign n7713 = n7712 ^ n224 ^ 1'b0 ;
  assign n7716 = n3194 & ~n3991 ;
  assign n7717 = ~n2515 & n7716 ;
  assign n7715 = n5995 ^ n2272 ^ 1'b0 ;
  assign n7718 = n7717 ^ n7715 ^ n4416 ;
  assign n7714 = ~n4229 & n6915 ;
  assign n7719 = n7718 ^ n7714 ^ 1'b0 ;
  assign n7720 = n7719 ^ n2387 ^ 1'b0 ;
  assign n7721 = ( n1528 & n2484 ) | ( n1528 & ~n7423 ) | ( n2484 & ~n7423 ) ;
  assign n7722 = n1896 ^ n105 ^ 1'b0 ;
  assign n7723 = n7722 ^ n2157 ^ 1'b0 ;
  assign n7724 = n2857 | n7723 ;
  assign n7725 = n2164 & ~n6858 ;
  assign n7726 = n5758 & n7725 ;
  assign n7727 = n5900 ^ n2260 ^ 1'b0 ;
  assign n7728 = n5678 & ~n7727 ;
  assign n7729 = n7728 ^ n4773 ^ 1'b0 ;
  assign n7730 = n7729 ^ n2496 ^ 1'b0 ;
  assign n7731 = n6172 ^ n3105 ^ 1'b0 ;
  assign n7732 = n3139 ^ n1226 ^ 1'b0 ;
  assign n7733 = n3235 & n7732 ;
  assign n7734 = n7733 ^ n316 ^ 1'b0 ;
  assign n7735 = n2794 ^ n884 ^ 1'b0 ;
  assign n7736 = n2389 ^ n1385 ^ n1140 ;
  assign n7737 = n7736 ^ n477 ^ 1'b0 ;
  assign n7738 = n1837 ^ n415 ^ 1'b0 ;
  assign n7739 = n4755 & n7738 ;
  assign n7740 = n7739 ^ n1534 ^ 1'b0 ;
  assign n7741 = ~n3081 & n7740 ;
  assign n7742 = n1758 | n2803 ;
  assign n7743 = n7742 ^ n49 ^ 1'b0 ;
  assign n7744 = ( n3886 & n6871 ) | ( n3886 & n7743 ) | ( n6871 & n7743 ) ;
  assign n7745 = n7741 & n7744 ;
  assign n7746 = n7745 ^ n3438 ^ 1'b0 ;
  assign n7749 = ~n1118 & n1912 ;
  assign n7747 = ~n131 & n968 ;
  assign n7748 = n2095 & ~n7747 ;
  assign n7750 = n7749 ^ n7748 ^ 1'b0 ;
  assign n7751 = ~n4466 & n7750 ;
  assign n7752 = n7751 ^ n4173 ^ 1'b0 ;
  assign n7753 = n5711 ^ n327 ^ n162 ;
  assign n7754 = n7238 ^ n1389 ^ 1'b0 ;
  assign n7755 = n5331 & ~n7754 ;
  assign n7756 = ~n812 & n3961 ;
  assign n7757 = n530 & ~n2376 ;
  assign n7758 = n3998 | n7757 ;
  assign n7759 = ( n56 & ~n1403 ) | ( n56 & n2877 ) | ( ~n1403 & n2877 ) ;
  assign n7760 = n7759 ^ n7685 ^ 1'b0 ;
  assign n7761 = n6653 & n7760 ;
  assign n7762 = n1439 ^ n1390 ^ 1'b0 ;
  assign n7763 = n1109 | n7762 ;
  assign n7764 = n7763 ^ n776 ^ 1'b0 ;
  assign n7765 = n1312 | n7764 ;
  assign n7766 = ( n997 & n3541 ) | ( n997 & n7765 ) | ( n3541 & n7765 ) ;
  assign n7767 = ~n1434 & n7766 ;
  assign n7768 = n744 & n7767 ;
  assign n7769 = ~n372 & n1398 ;
  assign n7770 = n372 & n7769 ;
  assign n7771 = n2583 ^ n2242 ^ n1504 ;
  assign n7772 = n7770 | n7771 ;
  assign n7773 = n7770 & ~n7772 ;
  assign n7774 = n376 & ~n4550 ;
  assign n7775 = n4550 & n7774 ;
  assign n7776 = n7775 ^ n5997 ^ n1300 ;
  assign n7777 = n5121 & ~n7396 ;
  assign n7778 = ~n5273 & n7777 ;
  assign n7779 = n5085 & ~n7778 ;
  assign n7784 = ( ~n1422 & n1542 ) | ( ~n1422 & n2637 ) | ( n1542 & n2637 ) ;
  assign n7780 = n1925 | n3079 ;
  assign n7781 = n7780 ^ n5288 ^ 1'b0 ;
  assign n7782 = n7781 ^ n6489 ^ n5285 ;
  assign n7783 = n291 | n7782 ;
  assign n7785 = n7784 ^ n7783 ^ 1'b0 ;
  assign n7786 = n726 & ~n7785 ;
  assign n7787 = n809 ^ n552 ^ n369 ;
  assign n7788 = ( n3530 & ~n7005 ) | ( n3530 & n7787 ) | ( ~n7005 & n7787 ) ;
  assign n7789 = n2689 & n3896 ;
  assign n7790 = n5906 | n7789 ;
  assign n7791 = n3367 | n7790 ;
  assign n7792 = ~n1122 & n5860 ;
  assign n7793 = n7792 ^ n1136 ^ 1'b0 ;
  assign n7794 = n1023 ^ n755 ^ 1'b0 ;
  assign n7795 = n7683 & n7794 ;
  assign n7796 = n1258 & ~n4464 ;
  assign n7797 = ~n2199 & n7796 ;
  assign n7798 = n150 & ~n7797 ;
  assign n7799 = n7506 ^ n5052 ^ 1'b0 ;
  assign n7800 = n1257 | n2161 ;
  assign n7801 = n7799 & n7800 ;
  assign n7802 = ~n7798 & n7801 ;
  assign n7803 = n4559 ^ n225 ^ 1'b0 ;
  assign n7804 = n3345 | n4991 ;
  assign n7805 = n7803 | n7804 ;
  assign n7806 = n3416 | n7805 ;
  assign n7807 = n3292 & n6488 ;
  assign n7808 = n6396 & n7807 ;
  assign n7809 = ~n1535 & n7808 ;
  assign n7810 = n1065 & n3589 ;
  assign n7811 = n1326 & n7810 ;
  assign n7812 = ~n3015 & n7811 ;
  assign n7813 = n7812 ^ n6765 ^ 1'b0 ;
  assign n7814 = n7813 ^ n412 ^ 1'b0 ;
  assign n7815 = n5145 ^ n1099 ^ 1'b0 ;
  assign n7816 = n3665 | n7815 ;
  assign n7817 = n3680 & ~n4346 ;
  assign n7818 = ~n2899 & n7817 ;
  assign n7819 = n3724 | n7818 ;
  assign n7820 = n4007 & ~n7819 ;
  assign n7821 = n307 | n7820 ;
  assign n7822 = n7821 ^ n199 ^ 1'b0 ;
  assign n7823 = n2677 ^ n1972 ^ 1'b0 ;
  assign n7824 = n6358 | n7823 ;
  assign n7825 = n5110 | n6796 ;
  assign n7826 = n4670 ^ n4425 ^ 1'b0 ;
  assign n7827 = n1907 | n7826 ;
  assign n7828 = n4512 | n4826 ;
  assign n7829 = n7828 ^ n7727 ^ 1'b0 ;
  assign n7830 = ~n671 & n1714 ;
  assign n7831 = ( n3011 & n5474 ) | ( n3011 & n7830 ) | ( n5474 & n7830 ) ;
  assign n7832 = ~n365 & n1431 ;
  assign n7833 = n4976 | n7832 ;
  assign n7834 = ~n1042 & n1816 ;
  assign n7835 = n40 & n7834 ;
  assign n7837 = n493 & ~n1010 ;
  assign n7836 = n2120 | n4061 ;
  assign n7838 = n7837 ^ n7836 ^ 1'b0 ;
  assign n7839 = ~n7835 & n7838 ;
  assign n7840 = n4837 & n7839 ;
  assign n7841 = n7840 ^ n820 ^ 1'b0 ;
  assign n7842 = n2039 ^ n1142 ^ 1'b0 ;
  assign n7843 = ~n5154 & n7842 ;
  assign n7844 = ( ~n1241 & n1401 ) | ( ~n1241 & n1994 ) | ( n1401 & n1994 ) ;
  assign n7845 = n4104 & ~n4368 ;
  assign n7846 = n7845 ^ n277 ^ 1'b0 ;
  assign n7847 = n3547 & ~n5404 ;
  assign n7848 = n4252 | n6548 ;
  assign n7849 = n3315 ^ n1237 ^ 1'b0 ;
  assign n7850 = n6620 | n7849 ;
  assign n7851 = n1480 & ~n3298 ;
  assign n7852 = n233 & n1182 ;
  assign n7853 = ~n233 & n7852 ;
  assign n7854 = n1480 | n7853 ;
  assign n7855 = n7854 ^ n767 ^ 1'b0 ;
  assign n7856 = n5982 ^ n1600 ^ 1'b0 ;
  assign n7857 = n7856 ^ n3139 ^ 1'b0 ;
  assign n7860 = n1199 & ~n2817 ;
  assign n7858 = n6029 & n7082 ;
  assign n7859 = n3111 & n7858 ;
  assign n7861 = n7860 ^ n7859 ^ n255 ;
  assign n7862 = ( ~n2861 & n5516 ) | ( ~n2861 & n6099 ) | ( n5516 & n6099 ) ;
  assign n7863 = n1639 ^ n445 ^ 1'b0 ;
  assign n7864 = ~n7862 & n7863 ;
  assign n7866 = ( n428 & n754 ) | ( n428 & ~n4894 ) | ( n754 & ~n4894 ) ;
  assign n7865 = n828 & n4359 ;
  assign n7867 = n7866 ^ n7865 ^ 1'b0 ;
  assign n7868 = n3576 & n7867 ;
  assign n7869 = ~n1663 & n7868 ;
  assign n7870 = n7803 | n7869 ;
  assign n7871 = n5141 | n7870 ;
  assign n7877 = n4474 & n4835 ;
  assign n7872 = n2630 ^ n1530 ^ 1'b0 ;
  assign n7873 = ~n1789 & n7872 ;
  assign n7874 = n7873 ^ n1252 ^ 1'b0 ;
  assign n7875 = n2675 & n7874 ;
  assign n7876 = n2411 & n7875 ;
  assign n7878 = n7877 ^ n7876 ^ 1'b0 ;
  assign n7879 = ~n1434 & n3173 ;
  assign n7880 = n5033 & ~n7879 ;
  assign n7881 = n2065 & ~n5721 ;
  assign n7882 = n7881 ^ n7663 ^ 1'b0 ;
  assign n7883 = n3745 ^ n627 ^ 1'b0 ;
  assign n7884 = n3115 | n7883 ;
  assign n7885 = n7882 | n7884 ;
  assign n7886 = n7880 | n7885 ;
  assign n7887 = n401 & ~n2094 ;
  assign n7888 = ~n1985 & n7887 ;
  assign n7889 = n7707 & n7888 ;
  assign n7890 = n4464 ^ n1771 ^ 1'b0 ;
  assign n7891 = ~n184 & n7890 ;
  assign n7892 = n1352 & n5378 ;
  assign n7893 = ~n7891 & n7892 ;
  assign n7894 = n2308 ^ n1251 ^ 1'b0 ;
  assign n7895 = ~n2743 & n7894 ;
  assign n7896 = ~n7893 & n7895 ;
  assign n7897 = n6219 & n7896 ;
  assign n7898 = ~n5823 & n7442 ;
  assign n7899 = ~n133 & n835 ;
  assign n7900 = ~n3052 & n3285 ;
  assign n7901 = n1398 | n2695 ;
  assign n7902 = n7900 | n7901 ;
  assign n7903 = n5406 ^ n2455 ^ 1'b0 ;
  assign n7904 = n2051 & ~n7903 ;
  assign n7905 = n7904 ^ n5576 ^ 1'b0 ;
  assign n7906 = n4432 & n7905 ;
  assign n7907 = n3874 | n5668 ;
  assign n7908 = ( n1744 & ~n2189 ) | ( n1744 & n4203 ) | ( ~n2189 & n4203 ) ;
  assign n7909 = n7908 ^ n340 ^ 1'b0 ;
  assign n7910 = n777 | n4180 ;
  assign n7911 = ~n7909 & n7910 ;
  assign n7912 = ~n5334 & n7911 ;
  assign n7913 = n7907 & n7912 ;
  assign n7914 = n2885 ^ n1435 ^ n311 ;
  assign n7915 = n6247 | n6589 ;
  assign n7916 = ( ~n2745 & n7092 ) | ( ~n2745 & n7703 ) | ( n7092 & n7703 ) ;
  assign n7917 = ( n1720 & n7915 ) | ( n1720 & n7916 ) | ( n7915 & n7916 ) ;
  assign n7918 = ~n69 & n3516 ;
  assign n7919 = n7918 ^ n892 ^ n396 ;
  assign n7920 = n216 & ~n2267 ;
  assign n7921 = n1783 & n7920 ;
  assign n7922 = n4105 ^ n1075 ^ 1'b0 ;
  assign n7923 = n7921 & ~n7922 ;
  assign n7924 = n7923 ^ n7165 ^ 1'b0 ;
  assign n7931 = n3724 | n4254 ;
  assign n7926 = n299 ^ n89 ^ 1'b0 ;
  assign n7927 = ~n450 & n2101 ;
  assign n7928 = n7927 ^ n2833 ^ 1'b0 ;
  assign n7929 = ~n7926 & n7928 ;
  assign n7930 = n5001 & ~n7929 ;
  assign n7925 = n598 & ~n4787 ;
  assign n7932 = n7931 ^ n7930 ^ n7925 ;
  assign n7933 = ~n302 & n4859 ;
  assign n7934 = n1769 ^ n305 ^ 1'b0 ;
  assign n7935 = ( ~n539 & n548 ) | ( ~n539 & n2058 ) | ( n548 & n2058 ) ;
  assign n7936 = n5485 ^ n1288 ^ 1'b0 ;
  assign n7937 = ( ~n647 & n5939 ) | ( ~n647 & n7936 ) | ( n5939 & n7936 ) ;
  assign n7938 = n2261 & ~n4398 ;
  assign n7939 = ~n6709 & n7938 ;
  assign n7940 = n414 & ~n6221 ;
  assign n7941 = n7170 ^ n130 ^ 1'b0 ;
  assign n7942 = n5714 ^ n4949 ^ 1'b0 ;
  assign n7943 = n2044 & n7942 ;
  assign n7944 = ~n1779 & n7943 ;
  assign n7945 = ~n3333 & n7944 ;
  assign n7946 = n2700 | n7945 ;
  assign n7947 = n463 & ~n7946 ;
  assign n7948 = n2199 ^ n1066 ^ n40 ;
  assign n7949 = n7948 ^ n5202 ^ 1'b0 ;
  assign n7950 = n4396 | n7949 ;
  assign n7951 = n2154 | n7950 ;
  assign n7952 = n344 | n433 ;
  assign n7953 = n2840 ^ n551 ^ n295 ;
  assign n7954 = n3245 & ~n4696 ;
  assign n7955 = ~n781 & n7954 ;
  assign n7956 = n5492 ^ n2588 ^ 1'b0 ;
  assign n7957 = n468 | n7956 ;
  assign n7958 = n2850 ^ n1418 ^ 1'b0 ;
  assign n7959 = n7135 | n7958 ;
  assign n7960 = n7959 ^ n7643 ^ 1'b0 ;
  assign n7961 = n1092 & ~n5270 ;
  assign n7962 = n2330 ^ n2060 ^ 1'b0 ;
  assign n7963 = n7962 ^ n3917 ^ 1'b0 ;
  assign n7964 = n7961 | n7963 ;
  assign n7965 = ~n3358 & n6372 ;
  assign n7966 = x5 & n6447 ;
  assign n7967 = n425 & n7966 ;
  assign n7968 = n5263 ^ n1534 ^ 1'b0 ;
  assign n7969 = ( ~n868 & n6479 ) | ( ~n868 & n7968 ) | ( n6479 & n7968 ) ;
  assign n7970 = ( ~n2978 & n5623 ) | ( ~n2978 & n7969 ) | ( n5623 & n7969 ) ;
  assign n7971 = n2425 & n7970 ;
  assign n7972 = n439 ^ n372 ^ 1'b0 ;
  assign n7973 = n978 | n7972 ;
  assign n7974 = x1 & ~n3774 ;
  assign n7975 = ~n7973 & n7974 ;
  assign n7976 = n33 | n7975 ;
  assign n7977 = n4122 & ~n7976 ;
  assign n7978 = n4917 ^ n4028 ^ 1'b0 ;
  assign n7979 = n4489 ^ n488 ^ n105 ;
  assign n7980 = n7104 ^ n6732 ^ 1'b0 ;
  assign n7981 = ~n7979 & n7980 ;
  assign n7982 = ~n402 & n2051 ;
  assign n7983 = n4587 ^ n122 ^ 1'b0 ;
  assign n7984 = ( ~n4213 & n7185 ) | ( ~n4213 & n7983 ) | ( n7185 & n7983 ) ;
  assign n7985 = n376 & n898 ;
  assign n7986 = n6059 & n7985 ;
  assign n7987 = n3897 & n7986 ;
  assign n7988 = n578 & n5410 ;
  assign n7989 = n7988 ^ n1231 ^ 1'b0 ;
  assign n7990 = n5118 ^ n1739 ^ 1'b0 ;
  assign n7991 = n2101 & n2398 ;
  assign n7992 = n5363 & n7991 ;
  assign n7993 = n7992 ^ n3867 ^ 1'b0 ;
  assign n7994 = n1103 | n7993 ;
  assign n7995 = n604 & n2090 ;
  assign n7996 = n7995 ^ n459 ^ 1'b0 ;
  assign n7997 = ( n1960 & n4903 ) | ( n1960 & n7145 ) | ( n4903 & n7145 ) ;
  assign n7998 = n7997 ^ n2732 ^ 1'b0 ;
  assign n7999 = ~n1069 & n2336 ;
  assign n8000 = n423 | n5805 ;
  assign n8001 = ~n4142 & n8000 ;
  assign n8002 = n1245 & ~n5041 ;
  assign n8003 = n8001 | n8002 ;
  assign n8004 = ~n1000 & n5031 ;
  assign n8005 = n6275 & n8004 ;
  assign n8006 = ~n7948 & n8005 ;
  assign n8007 = n8006 ^ n1323 ^ 1'b0 ;
  assign n8008 = ( n3652 & n4432 ) | ( n3652 & n6272 ) | ( n4432 & n6272 ) ;
  assign n8009 = n2336 ^ n625 ^ 1'b0 ;
  assign n8010 = n8009 ^ n6063 ^ 1'b0 ;
  assign n8011 = n4170 & ~n6878 ;
  assign n8012 = n7126 ^ n5028 ^ 1'b0 ;
  assign n8013 = n8012 ^ n7238 ^ 1'b0 ;
  assign n8014 = n6083 & ~n8013 ;
  assign n8015 = n597 | n1627 ;
  assign n8016 = n1695 | n8015 ;
  assign n8017 = ~n1018 & n8016 ;
  assign n8018 = n8017 ^ n1863 ^ 1'b0 ;
  assign n8019 = n7972 ^ n521 ^ 1'b0 ;
  assign n8020 = n1469 & n1847 ;
  assign n8021 = ~n5194 & n5841 ;
  assign n8022 = n8021 ^ n3166 ^ 1'b0 ;
  assign n8028 = n931 & ~n1245 ;
  assign n8029 = n1756 & n8028 ;
  assign n8026 = n690 & ~n1972 ;
  assign n8027 = n4688 & ~n8026 ;
  assign n8030 = n8029 ^ n8027 ^ n4260 ;
  assign n8031 = ~n7343 & n8030 ;
  assign n8023 = n1164 | n1336 ;
  assign n8024 = ~n5083 & n8023 ;
  assign n8025 = n6479 | n8024 ;
  assign n8032 = n8031 ^ n8025 ^ 1'b0 ;
  assign n8033 = ~n86 & n104 ;
  assign n8034 = n6740 ^ n4977 ^ n335 ;
  assign n8035 = ~n3831 & n8034 ;
  assign n8036 = n8035 ^ n1546 ^ 1'b0 ;
  assign n8037 = n924 & n7197 ;
  assign n8038 = ~n5030 & n8037 ;
  assign n8039 = n2736 & n8038 ;
  assign n8040 = ~n2242 & n2533 ;
  assign n8041 = ~n867 & n910 ;
  assign n8042 = ( n2859 & n8040 ) | ( n2859 & n8041 ) | ( n8040 & n8041 ) ;
  assign n8043 = n5649 & n6228 ;
  assign n8044 = n4218 & ~n6759 ;
  assign n8045 = ~n4218 & n8044 ;
  assign n8046 = n7530 ^ n695 ^ 1'b0 ;
  assign n8047 = ~n8045 & n8046 ;
  assign n8048 = n5979 ^ n4792 ^ 1'b0 ;
  assign n8049 = x6 & ~n8048 ;
  assign n8050 = n4537 ^ n1286 ^ 1'b0 ;
  assign n8051 = n7927 & ~n8050 ;
  assign n8052 = n6927 ^ n3160 ^ 1'b0 ;
  assign n8053 = n8051 & n8052 ;
  assign n8054 = ~n1329 & n3562 ;
  assign n8055 = ~n104 & n1857 ;
  assign n8056 = n4058 & n8055 ;
  assign n8057 = ~n8054 & n8056 ;
  assign n8058 = n229 & ~n8057 ;
  assign n8059 = n7430 ^ n548 ^ 1'b0 ;
  assign n8060 = n3552 | n8059 ;
  assign n8061 = ( ~n4116 & n8058 ) | ( ~n4116 & n8060 ) | ( n8058 & n8060 ) ;
  assign n8062 = ~n33 & n2674 ;
  assign n8063 = n5023 & ~n5182 ;
  assign n8064 = ~n4632 & n8063 ;
  assign n8065 = n5727 | n8064 ;
  assign n8066 = n8062 & ~n8065 ;
  assign n8067 = n1434 | n1789 ;
  assign n8068 = n8067 ^ n3403 ^ 1'b0 ;
  assign n8069 = n6020 ^ n2922 ^ 1'b0 ;
  assign n8070 = n8068 & n8069 ;
  assign n8071 = n8070 ^ n234 ^ 1'b0 ;
  assign n8072 = n371 | n4535 ;
  assign n8073 = ~n150 & n1688 ;
  assign n8074 = n926 & ~n8073 ;
  assign n8075 = n1542 | n8074 ;
  assign n8076 = n8075 ^ n5016 ^ 1'b0 ;
  assign n8077 = n2380 ^ n175 ^ 1'b0 ;
  assign n8078 = n5420 ^ n708 ^ 1'b0 ;
  assign n8079 = n6233 ^ n5059 ^ 1'b0 ;
  assign n8084 = n3406 ^ n802 ^ 1'b0 ;
  assign n8085 = n1050 ^ n316 ^ 1'b0 ;
  assign n8086 = n8084 & ~n8085 ;
  assign n8082 = ~n4235 & n5089 ;
  assign n8080 = n1369 ^ n627 ^ 1'b0 ;
  assign n8081 = ( n792 & ~n5523 ) | ( n792 & n8080 ) | ( ~n5523 & n8080 ) ;
  assign n8083 = n8082 ^ n8081 ^ 1'b0 ;
  assign n8087 = n8086 ^ n8083 ^ 1'b0 ;
  assign n8088 = n4814 & n8087 ;
  assign n8089 = n8088 ^ n1337 ^ 1'b0 ;
  assign n8090 = n1454 | n1700 ;
  assign n8091 = n160 | n8090 ;
  assign n8092 = n682 | n5800 ;
  assign n8093 = n8091 | n8092 ;
  assign n8094 = ~n167 & n5082 ;
  assign n8095 = n8094 ^ n2128 ^ 1'b0 ;
  assign n8096 = ~n726 & n6350 ;
  assign n8097 = n3762 & n8096 ;
  assign n8098 = n8097 ^ n3873 ^ 1'b0 ;
  assign n8099 = n8095 & n8098 ;
  assign n8100 = n4457 & n5785 ;
  assign n8101 = n505 & n3480 ;
  assign n8102 = n1408 ^ n1398 ^ 1'b0 ;
  assign n8103 = n8102 ^ n2662 ^ 1'b0 ;
  assign n8104 = n4993 & ~n8103 ;
  assign n8105 = n760 & n5317 ;
  assign n8106 = n7495 ^ n910 ^ 1'b0 ;
  assign n8107 = ~n8105 & n8106 ;
  assign n8108 = n261 | n5247 ;
  assign n8109 = n8108 ^ n772 ^ 1'b0 ;
  assign n8110 = n8109 ^ n2045 ^ 1'b0 ;
  assign n8111 = n283 | n8110 ;
  assign n8112 = ~n4696 & n8111 ;
  assign n8113 = n4696 & n8112 ;
  assign n8114 = n7707 | n8113 ;
  assign n8115 = n8113 & ~n8114 ;
  assign n8116 = n1374 & ~n1623 ;
  assign n8117 = n8116 ^ n3193 ^ 1'b0 ;
  assign n8118 = n2689 ^ n1477 ^ 1'b0 ;
  assign n8119 = n4537 ^ n2554 ^ 1'b0 ;
  assign n8120 = n8119 ^ n6028 ^ 1'b0 ;
  assign n8121 = n305 & n488 ;
  assign n8122 = n2780 & n8121 ;
  assign n8123 = n4005 ^ n280 ^ 1'b0 ;
  assign n8124 = n8122 | n8123 ;
  assign n8125 = n5569 | n8124 ;
  assign n8126 = n8120 | n8125 ;
  assign n8127 = n5328 ^ n695 ^ 1'b0 ;
  assign n8128 = n294 | n835 ;
  assign n8129 = n6731 ^ n2932 ^ 1'b0 ;
  assign n8130 = ~n4386 & n5982 ;
  assign n8131 = n2890 ^ n2114 ^ 1'b0 ;
  assign n8132 = n3770 & n8131 ;
  assign n8133 = n6127 ^ n543 ^ 1'b0 ;
  assign n8134 = ~n8132 & n8133 ;
  assign n8135 = n5336 ^ n1558 ^ n1081 ;
  assign n8136 = n3896 & n7041 ;
  assign n8137 = n6491 ^ n477 ^ 1'b0 ;
  assign n8138 = n3274 | n8137 ;
  assign n8139 = n6498 ^ n609 ^ 1'b0 ;
  assign n8140 = ~n323 & n7329 ;
  assign n8141 = n1367 & n8140 ;
  assign n8142 = n7187 | n7732 ;
  assign n8143 = n2238 | n4214 ;
  assign n8144 = n8143 ^ n4333 ^ 1'b0 ;
  assign n8145 = n5833 ^ n4083 ^ 1'b0 ;
  assign n8146 = n8145 ^ n1668 ^ 1'b0 ;
  assign n8147 = ~n8144 & n8146 ;
  assign n8148 = n2730 | n6553 ;
  assign n8150 = n5859 ^ n5032 ^ 1'b0 ;
  assign n8149 = n3314 | n7139 ;
  assign n8151 = n8150 ^ n8149 ^ 1'b0 ;
  assign n8152 = ( n1528 & ~n5422 ) | ( n1528 & n8151 ) | ( ~n5422 & n8151 ) ;
  assign n8153 = n3105 ^ n2697 ^ 1'b0 ;
  assign n8154 = n3131 & n4949 ;
  assign n8155 = n376 & ~n7498 ;
  assign n8156 = n5149 & n8155 ;
  assign n8157 = ~n2483 & n3207 ;
  assign n8158 = n2664 ^ n1116 ^ 1'b0 ;
  assign n8159 = n1243 & n8158 ;
  assign n8160 = n2691 & n2921 ;
  assign n8161 = n8160 ^ n2207 ^ 1'b0 ;
  assign n8162 = n8161 ^ n5940 ^ 1'b0 ;
  assign n8163 = ~n1490 & n8162 ;
  assign n8164 = n8163 ^ n2367 ^ 1'b0 ;
  assign n8165 = n8159 & ~n8164 ;
  assign n8166 = n8157 & ~n8165 ;
  assign n8167 = n2760 & n4059 ;
  assign n8168 = n8167 ^ n1297 ^ 1'b0 ;
  assign n8169 = n5834 ^ n1615 ^ 1'b0 ;
  assign n8170 = n4036 & ~n8169 ;
  assign n8171 = n8168 & n8170 ;
  assign n8172 = ~n3363 & n3584 ;
  assign n8173 = n219 | n8172 ;
  assign n8174 = n44 & n1837 ;
  assign n8179 = n806 & ~n2125 ;
  assign n8180 = n8179 ^ n5805 ^ 1'b0 ;
  assign n8181 = n1327 | n8180 ;
  assign n8182 = n8181 ^ n1670 ^ 1'b0 ;
  assign n8175 = n7588 ^ n1917 ^ 1'b0 ;
  assign n8176 = n4264 | n8175 ;
  assign n8177 = n8176 ^ n490 ^ 1'b0 ;
  assign n8178 = ~n6760 & n8177 ;
  assign n8183 = n8182 ^ n8178 ^ 1'b0 ;
  assign n8185 = n3457 & ~n4218 ;
  assign n8186 = n8185 ^ n1385 ^ 1'b0 ;
  assign n8184 = n961 & n6907 ;
  assign n8187 = n8186 ^ n8184 ^ 1'b0 ;
  assign n8188 = ( n832 & n4020 ) | ( n832 & ~n4461 ) | ( n4020 & ~n4461 ) ;
  assign n8189 = n1132 | n8188 ;
  assign n8190 = n8189 ^ n5426 ^ 1'b0 ;
  assign n8191 = n7586 ^ n7096 ^ 1'b0 ;
  assign n8192 = n8190 | n8191 ;
  assign n8193 = n6941 | n8064 ;
  assign n8194 = n8193 ^ n3202 ^ 1'b0 ;
  assign n8195 = n5300 & ~n8194 ;
  assign n8196 = n320 | n2152 ;
  assign n8197 = n8196 ^ n4028 ^ 1'b0 ;
  assign n8198 = n8197 ^ n4279 ^ 1'b0 ;
  assign n8199 = ( ~n640 & n2576 ) | ( ~n640 & n5755 ) | ( n2576 & n5755 ) ;
  assign n8200 = ~n987 & n3176 ;
  assign n8201 = ( n2628 & n3937 ) | ( n2628 & ~n5484 ) | ( n3937 & ~n5484 ) ;
  assign n8203 = n5937 ^ n4220 ^ 1'b0 ;
  assign n8204 = n1914 & ~n8203 ;
  assign n8205 = n132 & n809 ;
  assign n8206 = ~n121 & n8205 ;
  assign n8207 = ~n1145 & n8206 ;
  assign n8208 = n8204 & n8207 ;
  assign n8202 = n535 & ~n5135 ;
  assign n8209 = n8208 ^ n8202 ^ 1'b0 ;
  assign n8210 = n1308 & ~n8132 ;
  assign n8211 = n7422 & ~n8210 ;
  assign n8212 = n1469 & ~n5168 ;
  assign n8213 = ~n2252 & n2785 ;
  assign n8214 = n8213 ^ n2168 ^ 1'b0 ;
  assign n8215 = ~n3827 & n8214 ;
  assign n8216 = ~n104 & n470 ;
  assign n8217 = n1233 & ~n2619 ;
  assign n8218 = n1568 | n8217 ;
  assign n8219 = n3496 | n8218 ;
  assign n8220 = n2663 | n3409 ;
  assign n8221 = n5121 & n6029 ;
  assign n8222 = n8221 ^ n3415 ^ 1'b0 ;
  assign n8223 = ( n1161 & n3621 ) | ( n1161 & n8222 ) | ( n3621 & n8222 ) ;
  assign n8224 = ( n1241 & n2895 ) | ( n1241 & n8223 ) | ( n2895 & n8223 ) ;
  assign n8225 = n1378 | n6496 ;
  assign n8226 = ~n4390 & n6790 ;
  assign n8227 = ~n6110 & n8226 ;
  assign n8228 = n1505 & n8227 ;
  assign n8229 = n7941 ^ n3962 ^ 1'b0 ;
  assign n8230 = n3641 ^ n1978 ^ 1'b0 ;
  assign n8231 = n3508 & n3530 ;
  assign n8232 = n8231 ^ n1775 ^ 1'b0 ;
  assign n8233 = n209 & ~n2250 ;
  assign n8234 = n3680 & n8233 ;
  assign n8235 = ~n8232 & n8234 ;
  assign n8236 = ( n1770 & ~n8230 ) | ( n1770 & n8235 ) | ( ~n8230 & n8235 ) ;
  assign n8239 = n4537 ^ n3880 ^ n2195 ;
  assign n8240 = n8239 ^ n1187 ^ 1'b0 ;
  assign n8241 = n7879 & ~n8240 ;
  assign n8237 = ( n1891 & n3227 ) | ( n1891 & n7883 ) | ( n3227 & n7883 ) ;
  assign n8238 = n3272 | n8237 ;
  assign n8242 = n8241 ^ n8238 ^ 1'b0 ;
  assign n8243 = n4013 & ~n6919 ;
  assign n8244 = n1845 ^ n131 ^ 1'b0 ;
  assign n8245 = ~n2151 & n4540 ;
  assign n8246 = n8245 ^ n6589 ^ 1'b0 ;
  assign n8247 = n4599 ^ n2991 ^ 1'b0 ;
  assign n8248 = ~n397 & n8247 ;
  assign n8249 = n595 & n910 ;
  assign n8250 = n8249 ^ n8076 ^ 1'b0 ;
  assign n8251 = n8248 | n8250 ;
  assign n8252 = n4727 ^ n2382 ^ 1'b0 ;
  assign n8253 = n7475 ^ n6174 ^ 1'b0 ;
  assign n8254 = n1063 ^ n445 ^ 1'b0 ;
  assign n8255 = n8254 ^ n7448 ^ 1'b0 ;
  assign n8256 = n1761 & n8255 ;
  assign n8257 = ~n150 & n8256 ;
  assign n8258 = n5520 & n8257 ;
  assign n8259 = ~n5170 & n5756 ;
  assign n8260 = n3034 ^ n2923 ^ 1'b0 ;
  assign n8261 = ~n1454 & n8260 ;
  assign n8262 = n8261 ^ n6426 ^ 1'b0 ;
  assign n8263 = ~n2018 & n4670 ;
  assign n8264 = ~n4050 & n8263 ;
  assign n8265 = ~n2717 & n8264 ;
  assign n8266 = n7927 ^ n6427 ^ 1'b0 ;
  assign n8267 = ~n6930 & n8266 ;
  assign n8268 = n574 | n4537 ;
  assign n8269 = n3633 & ~n8268 ;
  assign n8270 = n286 | n6160 ;
  assign n8272 = n785 & ~n1306 ;
  assign n8273 = n570 & n8272 ;
  assign n8274 = n4470 & n8273 ;
  assign n8271 = n1867 | n4491 ;
  assign n8275 = n8274 ^ n8271 ^ 1'b0 ;
  assign n8276 = n8275 ^ n7952 ^ n1700 ;
  assign n8277 = n5673 & n8024 ;
  assign n8278 = ( n183 & ~n3229 ) | ( n183 & n6976 ) | ( ~n3229 & n6976 ) ;
  assign n8279 = n2166 ^ n356 ^ 1'b0 ;
  assign n8280 = n3487 & ~n8279 ;
  assign n8281 = n8280 ^ n1868 ^ 1'b0 ;
  assign n8282 = ( ~n1366 & n6575 ) | ( ~n1366 & n7717 ) | ( n6575 & n7717 ) ;
  assign n8283 = ~n2022 & n3066 ;
  assign n8284 = n1295 & ~n1918 ;
  assign n8285 = n8284 ^ n5459 ^ n2159 ;
  assign n8286 = n5865 & n8285 ;
  assign n8287 = ~n474 & n1968 ;
  assign n8288 = n8287 ^ n2860 ^ 1'b0 ;
  assign n8289 = ( ~n1422 & n3911 ) | ( ~n1422 & n7948 ) | ( n3911 & n7948 ) ;
  assign n8290 = n315 & n6500 ;
  assign n8291 = n1143 & n8290 ;
  assign n8292 = ( n4958 & n8289 ) | ( n4958 & n8291 ) | ( n8289 & n8291 ) ;
  assign n8293 = ~n2927 & n6988 ;
  assign n8294 = n946 | n1346 ;
  assign n8295 = n8294 ^ n271 ^ 1'b0 ;
  assign n8296 = n8295 ^ n5510 ^ n4613 ;
  assign n8299 = n3955 ^ n2623 ^ 1'b0 ;
  assign n8300 = n1202 & ~n8299 ;
  assign n8297 = n6269 ^ n3932 ^ 1'b0 ;
  assign n8298 = n1788 | n8297 ;
  assign n8301 = n8300 ^ n8298 ^ 1'b0 ;
  assign n8302 = n3827 | n7452 ;
  assign n8308 = ~n568 & n5602 ;
  assign n8303 = ( n63 & n606 ) | ( n63 & ~n1179 ) | ( n606 & ~n1179 ) ;
  assign n8304 = n4997 ^ n2641 ^ 1'b0 ;
  assign n8305 = n224 & n8304 ;
  assign n8306 = n8303 | n8305 ;
  assign n8307 = n1783 & ~n8306 ;
  assign n8309 = n8308 ^ n8307 ^ n4545 ;
  assign n8310 = n5342 ^ n3875 ^ 1'b0 ;
  assign n8311 = n2996 ^ n2267 ^ 1'b0 ;
  assign n8312 = n2097 & n2749 ;
  assign n8313 = n8311 & ~n8312 ;
  assign n8314 = n2747 & n8313 ;
  assign n8315 = n5997 ^ n4914 ^ n259 ;
  assign n8316 = n619 & ~n8315 ;
  assign n8317 = n7717 & n8316 ;
  assign n8318 = n492 & n4250 ;
  assign n8319 = ~n2154 & n8318 ;
  assign n8320 = n138 & n5900 ;
  assign n8321 = n8319 & n8320 ;
  assign n8322 = ~n5059 & n8055 ;
  assign n8323 = n4348 & n8322 ;
  assign n8324 = n8323 ^ n2492 ^ 1'b0 ;
  assign n8325 = ( n338 & n598 ) | ( n338 & ~n3867 ) | ( n598 & ~n3867 ) ;
  assign n8326 = ~n1141 & n8325 ;
  assign n8327 = n7338 ^ n5128 ^ n1660 ;
  assign n8328 = ~n987 & n1499 ;
  assign n8329 = n1937 & n2257 ;
  assign n8330 = ~n8328 & n8329 ;
  assign n8331 = n6452 ^ n1868 ^ n1365 ;
  assign n8332 = ~n1662 & n3817 ;
  assign n8333 = n8331 | n8332 ;
  assign n8334 = n8333 ^ n5027 ^ 1'b0 ;
  assign n8335 = n1485 ^ n189 ^ 1'b0 ;
  assign n8336 = n7396 | n8335 ;
  assign n8337 = n6991 & ~n8336 ;
  assign n8338 = n1857 ^ n220 ^ 1'b0 ;
  assign n8339 = n8337 & ~n8338 ;
  assign n8340 = n8339 ^ n1755 ^ 1'b0 ;
  assign n8341 = n8340 ^ n5607 ^ 1'b0 ;
  assign n8342 = n8273 ^ n5810 ^ n4324 ;
  assign n8343 = n4267 ^ n1124 ^ 1'b0 ;
  assign n8344 = n7176 & n8343 ;
  assign n8345 = ~n5583 & n7810 ;
  assign n8346 = n291 & n8345 ;
  assign n8347 = n5141 ^ n839 ^ 1'b0 ;
  assign n8348 = n8346 | n8347 ;
  assign n8349 = n8348 ^ n5030 ^ 1'b0 ;
  assign n8350 = n1743 & n5366 ;
  assign n8351 = n6878 ^ n1056 ^ 1'b0 ;
  assign n8352 = ( n835 & n1092 ) | ( n835 & ~n3382 ) | ( n1092 & ~n3382 ) ;
  assign n8353 = n8352 ^ n1633 ^ 1'b0 ;
  assign n8354 = ~n1714 & n8353 ;
  assign n8355 = n6730 ^ n4651 ^ n4297 ;
  assign n8356 = n1598 & n2306 ;
  assign n8357 = ~n8355 & n8356 ;
  assign n8358 = ~n560 & n5052 ;
  assign n8359 = n8358 ^ n2772 ^ 1'b0 ;
  assign n8360 = n5408 ^ n5161 ^ n138 ;
  assign n8361 = ~n6806 & n8360 ;
  assign n8362 = n2601 & n8361 ;
  assign n8363 = n5217 ^ n208 ^ 1'b0 ;
  assign n8364 = n8363 ^ n4676 ^ 1'b0 ;
  assign n8365 = n3424 & ~n8364 ;
  assign n8366 = n8365 ^ n8324 ^ 1'b0 ;
  assign n8367 = n471 & n996 ;
  assign n8368 = n2849 ^ n567 ^ 1'b0 ;
  assign n8369 = n8368 ^ n2356 ^ 1'b0 ;
  assign n8370 = ~n3781 & n8369 ;
  assign n8371 = n2662 & n8370 ;
  assign n8372 = n8371 ^ n6941 ^ 1'b0 ;
  assign n8373 = n2951 & n7179 ;
  assign n8374 = n1316 & n6408 ;
  assign n8375 = n8374 ^ n263 ^ 1'b0 ;
  assign n8376 = n5896 ^ n1624 ^ 1'b0 ;
  assign n8377 = n8375 | n8376 ;
  assign n8378 = n8377 ^ n7004 ^ 1'b0 ;
  assign n8379 = n4005 ^ n194 ^ 1'b0 ;
  assign n8380 = n910 | n8379 ;
  assign n8381 = n3549 ^ n2291 ^ 1'b0 ;
  assign n8382 = ~n536 & n561 ;
  assign n8383 = n8382 ^ n2735 ^ 1'b0 ;
  assign n8384 = n6311 ^ n1196 ^ 1'b0 ;
  assign n8385 = n588 | n8384 ;
  assign n8386 = n582 & ~n971 ;
  assign n8387 = n8386 ^ n4613 ^ 1'b0 ;
  assign n8388 = n3723 & n8387 ;
  assign n8389 = n2328 & ~n3518 ;
  assign n8390 = n8388 & n8389 ;
  assign n8391 = ~n8385 & n8390 ;
  assign n8392 = n8391 ^ n4993 ^ 1'b0 ;
  assign n8393 = n6888 ^ n1594 ^ 1'b0 ;
  assign n8394 = n914 & ~n7873 ;
  assign n8395 = ~n1847 & n8394 ;
  assign n8396 = n8395 ^ n2598 ^ 1'b0 ;
  assign n8402 = n5809 ^ n978 ^ n799 ;
  assign n8403 = n8402 ^ n3372 ^ 1'b0 ;
  assign n8397 = n4626 | n5152 ;
  assign n8398 = n2386 | n8247 ;
  assign n8399 = n8397 & ~n8398 ;
  assign n8400 = n8020 | n8399 ;
  assign n8401 = n4995 & ~n8400 ;
  assign n8404 = n8403 ^ n8401 ^ n1956 ;
  assign n8406 = n4422 ^ n224 ^ 1'b0 ;
  assign n8405 = n2641 | n2869 ;
  assign n8407 = n8406 ^ n8405 ^ 1'b0 ;
  assign n8408 = n8251 ^ n226 ^ 1'b0 ;
  assign n8409 = n2138 ^ n228 ^ 1'b0 ;
  assign n8410 = n7683 & ~n8409 ;
  assign n8411 = n8410 ^ n2588 ^ 1'b0 ;
  assign n8412 = n805 & ~n8217 ;
  assign n8413 = ( n1378 & n4977 ) | ( n1378 & n7527 ) | ( n4977 & n7527 ) ;
  assign n8414 = n3088 | n3214 ;
  assign n8415 = n5612 | n8414 ;
  assign n8416 = n2087 | n8415 ;
  assign n8417 = ( n98 & n1284 ) | ( n98 & n6149 ) | ( n1284 & n6149 ) ;
  assign n8418 = ~n2634 & n8417 ;
  assign n8419 = n8418 ^ n5396 ^ 1'b0 ;
  assign n8420 = n926 | n1233 ;
  assign n8421 = n1184 | n8420 ;
  assign n8422 = n4859 & n8421 ;
  assign n8423 = n8422 ^ n4406 ^ 1'b0 ;
  assign n8424 = n2304 ^ n2277 ^ 1'b0 ;
  assign n8425 = n6768 ^ n475 ^ 1'b0 ;
  assign n8426 = ( n2876 & n8424 ) | ( n2876 & n8425 ) | ( n8424 & n8425 ) ;
  assign n8427 = n1594 & n5450 ;
  assign n8431 = n3548 & n6756 ;
  assign n8432 = n8431 ^ n2811 ^ 1'b0 ;
  assign n8429 = n820 & n6133 ;
  assign n8430 = n5722 & n8429 ;
  assign n8428 = n5649 ^ n4185 ^ 1'b0 ;
  assign n8433 = n8432 ^ n8430 ^ n8428 ;
  assign n8434 = n8148 ^ n2321 ^ 1'b0 ;
  assign n8435 = n195 | n8434 ;
  assign n8436 = n2812 ^ n2753 ^ n1884 ;
  assign n8437 = n8436 ^ n1620 ^ 1'b0 ;
  assign n8438 = n5033 & n8437 ;
  assign n8440 = ~n574 & n4367 ;
  assign n8439 = ~n1657 & n2445 ;
  assign n8441 = n8440 ^ n8439 ^ 1'b0 ;
  assign n8442 = n6664 ^ n124 ^ 1'b0 ;
  assign n8443 = n6842 & ~n8442 ;
  assign n8444 = n1528 & ~n7657 ;
  assign n8445 = ~n8443 & n8444 ;
  assign n8446 = n3724 ^ n1386 ^ 1'b0 ;
  assign n8447 = n3584 ^ n856 ^ 1'b0 ;
  assign n8448 = n8447 ^ n2065 ^ n261 ;
  assign n8449 = n6628 | n8448 ;
  assign n8450 = n1711 & ~n2588 ;
  assign n8451 = n207 & n253 ;
  assign n8452 = n8451 ^ n7357 ^ 1'b0 ;
  assign n8453 = n6106 ^ n2066 ^ 1'b0 ;
  assign n8454 = n8453 ^ n5124 ^ 1'b0 ;
  assign n8455 = n2161 & ~n5538 ;
  assign n8456 = n1759 & n8455 ;
  assign n8457 = n5458 & ~n8456 ;
  assign n8458 = n2173 & ~n2367 ;
  assign n8459 = n965 & n8458 ;
  assign n8460 = ~n1057 & n8459 ;
  assign n8461 = n8460 ^ n4030 ^ 1'b0 ;
  assign n8462 = n3833 ^ n634 ^ 1'b0 ;
  assign n8463 = n2494 & n8462 ;
  assign n8464 = ~n1181 & n4476 ;
  assign n8465 = n8464 ^ n2095 ^ 1'b0 ;
  assign n8466 = n6758 | n8465 ;
  assign n8467 = n8466 ^ n5369 ^ 1'b0 ;
  assign n8468 = ~n3919 & n8467 ;
  assign n8473 = n5671 ^ n1035 ^ 1'b0 ;
  assign n8474 = n3962 | n8473 ;
  assign n8475 = n8474 ^ n4809 ^ 1'b0 ;
  assign n8469 = n1558 & ~n3303 ;
  assign n8470 = ~n1517 & n8469 ;
  assign n8471 = n7736 & ~n8470 ;
  assign n8472 = ~n7665 & n8471 ;
  assign n8476 = n8475 ^ n8472 ^ 1'b0 ;
  assign n8480 = n6006 ^ n3942 ^ 1'b0 ;
  assign n8477 = n1819 | n3259 ;
  assign n8478 = n8477 ^ n3926 ^ n2082 ;
  assign n8479 = n4347 & ~n8478 ;
  assign n8481 = n8480 ^ n8479 ^ 1'b0 ;
  assign n8482 = n3926 ^ n2321 ^ 1'b0 ;
  assign n8483 = ( n479 & n2645 ) | ( n479 & n8482 ) | ( n2645 & n8482 ) ;
  assign n8484 = n6783 & ~n7280 ;
  assign n8485 = ~n8483 & n8484 ;
  assign n8486 = n3919 ^ n1025 ^ 1'b0 ;
  assign n8487 = n1744 | n8486 ;
  assign n8488 = n7162 & ~n8487 ;
  assign n8489 = n8488 ^ n998 ^ 1'b0 ;
  assign n8490 = n2539 ^ n1845 ^ 1'b0 ;
  assign n8491 = n4007 ^ n2666 ^ 1'b0 ;
  assign n8492 = n1441 ^ n976 ^ 1'b0 ;
  assign n8493 = n5883 ^ n3529 ^ 1'b0 ;
  assign n8494 = n8492 & ~n8493 ;
  assign n8495 = n5302 ^ n184 ^ 1'b0 ;
  assign n8496 = n2675 ^ n35 ^ 1'b0 ;
  assign n8497 = n2072 & n8496 ;
  assign n8498 = n8497 ^ n974 ^ 1'b0 ;
  assign n8499 = n2014 & n8498 ;
  assign n8500 = n8499 ^ n331 ^ 1'b0 ;
  assign n8501 = n2473 & ~n8500 ;
  assign n8502 = ~n8495 & n8501 ;
  assign n8503 = n8323 ^ n1666 ^ 1'b0 ;
  assign n8504 = n2155 | n4097 ;
  assign n8505 = n746 | n8504 ;
  assign n8506 = ( n1204 & n6355 ) | ( n1204 & n8505 ) | ( n6355 & n8505 ) ;
  assign n8507 = n4121 ^ n861 ^ 1'b0 ;
  assign n8508 = ( n3223 & ~n3967 ) | ( n3223 & n7371 ) | ( ~n3967 & n7371 ) ;
  assign n8509 = n8508 ^ n622 ^ 1'b0 ;
  assign n8510 = n8507 & ~n8509 ;
  assign n8511 = n1531 | n4999 ;
  assign n8512 = n2446 & ~n8511 ;
  assign n8513 = ( ~n181 & n1688 ) | ( ~n181 & n8512 ) | ( n1688 & n8512 ) ;
  assign n8514 = ~n1771 & n8513 ;
  assign n8515 = n3078 & ~n8225 ;
  assign n8516 = n3124 & ~n7337 ;
  assign n8517 = n183 | n2253 ;
  assign n8518 = n8516 | n8517 ;
  assign n8519 = n2535 ^ n1502 ^ 1'b0 ;
  assign n8520 = n7164 ^ n6954 ^ 1'b0 ;
  assign n8521 = n8519 & n8520 ;
  assign n8522 = ~n667 & n2465 ;
  assign n8523 = ( ~n4094 & n7219 ) | ( ~n4094 & n8522 ) | ( n7219 & n8522 ) ;
  assign n8524 = n8523 ^ n7997 ^ 1'b0 ;
  assign n8525 = n6681 & n8524 ;
  assign n8526 = n6155 | n7391 ;
  assign n8527 = n5818 & ~n6576 ;
  assign n8528 = n2960 ^ n725 ^ 1'b0 ;
  assign n8529 = ~n4094 & n8528 ;
  assign n8531 = n5002 ^ n3080 ^ 1'b0 ;
  assign n8530 = n4575 & n7875 ;
  assign n8532 = n8531 ^ n8530 ^ 1'b0 ;
  assign n8533 = n395 | n2367 ;
  assign n8534 = n8533 ^ n560 ^ 1'b0 ;
  assign n8535 = ~n5016 & n8534 ;
  assign n8536 = n1930 & n8535 ;
  assign n8537 = ~n1143 & n1915 ;
  assign n8538 = n4081 & n8537 ;
  assign n8539 = n8538 ^ n386 ^ 1'b0 ;
  assign n8540 = ~n3035 & n8539 ;
  assign n8541 = ~n6450 & n8540 ;
  assign n8542 = n3631 & n8541 ;
  assign n8543 = n6576 | n7933 ;
  assign n8544 = ~n2989 & n7097 ;
  assign n8545 = n3270 & n8544 ;
  assign n8546 = n2673 | n8545 ;
  assign n8547 = n1300 | n8546 ;
  assign n8548 = n3277 | n5974 ;
  assign n8549 = n5976 ^ n1853 ^ 1'b0 ;
  assign n8550 = n1262 & n6223 ;
  assign n8551 = ( ~n5101 & n8549 ) | ( ~n5101 & n8550 ) | ( n8549 & n8550 ) ;
  assign n8552 = n5736 & ~n7490 ;
  assign n8553 = n6206 | n7729 ;
  assign n8554 = n4677 & ~n6411 ;
  assign n8555 = n7427 ^ n6569 ^ n2831 ;
  assign n8556 = n1884 & n3668 ;
  assign n8557 = n8556 ^ n6903 ^ 1'b0 ;
  assign n8558 = n2211 & ~n8557 ;
  assign n8559 = n7812 & n8558 ;
  assign n8560 = n441 & ~n802 ;
  assign n8561 = n8560 ^ n972 ^ 1'b0 ;
  assign n8562 = ~n8559 & n8561 ;
  assign n8563 = n1192 & ~n8562 ;
  assign n8564 = ~n1138 & n3186 ;
  assign n8565 = ~n4579 & n8564 ;
  assign n8566 = ( n456 & n726 ) | ( n456 & ~n5284 ) | ( n726 & ~n5284 ) ;
  assign n8567 = n2976 ^ n2273 ^ 1'b0 ;
  assign n8568 = n8567 ^ n5326 ^ 1'b0 ;
  assign n8569 = n3172 ^ n2789 ^ 1'b0 ;
  assign n8570 = n1345 & n8569 ;
  assign n8571 = ~n1161 & n8570 ;
  assign n8572 = ~n4646 & n8571 ;
  assign n8573 = n8572 ^ n6079 ^ n983 ;
  assign n8574 = n1544 & n1770 ;
  assign n8575 = n3146 & ~n5469 ;
  assign n8576 = n8575 ^ n4400 ^ 1'b0 ;
  assign n8577 = n8576 ^ n5721 ^ n1326 ;
  assign n8578 = n8574 & ~n8577 ;
  assign n8579 = ~n3655 & n8233 ;
  assign n8580 = n8579 ^ n4687 ^ 1'b0 ;
  assign n8581 = n2173 & ~n2549 ;
  assign n8582 = n7443 & n8581 ;
  assign n8583 = n8580 | n8582 ;
  assign n8584 = n8578 | n8583 ;
  assign n8585 = n3264 ^ n1568 ^ 1'b0 ;
  assign n8586 = n2854 & ~n8585 ;
  assign n8587 = n7016 & n8586 ;
  assign n8588 = n4293 & n8587 ;
  assign n8589 = n325 & ~n8588 ;
  assign n8590 = n1251 & ~n1639 ;
  assign n8591 = n8590 ^ n3770 ^ 1'b0 ;
  assign n8592 = n2275 | n8591 ;
  assign n8593 = n3210 | n6089 ;
  assign n8594 = n8593 ^ n6559 ^ 1'b0 ;
  assign n8595 = n1811 & ~n8396 ;
  assign n8596 = n1798 & ~n3619 ;
  assign n8597 = n4551 ^ n3379 ^ 1'b0 ;
  assign n8598 = n1897 | n8597 ;
  assign n8599 = n8596 & ~n8598 ;
  assign n8600 = n4276 & n5031 ;
  assign n8601 = ~n2359 & n2653 ;
  assign n8602 = ~n8497 & n8601 ;
  assign n8603 = n8602 ^ n3758 ^ 1'b0 ;
  assign n8604 = n6768 ^ n1566 ^ 1'b0 ;
  assign n8605 = n4402 ^ n4151 ^ 1'b0 ;
  assign n8606 = n8604 | n8605 ;
  assign n8607 = n8606 ^ n459 ^ 1'b0 ;
  assign n8608 = ~n3298 & n5001 ;
  assign n8609 = n5452 ^ n2365 ^ 1'b0 ;
  assign n8610 = n8608 & n8609 ;
  assign n8611 = n536 | n8610 ;
  assign n8612 = n6048 | n6238 ;
  assign n8613 = n8612 ^ n6647 ^ 1'b0 ;
  assign n8614 = n3488 ^ n3072 ^ 1'b0 ;
  assign n8615 = n4419 ^ n2266 ^ 1'b0 ;
  assign n8616 = ~n1300 & n5833 ;
  assign n8617 = n8616 ^ n3160 ^ 1'b0 ;
  assign n8618 = ~n8615 & n8617 ;
  assign n8619 = n1347 ^ n1141 ^ 1'b0 ;
  assign n8620 = n8619 ^ n6732 ^ 1'b0 ;
  assign n8621 = n8327 ^ n8018 ^ 1'b0 ;
  assign n8622 = n4884 ^ n2387 ^ 1'b0 ;
  assign n8623 = ~n2197 & n8622 ;
  assign n8624 = n8623 ^ n2190 ^ 1'b0 ;
  assign n8627 = n2570 | n5154 ;
  assign n8628 = n8627 ^ n5377 ^ 1'b0 ;
  assign n8625 = n8385 ^ n4537 ^ 1'b0 ;
  assign n8626 = ~n4698 & n8625 ;
  assign n8629 = n8628 ^ n8626 ^ 1'b0 ;
  assign n8630 = n4850 | n8287 ;
  assign n8631 = n6233 & ~n8630 ;
  assign n8632 = n2267 ^ n1832 ^ 1'b0 ;
  assign n8633 = n1877 & n8632 ;
  assign n8634 = n1560 ^ n433 ^ 1'b0 ;
  assign n8635 = ~n8633 & n8634 ;
  assign n8636 = n2662 & n8635 ;
  assign n8637 = n8636 ^ n6408 ^ 1'b0 ;
  assign n8638 = n2944 & n4100 ;
  assign n8639 = n8638 ^ n4849 ^ 1'b0 ;
  assign n8640 = n1331 | n8639 ;
  assign n8642 = n113 & ~n4149 ;
  assign n8643 = n8642 ^ n33 ^ 1'b0 ;
  assign n8641 = ~n1598 & n3891 ;
  assign n8644 = n8643 ^ n8641 ^ 1'b0 ;
  assign n8645 = n8644 ^ n8058 ^ 1'b0 ;
  assign n8646 = ( n2763 & ~n7236 ) | ( n2763 & n8645 ) | ( ~n7236 & n8645 ) ;
  assign n8647 = n2994 ^ n1235 ^ 1'b0 ;
  assign n8648 = n8647 ^ n488 ^ 1'b0 ;
  assign n8649 = n8648 ^ n857 ^ 1'b0 ;
  assign n8650 = n5432 & n8649 ;
  assign n8653 = n3424 ^ n1838 ^ n251 ;
  assign n8654 = n2623 | n4852 ;
  assign n8655 = n8653 & ~n8654 ;
  assign n8651 = n3838 & ~n5330 ;
  assign n8652 = n8651 ^ n3833 ^ 1'b0 ;
  assign n8656 = n8655 ^ n8652 ^ n3298 ;
  assign n8657 = n5083 ^ n369 ^ 1'b0 ;
  assign n8658 = n1190 & ~n8657 ;
  assign n8659 = ( n356 & n840 ) | ( n356 & n8055 ) | ( n840 & n8055 ) ;
  assign n8660 = n8659 ^ n7771 ^ 1'b0 ;
  assign n8661 = n8660 ^ n2138 ^ n1063 ;
  assign n8662 = ( n4489 & ~n8658 ) | ( n4489 & n8661 ) | ( ~n8658 & n8661 ) ;
  assign n8663 = n3052 & n8662 ;
  assign n8664 = n7054 ^ n2273 ^ 1'b0 ;
  assign n8665 = n6911 & ~n8664 ;
  assign n8666 = n2225 | n3574 ;
  assign n8667 = n7907 | n8666 ;
  assign n8668 = n4463 | n6196 ;
  assign n8669 = n8668 ^ n5690 ^ 1'b0 ;
  assign n8670 = ~n3033 & n8669 ;
  assign n8671 = n2218 & n8670 ;
  assign n8672 = n8671 ^ n6966 ^ 1'b0 ;
  assign n8673 = ~n3345 & n3660 ;
  assign n8674 = ~n6563 & n8673 ;
  assign n8675 = n2029 | n8674 ;
  assign n8676 = ~n43 & n2127 ;
  assign n8677 = ~n8049 & n8676 ;
  assign n8680 = n188 & ~n2616 ;
  assign n8678 = n4017 ^ n2914 ^ 1'b0 ;
  assign n8679 = n5806 | n8678 ;
  assign n8681 = n8680 ^ n8679 ^ n3745 ;
  assign n8683 = n551 & ~n6006 ;
  assign n8682 = n704 & ~n7280 ;
  assign n8684 = n8683 ^ n8682 ^ 1'b0 ;
  assign n8685 = n4229 & ~n7078 ;
  assign n8686 = n1096 | n8685 ;
  assign n8687 = ~n414 & n2290 ;
  assign n8688 = ~n3504 & n8687 ;
  assign n8689 = n2822 | n4975 ;
  assign n8692 = n579 & ~n1029 ;
  assign n8693 = n8692 ^ n304 ^ 1'b0 ;
  assign n8690 = n4478 | n5973 ;
  assign n8691 = n140 & ~n8690 ;
  assign n8694 = n8693 ^ n8691 ^ 1'b0 ;
  assign n8695 = n8694 ^ n4386 ^ 1'b0 ;
  assign n8696 = n2022 | n8695 ;
  assign n8697 = n8689 | n8696 ;
  assign n8700 = n968 & n4751 ;
  assign n8701 = n5163 ^ n2226 ^ 1'b0 ;
  assign n8702 = n8700 | n8701 ;
  assign n8703 = n3324 | n8702 ;
  assign n8698 = ~n401 & n2537 ;
  assign n8699 = n5982 & n8698 ;
  assign n8704 = n8703 ^ n8699 ^ 1'b0 ;
  assign n8705 = ~n2073 & n8328 ;
  assign n8706 = ~n3418 & n8204 ;
  assign n8707 = ~n262 & n4635 ;
  assign n8708 = n8706 & n8707 ;
  assign n8709 = n4442 | n4666 ;
  assign n8710 = n5814 & ~n8709 ;
  assign n8711 = n2806 & n4007 ;
  assign n8712 = ~n6759 & n8711 ;
  assign n8713 = n2925 & ~n5217 ;
  assign n8714 = n6947 & n8713 ;
  assign n8715 = n3085 & ~n8714 ;
  assign n8716 = ~n5293 & n5454 ;
  assign n8717 = n5554 ^ n854 ^ 1'b0 ;
  assign n8718 = ~n287 & n3851 ;
  assign n8719 = n1055 & n8718 ;
  assign n8720 = n4616 & ~n8719 ;
  assign n8721 = n2445 & n7467 ;
  assign n8722 = n5473 | n5757 ;
  assign n8723 = n617 & ~n8722 ;
  assign n8724 = ~n982 & n8723 ;
  assign n8725 = n2083 | n2139 ;
  assign n8726 = n8725 ^ n48 ^ 1'b0 ;
  assign n8727 = n8724 & n8726 ;
  assign n8728 = n2918 ^ n425 ^ 1'b0 ;
  assign n8730 = n1745 ^ n1016 ^ 1'b0 ;
  assign n8731 = ~n8122 & n8730 ;
  assign n8729 = n1715 & ~n4131 ;
  assign n8732 = n8731 ^ n8729 ^ 1'b0 ;
  assign n8733 = ~n8728 & n8732 ;
  assign n8734 = ~n1392 & n8733 ;
  assign n8735 = n6238 ^ n2780 ^ 1'b0 ;
  assign n8736 = n5123 & n5168 ;
  assign n8737 = n8736 ^ n5186 ^ 1'b0 ;
  assign n8738 = n2652 ^ n2446 ^ 1'b0 ;
  assign n8739 = n3536 ^ n2376 ^ 1'b0 ;
  assign n8740 = n8738 & ~n8739 ;
  assign n8741 = ~n2879 & n8740 ;
  assign n8742 = n3166 ^ n1155 ^ 1'b0 ;
  assign n8743 = n5246 | n8742 ;
  assign n8744 = n5151 & ~n8743 ;
  assign n8745 = n8744 ^ n4931 ^ 1'b0 ;
  assign n8746 = ~n2210 & n8745 ;
  assign n8747 = n8746 ^ n5388 ^ 1'b0 ;
  assign n8748 = n7556 ^ n6914 ^ 1'b0 ;
  assign n8749 = n2727 & n8748 ;
  assign n8750 = n8639 ^ n2924 ^ 1'b0 ;
  assign n8751 = ( n2277 & ~n4770 ) | ( n2277 & n6112 ) | ( ~n4770 & n6112 ) ;
  assign n8752 = n3936 ^ n3238 ^ n205 ;
  assign n8753 = n8752 ^ n6574 ^ 1'b0 ;
  assign n8754 = n8751 & n8753 ;
  assign n8756 = n833 & ~n1313 ;
  assign n8755 = n1464 & n4960 ;
  assign n8757 = n8756 ^ n8755 ^ 1'b0 ;
  assign n8758 = n5061 & n8757 ;
  assign n8759 = n1886 & ~n3680 ;
  assign n8760 = n835 & n1635 ;
  assign n8761 = ~n7589 & n8760 ;
  assign n8762 = n7377 ^ n5936 ^ 1'b0 ;
  assign n8763 = n8761 & ~n8762 ;
  assign n8764 = n7530 ^ n2446 ^ n150 ;
  assign n8765 = n8764 ^ n4321 ^ 1'b0 ;
  assign n8766 = n7022 & ~n8765 ;
  assign n8772 = ~n257 & n5769 ;
  assign n8773 = n8772 ^ n7109 ^ 1'b0 ;
  assign n8771 = n2850 & ~n4813 ;
  assign n8767 = n2260 ^ n331 ^ 1'b0 ;
  assign n8768 = n3827 & n8767 ;
  assign n8769 = ~n3096 & n8768 ;
  assign n8770 = n8769 ^ n6881 ^ 1'b0 ;
  assign n8774 = n8773 ^ n8771 ^ n8770 ;
  assign n8778 = n1365 & n3314 ;
  assign n8779 = n8778 ^ n2146 ^ x0 ;
  assign n8776 = n63 & n1353 ;
  assign n8775 = n398 & n7867 ;
  assign n8777 = n8776 ^ n8775 ^ 1'b0 ;
  assign n8780 = n8779 ^ n8777 ^ 1'b0 ;
  assign n8781 = n8061 & n8780 ;
  assign n8782 = n3389 ^ n2855 ^ n582 ;
  assign n8783 = n3990 ^ n2484 ^ 1'b0 ;
  assign n8784 = ~n7849 & n8783 ;
  assign n8787 = ~n2204 & n3428 ;
  assign n8785 = n6997 ^ n2244 ^ 1'b0 ;
  assign n8786 = n277 & ~n8785 ;
  assign n8788 = n8787 ^ n8786 ^ 1'b0 ;
  assign n8789 = n5526 & ~n7792 ;
  assign n8790 = ~n3255 & n6607 ;
  assign n8791 = n2624 & ~n4374 ;
  assign n8792 = n2178 & n8791 ;
  assign n8793 = n746 & n8792 ;
  assign n8794 = n1825 ^ n875 ^ 1'b0 ;
  assign n8795 = ~n8793 & n8794 ;
  assign n8796 = n8795 ^ n8494 ^ 1'b0 ;
  assign n8797 = n8790 & n8796 ;
  assign n8798 = n6193 ^ n4324 ^ 1'b0 ;
  assign n8799 = n4764 ^ n422 ^ 1'b0 ;
  assign n8800 = n2535 | n8799 ;
  assign n8801 = n3417 & ~n8800 ;
  assign n8802 = ( n5918 & n8330 ) | ( n5918 & n8801 ) | ( n8330 & n8801 ) ;
  assign n8803 = n1818 ^ n205 ^ 1'b0 ;
  assign n8804 = n322 & n477 ;
  assign n8805 = n8803 & n8804 ;
  assign n8806 = n8805 ^ n5861 ^ 1'b0 ;
  assign n8807 = n4024 | n7756 ;
  assign n8811 = ( n2429 & n2686 ) | ( n2429 & ~n4740 ) | ( n2686 & ~n4740 ) ;
  assign n8808 = n7628 ^ n2754 ^ 1'b0 ;
  assign n8809 = ~n125 & n8808 ;
  assign n8810 = n5990 & n8809 ;
  assign n8812 = n8811 ^ n8810 ^ 1'b0 ;
  assign n8813 = x9 & n152 ;
  assign n8814 = n8813 ^ n49 ^ 1'b0 ;
  assign n8815 = n8814 ^ n4720 ^ 1'b0 ;
  assign n8816 = ~n6846 & n8815 ;
  assign n8817 = n8816 ^ n5803 ^ 1'b0 ;
  assign n8818 = n1329 & n2113 ;
  assign n8819 = ~n2248 & n8818 ;
  assign n8820 = n8819 ^ n451 ^ 1'b0 ;
  assign n8821 = n2772 ^ n1445 ^ n1164 ;
  assign n8822 = ~n135 & n8821 ;
  assign n8823 = n8820 & n8822 ;
  assign n8824 = n6000 ^ n3790 ^ 1'b0 ;
  assign n8825 = n2039 ^ n1560 ^ 1'b0 ;
  assign n8826 = n8825 ^ n7672 ^ n623 ;
  assign n8827 = n1307 ^ n459 ^ 1'b0 ;
  assign n8828 = n3828 & ~n8827 ;
  assign n8829 = n8828 ^ n2451 ^ 1'b0 ;
  assign n8830 = ~n4427 & n8829 ;
  assign n8831 = n4519 ^ n3245 ^ n1637 ;
  assign n8832 = n8831 ^ n5229 ^ 1'b0 ;
  assign n8833 = ~n5555 & n8832 ;
  assign n8834 = n8833 ^ n861 ^ 1'b0 ;
  assign n8835 = n7124 ^ n1962 ^ 1'b0 ;
  assign n8836 = n5547 & n8835 ;
  assign n8837 = n3333 ^ n552 ^ 1'b0 ;
  assign n8838 = n3414 | n8837 ;
  assign n8839 = n1778 ^ n503 ^ 1'b0 ;
  assign n8840 = ~n1848 & n8839 ;
  assign n8841 = n8840 ^ n4578 ^ 1'b0 ;
  assign n8842 = n8841 ^ n8259 ^ n6891 ;
  assign n8843 = ( n17 & n2125 ) | ( n17 & ~n8109 ) | ( n2125 & ~n8109 ) ;
  assign n8844 = n8843 ^ n8715 ^ n905 ;
  assign n8845 = n3418 & ~n7605 ;
  assign n8846 = ~n714 & n3350 ;
  assign n8847 = n2648 & n8846 ;
  assign n8848 = n1128 & n1941 ;
  assign n8849 = n8847 & n8848 ;
  assign n8850 = n2940 | n8849 ;
  assign n8851 = n1723 & ~n3843 ;
  assign n8852 = n956 & n8851 ;
  assign n8853 = n8852 ^ n1497 ^ 1'b0 ;
  assign n8858 = n6028 ^ n2983 ^ 1'b0 ;
  assign n8854 = n1365 ^ n1023 ^ 1'b0 ;
  assign n8855 = n4702 & ~n8854 ;
  assign n8856 = n6067 & n8855 ;
  assign n8857 = n8856 ^ n3795 ^ 1'b0 ;
  assign n8859 = n8858 ^ n8857 ^ 1'b0 ;
  assign n8860 = n8853 & ~n8859 ;
  assign n8861 = n1944 & n2104 ;
  assign n8862 = ~n2087 & n8861 ;
  assign n8866 = ~n3160 & n3232 ;
  assign n8867 = n8866 ^ n1684 ^ 1'b0 ;
  assign n8864 = n4632 & ~n4785 ;
  assign n8865 = ~n3880 & n8864 ;
  assign n8868 = n8867 ^ n8865 ^ n2377 ;
  assign n8863 = n2808 & n3444 ;
  assign n8869 = n8868 ^ n8863 ^ n360 ;
  assign n8870 = n1898 | n8869 ;
  assign n8871 = n4345 & n8870 ;
  assign n8872 = n4091 & ~n8073 ;
  assign n8873 = n8872 ^ n214 ^ 1'b0 ;
  assign n8874 = n5124 ^ n4121 ^ n983 ;
  assign n8875 = ~n8873 & n8874 ;
  assign n8876 = n8875 ^ n1854 ^ 1'b0 ;
  assign n8877 = n60 | n1592 ;
  assign n8878 = n8877 ^ n3080 ^ 1'b0 ;
  assign n8879 = n208 | n489 ;
  assign n8881 = n431 & n2421 ;
  assign n8880 = n1539 & n1789 ;
  assign n8882 = n8881 ^ n8880 ^ 1'b0 ;
  assign n8883 = n8879 & n8882 ;
  assign n8884 = n1933 ^ n223 ^ 1'b0 ;
  assign n8885 = n146 | n3152 ;
  assign n8886 = n8885 ^ n5880 ^ n1993 ;
  assign n8887 = n8430 ^ n448 ^ 1'b0 ;
  assign n8888 = ~n8319 & n8887 ;
  assign n8889 = ~n7599 & n8888 ;
  assign n8890 = n8889 ^ n2755 ^ 1'b0 ;
  assign n8891 = n2946 | n8890 ;
  assign n8892 = n1286 | n7051 ;
  assign n8893 = n8892 ^ n7804 ^ 1'b0 ;
  assign n8894 = n1307 & n1389 ;
  assign n8895 = n4381 | n8894 ;
  assign n8896 = n8895 ^ n2238 ^ 1'b0 ;
  assign n8897 = n6161 & ~n8896 ;
  assign n8898 = n2937 & n8897 ;
  assign n8899 = ~n474 & n4039 ;
  assign n8900 = n8899 ^ n1765 ^ 1'b0 ;
  assign n8901 = n525 & ~n8900 ;
  assign n8902 = ~n5122 & n8901 ;
  assign n8903 = n4643 & n8902 ;
  assign n8904 = n1327 & n8506 ;
  assign n8905 = n6325 & n8904 ;
  assign n8906 = n304 & ~n850 ;
  assign n8907 = ~n2361 & n7798 ;
  assign n8908 = n279 & n2658 ;
  assign n8911 = n4222 ^ n1078 ^ 1'b0 ;
  assign n8909 = n395 | n7018 ;
  assign n8910 = n8909 ^ n4976 ^ 1'b0 ;
  assign n8912 = n8911 ^ n8910 ^ 1'b0 ;
  assign n8913 = n8908 & ~n8912 ;
  assign n8914 = n2204 | n5468 ;
  assign n8915 = n8914 ^ n4376 ^ 1'b0 ;
  assign n8916 = n8915 ^ n4755 ^ 1'b0 ;
  assign n8917 = n8916 ^ n3080 ^ 1'b0 ;
  assign n8918 = n8917 ^ n1871 ^ 1'b0 ;
  assign n8919 = n3143 ^ n115 ^ 1'b0 ;
  assign n8920 = n7981 ^ n1534 ^ 1'b0 ;
  assign n8921 = n2812 ^ n875 ^ 1'b0 ;
  assign n8922 = n3335 | n8921 ;
  assign n8923 = n8922 ^ n505 ^ 1'b0 ;
  assign n8924 = n3881 & ~n8923 ;
  assign n8931 = n1092 & n2326 ;
  assign n8932 = n13 | n8931 ;
  assign n8933 = n163 | n8932 ;
  assign n8925 = n3971 ^ n1271 ^ 1'b0 ;
  assign n8926 = n401 & n8925 ;
  assign n8927 = n8926 ^ n1465 ^ n1462 ;
  assign n8928 = n5828 ^ n2701 ^ n1276 ;
  assign n8929 = ~n1880 & n8928 ;
  assign n8930 = ~n8927 & n8929 ;
  assign n8934 = n8933 ^ n8930 ^ 1'b0 ;
  assign n8935 = n2614 & n3935 ;
  assign n8936 = ~n5324 & n8935 ;
  assign n8937 = n667 & ~n8936 ;
  assign n8938 = n4187 ^ n3252 ^ 1'b0 ;
  assign n8939 = n1816 | n8938 ;
  assign n8940 = n1217 & ~n2523 ;
  assign n8941 = ~n5954 & n8940 ;
  assign n8942 = n8939 & n8941 ;
  assign n8943 = n8942 ^ n8083 ^ 1'b0 ;
  assign n8944 = n7992 ^ n4278 ^ 1'b0 ;
  assign n8945 = n8944 ^ n3176 ^ 1'b0 ;
  assign n8946 = ~n2669 & n8874 ;
  assign n8947 = n1198 | n1418 ;
  assign n8948 = n8947 ^ n6110 ^ 1'b0 ;
  assign n8949 = n3135 | n8948 ;
  assign n8950 = n7360 & ~n8949 ;
  assign n8951 = n5535 ^ n2547 ^ 1'b0 ;
  assign n8952 = ~n5072 & n6978 ;
  assign n8953 = n5289 ^ n1349 ^ 1'b0 ;
  assign n8954 = ~n2920 & n8953 ;
  assign n8955 = n302 | n7837 ;
  assign n8956 = n8955 ^ n8376 ^ 1'b0 ;
  assign n8957 = n2152 & ~n8956 ;
  assign n8958 = n1111 | n5244 ;
  assign n8959 = ~n627 & n4275 ;
  assign n8960 = n3686 ^ n3308 ^ 1'b0 ;
  assign n8961 = n8960 ^ n6713 ^ 1'b0 ;
  assign n8962 = n8961 ^ n2594 ^ 1'b0 ;
  assign n8963 = n2902 | n6342 ;
  assign n8964 = n4576 ^ n3287 ^ 1'b0 ;
  assign n8965 = n5138 & ~n8964 ;
  assign n8967 = n2474 ^ n1753 ^ 1'b0 ;
  assign n8966 = n3361 ^ n1337 ^ 1'b0 ;
  assign n8968 = n8967 ^ n8966 ^ 1'b0 ;
  assign n8969 = ~n7155 & n8968 ;
  assign n8970 = n8969 ^ n1425 ^ 1'b0 ;
  assign n8971 = ( n1618 & ~n5216 ) | ( n1618 & n8970 ) | ( ~n5216 & n8970 ) ;
  assign n8972 = n1701 & ~n8634 ;
  assign n8973 = n7922 ^ n5212 ^ 1'b0 ;
  assign n8974 = n8973 ^ n6216 ^ n1586 ;
  assign n8975 = n1055 | n2242 ;
  assign n8976 = n8975 ^ n5759 ^ 1'b0 ;
  assign n8977 = n8976 ^ n4438 ^ 1'b0 ;
  assign n8978 = ~n3725 & n8559 ;
  assign n8979 = n835 & ~n5719 ;
  assign n8980 = n8979 ^ n6200 ^ 1'b0 ;
  assign n8981 = n5235 & ~n8448 ;
  assign n8982 = n1038 & n2261 ;
  assign n8983 = ~n1219 & n8982 ;
  assign n8984 = ~n2548 & n2609 ;
  assign n8985 = n8984 ^ n2217 ^ 1'b0 ;
  assign n8986 = ( ~n347 & n8983 ) | ( ~n347 & n8985 ) | ( n8983 & n8985 ) ;
  assign n8987 = n5865 & n8986 ;
  assign n8988 = n1868 & ~n8987 ;
  assign n8989 = ~n5809 & n8988 ;
  assign n8990 = n3591 & ~n8989 ;
  assign n8991 = n8990 ^ n6663 ^ 1'b0 ;
  assign n8992 = n3839 ^ n586 ^ 1'b0 ;
  assign n8993 = n8992 ^ n4561 ^ 1'b0 ;
  assign n8994 = ~n445 & n2130 ;
  assign n8995 = ~n292 & n8994 ;
  assign n8996 = n8995 ^ n6187 ^ 1'b0 ;
  assign n8997 = ~n8468 & n8996 ;
  assign n8998 = ( n2206 & ~n5970 ) | ( n2206 & n7278 ) | ( ~n5970 & n7278 ) ;
  assign n8999 = n2272 & n2932 ;
  assign n9000 = n8999 ^ n3095 ^ 1'b0 ;
  assign n9001 = n3193 ^ n2639 ^ 1'b0 ;
  assign n9002 = n1132 & ~n9001 ;
  assign n9003 = n3145 & n3504 ;
  assign n9004 = ~n6756 & n9003 ;
  assign n9005 = n4435 & ~n9004 ;
  assign n9006 = ~n9002 & n9005 ;
  assign n9007 = n7989 & ~n8266 ;
  assign n9008 = n1182 & n9007 ;
  assign n9009 = n1411 & ~n7627 ;
  assign n9010 = ~n112 & n2432 ;
  assign n9011 = n841 & ~n8254 ;
  assign n9012 = n9011 ^ n2952 ^ 1'b0 ;
  assign n9013 = n9010 & ~n9012 ;
  assign n9014 = n3520 & n9013 ;
  assign n9016 = n270 & n564 ;
  assign n9017 = n9016 ^ n6892 ^ 1'b0 ;
  assign n9015 = n6870 | n8700 ;
  assign n9018 = n9017 ^ n9015 ^ 1'b0 ;
  assign n9019 = n344 & ~n8598 ;
  assign n9020 = ~n6104 & n9019 ;
  assign n9021 = n9020 ^ n7012 ^ 1'b0 ;
  assign n9022 = n2303 & n9021 ;
  assign n9023 = n6110 ^ n3623 ^ 1'b0 ;
  assign n9024 = n9023 ^ n3232 ^ 1'b0 ;
  assign n9025 = n3715 & ~n8024 ;
  assign n9026 = ~n6842 & n9025 ;
  assign n9027 = n9026 ^ n2986 ^ 1'b0 ;
  assign n9028 = n6516 | n9027 ;
  assign n9029 = n6491 & ~n9028 ;
  assign n9030 = ~n1745 & n5139 ;
  assign n9031 = n6015 ^ n3293 ^ 1'b0 ;
  assign n9032 = ( n4034 & n4667 ) | ( n4034 & n7534 ) | ( n4667 & n7534 ) ;
  assign n9033 = n7806 & n9032 ;
  assign n9034 = ~n750 & n1069 ;
  assign n9035 = ~n2315 & n9034 ;
  assign n9036 = n9035 ^ n7526 ^ 1'b0 ;
  assign n9037 = n6554 ^ n1284 ^ 1'b0 ;
  assign n9038 = n9037 ^ n7753 ^ n3116 ;
  assign n9039 = n4160 | n5227 ;
  assign n9040 = ~n5656 & n9039 ;
  assign n9041 = ~n8129 & n9040 ;
  assign n9042 = n8934 ^ n2677 ^ 1'b0 ;
  assign n9043 = ~n6355 & n9042 ;
  assign n9044 = n4091 ^ n749 ^ 1'b0 ;
  assign n9045 = n6037 ^ n2019 ^ 1'b0 ;
  assign n9046 = n9045 ^ n3643 ^ n468 ;
  assign n9047 = ~n150 & n1065 ;
  assign n9048 = n3125 ^ n798 ^ 1'b0 ;
  assign n9049 = n7526 ^ n2384 ^ 1'b0 ;
  assign n9050 = n52 & ~n5756 ;
  assign n9051 = n9049 & n9050 ;
  assign n9052 = n8995 ^ n3552 ^ 1'b0 ;
  assign n9053 = ~n7897 & n9052 ;
  assign n9057 = n1241 ^ n790 ^ 1'b0 ;
  assign n9056 = n5240 ^ n3472 ^ 1'b0 ;
  assign n9054 = n734 ^ n188 ^ 1'b0 ;
  assign n9055 = n3715 & ~n9054 ;
  assign n9058 = n9057 ^ n9056 ^ n9055 ;
  assign n9059 = n6080 | n7778 ;
  assign n9060 = n205 | n5724 ;
  assign n9061 = n6000 & n8423 ;
  assign n9062 = n9061 ^ n4117 ^ 1'b0 ;
  assign n9063 = n2264 & n6903 ;
  assign n9064 = n7416 ^ n1938 ^ 1'b0 ;
  assign n9065 = n9063 & ~n9064 ;
  assign n9068 = n8399 ^ n1631 ^ 1'b0 ;
  assign n9066 = n1516 & n2159 ;
  assign n9067 = n9066 ^ n592 ^ 1'b0 ;
  assign n9069 = n9068 ^ n9067 ^ 1'b0 ;
  assign n9070 = ~n1574 & n6230 ;
  assign n9071 = n7931 ^ n607 ^ 1'b0 ;
  assign n9072 = n9071 ^ n694 ^ 1'b0 ;
  assign n9073 = n9072 ^ n4327 ^ 1'b0 ;
  assign n9074 = n6542 | n9073 ;
  assign n9075 = n4990 | n8243 ;
  assign n9076 = n6925 | n9075 ;
  assign n9077 = n3437 ^ n2002 ^ n1031 ;
  assign n9078 = n4086 ^ n1154 ^ 1'b0 ;
  assign n9079 = n4293 ^ n4252 ^ 1'b0 ;
  assign n9080 = n9078 & ~n9079 ;
  assign n9081 = ~n5654 & n9080 ;
  assign n9082 = n9081 ^ n7121 ^ 1'b0 ;
  assign n9083 = n1300 & n9082 ;
  assign n9084 = ~n1639 & n3544 ;
  assign n9085 = n582 & ~n7633 ;
  assign n9086 = ~n5281 & n6227 ;
  assign n9087 = ~n150 & n733 ;
  assign n9088 = ~n1674 & n9087 ;
  assign n9089 = n7498 | n9088 ;
  assign n9090 = ( n588 & ~n659 ) | ( n588 & n765 ) | ( ~n659 & n765 ) ;
  assign n9091 = ~n4007 & n9090 ;
  assign n9092 = n2769 & n4121 ;
  assign n9093 = n6972 ^ n3199 ^ 1'b0 ;
  assign n9094 = ~n9092 & n9093 ;
  assign n9095 = n5325 ^ n94 ^ 1'b0 ;
  assign n9096 = n115 | n162 ;
  assign n9097 = n9096 ^ n7288 ^ 1'b0 ;
  assign n9098 = n732 | n9097 ;
  assign n9099 = ~n387 & n1351 ;
  assign n9100 = n9099 ^ n5652 ^ 1'b0 ;
  assign n9101 = n795 | n9100 ;
  assign n9102 = n901 | n9101 ;
  assign n9103 = ~n3674 & n9102 ;
  assign n9104 = n9103 ^ n831 ^ 1'b0 ;
  assign n9105 = n922 & ~n4819 ;
  assign n9106 = ~n9104 & n9105 ;
  assign n9107 = ~n5649 & n8186 ;
  assign n9110 = n2236 & n3357 ;
  assign n9108 = n6854 ^ n1363 ^ 1'b0 ;
  assign n9109 = n9108 ^ n4290 ^ 1'b0 ;
  assign n9111 = n9110 ^ n9109 ^ 1'b0 ;
  assign n9112 = n885 ^ n411 ^ 1'b0 ;
  assign n9113 = n845 & n9112 ;
  assign n9114 = n4457 | n9113 ;
  assign n9115 = n2900 & n4787 ;
  assign n9116 = n9115 ^ n2927 ^ 1'b0 ;
  assign n9117 = ~n4328 & n9116 ;
  assign n9118 = n8122 | n9117 ;
  assign n9119 = n9118 ^ n2455 ^ 1'b0 ;
  assign n9120 = ~n2751 & n9119 ;
  assign n9121 = n6172 ^ n3797 ^ 1'b0 ;
  assign n9122 = n9121 ^ n2837 ^ 1'b0 ;
  assign n9123 = ~n1533 & n9122 ;
  assign n9124 = ~n9120 & n9123 ;
  assign n9125 = n9114 & ~n9124 ;
  assign n9126 = n9125 ^ n950 ^ 1'b0 ;
  assign n9134 = n884 | n4655 ;
  assign n9127 = ~n3173 & n6719 ;
  assign n9128 = n9127 ^ n105 ^ 1'b0 ;
  assign n9129 = n6157 ^ n2806 ^ n2787 ;
  assign n9130 = n9128 | n9129 ;
  assign n9131 = n6084 & ~n9130 ;
  assign n9132 = n4405 | n9131 ;
  assign n9133 = n9132 ^ n1639 ^ 1'b0 ;
  assign n9135 = n9134 ^ n9133 ^ 1'b0 ;
  assign n9136 = n5136 & n7830 ;
  assign n9137 = ( n2574 & n6114 ) | ( n2574 & n9136 ) | ( n6114 & n9136 ) ;
  assign n9138 = n434 & ~n2379 ;
  assign n9139 = ~n2933 & n9138 ;
  assign n9140 = n9139 ^ n6649 ^ 1'b0 ;
  assign n9141 = n2106 & ~n2225 ;
  assign n9142 = n9141 ^ n8731 ^ 1'b0 ;
  assign n9143 = ~n2790 & n9142 ;
  assign n9144 = n6997 ^ n2637 ^ 1'b0 ;
  assign n9145 = n845 & ~n9144 ;
  assign n9146 = n9145 ^ n3556 ^ 1'b0 ;
  assign n9147 = n2886 ^ n1141 ^ 1'b0 ;
  assign n9148 = n9147 ^ n3881 ^ 1'b0 ;
  assign n9150 = n466 & n3487 ;
  assign n9149 = ~n288 & n1668 ;
  assign n9151 = n9150 ^ n9149 ^ 1'b0 ;
  assign n9152 = n1832 | n9151 ;
  assign n9153 = n28 & ~n9152 ;
  assign n9154 = n4326 ^ n612 ^ 1'b0 ;
  assign n9155 = ~n2463 & n9154 ;
  assign n9156 = ~n9153 & n9155 ;
  assign n9157 = n9156 ^ n1743 ^ 1'b0 ;
  assign n9158 = n129 & n9157 ;
  assign n9159 = n1516 & ~n2197 ;
  assign n9160 = n7170 ^ n3167 ^ 1'b0 ;
  assign n9161 = n2653 & ~n9160 ;
  assign n9162 = n1029 & n9161 ;
  assign n9163 = n9159 & n9162 ;
  assign n9164 = n9163 ^ n978 ^ 1'b0 ;
  assign n9165 = n9158 & n9164 ;
  assign n9166 = n1764 & ~n1789 ;
  assign n9167 = n9166 ^ n2715 ^ n1772 ;
  assign n9168 = n1670 & ~n9167 ;
  assign n9169 = n7153 & n9168 ;
  assign n9170 = n4976 ^ n2478 ^ 1'b0 ;
  assign n9171 = n3408 | n5420 ;
  assign n9172 = n6994 & ~n9171 ;
  assign n9173 = ~n9122 & n9172 ;
  assign n9174 = n3364 ^ n2324 ^ 1'b0 ;
  assign n9175 = n1461 | n9174 ;
  assign n9176 = n445 | n9175 ;
  assign n9177 = n9176 ^ n2811 ^ 1'b0 ;
  assign n9178 = n706 & ~n2409 ;
  assign n9179 = n1416 & ~n2137 ;
  assign n9180 = n9179 ^ n4040 ^ 1'b0 ;
  assign n9181 = n7127 ^ n4163 ^ 1'b0 ;
  assign n9182 = ~n1208 & n9181 ;
  assign n9183 = n1033 ^ n1032 ^ 1'b0 ;
  assign n9184 = n7889 | n9183 ;
  assign n9185 = n183 | n5874 ;
  assign n9186 = n9185 ^ n1077 ^ 1'b0 ;
  assign n9187 = n3482 ^ n631 ^ 1'b0 ;
  assign n9188 = n1114 ^ n508 ^ 1'b0 ;
  assign n9189 = n6059 | n9188 ;
  assign n9190 = n9187 | n9189 ;
  assign n9191 = ~n9186 & n9190 ;
  assign n9192 = n708 & ~n4505 ;
  assign n9193 = n3011 ^ n390 ^ n13 ;
  assign n9194 = ~n8197 & n9193 ;
  assign n9195 = n9194 ^ n326 ^ 1'b0 ;
  assign n9196 = n8708 ^ n1252 ^ 1'b0 ;
  assign n9197 = ~n322 & n2915 ;
  assign n9198 = n5811 & n9197 ;
  assign n9199 = n2545 & n9198 ;
  assign n9200 = n6463 | n9199 ;
  assign n9201 = n9200 ^ n5513 ^ 1'b0 ;
  assign n9202 = n1900 | n3610 ;
  assign n9203 = n49 & ~n9202 ;
  assign n9204 = ( n3423 & ~n3564 ) | ( n3423 & n4912 ) | ( ~n3564 & n4912 ) ;
  assign n9205 = ~n5641 & n9204 ;
  assign n9206 = ~n88 & n7126 ;
  assign n9207 = n9206 ^ n6108 ^ 1'b0 ;
  assign n9208 = ( n120 & n2206 ) | ( n120 & ~n3774 ) | ( n2206 & ~n3774 ) ;
  assign n9209 = n1798 & n3064 ;
  assign n9210 = n9209 ^ n3501 ^ n3098 ;
  assign n9211 = n1318 & n9210 ;
  assign n9212 = n360 & n9211 ;
  assign n9213 = n592 | n1705 ;
  assign n9214 = n7683 & n9213 ;
  assign n9215 = n9214 ^ n390 ^ 1'b0 ;
  assign n9216 = n7159 ^ n3974 ^ 1'b0 ;
  assign n9218 = n4650 & ~n6491 ;
  assign n9219 = n9218 ^ n3676 ^ 1'b0 ;
  assign n9217 = n997 | n6256 ;
  assign n9220 = n9219 ^ n9217 ^ 1'b0 ;
  assign n9221 = n33 | n4294 ;
  assign n9222 = n6589 & ~n9221 ;
  assign n9223 = n9222 ^ n2637 ^ n1363 ;
  assign n9224 = ~n593 & n9223 ;
  assign n9225 = ~n7727 & n9224 ;
  assign n9226 = n2103 | n8395 ;
  assign n9227 = ~n3080 & n9226 ;
  assign n9228 = n2595 & n8608 ;
  assign n9229 = ~n3125 & n9228 ;
  assign n9230 = n1234 & n5213 ;
  assign n9231 = n9229 & n9230 ;
  assign n9232 = n2874 & n9231 ;
  assign n9235 = n644 & n6248 ;
  assign n9236 = n6934 & n8764 ;
  assign n9237 = ~n9235 & n9236 ;
  assign n9233 = ( n1900 & ~n4072 ) | ( n1900 & n6452 ) | ( ~n4072 & n6452 ) ;
  assign n9234 = n105 & n9233 ;
  assign n9238 = n9237 ^ n9234 ^ 1'b0 ;
  assign n9239 = n3530 | n4162 ;
  assign n9240 = n2185 ^ n2007 ^ 1'b0 ;
  assign n9241 = n9240 ^ n5864 ^ n841 ;
  assign n9242 = n7979 ^ n2807 ^ n390 ;
  assign n9243 = n1117 & n9242 ;
  assign n9244 = n5417 & n9243 ;
  assign n9245 = n7109 ^ n1534 ^ 1'b0 ;
  assign n9246 = ~n2894 & n2895 ;
  assign n9247 = n9246 ^ n177 ^ 1'b0 ;
  assign n9248 = n9247 ^ n3646 ^ n1161 ;
  assign n9249 = n3050 | n9248 ;
  assign n9250 = n6666 & ~n9249 ;
  assign n9251 = n605 & n754 ;
  assign n9252 = n2246 & ~n4573 ;
  assign n9253 = n676 & ~n9252 ;
  assign n9254 = ~n5086 & n7206 ;
  assign n9255 = n4925 & n8233 ;
  assign n9256 = n9255 ^ n7829 ^ 1'b0 ;
  assign n9257 = n6950 & ~n7897 ;
  assign n9258 = ~n1408 & n9257 ;
  assign n9259 = n61 | n2781 ;
  assign n9260 = n9259 ^ n551 ^ 1'b0 ;
  assign n9261 = ~n3262 & n3613 ;
  assign n9262 = n7119 ^ n4409 ^ 1'b0 ;
  assign n9263 = n9261 & n9262 ;
  assign n9264 = n3440 ^ n3223 ^ 1'b0 ;
  assign n9265 = n9264 ^ n729 ^ 1'b0 ;
  assign n9266 = n6751 | n9265 ;
  assign n9267 = n8685 ^ n8506 ^ 1'b0 ;
  assign n9268 = n8588 ^ n5711 ^ n5292 ;
  assign n9269 = n2968 ^ n776 ^ 1'b0 ;
  assign n9272 = n3314 ^ n2533 ^ n19 ;
  assign n9270 = n7881 ^ n582 ^ 1'b0 ;
  assign n9271 = n9270 ^ n6227 ^ 1'b0 ;
  assign n9273 = n9272 ^ n9271 ^ n3633 ;
  assign n9274 = n1839 | n3736 ;
  assign n9275 = n2265 | n9274 ;
  assign n9276 = n2569 | n9275 ;
  assign n9277 = n7757 ^ n4407 ^ 1'b0 ;
  assign n9278 = n996 & n4913 ;
  assign n9279 = n9278 ^ n4583 ^ 1'b0 ;
  assign n9280 = n8976 & ~n9279 ;
  assign n9281 = n9277 | n9280 ;
  assign n9282 = n4420 & ~n9281 ;
  assign n9283 = n8570 ^ n4782 ^ 1'b0 ;
  assign n9284 = n4581 | n9283 ;
  assign n9285 = n74 & ~n6722 ;
  assign n9286 = ~n1336 & n9285 ;
  assign n9287 = n9286 ^ n4278 ^ n3143 ;
  assign n9288 = n1969 & ~n3390 ;
  assign n9289 = n841 & n7766 ;
  assign n9290 = n805 | n9289 ;
  assign n9291 = n4058 ^ n1087 ^ 1'b0 ;
  assign n9292 = n9291 ^ n8470 ^ n3258 ;
  assign n9293 = n4566 ^ n2540 ^ 1'b0 ;
  assign n9294 = ( n622 & n2108 ) | ( n622 & ~n9293 ) | ( n2108 & ~n9293 ) ;
  assign n9295 = ~n8459 & n9294 ;
  assign n9296 = n506 & n9295 ;
  assign n9297 = n392 | n1832 ;
  assign n9298 = n392 & ~n9297 ;
  assign n9299 = n223 & ~n9298 ;
  assign n9300 = ~n223 & n9299 ;
  assign n9301 = n339 & n9300 ;
  assign n9302 = ~n578 & n9301 ;
  assign n9303 = n9296 & n9302 ;
  assign n9304 = n3044 & n4979 ;
  assign n9305 = n9304 ^ n6063 ^ 1'b0 ;
  assign n9306 = ~n9303 & n9305 ;
  assign n9307 = ~n7810 & n9306 ;
  assign n9308 = n749 | n7604 ;
  assign n9309 = n9308 ^ n2829 ^ 1'b0 ;
  assign n9310 = n73 & ~n1387 ;
  assign n9311 = n9310 ^ n2816 ^ 1'b0 ;
  assign n9312 = n9311 ^ n4179 ^ 1'b0 ;
  assign n9313 = n9312 ^ n5367 ^ 1'b0 ;
  assign n9314 = n9309 & ~n9313 ;
  assign n9315 = n1839 ^ n318 ^ 1'b0 ;
  assign n9316 = n4674 & n9315 ;
  assign n9317 = n2879 & ~n5810 ;
  assign n9322 = n2867 ^ n1092 ^ 1'b0 ;
  assign n9318 = n4433 & n5128 ;
  assign n9319 = n9318 ^ n7677 ^ 1'b0 ;
  assign n9320 = n3797 ^ n3619 ^ 1'b0 ;
  assign n9321 = n9319 | n9320 ;
  assign n9323 = n9322 ^ n9321 ^ 1'b0 ;
  assign n9324 = n506 ^ n105 ^ 1'b0 ;
  assign n9325 = ~n2932 & n9324 ;
  assign n9326 = n3255 ^ n3071 ^ 1'b0 ;
  assign n9327 = n5061 ^ n3820 ^ 1'b0 ;
  assign n9328 = n259 | n9327 ;
  assign n9329 = n5484 & ~n9328 ;
  assign n9330 = n881 & n9329 ;
  assign n9331 = n1571 & n5001 ;
  assign n9332 = n9331 ^ x5 ^ 1'b0 ;
  assign n9333 = n8510 & ~n9332 ;
  assign n9334 = n9333 ^ n3347 ^ 1'b0 ;
  assign n9335 = ( n5051 & n6551 ) | ( n5051 & n7321 ) | ( n6551 & n7321 ) ;
  assign n9336 = n267 & n6527 ;
  assign n9337 = n3361 & n4382 ;
  assign n9338 = ~n1956 & n3449 ;
  assign n9339 = n221 & n7945 ;
  assign n9340 = ~n7332 & n8943 ;
  assign n9341 = n9340 ^ n1449 ^ 1'b0 ;
  assign n9342 = n2806 | n3446 ;
  assign n9343 = n9342 ^ n668 ^ 1'b0 ;
  assign n9344 = n9343 ^ n7829 ^ n1764 ;
  assign n9345 = n5499 ^ n5057 ^ 1'b0 ;
  assign n9346 = n320 & n1136 ;
  assign n9347 = n2872 ^ n574 ^ 1'b0 ;
  assign n9348 = n1118 & n9347 ;
  assign n9349 = n9348 ^ n2282 ^ 1'b0 ;
  assign n9350 = n9346 & n9349 ;
  assign n9351 = n9350 ^ n870 ^ 1'b0 ;
  assign n9352 = n9345 | n9351 ;
  assign n9353 = n8054 | n9352 ;
  assign n9354 = n3432 ^ n948 ^ 1'b0 ;
  assign n9355 = n2401 | n9100 ;
  assign n9356 = n9354 & ~n9355 ;
  assign n9357 = n3111 & ~n3928 ;
  assign n9358 = ~n3145 & n9357 ;
  assign n9359 = n6699 ^ n1566 ^ 1'b0 ;
  assign n9360 = n9358 | n9359 ;
  assign n9361 = ~n49 & n2288 ;
  assign n9362 = n9360 | n9361 ;
  assign n9363 = n1728 & ~n9362 ;
  assign n9364 = n2403 & ~n8441 ;
  assign n9365 = n2655 & n3167 ;
  assign n9366 = n3135 | n9365 ;
  assign n9367 = n58 & ~n2048 ;
  assign n9368 = n9367 ^ n368 ^ 1'b0 ;
  assign n9369 = ( n5049 & ~n6423 ) | ( n5049 & n6674 ) | ( ~n6423 & n6674 ) ;
  assign n9372 = n1258 ^ n366 ^ 1'b0 ;
  assign n9373 = n9372 ^ n3827 ^ 1'b0 ;
  assign n9370 = n5262 ^ n2409 ^ 1'b0 ;
  assign n9371 = ~n1973 & n9370 ;
  assign n9374 = n9373 ^ n9371 ^ 1'b0 ;
  assign n9375 = ~n305 & n9374 ;
  assign n9376 = ( n2438 & ~n2799 ) | ( n2438 & n9375 ) | ( ~n2799 & n9375 ) ;
  assign n9377 = ~n2684 & n7989 ;
  assign n9378 = n2042 | n9377 ;
  assign n9379 = n3106 ^ n2821 ^ 1'b0 ;
  assign n9380 = n142 | n9379 ;
  assign n9381 = n8908 ^ n6809 ^ 1'b0 ;
  assign n9382 = n2292 ^ n2034 ^ 1'b0 ;
  assign n9383 = n2134 | n9382 ;
  assign n9384 = n4311 & n9383 ;
  assign n9385 = n8279 ^ n1109 ^ 1'b0 ;
  assign n9386 = n9384 & n9385 ;
  assign n9388 = ~n916 & n4745 ;
  assign n9387 = n311 & n8745 ;
  assign n9389 = n9388 ^ n9387 ^ 1'b0 ;
  assign n9390 = n854 | n9389 ;
  assign n9391 = n5217 & ~n5365 ;
  assign n9392 = n706 & ~n3236 ;
  assign n9393 = n9391 & n9392 ;
  assign n9394 = n2805 ^ n17 ^ 1'b0 ;
  assign n9395 = ~n5516 & n9394 ;
  assign n9396 = n9395 ^ n241 ^ 1'b0 ;
  assign n9397 = ~n878 & n9396 ;
  assign n9398 = n6200 & n9397 ;
  assign n9399 = ~n9022 & n9398 ;
  assign n9400 = n4242 & ~n5295 ;
  assign n9401 = n9400 ^ n3721 ^ 1'b0 ;
  assign n9402 = n4670 & n9401 ;
  assign n9403 = n9402 ^ n3579 ^ 1'b0 ;
  assign n9404 = ~n4919 & n9403 ;
  assign n9405 = n2438 ^ n692 ^ 1'b0 ;
  assign n9406 = n154 & n1853 ;
  assign n9407 = n9405 & n9406 ;
  assign n9408 = ~n688 & n9407 ;
  assign n9409 = n4484 | n9408 ;
  assign n9410 = n9409 ^ n8576 ^ 1'b0 ;
  assign n9411 = n9410 ^ n107 ^ 1'b0 ;
  assign n9412 = n2635 ^ n492 ^ 1'b0 ;
  assign n9413 = n6325 | n9412 ;
  assign n9414 = n9413 ^ n1789 ^ 1'b0 ;
  assign n9415 = n6392 ^ n2045 ^ 1'b0 ;
  assign n9416 = n5689 & n9415 ;
  assign n9417 = n9416 ^ n3818 ^ 1'b0 ;
  assign n9418 = n343 & ~n2240 ;
  assign n9419 = n9418 ^ n3415 ^ 1'b0 ;
  assign n9420 = n2833 ^ n2822 ^ 1'b0 ;
  assign n9421 = n978 & n9420 ;
  assign n9422 = n6688 ^ n3011 ^ 1'b0 ;
  assign n9423 = n8560 & ~n9422 ;
  assign n9424 = n846 | n3465 ;
  assign n9425 = ~n1337 & n9424 ;
  assign n9426 = ~n9423 & n9425 ;
  assign n9427 = n4596 | n4666 ;
  assign n9428 = ( n2897 & ~n7282 ) | ( n2897 & n8450 ) | ( ~n7282 & n8450 ) ;
  assign n9429 = n924 & n5606 ;
  assign n9430 = ~n493 & n9429 ;
  assign n9431 = n5638 ^ n5450 ^ 1'b0 ;
  assign n9432 = n2711 & n9431 ;
  assign n9433 = ~n269 & n9432 ;
  assign n9434 = n9433 ^ n2177 ^ 1'b0 ;
  assign n9435 = ~n2252 & n2338 ;
  assign n9436 = ~n6183 & n9435 ;
  assign n9437 = n9436 ^ n7241 ^ 1'b0 ;
  assign n9438 = n7904 & n8449 ;
  assign n9439 = n9438 ^ n2929 ^ 1'b0 ;
  assign n9440 = n2726 | n4158 ;
  assign n9441 = n1430 & ~n6396 ;
  assign n9442 = n2384 & ~n8974 ;
  assign n9443 = n2136 ^ n150 ^ 1'b0 ;
  assign n9444 = n135 | n9443 ;
  assign n9445 = n3370 & ~n9444 ;
  assign n9462 = ~n1884 & n6092 ;
  assign n9463 = ~n2207 & n9462 ;
  assign n9455 = n2097 & n2526 ;
  assign n9456 = n886 & ~n944 ;
  assign n9457 = ~n6568 & n9456 ;
  assign n9458 = n9457 ^ n3891 ^ 1'b0 ;
  assign n9459 = n265 | n9458 ;
  assign n9460 = n4379 & ~n9459 ;
  assign n9461 = n9455 & ~n9460 ;
  assign n9464 = n9463 ^ n9461 ^ n3363 ;
  assign n9446 = n43 & n4626 ;
  assign n9447 = n2408 & n9446 ;
  assign n9448 = n5022 ^ n1690 ^ 1'b0 ;
  assign n9449 = ~n4359 & n9448 ;
  assign n9450 = n9449 ^ n3958 ^ 1'b0 ;
  assign n9451 = ~n9447 & n9450 ;
  assign n9452 = ~n2491 & n5733 ;
  assign n9453 = ~n1905 & n9452 ;
  assign n9454 = n9451 & ~n9453 ;
  assign n9465 = n9464 ^ n9454 ^ 1'b0 ;
  assign n9466 = n2097 | n2818 ;
  assign n9467 = n9466 ^ n4436 ^ 1'b0 ;
  assign n9468 = ~n320 & n3950 ;
  assign n9469 = n434 & n3628 ;
  assign n9470 = n1455 & n9469 ;
  assign n9471 = n5992 | n9470 ;
  assign n9472 = n5541 & n9471 ;
  assign n9473 = n9472 ^ n8831 ^ 1'b0 ;
  assign n9474 = n4571 ^ n1107 ^ 1'b0 ;
  assign n9475 = ~n1066 & n9474 ;
  assign n9476 = n7967 & n9475 ;
  assign n9477 = n6210 ^ n2070 ^ 1'b0 ;
  assign n9478 = n8951 & n9477 ;
  assign n9479 = n2614 & n4174 ;
  assign n9480 = n9136 & n9479 ;
  assign n9481 = n9480 ^ n6940 ^ 1'b0 ;
  assign n9482 = n6910 ^ n4538 ^ 1'b0 ;
  assign n9483 = n5836 | n9482 ;
  assign n9484 = n4056 | n4087 ;
  assign n9485 = n5116 | n7010 ;
  assign n9486 = n8779 ^ n7125 ^ 1'b0 ;
  assign n9488 = n2292 & n3122 ;
  assign n9487 = n3720 | n6340 ;
  assign n9489 = n9488 ^ n9487 ^ 1'b0 ;
  assign n9490 = ~n793 & n1313 ;
  assign n9491 = n9490 ^ n2693 ^ 1'b0 ;
  assign n9492 = ~n1521 & n2555 ;
  assign n9493 = n9491 | n9492 ;
  assign n9494 = n2854 ^ n287 ^ 1'b0 ;
  assign n9495 = n2772 | n9494 ;
  assign n9498 = n987 | n5690 ;
  assign n9499 = n9498 ^ n5853 ^ 1'b0 ;
  assign n9496 = n4914 & n6127 ;
  assign n9497 = n9496 ^ n7841 ^ 1'b0 ;
  assign n9500 = n9499 ^ n9497 ^ n7626 ;
  assign n9501 = n4133 | n6040 ;
  assign n9502 = n9501 ^ n1726 ^ 1'b0 ;
  assign n9503 = n8428 ^ n8235 ^ n4540 ;
  assign n9504 = ~n3700 & n8831 ;
  assign n9505 = n9504 ^ n764 ^ 1'b0 ;
  assign n9506 = n8531 ^ n7390 ^ 1'b0 ;
  assign n9507 = n9505 | n9506 ;
  assign n9508 = n2664 ^ n1521 ^ 1'b0 ;
  assign n9509 = n1920 ^ n1312 ^ 1'b0 ;
  assign n9510 = ~n9508 & n9509 ;
  assign n9511 = n9510 ^ n3605 ^ 1'b0 ;
  assign n9512 = n1085 | n9511 ;
  assign n9513 = n9512 ^ n1944 ^ 1'b0 ;
  assign n9514 = n8273 | n9481 ;
  assign n9515 = n6241 & ~n9514 ;
  assign n9516 = n3881 ^ n3820 ^ 1'b0 ;
  assign n9517 = n2512 & ~n9516 ;
  assign n9518 = n1716 | n9517 ;
  assign n9519 = n4084 & n4260 ;
  assign n9520 = ~n1172 & n9519 ;
  assign n9521 = ~n9518 & n9520 ;
  assign n9522 = ( n397 & ~n441 ) | ( n397 & n5726 ) | ( ~n441 & n5726 ) ;
  assign n9523 = n9522 ^ n692 ^ 1'b0 ;
  assign n9528 = n4113 | n6651 ;
  assign n9524 = n2765 & n7322 ;
  assign n9525 = ~n406 & n9524 ;
  assign n9526 = n3874 ^ n1962 ^ 1'b0 ;
  assign n9527 = n9525 | n9526 ;
  assign n9529 = n9528 ^ n9527 ^ 1'b0 ;
  assign n9530 = ( ~n2310 & n4735 ) | ( ~n2310 & n9529 ) | ( n4735 & n9529 ) ;
  assign n9531 = n7056 ^ n528 ^ 1'b0 ;
  assign n9532 = ~n4363 & n9531 ;
  assign n9533 = ~n7955 & n9532 ;
  assign n9534 = n7825 & n9533 ;
  assign n9535 = n3125 ^ n356 ^ 1'b0 ;
  assign n9536 = n3303 ^ n2648 ^ 1'b0 ;
  assign n9537 = ~n7512 & n9536 ;
  assign n9538 = ~n9535 & n9537 ;
  assign n9539 = n3210 & n8703 ;
  assign n9540 = ~n27 & n2231 ;
  assign n9541 = ~n1349 & n9540 ;
  assign n9542 = ~n1770 & n9541 ;
  assign n9543 = n669 | n9542 ;
  assign n9544 = n7500 ^ n4489 ^ 1'b0 ;
  assign n9545 = n3537 | n5008 ;
  assign n9546 = n478 & ~n1455 ;
  assign n9547 = n9546 ^ n3489 ^ 1'b0 ;
  assign n9548 = n9383 | n9547 ;
  assign n9549 = n9545 | n9548 ;
  assign n9550 = n2902 | n9549 ;
  assign n9551 = ~n1677 & n8040 ;
  assign n9552 = ~n535 & n9551 ;
  assign n9553 = n1245 & n2266 ;
  assign n9554 = n2007 & n2405 ;
  assign n9555 = n5049 & n9554 ;
  assign n9556 = n2243 & ~n9555 ;
  assign n9557 = n4484 & n9556 ;
  assign n9558 = n1623 | n9557 ;
  assign n9559 = n4521 | n9558 ;
  assign n9560 = n896 & n3822 ;
  assign n9561 = n150 & n703 ;
  assign n9562 = n9561 ^ n1477 ^ 1'b0 ;
  assign n9564 = n620 & ~n1155 ;
  assign n9563 = n7337 ^ n144 ^ n115 ;
  assign n9565 = n9564 ^ n9563 ^ 1'b0 ;
  assign n9566 = n9562 | n9565 ;
  assign n9567 = n9566 ^ n1721 ^ n1705 ;
  assign n9568 = n1298 & n9567 ;
  assign n9569 = ~n1365 & n9568 ;
  assign n9570 = n7882 & ~n9569 ;
  assign n9571 = n1083 | n5497 ;
  assign n9572 = n9571 ^ n1456 ^ 1'b0 ;
  assign n9573 = n437 & ~n8169 ;
  assign n9574 = n2267 & n9573 ;
  assign n9582 = n4214 ^ n1434 ^ 1'b0 ;
  assign n9583 = n7694 & ~n9582 ;
  assign n9575 = n4229 | n4894 ;
  assign n9576 = n9575 ^ n5888 ^ 1'b0 ;
  assign n9577 = n1077 ^ n873 ^ 1'b0 ;
  assign n9578 = n9577 ^ n3078 ^ 1'b0 ;
  assign n9579 = n9578 ^ n617 ^ 1'b0 ;
  assign n9580 = ~n4364 & n9579 ;
  assign n9581 = n9576 & n9580 ;
  assign n9584 = n9583 ^ n9581 ^ 1'b0 ;
  assign n9585 = n2918 & n2996 ;
  assign n9586 = n3295 | n5518 ;
  assign n9587 = n3531 & n9586 ;
  assign n9588 = n9587 ^ n5841 ^ 1'b0 ;
  assign n9589 = n2440 & ~n9588 ;
  assign n9590 = n4677 & n5874 ;
  assign n9592 = n4390 | n6297 ;
  assign n9591 = n2576 & ~n9562 ;
  assign n9593 = n9592 ^ n9591 ^ n2384 ;
  assign n9594 = n3078 ^ n561 ^ 1'b0 ;
  assign n9595 = ~n4607 & n9594 ;
  assign n9596 = ~n940 & n9595 ;
  assign n9597 = ~n581 & n9596 ;
  assign n9598 = n318 & ~n6338 ;
  assign n9599 = n3080 & n6811 ;
  assign n9600 = n1937 & ~n5607 ;
  assign n9601 = ( n1669 & n4111 ) | ( n1669 & n9600 ) | ( n4111 & n9600 ) ;
  assign n9602 = n9121 ^ n6681 ^ 1'b0 ;
  assign n9603 = n2968 & ~n5247 ;
  assign n9604 = n9603 ^ n213 ^ 1'b0 ;
  assign n9605 = n57 & ~n2366 ;
  assign n9606 = n1673 & ~n9605 ;
  assign n9607 = n9606 ^ n6892 ^ 1'b0 ;
  assign n9608 = n5431 & n9607 ;
  assign n9609 = n1933 | n4235 ;
  assign n9610 = n6527 ^ n1121 ^ 1'b0 ;
  assign n9611 = n7256 & n9610 ;
  assign n9612 = ( ~n362 & n4439 ) | ( ~n362 & n9463 ) | ( n4439 & n9463 ) ;
  assign n9613 = n9612 ^ n9601 ^ 1'b0 ;
  assign n9614 = n4802 | n5137 ;
  assign n9615 = n9613 & ~n9614 ;
  assign n9616 = n4276 ^ n3943 ^ 1'b0 ;
  assign n9617 = n322 & ~n1961 ;
  assign n9619 = ~n1868 & n6709 ;
  assign n9620 = n9619 ^ n3242 ^ 1'b0 ;
  assign n9618 = n425 & n4602 ;
  assign n9621 = n9620 ^ n9618 ^ 1'b0 ;
  assign n9623 = n4061 ^ n1946 ^ 1'b0 ;
  assign n9622 = n890 & ~n2981 ;
  assign n9624 = n9623 ^ n9622 ^ 1'b0 ;
  assign n9625 = ( n9617 & n9621 ) | ( n9617 & n9624 ) | ( n9621 & n9624 ) ;
  assign n9626 = n5121 & n5168 ;
  assign n9627 = ~n1590 & n9626 ;
  assign n9628 = n7374 | n9627 ;
  assign n9629 = n9153 & ~n9628 ;
  assign n9630 = n3031 ^ n2926 ^ 1'b0 ;
  assign n9631 = n1627 & n9630 ;
  assign n9632 = n9543 & n9631 ;
  assign n9633 = n6198 & ~n8852 ;
  assign n9634 = n9633 ^ n3001 ^ 1'b0 ;
  assign n9635 = n1038 & ~n4086 ;
  assign n9636 = n9634 & n9635 ;
  assign n9637 = ~n1738 & n2206 ;
  assign n9638 = ~n1701 & n9637 ;
  assign n9639 = n5177 | n9638 ;
  assign n9640 = n2020 | n9414 ;
  assign n9641 = n8396 | n9640 ;
  assign n9642 = n354 & ~n3628 ;
  assign n9643 = ( ~n1181 & n4054 ) | ( ~n1181 & n9642 ) | ( n4054 & n9642 ) ;
  assign n9644 = n9643 ^ n6025 ^ 1'b0 ;
  assign n9645 = n749 & n9644 ;
  assign n9646 = n4709 | n7344 ;
  assign n9647 = n1553 | n9646 ;
  assign n9648 = n214 | n9647 ;
  assign n9649 = n2807 ^ n1045 ^ 1'b0 ;
  assign n9650 = n746 & n9649 ;
  assign n9651 = n225 | n9650 ;
  assign n9652 = ~n202 & n5360 ;
  assign n9653 = ( ~n465 & n3026 ) | ( ~n465 & n9652 ) | ( n3026 & n9652 ) ;
  assign n9654 = n9651 & n9653 ;
  assign n9655 = n9654 ^ n9293 ^ 1'b0 ;
  assign n9659 = n1213 & n1845 ;
  assign n9656 = n2288 | n6401 ;
  assign n9657 = n6225 & ~n9656 ;
  assign n9658 = n7607 | n9657 ;
  assign n9660 = n9659 ^ n9658 ^ 1'b0 ;
  assign n9661 = n4229 ^ n3414 ^ 1'b0 ;
  assign n9662 = ( n3974 & ~n9317 ) | ( n3974 & n9661 ) | ( ~n9317 & n9661 ) ;
  assign n9663 = ~n401 & n4546 ;
  assign n9664 = n326 & ~n2140 ;
  assign n9665 = ( n505 & ~n6356 ) | ( n505 & n6931 ) | ( ~n6356 & n6931 ) ;
  assign n9666 = n5662 & ~n7369 ;
  assign n9667 = ~n6711 & n9666 ;
  assign n9668 = ~n3437 & n6232 ;
  assign n9669 = n3199 & ~n5183 ;
  assign n9670 = n1337 & n9669 ;
  assign n9671 = n9670 ^ n1623 ^ 1'b0 ;
  assign n9672 = n4599 & n9671 ;
  assign n9673 = n3359 | n3578 ;
  assign n9674 = n249 & n9673 ;
  assign n9675 = n5346 ^ n2914 ^ 1'b0 ;
  assign n9676 = n5689 & n9675 ;
  assign n9677 = n270 & n6589 ;
  assign n9678 = n2023 | n9677 ;
  assign n9679 = n6419 ^ n5223 ^ 1'b0 ;
  assign n9680 = n9679 ^ n697 ^ 1'b0 ;
  assign n9681 = n1668 & ~n5048 ;
  assign n9682 = n9681 ^ n2815 ^ 1'b0 ;
  assign n9683 = ~n4122 & n9682 ;
  assign n9684 = n9680 & n9683 ;
  assign n9686 = ~n3877 & n5082 ;
  assign n9685 = n966 & ~n2227 ;
  assign n9687 = n9686 ^ n9685 ^ 1'b0 ;
  assign n9688 = n1264 & ~n1769 ;
  assign n9689 = n9688 ^ n5766 ^ n495 ;
  assign n9690 = n3238 | n7771 ;
  assign n9691 = n9689 | n9690 ;
  assign n9692 = n40 & ~n9691 ;
  assign n9693 = n9692 ^ n2219 ^ 1'b0 ;
  assign n9694 = n723 ^ n411 ^ 1'b0 ;
  assign n9695 = ~n6093 & n9694 ;
  assign n9696 = n9695 ^ n7601 ^ 1'b0 ;
  assign n9697 = n8187 ^ n6560 ^ 1'b0 ;
  assign n9698 = ( n1293 & ~n2930 ) | ( n1293 & n3082 ) | ( ~n2930 & n3082 ) ;
  assign n9699 = n372 | n3657 ;
  assign n9703 = n4837 ^ n2588 ^ 1'b0 ;
  assign n9700 = ( n1068 & n1723 ) | ( n1068 & n2399 ) | ( n1723 & n2399 ) ;
  assign n9701 = n5589 ^ n4561 ^ 1'b0 ;
  assign n9702 = n9700 & n9701 ;
  assign n9704 = n9703 ^ n9702 ^ 1'b0 ;
  assign n9705 = n5397 ^ n3438 ^ 1'b0 ;
  assign n9706 = n557 & ~n9705 ;
  assign n9707 = n4020 ^ n1453 ^ 1'b0 ;
  assign n9708 = ~n373 & n3680 ;
  assign n9709 = ~n9707 & n9708 ;
  assign n9710 = n7170 ^ n5639 ^ 1'b0 ;
  assign n9711 = n6556 ^ n577 ^ 1'b0 ;
  assign n9712 = ~n3315 & n9711 ;
  assign n9713 = n9712 ^ n1057 ^ 1'b0 ;
  assign n9714 = n164 | n9713 ;
  assign n9715 = n1582 | n2952 ;
  assign n9716 = ~n3301 & n9715 ;
  assign n9717 = n302 & n4707 ;
  assign n9718 = n1189 & n9717 ;
  assign n9719 = ~n9716 & n9718 ;
  assign n9720 = n121 & ~n4615 ;
  assign n9723 = n1182 | n1779 ;
  assign n9724 = n5805 & ~n9723 ;
  assign n9721 = ~n280 & n4528 ;
  assign n9722 = ~n1709 & n9721 ;
  assign n9725 = n9724 ^ n9722 ^ 1'b0 ;
  assign n9726 = ( n1600 & ~n9720 ) | ( n1600 & n9725 ) | ( ~n9720 & n9725 ) ;
  assign n9728 = n2367 & n4189 ;
  assign n9727 = n3756 & ~n7660 ;
  assign n9729 = n9728 ^ n9727 ^ 1'b0 ;
  assign n9730 = n4572 ^ n1742 ^ 1'b0 ;
  assign n9731 = n9730 ^ n562 ^ 1'b0 ;
  assign n9732 = n7475 ^ n3239 ^ 1'b0 ;
  assign n9733 = n3093 ^ n2347 ^ 1'b0 ;
  assign n9734 = n2104 & n2662 ;
  assign n9735 = n9734 ^ n1198 ^ 1'b0 ;
  assign n9736 = ~n360 & n2991 ;
  assign n9737 = n2861 & n9736 ;
  assign n9738 = n9737 ^ n1736 ^ 1'b0 ;
  assign n9739 = ~n6485 & n9738 ;
  assign n9740 = n1411 & n9739 ;
  assign n9741 = n9740 ^ n3526 ^ n2101 ;
  assign n9742 = n9735 & n9741 ;
  assign n9743 = n1361 & n9742 ;
  assign n9744 = n1523 ^ n1042 ^ n997 ;
  assign n9745 = n9744 ^ n3998 ^ 1'b0 ;
  assign n9746 = n5360 | n9745 ;
  assign n9747 = ~n1889 & n4256 ;
  assign n9748 = n9746 & n9747 ;
  assign n9749 = n9748 ^ n1618 ^ 1'b0 ;
  assign n9753 = n2771 ^ n35 ^ 1'b0 ;
  assign n9754 = n9753 ^ n2754 ^ 1'b0 ;
  assign n9750 = n5007 ^ n668 ^ 1'b0 ;
  assign n9751 = ~n997 & n9750 ;
  assign n9752 = n9751 ^ n880 ^ 1'b0 ;
  assign n9755 = n9754 ^ n9752 ^ 1'b0 ;
  assign n9756 = n1069 & ~n1219 ;
  assign n9757 = n9756 ^ n5080 ^ 1'b0 ;
  assign n9758 = n9755 | n9757 ;
  assign n9759 = n3639 ^ n2569 ^ 1'b0 ;
  assign n9760 = ~n225 & n9759 ;
  assign n9761 = n9760 ^ n4317 ^ 1'b0 ;
  assign n9762 = n4733 ^ n71 ^ 1'b0 ;
  assign n9763 = n9762 ^ n4335 ^ 1'b0 ;
  assign n9764 = n2900 & ~n3252 ;
  assign n9765 = n9763 & n9764 ;
  assign n9766 = ~n5382 & n5551 ;
  assign n9767 = n978 | n9766 ;
  assign n9768 = n5031 | n9767 ;
  assign n9769 = n9768 ^ n4256 ^ n669 ;
  assign n9774 = n2626 & ~n7486 ;
  assign n9775 = n2588 & n9774 ;
  assign n9770 = n622 & n3227 ;
  assign n9771 = n9770 ^ n4083 ^ 1'b0 ;
  assign n9772 = n2879 | n9771 ;
  assign n9773 = n9772 ^ n1109 ^ 1'b0 ;
  assign n9776 = n9775 ^ n9773 ^ 1'b0 ;
  assign n9777 = n233 & ~n3797 ;
  assign n9778 = n1479 & n4428 ;
  assign n9779 = ~n9770 & n9778 ;
  assign n9780 = n559 & n6094 ;
  assign n9781 = ( ~n3555 & n4484 ) | ( ~n3555 & n9780 ) | ( n4484 & n9780 ) ;
  assign n9782 = n9781 ^ n7922 ^ 1'b0 ;
  assign n9783 = n9779 | n9782 ;
  assign n9784 = ( n3027 & ~n3225 ) | ( n3027 & n9210 ) | ( ~n3225 & n9210 ) ;
  assign n9785 = n2438 | n7657 ;
  assign n9786 = n1301 & ~n9785 ;
  assign n9787 = n9786 ^ n6180 ^ 1'b0 ;
  assign n9788 = n3635 | n3820 ;
  assign n9789 = n2311 | n8974 ;
  assign n9790 = n3088 ^ n3031 ^ 1'b0 ;
  assign n9791 = ~n1971 & n7407 ;
  assign n9792 = n1889 & n9791 ;
  assign n9793 = n5227 & ~n9792 ;
  assign n9794 = n9793 ^ n9288 ^ 1'b0 ;
  assign n9795 = x2 | n880 ;
  assign n9796 = n9795 ^ n4982 ^ n30 ;
  assign n9797 = n9796 ^ n248 ^ 1'b0 ;
  assign n9798 = n9797 ^ n1204 ^ 1'b0 ;
  assign n9799 = n3379 | n9798 ;
  assign n9800 = n162 & ~n1592 ;
  assign n9801 = n365 & ~n9800 ;
  assign n9802 = n4464 & n9801 ;
  assign n9803 = ~n3693 & n9153 ;
  assign n9804 = ( n696 & ~n3191 ) | ( n696 & n9803 ) | ( ~n3191 & n9803 ) ;
  assign n9805 = n2101 & ~n6012 ;
  assign n9806 = ~n2363 & n9805 ;
  assign n9807 = x10 & ~n9806 ;
  assign n9808 = ~n5417 & n9807 ;
  assign n9809 = n2417 & ~n9808 ;
  assign n9810 = n9804 & n9809 ;
  assign n9811 = n2343 & ~n9810 ;
  assign n9812 = n9802 & n9811 ;
  assign n9813 = n2961 | n9361 ;
  assign n9814 = n9361 & ~n9813 ;
  assign n9815 = n9812 | n9814 ;
  assign n9816 = n6957 & ~n9815 ;
  assign n9817 = n957 & ~n6239 ;
  assign n9818 = n9817 ^ n805 ^ 1'b0 ;
  assign n9819 = n4578 | n9818 ;
  assign n9824 = n1668 & n4194 ;
  assign n9825 = n9824 ^ n5236 ^ 1'b0 ;
  assign n9822 = n1552 & ~n3946 ;
  assign n9823 = n6696 & n9822 ;
  assign n9820 = n1042 | n4883 ;
  assign n9821 = n9820 ^ n3258 ^ 1'b0 ;
  assign n9826 = n9825 ^ n9823 ^ n9821 ;
  assign n9827 = n6465 & n9826 ;
  assign n9828 = n5438 ^ n1829 ^ 1'b0 ;
  assign n9829 = n5189 | n9828 ;
  assign n9830 = n8217 | n9829 ;
  assign n9831 = n1639 & ~n9830 ;
  assign n9832 = n3788 & ~n9831 ;
  assign n9833 = ~n3859 & n5950 ;
  assign n9834 = n3631 & n5375 ;
  assign n9835 = n2046 & n9834 ;
  assign n9836 = n9835 ^ n7591 ^ n6907 ;
  assign n9837 = n5080 ^ n4254 ^ 1'b0 ;
  assign n9839 = n4551 ^ n1993 ^ 1'b0 ;
  assign n9838 = n357 | n3622 ;
  assign n9840 = n9839 ^ n9838 ^ 1'b0 ;
  assign n9841 = n6116 ^ n4651 ^ 1'b0 ;
  assign n9842 = n863 & ~n9841 ;
  assign n9843 = n9840 & ~n9842 ;
  assign n9844 = n1366 | n3113 ;
  assign n9845 = n9844 ^ n2549 ^ 1'b0 ;
  assign n9846 = ~n9843 & n9845 ;
  assign n9847 = n4395 ^ n2638 ^ 1'b0 ;
  assign n9848 = ~n4307 & n9847 ;
  assign n9849 = ~n1867 & n9848 ;
  assign n9850 = ~n9846 & n9849 ;
  assign n9851 = ( n511 & n1858 ) | ( n511 & n9080 ) | ( n1858 & n9080 ) ;
  assign n9852 = n374 | n1143 ;
  assign n9853 = n9852 ^ n983 ^ 1'b0 ;
  assign n9854 = n9851 | n9853 ;
  assign n9855 = n9854 ^ n5448 ^ 1'b0 ;
  assign n9862 = ~n3776 & n9577 ;
  assign n9856 = n6564 ^ n2134 ^ 1'b0 ;
  assign n9857 = ~n8099 & n9856 ;
  assign n9858 = n9857 ^ n8105 ^ 1'b0 ;
  assign n9859 = n2721 ^ n1868 ^ 1'b0 ;
  assign n9860 = n4041 & ~n9859 ;
  assign n9861 = n9858 & n9860 ;
  assign n9863 = n9862 ^ n9861 ^ 1'b0 ;
  assign n9864 = ~n822 & n4275 ;
  assign n9865 = n9864 ^ n395 ^ 1'b0 ;
  assign n9866 = n3050 | n9865 ;
  assign n9867 = n8792 & ~n9866 ;
  assign n9868 = n2791 | n3777 ;
  assign n9869 = n3651 | n4523 ;
  assign n9870 = n9869 ^ n3172 ^ 1'b0 ;
  assign n9871 = n9870 ^ n4810 ^ n782 ;
  assign n9872 = n6732 & n9871 ;
  assign n9873 = n9872 ^ n8500 ^ 1'b0 ;
  assign n9874 = ~n9868 & n9873 ;
  assign n9875 = n7099 ^ n4733 ^ n1032 ;
  assign n9876 = n1615 & ~n9875 ;
  assign n9877 = n9876 ^ n8857 ^ 1'b0 ;
  assign n9878 = n2532 | n9877 ;
  assign n9879 = n1486 & ~n3505 ;
  assign n9880 = n9879 ^ n1488 ^ 1'b0 ;
  assign n9882 = n4054 ^ n3290 ^ 1'b0 ;
  assign n9881 = n886 & ~n5607 ;
  assign n9883 = n9882 ^ n9881 ^ 1'b0 ;
  assign n9884 = n7778 ^ n6285 ^ n3229 ;
  assign n9885 = n5463 & ~n6586 ;
  assign n9886 = n917 & n9885 ;
  assign n9887 = n1705 ^ n1307 ^ 1'b0 ;
  assign n9888 = n5314 ^ n4474 ^ 1'b0 ;
  assign n9889 = n6972 & n9888 ;
  assign n9890 = n9889 ^ n829 ^ 1'b0 ;
  assign n9891 = n9887 | n9890 ;
  assign n9892 = n6971 ^ n2955 ^ n325 ;
  assign n9893 = ~n3617 & n9892 ;
  assign n9894 = n8926 ^ n6817 ^ 1'b0 ;
  assign n9895 = n1167 & n9894 ;
  assign n9896 = n5256 & n9895 ;
  assign n9897 = n9896 ^ n6925 ^ 1'b0 ;
  assign n9898 = n9624 & ~n9897 ;
  assign n9899 = n1742 & ~n3683 ;
  assign n9900 = n7333 ^ n2439 ^ 1'b0 ;
  assign n9901 = ~n9899 & n9900 ;
  assign n9903 = n1161 & n3473 ;
  assign n9904 = ~n162 & n9903 ;
  assign n9905 = n2894 & ~n9904 ;
  assign n9902 = n260 & n6238 ;
  assign n9906 = n9905 ^ n9902 ^ 1'b0 ;
  assign n9907 = n9906 ^ n5544 ^ 1'b0 ;
  assign n9908 = n120 & n3240 ;
  assign n9909 = n4053 ^ n2515 ^ 1'b0 ;
  assign n9910 = n1945 | n9909 ;
  assign n9921 = n7398 ^ n2086 ^ n497 ;
  assign n9911 = n4241 ^ n2956 ^ 1'b0 ;
  assign n9912 = n291 | n9911 ;
  assign n9913 = n9912 ^ n927 ^ 1'b0 ;
  assign n9914 = n9721 & n9913 ;
  assign n9915 = ~n4546 & n9914 ;
  assign n9916 = n9915 ^ n3687 ^ n2621 ;
  assign n9917 = n9916 ^ n40 ^ 1'b0 ;
  assign n9918 = ~n5124 & n9917 ;
  assign n9919 = ~n839 & n9918 ;
  assign n9920 = n8265 & ~n9919 ;
  assign n9922 = n9921 ^ n9920 ^ 1'b0 ;
  assign n9923 = ( n2408 & n4997 ) | ( n2408 & ~n6817 ) | ( n4997 & ~n6817 ) ;
  assign n9924 = n6729 & ~n7475 ;
  assign n9925 = ~n8915 & n9924 ;
  assign n9926 = ~n1976 & n2501 ;
  assign n9927 = n6033 & n9926 ;
  assign n9928 = n6671 ^ n3041 ^ 1'b0 ;
  assign n9929 = n931 | n9928 ;
  assign n9930 = n458 | n5403 ;
  assign n9931 = n3890 & ~n9930 ;
  assign n9932 = n9931 ^ n2894 ^ 1'b0 ;
  assign n9933 = n9336 & n9932 ;
  assign n9934 = n466 | n4546 ;
  assign n9935 = n1726 | n6464 ;
  assign n9936 = ( n3469 & ~n3903 ) | ( n3469 & n9935 ) | ( ~n3903 & n9935 ) ;
  assign n9937 = n4575 & ~n9936 ;
  assign n9938 = ~n5268 & n9937 ;
  assign n9939 = n3987 & ~n9938 ;
  assign n9940 = n3474 & n9939 ;
  assign n9941 = n4468 | n9189 ;
  assign n9942 = n7066 | n9941 ;
  assign n9943 = n9942 ^ n3115 ^ 1'b0 ;
  assign n9944 = ~n6065 & n8462 ;
  assign n9945 = ~n3186 & n9944 ;
  assign n9946 = ~n617 & n1323 ;
  assign n9947 = n3574 | n9946 ;
  assign n9948 = n9947 ^ n1932 ^ 1'b0 ;
  assign n9949 = n6106 ^ n304 ^ 1'b0 ;
  assign n9950 = n384 | n860 ;
  assign n9951 = n8093 ^ n7389 ^ 1'b0 ;
  assign n9952 = ~n9950 & n9951 ;
  assign n9953 = ( n56 & n9949 ) | ( n56 & n9952 ) | ( n9949 & n9952 ) ;
  assign n9954 = n1154 ^ n931 ^ 1'b0 ;
  assign n9955 = n3897 & n9954 ;
  assign n9958 = n2902 ^ n896 ^ 1'b0 ;
  assign n9959 = n6927 | n9958 ;
  assign n9956 = n3774 & ~n4013 ;
  assign n9957 = ~n975 & n9956 ;
  assign n9960 = n9959 ^ n9957 ^ 1'b0 ;
  assign n9961 = ~n5663 & n9960 ;
  assign n9962 = ( n2541 & n9955 ) | ( n2541 & ~n9961 ) | ( n9955 & ~n9961 ) ;
  assign n9963 = n7759 ^ n7651 ^ n3775 ;
  assign n9964 = n9963 ^ n2580 ^ 1'b0 ;
  assign n9965 = n697 & n9964 ;
  assign n9966 = n967 | n6160 ;
  assign n9967 = ( ~n31 & n6377 ) | ( ~n31 & n9966 ) | ( n6377 & n9966 ) ;
  assign n9968 = ( n1174 & n5473 ) | ( n1174 & ~n7589 ) | ( n5473 & ~n7589 ) ;
  assign n9969 = n9968 ^ n5077 ^ 1'b0 ;
  assign n9972 = ~n8180 & n8537 ;
  assign n9970 = n5546 ^ n49 ^ 1'b0 ;
  assign n9971 = n124 | n9970 ;
  assign n9973 = n9972 ^ n9971 ^ 1'b0 ;
  assign n9974 = ~n2330 & n8083 ;
  assign n9975 = n7280 ^ n4671 ^ 1'b0 ;
  assign n9976 = n5628 ^ n4873 ^ 1'b0 ;
  assign n9977 = ~n2008 & n9976 ;
  assign n9978 = n4905 ^ n2371 ^ 1'b0 ;
  assign n9979 = n5485 & ~n9978 ;
  assign n9980 = ~n5320 & n8539 ;
  assign n9981 = n9980 ^ n2986 ^ 1'b0 ;
  assign n9982 = n1471 | n9981 ;
  assign n9983 = n9982 ^ n8510 ^ 1'b0 ;
  assign n9984 = n2151 & ~n5812 ;
  assign n9985 = n7501 & ~n9984 ;
  assign n9986 = ~n6267 & n9985 ;
  assign n9987 = n9986 ^ n1021 ^ 1'b0 ;
  assign n9988 = n5128 ^ n3584 ^ 1'b0 ;
  assign n9989 = ~n9364 & n9988 ;
  assign n9990 = n4218 & n9989 ;
  assign n9991 = n6221 ^ n292 ^ 1'b0 ;
  assign n9992 = n395 & ~n9991 ;
  assign n9993 = n9992 ^ n6674 ^ 1'b0 ;
  assign n9994 = n9196 & ~n9993 ;
  assign n9995 = n1350 ^ n387 ^ 1'b0 ;
  assign n9996 = n6006 & ~n9995 ;
  assign n9997 = n1469 & ~n6766 ;
  assign n9998 = n3746 & n9997 ;
  assign n9999 = n9998 ^ n505 ^ 1'b0 ;
  assign n10000 = n267 & ~n9999 ;
  assign n10001 = n10000 ^ n4650 ^ n858 ;
  assign n10002 = n1347 & n2829 ;
  assign n10003 = n1173 & n1673 ;
  assign n10004 = ~n365 & n10003 ;
  assign n10005 = n2185 & ~n7193 ;
  assign n10006 = n6449 & n6790 ;
  assign n10007 = n10006 ^ n3305 ^ 1'b0 ;
  assign n10012 = n2377 | n3858 ;
  assign n10008 = n5744 ^ n296 ^ 1'b0 ;
  assign n10009 = n2637 & n4213 ;
  assign n10010 = n1138 & n10009 ;
  assign n10011 = n10008 & ~n10010 ;
  assign n10013 = n10012 ^ n10011 ^ 1'b0 ;
  assign n10014 = n3933 & ~n10013 ;
  assign n10015 = n7044 & n10014 ;
  assign n10016 = n5234 ^ n3030 ^ n283 ;
  assign n10017 = n3207 ^ n2787 ^ 1'b0 ;
  assign n10018 = n9266 | n10017 ;
  assign n10019 = ( n1993 & n4044 ) | ( n1993 & n8720 ) | ( n4044 & n8720 ) ;
  assign n10020 = n3576 & n9248 ;
  assign n10021 = ~n5235 & n10020 ;
  assign n10022 = ( ~n4446 & n9335 ) | ( ~n4446 & n10021 ) | ( n9335 & n10021 ) ;
  assign n10023 = n1607 & n2589 ;
  assign n10024 = n10023 ^ n4114 ^ 1'b0 ;
  assign n10025 = n6762 | n10024 ;
  assign n10026 = n8711 ^ n379 ^ 1'b0 ;
  assign n10027 = n7800 & n10026 ;
  assign n10028 = n10027 ^ n2602 ^ 1'b0 ;
  assign n10029 = ~n10025 & n10028 ;
  assign n10030 = n1839 ^ n1117 ^ 1'b0 ;
  assign n10031 = ~n559 & n10030 ;
  assign n10032 = n1699 & ~n7327 ;
  assign n10033 = n10032 ^ n4029 ^ 1'b0 ;
  assign n10034 = n1401 & ~n10033 ;
  assign n10035 = n1306 | n1366 ;
  assign n10036 = n10035 ^ n4666 ^ 1'b0 ;
  assign n10037 = n419 & ~n10036 ;
  assign n10038 = n1307 | n5179 ;
  assign n10039 = ( n6762 & n8874 ) | ( n6762 & n10038 ) | ( n8874 & n10038 ) ;
  assign n10040 = n8177 & n10039 ;
  assign n10041 = n2736 & n8985 ;
  assign n10042 = n2077 ^ n989 ^ 1'b0 ;
  assign n10043 = n5435 & n7878 ;
  assign n10044 = n10043 ^ n1674 ^ 1'b0 ;
  assign n10045 = n749 ^ n132 ^ 1'b0 ;
  assign n10046 = n126 | n714 ;
  assign n10047 = n10046 ^ n861 ^ 1'b0 ;
  assign n10049 = n4716 ^ n1526 ^ 1'b0 ;
  assign n10048 = ~n228 & n2118 ;
  assign n10050 = n10049 ^ n10048 ^ 1'b0 ;
  assign n10051 = n10047 | n10050 ;
  assign n10052 = n8884 ^ n437 ^ 1'b0 ;
  assign n10053 = ~n2041 & n10052 ;
  assign n10054 = n10053 ^ n1961 ^ 1'b0 ;
  assign n10055 = n5896 ^ n150 ^ 1'b0 ;
  assign n10056 = n7018 & n8453 ;
  assign n10057 = n5989 | n9919 ;
  assign n10058 = x6 & n521 ;
  assign n10059 = n10058 ^ n1351 ^ 1'b0 ;
  assign n10060 = n150 & ~n10059 ;
  assign n10061 = ( n1534 & ~n6622 ) | ( n1534 & n10060 ) | ( ~n6622 & n10060 ) ;
  assign n10063 = ( n2504 & n5085 ) | ( n2504 & n8586 ) | ( n5085 & n8586 ) ;
  assign n10064 = n10063 ^ n2336 ^ 1'b0 ;
  assign n10065 = n1535 | n10064 ;
  assign n10062 = ~n4119 & n6616 ;
  assign n10066 = n10065 ^ n10062 ^ 1'b0 ;
  assign n10067 = n2739 ^ n680 ^ x6 ;
  assign n10068 = n997 | n10067 ;
  assign n10069 = n8843 & ~n10068 ;
  assign n10070 = ( n7681 & ~n9361 ) | ( n7681 & n10069 ) | ( ~n9361 & n10069 ) ;
  assign n10071 = n9593 ^ n229 ^ 1'b0 ;
  assign n10072 = ~n451 & n1578 ;
  assign n10073 = n10072 ^ n320 ^ 1'b0 ;
  assign n10074 = n2214 ^ n2080 ^ 1'b0 ;
  assign n10075 = n1627 | n10074 ;
  assign n10076 = n6351 ^ n3968 ^ n3488 ;
  assign n10077 = n7627 ^ n3763 ^ 1'b0 ;
  assign n10078 = n9170 & ~n10077 ;
  assign n10079 = n4702 ^ n1819 ^ 1'b0 ;
  assign n10080 = n10079 ^ n9363 ^ 1'b0 ;
  assign n10081 = n423 & ~n10080 ;
  assign n10082 = n3314 ^ n2816 ^ 1'b0 ;
  assign n10083 = ~n2393 & n10082 ;
  assign n10084 = ( n4685 & n9233 ) | ( n4685 & n10083 ) | ( n9233 & n10083 ) ;
  assign n10085 = n1199 & ~n1465 ;
  assign n10086 = n10085 ^ n4572 ^ 1'b0 ;
  assign n10087 = n2163 ^ n1742 ^ 1'b0 ;
  assign n10088 = ~n1334 & n9611 ;
  assign n10089 = n10088 ^ n2265 ^ 1'b0 ;
  assign n10090 = n3239 ^ n1116 ^ 1'b0 ;
  assign n10091 = n1298 & ~n10090 ;
  assign n10092 = n10091 ^ n4280 ^ 1'b0 ;
  assign n10093 = n3214 | n9014 ;
  assign n10094 = n431 | n3197 ;
  assign n10095 = n10094 ^ n2779 ^ 1'b0 ;
  assign n10096 = n6869 & n10095 ;
  assign n10098 = ( n88 & ~n311 ) | ( n88 & n2427 ) | ( ~n311 & n2427 ) ;
  assign n10097 = ~n970 & n2489 ;
  assign n10099 = n10098 ^ n10097 ^ 1'b0 ;
  assign n10100 = n4275 & n10099 ;
  assign n10101 = ~n982 & n10100 ;
  assign n10102 = ( ~n3496 & n5982 ) | ( ~n3496 & n10101 ) | ( n5982 & n10101 ) ;
  assign n10103 = n10096 & ~n10102 ;
  assign n10104 = ~n4568 & n10103 ;
  assign n10105 = ~n1896 & n10104 ;
  assign n10106 = n5779 ^ n1734 ^ 1'b0 ;
  assign n10107 = n7771 ^ n5107 ^ 1'b0 ;
  assign n10108 = n10107 ^ n6182 ^ 1'b0 ;
  assign n10109 = n115 | n6079 ;
  assign n10110 = n10109 ^ n9204 ^ 1'b0 ;
  assign n10111 = ~n9088 & n10110 ;
  assign n10112 = ~n2628 & n4947 ;
  assign n10113 = n1497 & ~n10112 ;
  assign n10114 = n10113 ^ n7609 ^ 1'b0 ;
  assign n10115 = n3541 & ~n5260 ;
  assign n10116 = ~n4910 & n8781 ;
  assign n10117 = ~n10115 & n10116 ;
  assign n10118 = ( n1511 & n2994 ) | ( n1511 & n10117 ) | ( n2994 & n10117 ) ;
  assign n10119 = ~n127 & n6060 ;
  assign n10120 = n4735 & ~n9080 ;
  assign n10121 = n1111 ^ n1096 ^ 1'b0 ;
  assign n10122 = n4285 | n10121 ;
  assign n10123 = n1767 | n10122 ;
  assign n10124 = n9470 ^ n4104 ^ 1'b0 ;
  assign n10125 = n10124 ^ n4698 ^ 1'b0 ;
  assign n10126 = ~n4478 & n10125 ;
  assign n10127 = n3258 & ~n7380 ;
  assign n10128 = n10127 ^ n6450 ^ 1'b0 ;
  assign n10129 = n10128 ^ n9522 ^ n2277 ;
  assign n10130 = n822 | n1677 ;
  assign n10131 = n2658 | n10130 ;
  assign n10132 = n10131 ^ n5438 ^ 1'b0 ;
  assign n10133 = ~n1573 & n10132 ;
  assign n10134 = n5849 ^ n3647 ^ 1'b0 ;
  assign n10135 = ~n3207 & n4704 ;
  assign n10136 = n3569 | n9532 ;
  assign n10137 = n3268 & ~n3693 ;
  assign n10138 = n1080 & ~n9002 ;
  assign n10139 = n10138 ^ n6534 ^ 1'b0 ;
  assign n10140 = n1521 & n10139 ;
  assign n10141 = ~n3369 & n8120 ;
  assign n10142 = n3044 & ~n10141 ;
  assign n10143 = n9360 & n9698 ;
  assign n10144 = n2985 ^ n1275 ^ 1'b0 ;
  assign n10145 = n9292 & ~n10144 ;
  assign n10146 = n10066 ^ n3423 ^ 1'b0 ;
  assign n10147 = n1329 & ~n3507 ;
  assign n10148 = n535 & n2473 ;
  assign n10149 = n6575 & n10148 ;
  assign n10150 = ( n1505 & n10048 ) | ( n1505 & n10149 ) | ( n10048 & n10149 ) ;
  assign n10151 = n9163 ^ n1023 ^ 1'b0 ;
  assign n10152 = ~n7624 & n10151 ;
  assign n10153 = n2340 | n7977 ;
  assign n10154 = n7270 ^ n5364 ^ 1'b0 ;
  assign n10155 = n4907 ^ n3715 ^ 1'b0 ;
  assign n10156 = n10154 | n10155 ;
  assign n10157 = n1192 | n10156 ;
  assign n10158 = n1908 ^ n1600 ^ 1'b0 ;
  assign n10159 = n10158 ^ n7851 ^ 1'b0 ;
  assign n10160 = n10159 ^ n6408 ^ 1'b0 ;
  assign n10161 = n466 | n7459 ;
  assign n10162 = ~n2337 & n10161 ;
  assign n10163 = n1044 ^ n113 ^ 1'b0 ;
  assign n10164 = n221 & ~n10163 ;
  assign n10165 = n8159 ^ n5940 ^ 1'b0 ;
  assign n10166 = n10164 & ~n10165 ;
  assign n10167 = n204 & ~n4228 ;
  assign n10168 = n105 | n3197 ;
  assign n10169 = n4457 & ~n8708 ;
  assign n10170 = n10168 & n10169 ;
  assign n10171 = ~n1256 & n7567 ;
  assign n10172 = n2619 | n3122 ;
  assign n10173 = n10172 ^ n755 ^ 1'b0 ;
  assign n10174 = n6067 & ~n10173 ;
  assign n10175 = n10174 ^ n6525 ^ 1'b0 ;
  assign n10176 = n1726 | n4793 ;
  assign n10177 = n2092 & ~n10176 ;
  assign n10178 = n10175 & n10177 ;
  assign n10179 = n3533 & n6083 ;
  assign n10180 = n10179 ^ n1520 ^ 1'b0 ;
  assign n10181 = ( n3137 & ~n3670 ) | ( n3137 & n4000 ) | ( ~n3670 & n4000 ) ;
  assign n10182 = ( ~n5391 & n8865 ) | ( ~n5391 & n10181 ) | ( n8865 & n10181 ) ;
  assign n10183 = n6282 ^ n61 ^ 1'b0 ;
  assign n10184 = n910 | n10183 ;
  assign n10185 = n451 & ~n10184 ;
  assign n10186 = n1338 & ~n10185 ;
  assign n10187 = n6702 & n10186 ;
  assign n10188 = n6075 ^ n302 ^ 1'b0 ;
  assign n10189 = n7759 ^ n6441 ^ 1'b0 ;
  assign n10190 = ~n5902 & n9401 ;
  assign n10191 = n10190 ^ n3779 ^ 1'b0 ;
  assign n10192 = ~n3358 & n5375 ;
  assign n10193 = n551 & n10192 ;
  assign n10194 = ( n3695 & n4348 ) | ( n3695 & ~n9261 ) | ( n4348 & ~n9261 ) ;
  assign n10195 = n10194 ^ n8441 ^ 1'b0 ;
  assign n10196 = n96 & ~n898 ;
  assign n10197 = n5554 & n5995 ;
  assign n10198 = n365 & ~n3188 ;
  assign n10199 = n3285 | n4082 ;
  assign n10200 = ~n2267 & n10199 ;
  assign n10201 = ~n199 & n10200 ;
  assign n10202 = n6359 & ~n10201 ;
  assign n10203 = n9381 & n10202 ;
  assign n10204 = n919 & ~n7179 ;
  assign n10205 = n10204 ^ n4328 ^ 1'b0 ;
  assign n10206 = n5627 ^ n1530 ^ 1'b0 ;
  assign n10207 = ~n6931 & n10206 ;
  assign n10208 = n9938 ^ n3047 ^ 1'b0 ;
  assign n10209 = n8975 ^ n1939 ^ 1'b0 ;
  assign n10210 = n5786 & ~n10209 ;
  assign n10211 = n2227 | n4792 ;
  assign n10212 = ~n778 & n10211 ;
  assign n10213 = n8778 ^ n6950 ^ 1'b0 ;
  assign n10214 = n3011 ^ n382 ^ 1'b0 ;
  assign n10215 = ~n8459 & n10214 ;
  assign n10216 = n5080 ^ n2802 ^ 1'b0 ;
  assign n10217 = n10215 & ~n10216 ;
  assign n10218 = n5023 & n6278 ;
  assign n10219 = n6730 & n10218 ;
  assign n10220 = ~n10217 & n10219 ;
  assign n10221 = n8531 & ~n10220 ;
  assign n10222 = n3231 ^ n2243 ^ 1'b0 ;
  assign n10223 = n10222 ^ n8507 ^ 1'b0 ;
  assign n10224 = n10012 ^ n4521 ^ 1'b0 ;
  assign n10225 = n4537 & n10224 ;
  assign n10226 = n8655 ^ n6633 ^ 1'b0 ;
  assign n10227 = n3703 & n10226 ;
  assign n10228 = ~n7532 & n10227 ;
  assign n10229 = ~n388 & n7048 ;
  assign n10230 = ~n4053 & n10229 ;
  assign n10231 = n2460 | n5569 ;
  assign n10232 = n831 & ~n10231 ;
  assign n10233 = ~n6298 & n7600 ;
  assign n10234 = ~n3487 & n10233 ;
  assign n10235 = n3998 | n8331 ;
  assign n10236 = n8247 ^ n4688 ^ 1'b0 ;
  assign n10237 = ~n8470 & n10236 ;
  assign n10238 = n6716 & n10237 ;
  assign n10239 = n1432 | n5067 ;
  assign n10240 = ~n2062 & n6075 ;
  assign n10241 = n10240 ^ n7335 ^ 1'b0 ;
  assign n10242 = n8134 ^ n4444 ^ x10 ;
  assign n10243 = n2668 & ~n3369 ;
  assign n10244 = ~n2569 & n10243 ;
  assign n10245 = n8725 ^ n8282 ^ n1700 ;
  assign n10246 = ~n484 & n4536 ;
  assign n10247 = n10246 ^ n6006 ^ n4364 ;
  assign n10248 = ~n1152 & n10247 ;
  assign n10249 = ~n3062 & n9187 ;
  assign n10250 = n2282 ^ n680 ^ 1'b0 ;
  assign n10251 = ~n4359 & n10250 ;
  assign n10252 = ~n1238 & n1989 ;
  assign n10253 = ~n3510 & n10252 ;
  assign n10254 = ( ~x10 & n10251 ) | ( ~x10 & n10253 ) | ( n10251 & n10253 ) ;
  assign n10255 = n10254 ^ n5837 ^ 1'b0 ;
  assign n10256 = n1802 & ~n10255 ;
  assign n10257 = n4138 | n10256 ;
  assign n10258 = n543 & n721 ;
  assign n10259 = n5929 & n10258 ;
  assign n10261 = n4012 ^ n2387 ^ 1'b0 ;
  assign n10262 = n3851 & n10261 ;
  assign n10260 = ~n2726 & n5796 ;
  assign n10263 = n10262 ^ n10260 ^ 1'b0 ;
  assign n10264 = n2155 ^ n1750 ^ 1'b0 ;
  assign n10265 = n10264 ^ n6442 ^ 1'b0 ;
  assign n10266 = n7494 ^ n667 ^ 1'b0 ;
  assign n10267 = n3314 | n10266 ;
  assign n10268 = n6542 ^ n4539 ^ 1'b0 ;
  assign n10269 = n4754 ^ n4005 ^ n1984 ;
  assign n10270 = ~n3971 & n10269 ;
  assign n10271 = n10270 ^ n2848 ^ 1'b0 ;
  assign n10272 = n2919 | n9037 ;
  assign n10273 = n7294 & ~n10272 ;
  assign n10274 = n2855 & n10273 ;
  assign n10275 = ( n7960 & n8815 ) | ( n7960 & ~n9776 ) | ( n8815 & ~n9776 ) ;
  assign n10276 = n6871 & ~n7200 ;
  assign n10277 = n10276 ^ n8714 ^ 1'b0 ;
  assign n10278 = n146 & n2095 ;
  assign n10279 = n6492 ^ n592 ^ 1'b0 ;
  assign n10280 = n10278 | n10279 ;
  assign n10281 = n8342 ^ n4792 ^ 1'b0 ;
  assign n10282 = ( n342 & n463 ) | ( n342 & ~n5224 ) | ( n463 & ~n5224 ) ;
  assign n10283 = ~n1523 & n10282 ;
  assign n10284 = n1377 ^ n667 ^ 1'b0 ;
  assign n10285 = ~n4042 & n4588 ;
  assign n10286 = ~n4479 & n10285 ;
  assign n10287 = n3539 | n7627 ;
  assign n10288 = n4102 | n10287 ;
  assign n10289 = n3852 & ~n9321 ;
  assign n10290 = ~n85 & n4101 ;
  assign n10291 = n10290 ^ n4761 ^ 1'b0 ;
  assign n10292 = n83 & n10291 ;
  assign n10293 = ~n4095 & n10292 ;
  assign n10294 = n10293 ^ n6559 ^ 1'b0 ;
  assign n10295 = n3242 & n7391 ;
  assign n10296 = n7448 ^ n2028 ^ 1'b0 ;
  assign n10297 = ~n3434 & n10296 ;
  assign n10298 = ( n4666 & n4734 ) | ( n4666 & n7187 ) | ( n4734 & n7187 ) ;
  assign n10299 = ~n7969 & n10298 ;
  assign n10300 = n1144 & n3410 ;
  assign n10301 = n10300 ^ n2335 ^ 1'b0 ;
  assign n10302 = ~n10299 & n10301 ;
  assign n10303 = n4048 ^ n2225 ^ 1'b0 ;
  assign n10304 = n525 & ~n1419 ;
  assign n10305 = n3875 & n10304 ;
  assign n10306 = n4510 | n10305 ;
  assign n10307 = n9043 ^ n7237 ^ 1'b0 ;
  assign n10310 = n3028 & n3080 ;
  assign n10311 = n10310 ^ n1835 ^ 1'b0 ;
  assign n10308 = ~n205 & n2632 ;
  assign n10309 = n10308 ^ n4476 ^ 1'b0 ;
  assign n10312 = n10311 ^ n10309 ^ 1'b0 ;
  assign n10313 = n5001 & n10312 ;
  assign n10314 = ~n5606 & n10313 ;
  assign n10315 = n3716 ^ n844 ^ n25 ;
  assign n10316 = n7731 ^ n511 ^ 1'b0 ;
  assign n10317 = n1377 & n10316 ;
  assign n10319 = ( n167 & ~n533 ) | ( n167 & n2973 ) | ( ~n533 & n2973 ) ;
  assign n10320 = ( ~n1712 & n4537 ) | ( ~n1712 & n10319 ) | ( n4537 & n10319 ) ;
  assign n10318 = n3837 ^ n1363 ^ 1'b0 ;
  assign n10321 = n10320 ^ n10318 ^ 1'b0 ;
  assign n10322 = ~n1090 & n10000 ;
  assign n10323 = n3961 | n10322 ;
  assign n10324 = n9970 ^ n9371 ^ 1'b0 ;
  assign n10325 = n4280 & n10324 ;
  assign n10326 = n9535 & n10325 ;
  assign n10327 = n10326 ^ n3202 ^ 1'b0 ;
  assign n10328 = ~n987 & n3086 ;
  assign n10329 = n8062 & n10328 ;
  assign n10330 = n1449 & n4141 ;
  assign n10332 = n4632 & ~n4650 ;
  assign n10333 = n10332 ^ n575 ^ 1'b0 ;
  assign n10331 = n9047 | n9055 ;
  assign n10334 = n10333 ^ n10331 ^ 1'b0 ;
  assign n10335 = ~n10330 & n10334 ;
  assign n10338 = n619 | n7949 ;
  assign n10336 = n2444 ^ n1063 ^ 1'b0 ;
  assign n10337 = n8230 | n10336 ;
  assign n10339 = n10338 ^ n10337 ^ 1'b0 ;
  assign n10340 = n9258 | n10339 ;
  assign n10342 = n4014 ^ n1538 ^ 1'b0 ;
  assign n10341 = n4734 & ~n6441 ;
  assign n10343 = n10342 ^ n10341 ^ 1'b0 ;
  assign n10344 = n10239 ^ n2665 ^ 1'b0 ;
  assign n10345 = n8822 & ~n10344 ;
  assign n10346 = n5647 ^ n3212 ^ 1'b0 ;
  assign n10347 = n3369 | n10346 ;
  assign n10351 = n1264 & n2647 ;
  assign n10348 = n802 & ~n2228 ;
  assign n10349 = n8983 ^ n4029 ^ 1'b0 ;
  assign n10350 = ~n10348 & n10349 ;
  assign n10352 = n10351 ^ n10350 ^ 1'b0 ;
  assign n10353 = n3957 & n7668 ;
  assign n10354 = ~n10352 & n10353 ;
  assign n10356 = n6705 ^ n4899 ^ 1'b0 ;
  assign n10355 = ~n98 & n4166 ;
  assign n10357 = n10356 ^ n10355 ^ 1'b0 ;
  assign n10358 = n2318 ^ n2247 ^ 1'b0 ;
  assign n10359 = n3178 & ~n10358 ;
  assign n10360 = n10359 ^ n725 ^ 1'b0 ;
  assign n10361 = ~n10357 & n10360 ;
  assign n10362 = n509 ^ n430 ^ 1'b0 ;
  assign n10363 = n10362 ^ n8870 ^ n6216 ;
  assign n10364 = n2551 ^ n2173 ^ n722 ;
  assign n10365 = n10364 ^ n7908 ^ n5829 ;
  assign n10366 = ~n801 & n5084 ;
  assign n10367 = ~n113 & n3216 ;
  assign n10368 = ~n1504 & n4313 ;
  assign n10369 = n3114 ^ n1726 ^ 1'b0 ;
  assign n10370 = n10185 ^ n2268 ^ 1'b0 ;
  assign n10371 = n5215 & ~n10370 ;
  assign n10372 = n10371 ^ n4282 ^ 1'b0 ;
  assign n10373 = n6200 ^ n2252 ^ 1'b0 ;
  assign n10374 = n7679 & n10373 ;
  assign n10375 = n10372 & n10374 ;
  assign n10376 = n10375 ^ n3108 ^ 1'b0 ;
  assign n10377 = n5949 & ~n9771 ;
  assign n10378 = n473 | n6401 ;
  assign n10379 = ~n7823 & n10378 ;
  assign n10380 = n10377 | n10379 ;
  assign n10381 = n10380 ^ n8543 ^ 1'b0 ;
  assign n10384 = n795 | n4188 ;
  assign n10385 = n6326 | n10384 ;
  assign n10382 = ~n2492 & n6526 ;
  assign n10383 = n5654 & n10382 ;
  assign n10386 = n10385 ^ n10383 ^ 1'b0 ;
  assign n10387 = n7823 | n10386 ;
  assign n10388 = n6049 ^ n4353 ^ 1'b0 ;
  assign n10389 = n10388 ^ n302 ^ 1'b0 ;
  assign n10390 = n1876 & ~n9680 ;
  assign n10391 = n10390 ^ n4009 ^ 1'b0 ;
  assign n10392 = n9798 ^ n9483 ^ n2246 ;
  assign n10393 = n8441 | n10392 ;
  assign n10394 = n61 & ~n1910 ;
  assign n10395 = n10394 ^ n5257 ^ 1'b0 ;
  assign n10396 = ~n133 & n745 ;
  assign n10397 = n3823 & ~n10396 ;
  assign n10398 = n10395 | n10397 ;
  assign n10399 = n10398 ^ n8491 ^ 1'b0 ;
  assign n10402 = n695 ^ n152 ^ 1'b0 ;
  assign n10403 = ~n2415 & n10402 ;
  assign n10404 = n10403 ^ n4856 ^ 1'b0 ;
  assign n10400 = n2246 & ~n3021 ;
  assign n10401 = ~n3453 & n10400 ;
  assign n10405 = n10404 ^ n10401 ^ 1'b0 ;
  assign n10406 = n997 | n8625 ;
  assign n10407 = n6518 & ~n7958 ;
  assign n10408 = n497 | n6922 ;
  assign n10409 = n10408 ^ n5472 ^ 1'b0 ;
  assign n10410 = n5936 & n6552 ;
  assign n10411 = ~n10409 & n10410 ;
  assign n10412 = n5328 & ~n6258 ;
  assign n10413 = n7247 ^ n1416 ^ 1'b0 ;
  assign n10414 = n8689 & n10413 ;
  assign n10415 = ( n3729 & n4547 ) | ( n3729 & ~n10414 ) | ( n4547 & ~n10414 ) ;
  assign n10416 = n142 | n1918 ;
  assign n10417 = n3811 | n10416 ;
  assign n10418 = n5101 ^ n4489 ^ n3688 ;
  assign n10419 = n10418 ^ n2754 ^ 1'b0 ;
  assign n10420 = n10417 & ~n10419 ;
  assign n10421 = n6542 ^ n4814 ^ n2288 ;
  assign n10422 = n5334 ^ n406 ^ 1'b0 ;
  assign n10423 = n10421 & n10422 ;
  assign n10424 = n4814 & ~n10264 ;
  assign n10425 = n7981 & n10424 ;
  assign n10426 = n162 & n1284 ;
  assign n10427 = ~n248 & n701 ;
  assign n10428 = n6203 & n10427 ;
  assign n10429 = n1685 & ~n10428 ;
  assign n10430 = n4648 & n10429 ;
  assign n10431 = n2564 & n10430 ;
  assign n10432 = n6363 & ~n8847 ;
  assign n10433 = n911 | n7930 ;
  assign n10434 = ~n3295 & n3307 ;
  assign n10435 = n2494 & n8340 ;
  assign n10436 = ~n10434 & n10435 ;
  assign n10437 = n9322 ^ n4331 ^ 1'b0 ;
  assign n10438 = ~n124 & n695 ;
  assign n10439 = ( n2614 & n6590 ) | ( n2614 & n10438 ) | ( n6590 & n10438 ) ;
  assign n10440 = ~n1000 & n3982 ;
  assign n10441 = n4641 & n10440 ;
  assign n10442 = n4685 & ~n10441 ;
  assign n10443 = n10442 ^ n703 ^ 1'b0 ;
  assign n10444 = n1316 & n9170 ;
  assign n10445 = ~n6800 & n10444 ;
  assign n10446 = ~n184 & n3390 ;
  assign n10447 = ~n7781 & n10446 ;
  assign n10449 = ~n5645 & n8176 ;
  assign n10448 = n1025 & ~n5413 ;
  assign n10450 = n10449 ^ n10448 ^ 1'b0 ;
  assign n10451 = ~n5119 & n10450 ;
  assign n10452 = n9322 ^ n6358 ^ 1'b0 ;
  assign n10453 = n10452 ^ n7820 ^ 1'b0 ;
  assign n10454 = n2953 & n10453 ;
  assign n10455 = n10454 ^ n7059 ^ 1'b0 ;
  assign n10456 = n2721 & n10455 ;
  assign n10457 = ~n5821 & n10456 ;
  assign n10458 = n2390 & ~n3975 ;
  assign n10459 = n10458 ^ n9416 ^ 1'b0 ;
  assign n10460 = n2875 | n10459 ;
  assign n10461 = ~n326 & n10460 ;
  assign n10462 = n10461 ^ n6384 ^ 1'b0 ;
  assign n10463 = ~n378 & n2197 ;
  assign n10464 = n842 | n1003 ;
  assign n10465 = n1050 | n10464 ;
  assign n10466 = n10465 ^ n2730 ^ 1'b0 ;
  assign n10467 = n10466 ^ n10366 ^ n6758 ;
  assign n10468 = ~n10463 & n10467 ;
  assign n10469 = n4496 ^ n4472 ^ 1'b0 ;
  assign n10470 = ~n2776 & n10469 ;
  assign n10471 = n4665 ^ n2004 ^ 1'b0 ;
  assign n10472 = n1633 & n10471 ;
  assign n10473 = n502 & ~n10472 ;
  assign n10474 = n10473 ^ n3954 ^ 1'b0 ;
  assign n10475 = n1570 | n10474 ;
  assign n10476 = n4335 | n7316 ;
  assign n10477 = ( ~n2112 & n10475 ) | ( ~n2112 & n10476 ) | ( n10475 & n10476 ) ;
  assign n10478 = n2925 & n3930 ;
  assign n10479 = ~n2628 & n10478 ;
  assign n10480 = n10477 | n10479 ;
  assign n10481 = n6404 ^ n4875 ^ n4033 ;
  assign n10482 = n8862 ^ n214 ^ 1'b0 ;
  assign n10483 = n10481 & ~n10482 ;
  assign n10484 = n2571 ^ n1269 ^ n211 ;
  assign n10485 = n704 & n828 ;
  assign n10486 = n7981 ^ n2133 ^ 1'b0 ;
  assign n10487 = n10486 ^ n5229 ^ 1'b0 ;
  assign n10488 = n10485 & n10487 ;
  assign n10489 = n3343 & ~n6004 ;
  assign n10490 = n10314 ^ n2596 ^ 1'b0 ;
  assign n10491 = n179 | n10490 ;
  assign n10492 = n5773 & n6238 ;
  assign n10493 = ( ~n1620 & n5274 ) | ( ~n1620 & n10492 ) | ( n5274 & n10492 ) ;
  assign n10494 = n8494 ^ n3453 ^ 1'b0 ;
  assign n10495 = n2628 & ~n10494 ;
  assign n10496 = n778 | n5911 ;
  assign n10497 = n3450 | n10496 ;
  assign n10498 = n2112 | n10497 ;
  assign n10499 = n10498 ^ n3167 ^ 1'b0 ;
  assign n10500 = n3020 ^ n2572 ^ 1'b0 ;
  assign n10501 = n4001 & ~n10500 ;
  assign n10502 = n7282 ^ n2161 ^ 1'b0 ;
  assign n10503 = n795 | n10502 ;
  assign n10504 = n10503 ^ n2134 ^ 1'b0 ;
  assign n10505 = n10504 ^ n5799 ^ n3847 ;
  assign n10506 = n919 & n1355 ;
  assign n10507 = ~n488 & n10506 ;
  assign n10508 = n10507 ^ n3853 ^ n3259 ;
  assign n10509 = n729 & n1699 ;
  assign n10510 = ~n10508 & n10509 ;
  assign n10511 = ( n447 & ~n2806 ) | ( n447 & n4091 ) | ( ~n2806 & n4091 ) ;
  assign n10512 = n10511 ^ n8552 ^ 1'b0 ;
  assign n10513 = n9114 & ~n10512 ;
  assign n10514 = n10510 & n10513 ;
  assign n10515 = n978 & ~n9883 ;
  assign n10516 = n10515 ^ n8916 ^ 1'b0 ;
  assign n10520 = n7516 ^ n4051 ^ 1'b0 ;
  assign n10517 = n3990 | n6396 ;
  assign n10518 = n1789 | n10517 ;
  assign n10519 = n10518 ^ n9202 ^ 1'b0 ;
  assign n10521 = n10520 ^ n10519 ^ n1284 ;
  assign n10522 = n2442 & n5733 ;
  assign n10523 = ~n4578 & n5610 ;
  assign n10524 = n10523 ^ n9319 ^ 1'b0 ;
  assign n10525 = n557 & ~n894 ;
  assign n10526 = ~n4463 & n10525 ;
  assign n10527 = n282 & n10526 ;
  assign n10528 = n7964 ^ n7112 ^ n4671 ;
  assign n10529 = n213 | n4597 ;
  assign n10530 = n2393 ^ n1024 ^ 1'b0 ;
  assign n10531 = n5594 ^ n4902 ^ 1'b0 ;
  assign n10532 = n10531 ^ n10498 ^ 1'b0 ;
  assign n10533 = n10532 ^ n4111 ^ n738 ;
  assign n10534 = ~n3710 & n6215 ;
  assign n10535 = n2549 & ~n10463 ;
  assign n10536 = ~n1550 & n10535 ;
  assign n10537 = n3662 | n5637 ;
  assign n10538 = n10537 ^ n2901 ^ 1'b0 ;
  assign n10539 = n722 | n8815 ;
  assign n10540 = ~n1832 & n6635 ;
  assign n10541 = ~n4359 & n10540 ;
  assign n10542 = n10541 ^ n49 ^ 1'b0 ;
  assign n10543 = n10542 ^ n6756 ^ n1750 ;
  assign n10544 = n846 | n1513 ;
  assign n10545 = n2765 & n10544 ;
  assign n10546 = n1066 & ~n6774 ;
  assign n10547 = n10546 ^ n6988 ^ 1'b0 ;
  assign n10548 = ~n10232 & n10547 ;
  assign n10549 = n910 ^ n213 ^ 1'b0 ;
  assign n10550 = n10549 ^ n5757 ^ 1'b0 ;
  assign n10551 = n10550 ^ n4573 ^ 1'b0 ;
  assign n10552 = n7931 | n10551 ;
  assign n10553 = n10552 ^ n290 ^ 1'b0 ;
  assign n10554 = n69 & n2277 ;
  assign n10555 = n10554 ^ n4132 ^ 1'b0 ;
  assign n10556 = ~n5825 & n10555 ;
  assign n10557 = n841 | n1539 ;
  assign n10558 = n10556 | n10557 ;
  assign n10559 = n10553 & n10558 ;
  assign n10560 = n4637 ^ n3777 ^ n1987 ;
  assign n10561 = n4519 ^ n3110 ^ 1'b0 ;
  assign n10562 = ~n3753 & n10561 ;
  assign n10563 = ~n10117 & n10562 ;
  assign n10564 = ~n8635 & n10563 ;
  assign n10565 = n4366 | n7463 ;
  assign n10566 = n91 & ~n3299 ;
  assign n10567 = n473 & n10566 ;
  assign n10568 = n10567 ^ n495 ^ 1'b0 ;
  assign n10569 = n9083 & ~n10568 ;
  assign n10570 = n10569 ^ n5331 ^ 1'b0 ;
  assign n10574 = ~n1014 & n1814 ;
  assign n10575 = n9088 & n10574 ;
  assign n10579 = n770 | n6099 ;
  assign n10576 = n1010 & ~n4248 ;
  assign n10577 = n10576 ^ n3848 ^ 1'b0 ;
  assign n10578 = n6043 | n10577 ;
  assign n10580 = n10579 ^ n10578 ^ 1'b0 ;
  assign n10581 = ( ~n5684 & n10575 ) | ( ~n5684 & n10580 ) | ( n10575 & n10580 ) ;
  assign n10571 = ~n362 & n1721 ;
  assign n10572 = ~n9113 & n10571 ;
  assign n10573 = n598 & ~n10572 ;
  assign n10582 = n10581 ^ n10573 ^ 1'b0 ;
  assign n10583 = n4038 ^ n1809 ^ 1'b0 ;
  assign n10584 = ~n2946 & n10583 ;
  assign n10585 = ~n7174 & n10584 ;
  assign n10586 = n4446 | n10585 ;
  assign n10587 = ~n8745 & n8933 ;
  assign n10588 = n4787 & ~n6151 ;
  assign n10589 = n10588 ^ n3167 ^ 1'b0 ;
  assign n10590 = n832 & n10589 ;
  assign n10591 = n10590 ^ n8577 ^ 1'b0 ;
  assign n10592 = n1327 & n10591 ;
  assign n10593 = n6937 | n10592 ;
  assign n10594 = ~n5295 & n8451 ;
  assign n10595 = n10594 ^ n2772 ^ 1'b0 ;
  assign n10596 = n10595 ^ n8683 ^ 1'b0 ;
  assign n10597 = n10297 ^ n7702 ^ 1'b0 ;
  assign n10598 = n4671 & ~n10597 ;
  assign n10599 = n2134 & n7581 ;
  assign n10600 = n2719 & n10599 ;
  assign n10601 = n1802 ^ n439 ^ 1'b0 ;
  assign n10602 = n3298 ^ n995 ^ 1'b0 ;
  assign n10603 = ~n3050 & n10602 ;
  assign n10604 = ( n1951 & n5616 ) | ( n1951 & n10603 ) | ( n5616 & n10603 ) ;
  assign n10605 = ~n5286 & n10374 ;
  assign n10606 = ~n10604 & n10605 ;
  assign n10607 = n4989 ^ n1050 ^ 1'b0 ;
  assign n10608 = n7135 ^ n6868 ^ 1'b0 ;
  assign n10609 = n10607 & ~n10608 ;
  assign n10611 = n2419 | n7534 ;
  assign n10610 = n1510 ^ n67 ^ 1'b0 ;
  assign n10612 = n10611 ^ n10610 ^ 1'b0 ;
  assign n10615 = n2749 & n5435 ;
  assign n10616 = n10615 ^ n996 ^ 1'b0 ;
  assign n10613 = n489 ^ n299 ^ 1'b0 ;
  assign n10614 = n5008 | n10613 ;
  assign n10617 = n10616 ^ n10614 ^ 1'b0 ;
  assign n10618 = n214 & ~n10617 ;
  assign n10619 = n7520 ^ n4002 ^ 1'b0 ;
  assign n10620 = n3486 & n10619 ;
  assign n10621 = n9330 ^ n4550 ^ 1'b0 ;
  assign n10622 = ~n1615 & n10621 ;
  assign n10623 = n7972 ^ n2785 ^ 1'b0 ;
  assign n10624 = n571 | n10623 ;
  assign n10625 = n798 & n2211 ;
  assign n10626 = n4044 & n10625 ;
  assign n10627 = n10626 ^ n8230 ^ 1'b0 ;
  assign n10628 = n10624 | n10627 ;
  assign n10629 = n2440 ^ n1434 ^ 1'b0 ;
  assign n10630 = n1347 & ~n10629 ;
  assign n10631 = ~n1779 & n10630 ;
  assign n10632 = n10628 & n10631 ;
  assign n10636 = n1351 & ~n7490 ;
  assign n10637 = n2796 & n10636 ;
  assign n10633 = n565 ^ n552 ^ 1'b0 ;
  assign n10634 = ~n5383 & n10633 ;
  assign n10635 = n5297 | n10634 ;
  assign n10638 = n10637 ^ n10635 ^ n8578 ;
  assign n10639 = n749 & n9247 ;
  assign n10640 = n10639 ^ n2367 ^ 1'b0 ;
  assign n10641 = n10640 ^ n4020 ^ n4010 ;
  assign n10642 = n3049 | n9272 ;
  assign n10643 = n652 & n2331 ;
  assign n10644 = n10643 ^ n2794 ^ 1'b0 ;
  assign n10645 = ( ~n1383 & n7000 ) | ( ~n1383 & n10644 ) | ( n7000 & n10644 ) ;
  assign n10646 = n8608 & n9209 ;
  assign n10647 = ( n4108 & n10645 ) | ( n4108 & n10646 ) | ( n10645 & n10646 ) ;
  assign n10648 = n10642 & n10647 ;
  assign n10649 = ~n10641 & n10648 ;
  assign n10650 = n8029 ^ n6248 ^ 1'b0 ;
  assign n10651 = n10215 & ~n10650 ;
  assign n10652 = n10651 ^ n3449 ^ 1'b0 ;
  assign n10653 = ~n1085 & n4296 ;
  assign n10654 = n4372 ^ n902 ^ 1'b0 ;
  assign n10655 = n1895 & n7541 ;
  assign n10656 = n10654 & n10655 ;
  assign n10657 = ( n5866 & n7744 ) | ( n5866 & ~n8788 ) | ( n7744 & ~n8788 ) ;
  assign n10658 = n6367 & ~n8606 ;
  assign n10659 = n2883 ^ n2288 ^ 1'b0 ;
  assign n10660 = n7520 | n10659 ;
  assign n10661 = n6777 | n10660 ;
  assign n10662 = n10661 ^ n9277 ^ 1'b0 ;
  assign n10663 = n1666 & n2602 ;
  assign n10664 = n10663 ^ n2139 ^ 1'b0 ;
  assign n10665 = n5393 & n10664 ;
  assign n10666 = n8611 & n10665 ;
  assign n10667 = n3187 & n10666 ;
  assign n10668 = n7332 ^ n6832 ^ 1'b0 ;
  assign n10669 = n841 & ~n1205 ;
  assign n10670 = ~n6602 & n10669 ;
  assign n10671 = n10303 & ~n10670 ;
  assign n10672 = n10668 & n10671 ;
  assign n10673 = ( n2317 & n3917 ) | ( n2317 & ~n7552 ) | ( n3917 & ~n7552 ) ;
  assign n10674 = n6702 ^ n6591 ^ 1'b0 ;
  assign n10675 = ~n552 & n1374 ;
  assign n10676 = ( n3807 & n5277 ) | ( n3807 & n10675 ) | ( n5277 & n10675 ) ;
  assign n10677 = ~n8453 & n10676 ;
  assign n10678 = ~n4298 & n10677 ;
  assign n10680 = n4843 ^ n4644 ^ 1'b0 ;
  assign n10681 = ~n3663 & n10680 ;
  assign n10679 = n1914 & n8451 ;
  assign n10682 = n10681 ^ n10679 ^ 1'b0 ;
  assign n10683 = n119 | n6799 ;
  assign n10684 = n10683 ^ n6825 ^ 1'b0 ;
  assign n10685 = n249 & ~n8915 ;
  assign n10686 = n3721 & n10685 ;
  assign n10687 = n10686 ^ n2517 ^ n129 ;
  assign n10688 = n10687 ^ n4006 ^ x0 ;
  assign n10691 = n673 & n6947 ;
  assign n10689 = ( ~n204 & n216 ) | ( ~n204 & n5511 ) | ( n216 & n5511 ) ;
  assign n10690 = ~n1172 & n10689 ;
  assign n10692 = n10691 ^ n10690 ^ 1'b0 ;
  assign n10693 = n4034 ^ n604 ^ 1'b0 ;
  assign n10694 = n2404 & n10693 ;
  assign n10695 = n6045 | n10128 ;
  assign n10696 = ( ~n6042 & n10694 ) | ( ~n6042 & n10695 ) | ( n10694 & n10695 ) ;
  assign n10697 = n83 & n6635 ;
  assign n10698 = n6474 & n10697 ;
  assign n10699 = n4944 & ~n10698 ;
  assign n10700 = ~n9252 & n10699 ;
  assign n10701 = n10696 & n10700 ;
  assign n10702 = n6729 ^ n5222 ^ 1'b0 ;
  assign n10703 = n3201 | n10702 ;
  assign n10704 = n5367 & n8135 ;
  assign n10705 = n10704 ^ n5684 ^ 1'b0 ;
  assign n10706 = n8451 ^ n1507 ^ 1'b0 ;
  assign n10707 = n74 & n4226 ;
  assign n10708 = n10707 ^ n4077 ^ 1'b0 ;
  assign n10709 = n10708 ^ n6392 ^ 1'b0 ;
  assign n10710 = n10706 & n10709 ;
  assign n10711 = n5170 & n10710 ;
  assign n10712 = n2658 ^ n1050 ^ 1'b0 ;
  assign n10713 = ~n3075 & n10712 ;
  assign n10714 = n6777 | n8545 ;
  assign n10715 = n8103 | n10714 ;
  assign n10716 = n3341 & ~n10715 ;
  assign n10717 = n1040 | n2815 ;
  assign n10718 = n5613 ^ n688 ^ 1'b0 ;
  assign n10719 = ~n10717 & n10718 ;
  assign n10720 = n4250 & ~n4808 ;
  assign n10721 = n1667 & ~n8706 ;
  assign n10725 = n4954 ^ n3592 ^ 1'b0 ;
  assign n10726 = ~n5044 & n10725 ;
  assign n10722 = n874 ^ n136 ^ 1'b0 ;
  assign n10723 = n1732 & n10722 ;
  assign n10724 = ~n1010 & n10723 ;
  assign n10727 = n10726 ^ n10724 ^ 1'b0 ;
  assign n10728 = n10721 & ~n10727 ;
  assign n10729 = ~n5046 & n6035 ;
  assign n10730 = ~n2932 & n10729 ;
  assign n10731 = ( n115 & n4576 ) | ( n115 & n10730 ) | ( n4576 & n10730 ) ;
  assign n10732 = n6401 | n9765 ;
  assign n10733 = n9819 & ~n10732 ;
  assign n10734 = n3772 | n8414 ;
  assign n10735 = n10734 ^ n1099 ^ 1'b0 ;
  assign n10736 = n8550 | n9679 ;
  assign n10737 = n10736 ^ n1744 ^ 1'b0 ;
  assign n10738 = ( n2206 & ~n2763 ) | ( n2206 & n5834 ) | ( ~n2763 & n5834 ) ;
  assign n10739 = n10738 ^ n2262 ^ n1453 ;
  assign n10740 = ~n3054 & n5613 ;
  assign n10741 = n2539 & n10740 ;
  assign n10742 = n10741 ^ n5106 ^ 1'b0 ;
  assign n10743 = n10660 | n10742 ;
  assign n10744 = n7073 & n7916 ;
  assign n10745 = n10744 ^ n5968 ^ 1'b0 ;
  assign n10746 = n164 & n5689 ;
  assign n10747 = n10746 ^ n129 ^ 1'b0 ;
  assign n10748 = n10747 ^ n3592 ^ 1'b0 ;
  assign n10751 = n7741 | n8273 ;
  assign n10752 = n6238 & ~n10751 ;
  assign n10749 = n1816 ^ n732 ^ 1'b0 ;
  assign n10750 = n9388 | n10749 ;
  assign n10753 = n10752 ^ n10750 ^ 1'b0 ;
  assign n10754 = n314 | n4386 ;
  assign n10755 = ~n4419 & n10754 ;
  assign n10756 = ~n8850 & n10755 ;
  assign n10757 = ~n333 & n2614 ;
  assign n10758 = n10757 ^ n6229 ^ 1'b0 ;
  assign n10759 = n10758 ^ n4837 ^ 1'b0 ;
  assign n10760 = n4573 & n5692 ;
  assign n10761 = ~n822 & n10760 ;
  assign n10762 = ~n970 & n3507 ;
  assign n10763 = n2843 | n6210 ;
  assign n10764 = n10763 ^ n4159 ^ n3797 ;
  assign n10766 = n890 & n5227 ;
  assign n10765 = n664 | n8695 ;
  assign n10767 = n10766 ^ n10765 ^ 1'b0 ;
  assign n10768 = n307 & ~n2352 ;
  assign n10769 = ( n667 & n3998 ) | ( n667 & n10768 ) | ( n3998 & n10768 ) ;
  assign n10770 = n10769 ^ n9112 ^ n800 ;
  assign n10772 = n6351 ^ n5258 ^ n765 ;
  assign n10771 = n1720 & ~n4139 ;
  assign n10773 = n10772 ^ n10771 ^ 1'b0 ;
  assign n10774 = ~n5935 & n10773 ;
  assign n10775 = n5021 & n10726 ;
  assign n10776 = n10775 ^ n3012 ^ 1'b0 ;
  assign n10777 = n4675 ^ n798 ^ 1'b0 ;
  assign n10778 = n1768 & ~n10777 ;
  assign n10779 = n7696 & ~n10351 ;
  assign n10780 = ~n10778 & n10779 ;
  assign n10781 = n5202 ^ n600 ^ 1'b0 ;
  assign n10782 = n5773 & ~n10781 ;
  assign n10783 = n2962 ^ n2680 ^ 1'b0 ;
  assign n10784 = n1334 & n10783 ;
  assign n10785 = ( n3277 & ~n4248 ) | ( n3277 & n10281 ) | ( ~n4248 & n10281 ) ;
  assign n10786 = n5973 | n6805 ;
  assign n10787 = n10786 ^ n9502 ^ 1'b0 ;
  assign n10788 = n10787 ^ n8779 ^ 1'b0 ;
  assign n10789 = ~n1150 & n8516 ;
  assign n10790 = n10789 ^ n5071 ^ 1'b0 ;
  assign n10791 = n4005 & ~n10790 ;
  assign n10792 = n10791 ^ n2883 ^ 1'b0 ;
  assign n10793 = n368 | n6456 ;
  assign n10794 = n8840 ^ n7463 ^ 1'b0 ;
  assign n10795 = n10793 | n10794 ;
  assign n10796 = n6872 | n6991 ;
  assign n10797 = n292 & ~n6322 ;
  assign n10798 = n492 & ~n10797 ;
  assign n10799 = n10798 ^ n3423 ^ 1'b0 ;
  assign n10800 = ~n6410 & n10799 ;
  assign n10801 = n10800 ^ n1984 ^ 1'b0 ;
  assign n10802 = ~n261 & n1637 ;
  assign n10803 = ~n6984 & n10802 ;
  assign n10804 = n1329 & ~n3634 ;
  assign n10805 = n1580 & ~n10465 ;
  assign n10806 = n10804 & ~n10805 ;
  assign n10807 = n1109 & n10806 ;
  assign n10808 = n725 ^ n286 ^ 1'b0 ;
  assign n10809 = ~n2185 & n10808 ;
  assign n10810 = n1117 & n1484 ;
  assign n10811 = ~n667 & n10810 ;
  assign n10812 = n10811 ^ n8919 ^ 1'b0 ;
  assign n10813 = n4704 & ~n5511 ;
  assign n10814 = ~n6941 & n10813 ;
  assign n10815 = n7414 ^ n2519 ^ 1'b0 ;
  assign n10816 = ( n61 & ~n1743 ) | ( n61 & n6919 ) | ( ~n1743 & n6919 ) ;
  assign n10817 = ( n1047 & ~n3582 ) | ( n1047 & n4599 ) | ( ~n3582 & n4599 ) ;
  assign n10818 = n2751 | n10817 ;
  assign n10819 = ~n7393 & n10818 ;
  assign n10820 = n536 & ~n5736 ;
  assign n10821 = n3447 | n5308 ;
  assign n10822 = n5270 | n10821 ;
  assign n10823 = ( ~n1327 & n4768 ) | ( ~n1327 & n10822 ) | ( n4768 & n10822 ) ;
  assign n10824 = ~n6431 & n10823 ;
  assign n10825 = n10820 & n10824 ;
  assign n10828 = n169 & n209 ;
  assign n10826 = n1322 & n3424 ;
  assign n10827 = n4251 & n10826 ;
  assign n10829 = n10828 ^ n10827 ^ 1'b0 ;
  assign n10830 = ~n614 & n8773 ;
  assign n10831 = n3137 & n10830 ;
  assign n10832 = n7604 | n10831 ;
  assign n10833 = n5122 | n10575 ;
  assign n10834 = n2010 & ~n10833 ;
  assign n10835 = n454 & n5574 ;
  assign n10836 = n10835 ^ n3780 ^ 1'b0 ;
  assign n10837 = n9727 ^ n6456 ^ n127 ;
  assign n10838 = n7668 & n10837 ;
  assign n10839 = ~n10836 & n10838 ;
  assign n10843 = n3760 ^ n646 ^ 1'b0 ;
  assign n10844 = n253 & ~n10843 ;
  assign n10840 = n3954 ^ n2388 ^ n521 ;
  assign n10841 = n4104 & ~n10840 ;
  assign n10842 = n2225 & ~n10841 ;
  assign n10845 = n10844 ^ n10842 ^ 1'b0 ;
  assign n10846 = n10845 ^ n3240 ^ 1'b0 ;
  assign n10847 = n6959 & ~n10846 ;
  assign n10848 = n1045 & ~n2818 ;
  assign n10849 = n1283 & ~n6441 ;
  assign n10850 = n10849 ^ n7696 ^ 1'b0 ;
  assign n10851 = n150 ^ x11 ^ 1'b0 ;
  assign n10852 = n6289 ^ n1941 ^ 1'b0 ;
  assign n10853 = n1327 & ~n4214 ;
  assign n10854 = n6321 & n10853 ;
  assign n10855 = n10852 & n10854 ;
  assign n10856 = n5300 & ~n10855 ;
  assign n10859 = ~n671 & n5524 ;
  assign n10860 = ~n3854 & n10859 ;
  assign n10857 = n83 | n3833 ;
  assign n10858 = n8249 & n10857 ;
  assign n10861 = n10860 ^ n10858 ^ 1'b0 ;
  assign n10862 = n4991 ^ n1173 ^ n390 ;
  assign n10863 = ~n2244 & n2973 ;
  assign n10864 = n4999 | n6856 ;
  assign n10865 = n667 & n6187 ;
  assign n10866 = n10864 & n10865 ;
  assign n10867 = n7066 ^ n755 ^ 1'b0 ;
  assign n10868 = n10866 | n10867 ;
  assign n10869 = n1728 | n10015 ;
  assign n10870 = n10869 ^ n9716 ^ 1'b0 ;
  assign n10871 = n1631 ^ x5 ^ 1'b0 ;
  assign n10872 = n3327 | n10871 ;
  assign n10873 = n10872 ^ n1455 ^ n831 ;
  assign n10874 = n10873 ^ n188 ^ 1'b0 ;
  assign n10875 = n6637 | n10874 ;
  assign n10876 = n10875 ^ n6208 ^ 1'b0 ;
  assign n10877 = n5745 | n10876 ;
  assign n10878 = n10877 ^ n2435 ^ 1'b0 ;
  assign n10879 = ~n2678 & n10878 ;
  assign n10880 = n5895 & n10879 ;
  assign n10881 = n792 & n10880 ;
  assign n10882 = n6619 ^ n1437 ^ 1'b0 ;
  assign n10883 = n8446 ^ n774 ^ 1'b0 ;
  assign n10884 = n2754 & n10634 ;
  assign n10885 = n4296 | n10884 ;
  assign n10886 = ( n105 & n1741 ) | ( n105 & ~n1767 ) | ( n1741 & ~n1767 ) ;
  assign n10887 = n3023 ^ n1973 ^ 1'b0 ;
  assign n10888 = n1454 | n10887 ;
  assign n10889 = n241 & ~n10888 ;
  assign n10890 = n10889 ^ n873 ^ 1'b0 ;
  assign n10891 = ( n251 & ~n10475 ) | ( n251 & n10890 ) | ( ~n10475 & n10890 ) ;
  assign n10892 = ( n2588 & n4903 ) | ( n2588 & n8219 ) | ( n4903 & n8219 ) ;
  assign n10893 = n1422 | n2444 ;
  assign n10894 = n10893 ^ n3121 ^ n924 ;
  assign n10895 = n4568 ^ n4000 ^ 1'b0 ;
  assign n10896 = n2229 ^ n1010 ^ 1'b0 ;
  assign n10897 = ~n6304 & n10896 ;
  assign n10898 = n10897 ^ n10188 ^ 1'b0 ;
  assign n10899 = n9059 & n10898 ;
  assign n10900 = n10895 & n10899 ;
  assign n10901 = n7187 & ~n8312 ;
  assign n10902 = ~n5599 & n5870 ;
  assign n10903 = n165 & n2933 ;
  assign n10904 = ( n3745 & n5841 ) | ( n3745 & ~n7641 ) | ( n5841 & ~n7641 ) ;
  assign n10905 = ( ~n423 & n4993 ) | ( ~n423 & n10904 ) | ( n4993 & n10904 ) ;
  assign n10906 = n1707 & n3461 ;
  assign n10907 = n10906 ^ n9163 ^ 1'b0 ;
  assign n10908 = n9186 ^ n7922 ^ 1'b0 ;
  assign n10909 = n10908 ^ n7050 ^ 1'b0 ;
  assign n10910 = ( n971 & ~n1276 ) | ( n971 & n5548 ) | ( ~n1276 & n5548 ) ;
  assign n10911 = n9293 ^ n4278 ^ n48 ;
  assign n10912 = n8868 & n10911 ;
  assign n10913 = n10912 ^ n451 ^ 1'b0 ;
  assign n10914 = n10913 ^ n4567 ^ 1'b0 ;
  assign n10915 = ( ~n365 & n3333 ) | ( ~n365 & n3822 ) | ( n3333 & n3822 ) ;
  assign n10916 = n2063 & n10915 ;
  assign n10917 = n10916 ^ n2971 ^ 1'b0 ;
  assign n10918 = n924 & n10917 ;
  assign n10919 = n10918 ^ n4025 ^ 1'b0 ;
  assign n10929 = n8144 ^ n3142 ^ 1'b0 ;
  assign n10920 = n688 & n1561 ;
  assign n10921 = ~n1561 & n10920 ;
  assign n10922 = n7893 | n8227 ;
  assign n10923 = n10922 ^ n3584 ^ 1'b0 ;
  assign n10924 = n4823 & n10923 ;
  assign n10925 = ~n10923 & n10924 ;
  assign n10926 = n10921 | n10925 ;
  assign n10927 = n10921 & ~n10926 ;
  assign n10928 = ~n5566 & n10927 ;
  assign n10930 = n10929 ^ n10928 ^ 1'b0 ;
  assign n10931 = n10919 & ~n10930 ;
  assign n10932 = n5610 ^ n2895 ^ 1'b0 ;
  assign n10933 = ~n3740 & n10932 ;
  assign n10934 = n8144 & n9024 ;
  assign n10935 = n5397 & ~n10934 ;
  assign n10936 = n10767 & ~n10935 ;
  assign n10937 = ~n10933 & n10936 ;
  assign n10938 = n4381 ^ n56 ^ 1'b0 ;
  assign n10939 = n5612 | n10938 ;
  assign n10940 = n10939 ^ n4007 ^ 1'b0 ;
  assign n10941 = n4214 & n10940 ;
  assign n10942 = n577 & ~n10941 ;
  assign n10943 = n73 & n8091 ;
  assign n10944 = n1087 & n10943 ;
  assign n10945 = n8451 & ~n10944 ;
  assign n10946 = n10942 | n10945 ;
  assign n10947 = ~n5756 & n6496 ;
  assign n10948 = n4019 & n10947 ;
  assign n10949 = n4024 | n10948 ;
  assign n10950 = n4760 & ~n10949 ;
  assign n10951 = n692 | n9056 ;
  assign n10952 = n3958 ^ n3320 ^ n2087 ;
  assign n10953 = n283 | n2488 ;
  assign n10954 = n10953 ^ n3314 ^ 1'b0 ;
  assign n10955 = ~n10952 & n10954 ;
  assign n10956 = n2282 | n10955 ;
  assign n10957 = ~n8830 & n10956 ;
  assign n10958 = n2756 ^ n2324 ^ n1040 ;
  assign n10959 = n7191 ^ n3097 ^ 1'b0 ;
  assign n10960 = n4008 & ~n10935 ;
  assign n10961 = n10960 ^ n7881 ^ 1'b0 ;
  assign n10962 = n6291 ^ n177 ^ 1'b0 ;
  assign n10963 = n2987 & ~n6235 ;
  assign n10964 = n4618 | n10963 ;
  assign n10965 = n2496 & n5353 ;
  assign n10966 = n10965 ^ n692 ^ 1'b0 ;
  assign n10967 = n6866 & ~n10966 ;
  assign n10968 = ~n6857 & n8553 ;
  assign n10972 = n6617 & n10154 ;
  assign n10973 = n10972 ^ n1024 ^ 1'b0 ;
  assign n10969 = n6449 ^ n1971 ^ 1'b0 ;
  assign n10970 = n2129 & ~n10969 ;
  assign n10971 = n842 | n10970 ;
  assign n10974 = n10973 ^ n10971 ^ n6316 ;
  assign n10975 = n10974 ^ n3015 ^ 1'b0 ;
  assign n10976 = n1657 | n3012 ;
  assign n10977 = n3143 & n6287 ;
  assign n10978 = n10977 ^ n4954 ^ 1'b0 ;
  assign n10979 = n9677 & ~n10978 ;
  assign n10980 = n9873 & n10979 ;
  assign n10981 = n911 | n1928 ;
  assign n10982 = n911 & ~n10981 ;
  assign n10983 = n5268 & ~n10982 ;
  assign n10984 = ~n663 & n765 ;
  assign n10985 = ~n765 & n10984 ;
  assign n10986 = ~n330 & n782 ;
  assign n10987 = n330 & n10986 ;
  assign n10988 = n10985 | n10987 ;
  assign n10989 = n10985 & ~n10988 ;
  assign n10990 = ~n7171 & n10989 ;
  assign n10991 = n220 & ~n717 ;
  assign n10992 = ~n220 & n10991 ;
  assign n10993 = n4254 & ~n10992 ;
  assign n10994 = ( n10983 & ~n10990 ) | ( n10983 & n10993 ) | ( ~n10990 & n10993 ) ;
  assign n10996 = ( ~n142 & n1434 ) | ( ~n142 & n9995 ) | ( n1434 & n9995 ) ;
  assign n10995 = n7722 & ~n8660 ;
  assign n10997 = n10996 ^ n10995 ^ 1'b0 ;
  assign n10998 = ~n1150 & n5831 ;
  assign n10999 = ~n4554 & n9580 ;
  assign n11000 = n10999 ^ n4493 ^ 1'b0 ;
  assign n11001 = n6120 | n9891 ;
  assign n11004 = n2587 & ~n5874 ;
  assign n11005 = n11004 ^ n1237 ^ 1'b0 ;
  assign n11002 = n1761 & n3181 ;
  assign n11003 = n5346 & n11002 ;
  assign n11006 = n11005 ^ n11003 ^ 1'b0 ;
  assign n11007 = n796 ^ n790 ^ 1'b0 ;
  assign n11008 = n3626 | n11007 ;
  assign n11009 = n7943 ^ n1701 ^ n1485 ;
  assign n11010 = ~n10076 & n11009 ;
  assign n11011 = n11010 ^ n3592 ^ 1'b0 ;
  assign n11012 = n5652 | n10370 ;
  assign n11013 = n11012 ^ n8161 ^ 1'b0 ;
  assign n11014 = n3251 & n11013 ;
  assign n11015 = n1254 & ~n2038 ;
  assign n11016 = n11015 ^ n3402 ^ 1'b0 ;
  assign n11017 = n623 | n790 ;
  assign n11018 = n3647 & ~n11017 ;
  assign n11019 = n2787 | n11018 ;
  assign n11020 = n11016 & ~n11019 ;
  assign n11021 = n9290 ^ n4845 ^ 1'b0 ;
  assign n11022 = n5054 & ~n6383 ;
  assign n11023 = n11022 ^ n3449 ^ 1'b0 ;
  assign n11024 = n2247 & ~n3968 ;
  assign n11025 = n1212 & ~n11024 ;
  assign n11026 = n5045 & n11025 ;
  assign n11027 = n11026 ^ n9741 ^ 1'b0 ;
  assign n11029 = n2108 & ~n4290 ;
  assign n11030 = n11029 ^ n3318 ^ 1'b0 ;
  assign n11031 = n11030 ^ n7467 ^ 1'b0 ;
  assign n11032 = n892 | n11031 ;
  assign n11028 = ~n7482 & n9464 ;
  assign n11033 = n11032 ^ n11028 ^ 1'b0 ;
  assign n11034 = n10898 ^ n2190 ^ 1'b0 ;
  assign n11035 = n1832 ^ n627 ^ 1'b0 ;
  assign n11036 = ~n5760 & n9721 ;
  assign n11037 = n11036 ^ n4252 ^ 1'b0 ;
  assign n11038 = ~n6102 & n6617 ;
  assign n11044 = n1921 & ~n3194 ;
  assign n11039 = n2363 ^ n2017 ^ n1578 ;
  assign n11040 = n11039 ^ n4065 ^ 1'b0 ;
  assign n11041 = ~n1123 & n11040 ;
  assign n11042 = n7283 & n11041 ;
  assign n11043 = n11042 ^ n1770 ^ 1'b0 ;
  assign n11045 = n11044 ^ n11043 ^ 1'b0 ;
  assign n11046 = ~n326 & n11045 ;
  assign n11047 = n9808 & ~n10320 ;
  assign n11048 = n11047 ^ n2618 ^ 1'b0 ;
  assign n11049 = n3990 & n6560 ;
  assign n11050 = ( n1398 & n10486 ) | ( n1398 & ~n11049 ) | ( n10486 & ~n11049 ) ;
  assign n11051 = n6605 ^ n1771 ^ 1'b0 ;
  assign n11052 = n8647 & n11051 ;
  assign n11053 = ~n10526 & n11052 ;
  assign n11054 = n11053 ^ n8354 ^ 1'b0 ;
  assign n11055 = n8719 ^ n8650 ^ 1'b0 ;
  assign n11056 = n11055 ^ n4571 ^ 1'b0 ;
  assign n11060 = n2749 & n3378 ;
  assign n11061 = n11060 ^ n1164 ^ 1'b0 ;
  assign n11057 = ~n3045 & n3210 ;
  assign n11058 = ~n1462 & n11057 ;
  assign n11059 = n11058 ^ n8766 ^ n7590 ;
  assign n11062 = n11061 ^ n11059 ^ n98 ;
  assign n11063 = n657 & ~n8142 ;
  assign n11064 = ~n4229 & n6326 ;
  assign n11065 = n5303 | n9604 ;
  assign n11066 = n5586 ^ n2292 ^ 1'b0 ;
  assign n11067 = n957 & n6568 ;
  assign n11068 = n11067 ^ n4487 ^ 1'b0 ;
  assign n11069 = n5095 & ~n7675 ;
  assign n11070 = n11068 & ~n11069 ;
  assign n11071 = n261 & n4163 ;
  assign n11072 = n6409 & n11071 ;
  assign n11073 = ~n3205 & n5508 ;
  assign n11074 = n380 & n4259 ;
  assign n11075 = n11073 & ~n11074 ;
  assign n11076 = n11075 ^ n2291 ^ 1'b0 ;
  assign n11078 = n4025 ^ n3461 ^ 1'b0 ;
  assign n11079 = n9235 & ~n11078 ;
  assign n11077 = n4438 ^ n4248 ^ 1'b0 ;
  assign n11080 = n11079 ^ n11077 ^ 1'b0 ;
  assign n11081 = n11076 & n11080 ;
  assign n11082 = n7539 ^ n5454 ^ 1'b0 ;
  assign n11083 = n5898 | n11082 ;
  assign n11084 = n6670 & ~n7531 ;
  assign n11085 = n2467 & n11084 ;
  assign n11086 = n2243 | n8266 ;
  assign n11087 = n8354 & ~n11086 ;
  assign n11094 = n9137 ^ n8727 ^ 1'b0 ;
  assign n11088 = n4914 & n7046 ;
  assign n11089 = n10253 ^ n7123 ^ 1'b0 ;
  assign n11090 = ~n1647 & n11089 ;
  assign n11091 = n1569 & n11090 ;
  assign n11092 = n11091 ^ n2755 ^ 1'b0 ;
  assign n11093 = n11088 & ~n11092 ;
  assign n11095 = n11094 ^ n11093 ^ 1'b0 ;
  assign n11096 = n3236 | n7829 ;
  assign n11097 = n11096 ^ n4852 ^ 1'b0 ;
  assign n11098 = n7534 & ~n11097 ;
  assign n11099 = ~n4893 & n10063 ;
  assign n11100 = ~n9189 & n11099 ;
  assign n11101 = n9256 ^ n6969 ^ 1'b0 ;
  assign n11102 = n6734 | n11101 ;
  assign n11103 = n320 & ~n4054 ;
  assign n11104 = n4556 & ~n11103 ;
  assign n11105 = n7066 & n11104 ;
  assign n11106 = n4427 ^ n4344 ^ n4133 ;
  assign n11107 = n11106 ^ n4007 ^ 1'b0 ;
  assign n11108 = n11107 ^ n3131 ^ 1'b0 ;
  assign n11109 = n3272 | n11108 ;
  assign n11110 = n3536 ^ n2367 ^ 1'b0 ;
  assign n11111 = n2005 & ~n11110 ;
  assign n11112 = n6578 | n11111 ;
  assign n11113 = n11109 & n11112 ;
  assign n11114 = n2820 | n4641 ;
  assign n11115 = n334 | n11114 ;
  assign n11116 = n1196 | n4907 ;
  assign n11117 = n7703 & ~n11116 ;
  assign n11118 = n7153 ^ n5847 ^ 1'b0 ;
  assign n11119 = ( ~n1055 & n8443 ) | ( ~n1055 & n9958 ) | ( n8443 & n9958 ) ;
  assign n11121 = ( n309 & n3962 ) | ( n309 & ~n4374 ) | ( n3962 & ~n4374 ) ;
  assign n11120 = n5018 ^ n3646 ^ 1'b0 ;
  assign n11122 = n11121 ^ n11120 ^ n2522 ;
  assign n11123 = n6933 ^ n1389 ^ 1'b0 ;
  assign n11124 = n11123 ^ n286 ^ 1'b0 ;
  assign n11125 = n6506 & n11124 ;
  assign n11126 = ~n4801 & n11125 ;
  assign n11127 = n7358 & n11126 ;
  assign n11128 = n4012 & n8697 ;
  assign n11129 = n3416 & n11128 ;
  assign n11130 = n5526 ^ n163 ^ 1'b0 ;
  assign n11131 = n1356 | n11130 ;
  assign n11132 = n5834 | n7960 ;
  assign n11133 = n11132 ^ n690 ^ 1'b0 ;
  assign n11134 = n239 & ~n6872 ;
  assign n11135 = n11133 & n11134 ;
  assign n11136 = n5215 ^ n368 ^ 1'b0 ;
  assign n11137 = n11135 | n11136 ;
  assign n11138 = n1567 | n4164 ;
  assign n11139 = n2104 & n8338 ;
  assign n11140 = n3052 & n11139 ;
  assign n11141 = n6397 ^ n826 ^ 1'b0 ;
  assign n11142 = n11141 ^ n5543 ^ 1'b0 ;
  assign n11143 = n3469 & ~n8725 ;
  assign n11144 = n11143 ^ n445 ^ 1'b0 ;
  assign n11145 = ~n646 & n2377 ;
  assign n11146 = n11145 ^ n6699 ^ 1'b0 ;
  assign n11147 = ( n2527 & ~n8737 ) | ( n2527 & n11146 ) | ( ~n8737 & n11146 ) ;
  assign n11148 = n6609 & ~n8908 ;
  assign n11149 = n1363 & n1654 ;
  assign n11150 = n395 & n11149 ;
  assign n11151 = n11150 ^ n10575 ^ 1'b0 ;
  assign n11152 = ~n8018 & n11151 ;
  assign n11153 = ~n273 & n8503 ;
  assign n11154 = n11153 ^ n10038 ^ 1'b0 ;
  assign n11155 = n7537 ^ n4681 ^ 1'b0 ;
  assign n11160 = ~n2062 & n2660 ;
  assign n11156 = ~n4604 & n9371 ;
  assign n11157 = n11156 ^ n5394 ^ 1'b0 ;
  assign n11158 = n11157 ^ n1226 ^ 1'b0 ;
  assign n11159 = n5859 & n11158 ;
  assign n11161 = n11160 ^ n11159 ^ 1'b0 ;
  assign n11162 = ~n3738 & n11161 ;
  assign n11164 = n1461 ^ n1460 ^ 1'b0 ;
  assign n11163 = n5443 & n10752 ;
  assign n11165 = n11164 ^ n11163 ^ 1'b0 ;
  assign n11166 = n1534 ^ n978 ^ 1'b0 ;
  assign n11167 = n2758 & ~n2837 ;
  assign n11168 = n11167 ^ n4789 ^ n4537 ;
  assign n11169 = n2560 | n11168 ;
  assign n11170 = ~n2470 & n7054 ;
  assign n11171 = ~n2019 & n11170 ;
  assign n11172 = n9109 & n11171 ;
  assign n11173 = n11172 ^ n5914 ^ 1'b0 ;
  assign n11174 = ~n11169 & n11173 ;
  assign n11175 = n559 & ~n10087 ;
  assign n11176 = n11175 ^ n387 ^ 1'b0 ;
  assign n11177 = n1426 & n3751 ;
  assign n11178 = n3631 & n6179 ;
  assign n11179 = n11178 ^ n6957 ^ 1'b0 ;
  assign n11180 = n11179 ^ n8482 ^ 1'b0 ;
  assign n11181 = ~n222 & n4504 ;
  assign n11182 = n11181 ^ n9804 ^ 1'b0 ;
  assign n11183 = n4143 & ~n11182 ;
  assign n11184 = n4273 | n5273 ;
  assign n11185 = n4754 ^ n132 ^ 1'b0 ;
  assign n11186 = n7799 & ~n11185 ;
  assign n11187 = n11186 ^ n9199 ^ 1'b0 ;
  assign n11188 = n1730 & ~n3712 ;
  assign n11189 = n11188 ^ n9272 ^ 1'b0 ;
  assign n11190 = n11189 ^ n3927 ^ 1'b0 ;
  assign n11191 = n8463 & n11190 ;
  assign n11192 = n11191 ^ n770 ^ 1'b0 ;
  assign n11193 = n1277 ^ n108 ^ 1'b0 ;
  assign n11194 = n2458 & n11193 ;
  assign n11195 = ~n753 & n3306 ;
  assign n11196 = ~n503 & n11195 ;
  assign n11197 = n4478 | n11196 ;
  assign n11198 = n11197 ^ n8289 ^ 1'b0 ;
  assign n11199 = n2381 & ~n8456 ;
  assign n11200 = n1663 & ~n11199 ;
  assign n11201 = n11198 & n11200 ;
  assign n11202 = ( n2900 & n3746 ) | ( n2900 & n9605 ) | ( n3746 & n9605 ) ;
  assign n11203 = n8448 | n8599 ;
  assign n11204 = n6135 & ~n11203 ;
  assign n11205 = ( ~n4487 & n5217 ) | ( ~n4487 & n6831 ) | ( n5217 & n6831 ) ;
  assign n11206 = n5767 & ~n11205 ;
  assign n11207 = n404 & ~n8814 ;
  assign n11208 = n1939 & n11207 ;
  assign n11209 = n11208 ^ n5447 ^ 1'b0 ;
  assign n11210 = n3757 | n11209 ;
  assign n11211 = n11206 & ~n11210 ;
  assign n11214 = n1912 & n2108 ;
  assign n11212 = n3903 | n8336 ;
  assign n11213 = ~n1205 & n11212 ;
  assign n11215 = n11214 ^ n11213 ^ 1'b0 ;
  assign n11216 = n3616 & ~n11215 ;
  assign n11217 = ~n749 & n11216 ;
  assign n11219 = n5247 ^ n4767 ^ 1'b0 ;
  assign n11220 = ~n1650 & n11219 ;
  assign n11218 = n5682 & n7038 ;
  assign n11221 = n11220 ^ n11218 ^ n8512 ;
  assign n11222 = ( n6545 & ~n10703 ) | ( n6545 & n11221 ) | ( ~n10703 & n11221 ) ;
  assign n11223 = ( ~n326 & n3045 ) | ( ~n326 & n7763 ) | ( n3045 & n7763 ) ;
  assign n11224 = ~n311 & n2121 ;
  assign n11225 = n11224 ^ n2723 ^ 1'b0 ;
  assign n11226 = n2114 & ~n11225 ;
  assign n11227 = n11226 ^ n1984 ^ 1'b0 ;
  assign n11228 = ( n1785 & ~n10812 ) | ( n1785 & n11227 ) | ( ~n10812 & n11227 ) ;
  assign n11229 = n43 & n2192 ;
  assign n11230 = ~n1896 & n11229 ;
  assign n11231 = n2953 & n8086 ;
  assign n11232 = n11231 ^ n1121 ^ 1'b0 ;
  assign n11233 = n7909 ^ n7371 ^ 1'b0 ;
  assign n11234 = n6051 | n10841 ;
  assign n11235 = n11234 ^ n6405 ^ n2735 ;
  assign n11236 = n11235 ^ n7649 ^ 1'b0 ;
  assign n11237 = n11233 | n11236 ;
  assign n11238 = ~n2225 & n11237 ;
  assign n11239 = n4895 ^ n418 ^ 1'b0 ;
  assign n11240 = ~n10348 & n11239 ;
  assign n11241 = n3955 & n11240 ;
  assign n11242 = n2694 & n11241 ;
  assign n11243 = n466 & ~n11242 ;
  assign n11244 = n7691 ^ n76 ^ 1'b0 ;
  assign n11245 = n9962 ^ n2031 ^ 1'b0 ;
  assign n11246 = n7239 & ~n11245 ;
  assign n11247 = n1747 & ~n7767 ;
  assign n11248 = n11247 ^ n5982 ^ 1'b0 ;
  assign n11249 = n11248 ^ n5766 ^ 1'b0 ;
  assign n11250 = n1002 & ~n3009 ;
  assign n11251 = n11250 ^ n1068 ^ 1'b0 ;
  assign n11252 = n11251 ^ n10013 ^ 1'b0 ;
  assign n11253 = n11252 ^ n4599 ^ 1'b0 ;
  assign n11254 = n5702 ^ n2576 ^ 1'b0 ;
  assign n11255 = n9383 | n11254 ;
  assign n11256 = n1804 & n5613 ;
  assign n11257 = n10027 ^ n1845 ^ 1'b0 ;
  assign n11258 = n5388 | n8224 ;
  assign n11259 = ~n6356 & n7492 ;
  assign n11260 = n291 & n11259 ;
  assign n11261 = n4252 ^ n4010 ^ 1'b0 ;
  assign n11262 = n4885 ^ n2163 ^ 1'b0 ;
  assign n11263 = n309 | n11262 ;
  assign n11264 = n5618 & ~n11263 ;
  assign n11265 = n9421 | n11264 ;
  assign n11266 = n11261 & ~n11265 ;
  assign n11267 = n657 & n7155 ;
  assign n11268 = n11267 ^ n2120 ^ 1'b0 ;
  assign n11269 = n8403 ^ n5444 ^ 1'b0 ;
  assign n11270 = n11268 | n11269 ;
  assign n11271 = n8197 ^ n4379 ^ n1081 ;
  assign n11272 = n104 & ~n11271 ;
  assign n11273 = ~n5401 & n11272 ;
  assign n11274 = n4551 | n5260 ;
  assign n11275 = n2717 ^ n2275 ^ 1'b0 ;
  assign n11276 = n2680 | n11275 ;
  assign n11277 = n3145 ^ n620 ^ 1'b0 ;
  assign n11278 = ( ~n205 & n290 ) | ( ~n205 & n2291 ) | ( n290 & n2291 ) ;
  assign n11279 = ~n11277 & n11278 ;
  assign n11280 = ~n11276 & n11279 ;
  assign n11281 = ~n209 & n11280 ;
  assign n11282 = n5001 ^ n4583 ^ 1'b0 ;
  assign n11283 = n7741 & n11282 ;
  assign n11284 = n10719 & n11283 ;
  assign n11285 = n9254 & n11284 ;
  assign n11286 = n623 | n9717 ;
  assign n11287 = n9550 & ~n11286 ;
  assign n11288 = n2940 & ~n3359 ;
  assign n11289 = n11288 ^ n6231 ^ 1'b0 ;
  assign n11290 = n11289 ^ n8566 ^ 1'b0 ;
  assign n11291 = n6428 ^ n849 ^ n792 ;
  assign n11292 = n2472 & n11291 ;
  assign n11293 = n11292 ^ n8150 ^ 1'b0 ;
  assign n11294 = ~n9049 & n11293 ;
  assign n11295 = ~n311 & n339 ;
  assign n11296 = n3696 & n5309 ;
  assign n11297 = n11296 ^ n7791 ^ 1'b0 ;
  assign n11298 = n10237 ^ n1307 ^ 1'b0 ;
  assign n11299 = n4525 & n11298 ;
  assign n11300 = n2733 ^ n352 ^ 1'b0 ;
  assign n11301 = n518 ^ n362 ^ 1'b0 ;
  assign n11302 = n11300 | n11301 ;
  assign n11303 = n970 | n1491 ;
  assign n11304 = n11303 ^ n7327 ^ 1'b0 ;
  assign n11305 = n11304 ^ n6430 ^ n305 ;
  assign n11306 = ( n8211 & n11302 ) | ( n8211 & n11305 ) | ( n11302 & n11305 ) ;
  assign n11307 = ~n2460 & n9731 ;
  assign n11308 = n4357 & n11307 ;
  assign n11311 = n6350 ^ n1765 ^ 1'b0 ;
  assign n11312 = n3110 | n11311 ;
  assign n11309 = n5719 ^ n3902 ^ 1'b0 ;
  assign n11310 = n3470 & ~n11309 ;
  assign n11313 = n11312 ^ n11310 ^ 1'b0 ;
  assign n11314 = n5581 ^ n2373 ^ 1'b0 ;
  assign n11315 = n3853 & ~n10055 ;
  assign n11316 = ( n4270 & n10706 ) | ( n4270 & n11315 ) | ( n10706 & n11315 ) ;
  assign n11317 = n11316 ^ n4291 ^ 1'b0 ;
  assign n11318 = ~n5724 & n11317 ;
  assign n11319 = n9054 ^ n2956 ^ 1'b0 ;
  assign n11320 = n5880 | n11319 ;
  assign n11321 = ~n3150 & n11320 ;
  assign n11322 = n738 | n1087 ;
  assign n11323 = n302 & ~n4843 ;
  assign n11324 = ( n2489 & ~n3438 ) | ( n2489 & n4105 ) | ( ~n3438 & n4105 ) ;
  assign n11325 = n11324 ^ n1688 ^ 1'b0 ;
  assign n11326 = n1182 ^ n61 ^ 1'b0 ;
  assign n11327 = n3119 & ~n11326 ;
  assign n11328 = n3126 & n11327 ;
  assign n11329 = ~n2321 & n11328 ;
  assign n11330 = n9940 ^ n4578 ^ 1'b0 ;
  assign n11331 = ~n2803 & n11330 ;
  assign n11332 = n4153 | n5342 ;
  assign n11333 = n676 | n11332 ;
  assign n11334 = n11333 ^ n3583 ^ 1'b0 ;
  assign n11335 = n1770 & ~n2522 ;
  assign n11336 = n11335 ^ n4405 ^ 1'b0 ;
  assign n11337 = ~n2891 & n11336 ;
  assign n11338 = n395 & n11337 ;
  assign n11339 = n11338 ^ n4727 ^ n3418 ;
  assign n11340 = ~n125 & n459 ;
  assign n11341 = n11340 ^ n5168 ^ 1'b0 ;
  assign n11344 = n1271 ^ n749 ^ 1'b0 ;
  assign n11345 = ~n139 & n11344 ;
  assign n11342 = n8723 ^ n802 ^ 1'b0 ;
  assign n11343 = n4569 | n11342 ;
  assign n11346 = n11345 ^ n11343 ^ 1'b0 ;
  assign n11347 = ~n9958 & n10822 ;
  assign n11348 = n11347 ^ n1213 ^ 1'b0 ;
  assign n11349 = ~n1077 & n11348 ;
  assign n11351 = n288 | n2415 ;
  assign n11352 = n11351 ^ n3774 ^ 1'b0 ;
  assign n11350 = ~n140 & n3274 ;
  assign n11353 = n11352 ^ n11350 ^ 1'b0 ;
  assign n11355 = n1128 & n5074 ;
  assign n11354 = n3785 & n10472 ;
  assign n11356 = n11355 ^ n11354 ^ 1'b0 ;
  assign n11357 = n11356 ^ n6924 ^ 1'b0 ;
  assign n11358 = n1246 & ~n11357 ;
  assign n11359 = n7659 ^ n3290 ^ 1'b0 ;
  assign n11360 = n11359 ^ n6730 ^ 1'b0 ;
  assign n11361 = n9713 ^ n1897 ^ 1'b0 ;
  assign n11362 = ~n11360 & n11361 ;
  assign n11363 = n6424 | n10497 ;
  assign n11364 = n3226 & n4785 ;
  assign n11365 = n914 & n7685 ;
  assign n11366 = n4860 & n11365 ;
  assign n11367 = n497 & n2932 ;
  assign n11368 = n11055 & ~n11367 ;
  assign n11369 = n11368 ^ n5886 ^ 1'b0 ;
  assign n11370 = n533 ^ n266 ^ 1'b0 ;
  assign n11371 = ~n709 & n11370 ;
  assign n11372 = n11371 ^ n10556 ^ 1'b0 ;
  assign n11374 = ( ~n1089 & n3209 ) | ( ~n1089 & n10215 ) | ( n3209 & n10215 ) ;
  assign n11373 = n8820 & n9868 ;
  assign n11375 = n11374 ^ n11373 ^ 1'b0 ;
  assign n11376 = n3917 | n4119 ;
  assign n11377 = n11376 ^ n2361 ^ 1'b0 ;
  assign n11378 = n1611 ^ n1211 ^ 1'b0 ;
  assign n11379 = n2004 & n11378 ;
  assign n11380 = n11379 ^ n3166 ^ 1'b0 ;
  assign n11381 = n8235 & ~n11380 ;
  assign n11382 = n2145 & ~n11381 ;
  assign n11383 = ~n6215 & n11382 ;
  assign n11384 = n8756 | n11383 ;
  assign n11385 = n858 | n7655 ;
  assign n11386 = n11385 ^ n362 ^ 1'b0 ;
  assign n11387 = n11386 ^ n3382 ^ n2395 ;
  assign n11388 = n1161 | n6583 ;
  assign n11389 = ~n2610 & n7749 ;
  assign n11390 = n3886 & n6274 ;
  assign n11391 = n5037 ^ n43 ^ 1'b0 ;
  assign n11392 = ~n4346 & n11391 ;
  assign n11393 = n1207 | n11392 ;
  assign n11394 = n11393 ^ n5240 ^ 1'b0 ;
  assign n11395 = n1802 & n6230 ;
  assign n11396 = n11395 ^ n7718 ^ 1'b0 ;
  assign n11397 = ( n7307 & n8151 ) | ( n7307 & n10372 ) | ( n8151 & n10372 ) ;
  assign n11398 = n744 & n8195 ;
  assign n11399 = ~n744 & n11398 ;
  assign n11400 = n2954 ^ n2539 ^ 1'b0 ;
  assign n11401 = n4154 ^ n3353 ^ 1'b0 ;
  assign n11402 = n11400 & ~n11401 ;
  assign n11403 = n3110 ^ n1157 ^ 1'b0 ;
  assign n11404 = n2556 | n11403 ;
  assign n11405 = n11404 ^ n11164 ^ 1'b0 ;
  assign n11406 = n1422 & ~n7609 ;
  assign n11407 = n10121 | n11406 ;
  assign n11409 = n5246 ^ n1126 ^ 1'b0 ;
  assign n11410 = n2854 & ~n11409 ;
  assign n11411 = n11410 ^ n2855 ^ 1'b0 ;
  assign n11408 = n8883 & ~n11126 ;
  assign n11412 = n11411 ^ n11408 ^ 1'b0 ;
  assign n11413 = n5352 ^ n4814 ^ 1'b0 ;
  assign n11414 = ~n1461 & n11413 ;
  assign n11415 = n11414 ^ n5036 ^ 1'b0 ;
  assign n11416 = n4346 & n11415 ;
  assign n11417 = n6132 ^ n1064 ^ 1'b0 ;
  assign n11418 = n9104 & ~n10848 ;
  assign n11419 = n3664 ^ n2678 ^ 1'b0 ;
  assign n11420 = ~n1109 & n11419 ;
  assign n11421 = n661 & ~n11420 ;
  assign n11422 = n152 | n1280 ;
  assign n11423 = n3744 | n11422 ;
  assign n11424 = n11423 ^ n2272 ^ 1'b0 ;
  assign n11425 = ~n2359 & n11424 ;
  assign n11426 = n9441 | n11425 ;
  assign n11427 = n246 & ~n3351 ;
  assign n11428 = ( n1439 & n6039 ) | ( n1439 & ~n11427 ) | ( n6039 & ~n11427 ) ;
  assign n11429 = n5295 | n9434 ;
  assign n11430 = n667 & ~n9447 ;
  assign n11431 = ~n5145 & n11430 ;
  assign n11432 = n6526 ^ n733 ^ 1'b0 ;
  assign n11433 = ~n3762 & n11432 ;
  assign n11434 = n11433 ^ n7460 ^ 1'b0 ;
  assign n11435 = n5085 ^ n1416 ^ 1'b0 ;
  assign n11436 = n11264 ^ n4857 ^ 1'b0 ;
  assign n11437 = ~n806 & n968 ;
  assign n11438 = n5419 & ~n11437 ;
  assign n11439 = n9062 ^ n7949 ^ 1'b0 ;
  assign n11440 = ~n2046 & n7372 ;
  assign n11442 = ~n4593 & n8347 ;
  assign n11443 = n11442 ^ n5548 ^ n2145 ;
  assign n11441 = ~n630 & n9985 ;
  assign n11444 = n11443 ^ n11441 ^ 1'b0 ;
  assign n11445 = n11444 ^ n343 ^ 1'b0 ;
  assign n11446 = ( n2273 & ~n5394 ) | ( n2273 & n5402 ) | ( ~n5394 & n5402 ) ;
  assign n11447 = n1688 ^ n1369 ^ 1'b0 ;
  assign n11448 = n6856 & n7476 ;
  assign n11449 = n9330 & n11448 ;
  assign n11450 = n11449 ^ n10711 ^ 1'b0 ;
  assign n11451 = ~n1116 & n11450 ;
  assign n11452 = n2148 & ~n9088 ;
  assign n11453 = n1747 & ~n2522 ;
  assign n11454 = n1997 | n7583 ;
  assign n11455 = n8715 ^ n1210 ^ 1'b0 ;
  assign n11456 = n3657 ^ n2373 ^ n227 ;
  assign n11457 = n11456 ^ n8550 ^ n6498 ;
  assign n11458 = n4872 & ~n11457 ;
  assign n11459 = n9770 & n11458 ;
  assign n11460 = ~n11455 & n11459 ;
  assign n11461 = n1847 & ~n5971 ;
  assign n11462 = ~n3518 & n6566 ;
  assign n11463 = n3854 & n6421 ;
  assign n11464 = n11463 ^ n4294 ^ 1'b0 ;
  assign n11465 = n4881 ^ n3477 ^ 1'b0 ;
  assign n11466 = n11464 & n11465 ;
  assign n11467 = n854 | n861 ;
  assign n11468 = n1174 & ~n2143 ;
  assign n11469 = n4933 ^ n463 ^ n150 ;
  assign n11470 = n4716 & ~n11469 ;
  assign n11471 = n4222 & n11470 ;
  assign n11472 = n10146 & n11471 ;
  assign n11473 = n7899 & ~n11472 ;
  assign n11474 = n11473 ^ n4326 ^ 1'b0 ;
  assign n11475 = n77 & ~n2755 ;
  assign n11476 = n8684 & n11475 ;
  assign n11477 = n4910 & ~n8706 ;
  assign n11478 = n4464 | n10663 ;
  assign n11479 = n5431 | n11478 ;
  assign n11480 = n7010 & ~n11479 ;
  assign n11481 = n5663 ^ n3474 ^ n336 ;
  assign n11482 = ( ~n1237 & n2282 ) | ( ~n1237 & n11481 ) | ( n2282 & n11481 ) ;
  assign n11483 = n1520 ^ n723 ^ 1'b0 ;
  assign n11484 = ~n2658 & n6534 ;
  assign n11485 = n5783 ^ n5632 ^ 1'b0 ;
  assign n11486 = n1464 & ~n3466 ;
  assign n11487 = ~n685 & n7835 ;
  assign n11488 = n9289 ^ n8593 ^ 1'b0 ;
  assign n11489 = n7668 & ~n11488 ;
  assign n11490 = n3432 ^ n30 ^ 1'b0 ;
  assign n11491 = n2411 & ~n11490 ;
  assign n11492 = n288 | n3762 ;
  assign n11493 = n3762 & ~n11492 ;
  assign n11494 = n11491 & n11493 ;
  assign n11495 = ~n2726 & n11494 ;
  assign n11496 = ~n11494 & n11495 ;
  assign n11497 = n6392 ^ n6012 ^ n1469 ;
  assign n11498 = n3796 & ~n11497 ;
  assign n11499 = ~n1442 & n11498 ;
  assign n11500 = n5646 ^ n5018 ^ 1'b0 ;
  assign n11501 = n11500 ^ n6878 ^ 1'b0 ;
  assign n11502 = ~n5018 & n11501 ;
  assign n11503 = n6559 & n7524 ;
  assign n11504 = n4977 ^ n2417 ^ 1'b0 ;
  assign n11505 = n1202 | n4778 ;
  assign n11506 = n11505 ^ n6323 ^ 1'b0 ;
  assign n11507 = n1697 | n6586 ;
  assign n11508 = n4914 | n11507 ;
  assign n11509 = ~n3443 & n5082 ;
  assign n11510 = ~n356 & n11509 ;
  assign n11511 = n11510 ^ n1938 ^ 1'b0 ;
  assign n11512 = n5137 ^ n2821 ^ 1'b0 ;
  assign n11513 = ~n2498 & n11512 ;
  assign n11514 = n3779 & n11513 ;
  assign n11515 = n2580 ^ n522 ^ 1'b0 ;
  assign n11516 = n11515 ^ n1802 ^ 1'b0 ;
  assign n11517 = ~n4519 & n11516 ;
  assign n11518 = ( n704 & n2563 ) | ( n704 & ~n11517 ) | ( n2563 & ~n11517 ) ;
  assign n11521 = ~n1603 & n3787 ;
  assign n11522 = n9153 | n11521 ;
  assign n11523 = n11522 ^ n2137 ^ 1'b0 ;
  assign n11519 = n2632 ^ n1951 ^ 1'b0 ;
  assign n11520 = n1215 & ~n11519 ;
  assign n11524 = n11523 ^ n11520 ^ 1'b0 ;
  assign n11525 = n8857 & ~n11524 ;
  assign n11526 = n3191 & n4048 ;
  assign n11527 = n11526 ^ n4376 ^ 1'b0 ;
  assign n11528 = ~n7945 & n11527 ;
  assign n11529 = ~n11525 & n11528 ;
  assign n11530 = n5549 & ~n11529 ;
  assign n11531 = n10465 ^ n9470 ^ 1'b0 ;
  assign n11532 = n466 & ~n11531 ;
  assign n11533 = n3873 ^ n3118 ^ 1'b0 ;
  assign n11534 = n1995 & n4229 ;
  assign n11535 = n3822 | n4116 ;
  assign n11536 = n397 | n11535 ;
  assign n11537 = ~n3114 & n4576 ;
  assign n11538 = n3634 & n11537 ;
  assign n11539 = n9028 ^ n1709 ^ 1'b0 ;
  assign n11540 = ~n11538 & n11539 ;
  assign n11541 = ( n152 & n235 ) | ( n152 & n1739 ) | ( n235 & n1739 ) ;
  assign n11542 = n1104 & n2902 ;
  assign n11543 = ~n5989 & n11542 ;
  assign n11545 = ~n2178 & n2248 ;
  assign n11546 = n4726 & n11545 ;
  assign n11544 = n1002 & ~n4554 ;
  assign n11547 = n11546 ^ n11544 ^ 1'b0 ;
  assign n11548 = ~n4270 & n11547 ;
  assign n11549 = n4005 & n11548 ;
  assign n11550 = n6687 & n7508 ;
  assign n11551 = n1917 ^ n840 ^ 1'b0 ;
  assign n11552 = n5872 ^ n1652 ^ 1'b0 ;
  assign n11553 = ( n5417 & n7186 ) | ( n5417 & ~n11552 ) | ( n7186 & ~n11552 ) ;
  assign n11554 = n1745 | n3494 ;
  assign n11555 = ( n3400 & n11553 ) | ( n3400 & n11554 ) | ( n11553 & n11554 ) ;
  assign n11556 = n6989 ^ n2361 ^ 1'b0 ;
  assign n11557 = n9426 | n11556 ;
  assign n11558 = n7027 ^ n5829 ^ 1'b0 ;
  assign n11559 = n8889 | n11558 ;
  assign n11560 = n3218 & ~n3957 ;
  assign n11561 = ( n2857 & ~n6975 ) | ( n2857 & n9797 ) | ( ~n6975 & n9797 ) ;
  assign n11562 = n11561 ^ n8249 ^ n7877 ;
  assign n11563 = n10264 | n11562 ;
  assign n11564 = n559 & ~n989 ;
  assign n11565 = n2403 & n11249 ;
  assign n11566 = ~n9687 & n11565 ;
  assign n11567 = n11566 ^ n10601 ^ 1'b0 ;
  assign n11568 = n5141 & ~n5944 ;
  assign n11569 = n11568 ^ n3794 ^ 1'b0 ;
  assign n11570 = n3086 & ~n11569 ;
  assign n11571 = n11333 ^ n1688 ^ 1'b0 ;
  assign n11572 = ~n4211 & n11571 ;
  assign n11573 = n11572 ^ n5072 ^ 1'b0 ;
  assign n11575 = n582 | n4464 ;
  assign n11576 = n11575 ^ n746 ^ 1'b0 ;
  assign n11577 = n11576 ^ n277 ^ 1'b0 ;
  assign n11574 = n6458 ^ n431 ^ 1'b0 ;
  assign n11578 = n11577 ^ n11574 ^ n7154 ;
  assign n11579 = n11578 ^ n11184 ^ 1'b0 ;
  assign n11580 = ~n11573 & n11579 ;
  assign n11581 = n591 | n6841 ;
  assign n11582 = n5866 & ~n11581 ;
  assign n11583 = ~n1369 & n7476 ;
  assign n11584 = n10325 ^ n9741 ^ 1'b0 ;
  assign n11588 = n5217 ^ n4691 ^ 1'b0 ;
  assign n11585 = n4379 | n6931 ;
  assign n11586 = n6621 ^ n212 ^ 1'b0 ;
  assign n11587 = n11585 & ~n11586 ;
  assign n11589 = n11588 ^ n11587 ^ 1'b0 ;
  assign n11590 = ~n6946 & n11406 ;
  assign n11591 = n11590 ^ n2351 ^ 1'b0 ;
  assign n11592 = n2682 ^ n199 ^ 1'b0 ;
  assign n11593 = ~n8635 & n11592 ;
  assign n11594 = n376 & n3105 ;
  assign n11595 = n11594 ^ n6523 ^ 1'b0 ;
  assign n11596 = n1552 & n10079 ;
  assign n11597 = ~n565 & n11596 ;
  assign n11598 = n5182 | n11597 ;
  assign n11599 = n5367 | n11598 ;
  assign n11600 = n11599 ^ n4677 ^ 1'b0 ;
  assign n11601 = n5395 & ~n6027 ;
  assign n11602 = ~n3232 & n11601 ;
  assign n11603 = n5469 ^ n2366 ^ 1'b0 ;
  assign n11604 = n344 | n11603 ;
  assign n11605 = ( ~n4645 & n8776 ) | ( ~n4645 & n11604 ) | ( n8776 & n11604 ) ;
  assign n11606 = n4460 | n11605 ;
  assign n11607 = n11606 ^ n6216 ^ 1'b0 ;
  assign n11608 = n2891 | n3747 ;
  assign n11609 = n2154 | n2806 ;
  assign n11610 = n11609 ^ n7092 ^ 1'b0 ;
  assign n11611 = ~n2394 & n6669 ;
  assign n11612 = ~n7265 & n11611 ;
  assign n11613 = n5991 ^ n4256 ^ 1'b0 ;
  assign n11614 = n3072 ^ n2420 ^ n1770 ;
  assign n11615 = n3272 | n11614 ;
  assign n11616 = n11615 ^ n4436 ^ 1'b0 ;
  assign n11617 = n11616 ^ n7483 ^ 1'b0 ;
  assign n11618 = n6823 | n11617 ;
  assign n11619 = n7338 | n11618 ;
  assign n11620 = ~n3085 & n11619 ;
  assign n11621 = n11435 ^ n8475 ^ 1'b0 ;
  assign n11622 = n2362 ^ n1545 ^ 1'b0 ;
  assign n11623 = n11622 ^ n7589 ^ 1'b0 ;
  assign n11624 = n2399 & n11623 ;
  assign n11625 = n9063 ^ n3473 ^ 1'b0 ;
  assign n11627 = n6966 ^ n2130 ^ 1'b0 ;
  assign n11628 = n9892 ^ n914 ^ 1'b0 ;
  assign n11629 = n10374 & ~n11628 ;
  assign n11630 = n11627 & n11629 ;
  assign n11631 = n1476 & ~n11630 ;
  assign n11632 = n11631 ^ n1643 ^ 1'b0 ;
  assign n11626 = n1096 | n3372 ;
  assign n11633 = n11632 ^ n11626 ^ 1'b0 ;
  assign n11635 = ~n1254 & n3680 ;
  assign n11634 = n6598 & ~n11248 ;
  assign n11636 = n11635 ^ n11634 ^ 1'b0 ;
  assign n11637 = ~n1511 & n1561 ;
  assign n11638 = n2632 | n11637 ;
  assign n11639 = n2469 | n8963 ;
  assign n11640 = n11638 | n11639 ;
  assign n11641 = n8381 & ~n9915 ;
  assign n11642 = ~n6248 & n11641 ;
  assign n11643 = n4955 ^ x11 ^ 1'b0 ;
  assign n11644 = ~n4819 & n11643 ;
  assign n11646 = n7703 ^ n304 ^ 1'b0 ;
  assign n11647 = n2469 | n11646 ;
  assign n11648 = ( n1650 & ~n6401 ) | ( n1650 & n11647 ) | ( ~n6401 & n11647 ) ;
  assign n11645 = n2560 | n5706 ;
  assign n11649 = n11648 ^ n11645 ^ 1'b0 ;
  assign n11650 = n5077 & ~n11649 ;
  assign n11651 = ~n10692 & n11650 ;
  assign n11652 = n1210 & ~n3361 ;
  assign n11653 = n316 | n11652 ;
  assign n11654 = n1211 & ~n10362 ;
  assign n11655 = n11654 ^ n448 ^ 1'b0 ;
  assign n11656 = n7048 & n11655 ;
  assign n11657 = n6156 & ~n6229 ;
  assign n11658 = n2537 & n10863 ;
  assign n11659 = n11658 ^ n2541 ^ 1'b0 ;
  assign n11660 = n1323 ^ n270 ^ 1'b0 ;
  assign n11661 = n5264 | n11660 ;
  assign n11662 = n914 & n11661 ;
  assign n11663 = n5781 | n6625 ;
  assign n11664 = n7087 | n11663 ;
  assign n11665 = n1659 & n2102 ;
  assign n11666 = n3032 & n11665 ;
  assign n11667 = ( n2317 & n11664 ) | ( n2317 & n11666 ) | ( n11664 & n11666 ) ;
  assign n11668 = n4396 ^ n3236 ^ n1915 ;
  assign n11669 = n9955 & n11668 ;
  assign n11670 = n11669 ^ n1161 ^ 1'b0 ;
  assign n11671 = n870 & ~n11670 ;
  assign n11672 = ~n261 & n1254 ;
  assign n11673 = n11672 ^ n2778 ^ 1'b0 ;
  assign n11674 = n796 & n3903 ;
  assign n11675 = ~n1431 & n11674 ;
  assign n11676 = n11673 & n11675 ;
  assign n11677 = n2308 ^ n124 ^ 1'b0 ;
  assign n11678 = ~n2694 & n11677 ;
  assign n11679 = n7350 & n11678 ;
  assign n11680 = n11679 ^ n6212 ^ 1'b0 ;
  assign n11681 = ( n1394 & n6651 ) | ( n1394 & n6792 ) | ( n6651 & n6792 ) ;
  assign n11682 = ( n703 & ~n2632 ) | ( n703 & n2953 ) | ( ~n2632 & n2953 ) ;
  assign n11683 = n11682 ^ n667 ^ 1'b0 ;
  assign n11684 = n1927 & n11683 ;
  assign n11685 = n11684 ^ n4750 ^ 1'b0 ;
  assign n11686 = n11685 ^ n144 ^ 1'b0 ;
  assign n11687 = n11681 & n11686 ;
  assign n11688 = ~n11680 & n11687 ;
  assign n11689 = n10099 ^ n9194 ^ n753 ;
  assign n11690 = n11689 ^ n11483 ^ 1'b0 ;
  assign n11691 = n6748 | n7396 ;
  assign n11692 = n11671 & ~n11691 ;
  assign n11693 = n3864 & ~n11312 ;
  assign n11694 = n10620 ^ n7507 ^ n1664 ;
  assign n11695 = n11694 ^ n10475 ^ 1'b0 ;
  assign n11696 = n11693 & n11695 ;
  assign n11697 = ~n7583 & n8332 ;
  assign n11698 = n7695 ^ n996 ^ 1'b0 ;
  assign n11699 = n1939 ^ n1538 ^ 1'b0 ;
  assign n11700 = n2943 & n11699 ;
  assign n11701 = ~n1098 & n11700 ;
  assign n11702 = n4765 | n10780 ;
  assign n11704 = n2474 | n2489 ;
  assign n11703 = n5753 ^ n3882 ^ 1'b0 ;
  assign n11705 = n11704 ^ n11703 ^ 1'b0 ;
  assign n11710 = n2733 & n6419 ;
  assign n11707 = n1870 ^ n610 ^ 1'b0 ;
  assign n11708 = n1564 & n11707 ;
  assign n11709 = ~n3176 & n11708 ;
  assign n11711 = n11710 ^ n11709 ^ 1'b0 ;
  assign n11712 = n11711 ^ n910 ^ 1'b0 ;
  assign n11713 = n7616 & n11712 ;
  assign n11714 = n11713 ^ n8522 ^ 1'b0 ;
  assign n11706 = n477 & n3001 ;
  assign n11715 = n11714 ^ n11706 ^ 1'b0 ;
  assign n11716 = ~n183 & n3374 ;
  assign n11717 = n11716 ^ n11131 ^ 1'b0 ;
  assign n11718 = n5477 ^ n5020 ^ 1'b0 ;
  assign n11719 = n6176 | n11718 ;
  assign n11720 = n287 | n11719 ;
  assign n11721 = n7066 & ~n11720 ;
  assign n11722 = n3912 ^ n220 ^ 1'b0 ;
  assign n11723 = n4066 & ~n11722 ;
  assign n11724 = ( n2157 & n3646 ) | ( n2157 & ~n11723 ) | ( n3646 & ~n11723 ) ;
  assign n11725 = n1276 & ~n9481 ;
  assign n11726 = n3514 & n11725 ;
  assign n11727 = ~n8594 & n11726 ;
  assign n11728 = n5636 & n8747 ;
  assign n11729 = n10019 & n11728 ;
  assign n11730 = ~n1020 & n7900 ;
  assign n11731 = n11730 ^ n8230 ^ 1'b0 ;
  assign n11732 = n11731 ^ n790 ^ n479 ;
  assign n11733 = n8279 ^ n6168 ^ n675 ;
  assign n11734 = n737 & ~n1967 ;
  assign n11735 = n11733 & n11734 ;
  assign n11737 = n3345 & n8911 ;
  assign n11736 = n4289 | n7591 ;
  assign n11738 = n11737 ^ n11736 ^ 1'b0 ;
  assign n11739 = n61 | n6556 ;
  assign n11740 = n11738 | n11739 ;
  assign n11741 = n3939 ^ n1505 ^ n1363 ;
  assign n11742 = n7110 | n11383 ;
  assign n11743 = n11742 ^ n11585 ^ 1'b0 ;
  assign n11744 = n1235 & ~n6232 ;
  assign n11745 = n2137 | n4916 ;
  assign n11746 = n152 & ~n9016 ;
  assign n11747 = n11746 ^ n7765 ^ 1'b0 ;
  assign n11748 = n11747 ^ n9884 ^ 1'b0 ;
  assign n11749 = n9260 | n11748 ;
  assign n11750 = n9812 ^ n8776 ^ n8703 ;
  assign n11751 = ~n651 & n11572 ;
  assign n11752 = n5795 ^ n5256 ^ 1'b0 ;
  assign n11753 = n454 | n2769 ;
  assign n11754 = n11753 ^ n8279 ^ 1'b0 ;
  assign n11755 = n1600 ^ n844 ^ 1'b0 ;
  assign n11756 = x3 & ~n676 ;
  assign n11757 = ~n11755 & n11756 ;
  assign n11758 = ~n3531 & n7238 ;
  assign n11759 = ( n1558 & n11757 ) | ( n1558 & n11758 ) | ( n11757 & n11758 ) ;
  assign n11760 = n3796 & n7627 ;
  assign n11761 = n3062 ^ n1238 ^ 1'b0 ;
  assign n11762 = n952 | n11281 ;
  assign n11763 = n74 & ~n11762 ;
  assign n11764 = n2145 | n2906 ;
  assign n11765 = n5083 ^ n4098 ^ 1'b0 ;
  assign n11766 = ( ~n5247 & n6600 ) | ( ~n5247 & n11765 ) | ( n6600 & n11765 ) ;
  assign n11770 = ~n1657 & n8026 ;
  assign n11767 = ~n3674 & n7024 ;
  assign n11768 = n11767 ^ n2547 ^ 1'b0 ;
  assign n11769 = n315 & n11768 ;
  assign n11771 = n11770 ^ n11769 ^ 1'b0 ;
  assign n11772 = n2122 & n2723 ;
  assign n11773 = n8695 ^ n226 ^ 1'b0 ;
  assign n11774 = n11772 | n11773 ;
  assign n11775 = n568 & n5933 ;
  assign n11776 = n11775 ^ n5308 ^ 1'b0 ;
  assign n11777 = ~n4291 & n8661 ;
  assign n11778 = ~n163 & n6757 ;
  assign n11779 = n11300 ^ n1465 ^ n291 ;
  assign n11780 = ~n11778 & n11779 ;
  assign n11781 = ~n4340 & n11780 ;
  assign n11782 = n11777 & n11781 ;
  assign n11783 = n9346 ^ n5454 ^ n4222 ;
  assign n11784 = n10287 ^ n3646 ^ 1'b0 ;
  assign n11785 = n10145 ^ n1235 ^ 1'b0 ;
  assign n11786 = n11784 & n11785 ;
  assign n11787 = n3402 & n6607 ;
  assign n11788 = n4066 & n11787 ;
  assign n11789 = n11788 ^ n1305 ^ 1'b0 ;
  assign n11790 = ~n2564 & n7464 ;
  assign n11791 = n10996 & ~n11790 ;
  assign n11792 = n8018 | n8884 ;
  assign n11793 = n7044 & n7973 ;
  assign n11794 = n11792 & n11793 ;
  assign n11795 = n1584 ^ n115 ^ 1'b0 ;
  assign n11796 = ~n3172 & n5227 ;
  assign n11797 = n2350 | n3780 ;
  assign n11798 = n4460 & ~n11797 ;
  assign n11799 = n4665 ^ n479 ^ 1'b0 ;
  assign n11800 = ~n2971 & n11799 ;
  assign n11801 = ~n5890 & n11238 ;
  assign n11802 = n5869 ^ n3942 ^ n1887 ;
  assign n11803 = ~n4153 & n8940 ;
  assign n11804 = n11803 ^ n1945 ^ 1'b0 ;
  assign n11805 = n11802 | n11804 ;
  assign n11806 = ~n8563 & n11747 ;
  assign n11807 = ~n1902 & n11806 ;
  assign n11808 = n6289 & ~n11807 ;
  assign n11809 = n11808 ^ n6839 ^ 1'b0 ;
  assign n11810 = n7861 ^ n1454 ^ 1'b0 ;
  assign n11811 = n1548 & n11810 ;
  assign n11812 = n5430 | n8500 ;
  assign n11813 = n4240 ^ n3686 ^ 1'b0 ;
  assign n11814 = ~n2634 & n5529 ;
  assign n11815 = n4359 & n11814 ;
  assign n11816 = ( ~n671 & n2855 ) | ( ~n671 & n6765 ) | ( n2855 & n6765 ) ;
  assign n11817 = n11816 ^ n3574 ^ 1'b0 ;
  assign n11818 = n6940 & n11817 ;
  assign n11819 = n9670 & n10008 ;
  assign n11820 = ( n1307 & n3314 ) | ( n1307 & n10886 ) | ( n3314 & n10886 ) ;
  assign n11821 = n11820 ^ n1134 ^ 1'b0 ;
  assign n11822 = n11819 | n11821 ;
  assign n11823 = ~n592 & n2807 ;
  assign n11824 = ~n1079 & n11823 ;
  assign n11825 = n11264 ^ n1300 ^ 1'b0 ;
  assign n11826 = n11825 ^ n782 ^ 1'b0 ;
  assign n11827 = n11826 ^ n5212 ^ 1'b0 ;
  assign n11828 = n11827 ^ n291 ^ 1'b0 ;
  assign n11829 = n11824 | n11828 ;
  assign n11830 = n5748 & n6337 ;
  assign n11831 = ~n6714 & n11830 ;
  assign n11832 = n9868 ^ n7376 ^ 1'b0 ;
  assign n11833 = n1679 & ~n10811 ;
  assign n11834 = ~n81 & n11833 ;
  assign n11835 = n5369 ^ n3372 ^ 1'b0 ;
  assign n11836 = ~n11834 & n11835 ;
  assign n11840 = n1863 | n3708 ;
  assign n11837 = n3699 ^ n1497 ^ 1'b0 ;
  assign n11838 = ( n1069 & n3218 ) | ( n1069 & ~n8773 ) | ( n3218 & ~n8773 ) ;
  assign n11839 = n11837 & n11838 ;
  assign n11841 = n11840 ^ n11839 ^ n343 ;
  assign n11845 = n495 | n717 ;
  assign n11842 = n5293 | n10319 ;
  assign n11843 = n9557 & ~n11842 ;
  assign n11844 = n9459 & ~n11843 ;
  assign n11846 = n11845 ^ n11844 ^ 1'b0 ;
  assign n11847 = n1728 & ~n11846 ;
  assign n11848 = n488 & n2358 ;
  assign n11849 = n5647 | n7753 ;
  assign n11852 = n15 | n373 ;
  assign n11850 = ( ~n135 & n1381 ) | ( ~n135 & n11527 ) | ( n1381 & n11527 ) ;
  assign n11851 = ~n2359 & n11850 ;
  assign n11853 = n11852 ^ n11851 ^ 1'b0 ;
  assign n11854 = n6316 & n6609 ;
  assign n11855 = n10793 ^ n6282 ^ 1'b0 ;
  assign n11856 = ~n10979 & n11855 ;
  assign n11857 = ~n9406 & n11856 ;
  assign n11858 = ~n4827 & n6404 ;
  assign n11859 = n846 & ~n3583 ;
  assign n11860 = ( n3833 & n7605 ) | ( n3833 & ~n11859 ) | ( n7605 & ~n11859 ) ;
  assign n11861 = n1111 ^ n862 ^ 1'b0 ;
  assign n11862 = n3847 & ~n6467 ;
  assign n11863 = n559 & n1187 ;
  assign n11864 = n11616 | n11863 ;
  assign n11865 = n11864 ^ n6360 ^ 1'b0 ;
  assign n11866 = n7791 ^ n7604 ^ 1'b0 ;
  assign n11867 = ~n11865 & n11866 ;
  assign n11868 = n11867 ^ n10812 ^ n9505 ;
  assign n11869 = ( n2951 & ~n5330 ) | ( n2951 & n5470 ) | ( ~n5330 & n5470 ) ;
  assign n11870 = n8101 ^ n6943 ^ 1'b0 ;
  assign n11871 = n6373 | n7576 ;
  assign n11872 = n11870 | n11871 ;
  assign n11873 = ~n219 & n8133 ;
  assign n11874 = n163 & n4707 ;
  assign n11875 = n1608 & ~n4059 ;
  assign n11876 = ( n5211 & n8161 ) | ( n5211 & n11875 ) | ( n8161 & n11875 ) ;
  assign n11877 = n9208 ^ n2560 ^ 1'b0 ;
  assign n11878 = n11876 | n11877 ;
  assign n11879 = n11878 ^ n7940 ^ 1'b0 ;
  assign n11880 = n3861 ^ n3623 ^ 1'b0 ;
  assign n11881 = n10029 & ~n11880 ;
  assign n11882 = n11881 ^ n4461 ^ 1'b0 ;
  assign n11883 = n7486 | n11882 ;
  assign n11884 = n6081 ^ n3455 ^ 1'b0 ;
  assign n11889 = n10890 ^ n3343 ^ 1'b0 ;
  assign n11890 = n4244 & ~n11889 ;
  assign n11885 = n1144 | n5740 ;
  assign n11886 = ~n387 & n11885 ;
  assign n11887 = n11886 ^ n4401 ^ 1'b0 ;
  assign n11888 = n8960 & ~n11887 ;
  assign n11891 = n11890 ^ n11888 ^ 1'b0 ;
  assign n11895 = n7362 ^ n4918 ^ 1'b0 ;
  assign n11896 = n3254 & ~n11895 ;
  assign n11892 = ~n2610 & n4017 ;
  assign n11893 = n11892 ^ n2512 ^ 1'b0 ;
  assign n11894 = n5211 | n11893 ;
  assign n11897 = n11896 ^ n11894 ^ 1'b0 ;
  assign n11898 = n7237 & ~n11897 ;
  assign n11899 = ~n2098 & n7147 ;
  assign n11904 = n295 & ~n2773 ;
  assign n11905 = n11904 ^ n5344 ^ 1'b0 ;
  assign n11900 = n1200 & ~n3147 ;
  assign n11901 = n3080 | n11900 ;
  assign n11902 = n11901 ^ n5348 ^ 1'b0 ;
  assign n11903 = n2775 & n11902 ;
  assign n11906 = n11905 ^ n11903 ^ 1'b0 ;
  assign n11908 = n1695 ^ n1603 ^ n1582 ;
  assign n11909 = ~n4539 & n11908 ;
  assign n11910 = n11909 ^ n4148 ^ 1'b0 ;
  assign n11911 = n5874 | n11910 ;
  assign n11907 = ( n1382 & n6509 ) | ( n1382 & n11225 ) | ( n6509 & n11225 ) ;
  assign n11912 = n11911 ^ n11907 ^ 1'b0 ;
  assign n11913 = n3589 & ~n11912 ;
  assign n11914 = n9048 & n11913 ;
  assign n11916 = n6748 ^ n5137 ^ 1'b0 ;
  assign n11915 = n4267 & ~n11008 ;
  assign n11917 = n11916 ^ n11915 ^ 1'b0 ;
  assign n11918 = n8336 ^ n2941 ^ n255 ;
  assign n11920 = n6176 ^ n2352 ^ 1'b0 ;
  assign n11921 = n11920 ^ n1282 ^ 1'b0 ;
  assign n11922 = ~n1271 & n11921 ;
  assign n11919 = n4220 | n9852 ;
  assign n11923 = n11922 ^ n11919 ^ 1'b0 ;
  assign n11924 = n595 ^ n225 ^ 1'b0 ;
  assign n11925 = n2763 & n11924 ;
  assign n11926 = n2495 & n11925 ;
  assign n11927 = n11926 ^ n1543 ^ 1'b0 ;
  assign n11928 = n2812 & ~n11927 ;
  assign n11929 = n10201 & ~n11928 ;
  assign n11930 = n11929 ^ n4180 ^ 1'b0 ;
  assign n11931 = n52 & n11930 ;
  assign n11933 = ~n2853 & n10610 ;
  assign n11934 = n11933 ^ n4015 ^ 1'b0 ;
  assign n11932 = n6012 ^ n4916 ^ 1'b0 ;
  assign n11935 = n11934 ^ n11932 ^ n1568 ;
  assign n11936 = n9279 ^ n2055 ^ 1'b0 ;
  assign n11937 = n4153 | n11936 ;
  assign n11938 = ~n1712 & n4626 ;
  assign n11939 = ~n1224 & n3167 ;
  assign n11940 = n3835 ^ n588 ^ 1'b0 ;
  assign n11941 = n1580 & n7408 ;
  assign n11942 = ~n11712 & n11941 ;
  assign n11943 = n11940 | n11942 ;
  assign n11944 = n2128 & ~n11552 ;
  assign n11945 = n9792 & n11944 ;
  assign n11946 = ~n3797 & n11945 ;
  assign n11947 = n11946 ^ n11605 ^ n7344 ;
  assign n11948 = n7152 ^ n4177 ^ n828 ;
  assign n11949 = ~n414 & n2894 ;
  assign n11950 = ~n4486 & n11949 ;
  assign n11951 = n11950 ^ n9410 ^ 1'b0 ;
  assign n11953 = n8852 ^ n33 ^ 1'b0 ;
  assign n11954 = n3212 & n11953 ;
  assign n11952 = ~n1430 & n5776 ;
  assign n11955 = n11954 ^ n11952 ^ 1'b0 ;
  assign n11956 = n3041 | n11955 ;
  assign n11957 = ~n597 & n7499 ;
  assign n11958 = n11957 ^ n4729 ^ 1'b0 ;
  assign n11959 = n9592 ^ n3095 ^ 1'b0 ;
  assign n11960 = n1718 ^ n732 ^ 1'b0 ;
  assign n11961 = n2359 ^ n961 ^ 1'b0 ;
  assign n11963 = n799 & n1370 ;
  assign n11964 = n326 & n11963 ;
  assign n11962 = n302 & n7735 ;
  assign n11965 = n11964 ^ n11962 ^ 1'b0 ;
  assign n11966 = n6528 & n11965 ;
  assign n11967 = ~n11961 & n11966 ;
  assign n11968 = ~n3334 & n8554 ;
  assign n11969 = n886 & ~n1688 ;
  assign n11970 = n10891 ^ n5442 ^ 1'b0 ;
  assign n11971 = n5254 & ~n11970 ;
  assign n11972 = n2494 & ~n7382 ;
  assign n11973 = n9563 ^ n6180 ^ 1'b0 ;
  assign n11974 = n5326 | n11973 ;
  assign n11975 = n5282 & ~n11974 ;
  assign n11976 = n2802 ^ n630 ^ 1'b0 ;
  assign n11977 = ~n1083 & n11976 ;
  assign n11978 = n11977 ^ n10333 ^ 1'b0 ;
  assign n11979 = n4122 ^ n997 ^ 1'b0 ;
  assign n11980 = n11979 ^ n10674 ^ n765 ;
  assign n11981 = n6864 ^ n5292 ^ 1'b0 ;
  assign n11982 = n11981 ^ n1312 ^ 1'b0 ;
  assign n11983 = n74 & ~n369 ;
  assign n11984 = ~n74 & n11983 ;
  assign n11985 = n2403 | n3056 ;
  assign n11986 = n2403 & ~n11985 ;
  assign n11987 = n11986 ^ n3437 ^ 1'b0 ;
  assign n11988 = n11984 & n11987 ;
  assign n11989 = n7398 ^ n712 ^ 1'b0 ;
  assign n11990 = n11988 & n11989 ;
  assign n11991 = n11982 & n11990 ;
  assign n11992 = ~n11982 & n11991 ;
  assign n11993 = n11194 & ~n11992 ;
  assign n11994 = n10403 ^ n5490 ^ 1'b0 ;
  assign n11995 = ~n1386 & n11994 ;
  assign n11996 = n11995 ^ n10161 ^ n2427 ;
  assign n11997 = n10946 ^ n7877 ^ 1'b0 ;
  assign n11998 = ( n11993 & n11996 ) | ( n11993 & n11997 ) | ( n11996 & n11997 ) ;
  assign n11999 = ~n8660 & n10767 ;
  assign n12000 = ~n7000 & n9191 ;
  assign n12001 = n2859 | n3137 ;
  assign n12002 = n6732 | n12001 ;
  assign n12003 = ~n3565 & n12002 ;
  assign n12004 = n560 | n8771 ;
  assign n12005 = n8949 ^ n2840 ^ 1'b0 ;
  assign n12006 = n12005 ^ n5364 ^ 1'b0 ;
  assign n12007 = ( ~n1251 & n4935 ) | ( ~n1251 & n10246 ) | ( n4935 & n10246 ) ;
  assign n12008 = n7146 ^ n1507 ^ n1304 ;
  assign n12009 = n12008 ^ n11555 ^ 1'b0 ;
  assign n12010 = n8432 ^ n4831 ^ 1'b0 ;
  assign n12011 = n7391 & ~n12010 ;
  assign n12022 = ~n2244 & n6806 ;
  assign n12021 = n5213 | n6556 ;
  assign n12023 = n12022 ^ n12021 ^ 1'b0 ;
  assign n12019 = ~n5573 & n9023 ;
  assign n12020 = n12019 ^ n8181 ^ 1'b0 ;
  assign n12024 = n12023 ^ n12020 ^ 1'b0 ;
  assign n12016 = n1313 | n4116 ;
  assign n12014 = n5151 ^ n1750 ^ 1'b0 ;
  assign n12015 = n1142 & ~n12014 ;
  assign n12012 = x8 & n604 ;
  assign n12013 = ~n225 & n12012 ;
  assign n12017 = n12016 ^ n12015 ^ n12013 ;
  assign n12018 = n12017 ^ n7949 ^ n5783 ;
  assign n12025 = n12024 ^ n12018 ^ n9808 ;
  assign n12026 = n12025 ^ n6233 ^ 1'b0 ;
  assign n12027 = n1065 & ~n1469 ;
  assign n12028 = n12027 ^ n3040 ^ 1'b0 ;
  assign n12029 = n12028 ^ n4819 ^ 1'b0 ;
  assign n12030 = n8267 & n12029 ;
  assign n12031 = n2173 & n8904 ;
  assign n12032 = ~n11462 & n12031 ;
  assign n12033 = n4160 | n7643 ;
  assign n12034 = n12033 ^ n10411 ^ 1'b0 ;
  assign n12035 = n5865 | n8591 ;
  assign n12036 = n12035 ^ n10861 ^ 1'b0 ;
  assign n12037 = n58 & ~n10437 ;
  assign n12038 = n8440 | n11294 ;
  assign n12039 = n2444 ^ n2337 ^ 1'b0 ;
  assign n12040 = ~n5047 & n12039 ;
  assign n12041 = n5528 & n7823 ;
  assign n12042 = n5638 & ~n12041 ;
  assign n12043 = n12042 ^ n4618 ^ 1'b0 ;
  assign n12044 = ~n2291 & n6538 ;
  assign n12045 = ~n1050 & n12044 ;
  assign n12046 = n9511 | n12045 ;
  assign n12047 = n5393 ^ n3133 ^ n1354 ;
  assign n12048 = n6576 | n12047 ;
  assign n12049 = n12048 ^ n5138 ^ 1'b0 ;
  assign n12050 = n10694 ^ n8865 ^ 1'b0 ;
  assign n12051 = n7375 & ~n12050 ;
  assign n12052 = n5199 & n12051 ;
  assign n12053 = n12049 & ~n12052 ;
  assign n12054 = n1997 | n6065 ;
  assign n12055 = n1329 & ~n12054 ;
  assign n12056 = n3564 | n12055 ;
  assign n12057 = n9479 ^ n1334 ^ 1'b0 ;
  assign n12058 = ~n5458 & n12057 ;
  assign n12059 = ( n1764 & ~n1816 ) | ( n1764 & n6427 ) | ( ~n1816 & n6427 ) ;
  assign n12060 = n12059 ^ n4634 ^ 1'b0 ;
  assign n12061 = ~n1305 & n3660 ;
  assign n12062 = n12061 ^ n61 ^ 1'b0 ;
  assign n12063 = n3723 | n6575 ;
  assign n12064 = n12062 & ~n12063 ;
  assign n12065 = n12064 ^ n7515 ^ 1'b0 ;
  assign n12072 = ( n3013 & n3191 ) | ( n3013 & ~n5644 ) | ( n3191 & ~n5644 ) ;
  assign n12068 = n11423 ^ n4589 ^ 1'b0 ;
  assign n12069 = n9406 & ~n12068 ;
  assign n12066 = ~n5057 & n7170 ;
  assign n12067 = ~n5079 & n12066 ;
  assign n12070 = n12069 ^ n12067 ^ 1'b0 ;
  assign n12071 = n5745 | n12070 ;
  assign n12073 = n12072 ^ n12071 ^ 1'b0 ;
  assign n12074 = ~n183 & n1528 ;
  assign n12075 = ~n805 & n12074 ;
  assign n12076 = ~n3718 & n12075 ;
  assign n12077 = n12076 ^ n7978 ^ 1'b0 ;
  assign n12078 = n12073 & ~n12077 ;
  assign n12079 = n2146 ^ n1377 ^ 1'b0 ;
  assign n12080 = n6344 & ~n6542 ;
  assign n12081 = n12080 ^ n2980 ^ 1'b0 ;
  assign n12082 = n4540 | n10864 ;
  assign n12083 = n5697 ^ n1915 ^ 1'b0 ;
  assign n12084 = n1058 | n12083 ;
  assign n12085 = n3349 | n12084 ;
  assign n12086 = n2529 & ~n12085 ;
  assign n12087 = n3350 & ~n9322 ;
  assign n12088 = n12087 ^ n2991 ^ 1'b0 ;
  assign n12089 = n12088 ^ n2664 ^ 1'b0 ;
  assign n12090 = ~n1898 & n12089 ;
  assign n12091 = n7919 & ~n12090 ;
  assign n12092 = n934 | n1029 ;
  assign n12094 = n8215 ^ n6576 ^ 1'b0 ;
  assign n12093 = ~n1207 & n4001 ;
  assign n12095 = n12094 ^ n12093 ^ 1'b0 ;
  assign n12096 = ( n259 & n2618 ) | ( n259 & n5379 ) | ( n2618 & n5379 ) ;
  assign n12097 = n8998 & ~n12096 ;
  assign n12098 = ~n9933 & n12097 ;
  assign n12099 = n480 | n12098 ;
  assign n12100 = n3384 ^ n2749 ^ 1'b0 ;
  assign n12101 = ~n5759 & n12100 ;
  assign n12102 = n9410 ^ n4429 ^ 1'b0 ;
  assign n12103 = n212 & ~n12102 ;
  assign n12104 = n12103 ^ n3852 ^ 1'b0 ;
  assign n12105 = n1148 | n6401 ;
  assign n12106 = ( n181 & ~n11225 ) | ( n181 & n12105 ) | ( ~n11225 & n12105 ) ;
  assign n12107 = n2637 ^ n195 ^ 1'b0 ;
  assign n12108 = n4718 | n9508 ;
  assign n12109 = n1379 | n12108 ;
  assign n12110 = n1416 & n12109 ;
  assign n12111 = n12110 ^ n11253 ^ 1'b0 ;
  assign n12112 = n1047 & n12111 ;
  assign n12113 = ~n1451 & n12112 ;
  assign n12114 = n6797 ^ n5313 ^ 1'b0 ;
  assign n12116 = ~n1645 & n7448 ;
  assign n12115 = n11167 ^ n7033 ^ 1'b0 ;
  assign n12117 = n12116 ^ n12115 ^ 1'b0 ;
  assign n12118 = n4136 ^ n1329 ^ 1'b0 ;
  assign n12119 = n3442 | n12118 ;
  assign n12120 = n667 | n2433 ;
  assign n12121 = ~n8668 & n12120 ;
  assign n12122 = n12121 ^ n9436 ^ 1'b0 ;
  assign n12123 = n5663 | n9643 ;
  assign n12129 = n4960 ^ n4804 ^ 1'b0 ;
  assign n12130 = n2326 | n12129 ;
  assign n12131 = n4326 & ~n12130 ;
  assign n12124 = n1936 ^ n1245 ^ n415 ;
  assign n12125 = n5629 ^ n257 ^ 1'b0 ;
  assign n12126 = ( n2100 & ~n4111 ) | ( n2100 & n12125 ) | ( ~n4111 & n12125 ) ;
  assign n12127 = n12124 & ~n12126 ;
  assign n12128 = n12127 ^ n4859 ^ 1'b0 ;
  assign n12132 = n12131 ^ n12128 ^ 1'b0 ;
  assign n12133 = n5867 ^ n5587 ^ 1'b0 ;
  assign n12134 = n3284 | n11138 ;
  assign n12137 = n271 ^ n33 ^ 1'b0 ;
  assign n12135 = n1742 ^ n1353 ^ 1'b0 ;
  assign n12136 = n1146 | n12135 ;
  assign n12138 = n12137 ^ n12136 ^ 1'b0 ;
  assign n12139 = n7895 ^ n4797 ^ 1'b0 ;
  assign n12140 = n11938 | n12139 ;
  assign n12141 = n12140 ^ n3078 ^ 1'b0 ;
  assign n12142 = n11755 ^ n6347 ^ 1'b0 ;
  assign n12143 = n7687 & ~n12142 ;
  assign n12144 = n12143 ^ n183 ^ 1'b0 ;
  assign n12145 = ~n4218 & n11358 ;
  assign n12148 = n5463 ^ n1403 ^ 1'b0 ;
  assign n12149 = n9812 | n12148 ;
  assign n12146 = n924 & n8325 ;
  assign n12147 = ~n7743 & n12146 ;
  assign n12150 = n12149 ^ n12147 ^ 1'b0 ;
  assign n12151 = n1988 & ~n12150 ;
  assign n12152 = n12151 ^ n1141 ^ 1'b0 ;
  assign n12153 = n3686 ^ n331 ^ 1'b0 ;
  assign n12154 = n12152 & ~n12153 ;
  assign n12155 = n5663 ^ n2637 ^ 1'b0 ;
  assign n12156 = n11482 ^ n4719 ^ 1'b0 ;
  assign n12158 = n6671 ^ n1731 ^ 1'b0 ;
  assign n12159 = n2114 | n12158 ;
  assign n12157 = n2769 ^ n2630 ^ 1'b0 ;
  assign n12160 = n12159 ^ n12157 ^ 1'b0 ;
  assign n12161 = n5745 | n7354 ;
  assign n12162 = n12161 ^ n3472 ^ 1'b0 ;
  assign n12163 = n360 & ~n8188 ;
  assign n12164 = n12163 ^ n7079 ^ 1'b0 ;
  assign n12165 = ~n3724 & n12164 ;
  assign n12166 = n1842 | n11387 ;
  assign n12167 = ( n4093 & ~n6012 ) | ( n4093 & n6584 ) | ( ~n6012 & n6584 ) ;
  assign n12168 = n7460 & ~n12167 ;
  assign n12169 = n10963 ^ n967 ^ 1'b0 ;
  assign n12170 = n10900 | n12169 ;
  assign n12171 = n12170 ^ n2647 ^ 1'b0 ;
  assign n12172 = n9606 ^ n7778 ^ n5240 ;
  assign n12173 = n8068 & n12172 ;
  assign n12174 = n4855 & ~n12173 ;
  assign n12175 = ~n1374 & n12174 ;
  assign n12176 = n11318 ^ n3949 ^ 1'b0 ;
  assign n12177 = n8688 ^ n7588 ^ 1'b0 ;
  assign n12178 = n10066 ^ n1912 ^ 1'b0 ;
  assign n12179 = n12178 ^ n5385 ^ 1'b0 ;
  assign n12180 = n6307 & n6670 ;
  assign n12181 = n8797 ^ n4044 ^ 1'b0 ;
  assign n12182 = n2749 & n5681 ;
  assign n12183 = n1147 & n12182 ;
  assign n12184 = n12183 ^ n9580 ^ 1'b0 ;
  assign n12185 = n4340 & ~n12184 ;
  assign n12186 = n5549 ^ n3437 ^ 1'b0 ;
  assign n12187 = n12185 & ~n12186 ;
  assign n12188 = n2045 ^ n1118 ^ 1'b0 ;
  assign n12189 = n7922 & n12188 ;
  assign n12190 = n3355 ^ n331 ^ 1'b0 ;
  assign n12191 = n12190 ^ n747 ^ 1'b0 ;
  assign n12192 = n3992 & n12191 ;
  assign n12193 = n8037 & n12192 ;
  assign n12194 = n4088 & ~n5929 ;
  assign n12195 = n12193 & n12194 ;
  assign n12196 = n12195 ^ n5606 ^ n3072 ;
  assign n12197 = n4478 ^ n2040 ^ 1'b0 ;
  assign n12198 = ~n535 & n1507 ;
  assign n12199 = n3305 & n6056 ;
  assign n12200 = n1715 & n12199 ;
  assign n12201 = ~n4017 & n12200 ;
  assign n12202 = n5396 ^ n175 ^ 1'b0 ;
  assign n12205 = n8534 & n10720 ;
  assign n12206 = n12205 ^ n1538 ^ 1'b0 ;
  assign n12203 = n809 & ~n8168 ;
  assign n12204 = n12203 ^ n6198 ^ 1'b0 ;
  assign n12207 = n12206 ^ n12204 ^ 1'b0 ;
  assign n12208 = n12202 & ~n12207 ;
  assign n12212 = n806 & ~n6039 ;
  assign n12213 = n12212 ^ n886 ^ 1'b0 ;
  assign n12210 = n3490 & n7087 ;
  assign n12211 = n12210 ^ n2873 ^ 1'b0 ;
  assign n12214 = n12213 ^ n12211 ^ n45 ;
  assign n12209 = ~n447 & n11107 ;
  assign n12215 = n12214 ^ n12209 ^ n9252 ;
  assign n12216 = n4082 | n6074 ;
  assign n12217 = n12216 ^ n10682 ^ 1'b0 ;
  assign n12221 = n3873 & n4895 ;
  assign n12218 = n4675 ^ n1876 ^ 1'b0 ;
  assign n12219 = n12218 ^ n6430 ^ 1'b0 ;
  assign n12220 = ~n9364 & n12219 ;
  assign n12222 = n12221 ^ n12220 ^ 1'b0 ;
  assign n12224 = n6966 | n8580 ;
  assign n12223 = n1603 | n5363 ;
  assign n12225 = n12224 ^ n12223 ^ 1'b0 ;
  assign n12226 = ( n5908 & ~n9839 ) | ( n5908 & n9946 ) | ( ~n9839 & n9946 ) ;
  assign n12227 = n6608 | n12226 ;
  assign n12228 = n12227 ^ n6999 ^ 1'b0 ;
  assign n12229 = n6669 & n12228 ;
  assign n12230 = n12229 ^ n5981 ^ 1'b0 ;
  assign n12233 = n1667 ^ n497 ^ 1'b0 ;
  assign n12231 = ~n2139 & n3375 ;
  assign n12232 = n1161 | n12231 ;
  assign n12234 = n12233 ^ n12232 ^ 1'b0 ;
  assign n12235 = n5860 ^ n2040 ^ 1'b0 ;
  assign n12236 = n8580 | n12235 ;
  assign n12237 = n7544 ^ n5360 ^ n291 ;
  assign n12238 = n1590 | n8553 ;
  assign n12239 = n1121 | n1933 ;
  assign n12240 = ( n135 & ~n205 ) | ( n135 & n488 ) | ( ~n205 & n488 ) ;
  assign n12241 = n4511 & ~n12045 ;
  assign n12242 = ~n12240 & n12241 ;
  assign n12243 = ( n3584 & n7254 ) | ( n3584 & ~n12242 ) | ( n7254 & ~n12242 ) ;
  assign n12244 = ( ~n9716 & n12239 ) | ( ~n9716 & n12243 ) | ( n12239 & n12243 ) ;
  assign n12245 = n5141 & ~n5685 ;
  assign n12246 = ~n237 & n12245 ;
  assign n12247 = n562 | n2719 ;
  assign n12248 = n12246 & ~n12247 ;
  assign n12249 = ( ~n1462 & n1821 ) | ( ~n1462 & n3736 ) | ( n1821 & n3736 ) ;
  assign n12250 = n954 & n3935 ;
  assign n12251 = ~n4216 & n12250 ;
  assign n12252 = n12249 | n12251 ;
  assign n12253 = n12248 & ~n12252 ;
  assign n12254 = n2227 & n3279 ;
  assign n12255 = n5839 ^ n235 ^ 1'b0 ;
  assign n12256 = n135 | n12255 ;
  assign n12257 = n2549 | n8378 ;
  assign n12258 = n12256 & ~n12257 ;
  assign n12259 = n2350 ^ n1556 ^ 1'b0 ;
  assign n12260 = ~n3894 & n12259 ;
  assign n12261 = n6073 & ~n12260 ;
  assign n12262 = n12258 & n12261 ;
  assign n12263 = n8715 | n12262 ;
  assign n12264 = n12254 | n12263 ;
  assign n12265 = n4399 ^ n2010 ^ n372 ;
  assign n12266 = n12265 ^ n243 ^ 1'b0 ;
  assign n12267 = n1336 & n12266 ;
  assign n12268 = n12267 ^ n367 ^ 1'b0 ;
  assign n12269 = n1978 & n12268 ;
  assign n12270 = n12269 ^ n9497 ^ 1'b0 ;
  assign n12271 = n4852 ^ n4460 ^ 1'b0 ;
  assign n12272 = n2019 | n2785 ;
  assign n12273 = n6888 | n12272 ;
  assign n12274 = n12273 ^ n4136 ^ 1'b0 ;
  assign n12275 = ~n8940 & n10703 ;
  assign n12276 = ~n2326 & n10162 ;
  assign n12277 = ~n11221 & n12276 ;
  assign n12278 = n3479 & ~n12277 ;
  assign n12279 = n12275 & n12278 ;
  assign n12280 = ( n1677 & n3565 ) | ( n1677 & ~n6588 ) | ( n3565 & ~n6588 ) ;
  assign n12281 = n2048 | n12280 ;
  assign n12282 = n12281 ^ n8407 ^ 1'b0 ;
  assign n12283 = n1286 ^ n625 ^ 1'b0 ;
  assign n12284 = n4727 ^ n3933 ^ 1'b0 ;
  assign n12285 = n4135 | n12284 ;
  assign n12286 = n8919 ^ n4605 ^ 1'b0 ;
  assign n12287 = ~n2678 & n3284 ;
  assign n12288 = ~n12286 & n12287 ;
  assign n12289 = n1413 | n8675 ;
  assign n12290 = ~n447 & n1591 ;
  assign n12291 = n12290 ^ n9139 ^ 1'b0 ;
  assign n12293 = n2668 | n7261 ;
  assign n12292 = ~n654 & n9495 ;
  assign n12294 = n12293 ^ n12292 ^ n1336 ;
  assign n12295 = n4446 ^ n3374 ^ 1'b0 ;
  assign n12296 = n12077 & ~n12295 ;
  assign n12297 = n8273 & n12296 ;
  assign n12298 = n8976 ^ n2893 ^ 1'b0 ;
  assign n12299 = ( n659 & n1244 ) | ( n659 & ~n11852 ) | ( n1244 & ~n11852 ) ;
  assign n12300 = n12299 ^ n1505 ^ n376 ;
  assign n12301 = n4218 ^ n2758 ^ 1'b0 ;
  assign n12302 = n4990 ^ n1679 ^ 1'b0 ;
  assign n12303 = ~n3845 & n11172 ;
  assign n12304 = n12303 ^ n8552 ^ 1'b0 ;
  assign n12305 = n12302 | n12304 ;
  assign n12306 = n4977 ^ n2697 ^ 1'b0 ;
  assign n12307 = n793 | n12306 ;
  assign n12308 = n2143 & ~n9189 ;
  assign n12309 = ~n3982 & n12308 ;
  assign n12311 = n5681 ^ n541 ^ 1'b0 ;
  assign n12312 = n7725 & ~n12311 ;
  assign n12313 = n2773 ^ n2533 ^ 1'b0 ;
  assign n12314 = n12312 & ~n12313 ;
  assign n12310 = n1514 | n8759 ;
  assign n12315 = n12314 ^ n12310 ^ 1'b0 ;
  assign n12316 = ~n12309 & n12315 ;
  assign n12317 = n5451 & n12316 ;
  assign n12318 = n9264 ^ n3644 ^ 1'b0 ;
  assign n12319 = ~n1247 & n12318 ;
  assign n12320 = ~n1329 & n11009 ;
  assign n12321 = n12320 ^ n7416 ^ 1'b0 ;
  assign n12322 = ( n8844 & n9198 ) | ( n8844 & n9955 ) | ( n9198 & n9955 ) ;
  assign n12323 = ~n439 & n1944 ;
  assign n12324 = ~n8012 & n12323 ;
  assign n12325 = n6714 & n11305 ;
  assign n12326 = ~n12056 & n12325 ;
  assign n12327 = ( n533 & n541 ) | ( n533 & n2120 ) | ( n541 & n2120 ) ;
  assign n12328 = n12327 ^ n8130 ^ 1'b0 ;
  assign n12329 = n12328 ^ n5001 ^ 1'b0 ;
  assign n12330 = ~n8406 & n12329 ;
  assign n12331 = ~n1697 & n4492 ;
  assign n12332 = n4089 & n12331 ;
  assign n12333 = n12332 ^ n9381 ^ 1'b0 ;
  assign n12334 = n8105 & ~n9605 ;
  assign n12335 = n1177 & n12334 ;
  assign n12336 = n1703 | n12335 ;
  assign n12337 = n2927 | n12336 ;
  assign n12338 = n12337 ^ n4106 ^ 1'b0 ;
  assign n12339 = n5333 ^ n1724 ^ n91 ;
  assign n12340 = n12339 ^ n12155 ^ 1'b0 ;
  assign n12341 = n4984 ^ n3738 ^ n845 ;
  assign n12342 = n12341 ^ n2605 ^ 1'b0 ;
  assign n12343 = ~n1167 & n12342 ;
  assign n12344 = n3324 ^ n903 ^ 1'b0 ;
  assign n12345 = n3088 & n8308 ;
  assign n12346 = n1845 & ~n3779 ;
  assign n12347 = ~n12345 & n12346 ;
  assign n12348 = n5033 & n11087 ;
  assign n12349 = ~n6500 & n12348 ;
  assign n12350 = n3239 & n12349 ;
  assign n12352 = n825 | n1976 ;
  assign n12353 = n2989 & ~n12352 ;
  assign n12351 = n3153 | n4571 ;
  assign n12354 = n12353 ^ n12351 ^ 1'b0 ;
  assign n12355 = n2918 & ~n3202 ;
  assign n12356 = ~n4378 & n12355 ;
  assign n12357 = n7577 ^ n4104 ^ n3794 ;
  assign n12358 = ~n4311 & n12357 ;
  assign n12359 = n484 & ~n8201 ;
  assign n12360 = ~n746 & n12359 ;
  assign n12361 = n1877 ^ n122 ^ 1'b0 ;
  assign n12362 = ~n3054 & n6227 ;
  assign n12363 = n4589 & n12362 ;
  assign n12364 = n12363 ^ n940 ^ 1'b0 ;
  assign n12365 = n6447 | n8660 ;
  assign n12366 = n9286 ^ n6059 ^ x0 ;
  assign n12367 = n7135 ^ n6110 ^ 1'b0 ;
  assign n12368 = n8482 & n12367 ;
  assign n12369 = ( n2554 & ~n12366 ) | ( n2554 & n12368 ) | ( ~n12366 & n12368 ) ;
  assign n12370 = n11907 ^ n10840 ^ 1'b0 ;
  assign n12371 = n11120 & n12370 ;
  assign n12372 = n6106 ^ n562 ^ 1'b0 ;
  assign n12373 = ~n8222 & n12372 ;
  assign n12374 = ~n1530 & n12373 ;
  assign n12375 = n2122 & n7109 ;
  assign n12376 = ~n175 & n11064 ;
  assign n12377 = ~n4636 & n11170 ;
  assign n12378 = n2749 & ~n12377 ;
  assign n12379 = n6431 & n12378 ;
  assign n12380 = n1599 | n1705 ;
  assign n12381 = n12380 ^ n2465 ^ 1'b0 ;
  assign n12382 = n12379 | n12381 ;
  assign n12383 = n7185 ^ n3186 ^ n1264 ;
  assign n12384 = n7208 & n8441 ;
  assign n12385 = ~n7631 & n12384 ;
  assign n12386 = n11323 | n12385 ;
  assign n12387 = n12386 ^ n2915 ^ 1'b0 ;
  assign n12388 = ~n112 & n2438 ;
  assign n12389 = n12388 ^ n1049 ^ 1'b0 ;
  assign n12390 = ~n10357 & n12389 ;
  assign n12391 = ~n9766 & n12390 ;
  assign n12392 = n5052 & n6415 ;
  assign n12393 = n1269 ^ n773 ^ 1'b0 ;
  assign n12394 = n12393 ^ n7063 ^ 1'b0 ;
  assign n12395 = n12392 & ~n12394 ;
  assign n12399 = n1155 | n5865 ;
  assign n12400 = n12399 ^ n1863 ^ 1'b0 ;
  assign n12401 = n6474 & n8132 ;
  assign n12402 = n12401 ^ n121 ^ 1'b0 ;
  assign n12403 = n12402 ^ n10366 ^ n8539 ;
  assign n12404 = n12400 | n12403 ;
  assign n12396 = n4646 ^ n144 ^ 1'b0 ;
  assign n12397 = n9082 | n12396 ;
  assign n12398 = n2653 & ~n12397 ;
  assign n12405 = n12404 ^ n12398 ^ 1'b0 ;
  assign n12406 = n8629 & n8891 ;
  assign n12407 = n7674 | n10246 ;
  assign n12408 = n1854 & n3218 ;
  assign n12409 = n1760 & n3306 ;
  assign n12410 = n4993 ^ n4837 ^ 1'b0 ;
  assign n12411 = n12409 & n12410 ;
  assign n12412 = n8126 ^ n4519 ^ n2709 ;
  assign n12413 = n5348 & ~n12412 ;
  assign n12414 = n1663 & ~n8886 ;
  assign n12415 = n12414 ^ n1211 ^ 1'b0 ;
  assign n12416 = n27 | n9085 ;
  assign n12417 = n5706 & ~n12416 ;
  assign n12418 = n12417 ^ n4377 ^ 1'b0 ;
  assign n12419 = n10432 ^ n2044 ^ 1'b0 ;
  assign n12420 = n3735 & ~n12043 ;
  assign n12421 = ~n4435 & n12420 ;
  assign n12424 = n409 & ~n1591 ;
  assign n12422 = n695 & ~n6993 ;
  assign n12423 = n12422 ^ n10837 ^ n547 ;
  assign n12425 = n12424 ^ n12423 ^ n2505 ;
  assign n12426 = n6102 ^ n4040 ^ n3054 ;
  assign n12427 = n6271 | n12426 ;
  assign n12428 = n788 & ~n12427 ;
  assign n12429 = n2252 ^ n2070 ^ 1'b0 ;
  assign n12430 = n3502 & n12429 ;
  assign n12431 = ~n4389 & n10038 ;
  assign n12432 = n12431 ^ n8229 ^ 1'b0 ;
  assign n12433 = n12430 & ~n12432 ;
  assign n12434 = n4451 ^ n553 ^ 1'b0 ;
  assign n12435 = ~n7884 & n12434 ;
  assign n12436 = n12435 ^ n8000 ^ n1667 ;
  assign n12437 = n2671 ^ n2653 ^ 1'b0 ;
  assign n12438 = ~n12436 & n12437 ;
  assign n12439 = n4333 ^ n3006 ^ 1'b0 ;
  assign n12440 = n1191 & ~n12439 ;
  assign n12441 = ( ~n3928 & n4741 ) | ( ~n3928 & n12440 ) | ( n4741 & n12440 ) ;
  assign n12442 = ( n4731 & ~n5305 ) | ( n4731 & n7067 ) | ( ~n5305 & n7067 ) ;
  assign n12443 = n9423 & n12442 ;
  assign n12444 = ~n12441 & n12443 ;
  assign n12445 = n4576 & ~n5839 ;
  assign n12446 = ~n675 & n12445 ;
  assign n12447 = n3913 ^ n3003 ^ n753 ;
  assign n12448 = n1131 | n12447 ;
  assign n12449 = ~n1132 & n7053 ;
  assign n12450 = n10715 ^ n7170 ^ n2288 ;
  assign n12451 = n12449 | n12450 ;
  assign n12452 = n9286 ^ n3202 ^ 1'b0 ;
  assign n12453 = n5769 & n12452 ;
  assign n12454 = n6267 | n7405 ;
  assign n12455 = n12453 | n12454 ;
  assign n12456 = n9511 & n12455 ;
  assign n12457 = n11281 ^ n527 ^ 1'b0 ;
  assign n12458 = n6383 | n12457 ;
  assign n12459 = ~n1971 & n11001 ;
  assign n12460 = n5041 & n12459 ;
  assign n12461 = n11253 ^ n4645 ^ 1'b0 ;
  assign n12462 = n6781 & ~n11366 ;
  assign n12463 = n796 & n12462 ;
  assign n12464 = n3651 ^ n2328 ^ 1'b0 ;
  assign n12465 = n221 & ~n12464 ;
  assign n12466 = n12465 ^ n3571 ^ 1'b0 ;
  assign n12467 = n2359 ^ n957 ^ n541 ;
  assign n12468 = n12467 ^ n9343 ^ 1'b0 ;
  assign n12469 = n12468 ^ n8604 ^ 1'b0 ;
  assign n12470 = ~n6928 & n12469 ;
  assign n12471 = ~n6874 & n7530 ;
  assign n12472 = n3817 & n4279 ;
  assign n12473 = n7962 & n8077 ;
  assign n12474 = n12473 ^ n6554 ^ 1'b0 ;
  assign n12475 = ( n12471 & ~n12472 ) | ( n12471 & n12474 ) | ( ~n12472 & n12474 ) ;
  assign n12476 = n11525 ^ n2645 ^ 1'b0 ;
  assign n12477 = ~n12475 & n12476 ;
  assign n12478 = n9536 & n11668 ;
  assign n12479 = n1848 & n12478 ;
  assign n12480 = ~n3349 & n11491 ;
  assign n12481 = ~n10667 & n12480 ;
  assign n12482 = n12479 & n12481 ;
  assign n12483 = ( n479 & ~n3388 ) | ( n479 & n7029 ) | ( ~n3388 & n7029 ) ;
  assign n12484 = ( n372 & n403 ) | ( n372 & n5616 ) | ( n403 & n5616 ) ;
  assign n12485 = n12484 ^ n7932 ^ 1'b0 ;
  assign n12486 = n117 | n4696 ;
  assign n12487 = n12486 ^ n5554 ^ 1'b0 ;
  assign n12488 = n12487 ^ n7534 ^ 1'b0 ;
  assign n12489 = n4999 & ~n5391 ;
  assign n12490 = n12489 ^ n1469 ^ 1'b0 ;
  assign n12491 = n6385 & ~n7100 ;
  assign n12492 = ~n163 & n12491 ;
  assign n12493 = n1523 | n12492 ;
  assign n12494 = n3216 | n12493 ;
  assign n12495 = ( n1242 & n11390 ) | ( n1242 & n12494 ) | ( n11390 & n12494 ) ;
  assign n12496 = x2 & n3299 ;
  assign n12497 = n4764 ^ n4567 ^ 1'b0 ;
  assign n12498 = ~n5916 & n7209 ;
  assign n12499 = n12498 ^ n3678 ^ 1'b0 ;
  assign n12506 = n995 | n9804 ;
  assign n12507 = n12506 ^ n112 ^ 1'b0 ;
  assign n12508 = n4251 & ~n12507 ;
  assign n12509 = n11185 & n12508 ;
  assign n12500 = n4331 & ~n7986 ;
  assign n12501 = n5317 & n12500 ;
  assign n12502 = n12501 ^ n239 ^ 1'b0 ;
  assign n12503 = ~n540 & n2140 ;
  assign n12504 = ( n3232 & n12502 ) | ( n3232 & n12503 ) | ( n12502 & n12503 ) ;
  assign n12505 = n4583 & n12504 ;
  assign n12510 = n12509 ^ n12505 ^ 1'b0 ;
  assign n12511 = ~n1439 & n5114 ;
  assign n12512 = n12511 ^ n1674 ^ 1'b0 ;
  assign n12513 = ~n927 & n12512 ;
  assign n12514 = n12513 ^ n9698 ^ n253 ;
  assign n12515 = n646 | n815 ;
  assign n12516 = n12515 ^ n9293 ^ 1'b0 ;
  assign n12517 = n12514 | n12516 ;
  assign n12518 = n555 & ~n7137 ;
  assign n12519 = ( n229 & ~n8730 ) | ( n229 & n12518 ) | ( ~n8730 & n12518 ) ;
  assign n12520 = n1904 ^ n1460 ^ 1'b0 ;
  assign n12521 = ~n2055 & n10941 ;
  assign n12522 = ~n6119 & n7544 ;
  assign n12523 = n9874 & n12522 ;
  assign n12526 = n4819 & ~n4894 ;
  assign n12527 = ~n2388 & n7510 ;
  assign n12528 = ~n12526 & n12527 ;
  assign n12524 = n3638 & n5665 ;
  assign n12525 = n12524 ^ n4401 ^ 1'b0 ;
  assign n12529 = n12528 ^ n12525 ^ 1'b0 ;
  assign n12530 = ~n2444 & n3952 ;
  assign n12531 = n12529 & n12530 ;
  assign n12532 = ~n9525 & n11461 ;
  assign n12533 = n12532 ^ n6902 ^ 1'b0 ;
  assign n12534 = n891 | n3434 ;
  assign n12535 = n3172 ^ n2824 ^ 1'b0 ;
  assign n12539 = n959 & n1182 ;
  assign n12540 = n12539 ^ n591 ^ 1'b0 ;
  assign n12536 = ~n3672 & n8667 ;
  assign n12537 = n12536 ^ n2213 ^ 1'b0 ;
  assign n12538 = n6768 & n12537 ;
  assign n12541 = n12540 ^ n12538 ^ 1'b0 ;
  assign n12542 = n9212 | n12541 ;
  assign n12543 = n6593 & ~n12542 ;
  assign n12544 = ~n546 & n984 ;
  assign n12545 = n9836 | n12544 ;
  assign n12546 = n12545 ^ n4098 ^ 1'b0 ;
  assign n12547 = n10610 ^ n7649 ^ 1'b0 ;
  assign n12548 = ~n3657 & n7836 ;
  assign n12549 = n3388 ^ n1744 ^ 1'b0 ;
  assign n12550 = ~n5036 & n6804 ;
  assign n12551 = n12550 ^ n514 ^ 1'b0 ;
  assign n12552 = n12551 ^ n6036 ^ 1'b0 ;
  assign n12553 = n12549 & n12552 ;
  assign n12554 = ~n4765 & n8126 ;
  assign n12555 = ~n61 & n12554 ;
  assign n12556 = n5022 & n5857 ;
  assign n12557 = n12556 ^ n2595 ^ 1'b0 ;
  assign n12558 = n12557 ^ n10314 ^ 1'b0 ;
  assign n12559 = n4318 | n12558 ;
  assign n12560 = n7287 ^ n5863 ^ 1'b0 ;
  assign n12561 = n8200 | n12560 ;
  assign n12562 = n10269 & ~n12561 ;
  assign n12563 = n1918 & ~n6560 ;
  assign n12564 = n914 & n12563 ;
  assign n12565 = ~n5507 & n12564 ;
  assign n12566 = n3235 & ~n5607 ;
  assign n12567 = n5214 ^ n19 ^ 1'b0 ;
  assign n12568 = ( n3238 & n12236 ) | ( n3238 & n12567 ) | ( n12236 & n12567 ) ;
  assign n12569 = ~n473 & n533 ;
  assign n12570 = ~n533 & n12569 ;
  assign n12571 = n4902 | n12570 ;
  assign n12572 = n12571 ^ n2395 ^ 1'b0 ;
  assign n12573 = ~n4914 & n10403 ;
  assign n12574 = n12573 ^ n1337 ^ 1'b0 ;
  assign n12575 = ~n1226 & n12574 ;
  assign n12576 = n9463 ^ n6656 ^ 1'b0 ;
  assign n12577 = n12576 ^ n2915 ^ 1'b0 ;
  assign n12578 = n2150 & n12577 ;
  assign n12579 = ~n266 & n12578 ;
  assign n12580 = ( n8200 & n12575 ) | ( n8200 & n12579 ) | ( n12575 & n12579 ) ;
  assign n12581 = n3034 ^ n2856 ^ 1'b0 ;
  assign n12582 = ~n4116 & n12581 ;
  assign n12583 = n4017 & n12582 ;
  assign n12584 = n5266 ^ n2996 ^ 1'b0 ;
  assign n12585 = n12584 ^ n2721 ^ 1'b0 ;
  assign n12586 = n3842 | n5901 ;
  assign n12587 = n5564 & ~n7737 ;
  assign n12588 = n12587 ^ n1994 ^ 1'b0 ;
  assign n12591 = n10786 ^ n10665 ^ 1'b0 ;
  assign n12589 = n2655 | n4942 ;
  assign n12590 = n8761 | n12589 ;
  assign n12592 = n12591 ^ n12590 ^ 1'b0 ;
  assign n12593 = n10257 ^ n582 ^ 1'b0 ;
  assign n12594 = n9002 ^ n8399 ^ 1'b0 ;
  assign n12595 = n6366 | n12594 ;
  assign n12596 = n3794 ^ n2754 ^ 1'b0 ;
  assign n12597 = n12596 ^ n183 ^ 1'b0 ;
  assign n12598 = n12597 ^ n5281 ^ 1'b0 ;
  assign n12599 = n1951 ^ n934 ^ 1'b0 ;
  assign n12600 = n10767 ^ n7635 ^ 1'b0 ;
  assign n12601 = n6463 | n12600 ;
  assign n12602 = n12599 | n12601 ;
  assign n12603 = n1138 | n2199 ;
  assign n12604 = n2346 & ~n12603 ;
  assign n12605 = n8029 ^ n362 ^ 1'b0 ;
  assign n12606 = n2624 & ~n12605 ;
  assign n12607 = n12606 ^ n2576 ^ 1'b0 ;
  assign n12608 = n244 | n12607 ;
  assign n12609 = n8512 | n12608 ;
  assign n12610 = n12604 | n12609 ;
  assign n12611 = n12610 ^ n9621 ^ 1'b0 ;
  assign n12612 = n8284 ^ n5812 ^ 1'b0 ;
  assign n12613 = n4735 ^ n1437 ^ 1'b0 ;
  assign n12614 = n1592 | n12613 ;
  assign n12615 = n1434 | n4324 ;
  assign n12616 = n12615 ^ n1353 ^ 1'b0 ;
  assign n12617 = n12616 ^ n9912 ^ 1'b0 ;
  assign n12618 = ( n4626 & ~n6360 ) | ( n4626 & n12617 ) | ( ~n6360 & n12617 ) ;
  assign n12619 = n4945 ^ n3019 ^ n1693 ;
  assign n12620 = n12618 | n12619 ;
  assign n12621 = n5026 | n12620 ;
  assign n12622 = n12621 ^ n11295 ^ n3145 ;
  assign n12623 = n9781 ^ n7142 ^ 1'b0 ;
  assign n12624 = ~n260 & n1660 ;
  assign n12625 = n12624 ^ n2246 ^ 1'b0 ;
  assign n12626 = n12625 ^ n9072 ^ 1'b0 ;
  assign n12627 = n5510 | n8273 ;
  assign n12628 = n7479 & ~n12627 ;
  assign n12629 = n12628 ^ n1738 ^ 1'b0 ;
  assign n12630 = ~n10170 & n12629 ;
  assign n12631 = n11664 ^ n6566 ^ 1'b0 ;
  assign n12632 = n8510 & n12631 ;
  assign n12633 = n2405 | n3042 ;
  assign n12634 = ~n4167 & n10003 ;
  assign n12635 = n1731 & ~n12634 ;
  assign n12636 = ~n2723 & n11176 ;
  assign n12637 = ~n3802 & n11088 ;
  assign n12638 = n12637 ^ n6037 ^ n1985 ;
  assign n12640 = n865 & n9016 ;
  assign n12641 = n8247 & n12640 ;
  assign n12639 = n434 & n7736 ;
  assign n12642 = n12641 ^ n12639 ^ 1'b0 ;
  assign n12643 = n5226 | n12642 ;
  assign n12644 = n6768 & n10439 ;
  assign n12645 = n4170 ^ n3924 ^ 1'b0 ;
  assign n12646 = ~n2811 & n12645 ;
  assign n12647 = n8030 ^ n1476 ^ 1'b0 ;
  assign n12648 = n9089 | n12647 ;
  assign n12649 = n12224 & ~n12648 ;
  assign n12650 = n10264 ^ n5332 ^ 1'b0 ;
  assign n12651 = n12130 | n12650 ;
  assign n12652 = n1747 | n2382 ;
  assign n12653 = ~n1639 & n2408 ;
  assign n12654 = n2881 | n3019 ;
  assign n12655 = n2044 & ~n7019 ;
  assign n12656 = n8486 | n12655 ;
  assign n12657 = n634 | n12656 ;
  assign n12658 = n12654 | n12657 ;
  assign n12659 = ~n774 & n4510 ;
  assign n12660 = ~n9461 & n12659 ;
  assign n12661 = n61 | n1434 ;
  assign n12662 = n441 & n12661 ;
  assign n12667 = n2943 | n7322 ;
  assign n12663 = n175 | n228 ;
  assign n12664 = n511 | n12663 ;
  assign n12665 = n9170 | n9685 ;
  assign n12666 = n12664 & n12665 ;
  assign n12668 = n12667 ^ n12666 ^ 1'b0 ;
  assign n12669 = n9038 & ~n12668 ;
  assign n12670 = n9111 ^ n1424 ^ 1'b0 ;
  assign n12671 = n11271 | n12670 ;
  assign n12672 = n1976 ^ n749 ^ 1'b0 ;
  assign n12673 = ~n2273 & n12672 ;
  assign n12674 = n12673 ^ n5345 ^ 1'b0 ;
  assign n12675 = n8630 | n12674 ;
  assign n12676 = n6575 ^ n2136 ^ 1'b0 ;
  assign n12677 = ~n5154 & n12676 ;
  assign n12678 = n5191 & ~n12677 ;
  assign n12679 = ~n2030 & n10229 ;
  assign n12680 = n3011 | n4139 ;
  assign n12681 = n51 & ~n10121 ;
  assign n12682 = n9163 ^ n6413 ^ 1'b0 ;
  assign n12683 = n2079 & n2610 ;
  assign n12684 = ~n5085 & n5432 ;
  assign n12685 = n12684 ^ n786 ^ 1'b0 ;
  assign n12686 = n12685 ^ n5981 ^ n543 ;
  assign n12687 = n6700 & ~n12686 ;
  assign n12688 = ( n1854 & n7008 ) | ( n1854 & ~n12687 ) | ( n7008 & ~n12687 ) ;
  assign n12689 = n12688 ^ n1208 ^ 1'b0 ;
  assign n12690 = n2558 & n4085 ;
  assign n12691 = n3338 | n6525 ;
  assign n12692 = n9535 | n12691 ;
  assign n12693 = n8563 & n12692 ;
  assign n12694 = ( n1055 & n12690 ) | ( n1055 & n12693 ) | ( n12690 & n12693 ) ;
  assign n12695 = n10254 & ~n11276 ;
  assign n12696 = n10110 ^ n2562 ^ 1'b0 ;
  assign n12697 = ~n12695 & n12696 ;
  assign n12698 = n8322 & n12697 ;
  assign n12699 = n5403 | n7916 ;
  assign n12700 = ~n4235 & n12699 ;
  assign n12701 = n1688 | n3314 ;
  assign n12702 = n1078 & n12701 ;
  assign n12703 = n8482 ^ n4015 ^ 1'b0 ;
  assign n12704 = n12703 ^ n7430 ^ 1'b0 ;
  assign n12705 = n940 & n12187 ;
  assign n12706 = n2394 | n5016 ;
  assign n12707 = n2394 & ~n12706 ;
  assign n12708 = n354 & ~n12707 ;
  assign n12709 = ~n354 & n12708 ;
  assign n12710 = n2580 & n12709 ;
  assign n12711 = n7189 & ~n12710 ;
  assign n12712 = n12710 & n12711 ;
  assign n12713 = n5824 & n12501 ;
  assign n12714 = ~n5001 & n6950 ;
  assign n12715 = ~n9190 & n12714 ;
  assign n12716 = n3272 | n12715 ;
  assign n12717 = ( n155 & ~n1063 ) | ( n155 & n6035 ) | ( ~n1063 & n6035 ) ;
  assign n12718 = n12717 ^ n2377 ^ 1'b0 ;
  assign n12719 = ( ~n3017 & n3680 ) | ( ~n3017 & n6278 ) | ( n3680 & n6278 ) ;
  assign n12720 = ~n1774 & n12719 ;
  assign n12721 = ~n12718 & n12720 ;
  assign n12722 = ~n1514 & n11902 ;
  assign n12723 = n12721 & n12722 ;
  assign n12725 = n1949 | n2683 ;
  assign n12724 = n2929 | n7771 ;
  assign n12726 = n12725 ^ n12724 ^ 1'b0 ;
  assign n12727 = ~n9432 & n12726 ;
  assign n12728 = n3272 ^ n38 ^ 1'b0 ;
  assign n12729 = n7569 & ~n12728 ;
  assign n12730 = n5237 & n12729 ;
  assign n12731 = ~n4085 & n12730 ;
  assign n12732 = ~n1114 & n2724 ;
  assign n12733 = ( n7645 & n9589 ) | ( n7645 & n12732 ) | ( n9589 & n12732 ) ;
  assign n12734 = n4726 ^ n1240 ^ 1'b0 ;
  assign n12735 = ~n189 & n12734 ;
  assign n12736 = n5760 ^ n5412 ^ 1'b0 ;
  assign n12737 = n12736 ^ n3502 ^ 1'b0 ;
  assign n12738 = ~n7075 & n12737 ;
  assign n12739 = ~n899 & n6568 ;
  assign n12740 = n11469 & n12739 ;
  assign n12741 = n12056 & ~n12740 ;
  assign n12742 = n3187 & n12741 ;
  assign n12743 = n1747 & n2324 ;
  assign n12744 = n12743 ^ n3951 ^ 1'b0 ;
  assign n12745 = n6757 & ~n12450 ;
  assign n12746 = ~n12744 & n12745 ;
  assign n12747 = ( n910 & n4609 ) | ( n910 & ~n7660 ) | ( n4609 & ~n7660 ) ;
  assign n12752 = n4607 ^ n4403 ^ 1'b0 ;
  assign n12753 = n10299 & n12752 ;
  assign n12754 = ~n3962 & n12753 ;
  assign n12749 = n301 & ~n473 ;
  assign n12750 = n2619 & n12749 ;
  assign n12748 = n5890 | n12076 ;
  assign n12751 = n12750 ^ n12748 ^ 1'b0 ;
  assign n12755 = n12754 ^ n12751 ^ 1'b0 ;
  assign n12756 = n12673 ^ n3019 ^ 1'b0 ;
  assign n12757 = ~n8949 & n12756 ;
  assign n12758 = n12757 ^ n3377 ^ 1'b0 ;
  assign n12759 = n2904 ^ n896 ^ 1'b0 ;
  assign n12760 = n12759 ^ n5426 ^ 1'b0 ;
  assign n12761 = ~n5447 & n12760 ;
  assign n12762 = n12052 & n12761 ;
  assign n12763 = n6817 ^ n296 ^ 1'b0 ;
  assign n12764 = n10251 & ~n12763 ;
  assign n12765 = n5393 & ~n8062 ;
  assign n12766 = n2233 & n12765 ;
  assign n12767 = ( ~n9832 & n12764 ) | ( ~n9832 & n12766 ) | ( n12764 & n12766 ) ;
  assign n12768 = n1032 & n4313 ;
  assign n12769 = n12768 ^ n7133 ^ 1'b0 ;
  assign n12770 = ~n9745 & n12769 ;
  assign n12774 = n3424 & n3794 ;
  assign n12775 = ~n3891 & n12774 ;
  assign n12772 = n3942 | n4053 ;
  assign n12773 = n12772 ^ n378 ^ 1'b0 ;
  assign n12776 = n12775 ^ n12773 ^ 1'b0 ;
  assign n12771 = n2996 ^ n1353 ^ n401 ;
  assign n12777 = n12776 ^ n12771 ^ 1'b0 ;
  assign n12778 = ~n4956 & n10016 ;
  assign n12779 = n12778 ^ n12617 ^ 1'b0 ;
  assign n12780 = n874 & n6836 ;
  assign n12781 = n6869 & ~n12780 ;
  assign n12782 = n5949 | n6832 ;
  assign n12783 = ~n112 & n5844 ;
  assign n12784 = n2517 & n12783 ;
  assign n12785 = n5269 ^ n1271 ^ 1'b0 ;
  assign n12786 = n11678 & n12785 ;
  assign n12787 = n9288 & n12786 ;
  assign n12788 = n12787 ^ n6269 ^ 1'b0 ;
  assign n12789 = n4768 ^ n2869 ^ 1'b0 ;
  assign n12790 = n2567 & ~n12789 ;
  assign n12791 = n1395 & ~n6108 ;
  assign n12792 = n3371 ^ n995 ^ 1'b0 ;
  assign n12793 = n5513 & n12792 ;
  assign n12794 = n8913 & ~n12793 ;
  assign n12795 = n9915 ^ n452 ^ 1'b0 ;
  assign n12796 = ~n2413 & n12795 ;
  assign n12798 = n2860 | n3724 ;
  assign n12799 = n2435 & ~n12798 ;
  assign n12797 = n1652 & ~n9311 ;
  assign n12800 = n12799 ^ n12797 ^ 1'b0 ;
  assign n12801 = n6621 ^ n183 ^ 1'b0 ;
  assign n12802 = n12801 ^ n181 ^ 1'b0 ;
  assign n12803 = n3530 ^ n2014 ^ n564 ;
  assign n12804 = n12285 & n12803 ;
  assign n12805 = n9690 ^ n8487 ^ 1'b0 ;
  assign n12806 = n5493 ^ n4238 ^ 1'b0 ;
  assign n12807 = n4890 & ~n12806 ;
  assign n12808 = n12807 ^ n8599 ^ n6831 ;
  assign n12809 = ~n4884 & n12808 ;
  assign n12811 = n1740 & n6496 ;
  assign n12812 = n4289 & n12811 ;
  assign n12813 = n12812 ^ n7707 ^ n2195 ;
  assign n12810 = ~n3081 & n10616 ;
  assign n12814 = n12813 ^ n12810 ^ 1'b0 ;
  assign n12815 = ~n1398 & n9095 ;
  assign n12816 = ( n1252 & n4762 ) | ( n1252 & n9877 ) | ( n4762 & n9877 ) ;
  assign n12817 = n667 & ~n726 ;
  assign n12818 = n12817 ^ n4338 ^ 1'b0 ;
  assign n12819 = n4819 | n12818 ;
  assign n12820 = n5903 ^ n4446 ^ 1'b0 ;
  assign n12821 = n1918 & ~n12820 ;
  assign n12822 = ~n12819 & n12821 ;
  assign n12823 = n12822 ^ n1414 ^ 1'b0 ;
  assign n12824 = n5973 ^ n88 ^ 1'b0 ;
  assign n12825 = n12824 ^ n9447 ^ 1'b0 ;
  assign n12826 = n10544 ^ n3776 ^ 1'b0 ;
  assign n12827 = n8992 ^ n443 ^ 1'b0 ;
  assign n12828 = n11949 & ~n12827 ;
  assign n12829 = n12828 ^ n4125 ^ 1'b0 ;
  assign n12830 = n12829 ^ n3576 ^ 1'b0 ;
  assign n12831 = n1771 | n2807 ;
  assign n12832 = n12022 ^ n2719 ^ 1'b0 ;
  assign n12833 = n12831 & ~n12832 ;
  assign n12834 = ~n7289 & n8959 ;
  assign n12835 = n12834 ^ n6749 ^ 1'b0 ;
  assign n12836 = n4679 ^ n2202 ^ 1'b0 ;
  assign n12837 = ~n1744 & n6411 ;
  assign n12838 = ~n5084 & n11890 ;
  assign n12839 = n12838 ^ n3488 ^ 1'b0 ;
  assign n12840 = n4158 ^ n2808 ^ n1291 ;
  assign n12841 = n1318 & n12840 ;
  assign n12842 = n8827 & n12841 ;
  assign n12843 = n12842 ^ n8549 ^ 1'b0 ;
  assign n12844 = n12843 ^ n2317 ^ 1'b0 ;
  assign n12845 = n12839 & n12844 ;
  assign n12846 = n10782 & n12845 ;
  assign n12847 = n6383 & n12846 ;
  assign n12848 = n6203 ^ n5195 ^ 1'b0 ;
  assign n12849 = n8660 | n12848 ;
  assign n12850 = n12849 ^ n1293 ^ 1'b0 ;
  assign n12851 = n6102 & n12850 ;
  assign n12852 = n12851 ^ n8604 ^ 1'b0 ;
  assign n12853 = n5872 & ~n12852 ;
  assign n12854 = n5511 & n7298 ;
  assign n12855 = n3289 & ~n5145 ;
  assign n12856 = ~n12854 & n12855 ;
  assign n12857 = n12856 ^ n5324 ^ 1'b0 ;
  assign n12858 = n1703 | n12857 ;
  assign n12859 = n466 & n11124 ;
  assign n12860 = n4732 & n12859 ;
  assign n12861 = n2576 | n12860 ;
  assign n12862 = n1686 & ~n12861 ;
  assign n12863 = n12007 ^ n852 ^ 1'b0 ;
  assign n12864 = n12862 | n12863 ;
  assign n12865 = n885 | n12864 ;
  assign n12866 = ~n7655 & n12865 ;
  assign n12867 = ~n4787 & n12866 ;
  assign n12868 = n2605 ^ n1893 ^ 1'b0 ;
  assign n12869 = n12868 ^ n9159 ^ 1'b0 ;
  assign n12870 = ~n2680 & n12869 ;
  assign n12871 = n12634 & ~n12870 ;
  assign n12872 = n25 & ~n7030 ;
  assign n12873 = n1778 & n12872 ;
  assign n12874 = n10012 ^ n991 ^ 1'b0 ;
  assign n12875 = n4285 | n12874 ;
  assign n12876 = ~n257 & n7881 ;
  assign n12877 = n6408 & n12876 ;
  assign n12878 = n7131 | n12877 ;
  assign n12879 = ~n806 & n1895 ;
  assign n12880 = ~n140 & n788 ;
  assign n12881 = n12880 ^ n7562 ^ 1'b0 ;
  assign n12882 = n957 & n12881 ;
  assign n12883 = n10537 & n12882 ;
  assign n12884 = n5491 ^ n5099 ^ 1'b0 ;
  assign n12885 = n3657 | n12884 ;
  assign n12886 = n5076 & n9771 ;
  assign n12887 = ~n11428 & n12886 ;
  assign n12888 = n8144 & ~n12887 ;
  assign n12889 = n10320 & n12888 ;
  assign n12890 = n3165 ^ n3063 ^ 1'b0 ;
  assign n12891 = ( ~n2148 & n6771 ) | ( ~n2148 & n10349 ) | ( n6771 & n10349 ) ;
  assign n12892 = n12891 ^ n8553 ^ 1'b0 ;
  assign n12893 = ~n12890 & n12892 ;
  assign n12894 = n423 & n1991 ;
  assign n12895 = ~n125 & n5779 ;
  assign n12896 = ( ~n5348 & n12894 ) | ( ~n5348 & n12895 ) | ( n12894 & n12895 ) ;
  assign n12897 = n3212 & ~n9863 ;
  assign n12898 = n3049 ^ n1464 ^ 1'b0 ;
  assign n12899 = n342 & n12898 ;
  assign n12900 = ~n5126 & n8996 ;
  assign n12901 = n12900 ^ n2967 ^ 1'b0 ;
  assign n12902 = n12899 & n12901 ;
  assign n12903 = n12902 ^ n8189 ^ 1'b0 ;
  assign n12904 = n2895 ^ n167 ^ 1'b0 ;
  assign n12905 = n7515 | n12904 ;
  assign n12906 = n12905 ^ n7766 ^ 1'b0 ;
  assign n12907 = n3637 ^ n2806 ^ 1'b0 ;
  assign n12908 = n9346 & ~n12907 ;
  assign n12909 = n12908 ^ n10144 ^ 1'b0 ;
  assign n12910 = n12909 ^ n2760 ^ 1'b0 ;
  assign n12911 = n12906 | n12910 ;
  assign n12912 = ~n1055 & n2686 ;
  assign n12913 = n12912 ^ n368 ^ 1'b0 ;
  assign n12914 = n7590 & ~n9629 ;
  assign n12915 = ( n352 & ~n545 ) | ( n352 & n984 ) | ( ~n545 & n984 ) ;
  assign n12916 = n2708 | n12915 ;
  assign n12917 = n10290 ^ n7245 ^ 1'b0 ;
  assign n12918 = n4553 & n9717 ;
  assign n12919 = n3214 & n12918 ;
  assign n12920 = n12919 ^ n2884 ^ 1'b0 ;
  assign n12921 = n7500 & n10723 ;
  assign n12922 = n3760 & n8236 ;
  assign n12923 = n8757 | n12922 ;
  assign n12924 = n12923 ^ n3619 ^ 1'b0 ;
  assign n12925 = ( n12603 & n12921 ) | ( n12603 & n12924 ) | ( n12921 & n12924 ) ;
  assign n12926 = n2335 & ~n3809 ;
  assign n12927 = n1686 & n12926 ;
  assign n12928 = n9140 | n12927 ;
  assign n12929 = n12928 ^ n2199 ^ 1'b0 ;
  assign n12930 = n6247 ^ n1536 ^ 1'b0 ;
  assign n12931 = ~n8312 & n11107 ;
  assign n12932 = n1769 ^ n808 ^ 1'b0 ;
  assign n12933 = n3088 ^ n2207 ^ 1'b0 ;
  assign n12934 = n1723 & n12933 ;
  assign n12935 = n12934 ^ n3591 ^ n1558 ;
  assign n12936 = n3735 & ~n12935 ;
  assign n12937 = ~n12932 & n12936 ;
  assign n12938 = n11572 ^ n3033 ^ 1'b0 ;
  assign n12939 = n8241 ^ n1522 ^ 1'b0 ;
  assign n12940 = n11927 ^ n1726 ^ 1'b0 ;
  assign n12941 = n9186 | n12940 ;
  assign n12942 = n3353 & n12941 ;
  assign n12943 = n2802 & n10311 ;
  assign n12944 = n2771 | n12943 ;
  assign n12945 = ( n3476 & n6839 ) | ( n3476 & ~n11923 ) | ( n6839 & ~n11923 ) ;
  assign n12946 = n10911 ^ n9745 ^ 1'b0 ;
  assign n12947 = n1441 | n12946 ;
  assign n12948 = n9220 ^ n3449 ^ 1'b0 ;
  assign n12949 = n586 | n12948 ;
  assign n12950 = ~n3995 & n9540 ;
  assign n12951 = n10611 & ~n12950 ;
  assign n12952 = n12951 ^ n10611 ^ n171 ;
  assign n12953 = ~n3060 & n8023 ;
  assign n12954 = ~n8023 & n12953 ;
  assign n12955 = n995 | n12954 ;
  assign n12956 = n995 & ~n12955 ;
  assign n12957 = n10166 & ~n12956 ;
  assign n12960 = n144 | n4595 ;
  assign n12961 = n4595 & ~n12960 ;
  assign n12962 = n9650 & n12961 ;
  assign n12958 = n1779 | n4135 ;
  assign n12959 = n1779 & ~n12958 ;
  assign n12963 = n12962 ^ n12959 ^ 1'b0 ;
  assign n12964 = n12957 & ~n12963 ;
  assign n12965 = n253 & ~n1709 ;
  assign n12966 = n1620 | n12965 ;
  assign n12967 = n3331 ^ n1920 ^ 1'b0 ;
  assign n12968 = ~n948 & n7293 ;
  assign n12969 = n577 & n9094 ;
  assign n12970 = n5841 | n12432 ;
  assign n12971 = n8819 ^ n6969 ^ 1'b0 ;
  assign n12972 = n6378 & n12971 ;
  assign n12973 = n212 | n10684 ;
  assign n12974 = n12973 ^ n8058 ^ 1'b0 ;
  assign n12975 = ~n3598 & n9892 ;
  assign n12976 = n12975 ^ n2363 ^ 1'b0 ;
  assign n12977 = n12976 ^ n5360 ^ 1'b0 ;
  assign n12978 = n7997 & n9944 ;
  assign n12979 = ~n3565 & n12978 ;
  assign n12980 = n12979 ^ n10603 ^ 1'b0 ;
  assign n12981 = n4166 & n9579 ;
  assign n12982 = n5118 & ~n12981 ;
  assign n12983 = n7659 & n12982 ;
  assign n12984 = ( n7597 & n12980 ) | ( n7597 & ~n12983 ) | ( n12980 & ~n12983 ) ;
  assign n12985 = n3691 & n3944 ;
  assign n12986 = ~n3783 & n12985 ;
  assign n12987 = ( n10786 & n11363 ) | ( n10786 & ~n12152 ) | ( n11363 & ~n12152 ) ;
  assign n12989 = n6680 ^ n5332 ^ 1'b0 ;
  assign n12988 = n5412 ^ n4117 ^ 1'b0 ;
  assign n12990 = n12989 ^ n12988 ^ n8152 ;
  assign n12991 = ~n12693 & n12990 ;
  assign n12996 = n4510 & ~n5403 ;
  assign n12992 = n4422 | n4485 ;
  assign n12993 = n12992 ^ n518 ^ 1'b0 ;
  assign n12994 = n12993 ^ n3972 ^ 1'b0 ;
  assign n12995 = n12994 ^ n5284 ^ 1'b0 ;
  assign n12997 = n12996 ^ n12995 ^ 1'b0 ;
  assign n12998 = n459 & ~n12997 ;
  assign n12999 = n7734 ^ n7033 ^ 1'b0 ;
  assign n13000 = n12998 & ~n12999 ;
  assign n13007 = n4546 ^ n302 ^ 1'b0 ;
  assign n13001 = n4098 & n8820 ;
  assign n13002 = n13001 ^ n4990 ^ 1'b0 ;
  assign n13003 = n598 & n9219 ;
  assign n13004 = ~n13002 & n13003 ;
  assign n13005 = n12128 | n13004 ;
  assign n13006 = n13005 ^ n10270 ^ 1'b0 ;
  assign n13008 = n13007 ^ n13006 ^ n1726 ;
  assign n13009 = n3501 | n6697 ;
  assign n13010 = n13009 ^ n6542 ^ 1'b0 ;
  assign n13011 = n3422 & ~n3571 ;
  assign n13012 = ~n10913 & n13011 ;
  assign n13013 = n13012 ^ n2132 ^ 1'b0 ;
  assign n13014 = n2899 & n9353 ;
  assign n13015 = n4551 & n13014 ;
  assign n13016 = n11064 ^ n6457 ^ 1'b0 ;
  assign n13017 = ~n5419 & n13016 ;
  assign n13018 = n3823 ^ n2953 ^ 1'b0 ;
  assign n13019 = n10820 ^ n10298 ^ 1'b0 ;
  assign n13020 = n782 & ~n3301 ;
  assign n13021 = n4162 & n13020 ;
  assign n13022 = n13021 ^ n7523 ^ 1'b0 ;
  assign n13023 = n171 & ~n13022 ;
  assign n13024 = n5557 & n9026 ;
  assign n13025 = n1293 | n13024 ;
  assign n13026 = n13025 ^ n5399 ^ 1'b0 ;
  assign n13027 = n13026 ^ n3696 ^ 1'b0 ;
  assign n13028 = n6389 & ~n13027 ;
  assign n13029 = n13028 ^ n11694 ^ 1'b0 ;
  assign n13030 = n7482 | n13029 ;
  assign n13031 = n9049 ^ n4463 ^ 1'b0 ;
  assign n13032 = n219 & ~n5110 ;
  assign n13033 = ~n13031 & n13032 ;
  assign n13034 = n9641 & n13033 ;
  assign n13035 = n13034 ^ n4007 ^ 1'b0 ;
  assign n13036 = n4264 & ~n4679 ;
  assign n13037 = n12587 ^ n10118 ^ 1'b0 ;
  assign n13038 = n5936 ^ n1208 ^ 1'b0 ;
  assign n13039 = n11006 & ~n13038 ;
  assign n13040 = n3432 | n13039 ;
  assign n13041 = n13037 & n13040 ;
  assign n13042 = n11016 ^ n6719 ^ 1'b0 ;
  assign n13043 = n3902 | n13042 ;
  assign n13044 = n8693 | n13043 ;
  assign n13045 = n4183 ^ n1893 ^ 1'b0 ;
  assign n13046 = n13044 & n13045 ;
  assign n13047 = n219 | n2812 ;
  assign n13048 = n13047 ^ n1976 ^ 1'b0 ;
  assign n13049 = n5123 ^ n2384 ^ 1'b0 ;
  assign n13050 = n86 & n13049 ;
  assign n13051 = n2885 & ~n10383 ;
  assign n13052 = ~n13050 & n13051 ;
  assign n13053 = ~n13048 & n13052 ;
  assign n13058 = n1720 | n7546 ;
  assign n13059 = n13058 ^ n5903 ^ 1'b0 ;
  assign n13055 = n2560 & ~n4899 ;
  assign n13054 = n3568 & n3897 ;
  assign n13056 = n13055 ^ n13054 ^ 1'b0 ;
  assign n13057 = ~n6557 & n13056 ;
  assign n13060 = n13059 ^ n13057 ^ 1'b0 ;
  assign n13061 = ~n3839 & n4170 ;
  assign n13062 = n8319 ^ n3539 ^ 1'b0 ;
  assign n13063 = ~n2238 & n11402 ;
  assign n13064 = n8332 & n10083 ;
  assign n13065 = ~n12188 & n13064 ;
  assign n13066 = n179 | n13065 ;
  assign n13067 = n4027 ^ n1693 ^ 1'b0 ;
  assign n13068 = n3090 & ~n13067 ;
  assign n13069 = n13068 ^ n6350 ^ 1'b0 ;
  assign n13070 = n7720 & ~n13061 ;
  assign n13071 = ( n7091 & ~n9534 ) | ( n7091 & n13070 ) | ( ~n9534 & n13070 ) ;
  assign n13072 = n13069 & n13071 ;
  assign n13073 = n13072 ^ n3921 ^ 1'b0 ;
  assign n13074 = ~n320 & n8332 ;
  assign n13075 = n13074 ^ n995 ^ 1'b0 ;
  assign n13076 = n5801 ^ n3351 ^ 1'b0 ;
  assign n13077 = n10024 | n13076 ;
  assign n13078 = n8416 ^ n3361 ^ 1'b0 ;
  assign n13079 = n7864 & ~n13078 ;
  assign n13080 = n1802 | n6817 ;
  assign n13081 = n12582 ^ n3504 ^ 1'b0 ;
  assign n13082 = n11187 ^ n9094 ^ 1'b0 ;
  assign n13083 = n1205 ^ n717 ^ 1'b0 ;
  assign n13084 = n13083 ^ n10556 ^ 1'b0 ;
  assign n13085 = n5618 | n13084 ;
  assign n13086 = n3987 & ~n13085 ;
  assign n13087 = n2641 ^ n1035 ^ 1'b0 ;
  assign n13088 = n6527 & n13087 ;
  assign n13089 = ~n2758 & n13088 ;
  assign n13090 = n2914 & n4675 ;
  assign n13091 = n13090 ^ n6729 ^ 1'b0 ;
  assign n13092 = n159 & ~n13091 ;
  assign n13093 = n5695 ^ n873 ^ 1'b0 ;
  assign n13094 = ~n8989 & n13093 ;
  assign n13095 = n4973 & ~n9684 ;
  assign n13096 = n5497 | n11782 ;
  assign n13100 = n2700 | n11074 ;
  assign n13101 = n754 & ~n13100 ;
  assign n13097 = n1181 & ~n6878 ;
  assign n13098 = n6633 ^ n3942 ^ 1'b0 ;
  assign n13099 = n13097 & n13098 ;
  assign n13102 = n13101 ^ n13099 ^ 1'b0 ;
  assign n13103 = n6607 ^ n4133 ^ 1'b0 ;
  assign n13104 = ~n5450 & n7574 ;
  assign n13106 = n5039 ^ n3891 ^ 1'b0 ;
  assign n13105 = n11292 ^ n1956 ^ 1'b0 ;
  assign n13107 = n13106 ^ n13105 ^ 1'b0 ;
  assign n13108 = ~n13104 & n13107 ;
  assign n13109 = n10913 & ~n13108 ;
  assign n13110 = n13109 ^ n9505 ^ 1'b0 ;
  assign n13111 = ~n253 & n1169 ;
  assign n13112 = ( ~n1843 & n5508 ) | ( ~n1843 & n13111 ) | ( n5508 & n13111 ) ;
  assign n13113 = n5182 ^ n2282 ^ 1'b0 ;
  assign n13114 = n354 & n13113 ;
  assign n13115 = n6206 | n8147 ;
  assign n13116 = n509 & ~n11618 ;
  assign n13117 = n777 & n13116 ;
  assign n13119 = n796 | n11225 ;
  assign n13118 = n4774 & ~n5168 ;
  assign n13120 = n13119 ^ n13118 ^ n3001 ;
  assign n13121 = ~n4917 & n5375 ;
  assign n13122 = n13121 ^ n5254 ^ 1'b0 ;
  assign n13123 = n13122 ^ n10903 ^ n6343 ;
  assign n13124 = ( n1536 & ~n2504 ) | ( n1536 & n4718 ) | ( ~n2504 & n4718 ) ;
  assign n13125 = n11497 | n13124 ;
  assign n13126 = n3992 | n11861 ;
  assign n13127 = n10330 ^ n4709 ^ 1'b0 ;
  assign n13128 = n2403 & n13127 ;
  assign n13129 = n13128 ^ n420 ^ 1'b0 ;
  assign n13130 = n1385 & ~n4499 ;
  assign n13131 = n13130 ^ n8936 ^ n3224 ;
  assign n13132 = n6330 & ~n8259 ;
  assign n13133 = n13132 ^ n4913 ^ 1'b0 ;
  assign n13134 = ( n982 & ~n1205 ) | ( n982 & n5595 ) | ( ~n1205 & n5595 ) ;
  assign n13135 = ~n1657 & n1920 ;
  assign n13136 = ~n13134 & n13135 ;
  assign n13137 = n10933 & ~n13136 ;
  assign n13138 = n5219 ^ n886 ^ 1'b0 ;
  assign n13139 = ~n778 & n9060 ;
  assign n13140 = n13139 ^ n2883 ^ 1'b0 ;
  assign n13141 = n3488 & ~n10441 ;
  assign n13142 = n13141 ^ n5480 ^ 1'b0 ;
  assign n13143 = n9908 | n13142 ;
  assign n13144 = n568 & ~n7632 ;
  assign n13145 = n7077 ^ n3334 ^ 1'b0 ;
  assign n13146 = n6989 | n13145 ;
  assign n13149 = n2914 & n3827 ;
  assign n13150 = n13149 ^ n3591 ^ 1'b0 ;
  assign n13151 = n4010 | n4290 ;
  assign n13152 = n280 | n13151 ;
  assign n13153 = n13152 ^ n9646 ^ 1'b0 ;
  assign n13154 = n13150 | n13153 ;
  assign n13155 = n2314 ^ n528 ^ 1'b0 ;
  assign n13156 = n782 & n1900 ;
  assign n13157 = n13156 ^ n3270 ^ 1'b0 ;
  assign n13158 = n1495 & ~n13157 ;
  assign n13159 = ~n13155 & n13158 ;
  assign n13160 = n8948 & ~n13159 ;
  assign n13161 = n3710 & n13160 ;
  assign n13162 = n2340 | n13161 ;
  assign n13163 = n13162 ^ n7611 ^ 1'b0 ;
  assign n13164 = n13154 & n13163 ;
  assign n13147 = ~n1033 & n2588 ;
  assign n13148 = n8521 & ~n13147 ;
  assign n13165 = n13164 ^ n13148 ^ 1'b0 ;
  assign n13166 = n5328 ^ n880 ^ 1'b0 ;
  assign n13167 = n1830 | n13166 ;
  assign n13168 = n7160 ^ n144 ^ 1'b0 ;
  assign n13169 = ~n1538 & n6095 ;
  assign n13170 = ~n2767 & n13169 ;
  assign n13171 = n13170 ^ n1269 ^ 1'b0 ;
  assign n13172 = n688 | n4585 ;
  assign n13173 = n440 & n6926 ;
  assign n13175 = n541 & ~n1144 ;
  assign n13174 = n11637 ^ n1416 ^ 1'b0 ;
  assign n13176 = n13175 ^ n13174 ^ 1'b0 ;
  assign n13177 = n10911 ^ n4926 ^ 1'b0 ;
  assign n13178 = n7170 & n8403 ;
  assign n13179 = n5119 & n13178 ;
  assign n13180 = ~n7699 & n7765 ;
  assign n13181 = n1382 & ~n13180 ;
  assign n13182 = n4772 & ~n4942 ;
  assign n13183 = n1511 & n4757 ;
  assign n13184 = ( n478 & n1715 ) | ( n478 & n13183 ) | ( n1715 & n13183 ) ;
  assign n13185 = ~n5027 & n5049 ;
  assign n13186 = ~n191 & n1379 ;
  assign n13187 = n10703 & n13186 ;
  assign n13188 = n13187 ^ n4389 ^ 1'b0 ;
  assign n13189 = n8578 ^ n5188 ^ 1'b0 ;
  assign n13190 = n4511 & ~n13189 ;
  assign n13191 = n7647 & n13190 ;
  assign n13192 = n13191 ^ n2564 ^ 1'b0 ;
  assign n13193 = n1499 & n1528 ;
  assign n13194 = n13193 ^ n5501 ^ 1'b0 ;
  assign n13195 = n376 & n2941 ;
  assign n13196 = ~n2784 & n13195 ;
  assign n13197 = n13196 ^ n61 ^ 1'b0 ;
  assign n13198 = n3402 & n13197 ;
  assign n13199 = ~n2022 & n2085 ;
  assign n13200 = n2681 & n13199 ;
  assign n13201 = ~n942 & n13200 ;
  assign n13202 = n13198 | n13201 ;
  assign n13203 = ~n4088 & n9264 ;
  assign n13204 = n5997 & ~n12178 ;
  assign n13205 = n263 & n4712 ;
  assign n13206 = n13205 ^ n4858 ^ 1'b0 ;
  assign n13207 = n5458 | n13206 ;
  assign n13208 = n3995 ^ n2796 ^ 1'b0 ;
  assign n13209 = n9288 & n10376 ;
  assign n13210 = n13209 ^ n7007 ^ 1'b0 ;
  assign n13211 = n11041 ^ n10864 ^ 1'b0 ;
  assign n13212 = n12998 & n13211 ;
  assign n13213 = n13212 ^ n423 ^ 1'b0 ;
  assign n13214 = n13213 ^ n7696 ^ n2695 ;
  assign n13215 = n9336 ^ n6976 ^ 1'b0 ;
  assign n13216 = n13214 & n13215 ;
  assign n13217 = n11118 ^ n3114 ^ 1'b0 ;
  assign n13218 = ~n870 & n13217 ;
  assign n13219 = n758 | n11292 ;
  assign n13220 = ~n5717 & n13219 ;
  assign n13221 = n13220 ^ n10114 ^ 1'b0 ;
  assign n13222 = ~n9047 & n11477 ;
  assign n13223 = n13221 & n13222 ;
  assign n13224 = ~n12383 & n13223 ;
  assign n13228 = n119 | n4077 ;
  assign n13229 = n13228 ^ n112 ^ 1'b0 ;
  assign n13225 = n9536 ^ n6056 ^ 1'b0 ;
  assign n13226 = n8134 ^ n5296 ^ 1'b0 ;
  assign n13227 = n13225 | n13226 ;
  assign n13230 = n13229 ^ n13227 ^ 1'b0 ;
  assign n13231 = n10728 ^ n5390 ^ 1'b0 ;
  assign n13232 = ~n371 & n8537 ;
  assign n13233 = n13232 ^ n9493 ^ 1'b0 ;
  assign n13234 = n13233 ^ n3044 ^ 1'b0 ;
  assign n13235 = n699 & ~n805 ;
  assign n13236 = n7382 & n13235 ;
  assign n13237 = ( ~n362 & n2562 ) | ( ~n362 & n8838 ) | ( n2562 & n8838 ) ;
  assign n13238 = n5482 ^ n1729 ^ 1'b0 ;
  assign n13239 = n7297 & ~n13238 ;
  assign n13240 = n11058 & n13239 ;
  assign n13241 = n13240 ^ n839 ^ 1'b0 ;
  assign n13242 = ~n2019 & n13241 ;
  assign n13243 = n3044 & n10567 ;
  assign n13244 = n10209 ^ n1337 ^ 1'b0 ;
  assign n13245 = ~n13243 & n13244 ;
  assign n13246 = n8970 & n13245 ;
  assign n13247 = n8293 ^ n4506 ^ n3802 ;
  assign n13248 = n2565 & ~n9204 ;
  assign n13249 = ~n200 & n6924 ;
  assign n13251 = ~n1650 & n2394 ;
  assign n13250 = n1670 & ~n7621 ;
  assign n13252 = n13251 ^ n13250 ^ 1'b0 ;
  assign n13253 = n13252 ^ n12637 ^ 1'b0 ;
  assign n13254 = n903 & ~n13253 ;
  assign n13255 = n11831 ^ n7125 ^ 1'b0 ;
  assign n13256 = n6172 ^ n3035 ^ 1'b0 ;
  assign n13257 = ~n327 & n3574 ;
  assign n13258 = n6766 ^ n2533 ^ 1'b0 ;
  assign n13259 = n7705 & n13258 ;
  assign n13260 = n226 & ~n9317 ;
  assign n13261 = n13260 ^ n11909 ^ 1'b0 ;
  assign n13262 = ( n2680 & ~n5368 ) | ( n2680 & n5446 ) | ( ~n5368 & n5446 ) ;
  assign n13263 = n4505 & n10232 ;
  assign n13264 = n4302 & ~n5179 ;
  assign n13265 = n13264 ^ n3399 ^ 1'b0 ;
  assign n13266 = n9546 & ~n13265 ;
  assign n13267 = ~n8758 & n12103 ;
  assign n13268 = n13267 ^ n10231 ^ 1'b0 ;
  assign n13269 = n13266 & ~n13268 ;
  assign n13270 = ~n1083 & n2669 ;
  assign n13271 = n4419 & ~n9202 ;
  assign n13272 = n13271 ^ n10944 ^ 1'b0 ;
  assign n13273 = n9106 & ~n10900 ;
  assign n13274 = n13272 & ~n13273 ;
  assign n13275 = n2494 | n12336 ;
  assign n13276 = ~n12968 & n13275 ;
  assign n13277 = n7520 & n13276 ;
  assign n13278 = n31 | n6794 ;
  assign n13279 = n9682 | n13278 ;
  assign n13280 = ~n9779 & n13279 ;
  assign n13281 = n13280 ^ n11386 ^ 1'b0 ;
  assign n13282 = n9305 & ~n13281 ;
  assign n13283 = n4793 & n13282 ;
  assign n13284 = n11151 & ~n13283 ;
  assign n13285 = n13284 ^ n7598 ^ 1'b0 ;
  assign n13286 = n2336 & n10404 ;
  assign n13287 = n2022 & n13286 ;
  assign n13288 = n13287 ^ n5106 ^ n2749 ;
  assign n13289 = n13288 ^ n10093 ^ 1'b0 ;
  assign n13290 = n736 & ~n13289 ;
  assign n13291 = n5151 & ~n7285 ;
  assign n13292 = ~n13290 & n13291 ;
  assign n13293 = n13189 ^ n9031 ^ 1'b0 ;
  assign n13294 = n13293 ^ n6675 ^ 1'b0 ;
  assign n13295 = n1853 & ~n13294 ;
  assign n13296 = n8103 ^ n910 ^ 1'b0 ;
  assign n13297 = n7628 ^ n2520 ^ 1'b0 ;
  assign n13298 = ~n2791 & n13297 ;
  assign n13299 = ( n1576 & n5474 ) | ( n1576 & ~n12492 ) | ( n5474 & ~n12492 ) ;
  assign n13300 = n7660 | n13299 ;
  assign n13301 = n12901 | n13300 ;
  assign n13302 = n13298 & n13301 ;
  assign n13303 = n1014 | n9858 ;
  assign n13304 = ~n3740 & n7067 ;
  assign n13305 = n13304 ^ n13018 ^ 1'b0 ;
  assign n13306 = n5241 | n13305 ;
  assign n13307 = n9733 & ~n11951 ;
  assign n13308 = n13307 ^ n6797 ^ 1'b0 ;
  assign n13309 = n7767 ^ n2741 ^ n1834 ;
  assign n13310 = ~n8906 & n13309 ;
  assign n13311 = n13310 ^ n7050 ^ 1'b0 ;
  assign n13312 = n1731 & ~n1922 ;
  assign n13313 = ~n13311 & n13312 ;
  assign n13314 = n13313 ^ n11218 ^ 1'b0 ;
  assign n13315 = n2618 & n3418 ;
  assign n13316 = n3482 & n3881 ;
  assign n13317 = n13315 & n13316 ;
  assign n13318 = n1469 & ~n10466 ;
  assign n13319 = ~n5953 & n13318 ;
  assign n13320 = n13319 ^ n12594 ^ 1'b0 ;
  assign n13321 = n9557 ^ n5759 ^ 1'b0 ;
  assign n13322 = ~n474 & n13321 ;
  assign n13323 = x4 & n8961 ;
  assign n13324 = n4201 | n8645 ;
  assign n13325 = n13324 ^ n3235 ^ 1'b0 ;
  assign n13326 = n2531 & n6293 ;
  assign n13327 = ( ~n5311 & n6018 ) | ( ~n5311 & n13326 ) | ( n6018 & n13326 ) ;
  assign n13328 = n1730 ^ n315 ^ 1'b0 ;
  assign n13329 = n406 & n8500 ;
  assign n13330 = n13329 ^ n8441 ^ 1'b0 ;
  assign n13331 = n13111 ^ n3611 ^ 1'b0 ;
  assign n13332 = n13331 ^ n3647 ^ 1'b0 ;
  assign n13333 = n502 & ~n1235 ;
  assign n13334 = n13333 ^ n3858 ^ 1'b0 ;
  assign n13335 = n10892 & ~n13334 ;
  assign n13336 = n737 & ~n10003 ;
  assign n13337 = n2588 ^ n133 ^ 1'b0 ;
  assign n13338 = ( n6685 & n13336 ) | ( n6685 & n13337 ) | ( n13336 & n13337 ) ;
  assign n13339 = n8082 & ~n12755 ;
  assign n13340 = n13339 ^ n10895 ^ 1'b0 ;
  assign n13341 = n3050 ^ n2380 ^ 1'b0 ;
  assign n13342 = n5054 | n13341 ;
  assign n13343 = n302 & ~n13342 ;
  assign n13344 = n291 | n13343 ;
  assign n13345 = n13344 ^ n120 ^ 1'b0 ;
  assign n13346 = n9606 ^ n2921 ^ n2337 ;
  assign n13347 = n5757 ^ n3221 ^ 1'b0 ;
  assign n13348 = n27 & n13347 ;
  assign n13349 = n13348 ^ n8350 ^ 1'b0 ;
  assign n13350 = ~n5994 & n12789 ;
  assign n13351 = n3513 ^ n2640 ^ 1'b0 ;
  assign n13352 = n13351 ^ n3655 ^ 1'b0 ;
  assign n13353 = ~n938 & n13352 ;
  assign n13354 = n13353 ^ n12541 ^ 1'b0 ;
  assign n13355 = n5767 & n6723 ;
  assign n13356 = n13355 ^ n8728 ^ 1'b0 ;
  assign n13357 = n873 ^ n539 ^ 1'b0 ;
  assign n13358 = n1230 & ~n10492 ;
  assign n13359 = n6320 ^ n1518 ^ 1'b0 ;
  assign n13360 = n13359 ^ n12504 ^ 1'b0 ;
  assign n13361 = n6298 | n13360 ;
  assign n13362 = n10797 | n13130 ;
  assign n13363 = n13362 ^ n7765 ^ 1'b0 ;
  assign n13364 = n8779 & ~n13363 ;
  assign n13365 = ~n5425 & n10752 ;
  assign n13366 = ~n2176 & n13365 ;
  assign n13371 = ( n1691 & n2685 ) | ( n1691 & n12735 ) | ( n2685 & n12735 ) ;
  assign n13367 = n4782 ^ n3451 ^ 1'b0 ;
  assign n13368 = n4006 & n11383 ;
  assign n13369 = n13368 ^ n4201 ^ 1'b0 ;
  assign n13370 = ( n7134 & ~n13367 ) | ( n7134 & n13369 ) | ( ~n13367 & n13369 ) ;
  assign n13372 = n13371 ^ n13370 ^ 1'b0 ;
  assign n13373 = n8738 & ~n13372 ;
  assign n13374 = n1945 | n4214 ;
  assign n13375 = n968 & ~n13374 ;
  assign n13376 = n13375 ^ n11597 ^ 1'b0 ;
  assign n13377 = n6849 | n13376 ;
  assign n13378 = n6354 & ~n8644 ;
  assign n13379 = n13378 ^ n6955 ^ 1'b0 ;
  assign n13380 = n9323 | n10721 ;
  assign n13381 = n13380 ^ n7581 ^ 1'b0 ;
  assign n13382 = n1425 & ~n7635 ;
  assign n13383 = n2605 & n13382 ;
  assign n13384 = n6059 ^ n5108 ^ 1'b0 ;
  assign n13385 = n13383 | n13384 ;
  assign n13386 = n4921 & n13266 ;
  assign n13387 = n3998 ^ n627 ^ 1'b0 ;
  assign n13388 = n7075 | n13387 ;
  assign n13389 = n11430 ^ n2192 ^ 1'b0 ;
  assign n13390 = n13389 ^ n11223 ^ n5464 ;
  assign n13391 = n5080 & ~n10609 ;
  assign n13392 = n9233 & n9284 ;
  assign n13393 = n2470 ^ n1753 ^ 1'b0 ;
  assign n13394 = n13393 ^ n5071 ^ 1'b0 ;
  assign n13395 = ( n1723 & ~n5468 ) | ( n1723 & n13119 ) | ( ~n5468 & n13119 ) ;
  assign n13396 = n4792 ^ n1539 ^ 1'b0 ;
  assign n13397 = n798 & ~n13396 ;
  assign n13398 = ~n523 & n13397 ;
  assign n13399 = n13398 ^ n8677 ^ 1'b0 ;
  assign n13400 = n1471 | n7951 ;
  assign n13401 = n5052 & n10804 ;
  assign n13402 = ~n1968 & n13401 ;
  assign n13403 = n9405 ^ n1818 ^ 1'b0 ;
  assign n13404 = n13403 ^ n1839 ^ n850 ;
  assign n13405 = n1141 & ~n13404 ;
  assign n13406 = n13405 ^ n11206 ^ 1'b0 ;
  assign n13407 = n13402 | n13406 ;
  assign n13408 = n13152 & n13407 ;
  assign n13410 = n344 & ~n3791 ;
  assign n13411 = n13410 ^ n2682 ^ 1'b0 ;
  assign n13412 = n5658 & n13411 ;
  assign n13409 = n6707 & ~n12587 ;
  assign n13413 = n13412 ^ n13409 ^ 1'b0 ;
  assign n13414 = n7207 | n10370 ;
  assign n13415 = ~n2136 & n13414 ;
  assign n13416 = n1739 & ~n10489 ;
  assign n13417 = n13416 ^ n11999 ^ n5673 ;
  assign n13418 = n6473 & n7726 ;
  assign n13419 = n13418 ^ n12585 ^ 1'b0 ;
  assign n13420 = ( n5121 & n5406 ) | ( n5121 & n5722 ) | ( n5406 & n5722 ) ;
  assign n13421 = n13420 ^ n195 ^ 1'b0 ;
  assign n13422 = ~n1962 & n13421 ;
  assign n13423 = ~n989 & n2004 ;
  assign n13424 = n13423 ^ n2577 ^ 1'b0 ;
  assign n13425 = n6756 | n8042 ;
  assign n13426 = n10262 ^ n1772 ^ 1'b0 ;
  assign n13427 = n12669 & n13426 ;
  assign n13428 = n1353 | n6696 ;
  assign n13429 = n1915 | n13428 ;
  assign n13430 = n7534 & ~n13429 ;
  assign n13431 = n3388 ^ n502 ^ 1'b0 ;
  assign n13432 = n368 | n13431 ;
  assign n13433 = n13432 ^ n7484 ^ 1'b0 ;
  assign n13434 = n1988 & n13433 ;
  assign n13435 = n10897 ^ n3477 ^ 1'b0 ;
  assign n13436 = n5313 & ~n13435 ;
  assign n13437 = ( ~n415 & n848 ) | ( ~n415 & n3893 ) | ( n848 & n3893 ) ;
  assign n13438 = ~n6265 & n9785 ;
  assign n13439 = n5244 & ~n13438 ;
  assign n13440 = n13439 ^ n2849 ^ 1'b0 ;
  assign n13441 = n12695 ^ n3110 ^ 1'b0 ;
  assign n13442 = n683 & ~n3325 ;
  assign n13443 = n12865 ^ n11402 ^ n11097 ;
  assign n13444 = n1912 & n2085 ;
  assign n13445 = n844 | n4158 ;
  assign n13446 = n13444 & ~n13445 ;
  assign n13447 = n13446 ^ n2141 ^ 1'b0 ;
  assign n13448 = n336 & n4871 ;
  assign n13449 = n13448 ^ n2894 ^ 1'b0 ;
  assign n13450 = ~n8163 & n13449 ;
  assign n13451 = ~n3959 & n13450 ;
  assign n13452 = ( n1534 & n4960 ) | ( n1534 & n13451 ) | ( n4960 & n13451 ) ;
  assign n13453 = n1439 & ~n13452 ;
  assign n13454 = n5627 & n13453 ;
  assign n13455 = n11504 ^ n43 ^ 1'b0 ;
  assign n13456 = n4091 | n13455 ;
  assign n13457 = n8611 & ~n13456 ;
  assign n13458 = ~n5823 & n13457 ;
  assign n13459 = n9393 ^ n4677 ^ 1'b0 ;
  assign n13460 = n13270 & ~n13459 ;
  assign n13461 = n1513 & ~n6071 ;
  assign n13462 = n13461 ^ n926 ^ 1'b0 ;
  assign n13463 = n13462 ^ n12438 ^ 1'b0 ;
  assign n13464 = ( n1210 & ~n3871 ) | ( n1210 & n4408 ) | ( ~n3871 & n4408 ) ;
  assign n13465 = n2685 & n3041 ;
  assign n13466 = n2860 ^ n1732 ^ 1'b0 ;
  assign n13467 = n2885 | n13466 ;
  assign n13468 = n2486 | n13467 ;
  assign n13469 = n13465 | n13468 ;
  assign n13470 = n13469 ^ n561 ^ 1'b0 ;
  assign n13471 = ~n9274 & n11975 ;
  assign n13472 = n10161 ^ n7741 ^ 1'b0 ;
  assign n13473 = ~n8076 & n13472 ;
  assign n13474 = n4463 & ~n4696 ;
  assign n13475 = n1351 ^ n451 ^ 1'b0 ;
  assign n13476 = n13475 ^ n4977 ^ 1'b0 ;
  assign n13477 = n11678 & n13476 ;
  assign n13478 = ~n13232 & n13477 ;
  assign n13479 = n10497 ^ n1315 ^ 1'b0 ;
  assign n13480 = n4662 & n8420 ;
  assign n13481 = n13480 ^ n3341 ^ 1'b0 ;
  assign n13482 = n2316 & n3885 ;
  assign n13483 = n571 | n3705 ;
  assign n13484 = n511 | n13483 ;
  assign n13485 = n10217 & ~n13484 ;
  assign n13486 = ~n582 & n5152 ;
  assign n13487 = n13486 ^ n3526 ^ 1'b0 ;
  assign n13488 = n4538 ^ n2252 ^ 1'b0 ;
  assign n13489 = n13488 ^ n13106 ^ 1'b0 ;
  assign n13490 = n2197 ^ n2109 ^ n551 ;
  assign n13491 = n680 | n2031 ;
  assign n13492 = n2871 & ~n13491 ;
  assign n13493 = ~n2005 & n13492 ;
  assign n13494 = ( n9601 & n13490 ) | ( n9601 & ~n13493 ) | ( n13490 & ~n13493 ) ;
  assign n13495 = n318 ^ n138 ^ 1'b0 ;
  assign n13496 = n11778 & ~n13495 ;
  assign n13497 = x5 & ~n1999 ;
  assign n13498 = ~n13496 & n13497 ;
  assign n13499 = n12411 & ~n13498 ;
  assign n13500 = n13494 & n13499 ;
  assign n13501 = n6099 & ~n7556 ;
  assign n13502 = n10665 ^ n9946 ^ 1'b0 ;
  assign n13503 = n885 & ~n13502 ;
  assign n13506 = n3216 ^ n56 ^ 1'b0 ;
  assign n13507 = n5492 & ~n13506 ;
  assign n13504 = n220 & n1055 ;
  assign n13505 = ~n11547 & n13504 ;
  assign n13508 = n13507 ^ n13505 ^ n7176 ;
  assign n13509 = n3967 ^ n2041 ^ 1'b0 ;
  assign n13510 = n9109 | n13509 ;
  assign n13511 = n13510 ^ n6095 ^ 1'b0 ;
  assign n13512 = n3181 ^ n1783 ^ 1'b0 ;
  assign n13513 = ~n7075 & n13512 ;
  assign n13514 = n13513 ^ n9346 ^ 1'b0 ;
  assign n13515 = n4163 & n13514 ;
  assign n13516 = n2376 | n4140 ;
  assign n13517 = n6583 & ~n13516 ;
  assign n13518 = n13515 & ~n13517 ;
  assign n13519 = n13518 ^ n1714 ^ 1'b0 ;
  assign n13520 = n7384 & ~n13519 ;
  assign n13521 = n3390 ^ n2688 ^ 1'b0 ;
  assign n13522 = n2082 & n13521 ;
  assign n13523 = n13522 ^ n1767 ^ 1'b0 ;
  assign n13524 = n7321 ^ n6041 ^ 1'b0 ;
  assign n13525 = n7659 | n12380 ;
  assign n13526 = n13525 ^ n727 ^ 1'b0 ;
  assign n13527 = n13526 ^ n13521 ^ 1'b0 ;
  assign n13528 = n76 & ~n2604 ;
  assign n13529 = n7319 ^ n5906 ^ n883 ;
  assign n13530 = n7246 & ~n13529 ;
  assign n13531 = n13530 ^ n2596 ^ 1'b0 ;
  assign n13532 = n10428 ^ n804 ^ 1'b0 ;
  assign n13533 = ~n13531 & n13532 ;
  assign n13534 = n13533 ^ n5063 ^ 1'b0 ;
  assign n13535 = n13534 ^ n3906 ^ 1'b0 ;
  assign n13536 = n2598 ^ n1087 ^ 1'b0 ;
  assign n13537 = n706 & n13536 ;
  assign n13538 = n13537 ^ n3266 ^ 1'b0 ;
  assign n13539 = n4960 & ~n13538 ;
  assign n13544 = ~n5458 & n8180 ;
  assign n13540 = n8080 ^ n4085 ^ n3548 ;
  assign n13541 = n13540 ^ n9332 ^ n77 ;
  assign n13542 = n7058 & ~n13541 ;
  assign n13543 = ~n7494 & n13542 ;
  assign n13545 = n13544 ^ n13543 ^ 1'b0 ;
  assign n13546 = n904 ^ n488 ^ 1'b0 ;
  assign n13547 = ~n5866 & n13546 ;
  assign n13548 = n12485 & n13547 ;
  assign n13549 = n13548 ^ n6458 ^ 1'b0 ;
  assign n13550 = n974 & n7111 ;
  assign n13551 = n1724 ^ n160 ^ 1'b0 ;
  assign n13552 = ~n5188 & n13551 ;
  assign n13553 = ~n2888 & n13552 ;
  assign n13554 = n13553 ^ n5346 ^ 1'b0 ;
  assign n13555 = n4042 ^ n733 ^ 1'b0 ;
  assign n13556 = ~n8307 & n9740 ;
  assign n13557 = ~n790 & n13556 ;
  assign n13558 = n3504 ^ n20 ^ 1'b0 ;
  assign n13559 = ~n13557 & n13558 ;
  assign n13560 = ~n13555 & n13559 ;
  assign n13561 = n13554 & n13560 ;
  assign n13562 = n9915 ^ n2469 ^ 1'b0 ;
  assign n13563 = n4891 ^ n4185 ^ 1'b0 ;
  assign n13564 = n7621 | n13563 ;
  assign n13565 = n9008 | n13564 ;
  assign n13566 = n10956 | n13565 ;
  assign n13567 = n10589 & ~n12007 ;
  assign n13568 = n6314 & ~n13567 ;
  assign n13569 = ( ~n12686 & n13566 ) | ( ~n12686 & n13568 ) | ( n13566 & n13568 ) ;
  assign n13570 = ~n1204 & n4677 ;
  assign n13571 = n606 & n13570 ;
  assign n13572 = n3242 | n4982 ;
  assign n13573 = n13571 & ~n13572 ;
  assign n13574 = n12337 ^ n3293 ^ 1'b0 ;
  assign n13575 = n996 | n13574 ;
  assign n13578 = n10835 ^ n9089 ^ n3036 ;
  assign n13576 = n3918 ^ n1187 ^ 1'b0 ;
  assign n13577 = ~n10235 & n13576 ;
  assign n13579 = n13578 ^ n13577 ^ 1'b0 ;
  assign n13580 = n2662 & ~n8499 ;
  assign n13581 = n13380 | n13580 ;
  assign n13582 = n8432 ^ n4958 ^ 1'b0 ;
  assign n13583 = n13582 ^ n11438 ^ 1'b0 ;
  assign n13584 = n4027 | n7080 ;
  assign n13585 = n233 | n13584 ;
  assign n13586 = n3837 & ~n13585 ;
  assign n13588 = ~n2869 & n8549 ;
  assign n13587 = n3892 ^ n1726 ^ 1'b0 ;
  assign n13589 = n13588 ^ n13587 ^ 1'b0 ;
  assign n13590 = ~n826 & n13015 ;
  assign n13591 = n12514 ^ n8777 ^ 1'b0 ;
  assign n13592 = n3416 & ~n13591 ;
  assign n13593 = n1703 | n13134 ;
  assign n13594 = n13593 ^ n31 ^ 1'b0 ;
  assign n13595 = n612 & ~n13594 ;
  assign n13596 = n13595 ^ n2007 ^ 1'b0 ;
  assign n13597 = n5234 ^ n764 ^ 1'b0 ;
  assign n13598 = n6951 | n13597 ;
  assign n13599 = n3345 | n7833 ;
  assign n13600 = n6705 & n13599 ;
  assign n13601 = n13600 ^ n11622 ^ 1'b0 ;
  assign n13605 = n4632 ^ n1103 ^ 1'b0 ;
  assign n13602 = n4747 & ~n10475 ;
  assign n13603 = n13602 ^ n9090 ^ 1'b0 ;
  assign n13604 = n7824 | n13603 ;
  assign n13606 = n13605 ^ n13604 ^ 1'b0 ;
  assign n13607 = ~n3939 & n10873 ;
  assign n13608 = n1499 & ~n1538 ;
  assign n13609 = n5627 | n13608 ;
  assign n13610 = n3686 | n13609 ;
  assign n13611 = n12609 & ~n13610 ;
  assign n13612 = n13580 ^ n9753 ^ 1'b0 ;
  assign n13613 = n7564 ^ n492 ^ 1'b0 ;
  assign n13614 = n2476 ^ n732 ^ 1'b0 ;
  assign n13615 = n3158 | n11175 ;
  assign n13616 = n7717 ^ n1933 ^ 1'b0 ;
  assign n13617 = ~n5120 & n13616 ;
  assign n13618 = n9844 ^ n1159 ^ 1'b0 ;
  assign n13619 = n3617 & ~n11167 ;
  assign n13620 = n13618 & n13619 ;
  assign n13621 = ( ~n2287 & n7904 ) | ( ~n2287 & n8749 ) | ( n7904 & n8749 ) ;
  assign n13622 = ~n11021 & n13621 ;
  assign n13623 = ~n13069 & n13622 ;
  assign n13624 = n10076 ^ n7675 ^ 1'b0 ;
  assign n13625 = n5128 & ~n13624 ;
  assign n13626 = n239 & ~n4074 ;
  assign n13627 = n6907 ^ n124 ^ 1'b0 ;
  assign n13628 = n13626 & ~n13627 ;
  assign n13629 = n6578 ^ n682 ^ 1'b0 ;
  assign n13630 = ~n1109 & n13629 ;
  assign n13631 = n8445 & n11193 ;
  assign n13632 = n13631 ^ n7809 ^ 1'b0 ;
  assign n13633 = n4503 ^ n2177 ^ 1'b0 ;
  assign n13634 = ~n13632 & n13633 ;
  assign n13635 = ~n4025 & n5410 ;
  assign n13636 = n13635 ^ n7884 ^ 1'b0 ;
  assign n13637 = n5837 ^ n968 ^ 1'b0 ;
  assign n13638 = n6557 ^ n1861 ^ 1'b0 ;
  assign n13639 = n1915 | n10968 ;
  assign n13656 = n9202 ^ n8814 ^ 1'b0 ;
  assign n13657 = n2733 | n13656 ;
  assign n13654 = n4430 & ~n6176 ;
  assign n13655 = n6176 & n13654 ;
  assign n13658 = n13657 ^ n13655 ^ 1'b0 ;
  assign n13659 = n3794 & n13658 ;
  assign n13640 = n1877 ^ n1425 ^ 1'b0 ;
  assign n13641 = n974 & ~n12570 ;
  assign n13642 = ~n974 & n13641 ;
  assign n13643 = n849 & n13642 ;
  assign n13644 = ~n1072 & n13643 ;
  assign n13645 = ~n1386 & n13644 ;
  assign n13646 = ~n13640 & n13645 ;
  assign n13647 = n1254 & ~n1389 ;
  assign n13648 = ~n1254 & n13647 ;
  assign n13649 = n4324 | n13648 ;
  assign n13650 = n13648 & ~n13649 ;
  assign n13651 = n310 | n13650 ;
  assign n13652 = n13646 & ~n13651 ;
  assign n13653 = n4077 & ~n13652 ;
  assign n13660 = n13659 ^ n13653 ^ 1'b0 ;
  assign n13661 = n471 & ~n12746 ;
  assign n13662 = n1501 | n11434 ;
  assign n13663 = n13662 ^ n12338 ^ 1'b0 ;
  assign n13664 = n275 & n1853 ;
  assign n13665 = ~n6023 & n13664 ;
  assign n13666 = ~n3817 & n6275 ;
  assign n13667 = n4088 & n4146 ;
  assign n13668 = n13667 ^ n282 ^ 1'b0 ;
  assign n13669 = n8000 & ~n13668 ;
  assign n13670 = ~n13666 & n13669 ;
  assign n13671 = n7134 ^ n5334 ^ 1'b0 ;
  assign n13672 = n1439 & n13671 ;
  assign n13673 = n13672 ^ n10134 ^ 1'b0 ;
  assign n13674 = ~n610 & n3111 ;
  assign n13675 = n13674 ^ n3428 ^ 1'b0 ;
  assign n13676 = n13675 ^ n9008 ^ 1'b0 ;
  assign n13677 = ~n752 & n8790 ;
  assign n13678 = n11813 ^ n8346 ^ n7027 ;
  assign n13679 = ~n1864 & n2262 ;
  assign n13680 = n13679 ^ n1280 ^ 1'b0 ;
  assign n13681 = n5525 & n13680 ;
  assign n13682 = n13681 ^ n9606 ^ 1'b0 ;
  assign n13683 = n9676 & ~n13682 ;
  assign n13684 = ~n4395 & n13683 ;
  assign n13687 = ~n403 & n6911 ;
  assign n13685 = n12750 ^ n6396 ^ n4459 ;
  assign n13686 = ~n13495 & n13685 ;
  assign n13688 = n13687 ^ n13686 ^ 1'b0 ;
  assign n13689 = n4702 ^ n712 ^ 1'b0 ;
  assign n13690 = ~n11927 & n13689 ;
  assign n13691 = n1898 & ~n4093 ;
  assign n13692 = n8731 ^ n170 ^ 1'b0 ;
  assign n13693 = n5182 | n9151 ;
  assign n13694 = n7102 | n10199 ;
  assign n13695 = n56 & n5545 ;
  assign n13696 = n13695 ^ n9424 ^ 1'b0 ;
  assign n13697 = n8337 & n12502 ;
  assign n13698 = n11182 | n13697 ;
  assign n13699 = n5049 | n10059 ;
  assign n13700 = n13698 & ~n13699 ;
  assign n13701 = n6827 & n13700 ;
  assign n13702 = n7303 ^ n5903 ^ n3140 ;
  assign n13703 = n4153 | n13702 ;
  assign n13704 = n13703 ^ n1407 ^ 1'b0 ;
  assign n13705 = n8596 | n13704 ;
  assign n13706 = n7266 & ~n13705 ;
  assign n13707 = n10160 & ~n13706 ;
  assign n13708 = ~n395 & n3133 ;
  assign n13709 = n7333 ^ n3993 ^ 1'b0 ;
  assign n13710 = n13708 | n13709 ;
  assign n13711 = n5978 ^ n2358 ^ 1'b0 ;
  assign n13712 = n9821 & n13711 ;
  assign n13713 = n13712 ^ n3957 ^ 1'b0 ;
  assign n13714 = n13069 & n13713 ;
  assign n13715 = n5477 ^ n1533 ^ 1'b0 ;
  assign n13716 = n13715 ^ n7577 ^ n5845 ;
  assign n13717 = n13716 ^ n8737 ^ 1'b0 ;
  assign n13718 = n11893 | n13717 ;
  assign n13719 = n13718 ^ n13524 ^ 1'b0 ;
  assign n13720 = n3974 | n6886 ;
  assign n13721 = n2310 & ~n13720 ;
  assign n13722 = n13721 ^ n9331 ^ 1'b0 ;
  assign n13723 = n4167 | n13722 ;
  assign n13724 = n2619 & n5733 ;
  assign n13725 = n1312 | n3779 ;
  assign n13726 = n5187 | n13725 ;
  assign n13727 = n160 & ~n2881 ;
  assign n13728 = n13727 ^ n3560 ^ 1'b0 ;
  assign n13729 = n13728 ^ n2985 ^ 1'b0 ;
  assign n13730 = n13726 | n13729 ;
  assign n13731 = n3078 ^ n403 ^ 1'b0 ;
  assign n13732 = n13731 ^ n11981 ^ 1'b0 ;
  assign n13733 = n148 | n12967 ;
  assign n13734 = n3866 & ~n13733 ;
  assign n13735 = ~n1700 & n7322 ;
  assign n13736 = ~n2371 & n11274 ;
  assign n13737 = n2802 | n13210 ;
  assign n13738 = n6584 ^ n2243 ^ 1'b0 ;
  assign n13739 = n40 | n13738 ;
  assign n13740 = ( n6665 & ~n10479 ) | ( n6665 & n13739 ) | ( ~n10479 & n13739 ) ;
  assign n13741 = n4141 ^ n2736 ^ n2050 ;
  assign n13742 = n7841 | n13741 ;
  assign n13743 = n5726 & n8392 ;
  assign n13744 = n2512 & n6406 ;
  assign n13745 = n5477 | n8392 ;
  assign n13746 = n13745 ^ n5081 ^ 1'b0 ;
  assign n13747 = ~n13180 & n13746 ;
  assign n13748 = n13613 ^ n3367 ^ 1'b0 ;
  assign n13749 = n1728 | n8648 ;
  assign n13750 = n3101 & ~n13749 ;
  assign n13751 = n5058 ^ n4600 ^ 1'b0 ;
  assign n13752 = n851 | n11142 ;
  assign n13753 = n13752 ^ n4343 ^ 1'b0 ;
  assign n13754 = n13753 ^ n5511 ^ 1'b0 ;
  assign n13755 = n4409 ^ n1431 ^ 1'b0 ;
  assign n13756 = ( n8578 & n10881 ) | ( n8578 & ~n13163 ) | ( n10881 & ~n13163 ) ;
  assign n13757 = n8031 | n12076 ;
  assign n13758 = n9762 | n13757 ;
  assign n13759 = ~n7179 & n13758 ;
  assign n13760 = n13759 ^ n10832 ^ 1'b0 ;
  assign n13761 = n3502 | n11194 ;
  assign n13762 = n10331 ^ n415 ^ 1'b0 ;
  assign n13763 = n2799 & n9426 ;
  assign n13764 = n8436 & ~n12842 ;
  assign n13765 = n754 & n13764 ;
  assign n13766 = ~n10015 & n13050 ;
  assign n13767 = n13766 ^ n6247 ^ 1'b0 ;
  assign n13768 = ~n13765 & n13767 ;
  assign n13769 = n7360 & n13768 ;
  assign n13770 = n736 & ~n11208 ;
  assign n13771 = n342 & n13770 ;
  assign n13772 = n572 & n11043 ;
  assign n13773 = ~n8789 & n13772 ;
  assign n13774 = n13773 ^ n409 ^ 1'b0 ;
  assign n13775 = n1988 ^ n835 ^ 1'b0 ;
  assign n13776 = n4068 & ~n13775 ;
  assign n13777 = ( ~n4645 & n6550 ) | ( ~n4645 & n13776 ) | ( n6550 & n13776 ) ;
  assign n13778 = n13777 ^ n1568 ^ 1'b0 ;
  assign n13785 = n7169 ^ n5197 ^ n1177 ;
  assign n13779 = n3671 & n4474 ;
  assign n13780 = ~n4474 & n13779 ;
  assign n13781 = n1002 & ~n4220 ;
  assign n13782 = n4220 & n13781 ;
  assign n13783 = n3777 & ~n13782 ;
  assign n13784 = ~n13780 & n13783 ;
  assign n13786 = n13785 ^ n13784 ^ 1'b0 ;
  assign n13787 = n2850 ^ n2390 ^ n122 ;
  assign n13788 = n7416 ^ n710 ^ 1'b0 ;
  assign n13789 = n13787 | n13788 ;
  assign n13794 = n3693 | n5475 ;
  assign n13790 = n6099 ^ n5615 ^ 1'b0 ;
  assign n13791 = n13790 ^ n1413 ^ 1'b0 ;
  assign n13792 = n11189 & n13791 ;
  assign n13793 = n2073 & n13792 ;
  assign n13795 = n13794 ^ n13793 ^ 1'b0 ;
  assign n13796 = n737 & ~n4088 ;
  assign n13797 = n225 & n13796 ;
  assign n13798 = n3108 ^ n2233 ^ 1'b0 ;
  assign n13799 = n7069 & n13798 ;
  assign n13800 = n13797 & n13799 ;
  assign n13801 = ~n1484 & n2390 ;
  assign n13802 = n2547 & ~n4738 ;
  assign n13803 = n13801 | n13802 ;
  assign n13804 = n4917 & n5059 ;
  assign n13805 = n13804 ^ n9195 ^ 1'b0 ;
  assign n13806 = n2039 | n10976 ;
  assign n13807 = n7593 | n8000 ;
  assign n13808 = n13807 ^ n9375 ^ 1'b0 ;
  assign n13817 = n7211 ^ n722 ^ 1'b0 ;
  assign n13814 = n606 | n6185 ;
  assign n13815 = n606 & ~n13814 ;
  assign n13816 = n1644 & n13815 ;
  assign n13809 = n5857 ^ n1564 ^ 1'b0 ;
  assign n13810 = n3962 | n13809 ;
  assign n13811 = n13809 & ~n13810 ;
  assign n13812 = n622 | n13811 ;
  assign n13813 = n13811 & ~n13812 ;
  assign n13818 = n13817 ^ n13816 ^ n13813 ;
  assign n13819 = ~n5367 & n5673 ;
  assign n13820 = n13819 ^ n12550 ^ 1'b0 ;
  assign n13821 = n13122 ^ n6241 ^ 1'b0 ;
  assign n13822 = n13821 ^ n11468 ^ 1'b0 ;
  assign n13823 = ~n7634 & n13822 ;
  assign n13824 = n1660 & n10114 ;
  assign n13825 = n13824 ^ n13750 ^ 1'b0 ;
  assign n13826 = n2953 & n9511 ;
  assign n13827 = n11333 & n13826 ;
  assign n13828 = n11834 ^ n1063 ^ 1'b0 ;
  assign n13829 = ~n8139 & n8312 ;
  assign n13830 = ~n3197 & n3694 ;
  assign n13831 = ~n10620 & n13830 ;
  assign n13832 = ( n2584 & n2756 ) | ( n2584 & ~n13279 ) | ( n2756 & ~n13279 ) ;
  assign n13833 = n4228 ^ n1853 ^ 1'b0 ;
  assign n13834 = n1845 ^ n214 ^ 1'b0 ;
  assign n13835 = n13833 & ~n13834 ;
  assign n13836 = n12740 ^ n3207 ^ 1'b0 ;
  assign n13837 = n13836 ^ n10775 ^ 1'b0 ;
  assign n13838 = n1868 & n13837 ;
  assign n13839 = n851 & ~n13668 ;
  assign n13840 = n13839 ^ n7177 ^ n4079 ;
  assign n13841 = n1546 & n8023 ;
  assign n13842 = n4395 | n5832 ;
  assign n13843 = n12158 & ~n13842 ;
  assign n13844 = n2618 & ~n13843 ;
  assign n13845 = ~n10466 & n13844 ;
  assign n13846 = n13841 & n13845 ;
  assign n13847 = n1865 | n2948 ;
  assign n13848 = n13846 | n13847 ;
  assign n13849 = n13526 ^ n6479 ^ 1'b0 ;
  assign n13850 = n5759 | n6226 ;
  assign n13851 = n13850 ^ n1247 ^ 1'b0 ;
  assign n13852 = n8759 ^ n1126 ^ 1'b0 ;
  assign n13853 = n13852 ^ n3903 ^ 1'b0 ;
  assign n13854 = n7437 & n13853 ;
  assign n13855 = n10517 ^ n106 ^ 1'b0 ;
  assign n13856 = n6077 | n13855 ;
  assign n13857 = n2239 & ~n13856 ;
  assign n13858 = ~n3372 & n8399 ;
  assign n13859 = n8237 & n9336 ;
  assign n13860 = n13858 & n13859 ;
  assign n13861 = n1802 ^ n1050 ^ 1'b0 ;
  assign n13862 = n746 & n7382 ;
  assign n13863 = ~n10101 & n13002 ;
  assign n13864 = n5281 & ~n13070 ;
  assign n13865 = n4007 | n13864 ;
  assign n13866 = n8070 | n13865 ;
  assign n13867 = n19 | n1269 ;
  assign n13868 = n1448 & ~n13867 ;
  assign n13869 = n8284 | n13868 ;
  assign n13870 = n8103 ^ n5607 ^ 1'b0 ;
  assign n13871 = n11761 & ~n13870 ;
  assign n13872 = n9218 & n11378 ;
  assign n13873 = ~n6748 & n13872 ;
  assign n13874 = n13858 | n13873 ;
  assign n13875 = n3035 & n13874 ;
  assign n13876 = ~n470 & n1138 ;
  assign n13877 = n4674 & ~n13876 ;
  assign n13878 = n5242 & ~n13877 ;
  assign n13879 = n4119 & ~n5724 ;
  assign n13880 = n9776 ^ n422 ^ 1'b0 ;
  assign n13881 = n13879 & n13880 ;
  assign n13882 = n13881 ^ n11287 ^ 1'b0 ;
  assign n13883 = n13878 & n13882 ;
  assign n13884 = n1886 & n4765 ;
  assign n13885 = n8207 & n13884 ;
  assign n13886 = n2262 & ~n4745 ;
  assign n13887 = n10319 & n13886 ;
  assign n13888 = n9151 ^ n3116 ^ 1'b0 ;
  assign n13889 = n13887 | n13888 ;
  assign n13890 = n27 & ~n7618 ;
  assign n13891 = n13890 ^ n532 ^ 1'b0 ;
  assign n13892 = n2159 & n4690 ;
  assign n13893 = n13892 ^ n6632 ^ 1'b0 ;
  assign n13894 = n2950 | n10073 ;
  assign n13895 = n10670 & ~n13894 ;
  assign n13896 = ( n8461 & ~n11829 ) | ( n8461 & n12246 ) | ( ~n11829 & n12246 ) ;
  assign n13897 = n978 & ~n8716 ;
  assign n13898 = n4209 & n13897 ;
  assign n13899 = n1548 & n13898 ;
  assign n13900 = n12406 & ~n13207 ;
  assign n13901 = n11497 ^ n5442 ^ 1'b0 ;
  assign n13902 = n312 & ~n6621 ;
  assign n13903 = ~n6943 & n13902 ;
  assign n13904 = n13901 | n13903 ;
  assign n13905 = n10908 ^ n1543 ^ 1'b0 ;
  assign n13906 = n13905 ^ n2094 ^ 1'b0 ;
  assign n13907 = n10338 & n13906 ;
  assign n13910 = n5111 & ~n5788 ;
  assign n13908 = ~n3295 & n6226 ;
  assign n13909 = n13908 ^ n6769 ^ 1'b0 ;
  assign n13911 = n13910 ^ n13909 ^ n10181 ;
  assign n13912 = n3083 & ~n7848 ;
  assign n13913 = n7137 ^ n6924 ^ 1'b0 ;
  assign n13914 = n10003 ^ n5841 ^ 1'b0 ;
  assign n13915 = ~n8728 & n13914 ;
  assign n13916 = n10504 ^ n8942 ^ n2771 ;
  assign n13917 = n12409 & n13694 ;
  assign n13918 = ~n6701 & n13917 ;
  assign n13919 = n9685 ^ n7567 ^ 1'b0 ;
  assign n13921 = n1434 & n5365 ;
  assign n13920 = n5821 ^ n5365 ^ 1'b0 ;
  assign n13922 = n13921 ^ n13920 ^ 1'b0 ;
  assign n13923 = n13922 ^ n3448 ^ 1'b0 ;
  assign n13924 = ~n6275 & n13923 ;
  assign n13925 = n11839 ^ n2455 ^ 1'b0 ;
  assign n13926 = n3602 ^ n2872 ^ n1711 ;
  assign n13927 = n13404 ^ n6834 ^ n899 ;
  assign n13928 = n5139 ^ n3226 ^ 1'b0 ;
  assign n13929 = n625 & ~n13928 ;
  assign n13930 = ~n5368 & n13929 ;
  assign n13931 = n13930 ^ n11655 ^ 1'b0 ;
  assign n13932 = n13931 ^ n8543 ^ 1'b0 ;
  assign n13933 = ~n12671 & n13932 ;
  assign n13934 = ~n1327 & n3114 ;
  assign n13935 = n9744 ^ n3990 ^ 1'b0 ;
  assign n13936 = n9743 | n13935 ;
  assign n13937 = n11427 | n13936 ;
  assign n13938 = n13879 ^ n7377 ^ 1'b0 ;
  assign n13939 = n419 & ~n13938 ;
  assign n13940 = n125 | n1087 ;
  assign n13941 = n1289 | n13940 ;
  assign n13942 = ~n5348 & n13941 ;
  assign n13943 = ~n11927 & n13942 ;
  assign n13944 = ~n442 & n1382 ;
  assign n13945 = n298 & n2478 ;
  assign n13946 = ~n12733 & n13945 ;
  assign n13947 = n420 | n849 ;
  assign n13948 = ~n11729 & n13947 ;
  assign n13949 = n13948 ^ n8433 ^ 1'b0 ;
  assign n13950 = n4182 & n12854 ;
  assign n13951 = n13950 ^ n6805 ^ 1'b0 ;
  assign n13952 = n6730 ^ n768 ^ 1'b0 ;
  assign n13953 = n2228 | n13952 ;
  assign n13954 = n12172 ^ n4787 ^ 1'b0 ;
  assign n13955 = ~n13953 & n13954 ;
  assign n13956 = n13955 ^ n349 ^ 1'b0 ;
  assign n13957 = n3848 ^ n2574 ^ n2236 ;
  assign n13958 = n9109 ^ n1715 ^ 1'b0 ;
  assign n13959 = n3190 | n13958 ;
  assign n13960 = n13957 | n13959 ;
  assign n13961 = n466 & ~n3324 ;
  assign n13962 = n9667 | n11610 ;
  assign n13963 = n13961 | n13962 ;
  assign n13964 = n5861 | n13963 ;
  assign n13965 = ~n8174 & n13964 ;
  assign n13966 = n2662 | n5001 ;
  assign n13967 = n13966 ^ n6711 ^ 1'b0 ;
  assign n13968 = n3915 & n13967 ;
  assign n13969 = n10942 ^ n4037 ^ 1'b0 ;
  assign n13970 = n3822 & n13969 ;
  assign n13971 = n13970 ^ n9427 ^ 1'b0 ;
  assign n13972 = n11710 ^ n7813 ^ 1'b0 ;
  assign n13973 = n12249 | n13972 ;
  assign n13974 = n2660 & ~n13664 ;
  assign n13975 = n13974 ^ n3036 ^ 1'b0 ;
  assign n13976 = n1111 | n3301 ;
  assign n13977 = n1732 | n13976 ;
  assign n13978 = ~n4497 & n13977 ;
  assign n13979 = ~n13975 & n13978 ;
  assign n13980 = ( n1814 & n13973 ) | ( n1814 & ~n13979 ) | ( n13973 & ~n13979 ) ;
  assign n13981 = n13980 ^ n9636 ^ n4666 ;
  assign n13982 = n6398 ^ n4287 ^ 1'b0 ;
  assign n13983 = ~n6797 & n13982 ;
  assign n13984 = n13983 ^ n9133 ^ 1'b0 ;
  assign n13985 = n1208 ^ n140 ^ 1'b0 ;
  assign n13986 = n7593 ^ n115 ^ 1'b0 ;
  assign n13987 = ~n8862 & n13535 ;
  assign n13988 = n1851 & n13987 ;
  assign n13989 = ~n3753 & n7899 ;
  assign n13990 = n13989 ^ n2682 ^ 1'b0 ;
  assign n13991 = n10400 & ~n12921 ;
  assign n13992 = n4269 | n5367 ;
  assign n13993 = n61 | n2028 ;
  assign n13994 = n13992 | n13993 ;
  assign n13995 = ~n8801 & n13994 ;
  assign n14000 = n110 | n1838 ;
  assign n14001 = n14000 ^ n8880 ^ 1'b0 ;
  assign n13998 = n1336 ^ x9 ^ 1'b0 ;
  assign n13996 = n5393 ^ n2062 ^ n1522 ;
  assign n13997 = n3521 & ~n13996 ;
  assign n13999 = n13998 ^ n13997 ^ 1'b0 ;
  assign n14002 = n14001 ^ n13999 ^ 1'b0 ;
  assign n14003 = n13995 & ~n14002 ;
  assign n14004 = ~n3031 & n4012 ;
  assign n14005 = n878 & n14004 ;
  assign n14006 = ~n3095 & n14005 ;
  assign n14007 = n133 | n8391 ;
  assign n14008 = n13702 ^ n7943 ^ n6074 ;
  assign n14009 = n1369 & ~n14008 ;
  assign n14010 = n14007 & ~n14009 ;
  assign n14011 = n3158 | n11690 ;
  assign n14012 = n8322 ^ n968 ^ 1'b0 ;
  assign n14013 = n1469 & n8470 ;
  assign n14014 = n1252 & ~n10795 ;
  assign n14016 = n5362 ^ n1742 ^ 1'b0 ;
  assign n14017 = n4353 | n14016 ;
  assign n14018 = n1066 | n14017 ;
  assign n14019 = n14018 ^ n8490 ^ 1'b0 ;
  assign n14015 = n1422 & ~n11904 ;
  assign n14020 = n14019 ^ n14015 ^ 1'b0 ;
  assign n14021 = n14020 ^ n10533 ^ 1'b0 ;
  assign n14022 = n2796 | n14021 ;
  assign n14023 = n2927 | n14022 ;
  assign n14024 = n14014 | n14023 ;
  assign n14026 = n5107 ^ n4166 ^ 1'b0 ;
  assign n14027 = n4170 & ~n14026 ;
  assign n14025 = n1834 & n8860 ;
  assign n14028 = n14027 ^ n14025 ^ 1'b0 ;
  assign n14029 = n2560 | n10743 ;
  assign n14030 = n6586 ^ n1256 ^ 1'b0 ;
  assign n14031 = n3037 ^ n2131 ^ 1'b0 ;
  assign n14032 = ~n831 & n14031 ;
  assign n14036 = ~n6231 & n8658 ;
  assign n14037 = n4754 & n14036 ;
  assign n14033 = n7653 | n8161 ;
  assign n14034 = n8331 & ~n14033 ;
  assign n14035 = n2802 | n14034 ;
  assign n14038 = n14037 ^ n14035 ^ 1'b0 ;
  assign n14039 = n8230 & n13505 ;
  assign n14040 = n11763 ^ n10018 ^ 1'b0 ;
  assign n14041 = ~n6271 & n14040 ;
  assign n14042 = n4519 | n12511 ;
  assign n14043 = n5688 & n7321 ;
  assign n14044 = ~n5484 & n14043 ;
  assign n14045 = n4034 ^ n423 ^ 1'b0 ;
  assign n14046 = ~n4041 & n13547 ;
  assign n14047 = n1169 & n3942 ;
  assign n14048 = n14047 ^ n4420 ^ 1'b0 ;
  assign n14049 = n6607 & n14048 ;
  assign n14050 = n1832 | n14049 ;
  assign n14051 = n2574 & ~n12272 ;
  assign n14052 = n13582 & n14051 ;
  assign n14053 = n14052 ^ n5523 ^ 1'b0 ;
  assign n14054 = n14053 ^ n8695 ^ n8082 ;
  assign n14055 = n846 & ~n8305 ;
  assign n14056 = ~n14017 & n14055 ;
  assign n14057 = n14056 ^ n1395 ^ 1'b0 ;
  assign n14058 = n3201 ^ n3026 ^ n1024 ;
  assign n14059 = n6208 | n6518 ;
  assign n14060 = ~n14058 & n14059 ;
  assign n14061 = ~n3947 & n14060 ;
  assign n14062 = ~n9443 & n12422 ;
  assign n14063 = ~n8212 & n14062 ;
  assign n14064 = n14061 & ~n14063 ;
  assign n14065 = n10208 ^ n3512 ^ 1'b0 ;
  assign n14066 = ~n3550 & n14065 ;
  assign n14067 = n8885 ^ n7474 ^ 1'b0 ;
  assign n14068 = n3093 & ~n8478 ;
  assign n14069 = n6356 ^ n4712 ^ 1'b0 ;
  assign n14070 = n5828 & ~n12299 ;
  assign n14071 = n121 & n9153 ;
  assign n14072 = n6323 | n14071 ;
  assign n14073 = n14072 ^ n10195 ^ 1'b0 ;
  assign n14074 = n3756 & n4674 ;
  assign n14075 = n14074 ^ n12653 ^ 1'b0 ;
  assign n14076 = n4935 | n9707 ;
  assign n14077 = n978 & n3235 ;
  assign n14078 = n14076 & n14077 ;
  assign n14079 = n5454 ^ n3335 ^ 1'b0 ;
  assign n14080 = ~n5240 & n14079 ;
  assign n14081 = ( n1914 & n11217 ) | ( n1914 & n14080 ) | ( n11217 & n14080 ) ;
  assign n14082 = n10166 ^ n4895 ^ 1'b0 ;
  assign n14083 = n11897 & n14082 ;
  assign n14084 = n6644 | n10201 ;
  assign n14085 = n14084 ^ n3544 ^ 1'b0 ;
  assign n14086 = n7400 & n14085 ;
  assign n14087 = n5916 & ~n7105 ;
  assign n14088 = n14087 ^ n3383 ^ 1'b0 ;
  assign n14089 = n428 & n2308 ;
  assign n14090 = n2261 & ~n13124 ;
  assign n14091 = n14090 ^ n2802 ^ 1'b0 ;
  assign n14092 = n11140 & n14091 ;
  assign n14093 = n14092 ^ n2993 ^ 1'b0 ;
  assign n14094 = n10253 ^ n8068 ^ n7620 ;
  assign n14095 = ( ~n9730 & n11462 ) | ( ~n9730 & n14094 ) | ( n11462 & n14094 ) ;
  assign n14096 = n7808 | n11825 ;
  assign n14097 = n1645 & ~n14096 ;
  assign n14098 = n4965 | n12366 ;
  assign n14099 = x4 | n14098 ;
  assign n14100 = n2435 | n7611 ;
  assign n14101 = n14100 ^ n4001 ^ 1'b0 ;
  assign n14102 = n14099 & n14101 ;
  assign n14103 = n9612 & n14102 ;
  assign n14104 = n14097 & n14103 ;
  assign n14107 = n10917 ^ n362 ^ 1'b0 ;
  assign n14105 = n5660 ^ n1366 ^ 1'b0 ;
  assign n14106 = ~n5571 & n14105 ;
  assign n14108 = n14107 ^ n14106 ^ n9205 ;
  assign n14109 = n865 | n8138 ;
  assign n14110 = n11166 ^ n7695 ^ 1'b0 ;
  assign n14111 = n14109 & ~n14110 ;
  assign n14112 = n11274 ^ n536 ^ 1'b0 ;
  assign n14113 = n5067 & n14112 ;
  assign n14114 = n14113 ^ n13100 ^ 1'b0 ;
  assign n14115 = n8819 ^ n2719 ^ 1'b0 ;
  assign n14116 = n5329 & n12100 ;
  assign n14117 = n12249 ^ n12091 ^ 1'b0 ;
  assign n14118 = n5142 | n11194 ;
  assign n14119 = n3690 & ~n14118 ;
  assign n14120 = n14119 ^ n3818 ^ 1'b0 ;
  assign n14121 = n620 & ~n14120 ;
  assign n14122 = n14081 ^ n11726 ^ 1'b0 ;
  assign n14123 = n1310 & n5331 ;
  assign n14124 = n11220 & ~n14123 ;
  assign n14125 = ~n35 & n2581 ;
  assign n14126 = ( n3218 & n8738 ) | ( n3218 & ~n9036 ) | ( n8738 & ~n9036 ) ;
  assign n14127 = n11774 & ~n13925 ;
  assign n14128 = n11678 ^ n6997 ^ 1'b0 ;
  assign n14129 = n1564 & ~n14128 ;
  assign n14130 = ~n1556 & n5824 ;
  assign n14131 = n4550 & n14130 ;
  assign n14132 = ~n5759 & n14131 ;
  assign n14133 = n2060 & n7116 ;
  assign n14134 = n5497 & n14133 ;
  assign n14135 = n5191 & ~n8086 ;
  assign n14136 = n11426 ^ n7239 ^ 1'b0 ;
  assign n14137 = n8136 & ~n11740 ;
  assign n14138 = n9219 & ~n10580 ;
  assign n14139 = n10828 ^ n8485 ^ 1'b0 ;
  assign n14140 = n14138 & n14139 ;
  assign n14141 = n14140 ^ n11374 ^ 1'b0 ;
  assign n14142 = ~n8027 & n14141 ;
  assign n14143 = n6702 ^ n6124 ^ 1'b0 ;
  assign n14144 = ~n6131 & n14143 ;
  assign n14145 = ~n3331 & n14144 ;
  assign n14146 = n488 & n6765 ;
  assign n14147 = ~n9385 & n11980 ;
  assign n14148 = n738 & ~n14147 ;
  assign n14152 = n4024 ^ n316 ^ 1'b0 ;
  assign n14153 = n14152 ^ n4185 ^ 1'b0 ;
  assign n14154 = n574 | n14153 ;
  assign n14155 = n6004 & ~n14154 ;
  assign n14149 = n802 | n3574 ;
  assign n14150 = n11179 ^ n788 ^ 1'b0 ;
  assign n14151 = n14149 & n14150 ;
  assign n14156 = n14155 ^ n14151 ^ 1'b0 ;
  assign n14157 = ~n6135 & n14156 ;
  assign n14158 = n14157 ^ n2899 ^ 1'b0 ;
  assign n14159 = n1485 | n4951 ;
  assign n14160 = ( ~n437 & n3970 ) | ( ~n437 & n14159 ) | ( n3970 & n14159 ) ;
  assign n14161 = ~n264 & n7251 ;
  assign n14162 = n3678 & n6392 ;
  assign n14163 = n14162 ^ n5721 ^ 1'b0 ;
  assign n14164 = n10311 & ~n14163 ;
  assign n14165 = n1978 | n14164 ;
  assign n14166 = n7530 ^ n4276 ^ n2101 ;
  assign n14167 = n6342 ^ n5685 ^ 1'b0 ;
  assign n14168 = ~n919 & n3258 ;
  assign n14169 = n14168 ^ n7687 ^ 1'b0 ;
  assign n14170 = ~n1329 & n2409 ;
  assign n14171 = ~n2334 & n7456 ;
  assign n14172 = n3616 & ~n14171 ;
  assign n14173 = n14172 ^ n11521 ^ 1'b0 ;
  assign n14174 = n1946 & ~n12201 ;
  assign n14175 = n14174 ^ n7524 ^ 1'b0 ;
  assign n14176 = n122 | n1771 ;
  assign n14177 = n347 & ~n14176 ;
  assign n14178 = n2045 & ~n14177 ;
  assign n14179 = ~n2045 & n14178 ;
  assign n14180 = n5342 ^ n780 ^ 1'b0 ;
  assign n14181 = n14179 | n14180 ;
  assign n14182 = n14179 & ~n14181 ;
  assign n14185 = ~n5880 & n6224 ;
  assign n14186 = ~n6224 & n14185 ;
  assign n14183 = n4774 ^ n883 ^ 1'b0 ;
  assign n14184 = ~n13959 & n14183 ;
  assign n14187 = n14186 ^ n14184 ^ 1'b0 ;
  assign n14188 = ~n14182 & n14187 ;
  assign n14189 = n160 & n920 ;
  assign n14190 = ~n159 & n14189 ;
  assign n14191 = n14190 ^ n8667 ^ n2367 ;
  assign n14192 = ( n722 & ~n2663 ) | ( n722 & n5813 ) | ( ~n2663 & n5813 ) ;
  assign n14193 = ~n2260 & n14192 ;
  assign n14194 = n14191 & n14193 ;
  assign n14195 = ~n33 & n1668 ;
  assign n14196 = n14194 & n14195 ;
  assign n14197 = n533 & ~n3299 ;
  assign n14198 = n71 | n1852 ;
  assign n14199 = n1853 & ~n8074 ;
  assign n14200 = n14199 ^ n11542 ^ 1'b0 ;
  assign n14201 = n2359 & ~n14200 ;
  assign n14202 = n14201 ^ n1276 ^ 1'b0 ;
  assign n14203 = n14198 & ~n14202 ;
  assign n14204 = n121 & n14203 ;
  assign n14205 = n14204 ^ n3086 ^ 1'b0 ;
  assign n14208 = n8459 ^ n1685 ^ 1'b0 ;
  assign n14206 = n2262 ^ n1694 ^ 1'b0 ;
  assign n14207 = n14206 ^ n12070 ^ 1'b0 ;
  assign n14209 = n14208 ^ n14207 ^ 1'b0 ;
  assign n14210 = ~n14205 & n14209 ;
  assign n14211 = ~n3866 & n8021 ;
  assign n14212 = n14211 ^ n2409 ^ 1'b0 ;
  assign n14213 = n14212 ^ n2610 ^ 1'b0 ;
  assign n14216 = n8702 ^ n4433 ^ 1'b0 ;
  assign n14217 = n1464 & ~n14216 ;
  assign n14214 = n1276 ^ n1134 ^ 1'b0 ;
  assign n14215 = n6433 & n14214 ;
  assign n14218 = n14217 ^ n14215 ^ 1'b0 ;
  assign n14219 = n251 | n14218 ;
  assign n14220 = ~n8259 & n11865 ;
  assign n14226 = n6833 ^ n4138 ^ n2133 ;
  assign n14221 = n4738 ^ n3270 ^ 1'b0 ;
  assign n14222 = n11068 & n14221 ;
  assign n14223 = n8192 & n14222 ;
  assign n14224 = n7312 | n14223 ;
  assign n14225 = n14224 ^ n4014 ^ 1'b0 ;
  assign n14227 = n14226 ^ n14225 ^ 1'b0 ;
  assign n14228 = n3319 | n7784 ;
  assign n14229 = ~n10582 & n11388 ;
  assign n14230 = n4958 ^ n931 ^ 1'b0 ;
  assign n14231 = n4732 ^ n301 ^ 1'b0 ;
  assign n14232 = n6473 ^ n6409 ^ 1'b0 ;
  assign n14233 = n2549 & ~n14232 ;
  assign n14234 = n5540 ^ n1724 ^ n615 ;
  assign n14235 = n14234 ^ n4528 ^ n1790 ;
  assign n14236 = n48 | n14235 ;
  assign n14237 = n8922 ^ n4476 ^ 1'b0 ;
  assign n14240 = n1336 & n1370 ;
  assign n14241 = n14240 ^ n6777 ^ 1'b0 ;
  assign n14238 = n3746 | n4391 ;
  assign n14239 = n12079 | n14238 ;
  assign n14242 = n14241 ^ n14239 ^ 1'b0 ;
  assign n14243 = n6455 ^ n181 ^ 1'b0 ;
  assign n14244 = ( ~n1363 & n8299 ) | ( ~n1363 & n14243 ) | ( n8299 & n14243 ) ;
  assign n14245 = n3096 | n3384 ;
  assign n14246 = n1829 | n14245 ;
  assign n14247 = n8168 | n14246 ;
  assign n14248 = n4773 | n8150 ;
  assign n14249 = ~n9453 & n14248 ;
  assign n14250 = n11825 ^ n6057 ^ 1'b0 ;
  assign n14251 = n11356 | n14250 ;
  assign n14252 = n642 & ~n10479 ;
  assign n14253 = n4712 ^ n995 ^ n675 ;
  assign n14254 = n7967 & n14001 ;
  assign n14255 = ~n8413 & n9741 ;
  assign n14256 = n12634 ^ n428 ^ 1'b0 ;
  assign n14257 = ~n13234 & n14256 ;
  assign n14258 = n1568 & n14257 ;
  assign n14259 = n8211 ^ n4477 ^ n1109 ;
  assign n14260 = n14259 ^ n5779 ^ 1'b0 ;
  assign n14261 = n302 ^ x3 ^ 1'b0 ;
  assign n14262 = n4962 ^ n1114 ^ 1'b0 ;
  assign n14263 = n3171 & ~n8784 ;
  assign n14264 = ~n5008 & n14263 ;
  assign n14265 = n5714 & ~n14264 ;
  assign n14266 = n14265 ^ n7596 ^ 1'b0 ;
  assign n14267 = n5688 ^ n3082 ^ 1'b0 ;
  assign n14270 = ~n30 & n1365 ;
  assign n14271 = ~n9854 & n14270 ;
  assign n14272 = n14271 ^ n2455 ^ 1'b0 ;
  assign n14268 = n4380 | n6570 ;
  assign n14269 = ~n6476 & n14268 ;
  assign n14273 = n14272 ^ n14269 ^ 1'b0 ;
  assign n14274 = n14267 & n14273 ;
  assign n14275 = n246 & n4668 ;
  assign n14276 = n14275 ^ n5077 ^ 1'b0 ;
  assign n14277 = ~n4305 & n4543 ;
  assign n14278 = n11148 & n14277 ;
  assign n14279 = n14278 ^ n7686 ^ 1'b0 ;
  assign n14280 = ( x5 & n4088 ) | ( x5 & n6239 ) | ( n4088 & n6239 ) ;
  assign n14281 = ~n4942 & n11819 ;
  assign n14282 = n6095 ^ n4090 ^ 1'b0 ;
  assign n14283 = n2637 & ~n4228 ;
  assign n14284 = n14283 ^ n11774 ^ 1'b0 ;
  assign n14285 = ( n2761 & ~n7965 ) | ( n2761 & n14284 ) | ( ~n7965 & n14284 ) ;
  assign n14286 = n11497 ^ n3817 ^ 1'b0 ;
  assign n14287 = n10745 & ~n11511 ;
  assign n14288 = n10142 & n10774 ;
  assign n14289 = n3822 ^ n3298 ^ n3147 ;
  assign n14290 = ~n1392 & n14289 ;
  assign n14291 = n14288 & n14290 ;
  assign n14292 = n4460 & ~n5085 ;
  assign n14293 = n14291 & n14292 ;
  assign n14294 = n1284 | n2812 ;
  assign n14295 = n7492 | n14294 ;
  assign n14296 = n7389 & n12990 ;
  assign n14297 = n14296 ^ n5058 ^ 1'b0 ;
  assign n14298 = x8 & ~n14297 ;
  assign n14299 = n14298 ^ n4883 ^ 1'b0 ;
  assign n14300 = n2986 ^ n1870 ^ 1'b0 ;
  assign n14301 = n4529 | n14300 ;
  assign n14302 = n14301 ^ n3766 ^ 1'b0 ;
  assign n14306 = n2616 & ~n2948 ;
  assign n14303 = n3078 & ~n5199 ;
  assign n14304 = n14303 ^ n311 ^ 1'b0 ;
  assign n14305 = n14304 ^ n10582 ^ 1'b0 ;
  assign n14307 = n14306 ^ n14305 ^ n1449 ;
  assign n14308 = n2079 & n2769 ;
  assign n14309 = n2693 ^ n1078 ^ 1'b0 ;
  assign n14310 = n10264 | n14309 ;
  assign n14311 = n14308 & ~n14310 ;
  assign n14312 = n2549 & ~n12117 ;
  assign n14314 = ~n3693 & n5854 ;
  assign n14315 = n14314 ^ n5497 ^ 1'b0 ;
  assign n14313 = n6151 | n9291 ;
  assign n14316 = n14315 ^ n14313 ^ 1'b0 ;
  assign n14317 = n14316 ^ n11685 ^ 1'b0 ;
  assign n14318 = n212 & ~n5150 ;
  assign n14319 = n11451 & n11703 ;
  assign n14320 = n14318 & n14319 ;
  assign n14321 = n3678 & ~n6701 ;
  assign n14322 = n14321 ^ n10185 ^ 1'b0 ;
  assign n14323 = ~n1953 & n3568 ;
  assign n14324 = n14323 ^ n6048 ^ 1'b0 ;
  assign n14325 = n6827 ^ n5082 ^ n4542 ;
  assign n14326 = n14324 & ~n14325 ;
  assign n14327 = n2967 & n14326 ;
  assign n14328 = n12077 & n12821 ;
  assign n14329 = n14328 ^ n741 ^ 1'b0 ;
  assign n14330 = n3107 & ~n6891 ;
  assign n14331 = n1265 | n8001 ;
  assign n14332 = n14331 ^ n1461 ^ 1'b0 ;
  assign n14333 = n89 & n14332 ;
  assign n14334 = n8522 & n10769 ;
  assign n14335 = n2994 & n5293 ;
  assign n14337 = ~n518 & n4072 ;
  assign n14336 = ~n13875 & n14116 ;
  assign n14338 = n14337 ^ n14336 ^ 1'b0 ;
  assign n14339 = n4051 | n12614 ;
  assign n14340 = n12996 | n14339 ;
  assign n14341 = n4583 & ~n8102 ;
  assign n14342 = n5870 & ~n14341 ;
  assign n14343 = n4556 & ~n7219 ;
  assign n14344 = ~n4670 & n14343 ;
  assign n14345 = n4564 ^ n2073 ^ 1'b0 ;
  assign n14346 = n2857 | n14345 ;
  assign n14347 = n872 | n14346 ;
  assign n14348 = n14343 ^ n4022 ^ 1'b0 ;
  assign n14349 = n14348 ^ n3270 ^ 1'b0 ;
  assign n14350 = n14349 ^ n400 ^ 1'b0 ;
  assign n14351 = n13666 ^ n8715 ^ n5473 ;
  assign n14352 = n14351 ^ n1009 ^ 1'b0 ;
  assign n14353 = ~n11189 & n11206 ;
  assign n14354 = n14353 ^ n10376 ^ 1'b0 ;
  assign n14356 = n2374 ^ n2309 ^ 1'b0 ;
  assign n14355 = n8214 & n12199 ;
  assign n14357 = n14356 ^ n14355 ^ 1'b0 ;
  assign n14358 = n8082 & ~n14357 ;
  assign n14359 = ~n5103 & n14358 ;
  assign n14360 = n14359 ^ n1403 ^ 1'b0 ;
  assign n14361 = n3906 & ~n10579 ;
  assign n14362 = ~n7715 & n14361 ;
  assign n14364 = n7695 & n11704 ;
  assign n14365 = n14364 ^ n12608 ^ n9908 ;
  assign n14363 = n2914 & n3727 ;
  assign n14366 = n14365 ^ n14363 ^ 1'b0 ;
  assign n14367 = ~n4188 & n9977 ;
  assign n14368 = n14367 ^ n8619 ^ 1'b0 ;
  assign n14369 = n5660 | n6557 ;
  assign n14370 = n8946 & n10846 ;
  assign n14371 = n3195 & n14370 ;
  assign n14372 = ( n2185 & ~n14369 ) | ( n2185 & n14371 ) | ( ~n14369 & n14371 ) ;
  assign n14373 = n9645 ^ n588 ^ 1'b0 ;
  assign n14374 = n6291 ^ n1560 ^ 1'b0 ;
  assign n14375 = n6314 & n10642 ;
  assign n14376 = n8482 ^ n6996 ^ 1'b0 ;
  assign n14377 = n1887 & ~n7598 ;
  assign n14378 = ~n14376 & n14377 ;
  assign n14379 = ( n5513 & n14375 ) | ( n5513 & n14378 ) | ( n14375 & n14378 ) ;
  assign n14380 = n2478 & ~n10979 ;
  assign n14381 = n3109 | n14380 ;
  assign n14382 = n14381 ^ n9380 ^ 1'b0 ;
  assign n14383 = n2693 ^ n2529 ^ 1'b0 ;
  assign n14384 = n1242 & ~n14383 ;
  assign n14385 = n3541 ^ n548 ^ n362 ;
  assign n14386 = ~n7282 & n14385 ;
  assign n14387 = n6455 | n7187 ;
  assign n14388 = n10407 ^ n8275 ^ n7861 ;
  assign n14389 = n14388 ^ n3331 ^ 1'b0 ;
  assign n14390 = n10240 ^ n7784 ^ 1'b0 ;
  assign n14391 = n7134 ^ n5080 ^ 1'b0 ;
  assign n14392 = ~n1700 & n14391 ;
  assign n14393 = n2596 & n13018 ;
  assign n14394 = n14393 ^ n10012 ^ 1'b0 ;
  assign n14395 = n5144 & n10156 ;
  assign n14396 = n14395 ^ n360 ^ 1'b0 ;
  assign n14397 = ~n5636 & n6017 ;
  assign n14398 = ~n8645 & n14397 ;
  assign n14400 = n2012 | n3140 ;
  assign n14399 = n5360 & n6011 ;
  assign n14401 = n14400 ^ n14399 ^ 1'b0 ;
  assign n14402 = ( n6259 & ~n8521 ) | ( n6259 & n14401 ) | ( ~n8521 & n14401 ) ;
  assign n14403 = ~n1868 & n8011 ;
  assign n14404 = n11352 ^ n6124 ^ 1'b0 ;
  assign n14405 = ( n1413 & n5132 ) | ( n1413 & n9812 ) | ( n5132 & n9812 ) ;
  assign n14408 = n1416 & n5237 ;
  assign n14409 = ~n12816 & n14408 ;
  assign n14406 = n2771 & n10083 ;
  assign n14407 = n11498 | n14406 ;
  assign n14410 = n14409 ^ n14407 ^ 1'b0 ;
  assign n14411 = n12906 | n12949 ;
  assign n14412 = n14411 ^ n3280 ^ 1'b0 ;
  assign n14413 = n6345 ^ n4070 ^ 1'b0 ;
  assign n14414 = n14413 ^ n12836 ^ 1'b0 ;
  assign n14415 = n6394 | n14414 ;
  assign n14416 = n14415 ^ n155 ^ 1'b0 ;
  assign n14417 = n13290 ^ n10007 ^ 1'b0 ;
  assign n14418 = ~n1986 & n13881 ;
  assign n14419 = n14418 ^ n5572 ^ 1'b0 ;
  assign n14420 = n1469 & n14419 ;
  assign n14421 = n5708 & n11722 ;
  assign n14422 = ~n6764 & n14421 ;
  assign n14423 = n4121 ^ n1691 ^ 1'b0 ;
  assign n14427 = n3206 & ~n5731 ;
  assign n14428 = n14427 ^ n9304 ^ 1'b0 ;
  assign n14429 = n3107 & ~n6126 ;
  assign n14430 = ~n5684 & n14429 ;
  assign n14431 = ~n14428 & n14430 ;
  assign n14424 = n1772 & n6442 ;
  assign n14425 = n2650 & n12484 ;
  assign n14426 = n14424 | n14425 ;
  assign n14432 = n14431 ^ n14426 ^ 1'b0 ;
  assign n14433 = n14423 & ~n14432 ;
  assign n14434 = n6585 & ~n9316 ;
  assign n14435 = n14434 ^ n8832 ^ n4267 ;
  assign n14436 = n12022 ^ n5750 ^ 1'b0 ;
  assign n14437 = n4913 & ~n14436 ;
  assign n14438 = n6891 | n14437 ;
  assign n14439 = n8365 ^ n1775 ^ n1212 ;
  assign n14440 = n14439 ^ n4849 ^ n224 ;
  assign n14441 = ~n7104 & n14440 ;
  assign n14442 = n3724 ^ n1009 ^ 1'b0 ;
  assign n14443 = n6534 ^ n2517 ^ 1'b0 ;
  assign n14444 = n11938 | n14443 ;
  assign n14445 = n10259 ^ n2751 ^ 1'b0 ;
  assign n14446 = n11586 | n14445 ;
  assign n14447 = n2513 ^ n2395 ^ 1'b0 ;
  assign n14448 = n14446 & n14447 ;
  assign n14449 = n13833 ^ n6996 ^ 1'b0 ;
  assign n14450 = n8410 & n14449 ;
  assign n14451 = n1413 & ~n2403 ;
  assign n14452 = ( n4199 & n4533 ) | ( n4199 & n6578 ) | ( n4533 & n6578 ) ;
  assign n14453 = n14452 ^ n10239 ^ 1'b0 ;
  assign n14455 = ~n2771 & n5368 ;
  assign n14454 = n2235 & ~n12647 ;
  assign n14456 = n14455 ^ n14454 ^ 1'b0 ;
  assign n14457 = n14453 | n14456 ;
  assign n14458 = n14457 ^ n12179 ^ 1'b0 ;
  assign n14459 = n7014 ^ n5648 ^ n1927 ;
  assign n14460 = n12414 ^ n5779 ^ 1'b0 ;
  assign n14461 = n13902 ^ n839 ^ 1'b0 ;
  assign n14462 = n9779 | n14461 ;
  assign n14463 = n6229 & n11935 ;
  assign n14464 = n14462 & n14463 ;
  assign n14465 = n6102 & n13728 ;
  assign n14466 = n5815 | n12736 ;
  assign n14467 = n7685 & ~n9802 ;
  assign n14468 = ~n8005 & n14467 ;
  assign n14469 = n14466 | n14468 ;
  assign n14470 = n4457 ^ n1622 ^ 1'b0 ;
  assign n14471 = n14470 ^ n4068 ^ 1'b0 ;
  assign n14472 = n8098 & n14471 ;
  assign n14473 = n14472 ^ n2628 ^ 1'b0 ;
  assign n14474 = n2709 & ~n7486 ;
  assign n14475 = ( n4429 & ~n5877 ) | ( n4429 & n14474 ) | ( ~n5877 & n14474 ) ;
  assign n14476 = n4317 | n7830 ;
  assign n14477 = n4884 & ~n14476 ;
  assign n14478 = n619 & ~n2612 ;
  assign n14479 = n14478 ^ n8287 ^ 1'b0 ;
  assign n14480 = ~n14477 & n14479 ;
  assign n14481 = n5868 ^ n2894 ^ 1'b0 ;
  assign n14482 = n14481 ^ n6669 ^ 1'b0 ;
  assign n14483 = n136 | n14482 ;
  assign n14484 = ~n13336 & n14483 ;
  assign n14485 = n13040 ^ n5305 ^ 1'b0 ;
  assign n14486 = n13196 ^ n12322 ^ n11878 ;
  assign n14487 = n7996 ^ n31 ^ 1'b0 ;
  assign n14488 = n12461 ^ n2048 ^ 1'b0 ;
  assign n14489 = n10218 & n14488 ;
  assign n14490 = n14489 ^ n13707 ^ 1'b0 ;
  assign n14491 = n14487 | n14490 ;
  assign n14492 = n9535 ^ n861 ^ 1'b0 ;
  assign n14493 = n14492 ^ n7836 ^ 1'b0 ;
  assign n14494 = n3254 ^ n752 ^ 1'b0 ;
  assign n14495 = n12496 | n14494 ;
  assign n14496 = n10857 ^ x2 ^ 1'b0 ;
  assign n14497 = ~n8805 & n14496 ;
  assign n14498 = ( n13127 & n14183 ) | ( n13127 & n14497 ) | ( n14183 & n14497 ) ;
  assign n14499 = n14400 ^ n7476 ^ 1'b0 ;
  assign n14500 = ~n2502 & n14499 ;
  assign n14501 = n3618 | n13973 ;
  assign n14502 = n7528 | n14501 ;
  assign n14505 = n12563 ^ n5073 ^ 1'b0 ;
  assign n14506 = n14505 ^ n5662 ^ 1'b0 ;
  assign n14503 = n8924 ^ n2024 ^ 1'b0 ;
  assign n14504 = n14503 ^ n13568 ^ 1'b0 ;
  assign n14507 = n14506 ^ n14504 ^ 1'b0 ;
  assign n14509 = n8768 ^ n669 ^ 1'b0 ;
  assign n14508 = n598 & ~n2981 ;
  assign n14510 = n14509 ^ n14508 ^ 1'b0 ;
  assign n14511 = n14510 ^ n4569 ^ 1'b0 ;
  assign n14512 = n4489 & ~n9875 ;
  assign n14513 = n4187 & ~n14512 ;
  assign n14514 = ~n8212 & n14513 ;
  assign n14515 = ~n311 & n1818 ;
  assign n14516 = n858 & n14515 ;
  assign n14517 = n14516 ^ n9508 ^ 1'b0 ;
  assign n14518 = n2309 & n14517 ;
  assign n14519 = n6766 | n14518 ;
  assign n14520 = n829 & ~n11509 ;
  assign n14521 = n7219 ^ n1539 ^ n774 ;
  assign n14522 = n6833 | n14521 ;
  assign n14523 = n10211 & ~n14522 ;
  assign n14524 = n14523 ^ n231 ^ 1'b0 ;
  assign n14525 = n14520 | n14524 ;
  assign n14526 = n10049 ^ n7516 ^ 1'b0 ;
  assign n14527 = n3811 & ~n14526 ;
  assign n14528 = n2771 | n5213 ;
  assign n14529 = n1434 & ~n14528 ;
  assign n14530 = n12919 ^ n4596 ^ 1'b0 ;
  assign n14531 = ~n10711 & n14530 ;
  assign n14532 = n1419 & n14531 ;
  assign n14533 = ~n3361 & n3949 ;
  assign n14534 = n14533 ^ n2236 ^ 1'b0 ;
  assign n14535 = n5872 & ~n14534 ;
  assign n14536 = n5508 & n14535 ;
  assign n14537 = n4506 ^ n3548 ^ n163 ;
  assign n14538 = n5348 ^ n540 ^ 1'b0 ;
  assign n14539 = n2455 & n6185 ;
  assign n14540 = n14539 ^ n11553 ^ 1'b0 ;
  assign n14541 = n2036 & n3706 ;
  assign n14542 = n14541 ^ n752 ^ 1'b0 ;
  assign n14543 = n209 & n13345 ;
  assign n14544 = ~n3633 & n4175 ;
  assign n14545 = ~n5319 & n13346 ;
  assign n14546 = n14544 & n14545 ;
  assign n14547 = n9373 ^ n1187 ^ 1'b0 ;
  assign n14548 = ~n12528 & n14547 ;
  assign n14549 = n2711 & n14548 ;
  assign n14550 = n14549 ^ n9608 ^ 1'b0 ;
  assign n14551 = ~n3133 & n8040 ;
  assign n14552 = n14551 ^ n8136 ^ 1'b0 ;
  assign n14554 = n302 & n812 ;
  assign n14555 = n8554 & n14554 ;
  assign n14553 = n1584 | n13751 ;
  assign n14556 = n14555 ^ n14553 ^ 1'b0 ;
  assign n14557 = n144 ^ n83 ^ 1'b0 ;
  assign n14558 = ~n4570 & n14557 ;
  assign n14559 = n14558 ^ n14423 ^ n2955 ;
  assign n14560 = ~n541 & n7735 ;
  assign n14561 = n1983 & ~n13879 ;
  assign n14562 = ~n106 & n10720 ;
  assign n14563 = n14562 ^ n1715 ^ 1'b0 ;
  assign n14564 = n14563 ^ n8730 ^ n5099 ;
  assign n14565 = n1391 ^ n51 ^ 1'b0 ;
  assign n14566 = n10209 & ~n14565 ;
  assign n14567 = ~n3033 & n14566 ;
  assign n14568 = n14564 & n14567 ;
  assign n14570 = ( ~n2427 & n4082 ) | ( ~n2427 & n5893 ) | ( n4082 & n5893 ) ;
  assign n14571 = ( ~n4104 & n9906 ) | ( ~n4104 & n11423 ) | ( n9906 & n11423 ) ;
  assign n14572 = n2566 ^ n911 ^ 1'b0 ;
  assign n14573 = n8478 | n14572 ;
  assign n14574 = n14571 | n14573 ;
  assign n14575 = n14570 & ~n14574 ;
  assign n14569 = n12814 ^ n5167 ^ n2872 ;
  assign n14576 = n14575 ^ n14569 ^ 1'b0 ;
  assign n14577 = ~n9688 & n14576 ;
  assign n14578 = n11511 | n14577 ;
  assign n14579 = n13695 ^ n6670 ^ 1'b0 ;
  assign n14580 = n8663 & ~n12105 ;
  assign n14581 = n5490 & ~n9688 ;
  assign n14582 = ~n5145 & n14581 ;
  assign n14583 = ~n1694 & n4596 ;
  assign n14584 = ( n88 & n1420 ) | ( n88 & ~n11185 ) | ( n1420 & ~n11185 ) ;
  assign n14585 = n14583 & ~n14584 ;
  assign n14586 = ~n11668 & n14585 ;
  assign n14587 = n14586 ^ n6305 ^ n3993 ;
  assign n14588 = n4267 & ~n14587 ;
  assign n14589 = n14588 ^ n1422 ^ 1'b0 ;
  assign n14590 = n11726 ^ n669 ^ 1'b0 ;
  assign n14591 = n14589 | n14590 ;
  assign n14592 = n4066 & ~n14591 ;
  assign n14593 = n14592 ^ n3744 ^ 1'b0 ;
  assign n14594 = n12402 ^ n214 ^ 1'b0 ;
  assign n14595 = ~n13961 & n14594 ;
  assign n14596 = n11285 ^ n8863 ^ 1'b0 ;
  assign n14597 = n2732 ^ n2631 ^ 1'b0 ;
  assign n14598 = n11189 ^ n2958 ^ 1'b0 ;
  assign n14599 = n14598 ^ n8217 ^ 1'b0 ;
  assign n14600 = ~n12625 & n14599 ;
  assign n14601 = n10404 ^ n6618 ^ 1'b0 ;
  assign n14602 = ~n1580 & n5647 ;
  assign n14603 = n11056 & ~n14602 ;
  assign n14604 = n5628 & n8163 ;
  assign n14605 = n14604 ^ n2773 ^ 1'b0 ;
  assign n14606 = n1935 | n14605 ;
  assign n14607 = n8758 & ~n14606 ;
  assign n14608 = n9057 ^ n2859 ^ 1'b0 ;
  assign n14609 = n11838 ^ n3418 ^ 1'b0 ;
  assign n14610 = n8106 | n14609 ;
  assign n14611 = n14610 ^ n4760 ^ 1'b0 ;
  assign n14612 = n8022 ^ n1828 ^ 1'b0 ;
  assign n14613 = ~n3212 & n12301 ;
  assign n14614 = n694 & ~n13873 ;
  assign n14615 = n1922 | n8402 ;
  assign n14616 = n10348 & ~n14615 ;
  assign n14617 = n5493 & ~n7964 ;
  assign n14618 = n14617 ^ n1920 ^ 1'b0 ;
  assign n14619 = n5733 & ~n14618 ;
  assign n14620 = n6771 & n14619 ;
  assign n14621 = n489 & n8301 ;
  assign n14622 = n2451 & n14621 ;
  assign n14623 = n14622 ^ n9465 ^ 1'b0 ;
  assign n14624 = n440 & n14623 ;
  assign n14628 = n5016 | n5073 ;
  assign n14629 = n5073 & ~n14628 ;
  assign n14625 = n2686 & n3500 ;
  assign n14626 = ~n2686 & n14625 ;
  assign n14627 = n2664 | n14626 ;
  assign n14630 = n14629 ^ n14627 ^ 1'b0 ;
  assign n14631 = n1861 | n6138 ;
  assign n14632 = n1861 & ~n14631 ;
  assign n14633 = n14630 | n14632 ;
  assign n14634 = n14630 & ~n14633 ;
  assign n14635 = n7354 ^ n5441 ^ n1439 ;
  assign n14636 = n14635 ^ n10778 ^ 1'b0 ;
  assign n14637 = n6353 & ~n10209 ;
  assign n14638 = n3944 ^ n2327 ^ 1'b0 ;
  assign n14639 = n4263 & ~n14638 ;
  assign n14640 = n12563 & ~n14639 ;
  assign n14641 = n14637 & ~n14640 ;
  assign n14642 = n5431 & n14641 ;
  assign n14643 = n14642 ^ n6818 ^ 1'b0 ;
  assign n14644 = ~n5730 & n14643 ;
  assign n14645 = n8766 & ~n11277 ;
  assign n14646 = n14645 ^ n2046 ^ 1'b0 ;
  assign n14647 = n14646 ^ n723 ^ 1'b0 ;
  assign n14648 = ~n889 & n14647 ;
  assign n14649 = n13751 ^ n4848 ^ 1'b0 ;
  assign n14650 = n6777 ^ n1252 ^ 1'b0 ;
  assign n14651 = n14650 ^ n9769 ^ 1'b0 ;
  assign n14652 = n6711 & n14651 ;
  assign n14653 = ( n4037 & n6281 ) | ( n4037 & n6948 ) | ( n6281 & n6948 ) ;
  assign n14656 = ( n2618 & ~n3736 ) | ( n2618 & n7046 ) | ( ~n3736 & n7046 ) ;
  assign n14654 = n7147 ^ n3349 ^ 1'b0 ;
  assign n14655 = ~n7011 & n14654 ;
  assign n14657 = n14656 ^ n14655 ^ 1'b0 ;
  assign n14658 = n5744 & n8144 ;
  assign n14659 = n6259 ^ n5240 ^ 1'b0 ;
  assign n14660 = n14658 & ~n14659 ;
  assign n14661 = n14660 ^ n4545 ^ 1'b0 ;
  assign n14662 = n2549 & ~n14661 ;
  assign n14663 = n13198 ^ n4512 ^ 1'b0 ;
  assign n14664 = n2647 | n14663 ;
  assign n14665 = n14664 ^ n11547 ^ 1'b0 ;
  assign n14669 = ~n2128 & n12985 ;
  assign n14666 = n551 | n3227 ;
  assign n14667 = n14666 ^ n6904 ^ 1'b0 ;
  assign n14668 = n14667 ^ n8919 ^ 1'b0 ;
  assign n14670 = n14669 ^ n14668 ^ 1'b0 ;
  assign n14671 = n3915 ^ n2086 ^ 1'b0 ;
  assign n14672 = n133 | n14671 ;
  assign n14673 = ( n1010 & n7102 ) | ( n1010 & n14672 ) | ( n7102 & n14672 ) ;
  assign n14674 = n4651 & n14673 ;
  assign n14675 = n2915 | n11339 ;
  assign n14676 = n6773 & ~n7707 ;
  assign n14677 = n752 | n6455 ;
  assign n14678 = n14677 ^ n11327 ^ 1'b0 ;
  assign n14679 = n5725 & n14678 ;
  assign n14680 = n856 & ~n1675 ;
  assign n14681 = ~n2716 & n14680 ;
  assign n14682 = ~n4168 & n14681 ;
  assign n14683 = n9738 | n12011 ;
  assign n14684 = n14682 | n14683 ;
  assign n14685 = n1295 & ~n3417 ;
  assign n14686 = ( n6093 & n6193 ) | ( n6093 & n11199 ) | ( n6193 & n11199 ) ;
  assign n14687 = n12719 ^ n8416 ^ 1'b0 ;
  assign n14688 = n14687 ^ n7167 ^ 1'b0 ;
  assign n14689 = n12344 | n14688 ;
  assign n14690 = n6663 ^ n915 ^ 1'b0 ;
  assign n14691 = n6527 & n14690 ;
  assign n14692 = n14691 ^ n5598 ^ 1'b0 ;
  assign n14693 = n12233 & n14692 ;
  assign n14694 = n5212 & ~n10873 ;
  assign n14695 = n14694 ^ n4838 ^ 1'b0 ;
  assign n14696 = n13059 & ~n14695 ;
  assign n14697 = n1845 | n4367 ;
  assign n14698 = n209 & n513 ;
  assign n14699 = ~n209 & n14698 ;
  assign n14700 = n746 & n14699 ;
  assign n14701 = ~n14699 & n14700 ;
  assign n14702 = n3854 & n14701 ;
  assign n14703 = n3726 & ~n14702 ;
  assign n14704 = n7130 & n14471 ;
  assign n14705 = ~n14471 & n14704 ;
  assign n14706 = ( n298 & n14703 ) | ( n298 & ~n14705 ) | ( n14703 & ~n14705 ) ;
  assign n14707 = n4921 & n14164 ;
  assign n14708 = ~n12665 & n14707 ;
  assign n14709 = n314 | n4789 ;
  assign n14710 = x0 | n14709 ;
  assign n14711 = ~n5697 & n14710 ;
  assign n14712 = n10542 & n14711 ;
  assign n14714 = n3406 ^ n2219 ^ 1'b0 ;
  assign n14715 = n466 & ~n6799 ;
  assign n14716 = ~n14714 & n14715 ;
  assign n14713 = n9712 ^ n5402 ^ n3889 ;
  assign n14717 = n14716 ^ n14713 ^ 1'b0 ;
  assign n14718 = n4789 | n14717 ;
  assign n14719 = n2656 & ~n14718 ;
  assign n14720 = n14712 & n14719 ;
  assign n14721 = n7782 | n12466 ;
  assign n14722 = n14721 ^ n3323 ^ 1'b0 ;
  assign n14723 = ~n5699 & n13279 ;
  assign n14724 = n5258 & n14723 ;
  assign n14729 = n4576 & ~n10023 ;
  assign n14727 = n968 & n1980 ;
  assign n14728 = n3539 | n14727 ;
  assign n14725 = n8304 ^ n7763 ^ 1'b0 ;
  assign n14726 = n1643 | n14725 ;
  assign n14730 = n14729 ^ n14728 ^ n14726 ;
  assign n14731 = n4307 | n5382 ;
  assign n14733 = n8643 & ~n9408 ;
  assign n14734 = ~n2876 & n14733 ;
  assign n14732 = ~n2811 & n11758 ;
  assign n14735 = n14734 ^ n14732 ^ 1'b0 ;
  assign n14736 = ( n637 & n714 ) | ( n637 & ~n1337 ) | ( n714 & ~n1337 ) ;
  assign n14737 = n6854 & n14736 ;
  assign n14738 = n8406 ^ n5172 ^ n226 ;
  assign n14739 = ( n9844 & n14737 ) | ( n9844 & ~n14738 ) | ( n14737 & ~n14738 ) ;
  assign n14740 = n2494 & ~n5393 ;
  assign n14741 = n752 | n10342 ;
  assign n14742 = n2767 | n3886 ;
  assign n14743 = n1024 & ~n14742 ;
  assign n14744 = n651 & n3480 ;
  assign n14745 = n4449 | n14744 ;
  assign n14746 = n14743 & ~n14745 ;
  assign n14747 = n7676 & ~n13200 ;
  assign n14748 = ~x11 & n14747 ;
  assign n14749 = n6954 ^ n6543 ^ n6273 ;
  assign n14750 = ~n219 & n14749 ;
  assign n14751 = n7150 ^ n5369 ^ 1'b0 ;
  assign n14752 = n5901 & n14751 ;
  assign n14753 = ~n14750 & n14752 ;
  assign n14754 = n5464 & ~n8545 ;
  assign n14756 = n1285 & ~n1599 ;
  assign n14757 = ~n477 & n14756 ;
  assign n14758 = n2045 | n14757 ;
  assign n14759 = n14758 ^ n5940 ^ 1'b0 ;
  assign n14755 = n4977 & n6562 ;
  assign n14760 = n14759 ^ n14755 ^ 1'b0 ;
  assign n14761 = n5360 ^ n1878 ^ 1'b0 ;
  assign n14762 = n1504 & ~n12819 ;
  assign n14763 = ~n493 & n14762 ;
  assign n14764 = n12142 ^ n5911 ^ 1'b0 ;
  assign n14765 = ~n8173 & n14764 ;
  assign n14766 = ( n5057 & n7367 ) | ( n5057 & n8887 ) | ( n7367 & n8887 ) ;
  assign n14767 = ~n6827 & n14766 ;
  assign n14768 = ~n1087 & n14767 ;
  assign n14769 = n1196 | n14768 ;
  assign n14770 = n14769 ^ n2474 ^ 1'b0 ;
  assign n14771 = n1714 | n8141 ;
  assign n14772 = n5093 & ~n14771 ;
  assign n14773 = n3279 ^ n846 ^ 1'b0 ;
  assign n14774 = ( ~n8008 & n8647 ) | ( ~n8008 & n14773 ) | ( n8647 & n14773 ) ;
  assign n14775 = n1157 & ~n8269 ;
  assign n14776 = n1138 | n14775 ;
  assign n14777 = n746 & ~n9322 ;
  assign n14778 = n14777 ^ n1816 ^ 1'b0 ;
  assign n14779 = n296 | n14778 ;
  assign n14780 = n14779 ^ n11308 ^ 1'b0 ;
  assign n14781 = n6528 | n14780 ;
  assign n14782 = n14781 ^ n5114 ^ 1'b0 ;
  assign n14783 = n3019 ^ n2367 ^ 1'b0 ;
  assign n14784 = n1363 & ~n14783 ;
  assign n14785 = n1063 & n1750 ;
  assign n14786 = ~n831 & n14785 ;
  assign n14787 = ~n14784 & n14786 ;
  assign n14788 = n3539 ^ n260 ^ 1'b0 ;
  assign n14789 = ~n14787 & n14788 ;
  assign n14790 = n14789 ^ n14712 ^ 1'b0 ;
  assign n14791 = n5906 & ~n14381 ;
  assign n14792 = n5936 ^ n4645 ^ n181 ;
  assign n14793 = n9686 ^ n6162 ^ 1'b0 ;
  assign n14794 = n502 & n14793 ;
  assign n14795 = ~n4774 & n14794 ;
  assign n14796 = n1673 & ~n3594 ;
  assign n14797 = n2217 | n8827 ;
  assign n14798 = n43 | n14797 ;
  assign n14799 = n14798 ^ n5478 ^ 1'b0 ;
  assign n14800 = n6980 & n14799 ;
  assign n14801 = ~n14119 & n14800 ;
  assign n14802 = n14801 ^ n11469 ^ 1'b0 ;
  assign n14803 = n4343 ^ n2146 ^ 1'b0 ;
  assign n14804 = n14802 & n14803 ;
  assign n14805 = n2231 ^ n163 ^ 1'b0 ;
  assign n14806 = n12312 ^ n2358 ^ 1'b0 ;
  assign n14807 = n8663 & ~n14806 ;
  assign n14808 = ~n3744 & n14807 ;
  assign n14809 = n2507 & n3476 ;
  assign n14810 = n14809 ^ n10484 ^ 1'b0 ;
  assign n14811 = n11692 ^ n7293 ^ 1'b0 ;
  assign n14812 = n8858 & ~n14811 ;
  assign n14813 = n9049 ^ n5815 ^ 1'b0 ;
  assign n14814 = n14813 ^ n9743 ^ 1'b0 ;
  assign n14815 = n1566 | n14814 ;
  assign n14816 = ~n3845 & n11685 ;
  assign n14817 = ~n488 & n14816 ;
  assign n14818 = n7293 ^ n4001 ^ 1'b0 ;
  assign n14819 = n2351 & n13147 ;
  assign n14820 = n13251 ^ n8101 ^ 1'b0 ;
  assign n14821 = n4113 & n4933 ;
  assign n14822 = n11827 ^ n9248 ^ 1'b0 ;
  assign n14823 = n14821 & n14822 ;
  assign n14824 = ~n14820 & n14823 ;
  assign n14825 = n10854 ^ n571 ^ 1'b0 ;
  assign n14826 = n13532 ^ n11812 ^ 1'b0 ;
  assign n14827 = ~n14667 & n14826 ;
  assign n14828 = n12246 ^ n7825 ^ 1'b0 ;
  assign n14829 = n14828 ^ n2438 ^ 1'b0 ;
  assign n14831 = n2014 | n8652 ;
  assign n14830 = n5184 | n6632 ;
  assign n14832 = n14831 ^ n14830 ^ 1'b0 ;
  assign n14833 = n6526 ^ n1269 ^ 1'b0 ;
  assign n14834 = n253 & n2398 ;
  assign n14835 = ~n14833 & n14834 ;
  assign n14836 = n6020 & ~n14835 ;
  assign n14837 = n3611 & n14836 ;
  assign n14838 = n445 & ~n8258 ;
  assign n14839 = ( ~n2785 & n2943 ) | ( ~n2785 & n14838 ) | ( n2943 & n14838 ) ;
  assign n14840 = n1714 | n6059 ;
  assign n14841 = n3361 & ~n14840 ;
  assign n14842 = n14841 ^ n787 ^ 1'b0 ;
  assign n14843 = n220 & ~n590 ;
  assign n14844 = n778 & n14843 ;
  assign n14845 = ~n1576 & n14844 ;
  assign n14846 = n4313 ^ n2966 ^ 1'b0 ;
  assign n14847 = n12221 ^ n3299 ^ 1'b0 ;
  assign n14848 = ( ~n489 & n7588 ) | ( ~n489 & n14847 ) | ( n7588 & n14847 ) ;
  assign n14849 = n8986 ^ n2558 ^ 1'b0 ;
  assign n14850 = n14849 ^ n3476 ^ 1'b0 ;
  assign n14851 = n14848 & ~n14850 ;
  assign n14852 = n14851 ^ n2116 ^ 1'b0 ;
  assign n14853 = ~n14602 & n14852 ;
  assign n14854 = ~n1196 & n10857 ;
  assign n14855 = ~n764 & n14854 ;
  assign n14856 = n12261 & ~n14855 ;
  assign n14857 = n9341 ^ n1808 ^ 1'b0 ;
  assign n14862 = n6411 ^ n3909 ^ 1'b0 ;
  assign n14863 = n7657 | n14862 ;
  assign n14864 = n14863 ^ n5779 ^ 1'b0 ;
  assign n14865 = n5680 & n14864 ;
  assign n14866 = n9631 & ~n14865 ;
  assign n14858 = n3756 ^ n489 ^ 1'b0 ;
  assign n14859 = n14858 ^ n4303 ^ 1'b0 ;
  assign n14860 = ~n5480 & n14859 ;
  assign n14861 = ( n3796 & ~n11576 ) | ( n3796 & n14860 ) | ( ~n11576 & n14860 ) ;
  assign n14867 = n14866 ^ n14861 ^ 1'b0 ;
  assign n14868 = n1589 & n3635 ;
  assign n14869 = n7140 | n14868 ;
  assign n14870 = n14869 ^ n10809 ^ 1'b0 ;
  assign n14871 = n7960 & ~n10510 ;
  assign n14872 = ~n3734 & n14871 ;
  assign n14873 = n10853 | n13424 ;
  assign n14875 = ~n3647 & n9779 ;
  assign n14874 = n3881 & ~n11474 ;
  assign n14876 = n14875 ^ n14874 ^ 1'b0 ;
  assign n14877 = n14876 ^ n13320 ^ n10099 ;
  assign n14878 = ( n3612 & ~n5652 ) | ( n3612 & n14275 ) | ( ~n5652 & n14275 ) ;
  assign n14879 = n14878 ^ n8860 ^ 1'b0 ;
  assign n14880 = n2228 | n14879 ;
  assign n14882 = ~n295 & n1031 ;
  assign n14883 = n14882 ^ n1650 ^ 1'b0 ;
  assign n14884 = n13351 | n14883 ;
  assign n14881 = n12299 & n12780 ;
  assign n14885 = n14884 ^ n14881 ^ 1'b0 ;
  assign n14887 = ~n865 & n9873 ;
  assign n14886 = n7174 & ~n8402 ;
  assign n14888 = n14887 ^ n14886 ^ 1'b0 ;
  assign n14889 = ~n9319 & n14888 ;
  assign n14890 = n8506 ^ n8001 ^ 1'b0 ;
  assign n14891 = n35 & n8500 ;
  assign n14892 = n8894 & ~n11876 ;
  assign n14893 = n14138 & ~n14892 ;
  assign n14894 = ~n7335 & n14893 ;
  assign n14895 = n3971 ^ n3441 ^ 1'b0 ;
  assign n14896 = n4980 & n13726 ;
  assign n14897 = n14895 & n14896 ;
  assign n14898 = n14894 & n14897 ;
  assign n14899 = ~n11242 & n14898 ;
  assign n14900 = n1056 & n9741 ;
  assign n14901 = ~n7569 & n14900 ;
  assign n14902 = n14901 ^ n4169 ^ 1'b0 ;
  assign n14903 = n2698 & n11189 ;
  assign n14904 = ~n5349 & n14903 ;
  assign n14905 = n5022 | n12661 ;
  assign n14906 = n14905 ^ n13991 ^ 1'b0 ;
  assign n14907 = n11584 & ~n14906 ;
  assign n14908 = n83 & ~n12561 ;
  assign n14909 = n14908 ^ n8628 ^ 1'b0 ;
  assign n14910 = n6796 & n14909 ;
  assign n14911 = n13675 ^ n7480 ^ 1'b0 ;
  assign n14912 = n1073 & ~n12046 ;
  assign n14913 = ~n1591 & n14912 ;
  assign n14914 = n14911 & ~n14913 ;
  assign n14915 = n14914 ^ n7293 ^ 1'b0 ;
  assign n14916 = n6330 ^ n3400 ^ 1'b0 ;
  assign n14917 = n7300 ^ n3231 ^ 1'b0 ;
  assign n14918 = n3132 | n14917 ;
  assign n14919 = n12896 ^ n940 ^ 1'b0 ;
  assign n14920 = n7478 & ~n14919 ;
  assign n14921 = n5649 & n6067 ;
  assign n14922 = n403 & n14921 ;
  assign n14923 = ~n398 & n4857 ;
  assign n14924 = n1582 | n1592 ;
  assign n14925 = n14924 ^ n5161 ^ 1'b0 ;
  assign n14926 = n2747 | n4496 ;
  assign n14927 = n7464 & n12202 ;
  assign n14928 = n11214 & ~n13832 ;
  assign n14929 = n10340 | n13223 ;
  assign n14930 = n7137 & ~n14929 ;
  assign n14931 = ~n2480 & n5185 ;
  assign n14932 = n2108 & n5995 ;
  assign n14933 = n1781 | n3713 ;
  assign n14934 = ~n7152 & n7955 ;
  assign n14936 = n2705 ^ n510 ^ 1'b0 ;
  assign n14937 = n1191 & n14936 ;
  assign n14935 = n764 & n4837 ;
  assign n14938 = n14937 ^ n14935 ^ 1'b0 ;
  assign n14939 = n14938 ^ n10364 ^ 1'b0 ;
  assign n14940 = n5467 | n14939 ;
  assign n14941 = n43 | n14940 ;
  assign n14942 = n4776 ^ n40 ^ 1'b0 ;
  assign n14943 = n7171 | n14942 ;
  assign n14944 = n7708 | n14943 ;
  assign n14945 = n1430 & ~n2848 ;
  assign n14946 = ( n1050 & ~n4293 ) | ( n1050 & n13429 ) | ( ~n4293 & n13429 ) ;
  assign n14947 = n14945 & ~n14946 ;
  assign n14948 = n1946 & n4246 ;
  assign n14949 = ( n4117 & ~n4389 ) | ( n4117 & n14948 ) | ( ~n4389 & n14948 ) ;
  assign n14950 = n1588 & n14949 ;
  assign n14951 = n2812 & n2833 ;
  assign n14952 = ~n3416 & n14951 ;
  assign n14953 = n5082 ^ n4264 ^ 1'b0 ;
  assign n14954 = n9195 ^ n7933 ^ 1'b0 ;
  assign n14955 = n839 | n11628 ;
  assign n14956 = n3182 | n5743 ;
  assign n14957 = n5682 & ~n14956 ;
  assign n14958 = n12480 ^ n7105 ^ 1'b0 ;
  assign n14959 = ~n1237 & n4203 ;
  assign n14960 = n12597 ^ n4005 ^ 1'b0 ;
  assign n14961 = ~n2114 & n14960 ;
  assign n14962 = ~n3091 & n4780 ;
  assign n14963 = ~n1157 & n1700 ;
  assign n14964 = ~n4753 & n14963 ;
  assign n14965 = n7061 & n14964 ;
  assign n14966 = ~n14962 & n14965 ;
  assign n14967 = n3760 | n6040 ;
  assign n14968 = n3892 | n14967 ;
  assign n14969 = n14966 & n14968 ;
  assign n14970 = n12646 ^ n5234 ^ 1'b0 ;
  assign n14971 = ~n3113 & n14970 ;
  assign n14972 = ~n3106 & n14971 ;
  assign n14973 = n3985 & n14972 ;
  assign n14974 = n4504 ^ n3957 ^ 1'b0 ;
  assign n14975 = ~n1506 & n14974 ;
  assign n14976 = n14975 ^ n5897 ^ n5660 ;
  assign n14977 = n251 | n423 ;
  assign n14978 = ~n1199 & n14977 ;
  assign n14979 = n9574 & n14978 ;
  assign n14982 = n5256 & ~n10221 ;
  assign n14983 = n2146 & n14982 ;
  assign n14980 = n5348 ^ n831 ^ 1'b0 ;
  assign n14981 = n9247 & ~n14980 ;
  assign n14984 = n14983 ^ n14981 ^ 1'b0 ;
  assign n14985 = n5202 | n14984 ;
  assign n14986 = ~n1832 & n6258 ;
  assign n14987 = n4535 & n14986 ;
  assign n14988 = n14987 ^ n14419 ^ 1'b0 ;
  assign n14989 = n14988 ^ n12816 ^ 1'b0 ;
  assign n14990 = n8029 | n9436 ;
  assign n14991 = n14990 ^ n3864 ^ 1'b0 ;
  assign n14992 = n9499 | n14487 ;
  assign n14993 = ~n8643 & n14992 ;
  assign n14994 = ~x7 & n14993 ;
  assign n14995 = n1134 | n14668 ;
  assign n14996 = n1006 & ~n14995 ;
  assign n14997 = n2252 & n14996 ;
  assign n14998 = n5151 & n7730 ;
  assign n14999 = n14616 & n14998 ;
  assign n15000 = n8506 ^ n4038 ^ 1'b0 ;
  assign n15001 = n6598 & n15000 ;
  assign n15002 = n13871 ^ n4903 ^ 1'b0 ;
  assign n15003 = n8659 | n9868 ;
  assign n15004 = n10951 ^ n1049 ^ 1'b0 ;
  assign n15005 = n2313 & n15004 ;
  assign n15006 = n14749 ^ n11278 ^ 1'b0 ;
  assign n15007 = n9128 | n15006 ;
  assign n15008 = n3044 | n15007 ;
  assign n15009 = n1889 & n12850 ;
  assign n15010 = ~n4038 & n4463 ;
  assign n15011 = ( ~n1354 & n5010 ) | ( ~n1354 & n15010 ) | ( n5010 & n15010 ) ;
  assign n15012 = n5547 & ~n15011 ;
  assign n15013 = n15012 ^ n1434 ^ 1'b0 ;
  assign n15014 = n5513 & ~n12496 ;
  assign n15015 = n15014 ^ n3909 ^ 1'b0 ;
  assign n15016 = n3054 ^ n1839 ^ 1'b0 ;
  assign n15017 = n5095 & ~n13065 ;
  assign n15018 = ~n7652 & n15017 ;
  assign n15019 = n845 | n15018 ;
  assign n15020 = ~n2363 & n14813 ;
  assign n15021 = n7278 & ~n8541 ;
  assign n15022 = n6806 & n15021 ;
  assign n15023 = n3033 & n8625 ;
  assign n15024 = n10259 & ~n15023 ;
  assign n15025 = n302 & n15024 ;
  assign n15026 = ~n3392 & n4729 ;
  assign n15027 = n15026 ^ n7285 ^ 1'b0 ;
  assign n15028 = n3110 ^ n2517 ^ 1'b0 ;
  assign n15029 = n2576 & ~n15028 ;
  assign n15030 = n7523 ^ n6700 ^ 1'b0 ;
  assign n15031 = n1553 & ~n6410 ;
  assign n15032 = n8365 ^ n7549 ^ 1'b0 ;
  assign n15033 = n5267 ^ n3674 ^ 1'b0 ;
  assign n15034 = n4474 & n15033 ;
  assign n15035 = n15034 ^ n5632 ^ 1'b0 ;
  assign n15036 = n2779 ^ n1121 ^ 1'b0 ;
  assign n15037 = n15035 | n15036 ;
  assign n15038 = n8909 | n15037 ;
  assign n15040 = n4622 & ~n7349 ;
  assign n15041 = ~n1987 & n15040 ;
  assign n15042 = n302 & n15041 ;
  assign n15039 = n10365 & n11699 ;
  assign n15043 = n15042 ^ n15039 ^ 1'b0 ;
  assign n15044 = n6398 | n8024 ;
  assign n15045 = n15044 ^ n6083 ^ 1'b0 ;
  assign n15046 = n10239 ^ n7861 ^ 1'b0 ;
  assign n15047 = ~n2773 & n15046 ;
  assign n15048 = n15045 & n15047 ;
  assign n15049 = n9002 ^ n316 ^ 1'b0 ;
  assign n15050 = n15049 ^ n14923 ^ 1'b0 ;
  assign n15051 = n6250 & ~n7437 ;
  assign n15052 = n1973 & ~n15051 ;
  assign n15053 = n2028 ^ n1728 ^ 1'b0 ;
  assign n15054 = n3646 | n5418 ;
  assign n15055 = n13881 ^ n7792 ^ 1'b0 ;
  assign n15056 = n1141 & n2771 ;
  assign n15061 = n3612 ^ n40 ^ 1'b0 ;
  assign n15062 = ( n640 & n7936 ) | ( n640 & ~n15061 ) | ( n7936 & ~n15061 ) ;
  assign n15057 = n177 | n288 ;
  assign n15058 = n15057 ^ n904 ^ 1'b0 ;
  assign n15059 = n15058 ^ n1409 ^ 1'b0 ;
  assign n15060 = n4388 & ~n15059 ;
  assign n15063 = n15062 ^ n15060 ^ 1'b0 ;
  assign n15064 = n11909 | n15063 ;
  assign n15065 = n5837 & n11668 ;
  assign n15066 = n15065 ^ n10702 ^ 1'b0 ;
  assign n15067 = ~n5641 & n15066 ;
  assign n15068 = n5064 | n15067 ;
  assign n15069 = n13708 ^ n10554 ^ 1'b0 ;
  assign n15070 = ( n6981 & n15068 ) | ( n6981 & ~n15069 ) | ( n15068 & ~n15069 ) ;
  assign n15071 = n4576 & n12789 ;
  assign n15072 = n1371 & ~n12468 ;
  assign n15073 = n15072 ^ n5168 ^ 1'b0 ;
  assign n15074 = n8784 | n15073 ;
  assign n15075 = n244 & ~n15074 ;
  assign n15076 = n7768 ^ n219 ^ 1'b0 ;
  assign n15077 = n15076 ^ n6585 ^ 1'b0 ;
  assign n15078 = n1983 & n15077 ;
  assign n15079 = n10238 ^ n3618 ^ 1'b0 ;
  assign n15080 = n12173 | n15079 ;
  assign n15081 = n15080 ^ n403 ^ 1'b0 ;
  assign n15083 = n4077 ^ n493 ^ 1'b0 ;
  assign n15082 = n2670 & ~n11209 ;
  assign n15084 = n15083 ^ n15082 ^ 1'b0 ;
  assign n15085 = ~n1694 & n3403 ;
  assign n15086 = n15085 ^ n5685 ^ 1'b0 ;
  assign n15087 = n492 & ~n4714 ;
  assign n15088 = n3213 ^ n86 ^ 1'b0 ;
  assign n15089 = n15088 ^ n3335 ^ 1'b0 ;
  assign n15090 = n7388 | n15089 ;
  assign n15091 = n403 & n2505 ;
  assign n15092 = n15091 ^ n7019 ^ 1'b0 ;
  assign n15093 = n910 & n4007 ;
  assign n15094 = n15093 ^ n2073 ^ 1'b0 ;
  assign n15095 = ~n6638 & n15094 ;
  assign n15096 = n15095 ^ n3864 ^ 1'b0 ;
  assign n15097 = n15096 ^ n2548 ^ 1'b0 ;
  assign n15098 = n5517 & n15097 ;
  assign n15099 = n7277 ^ n3592 ^ 1'b0 ;
  assign n15100 = n6430 | n6804 ;
  assign n15101 = n15100 ^ n1877 ^ 1'b0 ;
  assign n15102 = n8719 | n15101 ;
  assign n15103 = ( ~n3683 & n12588 ) | ( ~n3683 & n15102 ) | ( n12588 & n15102 ) ;
  assign n15104 = n8960 | n15103 ;
  assign n15105 = n15104 ^ n8073 ^ 1'b0 ;
  assign n15106 = n5900 ^ n582 ^ 1'b0 ;
  assign n15107 = n6098 ^ n745 ^ 1'b0 ;
  assign n15108 = n5458 & n15107 ;
  assign n15109 = n4040 ^ n3867 ^ 1'b0 ;
  assign n15110 = n10084 & n15109 ;
  assign n15111 = ~n12344 & n15110 ;
  assign n15112 = n5321 & n15111 ;
  assign n15113 = n5814 ^ n3671 ^ n600 ;
  assign n15114 = n15113 ^ n11755 ^ 1'b0 ;
  assign n15115 = n15114 ^ n10152 ^ n2721 ;
  assign n15116 = n12788 & ~n12889 ;
  assign n15117 = n546 & n15116 ;
  assign n15121 = n5290 ^ n1918 ^ 1'b0 ;
  assign n15122 = n10454 & n15121 ;
  assign n15118 = n2195 | n6834 ;
  assign n15119 = n2610 & ~n15118 ;
  assign n15120 = n15119 ^ n5151 ^ 1'b0 ;
  assign n15123 = n15122 ^ n15120 ^ 1'b0 ;
  assign n15124 = n3382 ^ n3127 ^ 1'b0 ;
  assign n15125 = n12353 | n15124 ;
  assign n15126 = n12628 & ~n15125 ;
  assign n15127 = ( ~n7371 & n13233 ) | ( ~n7371 & n13912 ) | ( n13233 & n13912 ) ;
  assign n15128 = n3379 & n11221 ;
  assign n15129 = n12375 & ~n15128 ;
  assign n15130 = n251 | n7686 ;
  assign n15131 = n9151 & ~n10654 ;
  assign n15132 = ~n15130 & n15131 ;
  assign n15133 = n6498 ^ n1563 ^ 1'b0 ;
  assign n15135 = n7342 ^ n3792 ^ n1009 ;
  assign n15134 = ~n723 & n1257 ;
  assign n15136 = n15135 ^ n15134 ^ 1'b0 ;
  assign n15143 = n267 & ~n1454 ;
  assign n15144 = n15143 ^ n2061 ^ 1'b0 ;
  assign n15137 = ~n150 & n625 ;
  assign n15138 = ~n479 & n15137 ;
  assign n15139 = ~n12118 & n15138 ;
  assign n15140 = n15139 ^ n3035 ^ 1'b0 ;
  assign n15141 = n15140 ^ n13138 ^ 1'b0 ;
  assign n15142 = ~n1095 & n15141 ;
  assign n15145 = n15144 ^ n15142 ^ 1'b0 ;
  assign n15146 = n261 | n1794 ;
  assign n15147 = n3968 & ~n15146 ;
  assign n15148 = n15147 ^ n5766 ^ 1'b0 ;
  assign n15149 = n2384 & n15148 ;
  assign n15150 = n15149 ^ n10761 ^ 1'b0 ;
  assign n15152 = n1212 ^ n1000 ^ 1'b0 ;
  assign n15153 = ~n5557 & n15152 ;
  assign n15154 = n4084 & n9314 ;
  assign n15155 = ~n15153 & n15154 ;
  assign n15151 = n4747 ^ n51 ^ 1'b0 ;
  assign n15156 = n15155 ^ n15151 ^ 1'b0 ;
  assign n15157 = n7983 | n15156 ;
  assign n15158 = ~n3886 & n13354 ;
  assign n15159 = n7015 & n15158 ;
  assign n15162 = n9779 ^ n5982 ^ 1'b0 ;
  assign n15163 = n10910 | n15162 ;
  assign n15160 = n772 | n10448 ;
  assign n15161 = n7846 & ~n15160 ;
  assign n15164 = n15163 ^ n15161 ^ 1'b0 ;
  assign n15165 = n2356 | n4014 ;
  assign n15166 = n15165 ^ n2460 ^ 1'b0 ;
  assign n15167 = n15166 ^ n7372 ^ 1'b0 ;
  assign n15168 = n10430 | n15167 ;
  assign n15169 = n3054 | n5378 ;
  assign n15170 = n1900 & ~n15169 ;
  assign n15171 = ~n4538 & n4764 ;
  assign n15172 = n7015 & ~n15171 ;
  assign n15173 = n7675 | n15172 ;
  assign n15174 = n14213 | n15173 ;
  assign n15175 = n12028 ^ n3537 ^ n2390 ;
  assign n15176 = n8526 | n15175 ;
  assign n15177 = n15176 ^ n7989 ^ 1'b0 ;
  assign n15178 = n1288 & ~n15177 ;
  assign n15179 = ~n9488 & n10420 ;
  assign n15180 = ~n8232 & n15179 ;
  assign n15181 = n4167 ^ n2419 ^ 1'b0 ;
  assign n15182 = n3572 & ~n15181 ;
  assign n15183 = n15182 ^ n623 ^ 1'b0 ;
  assign n15184 = n121 & n4058 ;
  assign n15185 = n492 & ~n15184 ;
  assign n15186 = n15185 ^ n3323 ^ 1'b0 ;
  assign n15187 = n4704 & ~n15186 ;
  assign n15188 = n8937 ^ n7342 ^ n56 ;
  assign n15189 = n12392 ^ n3747 ^ 1'b0 ;
  assign n15190 = n9941 ^ n154 ^ 1'b0 ;
  assign n15191 = ( n2799 & n8735 ) | ( n2799 & n11160 ) | ( n8735 & n11160 ) ;
  assign n15192 = n2120 | n12904 ;
  assign n15193 = n11037 ^ n9210 ^ 1'b0 ;
  assign n15194 = n15168 ^ n7389 ^ 1'b0 ;
  assign n15195 = n11584 & ~n15194 ;
  assign n15196 = n8723 ^ n3112 ^ 1'b0 ;
  assign n15197 = ~n749 & n7881 ;
  assign n15198 = n15196 & n15197 ;
  assign n15199 = n9476 ^ n7846 ^ 1'b0 ;
  assign n15200 = ~n15198 & n15199 ;
  assign n15201 = n2588 | n4333 ;
  assign n15202 = n7844 ^ n1868 ^ 1'b0 ;
  assign n15203 = n15201 & n15202 ;
  assign n15204 = n15203 ^ n5288 ^ 1'b0 ;
  assign n15205 = n1267 | n15204 ;
  assign n15206 = ~n9110 & n15205 ;
  assign n15207 = n857 & n3694 ;
  assign n15208 = n15207 ^ n4621 ^ 1'b0 ;
  assign n15209 = n13274 | n15208 ;
  assign n15210 = n3958 | n8758 ;
  assign n15211 = n8005 & n12843 ;
  assign n15212 = n15211 ^ n33 ^ 1'b0 ;
  assign n15213 = n8324 | n15212 ;
  assign n15214 = n15213 ^ n3384 ^ n801 ;
  assign n15215 = n13061 ^ n12173 ^ 1'b0 ;
  assign n15216 = n5470 ^ n4485 ^ 1'b0 ;
  assign n15217 = n10973 & ~n15216 ;
  assign n15218 = n15215 & ~n15217 ;
  assign n15219 = n4226 ^ n495 ^ 1'b0 ;
  assign n15220 = n4832 & ~n15219 ;
  assign n15221 = n7423 & ~n10388 ;
  assign n15222 = n8023 ^ n4637 ^ 1'b0 ;
  assign n15223 = n2874 & ~n10980 ;
  assign n15224 = n6797 & n15223 ;
  assign n15225 = n4558 & ~n15224 ;
  assign n15226 = n15225 ^ n13827 ^ 1'b0 ;
  assign n15227 = n15119 ^ n1714 ^ 1'b0 ;
  assign n15228 = ~n12618 & n15227 ;
  assign n15229 = n1584 & ~n10189 ;
  assign n15230 = n14736 & n15229 ;
  assign n15234 = n7337 & ~n12487 ;
  assign n15231 = ~n593 & n3630 ;
  assign n15232 = n15231 ^ n10691 ^ 1'b0 ;
  assign n15233 = n6156 & ~n15232 ;
  assign n15235 = n15234 ^ n15233 ^ 1'b0 ;
  assign n15236 = n1897 | n5293 ;
  assign n15237 = n263 & ~n15236 ;
  assign n15238 = ~n13697 & n15237 ;
  assign n15239 = n211 | n908 ;
  assign n15240 = n15239 ^ n3445 ^ n165 ;
  assign n15241 = n4802 ^ n4082 ^ 1'b0 ;
  assign n15242 = n6898 ^ n2626 ^ 1'b0 ;
  assign n15243 = n884 & ~n15242 ;
  assign n15244 = ( ~n1741 & n15241 ) | ( ~n1741 & n15243 ) | ( n15241 & n15243 ) ;
  assign n15245 = n9056 | n14884 ;
  assign n15246 = n7316 & ~n15245 ;
  assign n15247 = n11211 ^ n2343 ^ 1'b0 ;
  assign n15248 = n14315 & ~n15247 ;
  assign n15249 = ~n10119 & n15248 ;
  assign n15250 = n15249 ^ n9049 ^ 1'b0 ;
  assign n15251 = n3564 & ~n4159 ;
  assign n15252 = ~n10616 & n15251 ;
  assign n15253 = n15252 ^ n6831 ^ 1'b0 ;
  assign n15254 = n3430 ^ n1693 ^ 1'b0 ;
  assign n15255 = n11098 ^ n311 ^ 1'b0 ;
  assign n15256 = n15254 & n15255 ;
  assign n15257 = n3064 | n7375 ;
  assign n15258 = n2964 ^ n150 ^ 1'b0 ;
  assign n15259 = n1991 & n15258 ;
  assign n15260 = n4248 ^ n3201 ^ n2427 ;
  assign n15261 = n9680 ^ n924 ^ 1'b0 ;
  assign n15262 = n12584 ^ n5058 ^ 1'b0 ;
  assign n15263 = ~n7384 & n8497 ;
  assign n15264 = n8842 | n10846 ;
  assign n15265 = n15264 ^ n4121 ^ 1'b0 ;
  assign n15266 = n12413 ^ n3974 ^ 1'b0 ;
  assign n15267 = n4845 & n15266 ;
  assign n15268 = ~n5286 & n10676 ;
  assign n15269 = n13458 ^ n3933 ^ 1'b0 ;
  assign n15270 = n12638 & ~n15269 ;
  assign n15271 = n1369 & n12023 ;
  assign n15272 = ~n431 & n1271 ;
  assign n15273 = n15272 ^ n10917 ^ 1'b0 ;
  assign n15274 = ~n12041 & n15273 ;
  assign n15275 = n1429 | n7546 ;
  assign n15276 = n5344 & ~n5695 ;
  assign n15277 = n15276 ^ n2172 ^ 1'b0 ;
  assign n15278 = n8879 & n15277 ;
  assign n15279 = ~n3686 & n4808 ;
  assign n15280 = n2733 | n15279 ;
  assign n15281 = n12402 & ~n15280 ;
  assign n15282 = n5584 ^ x11 ^ 1'b0 ;
  assign n15283 = ~n7119 & n15282 ;
  assign n15284 = n11768 & ~n12262 ;
  assign n15285 = ~n15283 & n15284 ;
  assign n15286 = n6131 | n15285 ;
  assign n15287 = n13524 & ~n15286 ;
  assign n15288 = n915 ^ n536 ^ 1'b0 ;
  assign n15289 = n1431 & n15288 ;
  assign n15290 = n5658 & ~n15289 ;
  assign n15291 = ~n3017 & n3386 ;
  assign n15292 = n2317 ^ n229 ^ 1'b0 ;
  assign n15293 = n6878 & ~n15292 ;
  assign n15294 = n14847 | n15293 ;
  assign n15295 = n8576 | n15294 ;
  assign n15296 = n10884 & n15295 ;
  assign n15297 = n15296 ^ n4745 ^ 1'b0 ;
  assign n15298 = n12487 | n15297 ;
  assign n15299 = ~n5641 & n11681 ;
  assign n15300 = n14511 ^ n12899 ^ n6189 ;
  assign n15301 = n9540 ^ n6771 ^ 1'b0 ;
  assign n15302 = ~n874 & n15301 ;
  assign n15303 = n12503 ^ n5663 ^ 1'b0 ;
  assign n15304 = n1576 & ~n15303 ;
  assign n15305 = n749 & n13087 ;
  assign n15306 = ~n15304 & n15305 ;
  assign n15307 = ~n15302 & n15306 ;
  assign n15308 = n1848 | n2812 ;
  assign n15309 = n3280 & ~n15308 ;
  assign n15310 = ~n6979 & n15309 ;
  assign n15311 = n2859 | n3560 ;
  assign n15312 = n15311 ^ n1510 ^ 1'b0 ;
  assign n15313 = n3054 & n15312 ;
  assign n15314 = n5254 & ~n7466 ;
  assign n15315 = n1609 & n15314 ;
  assign n15316 = n15315 ^ n5914 ^ 1'b0 ;
  assign n15317 = n2152 ^ n150 ^ 1'b0 ;
  assign n15318 = n15317 ^ n11572 ^ n835 ;
  assign n15319 = n15147 ^ n6729 ^ 1'b0 ;
  assign n15320 = ~n10716 & n15319 ;
  assign n15321 = ~n160 & n15320 ;
  assign n15322 = n12324 ^ n8971 ^ 1'b0 ;
  assign n15323 = n1930 ^ n1269 ^ 1'b0 ;
  assign n15324 = n229 | n15323 ;
  assign n15325 = n3592 & n6764 ;
  assign n15326 = ~n15324 & n15325 ;
  assign n15327 = n7442 ^ n2382 ^ 1'b0 ;
  assign n15328 = n214 & ~n15327 ;
  assign n15329 = ~n699 & n2045 ;
  assign n15330 = n15329 ^ n13462 ^ 1'b0 ;
  assign n15331 = n15330 ^ n1662 ^ 1'b0 ;
  assign n15332 = n8002 ^ n5633 ^ 1'b0 ;
  assign n15334 = n3555 ^ n582 ^ 1'b0 ;
  assign n15333 = n4738 & ~n7877 ;
  assign n15335 = n15334 ^ n15333 ^ 1'b0 ;
  assign n15336 = n15332 | n15335 ;
  assign n15337 = n4731 ^ n4448 ^ 1'b0 ;
  assign n15338 = n6613 ^ n4993 ^ 1'b0 ;
  assign n15339 = n7562 | n10389 ;
  assign n15340 = n12464 ^ n4816 ^ 1'b0 ;
  assign n15341 = n8106 & n15340 ;
  assign n15342 = n1445 ^ n1157 ^ 1'b0 ;
  assign n15343 = ( ~n1862 & n6701 ) | ( ~n1862 & n7843 ) | ( n6701 & n7843 ) ;
  assign n15344 = n15343 ^ n3958 ^ n2867 ;
  assign n15346 = n2886 & ~n3052 ;
  assign n15345 = ~n3594 & n5823 ;
  assign n15347 = n15346 ^ n15345 ^ 1'b0 ;
  assign n15350 = n1199 & n1814 ;
  assign n15351 = n15350 ^ x7 ^ 1'b0 ;
  assign n15348 = n20 & ~n11183 ;
  assign n15349 = n8661 & ~n15348 ;
  assign n15352 = n15351 ^ n15349 ^ 1'b0 ;
  assign n15353 = n12998 ^ n12407 ^ 1'b0 ;
  assign n15354 = n10119 | n15353 ;
  assign n15355 = n12965 ^ n8181 ^ 1'b0 ;
  assign n15356 = n15355 ^ n15263 ^ 1'b0 ;
  assign n15362 = n5658 & n6385 ;
  assign n15363 = n2020 & n15362 ;
  assign n15357 = n2808 & n4553 ;
  assign n15358 = n15357 ^ n1363 ^ 1'b0 ;
  assign n15359 = n5885 | n15358 ;
  assign n15360 = n13677 ^ n2351 ^ n1744 ;
  assign n15361 = ~n15359 & n15360 ;
  assign n15364 = n15363 ^ n15361 ^ 1'b0 ;
  assign n15365 = n1016 & ~n2408 ;
  assign n15369 = n8448 ^ n2517 ^ 1'b0 ;
  assign n15370 = n4871 & ~n15369 ;
  assign n15367 = n6556 ^ n121 ^ 1'b0 ;
  assign n15366 = n2652 & n6762 ;
  assign n15368 = n15367 ^ n15366 ^ 1'b0 ;
  assign n15371 = n15370 ^ n15368 ^ n1342 ;
  assign n15372 = ~n132 & n1943 ;
  assign n15373 = n5480 & n12765 ;
  assign n15374 = ~n15372 & n15373 ;
  assign n15376 = n10616 & ~n10736 ;
  assign n15375 = ~n1613 & n9122 ;
  assign n15377 = n15376 ^ n15375 ^ 1'b0 ;
  assign n15379 = ~n218 & n6122 ;
  assign n15380 = ~n5022 & n15379 ;
  assign n15381 = n15380 ^ n7665 ^ n2260 ;
  assign n15382 = n15381 ^ n5730 ^ 1'b0 ;
  assign n15383 = n7799 & n15382 ;
  assign n15384 = n15383 ^ n6103 ^ 1'b0 ;
  assign n15385 = ~n12576 & n15384 ;
  assign n15378 = ~n5320 & n8332 ;
  assign n15386 = n15385 ^ n15378 ^ 1'b0 ;
  assign n15387 = n3035 | n15386 ;
  assign n15388 = n2576 & n4677 ;
  assign n15389 = ~n3778 & n15388 ;
  assign n15390 = n1929 & n15389 ;
  assign n15391 = n5288 & n15390 ;
  assign n15392 = ~n11570 & n15391 ;
  assign n15393 = n2008 ^ n1548 ^ 1'b0 ;
  assign n15394 = n7008 ^ n2847 ^ n835 ;
  assign n15395 = ~n2679 & n9594 ;
  assign n15396 = n15394 & n15395 ;
  assign n15397 = n1004 ^ n131 ^ 1'b0 ;
  assign n15398 = ~n3992 & n15397 ;
  assign n15399 = n15398 ^ n14058 ^ 1'b0 ;
  assign n15400 = n4384 & n8904 ;
  assign n15401 = n4837 | n15400 ;
  assign n15402 = n2351 & ~n8268 ;
  assign n15403 = ~n6757 & n15402 ;
  assign n15404 = n3158 & n5767 ;
  assign n15405 = n5285 | n8730 ;
  assign n15406 = n4685 | n15405 ;
  assign n15407 = n15406 ^ n7107 ^ n2587 ;
  assign n15408 = n3450 & n13992 ;
  assign n15409 = n15408 ^ n4546 ^ 1'b0 ;
  assign n15410 = n3830 & ~n7280 ;
  assign n15411 = n15410 ^ n4199 ^ 1'b0 ;
  assign n15412 = n3522 & ~n7635 ;
  assign n15413 = n5030 ^ n2753 ^ 1'b0 ;
  assign n15414 = n4038 & n13393 ;
  assign n15415 = ~n15413 & n15414 ;
  assign n15416 = ( n694 & n8633 ) | ( n694 & ~n14639 ) | ( n8633 & ~n14639 ) ;
  assign n15417 = n15415 | n15416 ;
  assign n15418 = n9309 ^ n8987 ^ n2478 ;
  assign n15419 = n2170 | n15418 ;
  assign n15420 = n15419 ^ n11162 ^ 1'b0 ;
  assign n15421 = ( n2079 & ~n2460 ) | ( n2079 & n2924 ) | ( ~n2460 & n2924 ) ;
  assign n15422 = n445 | n15421 ;
  assign n15423 = n12718 | n15422 ;
  assign n15424 = n15423 ^ n4544 ^ 1'b0 ;
  assign n15425 = n3959 | n7153 ;
  assign n15426 = n15425 ^ n13342 ^ 1'b0 ;
  assign n15427 = n15426 ^ n15002 ^ 1'b0 ;
  assign n15428 = n5139 & ~n15201 ;
  assign n15429 = n15428 ^ n3777 ^ 1'b0 ;
  assign n15430 = n4719 ^ n1267 ^ 1'b0 ;
  assign n15431 = n5116 | n15430 ;
  assign n15432 = n9276 ^ n3258 ^ 1'b0 ;
  assign n15433 = ~n15431 & n15432 ;
  assign n15434 = n6876 & ~n8390 ;
  assign n15435 = n15434 ^ n2780 ^ 1'b0 ;
  assign n15436 = n8256 ^ n4350 ^ 1'b0 ;
  assign n15437 = n431 & ~n910 ;
  assign n15438 = n14353 ^ n214 ^ 1'b0 ;
  assign n15440 = n9366 | n9580 ;
  assign n15441 = n8402 ^ n2547 ^ 1'b0 ;
  assign n15442 = n15440 & ~n15441 ;
  assign n15439 = ~n5143 & n8685 ;
  assign n15443 = n15442 ^ n15439 ^ 1'b0 ;
  assign n15444 = n6911 ^ n1929 ^ n1574 ;
  assign n15445 = n7054 & ~n11105 ;
  assign n15446 = n15445 ^ n5274 ^ 1'b0 ;
  assign n15447 = n4875 | n15446 ;
  assign n15448 = n8157 ^ n27 ^ 1'b0 ;
  assign n15449 = ~n6189 & n10542 ;
  assign n15450 = n7048 ^ n5579 ^ 1'b0 ;
  assign n15451 = n15449 & ~n15450 ;
  assign n15453 = n5178 | n8312 ;
  assign n15454 = n968 | n15453 ;
  assign n15452 = n11922 & n12230 ;
  assign n15455 = n15454 ^ n15452 ^ 1'b0 ;
  assign n15456 = n4720 & n5673 ;
  assign n15457 = n15456 ^ n212 ^ 1'b0 ;
  assign n15458 = n1462 & n4980 ;
  assign n15459 = n4916 & n15458 ;
  assign n15460 = ~n1235 & n15459 ;
  assign n15461 = n15460 ^ n7467 ^ 1'b0 ;
  assign n15462 = n15457 | n15461 ;
  assign n15463 = n7771 ^ n5984 ^ 1'b0 ;
  assign n15464 = n8667 & n15463 ;
  assign n15465 = ~n564 & n15464 ;
  assign n15466 = n1743 | n12701 ;
  assign n15467 = n2574 | n15466 ;
  assign n15468 = n9724 & ~n15467 ;
  assign n15470 = n7066 ^ n2899 ^ 1'b0 ;
  assign n15469 = n1726 & n5463 ;
  assign n15471 = n15470 ^ n15469 ^ 1'b0 ;
  assign n15472 = n3361 & n3983 ;
  assign n15473 = n1454 & ~n15472 ;
  assign n15474 = n1385 ^ n560 ^ 1'b0 ;
  assign n15475 = ~n11523 & n15474 ;
  assign n15476 = n15475 ^ n6618 ^ 1'b0 ;
  assign n15477 = n7624 & n15476 ;
  assign n15478 = n4540 ^ n987 ^ n86 ;
  assign n15479 = n15477 | n15478 ;
  assign n15480 = n13589 ^ n2529 ^ 1'b0 ;
  assign n15481 = n2121 & n15480 ;
  assign n15482 = n5791 | n14539 ;
  assign n15483 = n1853 | n15482 ;
  assign n15484 = n4573 & n13165 ;
  assign n15485 = n914 | n1391 ;
  assign n15487 = n5378 ^ n577 ^ 1'b0 ;
  assign n15486 = n110 | n2923 ;
  assign n15488 = n15487 ^ n15486 ^ 1'b0 ;
  assign n15489 = n11911 ^ n3293 ^ 1'b0 ;
  assign n15491 = n6498 ^ n6352 ^ n770 ;
  assign n15490 = n489 | n5554 ;
  assign n15492 = n15491 ^ n15490 ^ 1'b0 ;
  assign n15493 = n15492 ^ n1791 ^ 1'b0 ;
  assign n15494 = n1016 & ~n3439 ;
  assign n15495 = n15494 ^ n14948 ^ 1'b0 ;
  assign n15496 = n3597 & ~n7282 ;
  assign n15497 = ~n9665 & n15496 ;
  assign n15498 = n6240 ^ n3682 ^ 1'b0 ;
  assign n15499 = ~n6566 & n15498 ;
  assign n15500 = n1631 & ~n1962 ;
  assign n15501 = n9912 & n15500 ;
  assign n15502 = n11563 ^ n8354 ^ 1'b0 ;
  assign n15503 = ~n2723 & n7739 ;
  assign n15504 = n5422 & n15503 ;
  assign n15505 = n344 & n15504 ;
  assign n15506 = n15505 ^ n7529 ^ 1'b0 ;
  assign n15507 = n8790 ^ n890 ^ 1'b0 ;
  assign n15508 = n2340 & ~n6895 ;
  assign n15509 = n4561 | n12109 ;
  assign n15510 = n11356 ^ n6018 ^ 1'b0 ;
  assign n15511 = ~n2403 & n15510 ;
  assign n15512 = n15511 ^ n6328 ^ 1'b0 ;
  assign n15513 = n5306 & n5949 ;
  assign n15514 = n12799 ^ n10816 ^ 1'b0 ;
  assign n15515 = n15514 ^ n4814 ^ n2465 ;
  assign n15518 = n91 & ~n2349 ;
  assign n15519 = n15518 ^ n4302 ^ 1'b0 ;
  assign n15516 = ~n1994 & n7047 ;
  assign n15517 = n11367 | n15516 ;
  assign n15520 = n15519 ^ n15517 ^ 1'b0 ;
  assign n15521 = n7346 ^ n6219 ^ n584 ;
  assign n15522 = n13327 ^ n11968 ^ n4881 ;
  assign n15523 = n3623 ^ n1711 ^ 1'b0 ;
  assign n15524 = n15523 ^ n10280 ^ 1'b0 ;
  assign n15525 = n12819 ^ n3536 ^ 1'b0 ;
  assign n15526 = n8700 ^ n6762 ^ 1'b0 ;
  assign n15527 = n6126 ^ n2406 ^ n2185 ;
  assign n15528 = n10853 | n11616 ;
  assign n15529 = n15527 & n15528 ;
  assign n15530 = n11920 ^ n8805 ^ 1'b0 ;
  assign n15531 = n3833 & ~n15530 ;
  assign n15532 = n2232 & n15531 ;
  assign n15533 = ( ~n395 & n15529 ) | ( ~n395 & n15532 ) | ( n15529 & n15532 ) ;
  assign n15536 = n7249 ^ n3334 ^ 1'b0 ;
  assign n15537 = ~n6949 & n15536 ;
  assign n15534 = n2113 & n5046 ;
  assign n15535 = n15171 & n15534 ;
  assign n15538 = n15537 ^ n15535 ^ n4347 ;
  assign n15539 = n1907 | n15538 ;
  assign n15540 = n6553 | n9844 ;
  assign n15541 = n7516 | n15540 ;
  assign n15542 = n1387 & n13323 ;
  assign n15543 = n15541 & n15542 ;
  assign n15544 = ~n14415 & n15543 ;
  assign n15545 = ~n4852 & n8053 ;
  assign n15546 = n1603 & n4301 ;
  assign n15547 = n6343 | n15546 ;
  assign n15548 = n3317 & n6601 ;
  assign n15549 = n1546 & n6773 ;
  assign n15550 = ~n14805 & n15549 ;
  assign n15555 = n5079 & n5493 ;
  assign n15556 = n2996 & n15555 ;
  assign n15551 = n4259 | n8385 ;
  assign n15552 = n15551 ^ n6605 ^ 1'b0 ;
  assign n15553 = n4377 & ~n15552 ;
  assign n15554 = n14371 & n15553 ;
  assign n15557 = n15556 ^ n15554 ^ n8354 ;
  assign n15558 = ~n570 & n3392 ;
  assign n15559 = n13609 ^ n13070 ^ n2240 ;
  assign n15560 = n3177 & n13507 ;
  assign n15561 = n15560 ^ n466 ^ 1'b0 ;
  assign n15562 = n15559 & n15561 ;
  assign n15563 = n2324 ^ n1223 ^ 1'b0 ;
  assign n15564 = n8165 & n15563 ;
  assign n15565 = n15564 ^ n5382 ^ 1'b0 ;
  assign n15566 = n2781 ^ n1582 ^ 1'b0 ;
  assign n15567 = n15565 & n15566 ;
  assign n15568 = n2419 & n3012 ;
  assign n15569 = n15568 ^ n5427 ^ 1'b0 ;
  assign n15570 = n15569 ^ n4147 ^ 1'b0 ;
  assign n15571 = n3674 | n15570 ;
  assign n15572 = n1510 ^ n1147 ^ 1'b0 ;
  assign n15573 = n10287 & ~n15572 ;
  assign n15574 = n15573 ^ n6036 ^ 1'b0 ;
  assign n15575 = ( n485 & n2157 ) | ( n485 & n15574 ) | ( n2157 & n15574 ) ;
  assign n15583 = n1169 & n2986 ;
  assign n15578 = n2091 & ~n3710 ;
  assign n15579 = n5319 | n15578 ;
  assign n15580 = n15579 ^ n6552 ^ 1'b0 ;
  assign n15581 = ~n910 & n15580 ;
  assign n15576 = ~n3852 & n9738 ;
  assign n15577 = n3936 | n15576 ;
  assign n15582 = n15581 ^ n15577 ^ 1'b0 ;
  assign n15584 = n15583 ^ n15582 ^ 1'b0 ;
  assign n15585 = n12050 ^ n1363 ^ 1'b0 ;
  assign n15586 = ~n2355 & n4754 ;
  assign n15587 = n11664 ^ n3967 ^ n1887 ;
  assign n15588 = n1346 & n15587 ;
  assign n15589 = n8330 | n14564 ;
  assign n15590 = n15589 ^ n3597 ^ 1'b0 ;
  assign n15591 = n557 & ~n4040 ;
  assign n15592 = ~n15590 & n15591 ;
  assign n15593 = n846 | n15592 ;
  assign n15594 = n7893 & ~n15593 ;
  assign n15596 = n205 | n347 ;
  assign n15597 = n9139 | n15596 ;
  assign n15595 = n1055 & ~n14884 ;
  assign n15598 = n15597 ^ n15595 ^ 1'b0 ;
  assign n15599 = n8142 | n9748 ;
  assign n15600 = n533 | n2358 ;
  assign n15601 = n5736 & n8933 ;
  assign n15602 = ~n15600 & n15601 ;
  assign n15603 = n2775 | n15602 ;
  assign n15604 = n3449 | n3746 ;
  assign n15605 = n15604 ^ n5541 ^ 1'b0 ;
  assign n15606 = ( ~n7718 & n14720 ) | ( ~n7718 & n15605 ) | ( n14720 & n15605 ) ;
  assign n15607 = n8568 ^ n4369 ^ 1'b0 ;
  assign n15608 = n8541 | n15607 ;
  assign n15609 = n15608 ^ n10596 ^ 1'b0 ;
  assign n15610 = n9471 ^ n4000 ^ 1'b0 ;
  assign n15611 = n5600 | n15610 ;
  assign n15612 = n6631 & ~n8005 ;
  assign n15613 = n4104 & n15612 ;
  assign n15614 = n13927 & n15613 ;
  assign n15615 = n10929 | n14094 ;
  assign n15616 = n15615 ^ n8465 ^ 1'b0 ;
  assign n15617 = n14828 ^ n10749 ^ 1'b0 ;
  assign n15618 = ( n5842 & ~n13909 ) | ( n5842 & n15415 ) | ( ~n13909 & n15415 ) ;
  assign n15619 = n3535 & ~n12759 ;
  assign n15620 = n1024 & n8210 ;
  assign n15621 = n3393 & n7018 ;
  assign n15622 = n15621 ^ n855 ^ 1'b0 ;
  assign n15623 = ( ~n3386 & n11968 ) | ( ~n3386 & n14450 ) | ( n11968 & n14450 ) ;
  assign n15624 = n13540 ^ n5302 ^ 1'b0 ;
  assign n15625 = n699 | n15624 ;
  assign n15626 = n15624 & ~n15625 ;
  assign n15627 = n10637 | n15626 ;
  assign n15628 = n6540 | n15627 ;
  assign n15629 = ~n4586 & n15628 ;
  assign n15630 = n15629 ^ n10087 ^ 1'b0 ;
  assign n15631 = n7375 & ~n15630 ;
  assign n15632 = n682 & ~n15631 ;
  assign n15634 = n1534 & ~n2525 ;
  assign n15633 = n1205 | n3891 ;
  assign n15635 = n15634 ^ n15633 ^ n12616 ;
  assign n15636 = n15632 & n15635 ;
  assign n15637 = n10166 & n11318 ;
  assign n15638 = n15637 ^ n5531 ^ 1'b0 ;
  assign n15639 = n15128 ^ n13806 ^ 1'b0 ;
  assign n15640 = n1745 & n4244 ;
  assign n15641 = n5403 & n15640 ;
  assign n15642 = n10687 ^ n6262 ^ 1'b0 ;
  assign n15643 = ~n15641 & n15642 ;
  assign n15644 = n15643 ^ n15404 ^ 1'b0 ;
  assign n15645 = n3140 & ~n4468 ;
  assign n15646 = ~n3450 & n15645 ;
  assign n15647 = ~n3913 & n9772 ;
  assign n15648 = n15647 ^ n8089 ^ 1'b0 ;
  assign n15649 = n9171 ^ n7516 ^ 1'b0 ;
  assign n15650 = n6206 & n9608 ;
  assign n15657 = n6574 ^ n376 ^ 1'b0 ;
  assign n15651 = n875 & ~n3467 ;
  assign n15652 = n130 & ~n311 ;
  assign n15653 = ~n15651 & n15652 ;
  assign n15654 = n6122 & ~n15653 ;
  assign n15655 = n451 & n15654 ;
  assign n15656 = n3903 & ~n15655 ;
  assign n15658 = n15657 ^ n15656 ^ 1'b0 ;
  assign n15659 = ~n15650 & n15658 ;
  assign n15660 = n12497 ^ n5741 ^ n1424 ;
  assign n15661 = n11688 & ~n15660 ;
  assign n15662 = n15554 ^ n6136 ^ 1'b0 ;
  assign n15663 = n9426 ^ n1434 ^ n465 ;
  assign n15664 = n4077 & ~n15663 ;
  assign n15665 = n3135 ^ n1249 ^ 1'b0 ;
  assign n15666 = n1750 ^ n1508 ^ 1'b0 ;
  assign n15667 = ~n4893 & n15666 ;
  assign n15670 = n9416 ^ n2498 ^ 1'b0 ;
  assign n15671 = n4263 & ~n15670 ;
  assign n15669 = ~n533 & n12526 ;
  assign n15672 = n15671 ^ n15669 ^ 1'b0 ;
  assign n15668 = n3935 | n7067 ;
  assign n15673 = n15672 ^ n15668 ^ 1'b0 ;
  assign n15674 = n15667 & ~n15673 ;
  assign n15675 = ~n7722 & n10269 ;
  assign n15676 = n3060 & n8570 ;
  assign n15677 = ~n796 & n4751 ;
  assign n15678 = n15676 & n15677 ;
  assign n15679 = n5250 | n15678 ;
  assign n15680 = n15675 | n15679 ;
  assign n15681 = ( ~n1510 & n11649 ) | ( ~n1510 & n15680 ) | ( n11649 & n15680 ) ;
  assign n15685 = n316 | n4725 ;
  assign n15686 = n15685 ^ n5727 ^ n3995 ;
  assign n15682 = n2290 & n5297 ;
  assign n15683 = n15682 ^ n13264 ^ 1'b0 ;
  assign n15684 = n5302 | n15683 ;
  assign n15687 = n15686 ^ n15684 ^ 1'b0 ;
  assign n15688 = ~n4473 & n13242 ;
  assign n15689 = n15688 ^ n2954 ^ 1'b0 ;
  assign n15690 = ~n2458 & n15467 ;
  assign n15691 = ~n1004 & n8534 ;
  assign n15692 = ( ~n192 & n9331 ) | ( ~n192 & n15691 ) | ( n9331 & n15691 ) ;
  assign n15693 = n703 & n15388 ;
  assign n15694 = n7659 & n15693 ;
  assign n15695 = n5027 & ~n15694 ;
  assign n15696 = n4030 & ~n15695 ;
  assign n15697 = ~n5847 & n15696 ;
  assign n15698 = n15692 & ~n15697 ;
  assign n15699 = n712 ^ n144 ^ 1'b0 ;
  assign n15700 = n7485 & n15699 ;
  assign n15701 = n1907 & n8831 ;
  assign n15702 = n15701 ^ n11683 ^ 1'b0 ;
  assign n15703 = n13402 ^ n10754 ^ n4317 ;
  assign n15704 = n9177 ^ n4969 ^ n4350 ;
  assign n15705 = n8414 & ~n15704 ;
  assign n15706 = n5410 ^ n3437 ^ 1'b0 ;
  assign n15707 = ~n1006 & n15706 ;
  assign n15708 = n15707 ^ n12231 ^ 1'b0 ;
  assign n15709 = n1154 & ~n14052 ;
  assign n15710 = n15709 ^ n15231 ^ 1'b0 ;
  assign n15711 = n15210 ^ n7647 ^ 1'b0 ;
  assign n15712 = n2445 & ~n15711 ;
  assign n15713 = n1276 & n2067 ;
  assign n15714 = n7593 & n15713 ;
  assign n15715 = n15714 ^ n2946 ^ 1'b0 ;
  assign n15716 = n8494 ^ n8412 ^ 1'b0 ;
  assign n15717 = n4085 & ~n11816 ;
  assign n15718 = n15717 ^ n6533 ^ 1'b0 ;
  assign n15719 = n2517 | n8000 ;
  assign n15720 = n3703 ^ n3428 ^ 1'b0 ;
  assign n15721 = n1329 & n15720 ;
  assign n15722 = n1387 | n12602 ;
  assign n15723 = n15721 & n15722 ;
  assign n15724 = n15653 ^ n2097 ^ 1'b0 ;
  assign n15725 = ~n3904 & n15724 ;
  assign n15726 = ~n7682 & n11234 ;
  assign n15727 = n15726 ^ n11722 ^ 1'b0 ;
  assign n15728 = n13079 & ~n15727 ;
  assign n15729 = n7785 ^ n1147 ^ 1'b0 ;
  assign n15730 = ~n4301 & n15729 ;
  assign n15731 = n5697 | n13668 ;
  assign n15732 = n12641 & ~n15731 ;
  assign n15733 = n15730 & ~n15732 ;
  assign n15734 = ~n15730 & n15733 ;
  assign n15735 = n4881 | n8630 ;
  assign n15736 = n15735 ^ n8233 ^ n3318 ;
  assign n15737 = n9296 ^ n2732 ^ 1'b0 ;
  assign n15738 = n3919 | n5634 ;
  assign n15739 = n9536 | n15738 ;
  assign n15740 = n1493 & n6296 ;
  assign n15741 = n9910 & ~n15740 ;
  assign n15742 = n15739 & n15741 ;
  assign n15743 = n8483 & n11737 ;
  assign n15744 = n2051 & n15743 ;
  assign n15745 = ~n7739 & n15744 ;
  assign n15746 = ( ~n4039 & n4381 ) | ( ~n4039 & n12673 ) | ( n4381 & n12673 ) ;
  assign n15747 = n10282 ^ n214 ^ 1'b0 ;
  assign n15748 = n12199 & ~n15747 ;
  assign n15749 = ~n15746 & n15748 ;
  assign n15750 = n1878 & n15749 ;
  assign n15751 = n5097 ^ n845 ^ 1'b0 ;
  assign n15752 = ( ~n4116 & n5260 ) | ( ~n4116 & n15751 ) | ( n5260 & n15751 ) ;
  assign n15753 = n15752 ^ n5151 ^ 1'b0 ;
  assign n15754 = n11529 | n15753 ;
  assign n15755 = n7657 ^ n5054 ^ 1'b0 ;
  assign n15756 = n15754 | n15755 ;
  assign n15757 = n6817 & ~n9171 ;
  assign n15758 = n13885 & ~n15757 ;
  assign n15759 = ~n5917 & n15758 ;
  assign n15760 = n2701 | n10844 ;
  assign n15761 = n1104 & ~n6228 ;
  assign n15764 = n4033 & n6196 ;
  assign n15762 = n515 | n6644 ;
  assign n15763 = n6743 | n15762 ;
  assign n15765 = n15764 ^ n15763 ^ 1'b0 ;
  assign n15766 = n100 | n2861 ;
  assign n15767 = n8647 & ~n15766 ;
  assign n15768 = n15767 ^ n3113 ^ 1'b0 ;
  assign n15769 = n9248 & ~n15768 ;
  assign n15770 = n15769 ^ n188 ^ 1'b0 ;
  assign n15771 = n13726 & ~n15770 ;
  assign n15772 = n4291 ^ n970 ^ 1'b0 ;
  assign n15773 = n11208 | n15772 ;
  assign n15774 = n15773 ^ n4931 ^ 1'b0 ;
  assign n15775 = ~n4028 & n15774 ;
  assign n15776 = n5179 ^ n1313 ^ n212 ;
  assign n15779 = n5242 & n11333 ;
  assign n15780 = n14094 & n15779 ;
  assign n15777 = n2456 & ~n7882 ;
  assign n15778 = ~n1205 & n15777 ;
  assign n15781 = n15780 ^ n15778 ^ 1'b0 ;
  assign n15782 = ~n3712 & n15781 ;
  assign n15783 = n15776 & ~n15782 ;
  assign n15784 = n2987 & n15783 ;
  assign n15786 = ~n4813 & n12582 ;
  assign n15787 = n4668 & n15786 ;
  assign n15785 = n7131 & ~n8392 ;
  assign n15788 = n15787 ^ n15785 ^ n326 ;
  assign n15789 = n5949 & n10296 ;
  assign n15790 = n13463 ^ n7795 ^ 1'b0 ;
  assign n15791 = n3114 & ~n3318 ;
  assign n15792 = ~n10513 & n15791 ;
  assign n15793 = n15792 ^ n458 ^ 1'b0 ;
  assign n15794 = n645 | n15793 ;
  assign n15795 = n15794 ^ n14784 ^ 1'b0 ;
  assign n15796 = n2624 ^ n164 ^ 1'b0 ;
  assign n15797 = n5144 ^ n2029 ^ 1'b0 ;
  assign n15798 = ~n15796 & n15797 ;
  assign n15799 = n15798 ^ n5743 ^ 1'b0 ;
  assign n15800 = n6038 | n10477 ;
  assign n15801 = n15800 ^ n3661 ^ 1'b0 ;
  assign n15802 = n150 & n3420 ;
  assign n15803 = n431 & n15802 ;
  assign n15804 = ~n3723 & n9804 ;
  assign n15805 = ( n390 & ~n8834 ) | ( n390 & n15130 ) | ( ~n8834 & n15130 ) ;
  assign n15806 = n3425 | n15805 ;
  assign n15807 = n15804 | n15806 ;
  assign n15808 = n15807 ^ n13 ^ 1'b0 ;
  assign n15809 = n15803 | n15808 ;
  assign n15810 = n1707 & ~n2070 ;
  assign n15811 = n408 & n15810 ;
  assign n15812 = n11832 | n15811 ;
  assign n15813 = n9110 & ~n15812 ;
  assign n15814 = n10215 & n11685 ;
  assign n15815 = n15814 ^ n5632 ^ 1'b0 ;
  assign n15818 = ( ~n825 & n1501 ) | ( ~n825 & n8328 ) | ( n1501 & n8328 ) ;
  assign n15817 = n9995 ^ n9716 ^ 1'b0 ;
  assign n15819 = n15818 ^ n15817 ^ 1'b0 ;
  assign n15816 = n6596 & ~n9037 ;
  assign n15820 = n15819 ^ n15816 ^ 1'b0 ;
  assign n15821 = ~n8452 & n15820 ;
  assign n15822 = n1935 & n15821 ;
  assign n15829 = n273 & ~n2002 ;
  assign n15823 = n4881 ^ n721 ^ 1'b0 ;
  assign n15824 = n1736 | n15823 ;
  assign n15825 = n7589 & ~n15824 ;
  assign n15826 = n7474 ^ n1326 ^ 1'b0 ;
  assign n15827 = n15826 ^ n1672 ^ 1'b0 ;
  assign n15828 = n15825 & ~n15827 ;
  assign n15830 = n15829 ^ n15828 ^ 1'b0 ;
  assign n15831 = ~n11691 & n15830 ;
  assign n15832 = n1103 & ~n11781 ;
  assign n15833 = n15832 ^ n7578 ^ 1'b0 ;
  assign n15834 = n826 ^ n200 ^ 1'b0 ;
  assign n15835 = ~n4384 & n11069 ;
  assign n15836 = ~n3483 & n15835 ;
  assign n15842 = n716 & n3102 ;
  assign n15838 = n1528 & ~n15803 ;
  assign n15839 = ~n9451 & n15838 ;
  assign n15840 = n15839 ^ n7800 ^ 1'b0 ;
  assign n15841 = n7566 | n15840 ;
  assign n15843 = n15842 ^ n15841 ^ 1'b0 ;
  assign n15837 = ~n9068 & n13019 ;
  assign n15844 = n15843 ^ n15837 ^ 1'b0 ;
  assign n15845 = n7857 | n15246 ;
  assign n15846 = n13927 ^ n1267 ^ 1'b0 ;
  assign n15847 = n15278 & n15846 ;
  assign n15860 = ~n874 & n13915 ;
  assign n15861 = n4032 & n15860 ;
  assign n15857 = ~n6108 & n13069 ;
  assign n15858 = n15857 ^ n2716 ^ 1'b0 ;
  assign n15859 = n3582 & n15858 ;
  assign n15862 = n15861 ^ n15859 ^ 1'b0 ;
  assign n15851 = n9229 ^ n1243 ^ 1'b0 ;
  assign n15852 = n15851 ^ n466 ^ 1'b0 ;
  assign n15853 = n6846 | n15852 ;
  assign n15854 = ~n106 & n15853 ;
  assign n15855 = n5026 & n15854 ;
  assign n15856 = n15855 ^ n7951 ^ 1'b0 ;
  assign n15848 = n1994 & n10147 ;
  assign n15849 = n12598 ^ n647 ^ 1'b0 ;
  assign n15850 = ~n15848 & n15849 ;
  assign n15863 = n15862 ^ n15856 ^ n15850 ;
  assign n15864 = n4480 | n8128 ;
  assign n15865 = n15864 ^ n14256 ^ 1'b0 ;
  assign n15866 = n10306 | n12007 ;
  assign n15867 = n7508 & ~n15866 ;
  assign n15868 = n7476 ^ n5250 ^ 1'b0 ;
  assign n15869 = ~n139 & n15868 ;
  assign n15870 = n8214 ^ n7759 ^ 1'b0 ;
  assign n15871 = n5842 ^ n5282 ^ 1'b0 ;
  assign n15872 = ~n4169 & n15871 ;
  assign n15873 = n15872 ^ n7290 ^ 1'b0 ;
  assign n15874 = n13358 ^ n8258 ^ 1'b0 ;
  assign n15875 = n1410 & ~n5584 ;
  assign n15876 = ~n10381 & n15875 ;
  assign n15877 = ~n6589 & n14736 ;
  assign n15878 = n15877 ^ n532 ^ 1'b0 ;
  assign n15879 = n15876 & ~n15878 ;
  assign n15880 = n13366 ^ n3813 ^ 1'b0 ;
  assign n15881 = n10156 & ~n15880 ;
  assign n15882 = ~n1249 & n1943 ;
  assign n15883 = n8331 ^ n7767 ^ 1'b0 ;
  assign n15884 = n6359 ^ n1234 ^ 1'b0 ;
  assign n15885 = ~n11845 & n15884 ;
  assign n15886 = n14897 ^ n831 ^ 1'b0 ;
  assign n15887 = n15885 & ~n15886 ;
  assign n15888 = n10400 ^ n10262 ^ 1'b0 ;
  assign n15889 = n6638 ^ n1493 ^ 1'b0 ;
  assign n15890 = n5810 | n10300 ;
  assign n15891 = n2536 | n14904 ;
  assign n15892 = n15017 | n15891 ;
  assign n15893 = n1136 & n11770 ;
  assign n15894 = n14733 ^ n9796 ^ 1'b0 ;
  assign n15896 = n5700 & n9139 ;
  assign n15895 = ~n1385 & n11088 ;
  assign n15897 = n15896 ^ n15895 ^ 1'b0 ;
  assign n15898 = n6229 | n15897 ;
  assign n15899 = n15894 & ~n15898 ;
  assign n15900 = n8513 & n15899 ;
  assign n15901 = n4169 | n6680 ;
  assign n15902 = n15901 ^ n6166 ^ 1'b0 ;
  assign n15903 = n1591 & n2847 ;
  assign n15904 = n15903 ^ n6089 ^ 1'b0 ;
  assign n15905 = n15904 ^ n8083 ^ 1'b0 ;
  assign n15906 = n4644 & n9102 ;
  assign n15907 = n14455 & n15906 ;
  assign n15908 = ~n11620 & n15907 ;
  assign n15909 = n15908 ^ n10544 ^ 1'b0 ;
  assign n15914 = n5317 ^ n1306 ^ 1'b0 ;
  assign n15915 = ( ~n286 & n400 ) | ( ~n286 & n15914 ) | ( n400 & n15914 ) ;
  assign n15911 = n2350 | n5976 ;
  assign n15912 = n3003 | n15911 ;
  assign n15910 = n1995 & ~n3560 ;
  assign n15913 = n15912 ^ n15910 ^ 1'b0 ;
  assign n15916 = n15915 ^ n15913 ^ 1'b0 ;
  assign n15917 = n10119 & n11897 ;
  assign n15918 = n12870 & n15917 ;
  assign n15919 = ~n4200 & n15918 ;
  assign n15920 = n5758 & ~n10497 ;
  assign n15922 = n1876 & ~n6037 ;
  assign n15921 = n9546 ^ n901 ^ 1'b0 ;
  assign n15923 = n15922 ^ n15921 ^ n15896 ;
  assign n15924 = n15923 ^ n6526 ^ 1'b0 ;
  assign n15925 = n15920 | n15924 ;
  assign n15926 = ( n4044 & ~n15919 ) | ( n4044 & n15925 ) | ( ~n15919 & n15925 ) ;
  assign n15927 = n11166 ^ n4328 ^ 1'b0 ;
  assign n15928 = n4563 & ~n15927 ;
  assign n15929 = n11299 ^ n2631 ^ 1'b0 ;
  assign n15930 = n1870 | n3410 ;
  assign n15931 = n14382 & n15930 ;
  assign n15936 = n7187 ^ n1842 ^ 1'b0 ;
  assign n15937 = ~n8830 & n15936 ;
  assign n15932 = n9229 ^ n6080 ^ n2151 ;
  assign n15933 = n6374 ^ n2843 ^ 1'b0 ;
  assign n15934 = n15932 & n15933 ;
  assign n15935 = n15934 ^ n13887 ^ 1'b0 ;
  assign n15938 = n15937 ^ n15935 ^ 1'b0 ;
  assign n15939 = n7687 & n13528 ;
  assign n15940 = n5080 ^ n1010 ^ 1'b0 ;
  assign n15941 = n11876 | n12824 ;
  assign n15942 = n15941 ^ n490 ^ 1'b0 ;
  assign n15943 = n15940 | n15942 ;
  assign n15944 = n4386 | n15943 ;
  assign n15945 = n15944 ^ n5293 ^ 1'b0 ;
  assign n15946 = ( n4351 & ~n8531 ) | ( n4351 & n12280 ) | ( ~n8531 & n12280 ) ;
  assign n15947 = n10542 ^ n4468 ^ 1'b0 ;
  assign n15948 = n15946 | n15947 ;
  assign n15949 = n8505 ^ n7249 ^ 1'b0 ;
  assign n15950 = n8486 | n15949 ;
  assign n15951 = n3825 | n5302 ;
  assign n15952 = n12608 & ~n15951 ;
  assign n15953 = n15952 ^ n14898 ^ 1'b0 ;
  assign n15954 = n5046 & n5195 ;
  assign n15955 = n15954 ^ n10161 ^ 1'b0 ;
  assign n15956 = n9208 & n15955 ;
  assign n15957 = n1918 ^ n1258 ^ 1'b0 ;
  assign n15958 = n5304 | n5954 ;
  assign n15959 = n8239 | n10452 ;
  assign n15960 = n15959 ^ n2875 ^ 1'b0 ;
  assign n15961 = n2767 | n12147 ;
  assign n15962 = n15961 ^ n12480 ^ 1'b0 ;
  assign n15963 = n15960 & ~n15962 ;
  assign n15964 = n12305 ^ n6305 ^ 1'b0 ;
  assign n15965 = n4829 & ~n5897 ;
  assign n15966 = n15965 ^ n10717 ^ 1'b0 ;
  assign n15967 = n15966 ^ n8770 ^ 1'b0 ;
  assign n15968 = n2937 | n6394 ;
  assign n15969 = n15968 ^ n11423 ^ 1'b0 ;
  assign n15970 = n774 & ~n15969 ;
  assign n15971 = n15970 ^ n1216 ^ 1'b0 ;
  assign n15972 = n14456 | n15971 ;
  assign n15973 = ( ~n5997 & n15967 ) | ( ~n5997 & n15972 ) | ( n15967 & n15972 ) ;
  assign n15974 = n15973 ^ n11050 ^ n1481 ;
  assign n15975 = n1411 | n5336 ;
  assign n15976 = ~n14309 & n15975 ;
  assign n15977 = n3723 | n11521 ;
  assign n15978 = n7657 & ~n15977 ;
  assign n15979 = n374 | n490 ;
  assign n15980 = n374 & ~n15979 ;
  assign n15981 = n15980 ^ n2317 ^ 1'b0 ;
  assign n15982 = n327 & ~n889 ;
  assign n15983 = ~n327 & n15982 ;
  assign n15984 = n1600 & n15983 ;
  assign n15985 = ~n4657 & n15984 ;
  assign n15986 = ~n15981 & n15985 ;
  assign n15987 = n15981 & n15986 ;
  assign n15988 = n12852 | n15987 ;
  assign n15989 = n14736 | n15988 ;
  assign n15990 = n15988 & ~n15989 ;
  assign n15991 = n12950 ^ n12461 ^ 1'b0 ;
  assign n15992 = n9179 & n15991 ;
  assign n15994 = n823 & n14401 ;
  assign n15995 = n15994 ^ n1329 ^ 1'b0 ;
  assign n15996 = n15995 ^ n7531 ^ 1'b0 ;
  assign n15993 = n2796 | n7123 ;
  assign n15997 = n15996 ^ n15993 ^ 1'b0 ;
  assign n15998 = n3331 & n13026 ;
  assign n15999 = n372 & n15998 ;
  assign n16000 = n15999 ^ n14308 ^ n7155 ;
  assign n16001 = n508 | n4143 ;
  assign n16002 = n16001 ^ n2603 ^ 1'b0 ;
  assign n16003 = n10152 | n14934 ;
  assign n16004 = n13021 ^ n3414 ^ 1'b0 ;
  assign n16005 = ~n4853 & n16004 ;
  assign n16006 = n16005 ^ n4253 ^ 1'b0 ;
  assign n16007 = n14944 ^ n2802 ^ 1'b0 ;
  assign n16008 = n16007 ^ n5551 ^ 1'b0 ;
  assign n16009 = n5359 ^ n4687 ^ 1'b0 ;
  assign n16010 = ~n3214 & n16009 ;
  assign n16011 = n10944 ^ n406 ^ 1'b0 ;
  assign n16012 = n1742 & ~n16011 ;
  assign n16015 = n1152 ^ n961 ^ n666 ;
  assign n16016 = ( ~n7758 & n9831 ) | ( ~n7758 & n16015 ) | ( n9831 & n16015 ) ;
  assign n16013 = n9249 | n15612 ;
  assign n16014 = n14276 & n16013 ;
  assign n16017 = n16016 ^ n16014 ^ 1'b0 ;
  assign n16018 = n3125 | n5329 ;
  assign n16019 = n4722 ^ n81 ^ 1'b0 ;
  assign n16020 = ( n676 & ~n4040 ) | ( n676 & n4151 ) | ( ~n4040 & n4151 ) ;
  assign n16021 = n5626 | n16020 ;
  assign n16022 = n8830 | n16021 ;
  assign n16023 = n15803 & ~n16022 ;
  assign n16024 = n5557 ^ n1534 ^ 1'b0 ;
  assign n16025 = n6653 & n16024 ;
  assign n16026 = n13947 ^ n2214 ^ 1'b0 ;
  assign n16027 = ~n9048 & n15907 ;
  assign n16028 = ~n5158 & n16027 ;
  assign n16029 = n2424 & ~n10259 ;
  assign n16030 = ~n3790 & n16029 ;
  assign n16031 = ~n7256 & n13328 ;
  assign n16032 = n12899 ^ n9332 ^ 1'b0 ;
  assign n16033 = n16032 ^ n1510 ^ 1'b0 ;
  assign n16034 = n8124 | n11802 ;
  assign n16035 = n1837 & ~n16034 ;
  assign n16036 = n1576 | n6942 ;
  assign n16037 = n9465 & ~n16036 ;
  assign n16038 = n16037 ^ n9145 ^ 1'b0 ;
  assign n16039 = n8036 | n16038 ;
  assign n16040 = n9857 ^ n6588 ^ 1'b0 ;
  assign n16041 = n15632 ^ n15582 ^ n15268 ;
  assign n16042 = n6433 ^ n2455 ^ 1'b0 ;
  assign n16043 = n568 & ~n8876 ;
  assign n16044 = n16043 ^ n15076 ^ 1'b0 ;
  assign n16045 = ~n265 & n4461 ;
  assign n16046 = n16045 ^ n3835 ^ 1'b0 ;
  assign n16047 = n7860 & ~n16046 ;
  assign n16048 = n401 & n6237 ;
  assign n16049 = n12069 & n16048 ;
  assign n16050 = ~n4046 & n16049 ;
  assign n16051 = n16050 ^ n1403 ^ 1'b0 ;
  assign n16052 = ~n4519 & n16051 ;
  assign n16061 = n9529 ^ n5888 ^ 1'b0 ;
  assign n16062 = n4607 | n16061 ;
  assign n16063 = n16062 ^ n7768 ^ n2521 ;
  assign n16054 = n4058 & n4369 ;
  assign n16055 = n1506 & n16054 ;
  assign n16056 = ( n2041 & ~n3073 ) | ( n2041 & n16055 ) | ( ~n3073 & n16055 ) ;
  assign n16053 = ( n2272 & n3194 ) | ( n2272 & n4745 ) | ( n3194 & n4745 ) ;
  assign n16057 = n16056 ^ n16053 ^ 1'b0 ;
  assign n16058 = n11862 | n16057 ;
  assign n16059 = n9818 | n16058 ;
  assign n16060 = ~n11083 & n16059 ;
  assign n16064 = n16063 ^ n16060 ^ 1'b0 ;
  assign n16065 = n6846 | n9634 ;
  assign n16066 = n3199 | n16065 ;
  assign n16067 = n1159 | n16066 ;
  assign n16068 = n14727 ^ n1083 ^ 1'b0 ;
  assign n16069 = ~n6245 & n6647 ;
  assign n16070 = n2460 | n16069 ;
  assign n16071 = n4384 & ~n14137 ;
  assign n16072 = n10388 & ~n10845 ;
  assign n16073 = ~n12224 & n16072 ;
  assign n16074 = n8168 & n9455 ;
  assign n16075 = n760 & n7271 ;
  assign n16076 = ~n451 & n16075 ;
  assign n16077 = ( n16033 & ~n16074 ) | ( n16033 & n16076 ) | ( ~n16074 & n16076 ) ;
  assign n16078 = n15045 ^ n4245 ^ 1'b0 ;
  assign n16079 = ~n6048 & n16078 ;
  assign n16080 = n142 | n4480 ;
  assign n16081 = n16079 | n16080 ;
  assign n16082 = n16081 ^ n15552 ^ 1'b0 ;
  assign n16083 = n15754 | n16082 ;
  assign n16084 = n10254 ^ n2891 ^ 1'b0 ;
  assign n16085 = n9095 & n16084 ;
  assign n16088 = n2753 | n10331 ;
  assign n16089 = n831 | n1063 ;
  assign n16090 = n11123 & ~n16089 ;
  assign n16091 = n16088 & n16090 ;
  assign n16086 = n7414 & ~n8356 ;
  assign n16087 = ~n3971 & n16086 ;
  assign n16092 = n16091 ^ n16087 ^ 1'b0 ;
  assign n16093 = n3655 ^ n2938 ^ 1'b0 ;
  assign n16094 = ~n1372 & n16093 ;
  assign n16095 = n2883 & ~n4229 ;
  assign n16096 = n16095 ^ n1297 ^ 1'b0 ;
  assign n16097 = n5520 | n16096 ;
  assign n16098 = n1020 & ~n16097 ;
  assign n16099 = n16094 | n16098 ;
  assign n16100 = n3818 & ~n6040 ;
  assign n16101 = n16100 ^ n7542 ^ 1'b0 ;
  assign n16102 = n15477 & n16101 ;
  assign n16103 = n16102 ^ n7151 ^ 1'b0 ;
  assign n16104 = n15341 & n16103 ;
  assign n16105 = ~n5873 & n10728 ;
  assign n16106 = n1567 & n16105 ;
  assign n16107 = ~n778 & n13454 ;
  assign n16108 = n1459 & ~n3839 ;
  assign n16117 = ~n2094 & n3790 ;
  assign n16114 = n11699 ^ n8012 ^ 1'b0 ;
  assign n16115 = n2833 & ~n16114 ;
  assign n16111 = n1036 & n2822 ;
  assign n16109 = n443 & n525 ;
  assign n16110 = n1257 & n16109 ;
  assign n16112 = n16111 ^ n16110 ^ 1'b0 ;
  assign n16113 = n1574 & ~n16112 ;
  assign n16116 = n16115 ^ n16113 ^ 1'b0 ;
  assign n16118 = n16117 ^ n16116 ^ 1'b0 ;
  assign n16120 = n515 & n1978 ;
  assign n16121 = n525 & n16120 ;
  assign n16122 = ~n525 & n16121 ;
  assign n16119 = ~n27 & n559 ;
  assign n16123 = n16122 ^ n16119 ^ 1'b0 ;
  assign n16124 = n5936 & n16123 ;
  assign n16125 = n6717 & n11542 ;
  assign n16126 = n16125 ^ n6103 ^ 1'b0 ;
  assign n16127 = n13631 ^ n8130 ^ n7251 ;
  assign n16128 = n16127 ^ n7731 ^ n31 ;
  assign n16129 = n9693 ^ n8029 ^ 1'b0 ;
  assign n16130 = n4755 & ~n15326 ;
  assign n16131 = n16130 ^ n682 ^ 1'b0 ;
  assign n16132 = n2358 & n12037 ;
  assign n16133 = n11936 & n16132 ;
  assign n16134 = n14880 ^ n6832 ^ 1'b0 ;
  assign n16135 = ~n15472 & n16134 ;
  assign n16136 = n3472 & n13485 ;
  assign n16137 = n15725 & n16136 ;
  assign n16138 = n3955 & ~n7918 ;
  assign n16139 = n8477 & n16138 ;
  assign n16140 = ~n5978 & n16139 ;
  assign n16141 = ~n3313 & n16140 ;
  assign n16142 = n4720 ^ n1956 ^ 1'b0 ;
  assign n16143 = n14675 ^ n11289 ^ 1'b0 ;
  assign n16144 = n3757 & n4468 ;
  assign n16145 = n16144 ^ n5880 ^ 1'b0 ;
  assign n16146 = n3531 | n16052 ;
  assign n16147 = n1506 & ~n9304 ;
  assign n16148 = n7124 ^ n1385 ^ 1'b0 ;
  assign n16149 = n10449 ^ n2426 ^ 1'b0 ;
  assign n16150 = n16148 & ~n16149 ;
  assign n16151 = n16150 ^ n3418 ^ 1'b0 ;
  assign n16152 = ~n6768 & n16151 ;
  assign n16153 = n6080 | n11954 ;
  assign n16154 = n3308 | n9491 ;
  assign n16155 = n8872 & ~n16154 ;
  assign n16156 = n11334 | n14820 ;
  assign n16157 = n16156 ^ n13941 ^ 1'b0 ;
  assign n16158 = ~n590 & n16157 ;
  assign n16159 = n16155 & n16158 ;
  assign n16160 = n15243 ^ n229 ^ 1'b0 ;
  assign n16161 = n12041 ^ n7151 ^ 1'b0 ;
  assign n16162 = n810 ^ n13 ^ 1'b0 ;
  assign n16163 = ~n16161 & n16162 ;
  assign n16165 = n2531 | n2645 ;
  assign n16166 = n1276 & ~n9304 ;
  assign n16167 = ~n16165 & n16166 ;
  assign n16164 = n9457 ^ n2000 ^ 1'b0 ;
  assign n16168 = n16167 ^ n16164 ^ 1'b0 ;
  assign n16169 = n2812 & n3592 ;
  assign n16170 = n3753 & ~n7156 ;
  assign n16171 = n7983 ^ n6756 ^ 1'b0 ;
  assign n16172 = n15680 ^ n9526 ^ 1'b0 ;
  assign n16173 = n4691 & n13980 ;
  assign n16174 = n8291 & ~n8719 ;
  assign n16175 = n16174 ^ n14249 ^ 1'b0 ;
  assign n16176 = n2637 ^ n1656 ^ 1'b0 ;
  assign n16177 = n4248 & n11077 ;
  assign n16178 = n13245 ^ n9585 ^ 1'b0 ;
  assign n16179 = ~n11238 & n16178 ;
  assign n16180 = n14217 ^ n9468 ^ 1'b0 ;
  assign n16181 = n1215 & n13741 ;
  assign n16182 = n3225 | n8843 ;
  assign n16183 = n16182 ^ n221 ^ 1'b0 ;
  assign n16184 = n25 & n16183 ;
  assign n16185 = n16184 ^ n4495 ^ 1'b0 ;
  assign n16186 = n11291 ^ n43 ^ 1'b0 ;
  assign n16187 = n16186 ^ n1718 ^ 1'b0 ;
  assign n16188 = ~n9413 & n16187 ;
  assign n16189 = n1442 ^ n1109 ^ 1'b0 ;
  assign n16190 = ~n442 & n16189 ;
  assign n16191 = n13776 & n16190 ;
  assign n16192 = n5124 & n16191 ;
  assign n16193 = n16188 | n16192 ;
  assign n16194 = n5399 & n16193 ;
  assign n16195 = ~n16185 & n16194 ;
  assign n16196 = ~n10424 & n13002 ;
  assign n16197 = n16196 ^ n8307 ^ 1'b0 ;
  assign n16198 = ~n4893 & n16197 ;
  assign n16199 = n667 & n16198 ;
  assign n16200 = n13430 ^ n4862 ^ 1'b0 ;
  assign n16201 = n7620 & n16200 ;
  assign n16202 = n10389 | n16201 ;
  assign n16203 = n11044 & n11576 ;
  assign n16204 = n3351 ^ n1121 ^ 1'b0 ;
  assign n16205 = n11390 | n16204 ;
  assign n16206 = n6678 & ~n16205 ;
  assign n16207 = ~n6993 & n14385 ;
  assign n16208 = n10220 ^ n1656 ^ 1'b0 ;
  assign n16209 = n16208 ^ n11572 ^ 1'b0 ;
  assign n16210 = n12094 ^ n1556 ^ 1'b0 ;
  assign n16211 = n16210 ^ n2739 ^ 1'b0 ;
  assign n16212 = n16211 ^ n5059 ^ 1'b0 ;
  assign n16213 = ~n11140 & n16212 ;
  assign n16214 = n5549 ^ n2411 ^ 1'b0 ;
  assign n16215 = ~n10527 & n16214 ;
  assign n16216 = n8151 ^ n5236 ^ 1'b0 ;
  assign n16217 = ( ~n2039 & n2695 ) | ( ~n2039 & n4862 ) | ( n2695 & n4862 ) ;
  assign n16218 = n2304 | n16217 ;
  assign n16219 = n16218 ^ n8478 ^ 1'b0 ;
  assign n16220 = n7994 ^ n5510 ^ n214 ;
  assign n16221 = n582 | n2779 ;
  assign n16222 = n3106 | n16221 ;
  assign n16223 = n8237 & ~n16222 ;
  assign n16224 = n16223 ^ n5311 ^ 1'b0 ;
  assign n16225 = n9889 & n13531 ;
  assign n16226 = n12551 & ~n13356 ;
  assign n16227 = n16225 & n16226 ;
  assign n16228 = n598 & ~n14724 ;
  assign n16229 = ~n598 & n16228 ;
  assign n16230 = n2543 & ~n12754 ;
  assign n16231 = n2709 ^ n1312 ^ 1'b0 ;
  assign n16232 = n5892 & ~n14330 ;
  assign n16233 = n3366 & n16232 ;
  assign n16239 = n5445 & n15059 ;
  assign n16234 = ~n600 & n6215 ;
  assign n16235 = n8275 ^ n211 ^ 1'b0 ;
  assign n16236 = n827 & ~n16235 ;
  assign n16237 = n16236 ^ n11556 ^ 1'b0 ;
  assign n16238 = n16234 & ~n16237 ;
  assign n16240 = n16239 ^ n16238 ^ 1'b0 ;
  assign n16243 = n13407 ^ n6930 ^ n4307 ;
  assign n16241 = n6311 | n12244 ;
  assign n16242 = n3753 | n16241 ;
  assign n16244 = n16243 ^ n16242 ^ 1'b0 ;
  assign n16245 = n265 & ~n9043 ;
  assign n16246 = n6027 & n12622 ;
  assign n16247 = ~n12347 & n16246 ;
  assign n16250 = ~n9447 & n15858 ;
  assign n16251 = n16250 ^ n978 ^ 1'b0 ;
  assign n16248 = n8432 ^ n8120 ^ 1'b0 ;
  assign n16249 = n2615 & n16248 ;
  assign n16252 = n16251 ^ n16249 ^ 1'b0 ;
  assign n16253 = n11649 | n16252 ;
  assign n16254 = n10579 ^ n9076 ^ 1'b0 ;
  assign n16255 = ~n11199 & n16254 ;
  assign n16256 = n10564 ^ n3998 ^ n873 ;
  assign n16257 = n3211 ^ n2130 ^ 1'b0 ;
  assign n16258 = ~n2048 & n2639 ;
  assign n16259 = n16258 ^ n76 ^ 1'b0 ;
  assign n16260 = n2610 & ~n16259 ;
  assign n16261 = n2336 & ~n6846 ;
  assign n16262 = n16261 ^ n6224 ^ 1'b0 ;
  assign n16263 = n14472 ^ n14240 ^ 1'b0 ;
  assign n16264 = n12413 | n16263 ;
  assign n16265 = n10976 | n16264 ;
  assign n16266 = n3971 | n10270 ;
  assign n16267 = n7779 & ~n16266 ;
  assign n16268 = n8216 | n8894 ;
  assign n16269 = ~n150 & n5023 ;
  assign n16270 = n16269 ^ n10149 ^ 1'b0 ;
  assign n16271 = ~n11613 & n16270 ;
  assign n16272 = n16271 ^ n5680 ^ 1'b0 ;
  assign n16273 = n8219 ^ n4840 ^ 1'b0 ;
  assign n16274 = n7155 & ~n16273 ;
  assign n16275 = n13534 | n16274 ;
  assign n16276 = n722 & ~n1794 ;
  assign n16277 = ~n722 & n16276 ;
  assign n16278 = n2875 & ~n16277 ;
  assign n16279 = n16278 ^ n1845 ^ 1'b0 ;
  assign n16280 = n11907 & ~n14612 ;
  assign n16281 = n12528 ^ n4079 ^ 1'b0 ;
  assign n16282 = n2833 & ~n13030 ;
  assign n16283 = ~n2458 & n10757 ;
  assign n16284 = n16283 ^ n11801 ^ 1'b0 ;
  assign n16287 = n8567 ^ n3818 ^ n2806 ;
  assign n16288 = n8998 ^ n7197 ^ 1'b0 ;
  assign n16289 = ~n16287 & n16288 ;
  assign n16285 = n2856 ^ n826 ^ 1'b0 ;
  assign n16286 = n16285 ^ n14215 ^ 1'b0 ;
  assign n16290 = n16289 ^ n16286 ^ 1'b0 ;
  assign n16291 = n15460 ^ n1047 ^ 1'b0 ;
  assign n16292 = n8980 ^ n6406 ^ 1'b0 ;
  assign n16293 = ~n316 & n16292 ;
  assign n16294 = n16293 ^ n14008 ^ n7999 ;
  assign n16298 = ~n4808 & n11710 ;
  assign n16296 = n3211 ^ n387 ^ 1'b0 ;
  assign n16295 = n9745 & n12115 ;
  assign n16297 = n16296 ^ n16295 ^ 1'b0 ;
  assign n16299 = n16298 ^ n16297 ^ 1'b0 ;
  assign n16300 = n584 | n12521 ;
  assign n16301 = n16300 ^ n14474 ^ 1'b0 ;
  assign n16302 = n6468 | n8363 ;
  assign n16303 = n6196 ^ n2879 ^ n2248 ;
  assign n16304 = ~n15940 & n16303 ;
  assign n16305 = n16304 ^ n5623 ^ 1'b0 ;
  assign n16306 = n8463 ^ n3957 ^ 1'b0 ;
  assign n16307 = ~n4169 & n6173 ;
  assign n16308 = n16307 ^ n8460 ^ 1'b0 ;
  assign n16309 = ( ~n1821 & n4364 ) | ( ~n1821 & n16308 ) | ( n4364 & n16308 ) ;
  assign n16310 = ( n4515 & ~n8720 ) | ( n4515 & n16309 ) | ( ~n8720 & n16309 ) ;
  assign n16311 = n11174 & n13050 ;
  assign n16312 = n16311 ^ n14502 ^ 1'b0 ;
  assign n16313 = n3162 & ~n16312 ;
  assign n16314 = n3386 & ~n8259 ;
  assign n16315 = n2442 | n12337 ;
  assign n16316 = n10614 ^ n6723 ^ 1'b0 ;
  assign n16317 = n7041 & n16316 ;
  assign n16318 = ~n13184 & n16317 ;
  assign n16319 = n2033 ^ n598 ^ 1'b0 ;
  assign n16320 = n2185 | n2567 ;
  assign n16321 = n754 & ~n6927 ;
  assign n16322 = n11927 & ~n16321 ;
  assign n16323 = n14144 ^ n8331 ^ 1'b0 ;
  assign n16324 = n2439 & ~n2790 ;
  assign n16325 = n16324 ^ n966 ^ 1'b0 ;
  assign n16326 = n2040 & ~n16325 ;
  assign n16327 = n16326 ^ n2552 ^ 1'b0 ;
  assign n16328 = n16323 & n16327 ;
  assign n16329 = n3867 & ~n9189 ;
  assign n16330 = n16329 ^ n4510 ^ 1'b0 ;
  assign n16331 = n342 & n2140 ;
  assign n16332 = ~n12784 & n16331 ;
  assign n16333 = n4218 | n12119 ;
  assign n16334 = n12789 & ~n16333 ;
  assign n16335 = n1566 | n13671 ;
  assign n16336 = n13106 ^ n5040 ^ 1'b0 ;
  assign n16337 = n16335 & n16336 ;
  assign n16338 = n2802 | n5492 ;
  assign n16339 = n1350 & ~n10105 ;
  assign n16340 = n16339 ^ n7578 ^ 1'b0 ;
  assign n16341 = n16340 ^ n3968 ^ 1'b0 ;
  assign n16342 = n15440 & n16341 ;
  assign n16343 = n48 & ~n285 ;
  assign n16344 = n16343 ^ n963 ^ 1'b0 ;
  assign n16345 = n16344 ^ n3698 ^ 1'b0 ;
  assign n16346 = n910 & n16345 ;
  assign n16347 = n9916 ^ n5654 ^ 1'b0 ;
  assign n16348 = n2085 & ~n16347 ;
  assign n16349 = ~n27 & n16348 ;
  assign n16350 = ~n9710 & n16349 ;
  assign n16351 = n3817 | n16350 ;
  assign n16352 = n130 & n1045 ;
  assign n16353 = n16352 ^ n466 ^ 1'b0 ;
  assign n16354 = n3968 | n16353 ;
  assign n16355 = n6296 | n16354 ;
  assign n16356 = ~n9288 & n16355 ;
  assign n16357 = n11360 & ~n15639 ;
  assign n16358 = ~n5719 & n16357 ;
  assign n16359 = n1401 & n7556 ;
  assign n16360 = ~n723 & n1745 ;
  assign n16361 = n8714 | n16360 ;
  assign n16362 = n16359 | n16361 ;
  assign n16363 = n8891 ^ n4370 ^ 1'b0 ;
  assign n16364 = n7907 | n16363 ;
  assign n16365 = n4526 | n5531 ;
  assign n16366 = ~n2719 & n8477 ;
  assign n16367 = n16366 ^ n3226 ^ 1'b0 ;
  assign n16368 = ~n5630 & n7019 ;
  assign n16369 = n16367 & n16368 ;
  assign n16370 = n16369 ^ n7089 ^ 1'b0 ;
  assign n16371 = ~n8838 & n16370 ;
  assign n16372 = n2275 & ~n6662 ;
  assign n16373 = n2056 & n16372 ;
  assign n16374 = n1184 & ~n9525 ;
  assign n16375 = ~n3644 & n16374 ;
  assign n16376 = n16373 & n16375 ;
  assign n16377 = n9693 ^ n1121 ^ 1'b0 ;
  assign n16378 = n701 & n4189 ;
  assign n16379 = n16378 ^ n7126 ^ 1'b0 ;
  assign n16380 = n9268 & ~n9526 ;
  assign n16381 = ~n16379 & n16380 ;
  assign n16382 = n5031 & n16381 ;
  assign n16383 = n3521 & ~n16382 ;
  assign n16384 = n16383 ^ n3221 ^ 1'b0 ;
  assign n16385 = ( n4087 & ~n13664 ) | ( n4087 & n16384 ) | ( ~n13664 & n16384 ) ;
  assign n16386 = n4657 ^ n575 ^ 1'b0 ;
  assign n16387 = n16386 ^ n459 ^ 1'b0 ;
  assign n16388 = n15511 ^ n5321 ^ 1'b0 ;
  assign n16389 = n16388 ^ n2178 ^ 1'b0 ;
  assign n16390 = n16387 & n16389 ;
  assign n16391 = n451 ^ n334 ^ 1'b0 ;
  assign n16392 = n16391 ^ n11504 ^ n4020 ;
  assign n16393 = n1094 & ~n15619 ;
  assign n16394 = ( n342 & ~n7940 ) | ( n342 & n9114 ) | ( ~n7940 & n9114 ) ;
  assign n16395 = ~n901 & n16394 ;
  assign n16396 = n5511 | n8001 ;
  assign n16397 = n13663 & ~n16396 ;
  assign n16398 = ~n2250 & n14675 ;
  assign n16399 = n6458 ^ n2108 ^ 1'b0 ;
  assign n16400 = ( n5958 & ~n7951 ) | ( n5958 & n16399 ) | ( ~n7951 & n16399 ) ;
  assign n16401 = n13580 & ~n16400 ;
  assign n16402 = ~n1848 & n5802 ;
  assign n16403 = n4400 & n16402 ;
  assign n16404 = n911 | n16403 ;
  assign n16405 = n9261 ^ n2496 ^ 1'b0 ;
  assign n16408 = n3601 & ~n8909 ;
  assign n16409 = ( ~n5209 & n6092 ) | ( ~n5209 & n16408 ) | ( n6092 & n16408 ) ;
  assign n16406 = ( n995 & n4090 ) | ( n995 & n11722 ) | ( n4090 & n11722 ) ;
  assign n16407 = n12337 | n16406 ;
  assign n16410 = n16409 ^ n16407 ^ n6662 ;
  assign n16411 = n11345 ^ n1235 ^ 1'b0 ;
  assign n16412 = n11169 ^ n1469 ^ 1'b0 ;
  assign n16413 = n3887 | n9049 ;
  assign n16414 = n1567 ^ n961 ^ 1'b0 ;
  assign n16415 = n16414 ^ n725 ^ 1'b0 ;
  assign n16416 = ~n2097 & n7449 ;
  assign n16417 = n3724 & n16416 ;
  assign n16418 = ( ~n1448 & n8357 ) | ( ~n1448 & n16417 ) | ( n8357 & n16417 ) ;
  assign n16419 = n8368 | n16418 ;
  assign n16420 = n5744 ^ n880 ^ 1'b0 ;
  assign n16421 = n8451 & ~n16420 ;
  assign n16422 = ~n4143 & n16421 ;
  assign n16423 = n914 & n6079 ;
  assign n16424 = ( n7729 & n10473 ) | ( n7729 & ~n16423 ) | ( n10473 & ~n16423 ) ;
  assign n16425 = n8950 ^ n8233 ^ 1'b0 ;
  assign n16426 = n16425 ^ n13529 ^ 1'b0 ;
  assign n16427 = n11313 ^ n6298 ^ 1'b0 ;
  assign n16428 = n12665 ^ n7262 ^ n249 ;
  assign n16429 = ~n2869 & n9624 ;
  assign n16430 = n12919 & n16429 ;
  assign n16431 = n16430 ^ n4422 ^ 1'b0 ;
  assign n16432 = n16431 ^ n4074 ^ 1'b0 ;
  assign n16433 = n2207 & ~n16432 ;
  assign n16434 = n1369 | n2532 ;
  assign n16435 = n16434 ^ n14318 ^ 1'b0 ;
  assign n16436 = n3636 & ~n14052 ;
  assign n16437 = n8745 ^ n1187 ^ 1'b0 ;
  assign n16438 = n1024 | n16437 ;
  assign n16439 = ( n2973 & n12913 ) | ( n2973 & ~n16438 ) | ( n12913 & ~n16438 ) ;
  assign n16440 = n15644 ^ n6542 ^ 1'b0 ;
  assign n16441 = n221 & n8801 ;
  assign n16442 = n16441 ^ n503 ^ 1'b0 ;
  assign n16443 = n10329 & ~n16442 ;
  assign n16444 = n16443 ^ n3917 ^ 1'b0 ;
  assign n16445 = ~n10249 & n16444 ;
  assign n16446 = n5760 | n16445 ;
  assign n16447 = n2848 | n16446 ;
  assign n16448 = n9199 | n11907 ;
  assign n16449 = n16448 ^ n15310 ^ 1'b0 ;
  assign n16450 = n4917 | n16449 ;
  assign n16451 = ~n778 & n7999 ;
  assign n16452 = n3486 & ~n16451 ;
  assign n16453 = n16452 ^ n3293 ^ 1'b0 ;
  assign n16461 = n9186 | n14977 ;
  assign n16460 = n5535 ^ n4046 ^ 1'b0 ;
  assign n16462 = n16461 ^ n16460 ^ 1'b0 ;
  assign n16454 = n5309 ^ n3265 ^ n1403 ;
  assign n16455 = ~n5724 & n16454 ;
  assign n16456 = n16455 ^ n4551 ^ n1608 ;
  assign n16457 = ~n1522 & n3715 ;
  assign n16458 = ~n1969 & n16457 ;
  assign n16459 = n16456 & ~n16458 ;
  assign n16463 = n16462 ^ n16459 ^ 1'b0 ;
  assign n16464 = n6193 ^ n1182 ^ 1'b0 ;
  assign n16465 = n16464 ^ n13951 ^ 1'b0 ;
  assign n16466 = n7398 ^ n1264 ^ 1'b0 ;
  assign n16467 = n695 | n5028 ;
  assign n16468 = n5618 ^ n3418 ^ 1'b0 ;
  assign n16469 = ~n6173 & n6516 ;
  assign n16470 = ~n14831 & n16469 ;
  assign n16471 = ( n5131 & n8508 ) | ( n5131 & n16358 ) | ( n8508 & n16358 ) ;
  assign n16472 = ~n14122 & n15099 ;
  assign n16473 = n3098 & ~n10362 ;
  assign n16476 = n4400 | n7621 ;
  assign n16477 = n892 & ~n16476 ;
  assign n16478 = ( n1437 & ~n1508 ) | ( n1437 & n4568 ) | ( ~n1508 & n4568 ) ;
  assign n16479 = ~n294 & n16478 ;
  assign n16480 = n12380 | n16479 ;
  assign n16481 = n16480 ^ n10964 ^ 1'b0 ;
  assign n16482 = ~n16477 & n16481 ;
  assign n16474 = n590 | n1247 ;
  assign n16475 = n15275 | n16474 ;
  assign n16483 = n16482 ^ n16475 ^ 1'b0 ;
  assign n16484 = n5445 ^ n412 ^ 1'b0 ;
  assign n16485 = n8543 & n16484 ;
  assign n16486 = ~n10004 & n16485 ;
  assign n16487 = n16486 ^ n8443 ^ 1'b0 ;
  assign n16488 = n5452 ^ n1679 ^ 1'b0 ;
  assign n16489 = ~n1164 & n16488 ;
  assign n16490 = ~n2875 & n16489 ;
  assign n16491 = n16490 ^ n360 ^ 1'b0 ;
  assign n16492 = n2981 | n6556 ;
  assign n16493 = n117 & ~n16492 ;
  assign n16494 = n5539 ^ n423 ^ 1'b0 ;
  assign n16495 = ~n16493 & n16494 ;
  assign n16496 = ( n6542 & ~n15905 ) | ( n6542 & n16495 ) | ( ~n15905 & n16495 ) ;
  assign n16498 = n219 | n3609 ;
  assign n16499 = n2140 | n16498 ;
  assign n16497 = n5489 | n11300 ;
  assign n16500 = n16499 ^ n16497 ^ n266 ;
  assign n16501 = n16500 ^ n5594 ^ 1'b0 ;
  assign n16502 = n15177 ^ n13290 ^ n3232 ;
  assign n16503 = n8675 & ~n16502 ;
  assign n16504 = n16503 ^ n8681 ^ 1'b0 ;
  assign n16505 = n12986 ^ n11582 ^ 1'b0 ;
  assign n16506 = ( ~n4519 & n9670 ) | ( ~n4519 & n14477 ) | ( n9670 & n14477 ) ;
  assign n16507 = ( ~n6456 & n12458 ) | ( ~n6456 & n16506 ) | ( n12458 & n16506 ) ;
  assign n16508 = n14977 ^ x11 ^ 1'b0 ;
  assign n16509 = n11978 & ~n14334 ;
  assign n16510 = n1863 & n6201 ;
  assign n16511 = ~n963 & n16510 ;
  assign n16512 = n15504 & n16511 ;
  assign n16513 = n1682 & ~n10063 ;
  assign n16514 = n16512 & ~n16513 ;
  assign n16515 = ~n541 & n9604 ;
  assign n16516 = n3361 & n8904 ;
  assign n16517 = ~n11462 & n15481 ;
  assign n16518 = n1590 & ~n7029 ;
  assign n16519 = ~n1187 & n3139 ;
  assign n16520 = ~n16518 & n16519 ;
  assign n16521 = n8189 ^ n1056 ^ 1'b0 ;
  assign n16523 = n12557 ^ n2193 ^ 1'b0 ;
  assign n16524 = n3261 & ~n16523 ;
  assign n16525 = n16524 ^ n6640 ^ 1'b0 ;
  assign n16522 = n1278 & ~n2168 ;
  assign n16526 = n16525 ^ n16522 ^ 1'b0 ;
  assign n16527 = n7848 ^ n2890 ^ 1'b0 ;
  assign n16528 = n8987 ^ n6979 ^ 1'b0 ;
  assign n16529 = n456 | n16528 ;
  assign n16530 = n16527 | n16529 ;
  assign n16531 = ~n3187 & n11362 ;
  assign n16532 = n16531 ^ n2173 ^ 1'b0 ;
  assign n16533 = ~n535 & n1081 ;
  assign n16534 = n16533 ^ n13855 ^ n6742 ;
  assign n16535 = ~n4666 & n10799 ;
  assign n16536 = n8279 ^ n6288 ^ 1'b0 ;
  assign n16537 = n15101 ^ n12284 ^ 1'b0 ;
  assign n16538 = n5076 & ~n16537 ;
  assign n16539 = n7503 ^ n4531 ^ n3097 ;
  assign n16540 = n3734 & n16539 ;
  assign n16541 = n16538 & ~n16540 ;
  assign n16542 = n16536 & n16541 ;
  assign n16543 = n8905 | n9334 ;
  assign n16544 = n2250 | n6754 ;
  assign n16545 = ~n2056 & n6604 ;
  assign n16546 = n10811 & n16545 ;
  assign n16547 = n10158 & ~n14560 ;
  assign n16548 = n9488 & n16547 ;
  assign n16549 = n16548 ^ n14027 ^ n105 ;
  assign n16550 = ( n9399 & n16546 ) | ( n9399 & n16549 ) | ( n16546 & n16549 ) ;
  assign n16551 = n15550 & ~n16550 ;
  assign n16552 = n1534 & n16551 ;
  assign n16553 = n3136 & ~n4782 ;
  assign n16554 = ~n6892 & n16553 ;
  assign n16555 = n16554 ^ n1451 ^ 1'b0 ;
  assign n16556 = n11771 ^ n11394 ^ 1'b0 ;
  assign n16557 = n7549 ^ n3583 ^ 1'b0 ;
  assign n16558 = ~n7803 & n16557 ;
  assign n16559 = n16558 ^ n5881 ^ 1'b0 ;
  assign n16560 = n5604 | n8586 ;
  assign n16561 = n6542 ^ n4106 ^ 1'b0 ;
  assign n16563 = n12380 ^ n1182 ^ 1'b0 ;
  assign n16564 = n16563 ^ n4229 ^ 1'b0 ;
  assign n16562 = n7761 & n8879 ;
  assign n16565 = n16564 ^ n16562 ^ n333 ;
  assign n16566 = ~n12158 & n16565 ;
  assign n16567 = n6808 ^ n461 ^ 1'b0 ;
  assign n16568 = n7581 & n16567 ;
  assign n16569 = n16568 ^ n16256 ^ 1'b0 ;
  assign n16570 = n184 | n16569 ;
  assign n16571 = n8521 ^ n5809 ^ n4982 ;
  assign n16572 = n10480 ^ n5929 ^ 1'b0 ;
  assign n16573 = n16571 & ~n16572 ;
  assign n16574 = ~n1024 & n16573 ;
  assign n16575 = n16574 ^ n9082 ^ 1'b0 ;
  assign n16576 = n16554 ^ n8820 ^ 1'b0 ;
  assign n16577 = n5259 | n6491 ;
  assign n16578 = ~n2940 & n10109 ;
  assign n16579 = ~n16577 & n16578 ;
  assign n16580 = n1124 & n2181 ;
  assign n16581 = n16580 ^ n4732 ^ 1'b0 ;
  assign n16582 = ~n1058 & n2648 ;
  assign n16583 = n2403 & n11925 ;
  assign n16584 = n16582 & n16583 ;
  assign n16585 = ~n1024 & n4463 ;
  assign n16586 = n16584 & n16585 ;
  assign n16587 = n16586 ^ n4174 ^ 1'b0 ;
  assign n16588 = ~n7614 & n16587 ;
  assign n16589 = ~n15951 & n16588 ;
  assign n16590 = ~n16581 & n16589 ;
  assign n16594 = n4173 & ~n7659 ;
  assign n16595 = ~n5678 & n16594 ;
  assign n16592 = n13424 ^ n2708 ^ 1'b0 ;
  assign n16593 = ~n8171 & n16592 ;
  assign n16591 = n10829 | n14318 ;
  assign n16596 = n16595 ^ n16593 ^ n16591 ;
  assign n16597 = ~n1014 & n11869 ;
  assign n16598 = n7952 & n13753 ;
  assign n16599 = n1246 & n3512 ;
  assign n16600 = n16599 ^ n5379 ^ 1'b0 ;
  assign n16601 = n16600 ^ n7384 ^ 1'b0 ;
  assign n16602 = n9002 & ~n16601 ;
  assign n16607 = n12535 ^ n6831 ^ 1'b0 ;
  assign n16603 = n15152 ^ n6067 ^ n2664 ;
  assign n16604 = n5055 ^ n855 ^ 1'b0 ;
  assign n16605 = n16604 ^ n4040 ^ 1'b0 ;
  assign n16606 = n16603 & ~n16605 ;
  assign n16608 = n16607 ^ n16606 ^ n2663 ;
  assign n16609 = ( n2771 & n12165 ) | ( n2771 & ~n13108 ) | ( n12165 & ~n13108 ) ;
  assign n16610 = n5865 ^ n2943 ^ 1'b0 ;
  assign n16611 = ~n3713 & n8801 ;
  assign n16612 = n16611 ^ n4367 ^ 1'b0 ;
  assign n16613 = n304 | n910 ;
  assign n16614 = n6584 | n16613 ;
  assign n16615 = n16614 ^ n1941 ^ 1'b0 ;
  assign n16616 = ~n12662 & n16615 ;
  assign n16617 = n6917 & n16616 ;
  assign n16618 = n11243 & n11860 ;
  assign n16619 = n16618 ^ n8812 ^ 1'b0 ;
  assign n16620 = n11511 | n16619 ;
  assign n16621 = n16620 ^ n12185 ^ 1'b0 ;
  assign n16622 = ~n4039 & n5348 ;
  assign n16623 = ~n4079 & n16622 ;
  assign n16624 = n9459 | n16623 ;
  assign n16625 = n16624 ^ n8327 ^ 1'b0 ;
  assign n16626 = n5329 | n16625 ;
  assign n16627 = n14999 | n16626 ;
  assign n16628 = n12589 ^ n227 ^ 1'b0 ;
  assign n16629 = n982 | n16628 ;
  assign n16630 = n16629 ^ n13888 ^ 1'b0 ;
  assign n16631 = n3536 & n5726 ;
  assign n16632 = ~n16630 & n16631 ;
  assign n16634 = n2669 & n3013 ;
  assign n16635 = n7061 & n16634 ;
  assign n16636 = n16635 ^ n1466 ^ 1'b0 ;
  assign n16633 = n5831 ^ n3944 ^ 1'b0 ;
  assign n16637 = n16636 ^ n16633 ^ 1'b0 ;
  assign n16639 = n4859 | n6617 ;
  assign n16638 = n1069 & ~n6335 ;
  assign n16640 = n16639 ^ n16638 ^ 1'b0 ;
  assign n16641 = n14733 ^ n4510 ^ 1'b0 ;
  assign n16642 = n9322 | n16641 ;
  assign n16643 = n15196 & ~n16642 ;
  assign n16644 = n16643 ^ n2914 ^ 1'b0 ;
  assign n16645 = n3364 & n13897 ;
  assign n16646 = n10724 & ~n12365 ;
  assign n16647 = n16646 ^ n16536 ^ 1'b0 ;
  assign n16651 = n16536 ^ n3519 ^ 1'b0 ;
  assign n16648 = ~n105 & n3339 ;
  assign n16649 = n10462 ^ n8425 ^ 1'b0 ;
  assign n16650 = n16648 | n16649 ;
  assign n16652 = n16651 ^ n16650 ^ 1'b0 ;
  assign n16653 = n11065 & n16652 ;
  assign n16654 = n9949 ^ n4468 ^ n2772 ;
  assign n16655 = ~n4248 & n11193 ;
  assign n16656 = n16654 & n16655 ;
  assign n16657 = n6236 ^ n451 ^ 1'b0 ;
  assign n16658 = n15254 | n16657 ;
  assign n16659 = n16656 & ~n16658 ;
  assign n16660 = n15620 & n16659 ;
  assign n16661 = n3580 | n10638 ;
  assign n16662 = n3518 | n9088 ;
  assign n16663 = n14094 & ~n16662 ;
  assign n16664 = n16663 ^ n4083 ^ 1'b0 ;
  assign n16665 = n10837 & ~n16664 ;
  assign n16666 = n390 & n4879 ;
  assign n16667 = n3779 & ~n6445 ;
  assign n16668 = n3762 | n16667 ;
  assign n16669 = n16668 ^ n1832 ^ 1'b0 ;
  assign n16670 = n4251 ^ n511 ^ 1'b0 ;
  assign n16671 = ~n4993 & n15659 ;
  assign n16672 = n6915 | n13623 ;
  assign n16673 = n11927 ^ n5733 ^ 1'b0 ;
  assign n16674 = ~n8327 & n16673 ;
  assign n16675 = ( n885 & n1812 ) | ( n885 & ~n3823 ) | ( n1812 & ~n3823 ) ;
  assign n16676 = n16675 ^ n15348 ^ 1'b0 ;
  assign n16677 = n8607 & ~n14798 ;
  assign n16678 = n2906 | n13864 ;
  assign n16681 = n5728 | n7405 ;
  assign n16679 = n15513 ^ n3137 ^ 1'b0 ;
  assign n16680 = n12773 | n16679 ;
  assign n16682 = n16681 ^ n16680 ^ n11656 ;
  assign n16683 = ~n1284 & n2313 ;
  assign n16684 = n13326 ^ n9867 ^ 1'b0 ;
  assign n16685 = n9233 & n16684 ;
  assign n16686 = n16683 & n16685 ;
  assign n16687 = ~n14895 & n15964 ;
  assign n16688 = n11035 & n16687 ;
  assign n16689 = n11800 & ~n15025 ;
  assign n16690 = n5251 ^ n1852 ^ 1'b0 ;
  assign n16691 = ~n10278 & n16690 ;
  assign n16692 = n16691 ^ n15737 ^ 1'b0 ;
  assign n16693 = ~n12197 & n16692 ;
  assign n16694 = n1699 & ~n15622 ;
  assign n16695 = n16694 ^ n16286 ^ 1'b0 ;
  assign n16696 = n6937 ^ n5044 ^ 1'b0 ;
  assign n16697 = n7335 ^ n459 ^ 1'b0 ;
  assign n16698 = n3393 & n14234 ;
  assign n16699 = n16697 & n16698 ;
  assign n16700 = n6604 & ~n16699 ;
  assign n16701 = n16696 & n16700 ;
  assign n16702 = n15134 ^ n11394 ^ 1'b0 ;
  assign n16703 = n2100 ^ n835 ^ 1'b0 ;
  assign n16704 = n13370 & n16703 ;
  assign n16705 = ~n14657 & n16704 ;
  assign n16706 = n16705 ^ n16335 ^ n468 ;
  assign n16707 = n11183 ^ n1099 ^ 1'b0 ;
  assign n16708 = n13061 ^ n2756 ^ 1'b0 ;
  assign n16709 = n1554 & n16708 ;
  assign n16710 = n13254 ^ n12621 ^ 1'b0 ;
  assign n16711 = n16709 & n16710 ;
  assign n16712 = ~n3139 & n4687 ;
  assign n16713 = n16712 ^ n16130 ^ 1'b0 ;
  assign n16714 = n4365 | n16363 ;
  assign n16715 = n16640 ^ n12694 ^ 1'b0 ;
  assign n16716 = n16714 | n16715 ;
  assign n16717 = n9530 ^ n695 ^ 1'b0 ;
  assign n16718 = n6578 & n16717 ;
  assign n16719 = n1211 ^ n49 ^ 1'b0 ;
  assign n16720 = n9935 & ~n16719 ;
  assign n16721 = n9941 & ~n16720 ;
  assign n16724 = n4405 ^ n3299 ^ 1'b0 ;
  assign n16725 = n1090 & ~n16724 ;
  assign n16722 = n6931 | n11314 ;
  assign n16723 = n1473 & ~n16722 ;
  assign n16726 = n16725 ^ n16723 ^ 1'b0 ;
  assign n16727 = n9891 ^ n7220 ^ 1'b0 ;
  assign n16728 = n7357 & n15332 ;
  assign n16729 = n8163 & n16728 ;
  assign n16730 = n5067 & ~n7038 ;
  assign n16731 = n11776 | n16730 ;
  assign n16732 = n15298 ^ n1896 ^ n1703 ;
  assign n16733 = ~n590 & n8811 ;
  assign n16734 = ~n120 & n4740 ;
  assign n16735 = n16734 ^ n8481 ^ 1'b0 ;
  assign n16736 = n3250 | n16735 ;
  assign n16737 = n4329 & ~n14071 ;
  assign n16738 = n16737 ^ n2837 ^ 1'b0 ;
  assign n16739 = n8157 ^ n6878 ^ 1'b0 ;
  assign n16740 = n9698 | n16739 ;
  assign n16742 = n4504 & n13444 ;
  assign n16743 = n16742 ^ n582 ^ 1'b0 ;
  assign n16741 = n8770 & ~n14694 ;
  assign n16744 = n16743 ^ n16741 ^ 1'b0 ;
  assign n16745 = ~n13313 & n16744 ;
  assign n16746 = n7744 & n16745 ;
  assign n16747 = ~n12288 & n16746 ;
  assign n16748 = n14865 ^ n150 ^ 1'b0 ;
  assign n16749 = ~n16747 & n16748 ;
  assign n16752 = n13593 ^ n2843 ^ 1'b0 ;
  assign n16753 = n546 | n16752 ;
  assign n16750 = n43 & ~n2460 ;
  assign n16751 = ~n1889 & n16750 ;
  assign n16754 = n16753 ^ n16751 ^ 1'b0 ;
  assign n16755 = n6003 & ~n6166 ;
  assign n16756 = n9457 & n16755 ;
  assign n16757 = n16756 ^ n3748 ^ 1'b0 ;
  assign n16758 = n8216 ^ n6742 ^ 1'b0 ;
  assign n16759 = n1580 & n7602 ;
  assign n16760 = ~n16565 & n16759 ;
  assign n16761 = n16760 ^ n14352 ^ 1'b0 ;
  assign n16762 = ~n2634 & n16761 ;
  assign n16763 = n646 | n16088 ;
  assign n16764 = n5725 | n16763 ;
  assign n16765 = n577 ^ n296 ^ 1'b0 ;
  assign n16766 = n968 & n2693 ;
  assign n16767 = ~n2693 & n16766 ;
  assign n16768 = ( n2257 & n11009 ) | ( n2257 & ~n16213 ) | ( n11009 & ~n16213 ) ;
  assign n16776 = ( n666 & n2753 ) | ( n666 & ~n6660 ) | ( n2753 & ~n6660 ) ;
  assign n16777 = n16776 ^ n3095 ^ 1'b0 ;
  assign n16778 = n16777 ^ n4017 ^ 1'b0 ;
  assign n16779 = n2885 & n16778 ;
  assign n16780 = n16779 ^ n8275 ^ 1'b0 ;
  assign n16781 = ( ~n1543 & n2101 ) | ( ~n1543 & n3622 ) | ( n2101 & n3622 ) ;
  assign n16782 = n16781 ^ n3974 ^ 1'b0 ;
  assign n16783 = n6473 & n16782 ;
  assign n16784 = n5267 & n16783 ;
  assign n16785 = n16784 ^ n14502 ^ 1'b0 ;
  assign n16786 = n16780 | n16785 ;
  assign n16769 = ~n5064 & n5684 ;
  assign n16770 = n16769 ^ n9584 ^ 1'b0 ;
  assign n16771 = n12718 ^ n4707 ^ 1'b0 ;
  assign n16772 = n1785 & n16771 ;
  assign n16773 = n16772 ^ n4537 ^ 1'b0 ;
  assign n16774 = ~n1783 & n16773 ;
  assign n16775 = n16770 & n16774 ;
  assign n16787 = n16786 ^ n16775 ^ 1'b0 ;
  assign n16788 = n3042 & ~n5340 ;
  assign n16789 = ~n8003 & n16788 ;
  assign n16790 = ~n3795 & n16789 ;
  assign n16791 = n8342 & ~n16790 ;
  assign n16792 = n1265 ^ n1202 ^ 1'b0 ;
  assign n16793 = n5523 | n13573 ;
  assign n16794 = n8985 & n10826 ;
  assign n16795 = ~n2286 & n16794 ;
  assign n16796 = n1453 | n16795 ;
  assign n16797 = ~n116 & n3060 ;
  assign n16798 = n116 & n16797 ;
  assign n16799 = n3851 & ~n16798 ;
  assign n16800 = ~n16796 & n16799 ;
  assign n16801 = n9557 ^ n7685 ^ 1'b0 ;
  assign n16802 = n10484 & ~n16801 ;
  assign n16803 = n14499 ^ n4832 ^ 1'b0 ;
  assign n16804 = n16803 ^ n5016 ^ 1'b0 ;
  assign n16805 = ~n1853 & n2675 ;
  assign n16806 = n16805 ^ n13447 ^ 1'b0 ;
  assign n16807 = n16806 ^ n1717 ^ 1'b0 ;
  assign n16808 = n451 & ~n16807 ;
  assign n16809 = n5768 & ~n6218 ;
  assign n16810 = ( n1582 & n3704 ) | ( n1582 & ~n16809 ) | ( n3704 & ~n16809 ) ;
  assign n16811 = n2346 & ~n6591 ;
  assign n16812 = n3040 ^ n2678 ^ 1'b0 ;
  assign n16813 = ~n7812 & n16812 ;
  assign n16814 = n13578 ^ n12219 ^ 1'b0 ;
  assign n16815 = ~n6071 & n16814 ;
  assign n16816 = n16813 & n16815 ;
  assign n16817 = n16816 ^ n8876 ^ 1'b0 ;
  assign n16818 = n7259 & ~n7967 ;
  assign n16819 = n8225 & n16818 ;
  assign n16820 = n6763 | n16819 ;
  assign n16821 = n13416 | n15442 ;
  assign n16822 = n9397 ^ n6318 ^ 1'b0 ;
  assign n16823 = ~n16477 & n16822 ;
  assign n16824 = n8899 ^ n7389 ^ n3350 ;
  assign n16825 = n3414 & n16824 ;
  assign n16826 = ~n1103 & n11840 ;
  assign n16827 = n15768 & n16826 ;
  assign n16828 = n16734 ^ n8299 ^ 1'b0 ;
  assign n16829 = ~n7626 & n16828 ;
  assign n16830 = n2092 | n16654 ;
  assign n16831 = n16830 ^ n1018 ^ 1'b0 ;
  assign n16832 = n9231 ^ n1323 ^ x5 ;
  assign n16833 = n6622 | n16832 ;
  assign n16834 = n16833 ^ n2272 ^ 1'b0 ;
  assign n16835 = ~n16831 & n16834 ;
  assign n16836 = n2283 | n5671 ;
  assign n16837 = n1212 & ~n16836 ;
  assign n16838 = n16837 ^ n13891 ^ n12877 ;
  assign n16839 = n404 & n13193 ;
  assign n16840 = n6836 & n16839 ;
  assign n16841 = n2275 & ~n3384 ;
  assign n16842 = n6080 & ~n16841 ;
  assign n16843 = n7164 ^ n6681 ^ 1'b0 ;
  assign n16844 = n2034 & ~n3670 ;
  assign n16845 = n8312 ^ n5165 ^ 1'b0 ;
  assign n16846 = n15563 & ~n16845 ;
  assign n16847 = n16846 ^ n6411 ^ n1430 ;
  assign n16848 = n3243 | n10553 ;
  assign n16849 = n16848 ^ n6296 ^ 1'b0 ;
  assign n16850 = n4928 ^ n968 ^ 1'b0 ;
  assign n16851 = n5915 ^ n722 ^ 1'b0 ;
  assign n16852 = n16851 ^ n10093 ^ 1'b0 ;
  assign n16853 = n6604 & n16852 ;
  assign n16854 = n8026 & n8413 ;
  assign n16855 = ~n5986 & n9799 ;
  assign n16856 = n10825 & n16855 ;
  assign n16857 = n16197 ^ n6747 ^ 1'b0 ;
  assign n16858 = n10231 | n16857 ;
  assign n16859 = n15054 | n16858 ;
  assign n16860 = n14510 ^ n7071 ^ n597 ;
  assign n16861 = ~n673 & n2926 ;
  assign n16862 = n16861 ^ n3562 ^ 1'b0 ;
  assign n16863 = n16860 & n16862 ;
  assign n16864 = n1355 & ~n11782 ;
  assign n16865 = n16864 ^ n4681 ^ 1'b0 ;
  assign n16866 = n1578 & n10317 ;
  assign n16867 = n16866 ^ n255 ^ 1'b0 ;
  assign n16868 = n15050 & n16867 ;
  assign n16869 = n4294 & n16868 ;
  assign n16870 = n7846 ^ n2812 ^ n1182 ;
  assign n16871 = n5970 & n16870 ;
  assign n16872 = ~n861 & n3890 ;
  assign n16873 = n2445 & ~n12284 ;
  assign n16874 = n16873 ^ n10404 ^ 1'b0 ;
  assign n16875 = n16874 ^ n11238 ^ 1'b0 ;
  assign n16876 = ~n16872 & n16875 ;
  assign n16877 = ~n13089 & n16876 ;
  assign n16878 = ~n16871 & n16877 ;
  assign n16879 = n13697 ^ n3768 ^ 1'b0 ;
  assign n16880 = n5152 | n16879 ;
  assign n16881 = n4160 ^ n3276 ^ 1'b0 ;
  assign n16882 = n9325 ^ n83 ^ 1'b0 ;
  assign n16883 = n1466 & n13585 ;
  assign n16884 = n3155 | n7849 ;
  assign n16885 = n14744 ^ n11035 ^ 1'b0 ;
  assign n16886 = ~n16884 & n16885 ;
  assign n16887 = ~n11360 & n16886 ;
  assign n16888 = ( n1724 & n7804 ) | ( n1724 & n9368 ) | ( n7804 & n9368 ) ;
  assign n16889 = n8960 ^ n5710 ^ 1'b0 ;
  assign n16890 = n1395 & ~n8076 ;
  assign n16891 = ~n3139 & n8933 ;
  assign n16892 = n14008 ^ n3583 ^ 1'b0 ;
  assign n16893 = n16891 | n16892 ;
  assign n16894 = n931 & ~n16893 ;
  assign n16895 = n2794 ^ n133 ^ 1'b0 ;
  assign n16896 = ~n1143 & n16895 ;
  assign n16900 = n2039 | n3438 ;
  assign n16901 = n6084 | n16900 ;
  assign n16902 = n16901 ^ n1993 ^ 1'b0 ;
  assign n16903 = ( ~n2570 & n6542 ) | ( ~n2570 & n16902 ) | ( n6542 & n16902 ) ;
  assign n16904 = ~n6651 & n16903 ;
  assign n16905 = n16904 ^ n2605 ^ 1'b0 ;
  assign n16897 = n9113 ^ n5184 ^ 1'b0 ;
  assign n16898 = n6065 | n16897 ;
  assign n16899 = n12458 | n16898 ;
  assign n16906 = n16905 ^ n16899 ^ 1'b0 ;
  assign n16907 = n16896 & n16906 ;
  assign n16908 = n15016 & n16907 ;
  assign n16909 = n9689 ^ n2427 ^ 1'b0 ;
  assign n16910 = ~n1726 & n3736 ;
  assign n16911 = n1989 | n16910 ;
  assign n16912 = n16911 ^ n16669 ^ 1'b0 ;
  assign n16913 = n16912 ^ n11771 ^ 1'b0 ;
  assign n16914 = n16913 ^ n13600 ^ 1'b0 ;
  assign n16915 = n16909 & ~n16914 ;
  assign n16916 = n3705 | n11041 ;
  assign n16917 = n6048 & n7348 ;
  assign n16918 = ~n6915 & n16917 ;
  assign n16919 = n56 & n2448 ;
  assign n16920 = n16919 ^ n3372 ^ 1'b0 ;
  assign n16921 = n16920 ^ n1283 ^ 1'b0 ;
  assign n16922 = n8761 & n16921 ;
  assign n16923 = n16657 ^ n1569 ^ 1'b0 ;
  assign n16924 = n16923 ^ n10491 ^ 1'b0 ;
  assign n16925 = n3264 & n3361 ;
  assign n16926 = n9922 ^ n1745 ^ 1'b0 ;
  assign n16927 = n16926 ^ n12496 ^ 1'b0 ;
  assign n16928 = ~n16925 & n16927 ;
  assign n16929 = ~n2155 & n10459 ;
  assign n16930 = n16929 ^ n14749 ^ 1'b0 ;
  assign n16931 = n16096 | n16930 ;
  assign n16932 = n9513 | n16931 ;
  assign n16933 = n4563 | n16932 ;
  assign n16934 = n1717 | n7170 ;
  assign n16935 = n16934 ^ n5959 ^ 1'b0 ;
  assign n16936 = n4254 & ~n16935 ;
  assign n16937 = n6644 ^ n1152 ^ 1'b0 ;
  assign n16938 = n1825 & n16937 ;
  assign n16939 = n16938 ^ n6925 ^ 1'b0 ;
  assign n16940 = n5348 ^ n488 ^ 1'b0 ;
  assign n16942 = n7316 & n10237 ;
  assign n16941 = n1007 & n3674 ;
  assign n16943 = n16942 ^ n16941 ^ n7756 ;
  assign n16944 = n16943 ^ n8097 ^ 1'b0 ;
  assign n16945 = n16940 & n16944 ;
  assign n16946 = n15915 ^ n15707 ^ 1'b0 ;
  assign n16947 = n11309 ^ n8537 ^ 1'b0 ;
  assign n16948 = n5209 & ~n6316 ;
  assign n16949 = n16948 ^ n456 ^ 1'b0 ;
  assign n16950 = n1235 & n16949 ;
  assign n16951 = n4599 & n6785 ;
  assign n16952 = n8919 ^ n3219 ^ 1'b0 ;
  assign n16953 = n6656 & n16952 ;
  assign n16954 = n16953 ^ n1491 ^ 1'b0 ;
  assign n16955 = n10840 & ~n15075 ;
  assign n16956 = n16955 ^ n16391 ^ 1'b0 ;
  assign n16957 = n9808 ^ n2883 ^ 1'b0 ;
  assign n16958 = n9274 ^ n2070 ^ 1'b0 ;
  assign n16959 = ~n16957 & n16958 ;
  assign n16960 = ~n8720 & n11701 ;
  assign n16961 = n13 & n5069 ;
  assign n16962 = n12518 & n16961 ;
  assign n16963 = n10610 ^ n9161 ^ n368 ;
  assign n16964 = n15777 ^ n3442 ^ 1'b0 ;
  assign n16965 = ~n1652 & n16964 ;
  assign n16966 = ~n269 & n16965 ;
  assign n16967 = n432 & n5274 ;
  assign n16968 = n16967 ^ n2826 ^ 1'b0 ;
  assign n16969 = n4804 | n16968 ;
  assign n16970 = n1371 & n12153 ;
  assign n16971 = n16970 ^ n3529 ^ 1'b0 ;
  assign n16972 = n1695 & n16971 ;
  assign n16973 = n3867 & ~n12201 ;
  assign n16974 = n16972 & n16973 ;
  assign n16975 = n16974 ^ n16740 ^ n1812 ;
  assign n16976 = n14301 ^ n205 ^ 1'b0 ;
  assign n16977 = n609 & ~n835 ;
  assign n16978 = n5930 & n16977 ;
  assign n16979 = n16978 ^ n11627 ^ 1'b0 ;
  assign n16980 = n7170 & n16979 ;
  assign n16981 = ~n9087 & n9266 ;
  assign n16982 = ~n2382 & n9720 ;
  assign n16983 = n16981 & n16982 ;
  assign n16984 = n4146 & ~n5005 ;
  assign n16985 = n5990 ^ n4495 ^ 1'b0 ;
  assign n16986 = ( n14478 & n16801 ) | ( n14478 & ~n16985 ) | ( n16801 & ~n16985 ) ;
  assign n16987 = ~n5497 & n16986 ;
  assign n16988 = n2355 & n3713 ;
  assign n16989 = n365 & ~n11469 ;
  assign n16990 = n16989 ^ n3462 ^ 1'b0 ;
  assign n16991 = ~n16988 & n16990 ;
  assign n16992 = n259 & n16991 ;
  assign n16994 = n3738 ^ n3412 ^ 1'b0 ;
  assign n16995 = n1968 & n16994 ;
  assign n16993 = n5967 & n14420 ;
  assign n16996 = n16995 ^ n16993 ^ 1'b0 ;
  assign n16997 = n10400 ^ n9288 ^ 1'b0 ;
  assign n16998 = n2529 | n16997 ;
  assign n16999 = n3859 & ~n16998 ;
  assign n17000 = ~n5513 & n16268 ;
  assign n17001 = n809 | n11027 ;
  assign n17002 = n10893 ^ n135 ^ 1'b0 ;
  assign n17003 = n266 | n1136 ;
  assign n17004 = n13251 & ~n17003 ;
  assign n17005 = n17004 ^ n1438 ^ 1'b0 ;
  assign n17006 = n10621 ^ n2290 ^ 1'b0 ;
  assign n17007 = ~n2584 & n17006 ;
  assign n17008 = ~n1390 & n4612 ;
  assign n17009 = ~n14350 & n17008 ;
  assign n17010 = ~n1118 & n17009 ;
  assign n17011 = n13203 & n16876 ;
  assign n17012 = n16884 ^ n14375 ^ 1'b0 ;
  assign n17013 = ~n14348 & n14937 ;
  assign n17014 = n7126 ^ n1960 ^ 1'b0 ;
  assign n17015 = ( n582 & n4788 ) | ( n582 & n6311 ) | ( n4788 & n6311 ) ;
  assign n17016 = n13285 & ~n15196 ;
  assign n17017 = n5890 & n17016 ;
  assign n17018 = n2087 & n5921 ;
  assign n17019 = n17017 & n17018 ;
  assign n17020 = n17019 ^ n1288 ^ 1'b0 ;
  assign n17021 = n5813 | n17020 ;
  assign n17022 = n7708 ^ n1635 ^ 1'b0 ;
  assign n17023 = n17022 ^ n14883 ^ n376 ;
  assign n17024 = n16373 ^ n263 ^ 1'b0 ;
  assign n17025 = n8376 ^ n6591 ^ n192 ;
  assign n17026 = n10670 ^ n263 ^ 1'b0 ;
  assign n17027 = n8414 & n17026 ;
  assign n17028 = n17025 & ~n17027 ;
  assign n17029 = n3775 & n7107 ;
  assign n17030 = n17029 ^ n4981 ^ 1'b0 ;
  assign n17031 = ~n9424 & n17030 ;
  assign n17032 = n17031 ^ n11805 ^ 1'b0 ;
  assign n17033 = n12214 & n17032 ;
  assign n17034 = n17028 & n17033 ;
  assign n17035 = n1312 & n4846 ;
  assign n17036 = n17035 ^ n11189 ^ 1'b0 ;
  assign n17037 = n12412 ^ n1068 ^ 1'b0 ;
  assign n17038 = ~n17036 & n17037 ;
  assign n17039 = ~n77 & n241 ;
  assign n17040 = n17039 ^ n8693 ^ 1'b0 ;
  assign n17041 = ~n2950 & n3248 ;
  assign n17042 = ~n10031 & n17041 ;
  assign n17043 = n12740 ^ n2092 ^ 1'b0 ;
  assign n17044 = n582 & n10288 ;
  assign n17045 = n8139 ^ n3068 ^ 1'b0 ;
  assign n17046 = n270 & ~n13375 ;
  assign n17047 = ~n8683 & n17046 ;
  assign n17048 = n576 & n7958 ;
  assign n17049 = n17048 ^ n9281 ^ 1'b0 ;
  assign n17050 = ~n17047 & n17049 ;
  assign n17051 = n183 | n5139 ;
  assign n17052 = n6079 & n17051 ;
  assign n17053 = n17052 ^ n14053 ^ 1'b0 ;
  assign n17054 = n17050 & ~n17053 ;
  assign n17055 = n15147 ^ n7382 ^ 1'b0 ;
  assign n17056 = n11400 & n17055 ;
  assign n17057 = n2332 & n17056 ;
  assign n17058 = ~n451 & n6740 ;
  assign n17059 = n17058 ^ n8182 ^ 1'b0 ;
  assign n17060 = ~n10342 & n11479 ;
  assign n17061 = n17059 & n17060 ;
  assign n17062 = n2228 ^ n51 ^ 1'b0 ;
  assign n17063 = n16758 & n17062 ;
  assign n17064 = ~n2955 & n11070 ;
  assign n17065 = ~n6935 & n7924 ;
  assign n17066 = n17065 ^ n12664 ^ 1'b0 ;
  assign n17067 = n11266 ^ n8637 ^ 1'b0 ;
  assign n17068 = n16511 | n17067 ;
  assign n17069 = n1258 & n1484 ;
  assign n17070 = n17069 ^ n2030 ^ 1'b0 ;
  assign n17071 = ~n1792 & n11710 ;
  assign n17072 = n17071 ^ n4914 ^ 1'b0 ;
  assign n17073 = n1868 & ~n17072 ;
  assign n17074 = n17073 ^ n9526 ^ 1'b0 ;
  assign n17075 = n7873 ^ n2387 ^ 1'b0 ;
  assign n17076 = n2340 | n17075 ;
  assign n17077 = n17076 ^ n14790 ^ 1'b0 ;
  assign n17078 = n17077 ^ n7242 ^ n1077 ;
  assign n17079 = ~n4087 & n17078 ;
  assign n17080 = n7194 & ~n10196 ;
  assign n17081 = n14694 ^ n9769 ^ 1'b0 ;
  assign n17082 = ~n841 & n2686 ;
  assign n17083 = n17082 ^ n884 ^ 1'b0 ;
  assign n17084 = ~n6589 & n17083 ;
  assign n17085 = n10686 | n17084 ;
  assign n17086 = ~n5592 & n9057 ;
  assign n17087 = n12625 ^ n1271 ^ 1'b0 ;
  assign n17088 = n17087 ^ n11797 ^ 1'b0 ;
  assign n17089 = n17088 ^ n924 ^ 1'b0 ;
  assign n17090 = n10126 & ~n17089 ;
  assign n17091 = n9056 ^ n6084 ^ 1'b0 ;
  assign n17092 = ~n13717 & n17091 ;
  assign n17093 = n5081 & n6866 ;
  assign n17094 = n17093 ^ n8909 ^ 1'b0 ;
  assign n17095 = ( n10584 & ~n13994 ) | ( n10584 & n17094 ) | ( ~n13994 & n17094 ) ;
  assign n17096 = n2048 | n2062 ;
  assign n17097 = n3166 | n17096 ;
  assign n17098 = ( n8061 & n13922 ) | ( n8061 & ~n17097 ) | ( n13922 & ~n17097 ) ;
  assign n17099 = n5086 & ~n10768 ;
  assign n17100 = n17099 ^ n1883 ^ 1'b0 ;
  assign n17101 = n5081 ^ n1783 ^ 1'b0 ;
  assign n17102 = n9280 | n17101 ;
  assign n17103 = n13349 & ~n14268 ;
  assign n17104 = n5072 | n16353 ;
  assign n17105 = n5253 | n17104 ;
  assign n17106 = n17105 ^ n4740 ^ 1'b0 ;
  assign n17107 = n841 | n3335 ;
  assign n17108 = n302 & ~n17107 ;
  assign n17109 = ~n5663 & n17108 ;
  assign n17110 = n8612 & n17109 ;
  assign n17111 = n7941 ^ n7316 ^ 1'b0 ;
  assign n17112 = ~n17110 & n17111 ;
  assign n17113 = n13283 ^ n61 ^ 1'b0 ;
  assign n17114 = n12972 & n17113 ;
  assign n17115 = n401 & ~n4823 ;
  assign n17116 = n17115 ^ n5176 ^ 1'b0 ;
  assign n17117 = ~n4197 & n17116 ;
  assign n17118 = n17114 | n17117 ;
  assign n17119 = n17112 & ~n17118 ;
  assign n17120 = n10124 & n17119 ;
  assign n17121 = n10488 & ~n17120 ;
  assign n17122 = ( ~n2717 & n12415 ) | ( ~n2717 & n13664 ) | ( n12415 & n13664 ) ;
  assign n17123 = ~n4937 & n9117 ;
  assign n17124 = n3461 & ~n17123 ;
  assign n17125 = n7382 | n9904 ;
  assign n17126 = n12784 & ~n17125 ;
  assign n17127 = n13283 ^ n8958 ^ 1'b0 ;
  assign n17128 = n10003 & n17127 ;
  assign n17129 = n3682 & ~n6623 ;
  assign n17130 = n14039 ^ n10041 ^ n7095 ;
  assign n17131 = ~n181 & n17130 ;
  assign n17132 = n12363 ^ n1493 ^ n88 ;
  assign n17133 = n13767 ^ n5484 ^ n3073 ;
  assign n17134 = ~n4290 & n17133 ;
  assign n17135 = ~n1167 & n1667 ;
  assign n17136 = n12389 ^ n10441 ^ 1'b0 ;
  assign n17137 = n17136 ^ n9953 ^ 1'b0 ;
  assign n17138 = n17135 & n17137 ;
  assign n17139 = ~n7482 & n17138 ;
  assign n17140 = n12677 ^ n1666 ^ 1'b0 ;
  assign n17141 = n9929 ^ n1788 ^ 1'b0 ;
  assign n17142 = ~n3003 & n6291 ;
  assign n17143 = n17142 ^ n1841 ^ 1'b0 ;
  assign n17144 = n10601 & ~n17143 ;
  assign n17145 = ( n8448 & ~n17141 ) | ( n8448 & n17144 ) | ( ~n17141 & n17144 ) ;
  assign n17146 = n8054 ^ n1669 ^ 1'b0 ;
  assign n17147 = ~n8830 & n10642 ;
  assign n17148 = ~n16303 & n17147 ;
  assign n17149 = n4587 & ~n6479 ;
  assign n17150 = n2498 & n17149 ;
  assign n17151 = n11946 ^ n7397 ^ 1'b0 ;
  assign n17152 = n17151 ^ n4675 ^ 1'b0 ;
  assign n17153 = ~n15080 & n17152 ;
  assign n17154 = n2507 & n16314 ;
  assign n17155 = n3724 & n17154 ;
  assign n17156 = n1385 & ~n15387 ;
  assign n17157 = n1381 & n2377 ;
  assign n17158 = n7965 ^ n307 ^ 1'b0 ;
  assign n17159 = n3966 | n17158 ;
  assign n17160 = n17159 ^ n3951 ^ 1'b0 ;
  assign n17161 = ~n3912 & n7303 ;
  assign n17162 = n801 & n17161 ;
  assign n17163 = n6281 & ~n17162 ;
  assign n17164 = n17163 ^ n14668 ^ 1'b0 ;
  assign n17165 = ~n2583 & n7529 ;
  assign n17166 = n16409 ^ n58 ^ 1'b0 ;
  assign n17167 = ~n433 & n17166 ;
  assign n17168 = n17167 ^ n3716 ^ 1'b0 ;
  assign n17169 = n8177 & n17168 ;
  assign n17170 = ( ~n54 & n1312 ) | ( ~n54 & n1568 ) | ( n1312 & n1568 ) ;
  assign n17171 = n16772 | n17170 ;
  assign n17172 = n5181 & ~n9519 ;
  assign n17173 = n4079 & ~n17172 ;
  assign n17174 = n15879 & n17173 ;
  assign n17175 = n6550 ^ n49 ^ 1'b0 ;
  assign n17176 = n16386 ^ n3459 ^ n1327 ;
  assign n17177 = n17176 ^ n10877 ^ 1'b0 ;
  assign n17178 = ~n7463 & n9112 ;
  assign n17179 = n17178 ^ n4639 ^ 1'b0 ;
  assign n17180 = n17177 | n17179 ;
  assign n17181 = ( n2531 & n4446 ) | ( n2531 & ~n6680 ) | ( n4446 & ~n6680 ) ;
  assign n17182 = n17181 ^ n12701 ^ n3280 ;
  assign n17183 = n13697 & ~n17182 ;
  assign n17184 = n14751 ^ n3371 ^ 1'b0 ;
  assign n17185 = ( ~n1878 & n1914 ) | ( ~n1878 & n10381 ) | ( n1914 & n10381 ) ;
  assign n17186 = n10489 ^ n304 ^ 1'b0 ;
  assign n17187 = n3113 | n17186 ;
  assign n17190 = n15537 ^ n1189 ^ 1'b0 ;
  assign n17191 = n17190 ^ n13185 ^ 1'b0 ;
  assign n17188 = n11073 & ~n14529 ;
  assign n17189 = n17188 ^ n870 ^ 1'b0 ;
  assign n17192 = n17191 ^ n17189 ^ 1'b0 ;
  assign n17193 = n10621 & n17192 ;
  assign n17194 = n1745 | n4765 ;
  assign n17195 = n17194 ^ n8852 ^ 1'b0 ;
  assign n17196 = n747 | n17195 ;
  assign n17197 = n8186 | n17196 ;
  assign n17198 = n8523 & n17197 ;
  assign n17199 = n1842 & n3759 ;
  assign n17200 = n1745 & ~n3181 ;
  assign n17201 = ~n3744 & n17200 ;
  assign n17202 = n3833 & ~n8138 ;
  assign n17203 = ~n8087 & n17202 ;
  assign n17204 = n5881 & ~n6656 ;
  assign n17205 = n1660 & ~n3618 ;
  assign n17206 = n17205 ^ n10076 ^ 1'b0 ;
  assign n17207 = n4903 & n17206 ;
  assign n17208 = ~n108 & n8710 ;
  assign n17219 = ~n3003 & n7322 ;
  assign n17209 = n315 & ~n1295 ;
  assign n17210 = ~n10758 & n17209 ;
  assign n17211 = n4187 & n17210 ;
  assign n17212 = n3823 ^ n856 ^ 1'b0 ;
  assign n17213 = ~n9444 & n17212 ;
  assign n17214 = n448 & ~n15389 ;
  assign n17215 = n17213 & n17214 ;
  assign n17216 = n17215 ^ n478 ^ 1'b0 ;
  assign n17217 = n11034 | n17216 ;
  assign n17218 = n17211 | n17217 ;
  assign n17220 = n17219 ^ n17218 ^ 1'b0 ;
  assign n17221 = n1958 | n10477 ;
  assign n17222 = n4735 & n17221 ;
  assign n17223 = n6437 & n17222 ;
  assign n17224 = n17223 ^ n8239 ^ 1'b0 ;
  assign n17225 = ~n188 & n579 ;
  assign n17226 = n17224 & n17225 ;
  assign n17227 = ~n4434 & n8037 ;
  assign n17228 = n17227 ^ n1069 ^ 1'b0 ;
  assign n17229 = ( ~n1223 & n4550 ) | ( ~n1223 & n12583 ) | ( n4550 & n12583 ) ;
  assign n17230 = n17229 ^ n6396 ^ 1'b0 ;
  assign n17231 = ~n4698 & n15651 ;
  assign n17232 = n14128 | n17231 ;
  assign n17233 = ~n2639 & n8359 ;
  assign n17234 = n3584 ^ n1481 ^ 1'b0 ;
  assign n17235 = n9405 & ~n17234 ;
  assign n17236 = n4619 & n7233 ;
  assign n17237 = n8026 & n17236 ;
  assign n17238 = n5801 | n6461 ;
  assign n17239 = n17238 ^ n10890 ^ 1'b0 ;
  assign n17240 = n10675 & ~n17239 ;
  assign n17241 = n17240 ^ n1904 ^ 1'b0 ;
  assign n17242 = n17241 ^ n7836 ^ 1'b0 ;
  assign n17245 = n3891 | n12287 ;
  assign n17243 = ~n1307 & n4016 ;
  assign n17244 = n17243 ^ n13545 ^ 1'b0 ;
  assign n17246 = n17245 ^ n17244 ^ n14200 ;
  assign n17247 = n12314 ^ n1109 ^ 1'b0 ;
  assign n17248 = n9564 & ~n17247 ;
  assign n17249 = n13925 | n17248 ;
  assign n17250 = n1161 | n7967 ;
  assign n17251 = n7326 & ~n17250 ;
  assign n17252 = n14456 | n17251 ;
  assign n17253 = n17252 ^ n13583 ^ 1'b0 ;
  assign n17254 = n229 & n12150 ;
  assign n17255 = n2833 & n5003 ;
  assign n17256 = n17255 ^ n8057 ^ 1'b0 ;
  assign n17257 = ( n7562 & n13758 ) | ( n7562 & n17256 ) | ( n13758 & n17256 ) ;
  assign n17258 = n12162 & ~n17257 ;
  assign n17259 = n7022 & ~n12305 ;
  assign n17260 = n15325 ^ n7961 ^ 1'b0 ;
  assign n17261 = n17260 ^ n9825 ^ 1'b0 ;
  assign n17262 = ~n15190 & n17261 ;
  assign n17263 = n17262 ^ n13041 ^ 1'b0 ;
  assign n17264 = n11243 & ~n17263 ;
  assign n17265 = ~n1212 & n10590 ;
  assign n17266 = ( n10696 & ~n15279 ) | ( n10696 & n17265 ) | ( ~n15279 & n17265 ) ;
  assign n17267 = n16012 ^ n12625 ^ 1'b0 ;
  assign n17268 = n14122 | n17267 ;
  assign n17269 = n2873 & ~n14663 ;
  assign n17270 = n3375 & n17269 ;
  assign n17271 = ~n61 & n17270 ;
  assign n17272 = n17271 ^ n17118 ^ 1'b0 ;
  assign n17273 = n8263 ^ n3690 ^ 1'b0 ;
  assign n17274 = n1029 & ~n17273 ;
  assign n17275 = ( n4201 & n4616 ) | ( n4201 & ~n7383 ) | ( n4616 & ~n7383 ) ;
  assign n17276 = n17275 ^ n8355 ^ n209 ;
  assign n17277 = n760 & n17276 ;
  assign n17278 = n17277 ^ n8034 ^ 1'b0 ;
  assign n17283 = n6102 ^ n5587 ^ n1809 ;
  assign n17284 = n17283 ^ n5444 ^ 1'b0 ;
  assign n17279 = n2943 & ~n13238 ;
  assign n17280 = n8456 & n17279 ;
  assign n17281 = ( ~n9507 & n14024 ) | ( ~n9507 & n17280 ) | ( n14024 & n17280 ) ;
  assign n17282 = ~n16337 & n17281 ;
  assign n17285 = n17284 ^ n17282 ^ 1'b0 ;
  assign n17286 = n8315 ^ n7589 ^ 1'b0 ;
  assign n17287 = n3099 & ~n17286 ;
  assign n17289 = ~n7787 & n10592 ;
  assign n17290 = n17289 ^ n12718 ^ 1'b0 ;
  assign n17288 = n841 & ~n5526 ;
  assign n17291 = n17290 ^ n17288 ^ 1'b0 ;
  assign n17292 = n10414 & n14099 ;
  assign n17293 = ~n17291 & n17292 ;
  assign n17294 = n12417 ^ n1031 ^ 1'b0 ;
  assign n17295 = n5821 | n17294 ;
  assign n17296 = ~n5893 & n7418 ;
  assign n17297 = n218 & n17296 ;
  assign n17298 = n17297 ^ n2101 ^ 1'b0 ;
  assign n17299 = n4920 & n6925 ;
  assign n17300 = ~n11909 & n17299 ;
  assign n17301 = n8399 ^ n4956 ^ n3646 ;
  assign n17302 = n17300 | n17301 ;
  assign n17303 = n17298 | n17302 ;
  assign n17304 = n1889 | n9797 ;
  assign n17305 = n16046 | n17304 ;
  assign n17306 = n17305 ^ n5420 ^ 1'b0 ;
  assign n17307 = n1712 & ~n3705 ;
  assign n17308 = ~n2101 & n17307 ;
  assign n17309 = n11052 | n17308 ;
  assign n17310 = n2807 | n10717 ;
  assign n17311 = n17310 ^ n4817 ^ 1'b0 ;
  assign n17312 = n17309 & n17311 ;
  assign n17313 = n3877 ^ n2694 ^ 1'b0 ;
  assign n17314 = n7879 | n12171 ;
  assign n17315 = n6039 ^ n4572 ^ 1'b0 ;
  assign n17316 = ~n1073 & n17315 ;
  assign n17317 = ~n4935 & n17316 ;
  assign n17318 = n17317 ^ n307 ^ 1'b0 ;
  assign n17319 = n17318 ^ n4425 ^ 1'b0 ;
  assign n17320 = n4335 ^ n2588 ^ 1'b0 ;
  assign n17321 = n8792 & ~n17320 ;
  assign n17322 = n17319 & ~n17321 ;
  assign n17323 = n17322 ^ n15582 ^ 1'b0 ;
  assign n17324 = n7967 ^ n1765 ^ 1'b0 ;
  assign n17325 = ( ~n5277 & n7562 ) | ( ~n5277 & n17324 ) | ( n7562 & n17324 ) ;
  assign n17326 = ~n1685 & n17325 ;
  assign n17327 = n8246 & ~n17326 ;
  assign n17328 = n15643 ^ n5695 ^ 1'b0 ;
  assign n17329 = n10212 & ~n17328 ;
  assign n17330 = n17329 ^ n14546 ^ n4781 ;
  assign n17331 = n9276 ^ n1293 ^ 1'b0 ;
  assign n17332 = ~n445 & n3012 ;
  assign n17333 = n17332 ^ n14883 ^ 1'b0 ;
  assign n17334 = n1073 & ~n1176 ;
  assign n17335 = n17334 ^ n1573 ^ 1'b0 ;
  assign n17336 = ~n14560 & n17335 ;
  assign n17337 = n16193 ^ n3489 ^ n132 ;
  assign n17338 = n17337 ^ n8134 ^ 1'b0 ;
  assign n17339 = n220 | n9777 ;
  assign n17340 = n1914 & ~n6865 ;
  assign n17341 = n17340 ^ n3334 ^ 1'b0 ;
  assign n17342 = n1269 | n17341 ;
  assign n17343 = n17342 ^ n14425 ^ 1'b0 ;
  assign n17344 = n1539 | n15905 ;
  assign n17345 = n17344 ^ n4173 ^ 1'b0 ;
  assign n17346 = n1584 & ~n2283 ;
  assign n17347 = n17346 ^ n12989 ^ 1'b0 ;
  assign n17348 = n15061 & n17347 ;
  assign n17349 = n5383 ^ n1023 ^ 1'b0 ;
  assign n17350 = n7715 & n17349 ;
  assign n17351 = n2925 & n17350 ;
  assign n17352 = n17351 ^ n12908 ^ 1'b0 ;
  assign n17353 = n2807 & ~n13790 ;
  assign n17354 = n17353 ^ n4946 ^ n4345 ;
  assign n17355 = n16388 & ~n17354 ;
  assign n17356 = n7105 | n9623 ;
  assign n17357 = n16599 & ~n17356 ;
  assign n17358 = n14385 ^ n135 ^ 1'b0 ;
  assign n17359 = n3595 | n17358 ;
  assign n17360 = n7329 | n17359 ;
  assign n17361 = n8503 ^ n4641 ^ n2321 ;
  assign n17362 = n17361 ^ n12406 ^ 1'b0 ;
  assign n17363 = n5214 | n17362 ;
  assign n17364 = n9451 ^ n2995 ^ 1'b0 ;
  assign n17365 = n3558 & n17364 ;
  assign n17366 = ~n3775 & n17365 ;
  assign n17367 = n11529 | n17366 ;
  assign n17368 = ~n1215 & n2067 ;
  assign n17369 = n8960 ^ n1336 ^ n133 ;
  assign n17370 = n4408 ^ n4155 ^ 1'b0 ;
  assign n17371 = n14741 | n17370 ;
  assign n17372 = n17369 | n17371 ;
  assign n17373 = ( ~n9399 & n10315 ) | ( ~n9399 & n17372 ) | ( n10315 & n17372 ) ;
  assign n17374 = x6 & n17373 ;
  assign n17375 = n17374 ^ n572 ^ 1'b0 ;
  assign n17376 = n6926 | n15273 ;
  assign n17377 = n17376 ^ n7739 ^ 1'b0 ;
  assign n17378 = ~n4402 & n10146 ;
  assign n17379 = n16999 ^ n845 ^ n395 ;
  assign n17380 = n9941 ^ n4790 ^ n1386 ;
  assign n17381 = n3899 & ~n8071 ;
  assign n17382 = n17380 & n17381 ;
  assign n17383 = n5219 & ~n17382 ;
  assign n17384 = n13638 ^ n12299 ^ 1'b0 ;
  assign n17385 = n11308 ^ n11217 ^ 1'b0 ;
  assign n17386 = n13134 ^ n6925 ^ 1'b0 ;
  assign n17387 = ~n17245 & n17386 ;
  assign n17388 = n10524 & ~n12705 ;
  assign n17389 = n1283 & ~n2653 ;
  assign n17390 = n17389 ^ n5580 ^ 1'b0 ;
  assign n17391 = n2634 ^ n2389 ^ n547 ;
  assign n17392 = n14264 | n17391 ;
  assign n17393 = n3334 & ~n17392 ;
  assign n17394 = ~n13743 & n17393 ;
  assign n17395 = n1050 | n3935 ;
  assign n17397 = n437 & ~n8393 ;
  assign n17398 = n17397 ^ n13308 ^ 1'b0 ;
  assign n17396 = n4083 & n16986 ;
  assign n17399 = n17398 ^ n17396 ^ 1'b0 ;
  assign n17400 = ~n8241 & n13023 ;
  assign n17401 = ( ~n505 & n4382 ) | ( ~n505 & n5719 ) | ( n4382 & n5719 ) ;
  assign n17402 = n17401 ^ n13371 ^ n6455 ;
  assign n17407 = n10743 | n17108 ;
  assign n17408 = n17407 ^ n36 ^ 1'b0 ;
  assign n17403 = n5648 ^ n4691 ^ n4279 ;
  assign n17404 = n17403 ^ n4886 ^ n2132 ;
  assign n17405 = n16861 ^ n12849 ^ 1'b0 ;
  assign n17406 = ~n17404 & n17405 ;
  assign n17409 = n17408 ^ n17406 ^ 1'b0 ;
  assign n17410 = ~n959 & n7997 ;
  assign n17411 = n11479 & ~n14006 ;
  assign n17412 = n5727 & ~n9014 ;
  assign n17413 = n1321 & ~n12769 ;
  assign n17414 = n17413 ^ n13980 ^ 1'b0 ;
  assign n17415 = n13379 | n17414 ;
  assign n17416 = n344 & n1983 ;
  assign n17417 = n9651 ^ n3266 ^ n2796 ;
  assign n17418 = n9570 | n17417 ;
  assign n17419 = ~n1962 & n4401 ;
  assign n17420 = n15472 & n17419 ;
  assign n17421 = n5158 | n8347 ;
  assign n17428 = n4173 ^ n1568 ^ 1'b0 ;
  assign n17426 = n13251 ^ n3190 ^ n2618 ;
  assign n17425 = n5645 | n15929 ;
  assign n17427 = n17426 ^ n17425 ^ 1'b0 ;
  assign n17422 = n1933 ^ n459 ^ 1'b0 ;
  assign n17423 = n3611 ^ n1471 ^ 1'b0 ;
  assign n17424 = n17422 & ~n17423 ;
  assign n17429 = n17428 ^ n17427 ^ n17424 ;
  assign n17430 = n8225 ^ n1344 ^ 1'b0 ;
  assign n17431 = n11371 & ~n17430 ;
  assign n17432 = n1276 | n12750 ;
  assign n17433 = n2555 ^ n27 ^ 1'b0 ;
  assign n17434 = ~n2386 & n3700 ;
  assign n17435 = n423 | n17434 ;
  assign n17436 = n5667 & ~n17435 ;
  assign n17437 = n17436 ^ n11098 ^ 1'b0 ;
  assign n17438 = n5791 | n6968 ;
  assign n17439 = n17438 ^ n2087 ^ 1'b0 ;
  assign n17440 = n8350 & n17439 ;
  assign n17441 = n17440 ^ n15144 ^ 1'b0 ;
  assign n17442 = ~n1566 & n2632 ;
  assign n17443 = ~n2632 & n17442 ;
  assign n17444 = n522 | n899 ;
  assign n17445 = n522 & ~n17444 ;
  assign n17446 = n5658 & n6756 ;
  assign n17447 = n17445 & n17446 ;
  assign n17448 = ~n17443 & n17447 ;
  assign n17449 = n11274 ^ n1060 ^ 1'b0 ;
  assign n17450 = n17449 ^ n8390 ^ 1'b0 ;
  assign n17451 = n17450 ^ n17052 ^ n1432 ;
  assign n17452 = ~n15596 & n17451 ;
  assign n17453 = n17 & n17452 ;
  assign n17454 = n5870 | n5997 ;
  assign n17455 = n17454 ^ n17061 ^ 1'b0 ;
  assign n17456 = n10870 ^ n1922 ^ 1'b0 ;
  assign n17457 = n16913 | n17456 ;
  assign n17458 = n557 & ~n6219 ;
  assign n17459 = n17458 ^ n5047 ^ 1'b0 ;
  assign n17460 = n327 & n17459 ;
  assign n17461 = n6678 & n17460 ;
  assign n17462 = n11552 | n14748 ;
  assign n17463 = n17462 ^ n16371 ^ 1'b0 ;
  assign n17466 = n3669 & ~n5803 ;
  assign n17467 = ~n10562 & n17466 ;
  assign n17464 = n1712 & ~n6082 ;
  assign n17465 = n1454 & n17464 ;
  assign n17468 = n17467 ^ n17465 ^ 1'b0 ;
  assign n17469 = n1450 & n2764 ;
  assign n17470 = n17469 ^ n6067 ^ 1'b0 ;
  assign n17471 = n17470 ^ n13337 ^ n8643 ;
  assign n17472 = ( n978 & n6277 ) | ( n978 & n17471 ) | ( n6277 & n17471 ) ;
  assign n17473 = n4070 & n7391 ;
  assign n17474 = ~n17472 & n17473 ;
  assign n17475 = n400 & n12338 ;
  assign n17476 = ~n12134 & n17475 ;
  assign n17477 = ~n5008 & n6876 ;
  assign n17479 = n5395 & n5662 ;
  assign n17478 = n2829 & n4986 ;
  assign n17480 = n17479 ^ n17478 ^ 1'b0 ;
  assign n17481 = n10610 & ~n17480 ;
  assign n17482 = ( ~n154 & n982 ) | ( ~n154 & n4135 ) | ( n982 & n4135 ) ;
  assign n17483 = ~n8124 & n17482 ;
  assign n17484 = n17483 ^ n9218 ^ 1'b0 ;
  assign n17485 = n17481 & ~n17484 ;
  assign n17486 = n17477 & n17485 ;
  assign n17487 = n14823 | n17066 ;
  assign n17488 = n2906 | n7034 ;
  assign n17489 = n6442 | n17488 ;
  assign n17490 = n4173 | n17489 ;
  assign n17491 = ~n280 & n1882 ;
  assign n17492 = n12240 ^ n5078 ^ 1'b0 ;
  assign n17493 = n10527 & ~n17492 ;
  assign n17494 = ( ~n6206 & n17491 ) | ( ~n6206 & n17493 ) | ( n17491 & n17493 ) ;
  assign n17495 = n989 ^ n86 ^ 1'b0 ;
  assign n17496 = n17494 & n17495 ;
  assign n17497 = n2213 & n17496 ;
  assign n17498 = n2118 & n8577 ;
  assign n17499 = n3760 & n17498 ;
  assign n17500 = n17499 ^ n1774 ^ 1'b0 ;
  assign n17501 = n1453 & ~n3964 ;
  assign n17502 = ~n3881 & n17501 ;
  assign n17503 = n15467 & ~n17502 ;
  assign n17504 = n13115 ^ n753 ^ 1'b0 ;
  assign n17505 = ~n17072 & n17504 ;
  assign n17506 = ~n15008 & n17505 ;
  assign n17508 = n2549 & ~n2987 ;
  assign n17507 = ( n2397 & ~n2543 ) | ( n2397 & n10915 ) | ( ~n2543 & n10915 ) ;
  assign n17509 = n17508 ^ n17507 ^ n2476 ;
  assign n17510 = ~n5967 & n9151 ;
  assign n17511 = n4977 & n12705 ;
  assign n17512 = n4002 & n12520 ;
  assign n17513 = n17512 ^ n13136 ^ 1'b0 ;
  assign n17514 = n1546 & ~n8224 ;
  assign n17515 = n8448 ^ n6594 ^ n4553 ;
  assign n17516 = ( n5223 & n11553 ) | ( n5223 & ~n17515 ) | ( n11553 & ~n17515 ) ;
  assign n17517 = n3030 & ~n10284 ;
  assign n17518 = n12576 & n17517 ;
  assign n17521 = ~n152 & n388 ;
  assign n17522 = n152 & n17521 ;
  assign n17523 = n418 & ~n1174 ;
  assign n17524 = n17522 & n17523 ;
  assign n17525 = n17524 ^ n2571 ^ 1'b0 ;
  assign n17519 = n3896 & ~n13032 ;
  assign n17520 = n13032 & n17519 ;
  assign n17526 = n17525 ^ n17520 ^ n1592 ;
  assign n17527 = n8110 ^ n5898 ^ 1'b0 ;
  assign n17528 = n17527 ^ n2570 ^ 1'b0 ;
  assign n17529 = n17528 ^ n11727 ^ n9222 ;
  assign n17530 = n17529 ^ n15939 ^ 1'b0 ;
  assign n17531 = n4287 | n17530 ;
  assign n17532 = ~n8908 & n11423 ;
  assign n17533 = n6878 | n17532 ;
  assign n17534 = n2628 & ~n4688 ;
  assign n17535 = ~n17533 & n17534 ;
  assign n17536 = n3218 & ~n9319 ;
  assign n17537 = n17536 ^ n1196 ^ 1'b0 ;
  assign n17540 = n2050 & ~n4858 ;
  assign n17538 = ~n2212 & n3058 ;
  assign n17539 = ~n7005 & n17538 ;
  assign n17541 = n17540 ^ n17539 ^ 1'b0 ;
  assign n17542 = n17537 & n17541 ;
  assign n17543 = n17542 ^ n4799 ^ 1'b0 ;
  assign n17544 = ~n1063 & n14497 ;
  assign n17545 = n6200 ^ n3334 ^ 1'b0 ;
  assign n17546 = n10117 | n17545 ;
  assign n17547 = n13162 ^ n4535 ^ 1'b0 ;
  assign n17548 = ~n7179 & n17547 ;
  assign n17549 = n9779 | n17548 ;
  assign n17550 = n7641 & ~n14458 ;
  assign n17551 = ~n13878 & n17550 ;
  assign n17553 = n6091 | n10638 ;
  assign n17552 = ~n219 & n733 ;
  assign n17554 = n17553 ^ n17552 ^ n924 ;
  assign n17555 = n891 ^ n500 ^ 1'b0 ;
  assign n17556 = n17555 ^ n5823 ^ 1'b0 ;
  assign n17557 = n2583 | n17556 ;
  assign n17558 = n10749 ^ n2081 ^ 1'b0 ;
  assign n17559 = n7421 & ~n7558 ;
  assign n17560 = ( n3863 & n4856 ) | ( n3863 & ~n17559 ) | ( n4856 & ~n17559 ) ;
  assign n17561 = n6927 & n7058 ;
  assign n17562 = n14020 & ~n17561 ;
  assign n17563 = n4183 & n17562 ;
  assign n17564 = n9995 ^ n5331 ^ 1'b0 ;
  assign n17565 = ~n2547 & n4801 ;
  assign n17566 = n17565 ^ n2478 ^ 1'b0 ;
  assign n17567 = n17566 ^ n16760 ^ n4299 ;
  assign n17568 = ~n2136 & n6229 ;
  assign n17569 = n5321 & n17568 ;
  assign n17570 = n15811 ^ n6902 ^ 1'b0 ;
  assign n17571 = n17569 | n17570 ;
  assign n17572 = n1705 & n3896 ;
  assign n17573 = n17572 ^ n5276 ^ 1'b0 ;
  assign n17574 = n10404 ^ n873 ^ 1'b0 ;
  assign n17575 = n7139 | n17574 ;
  assign n17576 = ~n331 & n10403 ;
  assign n17577 = n17575 & n17576 ;
  assign n17578 = n6182 & n14325 ;
  assign n17579 = ( n2515 & ~n4123 ) | ( n2515 & n17578 ) | ( ~n4123 & n17578 ) ;
  assign n17580 = n8438 | n9245 ;
  assign n17581 = n3042 | n5656 ;
  assign n17582 = n16408 | n17581 ;
  assign n17583 = n17582 ^ n15925 ^ n5151 ;
  assign n17585 = n6813 ^ n1073 ^ 1'b0 ;
  assign n17584 = n2956 & n8007 ;
  assign n17586 = n17585 ^ n17584 ^ n8208 ;
  assign n17587 = ~n530 & n16959 ;
  assign n17588 = n14895 ^ n6035 ^ 1'b0 ;
  assign n17589 = n1988 & ~n2175 ;
  assign n17590 = n17589 ^ n2189 ^ 1'b0 ;
  assign n17591 = n9580 & n17590 ;
  assign n17592 = n17591 ^ n10851 ^ 1'b0 ;
  assign n17593 = ( n7599 & ~n17588 ) | ( n7599 & n17592 ) | ( ~n17588 & n17592 ) ;
  assign n17594 = n17593 ^ n1172 ^ 1'b0 ;
  assign n17595 = n5189 | n13274 ;
  assign n17596 = n17594 & ~n17595 ;
  assign n17597 = ~n3287 & n5399 ;
  assign n17598 = n17597 ^ n14672 ^ 1'b0 ;
  assign n17599 = n9403 ^ n2275 ^ 1'b0 ;
  assign n17600 = ~n6775 & n17599 ;
  assign n17601 = n17598 & n17600 ;
  assign n17602 = n16296 ^ n3584 ^ 1'b0 ;
  assign n17603 = ~n5743 & n17602 ;
  assign n17604 = n17603 ^ n8915 ^ 1'b0 ;
  assign n17610 = n4235 & n6880 ;
  assign n17609 = n878 | n8655 ;
  assign n17611 = n17610 ^ n17609 ^ 1'b0 ;
  assign n17605 = n6446 ^ n3738 ^ 1'b0 ;
  assign n17606 = ~n183 & n17605 ;
  assign n17607 = n17606 ^ n10295 ^ 1'b0 ;
  assign n17608 = n13708 | n17607 ;
  assign n17612 = n17611 ^ n17608 ^ 1'b0 ;
  assign n17613 = n10897 ^ n10579 ^ 1'b0 ;
  assign n17614 = ~n2031 & n17613 ;
  assign n17615 = n17614 ^ n966 ^ 1'b0 ;
  assign n17616 = ~n10406 & n14027 ;
  assign n17617 = n2588 & ~n14369 ;
  assign n17618 = n17617 ^ n12231 ^ 1'b0 ;
  assign n17619 = n7364 | n10550 ;
  assign n17620 = n10598 | n17619 ;
  assign n17621 = n17620 ^ n11870 ^ n513 ;
  assign n17622 = n2262 | n17621 ;
  assign n17623 = n2473 & ~n10063 ;
  assign n17624 = n17623 ^ n6498 ^ 1'b0 ;
  assign n17625 = n2614 & n10101 ;
  assign n17626 = ~n6950 & n17625 ;
  assign n17627 = n3367 | n16891 ;
  assign n17628 = n2007 & n3226 ;
  assign n17629 = n17628 ^ n2986 ^ 1'b0 ;
  assign n17630 = ( n340 & n7082 ) | ( n340 & ~n12049 ) | ( n7082 & ~n12049 ) ;
  assign n17631 = n17630 ^ n13555 ^ n3618 ;
  assign n17632 = ( n5562 & n11000 ) | ( n5562 & ~n17631 ) | ( n11000 & ~n17631 ) ;
  assign n17633 = n17629 & ~n17632 ;
  assign n17634 = ~n17627 & n17633 ;
  assign n17635 = n15691 ^ n12665 ^ 1'b0 ;
  assign n17636 = ~n2343 & n7359 ;
  assign n17637 = n17636 ^ n13451 ^ 1'b0 ;
  assign n17638 = n4484 & n13386 ;
  assign n17639 = n16409 ^ n8747 ^ 1'b0 ;
  assign n17640 = n5869 ^ n1038 ^ 1'b0 ;
  assign n17641 = n6302 | n9523 ;
  assign n17642 = n8967 & ~n17641 ;
  assign n17643 = ~n3763 & n6074 ;
  assign n17644 = n3017 | n16403 ;
  assign n17645 = n5860 | n16801 ;
  assign n17646 = n17644 & ~n17645 ;
  assign n17647 = n17646 ^ n2131 ^ 1'b0 ;
  assign n17648 = n6201 & ~n13751 ;
  assign n17649 = ( n1221 & ~n2732 ) | ( n1221 & n16204 ) | ( ~n2732 & n16204 ) ;
  assign n17650 = n14483 ^ n8407 ^ 1'b0 ;
  assign n17651 = ~n7030 & n17650 ;
  assign n17652 = ~n17649 & n17651 ;
  assign n17653 = n6275 ^ n3379 ^ 1'b0 ;
  assign n17654 = n783 | n9388 ;
  assign n17655 = n17653 & ~n17654 ;
  assign n17656 = n753 | n10908 ;
  assign n17657 = n582 & ~n3305 ;
  assign n17658 = ( n4916 & ~n9883 ) | ( n4916 & n11632 ) | ( ~n9883 & n11632 ) ;
  assign n17659 = ~n9746 & n14922 ;
  assign n17660 = n12979 | n17659 ;
  assign n17661 = n9553 | n17660 ;
  assign n17662 = n6870 | n12821 ;
  assign n17663 = n17662 ^ n15271 ^ 1'b0 ;
  assign n17664 = n15681 & n17663 ;
  assign n17665 = n3616 ^ n220 ^ 1'b0 ;
  assign n17666 = n7899 & n15246 ;
  assign n17667 = n4816 ^ n4398 ^ 1'b0 ;
  assign n17668 = ~n4655 & n17667 ;
  assign n17669 = ~n6687 & n17668 ;
  assign n17670 = n14937 ^ n7899 ^ 1'b0 ;
  assign n17671 = ~n4159 & n4590 ;
  assign n17672 = n4578 ^ n419 ^ 1'b0 ;
  assign n17673 = n17671 & ~n17672 ;
  assign n17675 = n10964 & n14728 ;
  assign n17674 = ~n5242 & n5675 ;
  assign n17676 = n17675 ^ n17674 ^ 1'b0 ;
  assign n17677 = n8960 | n17676 ;
  assign n17678 = ( n4932 & n13066 ) | ( n4932 & n17677 ) | ( n13066 & n17677 ) ;
  assign n17679 = n3964 & ~n13541 ;
  assign n17680 = n5189 ^ n3535 ^ 1'b0 ;
  assign n17681 = n9594 & n10005 ;
  assign n17682 = n4995 | n7949 ;
  assign n17683 = n3958 | n17682 ;
  assign n17684 = n768 & n7491 ;
  assign n17685 = n6210 ^ n110 ^ 1'b0 ;
  assign n17686 = n8285 & n11255 ;
  assign n17687 = n17686 ^ n6542 ^ n1140 ;
  assign n17688 = n17685 & ~n17687 ;
  assign n17689 = ~n1260 & n6393 ;
  assign n17690 = n6099 & ~n17689 ;
  assign n17691 = n2719 & n17690 ;
  assign n17692 = n2154 ^ n1983 ^ 1'b0 ;
  assign n17693 = n16442 & ~n17692 ;
  assign n17694 = ~n5937 & n7076 ;
  assign n17695 = ( n2421 & n2796 ) | ( n2421 & n9928 ) | ( n2796 & n9928 ) ;
  assign n17696 = n3946 ^ n1771 ^ 1'b0 ;
  assign n17697 = n10126 ^ n6267 ^ 1'b0 ;
  assign n17698 = ( n7975 & ~n14773 ) | ( n7975 & n17697 ) | ( ~n14773 & n17697 ) ;
  assign n17699 = ~n468 & n3166 ;
  assign n17700 = ~n8552 & n17699 ;
  assign n17701 = n17700 ^ n4570 ^ 1'b0 ;
  assign n17702 = n17701 ^ n7601 ^ 1'b0 ;
  assign n17703 = n8702 ^ n4250 ^ 1'b0 ;
  assign n17704 = n1132 & n17703 ;
  assign n17705 = n17704 ^ n14362 ^ 1'b0 ;
  assign n17706 = n17608 & ~n17705 ;
  assign n17707 = ~n401 & n7099 ;
  assign n17708 = n17707 ^ n4381 ^ 1'b0 ;
  assign n17709 = ~n16263 & n17708 ;
  assign n17710 = n995 | n6082 ;
  assign n17711 = n17710 ^ n11737 ^ 1'b0 ;
  assign n17712 = n9694 & ~n17711 ;
  assign n17713 = n4886 | n17712 ;
  assign n17714 = n2163 & ~n17713 ;
  assign n17715 = n17714 ^ n3488 ^ 1'b0 ;
  assign n17719 = n6722 ^ n6036 ^ 1'b0 ;
  assign n17720 = ~n4141 & n17719 ;
  assign n17718 = n6080 & n7955 ;
  assign n17716 = n1845 & ~n10606 ;
  assign n17717 = n3618 & n17716 ;
  assign n17721 = n17720 ^ n17718 ^ n17717 ;
  assign n17722 = n12231 ^ n3317 ^ 1'b0 ;
  assign n17723 = n2940 & ~n17722 ;
  assign n17724 = n11699 & n17723 ;
  assign n17725 = n1603 & n17724 ;
  assign n17726 = n4770 & ~n17725 ;
  assign n17727 = n17726 ^ n6431 ^ 1'b0 ;
  assign n17728 = n3992 & ~n17403 ;
  assign n17729 = n17728 ^ n16319 ^ 1'b0 ;
  assign n17730 = ~n9592 & n9959 ;
  assign n17731 = n17730 ^ n14493 ^ 1'b0 ;
  assign n17732 = n7008 | n15538 ;
  assign n17733 = n1938 & n15569 ;
  assign n17734 = n2376 & n17733 ;
  assign n17735 = n17732 & n17734 ;
  assign n17736 = n13355 ^ n7421 ^ 1'b0 ;
  assign n17737 = n366 | n17736 ;
  assign n17738 = n17737 ^ n8236 ^ 1'b0 ;
  assign n17739 = n17735 & ~n17738 ;
  assign n17742 = n2090 ^ n2074 ^ n148 ;
  assign n17740 = ~n366 & n972 ;
  assign n17741 = n6367 & n17740 ;
  assign n17743 = n17742 ^ n17741 ^ n16633 ;
  assign n17744 = n4659 ^ n894 ^ 1'b0 ;
  assign n17745 = n615 & ~n7931 ;
  assign n17746 = n17744 & ~n17745 ;
  assign n17747 = n6585 ^ n334 ^ n312 ;
  assign n17748 = ~n6697 & n8795 ;
  assign n17749 = n15878 & n17748 ;
  assign n17750 = n17749 ^ n15017 ^ 1'b0 ;
  assign n17751 = n189 | n17750 ;
  assign n17758 = n724 | n3958 ;
  assign n17759 = n1251 | n17758 ;
  assign n17752 = n17310 ^ n996 ^ 1'b0 ;
  assign n17753 = n10321 | n17752 ;
  assign n17754 = n12915 ^ n5939 ^ 1'b0 ;
  assign n17755 = n8532 & n17754 ;
  assign n17756 = n17753 & n17755 ;
  assign n17757 = n2106 & ~n17756 ;
  assign n17760 = n17759 ^ n17757 ^ 1'b0 ;
  assign n17761 = n5524 & n9010 ;
  assign n17762 = n17761 ^ n8011 ^ 1'b0 ;
  assign n17763 = n17762 ^ n717 ^ 1'b0 ;
  assign n17765 = n2248 & n8233 ;
  assign n17766 = n17765 ^ n4744 ^ 1'b0 ;
  assign n17764 = n956 | n1987 ;
  assign n17767 = n17766 ^ n17764 ^ 1'b0 ;
  assign n17768 = n3601 & n9417 ;
  assign n17769 = n13832 & n17768 ;
  assign n17770 = n17118 ^ n11523 ^ n4720 ;
  assign n17771 = n2565 & n2833 ;
  assign n17772 = ~n6844 & n10720 ;
  assign n17773 = ~n17771 & n17772 ;
  assign n17774 = n5524 & n7785 ;
  assign n17775 = n6004 | n6749 ;
  assign n17776 = ~n2415 & n5185 ;
  assign n17777 = n8674 & n17776 ;
  assign n17778 = ~n7549 & n8834 ;
  assign n17779 = n17777 & ~n17778 ;
  assign n17780 = n15019 & ~n16613 ;
  assign n17781 = n17780 ^ n13018 ^ 1'b0 ;
  assign n17782 = n17781 ^ n453 ^ 1'b0 ;
  assign n17783 = n345 & ~n17782 ;
  assign n17784 = n482 & ~n13238 ;
  assign n17785 = n11232 & n17784 ;
  assign n17786 = n12380 ^ n8702 ^ 1'b0 ;
  assign n17787 = ~n1928 & n17786 ;
  assign n17788 = n1434 ^ n497 ^ 1'b0 ;
  assign n17789 = n3891 & ~n17788 ;
  assign n17790 = n14039 ^ n5954 ^ 1'b0 ;
  assign n17793 = n1730 & n2438 ;
  assign n17794 = n17793 ^ n3015 ^ 1'b0 ;
  assign n17791 = n2656 & ~n6620 ;
  assign n17792 = n8154 & n17791 ;
  assign n17795 = n17794 ^ n17792 ^ n10146 ;
  assign n17796 = n14749 | n17795 ;
  assign n17797 = n17790 & ~n17796 ;
  assign n17798 = ~n2754 & n2772 ;
  assign n17799 = n1984 | n7765 ;
  assign n17800 = ( n4368 & n4698 ) | ( n4368 & n17799 ) | ( n4698 & n17799 ) ;
  assign n17802 = ~n9616 & n11554 ;
  assign n17801 = n445 | n459 ;
  assign n17803 = n17802 ^ n17801 ^ 1'b0 ;
  assign n17804 = ~n12393 & n17803 ;
  assign n17805 = n6885 ^ n4457 ^ 1'b0 ;
  assign n17806 = n3990 | n12225 ;
  assign n17807 = n1163 & ~n10852 ;
  assign n17808 = n9210 & ~n13390 ;
  assign n17809 = n17808 ^ n188 ^ 1'b0 ;
  assign n17814 = n3339 ^ n2121 ^ 1'b0 ;
  assign n17815 = n9193 & n17814 ;
  assign n17810 = n9923 ^ n3800 ^ 1'b0 ;
  assign n17811 = ~n3514 & n12549 ;
  assign n17812 = n17811 ^ n6972 ^ 1'b0 ;
  assign n17813 = n17810 | n17812 ;
  assign n17816 = n17815 ^ n17813 ^ 1'b0 ;
  assign n17817 = n974 & n2404 ;
  assign n17818 = n17817 ^ n225 ^ 1'b0 ;
  assign n17819 = n515 | n17818 ;
  assign n17820 = n6353 | n17819 ;
  assign n17821 = n695 & ~n7630 ;
  assign n17822 = n1182 & ~n1381 ;
  assign n17823 = ~n1811 & n6080 ;
  assign n17824 = n17823 ^ n3437 ^ 1'b0 ;
  assign n17825 = n17822 & ~n17824 ;
  assign n17826 = n14694 ^ n12990 ^ 1'b0 ;
  assign n17827 = n15203 | n17826 ;
  assign n17828 = n11005 ^ n5183 ^ 1'b0 ;
  assign n17829 = n8949 ^ n17 ^ 1'b0 ;
  assign n17830 = n16192 ^ n6644 ^ 1'b0 ;
  assign n17831 = ~n5202 & n17830 ;
  assign n17832 = n17829 & n17831 ;
  assign n17833 = n515 & n17832 ;
  assign n17834 = ~n4608 & n17833 ;
  assign n17835 = n3892 & ~n17142 ;
  assign n17836 = ~n318 & n17835 ;
  assign n17837 = n6820 | n17836 ;
  assign n17838 = n16407 | n17837 ;
  assign n17839 = n10766 & ~n17838 ;
  assign n17840 = ~n1192 & n12637 ;
  assign n17841 = ( n6208 & ~n13523 ) | ( n6208 & n17840 ) | ( ~n13523 & n17840 ) ;
  assign n17842 = n919 | n3388 ;
  assign n17843 = n9933 | n17842 ;
  assign n17848 = n14875 ^ n10404 ^ n1582 ;
  assign n17844 = n4427 & ~n7106 ;
  assign n17845 = n17844 ^ n989 ^ 1'b0 ;
  assign n17846 = n17845 ^ n12251 ^ n724 ;
  assign n17847 = n10752 & ~n17846 ;
  assign n17849 = n17848 ^ n17847 ^ 1'b0 ;
  assign n17850 = n17843 & n17849 ;
  assign n17851 = n12757 ^ n69 ^ 1'b0 ;
  assign n17852 = n6527 & ~n17851 ;
  assign n17853 = n17852 ^ n565 ^ 1'b0 ;
  assign n17854 = n10911 ^ n3212 ^ 1'b0 ;
  assign n17855 = n5562 & n17854 ;
  assign n17856 = n17855 ^ n10937 ^ 1'b0 ;
  assign n17857 = n12337 | n17856 ;
  assign n17858 = n12346 | n17857 ;
  assign n17859 = ( n1174 & n3085 ) | ( n1174 & ~n13986 ) | ( n3085 & ~n13986 ) ;
  assign n17860 = n5747 & ~n10298 ;
  assign n17861 = ~n2272 & n5461 ;
  assign n17862 = n17861 ^ n14889 ^ 1'b0 ;
  assign n17863 = n2267 & n8274 ;
  assign n17864 = ~n2755 & n17863 ;
  assign n17865 = n9867 ^ n1812 ^ 1'b0 ;
  assign n17866 = n7877 & n17865 ;
  assign n17867 = n11913 & n17866 ;
  assign n17868 = ~n10592 & n17867 ;
  assign n17869 = ~n1962 & n17734 ;
  assign n17875 = n11046 & ~n11733 ;
  assign n17876 = ~n12766 & n17875 ;
  assign n17870 = ~n2751 & n3199 ;
  assign n17871 = n890 & n17870 ;
  assign n17872 = n9136 ^ n421 ^ 1'b0 ;
  assign n17873 = n4012 & ~n17872 ;
  assign n17874 = n17871 | n17873 ;
  assign n17877 = n17876 ^ n17874 ^ 1'b0 ;
  assign n17878 = n2085 & n17877 ;
  assign n17879 = n17878 ^ n17607 ^ n1369 ;
  assign n17880 = ( n1639 & n2321 ) | ( n1639 & n4523 ) | ( n2321 & n4523 ) ;
  assign n17881 = n17880 ^ n10087 ^ 1'b0 ;
  assign n17882 = n6698 ^ n1050 ^ 1'b0 ;
  assign n17883 = n2137 & ~n3574 ;
  assign n17884 = n13351 & n17883 ;
  assign n17885 = ~n17882 & n17884 ;
  assign n17886 = n17885 ^ n11582 ^ n4944 ;
  assign n17887 = n5524 ^ n3825 ^ 1'b0 ;
  assign n17888 = n12218 | n17887 ;
  assign n17889 = ~n2520 & n5096 ;
  assign n17890 = n10158 & n17889 ;
  assign n17891 = n17890 ^ n477 ^ 1'b0 ;
  assign n17892 = ~n700 & n17753 ;
  assign n17893 = x1 | n6566 ;
  assign n17894 = n15272 ^ n6901 ^ 1'b0 ;
  assign n17895 = n2232 & n17894 ;
  assign n17896 = n17895 ^ n10536 ^ 1'b0 ;
  assign n17897 = n1734 & ~n17896 ;
  assign n17898 = n3418 ^ n1312 ^ 1'b0 ;
  assign n17899 = n11189 & ~n17898 ;
  assign n17900 = ( ~n3676 & n8724 ) | ( ~n3676 & n17899 ) | ( n8724 & n17899 ) ;
  assign n17901 = n17647 & n17900 ;
  assign n17902 = ~n926 & n12050 ;
  assign n17903 = ~n623 & n10237 ;
  assign n17904 = n17903 ^ n15841 ^ 1'b0 ;
  assign n17909 = ( n1278 & ~n17084 ) | ( n1278 & n17829 ) | ( ~n17084 & n17829 ) ;
  assign n17910 = n736 & n17909 ;
  assign n17911 = ~n17909 & n17910 ;
  assign n17905 = n8331 ^ n898 ^ 1'b0 ;
  assign n17906 = n727 & n17905 ;
  assign n17907 = ~n5747 & n17906 ;
  assign n17908 = ~n7187 & n17907 ;
  assign n17912 = n17911 ^ n17908 ^ 1'b0 ;
  assign n17913 = n17912 ^ n6353 ^ 1'b0 ;
  assign n17914 = n1435 & ~n1747 ;
  assign n17915 = ~n13077 & n17914 ;
  assign n17916 = n11406 & ~n17915 ;
  assign n17917 = n17916 ^ n782 ^ 1'b0 ;
  assign n17921 = ~n1688 & n4194 ;
  assign n17918 = n4246 & n7277 ;
  assign n17919 = n17918 ^ n218 ^ 1'b0 ;
  assign n17920 = ~n6762 & n17919 ;
  assign n17922 = n17921 ^ n17920 ^ 1'b0 ;
  assign n17923 = n863 & n7493 ;
  assign n17924 = n17923 ^ n13523 ^ 1'b0 ;
  assign n17925 = n9233 ^ n6423 ^ 1'b0 ;
  assign n17926 = n17924 & ~n17925 ;
  assign n17927 = n4512 ^ n3623 ^ 1'b0 ;
  assign n17928 = n17662 & n17927 ;
  assign n17929 = ~n758 & n17928 ;
  assign n17930 = n2114 & n16770 ;
  assign n17931 = n17930 ^ n588 ^ 1'b0 ;
  assign n17932 = n3129 & n8249 ;
  assign n17933 = n2267 ^ n481 ^ 1'b0 ;
  assign n17934 = ~n11094 & n17933 ;
  assign n17935 = n16485 ^ n6827 ^ 1'b0 ;
  assign n17936 = ~n13566 & n17935 ;
  assign n17937 = n2367 ^ n1083 ^ 1'b0 ;
  assign n17938 = n2637 & ~n3571 ;
  assign n17939 = n1584 | n17938 ;
  assign n17940 = ~n4123 & n11523 ;
  assign n17941 = n6428 ^ n5636 ^ 1'b0 ;
  assign n17942 = ~n12867 & n17941 ;
  assign n17943 = n17942 ^ n12927 ^ 1'b0 ;
  assign n17944 = n8222 | n14635 ;
  assign n17945 = n17944 ^ n17266 ^ 1'b0 ;
  assign n17946 = ( n225 & n607 ) | ( n225 & ~n12450 ) | ( n607 & ~n12450 ) ;
  assign n17947 = n49 & n2462 ;
  assign n17948 = ~n2462 & n17947 ;
  assign n17949 = n17948 ^ n10950 ^ 1'b0 ;
  assign n17950 = n192 & ~n10330 ;
  assign n17951 = n10330 & n17950 ;
  assign n17952 = n765 | n17951 ;
  assign n17953 = n765 & ~n17952 ;
  assign n17954 = ~n2175 & n3871 ;
  assign n17955 = n2175 & n17954 ;
  assign n17956 = n3019 & ~n17955 ;
  assign n17957 = ~n3019 & n17956 ;
  assign n17958 = n17957 ^ n5184 ^ 1'b0 ;
  assign n17959 = n17953 | n17958 ;
  assign n17960 = n17949 & ~n17959 ;
  assign n17961 = ~n17949 & n17960 ;
  assign n17962 = ~n10601 & n15636 ;
  assign n17963 = ~n5150 & n12733 ;
  assign n17964 = ( ~n7871 & n12401 ) | ( ~n7871 & n14828 ) | ( n12401 & n14828 ) ;
  assign n17965 = n17964 ^ n1432 ^ 1'b0 ;
  assign n17966 = ( n4267 & n6949 ) | ( n4267 & ~n15914 ) | ( n6949 & ~n15914 ) ;
  assign n17967 = n17409 ^ n14653 ^ 1'b0 ;
  assign n17968 = n3804 | n17967 ;
  assign n17969 = n3111 | n11934 ;
  assign n17970 = n8091 ^ n4466 ^ 1'b0 ;
  assign n17971 = ~n3312 & n17970 ;
  assign n17972 = n17971 ^ n667 ^ 1'b0 ;
  assign n17973 = n2408 & ~n12345 ;
  assign n17974 = n17973 ^ n1327 ^ 1'b0 ;
  assign n17975 = n1383 & ~n16112 ;
  assign n17976 = n11146 & ~n17272 ;
  assign n17977 = n17976 ^ n12150 ^ 1'b0 ;
  assign n17978 = n17975 | n17977 ;
  assign n17979 = n8002 ^ n2541 ^ 1'b0 ;
  assign n17980 = ~n3545 & n17979 ;
  assign n17981 = n3766 & n17915 ;
  assign n17982 = n9676 | n15105 ;
  assign n17983 = n16410 ^ n309 ^ 1'b0 ;
  assign n17984 = n1343 & ~n6015 ;
  assign n17985 = n5765 | n8405 ;
  assign n17986 = n10425 | n17985 ;
  assign n17987 = n2578 & n17449 ;
  assign n17988 = n12513 ^ n1385 ^ 1'b0 ;
  assign n17989 = n8449 & ~n17988 ;
  assign n17990 = n17989 ^ n2031 ^ 1'b0 ;
  assign n17991 = n6342 | n8966 ;
  assign n17992 = n17265 | n17991 ;
  assign n17993 = n4020 ^ n3110 ^ 1'b0 ;
  assign n17994 = ( n1967 & n6675 ) | ( n1967 & ~n17993 ) | ( n6675 & ~n17993 ) ;
  assign n17995 = n3040 | n17994 ;
  assign n17996 = n17995 ^ n14487 ^ 1'b0 ;
  assign n17997 = n1912 & ~n17235 ;
  assign n17998 = ~n331 & n17997 ;
  assign n17999 = n1720 ^ n1591 ^ x3 ;
  assign n18000 = n17999 ^ n9693 ^ 1'b0 ;
  assign n18001 = ~n14720 & n18000 ;
  assign n18002 = n1988 & ~n18001 ;
  assign n18003 = ~n4618 & n13626 ;
  assign n18004 = n14428 | n18003 ;
  assign n18005 = n15596 ^ n7350 ^ n6846 ;
  assign n18006 = n16137 & ~n18005 ;
  assign n18007 = n6601 & ~n9657 ;
  assign n18008 = n7052 ^ n2407 ^ 1'b0 ;
  assign n18009 = n11875 & ~n18008 ;
  assign n18010 = n18009 ^ n1325 ^ 1'b0 ;
  assign n18011 = ( ~n1912 & n4949 ) | ( ~n1912 & n5058 ) | ( n4949 & n5058 ) ;
  assign n18012 = ~n10087 & n18011 ;
  assign n18013 = n18012 ^ n752 ^ 1'b0 ;
  assign n18014 = n914 & n7112 ;
  assign n18015 = n4105 ^ n3891 ^ n481 ;
  assign n18016 = n18015 ^ n1918 ^ 1'b0 ;
  assign n18017 = ( n857 & n5061 ) | ( n857 & n6538 ) | ( n5061 & n6538 ) ;
  assign n18018 = n12871 ^ n4086 ^ 1'b0 ;
  assign n18019 = n3477 | n11913 ;
  assign n18020 = n3526 ^ n2246 ^ 1'b0 ;
  assign n18021 = n18020 ^ n12865 ^ n3056 ;
  assign n18022 = n9696 ^ n7596 ^ n5459 ;
  assign n18023 = n18022 ^ n11675 ^ 1'b0 ;
  assign n18024 = n1631 & n18023 ;
  assign n18025 = n14968 ^ n8403 ^ 1'b0 ;
  assign n18026 = n1828 & n8883 ;
  assign n18027 = n14989 & n18026 ;
  assign n18031 = ~n2527 & n7234 ;
  assign n18028 = n1726 & n10723 ;
  assign n18029 = n18028 ^ n3635 ^ 1'b0 ;
  assign n18030 = n1469 & ~n18029 ;
  assign n18032 = n18031 ^ n18030 ^ 1'b0 ;
  assign n18033 = n14478 & n18032 ;
  assign n18034 = n15659 ^ n3090 ^ 1'b0 ;
  assign n18035 = n16629 ^ n5897 ^ 1'b0 ;
  assign n18036 = n1707 & n2807 ;
  assign n18037 = n16847 & ~n18036 ;
  assign n18038 = ~n302 & n16518 ;
  assign n18039 = n1741 & n18038 ;
  assign n18040 = n4039 & ~n5626 ;
  assign n18041 = n12755 ^ n4250 ^ 1'b0 ;
  assign n18042 = n18040 & n18041 ;
  assign n18044 = n13397 ^ n667 ^ 1'b0 ;
  assign n18045 = ~n7767 & n18044 ;
  assign n18046 = n18045 ^ n6344 ^ 1'b0 ;
  assign n18047 = n4526 | n18046 ;
  assign n18048 = n18047 ^ n727 ^ 1'b0 ;
  assign n18043 = n2765 & ~n10378 ;
  assign n18049 = n18048 ^ n18043 ^ 1'b0 ;
  assign n18050 = n10752 ^ n7027 ^ 1'b0 ;
  assign n18051 = n6982 & ~n8292 ;
  assign n18052 = n7259 & ~n17863 ;
  assign n18053 = n3107 ^ n283 ^ 1'b0 ;
  assign n18054 = n18053 ^ n11676 ^ 1'b0 ;
  assign n18055 = n506 | n18054 ;
  assign n18056 = n14010 & n14087 ;
  assign n18057 = n18056 ^ n3179 ^ 1'b0 ;
  assign n18058 = n11296 | n18057 ;
  assign n18059 = n18058 ^ n2758 ^ 1'b0 ;
  assign n18066 = ( n1975 & n5285 ) | ( n1975 & ~n6096 ) | ( n5285 & ~n6096 ) ;
  assign n18067 = ( ~n4365 & n6275 ) | ( ~n4365 & n18066 ) | ( n6275 & n18066 ) ;
  assign n18068 = n6217 ^ n4376 ^ 1'b0 ;
  assign n18069 = ~n18067 & n18068 ;
  assign n18060 = n505 & n5045 ;
  assign n18061 = n4088 & ~n9829 ;
  assign n18062 = n18061 ^ n8885 ^ 1'b0 ;
  assign n18063 = n11979 & ~n18062 ;
  assign n18064 = n18063 ^ n5916 ^ 1'b0 ;
  assign n18065 = n18060 & ~n18064 ;
  assign n18070 = n18069 ^ n18065 ^ 1'b0 ;
  assign n18071 = n10178 ^ n74 ^ 1'b0 ;
  assign n18072 = ~n4276 & n18071 ;
  assign n18073 = n18072 ^ n2958 ^ 1'b0 ;
  assign n18074 = n3944 & n7823 ;
  assign n18075 = n18074 ^ n2778 ^ 1'b0 ;
  assign n18076 = ~n18073 & n18075 ;
  assign n18077 = n13050 ^ n6081 ^ 1'b0 ;
  assign n18078 = n14003 ^ n241 ^ 1'b0 ;
  assign n18079 = ~n805 & n5906 ;
  assign n18080 = n18079 ^ n1392 ^ 1'b0 ;
  assign n18081 = ( ~n11371 & n11717 ) | ( ~n11371 & n18080 ) | ( n11717 & n18080 ) ;
  assign n18082 = n17365 & n18081 ;
  assign n18083 = n18078 & n18082 ;
  assign n18084 = ~n18077 & n18083 ;
  assign n18085 = n10751 ^ n3805 ^ 1'b0 ;
  assign n18086 = n14208 & ~n18085 ;
  assign n18087 = n18086 ^ n14031 ^ 1'b0 ;
  assign n18088 = n611 & ~n16697 ;
  assign n18089 = n18088 ^ n7810 ^ 1'b0 ;
  assign n18090 = n16303 ^ n6781 ^ 1'b0 ;
  assign n18091 = ~n2394 & n18090 ;
  assign n18092 = n14275 | n15561 ;
  assign n18093 = n2010 ^ n1897 ^ 1'b0 ;
  assign n18094 = n15695 ^ n2136 ^ 1'b0 ;
  assign n18095 = ~n9291 & n18094 ;
  assign n18096 = n18093 & ~n18095 ;
  assign n18097 = ~n8957 & n18096 ;
  assign n18098 = n18097 ^ n5201 ^ 1'b0 ;
  assign n18099 = n12636 | n18098 ;
  assign n18100 = n11657 ^ n4532 ^ 1'b0 ;
  assign n18101 = n4271 & n9373 ;
  assign n18102 = n18101 ^ n8926 ^ n8211 ;
  assign n18103 = n18102 ^ n12667 ^ 1'b0 ;
  assign n18104 = n16274 & ~n18103 ;
  assign n18105 = n15273 ^ n9715 ^ 1'b0 ;
  assign n18106 = n269 | n18105 ;
  assign n18107 = n18106 ^ n5606 ^ 1'b0 ;
  assign n18108 = n8061 & n18107 ;
  assign n18109 = ~n1845 & n6748 ;
  assign n18110 = n17420 & n18109 ;
  assign n18111 = n2203 | n16667 ;
  assign n18112 = ~n11742 & n16527 ;
  assign n18113 = n14264 & n18112 ;
  assign n18114 = n11447 & ~n18113 ;
  assign n18115 = ( n10156 & ~n18111 ) | ( n10156 & n18114 ) | ( ~n18111 & n18114 ) ;
  assign n18116 = n9693 ^ n4313 ^ 1'b0 ;
  assign n18117 = n13532 & n18116 ;
  assign n18123 = n1615 ^ n167 ^ 1'b0 ;
  assign n18124 = n5365 & n18123 ;
  assign n18120 = n8117 & n16066 ;
  assign n18121 = ~n5109 & n18120 ;
  assign n18122 = n758 & ~n18121 ;
  assign n18118 = n4944 ^ n3489 ^ 1'b0 ;
  assign n18119 = n14497 & n18118 ;
  assign n18125 = n18124 ^ n18122 ^ n18119 ;
  assign n18126 = n3064 & n9274 ;
  assign n18127 = ( ~n4053 & n6320 ) | ( ~n4053 & n12303 ) | ( n6320 & n12303 ) ;
  assign n18128 = n8915 ^ n8111 ^ n183 ;
  assign n18129 = n484 & ~n18128 ;
  assign n18130 = n18129 ^ n8174 ^ 1'b0 ;
  assign n18131 = n18127 & ~n18130 ;
  assign n18132 = n18131 ^ n13538 ^ 1'b0 ;
  assign n18133 = n567 & ~n8161 ;
  assign n18134 = n18133 ^ n6539 ^ 1'b0 ;
  assign n18135 = n3928 ^ n2433 ^ 1'b0 ;
  assign n18136 = n17656 | n18135 ;
  assign n18137 = n2381 & n2824 ;
  assign n18138 = n18137 ^ n441 ^ 1'b0 ;
  assign n18139 = n16006 ^ n3094 ^ 1'b0 ;
  assign n18140 = n15385 & n18139 ;
  assign n18142 = n3937 | n8690 ;
  assign n18141 = n1476 & ~n1812 ;
  assign n18143 = n18142 ^ n18141 ^ 1'b0 ;
  assign n18144 = n714 | n18143 ;
  assign n18145 = n9779 ^ n3647 ^ 1'b0 ;
  assign n18146 = ~n2387 & n18145 ;
  assign n18147 = n5406 | n14316 ;
  assign n18148 = n2719 | n9835 ;
  assign n18149 = n2940 & ~n18148 ;
  assign n18150 = n3374 & ~n9045 ;
  assign n18151 = n18150 ^ n7335 ^ 1'b0 ;
  assign n18152 = ~n2095 & n18151 ;
  assign n18153 = ~n6893 & n7590 ;
  assign n18154 = ~n4222 & n18153 ;
  assign n18155 = ~n7067 & n11520 ;
  assign n18156 = n15095 & n18155 ;
  assign n18157 = n18156 ^ n13534 ^ 1'b0 ;
  assign n18158 = ~n18154 & n18157 ;
  assign n18160 = n4269 | n4924 ;
  assign n18161 = n18160 ^ n1381 ^ 1'b0 ;
  assign n18159 = n9540 & n10086 ;
  assign n18162 = n18161 ^ n18159 ^ 1'b0 ;
  assign n18163 = n17635 ^ n13146 ^ 1'b0 ;
  assign n18164 = ~n11893 & n18163 ;
  assign n18165 = n1075 | n7558 ;
  assign n18166 = n14670 | n18165 ;
  assign n18167 = n13861 ^ n2176 ^ n1374 ;
  assign n18168 = n1732 & ~n18167 ;
  assign n18169 = n18168 ^ n8891 ^ 1'b0 ;
  assign n18170 = n4241 & n17373 ;
  assign n18171 = ~n15612 & n18170 ;
  assign n18172 = n4201 | n6997 ;
  assign n18173 = n18172 ^ n12832 ^ 1'b0 ;
  assign n18174 = n3505 ^ n1868 ^ 1'b0 ;
  assign n18175 = n2634 & ~n18174 ;
  assign n18176 = ~n265 & n18175 ;
  assign n18177 = n18176 ^ n7735 ^ 1'b0 ;
  assign n18178 = ~n10890 & n18177 ;
  assign n18179 = n1862 ^ n1548 ^ 1'b0 ;
  assign n18180 = ~n7643 & n18179 ;
  assign n18181 = n18180 ^ n6193 ^ 1'b0 ;
  assign n18182 = ~n8752 & n11360 ;
  assign n18183 = ~n5161 & n18182 ;
  assign n18184 = n712 & n13774 ;
  assign n18185 = n10476 | n18184 ;
  assign n18186 = ~n8480 & n14428 ;
  assign n18189 = n14669 ^ n12397 ^ 1'b0 ;
  assign n18190 = n3998 & n18189 ;
  assign n18191 = n18190 ^ n11857 ^ n805 ;
  assign n18187 = n7471 & ~n9605 ;
  assign n18188 = n211 | n18187 ;
  assign n18192 = n18191 ^ n18188 ^ 1'b0 ;
  assign n18193 = n619 & n10029 ;
  assign n18194 = n16595 & n18193 ;
  assign n18195 = ~n9987 & n14868 ;
  assign n18196 = n8944 & ~n10667 ;
  assign n18197 = ~n18195 & n18196 ;
  assign n18199 = ( ~n6067 & n9421 ) | ( ~n6067 & n12756 ) | ( n9421 & n12756 ) ;
  assign n18198 = n1306 | n12035 ;
  assign n18200 = n18199 ^ n18198 ^ n8029 ;
  assign n18201 = ~n1223 & n6371 ;
  assign n18202 = n18201 ^ n4624 ^ 1'b0 ;
  assign n18203 = n4700 & ~n8639 ;
  assign n18204 = n17806 & n18203 ;
  assign n18205 = n18202 & n18204 ;
  assign n18206 = n17008 ^ n4995 ^ 1'b0 ;
  assign n18207 = n11476 | n18206 ;
  assign n18208 = n4250 & ~n11119 ;
  assign n18209 = ( n246 & ~n1345 ) | ( n246 & n4627 ) | ( ~n1345 & n4627 ) ;
  assign n18210 = n17259 | n18209 ;
  assign n18211 = n152 & ~n12891 ;
  assign n18212 = n10352 ^ n8233 ^ 1'b0 ;
  assign n18213 = n18211 & n18212 ;
  assign n18214 = n9187 & n12724 ;
  assign n18215 = ~n2145 & n18214 ;
  assign n18216 = n5249 & ~n5660 ;
  assign n18217 = n18215 & n18216 ;
  assign n18218 = n9158 ^ n5885 ^ 1'b0 ;
  assign n18219 = n18218 ^ n8883 ^ 1'b0 ;
  assign n18220 = n18217 | n18219 ;
  assign n18222 = n817 & n1658 ;
  assign n18223 = n18222 ^ n13018 ^ 1'b0 ;
  assign n18224 = n6454 ^ n5481 ^ 1'b0 ;
  assign n18225 = ~n18223 & n18224 ;
  assign n18221 = n7319 & ~n8785 ;
  assign n18226 = n18225 ^ n18221 ^ 1'b0 ;
  assign n18227 = ~n3227 & n7053 ;
  assign n18228 = n4434 ^ n194 ^ 1'b0 ;
  assign n18229 = ~n5244 & n18228 ;
  assign n18230 = n1962 | n6593 ;
  assign n18231 = n18230 ^ n4420 ^ 1'b0 ;
  assign n18232 = n3198 & ~n9720 ;
  assign n18233 = n8823 ^ n1014 ^ 1'b0 ;
  assign n18234 = n18232 & n18233 ;
  assign n18235 = ~n18231 & n18234 ;
  assign n18236 = ~n16073 & n18235 ;
  assign n18237 = n8157 & n9721 ;
  assign n18238 = n18237 ^ n6701 ^ 1'b0 ;
  assign n18239 = n12793 & n18238 ;
  assign n18240 = n18239 ^ n1244 ^ 1'b0 ;
  assign n18241 = ~n956 & n3226 ;
  assign n18242 = ~n7147 & n18241 ;
  assign n18243 = n4038 & ~n7153 ;
  assign n18244 = n18243 ^ n16709 ^ 1'b0 ;
  assign n18245 = n10792 & ~n18244 ;
  assign n18246 = n10003 ^ n493 ^ 1'b0 ;
  assign n18247 = n1291 | n3827 ;
  assign n18248 = n12379 & ~n18247 ;
  assign n18249 = n12752 ^ n3556 ^ n2682 ;
  assign n18250 = ~n2614 & n17709 ;
  assign n18251 = n2671 & n7897 ;
  assign n18252 = ~n11699 & n18251 ;
  assign n18255 = n3510 ^ n2541 ^ 1'b0 ;
  assign n18253 = n9390 | n9854 ;
  assign n18254 = n1506 & ~n18253 ;
  assign n18256 = n18255 ^ n18254 ^ 1'b0 ;
  assign n18257 = ~n2304 & n16463 ;
  assign n18258 = n1161 & n18257 ;
  assign n18259 = ~n4143 & n4483 ;
  assign n18260 = n18259 ^ n9621 ^ 1'b0 ;
  assign n18261 = n13163 & n18260 ;
  assign n18262 = n1582 | n6904 ;
  assign n18263 = n3339 | n18262 ;
  assign n18264 = ~n17938 & n18263 ;
  assign n18265 = ~n11377 & n11451 ;
  assign n18266 = n2802 & n18265 ;
  assign n18267 = n13848 & ~n18266 ;
  assign n18268 = n18267 ^ n10118 ^ 1'b0 ;
  assign n18269 = n2193 & n5123 ;
  assign n18270 = n18269 ^ n3643 ^ 1'b0 ;
  assign n18271 = n11691 | n11898 ;
  assign n18272 = n13632 ^ n8273 ^ 1'b0 ;
  assign n18273 = n5463 ^ n4028 ^ 1'b0 ;
  assign n18274 = n18273 ^ n3867 ^ 1'b0 ;
  assign n18275 = n4554 | n17087 ;
  assign n18276 = n18275 ^ n6903 ^ 1'b0 ;
  assign n18279 = n14932 ^ n6813 ^ 1'b0 ;
  assign n18280 = n5747 | n18279 ;
  assign n18277 = n7259 & ~n16069 ;
  assign n18278 = ~n5803 & n18277 ;
  assign n18281 = n18280 ^ n18278 ^ 1'b0 ;
  assign n18282 = n2683 | n14744 ;
  assign n18283 = n8070 & n18282 ;
  assign n18284 = n13685 ^ n334 ^ 1'b0 ;
  assign n18285 = ~n1911 & n18284 ;
  assign n18286 = ~n4808 & n18285 ;
  assign n18287 = ~n3882 & n18286 ;
  assign n18288 = ~n11947 & n18287 ;
  assign n18289 = n13393 & ~n15771 ;
  assign n18290 = n12974 ^ n634 ^ 1'b0 ;
  assign n18291 = n18290 ^ n13059 ^ n2267 ;
  assign n18292 = n150 | n2070 ;
  assign n18293 = ~n6048 & n18292 ;
  assign n18294 = ~n7967 & n9701 ;
  assign n18295 = ~n7908 & n18294 ;
  assign n18296 = n4066 & ~n18295 ;
  assign n18297 = ~n18293 & n18296 ;
  assign n18298 = n8600 | n18297 ;
  assign n18299 = n18298 ^ n2365 ^ 1'b0 ;
  assign n18301 = n7054 & ~n7810 ;
  assign n18302 = n5609 & ~n18301 ;
  assign n18303 = n8420 & n18302 ;
  assign n18300 = ~n1897 & n12390 ;
  assign n18304 = n18303 ^ n18300 ^ 1'b0 ;
  assign n18305 = n1069 & n4116 ;
  assign n18306 = n10832 ^ n5739 ^ 1'b0 ;
  assign n18307 = n16828 & n18306 ;
  assign n18308 = ( ~n10191 & n18305 ) | ( ~n10191 & n18307 ) | ( n18305 & n18307 ) ;
  assign n18309 = ( n8886 & ~n14150 ) | ( n8886 & n16328 ) | ( ~n14150 & n16328 ) ;
  assign n18310 = n7155 ^ n3090 ^ 1'b0 ;
  assign n18311 = n360 | n5027 ;
  assign n18312 = n18310 & ~n18311 ;
  assign n18313 = n1306 | n7329 ;
  assign n18314 = n18312 | n18313 ;
  assign n18315 = n18199 & ~n18314 ;
  assign n18316 = n12406 ^ n6237 ^ 1'b0 ;
  assign n18317 = n18315 | n18316 ;
  assign n18321 = n2460 ^ n2377 ^ 1'b0 ;
  assign n18318 = n2668 & n3080 ;
  assign n18319 = n18318 ^ n6250 ^ 1'b0 ;
  assign n18320 = n4720 & ~n18319 ;
  assign n18322 = n18321 ^ n18320 ^ 1'b0 ;
  assign n18323 = ~n6857 & n11190 ;
  assign n18324 = n18323 ^ n5736 ^ 1'b0 ;
  assign n18325 = n564 & ~n12687 ;
  assign n18326 = ~n4551 & n18325 ;
  assign n18327 = n18324 & n18326 ;
  assign n18328 = n214 & n5355 ;
  assign n18329 = n15115 & n18328 ;
  assign n18330 = ( ~n365 & n2698 ) | ( ~n365 & n11190 ) | ( n2698 & n11190 ) ;
  assign n18331 = ~n7155 & n18330 ;
  assign n18332 = n18331 ^ n16013 ^ 1'b0 ;
  assign n18333 = n458 | n6144 ;
  assign n18334 = n5163 & ~n18333 ;
  assign n18335 = n18334 ^ n11685 ^ 1'b0 ;
  assign n18336 = n11409 | n12677 ;
  assign n18337 = n12666 & ~n18336 ;
  assign n18338 = n18337 ^ n3827 ^ 1'b0 ;
  assign n18341 = n2940 & n6991 ;
  assign n18342 = n3734 & n18341 ;
  assign n18339 = n6392 ^ n3970 ^ 1'b0 ;
  assign n18340 = n13122 | n18339 ;
  assign n18343 = n18342 ^ n18340 ^ n4665 ;
  assign n18344 = n16994 & ~n17203 ;
  assign n18345 = ~n16994 & n18344 ;
  assign n18351 = n2986 & ~n3133 ;
  assign n18346 = ~n1050 & n7495 ;
  assign n18347 = n18346 ^ n2239 ^ 1'b0 ;
  assign n18348 = n1763 | n18347 ;
  assign n18349 = n10826 ^ n2637 ^ 1'b0 ;
  assign n18350 = n18348 & n18349 ;
  assign n18352 = n18351 ^ n18350 ^ 1'b0 ;
  assign n18353 = n9205 ^ n3187 ^ 1'b0 ;
  assign n18354 = n7979 | n15843 ;
  assign n18355 = n18354 ^ n4311 ^ 1'b0 ;
  assign n18356 = ~n2762 & n2986 ;
  assign n18357 = ~n18355 & n18356 ;
  assign n18358 = n11058 ^ n6839 ^ 1'b0 ;
  assign n18359 = n640 | n18358 ;
  assign n18360 = n15066 & ~n18359 ;
  assign n18361 = n2116 ^ n1818 ^ 1'b0 ;
  assign n18362 = ~n16633 & n18361 ;
  assign n18363 = ( n2095 & n6040 ) | ( n2095 & n18362 ) | ( n6040 & n18362 ) ;
  assign n18364 = n18363 ^ n4079 ^ 1'b0 ;
  assign n18365 = n7241 & ~n10298 ;
  assign n18366 = ~n4448 & n18365 ;
  assign n18367 = n18366 ^ n8253 ^ 1'b0 ;
  assign n18368 = n18367 ^ n6846 ^ n1187 ;
  assign n18369 = n3066 & ~n17191 ;
  assign n18370 = n4690 & ~n11524 ;
  assign n18371 = n18370 ^ x11 ^ 1'b0 ;
  assign n18372 = n13298 & ~n18371 ;
  assign n18373 = n6375 & n12638 ;
  assign n18374 = n2504 & n18373 ;
  assign n18375 = n11452 ^ n7710 ^ 1'b0 ;
  assign n18376 = ~n6482 & n18375 ;
  assign n18377 = n18376 ^ n9574 ^ 1'b0 ;
  assign n18378 = n8806 & ~n18377 ;
  assign n18379 = n7164 & n14714 ;
  assign n18380 = n13152 ^ n9703 ^ 1'b0 ;
  assign n18381 = n18380 ^ n14337 ^ 1'b0 ;
  assign n18382 = n1973 ^ n1663 ^ n745 ;
  assign n18383 = n18382 ^ n3044 ^ 1'b0 ;
  assign n18384 = ~n3153 & n18383 ;
  assign n18385 = n18384 ^ n5779 ^ 1'b0 ;
  assign n18386 = n492 & ~n4434 ;
  assign n18387 = n11925 ^ n9291 ^ 1'b0 ;
  assign n18388 = n358 & ~n18387 ;
  assign n18389 = ( ~n255 & n5769 ) | ( ~n255 & n10866 ) | ( n5769 & n10866 ) ;
  assign n18390 = n18389 ^ n7078 ^ 1'b0 ;
  assign n18391 = n706 & n2390 ;
  assign n18392 = ~n2587 & n18391 ;
  assign n18393 = n13520 ^ n7645 ^ 1'b0 ;
  assign n18394 = ~n2356 & n11588 ;
  assign n18395 = n18394 ^ n12909 ^ 1'b0 ;
  assign n18396 = n18393 & n18395 ;
  assign n18397 = n18392 | n18396 ;
  assign n18398 = n18397 ^ n663 ^ 1'b0 ;
  assign n18399 = n8334 & n12938 ;
  assign n18400 = n61 | n7167 ;
  assign n18401 = n18400 ^ n15246 ^ 1'b0 ;
  assign n18402 = n18401 ^ n11318 ^ 1'b0 ;
  assign n18403 = n16793 ^ n179 ^ 1'b0 ;
  assign n18404 = n18402 | n18403 ;
  assign n18405 = n905 & n9657 ;
  assign n18406 = n6419 ^ n3738 ^ 1'b0 ;
  assign n18407 = n18405 & ~n18406 ;
  assign n18408 = n4365 & n5833 ;
  assign n18409 = n4712 & n18408 ;
  assign n18410 = n13521 & ~n18409 ;
  assign n18411 = n7972 & n13537 ;
  assign n18412 = n17864 ^ n14437 ^ 1'b0 ;
  assign n18413 = ~n8347 & n18412 ;
  assign n18414 = n13941 ^ n10492 ^ 1'b0 ;
  assign n18415 = n1790 ^ n584 ^ n257 ;
  assign n18416 = n1810 & n2874 ;
  assign n18417 = ~n1658 & n18416 ;
  assign n18418 = n790 & ~n18417 ;
  assign n18419 = ( ~n3985 & n17401 ) | ( ~n3985 & n18418 ) | ( n17401 & n18418 ) ;
  assign n18420 = n18415 & ~n18419 ;
  assign n18421 = n12756 & n13381 ;
  assign n18422 = n18421 ^ n846 ^ 1'b0 ;
  assign n18423 = ~n17532 & n18422 ;
  assign n18425 = n318 | n749 ;
  assign n18424 = ( n344 & n11196 ) | ( n344 & ~n12890 ) | ( n11196 & ~n12890 ) ;
  assign n18426 = n18425 ^ n18424 ^ n9187 ;
  assign n18427 = n13337 & n18426 ;
  assign n18428 = n18427 ^ n7921 ^ 1'b0 ;
  assign n18429 = n297 & n18428 ;
  assign n18430 = n9284 ^ n3939 ^ 1'b0 ;
  assign n18431 = n10249 ^ n3181 ^ 1'b0 ;
  assign n18432 = n3611 & n16796 ;
  assign n18433 = ~n18431 & n18432 ;
  assign n18434 = n15904 & ~n17788 ;
  assign n18435 = n18434 ^ n11971 ^ 1'b0 ;
  assign n18436 = ~n1883 & n7881 ;
  assign n18437 = ~n1802 & n18436 ;
  assign n18438 = n18011 | n18437 ;
  assign n18439 = ~n18435 & n18438 ;
  assign n18440 = n2998 & n8738 ;
  assign n18441 = n5293 & n18440 ;
  assign n18442 = n5190 | n18441 ;
  assign n18443 = ~n3746 & n17476 ;
  assign n18444 = n3207 & n7125 ;
  assign n18445 = n9215 & n18444 ;
  assign n18446 = n4461 | n18445 ;
  assign n18447 = n16184 ^ n9286 ^ n28 ;
  assign n18448 = n18447 ^ n14068 ^ 1'b0 ;
  assign n18449 = n18446 & n18448 ;
  assign n18450 = n14896 ^ n10480 ^ 1'b0 ;
  assign n18451 = ( n849 & ~n5139 ) | ( n849 & n12006 ) | ( ~n5139 & n12006 ) ;
  assign n18452 = ( ~n14865 & n16507 ) | ( ~n14865 & n18451 ) | ( n16507 & n18451 ) ;
  assign n18453 = n15363 ^ n2994 ^ 1'b0 ;
  assign n18454 = n3592 & ~n15119 ;
  assign n18455 = n199 | n3440 ;
  assign n18456 = n9700 ^ n872 ^ 1'b0 ;
  assign n18457 = n4002 & ~n5089 ;
  assign n18458 = n4760 & n18457 ;
  assign n18459 = n18456 & ~n18458 ;
  assign n18460 = n2178 & n18459 ;
  assign n18462 = n8449 ^ n2338 ^ 1'b0 ;
  assign n18463 = ~n9047 & n18462 ;
  assign n18464 = n8148 & n18463 ;
  assign n18461 = n229 | n8731 ;
  assign n18465 = n18464 ^ n18461 ^ 1'b0 ;
  assign n18466 = n7972 ^ n7516 ^ 1'b0 ;
  assign n18467 = n18466 ^ n18199 ^ 1'b0 ;
  assign n18468 = n13314 & ~n18467 ;
  assign n18469 = n3781 | n10000 ;
  assign n18470 = n7089 & n18469 ;
  assign n18471 = n2666 & n10365 ;
  assign n18472 = n18471 ^ n3985 ^ 1'b0 ;
  assign n18473 = n10393 & ~n11339 ;
  assign n18474 = n14667 ^ n11645 ^ 1'b0 ;
  assign n18475 = n18474 ^ n14059 ^ n4142 ;
  assign n18476 = n1955 | n9128 ;
  assign n18477 = n18476 ^ n18313 ^ 1'b0 ;
  assign n18478 = n3993 | n13375 ;
  assign n18479 = n6228 & ~n18478 ;
  assign n18480 = n3762 | n18479 ;
  assign n18481 = n2319 ^ n1371 ^ 1'b0 ;
  assign n18482 = n14883 ^ n6802 ^ 1'b0 ;
  assign n18483 = n8806 & ~n18482 ;
  assign n18484 = n18481 & n18483 ;
  assign n18485 = n18484 ^ n13809 ^ 1'b0 ;
  assign n18486 = n277 & ~n1414 ;
  assign n18487 = n1876 & n18486 ;
  assign n18488 = n18487 ^ n1679 ^ 1'b0 ;
  assign n18489 = n2336 | n13329 ;
  assign n18490 = n307 & ~n1042 ;
  assign n18491 = n3514 | n18490 ;
  assign n18492 = n18491 ^ n515 ^ 1'b0 ;
  assign n18493 = n6864 ^ n5824 ^ 1'b0 ;
  assign n18494 = n18493 ^ n446 ^ 1'b0 ;
  assign n18495 = n8118 & ~n16057 ;
  assign n18496 = n18494 & n18495 ;
  assign n18497 = n18496 ^ n9078 ^ 1'b0 ;
  assign n18498 = n18492 | n18497 ;
  assign n18499 = ~n7620 & n11477 ;
  assign n18500 = ( n15342 & n18498 ) | ( n15342 & ~n18499 ) | ( n18498 & ~n18499 ) ;
  assign n18501 = n17980 ^ n13000 ^ 1'b0 ;
  assign n18502 = ~n15386 & n18501 ;
  assign n18503 = n6038 | n18348 ;
  assign n18504 = n13685 ^ n11194 ^ 1'b0 ;
  assign n18505 = n18503 | n18504 ;
  assign n18506 = ( n2216 & n4823 ) | ( n2216 & ~n14883 ) | ( n4823 & ~n14883 ) ;
  assign n18507 = n9685 ^ n6678 ^ 1'b0 ;
  assign n18508 = n14029 ^ n5484 ^ 1'b0 ;
  assign n18509 = n2694 ^ n1880 ^ 1'b0 ;
  assign n18510 = n18509 ^ n7541 ^ 1'b0 ;
  assign n18511 = ~n4497 & n5393 ;
  assign n18512 = ~n7377 & n18511 ;
  assign n18513 = n18512 ^ n188 ^ 1'b0 ;
  assign n18514 = n5163 & ~n18513 ;
  assign n18518 = n1306 & ~n5890 ;
  assign n18519 = ~n782 & n18518 ;
  assign n18515 = n1884 | n16050 ;
  assign n18516 = n14795 & n18515 ;
  assign n18517 = n7613 & n18516 ;
  assign n18520 = n18519 ^ n18517 ^ 1'b0 ;
  assign n18521 = n13 | n9056 ;
  assign n18522 = n3255 & ~n18521 ;
  assign n18523 = n18522 ^ n11795 ^ n7724 ;
  assign n18524 = n8639 ^ n387 ^ 1'b0 ;
  assign n18525 = ~n609 & n18524 ;
  assign n18526 = n10059 & n18525 ;
  assign n18527 = n1105 & ~n18526 ;
  assign n18528 = n18527 ^ n3580 ^ 1'b0 ;
  assign n18529 = n3674 & ~n18528 ;
  assign n18530 = n9116 ^ n7741 ^ 1'b0 ;
  assign n18531 = n205 & n225 ;
  assign n18532 = n1075 & ~n18531 ;
  assign n18533 = n18519 & ~n18532 ;
  assign n18534 = n774 & n10112 ;
  assign n18535 = n1915 & ~n6190 ;
  assign n18536 = n8262 | n18535 ;
  assign n18537 = n18534 & ~n18536 ;
  assign n18538 = n2100 | n18537 ;
  assign n18539 = n3049 & ~n8173 ;
  assign n18540 = n18539 ^ n3726 ^ 1'b0 ;
  assign n18541 = n8269 ^ n351 ^ 1'b0 ;
  assign n18542 = n18540 & ~n18541 ;
  assign n18543 = n2989 ^ n1863 ^ 1'b0 ;
  assign n18544 = n1884 | n18543 ;
  assign n18545 = n8176 | n8976 ;
  assign n18546 = n18544 | n18545 ;
  assign n18547 = n18546 ^ n8894 ^ 1'b0 ;
  assign n18548 = n18547 ^ n10277 ^ n1112 ;
  assign n18549 = n18548 ^ n2155 ^ 1'b0 ;
  assign n18550 = n250 & ~n12095 ;
  assign n18551 = n15635 ^ n15364 ^ 1'b0 ;
  assign n18552 = n16536 ^ n10531 ^ 1'b0 ;
  assign n18553 = ~n2081 & n18552 ;
  assign n18554 = n18553 ^ n896 ^ 1'b0 ;
  assign n18555 = n12013 ^ n2248 ^ 1'b0 ;
  assign n18556 = n1230 & ~n18555 ;
  assign n18557 = ~n15359 & n16135 ;
  assign n18558 = n18557 ^ n423 ^ 1'b0 ;
  assign n18559 = n4153 | n18395 ;
  assign n18560 = n2852 & n16012 ;
  assign n18561 = n10572 | n14818 ;
  assign n18562 = n13035 ^ n6683 ^ 1'b0 ;
  assign n18563 = n3282 ^ n2820 ^ 1'b0 ;
  assign n18564 = n18563 ^ n6699 ^ 1'b0 ;
  assign n18565 = n144 | n18080 ;
  assign n18574 = ~n6316 & n9464 ;
  assign n18575 = n4333 & n18574 ;
  assign n18576 = n18575 ^ n1366 ^ 1'b0 ;
  assign n18566 = n6442 & n10287 ;
  assign n18567 = n1378 & ~n3272 ;
  assign n18568 = n1099 | n1785 ;
  assign n18569 = n18568 ^ n5269 ^ 1'b0 ;
  assign n18570 = ~n6100 & n18569 ;
  assign n18571 = n18570 ^ n14518 ^ 1'b0 ;
  assign n18572 = n18567 & n18571 ;
  assign n18573 = ( n10956 & ~n18566 ) | ( n10956 & n18572 ) | ( ~n18566 & n18572 ) ;
  assign n18577 = n18576 ^ n18573 ^ 1'b0 ;
  assign n18578 = n10066 & n18577 ;
  assign n18579 = n732 ^ n604 ^ 1'b0 ;
  assign n18580 = n15147 & n18579 ;
  assign n18581 = ~n13526 & n18580 ;
  assign n18582 = n18581 ^ n7076 ^ 1'b0 ;
  assign n18583 = n18578 & n18582 ;
  assign n18584 = ~n5497 & n10751 ;
  assign n18585 = n18584 ^ n8020 ^ 1'b0 ;
  assign n18586 = n3838 ^ n1036 ^ 1'b0 ;
  assign n18587 = n903 & ~n18586 ;
  assign n18588 = ( ~n2495 & n3919 ) | ( ~n2495 & n18587 ) | ( n3919 & n18587 ) ;
  assign n18589 = n12865 ^ n205 ^ 1'b0 ;
  assign n18590 = ~n4989 & n14429 ;
  assign n18591 = n18590 ^ n249 ^ 1'b0 ;
  assign n18592 = ~n1159 & n1731 ;
  assign n18593 = n18592 ^ n15515 ^ 1'b0 ;
  assign n18594 = ( ~n5607 & n9779 ) | ( ~n5607 & n14642 ) | ( n9779 & n14642 ) ;
  assign n18595 = n6783 ^ n3787 ^ 1'b0 ;
  assign n18596 = n810 & n18595 ;
  assign n18597 = n18596 ^ n7086 ^ 1'b0 ;
  assign n18598 = ~n56 & n14558 ;
  assign n18599 = ~n12330 & n18598 ;
  assign n18600 = ~n12725 & n17348 ;
  assign n18601 = n3414 | n11909 ;
  assign n18602 = n13040 & ~n18601 ;
  assign n18603 = n10093 ^ n5881 ^ 1'b0 ;
  assign n18604 = n7169 ^ n5111 ^ 1'b0 ;
  assign n18605 = n13042 | n18604 ;
  assign n18606 = n2893 & ~n18605 ;
  assign n18607 = ~n13685 & n18606 ;
  assign n18608 = n4875 ^ n983 ^ 1'b0 ;
  assign n18609 = n3845 | n11904 ;
  assign n18610 = n2425 | n18609 ;
  assign n18611 = ~n4983 & n7081 ;
  assign n18612 = n18611 ^ n4952 ^ 1'b0 ;
  assign n18616 = n2626 ^ n2600 ^ 1'b0 ;
  assign n18617 = n333 | n4435 ;
  assign n18618 = n18616 & n18617 ;
  assign n18619 = ~n4921 & n18618 ;
  assign n18613 = n11673 ^ n3272 ^ n519 ;
  assign n18614 = ~n7964 & n18613 ;
  assign n18615 = ~n8868 & n18614 ;
  assign n18620 = n18619 ^ n18615 ^ 1'b0 ;
  assign n18621 = ~n1159 & n1845 ;
  assign n18622 = n3472 | n18621 ;
  assign n18623 = n3359 | n5538 ;
  assign n18624 = n13134 | n18623 ;
  assign n18625 = n11535 & ~n18624 ;
  assign n18630 = ~n1241 & n12074 ;
  assign n18631 = ~n398 & n18630 ;
  assign n18632 = ~n5257 & n14611 ;
  assign n18633 = n18631 & n18632 ;
  assign n18626 = n13042 ^ n12994 ^ n7437 ;
  assign n18627 = n18626 ^ n4091 ^ 1'b0 ;
  assign n18628 = ~n2146 & n18627 ;
  assign n18629 = ~n4784 & n18628 ;
  assign n18634 = n18633 ^ n18629 ^ 1'b0 ;
  assign n18635 = n799 & ~n3372 ;
  assign n18636 = ~n1054 & n18635 ;
  assign n18637 = n11086 ^ n10298 ^ 1'b0 ;
  assign n18641 = ( n1299 & ~n2181 ) | ( n1299 & n4837 ) | ( ~n2181 & n4837 ) ;
  assign n18642 = n1071 & ~n18641 ;
  assign n18638 = ~n466 & n2628 ;
  assign n18639 = n4222 & n18638 ;
  assign n18640 = ( n269 & n6554 ) | ( n269 & ~n18639 ) | ( n6554 & ~n18639 ) ;
  assign n18643 = n18642 ^ n18640 ^ n1570 ;
  assign n18644 = n4136 & n17487 ;
  assign n18645 = n18644 ^ n4599 ^ 1'b0 ;
  assign n18647 = n4388 ^ n4157 ^ 1'b0 ;
  assign n18646 = n11322 & ~n14415 ;
  assign n18648 = n18647 ^ n18646 ^ 1'b0 ;
  assign n18649 = n18648 ^ n12271 ^ 1'b0 ;
  assign n18650 = n8292 | n18649 ;
  assign n18651 = n18650 ^ n723 ^ 1'b0 ;
  assign n18652 = ( n11416 & ~n12466 ) | ( n11416 & n18651 ) | ( ~n12466 & n18651 ) ;
  assign n18653 = n7126 ^ n4698 ^ 1'b0 ;
  assign n18654 = n18653 ^ n10698 ^ 1'b0 ;
  assign n18655 = n738 & n1192 ;
  assign n18656 = ~n1192 & n18655 ;
  assign n18657 = n4389 & ~n18656 ;
  assign n18658 = n14148 & ~n18657 ;
  assign n18659 = n842 & n18658 ;
  assign n18660 = ( n345 & n5443 ) | ( n345 & n9241 ) | ( n5443 & n9241 ) ;
  assign n18661 = n4960 ^ n3706 ^ 1'b0 ;
  assign n18662 = n10423 & n18661 ;
  assign n18663 = ~n18660 & n18662 ;
  assign n18664 = n18663 ^ n15635 ^ 1'b0 ;
  assign n18665 = n17260 ^ n1526 ^ 1'b0 ;
  assign n18666 = ~n6189 & n7139 ;
  assign n18667 = ~n695 & n18666 ;
  assign n18668 = n5778 & n9780 ;
  assign n18669 = ~n7137 & n18668 ;
  assign n18670 = n6111 & n18669 ;
  assign n18671 = n12458 ^ n9023 ^ n1908 ;
  assign n18672 = n11502 & ~n12332 ;
  assign n18673 = ~n666 & n10083 ;
  assign n18674 = n56 | n2833 ;
  assign n18675 = n5997 ^ n5067 ^ n4113 ;
  assign n18676 = n18674 | n18675 ;
  assign n18677 = ( x8 & n16872 ) | ( x8 & ~n18085 ) | ( n16872 & ~n18085 ) ;
  assign n18678 = ~n967 & n3486 ;
  assign n18679 = n5179 ^ n2502 ^ 1'b0 ;
  assign n18680 = n3150 | n18679 ;
  assign n18681 = n25 | n18680 ;
  assign n18682 = n1217 & n1278 ;
  assign n18683 = n3382 & n18682 ;
  assign n18684 = n14190 ^ n1134 ^ 1'b0 ;
  assign n18685 = ~n18683 & n18684 ;
  assign n18686 = ~n2397 & n3611 ;
  assign n18687 = ~n3611 & n18686 ;
  assign n18688 = n107 & n734 ;
  assign n18689 = ~n734 & n18688 ;
  assign n18690 = n1126 | n18689 ;
  assign n18691 = n18689 & ~n18690 ;
  assign n18692 = n169 | n18691 ;
  assign n18693 = n169 & ~n18692 ;
  assign n18694 = n18687 | n18693 ;
  assign n18695 = n18687 & ~n18694 ;
  assign n18696 = ( ~n5167 & n9736 ) | ( ~n5167 & n9848 ) | ( n9736 & n9848 ) ;
  assign n18697 = n13179 ^ n6351 ^ 1'b0 ;
  assign n18698 = n18696 & ~n18697 ;
  assign n18699 = ~n12773 & n18698 ;
  assign n18702 = n1943 & n7635 ;
  assign n18701 = ~n4560 & n12072 ;
  assign n18703 = n18702 ^ n18701 ^ 1'b0 ;
  assign n18700 = n10322 ^ n3262 ^ 1'b0 ;
  assign n18704 = n18703 ^ n18700 ^ 1'b0 ;
  assign n18705 = n1700 & n4928 ;
  assign n18706 = n18705 ^ n989 ^ 1'b0 ;
  assign n18707 = n12005 | n18706 ;
  assign n18708 = n11527 & n18707 ;
  assign n18709 = n18708 ^ n12680 ^ n11703 ;
  assign n18711 = n1141 & ~n7679 ;
  assign n18710 = n5809 & n15322 ;
  assign n18712 = n18711 ^ n18710 ^ 1'b0 ;
  assign n18713 = n2508 & n6609 ;
  assign n18714 = n18713 ^ n16693 ^ 1'b0 ;
  assign n18715 = n2117 & ~n6262 ;
  assign n18716 = ~n15677 & n18715 ;
  assign n18717 = n13210 | n18716 ;
  assign n18718 = n18717 ^ n9289 ^ 1'b0 ;
  assign n18719 = n6406 & n18718 ;
  assign n18720 = n4909 & ~n6339 ;
  assign n18721 = n18720 ^ n5525 ^ 1'b0 ;
  assign n18722 = n8166 | n10173 ;
  assign n18723 = n18722 ^ n7750 ^ 1'b0 ;
  assign n18724 = n18723 ^ n14741 ^ 1'b0 ;
  assign n18725 = n423 | n18724 ;
  assign n18726 = n6350 ^ n4315 ^ 1'b0 ;
  assign n18727 = ( ~n4814 & n15799 ) | ( ~n4814 & n18726 ) | ( n15799 & n18726 ) ;
  assign n18728 = n18727 ^ n7997 ^ 1'b0 ;
  assign n18729 = ~n18725 & n18728 ;
  assign n18730 = n83 & ~n13394 ;
  assign n18731 = ~n5995 & n18730 ;
  assign n18732 = n5146 & ~n18731 ;
  assign n18733 = n1896 | n10443 ;
  assign n18734 = n18733 ^ n8950 ^ 1'b0 ;
  assign n18735 = ~n3430 & n6534 ;
  assign n18736 = ( ~n5313 & n18734 ) | ( ~n5313 & n18735 ) | ( n18734 & n18735 ) ;
  assign n18737 = n12488 ^ n192 ^ 1'b0 ;
  assign n18738 = n13841 & ~n18737 ;
  assign n18739 = n6027 | n13443 ;
  assign n18740 = n9988 & n11025 ;
  assign n18741 = ~n5788 & n11616 ;
  assign n18742 = n9530 | n14523 ;
  assign n18743 = n2133 & ~n18742 ;
  assign n18745 = n2426 & n6259 ;
  assign n18746 = ~n212 & n18745 ;
  assign n18744 = n17008 ^ n13715 ^ n3372 ;
  assign n18747 = n18746 ^ n18744 ^ 1'b0 ;
  assign n18748 = ~n15367 & n18747 ;
  assign n18749 = n862 & n7541 ;
  assign n18750 = n5849 & ~n6291 ;
  assign n18751 = ~n18749 & n18750 ;
  assign n18752 = n8436 & ~n18751 ;
  assign n18753 = n16491 & n18752 ;
  assign n18754 = n9839 ^ n5123 ^ 1'b0 ;
  assign n18755 = n12604 ^ n806 ^ 1'b0 ;
  assign n18756 = n18755 ^ n6347 ^ 1'b0 ;
  assign n18757 = n9588 & n18756 ;
  assign n18758 = ~n4797 & n8124 ;
  assign n18759 = ~n4687 & n18758 ;
  assign n18760 = n2029 & n11599 ;
  assign n18761 = n16289 ^ n12149 ^ n6764 ;
  assign n18762 = n9867 ^ n7844 ^ 1'b0 ;
  assign n18763 = n2708 | n18762 ;
  assign n18764 = ~n2403 & n18763 ;
  assign n18765 = n6280 | n6311 ;
  assign n18766 = n1576 | n18765 ;
  assign n18767 = n18766 ^ n12022 ^ n4712 ;
  assign n18768 = n2900 & ~n11826 ;
  assign n18769 = n1654 & n7686 ;
  assign n18770 = ~n5405 & n18769 ;
  assign n18773 = n6127 | n13495 ;
  assign n18771 = n5967 & n18451 ;
  assign n18772 = ~n6020 & n18771 ;
  assign n18774 = n18773 ^ n18772 ^ 1'b0 ;
  assign n18776 = ~n959 & n1056 ;
  assign n18777 = ~n9102 & n18776 ;
  assign n18775 = ~n4999 & n15312 ;
  assign n18778 = n18777 ^ n18775 ^ 1'b0 ;
  assign n18781 = n33 | n5638 ;
  assign n18779 = n6435 ^ n2975 ^ 1'b0 ;
  assign n18780 = n3687 | n18779 ;
  assign n18782 = n18781 ^ n18780 ^ 1'b0 ;
  assign n18783 = n5406 ^ n3847 ^ 1'b0 ;
  assign n18784 = n18783 ^ n2899 ^ n612 ;
  assign n18785 = n412 & ~n13887 ;
  assign n18786 = n8097 & n18785 ;
  assign n18787 = n2910 & ~n3080 ;
  assign n18788 = n18787 ^ n60 ^ 1'b0 ;
  assign n18789 = n18788 ^ n4324 ^ 1'b0 ;
  assign n18790 = n11404 | n18789 ;
  assign n18791 = ~n822 & n1182 ;
  assign n18792 = n18791 ^ n12535 ^ 1'b0 ;
  assign n18793 = ( n2891 & ~n18790 ) | ( n2891 & n18792 ) | ( ~n18790 & n18792 ) ;
  assign n18794 = n781 & n11543 ;
  assign n18795 = n1763 | n3738 ;
  assign n18796 = n5235 | n18795 ;
  assign n18797 = ( n8924 & n9388 ) | ( n8924 & ~n12000 ) | ( n9388 & ~n12000 ) ;
  assign n18799 = ~n296 & n1715 ;
  assign n18798 = n4344 | n5779 ;
  assign n18800 = n18799 ^ n18798 ^ 1'b0 ;
  assign n18801 = ~n18797 & n18800 ;
  assign n18802 = ~n3595 & n5982 ;
  assign n18803 = n18802 ^ n908 ^ 1'b0 ;
  assign n18804 = n10023 & n13687 ;
  assign n18805 = n7044 ^ n6410 ^ 1'b0 ;
  assign n18806 = n4174 & n18805 ;
  assign n18807 = ~n15119 & n18806 ;
  assign n18808 = n3817 & n5929 ;
  assign n18809 = n1363 & n18808 ;
  assign n18810 = n11613 | n18809 ;
  assign n18811 = n7839 ^ n4740 ^ 1'b0 ;
  assign n18812 = n801 & n18558 ;
  assign n18813 = n3343 & ~n6699 ;
  assign n18814 = n1504 & ~n11857 ;
  assign n18815 = ~n18813 & n18814 ;
  assign n18819 = n3891 & ~n9071 ;
  assign n18820 = n18819 ^ n5222 ^ 1'b0 ;
  assign n18818 = n5345 & n11527 ;
  assign n18821 = n18820 ^ n18818 ^ 1'b0 ;
  assign n18816 = ~n1069 & n10851 ;
  assign n18817 = ~n14744 & n18816 ;
  assign n18822 = n18821 ^ n18817 ^ 1'b0 ;
  assign n18823 = n4643 & ~n18822 ;
  assign n18824 = n15893 ^ n12747 ^ 1'b0 ;
  assign n18825 = n16920 ^ n1042 ^ 1'b0 ;
  assign n18826 = n2721 & ~n18825 ;
  assign n18827 = ~n12537 & n18826 ;
  assign n18830 = n15946 ^ n6362 ^ 1'b0 ;
  assign n18831 = n18830 ^ n14471 ^ 1'b0 ;
  assign n18828 = ( n2533 & n7558 ) | ( n2533 & ~n10396 ) | ( n7558 & ~n10396 ) ;
  assign n18829 = n11744 | n18828 ;
  assign n18832 = n18831 ^ n18829 ^ 1'b0 ;
  assign n18833 = n18832 ^ n7953 ^ 1'b0 ;
  assign n18834 = n15400 ^ n9596 ^ 1'b0 ;
  assign n18835 = n5422 | n18834 ;
  assign n18836 = n18835 ^ n5586 ^ 1'b0 ;
  assign n18837 = n3361 & ~n9906 ;
  assign n18838 = n8068 ^ n7542 ^ 1'b0 ;
  assign n18839 = n998 & n9156 ;
  assign n18840 = n1853 & n18839 ;
  assign n18841 = n18838 & n18840 ;
  assign n18842 = n5517 ^ n1145 ^ 1'b0 ;
  assign n18843 = n15318 & ~n18842 ;
  assign n18844 = ~n6029 & n18843 ;
  assign n18845 = n14092 ^ n8665 ^ n6030 ;
  assign n18846 = n18845 ^ n12067 ^ 1'b0 ;
  assign n18847 = ( n514 & n15205 ) | ( n514 & n15912 ) | ( n15205 & n15912 ) ;
  assign n18848 = n4046 & ~n9002 ;
  assign n18849 = ( n1853 & n3484 ) | ( n1853 & n13375 ) | ( n3484 & n13375 ) ;
  assign n18850 = n5001 & n12558 ;
  assign n18851 = ( n9389 & ~n18849 ) | ( n9389 & n18850 ) | ( ~n18849 & n18850 ) ;
  assign n18852 = n18851 ^ n7360 ^ 1'b0 ;
  assign n18853 = n3110 | n18852 ;
  assign n18854 = n17749 & ~n18853 ;
  assign n18855 = n13538 ^ n6806 ^ 1'b0 ;
  assign n18856 = n817 | n18855 ;
  assign n18857 = n5329 | n12424 ;
  assign n18858 = n15885 | n18857 ;
  assign n18859 = n13264 ^ n10079 ^ 1'b0 ;
  assign n18860 = n18859 ^ n13871 ^ 1'b0 ;
  assign n18861 = n15596 ^ n2545 ^ 1'b0 ;
  assign n18862 = ~n2318 & n5154 ;
  assign n18863 = n15137 & n18862 ;
  assign n18864 = n18861 & n18863 ;
  assign n18866 = n1764 & ~n3039 ;
  assign n18865 = n3903 & n14250 ;
  assign n18867 = n18866 ^ n18865 ^ 1'b0 ;
  assign n18868 = n3848 & ~n5956 ;
  assign n18869 = n4885 & n18868 ;
  assign n18870 = n18869 ^ n10513 ^ 1'b0 ;
  assign n18871 = n18711 ^ n10811 ^ n6278 ;
  assign n18872 = n14493 & n18871 ;
  assign n18873 = n622 | n9153 ;
  assign n18874 = n18232 ^ n2753 ^ 1'b0 ;
  assign n18875 = n18873 | n18874 ;
  assign n18876 = n15029 ^ n754 ^ 1'b0 ;
  assign n18877 = ~n18875 & n18876 ;
  assign n18878 = ~n18872 & n18877 ;
  assign n18879 = n5823 & n17491 ;
  assign n18880 = n18879 ^ n5516 ^ 1'b0 ;
  assign n18881 = ~n5880 & n18880 ;
  assign n18882 = n18881 ^ n7693 ^ n5999 ;
  assign n18883 = ~n2202 & n8901 ;
  assign n18884 = n7247 & ~n18883 ;
  assign n18885 = ( n459 & n1052 ) | ( n459 & n5470 ) | ( n1052 & n5470 ) ;
  assign n18886 = n18885 ^ n1021 ^ 1'b0 ;
  assign n18887 = n14583 & n18886 ;
  assign n18888 = n1721 | n9503 ;
  assign n18889 = n18887 & n18888 ;
  assign n18890 = n12525 & ~n17024 ;
  assign n18891 = n7581 ^ n2112 ^ 1'b0 ;
  assign n18892 = n309 | n18891 ;
  assign n18893 = ~n2056 & n6250 ;
  assign n18894 = n18893 ^ n11902 ^ 1'b0 ;
  assign n18895 = n14753 | n18179 ;
  assign n18896 = n6009 & ~n16870 ;
  assign n18897 = n18896 ^ n608 ^ 1'b0 ;
  assign n18898 = ( n387 & n1603 ) | ( n387 & n2368 ) | ( n1603 & n2368 ) ;
  assign n18899 = n9383 | n18898 ;
  assign n18900 = n5036 & ~n18899 ;
  assign n18901 = n1682 | n3687 ;
  assign n18902 = n18901 ^ n18706 ^ 1'b0 ;
  assign n18903 = n12671 ^ n1199 ^ 1'b0 ;
  assign n18904 = n130 & ~n12703 ;
  assign n18905 = ~n18903 & n18904 ;
  assign n18906 = n15478 ^ n5760 ^ 1'b0 ;
  assign n18907 = n18906 ^ n150 ^ 1'b0 ;
  assign n18908 = n11456 ^ n9305 ^ n2614 ;
  assign n18909 = n18908 ^ n9363 ^ 1'b0 ;
  assign n18910 = ~n5466 & n18909 ;
  assign n18911 = n16419 ^ n14123 ^ n4357 ;
  assign n18912 = n8783 & n18911 ;
  assign n18913 = n989 & ~n9917 ;
  assign n18914 = n13544 ^ n9964 ^ 1'b0 ;
  assign n18915 = n18914 ^ n3876 ^ 1'b0 ;
  assign n18916 = n2634 | n11252 ;
  assign n18917 = n18915 | n18916 ;
  assign n18918 = ~n1852 & n6878 ;
  assign n18919 = n17629 ^ n9343 ^ n8391 ;
  assign n18920 = n16431 & n18234 ;
  assign n18921 = ( n6430 & n10476 ) | ( n6430 & n18920 ) | ( n10476 & n18920 ) ;
  assign n18922 = n7188 | n18921 ;
  assign n18923 = n18919 & ~n18922 ;
  assign n18924 = n8832 & n11445 ;
  assign n18925 = ~n16286 & n18924 ;
  assign n18926 = n8081 ^ n4976 ^ 1'b0 ;
  assign n18927 = ~n8635 & n18926 ;
  assign n18928 = n4947 ^ n3672 ^ n1326 ;
  assign n18929 = n4398 & n18928 ;
  assign n18930 = n14164 & n18222 ;
  assign n18931 = ~n590 & n1800 ;
  assign n18932 = n15547 & n18931 ;
  assign n18933 = n885 & n6989 ;
  assign n18934 = n18932 & n18933 ;
  assign n18935 = n1980 & ~n4572 ;
  assign n18936 = n602 & n18935 ;
  assign n18937 = n9018 | n10149 ;
  assign n18938 = n18936 & ~n18937 ;
  assign n18939 = n12016 ^ n10351 ^ n6213 ;
  assign n18940 = ~n17323 & n18939 ;
  assign n18941 = n12430 ^ n5443 ^ 1'b0 ;
  assign n18942 = n11846 | n15619 ;
  assign n18943 = n18941 | n18942 ;
  assign n18944 = ( n2944 & n5247 ) | ( n2944 & ~n15442 ) | ( n5247 & ~n15442 ) ;
  assign n18945 = n3791 & n4864 ;
  assign n18946 = ~n18944 & n18945 ;
  assign n18947 = n18946 ^ n16954 ^ 1'b0 ;
  assign n18948 = n3881 & ~n18947 ;
  assign n18951 = ~n450 & n5945 ;
  assign n18949 = n379 & n8788 ;
  assign n18950 = ~n132 & n18949 ;
  assign n18952 = n18951 ^ n18950 ^ 1'b0 ;
  assign n18953 = n6291 | n18952 ;
  assign n18954 = n6663 & ~n18953 ;
  assign n18955 = n7734 & n16630 ;
  assign n18956 = ( ~n4506 & n6945 ) | ( ~n4506 & n18315 ) | ( n6945 & n18315 ) ;
  assign n18957 = n11025 | n16743 ;
  assign n18958 = n12299 ^ n4856 ^ 1'b0 ;
  assign n18959 = n8730 | n18958 ;
  assign n18960 = n18959 ^ n3379 ^ 1'b0 ;
  assign n18961 = n7092 ^ n1199 ^ 1'b0 ;
  assign n18962 = ( n3049 & ~n16896 ) | ( n3049 & n18961 ) | ( ~n16896 & n18961 ) ;
  assign n18963 = n2808 & ~n7462 ;
  assign n18964 = ( n6553 & ~n18962 ) | ( n6553 & n18963 ) | ( ~n18962 & n18963 ) ;
  assign n18965 = n1947 & ~n18964 ;
  assign n18966 = n1758 | n7146 ;
  assign n18967 = ~n5300 & n9170 ;
  assign n18968 = n18967 ^ n5165 ^ 1'b0 ;
  assign n18969 = n2634 & n18968 ;
  assign n18970 = n18969 ^ n10549 ^ 1'b0 ;
  assign n18971 = n10702 | n18970 ;
  assign n18972 = n2900 & ~n13021 ;
  assign n18973 = ~n3838 & n18972 ;
  assign n18974 = n18973 ^ n1562 ^ 1'b0 ;
  assign n18975 = n14405 & n18974 ;
  assign n18976 = n2077 & n4690 ;
  assign n18977 = n18976 ^ n11327 ^ 1'b0 ;
  assign n18978 = n1143 | n4745 ;
  assign n18979 = n18977 | n18978 ;
  assign n18980 = n18975 | n18979 ;
  assign n18981 = ( n4767 & n6294 ) | ( n4767 & n11826 ) | ( n6294 & n11826 ) ;
  assign n18982 = n7685 | n18981 ;
  assign n18983 = n8979 ^ n2091 ^ 1'b0 ;
  assign n18984 = ~n334 & n18983 ;
  assign n18985 = n18984 ^ n16421 ^ 1'b0 ;
  assign n18986 = n441 & n18985 ;
  assign n18987 = n3476 & n18986 ;
  assign n18988 = n18987 ^ n17528 ^ 1'b0 ;
  assign n18989 = n17297 ^ n456 ^ 1'b0 ;
  assign n18990 = n18004 ^ n2093 ^ 1'b0 ;
  assign n18991 = n10253 ^ n28 ^ 1'b0 ;
  assign n18992 = n883 | n6296 ;
  assign n18993 = n5719 | n14330 ;
  assign n18994 = n1924 & ~n18993 ;
  assign n18995 = ( n8863 & ~n11240 ) | ( n8863 & n14766 ) | ( ~n11240 & n14766 ) ;
  assign n18996 = n179 & n15854 ;
  assign n18997 = ( n810 & n6723 ) | ( n810 & n7747 ) | ( n6723 & n7747 ) ;
  assign n18998 = n18997 ^ n7895 ^ 1'b0 ;
  assign n18999 = ( n3054 & n12990 ) | ( n3054 & n18998 ) | ( n12990 & n18998 ) ;
  assign n19000 = n14979 ^ n3446 ^ 1'b0 ;
  assign n19001 = n13040 | n19000 ;
  assign n19002 = n6589 ^ n2943 ^ n1915 ;
  assign n19003 = n19002 ^ n6161 ^ 1'b0 ;
  assign n19004 = ( n5584 & n6397 ) | ( n5584 & ~n19003 ) | ( n6397 & ~n19003 ) ;
  assign n19005 = n13887 ^ n4185 ^ 1'b0 ;
  assign n19006 = n1736 | n19005 ;
  assign n19007 = n1293 | n13279 ;
  assign n19008 = ( n10530 & n10846 ) | ( n10530 & ~n19007 ) | ( n10846 & ~n19007 ) ;
  assign n19009 = n13346 & ~n19008 ;
  assign n19010 = ~n9698 & n19009 ;
  assign n19011 = n10223 & ~n14248 ;
  assign n19012 = n19010 & n19011 ;
  assign n19013 = n19012 ^ n1200 ^ 1'b0 ;
  assign n19014 = n15388 ^ n4010 ^ 1'b0 ;
  assign n19015 = n8287 & ~n19014 ;
  assign n19016 = n19015 ^ n13985 ^ 1'b0 ;
  assign n19017 = n4208 & ~n9563 ;
  assign n19018 = ~n11787 & n19017 ;
  assign n19019 = n7725 | n19018 ;
  assign n19020 = n9068 ^ n936 ^ 1'b0 ;
  assign n19021 = n5518 & ~n19020 ;
  assign n19022 = ~n5755 & n19021 ;
  assign n19023 = n10796 | n19022 ;
  assign n19024 = n19019 & ~n19023 ;
  assign n19025 = n15007 ^ n5998 ^ 1'b0 ;
  assign n19026 = n18662 & n19025 ;
  assign n19027 = n19026 ^ n5128 ^ 1'b0 ;
  assign n19028 = n9605 ^ n2539 ^ 1'b0 ;
  assign n19029 = n9641 & ~n12829 ;
  assign n19030 = n19029 ^ n6350 ^ 1'b0 ;
  assign n19031 = n14462 ^ n515 ^ 1'b0 ;
  assign n19032 = n19030 & n19031 ;
  assign n19033 = n13350 & n19032 ;
  assign n19034 = n13802 & n19033 ;
  assign n19035 = n12695 ^ n1674 ^ 1'b0 ;
  assign n19036 = ~n12332 & n19035 ;
  assign n19037 = n6111 | n16321 ;
  assign n19038 = n16382 ^ n12261 ^ 1'b0 ;
  assign n19039 = n12380 ^ n7549 ^ 1'b0 ;
  assign n19040 = n3833 & ~n19039 ;
  assign n19044 = ~n40 & n826 ;
  assign n19043 = ~n666 & n12472 ;
  assign n19045 = n19044 ^ n19043 ^ 1'b0 ;
  assign n19041 = ~n5825 & n8278 ;
  assign n19042 = n19041 ^ n18744 ^ 1'b0 ;
  assign n19046 = n19045 ^ n19042 ^ 1'b0 ;
  assign n19049 = n261 & ~n8949 ;
  assign n19050 = n1079 & n19049 ;
  assign n19047 = n6182 ^ n543 ^ 1'b0 ;
  assign n19048 = n5304 & n19047 ;
  assign n19051 = n19050 ^ n19048 ^ 1'b0 ;
  assign n19052 = n10085 & n19051 ;
  assign n19053 = ~n14731 & n19052 ;
  assign n19054 = n19053 ^ n12625 ^ n7523 ;
  assign n19055 = ~n1918 & n17946 ;
  assign n19056 = n18603 & n19055 ;
  assign n19057 = n10549 ^ n2533 ^ 1'b0 ;
  assign n19058 = n7458 & n19057 ;
  assign n19059 = n19058 ^ n2914 ^ 1'b0 ;
  assign n19060 = ~n11074 & n19059 ;
  assign n19061 = n10797 & n15355 ;
  assign n19062 = n13004 & ~n19061 ;
  assign n19063 = n19062 ^ n3320 ^ n1134 ;
  assign n19064 = ~n8147 & n11411 ;
  assign n19065 = n9703 & n19064 ;
  assign n19066 = n19065 ^ n16236 ^ 1'b0 ;
  assign n19067 = n19066 ^ n8872 ^ 1'b0 ;
  assign n19068 = ~n12514 & n15388 ;
  assign n19069 = n19068 ^ n3933 ^ 1'b0 ;
  assign n19070 = ( ~n10162 & n11593 ) | ( ~n10162 & n19069 ) | ( n11593 & n19069 ) ;
  assign n19071 = n11033 & ~n19070 ;
  assign n19072 = n19071 ^ n5940 ^ 1'b0 ;
  assign n19073 = n12039 | n12911 ;
  assign n19074 = n16491 ^ n15716 ^ 1'b0 ;
  assign n19075 = n4484 ^ n1450 ^ 1'b0 ;
  assign n19076 = n905 | n19075 ;
  assign n19077 = n649 & ~n5352 ;
  assign n19078 = n3708 & n19077 ;
  assign n19079 = n4100 | n4515 ;
  assign n19080 = n4241 & ~n10354 ;
  assign n19081 = n19080 ^ n9004 ^ 1'b0 ;
  assign n19082 = n3461 ^ n1441 ^ 1'b0 ;
  assign n19083 = n7520 & ~n19082 ;
  assign n19084 = n16379 & ~n19083 ;
  assign n19085 = n802 & n4525 ;
  assign n19086 = n3947 ^ n419 ^ 1'b0 ;
  assign n19089 = n18903 ^ n5149 ^ 1'b0 ;
  assign n19090 = n3169 | n19089 ;
  assign n19091 = ~n6096 & n8630 ;
  assign n19092 = n19091 ^ n5393 ^ 1'b0 ;
  assign n19093 = n19090 | n19092 ;
  assign n19087 = ~n2382 & n5001 ;
  assign n19088 = n19087 ^ n18093 ^ 1'b0 ;
  assign n19094 = n19093 ^ n19088 ^ 1'b0 ;
  assign n19095 = n8403 ^ n3442 ^ 1'b0 ;
  assign n19096 = ( n4646 & ~n6941 ) | ( n4646 & n10628 ) | ( ~n6941 & n10628 ) ;
  assign n19097 = n19096 ^ n5508 ^ 1'b0 ;
  assign n19098 = n13566 | n17919 ;
  assign n19099 = n2353 & ~n3927 ;
  assign n19100 = n19099 ^ n959 ^ 1'b0 ;
  assign n19101 = n707 | n10537 ;
  assign n19102 = n19101 ^ n10944 ^ 1'b0 ;
  assign n19103 = n16450 ^ n10114 ^ 1'b0 ;
  assign n19104 = n4567 | n19103 ;
  assign n19105 = n19102 & n19104 ;
  assign n19106 = ~n2652 & n6001 ;
  assign n19107 = n19106 ^ n13638 ^ 1'b0 ;
  assign n19108 = n15976 & n19060 ;
  assign n19109 = n19108 ^ n4681 ^ n1918 ;
  assign n19110 = ~n5214 & n8275 ;
  assign n19111 = n2356 ^ n2332 ^ 1'b0 ;
  assign n19112 = n493 & n19111 ;
  assign n19113 = n2640 | n19112 ;
  assign n19114 = n1554 & n19113 ;
  assign n19115 = n10262 & n19114 ;
  assign n19116 = ( n1144 & n19110 ) | ( n1144 & n19115 ) | ( n19110 & n19115 ) ;
  assign n19117 = n15566 ^ n7875 ^ n1905 ;
  assign n19118 = n7338 ^ n6189 ^ 1'b0 ;
  assign n19119 = n19117 | n19118 ;
  assign n19120 = n19119 ^ n14712 ^ 1'b0 ;
  assign n19121 = n120 & ~n211 ;
  assign n19122 = ~n120 & n19121 ;
  assign n19123 = n640 | n19122 ;
  assign n19124 = n19122 & ~n19123 ;
  assign n19125 = n4725 & ~n19124 ;
  assign n19126 = ~n4725 & n19125 ;
  assign n19127 = n13350 ^ n9768 ^ 1'b0 ;
  assign n19128 = n13050 & n19127 ;
  assign n19129 = n14068 ^ n7121 ^ 1'b0 ;
  assign n19130 = n14126 ^ n7358 ^ 1'b0 ;
  assign n19131 = n4010 | n19130 ;
  assign n19132 = n2158 ^ n2029 ^ 1'b0 ;
  assign n19133 = ~n13124 & n19132 ;
  assign n19134 = n3223 & n19133 ;
  assign n19135 = ~n3867 & n19134 ;
  assign n19136 = ( n1767 & ~n7618 ) | ( n1767 & n19135 ) | ( ~n7618 & n19135 ) ;
  assign n19142 = n5259 | n14758 ;
  assign n19137 = x2 & n285 ;
  assign n19138 = ~n285 & n19137 ;
  assign n19139 = n1192 & ~n4819 ;
  assign n19140 = ~n1192 & n19139 ;
  assign n19141 = n19138 | n19140 ;
  assign n19143 = n19142 ^ n19141 ^ 1'b0 ;
  assign n19144 = n5458 ^ n5059 ^ 1'b0 ;
  assign n19145 = n8779 ^ n1267 ^ 1'b0 ;
  assign n19146 = n3409 | n19145 ;
  assign n19147 = n19146 ^ n7894 ^ 1'b0 ;
  assign n19148 = n19144 & ~n19147 ;
  assign n19149 = n19148 ^ n11547 ^ 1'b0 ;
  assign n19150 = n5859 ^ n296 ^ 1'b0 ;
  assign n19151 = ~n1908 & n19150 ;
  assign n19152 = n18519 | n19151 ;
  assign n19153 = n6988 & ~n19152 ;
  assign n19154 = n2382 | n12717 ;
  assign n19155 = n5811 & ~n19154 ;
  assign n19156 = ~n9434 & n10388 ;
  assign n19157 = n19155 & n19156 ;
  assign n19158 = n19157 ^ n901 ^ 1'b0 ;
  assign n19159 = n19110 ^ n878 ^ 1'b0 ;
  assign n19160 = n15316 ^ n5073 ^ n944 ;
  assign n19161 = n16555 ^ n3998 ^ 1'b0 ;
  assign n19162 = n7335 ^ n6697 ^ 1'b0 ;
  assign n19163 = ~n8297 & n19162 ;
  assign n19164 = n4738 | n19163 ;
  assign n19165 = n3843 | n10552 ;
  assign n19166 = n4074 ^ n3634 ^ 1'b0 ;
  assign n19167 = ~n11474 & n19166 ;
  assign n19168 = n19167 ^ n13 ^ 1'b0 ;
  assign n19169 = ~n19165 & n19168 ;
  assign n19170 = n19169 ^ n2219 ^ 1'b0 ;
  assign n19171 = n19170 ^ n12804 ^ 1'b0 ;
  assign n19172 = n19164 & n19171 ;
  assign n19173 = n10300 ^ n6004 ^ 1'b0 ;
  assign n19174 = n1173 | n1714 ;
  assign n19175 = n4747 | n19174 ;
  assign n19176 = n19175 ^ n244 ^ 1'b0 ;
  assign n19177 = n3449 | n19176 ;
  assign n19178 = n19177 ^ n2975 ^ 1'b0 ;
  assign n19179 = n2685 | n3889 ;
  assign n19180 = n1895 | n19179 ;
  assign n19181 = n1217 & ~n17871 ;
  assign n19182 = n19181 ^ n5458 ^ 1'b0 ;
  assign n19183 = n11294 & ~n19182 ;
  assign n19184 = ~n19180 & n19183 ;
  assign n19187 = n16111 ^ n8355 ^ 1'b0 ;
  assign n19185 = n2764 & ~n3492 ;
  assign n19186 = n5037 & n19185 ;
  assign n19188 = n19187 ^ n19186 ^ n3759 ;
  assign n19189 = ~n8553 & n18454 ;
  assign n19190 = n17829 ^ n9464 ^ n8259 ;
  assign n19191 = n16295 | n17971 ;
  assign n19192 = n5997 ^ n1781 ^ 1'b0 ;
  assign n19193 = n2694 | n6892 ;
  assign n19194 = n17818 ^ n4964 ^ 1'b0 ;
  assign n19195 = n8608 & ~n19194 ;
  assign n19196 = n5503 & n10394 ;
  assign n19197 = n19195 & ~n19196 ;
  assign n19198 = n19193 & n19197 ;
  assign n19199 = n19198 ^ n5973 ^ 1'b0 ;
  assign n19200 = n19192 & ~n19199 ;
  assign n19202 = ~n261 & n7247 ;
  assign n19203 = n9868 & n19202 ;
  assign n19201 = ~n764 & n6427 ;
  assign n19204 = n19203 ^ n19201 ^ 1'b0 ;
  assign n19205 = n7355 & ~n19204 ;
  assign n19206 = n19205 ^ n4504 ^ 1'b0 ;
  assign n19207 = ( n782 & n4018 ) | ( n782 & ~n5001 ) | ( n4018 & ~n5001 ) ;
  assign n19208 = n19207 ^ n4742 ^ 1'b0 ;
  assign n19209 = n9867 | n17753 ;
  assign n19210 = n19209 ^ n12654 ^ 1'b0 ;
  assign n19211 = n3939 & ~n14047 ;
  assign n19212 = ~n19210 & n19211 ;
  assign n19213 = n18743 ^ n2581 ^ 1'b0 ;
  assign n19214 = n12319 & n19213 ;
  assign n19215 = ( n188 & n2641 ) | ( n188 & n7140 ) | ( n2641 & n7140 ) ;
  assign n19216 = n19215 ^ n1806 ^ 1'b0 ;
  assign n19217 = n6762 ^ n3849 ^ 1'b0 ;
  assign n19218 = n15287 | n19217 ;
  assign n19219 = n8967 & ~n14327 ;
  assign n19220 = x11 & n1476 ;
  assign n19221 = n7848 | n17683 ;
  assign n19222 = n827 & ~n2395 ;
  assign n19223 = n6226 & ~n10428 ;
  assign n19224 = ~n19222 & n19223 ;
  assign n19225 = n19224 ^ n7647 ^ 1'b0 ;
  assign n19226 = n19225 ^ n14261 ^ 1'b0 ;
  assign n19227 = n18648 | n19226 ;
  assign n19228 = n19227 ^ n9957 ^ 1'b0 ;
  assign n19229 = n919 & ~n1211 ;
  assign n19230 = n1491 | n10528 ;
  assign n19231 = n4720 | n19230 ;
  assign n19232 = n6881 | n7003 ;
  assign n19233 = n6655 & ~n19232 ;
  assign n19234 = n6876 & ~n7136 ;
  assign n19235 = n7917 ^ n790 ^ 1'b0 ;
  assign n19236 = ~n1031 & n7919 ;
  assign n19237 = n14676 & n19236 ;
  assign n19238 = n2522 | n12731 ;
  assign n19239 = n1365 & ~n19170 ;
  assign n19240 = n12993 & n19239 ;
  assign n19241 = ~n3412 & n4497 ;
  assign n19242 = n7582 & n19241 ;
  assign n19243 = n19242 ^ n7824 ^ 1'b0 ;
  assign n19244 = n14369 | n16111 ;
  assign n19245 = n19244 ^ n49 ^ 1'b0 ;
  assign n19246 = n6947 | n19245 ;
  assign n19247 = n135 | n379 ;
  assign n19248 = n16833 ^ n14602 ^ 1'b0 ;
  assign n19249 = n209 & ~n3245 ;
  assign n19250 = ~n3327 & n11278 ;
  assign n19251 = ~n19249 & n19250 ;
  assign n19252 = n12950 | n15544 ;
  assign n19253 = n3488 & ~n9047 ;
  assign n19254 = n10888 & n19253 ;
  assign n19255 = n757 | n5874 ;
  assign n19256 = n15811 ^ n10041 ^ 1'b0 ;
  assign n19257 = n19256 ^ n1745 ^ 1'b0 ;
  assign n19258 = n2588 & ~n5885 ;
  assign n19259 = n19258 ^ n666 ^ 1'b0 ;
  assign n19260 = n5645 ^ n3072 ^ 1'b0 ;
  assign n19261 = n19259 & ~n19260 ;
  assign n19262 = n10786 ^ n6353 ^ n1267 ;
  assign n19263 = ( n11322 & ~n17050 ) | ( n11322 & n19262 ) | ( ~n17050 & n19262 ) ;
  assign n19264 = n8789 ^ n1430 ^ 1'b0 ;
  assign n19265 = n16028 & n19264 ;
  assign n19267 = n10300 ^ n5505 ^ 1'b0 ;
  assign n19266 = ~n1235 & n7873 ;
  assign n19268 = n19267 ^ n19266 ^ 1'b0 ;
  assign n19269 = n15887 ^ n13281 ^ 1'b0 ;
  assign n19270 = n12604 ^ n2006 ^ 1'b0 ;
  assign n19271 = ( n2634 & n5077 ) | ( n2634 & n11927 ) | ( n5077 & n11927 ) ;
  assign n19272 = n2505 & n18641 ;
  assign n19273 = ~n150 & n19272 ;
  assign n19274 = n19271 | n19273 ;
  assign n19275 = n19274 ^ n459 ^ 1'b0 ;
  assign n19279 = n2058 & ~n3676 ;
  assign n19276 = n760 & ~n12501 ;
  assign n19277 = n1574 & n19276 ;
  assign n19278 = n19277 ^ n7082 ^ n2778 ;
  assign n19280 = n19279 ^ n19278 ^ n11793 ;
  assign n19281 = n19280 ^ n18808 ^ 1'b0 ;
  assign n19282 = n828 & ~n10121 ;
  assign n19283 = n19282 ^ n4993 ^ 1'b0 ;
  assign n19284 = n17318 ^ n9440 ^ 1'b0 ;
  assign n19285 = ~n19283 & n19284 ;
  assign n19286 = ~n18135 & n19285 ;
  assign n19287 = n1093 & n19286 ;
  assign n19288 = n4615 | n9863 ;
  assign n19289 = n3462 ^ n1933 ^ 1'b0 ;
  assign n19290 = n528 ^ n463 ^ 1'b0 ;
  assign n19291 = n3740 ^ n2405 ^ 1'b0 ;
  assign n19292 = n8407 & ~n19291 ;
  assign n19293 = n19290 & n19292 ;
  assign n19294 = n963 ^ n188 ^ 1'b0 ;
  assign n19295 = n8071 | n19294 ;
  assign n19296 = n19295 ^ n9522 ^ 1'b0 ;
  assign n19297 = ~n1023 & n19296 ;
  assign n19298 = n2317 | n19005 ;
  assign n19299 = n19298 ^ n10507 ^ 1'b0 ;
  assign n19300 = n19297 | n19299 ;
  assign n19301 = n3372 | n15692 ;
  assign n19302 = n19301 ^ n8680 ^ 1'b0 ;
  assign n19303 = n19302 ^ n2614 ^ 1'b0 ;
  assign n19304 = n1546 & ~n19303 ;
  assign n19305 = n6647 ^ n1717 ^ 1'b0 ;
  assign n19306 = n2129 | n11797 ;
  assign n19307 = n19306 ^ n6282 ^ 1'b0 ;
  assign n19308 = n19305 | n19307 ;
  assign n19309 = n9688 ^ n666 ^ 1'b0 ;
  assign n19310 = n277 & n19309 ;
  assign n19311 = n12995 ^ n6342 ^ 1'b0 ;
  assign n19314 = n5188 | n15824 ;
  assign n19315 = n16162 | n19314 ;
  assign n19312 = n3770 | n12007 ;
  assign n19313 = n19312 ^ n13108 ^ n6722 ;
  assign n19316 = n19315 ^ n19313 ^ 1'b0 ;
  assign n19317 = n15844 & ~n19316 ;
  assign n19318 = n18834 ^ n16305 ^ 1'b0 ;
  assign n19319 = n1356 | n13068 ;
  assign n19320 = n2334 & n19319 ;
  assign n19321 = n19320 ^ n10286 ^ 1'b0 ;
  assign n19322 = n19052 ^ n6699 ^ 1'b0 ;
  assign n19323 = n6820 ^ n1853 ^ 1'b0 ;
  assign n19324 = ~n1771 & n19323 ;
  assign n19325 = ~n931 & n19324 ;
  assign n19326 = ~n1771 & n4386 ;
  assign n19327 = n19326 ^ n18963 ^ 1'b0 ;
  assign n19330 = n2614 ^ n813 ^ 1'b0 ;
  assign n19328 = n8172 ^ n4935 ^ 1'b0 ;
  assign n19329 = ~n10698 & n19328 ;
  assign n19331 = n19330 ^ n19329 ^ 1'b0 ;
  assign n19332 = n10611 & ~n19331 ;
  assign n19333 = n13486 ^ n8779 ^ 1'b0 ;
  assign n19334 = ~n10299 & n19333 ;
  assign n19335 = n19332 & n19334 ;
  assign n19336 = ~n5505 & n19335 ;
  assign n19337 = n98 | n17538 ;
  assign n19338 = n17026 | n19337 ;
  assign n19339 = n19338 ^ n8336 ^ 1'b0 ;
  assign n19340 = n19339 ^ n7256 ^ 1'b0 ;
  assign n19341 = ~n11524 & n19340 ;
  assign n19342 = n5570 & n11355 ;
  assign n19343 = ~n4540 & n19342 ;
  assign n19344 = n4231 & n19343 ;
  assign n19345 = n19344 ^ n16126 ^ n13098 ;
  assign n19346 = ~n4883 & n7020 ;
  assign n19347 = n19346 ^ n2202 ^ 1'b0 ;
  assign n19348 = n11852 | n19347 ;
  assign n19349 = ~n14226 & n19348 ;
  assign n19350 = n2317 & ~n5338 ;
  assign n19351 = n19350 ^ n10253 ^ 1'b0 ;
  assign n19352 = n3780 & n19351 ;
  assign n19353 = n15417 & n19352 ;
  assign n19354 = n1943 | n16721 ;
  assign n19355 = ~n1781 & n4329 ;
  assign n19356 = n19355 ^ n2082 ^ 1'b0 ;
  assign n19357 = n8291 | n9995 ;
  assign n19358 = n27 | n19357 ;
  assign n19359 = n12586 & ~n13927 ;
  assign n19360 = n88 & n9564 ;
  assign n19361 = n2539 & ~n19360 ;
  assign n19362 = n7116 & n19361 ;
  assign n19363 = n2124 ^ n1178 ^ 1'b0 ;
  assign n19364 = n19363 ^ n6219 ^ 1'b0 ;
  assign n19365 = n6804 ^ n4139 ^ n2555 ;
  assign n19366 = n19365 ^ n2388 ^ 1'b0 ;
  assign n19367 = n19364 & ~n19366 ;
  assign n19369 = n5544 & ~n5642 ;
  assign n19368 = ( ~n7188 & n13032 ) | ( ~n7188 & n15569 ) | ( n13032 & n15569 ) ;
  assign n19370 = n19369 ^ n19368 ^ 1'b0 ;
  assign n19371 = n11757 ^ n3695 ^ 1'b0 ;
  assign n19372 = ( n8704 & ~n13127 ) | ( n8704 & n19371 ) | ( ~n13127 & n19371 ) ;
  assign n19373 = n299 & n5491 ;
  assign n19374 = n19373 ^ n16028 ^ 1'b0 ;
  assign n19375 = n6660 ^ n1694 ^ 1'b0 ;
  assign n19376 = ~n16663 & n19375 ;
  assign n19377 = n1241 & ~n1875 ;
  assign n19378 = n6915 ^ n6248 ^ 1'b0 ;
  assign n19379 = n2612 | n6138 ;
  assign n19380 = n43 | n19379 ;
  assign n19381 = n1908 & n19380 ;
  assign n19382 = n19381 ^ n6009 ^ 1'b0 ;
  assign n19383 = n1096 & ~n19382 ;
  assign n19384 = ~n1293 & n6047 ;
  assign n19385 = n19384 ^ n8443 ^ 1'b0 ;
  assign n19386 = n8812 ^ n2762 ^ 1'b0 ;
  assign n19387 = n1040 ^ n696 ^ 1'b0 ;
  assign n19388 = n2349 | n19387 ;
  assign n19389 = n14560 & ~n19388 ;
  assign n19390 = n19389 ^ n10946 ^ n1562 ;
  assign n19391 = n12233 & ~n17509 ;
  assign n19392 = n19391 ^ n5078 ^ 1'b0 ;
  assign n19393 = ( n147 & n1837 ) | ( n147 & ~n2926 ) | ( n1837 & ~n2926 ) ;
  assign n19394 = n8855 & ~n19393 ;
  assign n19395 = n16185 & ~n17658 ;
  assign n19396 = n9150 | n10259 ;
  assign n19398 = n4376 | n6470 ;
  assign n19399 = n19398 ^ n3459 ^ 1'b0 ;
  assign n19400 = n19399 ^ n14006 ^ n8436 ;
  assign n19397 = n3759 ^ n3008 ^ 1'b0 ;
  assign n19401 = n19400 ^ n19397 ^ 1'b0 ;
  assign n19402 = n15301 ^ n5130 ^ n1235 ;
  assign n19403 = n2108 & n3186 ;
  assign n19404 = n19403 ^ n3926 ^ 1'b0 ;
  assign n19405 = n19404 ^ n17108 ^ 1'b0 ;
  assign n19406 = n19402 | n19405 ;
  assign n19407 = n7624 & n11404 ;
  assign n19408 = n36 & ~n3543 ;
  assign n19409 = n8019 & ~n19408 ;
  assign n19410 = n511 | n19409 ;
  assign n19411 = n19410 ^ n18861 ^ 1'b0 ;
  assign n19412 = ( n2384 & ~n6512 ) | ( n2384 & n19411 ) | ( ~n6512 & n19411 ) ;
  assign n19413 = n11727 | n15232 ;
  assign n19414 = n19413 ^ n4858 ^ 1'b0 ;
  assign n19415 = n8946 ^ n1469 ^ 1'b0 ;
  assign n19416 = ~n9085 & n19415 ;
  assign n19417 = n7589 ^ n4221 ^ 1'b0 ;
  assign n19418 = n1851 | n19417 ;
  assign n19419 = n19416 & n19418 ;
  assign n19420 = n610 ^ n74 ^ 1'b0 ;
  assign n19421 = n3085 | n19420 ;
  assign n19422 = n19421 ^ n2583 ^ 1'b0 ;
  assign n19423 = n4053 ^ n3522 ^ n722 ;
  assign n19424 = n11759 & ~n19423 ;
  assign n19425 = n13189 & n19424 ;
  assign n19426 = n4477 | n9668 ;
  assign n19427 = n19426 ^ n15946 ^ 1'b0 ;
  assign n19428 = n13507 ^ n4171 ^ 1'b0 ;
  assign n19429 = ~n19427 & n19428 ;
  assign n19430 = n19429 ^ n18222 ^ 1'b0 ;
  assign n19431 = n9321 ^ n4207 ^ 1'b0 ;
  assign n19432 = n11243 & ~n19431 ;
  assign n19433 = n8061 & ~n10728 ;
  assign n19434 = n19433 ^ n17891 ^ n9720 ;
  assign n19435 = n1510 & ~n3840 ;
  assign n19436 = n2024 & n19435 ;
  assign n19437 = n19434 & ~n19436 ;
  assign n19438 = n19437 ^ n7062 ^ n3441 ;
  assign n19439 = ( n1104 & n19432 ) | ( n1104 & n19438 ) | ( n19432 & n19438 ) ;
  assign n19440 = ~n10498 & n12625 ;
  assign n19441 = ~n3240 & n11961 ;
  assign n19442 = ~n17032 & n19441 ;
  assign n19443 = n14670 ^ n10085 ^ 1'b0 ;
  assign n19444 = ~n10170 & n19443 ;
  assign n19445 = n19444 ^ n16490 ^ 1'b0 ;
  assign n19446 = n7967 | n14009 ;
  assign n19447 = n19446 ^ n17070 ^ 1'b0 ;
  assign n19448 = n17404 | n19447 ;
  assign n19450 = ( n551 & ~n2155 ) | ( n551 & n10778 ) | ( ~n2155 & n10778 ) ;
  assign n19451 = ~n8915 & n19450 ;
  assign n19449 = n12546 ^ n8222 ^ 1'b0 ;
  assign n19452 = n19451 ^ n19449 ^ 1'b0 ;
  assign n19453 = ~n717 & n12408 ;
  assign n19454 = n8000 & n9604 ;
  assign n19455 = ~n9091 & n19454 ;
  assign n19456 = ~n8269 & n19455 ;
  assign n19457 = n10752 ^ n1217 ^ 1'b0 ;
  assign n19458 = n19456 & n19457 ;
  assign n19459 = n7523 ^ n5015 ^ 1'b0 ;
  assign n19460 = ~n18626 & n19459 ;
  assign n19461 = n18510 & n19460 ;
  assign n19462 = ~n997 & n1000 ;
  assign n19463 = n19462 ^ n3437 ^ 1'b0 ;
  assign n19464 = n12996 ^ n7658 ^ 1'b0 ;
  assign n19465 = ( ~n12147 & n19463 ) | ( ~n12147 & n19464 ) | ( n19463 & n19464 ) ;
  assign n19466 = n19465 ^ n14593 ^ 1'b0 ;
  assign n19468 = ( n142 & n9249 ) | ( n142 & ~n15119 ) | ( n9249 & ~n15119 ) ;
  assign n19467 = n3258 & n3582 ;
  assign n19469 = n19468 ^ n19467 ^ 1'b0 ;
  assign n19470 = n255 & ~n18184 ;
  assign n19471 = n7062 & n19470 ;
  assign n19472 = ~n5353 & n8973 ;
  assign n19473 = n19472 ^ n12549 ^ n9080 ;
  assign n19474 = ~n17023 & n18915 ;
  assign n19475 = ~n19339 & n19474 ;
  assign n19476 = n15240 ^ n10196 ^ 1'b0 ;
  assign n19477 = ~n19475 & n19476 ;
  assign n19478 = n17298 ^ n6406 ^ 1'b0 ;
  assign n19479 = ( n2054 & n3370 ) | ( n2054 & ~n8303 ) | ( n3370 & ~n8303 ) ;
  assign n19480 = ~n5767 & n19479 ;
  assign n19481 = n11109 | n19480 ;
  assign n19482 = n19481 ^ n1430 ^ 1'b0 ;
  assign n19483 = n4038 & ~n19482 ;
  assign n19484 = n19483 ^ n16391 ^ 1'b0 ;
  assign n19485 = n3915 | n19484 ;
  assign n19486 = n14114 ^ n8350 ^ 1'b0 ;
  assign n19487 = n6201 ^ n2587 ^ 1'b0 ;
  assign n19488 = ~n1096 & n19487 ;
  assign n19489 = n8206 & n19488 ;
  assign n19490 = n6096 | n8315 ;
  assign n19491 = n19489 | n19490 ;
  assign n19492 = n11079 & n17610 ;
  assign n19493 = ~n8771 & n18900 ;
  assign n19494 = n4726 & ~n16861 ;
  assign n19495 = ~n12002 & n19494 ;
  assign n19496 = n2808 & n10065 ;
  assign n19497 = n12612 | n19496 ;
  assign n19498 = n19165 & ~n19497 ;
  assign n19499 = n6522 & n15043 ;
  assign n19500 = n15882 ^ n9208 ^ 1'b0 ;
  assign n19501 = n2944 & n5401 ;
  assign n19502 = n19501 ^ n7297 ^ 1'b0 ;
  assign n19503 = n6888 | n13910 ;
  assign n19504 = ~n18124 & n19503 ;
  assign n19505 = n18048 ^ n978 ^ 1'b0 ;
  assign n19506 = ~n19504 & n19505 ;
  assign n19507 = n19506 ^ n5186 ^ 1'b0 ;
  assign n19508 = n11261 ^ n7651 ^ 1'b0 ;
  assign n19509 = n6128 & ~n19508 ;
  assign n19510 = ~n14663 & n19509 ;
  assign n19511 = n6749 & n19510 ;
  assign n19512 = n19511 ^ n12003 ^ 1'b0 ;
  assign n19513 = n19512 ^ n17380 ^ n8635 ;
  assign n19514 = n666 & n19513 ;
  assign n19515 = n8608 ^ n3730 ^ 1'b0 ;
  assign n19516 = n6635 & n9842 ;
  assign n19517 = ~n3243 & n19516 ;
  assign n19518 = n19517 ^ n13520 ^ 1'b0 ;
  assign n19519 = n13432 ^ n11409 ^ 1'b0 ;
  assign n19520 = ~n162 & n2918 ;
  assign n19521 = n1821 ^ n1504 ^ 1'b0 ;
  assign n19522 = n18958 | n19521 ;
  assign n19523 = n19520 | n19522 ;
  assign n19524 = n459 & ~n3974 ;
  assign n19525 = ( n4082 & ~n13850 ) | ( n4082 & n19524 ) | ( ~n13850 & n19524 ) ;
  assign n19526 = ( n1880 & n2192 ) | ( n1880 & ~n8181 ) | ( n2192 & ~n8181 ) ;
  assign n19527 = ~n3036 & n15319 ;
  assign n19528 = n19527 ^ n8165 ^ 1'b0 ;
  assign n19529 = n19526 | n19528 ;
  assign n19532 = n18328 & n18941 ;
  assign n19533 = n19532 ^ n98 ^ 1'b0 ;
  assign n19534 = n1962 & n19533 ;
  assign n19535 = ( ~n1993 & n15142 ) | ( ~n1993 & n19534 ) | ( n15142 & n19534 ) ;
  assign n19530 = n10403 ^ n5890 ^ n3892 ;
  assign n19531 = n13181 & ~n19530 ;
  assign n19536 = n19535 ^ n19531 ^ 1'b0 ;
  assign n19537 = ( n10898 & ~n13232 ) | ( n10898 & n14272 ) | ( ~n13232 & n14272 ) ;
  assign n19538 = n17829 | n19537 ;
  assign n19539 = ~n1653 & n6449 ;
  assign n19540 = n10730 & n19539 ;
  assign n19541 = n19540 ^ n8229 ^ 1'b0 ;
  assign n19542 = n7164 & ~n19541 ;
  assign n19543 = n11251 | n14573 ;
  assign n19544 = ~n3853 & n18347 ;
  assign n19545 = n2130 & ~n2525 ;
  assign n19546 = n19545 ^ n296 ^ 1'b0 ;
  assign n19547 = n9650 & n19546 ;
  assign n19548 = ~n7036 & n19547 ;
  assign n19549 = n10039 & ~n19548 ;
  assign n19550 = ~n19257 & n19549 ;
  assign n19551 = n142 & ~n13004 ;
  assign n19552 = n10420 ^ n5651 ^ n3277 ;
  assign n19553 = n10161 & n14665 ;
  assign n19554 = n19552 & n19553 ;
  assign n19555 = n15348 ^ n2645 ^ 1'b0 ;
  assign n19556 = n3372 | n4017 ;
  assign n19557 = n19556 ^ n1411 ^ 1'b0 ;
  assign n19558 = n14728 & n19557 ;
  assign n19559 = ~n19555 & n19558 ;
  assign n19560 = ~n16690 & n19559 ;
  assign n19561 = ~n423 & n854 ;
  assign n19562 = n4236 & n19561 ;
  assign n19563 = n1522 & n19562 ;
  assign n19564 = n94 & ~n19563 ;
  assign n19565 = ~n1437 & n12640 ;
  assign n19566 = n6124 & n19565 ;
  assign n19567 = n6937 ^ n1469 ^ 1'b0 ;
  assign n19568 = n19566 | n19567 ;
  assign n19569 = ( ~n8647 & n9687 ) | ( ~n8647 & n10209 ) | ( n9687 & n10209 ) ;
  assign n19570 = n12690 ^ n11829 ^ 1'b0 ;
  assign n19571 = n9611 | n19570 ;
  assign n19572 = n16129 ^ n3930 ^ 1'b0 ;
  assign n19573 = n11890 & n19572 ;
  assign n19574 = n19195 ^ n16546 ^ n1943 ;
  assign n19575 = n2919 | n19574 ;
  assign n19576 = n11356 | n19575 ;
  assign n19577 = n14498 ^ n6749 ^ 1'b0 ;
  assign n19578 = n4817 & ~n19577 ;
  assign n19579 = n19578 ^ n9760 ^ 1'b0 ;
  assign n19580 = n2170 | n7829 ;
  assign n19581 = n19580 ^ n6509 ^ 1'b0 ;
  assign n19582 = n6458 ^ n1090 ^ 1'b0 ;
  assign n19583 = ~n16678 & n19582 ;
  assign n19584 = n19583 ^ n13201 ^ 1'b0 ;
  assign n19585 = n19584 ^ n5880 ^ 1'b0 ;
  assign n19586 = n5516 | n19585 ;
  assign n19587 = ( ~n401 & n14835 ) | ( ~n401 & n17077 ) | ( n14835 & n17077 ) ;
  assign n19588 = n15317 & ~n16853 ;
  assign n19589 = n395 & ~n12380 ;
  assign n19590 = n19589 ^ n3300 ^ 1'b0 ;
  assign n19591 = ( n631 & ~n14735 ) | ( n631 & n19590 ) | ( ~n14735 & n19590 ) ;
  assign n19592 = n4128 & n8082 ;
  assign n19593 = n9006 & n19592 ;
  assign n19594 = n2749 & n13901 ;
  assign n19595 = n19594 ^ n2185 ^ 1'b0 ;
  assign n19596 = n19595 ^ n6311 ^ 1'b0 ;
  assign n19597 = n16600 | n19596 ;
  assign n19598 = n19593 & ~n19597 ;
  assign n19599 = n10747 ^ n9773 ^ 1'b0 ;
  assign n19600 = n19568 & n19599 ;
  assign n19601 = ~n5812 & n9831 ;
  assign n19602 = n11440 & n14842 ;
  assign n19603 = n7569 & n13744 ;
  assign n19604 = n6494 ^ n972 ^ 1'b0 ;
  assign n19605 = n4547 & ~n19604 ;
  assign n19606 = n11009 & n19605 ;
  assign n19607 = ~n8246 & n19606 ;
  assign n19608 = ~n1588 & n5616 ;
  assign n19609 = n11618 & n15854 ;
  assign n19610 = n8058 ^ n7233 ^ n4629 ;
  assign n19611 = n19610 ^ n4241 ^ 1'b0 ;
  assign n19612 = n11932 ^ n9542 ^ n5990 ;
  assign n19613 = ~n16016 & n19612 ;
  assign n19614 = n3936 ^ n1756 ^ 1'b0 ;
  assign n19615 = ~n8180 & n19614 ;
  assign n19617 = n1654 | n8553 ;
  assign n19616 = n640 | n10626 ;
  assign n19618 = n19617 ^ n19616 ^ 1'b0 ;
  assign n19619 = n1325 | n19618 ;
  assign n19620 = n19619 ^ n3785 ^ 1'b0 ;
  assign n19621 = n18351 | n19620 ;
  assign n19622 = ~n541 & n5048 ;
  assign n19623 = ~n19621 & n19622 ;
  assign n19624 = n14744 & n19623 ;
  assign n19625 = n3734 | n13130 ;
  assign n19626 = n19625 ^ n870 ^ 1'b0 ;
  assign n19627 = n2012 ^ n1716 ^ 1'b0 ;
  assign n19628 = n19627 ^ n6102 ^ 1'b0 ;
  assign n19629 = n14951 & ~n19628 ;
  assign n19630 = n19629 ^ n2802 ^ 1'b0 ;
  assign n19631 = n9864 & ~n19630 ;
  assign n19632 = ~n7040 & n15049 ;
  assign n19633 = n19632 ^ n12058 ^ n1196 ;
  assign n19634 = ~n8461 & n19633 ;
  assign n19635 = n15460 ^ n14978 ^ 1'b0 ;
  assign n19638 = n6704 | n6889 ;
  assign n19636 = ~n5893 & n9663 ;
  assign n19637 = ~n17226 & n19636 ;
  assign n19639 = n19638 ^ n19637 ^ 1'b0 ;
  assign n19640 = n17723 | n19639 ;
  assign n19641 = n4969 ^ n3738 ^ 1'b0 ;
  assign n19642 = ~n10264 & n19641 ;
  assign n19643 = n19642 ^ n3393 ^ 1'b0 ;
  assign n19644 = n14582 ^ n7591 ^ 1'b0 ;
  assign n19646 = n5139 & ~n8604 ;
  assign n19647 = ~n3158 & n19646 ;
  assign n19645 = n5063 ^ n3465 ^ n1178 ;
  assign n19648 = n19647 ^ n19645 ^ 1'b0 ;
  assign n19649 = n4583 & n8689 ;
  assign n19650 = n19648 & n19649 ;
  assign n19651 = ( n5008 & ~n6980 ) | ( n5008 & n9024 ) | ( ~n6980 & n9024 ) ;
  assign n19652 = n61 & n1033 ;
  assign n19653 = ~n19651 & n19652 ;
  assign n19654 = n14785 & ~n16509 ;
  assign n19655 = n19654 ^ n16220 ^ 1'b0 ;
  assign n19657 = n6450 ^ n2376 ^ 1'b0 ;
  assign n19658 = n13026 & n19657 ;
  assign n19659 = n19658 ^ n1050 ^ 1'b0 ;
  assign n19656 = n439 & ~n12667 ;
  assign n19660 = n19659 ^ n19656 ^ 1'b0 ;
  assign n19661 = n17105 | n19660 ;
  assign n19662 = n4635 ^ n2177 ^ 1'b0 ;
  assign n19663 = n4436 & ~n4850 ;
  assign n19664 = ( n4143 & n11719 ) | ( n4143 & n19663 ) | ( n11719 & n19663 ) ;
  assign n19665 = n5953 | n12405 ;
  assign n19666 = n3687 | n19665 ;
  assign n19667 = n5592 | n19666 ;
  assign n19670 = n770 ^ n687 ^ 1'b0 ;
  assign n19671 = n18301 | n19670 ;
  assign n19668 = n16943 ^ n5685 ^ 1'b0 ;
  assign n19669 = n443 | n19668 ;
  assign n19672 = n19671 ^ n19669 ^ n6894 ;
  assign n19673 = n10971 & ~n15184 ;
  assign n19674 = n2238 & n19673 ;
  assign n19675 = n10211 & n16319 ;
  assign n19676 = n7266 | n8124 ;
  assign n19677 = n19676 ^ n12357 ^ 1'b0 ;
  assign n19678 = n1202 & ~n7696 ;
  assign n19679 = ~n12503 & n19678 ;
  assign n19680 = n1590 | n19679 ;
  assign n19681 = n2893 & n19680 ;
  assign n19682 = n18220 ^ n16283 ^ 1'b0 ;
  assign n19683 = n12847 | n19682 ;
  assign n19684 = n5067 & n5123 ;
  assign n19685 = n19684 ^ n3652 ^ 1'b0 ;
  assign n19686 = n7109 ^ n243 ^ 1'b0 ;
  assign n19687 = ~n10057 & n19686 ;
  assign n19688 = n774 & n7042 ;
  assign n19689 = n7908 & n19688 ;
  assign n19690 = n1057 & n19689 ;
  assign n19691 = n16460 ^ n13311 ^ 1'b0 ;
  assign n19692 = n19691 ^ n2236 ^ 1'b0 ;
  assign n19693 = n19690 | n19692 ;
  assign n19695 = ~n2602 & n16270 ;
  assign n19696 = n19695 ^ n3484 ^ 1'b0 ;
  assign n19694 = n12074 & ~n15420 ;
  assign n19697 = n19696 ^ n19694 ^ 1'b0 ;
  assign n19698 = ~n9358 & n19697 ;
  assign n19699 = n19698 ^ n4762 ^ 1'b0 ;
  assign n19700 = n942 ^ n752 ^ 1'b0 ;
  assign n19701 = n4930 & ~n19700 ;
  assign n19702 = n6037 ^ n2852 ^ 1'b0 ;
  assign n19703 = ( n3320 & ~n4374 ) | ( n3320 & n8685 ) | ( ~n4374 & n8685 ) ;
  assign n19704 = n5468 ^ n1600 ^ 1'b0 ;
  assign n19705 = n6314 & ~n19704 ;
  assign n19706 = n8973 ^ n3440 ^ 1'b0 ;
  assign n19707 = n7690 & ~n19706 ;
  assign n19708 = n19707 ^ n11407 ^ 1'b0 ;
  assign n19709 = ~n19705 & n19708 ;
  assign n19710 = n19709 ^ n4102 ^ 1'b0 ;
  assign n19711 = ~n2388 & n6716 ;
  assign n19712 = ~n3987 & n19711 ;
  assign n19713 = n17118 ^ n5057 ^ 1'b0 ;
  assign n19714 = n5857 & ~n6042 ;
  assign n19715 = n5304 & ~n6806 ;
  assign n19716 = n19714 & n19715 ;
  assign n19717 = n2247 & ~n19716 ;
  assign n19718 = ~n3125 & n19717 ;
  assign n19720 = n5052 | n13562 ;
  assign n19719 = ~n5981 & n6250 ;
  assign n19721 = n19720 ^ n19719 ^ 1'b0 ;
  assign n19722 = ~n5641 & n5765 ;
  assign n19723 = n19722 ^ n2349 ^ 1'b0 ;
  assign n19724 = ~n6583 & n14561 ;
  assign n19725 = ~n1080 & n19724 ;
  assign n19726 = n14662 ^ n5378 ^ 1'b0 ;
  assign n19727 = n10913 & ~n16225 ;
  assign n19728 = n1964 & ~n9833 ;
  assign n19729 = n19726 & n19728 ;
  assign n19730 = n18297 ^ n7633 ^ 1'b0 ;
  assign n19731 = ~n5468 & n19730 ;
  assign n19732 = n19731 ^ n10910 ^ 1'b0 ;
  assign n19733 = n15265 ^ n6600 ^ 1'b0 ;
  assign n19734 = n1038 & n19733 ;
  assign n19735 = n5141 & n9736 ;
  assign n19736 = ~n9067 & n19735 ;
  assign n19737 = n11243 | n19736 ;
  assign n19738 = n16161 | n18635 ;
  assign n19739 = ( n2423 & n11363 ) | ( n2423 & ~n15413 ) | ( n11363 & ~n15413 ) ;
  assign n19740 = ( n4422 & ~n14196 ) | ( n4422 & n19739 ) | ( ~n14196 & n19739 ) ;
  assign n19741 = n18933 ^ n9256 ^ n7133 ;
  assign n19742 = n11162 & ~n19741 ;
  assign n19743 = n19742 ^ n4969 ^ 1'b0 ;
  assign n19744 = n19743 ^ n16565 ^ 1'b0 ;
  assign n19745 = n11960 ^ n1466 ^ 1'b0 ;
  assign n19746 = n7685 ^ n7243 ^ 1'b0 ;
  assign n19747 = ~n4301 & n19746 ;
  assign n19748 = n16784 | n19747 ;
  assign n19749 = n1199 | n19748 ;
  assign n19750 = n4902 | n11724 ;
  assign n19751 = n9832 ^ n1747 ^ 1'b0 ;
  assign n19752 = ( n1615 & ~n9929 ) | ( n1615 & n19751 ) | ( ~n9929 & n19751 ) ;
  assign n19753 = n12274 & ~n16398 ;
  assign n19754 = n11969 ^ n2938 ^ 1'b0 ;
  assign n19755 = n2771 ^ n1344 ^ 1'b0 ;
  assign n19756 = n19755 ^ n18135 ^ 1'b0 ;
  assign n19757 = ~n1040 & n1852 ;
  assign n19758 = n3198 & ~n13747 ;
  assign n19759 = n19758 ^ n6345 ^ 1'b0 ;
  assign n19760 = ( ~n2226 & n6096 ) | ( ~n2226 & n8265 ) | ( n6096 & n8265 ) ;
  assign n19761 = n3833 & ~n7827 ;
  assign n19762 = ~n7016 & n19761 ;
  assign n19763 = n18587 ^ n16206 ^ 1'b0 ;
  assign n19764 = n19762 | n19763 ;
  assign n19765 = n1434 | n4893 ;
  assign n19766 = n11107 | n19765 ;
  assign n19767 = n14825 & ~n19766 ;
  assign n19768 = n10170 ^ n7621 ^ 1'b0 ;
  assign n19769 = ~n14739 & n19768 ;
  assign n19770 = n8376 ^ n7414 ^ 1'b0 ;
  assign n19771 = n12389 & n19770 ;
  assign n19772 = n4034 ^ n432 ^ 1'b0 ;
  assign n19773 = ( n7627 & ~n19771 ) | ( n7627 & n19772 ) | ( ~n19771 & n19772 ) ;
  assign n19774 = ( n1469 & n12471 ) | ( n1469 & n19773 ) | ( n12471 & n19773 ) ;
  assign n19775 = ( n677 & ~n2526 ) | ( n677 & n19774 ) | ( ~n2526 & n19774 ) ;
  assign n19776 = ~n3050 & n8919 ;
  assign n19777 = n6262 & n6527 ;
  assign n19778 = n19777 ^ n9071 ^ 1'b0 ;
  assign n19779 = n588 | n10682 ;
  assign n19780 = n19779 ^ n17113 ^ 1'b0 ;
  assign n19786 = n7063 ^ n2796 ^ 1'b0 ;
  assign n19781 = ~n4757 & n14963 ;
  assign n19782 = n1800 & n19781 ;
  assign n19783 = ~n12643 & n19782 ;
  assign n19784 = n19783 ^ n11098 ^ 1'b0 ;
  assign n19785 = n1025 & n19784 ;
  assign n19787 = n19786 ^ n19785 ^ 1'b0 ;
  assign n19788 = n3300 | n12847 ;
  assign n19789 = n6866 ^ n4340 ^ 1'b0 ;
  assign n19790 = n16561 & n19144 ;
  assign n19791 = ~n6993 & n19790 ;
  assign n19792 = n11230 ^ n8130 ^ 1'b0 ;
  assign n19793 = n1016 & n19792 ;
  assign n19794 = n6975 | n19793 ;
  assign n19795 = n19794 ^ n10663 ^ 1'b0 ;
  assign n19796 = n14867 ^ n5699 ^ 1'b0 ;
  assign n19797 = ( n3132 & n3874 ) | ( n3132 & n7042 ) | ( n3874 & n7042 ) ;
  assign n19798 = n19797 ^ n9645 ^ n9437 ;
  assign n19799 = n19798 ^ n13056 ^ 1'b0 ;
  assign n19800 = n11595 ^ n8870 ^ 1'b0 ;
  assign n19801 = n1269 & n19800 ;
  assign n19802 = n9192 ^ n1260 ^ 1'b0 ;
  assign n19803 = n10769 ^ n1360 ^ 1'b0 ;
  assign n19804 = n4027 | n19803 ;
  assign n19805 = n3086 ^ n1326 ^ 1'b0 ;
  assign n19806 = n8608 & ~n19805 ;
  assign n19807 = n17388 & n19806 ;
  assign n19808 = n7485 ^ n326 ^ 1'b0 ;
  assign n19809 = n13290 | n19808 ;
  assign n19810 = n13257 ^ n7895 ^ n2691 ;
  assign n19811 = ~n1571 & n12289 ;
  assign n19812 = n15951 ^ n8118 ^ 1'b0 ;
  assign n19813 = n8301 & ~n19812 ;
  assign n19814 = n209 & ~n414 ;
  assign n19815 = n19814 ^ n3638 ^ 1'b0 ;
  assign n19816 = n8165 & n19815 ;
  assign n19817 = n7935 ^ n5604 ^ 1'b0 ;
  assign n19818 = n229 | n19817 ;
  assign n19819 = n19818 ^ n7479 ^ 1'b0 ;
  assign n19820 = n6907 & n19819 ;
  assign n19821 = n15165 ^ n9842 ^ n681 ;
  assign n19822 = n19821 ^ n15782 ^ 1'b0 ;
  assign n19823 = n8965 & n19822 ;
  assign n19824 = n19823 ^ n14152 ^ 1'b0 ;
  assign n19825 = n4528 & n8531 ;
  assign n19826 = ~n910 & n19825 ;
  assign n19827 = n1431 ^ n1114 ^ 1'b0 ;
  assign n19828 = n19827 ^ n15533 ^ n15049 ;
  assign n19829 = ~n3121 & n16016 ;
  assign n19830 = n9267 ^ n6302 ^ 1'b0 ;
  assign n19833 = n1528 & n4040 ;
  assign n19834 = n19833 ^ n264 ^ 1'b0 ;
  assign n19835 = n19834 ^ n7268 ^ 1'b0 ;
  assign n19832 = n2770 ^ n100 ^ 1'b0 ;
  assign n19831 = ~n40 & n1141 ;
  assign n19836 = n19835 ^ n19832 ^ n19831 ;
  assign n19837 = n9288 ^ n5658 ^ 1'b0 ;
  assign n19838 = n19837 ^ n13992 ^ 1'b0 ;
  assign n19839 = n7240 & n19838 ;
  assign n19842 = n17711 ^ n2010 ^ 1'b0 ;
  assign n19840 = n88 & n11841 ;
  assign n19841 = ( n13496 & ~n16854 ) | ( n13496 & n19840 ) | ( ~n16854 & n19840 ) ;
  assign n19843 = n19842 ^ n19841 ^ 1'b0 ;
  assign n19844 = n423 | n1167 ;
  assign n19845 = ~n17470 & n19844 ;
  assign n19846 = n19845 ^ n13726 ^ 1'b0 ;
  assign n19847 = n6858 ^ n1730 ^ n220 ;
  assign n19848 = n3112 & ~n11723 ;
  assign n19849 = n19848 ^ n10298 ^ 1'b0 ;
  assign n19850 = n2961 | n3981 ;
  assign n19851 = n33 & ~n19850 ;
  assign n19852 = n9026 | n19851 ;
  assign n19853 = n4331 | n19852 ;
  assign n19854 = ~n10713 & n19853 ;
  assign n19855 = n999 | n2332 ;
  assign n19856 = n999 & ~n19855 ;
  assign n19857 = ~n105 & n19856 ;
  assign n19858 = n4034 & n19857 ;
  assign n19859 = n12962 & ~n19858 ;
  assign n19860 = ~n17899 & n19859 ;
  assign n19861 = n19860 ^ n15567 ^ 1'b0 ;
  assign n19862 = n49 & n239 ;
  assign n19863 = ~n239 & n19862 ;
  assign n19864 = n7765 | n19863 ;
  assign n19865 = n19863 & ~n19864 ;
  assign n19866 = n840 | n1210 ;
  assign n19867 = n1210 & ~n19866 ;
  assign n19868 = n15685 & ~n19867 ;
  assign n19869 = n19865 & n19868 ;
  assign n19870 = n5715 | n19869 ;
  assign n19871 = n5715 & ~n19870 ;
  assign n19872 = n19861 & ~n19871 ;
  assign n19873 = ~n19861 & n19872 ;
  assign n19874 = n10759 | n19873 ;
  assign n19875 = n19873 & ~n19874 ;
  assign n19876 = n12441 ^ n10675 ^ n4442 ;
  assign n19877 = ~n2640 & n13212 ;
  assign n19878 = ~n3759 & n19877 ;
  assign n19879 = n19876 & ~n19878 ;
  assign n19880 = ( ~n9770 & n19368 ) | ( ~n9770 & n19879 ) | ( n19368 & n19879 ) ;
  assign n19881 = n8656 | n12906 ;
  assign n19882 = n2381 | n15521 ;
  assign n19883 = ~n3110 & n8408 ;
  assign n19884 = n19883 ^ n10368 ^ 1'b0 ;
  assign n19885 = n6781 & n11499 ;
  assign n19886 = ~n2754 & n19885 ;
  assign n19887 = n302 & ~n3716 ;
  assign n19888 = n19887 ^ n15144 ^ 1'b0 ;
  assign n19889 = ( n4710 & n8907 ) | ( n4710 & ~n19888 ) | ( n8907 & ~n19888 ) ;
  assign n19890 = n19889 ^ n19069 ^ 1'b0 ;
  assign n19891 = ~n2159 & n4555 ;
  assign n19892 = n18803 ^ n14225 ^ 1'b0 ;
  assign n19893 = n9731 ^ n3019 ^ 1'b0 ;
  assign n19894 = n19893 ^ n9726 ^ 1'b0 ;
  assign n19895 = n12226 | n19894 ;
  assign n19896 = n1723 & n11374 ;
  assign n19897 = n2998 & n3173 ;
  assign n19898 = n446 & ~n5727 ;
  assign n19899 = ~n2090 & n19898 ;
  assign n19900 = ~n17823 & n19899 ;
  assign n19901 = ~n19897 & n19900 ;
  assign n19902 = n3647 & n19901 ;
  assign n19903 = n817 | n4540 ;
  assign n19904 = ~n11353 & n19903 ;
  assign n19905 = n19904 ^ n13062 ^ 1'b0 ;
  assign n19906 = n3072 ^ n2873 ^ 1'b0 ;
  assign n19907 = n17583 ^ n15293 ^ 1'b0 ;
  assign n19908 = n7020 & n9271 ;
  assign n19909 = ~n1170 & n3483 ;
  assign n19910 = n2225 & n8908 ;
  assign n19911 = n3031 ^ n1905 ^ 1'b0 ;
  assign n19912 = ( n5886 & n10102 ) | ( n5886 & n11404 ) | ( n10102 & n11404 ) ;
  assign n19913 = n19912 ^ n10420 ^ 1'b0 ;
  assign n19914 = n19913 ^ n17481 ^ 1'b0 ;
  assign n19915 = n19911 | n19914 ;
  assign n19916 = ~n12197 & n16627 ;
  assign n19917 = n4238 | n4276 ;
  assign n19918 = n19917 ^ n10193 ^ 1'b0 ;
  assign n19919 = n16506 ^ n9254 ^ 1'b0 ;
  assign n19920 = n12260 ^ n2441 ^ 1'b0 ;
  assign n19921 = ( ~n4622 & n6861 ) | ( ~n4622 & n19920 ) | ( n6861 & n19920 ) ;
  assign n19922 = n2787 | n15035 ;
  assign n19923 = n7207 | n19922 ;
  assign n19924 = n12617 & n19923 ;
  assign n19925 = ~n19921 & n19924 ;
  assign n19926 = n3891 & n15424 ;
  assign n19927 = n5305 & ~n17774 ;
  assign n19928 = n1079 & n1321 ;
  assign n19929 = n19928 ^ n7118 ^ 1'b0 ;
  assign n19930 = n3514 | n3665 ;
  assign n19931 = ~n8251 & n9746 ;
  assign n19932 = n19931 ^ n12776 ^ n6213 ;
  assign n19933 = n5473 & n9331 ;
  assign n19934 = ( n8233 & n14506 ) | ( n8233 & ~n19933 ) | ( n14506 & ~n19933 ) ;
  assign n19935 = n19934 ^ n1944 ^ 1'b0 ;
  assign n19936 = n5867 & ~n10073 ;
  assign n19937 = n150 & n19936 ;
  assign n19938 = ~n961 & n6548 ;
  assign n19939 = n19938 ^ n1685 ^ 1'b0 ;
  assign n19940 = n12409 & n19939 ;
  assign n19941 = n19940 ^ n19762 ^ 1'b0 ;
  assign n19942 = n1192 & n14842 ;
  assign n19943 = n16249 ^ n1652 ^ 1'b0 ;
  assign n19944 = ~n983 & n6337 ;
  assign n19945 = n19944 ^ n1510 ^ 1'b0 ;
  assign n19946 = n19945 ^ n4296 ^ 1'b0 ;
  assign n19947 = n2775 & n19946 ;
  assign n19948 = n10620 & n13599 ;
  assign n19949 = n19948 ^ n12921 ^ 1'b0 ;
  assign n19950 = n1062 | n1418 ;
  assign n19951 = n1062 & ~n19950 ;
  assign n19952 = n220 & n19951 ;
  assign n19953 = n12799 | n19952 ;
  assign n19954 = n12799 & ~n19953 ;
  assign n19955 = n4863 & ~n19954 ;
  assign n19956 = n19954 & n19955 ;
  assign n19957 = n19956 ^ n18493 ^ 1'b0 ;
  assign n19958 = n18700 & n19957 ;
  assign n19959 = n7554 ^ n3665 ^ 1'b0 ;
  assign n19960 = n19959 ^ n944 ^ 1'b0 ;
  assign n19961 = n2403 & ~n19960 ;
  assign n19962 = n522 & ~n4760 ;
  assign n19963 = ~n5323 & n19962 ;
  assign n19964 = n11761 & ~n19963 ;
  assign n19965 = n1834 | n4327 ;
  assign n19966 = n5936 | n19965 ;
  assign n19967 = n19966 ^ n15492 ^ n4879 ;
  assign n19968 = n4276 | n19967 ;
  assign n19969 = n17674 & ~n19968 ;
  assign n19970 = n5755 & ~n9090 ;
  assign n19971 = n4004 | n14008 ;
  assign n19972 = n13739 & ~n19971 ;
  assign n19973 = n19972 ^ n9322 ^ n7802 ;
  assign n19974 = ~n19970 & n19973 ;
  assign n19975 = n19974 ^ n15155 ^ 1'b0 ;
  assign n19976 = n13063 & n19975 ;
  assign n19977 = n8037 & ~n15635 ;
  assign n19978 = n19977 ^ n15367 ^ 1'b0 ;
  assign n19979 = ~n2468 & n5912 ;
  assign n19980 = n19978 & n19979 ;
  assign n19981 = n13390 & n18041 ;
  assign n19982 = ~n6942 & n9941 ;
  assign n19983 = n19982 ^ n9441 ^ 1'b0 ;
  assign n19984 = n10839 ^ n9754 ^ 1'b0 ;
  assign n19985 = n15152 ^ n8659 ^ n6028 ;
  assign n19986 = ~n959 & n7410 ;
  assign n19987 = n19985 & n19986 ;
  assign n19988 = ~n8660 & n14733 ;
  assign n19989 = n19988 ^ n12057 ^ 1'b0 ;
  assign n19990 = n12690 ^ n10505 ^ 1'b0 ;
  assign n19991 = n8823 & ~n19990 ;
  assign n19992 = n16453 ^ n3259 ^ n2079 ;
  assign n19993 = n8478 & ~n9492 ;
  assign n19994 = ( n7197 & n13042 ) | ( n7197 & ~n19746 ) | ( n13042 & ~n19746 ) ;
  assign n19995 = ~n6077 & n19994 ;
  assign n19996 = n8071 | n19995 ;
  assign n19997 = n19996 ^ n6981 ^ n5869 ;
  assign n19998 = n16791 & n19997 ;
  assign n19999 = ~n8809 & n19998 ;
  assign n20000 = n970 | n19999 ;
  assign n20001 = n19993 | n20000 ;
  assign n20002 = n7220 ^ n5850 ^ 1'b0 ;
  assign n20003 = n14558 ^ n1285 ^ 1'b0 ;
  assign n20004 = n20002 | n20003 ;
  assign n20005 = n17107 ^ n1387 ^ 1'b0 ;
  assign n20006 = n20005 ^ n1422 ^ 1'b0 ;
  assign n20007 = n20006 ^ n12656 ^ n12084 ;
  assign n20008 = n15882 ^ n3135 ^ 1'b0 ;
  assign n20009 = n4508 & ~n6533 ;
  assign n20010 = n11681 | n12447 ;
  assign n20011 = ~n20009 & n20010 ;
  assign n20013 = ( n3646 & n4229 ) | ( n3646 & ~n17502 ) | ( n4229 & ~n17502 ) ;
  assign n20012 = n11221 & ~n16405 ;
  assign n20014 = n20013 ^ n20012 ^ 1'b0 ;
  assign n20015 = n5518 & ~n6161 ;
  assign n20016 = n10065 | n20015 ;
  assign n20017 = ( n4086 & n16314 ) | ( n4086 & n20016 ) | ( n16314 & n20016 ) ;
  assign n20018 = n14102 & n20017 ;
  assign n20019 = ~n20014 & n20018 ;
  assign n20020 = n14027 ^ n8070 ^ 1'b0 ;
  assign n20021 = ( ~n1574 & n6450 ) | ( ~n1574 & n7970 ) | ( n6450 & n7970 ) ;
  assign n20022 = ~n19468 & n20021 ;
  assign n20023 = n8684 ^ n5345 ^ 1'b0 ;
  assign n20024 = n11876 & ~n20023 ;
  assign n20025 = n11906 ^ n9507 ^ 1'b0 ;
  assign n20026 = n10501 | n18422 ;
  assign n20027 = n8420 ^ n5049 ^ n2469 ;
  assign n20029 = n6433 ^ n1546 ^ 1'b0 ;
  assign n20028 = n6999 & ~n11392 ;
  assign n20030 = n20029 ^ n20028 ^ 1'b0 ;
  assign n20044 = ~n7802 & n19808 ;
  assign n20031 = n220 & ~n567 ;
  assign n20032 = ~n1267 & n20031 ;
  assign n20033 = n1010 & ~n12993 ;
  assign n20034 = n20033 ^ n179 ^ 1'b0 ;
  assign n20035 = n7568 ^ n6743 ^ 1'b0 ;
  assign n20036 = n305 & n13694 ;
  assign n20037 = n9925 & n20036 ;
  assign n20038 = n11209 ^ n6121 ^ n1679 ;
  assign n20039 = n14499 & ~n20038 ;
  assign n20040 = ~n20037 & n20039 ;
  assign n20041 = ~n20035 & n20040 ;
  assign n20042 = ( n11563 & n20034 ) | ( n11563 & n20041 ) | ( n20034 & n20041 ) ;
  assign n20043 = n20032 | n20042 ;
  assign n20045 = n20044 ^ n20043 ^ 1'b0 ;
  assign n20046 = n20045 ^ n16409 ^ 1'b0 ;
  assign n20047 = n16820 ^ n7042 ^ 1'b0 ;
  assign n20048 = n12563 ^ n7355 ^ 1'b0 ;
  assign n20049 = n20048 ^ n4945 ^ 1'b0 ;
  assign n20050 = ~n1003 & n20049 ;
  assign n20051 = n5606 | n20050 ;
  assign n20057 = n406 & ~n1014 ;
  assign n20058 = ~n406 & n20057 ;
  assign n20055 = n1752 & n3797 ;
  assign n20056 = ~n5872 & n20055 ;
  assign n20052 = n1258 & n4685 ;
  assign n20053 = ~n1258 & n20052 ;
  assign n20054 = n4982 & n20053 ;
  assign n20059 = n20058 ^ n20056 ^ n20054 ;
  assign n20060 = ~n4153 & n5368 ;
  assign n20061 = n774 | n2923 ;
  assign n20062 = n2179 | n3847 ;
  assign n20063 = n20062 ^ n9906 ^ 1'b0 ;
  assign n20064 = n20061 & n20063 ;
  assign n20065 = n13326 & n20064 ;
  assign n20067 = n14663 ^ n2943 ^ 1'b0 ;
  assign n20068 = n15869 & n20067 ;
  assign n20066 = n1093 | n9074 ;
  assign n20069 = n20068 ^ n20066 ^ 1'b0 ;
  assign n20070 = ~n4626 & n11604 ;
  assign n20071 = n13819 ^ n2852 ^ 1'b0 ;
  assign n20072 = n20071 ^ n1648 ^ 1'b0 ;
  assign n20073 = n11622 & ~n20072 ;
  assign n20074 = n3301 ^ n2799 ^ 1'b0 ;
  assign n20075 = n6533 & ~n20074 ;
  assign n20076 = ~n3011 & n11971 ;
  assign n20077 = n7702 & n20076 ;
  assign n20078 = n7164 ^ n3227 ^ 1'b0 ;
  assign n20079 = ~n4059 & n7556 ;
  assign n20080 = n908 & n20079 ;
  assign n20081 = n7311 | n20080 ;
  assign n20082 = n20081 ^ n19821 ^ 1'b0 ;
  assign n20083 = ( n6296 & n9929 ) | ( n6296 & n13583 ) | ( n9929 & n13583 ) ;
  assign n20084 = n15862 ^ n9057 ^ 1'b0 ;
  assign n20085 = ~n6857 & n8499 ;
  assign n20086 = ~n8499 & n20085 ;
  assign n20087 = n13018 & ~n20086 ;
  assign n20088 = n20086 & n20087 ;
  assign n20089 = n688 | n18074 ;
  assign n20090 = n16436 & ~n20089 ;
  assign n20091 = n16940 & ~n18405 ;
  assign n20092 = n20091 ^ n6215 ^ n5973 ;
  assign n20093 = n18522 ^ n4149 ^ 1'b0 ;
  assign n20094 = n20093 ^ n11222 ^ 1'b0 ;
  assign n20095 = n14184 | n20094 ;
  assign n20096 = n3531 | n5126 ;
  assign n20097 = n20095 & ~n20096 ;
  assign n20098 = n4735 & ~n13456 ;
  assign n20099 = n20098 ^ n2488 ^ 1'b0 ;
  assign n20100 = n8507 & n8635 ;
  assign n20101 = ~n4747 & n20100 ;
  assign n20102 = ( ~n1516 & n2605 ) | ( ~n1516 & n6945 ) | ( n2605 & n6945 ) ;
  assign n20103 = n4902 | n20102 ;
  assign n20104 = n20103 ^ n7713 ^ 1'b0 ;
  assign n20105 = n20101 & ~n20104 ;
  assign n20106 = n16407 & ~n20105 ;
  assign n20107 = n20106 ^ n15634 ^ 1'b0 ;
  assign n20108 = n18021 & n20107 ;
  assign n20109 = n11469 ^ n9057 ^ 1'b0 ;
  assign n20110 = n5840 | n20109 ;
  assign n20111 = n20110 ^ n7589 ^ 1'b0 ;
  assign n20112 = n11327 & ~n20111 ;
  assign n20113 = n9858 ^ n4862 ^ 1'b0 ;
  assign n20114 = n20113 ^ n20030 ^ n944 ;
  assign n20115 = n17172 ^ n14254 ^ 1'b0 ;
  assign n20116 = n7601 & ~n20115 ;
  assign n20117 = n162 & n668 ;
  assign n20118 = n7718 ^ n6397 ^ 1'b0 ;
  assign n20119 = n2513 | n20118 ;
  assign n20120 = ~n18292 & n20119 ;
  assign n20121 = n7627 ^ n2821 ^ 1'b0 ;
  assign n20122 = n8880 | n20121 ;
  assign n20123 = n10946 ^ n6672 ^ 1'b0 ;
  assign n20124 = n881 | n15596 ;
  assign n20125 = n4529 & ~n20124 ;
  assign n20127 = n17428 ^ n2317 ^ n1657 ;
  assign n20126 = n11880 | n16400 ;
  assign n20128 = n20127 ^ n20126 ^ 1'b0 ;
  assign n20129 = ~n8332 & n20128 ;
  assign n20130 = n20129 ^ n18301 ^ 1'b0 ;
  assign n20131 = n20125 & n20130 ;
  assign n20135 = n7830 & n11850 ;
  assign n20136 = n20135 ^ n1726 ^ 1'b0 ;
  assign n20132 = n11850 ^ n1119 ^ 1'b0 ;
  assign n20133 = ~n19933 & n20132 ;
  assign n20134 = ~n16650 & n20133 ;
  assign n20137 = n20136 ^ n20134 ^ 1'b0 ;
  assign n20138 = n13196 ^ n2912 ^ 1'b0 ;
  assign n20139 = ( n905 & n996 ) | ( n905 & ~n5256 ) | ( n996 & ~n5256 ) ;
  assign n20140 = n372 & n7568 ;
  assign n20141 = n9098 ^ n7314 ^ 1'b0 ;
  assign n20142 = n16221 ^ n14901 ^ 1'b0 ;
  assign n20147 = n5936 | n6461 ;
  assign n20144 = n2316 | n4925 ;
  assign n20145 = n6941 & ~n20144 ;
  assign n20143 = n7263 ^ n6910 ^ 1'b0 ;
  assign n20146 = n20145 ^ n20143 ^ n6291 ;
  assign n20148 = n20147 ^ n20146 ^ n8539 ;
  assign n20149 = ~n312 & n2268 ;
  assign n20150 = n20149 ^ n11517 ^ n2452 ;
  assign n20151 = n11458 ^ n5375 ^ 1'b0 ;
  assign n20152 = n306 & ~n6818 ;
  assign n20153 = ~n16782 & n20152 ;
  assign n20154 = n5741 & ~n20153 ;
  assign n20155 = n17183 ^ n10199 ^ n2061 ;
  assign n20157 = n4141 & ~n7830 ;
  assign n20158 = ( ~n1883 & n13458 ) | ( ~n1883 & n20157 ) | ( n13458 & n20157 ) ;
  assign n20156 = ~n7131 & n8239 ;
  assign n20159 = n20158 ^ n20156 ^ 1'b0 ;
  assign n20160 = ~n5514 & n12726 ;
  assign n20161 = n20159 & n20160 ;
  assign n20162 = n19118 | n20161 ;
  assign n20167 = n152 & ~n7983 ;
  assign n20168 = n6680 & n20167 ;
  assign n20169 = n20168 ^ n7601 ^ n6813 ;
  assign n20164 = n5329 | n6442 ;
  assign n20165 = n2120 | n20164 ;
  assign n20163 = ( n2980 & ~n6172 ) | ( n2980 & n12789 ) | ( ~n6172 & n12789 ) ;
  assign n20166 = n20165 ^ n20163 ^ 1'b0 ;
  assign n20170 = n20169 ^ n20166 ^ 1'b0 ;
  assign n20171 = n10488 & n20170 ;
  assign n20172 = n8679 & n12059 ;
  assign n20173 = n7080 | n9704 ;
  assign n20174 = n4390 & ~n20173 ;
  assign n20175 = n20174 ^ n11797 ^ 1'b0 ;
  assign n20176 = n17583 ^ n2732 ^ 1'b0 ;
  assign n20177 = ~n1701 & n6940 ;
  assign n20184 = n14863 ^ n7627 ^ n5401 ;
  assign n20178 = n1673 ^ n58 ^ 1'b0 ;
  assign n20179 = n5323 & n20178 ;
  assign n20180 = n5236 & n20179 ;
  assign n20181 = ~n5236 & n20180 ;
  assign n20182 = ~n8254 & n20181 ;
  assign n20183 = n20182 ^ n15018 ^ 1'b0 ;
  assign n20185 = n20184 ^ n20183 ^ n9889 ;
  assign n20186 = ~n1413 & n11527 ;
  assign n20187 = ~n9733 & n20186 ;
  assign n20188 = n20187 ^ n4964 ^ 1'b0 ;
  assign n20189 = n2330 & ~n20188 ;
  assign n20190 = n105 | n15995 ;
  assign n20191 = n11271 & ~n20190 ;
  assign n20192 = n20191 ^ n16004 ^ n9426 ;
  assign n20193 = n20192 ^ n655 ^ 1'b0 ;
  assign n20194 = n40 | n15007 ;
  assign n20195 = n20194 ^ n7746 ^ 1'b0 ;
  assign n20196 = n14696 & ~n20195 ;
  assign n20197 = n20196 ^ n18869 ^ 1'b0 ;
  assign n20198 = ~n9133 & n20197 ;
  assign n20199 = n7904 ^ n5860 ^ 1'b0 ;
  assign n20200 = n20199 ^ n1114 ^ 1'b0 ;
  assign n20201 = n5268 & ~n20200 ;
  assign n20202 = n20201 ^ n862 ^ 1'b0 ;
  assign n20203 = n13801 & n20202 ;
  assign n20204 = ~n1830 & n20203 ;
  assign n20205 = n15724 & n20101 ;
  assign n20206 = x0 & n9150 ;
  assign n20207 = n20206 ^ n3227 ^ 1'b0 ;
  assign n20208 = n20207 ^ n18062 ^ n1821 ;
  assign n20209 = n6437 & n20208 ;
  assign n20215 = ~n311 & n5054 ;
  assign n20216 = ~n2222 & n20215 ;
  assign n20217 = n819 & ~n4935 ;
  assign n20218 = n20216 & n20217 ;
  assign n20213 = n961 | n10076 ;
  assign n20214 = n5010 | n20213 ;
  assign n20219 = n20218 ^ n20214 ^ 1'b0 ;
  assign n20210 = n13845 & n16448 ;
  assign n20211 = n20210 ^ n11680 ^ 1'b0 ;
  assign n20212 = n17741 | n20211 ;
  assign n20220 = n20219 ^ n20212 ^ 1'b0 ;
  assign n20221 = n592 | n10624 ;
  assign n20222 = ~n1469 & n15527 ;
  assign n20223 = ~n10910 & n15594 ;
  assign n20224 = ~n13031 & n20223 ;
  assign n20225 = n20224 ^ n1099 ^ 1'b0 ;
  assign n20226 = n14823 ^ n12943 ^ 1'b0 ;
  assign n20227 = n1066 | n20226 ;
  assign n20228 = n6576 | n20227 ;
  assign n20229 = ~n11202 & n14387 ;
  assign n20232 = ~n14200 & n15330 ;
  assign n20231 = n600 | n1958 ;
  assign n20233 = n20232 ^ n20231 ^ 1'b0 ;
  assign n20230 = n11855 ^ n1838 ^ 1'b0 ;
  assign n20234 = n20233 ^ n20230 ^ 1'b0 ;
  assign n20235 = n13028 & ~n13702 ;
  assign n20236 = n10392 & n20235 ;
  assign n20237 = n2275 & ~n20236 ;
  assign n20238 = n4624 & n17883 ;
  assign n20239 = n20238 ^ n8397 ^ 1'b0 ;
  assign n20240 = n8976 ^ n4631 ^ 1'b0 ;
  assign n20241 = ~n10711 & n14131 ;
  assign n20242 = n4802 & n7303 ;
  assign n20243 = n58 & n2303 ;
  assign n20244 = ~n1349 & n20243 ;
  assign n20245 = n20242 & n20244 ;
  assign n20246 = n20241 | n20245 ;
  assign n20247 = n20240 & ~n20246 ;
  assign n20248 = n16548 ^ n5747 ^ 1'b0 ;
  assign n20249 = n3030 & ~n20248 ;
  assign n20250 = n5438 & ~n7655 ;
  assign n20251 = ( n6293 & n11613 ) | ( n6293 & n20250 ) | ( n11613 & n20250 ) ;
  assign n20252 = n17075 & ~n20251 ;
  assign n20253 = n3264 ^ n371 ^ 1'b0 ;
  assign n20254 = n2998 & ~n20253 ;
  assign n20255 = n20254 ^ n9284 ^ 1'b0 ;
  assign n20256 = ~n4188 & n4903 ;
  assign n20257 = n20256 ^ n4170 ^ 1'b0 ;
  assign n20258 = n13507 & ~n20257 ;
  assign n20259 = n774 & ~n16673 ;
  assign n20260 = n7614 & ~n9707 ;
  assign n20261 = n19409 ^ n188 ^ 1'b0 ;
  assign n20262 = ~n20260 & n20261 ;
  assign n20263 = ~n3970 & n20262 ;
  assign n20264 = n3628 & n7906 ;
  assign n20265 = n20264 ^ n9050 ^ 1'b0 ;
  assign n20266 = ~n16597 & n20265 ;
  assign n20267 = n6273 | n11035 ;
  assign n20268 = n1271 & ~n20267 ;
  assign n20269 = n20266 & ~n20268 ;
  assign n20270 = n20269 ^ n16285 ^ 1'b0 ;
  assign n20271 = n11141 & n18276 ;
  assign n20272 = n8064 ^ n2420 ^ n1941 ;
  assign n20273 = n5067 & n20272 ;
  assign n20274 = n20273 ^ n7238 ^ 1'b0 ;
  assign n20275 = n4252 & n9832 ;
  assign n20276 = n20274 & n20275 ;
  assign n20277 = n14853 ^ n2163 ^ 1'b0 ;
  assign n20278 = n19685 ^ n12578 ^ 1'b0 ;
  assign n20279 = n7493 ^ n1802 ^ 1'b0 ;
  assign n20280 = n20279 ^ n19980 ^ 1'b0 ;
  assign n20281 = n16066 ^ n77 ^ 1'b0 ;
  assign n20282 = ( n919 & n10484 ) | ( n919 & n20281 ) | ( n10484 & n20281 ) ;
  assign n20283 = n5851 & ~n16018 ;
  assign n20284 = n1050 & ~n1437 ;
  assign n20285 = n20284 ^ n5377 ^ 1'b0 ;
  assign n20286 = n4208 & n13026 ;
  assign n20287 = ( ~n12704 & n20285 ) | ( ~n12704 & n20286 ) | ( n20285 & n20286 ) ;
  assign n20288 = n11457 & ~n18746 ;
  assign n20289 = n3062 & n7643 ;
  assign n20290 = n9825 ^ n6165 ^ 1'b0 ;
  assign n20291 = n20290 ^ n205 ^ 1'b0 ;
  assign n20292 = n7816 & n16975 ;
  assign n20293 = n3558 & n18209 ;
  assign n20294 = n20293 ^ n9795 ^ 1'b0 ;
  assign n20295 = n10882 & ~n12842 ;
  assign n20296 = n4773 | n9035 ;
  assign n20297 = ( ~n2883 & n7558 ) | ( ~n2883 & n11817 ) | ( n7558 & n11817 ) ;
  assign n20298 = n13832 ^ n9232 ^ 1'b0 ;
  assign n20299 = n20298 ^ n17100 ^ n13176 ;
  assign n20300 = n2120 | n5456 ;
  assign n20301 = n20300 ^ n13881 ^ 1'b0 ;
  assign n20302 = n13513 ^ n9946 ^ n5775 ;
  assign n20303 = n20302 ^ n5781 ^ 1'b0 ;
  assign n20304 = n15358 ^ n2444 ^ 1'b0 ;
  assign n20305 = n7447 & n20304 ;
  assign n20306 = n20305 ^ n1029 ^ 1'b0 ;
  assign n20307 = n20303 & ~n20306 ;
  assign n20308 = ( n5946 & n6473 ) | ( n5946 & n14904 ) | ( n6473 & n14904 ) ;
  assign n20309 = n10470 ^ n25 ^ 1'b0 ;
  assign n20310 = n8307 ^ n2796 ^ n805 ;
  assign n20311 = n612 & n20310 ;
  assign n20312 = ~n1167 & n8324 ;
  assign n20313 = n5750 & n7666 ;
  assign n20314 = n687 & ~n12282 ;
  assign n20315 = n20314 ^ n5461 ^ 1'b0 ;
  assign n20316 = n20313 & ~n20315 ;
  assign n20317 = ~n20312 & n20316 ;
  assign n20318 = ~n1700 & n9092 ;
  assign n20319 = n9449 ^ n1535 ^ 1'b0 ;
  assign n20320 = n20319 ^ n17604 ^ n2656 ;
  assign n20321 = n6951 ^ n3480 ^ 1'b0 ;
  assign n20322 = n2845 & n20321 ;
  assign n20323 = ~n4481 & n20322 ;
  assign n20324 = n1181 | n13438 ;
  assign n20325 = n20324 ^ n5021 ^ 1'b0 ;
  assign n20326 = ( n6870 & n19421 ) | ( n6870 & n20325 ) | ( n19421 & n20325 ) ;
  assign n20327 = n9416 & n20326 ;
  assign n20328 = n19602 ^ n18032 ^ 1'b0 ;
  assign n20329 = n11258 ^ n755 ^ 1'b0 ;
  assign n20331 = n365 & ~n856 ;
  assign n20332 = ~n2472 & n20331 ;
  assign n20330 = n3809 & n6998 ;
  assign n20333 = n20332 ^ n20330 ^ n3512 ;
  assign n20334 = n11913 | n20333 ;
  assign n20335 = n20334 ^ n6620 ^ 1'b0 ;
  assign n20336 = n7695 | n8327 ;
  assign n20338 = n5575 | n6569 ;
  assign n20339 = n20338 ^ n6681 ^ 1'b0 ;
  assign n20340 = ~n417 & n20339 ;
  assign n20337 = n302 & ~n5336 ;
  assign n20341 = n20340 ^ n20337 ^ n18462 ;
  assign n20342 = n5956 | n12187 ;
  assign n20343 = n302 & ~n15653 ;
  assign n20344 = n20343 ^ n2034 ^ 1'b0 ;
  assign n20345 = n20344 ^ n823 ^ 1'b0 ;
  assign n20346 = ~n3901 & n5444 ;
  assign n20347 = n10193 ^ n6590 ^ 1'b0 ;
  assign n20348 = n20093 ^ n1697 ^ 1'b0 ;
  assign n20349 = ~n6387 & n20348 ;
  assign n20350 = n20349 ^ n1778 ^ 1'b0 ;
  assign n20351 = n20350 ^ n5755 ^ 1'b0 ;
  assign n20352 = ( ~n1379 & n8321 ) | ( ~n1379 & n17784 ) | ( n8321 & n17784 ) ;
  assign n20353 = n11174 & ~n11834 ;
  assign n20354 = n20353 ^ n13189 ^ 1'b0 ;
  assign n20355 = ( n10738 & n20352 ) | ( n10738 & n20354 ) | ( n20352 & n20354 ) ;
  assign n20356 = n3050 | n20355 ;
  assign n20357 = n10917 | n20356 ;
  assign n20358 = n4977 & n7164 ;
  assign n20359 = n20358 ^ n15325 ^ 1'b0 ;
  assign n20360 = n5027 | n20359 ;
  assign n20361 = n20360 ^ n10736 ^ 1'b0 ;
  assign n20362 = n20361 ^ n3939 ^ 1'b0 ;
  assign n20363 = n18414 & ~n20362 ;
  assign n20364 = n7273 ^ n1546 ^ 1'b0 ;
  assign n20365 = n6756 & ~n20364 ;
  assign n20366 = n12649 & n20365 ;
  assign n20367 = n8062 ^ n737 ^ 1'b0 ;
  assign n20368 = ( n2218 & ~n18439 ) | ( n2218 & n20367 ) | ( ~n18439 & n20367 ) ;
  assign n20369 = n3335 & ~n9670 ;
  assign n20370 = ~n5747 & n20369 ;
  assign n20371 = n1745 & ~n8043 ;
  assign n20372 = n14134 & n20371 ;
  assign n20373 = ( n6028 & ~n20370 ) | ( n6028 & n20372 ) | ( ~n20370 & n20372 ) ;
  assign n20374 = n1655 & ~n5755 ;
  assign n20375 = n4369 ^ n83 ^ 1'b0 ;
  assign n20376 = n20374 | n20375 ;
  assign n20377 = n12990 ^ n2872 ^ 1'b0 ;
  assign n20378 = n11934 & ~n20377 ;
  assign n20379 = n7964 ^ n4824 ^ 1'b0 ;
  assign n20380 = n3933 & ~n17636 ;
  assign n20381 = n8328 ^ x6 ^ 1'b0 ;
  assign n20382 = n11477 & n20381 ;
  assign n20384 = n18799 ^ n3560 ^ 1'b0 ;
  assign n20385 = n3548 & n20384 ;
  assign n20383 = n13596 ^ n12693 ^ 1'b0 ;
  assign n20386 = n20385 ^ n20383 ^ n1422 ;
  assign n20387 = ~n6982 & n19989 ;
  assign n20388 = n20387 ^ n15171 ^ 1'b0 ;
  assign n20389 = n7933 ^ n7602 ^ 1'b0 ;
  assign n20390 = n15643 & ~n20389 ;
  assign n20391 = n5811 ^ n382 ^ 1'b0 ;
  assign n20392 = ( n4991 & n6817 ) | ( n4991 & ~n13721 ) | ( n6817 & ~n13721 ) ;
  assign n20393 = ~n1449 & n1839 ;
  assign n20394 = n20392 & ~n20393 ;
  assign n20395 = n8084 ^ n6535 ^ 1'b0 ;
  assign n20400 = n12565 ^ n10168 ^ n9312 ;
  assign n20396 = n16406 ^ n16165 ^ 1'b0 ;
  assign n20397 = ~n1466 & n20396 ;
  assign n20398 = n4036 & ~n10934 ;
  assign n20399 = ~n20397 & n20398 ;
  assign n20401 = n20400 ^ n20399 ^ 1'b0 ;
  assign n20402 = n12158 ^ n11981 ^ 1'b0 ;
  assign n20403 = n9972 & ~n20402 ;
  assign n20404 = n5383 ^ n1653 ^ 1'b0 ;
  assign n20405 = n1377 | n20404 ;
  assign n20406 = ( ~n777 & n20403 ) | ( ~n777 & n20405 ) | ( n20403 & n20405 ) ;
  assign n20407 = n5273 & ~n6393 ;
  assign n20408 = n5425 | n11483 ;
  assign n20409 = n16926 & n20408 ;
  assign n20410 = n20409 ^ n5836 ^ 1'b0 ;
  assign n20411 = n20410 ^ n8869 ^ n7162 ;
  assign n20412 = n1853 & ~n2152 ;
  assign n20413 = ~n5380 & n13969 ;
  assign n20414 = n20413 ^ n7475 ^ 1'b0 ;
  assign n20415 = n13521 & n19832 ;
  assign n20416 = n15491 ^ n7480 ^ 1'b0 ;
  assign n20417 = n667 & ~n20416 ;
  assign n20418 = n6774 & ~n14778 ;
  assign n20419 = n11140 | n12049 ;
  assign n20420 = n20419 ^ n6248 ^ 1'b0 ;
  assign n20421 = ~n9865 & n20420 ;
  assign n20422 = n20421 ^ n18900 ^ 1'b0 ;
  assign n20423 = n2660 | n9323 ;
  assign n20424 = n409 & ~n2002 ;
  assign n20425 = n20424 ^ n1841 ^ 1'b0 ;
  assign n20426 = n20423 | n20425 ;
  assign n20427 = n13573 ^ n5194 ^ 1'b0 ;
  assign n20428 = ~n11602 & n20427 ;
  assign n20429 = n1056 & n11703 ;
  assign n20430 = ( n631 & ~n14111 ) | ( n631 & n20429 ) | ( ~n14111 & n20429 ) ;
  assign n20431 = n7451 & n9447 ;
  assign n20432 = n11999 & n20431 ;
  assign n20433 = ~n961 & n20432 ;
  assign n20434 = n20433 ^ n19667 ^ 1'b0 ;
  assign n20435 = n20430 & ~n20434 ;
  assign n20436 = n13561 | n13990 ;
  assign n20437 = n20436 ^ n9803 ^ 1'b0 ;
  assign n20438 = n18244 ^ n625 ^ 1'b0 ;
  assign n20439 = n6498 ^ n782 ^ 1'b0 ;
  assign n20440 = n12839 & n20439 ;
  assign n20441 = n20440 ^ n19331 ^ n3226 ;
  assign n20442 = n10359 ^ n9534 ^ 1'b0 ;
  assign n20443 = ~n5285 & n20442 ;
  assign n20444 = n20443 ^ n3040 ^ 1'b0 ;
  assign n20445 = n20405 ^ n1590 ^ 1'b0 ;
  assign n20446 = n2961 | n6472 ;
  assign n20447 = n20446 ^ n5787 ^ 1'b0 ;
  assign n20448 = n1376 | n20447 ;
  assign n20449 = n1157 & ~n19982 ;
  assign n20450 = n20449 ^ n10686 ^ 1'b0 ;
  assign n20451 = n20450 ^ n16777 ^ 1'b0 ;
  assign n20452 = ~n796 & n2796 ;
  assign n20453 = n5561 ^ n5201 ^ 1'b0 ;
  assign n20454 = ~n7958 & n10090 ;
  assign n20456 = n1249 | n2473 ;
  assign n20457 = n1538 & ~n20456 ;
  assign n20458 = n2053 & ~n20457 ;
  assign n20459 = n9124 | n20458 ;
  assign n20460 = n20459 ^ n6274 ^ 1'b0 ;
  assign n20455 = n6095 & ~n6641 ;
  assign n20461 = n20460 ^ n20455 ^ 1'b0 ;
  assign n20462 = ~n18333 & n20461 ;
  assign n20463 = ~n12967 & n16490 ;
  assign n20464 = n9112 ^ n4381 ^ 1'b0 ;
  assign n20465 = n16712 | n20464 ;
  assign n20466 = n2432 & ~n17939 ;
  assign n20467 = ~n7080 & n20466 ;
  assign n20468 = ~n275 & n20467 ;
  assign n20469 = n16747 & n20468 ;
  assign n20470 = n15034 ^ n10423 ^ 1'b0 ;
  assign n20471 = n5176 & n20470 ;
  assign n20472 = n17873 ^ n10962 ^ 1'b0 ;
  assign n20473 = n20471 & n20472 ;
  assign n20474 = n20469 & n20473 ;
  assign n20475 = n10443 & ~n17027 ;
  assign n20476 = n2208 & ~n11790 ;
  assign n20477 = ~n2616 & n10092 ;
  assign n20478 = n16167 ^ n2048 ^ 1'b0 ;
  assign n20479 = ~n20477 & n20478 ;
  assign n20480 = n14768 ^ n13826 ^ 1'b0 ;
  assign n20481 = ~n11360 & n20480 ;
  assign n20482 = n1745 ^ n1647 ^ 1'b0 ;
  assign n20483 = n2353 & ~n20482 ;
  assign n20484 = n654 & n19999 ;
  assign n20485 = n6100 ^ n1705 ^ 1'b0 ;
  assign n20486 = n2246 ^ n944 ^ 1'b0 ;
  assign n20487 = n6723 | n20486 ;
  assign n20488 = n10638 ^ n5412 ^ 1'b0 ;
  assign n20489 = n20488 ^ n1837 ^ n60 ;
  assign n20490 = n20489 ^ n13155 ^ 1'b0 ;
  assign n20491 = ~n20487 & n20490 ;
  assign n20492 = n6258 ^ n2486 ^ n192 ;
  assign n20493 = n4711 & n10099 ;
  assign n20494 = ~n20492 & n20493 ;
  assign n20495 = n11386 & ~n12695 ;
  assign n20496 = n6568 & n20495 ;
  assign n20497 = n7369 | n20496 ;
  assign n20498 = n1845 | n20497 ;
  assign n20499 = ~n10618 & n20498 ;
  assign n20500 = n20499 ^ n9110 ^ n8728 ;
  assign n20501 = n2443 ^ n1414 ^ 1'b0 ;
  assign n20502 = n48 & ~n2498 ;
  assign n20503 = n2498 & n20502 ;
  assign n20504 = n5654 ^ n3643 ^ 1'b0 ;
  assign n20505 = n91 | n4543 ;
  assign n20506 = n1867 | n20505 ;
  assign n20507 = n8483 & n20506 ;
  assign n20508 = n8043 ^ n6083 ^ 1'b0 ;
  assign n20509 = n3738 | n20508 ;
  assign n20510 = n20509 ^ n18095 ^ n12873 ;
  assign n20511 = n10438 ^ n1884 ^ 1'b0 ;
  assign n20512 = n2387 & n20511 ;
  assign n20513 = n16252 ^ n9716 ^ 1'b0 ;
  assign n20514 = n20512 & n20513 ;
  assign n20515 = n20514 ^ n18528 ^ 1'b0 ;
  assign n20516 = n61 & ~n20515 ;
  assign n20518 = n983 & ~n3032 ;
  assign n20519 = n14736 | n20518 ;
  assign n20520 = n20519 ^ n12550 ^ 1'b0 ;
  assign n20517 = n7452 ^ n2657 ^ 1'b0 ;
  assign n20521 = n20520 ^ n20517 ^ 1'b0 ;
  assign n20522 = ( n417 & n1742 ) | ( n417 & n7187 ) | ( n1742 & n7187 ) ;
  assign n20523 = ~n5438 & n20522 ;
  assign n20524 = ~n20521 & n20523 ;
  assign n20525 = n694 | n3335 ;
  assign n20526 = n10726 & n20525 ;
  assign n20527 = n2317 | n14884 ;
  assign n20528 = n7554 ^ n1307 ^ 1'b0 ;
  assign n20529 = n1035 ^ n288 ^ 1'b0 ;
  assign n20530 = n1981 & ~n20529 ;
  assign n20531 = n20530 ^ n9725 ^ 1'b0 ;
  assign n20532 = n11447 ^ n5303 ^ 1'b0 ;
  assign n20533 = n19312 & ~n20532 ;
  assign n20534 = n910 & n2199 ;
  assign n20535 = n20534 ^ n11685 ^ 1'b0 ;
  assign n20536 = n13167 | n20535 ;
  assign n20537 = n20533 | n20536 ;
  assign n20539 = n1546 | n6185 ;
  assign n20538 = n2363 | n10424 ;
  assign n20540 = n20539 ^ n20538 ^ 1'b0 ;
  assign n20541 = n16651 ^ n1546 ^ 1'b0 ;
  assign n20542 = n20540 | n20541 ;
  assign n20543 = ~n10445 & n18735 ;
  assign n20547 = n3042 ^ n2856 ^ 1'b0 ;
  assign n20544 = n1601 & n3962 ;
  assign n20545 = n20544 ^ n13200 ^ 1'b0 ;
  assign n20546 = n20545 ^ n6330 ^ n448 ;
  assign n20548 = n20547 ^ n20546 ^ 1'b0 ;
  assign n20549 = n12740 & ~n14810 ;
  assign n20550 = n8898 & n20549 ;
  assign n20551 = n7544 & ~n19889 ;
  assign n20552 = n20550 & n20551 ;
  assign n20553 = ~n2270 & n9248 ;
  assign n20554 = n11850 & ~n13706 ;
  assign n20555 = n16353 & n20554 ;
  assign n20556 = n20555 ^ n10852 ^ 1'b0 ;
  assign n20557 = n20556 ^ n20017 ^ n4914 ;
  assign n20558 = n11789 & ~n20545 ;
  assign n20559 = n2877 ^ n1083 ^ 1'b0 ;
  assign n20560 = n7170 & n10257 ;
  assign n20561 = n20559 & n20560 ;
  assign n20562 = n4164 & ~n20561 ;
  assign n20563 = n1590 & n2020 ;
  assign n20564 = n11512 & ~n20203 ;
  assign n20565 = n2537 & ~n5480 ;
  assign n20566 = ~n89 & n20565 ;
  assign n20567 = n12603 ^ n7132 ^ 1'b0 ;
  assign n20568 = n1451 & n19524 ;
  assign n20569 = ~n20567 & n20568 ;
  assign n20570 = n5893 & n6429 ;
  assign n20571 = n8553 ^ n7782 ^ n6832 ;
  assign n20572 = n20571 ^ n15867 ^ n6003 ;
  assign n20573 = n10330 ^ n931 ^ 1'b0 ;
  assign n20574 = ~n2161 & n20573 ;
  assign n20575 = n4914 & ~n9212 ;
  assign n20576 = n20574 & n20575 ;
  assign n20577 = ~n5231 & n8497 ;
  assign n20578 = n9378 & n12390 ;
  assign n20579 = ~n20577 & n20578 ;
  assign n20580 = n15234 | n20579 ;
  assign n20581 = ~n2146 & n4088 ;
  assign n20582 = n2820 & n20581 ;
  assign n20584 = ~n11209 & n18179 ;
  assign n20583 = n1018 | n3979 ;
  assign n20585 = n20584 ^ n20583 ^ 1'b0 ;
  assign n20586 = n20573 & n20585 ;
  assign n20587 = n20586 ^ n316 ^ 1'b0 ;
  assign n20588 = n3434 & ~n15238 ;
  assign n20589 = n1948 | n2828 ;
  assign n20590 = n15748 | n20589 ;
  assign n20591 = n13685 & ~n14871 ;
  assign n20592 = n2492 & n3933 ;
  assign n20593 = n125 | n4685 ;
  assign n20594 = n798 | n20593 ;
  assign n20595 = n15177 ^ n14256 ^ n738 ;
  assign n20596 = ~n13614 & n15404 ;
  assign n20597 = n14611 ^ n11109 ^ 1'b0 ;
  assign n20598 = ~n2179 & n6281 ;
  assign n20599 = n10354 ^ n7266 ^ 1'b0 ;
  assign n20600 = n20598 & n20599 ;
  assign n20601 = n20600 ^ n11414 ^ 1'b0 ;
  assign n20602 = ~n2547 & n20601 ;
  assign n20603 = n19222 ^ n3928 ^ 1'b0 ;
  assign n20604 = ~n983 & n3924 ;
  assign n20605 = n20604 ^ n5626 ^ 1'b0 ;
  assign n20610 = n5607 ^ n1413 ^ 1'b0 ;
  assign n20611 = n19627 & n20610 ;
  assign n20606 = n2765 & ~n6794 ;
  assign n20607 = n20606 ^ n5902 ^ n5128 ;
  assign n20608 = n5145 & ~n20607 ;
  assign n20609 = n17834 & ~n20608 ;
  assign n20612 = n20611 ^ n20609 ^ 1'b0 ;
  assign n20613 = n6844 | n13257 ;
  assign n20614 = n8411 & ~n14378 ;
  assign n20615 = ~n3039 & n13375 ;
  assign n20616 = n4005 ^ n2873 ^ 1'b0 ;
  assign n20617 = n20616 ^ n1804 ^ 1'b0 ;
  assign n20618 = n1182 & ~n20617 ;
  assign n20619 = n2978 & n20618 ;
  assign n20620 = n11256 ^ n4832 ^ 1'b0 ;
  assign n20621 = ( n6749 & n20619 ) | ( n6749 & ~n20620 ) | ( n20619 & ~n20620 ) ;
  assign n20622 = n6630 | n17181 ;
  assign n20623 = n559 | n20622 ;
  assign n20624 = n7413 & ~n9905 ;
  assign n20625 = n20624 ^ n6012 ^ 1'b0 ;
  assign n20626 = n447 & n20625 ;
  assign n20627 = n20626 ^ n7051 ^ 1'b0 ;
  assign n20628 = ( n810 & n5058 ) | ( n810 & n7655 ) | ( n5058 & n7655 ) ;
  assign n20629 = n5733 & ~n20370 ;
  assign n20630 = ~n20628 & n20629 ;
  assign n20631 = ( n2427 & n10728 ) | ( n2427 & ~n15492 ) | ( n10728 & ~n15492 ) ;
  assign n20632 = n1323 | n20631 ;
  assign n20634 = n4725 | n4937 ;
  assign n20633 = n3661 & n18405 ;
  assign n20635 = n20634 ^ n20633 ^ 1'b0 ;
  assign n20636 = ( n4519 & n5368 ) | ( n4519 & n5524 ) | ( n5368 & n5524 ) ;
  assign n20637 = n20636 ^ n17622 ^ n14038 ;
  assign n20638 = n14875 & n15768 ;
  assign n20639 = n5306 ^ n3572 ^ 1'b0 ;
  assign n20640 = n2840 & ~n11742 ;
  assign n20641 = n347 & ~n11234 ;
  assign n20642 = n8393 & n11313 ;
  assign n20643 = n1069 & ~n20642 ;
  assign n20644 = n7342 ^ n6283 ^ 1'b0 ;
  assign n20645 = ~n5759 & n10665 ;
  assign n20646 = ~n1769 & n20645 ;
  assign n20647 = ~n20644 & n20646 ;
  assign n20648 = n5039 | n7296 ;
  assign n20649 = n20648 ^ n5444 ^ n2030 ;
  assign n20650 = n3314 & n12562 ;
  assign n20651 = n20650 ^ n5823 ^ 1'b0 ;
  assign n20652 = ~n2154 & n20651 ;
  assign n20653 = ~n20649 & n20652 ;
  assign n20654 = n6646 & n9209 ;
  assign n20655 = n8482 & ~n20654 ;
  assign n20656 = n13612 | n17166 ;
  assign n20657 = n20656 ^ n10872 ^ 1'b0 ;
  assign n20658 = n20657 ^ n8643 ^ n2661 ;
  assign n20661 = ~n1223 & n7997 ;
  assign n20662 = ~n5850 & n20661 ;
  assign n20663 = ~n3325 & n6082 ;
  assign n20664 = ~n1293 & n20663 ;
  assign n20665 = n20662 & n20664 ;
  assign n20666 = n3030 & ~n20665 ;
  assign n20667 = n15137 & ~n20666 ;
  assign n20659 = n8258 | n9680 ;
  assign n20660 = n6331 | n20659 ;
  assign n20668 = n20667 ^ n20660 ^ 1'b0 ;
  assign n20669 = n20668 ^ n11233 ^ 1'b0 ;
  assign n20670 = n17162 ^ n12773 ^ n6550 ;
  assign n20671 = ~n20669 & n20670 ;
  assign n20672 = ~n6722 & n9372 ;
  assign n20673 = n12622 ^ n1428 ^ 1'b0 ;
  assign n20674 = ~n12045 & n12145 ;
  assign n20675 = n13449 ^ n12239 ^ 1'b0 ;
  assign n20676 = n5449 ^ n2864 ^ 1'b0 ;
  assign n20677 = n7919 ^ n7556 ^ 1'b0 ;
  assign n20678 = n3198 & ~n20677 ;
  assign n20679 = n20678 ^ n13934 ^ 1'b0 ;
  assign n20680 = n417 & n8083 ;
  assign n20681 = ~n13320 & n20680 ;
  assign n20682 = n20681 ^ n4660 ^ 1'b0 ;
  assign n20685 = n4440 & n10164 ;
  assign n20683 = n3070 & ~n3937 ;
  assign n20684 = n20683 ^ n13251 ^ 1'b0 ;
  assign n20686 = n20685 ^ n20684 ^ 1'b0 ;
  assign n20687 = n15460 ^ n5117 ^ 1'b0 ;
  assign n20688 = n7132 & n7686 ;
  assign n20689 = n3867 & n20688 ;
  assign n20690 = n6291 & n12327 ;
  assign n20691 = n10652 ^ n3748 ^ 1'b0 ;
  assign n20692 = ~n2623 & n20691 ;
  assign n20693 = n20690 & n20692 ;
  assign n20694 = n20693 ^ n17632 ^ 1'b0 ;
  assign n20695 = ~n20689 & n20694 ;
  assign n20696 = ~n1539 & n10749 ;
  assign n20697 = n20696 ^ n4370 ^ 1'b0 ;
  assign n20698 = n10737 & ~n20697 ;
  assign n20699 = n20698 ^ n12996 ^ 1'b0 ;
  assign n20700 = n1029 ^ n448 ^ 1'b0 ;
  assign n20703 = n10118 ^ n6808 ^ 1'b0 ;
  assign n20704 = n2432 & ~n20703 ;
  assign n20701 = ~n578 & n5167 ;
  assign n20702 = n12173 & n20701 ;
  assign n20705 = n20704 ^ n20702 ^ 1'b0 ;
  assign n20706 = n20700 & ~n20705 ;
  assign n20707 = n17615 ^ n514 ^ 1'b0 ;
  assign n20708 = n870 | n3412 ;
  assign n20709 = n5073 & ~n20708 ;
  assign n20710 = n20709 ^ n15513 ^ 1'b0 ;
  assign n20711 = n20707 | n20710 ;
  assign n20712 = n17717 | n20711 ;
  assign n20713 = n17779 & ~n20712 ;
  assign n20714 = n18255 ^ n1738 ^ n609 ;
  assign n20715 = n10021 ^ n510 ^ 1'b0 ;
  assign n20716 = n694 & n20715 ;
  assign n20717 = ~n11312 & n20716 ;
  assign n20718 = n20717 ^ n5236 ^ 1'b0 ;
  assign n20719 = n2799 & ~n16478 ;
  assign n20720 = n20719 ^ n16491 ^ 1'b0 ;
  assign n20721 = n4378 & ~n20720 ;
  assign n20722 = n478 & ~n682 ;
  assign n20723 = ~n2796 & n3992 ;
  assign n20724 = n6360 & ~n20723 ;
  assign n20725 = n20722 | n20724 ;
  assign n20726 = n9569 ^ n7443 ^ 1'b0 ;
  assign n20727 = n20726 ^ n11008 ^ n4346 ;
  assign n20728 = n20725 & ~n20727 ;
  assign n20729 = n963 & n10133 ;
  assign n20730 = n13367 & n20729 ;
  assign n20731 = ~n3726 & n20730 ;
  assign n20732 = n4701 & ~n15468 ;
  assign n20733 = ~n6492 & n20732 ;
  assign n20734 = n3566 | n18317 ;
  assign n20735 = n20733 | n20734 ;
  assign n20736 = n5241 ^ n1136 ^ 1'b0 ;
  assign n20737 = ~n16719 & n20736 ;
  assign n20738 = n20737 ^ n17115 ^ 1'b0 ;
  assign n20739 = ~n676 & n7413 ;
  assign n20740 = n20739 ^ n17629 ^ 1'b0 ;
  assign n20741 = ~n3135 & n20740 ;
  assign n20742 = n10264 & n20741 ;
  assign n20743 = n18961 ^ n4341 ^ 1'b0 ;
  assign n20744 = n15393 & ~n20743 ;
  assign n20745 = n296 & n20744 ;
  assign n20746 = n14749 ^ n3618 ^ 1'b0 ;
  assign n20747 = ~n17268 & n20746 ;
  assign n20748 = n1428 & ~n6608 ;
  assign n20749 = n6608 & n20748 ;
  assign n20750 = n16112 & ~n20749 ;
  assign n20751 = n20750 ^ n6331 ^ 1'b0 ;
  assign n20752 = n1098 & n20514 ;
  assign n20753 = n20752 ^ n2610 ^ 1'b0 ;
  assign n20754 = ~n3146 & n8033 ;
  assign n20755 = n8876 & n20754 ;
  assign n20756 = n20755 ^ n2583 ^ 1'b0 ;
  assign n20757 = n10538 & ~n17209 ;
  assign n20758 = n6578 | n13403 ;
  assign n20759 = n20758 ^ n1520 ^ 1'b0 ;
  assign n20760 = ~n16961 & n20759 ;
  assign n20761 = n14716 ^ n202 ^ 1'b0 ;
  assign n20762 = n2798 ^ n1138 ^ 1'b0 ;
  assign n20763 = n8926 & n20762 ;
  assign n20764 = ~n1434 & n4732 ;
  assign n20765 = n20764 ^ n7086 ^ 1'b0 ;
  assign n20766 = n20763 & n20765 ;
  assign n20767 = n4558 ^ n1238 ^ 1'b0 ;
  assign n20768 = n13554 | n20767 ;
  assign n20769 = n1090 & n3886 ;
  assign n20770 = ( n3245 & ~n9540 ) | ( n3245 & n20769 ) | ( ~n9540 & n20769 ) ;
  assign n20771 = n11412 | n18973 ;
  assign n20772 = n20771 ^ n15177 ^ 1'b0 ;
  assign n20773 = n14904 & n20772 ;
  assign n20774 = n13724 & n15649 ;
  assign n20775 = n1715 & ~n9216 ;
  assign n20776 = n20775 ^ n15760 ^ 1'b0 ;
  assign n20777 = ~n7719 & n10099 ;
  assign n20778 = n20777 ^ n9481 ^ 1'b0 ;
  assign n20779 = n20778 ^ n2421 ^ 1'b0 ;
  assign n20780 = n9389 & ~n20779 ;
  assign n20781 = n9605 ^ n2548 ^ 1'b0 ;
  assign n20782 = n20756 ^ n11931 ^ 1'b0 ;
  assign n20783 = ~n8135 & n20782 ;
  assign n20784 = n4336 ^ n368 ^ 1'b0 ;
  assign n20785 = n412 & n20784 ;
  assign n20786 = n20785 ^ n1469 ^ 1'b0 ;
  assign n20787 = ~n4785 & n18181 ;
  assign n20788 = n11535 ^ n255 ^ 1'b0 ;
  assign n20789 = ~n9028 & n17572 ;
  assign n20790 = ~n1561 & n1853 ;
  assign n20791 = n12525 & n20790 ;
  assign n20792 = ~n1422 & n3068 ;
  assign n20793 = n852 & n20792 ;
  assign n20794 = n4325 & n10123 ;
  assign n20795 = n20793 & n20794 ;
  assign n20796 = n6065 | n11273 ;
  assign n20797 = n4845 ^ n4626 ^ 1'b0 ;
  assign n20798 = n4667 & ~n20797 ;
  assign n20799 = ~n446 & n20798 ;
  assign n20800 = n20796 & ~n20799 ;
  assign n20801 = n20795 & n20800 ;
  assign n20802 = n3293 ^ n3123 ^ 1'b0 ;
  assign n20803 = n20802 ^ n1003 ^ 1'b0 ;
  assign n20804 = n20803 ^ n20048 ^ 1'b0 ;
  assign n20805 = ~n10510 & n20804 ;
  assign n20806 = n1081 | n19663 ;
  assign n20809 = ~n7265 & n8754 ;
  assign n20807 = n7914 & ~n20403 ;
  assign n20808 = n20807 ^ n2175 ^ 1'b0 ;
  assign n20810 = n20809 ^ n20808 ^ n8252 ;
  assign n20811 = n2257 & ~n10948 ;
  assign n20812 = n18494 & n20811 ;
  assign n20813 = n6870 | n15961 ;
  assign n20814 = n20813 ^ n10565 ^ 1'b0 ;
  assign n20815 = ( n11452 & n20812 ) | ( n11452 & n20814 ) | ( n20812 & n20814 ) ;
  assign n20816 = n20810 & ~n20815 ;
  assign n20817 = ~n9908 & n17204 ;
  assign n20818 = n1889 | n2019 ;
  assign n20819 = n20818 ^ n4677 ^ 1'b0 ;
  assign n20820 = n11908 ^ n11308 ^ 1'b0 ;
  assign n20821 = n20820 ^ n11412 ^ 1'b0 ;
  assign n20822 = ~n5010 & n10513 ;
  assign n20823 = n1454 & n20822 ;
  assign n20824 = n2359 | n4483 ;
  assign n20825 = ~n4403 & n16361 ;
  assign n20826 = ~n20824 & n20825 ;
  assign n20827 = n11189 & ~n11605 ;
  assign n20828 = n18445 & n20827 ;
  assign n20829 = ~n17700 & n20828 ;
  assign n20830 = n2046 | n8346 ;
  assign n20831 = n10394 | n20830 ;
  assign n20832 = ~n16949 & n20831 ;
  assign n20833 = ~n9889 & n14751 ;
  assign n20837 = ( n851 & n1912 ) | ( n851 & n2240 ) | ( n1912 & n2240 ) ;
  assign n20838 = n9136 & ~n10300 ;
  assign n20839 = n3646 ^ n1035 ^ 1'b0 ;
  assign n20840 = n20838 | n20839 ;
  assign n20841 = n20837 | n20840 ;
  assign n20842 = n16699 & ~n20841 ;
  assign n20834 = n13475 ^ n8821 ^ 1'b0 ;
  assign n20835 = ~n11585 & n20834 ;
  assign n20836 = n12480 & n20835 ;
  assign n20843 = n20842 ^ n20836 ^ 1'b0 ;
  assign n20844 = n9290 & ~n14242 ;
  assign n20845 = n6110 ^ n5151 ^ n1914 ;
  assign n20846 = n20845 ^ n4683 ^ n2388 ;
  assign n20847 = n3366 | n9287 ;
  assign n20848 = n14877 & ~n20847 ;
  assign n20849 = n18806 ^ n14848 ^ n7041 ;
  assign n20850 = n1009 | n6842 ;
  assign n20851 = n17588 & ~n20850 ;
  assign n20852 = n2743 & n7910 ;
  assign n20853 = n3193 & n20852 ;
  assign n20854 = n20853 ^ n4533 ^ 1'b0 ;
  assign n20855 = n8427 & n20854 ;
  assign n20856 = n17341 | n20855 ;
  assign n20857 = n299 & ~n11169 ;
  assign n20858 = n20857 ^ n10915 ^ 1'b0 ;
  assign n20859 = n2134 & ~n20858 ;
  assign n20860 = ~n19101 & n20859 ;
  assign n20861 = n11527 & ~n18779 ;
  assign n20862 = n20860 & n20861 ;
  assign n20863 = n3335 ^ n3285 ^ 1'b0 ;
  assign n20864 = n6874 | n20863 ;
  assign n20865 = n1340 & n15578 ;
  assign n20866 = n20864 & n20865 ;
  assign n20867 = n20866 ^ n10251 ^ n8665 ;
  assign n20869 = n3501 ^ n2574 ^ 1'b0 ;
  assign n20868 = ~n74 & n5685 ;
  assign n20870 = n20869 ^ n20868 ^ 1'b0 ;
  assign n20871 = n12553 ^ n2197 ^ 1'b0 ;
  assign n20872 = ~n20870 & n20871 ;
  assign n20873 = n20872 ^ n2664 ^ 1'b0 ;
  assign n20874 = n2547 & ~n20873 ;
  assign n20875 = n226 & ~n651 ;
  assign n20876 = n13736 | n20875 ;
  assign n20877 = n9204 & ~n20876 ;
  assign n20878 = n6162 | n11276 ;
  assign n20879 = n9576 | n20878 ;
  assign n20880 = n6366 ^ n3891 ^ 1'b0 ;
  assign n20881 = n5023 & ~n20880 ;
  assign n20882 = n3802 | n11035 ;
  assign n20883 = n74 & ~n6174 ;
  assign n20884 = ~n74 & n20883 ;
  assign n20885 = n6102 & ~n20884 ;
  assign n20886 = n21 | n35 ;
  assign n20887 = n35 & ~n20886 ;
  assign n20888 = n1196 | n20887 ;
  assign n20889 = n20887 & ~n20888 ;
  assign n20890 = n25 & n79 ;
  assign n20891 = ~n79 & n20890 ;
  assign n20892 = n57 & ~n20891 ;
  assign n20893 = n20891 & n20892 ;
  assign n20894 = n358 & ~n2170 ;
  assign n20895 = n2170 & n20894 ;
  assign n20896 = n3235 & ~n20895 ;
  assign n20897 = n20895 & n20896 ;
  assign n20898 = n20893 | n20897 ;
  assign n20899 = n20889 & ~n20898 ;
  assign n20900 = n20885 | n20899 ;
  assign n20901 = n1016 | n20900 ;
  assign n20902 = n19921 ^ n11088 ^ 1'b0 ;
  assign n20903 = n20520 ^ n3289 ^ 1'b0 ;
  assign n20904 = n3361 | n20903 ;
  assign n20905 = n3760 | n20904 ;
  assign n20906 = n6832 & ~n20905 ;
  assign n20907 = n254 & n1648 ;
  assign n20908 = n6328 | n13449 ;
  assign n20909 = n1329 & n20908 ;
  assign n20910 = n7605 & n16795 ;
  assign n20911 = ~n20909 & n20910 ;
  assign n20912 = n20272 ^ n17166 ^ 1'b0 ;
  assign n20913 = n8534 & ~n19555 ;
  assign n20914 = n749 & ~n17167 ;
  assign n20915 = n20914 ^ n1269 ^ 1'b0 ;
  assign n20916 = n8710 ^ n2330 ^ 1'b0 ;
  assign n20920 = x6 & n3044 ;
  assign n20917 = n4142 ^ n2822 ^ 1'b0 ;
  assign n20918 = n20917 ^ n11152 ^ 1'b0 ;
  assign n20919 = n4267 & ~n20918 ;
  assign n20921 = n20920 ^ n20919 ^ 1'b0 ;
  assign n20922 = ~n6332 & n20921 ;
  assign n20923 = n11553 ^ n10231 ^ 1'b0 ;
  assign n20924 = n20848 ^ n17855 ^ 1'b0 ;
  assign n20925 = n4970 | n13869 ;
  assign n20926 = n14053 ^ n1109 ^ 1'b0 ;
  assign n20927 = n20925 | n20926 ;
  assign n20928 = n3562 ^ n1306 ^ 1'b0 ;
  assign n20929 = n2815 & n10753 ;
  assign n20930 = n20929 ^ n3657 ^ 1'b0 ;
  assign n20931 = n20930 ^ n2380 ^ 1'b0 ;
  assign n20932 = n2065 & ~n4063 ;
  assign n20933 = n20370 & n20932 ;
  assign n20934 = n31 | n20933 ;
  assign n20935 = n20934 ^ n10254 ^ 1'b0 ;
  assign n20936 = n8410 ^ n6681 ^ 1'b0 ;
  assign n20937 = n1052 & n17131 ;
  assign n20938 = ~n18363 & n20937 ;
  assign n20939 = n20938 ^ n15700 ^ 1'b0 ;
  assign n20940 = n20936 & ~n20939 ;
  assign n20942 = n1190 & ~n9241 ;
  assign n20943 = n20942 ^ n19193 ^ 1'b0 ;
  assign n20941 = ~n5906 & n17011 ;
  assign n20944 = n20943 ^ n20941 ^ 1'b0 ;
  assign n20945 = n6124 ^ n2460 ^ 1'b0 ;
  assign n20946 = n20944 & n20945 ;
  assign n20947 = n18685 ^ n18417 ^ 1'b0 ;
  assign n20948 = n806 & n11315 ;
  assign n20949 = ~n19935 & n20948 ;
  assign n20950 = n2161 & ~n14095 ;
  assign n20951 = n20950 ^ n16046 ^ 1'b0 ;
  assign n20952 = ~n916 & n13429 ;
  assign n20953 = ~n3023 & n20952 ;
  assign n20954 = n20953 ^ n993 ^ 1'b0 ;
  assign n20956 = ~n8378 & n15268 ;
  assign n20955 = ~n3682 & n14404 ;
  assign n20957 = n20956 ^ n20955 ^ 1'b0 ;
  assign n20958 = ~n390 & n1568 ;
  assign n20959 = ~n16208 & n20958 ;
  assign n20960 = n12995 | n20959 ;
  assign n20961 = n11035 & n17934 ;
  assign n20962 = ~n1999 & n12236 ;
  assign n20963 = n2469 & n20962 ;
  assign n20964 = n20963 ^ n14173 ^ n3664 ;
  assign n20965 = ~n2151 & n6833 ;
  assign n20966 = n8347 ^ n3389 ^ 1'b0 ;
  assign n20967 = ~n20965 & n20966 ;
  assign n20969 = n11283 & n18415 ;
  assign n20968 = n2118 | n18239 ;
  assign n20970 = n20969 ^ n20968 ^ 1'b0 ;
  assign n20971 = n3894 | n10099 ;
  assign n20972 = n4376 & ~n20971 ;
  assign n20973 = n12342 ^ n7031 ^ 1'b0 ;
  assign n20974 = n11030 & ~n20973 ;
  assign n20977 = n5128 & n8105 ;
  assign n20978 = n20977 ^ n829 ^ 1'b0 ;
  assign n20979 = n1211 | n20978 ;
  assign n20980 = n20979 ^ n2595 ^ 1'b0 ;
  assign n20975 = n12123 ^ n7686 ^ 1'b0 ;
  assign n20976 = n659 | n20975 ;
  assign n20981 = n20980 ^ n20976 ^ 1'b0 ;
  assign n20982 = n20974 & n20981 ;
  assign n20983 = n7639 ^ n2028 ^ 1'b0 ;
  assign n20984 = ~n1379 & n16876 ;
  assign n20985 = n17036 ^ n3756 ^ 1'b0 ;
  assign n20986 = n209 & ~n1571 ;
  assign n20987 = n20986 ^ n15569 ^ 1'b0 ;
  assign n20988 = n13087 & ~n20987 ;
  assign n20989 = n1469 | n16150 ;
  assign n20990 = n4174 ^ n1711 ^ n819 ;
  assign n20991 = ~n7787 & n12626 ;
  assign n20992 = n20991 ^ n5033 ^ 1'b0 ;
  assign n20993 = n20990 & ~n20992 ;
  assign n20994 = ~n10381 & n20993 ;
  assign n20995 = n10651 ^ n3731 ^ 1'b0 ;
  assign n20996 = n13202 ^ n7877 ^ n5185 ;
  assign n20997 = n16750 | n20996 ;
  assign n20998 = n20997 ^ n6371 ^ n861 ;
  assign n20999 = n12653 | n15007 ;
  assign n21000 = n20999 ^ n6578 ^ 1'b0 ;
  assign n21001 = n8777 & ~n21000 ;
  assign n21002 = n959 & ~n9361 ;
  assign n21003 = n8930 & n21002 ;
  assign n21004 = n21003 ^ n16033 ^ 1'b0 ;
  assign n21005 = n3940 & ~n16695 ;
  assign n21008 = n2813 | n13383 ;
  assign n21009 = ( ~n10729 & n12059 ) | ( ~n10729 & n21008 ) | ( n12059 & n21008 ) ;
  assign n21006 = n16144 ^ n5022 ^ 1'b0 ;
  assign n21007 = ~n234 & n21006 ;
  assign n21010 = n21009 ^ n21007 ^ 1'b0 ;
  assign n21011 = n1875 & ~n17323 ;
  assign n21012 = n4296 | n7833 ;
  assign n21013 = n10532 & ~n21012 ;
  assign n21014 = n9063 ^ n7252 ^ 1'b0 ;
  assign n21015 = ~n10895 & n21014 ;
  assign n21017 = n2492 & ~n12479 ;
  assign n21016 = n15137 & ~n18777 ;
  assign n21018 = n21017 ^ n21016 ^ 1'b0 ;
  assign n21019 = ( n17775 & n21015 ) | ( n17775 & ~n21018 ) | ( n21015 & ~n21018 ) ;
  assign n21020 = n2656 & ~n13921 ;
  assign n21021 = n6345 & n21020 ;
  assign n21022 = n12280 & ~n21021 ;
  assign n21023 = n21022 ^ n4111 ^ 1'b0 ;
  assign n21024 = n10536 ^ n1205 ^ 1'b0 ;
  assign n21025 = n1378 | n5036 ;
  assign n21026 = n21025 ^ n11692 ^ 1'b0 ;
  assign n21027 = n14472 ^ n1434 ^ 1'b0 ;
  assign n21028 = ( n2134 & n6591 ) | ( n2134 & ~n7848 ) | ( n6591 & ~n7848 ) ;
  assign n21029 = n4605 & n15605 ;
  assign n21030 = ( ~n3906 & n10596 ) | ( ~n3906 & n21029 ) | ( n10596 & n21029 ) ;
  assign n21031 = n9936 ^ n1724 ^ 1'b0 ;
  assign n21032 = n21031 ^ n19273 ^ 1'b0 ;
  assign n21033 = n205 & ~n21032 ;
  assign n21034 = n21030 & n21033 ;
  assign n21037 = n17693 ^ n5844 ^ 1'b0 ;
  assign n21035 = n12656 ^ n10720 ^ 1'b0 ;
  assign n21036 = n2756 & ~n21035 ;
  assign n21038 = n21037 ^ n21036 ^ 1'b0 ;
  assign n21039 = ~n304 & n9058 ;
  assign n21040 = n21039 ^ n1829 ^ 1'b0 ;
  assign n21041 = n21040 ^ n5369 ^ 1'b0 ;
  assign n21042 = ~n10568 & n21041 ;
  assign n21043 = ~n9981 & n12153 ;
  assign n21044 = n2103 & n21043 ;
  assign n21045 = n21044 ^ n10805 ^ n6675 ;
  assign n21046 = ~n21042 & n21045 ;
  assign n21047 = n10504 | n21046 ;
  assign n21049 = ( n3919 & n5147 ) | ( n3919 & n7513 ) | ( n5147 & n7513 ) ;
  assign n21048 = ~n6337 & n7624 ;
  assign n21050 = n21049 ^ n21048 ^ 1'b0 ;
  assign n21051 = n9069 ^ n3753 ^ 1'b0 ;
  assign n21052 = n3437 & ~n21051 ;
  assign n21053 = n6156 & n7544 ;
  assign n21054 = n6102 & n21053 ;
  assign n21055 = n9899 | n21054 ;
  assign n21056 = n21052 | n21055 ;
  assign n21057 = n1528 & n21056 ;
  assign n21058 = ~n1497 & n21057 ;
  assign n21059 = n4438 | n18014 ;
  assign n21060 = ( n6975 & ~n7653 ) | ( n6975 & n15682 ) | ( ~n7653 & n15682 ) ;
  assign n21061 = n3774 & ~n21060 ;
  assign n21062 = n21061 ^ n3992 ^ 1'b0 ;
  assign n21068 = n15819 ^ n5829 ^ 1'b0 ;
  assign n21063 = n5010 & n13852 ;
  assign n21064 = n21063 ^ n17538 ^ 1'b0 ;
  assign n21065 = n21064 ^ n1095 ^ 1'b0 ;
  assign n21066 = ~n14746 & n21065 ;
  assign n21067 = n1876 & ~n21066 ;
  assign n21069 = n21068 ^ n21067 ^ 1'b0 ;
  assign n21070 = n12950 & n14249 ;
  assign n21071 = ~n21069 & n21070 ;
  assign n21072 = n1747 & n5676 ;
  assign n21073 = n21072 ^ n10831 ^ 1'b0 ;
  assign n21074 = n6024 | n21073 ;
  assign n21075 = n21074 ^ n13832 ^ 1'b0 ;
  assign n21076 = n18066 | n21075 ;
  assign n21079 = n5132 ^ n3820 ^ 1'b0 ;
  assign n21077 = n8380 & ~n9274 ;
  assign n21078 = n11909 & ~n21077 ;
  assign n21080 = n21079 ^ n21078 ^ 1'b0 ;
  assign n21081 = n7199 & n9072 ;
  assign n21082 = n15771 & n21081 ;
  assign n21083 = n21080 & n21082 ;
  assign n21084 = n5492 & ~n21083 ;
  assign n21085 = n8152 ^ n3226 ^ 1'b0 ;
  assign n21086 = n13900 & n21085 ;
  assign n21087 = n3791 | n11005 ;
  assign n21088 = n21087 ^ n13231 ^ 1'b0 ;
  assign n21089 = n484 & n21088 ;
  assign n21090 = n14126 ^ n9736 ^ 1'b0 ;
  assign n21091 = n3338 & ~n11714 ;
  assign n21092 = n21090 | n21091 ;
  assign n21094 = n7448 & n19051 ;
  assign n21093 = n1078 & n19057 ;
  assign n21095 = n21094 ^ n21093 ^ 1'b0 ;
  assign n21096 = n2684 & ~n5612 ;
  assign n21097 = n2556 & n21096 ;
  assign n21098 = ( ~n12126 & n20689 ) | ( ~n12126 & n21097 ) | ( n20689 & n21097 ) ;
  assign n21099 = n5405 & ~n21098 ;
  assign n21100 = ~n13376 & n21099 ;
  assign n21101 = ( n5736 & ~n8332 ) | ( n5736 & n18456 ) | ( ~n8332 & n18456 ) ;
  assign n21102 = ( n15110 & n21100 ) | ( n15110 & n21101 ) | ( n21100 & n21101 ) ;
  assign n21103 = n968 & ~n1539 ;
  assign n21104 = n21103 ^ n2767 ^ 1'b0 ;
  assign n21105 = n522 ^ n318 ^ 1'b0 ;
  assign n21106 = n7414 & ~n10177 ;
  assign n21107 = ~n1408 & n21106 ;
  assign n21108 = ( ~n7261 & n21105 ) | ( ~n7261 & n21107 ) | ( n21105 & n21107 ) ;
  assign n21109 = n6749 & ~n20682 ;
  assign n21110 = n8591 ^ n5385 ^ 1'b0 ;
  assign n21111 = n9772 & ~n21110 ;
  assign n21112 = ~n2101 & n21111 ;
  assign n21113 = ~n9766 & n12622 ;
  assign n21114 = n21112 & n21113 ;
  assign n21115 = ( ~n3674 & n9584 ) | ( ~n3674 & n10550 ) | ( n9584 & n10550 ) ;
  assign n21116 = ~n3731 & n18393 ;
  assign n21117 = n4977 & n7027 ;
  assign n21118 = n9173 ^ n3403 ^ 1'b0 ;
  assign n21119 = n5034 & ~n21118 ;
  assign n21120 = ~n5663 & n11358 ;
  assign n21121 = n21120 ^ n10235 ^ 1'b0 ;
  assign n21123 = n3992 ^ n371 ^ 1'b0 ;
  assign n21124 = n3887 | n21123 ;
  assign n21122 = n5010 & n12222 ;
  assign n21125 = n21124 ^ n21122 ^ 1'b0 ;
  assign n21126 = n21125 ^ n1460 ^ 1'b0 ;
  assign n21127 = n10106 ^ n835 ^ 1'b0 ;
  assign n21128 = n3915 | n21127 ;
  assign n21129 = n3915 & ~n21128 ;
  assign n21130 = n150 | n8084 ;
  assign n21131 = n21130 ^ n12441 ^ n6124 ;
  assign n21132 = n7042 ^ n2847 ^ n1445 ;
  assign n21133 = ( n2248 & ~n4537 ) | ( n2248 & n21132 ) | ( ~n4537 & n21132 ) ;
  assign n21134 = n5073 ^ n474 ^ 1'b0 ;
  assign n21135 = n4788 | n19377 ;
  assign n21136 = n4962 ^ n1659 ^ 1'b0 ;
  assign n21137 = n21135 | n21136 ;
  assign n21138 = n17027 ^ n12177 ^ 1'b0 ;
  assign n21139 = n19228 | n21138 ;
  assign n21140 = n6213 & ~n16020 ;
  assign n21141 = n10137 & ~n21140 ;
  assign n21142 = n21141 ^ n12889 ^ 1'b0 ;
  assign n21143 = n18788 ^ n17178 ^ 1'b0 ;
  assign n21144 = n12284 | n21143 ;
  assign n21145 = n20131 ^ n5733 ^ 1'b0 ;
  assign n21146 = n17224 ^ n11791 ^ 1'b0 ;
  assign n21147 = n10134 & n21146 ;
  assign n21148 = n10177 & n21147 ;
  assign n21149 = n8553 | n15945 ;
  assign n21150 = n4168 & ~n6982 ;
  assign n21151 = ~n15411 & n21150 ;
  assign n21152 = n16578 ^ n13354 ^ n13279 ;
  assign n21153 = n19826 | n21152 ;
  assign n21154 = ( n7349 & n7808 ) | ( n7349 & n18735 ) | ( n7808 & n18735 ) ;
  assign n21155 = ( ~n541 & n1103 ) | ( ~n541 & n3300 ) | ( n1103 & n3300 ) ;
  assign n21156 = n21155 ^ n1304 ^ 1'b0 ;
  assign n21157 = n16657 ^ n2228 ^ 1'b0 ;
  assign n21158 = ~n21156 & n21157 ;
  assign n21159 = n3687 ^ n1786 ^ 1'b0 ;
  assign n21160 = n10385 & n21159 ;
  assign n21161 = n19556 ^ n5857 ^ n5592 ;
  assign n21162 = n21161 ^ n9753 ^ n4203 ;
  assign n21163 = ~n1865 & n14177 ;
  assign n21164 = ~n262 & n5332 ;
  assign n21165 = n21163 & n21164 ;
  assign n21166 = n18192 | n21165 ;
  assign n21173 = n8062 ^ n7076 ^ 1'b0 ;
  assign n21167 = n339 & n7927 ;
  assign n21168 = n4413 & n21167 ;
  assign n21169 = n21168 ^ n5872 ^ 1'b0 ;
  assign n21170 = n10168 | n21169 ;
  assign n21171 = n6460 | n15089 ;
  assign n21172 = ~n21170 & n21171 ;
  assign n21174 = n21173 ^ n21172 ^ 1'b0 ;
  assign n21175 = n17100 & ~n20378 ;
  assign n21176 = n5375 ^ n2981 ^ 1'b0 ;
  assign n21177 = ~n2588 & n21176 ;
  assign n21178 = n21177 ^ n749 ^ 1'b0 ;
  assign n21179 = n13016 & ~n21178 ;
  assign n21180 = n5402 & n12120 ;
  assign n21181 = n21180 ^ n17099 ^ 1'b0 ;
  assign n21182 = n1177 & ~n8573 ;
  assign n21183 = ( ~n1853 & n9970 ) | ( ~n1853 & n18961 ) | ( n9970 & n18961 ) ;
  assign n21184 = n4059 ^ n3726 ^ 1'b0 ;
  assign n21185 = n21184 ^ n949 ^ 1'b0 ;
  assign n21186 = n8712 & n21185 ;
  assign n21187 = ( n6351 & n21183 ) | ( n6351 & n21186 ) | ( n21183 & n21186 ) ;
  assign n21188 = ~n908 & n21187 ;
  assign n21189 = ~n4331 & n21188 ;
  assign n21190 = n21189 ^ n7075 ^ 1'b0 ;
  assign n21191 = n4805 & n21190 ;
  assign n21192 = n277 | n3054 ;
  assign n21193 = n21192 ^ n11378 ^ 1'b0 ;
  assign n21194 = n11364 | n21193 ;
  assign n21195 = ( ~n7452 & n10349 ) | ( ~n7452 & n18292 ) | ( n10349 & n18292 ) ;
  assign n21199 = n11711 ^ n4328 ^ 1'b0 ;
  assign n21200 = n16607 | n21199 ;
  assign n21196 = n13831 ^ n2494 ^ 1'b0 ;
  assign n21197 = n12361 & ~n21196 ;
  assign n21198 = n2940 & n21197 ;
  assign n21201 = n21200 ^ n21198 ^ 1'b0 ;
  assign n21202 = n7375 ^ n2706 ^ 1'b0 ;
  assign n21203 = n5332 & ~n21202 ;
  assign n21204 = n7604 ^ n3745 ^ 1'b0 ;
  assign n21205 = n6808 | n18707 ;
  assign n21206 = n1550 & ~n21205 ;
  assign n21207 = ~n9660 & n21206 ;
  assign n21208 = n12701 ^ n12501 ^ 1'b0 ;
  assign n21209 = n15951 ^ n7965 ^ 1'b0 ;
  assign n21210 = n9616 ^ n9388 ^ 1'b0 ;
  assign n21211 = n2370 & n9943 ;
  assign n21212 = n4048 | n21211 ;
  assign n21213 = n21212 ^ n1902 ^ 1'b0 ;
  assign n21214 = ~n11906 & n21213 ;
  assign n21215 = n3611 & n12496 ;
  assign n21216 = n17393 ^ n4368 ^ 1'b0 ;
  assign n21217 = n7973 ^ n6968 ^ 1'b0 ;
  assign n21218 = ( ~n13794 & n18519 ) | ( ~n13794 & n21217 ) | ( n18519 & n21217 ) ;
  assign n21219 = n3199 | n20191 ;
  assign n21220 = n7361 | n9222 ;
  assign n21221 = n21220 ^ n6410 ^ 1'b0 ;
  assign n21222 = n4226 | n21221 ;
  assign n21223 = n8782 | n21222 ;
  assign n21224 = n1327 & n16253 ;
  assign n21225 = ~n10265 & n21224 ;
  assign n21226 = n6348 & ~n8723 ;
  assign n21227 = n640 & ~n5881 ;
  assign n21228 = n5167 ^ n2812 ^ 1'b0 ;
  assign n21229 = n1260 | n21228 ;
  assign n21230 = n3482 ^ n438 ^ 1'b0 ;
  assign n21231 = n4857 & n21230 ;
  assign n21232 = n21229 & n21231 ;
  assign n21233 = n6136 & ~n21232 ;
  assign n21234 = n7621 | n17172 ;
  assign n21235 = n13487 | n21234 ;
  assign n21236 = n7795 & n9589 ;
  assign n21237 = n2062 & n5936 ;
  assign n21238 = ~n10978 & n18941 ;
  assign n21239 = n21237 & n21238 ;
  assign n21240 = n11645 | n13402 ;
  assign n21241 = n3035 & ~n21240 ;
  assign n21242 = ( n1163 & n21239 ) | ( n1163 & n21241 ) | ( n21239 & n21241 ) ;
  assign n21243 = ~n6893 & n10603 ;
  assign n21244 = n15444 ^ n6640 ^ 1'b0 ;
  assign n21245 = n3400 ^ n2772 ^ 1'b0 ;
  assign n21246 = n21245 ^ n19846 ^ 1'b0 ;
  assign n21248 = n1182 & n1275 ;
  assign n21249 = n7045 & n21248 ;
  assign n21247 = n6051 | n7839 ;
  assign n21250 = n21249 ^ n21247 ^ 1'b0 ;
  assign n21251 = n3502 ^ n1385 ^ 1'b0 ;
  assign n21252 = ~n2773 & n21251 ;
  assign n21253 = n21252 ^ n5555 ^ 1'b0 ;
  assign n21254 = n21253 ^ n18889 ^ 1'b0 ;
  assign n21256 = n4746 ^ n875 ^ 1'b0 ;
  assign n21255 = n15633 ^ n3971 ^ 1'b0 ;
  assign n21257 = n21256 ^ n21255 ^ n10769 ;
  assign n21261 = n5748 | n6831 ;
  assign n21259 = n4939 | n11852 ;
  assign n21258 = ~n4960 & n5875 ;
  assign n21260 = n21259 ^ n21258 ^ 1'b0 ;
  assign n21262 = n21261 ^ n21260 ^ 1'b0 ;
  assign n21263 = n9111 & ~n21262 ;
  assign n21264 = ~n5147 & n21049 ;
  assign n21265 = ~n8166 & n21264 ;
  assign n21266 = n21265 ^ n12426 ^ n2615 ;
  assign n21267 = ~n1143 & n11435 ;
  assign n21268 = n15293 & n21267 ;
  assign n21269 = n15407 ^ n6155 ^ n875 ;
  assign n21270 = n6771 ^ n5107 ^ 1'b0 ;
  assign n21271 = ~n14841 & n21270 ;
  assign n21272 = n21271 ^ n16588 ^ n1853 ;
  assign n21273 = n15523 & n19281 ;
  assign n21274 = n21273 ^ n2492 ^ 1'b0 ;
  assign n21275 = n4103 | n19226 ;
  assign n21276 = n5905 & ~n21275 ;
  assign n21277 = ~n1637 & n19267 ;
  assign n21278 = n3464 | n21277 ;
  assign n21279 = n21278 ^ n2288 ^ 1'b0 ;
  assign n21280 = n21279 ^ n14841 ^ 1'b0 ;
  assign n21281 = n14896 & ~n21280 ;
  assign n21282 = n17883 ^ n6445 ^ 1'b0 ;
  assign n21283 = n8773 & ~n21282 ;
  assign n21284 = n21283 ^ n15966 ^ n11414 ;
  assign n21285 = n419 | n4145 ;
  assign n21286 = n19341 ^ n1045 ^ 1'b0 ;
  assign n21287 = n1786 | n7259 ;
  assign n21288 = n2388 | n2492 ;
  assign n21289 = n8658 | n21288 ;
  assign n21290 = n16120 & n21289 ;
  assign n21291 = ~n4890 & n21290 ;
  assign n21292 = n21287 | n21291 ;
  assign n21293 = ~n1576 & n5880 ;
  assign n21294 = n21293 ^ n8745 ^ 1'b0 ;
  assign n21295 = n3674 | n12715 ;
  assign n21296 = n8080 & ~n15459 ;
  assign n21297 = n16073 & n21296 ;
  assign n21298 = ~n3955 & n9928 ;
  assign n21299 = n8223 & n11735 ;
  assign n21300 = n18548 ^ n6310 ^ 1'b0 ;
  assign n21301 = n3732 & ~n12288 ;
  assign n21302 = n11620 ^ n1969 ^ 1'b0 ;
  assign n21303 = n5644 | n21302 ;
  assign n21304 = ~n3923 & n21303 ;
  assign n21305 = n21304 ^ n2309 ^ 1'b0 ;
  assign n21306 = n5684 & n10908 ;
  assign n21307 = n3111 ^ n968 ^ 1'b0 ;
  assign n21308 = n2909 & n15236 ;
  assign n21309 = n4474 ^ n1056 ^ 1'b0 ;
  assign n21310 = n18864 | n21309 ;
  assign n21311 = n21308 & ~n21310 ;
  assign n21312 = ~n4785 & n5662 ;
  assign n21313 = ~n1304 & n21312 ;
  assign n21319 = ~n144 & n7761 ;
  assign n21314 = n5393 & ~n11560 ;
  assign n21315 = n21314 ^ n7184 ^ 1'b0 ;
  assign n21316 = n1403 | n4447 ;
  assign n21317 = n21316 ^ n8171 ^ 1'b0 ;
  assign n21318 = ( n3535 & n21315 ) | ( n3535 & n21317 ) | ( n21315 & n21317 ) ;
  assign n21320 = n21319 ^ n21318 ^ n1810 ;
  assign n21321 = ( n14750 & n21313 ) | ( n14750 & ~n21320 ) | ( n21313 & ~n21320 ) ;
  assign n21322 = n1454 | n9153 ;
  assign n21323 = n21322 ^ n3080 ^ 1'b0 ;
  assign n21324 = n3461 & n4335 ;
  assign n21325 = n14052 ^ n11077 ^ n2833 ;
  assign n21326 = n21325 ^ n12913 ^ 1'b0 ;
  assign n21327 = n21324 & ~n21326 ;
  assign n21328 = n21327 ^ n1215 ^ 1'b0 ;
  assign n21329 = n1245 & n3400 ;
  assign n21330 = n21329 ^ n3828 ^ n1307 ;
  assign n21331 = n6456 ^ n3848 ^ n2428 ;
  assign n21332 = n9272 ^ n2666 ^ 1'b0 ;
  assign n21333 = n1796 | n21332 ;
  assign n21334 = ~n16750 & n21333 ;
  assign n21335 = n6486 | n7154 ;
  assign n21336 = n21334 & n21335 ;
  assign n21337 = ~n2893 & n21336 ;
  assign n21338 = n2899 & n11052 ;
  assign n21339 = n21338 ^ n5145 ^ 1'b0 ;
  assign n21340 = n545 & ~n21339 ;
  assign n21341 = n21337 & n21340 ;
  assign n21342 = n576 & ~n21341 ;
  assign n21343 = n21331 & n21342 ;
  assign n21344 = n3574 | n7975 ;
  assign n21345 = n551 & n21344 ;
  assign n21346 = n21345 ^ n8163 ^ 1'b0 ;
  assign n21347 = n61 & ~n2790 ;
  assign n21348 = ~n11469 & n18043 ;
  assign n21349 = n21348 ^ n10572 ^ 1'b0 ;
  assign n21350 = n15161 | n21349 ;
  assign n21351 = n18912 & n21350 ;
  assign n21352 = n974 ^ n948 ^ 1'b0 ;
  assign n21353 = n3885 & ~n21352 ;
  assign n21354 = n9534 ^ n9085 ^ 1'b0 ;
  assign n21355 = n1234 & n21354 ;
  assign n21356 = n21353 & n21355 ;
  assign n21357 = n21356 ^ n11359 ^ 1'b0 ;
  assign n21358 = n1663 & ~n2481 ;
  assign n21359 = n2481 & n21358 ;
  assign n21360 = n3090 & n21359 ;
  assign n21361 = ~n7027 & n21360 ;
  assign n21362 = ~n6043 & n21361 ;
  assign n21363 = n21362 ^ n4468 ^ 1'b0 ;
  assign n21364 = n21363 ^ n16639 ^ 1'b0 ;
  assign n21365 = n1502 & ~n21364 ;
  assign n21366 = n965 | n8555 ;
  assign n21367 = n18283 & n21366 ;
  assign n21368 = ~n796 & n21367 ;
  assign n21369 = n14088 ^ n4937 ^ 1'b0 ;
  assign n21370 = n12123 ^ n4579 ^ 1'b0 ;
  assign n21371 = ~n7771 & n21370 ;
  assign n21372 = n16113 & n21371 ;
  assign n21373 = ~n17964 & n21372 ;
  assign n21374 = n21373 ^ n15023 ^ 1'b0 ;
  assign n21375 = ~n1161 & n21374 ;
  assign n21376 = n15614 ^ n12218 ^ 1'b0 ;
  assign n21377 = ~n899 & n7981 ;
  assign n21378 = n21377 ^ n4824 ^ 1'b0 ;
  assign n21379 = n21378 ^ n6880 ^ 1'b0 ;
  assign n21380 = n20108 ^ n15389 ^ 1'b0 ;
  assign n21381 = n13117 | n21380 ;
  assign n21382 = n3012 | n4698 ;
  assign n21383 = n21382 ^ n20689 ^ n9780 ;
  assign n21387 = ( ~n1944 & n6545 ) | ( ~n1944 & n8721 ) | ( n6545 & n8721 ) ;
  assign n21384 = n6491 ^ n135 ^ 1'b0 ;
  assign n21385 = ~n2380 & n21384 ;
  assign n21386 = n4335 & n21385 ;
  assign n21388 = n21387 ^ n21386 ^ 1'b0 ;
  assign n21389 = n1419 & n7669 ;
  assign n21390 = n1479 & ~n6572 ;
  assign n21391 = n4787 & n7626 ;
  assign n21392 = n1439 & ~n5954 ;
  assign n21393 = ~n2143 & n21392 ;
  assign n21394 = n21391 & ~n21393 ;
  assign n21395 = ~n21390 & n21394 ;
  assign n21396 = n6766 | n21395 ;
  assign n21397 = n1306 & ~n21396 ;
  assign n21398 = n5141 ^ n4077 ^ 1'b0 ;
  assign n21399 = n21398 ^ n1083 ^ 1'b0 ;
  assign n21400 = n3232 & ~n21399 ;
  assign n21401 = n6738 & n6871 ;
  assign n21402 = n21401 ^ n8979 ^ 1'b0 ;
  assign n21403 = n4054 | n5292 ;
  assign n21404 = n21402 | n21403 ;
  assign n21406 = n15807 ^ n12211 ^ 1'b0 ;
  assign n21407 = n6114 | n21406 ;
  assign n21405 = ~n11209 & n16062 ;
  assign n21408 = n21407 ^ n21405 ^ n12878 ;
  assign n21409 = n8584 & n16301 ;
  assign n21410 = n3552 | n7676 ;
  assign n21411 = ( n2366 & n20009 ) | ( n2366 & ~n21410 ) | ( n20009 & ~n21410 ) ;
  assign n21412 = n8051 | n21411 ;
  assign n21413 = n541 & n839 ;
  assign n21414 = ~n5744 & n9189 ;
  assign n21415 = n8072 | n18973 ;
  assign n21416 = n21415 ^ n1981 ^ 1'b0 ;
  assign n21417 = n12694 ^ n9938 ^ 1'b0 ;
  assign n21418 = n11810 ^ n4002 ^ 1'b0 ;
  assign n21419 = n7027 & ~n16010 ;
  assign n21420 = ( n611 & n21418 ) | ( n611 & n21419 ) | ( n21418 & n21419 ) ;
  assign n21421 = n1897 | n5001 ;
  assign n21422 = n21421 ^ n3408 ^ 1'b0 ;
  assign n21423 = ~n4159 & n12369 ;
  assign n21424 = n21423 ^ n13998 ^ 1'b0 ;
  assign n21425 = n15821 ^ n6147 ^ 1'b0 ;
  assign n21426 = n9938 & ~n21425 ;
  assign n21427 = n7749 ^ n2813 ^ 1'b0 ;
  assign n21428 = n21427 ^ n2120 ^ n749 ;
  assign n21429 = ~n16004 & n21428 ;
  assign n21430 = n20498 & n21429 ;
  assign n21431 = ~n3411 & n21430 ;
  assign n21432 = n3465 ^ n69 ^ 1'b0 ;
  assign n21433 = n21432 ^ n10790 ^ n559 ;
  assign n21434 = n21433 ^ n16160 ^ n9832 ;
  assign n21435 = n21434 ^ n20603 ^ 1'b0 ;
  assign n21436 = n5755 ^ n3410 ^ 1'b0 ;
  assign n21437 = n14845 & ~n21436 ;
  assign n21438 = n21437 ^ n19705 ^ 1'b0 ;
  assign n21439 = n1346 & n19611 ;
  assign n21440 = ( n1231 & n3584 ) | ( n1231 & n19798 ) | ( n3584 & n19798 ) ;
  assign n21441 = n2522 ^ n1657 ^ 1'b0 ;
  assign n21442 = n5380 & ~n21441 ;
  assign n21443 = n21442 ^ n13913 ^ 1'b0 ;
  assign n21444 = n7686 | n21287 ;
  assign n21445 = n11225 ^ n5493 ^ 1'b0 ;
  assign n21446 = ~n17243 & n21445 ;
  assign n21447 = n21446 ^ n9995 ^ 1'b0 ;
  assign n21448 = n5649 & n21447 ;
  assign n21449 = n21448 ^ n3513 ^ 1'b0 ;
  assign n21450 = ~n21444 & n21449 ;
  assign n21451 = n2521 & n21450 ;
  assign n21452 = ( n13450 & n17650 ) | ( n13450 & n21451 ) | ( n17650 & n21451 ) ;
  assign n21453 = n21452 ^ n12024 ^ 1'b0 ;
  assign n21454 = n18923 ^ n372 ^ 1'b0 ;
  assign n21455 = ~n4275 & n12168 ;
  assign n21456 = n21455 ^ n17575 ^ 1'b0 ;
  assign n21457 = ~n10445 & n21456 ;
  assign n21458 = n3847 ^ n1020 ^ 1'b0 ;
  assign n21459 = n1116 & ~n21458 ;
  assign n21460 = n3462 ^ n2233 ^ 1'b0 ;
  assign n21461 = n4366 & n21460 ;
  assign n21462 = n21461 ^ n17620 ^ 1'b0 ;
  assign n21463 = n21459 & ~n21462 ;
  assign n21464 = n8183 & n21463 ;
  assign n21465 = n3535 & n5517 ;
  assign n21466 = n21465 ^ n10270 ^ 1'b0 ;
  assign n21467 = n21466 ^ n12851 ^ n3390 ;
  assign n21468 = ( n3320 & n9270 ) | ( n3320 & ~n12377 ) | ( n9270 & ~n12377 ) ;
  assign n21469 = n1157 | n21468 ;
  assign n21470 = n16167 ^ n1723 ^ 1'b0 ;
  assign n21471 = n20123 ^ n5081 ^ 1'b0 ;
  assign n21472 = ~n8710 & n21471 ;
  assign n21473 = n1045 & ~n1972 ;
  assign n21474 = n16957 & n21473 ;
  assign n21475 = n4053 | n10322 ;
  assign n21476 = n3818 | n21475 ;
  assign n21477 = n8980 ^ n403 ^ 1'b0 ;
  assign n21478 = n6000 & n21477 ;
  assign n21479 = n21478 ^ n1029 ^ 1'b0 ;
  assign n21480 = n214 & ~n21479 ;
  assign n21481 = ~n8702 & n21480 ;
  assign n21482 = n21481 ^ n5080 ^ 1'b0 ;
  assign n21483 = n5010 | n10056 ;
  assign n21484 = n16793 & ~n21483 ;
  assign n21485 = n6895 & n8584 ;
  assign n21486 = n5886 ^ n611 ^ 1'b0 ;
  assign n21487 = n588 | n2082 ;
  assign n21488 = ~n664 & n9766 ;
  assign n21489 = n745 | n10173 ;
  assign n21490 = n1300 | n6584 ;
  assign n21491 = n16924 & ~n21490 ;
  assign n21492 = n6553 ^ n725 ^ 1'b0 ;
  assign n21493 = n18823 & ~n21492 ;
  assign n21494 = n12673 ^ n1326 ^ 1'b0 ;
  assign n21495 = n21493 & ~n21494 ;
  assign n21497 = n11052 ^ n3238 ^ 1'b0 ;
  assign n21498 = n8874 & n21497 ;
  assign n21496 = n20615 ^ n7160 ^ 1'b0 ;
  assign n21499 = n21498 ^ n21496 ^ 1'b0 ;
  assign n21500 = ( n5364 & ~n8034 ) | ( n5364 & n10705 ) | ( ~n8034 & n10705 ) ;
  assign n21501 = n14668 & ~n21500 ;
  assign n21502 = ~n4581 & n12875 ;
  assign n21503 = n3706 & n7549 ;
  assign n21504 = n21503 ^ n623 ^ 1'b0 ;
  assign n21505 = n21504 ^ n2697 ^ 1'b0 ;
  assign n21506 = n18511 ^ n16933 ^ 1'b0 ;
  assign n21507 = ( n74 & ~n7268 ) | ( n74 & n16536 ) | ( ~n7268 & n16536 ) ;
  assign n21508 = n21507 ^ n11543 ^ n802 ;
  assign n21509 = n10787 ^ n2872 ^ 1'b0 ;
  assign n21510 = n8260 ^ n3738 ^ 1'b0 ;
  assign n21511 = n17583 & ~n21510 ;
  assign n21512 = n13218 ^ n806 ^ 1'b0 ;
  assign n21513 = ~n11037 & n20802 ;
  assign n21514 = n21513 ^ n9598 ^ 1'b0 ;
  assign n21515 = n12337 ^ n10945 ^ n2134 ;
  assign n21516 = n21515 ^ n93 ^ 1'b0 ;
  assign n21517 = n10703 & n20403 ;
  assign n21518 = ~n5001 & n21517 ;
  assign n21519 = n21518 ^ n7164 ^ 1'b0 ;
  assign n21520 = n1829 & ~n21519 ;
  assign n21521 = n19525 & n21520 ;
  assign n21522 = ~n21516 & n21521 ;
  assign n21523 = ~n11918 & n12240 ;
  assign n21524 = n5155 & ~n12544 ;
  assign n21525 = n21523 & n21524 ;
  assign n21526 = n3488 | n13147 ;
  assign n21527 = n7799 | n21526 ;
  assign n21528 = n768 & ~n21009 ;
  assign n21529 = n16623 & n21528 ;
  assign n21530 = n8633 & ~n14180 ;
  assign n21531 = ~n1570 & n21530 ;
  assign n21532 = n21531 ^ n5751 ^ 1'b0 ;
  assign n21533 = n3892 | n7137 ;
  assign n21534 = n21533 ^ n15714 ^ 1'b0 ;
  assign n21535 = ~n6283 & n14694 ;
  assign n21536 = n21535 ^ n6212 ^ n821 ;
  assign n21537 = ~n3445 & n21536 ;
  assign n21538 = n21534 & ~n21537 ;
  assign n21539 = ~n21532 & n21538 ;
  assign n21540 = n4850 ^ n225 ^ 1'b0 ;
  assign n21541 = n12661 | n21540 ;
  assign n21542 = n4949 | n21541 ;
  assign n21543 = n15960 & ~n19902 ;
  assign n21544 = n5418 & n21543 ;
  assign n21545 = n10300 ^ n3093 ^ 1'b0 ;
  assign n21546 = n21545 ^ n1434 ^ 1'b0 ;
  assign n21547 = n1161 | n1342 ;
  assign n21548 = n17377 | n21547 ;
  assign n21549 = n21548 ^ n10897 ^ n5276 ;
  assign n21550 = ~n10582 & n10589 ;
  assign n21551 = ~n21549 & n21550 ;
  assign n21552 = n5648 ^ n2545 ^ 1'b0 ;
  assign n21553 = n5695 | n7377 ;
  assign n21554 = n179 & ~n21553 ;
  assign n21555 = n4075 ^ n1277 ^ 1'b0 ;
  assign n21556 = n3531 & n21555 ;
  assign n21557 = n6474 ^ n518 ^ 1'b0 ;
  assign n21558 = n21557 ^ n1845 ^ 1'b0 ;
  assign n21559 = n7126 & ~n21558 ;
  assign n21560 = n7889 & n21559 ;
  assign n21561 = n4470 & n6339 ;
  assign n21562 = n21561 ^ n5646 ^ 1'b0 ;
  assign n21563 = n1205 | n6818 ;
  assign n21564 = n4801 | n21563 ;
  assign n21565 = n21564 ^ n3393 ^ n1920 ;
  assign n21566 = n11338 ^ n11277 ^ 1'b0 ;
  assign n21567 = ~n6155 & n7877 ;
  assign n21568 = n1313 & n21567 ;
  assign n21569 = ~n21566 & n21568 ;
  assign n21570 = n21565 | n21569 ;
  assign n21571 = n3107 & ~n21570 ;
  assign n21572 = n1419 ^ n393 ^ 1'b0 ;
  assign n21573 = n4714 & n21572 ;
  assign n21574 = ~n4400 & n21573 ;
  assign n21575 = n4856 & n21574 ;
  assign n21576 = ~n4804 & n21575 ;
  assign n21577 = n892 & n12713 ;
  assign n21578 = ~n2405 & n21577 ;
  assign n21579 = n21578 ^ n18740 ^ 1'b0 ;
  assign n21580 = n21579 ^ n1861 ^ 1'b0 ;
  assign n21581 = n21467 & n21580 ;
  assign n21582 = ~n17325 & n18347 ;
  assign n21583 = n16021 ^ n15619 ^ n6903 ;
  assign n21584 = ( n315 & ~n8049 ) | ( n315 & n21583 ) | ( ~n8049 & n21583 ) ;
  assign n21586 = n2381 & n13407 ;
  assign n21585 = n15368 | n16016 ;
  assign n21587 = n21586 ^ n21585 ^ 1'b0 ;
  assign n21591 = n9913 ^ n9268 ^ n8702 ;
  assign n21588 = n3574 | n7151 ;
  assign n21589 = n21588 ^ n5136 ^ 1'b0 ;
  assign n21590 = ~n19050 & n21589 ;
  assign n21592 = n21591 ^ n21590 ^ 1'b0 ;
  assign n21593 = ~n3099 & n5209 ;
  assign n21594 = n1264 & n21593 ;
  assign n21595 = n790 & n1254 ;
  assign n21596 = n21595 ^ n19802 ^ 1'b0 ;
  assign n21598 = n9571 & ~n13341 ;
  assign n21597 = n2399 ^ n2050 ^ 1'b0 ;
  assign n21599 = n21598 ^ n21597 ^ 1'b0 ;
  assign n21600 = n4213 | n20177 ;
  assign n21601 = ~n13990 & n15289 ;
  assign n21602 = n21601 ^ n16697 ^ 1'b0 ;
  assign n21603 = ~n14244 & n19458 ;
  assign n21604 = n21603 ^ n10426 ^ 1'b0 ;
  assign n21606 = n21398 ^ n6895 ^ 1'b0 ;
  assign n21605 = ~n2567 & n7536 ;
  assign n21607 = n21606 ^ n21605 ^ 1'b0 ;
  assign n21608 = n19356 ^ n15752 ^ 1'b0 ;
  assign n21611 = n4564 & n13157 ;
  assign n21609 = ~n11227 & n11454 ;
  assign n21610 = n10467 & n21609 ;
  assign n21612 = n21611 ^ n21610 ^ n7589 ;
  assign n21616 = n5513 ^ n1325 ^ 1'b0 ;
  assign n21613 = n11007 ^ n7735 ^ 1'b0 ;
  assign n21614 = n404 | n21613 ;
  assign n21615 = n8441 | n21614 ;
  assign n21617 = n21616 ^ n21615 ^ n214 ;
  assign n21618 = n4038 ^ n315 ^ 1'b0 ;
  assign n21619 = ( ~n8871 & n15051 ) | ( ~n8871 & n15699 ) | ( n15051 & n15699 ) ;
  assign n21620 = n13293 ^ n5573 ^ 1'b0 ;
  assign n21621 = ~n21619 & n21620 ;
  assign n21622 = n11180 & n21621 ;
  assign n21623 = n21618 & n21622 ;
  assign n21624 = n5201 | n21623 ;
  assign n21625 = n792 | n7466 ;
  assign n21626 = n21625 ^ n18579 ^ 1'b0 ;
  assign n21627 = n15423 ^ n15008 ^ 1'b0 ;
  assign n21628 = n10050 | n21627 ;
  assign n21629 = n5077 & ~n6375 ;
  assign n21630 = ~n6576 & n8338 ;
  assign n21631 = ( n4005 & n21629 ) | ( n4005 & n21630 ) | ( n21629 & n21630 ) ;
  assign n21632 = n21631 ^ n20268 ^ n3402 ;
  assign n21634 = ( n2172 & ~n3165 ) | ( n2172 & n8363 ) | ( ~n3165 & n8363 ) ;
  assign n21635 = n3355 | n21634 ;
  assign n21636 = n1594 | n21635 ;
  assign n21633 = n7718 & ~n14988 ;
  assign n21637 = n21636 ^ n21633 ^ 1'b0 ;
  assign n21638 = n19746 & n20001 ;
  assign n21639 = n3095 | n5637 ;
  assign n21640 = n7986 & ~n21639 ;
  assign n21641 = n4245 & n21640 ;
  assign n21642 = n6057 & n11249 ;
  assign n21643 = n61 & n21642 ;
  assign n21644 = n8347 & ~n18799 ;
  assign n21651 = ( n9122 & n9697 ) | ( n9122 & n14123 ) | ( n9697 & n14123 ) ;
  assign n21649 = n20559 ^ n2032 ^ 1'b0 ;
  assign n21647 = n6176 | n9485 ;
  assign n21645 = n3050 | n16709 ;
  assign n21646 = ~n13173 & n21645 ;
  assign n21648 = n21647 ^ n21646 ^ 1'b0 ;
  assign n21650 = n21649 ^ n21648 ^ n1700 ;
  assign n21652 = n21651 ^ n21650 ^ 1'b0 ;
  assign n21653 = ( n3472 & ~n10910 ) | ( n3472 & n12994 ) | ( ~n10910 & n12994 ) ;
  assign n21654 = n12919 ^ n7771 ^ 1'b0 ;
  assign n21655 = n21653 & n21654 ;
  assign n21656 = ~n533 & n14710 ;
  assign n21657 = n6537 & n21656 ;
  assign n21658 = n9970 | n17500 ;
  assign n21659 = n21657 & ~n21658 ;
  assign n21660 = n14032 & n17418 ;
  assign n21661 = n17554 & ~n21660 ;
  assign n21662 = n16831 & n21661 ;
  assign n21663 = n17880 ^ n2549 ^ 1'b0 ;
  assign n21664 = n21663 ^ n12594 ^ 1'b0 ;
  assign n21665 = ( n7242 & ~n10866 ) | ( n7242 & n21664 ) | ( ~n10866 & n21664 ) ;
  assign n21666 = ~n518 & n4912 ;
  assign n21667 = n18939 ^ n12847 ^ 1'b0 ;
  assign n21668 = n21666 & n21667 ;
  assign n21669 = n1521 | n21244 ;
  assign n21670 = n21669 ^ n17025 ^ 1'b0 ;
  assign n21671 = n17714 & ~n21228 ;
  assign n21672 = ~n5349 & n21671 ;
  assign n21673 = n14646 ^ n3972 ^ 1'b0 ;
  assign n21674 = n21 | n21673 ;
  assign n21675 = n21674 ^ n8061 ^ 1'b0 ;
  assign n21676 = n18731 ^ n11157 ^ 1'b0 ;
  assign n21677 = ( n924 & ~n16407 ) | ( n924 & n18005 ) | ( ~n16407 & n18005 ) ;
  assign n21678 = n21676 & n21677 ;
  assign n21679 = ~n508 & n4061 ;
  assign n21680 = n11514 | n21679 ;
  assign n21681 = ~n6885 & n14066 ;
  assign n21682 = n2603 & ~n5981 ;
  assign n21683 = n21682 ^ n21189 ^ 1'b0 ;
  assign n21684 = n7045 | n21652 ;
  assign n21685 = n18199 & ~n21684 ;
  assign n21686 = n2284 & ~n6727 ;
  assign n21687 = n6727 & n21686 ;
  assign n21688 = n21687 ^ n14829 ^ 1'b0 ;
  assign n21689 = n21688 ^ n13480 ^ 1'b0 ;
  assign n21690 = n6060 & ~n21689 ;
  assign n21691 = n1414 & ~n3996 ;
  assign n21692 = n3996 & n21691 ;
  assign n21696 = n1726 & ~n3369 ;
  assign n21697 = ~n1726 & n21696 ;
  assign n21698 = ~n7273 & n21697 ;
  assign n21693 = n1256 & ~n1430 ;
  assign n21694 = ~n1256 & n21693 ;
  assign n21695 = n11214 & ~n21694 ;
  assign n21699 = n21698 ^ n21695 ^ 1'b0 ;
  assign n21700 = n4171 | n21699 ;
  assign n21701 = n21692 & ~n21700 ;
  assign n21702 = n18636 ^ n1261 ^ n376 ;
  assign n21703 = n20679 ^ n7062 ^ 1'b0 ;
  assign n21704 = n16871 & n21703 ;
  assign n21705 = n11815 ^ n5059 ^ 1'b0 ;
  assign n21706 = ~n10270 & n12897 ;
  assign n21707 = ~n20295 & n21706 ;
  assign n21708 = n1533 | n6465 ;
  assign n21709 = n7810 & ~n21708 ;
  assign n21710 = n19949 & ~n21709 ;
  assign n21711 = n21710 ^ n11106 ^ 1'b0 ;
  assign n21712 = n5269 ^ n2987 ^ n374 ;
  assign n21713 = ~n12784 & n14014 ;
  assign n21714 = ~n21712 & n21713 ;
  assign n21715 = n2980 | n7659 ;
  assign n21716 = n21714 & ~n21715 ;
  assign n21717 = n11172 ^ n8012 ^ n88 ;
  assign n21718 = n21717 ^ n12908 ^ 1'b0 ;
  assign n21719 = n21718 ^ n17720 ^ 1'b0 ;
  assign n21722 = n4940 & ~n7362 ;
  assign n21723 = ~n16703 & n21722 ;
  assign n21724 = n387 & ~n21723 ;
  assign n21720 = n15200 & n15488 ;
  assign n21721 = n343 | n21720 ;
  assign n21725 = n21724 ^ n21721 ^ 1'b0 ;
  assign n21726 = n415 | n7287 ;
  assign n21727 = n13934 & ~n21726 ;
  assign n21728 = n16978 ^ n5979 ^ 1'b0 ;
  assign n21729 = n15283 & ~n21728 ;
  assign n21730 = n5078 & n21729 ;
  assign n21731 = n6664 & n18317 ;
  assign n21732 = n7579 | n9812 ;
  assign n21733 = n16089 & ~n21732 ;
  assign n21734 = n15062 | n21733 ;
  assign n21735 = n5675 | n21734 ;
  assign n21736 = n1852 | n2066 ;
  assign n21737 = n21736 ^ n14082 ^ 1'b0 ;
  assign n21738 = n14362 | n21737 ;
  assign n21739 = n7877 | n14895 ;
  assign n21740 = n12757 & n16234 ;
  assign n21741 = ~n4639 & n21740 ;
  assign n21742 = n21741 ^ n20002 ^ 1'b0 ;
  assign n21743 = n21739 | n21742 ;
  assign n21744 = n7818 | n16891 ;
  assign n21745 = n20367 ^ n14152 ^ 1'b0 ;
  assign n21746 = n14760 | n21745 ;
  assign n21747 = ~n13157 & n13640 ;
  assign n21748 = n7128 ^ n2915 ^ 1'b0 ;
  assign n21749 = n21748 ^ n733 ^ 1'b0 ;
  assign n21752 = n506 | n3507 ;
  assign n21753 = n506 & ~n21752 ;
  assign n21754 = n16277 | n21753 ;
  assign n21755 = n16277 & ~n21754 ;
  assign n21756 = n21755 ^ n17051 ^ 1'b0 ;
  assign n21750 = n1389 | n6166 ;
  assign n21751 = n21750 ^ n9720 ^ 1'b0 ;
  assign n21757 = n21756 ^ n21751 ^ n17696 ;
  assign n21758 = ~n9477 & n18811 ;
  assign n21759 = n16094 ^ n1816 ^ 1'b0 ;
  assign n21760 = n4657 & n21759 ;
  assign n21761 = n4317 & n21760 ;
  assign n21763 = n9254 | n10890 ;
  assign n21764 = n21763 ^ n758 ^ 1'b0 ;
  assign n21762 = n663 | n10274 ;
  assign n21765 = n21764 ^ n21762 ^ 1'b0 ;
  assign n21766 = n6092 & ~n6931 ;
  assign n21767 = n8258 & n21766 ;
  assign n21768 = ~n1622 & n9685 ;
  assign n21769 = ~n9674 & n21768 ;
  assign n21770 = ~n19245 & n21769 ;
  assign n21771 = ~n21767 & n21770 ;
  assign n21772 = ~n21765 & n21771 ;
  assign n21773 = ~n1566 & n1726 ;
  assign n21774 = n21773 ^ n9002 ^ n7570 ;
  assign n21775 = n2812 | n21774 ;
  assign n21776 = n21775 ^ n16629 ^ n12559 ;
  assign n21777 = n21776 ^ n4048 ^ 1'b0 ;
  assign n21778 = ( n3776 & n11504 ) | ( n3776 & ~n16780 ) | ( n11504 & ~n16780 ) ;
  assign n21779 = n4298 | n11630 ;
  assign n21780 = ~n16790 & n20366 ;
  assign n21781 = n3572 & n8721 ;
  assign n21782 = n16982 ^ n15103 ^ n831 ;
  assign n21783 = ~n8355 & n8366 ;
  assign n21784 = n21783 ^ n2045 ^ 1'b0 ;
  assign n21785 = n15819 ^ n11442 ^ 1'b0 ;
  assign n21786 = n21784 | n21785 ;
  assign n21787 = n9883 | n21786 ;
  assign n21788 = n21787 ^ n17677 ^ 1'b0 ;
  assign n21789 = n8057 | n21788 ;
  assign n21790 = n8514 ^ n1460 ^ 1'b0 ;
  assign n21791 = n2024 & n21790 ;
  assign n21792 = n15565 & n17224 ;
  assign n21793 = ~n5495 & n21792 ;
  assign n21794 = n7965 & n21793 ;
  assign n21795 = ( n3715 & n3911 ) | ( n3715 & n7007 ) | ( n3911 & n7007 ) ;
  assign n21796 = n21795 ^ n8893 ^ 1'b0 ;
  assign n21797 = ~n5704 & n21796 ;
  assign n21798 = ~n4364 & n14052 ;
  assign n21799 = ~n3412 & n5147 ;
  assign n21800 = n2987 & n21799 ;
  assign n21801 = n20065 ^ n4489 ^ 1'b0 ;
  assign n21802 = n11678 ^ n6989 ^ 1'b0 ;
  assign n21803 = n15207 ^ n11880 ^ 1'b0 ;
  assign n21804 = ~n7881 & n21803 ;
  assign n21805 = n19681 ^ n1075 ^ n931 ;
  assign n21806 = n11355 & n21681 ;
  assign n21807 = ~n4671 & n18416 ;
  assign n21808 = n1812 & n21807 ;
  assign n21809 = n13040 & ~n21808 ;
  assign n21810 = ~n10209 & n18576 ;
  assign n21811 = n83 | n13152 ;
  assign n21812 = n21810 & ~n21811 ;
  assign n21813 = ~n3299 & n7048 ;
  assign n21814 = n21813 ^ n8328 ^ 1'b0 ;
  assign n21815 = n6469 | n6919 ;
  assign n21816 = n8553 | n21815 ;
  assign n21817 = n21814 & n21816 ;
  assign n21818 = n21817 ^ n4149 ^ 1'b0 ;
  assign n21819 = n9624 | n16336 ;
  assign n21820 = n1853 & ~n3442 ;
  assign n21821 = n2460 & ~n11838 ;
  assign n21822 = ~n2647 & n20520 ;
  assign n21823 = n3638 ^ n1327 ^ 1'b0 ;
  assign n21824 = n21823 ^ n1695 ^ 1'b0 ;
  assign n21825 = n11274 & ~n21824 ;
  assign n21826 = n21779 ^ n21581 ^ 1'b0 ;
  assign n21827 = n12142 ^ n10314 ^ 1'b0 ;
  assign n21828 = ~n1081 & n21827 ;
  assign n21829 = n619 & n21828 ;
  assign n21830 = n3443 & n21829 ;
  assign n21831 = n7602 ^ n3876 ^ 1'b0 ;
  assign n21832 = n5880 ^ n2641 ^ 1'b0 ;
  assign n21833 = n21831 | n21832 ;
  assign n21834 = ~n21621 & n21833 ;
  assign n21842 = n16131 ^ n9241 ^ 1'b0 ;
  assign n21843 = n2120 | n21842 ;
  assign n21838 = n4681 ^ n69 ^ 1'b0 ;
  assign n21839 = n21838 ^ n6984 ^ n1052 ;
  assign n21835 = n12379 ^ n9652 ^ 1'b0 ;
  assign n21836 = n21611 ^ n3102 ^ 1'b0 ;
  assign n21837 = ~n21835 & n21836 ;
  assign n21840 = n21839 ^ n21837 ^ 1'b0 ;
  assign n21841 = ~n3004 & n21840 ;
  assign n21844 = n21843 ^ n21841 ^ 1'b0 ;
  assign n21845 = n631 & n8655 ;
  assign n21846 = ( n3605 & ~n12168 ) | ( n3605 & n21845 ) | ( ~n12168 & n21845 ) ;
  assign n21847 = n3160 & n6274 ;
  assign n21848 = n6235 | n21847 ;
  assign n21849 = n1564 & ~n14749 ;
  assign n21850 = ~n1688 & n21849 ;
  assign n21851 = n5229 | n21221 ;
  assign n21852 = n21850 | n21851 ;
  assign n21853 = ~n7293 & n20030 ;
  assign n21854 = n10586 & ~n18418 ;
  assign n21855 = n21854 ^ n5744 ^ 1'b0 ;
  assign n21856 = n1118 & ~n4897 ;
  assign n21857 = n1199 & n21856 ;
  assign n21858 = n21857 ^ n13538 ^ n9189 ;
  assign n21859 = n7425 | n20453 ;
  assign n21860 = n21859 ^ n17270 ^ 1'b0 ;
  assign n21861 = n21858 | n21860 ;
  assign n21862 = n16884 ^ n4201 ^ 1'b0 ;
  assign n21863 = n4254 & n21862 ;
  assign n21864 = n5037 ^ n4690 ^ 1'b0 ;
  assign n21865 = n21863 & ~n21864 ;
  assign n21866 = n21865 ^ n9709 ^ 1'b0 ;
  assign n21867 = n9570 | n21866 ;
  assign n21868 = n6528 & ~n21867 ;
  assign n21869 = n11430 & n21868 ;
  assign n21870 = n3626 & ~n6417 ;
  assign n21871 = ~n4004 & n21870 ;
  assign n21872 = ~n2309 & n21871 ;
  assign n21873 = ~n5744 & n12893 ;
  assign n21874 = n21873 ^ n1747 ^ 1'b0 ;
  assign n21875 = ( ~n2287 & n5469 ) | ( ~n2287 & n17162 ) | ( n5469 & n17162 ) ;
  assign n21876 = n5489 & ~n18503 ;
  assign n21877 = ~n21348 & n21876 ;
  assign n21878 = n10607 & n21877 ;
  assign n21879 = n16479 ^ n4885 ^ 1'b0 ;
  assign n21880 = n21879 ^ n11887 ^ n2555 ;
  assign n21881 = n21880 ^ n10162 ^ 1'b0 ;
  assign n21882 = n7624 & n11159 ;
  assign n21883 = n4555 | n11664 ;
  assign n21884 = ( n1307 & n5412 ) | ( n1307 & ~n10052 ) | ( n5412 & ~n10052 ) ;
  assign n21885 = n14262 | n21884 ;
  assign n21886 = n15697 ^ n344 ^ 1'b0 ;
  assign n21887 = n835 & n2377 ;
  assign n21888 = n21887 ^ n9950 ^ 1'b0 ;
  assign n21889 = n21888 ^ n2351 ^ 1'b0 ;
  assign n21890 = n8009 ^ n1392 ^ 1'b0 ;
  assign n21891 = n6522 & n6764 ;
  assign n21892 = n21891 ^ n9063 ^ 1'b0 ;
  assign n21893 = n15556 ^ n11449 ^ 1'b0 ;
  assign n21894 = n1553 ^ n261 ^ 1'b0 ;
  assign n21895 = ~n5685 & n15605 ;
  assign n21896 = n21895 ^ n7843 ^ 1'b0 ;
  assign n21897 = n13205 ^ n7877 ^ n6866 ;
  assign n21898 = n15622 | n19818 ;
  assign n21899 = n17465 & ~n21898 ;
  assign n21900 = ( n13024 & n16581 ) | ( n13024 & ~n17725 ) | ( n16581 & ~n17725 ) ;
  assign n21903 = n1381 ^ n1094 ^ n266 ;
  assign n21904 = ~n6671 & n21903 ;
  assign n21901 = ~n4672 & n19688 ;
  assign n21902 = n21901 ^ n12078 ^ 1'b0 ;
  assign n21905 = n21904 ^ n21902 ^ n10039 ;
  assign n21906 = n6598 | n10929 ;
  assign n21907 = n21906 ^ n10795 ^ 1'b0 ;
  assign n21908 = n21907 ^ n2397 ^ 1'b0 ;
  assign n21909 = n8662 & n21908 ;
  assign n21910 = n9696 ^ n1269 ^ 1'b0 ;
  assign n21911 = ~n3923 & n21910 ;
  assign n21912 = n8792 ^ n5990 ^ 1'b0 ;
  assign n21913 = n16998 ^ n8960 ^ 1'b0 ;
  assign n21914 = n6626 ^ n6104 ^ 1'b0 ;
  assign n21915 = n5665 & n21914 ;
  assign n21916 = ~n10632 & n14744 ;
  assign n21917 = n8737 & ~n21916 ;
  assign n21918 = ~n21915 & n21917 ;
  assign n21919 = n2284 | n21918 ;
  assign n21920 = n545 & n5268 ;
  assign n21921 = ~n21919 & n21920 ;
  assign n21922 = n10047 | n21921 ;
  assign n21923 = n21922 ^ n5249 ^ 1'b0 ;
  assign n21927 = n1353 | n3549 ;
  assign n21928 = n21927 ^ n517 ^ 1'b0 ;
  assign n21929 = n21928 ^ n3849 ^ 1'b0 ;
  assign n21930 = ~n887 & n21929 ;
  assign n21924 = n8388 ^ n1637 ^ n1367 ;
  assign n21925 = n21924 ^ n12466 ^ 1'b0 ;
  assign n21926 = n898 & n21925 ;
  assign n21931 = n21930 ^ n21926 ^ n6841 ;
  assign n21932 = n2252 & n8070 ;
  assign n21936 = n8883 & ~n9354 ;
  assign n21933 = n1439 ^ n1344 ^ 1'b0 ;
  assign n21934 = n740 | n21933 ;
  assign n21935 = n21934 ^ n10656 ^ 1'b0 ;
  assign n21937 = n21936 ^ n21935 ^ 1'b0 ;
  assign n21938 = n67 | n21937 ;
  assign n21939 = ( n378 & ~n1772 ) | ( n378 & n6147 ) | ( ~n1772 & n6147 ) ;
  assign n21940 = n9908 & n21939 ;
  assign n21941 = n1563 | n5348 ;
  assign n21942 = n1540 & ~n6759 ;
  assign n21943 = n21942 ^ n9777 ^ 1'b0 ;
  assign n21944 = n21941 & ~n21943 ;
  assign n21945 = n4457 & n11058 ;
  assign n21946 = ~n3011 & n7856 ;
  assign n21947 = n21946 ^ n542 ^ 1'b0 ;
  assign n21948 = n15598 ^ n10956 ^ 1'b0 ;
  assign n21949 = n21947 & ~n21948 ;
  assign n21950 = ~n21945 & n21949 ;
  assign n21951 = n3352 ^ n2772 ^ 1'b0 ;
  assign n21952 = n11509 & n21951 ;
  assign n21953 = n4596 ^ n911 ^ 1'b0 ;
  assign n21954 = n9213 & ~n16048 ;
  assign n21955 = n21954 ^ n1391 ^ 1'b0 ;
  assign n21956 = ~n934 & n21955 ;
  assign n21957 = n13941 & ~n21956 ;
  assign n21958 = n21957 ^ n11252 ^ n4778 ;
  assign n21959 = n2813 & n14828 ;
  assign n21960 = n21958 & n21959 ;
  assign n21961 = n17083 ^ n7360 ^ 1'b0 ;
  assign n21962 = n21961 ^ n4369 ^ n2991 ;
  assign n21963 = n4422 | n4556 ;
  assign n21964 = n21963 ^ n920 ^ 1'b0 ;
  assign n21965 = n4405 | n16445 ;
  assign n21966 = n1111 | n5861 ;
  assign n21967 = n88 & ~n21966 ;
  assign n21968 = n727 | n21967 ;
  assign n21969 = n6184 & ~n21968 ;
  assign n21970 = ~n16387 & n17637 ;
  assign n21971 = n2671 & n17999 ;
  assign n21972 = ~n17999 & n21971 ;
  assign n21973 = n21972 ^ n7156 ^ 1'b0 ;
  assign n21974 = n4677 & ~n13617 ;
  assign n21975 = ~n4677 & n21974 ;
  assign n21976 = n5073 | n21975 ;
  assign n21977 = n5073 & ~n21976 ;
  assign n21978 = n21973 | n21977 ;
  assign n21979 = n21978 ^ n4051 ^ 1'b0 ;
  assign n21980 = ( n4939 & n13324 ) | ( n4939 & ~n21979 ) | ( n13324 & ~n21979 ) ;
  assign n21981 = n5749 ^ n5145 ^ 1'b0 ;
  assign n21982 = n21981 ^ n8454 ^ 1'b0 ;
  assign n21983 = n9689 | n11809 ;
  assign n21984 = n21982 & ~n21983 ;
  assign n21985 = n5990 & ~n20654 ;
  assign n21986 = n6408 ^ n5031 ^ 1'b0 ;
  assign n21987 = n2082 & ~n21986 ;
  assign n21988 = n530 & ~n7034 ;
  assign n21989 = n21988 ^ n11811 ^ 1'b0 ;
  assign n21990 = n1154 & n16299 ;
  assign n21991 = n11411 & n20829 ;
  assign n21992 = ~n936 & n21991 ;
  assign n21993 = n2912 & ~n21893 ;
  assign n21994 = n4753 & n12202 ;
  assign n21995 = n21994 ^ n1542 ^ 1'b0 ;
  assign n21996 = n12533 ^ n8061 ^ n492 ;
  assign n21997 = n3393 & ~n8891 ;
  assign n21998 = n4497 & n21997 ;
  assign n21999 = n15614 & ~n21998 ;
  assign n22000 = n21996 & n21999 ;
  assign n22001 = ~n695 & n18707 ;
  assign n22002 = n20299 ^ n11162 ^ 1'b0 ;
  assign n22003 = ~n2446 & n16720 ;
  assign n22004 = n15975 & n22003 ;
  assign n22005 = n10161 ^ n7835 ^ n1445 ;
  assign n22006 = n2314 & ~n2673 ;
  assign n22007 = n22005 & n22006 ;
  assign n22008 = n20290 | n22007 ;
  assign n22009 = n22008 ^ n5188 ^ 1'b0 ;
  assign n22010 = n3169 ^ n2852 ^ 1'b0 ;
  assign n22011 = n22010 ^ n1650 ^ 1'b0 ;
  assign n22012 = ~n2689 & n22011 ;
  assign n22013 = n45 & ~n3416 ;
  assign n22014 = n22012 & n22013 ;
  assign n22015 = ~n16782 & n22014 ;
  assign n22017 = n3758 ^ n115 ^ 1'b0 ;
  assign n22016 = n2145 & ~n2242 ;
  assign n22018 = n22017 ^ n22016 ^ 1'b0 ;
  assign n22019 = n12003 & ~n22018 ;
  assign n22020 = ~n15067 & n22019 ;
  assign n22021 = n8831 | n22020 ;
  assign n22022 = n20034 ^ n10012 ^ 1'b0 ;
  assign n22023 = n2004 & n22022 ;
  assign n22024 = n22023 ^ n86 ^ 1'b0 ;
  assign n22025 = ~n9184 & n22024 ;
  assign n22026 = ~n15511 & n22025 ;
  assign n22027 = n22026 ^ n3610 ^ 1'b0 ;
  assign n22028 = ~n20234 & n21175 ;
  assign n22029 = ( ~n513 & n535 ) | ( ~n513 & n5618 ) | ( n535 & n5618 ) ;
  assign n22030 = n14428 & ~n22029 ;
  assign n22031 = ~n4757 & n22030 ;
  assign n22032 = n3071 & n6732 ;
  assign n22033 = ~n1217 & n22032 ;
  assign n22034 = n13897 & ~n19552 ;
  assign n22035 = n11217 ^ n10834 ^ 1'b0 ;
  assign n22036 = n22035 ^ n20220 ^ 1'b0 ;
  assign n22037 = x11 & n16132 ;
  assign n22038 = n17408 ^ n16334 ^ 1'b0 ;
  assign n22039 = n16790 | n22038 ;
  assign n22040 = n6271 | n13684 ;
  assign n22041 = n1128 | n6543 ;
  assign n22043 = n8182 ^ n7784 ^ 1'b0 ;
  assign n22044 = n3756 & ~n22043 ;
  assign n22045 = n695 & n22044 ;
  assign n22046 = ~n10829 & n22045 ;
  assign n22042 = n4974 ^ n3270 ^ 1'b0 ;
  assign n22047 = n22046 ^ n22042 ^ n9202 ;
  assign n22048 = n4348 & n17221 ;
  assign n22049 = n667 | n1786 ;
  assign n22050 = n9502 | n22049 ;
  assign n22051 = n5856 ^ n1828 ^ 1'b0 ;
  assign n22052 = n8580 ^ n458 ^ 1'b0 ;
  assign n22053 = n7718 & n22052 ;
  assign n22054 = ~n2721 & n22053 ;
  assign n22059 = ( ~n1755 & n4335 ) | ( ~n1755 & n4832 ) | ( n4335 & n4832 ) ;
  assign n22060 = ~n15928 & n22059 ;
  assign n22055 = n2445 & ~n7526 ;
  assign n22056 = ~n10099 & n22055 ;
  assign n22057 = n8110 & ~n22056 ;
  assign n22058 = n9843 | n22057 ;
  assign n22061 = n22060 ^ n22058 ^ 1'b0 ;
  assign n22062 = ~n4438 & n22061 ;
  assign n22063 = n22062 ^ n12860 ^ 1'b0 ;
  assign n22067 = n5474 | n12529 ;
  assign n22064 = n1971 | n8815 ;
  assign n22065 = n22064 ^ n5810 ^ 1'b0 ;
  assign n22066 = n8460 | n22065 ;
  assign n22068 = n22067 ^ n22066 ^ 1'b0 ;
  assign n22069 = n11931 ^ n704 ^ 1'b0 ;
  assign n22070 = ~n4529 & n22069 ;
  assign n22071 = n384 | n1094 ;
  assign n22072 = n4182 ^ n2615 ^ 1'b0 ;
  assign n22073 = n489 & n22072 ;
  assign n22074 = n22073 ^ n6688 ^ 1'b0 ;
  assign n22075 = n22071 | n22074 ;
  assign n22076 = n11023 & ~n22075 ;
  assign n22077 = n22076 ^ n11620 ^ 1'b0 ;
  assign n22079 = n9657 | n13042 ;
  assign n22080 = n5632 & ~n22079 ;
  assign n22078 = n15098 & n16675 ;
  assign n22081 = n22080 ^ n22078 ^ 1'b0 ;
  assign n22082 = n10057 ^ n5132 ^ n3127 ;
  assign n22083 = ( n7527 & ~n11384 ) | ( n7527 & n22082 ) | ( ~n11384 & n22082 ) ;
  assign n22084 = n14573 ^ n1144 ^ 1'b0 ;
  assign n22085 = ~n3345 & n22084 ;
  assign n22086 = n22083 & n22085 ;
  assign n22087 = ( n9509 & ~n12233 ) | ( n9509 & n17975 ) | ( ~n12233 & n17975 ) ;
  assign n22088 = n19064 ^ n8043 ^ n5114 ;
  assign n22089 = n22088 ^ n4645 ^ 1'b0 ;
  assign n22090 = ~n22087 & n22089 ;
  assign n22091 = n18856 ^ n8773 ^ 1'b0 ;
  assign n22092 = ~n3950 & n5938 ;
  assign n22093 = n22092 ^ n15119 ^ 1'b0 ;
  assign n22094 = n1821 & n22093 ;
  assign n22095 = n8917 & ~n22094 ;
  assign n22096 = n4063 | n5747 ;
  assign n22097 = n849 | n22096 ;
  assign n22098 = ~n10543 & n12625 ;
  assign n22099 = n14957 ^ n5652 ^ n802 ;
  assign n22101 = n14509 ^ n9203 ^ 1'b0 ;
  assign n22100 = n7973 & ~n11397 ;
  assign n22102 = n22101 ^ n22100 ^ 1'b0 ;
  assign n22103 = n13147 ^ n8764 ^ n5863 ;
  assign n22104 = ~n10098 & n22103 ;
  assign n22105 = n22104 ^ n1868 ^ 1'b0 ;
  assign n22106 = ~n5226 & n21109 ;
  assign n22107 = n545 & ~n1410 ;
  assign n22108 = n22107 ^ n15582 ^ 1'b0 ;
  assign n22109 = n1657 | n10213 ;
  assign n22110 = n22109 ^ n20919 ^ 1'b0 ;
  assign n22112 = n1804 & ~n10300 ;
  assign n22113 = n2108 & ~n22112 ;
  assign n22111 = ~n9270 & n12659 ;
  assign n22114 = n22113 ^ n22111 ^ 1'b0 ;
  assign n22115 = n16945 ^ n3224 ^ 1'b0 ;
  assign n22116 = ~n8803 & n8885 ;
  assign n22117 = ~n7335 & n22116 ;
  assign n22118 = n7474 & ~n22117 ;
  assign n22119 = ~n19256 & n22118 ;
  assign n22120 = n1006 | n16838 ;
  assign n22121 = n7025 | n22120 ;
  assign n22122 = n19249 ^ n16284 ^ 1'b0 ;
  assign n22123 = n5047 | n22122 ;
  assign n22124 = n9254 ^ n4335 ^ 1'b0 ;
  assign n22125 = n2663 ^ n451 ^ 1'b0 ;
  assign n22126 = n22125 ^ n14714 ^ 1'b0 ;
  assign n22127 = ( n1714 & n11793 ) | ( n1714 & n22126 ) | ( n11793 & n22126 ) ;
  assign n22128 = n492 & n6398 ;
  assign n22130 = n7119 ^ n2324 ^ n459 ;
  assign n22131 = n22130 ^ n8041 ^ 1'b0 ;
  assign n22132 = n884 & n10230 ;
  assign n22133 = ~n22131 & n22132 ;
  assign n22129 = n10075 & ~n13205 ;
  assign n22134 = n22133 ^ n22129 ^ 1'b0 ;
  assign n22135 = n3626 | n10178 ;
  assign n22136 = n22135 ^ n13123 ^ 1'b0 ;
  assign n22137 = ~n10528 & n22136 ;
  assign n22138 = n22137 ^ n4676 ^ 1'b0 ;
  assign n22139 = n7444 ^ n1967 ^ 1'b0 ;
  assign n22140 = n14892 | n22139 ;
  assign n22141 = n18135 & ~n18589 ;
  assign n22142 = n1438 | n9311 ;
  assign n22143 = n21410 | n22142 ;
  assign n22144 = n19271 ^ n1098 ^ 1'b0 ;
  assign n22146 = n9016 ^ n6771 ^ n4675 ;
  assign n22145 = n3730 & n15519 ;
  assign n22147 = n22146 ^ n22145 ^ 1'b0 ;
  assign n22148 = n6278 & n22147 ;
  assign n22149 = n22148 ^ n5394 ^ 1'b0 ;
  assign n22150 = n4591 & n22149 ;
  assign n22151 = ~n19930 & n22150 ;
  assign n22152 = ~n1688 & n22151 ;
  assign n22153 = ~n805 & n11166 ;
  assign n22154 = n16144 & ~n16502 ;
  assign n22155 = n22153 & n22154 ;
  assign n22156 = n22155 ^ n9020 ^ 1'b0 ;
  assign n22157 = n7234 ^ n1539 ^ 1'b0 ;
  assign n22158 = n7099 ^ n205 ^ 1'b0 ;
  assign n22159 = n22158 ^ n1588 ^ 1'b0 ;
  assign n22160 = ~n10092 & n22159 ;
  assign n22161 = ~n4894 & n22160 ;
  assign n22162 = ~n13380 & n22161 ;
  assign n22163 = ~n22157 & n22162 ;
  assign n22171 = n2787 ^ n1422 ^ 1'b0 ;
  assign n22172 = n11995 & ~n22171 ;
  assign n22173 = n2486 & n22172 ;
  assign n22170 = n91 & ~n5377 ;
  assign n22174 = n22173 ^ n22170 ^ 1'b0 ;
  assign n22164 = n3618 | n4285 ;
  assign n22165 = n22164 ^ n6080 ^ 1'b0 ;
  assign n22166 = n8559 | n22165 ;
  assign n22167 = n22166 ^ n10241 ^ 1'b0 ;
  assign n22168 = n2935 | n22167 ;
  assign n22169 = n5874 | n22168 ;
  assign n22175 = n22174 ^ n22169 ^ 1'b0 ;
  assign n22176 = n1882 & n3580 ;
  assign n22177 = ~n4264 & n22176 ;
  assign n22178 = n22177 ^ n8322 ^ 1'b0 ;
  assign n22179 = ~n17345 & n22178 ;
  assign n22180 = n7836 ^ n5395 ^ 1'b0 ;
  assign n22181 = ( x6 & ~n12593 ) | ( x6 & n16903 ) | ( ~n12593 & n16903 ) ;
  assign n22182 = n4660 | n20667 ;
  assign n22183 = n15550 ^ n382 ^ 1'b0 ;
  assign n22184 = n21092 ^ n88 ^ 1'b0 ;
  assign n22185 = n1223 | n7448 ;
  assign n22186 = n22185 ^ n4340 ^ 1'b0 ;
  assign n22187 = ~n12307 & n22186 ;
  assign n22188 = n15372 ^ n11948 ^ n7645 ;
  assign n22189 = n22188 ^ n6841 ^ 1'b0 ;
  assign n22190 = n3924 & ~n12637 ;
  assign n22191 = n4432 ^ n328 ^ 1'b0 ;
  assign n22192 = n6966 & n22191 ;
  assign n22193 = n7597 | n22192 ;
  assign n22194 = n22193 ^ n21621 ^ n14575 ;
  assign n22195 = ~n1083 & n5417 ;
  assign n22196 = n1083 & n22195 ;
  assign n22197 = ~n7752 & n22196 ;
  assign n22198 = n18312 & n22197 ;
  assign n22199 = n15896 & n22198 ;
  assign n22200 = n2440 & n8863 ;
  assign n22201 = n22200 ^ n5574 ^ 1'b0 ;
  assign n22202 = ( n6333 & n7655 ) | ( n6333 & ~n22201 ) | ( n7655 & ~n22201 ) ;
  assign n22203 = n5992 ^ n1454 ^ 1'b0 ;
  assign n22204 = ~n12891 & n22203 ;
  assign n22205 = ~n5950 & n8365 ;
  assign n22206 = n10956 ^ n9444 ^ 1'b0 ;
  assign n22207 = n17766 ^ n749 ^ 1'b0 ;
  assign n22208 = n5445 ^ n3129 ^ 1'b0 ;
  assign n22209 = n12260 & ~n22208 ;
  assign n22210 = n22209 ^ n1821 ^ 1'b0 ;
  assign n22211 = ~n10171 & n22210 ;
  assign n22212 = x11 | n9250 ;
  assign n22213 = n4173 ^ n3444 ^ 1'b0 ;
  assign n22214 = n19821 & n22213 ;
  assign n22215 = n22214 ^ n14656 ^ 1'b0 ;
  assign n22216 = ~n5831 & n22215 ;
  assign n22217 = n13495 ^ n150 ^ 1'b0 ;
  assign n22218 = n552 & ~n20496 ;
  assign n22219 = ~n15898 & n22218 ;
  assign n22220 = n4960 & n22219 ;
  assign n22221 = n22217 & ~n22220 ;
  assign n22222 = n10342 ^ n8944 ^ 1'b0 ;
  assign n22223 = n9155 ^ n5680 ^ 1'b0 ;
  assign n22224 = n183 | n22223 ;
  assign n22225 = n1548 | n22224 ;
  assign n22226 = n22222 | n22225 ;
  assign n22227 = n22226 ^ n6442 ^ 1'b0 ;
  assign n22228 = n22221 | n22227 ;
  assign n22229 = n6481 & n17566 ;
  assign n22230 = n22228 & n22229 ;
  assign n22231 = n15109 ^ n1251 ^ 1'b0 ;
  assign n22232 = n11854 ^ n571 ^ 1'b0 ;
  assign n22233 = n22231 | n22232 ;
  assign n22234 = n20127 ^ n8322 ^ 1'b0 ;
  assign n22235 = n10771 & ~n22234 ;
  assign n22236 = ~n848 & n2236 ;
  assign n22237 = n12231 | n12994 ;
  assign n22238 = n6831 ^ n1483 ^ 1'b0 ;
  assign n22239 = ~n6914 & n22238 ;
  assign n22240 = n22239 ^ n11801 ^ 1'b0 ;
  assign n22241 = ~n1594 & n4733 ;
  assign n22242 = ~n10217 & n22241 ;
  assign n22243 = n17128 & n22242 ;
  assign n22244 = ~n1663 & n13318 ;
  assign n22245 = n22244 ^ n16318 ^ 1'b0 ;
  assign n22246 = ~n9585 & n22245 ;
  assign n22247 = ~n1369 & n22246 ;
  assign n22248 = n22247 ^ n9436 ^ 1'b0 ;
  assign n22249 = n11477 & ~n17784 ;
  assign n22250 = ~n1327 & n2975 ;
  assign n22251 = n13571 ^ n4113 ^ 1'b0 ;
  assign n22252 = n8756 ^ n452 ^ 1'b0 ;
  assign n22253 = n20617 | n22252 ;
  assign n22254 = n22251 | n22253 ;
  assign n22255 = n9864 & n9964 ;
  assign n22256 = n22255 ^ n2095 ^ 1'b0 ;
  assign n22257 = n9684 & ~n14932 ;
  assign n22258 = n6000 & n7297 ;
  assign n22259 = n22257 & n22258 ;
  assign n22260 = ~n5352 & n11318 ;
  assign n22261 = n14387 ^ n6864 ^ 1'b0 ;
  assign n22262 = n7480 | n9966 ;
  assign n22263 = ~n12134 & n22262 ;
  assign n22264 = n22263 ^ n4748 ^ 1'b0 ;
  assign n22265 = n8595 & n22264 ;
  assign n22266 = ~n16793 & n16971 ;
  assign n22267 = n11964 ^ n2195 ^ 1'b0 ;
  assign n22268 = n16028 ^ n11538 ^ 1'b0 ;
  assign n22269 = ( n630 & n14685 ) | ( n630 & ~n22268 ) | ( n14685 & ~n22268 ) ;
  assign n22270 = n4685 & ~n7062 ;
  assign n22271 = n5302 & n22270 ;
  assign n22272 = n9196 ^ n5555 ^ 1'b0 ;
  assign n22273 = n22272 ^ n12897 ^ 1'b0 ;
  assign n22274 = n1282 & n22273 ;
  assign n22275 = n4595 | n22218 ;
  assign n22276 = n22275 ^ n8549 ^ 1'b0 ;
  assign n22277 = ~n22274 & n22276 ;
  assign n22278 = n10084 & ~n19818 ;
  assign n22279 = n16364 ^ n11968 ^ n9899 ;
  assign n22280 = ~n668 & n2029 ;
  assign n22281 = n6454 & n22280 ;
  assign n22282 = ~n2395 & n10393 ;
  assign n22283 = n749 & n22282 ;
  assign n22284 = n22283 ^ n14768 ^ n302 ;
  assign n22285 = n18975 ^ n14369 ^ n19 ;
  assign n22286 = n11442 ^ n5329 ^ n2049 ;
  assign n22287 = n22286 ^ n5382 ^ 1'b0 ;
  assign n22288 = n1095 | n22287 ;
  assign n22289 = n19767 | n22288 ;
  assign n22290 = n7917 | n22158 ;
  assign n22291 = n22289 & ~n22290 ;
  assign n22292 = n1490 & ~n3674 ;
  assign n22293 = ( n5564 & n10366 ) | ( n5564 & n22292 ) | ( n10366 & n22292 ) ;
  assign n22294 = n2668 & n22293 ;
  assign n22295 = n22294 ^ n7734 ^ 1'b0 ;
  assign n22296 = n22295 ^ n758 ^ 1'b0 ;
  assign n22297 = n11936 ^ n4409 ^ n3699 ;
  assign n22298 = ~n22296 & n22297 ;
  assign n22299 = n22298 ^ n14091 ^ 1'b0 ;
  assign n22300 = ~n2787 & n7918 ;
  assign n22301 = n4694 | n15091 ;
  assign n22302 = n22300 | n22301 ;
  assign n22303 = ( n11409 & ~n13685 ) | ( n11409 & n20048 ) | ( ~n13685 & n20048 ) ;
  assign n22304 = ~n1783 & n11327 ;
  assign n22305 = n22304 ^ n9687 ^ 1'b0 ;
  assign n22306 = n555 & ~n4439 ;
  assign n22307 = n2110 | n12732 ;
  assign n22308 = n22306 & ~n22307 ;
  assign n22309 = n6979 & ~n22308 ;
  assign n22310 = n22309 ^ n3262 ^ 1'b0 ;
  assign n22311 = n7358 ^ n5001 ^ n2761 ;
  assign n22312 = n22311 ^ n12185 ^ 1'b0 ;
  assign n22313 = n17449 ^ n7739 ^ n149 ;
  assign n22314 = ( n7469 & n9694 ) | ( n7469 & n15459 ) | ( n9694 & n15459 ) ;
  assign n22315 = n16576 & ~n22314 ;
  assign n22316 = n22313 & n22315 ;
  assign n22317 = ~n1858 & n1984 ;
  assign n22318 = n22317 ^ n16150 ^ 1'b0 ;
  assign n22319 = n11458 & n16857 ;
  assign n22320 = n1040 | n16719 ;
  assign n22321 = n22320 ^ n5514 ^ 1'b0 ;
  assign n22322 = n15023 & ~n19534 ;
  assign n22323 = n22322 ^ n18024 ^ 1'b0 ;
  assign n22324 = ~n2181 & n3178 ;
  assign n22325 = n11577 & n22324 ;
  assign n22326 = ( ~n917 & n9391 ) | ( ~n917 & n22325 ) | ( n9391 & n22325 ) ;
  assign n22327 = n22326 ^ n9559 ^ 1'b0 ;
  assign n22328 = n4080 | n22327 ;
  assign n22329 = n11230 | n13110 ;
  assign n22330 = n17799 | n22329 ;
  assign n22331 = n740 | n881 ;
  assign n22332 = n21912 & ~n22331 ;
  assign n22333 = n22332 ^ n5831 ^ n2527 ;
  assign n22334 = n22333 ^ n18167 ^ 1'b0 ;
  assign n22335 = n22330 & n22334 ;
  assign n22336 = n19060 ^ n13337 ^ 1'b0 ;
  assign n22337 = n5314 & n22336 ;
  assign n22338 = n22337 ^ n6069 ^ 1'b0 ;
  assign n22341 = n9580 & ~n16823 ;
  assign n22339 = n10218 ^ n4952 ^ 1'b0 ;
  assign n22340 = n9117 & n22339 ;
  assign n22342 = n22341 ^ n22340 ^ 1'b0 ;
  assign n22343 = n14046 ^ n1828 ^ 1'b0 ;
  assign n22344 = n9455 ^ n1265 ^ 1'b0 ;
  assign n22345 = n22344 ^ n11995 ^ 1'b0 ;
  assign n22346 = n362 & ~n5508 ;
  assign n22347 = ~n10191 & n22346 ;
  assign n22348 = n6589 | n22347 ;
  assign n22349 = n10945 | n22348 ;
  assign n22350 = n22345 & n22349 ;
  assign n22351 = n6593 | n21305 ;
  assign n22353 = ( n2850 & n3056 ) | ( n2850 & n9224 ) | ( n3056 & n9224 ) ;
  assign n22352 = ~n5149 & n11690 ;
  assign n22354 = n22353 ^ n22352 ^ 1'b0 ;
  assign n22356 = n1370 & ~n4287 ;
  assign n22355 = n15487 | n15512 ;
  assign n22357 = n22356 ^ n22355 ^ 1'b0 ;
  assign n22358 = n2206 & n12550 ;
  assign n22359 = n8023 & n13477 ;
  assign n22360 = n22359 ^ n7001 ^ 1'b0 ;
  assign n22361 = n2968 & n4006 ;
  assign n22362 = n22361 ^ n9848 ^ 1'b0 ;
  assign n22363 = n4423 & n13600 ;
  assign n22364 = n22363 ^ n7934 ^ 1'b0 ;
  assign n22365 = ~n11742 & n22364 ;
  assign n22366 = n22365 ^ n9698 ^ 1'b0 ;
  assign n22367 = n7572 ^ n7342 ^ 1'b0 ;
  assign n22368 = n1293 | n22367 ;
  assign n22369 = n22368 ^ n20050 ^ 1'b0 ;
  assign n22370 = n14589 | n22369 ;
  assign n22371 = ( n224 & n20810 ) | ( n224 & ~n22370 ) | ( n20810 & ~n22370 ) ;
  assign n22372 = n22371 ^ n9391 ^ 1'b0 ;
  assign n22373 = n8487 & ~n9360 ;
  assign n22374 = n4087 & ~n22373 ;
  assign n22375 = n508 | n5700 ;
  assign n22376 = n7357 | n22375 ;
  assign n22377 = n6267 & n22376 ;
  assign n22378 = n311 | n2604 ;
  assign n22379 = n22378 ^ n13342 ^ 1'b0 ;
  assign n22380 = n22379 ^ n649 ^ 1'b0 ;
  assign n22381 = ~n9779 & n22380 ;
  assign n22388 = ~n1109 & n4407 ;
  assign n22389 = n22388 ^ n1372 ^ 1'b0 ;
  assign n22390 = ~n6633 & n22389 ;
  assign n22391 = ~n2628 & n22390 ;
  assign n22392 = ~n15023 & n22391 ;
  assign n22382 = ( ~n2631 & n7076 ) | ( ~n2631 & n11751 ) | ( n7076 & n11751 ) ;
  assign n22383 = n1276 & n4311 ;
  assign n22384 = n22383 ^ n2584 ^ 1'b0 ;
  assign n22385 = n6762 & n22384 ;
  assign n22386 = n22385 ^ n2202 ^ 1'b0 ;
  assign n22387 = n22382 | n22386 ;
  assign n22393 = n22392 ^ n22387 ^ 1'b0 ;
  assign n22394 = n14032 ^ n10449 ^ 1'b0 ;
  assign n22395 = ~n7128 & n9523 ;
  assign n22396 = n17305 ^ n3417 ^ 1'b0 ;
  assign n22397 = ( n425 & ~n5453 ) | ( n425 & n22396 ) | ( ~n5453 & n22396 ) ;
  assign n22398 = n19389 ^ n1050 ^ 1'b0 ;
  assign n22399 = n261 ^ n140 ^ 1'b0 ;
  assign n22400 = n3600 & n22399 ;
  assign n22401 = n22400 ^ n7924 ^ 1'b0 ;
  assign n22402 = n3762 & n6856 ;
  assign n22403 = ~n6856 & n22402 ;
  assign n22404 = ~n515 & n22403 ;
  assign n22405 = n22404 ^ n8003 ^ 1'b0 ;
  assign n22406 = n20408 ^ n7953 ^ 1'b0 ;
  assign n22407 = n1130 & ~n11964 ;
  assign n22408 = n3726 & n22407 ;
  assign n22409 = n22408 ^ n12163 ^ 1'b0 ;
  assign n22410 = n14068 & n16132 ;
  assign n22411 = ~n21046 & n22410 ;
  assign n22412 = n901 & ~n5448 ;
  assign n22413 = ~n7583 & n13547 ;
  assign n22414 = n5364 ^ n3800 ^ 1'b0 ;
  assign n22415 = ~n12789 & n22414 ;
  assign n22416 = n9860 & ~n14159 ;
  assign n22417 = n2656 & n4251 ;
  assign n22418 = n7721 | n21611 ;
  assign n22419 = n15737 & ~n22418 ;
  assign n22420 = n16528 & n22419 ;
  assign n22421 = n8967 ^ n3514 ^ 1'b0 ;
  assign n22422 = n22421 ^ n11904 ^ 1'b0 ;
  assign n22423 = n9574 | n22422 ;
  assign n22424 = n22423 ^ n11927 ^ 1'b0 ;
  assign n22425 = ~n9648 & n10251 ;
  assign n22426 = n2181 | n17538 ;
  assign n22427 = n22426 ^ n4707 ^ 1'b0 ;
  assign n22428 = n22427 ^ n10904 ^ n3330 ;
  assign n22429 = n13899 | n22428 ;
  assign n22430 = n22425 & ~n22429 ;
  assign n22431 = n5880 ^ n1434 ^ 1'b0 ;
  assign n22432 = ~n9270 & n10300 ;
  assign n22433 = n22432 ^ n150 ^ 1'b0 ;
  assign n22434 = n3962 & ~n16359 ;
  assign n22435 = ~n5662 & n22434 ;
  assign n22436 = n1221 | n6736 ;
  assign n22437 = n22436 ^ n20920 ^ 1'b0 ;
  assign n22438 = ~n15306 & n22437 ;
  assign n22439 = n1327 & n6839 ;
  assign n22440 = n22439 ^ n9550 ^ 1'b0 ;
  assign n22441 = n8750 | n22440 ;
  assign n22442 = n6081 | n22441 ;
  assign n22443 = n22442 ^ n5668 ^ n1064 ;
  assign n22444 = ~n17352 & n22443 ;
  assign n22445 = ~n22438 & n22444 ;
  assign n22446 = n22435 | n22445 ;
  assign n22447 = n10603 | n22446 ;
  assign n22448 = ~n3313 & n6984 ;
  assign n22449 = ~n9631 & n22448 ;
  assign n22450 = n3027 & n22449 ;
  assign n22451 = ~n7741 & n8186 ;
  assign n22452 = n9121 & ~n9724 ;
  assign n22453 = ~n7140 & n22452 ;
  assign n22454 = n7492 & n16425 ;
  assign n22455 = n13566 & n22454 ;
  assign n22456 = n22455 ^ n13503 ^ 1'b0 ;
  assign n22462 = n5965 & n8844 ;
  assign n22463 = n22462 ^ n5897 ^ 1'b0 ;
  assign n22459 = n14523 ^ n10963 ^ 1'b0 ;
  assign n22460 = ~n8884 & n22459 ;
  assign n22458 = ~n20136 & n21564 ;
  assign n22461 = n22460 ^ n22458 ^ 1'b0 ;
  assign n22464 = n22463 ^ n22461 ^ 1'b0 ;
  assign n22457 = n2962 & ~n4776 ;
  assign n22465 = n22464 ^ n22457 ^ 1'b0 ;
  assign n22466 = n11837 ^ n1531 ^ 1'b0 ;
  assign n22467 = n3449 ^ n695 ^ 1'b0 ;
  assign n22468 = n22467 ^ n7199 ^ 1'b0 ;
  assign n22469 = n5695 | n22468 ;
  assign n22470 = n9583 | n22469 ;
  assign n22471 = n22470 ^ n4121 ^ 1'b0 ;
  assign n22472 = n4169 ^ n1598 ^ 1'b0 ;
  assign n22473 = ~n3386 & n22472 ;
  assign n22474 = n2138 & n22473 ;
  assign n22475 = ~n2812 & n20653 ;
  assign n22476 = n18897 & n22475 ;
  assign n22477 = ~n959 & n4136 ;
  assign n22478 = n22477 ^ n5375 ^ 1'b0 ;
  assign n22479 = n1551 ^ n676 ^ 1'b0 ;
  assign n22480 = n5293 | n22479 ;
  assign n22481 = n22480 ^ n4945 ^ 1'b0 ;
  assign n22482 = n8147 & n22481 ;
  assign n22483 = n1620 & n1744 ;
  assign n22484 = ~n3315 & n22483 ;
  assign n22485 = n10601 ^ n3820 ^ 1'b0 ;
  assign n22486 = n12056 & ~n22485 ;
  assign n22487 = n1516 & n9873 ;
  assign n22488 = n8368 & n22487 ;
  assign n22491 = n1551 & n15137 ;
  assign n22492 = n22491 ^ n10610 ^ 1'b0 ;
  assign n22493 = n20625 ^ n2324 ^ 1'b0 ;
  assign n22494 = n22492 & ~n22493 ;
  assign n22489 = n4698 | n7664 ;
  assign n22490 = ~n19540 & n22489 ;
  assign n22495 = n22494 ^ n22490 ^ 1'b0 ;
  assign n22496 = ~n4512 & n21121 ;
  assign n22497 = n22496 ^ n372 ^ 1'b0 ;
  assign n22498 = n6672 | n11887 ;
  assign n22499 = n22498 ^ n588 ^ 1'b0 ;
  assign n22500 = n2048 | n17170 ;
  assign n22501 = n22499 & ~n22500 ;
  assign n22502 = n2029 & ~n16286 ;
  assign n22503 = ~n11834 & n22502 ;
  assign n22504 = n22503 ^ x11 ^ 1'b0 ;
  assign n22505 = n1340 & n11480 ;
  assign n22506 = ~n266 & n22505 ;
  assign n22507 = ~n884 & n3280 ;
  assign n22508 = n22506 | n22507 ;
  assign n22509 = n12602 | n22508 ;
  assign n22510 = ~n16010 & n19026 ;
  assign n22511 = n22510 ^ n16720 ^ 1'b0 ;
  assign n22512 = n3078 | n4685 ;
  assign n22513 = n22512 ^ n6185 ^ 1'b0 ;
  assign n22514 = n17 & ~n22513 ;
  assign n22515 = n13345 ^ n9929 ^ 1'b0 ;
  assign n22516 = n14353 ^ n13877 ^ n6613 ;
  assign n22517 = n18421 ^ n10782 ^ 1'b0 ;
  assign n22518 = ~n4543 & n11360 ;
  assign n22519 = n1426 & n22518 ;
  assign n22520 = ( n69 & ~n15597 ) | ( n69 & n22519 ) | ( ~n15597 & n22519 ) ;
  assign n22521 = n8825 & ~n22520 ;
  assign n22522 = ~n16144 & n22521 ;
  assign n22523 = n18100 ^ n6699 ^ n6161 ;
  assign n22524 = n13462 ^ n7865 ^ 1'b0 ;
  assign n22525 = n22524 ^ n20340 ^ n14580 ;
  assign n22526 = ~n5393 & n7665 ;
  assign n22527 = n14938 | n22526 ;
  assign n22528 = n22527 ^ n6206 ^ 1'b0 ;
  assign n22529 = n1686 | n22528 ;
  assign n22530 = n22529 ^ n1505 ^ 1'b0 ;
  assign n22531 = n160 & ~n20835 ;
  assign n22532 = n1275 & ~n19566 ;
  assign n22533 = ~n22531 & n22532 ;
  assign n22534 = n4132 & n20344 ;
  assign n22535 = ( n4452 & n10953 ) | ( n4452 & n22534 ) | ( n10953 & n22534 ) ;
  assign n22536 = n16020 ^ n15473 ^ 1'b0 ;
  assign n22537 = n9754 & ~n22536 ;
  assign n22538 = n6195 ^ n3813 ^ 1'b0 ;
  assign n22539 = n15590 & ~n22538 ;
  assign n22540 = n2455 & n22539 ;
  assign n22541 = n5775 ^ n3017 ^ 1'b0 ;
  assign n22542 = n13219 & ~n21399 ;
  assign n22543 = n22541 & n22542 ;
  assign n22544 = ~n6759 & n7236 ;
  assign n22545 = n22544 ^ n9770 ^ 1'b0 ;
  assign n22546 = n16464 & ~n22545 ;
  assign n22547 = n22546 ^ n20082 ^ 1'b0 ;
  assign n22548 = ~n9593 & n15045 ;
  assign n22549 = n22548 ^ n14364 ^ n4102 ;
  assign n22550 = n2343 & n3220 ;
  assign n22551 = n2922 & ~n22550 ;
  assign n22552 = n22551 ^ n15863 ^ 1'b0 ;
  assign n22553 = n22552 ^ n13201 ^ 1'b0 ;
  assign n22554 = ~n2872 & n3621 ;
  assign n22555 = n22554 ^ n7130 ^ 1'b0 ;
  assign n22556 = n22555 ^ n8291 ^ 1'b0 ;
  assign n22557 = n1615 & n22556 ;
  assign n22558 = n3414 & n22557 ;
  assign n22559 = n4951 & ~n22558 ;
  assign n22560 = n2605 & n22559 ;
  assign n22562 = n2346 & ~n16340 ;
  assign n22563 = n8392 & n22562 ;
  assign n22561 = n3558 | n6865 ;
  assign n22564 = n22563 ^ n22561 ^ 1'b0 ;
  assign n22566 = n5336 | n16751 ;
  assign n22567 = n13593 ^ n5797 ^ n1109 ;
  assign n22568 = n22566 | n22567 ;
  assign n22569 = n22568 ^ n841 ^ 1'b0 ;
  assign n22570 = n15062 | n22569 ;
  assign n22571 = n22570 ^ n11205 ^ 1'b0 ;
  assign n22565 = n18438 ^ n17363 ^ 1'b0 ;
  assign n22572 = n22571 ^ n22565 ^ n3395 ;
  assign n22573 = n1217 & ~n3574 ;
  assign n22574 = n4143 & n22573 ;
  assign n22575 = n22574 ^ n11533 ^ n609 ;
  assign n22576 = n5418 | n22575 ;
  assign n22577 = n6274 & ~n14450 ;
  assign n22578 = n13857 | n22577 ;
  assign n22579 = n7265 | n22578 ;
  assign n22580 = n4251 & ~n16393 ;
  assign n22581 = n2005 & ~n3017 ;
  assign n22582 = n11155 & n14126 ;
  assign n22583 = n22582 ^ n5353 ^ 1'b0 ;
  assign n22584 = n22581 & n22583 ;
  assign n22585 = n1538 ^ n277 ^ 1'b0 ;
  assign n22586 = n22585 ^ n13326 ^ n6177 ;
  assign n22587 = n22586 ^ n10454 ^ 1'b0 ;
  assign n22588 = n22587 ^ n8005 ^ 1'b0 ;
  assign n22589 = n12320 & n12460 ;
  assign n22590 = n22589 ^ n1984 ^ 1'b0 ;
  assign n22591 = ~n4693 & n12183 ;
  assign n22592 = n22591 ^ n12843 ^ 1'b0 ;
  assign n22593 = n22592 ^ n19400 ^ 1'b0 ;
  assign n22594 = n4780 ^ n1539 ^ 1'b0 ;
  assign n22596 = ~n792 & n8460 ;
  assign n22595 = n5664 | n9687 ;
  assign n22597 = n22596 ^ n22595 ^ 1'b0 ;
  assign n22600 = ~n792 & n5311 ;
  assign n22601 = ( n7234 & ~n7405 ) | ( n7234 & n22600 ) | ( ~n7405 & n22600 ) ;
  assign n22602 = n11009 & n22601 ;
  assign n22603 = n6895 & n22602 ;
  assign n22598 = n8362 ^ n1497 ^ 1'b0 ;
  assign n22599 = n22598 ^ n2666 ^ n1242 ;
  assign n22604 = n22603 ^ n22599 ^ n6761 ;
  assign n22605 = n5070 ^ n522 ^ 1'b0 ;
  assign n22606 = ~n15230 & n22605 ;
  assign n22607 = n6160 ^ n3655 ^ 1'b0 ;
  assign n22608 = ~n2771 & n22607 ;
  assign n22609 = n6975 & n22608 ;
  assign n22610 = n22609 ^ n1230 ^ 1'b0 ;
  assign n22611 = ~n1493 & n22610 ;
  assign n22612 = n16823 ^ n12693 ^ 1'b0 ;
  assign n22613 = n10140 ^ n4832 ^ 1'b0 ;
  assign n22614 = n22613 ^ n7630 ^ n4357 ;
  assign n22615 = n14177 ^ n9072 ^ 1'b0 ;
  assign n22616 = ( ~n5594 & n13393 ) | ( ~n5594 & n22615 ) | ( n13393 & n22615 ) ;
  assign n22617 = n15202 ^ n13964 ^ 1'b0 ;
  assign n22618 = n2796 & n22617 ;
  assign n22619 = ~n5139 & n10129 ;
  assign n22620 = n4095 | n22619 ;
  assign n22621 = n22618 | n22620 ;
  assign n22622 = n5564 & n18353 ;
  assign n22623 = n15206 ^ n10895 ^ 1'b0 ;
  assign n22624 = n3556 & n5057 ;
  assign n22625 = n7583 & n22624 ;
  assign n22626 = n9339 ^ n4518 ^ 1'b0 ;
  assign n22627 = n1530 & ~n22626 ;
  assign n22628 = ~n10759 & n16184 ;
  assign n22629 = ~n15940 & n19224 ;
  assign n22630 = n16217 & ~n22629 ;
  assign n22631 = n4291 ^ n716 ^ 1'b0 ;
  assign n22632 = n2631 & n22631 ;
  assign n22633 = ~n8230 & n22632 ;
  assign n22634 = n2519 & n22633 ;
  assign n22635 = ~n13044 & n22634 ;
  assign n22636 = ~n3838 & n7197 ;
  assign n22637 = n3959 | n8572 ;
  assign n22638 = n4329 & ~n22637 ;
  assign n22639 = n11437 | n12239 ;
  assign n22640 = n13096 | n22639 ;
  assign n22641 = n1347 & ~n5185 ;
  assign n22642 = n14602 | n22641 ;
  assign n22643 = ~n5115 & n12280 ;
  assign n22644 = n22642 & n22643 ;
  assign n22645 = n22644 ^ n983 ^ 1'b0 ;
  assign n22646 = ( n6216 & n6910 ) | ( n6216 & ~n15590 ) | ( n6910 & ~n15590 ) ;
  assign n22647 = n20254 ^ n1313 ^ 1'b0 ;
  assign n22648 = ~n22646 & n22647 ;
  assign n22649 = n4831 | n9124 ;
  assign n22650 = n22649 ^ n3212 ^ 1'b0 ;
  assign n22651 = n22650 ^ n1877 ^ 1'b0 ;
  assign n22652 = n22651 ^ n902 ^ 1'b0 ;
  assign n22653 = ~n14616 & n22652 ;
  assign n22654 = ( ~n170 & n7457 ) | ( ~n170 & n22653 ) | ( n7457 & n22653 ) ;
  assign n22655 = n19611 ^ n16310 ^ 1'b0 ;
  assign n22656 = n22654 & ~n22655 ;
  assign n22657 = n312 | n1514 ;
  assign n22658 = n22657 ^ n5693 ^ 1'b0 ;
  assign n22659 = n3502 & ~n5100 ;
  assign n22660 = n22658 & n22659 ;
  assign n22661 = ~n5267 & n22660 ;
  assign n22662 = n3194 & n22661 ;
  assign n22663 = ~n16555 & n22624 ;
  assign n22664 = n4142 & ~n22663 ;
  assign n22665 = ~n5748 & n22664 ;
  assign n22666 = n1870 | n8665 ;
  assign n22667 = n22666 ^ n13370 ^ 1'b0 ;
  assign n22668 = ( ~n547 & n14429 ) | ( ~n547 & n22629 ) | ( n14429 & n22629 ) ;
  assign n22669 = ~n2943 & n22668 ;
  assign n22670 = n9150 & n15094 ;
  assign n22671 = n13860 | n18996 ;
  assign n22672 = n1884 & n2287 ;
  assign n22673 = ~n5269 & n8103 ;
  assign n22674 = n22673 ^ n4135 ^ 1'b0 ;
  assign n22675 = n22624 ^ n19281 ^ 1'b0 ;
  assign n22676 = n9518 ^ n1066 ^ 1'b0 ;
  assign n22677 = ~n15634 & n22676 ;
  assign n22678 = ~n16313 & n22677 ;
  assign n22679 = n9150 & n11458 ;
  assign n22680 = n15459 & ~n22679 ;
  assign n22681 = ( n2321 & n3395 ) | ( n2321 & n6239 ) | ( n3395 & n6239 ) ;
  assign n22684 = n9690 | n15612 ;
  assign n22683 = n2772 & ~n11649 ;
  assign n22685 = n22684 ^ n22683 ^ 1'b0 ;
  assign n22686 = n3665 & ~n22685 ;
  assign n22682 = n11021 | n15853 ;
  assign n22687 = n22686 ^ n22682 ^ 1'b0 ;
  assign n22688 = n6043 ^ n3006 ^ 1'b0 ;
  assign n22689 = n8516 & ~n22688 ;
  assign n22690 = ~n3327 & n10809 ;
  assign n22691 = ~n1165 & n22690 ;
  assign n22692 = n22689 & ~n22691 ;
  assign n22693 = ~n13626 & n22692 ;
  assign n22694 = ~n749 & n4479 ;
  assign n22695 = n81 | n22694 ;
  assign n22696 = n11276 ^ n6943 ^ 1'b0 ;
  assign n22697 = ~n8803 & n22696 ;
  assign n22698 = n220 | n5166 ;
  assign n22699 = n7666 & ~n22698 ;
  assign n22700 = ~n20168 & n22699 ;
  assign n22701 = n22697 & ~n22700 ;
  assign n22702 = n77 & n6472 ;
  assign n22703 = n5364 | n10423 ;
  assign n22704 = n16032 ^ n6726 ^ 1'b0 ;
  assign n22705 = ~n8619 & n22704 ;
  assign n22706 = n22705 ^ n6559 ^ 1'b0 ;
  assign n22707 = n8909 & n16876 ;
  assign n22708 = n7961 & n22707 ;
  assign n22709 = ~n7767 & n11681 ;
  assign n22710 = ~n4947 & n22709 ;
  assign n22711 = ~n5747 & n22710 ;
  assign n22712 = n2978 ^ n2467 ^ n1085 ;
  assign n22713 = n6075 ^ n725 ^ 1'b0 ;
  assign n22714 = n22712 & n22713 ;
  assign n22715 = n22714 ^ n15370 ^ 1'b0 ;
  assign n22716 = ~n5695 & n22715 ;
  assign n22717 = n22716 ^ n17449 ^ 1'b0 ;
  assign n22719 = ~n12336 & n12634 ;
  assign n22720 = n22719 ^ n15569 ^ 1'b0 ;
  assign n22721 = n4044 & ~n22720 ;
  assign n22722 = ~n4044 & n22721 ;
  assign n22718 = ~n6628 & n7444 ;
  assign n22723 = n22722 ^ n22718 ^ 1'b0 ;
  assign n22724 = ~n1155 & n22723 ;
  assign n22726 = n8838 ^ n6261 ^ n6229 ;
  assign n22725 = n10851 & ~n20659 ;
  assign n22727 = n22726 ^ n22725 ^ 1'b0 ;
  assign n22728 = n3386 | n17484 ;
  assign n22729 = n16880 | n22728 ;
  assign n22730 = n1464 | n22729 ;
  assign n22731 = n9784 & n12433 ;
  assign n22732 = ~n9784 & n22731 ;
  assign n22733 = n1944 | n22732 ;
  assign n22734 = n10783 & ~n22733 ;
  assign n22735 = n22733 & n22734 ;
  assign n22736 = n8129 ^ n1567 ^ 1'b0 ;
  assign n22737 = n18218 ^ n5656 ^ 1'b0 ;
  assign n22738 = n22737 ^ n3738 ^ 1'b0 ;
  assign n22739 = n6783 ^ n5773 ^ 1'b0 ;
  assign n22740 = ( n5637 & n16603 ) | ( n5637 & n22739 ) | ( n16603 & n22739 ) ;
  assign n22741 = n91 | n22740 ;
  assign n22742 = n22741 ^ n4978 ^ 1'b0 ;
  assign n22743 = n7471 | n22742 ;
  assign n22744 = n22743 ^ n6154 ^ 1'b0 ;
  assign n22745 = n1914 & ~n19028 ;
  assign n22746 = n22744 & n22745 ;
  assign n22747 = n22746 ^ n3042 ^ 1'b0 ;
  assign n22748 = n22738 & n22747 ;
  assign n22749 = ( n2137 & ~n6874 ) | ( n2137 & n8710 ) | ( ~n6874 & n8710 ) ;
  assign n22750 = ~n4533 & n8887 ;
  assign n22751 = n22750 ^ n4790 ^ 1'b0 ;
  assign n22752 = n22751 ^ n18129 ^ 1'b0 ;
  assign n22753 = ~n365 & n22752 ;
  assign n22754 = n9848 ^ n9667 ^ 1'b0 ;
  assign n22755 = n19019 | n22754 ;
  assign n22756 = ~n15308 & n22755 ;
  assign n22757 = n1182 & ~n4732 ;
  assign n22758 = ~n10023 & n12185 ;
  assign n22759 = ~n22757 & n22758 ;
  assign n22760 = n365 & n3213 ;
  assign n22761 = ~n12582 & n22760 ;
  assign n22762 = n793 | n22761 ;
  assign n22763 = n22759 & ~n22762 ;
  assign n22764 = n5893 ^ n2594 ^ 1'b0 ;
  assign n22765 = ~n3165 & n12050 ;
  assign n22766 = n1645 & n22765 ;
  assign n22767 = n18310 ^ n11648 ^ 1'b0 ;
  assign n22768 = ( ~n15847 & n22766 ) | ( ~n15847 & n22767 ) | ( n22766 & n22767 ) ;
  assign n22769 = n18833 ^ n15261 ^ 1'b0 ;
  assign n22771 = n1832 | n15424 ;
  assign n22770 = n8740 ^ n3977 ^ 1'b0 ;
  assign n22772 = n22771 ^ n22770 ^ n5119 ;
  assign n22773 = n8030 ^ n6663 ^ n5474 ;
  assign n22774 = n17193 ^ n12893 ^ 1'b0 ;
  assign n22775 = n22773 & ~n22774 ;
  assign n22776 = n10237 ^ n7727 ^ 1'b0 ;
  assign n22777 = n16824 & ~n22776 ;
  assign n22778 = n12141 & ~n13454 ;
  assign n22779 = ~n183 & n10205 ;
  assign n22780 = n15005 ^ n2079 ^ 1'b0 ;
  assign n22781 = n15138 ^ n9584 ^ n241 ;
  assign n22782 = n6572 & ~n22781 ;
  assign n22783 = n22448 ^ n19632 ^ 1'b0 ;
  assign n22784 = ( n23 & n2739 ) | ( n23 & n9962 ) | ( n2739 & n9962 ) ;
  assign n22785 = n22784 ^ n3891 ^ 1'b0 ;
  assign n22786 = ~n22783 & n22785 ;
  assign n22787 = n6045 | n15944 ;
  assign n22788 = n8136 & n10945 ;
  assign n22789 = n22788 ^ n11621 ^ 1'b0 ;
  assign n22790 = ~n431 & n4157 ;
  assign n22791 = ~n1732 & n22790 ;
  assign n22792 = n11144 | n22791 ;
  assign n22793 = n22418 ^ n4754 ^ 1'b0 ;
  assign n22794 = n453 & ~n12849 ;
  assign n22795 = n22794 ^ n2272 ^ 1'b0 ;
  assign n22796 = n3220 | n7958 ;
  assign n22797 = n11875 & ~n22796 ;
  assign n22798 = n8266 & n22797 ;
  assign n22799 = n16463 | n20257 ;
  assign n22800 = ( ~n20442 & n22798 ) | ( ~n20442 & n22799 ) | ( n22798 & n22799 ) ;
  assign n22801 = n4865 ^ n1226 ^ 1'b0 ;
  assign n22802 = n8012 | n22801 ;
  assign n22803 = n22802 ^ n7531 ^ 1'b0 ;
  assign n22804 = n7606 & ~n11366 ;
  assign n22805 = n9915 ^ n88 ^ 1'b0 ;
  assign n22806 = n22805 ^ n17994 ^ 1'b0 ;
  assign n22807 = n19842 | n22806 ;
  assign n22808 = n16462 & ~n22807 ;
  assign n22809 = ~n404 & n7197 ;
  assign n22810 = n22809 ^ n2227 ^ 1'b0 ;
  assign n22811 = n5773 & n16150 ;
  assign n22812 = ~n12592 & n22811 ;
  assign n22813 = n5944 & n14897 ;
  assign n22814 = ~n13626 & n22813 ;
  assign n22815 = n18009 ^ n16110 ^ 1'b0 ;
  assign n22816 = n22814 | n22815 ;
  assign n22817 = n21769 ^ n3833 ^ 1'b0 ;
  assign n22818 = n402 | n22817 ;
  assign n22819 = ~n12173 & n18301 ;
  assign n22820 = n22819 ^ n17569 ^ 1'b0 ;
  assign n22821 = n18362 ^ n5443 ^ 1'b0 ;
  assign n22822 = n18126 & ~n22821 ;
  assign n22823 = ( n8120 & n21621 ) | ( n8120 & ~n22822 ) | ( n21621 & ~n22822 ) ;
  assign n22824 = n21767 ^ n260 ^ 1'b0 ;
  assign n22825 = n2769 | n22824 ;
  assign n22826 = n2789 & ~n22825 ;
  assign n22827 = n1814 & n9146 ;
  assign n22828 = n22384 ^ n14780 ^ n11222 ;
  assign n22829 = ~n1155 & n9290 ;
  assign n22830 = ~n3715 & n22829 ;
  assign n22831 = n1194 & ~n4760 ;
  assign n22832 = n22262 ^ n17692 ^ 1'b0 ;
  assign n22833 = n12513 & ~n22832 ;
  assign n22834 = ~n9393 & n13797 ;
  assign n22835 = n14259 | n22834 ;
  assign n22836 = n422 | n22835 ;
  assign n22837 = ( n4720 & n15062 ) | ( n4720 & ~n21042 ) | ( n15062 & ~n21042 ) ;
  assign n22838 = n2202 & n22837 ;
  assign n22839 = ~n11006 & n22838 ;
  assign n22840 = n22059 ^ n19026 ^ 1'b0 ;
  assign n22841 = n20128 ^ n2989 ^ 1'b0 ;
  assign n22842 = n10059 ^ n5391 ^ 1'b0 ;
  assign n22843 = ~n9344 & n22842 ;
  assign n22844 = n15796 & n22843 ;
  assign n22845 = n22844 ^ n877 ^ 1'b0 ;
  assign n22846 = n5748 & n22845 ;
  assign n22847 = n2437 | n16729 ;
  assign n22848 = n11946 ^ n8263 ^ n5130 ;
  assign n22849 = ~n15043 & n17537 ;
  assign n22850 = n22849 ^ n18571 ^ 1'b0 ;
  assign n22851 = ~n4937 & n18786 ;
  assign n22852 = n12586 ^ n11081 ^ 1'b0 ;
  assign n22853 = n15299 & n22852 ;
  assign n22854 = n16197 ^ n2053 ^ 1'b0 ;
  assign n22855 = n2650 | n9049 ;
  assign n22856 = ~n6045 & n14059 ;
  assign n22857 = n7015 ^ n6256 ^ 1'b0 ;
  assign n22858 = n22857 ^ n12655 ^ 1'b0 ;
  assign n22859 = n22858 ^ n10368 ^ 1'b0 ;
  assign n22860 = ( n4481 & ~n7981 ) | ( n4481 & n13002 ) | ( ~n7981 & n13002 ) ;
  assign n22861 = n14552 & n22860 ;
  assign n22862 = ~n3058 & n22861 ;
  assign n22863 = n1045 ^ n408 ^ 1'b0 ;
  assign n22864 = n3240 | n10783 ;
  assign n22865 = n5131 & n15624 ;
  assign n22866 = n22865 ^ n6350 ^ 1'b0 ;
  assign n22867 = n21810 | n22866 ;
  assign n22868 = n2231 | n22867 ;
  assign n22869 = n2078 & n6527 ;
  assign n22870 = n8652 | n13342 ;
  assign n22871 = n7568 ^ n2772 ^ 1'b0 ;
  assign n22872 = n16681 | n22871 ;
  assign n22873 = ~n6635 & n9102 ;
  assign n22874 = n22873 ^ n5150 ^ 1'b0 ;
  assign n22875 = n14969 | n22874 ;
  assign n22876 = n7529 | n12484 ;
  assign n22877 = n12717 & ~n22876 ;
  assign n22878 = ~n15497 & n17364 ;
  assign n22879 = n22878 ^ n8153 ^ 1'b0 ;
  assign n22880 = n22879 ^ n4105 ^ 1'b0 ;
  assign n22881 = n200 & ~n22880 ;
  assign n22882 = n2355 | n3520 ;
  assign n22883 = n7616 ^ n7014 ^ 1'b0 ;
  assign n22884 = n1018 | n22883 ;
  assign n22885 = n22884 ^ n1300 ^ 1'b0 ;
  assign n22886 = ~n9970 & n22885 ;
  assign n22887 = n22886 ^ n20366 ^ n11034 ;
  assign n22888 = n267 & n10783 ;
  assign n22889 = n3623 & n22888 ;
  assign n22890 = n22889 ^ n5005 ^ 1'b0 ;
  assign n22891 = n11453 | n18928 ;
  assign n22892 = n22891 ^ n3343 ^ 1'b0 ;
  assign n22893 = n5755 | n22892 ;
  assign n22894 = n12082 ^ n7412 ^ 1'b0 ;
  assign n22895 = n1690 & ~n4318 ;
  assign n22896 = n11874 ^ n858 ^ 1'b0 ;
  assign n22901 = n710 | n7191 ;
  assign n22897 = n8474 | n13491 ;
  assign n22898 = n7893 & ~n22897 ;
  assign n22899 = n8996 & ~n22898 ;
  assign n22900 = n20381 & n22899 ;
  assign n22902 = n22901 ^ n22900 ^ n6640 ;
  assign n22903 = n10908 ^ n5896 ^ 1'b0 ;
  assign n22904 = n4357 ^ n1435 ^ 1'b0 ;
  assign n22905 = ~n22903 & n22904 ;
  assign n22906 = ~n757 & n2664 ;
  assign n22907 = ~n9769 & n13108 ;
  assign n22908 = n22907 ^ n4302 ^ n1847 ;
  assign n22909 = ( n2386 & n3063 ) | ( n2386 & n4688 ) | ( n3063 & n4688 ) ;
  assign n22910 = n22909 ^ n7476 ^ 1'b0 ;
  assign n22911 = n22908 & n22910 ;
  assign n22912 = n17061 ^ n3231 ^ 1'b0 ;
  assign n22913 = n52 & n22912 ;
  assign n22914 = n3791 & ~n4988 ;
  assign n22915 = n16651 ^ n668 ^ 1'b0 ;
  assign n22916 = n22914 & ~n22915 ;
  assign n22917 = n22916 ^ n16003 ^ 1'b0 ;
  assign n22918 = n4999 ^ n2205 ^ 1'b0 ;
  assign n22919 = n19884 & n22918 ;
  assign n22920 = n8951 ^ n1306 ^ 1'b0 ;
  assign n22921 = n7151 | n21353 ;
  assign n22922 = n10864 | n16382 ;
  assign n22923 = n3768 & ~n22922 ;
  assign n22924 = ~n14115 & n22923 ;
  assign n22925 = ( n918 & ~n3178 ) | ( n918 & n21857 ) | ( ~n3178 & n21857 ) ;
  assign n22928 = n12899 ^ n10544 ^ 1'b0 ;
  assign n22929 = n3943 | n22928 ;
  assign n22930 = n21518 | n22929 ;
  assign n22926 = n3630 & n3851 ;
  assign n22927 = n22926 ^ n10436 ^ 1'b0 ;
  assign n22931 = n22930 ^ n22927 ^ 1'b0 ;
  assign n22932 = n10492 & n19142 ;
  assign n22933 = n22932 ^ n922 ^ 1'b0 ;
  assign n22934 = n4344 & n22933 ;
  assign n22935 = ~n886 & n5562 ;
  assign n22937 = n4231 ^ n61 ^ 1'b0 ;
  assign n22936 = n1469 | n2833 ;
  assign n22938 = n22937 ^ n22936 ^ n9397 ;
  assign n22939 = n9535 ^ n40 ^ 1'b0 ;
  assign n22940 = n22939 ^ n3959 ^ 1'b0 ;
  assign n22941 = n6891 & n22940 ;
  assign n22945 = n15961 ^ n15716 ^ 1'b0 ;
  assign n22946 = n4774 & ~n22945 ;
  assign n22942 = n495 & ~n4862 ;
  assign n22943 = n4504 ^ n2335 ^ 1'b0 ;
  assign n22944 = n22942 | n22943 ;
  assign n22947 = n22946 ^ n22944 ^ 1'b0 ;
  assign n22948 = n1819 | n2758 ;
  assign n22949 = n873 | n22948 ;
  assign n22950 = n22947 | n22949 ;
  assign n22951 = n14094 | n20908 ;
  assign n22952 = n22951 ^ n6645 ^ 1'b0 ;
  assign n22953 = n22952 ^ n221 ^ 1'b0 ;
  assign n22954 = n1289 & n8628 ;
  assign n22955 = n22954 ^ n15952 ^ 1'b0 ;
  assign n22956 = n17423 & n22955 ;
  assign n22963 = n7673 ^ n205 ^ 1'b0 ;
  assign n22958 = ~n4312 & n4734 ;
  assign n22959 = n22958 ^ n2086 ^ 1'b0 ;
  assign n22957 = ~n1994 & n9839 ;
  assign n22960 = n22959 ^ n22957 ^ 1'b0 ;
  assign n22961 = n22960 ^ n15400 ^ n2492 ;
  assign n22962 = n22879 & n22961 ;
  assign n22964 = n22963 ^ n22962 ^ 1'b0 ;
  assign n22965 = n4501 & n6526 ;
  assign n22966 = n22965 ^ n9208 ^ 1'b0 ;
  assign n22967 = n15454 ^ n2806 ^ 1'b0 ;
  assign n22968 = n22966 | n22967 ;
  assign n22969 = ( ~n614 & n7269 ) | ( ~n614 & n8026 ) | ( n7269 & n8026 ) ;
  assign n22970 = n6509 & n22969 ;
  assign n22971 = n22970 ^ n9992 ^ 1'b0 ;
  assign n22972 = n14057 ^ n13517 ^ 1'b0 ;
  assign n22973 = n338 & ~n2236 ;
  assign n22974 = n22973 ^ n795 ^ 1'b0 ;
  assign n22975 = n1337 | n6291 ;
  assign n22976 = n1337 & ~n22975 ;
  assign n22977 = n22974 & ~n22976 ;
  assign n22978 = ~n22974 & n22977 ;
  assign n22979 = n20646 ^ n6415 ^ 1'b0 ;
  assign n22980 = n6861 & ~n9899 ;
  assign n22981 = n14316 ^ n2313 ^ n1038 ;
  assign n22982 = n22981 ^ n1142 ^ 1'b0 ;
  assign n22983 = ~n1367 & n7934 ;
  assign n22984 = n22983 ^ n1355 ^ 1'b0 ;
  assign n22985 = n15807 & n22984 ;
  assign n22986 = n15969 ^ n14512 ^ 1'b0 ;
  assign n22987 = n7997 & ~n22986 ;
  assign n22988 = n22987 ^ n16888 ^ 1'b0 ;
  assign n22989 = n17697 ^ n14670 ^ 1'b0 ;
  assign n22990 = n11363 & ~n22989 ;
  assign n22991 = ( n3082 & ~n22988 ) | ( n3082 & n22990 ) | ( ~n22988 & n22990 ) ;
  assign n22992 = ( n1432 & ~n6330 ) | ( n1432 & n13883 ) | ( ~n6330 & n13883 ) ;
  assign n22993 = n22992 ^ n2596 ^ 1'b0 ;
  assign n22994 = n22236 & ~n22993 ;
  assign n22995 = ~n5290 & n17321 ;
  assign n22996 = n13986 ^ n2352 ^ 1'b0 ;
  assign n22997 = ~n2452 & n16749 ;
  assign n22998 = ~n4250 & n22997 ;
  assign n22999 = n7893 ^ n5414 ^ 1'b0 ;
  assign n23000 = n3833 ^ n1329 ^ 1'b0 ;
  assign n23001 = n762 | n23000 ;
  assign n23002 = n23001 ^ n18884 ^ 1'b0 ;
  assign n23003 = n22999 & ~n23002 ;
  assign n23004 = n9170 | n17427 ;
  assign n23005 = n23004 ^ n17836 ^ 1'b0 ;
  assign n23006 = n17108 ^ n5433 ^ n209 ;
  assign n23007 = n23006 ^ n8945 ^ 1'b0 ;
  assign n23008 = n3372 | n23007 ;
  assign n23009 = n5399 & n13131 ;
  assign n23010 = n23008 & n23009 ;
  assign n23011 = n15088 ^ n7314 ^ 1'b0 ;
  assign n23012 = n9256 & ~n9850 ;
  assign n23013 = ~n11502 & n23012 ;
  assign n23014 = n23011 & ~n23013 ;
  assign n23015 = n23014 ^ n753 ^ 1'b0 ;
  assign n23016 = n3012 | n6239 ;
  assign n23017 = ~n14817 & n23016 ;
  assign n23018 = n9421 | n12799 ;
  assign n23019 = n23018 ^ n15803 ^ 1'b0 ;
  assign n23020 = n3651 & ~n9928 ;
  assign n23021 = n20340 ^ n10423 ^ n1044 ;
  assign n23022 = ( n7379 & n23020 ) | ( n7379 & ~n23021 ) | ( n23020 & ~n23021 ) ;
  assign n23023 = n23019 & n23022 ;
  assign n23024 = n18114 ^ n2610 ^ 1'b0 ;
  assign n23025 = ~n4395 & n23024 ;
  assign n23026 = n10632 | n13436 ;
  assign n23027 = n8529 & ~n23026 ;
  assign n23028 = n21079 & n23027 ;
  assign n23029 = n23028 ^ n6028 ^ 1'b0 ;
  assign n23030 = ~n15113 & n23029 ;
  assign n23031 = n4279 & ~n11090 ;
  assign n23032 = n4348 | n5697 ;
  assign n23033 = n6910 | n23032 ;
  assign n23034 = n1481 ^ n1157 ^ 1'b0 ;
  assign n23035 = ~n56 & n23034 ;
  assign n23036 = ~n8971 & n23035 ;
  assign n23037 = n23036 ^ n8978 ^ 1'b0 ;
  assign n23038 = n11532 | n23037 ;
  assign n23039 = n4218 | n9139 ;
  assign n23040 = ( n1416 & ~n21950 ) | ( n1416 & n23039 ) | ( ~n21950 & n23039 ) ;
  assign n23041 = n9688 | n12155 ;
  assign n23042 = n7554 | n23041 ;
  assign n23047 = n13685 ^ n2081 ^ 1'b0 ;
  assign n23048 = n1090 & ~n23047 ;
  assign n23049 = n315 & ~n974 ;
  assign n23050 = ~n8072 & n23049 ;
  assign n23051 = ~n23048 & n23050 ;
  assign n23043 = n11955 ^ n3943 ^ 1'b0 ;
  assign n23044 = n23043 ^ n3911 ^ 1'b0 ;
  assign n23045 = n7679 | n23044 ;
  assign n23046 = n12699 & n23045 ;
  assign n23052 = n23051 ^ n23046 ^ 1'b0 ;
  assign n23053 = ( ~n466 & n11726 ) | ( ~n466 & n22624 ) | ( n11726 & n22624 ) ;
  assign n23054 = n835 & n7040 ;
  assign n23055 = n1981 & ~n19681 ;
  assign n23056 = n2930 | n4139 ;
  assign n23057 = n23056 ^ n5188 ^ 1'b0 ;
  assign n23058 = n23057 ^ n12849 ^ 1'b0 ;
  assign n23059 = n27 & n23058 ;
  assign n23060 = n11292 & n23059 ;
  assign n23061 = n10604 & ~n21329 ;
  assign n23062 = n23061 ^ n2400 ^ 1'b0 ;
  assign n23064 = n5367 & ~n15527 ;
  assign n23065 = n23064 ^ n9536 ^ 1'b0 ;
  assign n23063 = n12922 ^ n7165 ^ 1'b0 ;
  assign n23066 = n23065 ^ n23063 ^ 1'b0 ;
  assign n23067 = ( n15185 & n17860 ) | ( n15185 & ~n23066 ) | ( n17860 & ~n23066 ) ;
  assign n23068 = n3591 & n8082 ;
  assign n23069 = n188 & n23068 ;
  assign n23070 = n13262 & ~n23069 ;
  assign n23071 = ~n20340 & n23070 ;
  assign n23072 = n13340 ^ n209 ^ 1'b0 ;
  assign n23073 = n18530 | n23072 ;
  assign n23074 = n4002 | n9312 ;
  assign n23075 = n10760 ^ n564 ^ 1'b0 ;
  assign n23076 = n23075 ^ n1701 ^ 1'b0 ;
  assign n23077 = n4131 & ~n7020 ;
  assign n23078 = n5410 ^ n2717 ^ 1'b0 ;
  assign n23079 = n23078 ^ n20065 ^ 1'b0 ;
  assign n23080 = n20866 | n23079 ;
  assign n23081 = n7475 ^ n113 ^ 1'b0 ;
  assign n23082 = n23081 ^ n14250 ^ 1'b0 ;
  assign n23083 = n6583 | n13471 ;
  assign n23084 = n23083 ^ n18122 ^ 1'b0 ;
  assign n23085 = n14356 ^ n14075 ^ 1'b0 ;
  assign n23086 = ~n1538 & n7257 ;
  assign n23087 = n23086 ^ n20798 ^ 1'b0 ;
  assign n23088 = n23085 & ~n23087 ;
  assign n23089 = n1269 & n12458 ;
  assign n23090 = n17185 ^ n7073 ^ 1'b0 ;
  assign n23091 = n8403 ^ n283 ^ 1'b0 ;
  assign n23092 = n1867 | n23091 ;
  assign n23093 = ~n646 & n4195 ;
  assign n23094 = ( n18598 & n23092 ) | ( n18598 & n23093 ) | ( n23092 & n23093 ) ;
  assign n23095 = n9358 ^ n3186 ^ 1'b0 ;
  assign n23096 = n19834 | n23095 ;
  assign n23097 = n8128 & ~n23096 ;
  assign n23098 = n9564 & ~n23097 ;
  assign n23099 = n23098 ^ n20242 ^ 1'b0 ;
  assign n23100 = n23099 ^ n1941 ^ 1'b0 ;
  assign n23101 = n4037 ^ n1163 ^ 1'b0 ;
  assign n23102 = n23101 ^ n17607 ^ n9323 ;
  assign n23103 = n1694 | n23102 ;
  assign n23104 = n23103 ^ n12024 ^ 1'b0 ;
  assign n23105 = ~n2843 & n17032 ;
  assign n23106 = n19372 & n23105 ;
  assign n23107 = n798 | n16478 ;
  assign n23108 = n5453 | n23107 ;
  assign n23109 = n23108 ^ n5809 ^ 1'b0 ;
  assign n23110 = n17110 ^ n12340 ^ 1'b0 ;
  assign n23111 = n1178 & n3537 ;
  assign n23112 = n23111 ^ n5814 ^ 1'b0 ;
  assign n23113 = n11727 ^ n3095 ^ 1'b0 ;
  assign n23114 = n23112 & n23113 ;
  assign n23115 = n23114 ^ n17102 ^ 1'b0 ;
  assign n23116 = ~n1456 & n16430 ;
  assign n23117 = n6070 | n14622 ;
  assign n23118 = n21849 ^ n7611 ^ n3118 ;
  assign n23119 = n23118 ^ n3438 ^ 1'b0 ;
  assign n23120 = n513 & ~n23119 ;
  assign n23121 = n4639 ^ n2134 ^ 1'b0 ;
  assign n23122 = n23120 & ~n23121 ;
  assign n23123 = n7648 ^ n5054 ^ 1'b0 ;
  assign n23124 = n10855 ^ n8553 ^ 1'b0 ;
  assign n23125 = n2290 & n3887 ;
  assign n23126 = n23125 ^ n3079 ^ 1'b0 ;
  assign n23127 = ~n6527 & n23126 ;
  assign n23128 = n23127 ^ n7383 ^ 1'b0 ;
  assign n23129 = ~n11582 & n23128 ;
  assign n23130 = ~n1772 & n23129 ;
  assign n23131 = n7106 & n8452 ;
  assign n23132 = n3968 | n23131 ;
  assign n23133 = n23132 ^ n8721 ^ 1'b0 ;
  assign n23134 = n23133 ^ n5651 ^ 1'b0 ;
  assign n23136 = n860 | n2195 ;
  assign n23137 = n23136 ^ n631 ^ 1'b0 ;
  assign n23138 = ~n15618 & n23137 ;
  assign n23135 = n3209 | n14636 ;
  assign n23139 = n23138 ^ n23135 ^ 1'b0 ;
  assign n23140 = n23139 ^ n6672 ^ n5953 ;
  assign n23141 = n10430 | n11661 ;
  assign n23142 = n23141 ^ n105 ^ 1'b0 ;
  assign n23143 = n3903 & n23142 ;
  assign n23144 = n1506 | n7284 ;
  assign n23145 = n23144 ^ n17702 ^ 1'b0 ;
  assign n23146 = n2199 & n8061 ;
  assign n23147 = n23146 ^ n22389 ^ 1'b0 ;
  assign n23148 = n844 | n6230 ;
  assign n23149 = n8646 ^ n2489 ^ 1'b0 ;
  assign n23150 = ~n12464 & n23149 ;
  assign n23151 = n20592 & n23150 ;
  assign n23152 = n4009 | n13543 ;
  assign n23153 = n13739 | n21715 ;
  assign n23154 = n23152 & ~n23153 ;
  assign n23155 = n17190 ^ n6713 ^ 1'b0 ;
  assign n23156 = n4958 | n20644 ;
  assign n23157 = ~n22869 & n23156 ;
  assign n23158 = n23157 ^ n7833 ^ 1'b0 ;
  assign n23159 = n9792 | n14095 ;
  assign n23160 = n6129 | n23159 ;
  assign n23161 = n2610 | n17013 ;
  assign n23162 = n7915 & ~n23161 ;
  assign n23163 = n2391 & ~n3843 ;
  assign n23164 = n1141 & n17903 ;
  assign n23165 = n5936 | n18763 ;
  assign n23166 = n14812 & n18412 ;
  assign n23167 = n1329 & ~n14500 ;
  assign n23168 = n23167 ^ n8291 ^ 1'b0 ;
  assign n23169 = n15007 | n23168 ;
  assign n23170 = ( ~n11058 & n17871 ) | ( ~n11058 & n19273 ) | ( n17871 & n19273 ) ;
  assign n23171 = n20835 ^ n5589 ^ 1'b0 ;
  assign n23172 = n20726 & ~n23171 ;
  assign n23173 = n1700 & n10721 ;
  assign n23174 = n19182 ^ n10348 ^ 1'b0 ;
  assign n23175 = n11777 & n23174 ;
  assign n23176 = n5041 | n18996 ;
  assign n23177 = n8714 | n20002 ;
  assign n23178 = n4799 | n23177 ;
  assign n23179 = n23178 ^ n9388 ^ n2962 ;
  assign n23180 = n1282 & n2101 ;
  assign n23181 = n3861 & n23180 ;
  assign n23182 = n23181 ^ n4945 ^ 1'b0 ;
  assign n23187 = ~n1848 & n12786 ;
  assign n23188 = n5815 & n23187 ;
  assign n23189 = n23188 ^ n5289 ^ 1'b0 ;
  assign n23183 = n10076 ^ n5810 ^ 1'b0 ;
  assign n23184 = n23183 ^ n901 ^ 1'b0 ;
  assign n23185 = ~n567 & n23184 ;
  assign n23186 = n7585 & n23185 ;
  assign n23190 = n23189 ^ n23186 ^ 1'b0 ;
  assign n23191 = n12513 ^ n5329 ^ 1'b0 ;
  assign n23192 = n23190 | n23191 ;
  assign n23193 = n6889 & n12603 ;
  assign n23194 = n2832 & n8027 ;
  assign n23195 = n17684 ^ n10212 ^ n2694 ;
  assign n23196 = n14937 ^ n2284 ^ 1'b0 ;
  assign n23197 = n7589 | n20202 ;
  assign n23198 = n4938 & ~n23197 ;
  assign n23199 = n4276 & ~n8554 ;
  assign n23200 = n23199 ^ n12740 ^ 1'b0 ;
  assign n23201 = ~n1207 & n2090 ;
  assign n23202 = ~n9577 & n23201 ;
  assign n23203 = n8735 | n13739 ;
  assign n23204 = n14675 & n18307 ;
  assign n23205 = ( n23202 & n23203 ) | ( n23202 & ~n23204 ) | ( n23203 & ~n23204 ) ;
  assign n23206 = n5857 ^ n477 ^ 1'b0 ;
  assign n23207 = n8410 & n23206 ;
  assign n23208 = n23207 ^ n17070 ^ 1'b0 ;
  assign n23209 = n23208 ^ n18806 ^ 1'b0 ;
  assign n23210 = n7604 ^ n5137 ^ 1'b0 ;
  assign n23211 = n23209 & ~n23210 ;
  assign n23212 = n6296 | n17011 ;
  assign n23213 = n4550 & ~n23212 ;
  assign n23214 = ~n8944 & n20055 ;
  assign n23215 = ~n4784 & n9586 ;
  assign n23216 = ~n23214 & n23215 ;
  assign n23217 = n1848 & ~n23216 ;
  assign n23218 = n27 & n1701 ;
  assign n23219 = n23218 ^ n5012 ^ 1'b0 ;
  assign n23220 = n768 | n23219 ;
  assign n23221 = n19836 ^ n14200 ^ n7384 ;
  assign n23222 = n972 & n23221 ;
  assign n23223 = ~n2254 & n11515 ;
  assign n23224 = n23223 ^ n12072 ^ n2146 ;
  assign n23225 = n5469 | n23224 ;
  assign n23226 = n5358 | n15856 ;
  assign n23227 = n9245 | n23226 ;
  assign n23228 = n23227 ^ n2872 ^ 1'b0 ;
  assign n23229 = n5073 & ~n23228 ;
  assign n23230 = n19696 | n23229 ;
  assign n23231 = n23230 ^ n12292 ^ 1'b0 ;
  assign n23232 = n17050 ^ n12967 ^ 1'b0 ;
  assign n23233 = n839 & n8161 ;
  assign n23234 = n15076 ^ n11064 ^ 1'b0 ;
  assign n23235 = n23233 & n23234 ;
  assign n23236 = n23235 ^ n6680 ^ 1'b0 ;
  assign n23237 = n12292 | n23236 ;
  assign n23238 = ~n899 & n5646 ;
  assign n23239 = n20296 ^ n6343 ^ 1'b0 ;
  assign n23240 = n5809 & ~n23239 ;
  assign n23241 = ~n1675 & n18146 ;
  assign n23242 = n23241 ^ n13721 ^ 1'b0 ;
  assign n23243 = n10008 ^ n7660 ^ 1'b0 ;
  assign n23244 = n18270 ^ n5885 ^ 1'b0 ;
  assign n23246 = ( n7830 & n14710 ) | ( n7830 & n18545 ) | ( n14710 & n18545 ) ;
  assign n23245 = n10085 & n17256 ;
  assign n23247 = n23246 ^ n23245 ^ 1'b0 ;
  assign n23248 = n640 | n965 ;
  assign n23249 = n23248 ^ n184 ^ 1'b0 ;
  assign n23250 = n4245 ^ n2203 ^ 1'b0 ;
  assign n23251 = n20775 & n23250 ;
  assign n23252 = n959 & n4117 ;
  assign n23253 = ~n9146 & n23252 ;
  assign n23254 = n9395 ^ n135 ^ 1'b0 ;
  assign n23255 = n23253 | n23254 ;
  assign n23256 = n23251 | n23255 ;
  assign n23257 = n18194 ^ n11961 ^ 1'b0 ;
  assign n23258 = n7591 | n23257 ;
  assign n23259 = n23258 ^ n33 ^ 1'b0 ;
  assign n23260 = ~n205 & n23259 ;
  assign n23261 = n528 & n7372 ;
  assign n23262 = n23261 ^ n17352 ^ 1'b0 ;
  assign n23263 = n1327 & ~n23262 ;
  assign n23264 = n12591 ^ n1946 ^ n503 ;
  assign n23265 = n23264 ^ n438 ^ 1'b0 ;
  assign n23266 = ~n2762 & n23265 ;
  assign n23272 = n15292 ^ n6523 ^ n2905 ;
  assign n23267 = n4645 ^ n800 ^ 1'b0 ;
  assign n23268 = n7691 ^ n7427 ^ 1'b0 ;
  assign n23269 = n23267 & ~n23268 ;
  assign n23270 = n23269 ^ n6179 ^ 1'b0 ;
  assign n23271 = n179 & n23270 ;
  assign n23273 = n23272 ^ n23271 ^ n23057 ;
  assign n23274 = n924 & n2374 ;
  assign n23275 = n23274 ^ n7112 ^ n825 ;
  assign n23276 = n23275 ^ n982 ^ 1'b0 ;
  assign n23277 = n23276 ^ n3646 ^ 1'b0 ;
  assign n23278 = ~n23039 & n23277 ;
  assign n23279 = n6741 | n9018 ;
  assign n23280 = n10845 & ~n23279 ;
  assign n23281 = n10855 & ~n23280 ;
  assign n23282 = n669 & ~n23281 ;
  assign n23283 = n23282 ^ n7601 ^ 1'b0 ;
  assign n23284 = n11506 ^ n5279 ^ 1'b0 ;
  assign n23285 = n23283 | n23284 ;
  assign n23286 = n5609 | n6518 ;
  assign n23287 = ~n6817 & n23286 ;
  assign n23288 = n23287 ^ n14067 ^ 1'b0 ;
  assign n23289 = n2031 ^ n910 ^ 1'b0 ;
  assign n23290 = n4209 & ~n18060 ;
  assign n23291 = ( ~n14318 & n19521 ) | ( ~n14318 & n23290 ) | ( n19521 & n23290 ) ;
  assign n23292 = n19338 ^ n3541 ^ 1'b0 ;
  assign n23293 = n1212 & n23292 ;
  assign n23294 = n23293 ^ n18390 ^ 1'b0 ;
  assign n23295 = n6904 | n19520 ;
  assign n23296 = n1863 & n23295 ;
  assign n23297 = n23296 ^ n5146 ^ 1'b0 ;
  assign n23298 = n8905 ^ n805 ^ 1'b0 ;
  assign n23299 = n6711 | n23298 ;
  assign n23300 = n1853 & ~n19762 ;
  assign n23301 = n23300 ^ n13389 ^ 1'b0 ;
  assign n23302 = n13719 ^ n1918 ^ 1'b0 ;
  assign n23303 = n1204 & ~n23302 ;
  assign n23304 = n167 | n9779 ;
  assign n23305 = n2706 & n11931 ;
  assign n23306 = ~n23304 & n23305 ;
  assign n23307 = n3939 ^ n1242 ^ n439 ;
  assign n23308 = n22901 ^ n1658 ^ 1'b0 ;
  assign n23309 = n23307 | n23308 ;
  assign n23310 = n9958 ^ n7731 ^ 1'b0 ;
  assign n23311 = n23309 | n23310 ;
  assign n23312 = n21611 ^ n4691 ^ 1'b0 ;
  assign n23313 = n12666 & n23312 ;
  assign n23314 = ( n1430 & ~n6408 ) | ( n1430 & n6435 ) | ( ~n6408 & n6435 ) ;
  assign n23315 = n14892 ^ n105 ^ 1'b0 ;
  assign n23316 = n23315 ^ n18725 ^ 1'b0 ;
  assign n23324 = x5 & ~n330 ;
  assign n23317 = ~n1843 & n1852 ;
  assign n23318 = ( n2053 & n2205 ) | ( n2053 & n23317 ) | ( n2205 & n23317 ) ;
  assign n23319 = n23318 ^ n2033 ^ 1'b0 ;
  assign n23320 = ~n4550 & n23319 ;
  assign n23321 = n2833 & n23320 ;
  assign n23322 = n7206 & n23321 ;
  assign n23323 = n13934 | n23322 ;
  assign n23325 = n23324 ^ n23323 ^ 1'b0 ;
  assign n23326 = n5093 ^ n4877 ^ 1'b0 ;
  assign n23327 = n6713 | n23326 ;
  assign n23328 = n74 & n7883 ;
  assign n23329 = ( n5961 & n6102 ) | ( n5961 & ~n7167 ) | ( n6102 & ~n7167 ) ;
  assign n23330 = n5047 | n8612 ;
  assign n23331 = n23330 ^ n7048 ^ n6296 ;
  assign n23332 = n23331 ^ n17301 ^ 1'b0 ;
  assign n23333 = n2304 | n23332 ;
  assign n23334 = n23333 ^ n2602 ^ 1'b0 ;
  assign n23335 = n6542 | n23334 ;
  assign n23336 = n1251 & ~n20009 ;
  assign n23337 = n7791 ^ n4810 ^ 1'b0 ;
  assign n23338 = n14121 ^ n2746 ^ 1'b0 ;
  assign n23339 = ~n10001 & n23338 ;
  assign n23340 = n23337 | n23339 ;
  assign n23341 = ~n2189 & n5174 ;
  assign n23342 = ~n12935 & n15699 ;
  assign n23343 = n23341 & n23342 ;
  assign n23344 = n1312 & ~n23343 ;
  assign n23345 = n9714 ^ n1707 ^ 1'b0 ;
  assign n23346 = ~n13998 & n23345 ;
  assign n23347 = n23344 & n23346 ;
  assign n23348 = n10950 & n23347 ;
  assign n23349 = n20445 & n21235 ;
  assign n23350 = n23349 ^ n8995 ^ 1'b0 ;
  assign n23351 = n5652 | n11336 ;
  assign n23352 = n23351 ^ n10637 ^ 1'b0 ;
  assign n23353 = ~n4137 & n6764 ;
  assign n23354 = n4312 ^ n1300 ^ 1'b0 ;
  assign n23355 = n16988 | n23354 ;
  assign n23356 = ( ~n9292 & n20252 ) | ( ~n9292 & n23355 ) | ( n20252 & n23355 ) ;
  assign n23357 = n18994 ^ n13031 ^ 1'b0 ;
  assign n23358 = ~n8338 & n23357 ;
  assign n23359 = n22616 ^ n10209 ^ 1'b0 ;
  assign n23360 = n13288 & n19777 ;
  assign n23361 = n1993 & n23360 ;
  assign n23362 = n1191 & n23361 ;
  assign n23363 = n10845 ^ n10404 ^ 1'b0 ;
  assign n23364 = n19489 ^ n8007 ^ 1'b0 ;
  assign n23365 = ~n23363 & n23364 ;
  assign n23366 = n21751 & n23365 ;
  assign n23367 = n23366 ^ n5249 ^ 1'b0 ;
  assign n23368 = n23367 ^ n7299 ^ 1'b0 ;
  assign n23369 = n23362 | n23368 ;
  assign n23370 = n6552 & ~n15467 ;
  assign n23373 = ( n2877 & ~n9884 ) | ( n2877 & n11772 ) | ( ~n9884 & n11772 ) ;
  assign n23371 = n21532 ^ n13359 ^ 1'b0 ;
  assign n23372 = n8931 | n23371 ;
  assign n23374 = n23373 ^ n23372 ^ 1'b0 ;
  assign n23375 = n8387 & ~n23374 ;
  assign n23376 = ~n2041 & n21079 ;
  assign n23377 = n23376 ^ n21884 ^ 1'b0 ;
  assign n23378 = n10626 | n23377 ;
  assign n23379 = n9245 | n23378 ;
  assign n23380 = ~n4559 & n8214 ;
  assign n23381 = n13213 ^ n1811 ^ 1'b0 ;
  assign n23382 = n3867 | n7627 ;
  assign n23383 = n1520 & ~n23382 ;
  assign n23384 = n12673 ^ n2435 ^ 1'b0 ;
  assign n23385 = n13303 & ~n23384 ;
  assign n23386 = n11099 & ~n19832 ;
  assign n23387 = n6408 & n23386 ;
  assign n23388 = n3177 & ~n4229 ;
  assign n23389 = ~n10804 & n23388 ;
  assign n23390 = ~n4668 & n23389 ;
  assign n23391 = ~n13061 & n23390 ;
  assign n23392 = n22714 ^ n3906 ^ 1'b0 ;
  assign n23393 = ~n4855 & n9855 ;
  assign n23394 = n7484 ^ n1351 ^ 1'b0 ;
  assign n23395 = n2109 | n23394 ;
  assign n23396 = n23395 ^ n8909 ^ 1'b0 ;
  assign n23397 = n1469 | n23396 ;
  assign n23398 = ( n714 & n9848 ) | ( n714 & ~n16458 ) | ( n9848 & ~n16458 ) ;
  assign n23399 = n23398 ^ n966 ^ 1'b0 ;
  assign n23400 = n12575 ^ n4056 ^ 1'b0 ;
  assign n23401 = n6383 ^ n1857 ^ 1'b0 ;
  assign n23402 = ~n16096 & n23401 ;
  assign n23403 = n13167 & n23402 ;
  assign n23404 = n8613 | n23008 ;
  assign n23405 = n23403 & n23404 ;
  assign n23409 = ~n1329 & n1476 ;
  assign n23410 = ~n1476 & n23409 ;
  assign n23406 = ~n5758 & n14509 ;
  assign n23407 = n5758 & n23406 ;
  assign n23408 = n1080 & ~n23407 ;
  assign n23411 = n23410 ^ n23408 ^ 1'b0 ;
  assign n23412 = n1200 & n2199 ;
  assign n23413 = ~n1200 & n23412 ;
  assign n23414 = n1495 & n23413 ;
  assign n23415 = ~n2730 & n23414 ;
  assign n23416 = n548 & n23415 ;
  assign n23417 = n8970 | n23416 ;
  assign n23418 = n11117 & n23417 ;
  assign n23419 = n10383 & n23418 ;
  assign n23420 = n13335 & ~n23419 ;
  assign n23421 = ~n23411 & n23420 ;
  assign n23422 = n448 & ~n4466 ;
  assign n23423 = ~n6027 & n23422 ;
  assign n23424 = n12856 | n23423 ;
  assign n23425 = n1521 & ~n12897 ;
  assign n23426 = n9873 ^ n192 ^ 1'b0 ;
  assign n23427 = n1454 | n2353 ;
  assign n23428 = ( n2610 & n23426 ) | ( n2610 & ~n23427 ) | ( n23426 & ~n23427 ) ;
  assign n23429 = ~n16604 & n16867 ;
  assign n23430 = n16343 & n23429 ;
  assign n23431 = n20216 ^ n9651 ^ n144 ;
  assign n23432 = n14824 & n23431 ;
  assign n23433 = n5610 | n6159 ;
  assign n23434 = n6551 & n23433 ;
  assign n23435 = ~n18933 & n23434 ;
  assign n23436 = n4860 ^ n1941 ^ 1'b0 ;
  assign n23437 = n23435 | n23436 ;
  assign n23438 = ~n7830 & n8260 ;
  assign n23439 = n15232 ^ n10158 ^ 1'b0 ;
  assign n23440 = ~n19498 & n23439 ;
  assign n23441 = n23438 & n23440 ;
  assign n23442 = n1551 & ~n3886 ;
  assign n23443 = n23442 ^ n6012 ^ 1'b0 ;
  assign n23444 = ( n924 & ~n17528 ) | ( n924 & n23443 ) | ( ~n17528 & n23443 ) ;
  assign n23445 = n6323 ^ n365 ^ 1'b0 ;
  assign n23446 = ~n13201 & n23445 ;
  assign n23447 = n3438 | n16474 ;
  assign n23448 = n23447 ^ n7861 ^ 1'b0 ;
  assign n23449 = ( n6802 & n20414 ) | ( n6802 & ~n23448 ) | ( n20414 & ~n23448 ) ;
  assign n23450 = ~n5037 & n23449 ;
  assign n23451 = n23450 ^ n3721 ^ 1'b0 ;
  assign n23453 = n8931 ^ n3833 ^ 1'b0 ;
  assign n23454 = ( n9365 & n18716 ) | ( n9365 & n23453 ) | ( n18716 & n23453 ) ;
  assign n23452 = n4504 & ~n11353 ;
  assign n23455 = n23454 ^ n23452 ^ 1'b0 ;
  assign n23456 = n9732 ^ n4595 ^ n3966 ;
  assign n23457 = n17318 | n23456 ;
  assign n23458 = ~n489 & n11518 ;
  assign n23459 = ~n949 & n23458 ;
  assign n23460 = n6961 & ~n23459 ;
  assign n23461 = n14287 & n23460 ;
  assign n23463 = n1845 | n4750 ;
  assign n23464 = n4750 & ~n23463 ;
  assign n23465 = n18567 ^ n17189 ^ 1'b0 ;
  assign n23466 = ~n23464 & n23465 ;
  assign n23467 = n23466 ^ n3626 ^ 1'b0 ;
  assign n23462 = n7372 & ~n19757 ;
  assign n23468 = n23467 ^ n23462 ^ 1'b0 ;
  assign n23469 = n15764 ^ n7493 ^ 1'b0 ;
  assign n23470 = n9894 & ~n23469 ;
  assign n23471 = n2113 & n23470 ;
  assign n23472 = n7063 & n23471 ;
  assign n23473 = ~n1369 & n12106 ;
  assign n23474 = ~n14215 & n17256 ;
  assign n23475 = n9674 & ~n13108 ;
  assign n23476 = n23475 ^ n22846 ^ 1'b0 ;
  assign n23477 = n378 & ~n7402 ;
  assign n23478 = n23477 ^ n6796 ^ 1'b0 ;
  assign n23479 = n5965 ^ n4583 ^ 1'b0 ;
  assign n23480 = ~n454 & n23479 ;
  assign n23481 = n9244 ^ n6411 ^ 1'b0 ;
  assign n23482 = n644 & n13992 ;
  assign n23483 = n6261 & ~n22718 ;
  assign n23484 = ( n3011 & n23482 ) | ( n3011 & n23483 ) | ( n23482 & n23483 ) ;
  assign n23485 = n2094 | n3708 ;
  assign n23486 = n23485 ^ n615 ^ 1'b0 ;
  assign n23487 = n23486 ^ n14315 ^ 1'b0 ;
  assign n23488 = ~n13843 & n23487 ;
  assign n23489 = n10708 ^ n2864 ^ 1'b0 ;
  assign n23490 = n23488 & ~n23489 ;
  assign n23491 = n18538 & ~n23490 ;
  assign n23492 = ~n18770 & n18778 ;
  assign n23493 = ~n23491 & n23492 ;
  assign n23494 = n625 & n2886 ;
  assign n23495 = n2288 & n23494 ;
  assign n23496 = n5658 | n23495 ;
  assign n23497 = n23496 ^ n22499 ^ 1'b0 ;
  assign n23498 = n7007 | n23497 ;
  assign n23499 = n23498 ^ n21449 ^ 1'b0 ;
  assign n23500 = n23493 | n23499 ;
  assign n23502 = ~n1582 & n1744 ;
  assign n23503 = ~n1744 & n23502 ;
  assign n23501 = n2539 | n7735 ;
  assign n23504 = n23503 ^ n23501 ^ 1'b0 ;
  assign n23505 = n1590 & n23504 ;
  assign n23506 = ~n2463 & n9505 ;
  assign n23507 = n2186 & ~n23506 ;
  assign n23508 = n12951 & n23507 ;
  assign n23509 = n7753 | n12455 ;
  assign n23510 = ( n1944 & n4741 ) | ( n1944 & ~n23509 ) | ( n4741 & ~n23509 ) ;
  assign n23511 = n20911 | n23510 ;
  assign n23512 = n23511 ^ n22966 ^ 1'b0 ;
  assign n23513 = n13361 | n23512 ;
  assign n23514 = n23513 ^ n10735 ^ 1'b0 ;
  assign n23515 = n908 | n14425 ;
  assign n23516 = n6224 | n23515 ;
  assign n23517 = ~n17976 & n23516 ;
  assign n23518 = ( ~n1853 & n7265 ) | ( ~n1853 & n23517 ) | ( n7265 & n23517 ) ;
  assign n23519 = n724 | n7046 ;
  assign n23520 = n23519 ^ n12551 ^ 1'b0 ;
  assign n23521 = ~n6779 & n7100 ;
  assign n23522 = n14426 & n23521 ;
  assign n23523 = ~n23520 & n23522 ;
  assign n23524 = n23207 & n23523 ;
  assign n23525 = n2929 & ~n8975 ;
  assign n23526 = n15559 ^ n3993 ^ 1'b0 ;
  assign n23527 = n6568 | n23526 ;
  assign n23528 = n21878 ^ n10612 ^ 1'b0 ;
  assign n23529 = ~n23527 & n23528 ;
  assign n23530 = n15796 ^ n13879 ^ 1'b0 ;
  assign n23531 = n23530 ^ n17303 ^ 1'b0 ;
  assign n23532 = n3133 & n22601 ;
  assign n23533 = n11123 ^ n8549 ^ 1'b0 ;
  assign n23534 = n23533 ^ n6866 ^ 1'b0 ;
  assign n23535 = n13613 & ~n18268 ;
  assign n23536 = n23534 & n23535 ;
  assign n23537 = n23532 & ~n23536 ;
  assign n23538 = n6296 & ~n19755 ;
  assign n23539 = n23538 ^ n9210 ^ 1'b0 ;
  assign n23540 = n4568 & n9877 ;
  assign n23543 = ~n4849 & n14949 ;
  assign n23541 = n8660 ^ n6335 ^ n254 ;
  assign n23542 = n8710 | n23541 ;
  assign n23544 = n23543 ^ n23542 ^ 1'b0 ;
  assign n23545 = n12804 ^ n12271 ^ 1'b0 ;
  assign n23546 = n14867 & n23545 ;
  assign n23547 = n23546 ^ n2853 ^ 1'b0 ;
  assign n23548 = n985 & n9264 ;
  assign n23549 = n23548 ^ n2719 ^ 1'b0 ;
  assign n23556 = ~n5731 & n12799 ;
  assign n23550 = n5397 & ~n20969 ;
  assign n23551 = ~n3271 & n8040 ;
  assign n23552 = ~n5463 & n23551 ;
  assign n23553 = n23552 ^ n8497 ^ n6001 ;
  assign n23554 = n23553 ^ n13855 ^ 1'b0 ;
  assign n23555 = n23550 | n23554 ;
  assign n23557 = n23556 ^ n23555 ^ 1'b0 ;
  assign n23559 = n15590 ^ n9323 ^ 1'b0 ;
  assign n23560 = n7781 & ~n23559 ;
  assign n23558 = ( n3858 & n4097 ) | ( n3858 & ~n4194 ) | ( n4097 & ~n4194 ) ;
  assign n23561 = n23560 ^ n23558 ^ 1'b0 ;
  assign n23562 = ~n9983 & n23561 ;
  assign n23563 = n23562 ^ n21259 ^ 1'b0 ;
  assign n23564 = n18435 ^ n9608 ^ 1'b0 ;
  assign n23565 = n11064 | n18902 ;
  assign n23566 = n5961 & ~n23565 ;
  assign n23567 = ~n602 & n12496 ;
  assign n23568 = n695 & n23444 ;
  assign n23570 = n4351 | n5313 ;
  assign n23569 = n17873 ^ n4945 ^ 1'b0 ;
  assign n23571 = n23570 ^ n23569 ^ 1'b0 ;
  assign n23572 = n3818 & ~n9771 ;
  assign n23573 = n20060 & ~n23572 ;
  assign n23574 = n13080 & n20954 ;
  assign n23575 = ~n23573 & n23574 ;
  assign n23576 = n3090 & ~n14047 ;
  assign n23577 = n23576 ^ n2324 ^ 1'b0 ;
  assign n23578 = n23577 ^ n23286 ^ 1'b0 ;
  assign n23579 = ~n3772 & n23578 ;
  assign n23580 = n23579 ^ n28 ^ 1'b0 ;
  assign n23581 = n12281 ^ n8003 ^ 1'b0 ;
  assign n23582 = ~n22658 & n23581 ;
  assign n23583 = n2225 & ~n4408 ;
  assign n23584 = n23583 ^ n620 ^ 1'b0 ;
  assign n23585 = ~n2510 & n23584 ;
  assign n23586 = n20539 ^ n17718 ^ 1'b0 ;
  assign n23587 = n3536 & n17065 ;
  assign n23588 = ~n4833 & n16010 ;
  assign n23592 = n15114 ^ n4685 ^ n3494 ;
  assign n23589 = n7904 & ~n18291 ;
  assign n23590 = n453 & n23589 ;
  assign n23591 = n19551 & ~n23590 ;
  assign n23593 = n23592 ^ n23591 ^ 1'b0 ;
  assign n23594 = ~n51 & n15771 ;
  assign n23595 = n23594 ^ n2336 ^ 1'b0 ;
  assign n23596 = n12989 ^ n7830 ^ 1'b0 ;
  assign n23597 = n23595 | n23596 ;
  assign n23598 = n1395 & n14227 ;
  assign n23599 = n12690 & ~n18683 ;
  assign n23600 = n3674 | n19663 ;
  assign n23601 = n23600 ^ n22101 ^ 1'b0 ;
  assign n23602 = ~n328 & n23601 ;
  assign n23603 = n23602 ^ n11182 ^ 1'b0 ;
  assign n23604 = n14177 | n23603 ;
  assign n23605 = n3428 ^ n961 ^ 1'b0 ;
  assign n23606 = ( n14275 & ~n14525 ) | ( n14275 & n23605 ) | ( ~n14525 & n23605 ) ;
  assign n23607 = n23606 ^ n5364 ^ 1'b0 ;
  assign n23608 = n956 | n11021 ;
  assign n23609 = n23608 ^ n3854 ^ 1'b0 ;
  assign n23610 = n5385 & ~n23609 ;
  assign n23611 = n8230 | n17362 ;
  assign n23612 = n8446 & n11477 ;
  assign n23613 = n2114 | n2745 ;
  assign n23614 = n23613 ^ n773 ^ 1'b0 ;
  assign n23615 = n21888 & ~n23614 ;
  assign n23616 = n23615 ^ n9499 ^ 1'b0 ;
  assign n23617 = n7493 ^ n5253 ^ n3849 ;
  assign n23618 = ~n5284 & n6667 ;
  assign n23619 = n23618 ^ n3414 ^ 1'b0 ;
  assign n23620 = ~n592 & n4105 ;
  assign n23621 = ( n11206 & ~n15252 ) | ( n11206 & n23620 ) | ( ~n15252 & n23620 ) ;
  assign n23622 = n19889 ^ n15075 ^ 1'b0 ;
  assign n23623 = n23621 & n23622 ;
  assign n23624 = ~n3996 & n4720 ;
  assign n23625 = n3054 | n9216 ;
  assign n23629 = ~n6857 & n9022 ;
  assign n23630 = ~n22286 & n23629 ;
  assign n23626 = ~n506 & n12526 ;
  assign n23627 = ~n20716 & n23626 ;
  assign n23628 = n5647 & ~n23627 ;
  assign n23631 = n23630 ^ n23628 ^ 1'b0 ;
  assign n23632 = ~n18919 & n23156 ;
  assign n23634 = n6585 ^ n792 ^ 1'b0 ;
  assign n23635 = ~n638 & n23634 ;
  assign n23633 = n22073 ^ n1476 ^ 1'b0 ;
  assign n23636 = n23635 ^ n23633 ^ 1'b0 ;
  assign n23637 = n20919 & ~n23636 ;
  assign n23638 = n23632 & n23637 ;
  assign n23639 = n20525 ^ n4293 ^ 1'b0 ;
  assign n23641 = n9000 & n14275 ;
  assign n23642 = n8497 ^ n889 ^ 1'b0 ;
  assign n23643 = n88 | n23642 ;
  assign n23644 = n23641 | n23643 ;
  assign n23640 = x1 & ~n18132 ;
  assign n23645 = n23644 ^ n23640 ^ 1'b0 ;
  assign n23646 = n21268 | n23645 ;
  assign n23647 = n3307 ^ x0 ^ 1'b0 ;
  assign n23648 = ~x6 & n23647 ;
  assign n23649 = ( n2277 & n20325 ) | ( n2277 & n23648 ) | ( n20325 & n23648 ) ;
  assign n23655 = n15885 ^ n2494 ^ 1'b0 ;
  assign n23650 = ( n1517 & n7083 ) | ( n1517 & n14787 ) | ( n7083 & n14787 ) ;
  assign n23651 = n7955 & ~n20604 ;
  assign n23652 = n12713 & n23651 ;
  assign n23653 = n23652 ^ n4005 ^ 1'b0 ;
  assign n23654 = ( n8436 & n23650 ) | ( n8436 & n23653 ) | ( n23650 & n23653 ) ;
  assign n23656 = n23655 ^ n23654 ^ 1'b0 ;
  assign n23657 = n4470 ^ n4366 ^ 1'b0 ;
  assign n23658 = ~n1436 & n23657 ;
  assign n23659 = n23658 ^ n13597 ^ 1'b0 ;
  assign n23660 = ~n5511 & n17513 ;
  assign n23661 = n4139 & n23660 ;
  assign n23662 = n2494 & n2974 ;
  assign n23663 = n23662 ^ n4349 ^ 1'b0 ;
  assign n23664 = n12988 & ~n16137 ;
  assign n23665 = ~n2147 & n6945 ;
  assign n23666 = n11768 ^ n10819 ^ 1'b0 ;
  assign n23667 = n14652 ^ n6839 ^ 1'b0 ;
  assign n23668 = n23667 ^ n9630 ^ 1'b0 ;
  assign n23671 = n3639 ^ n2802 ^ 1'b0 ;
  assign n23672 = n20050 & ~n23671 ;
  assign n23669 = n667 & ~n10181 ;
  assign n23670 = n23669 ^ n7802 ^ 1'b0 ;
  assign n23673 = n23672 ^ n23670 ^ n11795 ;
  assign n23674 = ( n11447 & ~n15784 ) | ( n11447 & n23673 ) | ( ~n15784 & n23673 ) ;
  assign n23675 = ~n7806 & n9346 ;
  assign n23676 = n12981 | n23675 ;
  assign n23677 = n10331 | n23676 ;
  assign n23678 = n23677 ^ n2202 ^ 1'b0 ;
  assign n23679 = n11389 & n23678 ;
  assign n23680 = ~n20032 & n23679 ;
  assign n23681 = n915 | n1369 ;
  assign n23682 = n7270 & ~n23681 ;
  assign n23685 = n8373 & ~n13891 ;
  assign n23683 = ( n12696 & n15557 ) | ( n12696 & n16683 ) | ( n15557 & n16683 ) ;
  assign n23684 = n10121 | n23683 ;
  assign n23686 = n23685 ^ n23684 ^ 1'b0 ;
  assign n23687 = n18477 ^ n14038 ^ 1'b0 ;
  assign n23688 = ~n10309 & n23687 ;
  assign n23689 = n18685 & n23688 ;
  assign n23690 = n23689 ^ n5591 ^ 1'b0 ;
  assign n23691 = n17181 ^ n14887 ^ 1'b0 ;
  assign n23692 = ~n49 & n20144 ;
  assign n23693 = n2721 ^ n131 ^ 1'b0 ;
  assign n23694 = ( ~n8181 & n13358 ) | ( ~n8181 & n23693 ) | ( n13358 & n23693 ) ;
  assign n23695 = n23694 ^ n5107 ^ 1'b0 ;
  assign n23696 = n3218 | n8598 ;
  assign n23697 = n1618 & ~n9260 ;
  assign n23698 = n11021 & n23697 ;
  assign n23699 = ( ~n627 & n6271 ) | ( ~n627 & n15660 ) | ( n6271 & n15660 ) ;
  assign n23700 = ~n23698 & n23699 ;
  assign n23710 = n7926 | n9748 ;
  assign n23711 = n8258 & ~n23710 ;
  assign n23701 = n12807 ^ n12422 ^ n5204 ;
  assign n23702 = n6333 ^ n207 ^ 1'b0 ;
  assign n23703 = n4018 | n23702 ;
  assign n23704 = n2202 & n14728 ;
  assign n23705 = n5791 & n23704 ;
  assign n23706 = n8020 | n23705 ;
  assign n23707 = n23703 & ~n23706 ;
  assign n23708 = n23707 ^ n6538 ^ n5099 ;
  assign n23709 = n23701 & n23708 ;
  assign n23712 = n23711 ^ n23709 ^ 1'b0 ;
  assign n23714 = n4378 ^ n2580 ^ 1'b0 ;
  assign n23713 = n4837 & ~n18513 ;
  assign n23715 = n23714 ^ n23713 ^ 1'b0 ;
  assign n23716 = n14739 ^ n4139 ^ 1'b0 ;
  assign n23717 = n9024 ^ n4567 ^ 1'b0 ;
  assign n23718 = n5046 & ~n14220 ;
  assign n23719 = n20667 ^ n14358 ^ 1'b0 ;
  assign n23720 = n9928 ^ n3132 ^ 1'b0 ;
  assign n23722 = ~n169 & n982 ;
  assign n23723 = n4068 & n8287 ;
  assign n23724 = n5795 & n23723 ;
  assign n23725 = ( ~n9022 & n23722 ) | ( ~n9022 & n23724 ) | ( n23722 & n23724 ) ;
  assign n23721 = n11199 ^ n9908 ^ n4575 ;
  assign n23726 = n23725 ^ n23721 ^ n16941 ;
  assign n23727 = n5194 & n10854 ;
  assign n23728 = n4200 & n23727 ;
  assign n23729 = n23728 ^ n1029 ^ 1'b0 ;
  assign n23730 = n4259 & ~n20067 ;
  assign n23731 = n4009 & ~n23730 ;
  assign n23733 = ~n9117 & n15777 ;
  assign n23732 = ~n7786 & n16190 ;
  assign n23734 = n23733 ^ n23732 ^ 1'b0 ;
  assign n23737 = n10751 ^ n5344 ^ 1'b0 ;
  assign n23738 = n1497 & ~n23737 ;
  assign n23735 = ~n911 & n3147 ;
  assign n23736 = n23735 ^ n9481 ^ 1'b0 ;
  assign n23739 = n23738 ^ n23736 ^ n2445 ;
  assign n23740 = ~n11295 & n20954 ;
  assign n23741 = n23740 ^ n2148 ^ 1'b0 ;
  assign n23742 = n15376 | n22769 ;
  assign n23743 = n19225 ^ n8080 ^ 1'b0 ;
  assign n23744 = ( n6035 & n7263 ) | ( n6035 & n23743 ) | ( n7263 & n23743 ) ;
  assign n23745 = n10257 & n11731 ;
  assign n23746 = n23745 ^ n5984 ^ 1'b0 ;
  assign n23747 = n20607 & n23746 ;
  assign n23748 = ~n9321 & n10207 ;
  assign n23749 = ~n6594 & n23748 ;
  assign n23750 = n1207 | n6584 ;
  assign n23751 = n23750 ^ n5586 ^ 1'b0 ;
  assign n23752 = ~n10846 & n23751 ;
  assign n23753 = n23749 & n23752 ;
  assign n23754 = n8598 & ~n19215 ;
  assign n23755 = ~n4613 & n23754 ;
  assign n23756 = n23755 ^ n10793 ^ 1'b0 ;
  assign n23757 = n23756 ^ n4748 ^ 1'b0 ;
  assign n23758 = n23757 ^ n12561 ^ n10919 ;
  assign n23759 = n3937 | n4132 ;
  assign n23760 = n23759 ^ n6954 ^ 1'b0 ;
  assign n23761 = n155 & n23760 ;
  assign n23762 = n3025 & n23761 ;
  assign n23763 = n23758 & n23762 ;
  assign n23764 = n23753 & n23763 ;
  assign n23765 = n4533 & ~n5234 ;
  assign n23766 = n6179 & ~n14343 ;
  assign n23767 = n4326 & n23766 ;
  assign n23768 = ~n23765 & n23767 ;
  assign n23773 = n15765 ^ n1336 ^ 1'b0 ;
  assign n23774 = n11770 & n23773 ;
  assign n23775 = n14512 | n23774 ;
  assign n23769 = n6827 & ~n21583 ;
  assign n23770 = n23769 ^ n3565 ^ 1'b0 ;
  assign n23771 = n1408 & n17493 ;
  assign n23772 = ( ~n1212 & n23770 ) | ( ~n1212 & n23771 ) | ( n23770 & n23771 ) ;
  assign n23776 = n23775 ^ n23772 ^ 1'b0 ;
  assign n23777 = n7531 | n23776 ;
  assign n23778 = n10527 & n23023 ;
  assign n23779 = n5730 | n15011 ;
  assign n23780 = n6937 | n9290 ;
  assign n23781 = ~n19438 & n23780 ;
  assign n23782 = n10042 | n10745 ;
  assign n23783 = n6155 | n23782 ;
  assign n23784 = n387 & n8084 ;
  assign n23785 = n19421 & n23784 ;
  assign n23786 = ( n67 & n4519 ) | ( n67 & ~n23785 ) | ( n4519 & ~n23785 ) ;
  assign n23787 = n6891 ^ n5320 ^ 1'b0 ;
  assign n23788 = ~n23786 & n23787 ;
  assign n23789 = ~n4831 & n7170 ;
  assign n23790 = n23789 ^ n3539 ^ 1'b0 ;
  assign n23791 = n11454 ^ n9827 ^ 1'b0 ;
  assign n23792 = ( ~n20533 & n23790 ) | ( ~n20533 & n23791 ) | ( n23790 & n23791 ) ;
  assign n23793 = ( n159 & n737 ) | ( n159 & ~n6589 ) | ( n737 & ~n6589 ) ;
  assign n23794 = n23793 ^ n4089 ^ n1419 ;
  assign n23795 = n659 & ~n13998 ;
  assign n23797 = n4001 | n13404 ;
  assign n23798 = ( ~n2036 & n4510 ) | ( ~n2036 & n23797 ) | ( n4510 & n23797 ) ;
  assign n23796 = ~n5369 & n23449 ;
  assign n23799 = n23798 ^ n23796 ^ 1'b0 ;
  assign n23800 = n22285 ^ n7335 ^ 1'b0 ;
  assign n23801 = n6794 & ~n23800 ;
  assign n23802 = n6738 & n11384 ;
  assign n23803 = n4655 & n23802 ;
  assign n23804 = n652 ^ n625 ^ 1'b0 ;
  assign n23805 = ~n23803 & n23804 ;
  assign n23806 = n11954 ^ n8821 ^ 1'b0 ;
  assign n23807 = n1092 & ~n23806 ;
  assign n23808 = n23807 ^ n2621 ^ 1'b0 ;
  assign n23809 = n23808 ^ n2899 ^ 1'b0 ;
  assign n23810 = ~n2032 & n23809 ;
  assign n23811 = n8197 | n23810 ;
  assign n23812 = n1649 | n16501 ;
  assign n23813 = n23811 & n23812 ;
  assign n23814 = n23813 ^ n10361 ^ 1'b0 ;
  assign n23815 = n931 & ~n11380 ;
  assign n23816 = n23815 ^ n2417 ^ 1'b0 ;
  assign n23817 = n23816 ^ n3483 ^ 1'b0 ;
  assign n23818 = n9664 & n15342 ;
  assign n23819 = n23817 & n23818 ;
  assign n23820 = ~n19472 & n19494 ;
  assign n23821 = ~n10508 & n23820 ;
  assign n23822 = n1352 | n23821 ;
  assign n23823 = ~n2735 & n4311 ;
  assign n23824 = n23823 ^ n17403 ^ 1'b0 ;
  assign n23825 = n23824 ^ n6797 ^ 1'b0 ;
  assign n23826 = n9002 ^ n648 ^ 1'b0 ;
  assign n23827 = n13176 ^ n2131 ^ 1'b0 ;
  assign n23828 = n23827 ^ n13871 ^ 1'b0 ;
  assign n23829 = n1205 & ~n17191 ;
  assign n23830 = n4030 ^ n1205 ^ 1'b0 ;
  assign n23831 = ( n699 & ~n3919 ) | ( n699 & n17178 ) | ( ~n3919 & n17178 ) ;
  assign n23832 = ~n13245 & n23831 ;
  assign n23833 = n3349 & n12817 ;
  assign n23834 = n9912 ^ n8194 ^ n4145 ;
  assign n23835 = n9249 ^ n4986 ^ 1'b0 ;
  assign n23836 = n1867 | n23835 ;
  assign n23837 = n2738 & ~n23836 ;
  assign n23838 = n23837 ^ n787 ^ 1'b0 ;
  assign n23839 = n23834 & n23838 ;
  assign n23840 = n19892 ^ n9754 ^ 1'b0 ;
  assign n23841 = ~n23839 & n23840 ;
  assign n23842 = n2796 & n11759 ;
  assign n23843 = n23842 ^ n15519 ^ 1'b0 ;
  assign n23844 = n14368 & ~n16809 ;
  assign n23845 = n23843 & n23844 ;
  assign n23846 = n5692 & ~n13968 ;
  assign n23847 = n23846 ^ n18876 ^ 1'b0 ;
  assign n23848 = ~n1935 & n7016 ;
  assign n23849 = n23848 ^ n16144 ^ 1'b0 ;
  assign n23850 = n16174 ^ n12030 ^ 1'b0 ;
  assign n23851 = ~n20608 & n23850 ;
  assign n23852 = ( n6500 & n12084 ) | ( n6500 & n16055 ) | ( n12084 & n16055 ) ;
  assign n23856 = n924 & ~n1054 ;
  assign n23853 = n5580 | n6255 ;
  assign n23854 = n23853 ^ n15818 ^ 1'b0 ;
  assign n23855 = n3906 & ~n23854 ;
  assign n23857 = n23856 ^ n23855 ^ 1'b0 ;
  assign n23858 = n23852 | n23857 ;
  assign n23859 = n6472 & ~n23858 ;
  assign n23860 = n3239 & n5165 ;
  assign n23861 = ~n23859 & n23860 ;
  assign n23862 = n2785 & ~n12832 ;
  assign n23863 = n2905 | n20833 ;
  assign n23864 = n23863 ^ n2465 ^ 1'b0 ;
  assign n23865 = ~n611 & n8928 ;
  assign n23866 = n23865 ^ n2403 ^ 1'b0 ;
  assign n23867 = n16702 & n23866 ;
  assign n23868 = n8893 ^ n1573 ^ 1'b0 ;
  assign n23869 = n23868 ^ n4418 ^ 1'b0 ;
  assign n23870 = ~n5638 & n8745 ;
  assign n23871 = n23870 ^ n7023 ^ 1'b0 ;
  assign n23872 = n23871 ^ n13119 ^ 1'b0 ;
  assign n23873 = n23872 ^ n13789 ^ n3902 ;
  assign n23874 = ~n5001 & n7185 ;
  assign n23877 = n667 & n7160 ;
  assign n23875 = n9944 ^ n6200 ^ n86 ;
  assign n23876 = n14217 & ~n23875 ;
  assign n23878 = n23877 ^ n23876 ^ 1'b0 ;
  assign n23879 = ~n7396 & n23459 ;
  assign n23880 = n12475 ^ n4646 ^ 1'b0 ;
  assign n23881 = n309 | n4698 ;
  assign n23882 = n23880 & ~n23881 ;
  assign n23883 = n1329 & n5475 ;
  assign n23884 = ( n3064 & n9279 ) | ( n3064 & ~n23883 ) | ( n9279 & ~n23883 ) ;
  assign n23885 = n23884 ^ n2532 ^ 1'b0 ;
  assign n23886 = n6528 & ~n23885 ;
  assign n23887 = n23886 ^ n4132 ^ 1'b0 ;
  assign n23888 = n2140 | n23887 ;
  assign n23889 = n14198 ^ n10935 ^ 1'b0 ;
  assign n23892 = n20127 ^ n6904 ^ 1'b0 ;
  assign n23890 = n12389 & n13318 ;
  assign n23891 = n23890 ^ n14297 ^ 1'b0 ;
  assign n23893 = n23892 ^ n23891 ^ 1'b0 ;
  assign n23894 = n16725 & ~n23893 ;
  assign n23895 = n2899 & n3630 ;
  assign n23896 = n23895 ^ n13422 ^ 1'b0 ;
  assign n23897 = ( n942 & n11123 ) | ( n942 & ~n15076 ) | ( n11123 & ~n15076 ) ;
  assign n23898 = n23897 ^ n20068 ^ n3713 ;
  assign n23899 = n23898 ^ n14177 ^ 1'b0 ;
  assign n23900 = n2847 & n4645 ;
  assign n23901 = n6119 & n23900 ;
  assign n23902 = n4422 | n23901 ;
  assign n23903 = n1853 & ~n23306 ;
  assign n23904 = n3040 & n23903 ;
  assign n23905 = n7522 ^ n4903 ^ 1'b0 ;
  assign n23906 = n14362 ^ n7033 ^ 1'b0 ;
  assign n23907 = n18732 & n23906 ;
  assign n23908 = n1598 & ~n3510 ;
  assign n23909 = n23908 ^ n11407 ^ 1'b0 ;
  assign n23910 = n14417 ^ n98 ^ 1'b0 ;
  assign n23911 = n16925 ^ n13589 ^ 1'b0 ;
  assign n23912 = ( n36 & ~n11214 ) | ( n36 & n21469 ) | ( ~n11214 & n21469 ) ;
  assign n23913 = n9258 ^ n642 ^ 1'b0 ;
  assign n23914 = ~n5149 & n5445 ;
  assign n23915 = n6912 & n23914 ;
  assign n23916 = n2211 & ~n23915 ;
  assign n23917 = n4332 ^ n2068 ^ 1'b0 ;
  assign n23918 = n7023 ^ n5328 ^ 1'b0 ;
  assign n23919 = n13174 | n23918 ;
  assign n23920 = n1511 ^ n1223 ^ 1'b0 ;
  assign n23921 = n2925 & ~n7601 ;
  assign n23922 = ~n5676 & n23921 ;
  assign n23923 = n23920 & ~n23922 ;
  assign n23924 = n23923 ^ n13578 ^ 1'b0 ;
  assign n23925 = n23919 | n23924 ;
  assign n23926 = n22274 ^ n17320 ^ 1'b0 ;
  assign n23927 = n347 | n2619 ;
  assign n23928 = n23927 ^ n18393 ^ 1'b0 ;
  assign n23929 = n21334 & n23928 ;
  assign n23930 = n2094 | n6838 ;
  assign n23931 = n23930 ^ n6980 ^ 1'b0 ;
  assign n23932 = n14575 ^ n4136 ^ 1'b0 ;
  assign n23933 = n23932 ^ n14753 ^ 1'b0 ;
  assign n23934 = n23931 & ~n23933 ;
  assign n23935 = n562 | n2260 ;
  assign n23936 = n9111 | n23935 ;
  assign n23937 = n4253 | n8171 ;
  assign n23938 = n23937 ^ n12695 ^ 1'b0 ;
  assign n23939 = n9033 & n23938 ;
  assign n23940 = n23936 & n23939 ;
  assign n23941 = ~n3233 & n23940 ;
  assign n23942 = n20228 ^ n11046 ^ 1'b0 ;
  assign n23943 = ~n23941 & n23942 ;
  assign n23944 = n2550 & n4949 ;
  assign n23945 = n23944 ^ n19074 ^ n2350 ;
  assign n23948 = n18232 ^ n1771 ^ 1'b0 ;
  assign n23946 = n7648 ^ n5684 ^ 1'b0 ;
  assign n23947 = n1165 & ~n23946 ;
  assign n23949 = n23948 ^ n23947 ^ 1'b0 ;
  assign n23950 = ( ~n796 & n3724 ) | ( ~n796 & n23949 ) | ( n3724 & n23949 ) ;
  assign n23951 = n23950 ^ n9765 ^ 1'b0 ;
  assign n23952 = n17251 ^ n8109 ^ n1540 ;
  assign n23953 = n13056 ^ n10701 ^ 1'b0 ;
  assign n23954 = n23953 ^ n8313 ^ n936 ;
  assign n23955 = n8270 | n12849 ;
  assign n23956 = n23092 & ~n23955 ;
  assign n23957 = n23956 ^ n6179 ^ 1'b0 ;
  assign n23958 = ~n1083 & n10500 ;
  assign n23959 = n5175 & n23958 ;
  assign n23960 = ~n2682 & n23959 ;
  assign n23961 = n5522 ^ n3826 ^ n3261 ;
  assign n23962 = ~n7741 & n7899 ;
  assign n23963 = n23962 ^ n19278 ^ 1'b0 ;
  assign n23964 = ~n17052 & n23963 ;
  assign n23965 = n23964 ^ n5123 ^ 1'b0 ;
  assign n23966 = n8670 & ~n10223 ;
  assign n23967 = n4712 | n23966 ;
  assign n23968 = n23967 ^ n18873 ^ 1'b0 ;
  assign n23969 = n19546 ^ n16923 ^ n508 ;
  assign n23970 = n21420 | n23969 ;
  assign n23971 = n10592 | n23970 ;
  assign n23972 = n16317 ^ n12614 ^ 1'b0 ;
  assign n23973 = n9274 | n23972 ;
  assign n23974 = n18830 | n23746 ;
  assign n23975 = n23746 & ~n23974 ;
  assign n23976 = n703 & ~n1571 ;
  assign n23977 = n23976 ^ n13062 ^ 1'b0 ;
  assign n23978 = ( n7884 & n11534 ) | ( n7884 & n23977 ) | ( n11534 & n23977 ) ;
  assign n24001 = n785 & n2206 ;
  assign n24002 = ~n2206 & n24001 ;
  assign n24003 = n24002 ^ n574 ^ 1'b0 ;
  assign n23979 = n559 & ~n2205 ;
  assign n23980 = ~n559 & n23979 ;
  assign n23981 = n1401 | n1499 ;
  assign n23982 = n490 | n878 ;
  assign n23983 = n490 & ~n23982 ;
  assign n23984 = n988 | n23983 ;
  assign n23985 = n23983 & ~n23984 ;
  assign n23986 = ~n23981 & n23985 ;
  assign n23987 = n588 | n724 ;
  assign n23988 = n588 & ~n23987 ;
  assign n23989 = n23988 ^ n214 ^ 1'b0 ;
  assign n23990 = n23986 & ~n23989 ;
  assign n23991 = n135 & n23990 ;
  assign n23992 = n1845 & ~n23991 ;
  assign n23993 = n23980 & n23992 ;
  assign n23994 = n902 & ~n2872 ;
  assign n23995 = ~n902 & n23994 ;
  assign n23996 = n1285 & n3607 ;
  assign n23997 = n23996 ^ n16236 ^ 1'b0 ;
  assign n23998 = ~n23995 & n23997 ;
  assign n23999 = n23995 & n23998 ;
  assign n24000 = n23993 | n23999 ;
  assign n24004 = n24003 ^ n24000 ^ 1'b0 ;
  assign n24005 = n5918 & n10586 ;
  assign n24006 = n24005 ^ n749 ^ 1'b0 ;
  assign n24007 = ( ~n10805 & n16055 ) | ( ~n10805 & n24006 ) | ( n16055 & n24006 ) ;
  assign n24008 = n11813 ^ n2332 ^ 1'b0 ;
  assign n24009 = n24008 ^ n2328 ^ 1'b0 ;
  assign n24010 = ~n1747 & n4026 ;
  assign n24011 = ~n16197 & n24010 ;
  assign n24012 = n15532 & ~n19836 ;
  assign n24013 = n24012 ^ n21559 ^ 1'b0 ;
  assign n24015 = ~n1109 & n4182 ;
  assign n24014 = n675 | n23490 ;
  assign n24016 = n24015 ^ n24014 ^ n14309 ;
  assign n24017 = n15671 & n22013 ;
  assign n24018 = n582 | n10724 ;
  assign n24019 = n655 | n24018 ;
  assign n24020 = n23329 ^ n2923 ^ 1'b0 ;
  assign n24021 = n1246 & n7154 ;
  assign n24022 = n8258 & n24021 ;
  assign n24023 = n24022 ^ n7156 ^ 1'b0 ;
  assign n24024 = n970 | n1456 ;
  assign n24025 = n24023 & ~n24024 ;
  assign n24026 = n12393 | n20525 ;
  assign n24027 = n24026 ^ n3413 ^ 1'b0 ;
  assign n24028 = n5505 & n24027 ;
  assign n24029 = n24028 ^ n11374 ^ 1'b0 ;
  assign n24030 = ( n3037 & n3547 ) | ( n3037 & ~n4782 ) | ( n3547 & ~n4782 ) ;
  assign n24031 = n3520 ^ n3479 ^ 1'b0 ;
  assign n24032 = ~n21981 & n24031 ;
  assign n24033 = ~n506 & n7233 ;
  assign n24034 = n24033 ^ n920 ^ 1'b0 ;
  assign n24035 = ~n4082 & n24034 ;
  assign n24036 = ( n7312 & ~n8448 ) | ( n7312 & n13741 ) | ( ~n8448 & n13741 ) ;
  assign n24037 = n24035 & n24036 ;
  assign n24038 = n24037 ^ n4624 ^ 1'b0 ;
  assign n24039 = n13274 ^ n13046 ^ n7057 ;
  assign n24043 = ~n8042 & n21271 ;
  assign n24044 = n24043 ^ n8989 ^ 1'b0 ;
  assign n24040 = ~n4871 & n9540 ;
  assign n24041 = n12337 | n24040 ;
  assign n24042 = ~n38 & n24041 ;
  assign n24045 = n24044 ^ n24042 ^ 1'b0 ;
  assign n24046 = n6522 & ~n17535 ;
  assign n24047 = n4599 ^ n2228 ^ 1'b0 ;
  assign n24048 = n8173 ^ n1327 ^ 1'b0 ;
  assign n24049 = n3023 & ~n20364 ;
  assign n24050 = n2923 & n15554 ;
  assign n24051 = n16010 ^ n8216 ^ 1'b0 ;
  assign n24052 = ~n19151 & n24051 ;
  assign n24053 = n24052 ^ n5279 ^ 1'b0 ;
  assign n24054 = n1546 & ~n3907 ;
  assign n24055 = n24054 ^ n17035 ^ 1'b0 ;
  assign n24056 = n1422 & ~n3102 ;
  assign n24057 = ~n600 & n24056 ;
  assign n24058 = n20463 ^ n4209 ^ 1'b0 ;
  assign n24059 = n4197 | n24058 ;
  assign n24060 = n2522 | n24059 ;
  assign n24061 = n2101 | n24060 ;
  assign n24062 = n1276 & n20302 ;
  assign n24063 = n24062 ^ n6610 ^ 1'b0 ;
  assign n24064 = ~n3231 & n21849 ;
  assign n24065 = ~n5036 & n24064 ;
  assign n24066 = n4785 & ~n24065 ;
  assign n24067 = n12297 ^ n5395 ^ 1'b0 ;
  assign n24068 = n2812 & ~n5626 ;
  assign n24069 = n24068 ^ n11661 ^ 1'b0 ;
  assign n24070 = n2155 | n8043 ;
  assign n24071 = n24070 ^ n9373 ^ 1'b0 ;
  assign n24072 = ~n52 & n24071 ;
  assign n24073 = n10554 ^ n2630 ^ 1'b0 ;
  assign n24074 = ( n14497 & n20347 ) | ( n14497 & n24073 ) | ( n20347 & n24073 ) ;
  assign n24075 = n8163 ^ n5459 ^ 1'b0 ;
  assign n24076 = n15343 | n24075 ;
  assign n24077 = n4109 | n8314 ;
  assign n24078 = n15548 & ~n24077 ;
  assign n24079 = n9720 ^ n8685 ^ 1'b0 ;
  assign n24080 = n24079 ^ n2417 ^ 1'b0 ;
  assign n24081 = n5138 & n24080 ;
  assign n24082 = n2859 | n9787 ;
  assign n24083 = n6330 ^ n54 ^ 1'b0 ;
  assign n24084 = ~n10542 & n24083 ;
  assign n24085 = ~n8694 & n24084 ;
  assign n24086 = n24085 ^ n1477 ^ 1'b0 ;
  assign n24087 = n10910 ^ n3070 ^ 1'b0 ;
  assign n24088 = n6110 | n24087 ;
  assign n24089 = n24088 ^ n1068 ^ 1'b0 ;
  assign n24090 = n17592 ^ n3611 ^ 1'b0 ;
  assign n24091 = n24089 & ~n24090 ;
  assign n24093 = n7152 & ~n9332 ;
  assign n24092 = n330 | n13668 ;
  assign n24094 = n24093 ^ n24092 ^ n1298 ;
  assign n24095 = n15008 ^ n6321 ^ 1'b0 ;
  assign n24096 = n24094 & ~n24095 ;
  assign n24097 = n6748 ^ n4429 ^ 1'b0 ;
  assign n24098 = n9905 ^ n4970 ^ 1'b0 ;
  assign n24099 = ~n18187 & n24098 ;
  assign n24104 = n3019 & n9896 ;
  assign n24100 = n10568 | n11956 ;
  assign n24101 = x5 | n24100 ;
  assign n24102 = ( n5041 & n12860 ) | ( n5041 & n24101 ) | ( n12860 & n24101 ) ;
  assign n24103 = n1853 & ~n24102 ;
  assign n24105 = n24104 ^ n24103 ^ 1'b0 ;
  assign n24106 = n3970 & ~n6271 ;
  assign n24107 = ~n6201 & n6622 ;
  assign n24108 = ( n197 & n24106 ) | ( n197 & ~n24107 ) | ( n24106 & ~n24107 ) ;
  assign n24109 = n24108 ^ n2846 ^ 1'b0 ;
  assign n24110 = n16598 ^ n11759 ^ 1'b0 ;
  assign n24111 = n8296 & ~n24110 ;
  assign n24112 = n24111 ^ n1405 ^ 1'b0 ;
  assign n24113 = n24112 ^ n3325 ^ 1'b0 ;
  assign n24114 = n2222 & n24113 ;
  assign n24115 = n15562 ^ n7842 ^ n6799 ;
  assign n24116 = n4519 | n12081 ;
  assign n24117 = n1490 ^ n571 ^ 1'b0 ;
  assign n24118 = n16356 & ~n24117 ;
  assign n24119 = n4224 | n24118 ;
  assign n24120 = n13745 | n24119 ;
  assign n24121 = ~n5607 & n16791 ;
  assign n24122 = n24121 ^ n1313 ^ 1'b0 ;
  assign n24123 = n2781 ^ n1615 ^ 1'b0 ;
  assign n24124 = n171 & ~n23749 ;
  assign n24125 = n3235 & n9699 ;
  assign n24126 = n10115 ^ n9673 ^ n6593 ;
  assign n24127 = n2355 & n6613 ;
  assign n24128 = n1567 | n24127 ;
  assign n24129 = n20517 & ~n21500 ;
  assign n24130 = ~n1464 & n24129 ;
  assign n24137 = n7110 & ~n11020 ;
  assign n24133 = ~n6441 & n13063 ;
  assign n24134 = ~n7358 & n24133 ;
  assign n24131 = n3635 ^ n2267 ^ 1'b0 ;
  assign n24132 = n15117 & ~n24131 ;
  assign n24135 = n24134 ^ n24132 ^ 1'b0 ;
  assign n24136 = n15915 | n24135 ;
  assign n24138 = n24137 ^ n24136 ^ 1'b0 ;
  assign n24139 = n19879 & ~n24138 ;
  assign n24140 = n21461 ^ n14604 ^ n8201 ;
  assign n24141 = n22083 ^ n21315 ^ 1'b0 ;
  assign n24142 = n15435 ^ n7086 ^ 1'b0 ;
  assign n24143 = ~n12812 & n24142 ;
  assign n24144 = n8134 & n10175 ;
  assign n24145 = n19409 ^ n938 ^ 1'b0 ;
  assign n24146 = n21 & n4079 ;
  assign n24147 = n11296 ^ n8499 ^ 1'b0 ;
  assign n24148 = n6048 | n24147 ;
  assign n24149 = n24148 ^ n5707 ^ 1'b0 ;
  assign n24150 = n24149 ^ n17013 ^ 1'b0 ;
  assign n24151 = n11306 & ~n19822 ;
  assign n24152 = n3449 | n17843 ;
  assign n24153 = n12458 | n16458 ;
  assign n24154 = n6750 ^ n6429 ^ 1'b0 ;
  assign n24155 = n221 & ~n4691 ;
  assign n24156 = n10937 | n24155 ;
  assign n24157 = n24156 ^ n12632 ^ 1'b0 ;
  assign n24158 = n1601 & n12363 ;
  assign n24159 = n24157 & n24158 ;
  assign n24160 = n2146 ^ n1531 ^ 1'b0 ;
  assign n24161 = n1327 & n5615 ;
  assign n24162 = n24161 ^ n6805 ^ 1'b0 ;
  assign n24163 = n24162 ^ n19387 ^ 1'b0 ;
  assign n24164 = n5420 & ~n24163 ;
  assign n24165 = ~n24160 & n24164 ;
  assign n24166 = n24159 & n24165 ;
  assign n24167 = n22633 ^ n22249 ^ 1'b0 ;
  assign n24168 = ~n13618 & n16249 ;
  assign n24169 = n16591 | n19385 ;
  assign n24170 = ~n5546 & n24169 ;
  assign n24171 = n1413 | n7823 ;
  assign n24172 = n24171 ^ n10546 ^ 1'b0 ;
  assign n24173 = n5348 & ~n24172 ;
  assign n24174 = n9231 ^ n9170 ^ 1'b0 ;
  assign n24175 = n3867 ^ n619 ^ 1'b0 ;
  assign n24176 = n963 & n12879 ;
  assign n24177 = n1941 & n24176 ;
  assign n24178 = ~n2041 & n7238 ;
  assign n24179 = n3412 & n24178 ;
  assign n24180 = n18255 & n24179 ;
  assign n24181 = n15177 & n24180 ;
  assign n24182 = n24181 ^ n3351 ^ 1'b0 ;
  assign n24183 = ~n20350 & n24182 ;
  assign n24185 = n20029 | n21402 ;
  assign n24184 = n5458 | n15495 ;
  assign n24186 = n24185 ^ n24184 ^ 1'b0 ;
  assign n24187 = n4085 & n14200 ;
  assign n24188 = n24187 ^ n12070 ^ 1'b0 ;
  assign n24189 = n24188 ^ n17493 ^ n8166 ;
  assign n24190 = n3721 | n11366 ;
  assign n24191 = n11153 & ~n24190 ;
  assign n24192 = n21786 ^ n13340 ^ n3858 ;
  assign n24193 = ~n627 & n2754 ;
  assign n24194 = n5988 & n24193 ;
  assign n24195 = n3867 & ~n24194 ;
  assign n24196 = ~n14426 & n24195 ;
  assign n24197 = n12393 ^ n255 ^ 1'b0 ;
  assign n24198 = n12919 | n15470 ;
  assign n24199 = n24198 ^ n15089 ^ 1'b0 ;
  assign n24200 = n17673 & ~n24199 ;
  assign n24201 = n24200 ^ n9192 ^ 1'b0 ;
  assign n24202 = n24197 & ~n24201 ;
  assign n24203 = n9377 ^ n7798 ^ 1'b0 ;
  assign n24205 = n14602 ^ n7581 ^ 1'b0 ;
  assign n24206 = n6842 & ~n10263 ;
  assign n24207 = ~n24205 & n24206 ;
  assign n24208 = n8519 & ~n24207 ;
  assign n24204 = n9964 & n15231 ;
  assign n24209 = n24208 ^ n24204 ^ 1'b0 ;
  assign n24214 = ~n9912 & n11371 ;
  assign n24210 = n8743 | n9508 ;
  assign n24211 = n24210 ^ n4082 ^ 1'b0 ;
  assign n24212 = n8287 & ~n24211 ;
  assign n24213 = n24212 ^ n1853 ^ 1'b0 ;
  assign n24215 = n24214 ^ n24213 ^ n9963 ;
  assign n24216 = n24215 ^ n16173 ^ 1'b0 ;
  assign n24219 = n4416 & n7010 ;
  assign n24217 = n7219 ^ n6388 ^ 1'b0 ;
  assign n24218 = ~n4164 & n24217 ;
  assign n24220 = n24219 ^ n24218 ^ 1'b0 ;
  assign n24221 = n24220 ^ n23379 ^ n6638 ;
  assign n24222 = n7713 ^ n1413 ^ 1'b0 ;
  assign n24223 = n4532 & n9652 ;
  assign n24224 = n24223 ^ n5867 ^ 1'b0 ;
  assign n24225 = n24224 ^ n20065 ^ 1'b0 ;
  assign n24226 = ~n4147 & n24225 ;
  assign n24227 = n18486 & ~n21720 ;
  assign n24228 = n24227 ^ n8768 ^ 1'b0 ;
  assign n24229 = n24228 ^ n24131 ^ 1'b0 ;
  assign n24230 = n11345 & ~n24229 ;
  assign n24231 = n3413 & n13885 ;
  assign n24232 = n8962 | n19363 ;
  assign n24233 = n22779 | n24232 ;
  assign n24234 = n15045 ^ n8313 ^ n4967 ;
  assign n24235 = ~n11883 & n15230 ;
  assign n24236 = n24235 ^ n5821 ^ 1'b0 ;
  assign n24237 = n12550 ^ n2206 ^ 1'b0 ;
  assign n24238 = n7308 & n24237 ;
  assign n24239 = n19638 ^ n11002 ^ 1'b0 ;
  assign n24240 = n16297 & n24239 ;
  assign n24241 = n1267 | n14787 ;
  assign n24242 = n1267 & ~n24241 ;
  assign n24243 = n24242 ^ n15363 ^ 1'b0 ;
  assign n24244 = n18757 ^ n14954 ^ 1'b0 ;
  assign n24245 = n11050 & ~n24244 ;
  assign n24246 = ( n4328 & n24243 ) | ( n4328 & n24245 ) | ( n24243 & n24245 ) ;
  assign n24247 = n474 & ~n22638 ;
  assign n24248 = n3893 & ~n4066 ;
  assign n24249 = n20499 ^ n10858 ^ 1'b0 ;
  assign n24250 = ~n19632 & n24249 ;
  assign n24251 = n24250 ^ n5686 ^ 1'b0 ;
  assign n24252 = n24248 | n24251 ;
  assign n24253 = n4264 & ~n12884 ;
  assign n24254 = n5059 ^ n1205 ^ 1'b0 ;
  assign n24255 = n14968 & ~n24254 ;
  assign n24256 = n24255 ^ n8399 ^ 1'b0 ;
  assign n24257 = n24256 ^ n8375 ^ 1'b0 ;
  assign n24258 = ~n24253 & n24257 ;
  assign n24259 = n24258 ^ n20203 ^ n13228 ;
  assign n24260 = n1049 & n24259 ;
  assign n24261 = n7469 ^ n4318 ^ 1'b0 ;
  assign n24262 = n17999 ^ n11458 ^ 1'b0 ;
  assign n24263 = ( n401 & ~n1104 ) | ( n401 & n19494 ) | ( ~n1104 & n19494 ) ;
  assign n24264 = n7968 & n9746 ;
  assign n24265 = n24263 & ~n24264 ;
  assign n24266 = ~n2363 & n8758 ;
  assign n24267 = n11312 | n24266 ;
  assign n24268 = n24267 ^ n250 ^ 1'b0 ;
  assign n24269 = ( n5010 & ~n8551 ) | ( n5010 & n24073 ) | ( ~n8551 & n24073 ) ;
  assign n24270 = n6566 | n20987 ;
  assign n24271 = n24269 | n24270 ;
  assign n24272 = n18926 ^ n584 ^ 1'b0 ;
  assign n24273 = n24271 & ~n24272 ;
  assign n24274 = ~n1167 & n24273 ;
  assign n24275 = n24274 ^ n17318 ^ 1'b0 ;
  assign n24276 = n14001 ^ n8281 ^ 1'b0 ;
  assign n24277 = n15461 & ~n24276 ;
  assign n24278 = n6110 ^ n1877 ^ 1'b0 ;
  assign n24279 = n790 & ~n24278 ;
  assign n24280 = ~n899 & n3420 ;
  assign n24281 = ( n667 & n4659 ) | ( n667 & ~n23181 ) | ( n4659 & ~n23181 ) ;
  assign n24282 = n3761 | n24281 ;
  assign n24283 = n22660 ^ n18683 ^ 1'b0 ;
  assign n24284 = n24283 ^ n11489 ^ 1'b0 ;
  assign n24285 = n3772 ^ n3480 ^ 1'b0 ;
  assign n24286 = n15944 & n24285 ;
  assign n24287 = ~x11 & n8893 ;
  assign n24288 = n24287 ^ n9584 ^ n9348 ;
  assign n24289 = ~n19315 & n24288 ;
  assign n24290 = ~n9100 & n13481 ;
  assign n24291 = ( n7499 & ~n24288 ) | ( n7499 & n24290 ) | ( ~n24288 & n24290 ) ;
  assign n24292 = n17142 ^ n1742 ^ 1'b0 ;
  assign n24293 = ~n13597 & n24292 ;
  assign n24294 = n24293 ^ n15397 ^ 1'b0 ;
  assign n24295 = ( n16718 & ~n17271 ) | ( n16718 & n24294 ) | ( ~n17271 & n24294 ) ;
  assign n24296 = n6796 | n8292 ;
  assign n24297 = n24296 ^ n2685 ^ 1'b0 ;
  assign n24298 = n23772 ^ n2586 ^ 1'b0 ;
  assign n24299 = n1036 | n24298 ;
  assign n24300 = n3071 ^ n1819 ^ 1'b0 ;
  assign n24301 = n24300 ^ n19840 ^ n1020 ;
  assign n24302 = n5652 ^ n5477 ^ 1'b0 ;
  assign n24303 = ( n11240 & n13951 ) | ( n11240 & n20518 ) | ( n13951 & n20518 ) ;
  assign n24304 = n22341 ^ n9763 ^ 1'b0 ;
  assign n24305 = ~n11056 & n24304 ;
  assign n24306 = n24303 | n24305 ;
  assign n24307 = n24306 ^ n4734 ^ 1'b0 ;
  assign n24308 = n17134 & n18122 ;
  assign n24309 = n8693 & n8883 ;
  assign n24310 = n8660 ^ n1329 ^ 1'b0 ;
  assign n24311 = n5453 | n24310 ;
  assign n24312 = ( ~n1217 & n24309 ) | ( ~n1217 & n24311 ) | ( n24309 & n24311 ) ;
  assign n24313 = ~n16606 & n17079 ;
  assign n24314 = n4433 & ~n4965 ;
  assign n24315 = ~n19780 & n24314 ;
  assign n24316 = n22160 ^ n18879 ^ n11499 ;
  assign n24317 = n24316 ^ n3472 ^ 1'b0 ;
  assign n24318 = n18289 ^ n6758 ^ 1'b0 ;
  assign n24319 = n16788 ^ n790 ^ 1'b0 ;
  assign n24320 = n17662 & ~n24319 ;
  assign n24321 = ~n14030 & n24320 ;
  assign n24322 = n24318 & n24321 ;
  assign n24323 = ~n11723 & n19155 ;
  assign n24324 = ( n6520 & ~n16343 ) | ( n6520 & n24323 ) | ( ~n16343 & n24323 ) ;
  assign n24325 = ~n1582 & n1732 ;
  assign n24326 = n24325 ^ n2588 ^ 1'b0 ;
  assign n24327 = n13410 ^ n2730 ^ 1'b0 ;
  assign n24328 = n844 | n24327 ;
  assign n24329 = ( n3444 & ~n24326 ) | ( n3444 & n24328 ) | ( ~n24326 & n24328 ) ;
  assign n24330 = n9578 | n18236 ;
  assign n24331 = n1506 & n2518 ;
  assign n24332 = n24331 ^ n14988 ^ 1'b0 ;
  assign n24333 = n22293 ^ n1664 ^ 1'b0 ;
  assign n24334 = n3166 & ~n24333 ;
  assign n24335 = n738 & n3858 ;
  assign n24336 = n24334 | n24335 ;
  assign n24337 = ~n3665 & n7910 ;
  assign n24338 = n4372 & n24337 ;
  assign n24339 = n16292 & ~n24338 ;
  assign n24340 = ~n2484 & n15342 ;
  assign n24341 = ~n24339 & n24340 ;
  assign n24342 = n4835 & ~n5762 ;
  assign n24343 = n12236 ^ n6359 ^ 1'b0 ;
  assign n24344 = n23838 & ~n24343 ;
  assign n24345 = n24344 ^ n15244 ^ 1'b0 ;
  assign n24346 = n8267 ^ n5109 ^ 1'b0 ;
  assign n24347 = n24346 ^ n4618 ^ 1'b0 ;
  assign n24348 = ~n2769 & n24347 ;
  assign n24349 = n644 & ~n22801 ;
  assign n24350 = n11551 & n24349 ;
  assign n24359 = ~n228 & n1071 ;
  assign n24360 = ~n1071 & n24359 ;
  assign n24356 = n1510 & n3212 ;
  assign n24357 = ~n1510 & n24356 ;
  assign n24358 = n10881 | n24357 ;
  assign n24361 = n24360 ^ n24358 ^ 1'b0 ;
  assign n24351 = n9302 & n12015 ;
  assign n24352 = n1611 | n24351 ;
  assign n24353 = n24351 & ~n24352 ;
  assign n24354 = n24353 ^ n8406 ^ 1'b0 ;
  assign n24355 = n9023 & n24354 ;
  assign n24362 = n24361 ^ n24355 ^ n13523 ;
  assign n24363 = n16508 & n19645 ;
  assign n24364 = ~n4765 & n5259 ;
  assign n24365 = n24364 ^ n7405 ^ 1'b0 ;
  assign n24366 = n6979 & n24365 ;
  assign n24367 = n1014 & n24366 ;
  assign n24368 = ( n328 & ~n1988 ) | ( n328 & n11768 ) | ( ~n1988 & n11768 ) ;
  assign n24369 = n8229 & n24368 ;
  assign n24370 = n13481 & n24369 ;
  assign n24371 = n7918 | n13055 ;
  assign n24372 = n24370 & ~n24371 ;
  assign n24373 = n188 & ~n997 ;
  assign n24374 = ~n188 & n24373 ;
  assign n24375 = n1771 & ~n24374 ;
  assign n24376 = n20403 ^ n9441 ^ 1'b0 ;
  assign n24377 = n11885 & ~n24376 ;
  assign n24378 = n24375 | n24377 ;
  assign n24379 = n3470 & ~n16359 ;
  assign n24380 = n24379 ^ n3257 ^ 1'b0 ;
  assign n24381 = ~n21395 & n24380 ;
  assign n24382 = ~n1210 & n16369 ;
  assign n24383 = n10023 | n10189 ;
  assign n24384 = n17632 ^ n2523 ^ 1'b0 ;
  assign n24385 = n6838 | n9713 ;
  assign n24386 = n24271 ^ n6993 ^ 1'b0 ;
  assign n24387 = ~n8235 & n17477 ;
  assign n24388 = ~n1152 & n24387 ;
  assign n24389 = n16400 & n24388 ;
  assign n24391 = n4635 ^ n4084 ^ n316 ;
  assign n24392 = ( ~n835 & n15406 ) | ( ~n835 & n24391 ) | ( n15406 & n24391 ) ;
  assign n24390 = n4666 | n11381 ;
  assign n24393 = n24392 ^ n24390 ^ 1'b0 ;
  assign n24394 = ~n2929 & n5177 ;
  assign n24395 = ~n12168 & n24394 ;
  assign n24396 = n438 & n790 ;
  assign n24397 = n13769 & ~n21618 ;
  assign n24398 = n1742 & ~n10023 ;
  assign n24399 = n24398 ^ n4346 ^ 1'b0 ;
  assign n24400 = n20015 & ~n24399 ;
  assign n24401 = n8357 ^ n4263 ^ 1'b0 ;
  assign n24402 = n23670 ^ n7034 ^ 1'b0 ;
  assign n24403 = n24401 & ~n24402 ;
  assign n24404 = ~n3388 & n4780 ;
  assign n24405 = n24404 ^ n5363 ^ 1'b0 ;
  assign n24406 = n642 | n24405 ;
  assign n24407 = n17718 & n24406 ;
  assign n24408 = n24407 ^ n10562 ^ n86 ;
  assign n24409 = n5200 & ~n7589 ;
  assign n24410 = ~n6925 & n24409 ;
  assign n24411 = n17019 ^ n13329 ^ 1'b0 ;
  assign n24412 = n4528 & n24411 ;
  assign n24413 = n4835 ^ n1377 ^ n138 ;
  assign n24414 = n1521 & n24413 ;
  assign n24415 = ~n10218 & n24414 ;
  assign n24416 = n367 | n24415 ;
  assign n24417 = n24412 | n24416 ;
  assign n24419 = n7679 ^ n1038 ^ 1'b0 ;
  assign n24418 = n7747 | n14569 ;
  assign n24420 = n24419 ^ n24418 ^ 1'b0 ;
  assign n24421 = ~n21890 & n21956 ;
  assign n24422 = ( n4875 & n15897 ) | ( n4875 & ~n24421 ) | ( n15897 & ~n24421 ) ;
  assign n24423 = n4645 & n6516 ;
  assign n24424 = n24423 ^ n19913 ^ 1'b0 ;
  assign n24425 = n15651 & n24424 ;
  assign n24426 = n7978 ^ n3358 ^ 1'b0 ;
  assign n24427 = n208 & ~n582 ;
  assign n24428 = n24427 ^ n2708 ^ 1'b0 ;
  assign n24429 = n24428 ^ n1896 ^ 1'b0 ;
  assign n24430 = n11304 | n24429 ;
  assign n24431 = n2630 & n5824 ;
  assign n24432 = n24431 ^ n461 ^ 1'b0 ;
  assign n24433 = n10367 ^ n8145 ^ 1'b0 ;
  assign n24434 = n1025 & ~n2391 ;
  assign n24435 = n20294 ^ n8118 ^ 1'b0 ;
  assign n24436 = n24434 & n24435 ;
  assign n24438 = n5708 & n12875 ;
  assign n24437 = n5886 & ~n22420 ;
  assign n24439 = n24438 ^ n24437 ^ 1'b0 ;
  assign n24440 = n1109 & ~n24439 ;
  assign n24441 = n14861 & ~n23936 ;
  assign n24442 = n1823 & ~n10356 ;
  assign n24443 = n8798 & ~n24442 ;
  assign n24444 = n23 & ~n21187 ;
  assign n24445 = n19880 & ~n24444 ;
  assign n24446 = n24445 ^ n5564 ^ 1'b0 ;
  assign n24447 = n12496 & n13040 ;
  assign n24448 = n24447 ^ n74 ^ 1'b0 ;
  assign n24449 = n9593 ^ n2637 ^ 1'b0 ;
  assign n24450 = n14073 | n24449 ;
  assign n24451 = n15707 ^ n14989 ^ n14031 ;
  assign n24452 = n10278 ^ n8731 ^ 1'b0 ;
  assign n24455 = ( n3935 & n5235 ) | ( n3935 & ~n21591 ) | ( n5235 & ~n21591 ) ;
  assign n24453 = n15330 ^ n4621 ^ 1'b0 ;
  assign n24454 = ~n9967 & n24453 ;
  assign n24456 = n24455 ^ n24454 ^ 1'b0 ;
  assign n24457 = n1216 & n23314 ;
  assign n24458 = n24457 ^ n21331 ^ 1'b0 ;
  assign n24459 = n2816 ^ n1143 ^ 1'b0 ;
  assign n24462 = n17418 | n19343 ;
  assign n24463 = n14201 & ~n24462 ;
  assign n24460 = ~n6813 & n21870 ;
  assign n24461 = n21739 & n24460 ;
  assign n24464 = n24463 ^ n24461 ^ 1'b0 ;
  assign n24465 = ~n924 & n10740 ;
  assign n24466 = n24465 ^ n16786 ^ n6124 ;
  assign n24467 = n21717 ^ n6002 ^ 1'b0 ;
  assign n24468 = n8197 ^ n7456 ^ n6262 ;
  assign n24469 = n24467 & ~n24468 ;
  assign n24470 = n6869 | n18626 ;
  assign n24471 = ~n11176 & n12165 ;
  assign n24472 = n1090 & ~n6554 ;
  assign n24473 = ~n1045 & n24472 ;
  assign n24474 = n24473 ^ n16889 ^ n316 ;
  assign n24475 = n13114 ^ n115 ^ 1'b0 ;
  assign n24476 = x6 & ~n15512 ;
  assign n24477 = n24476 ^ n23749 ^ 1'b0 ;
  assign n24478 = n15766 ^ n7943 ^ n1204 ;
  assign n24479 = n3757 & ~n9748 ;
  assign n24480 = n24478 & n24479 ;
  assign n24481 = n24480 ^ n5895 ^ 1'b0 ;
  assign n24482 = n19680 & ~n24481 ;
  assign n24483 = ~n334 & n24482 ;
  assign n24484 = n61 | n16976 ;
  assign n24485 = n16410 | n24484 ;
  assign n24486 = ~n11251 & n15278 ;
  assign n24487 = n15273 ^ n14061 ^ n6100 ;
  assign n24488 = n368 | n5853 ;
  assign n24489 = n8352 | n24488 ;
  assign n24490 = n24489 ^ n5032 ^ 1'b0 ;
  assign n24491 = n11320 | n24490 ;
  assign n24492 = n24491 ^ n14206 ^ 1'b0 ;
  assign n24493 = ~n5768 & n24492 ;
  assign n24494 = n5813 ^ n1609 ^ 1'b0 ;
  assign n24495 = n3406 & ~n7767 ;
  assign n24496 = n9219 ^ n2619 ^ 1'b0 ;
  assign n24497 = ~n4024 & n24496 ;
  assign n24498 = ~n4931 & n8922 ;
  assign n24499 = n10595 ^ n9672 ^ 1'b0 ;
  assign n24500 = n20218 ^ n1576 ^ 1'b0 ;
  assign n24501 = ~n4519 & n24500 ;
  assign n24502 = ~n15322 & n24501 ;
  assign n24503 = n1010 & ~n2304 ;
  assign n24504 = n13794 & n24503 ;
  assign n24505 = n15519 ^ n1110 ^ 1'b0 ;
  assign n24506 = n1962 & ~n8099 ;
  assign n24507 = n327 & n24506 ;
  assign n24511 = ~n4993 & n19299 ;
  assign n24508 = n17162 ^ n2188 ^ 1'b0 ;
  assign n24509 = n952 | n24508 ;
  assign n24510 = n20819 & ~n24509 ;
  assign n24512 = n24511 ^ n24510 ^ n2735 ;
  assign n24513 = n24507 | n24512 ;
  assign n24517 = n9432 & n18808 ;
  assign n24514 = n2574 & ~n5051 ;
  assign n24515 = n6435 ^ n1187 ^ 1'b0 ;
  assign n24516 = n24514 & ~n24515 ;
  assign n24518 = n24517 ^ n24516 ^ 1'b0 ;
  assign n24519 = n9022 & ~n24518 ;
  assign n24520 = n24519 ^ n13990 ^ 1'b0 ;
  assign n24521 = n4113 & n6526 ;
  assign n24522 = n2552 & n15858 ;
  assign n24523 = ~n466 & n24522 ;
  assign n24524 = ~n21062 & n24523 ;
  assign n24525 = n666 | n18336 ;
  assign n24526 = n24525 ^ n10277 ^ 1'b0 ;
  assign n24528 = n9799 ^ n367 ^ 1'b0 ;
  assign n24529 = ~n15796 & n24528 ;
  assign n24530 = n19888 & n24529 ;
  assign n24531 = n24530 ^ n16050 ^ 1'b0 ;
  assign n24527 = ~n421 & n16343 ;
  assign n24532 = n24531 ^ n24527 ^ 1'b0 ;
  assign n24533 = n11314 ^ n6808 ^ 1'b0 ;
  assign n24534 = ~n7697 & n8031 ;
  assign n24535 = n5200 & ~n22864 ;
  assign n24536 = n4926 & n24535 ;
  assign n24537 = n774 | n24536 ;
  assign n24538 = n3303 & ~n24537 ;
  assign n24539 = n2118 & ~n23271 ;
  assign n24540 = n8482 ^ n4969 ^ 1'b0 ;
  assign n24541 = n3435 & ~n24540 ;
  assign n24542 = n16101 & n21083 ;
  assign n24543 = n390 | n1714 ;
  assign n24544 = n14138 & ~n24543 ;
  assign n24545 = n2317 & n21723 ;
  assign n24546 = n10901 ^ n6601 ^ 1'b0 ;
  assign n24547 = n4931 & n24546 ;
  assign n24548 = n4088 & n24547 ;
  assign n24549 = n12341 | n24548 ;
  assign n24550 = ~n2363 & n15442 ;
  assign n24551 = ~n9045 & n17350 ;
  assign n24552 = ~n4149 & n8924 ;
  assign n24553 = n24552 ^ n10342 ^ 1'b0 ;
  assign n24556 = n6079 & n7806 ;
  assign n24557 = n24556 ^ n17182 ^ 1'b0 ;
  assign n24558 = n24557 ^ n4430 ^ n3489 ;
  assign n24554 = n968 & ~n7326 ;
  assign n24555 = n311 & n24554 ;
  assign n24559 = n24558 ^ n24555 ^ 1'b0 ;
  assign n24560 = n106 | n671 ;
  assign n24561 = n6530 | n24560 ;
  assign n24565 = n2785 & ~n6003 ;
  assign n24562 = ~n8009 & n11779 ;
  assign n24563 = n24562 ^ n7346 ^ 1'b0 ;
  assign n24564 = ~n12995 & n24563 ;
  assign n24566 = n24565 ^ n24564 ^ 1'b0 ;
  assign n24567 = n24566 ^ n2885 ^ 1'b0 ;
  assign n24568 = ~n11472 & n24567 ;
  assign n24569 = n21596 ^ n11918 ^ 1'b0 ;
  assign n24570 = n24568 & n24569 ;
  assign n24571 = n5870 & n18252 ;
  assign n24572 = n1636 & n13069 ;
  assign n24573 = n12825 & n24572 ;
  assign n24574 = ( n9432 & n11946 ) | ( n9432 & ~n24573 ) | ( n11946 & ~n24573 ) ;
  assign n24575 = n10728 ^ n349 ^ 1'b0 ;
  assign n24576 = ~n2893 & n24575 ;
  assign n24577 = ~n1586 & n24576 ;
  assign n24578 = n24577 ^ n13028 ^ 1'b0 ;
  assign n24579 = n9170 ^ n5420 ^ 1'b0 ;
  assign n24580 = n24578 | n24579 ;
  assign n24581 = n10144 | n16493 ;
  assign n24582 = n4135 | n24581 ;
  assign n24583 = n7958 & ~n24582 ;
  assign n24584 = n9010 & ~n24583 ;
  assign n24585 = ~n12050 & n24584 ;
  assign n24586 = n24580 | n24585 ;
  assign n24587 = n24586 ^ n4207 ^ 1'b0 ;
  assign n24588 = n24574 & n24587 ;
  assign n24589 = n2362 & ~n4960 ;
  assign n24590 = ( n85 & ~n695 ) | ( n85 & n24589 ) | ( ~n695 & n24589 ) ;
  assign n24591 = n23253 ^ n19752 ^ 1'b0 ;
  assign n24592 = n7054 & ~n24591 ;
  assign n24593 = n18801 & n22920 ;
  assign n24594 = n14423 & n16701 ;
  assign n24595 = n8334 | n17465 ;
  assign n24596 = n873 & ~n24595 ;
  assign n24597 = ~n24594 & n24596 ;
  assign n24598 = n11972 & n21559 ;
  assign n24599 = ~n10318 & n24598 ;
  assign n24600 = n24149 ^ n12922 ^ 1'b0 ;
  assign n24601 = ~n16544 & n22039 ;
  assign n24604 = n138 & n1542 ;
  assign n24605 = ~n1542 & n24604 ;
  assign n24606 = n2382 | n24605 ;
  assign n24607 = n2382 & ~n24606 ;
  assign n24608 = n3446 | n24607 ;
  assign n24609 = n24607 & ~n24608 ;
  assign n24602 = n2275 ^ n2267 ^ n74 ;
  assign n24603 = n12128 | n24602 ;
  assign n24610 = n24609 ^ n24603 ^ n20075 ;
  assign n24611 = n312 & n4309 ;
  assign n24612 = ~n9038 & n24611 ;
  assign n24613 = n11875 ^ n10706 ^ 1'b0 ;
  assign n24614 = ~n19372 & n24613 ;
  assign n24615 = ~n2349 & n18134 ;
  assign n24616 = n24615 ^ n21048 ^ 1'b0 ;
  assign n24617 = n14081 & n24616 ;
  assign n24618 = ( n1976 & n2755 ) | ( n1976 & ~n16283 ) | ( n2755 & ~n16283 ) ;
  assign n24619 = n21124 & ~n24618 ;
  assign n24620 = n4189 & ~n23892 ;
  assign n24621 = ( n120 & n944 ) | ( n120 & ~n3622 ) | ( n944 & ~n3622 ) ;
  assign n24622 = n24620 & ~n24621 ;
  assign n24623 = n2891 | n5660 ;
  assign n24624 = n4859 | n24623 ;
  assign n24625 = n7814 & n24624 ;
  assign n24626 = ~n4394 & n6057 ;
  assign n24627 = n6570 & ~n24626 ;
  assign n24628 = n24625 & n24627 ;
  assign n24629 = ~n2798 & n12692 ;
  assign n24630 = n24629 ^ n4888 ^ 1'b0 ;
  assign n24631 = n13397 ^ n2645 ^ 1'b0 ;
  assign n24632 = ~n4351 & n24631 ;
  assign n24633 = n12700 & ~n24632 ;
  assign n24634 = n12380 | n12559 ;
  assign n24635 = n24634 ^ n5538 ^ 1'b0 ;
  assign n24637 = n7142 & n15531 ;
  assign n24636 = n12338 & n18421 ;
  assign n24638 = n24637 ^ n24636 ^ 1'b0 ;
  assign n24639 = n5823 & ~n18418 ;
  assign n24640 = n24639 ^ n9927 ^ 1'b0 ;
  assign n24641 = n942 | n23981 ;
  assign n24642 = n24641 ^ n2649 ^ 1'b0 ;
  assign n24643 = n24642 ^ n20383 ^ 1'b0 ;
  assign n24644 = n279 & ~n9493 ;
  assign n24645 = n24644 ^ n345 ^ 1'b0 ;
  assign n24646 = n24645 ^ n7965 ^ 1'b0 ;
  assign n24647 = n4357 & ~n23510 ;
  assign n24648 = ( n9031 & n18869 ) | ( n9031 & ~n21313 ) | ( n18869 & ~n21313 ) ;
  assign n24649 = n2976 & ~n15495 ;
  assign n24650 = n24649 ^ n8993 ^ 1'b0 ;
  assign n24651 = ~n2403 & n24650 ;
  assign n24652 = ~n1062 & n9721 ;
  assign n24653 = n23373 & n24652 ;
  assign n24654 = n16379 ^ n14194 ^ 1'b0 ;
  assign n24655 = n7146 & n24654 ;
  assign n24656 = n6074 & n14088 ;
  assign n24657 = n1286 | n15897 ;
  assign n24658 = ~n9325 & n21297 ;
  assign n24659 = n17439 ^ n162 ^ 1'b0 ;
  assign n24660 = ( n1315 & n15360 ) | ( n1315 & ~n24659 ) | ( n15360 & ~n24659 ) ;
  assign n24662 = n5042 ^ n4472 ^ 1'b0 ;
  assign n24663 = n5405 & n24662 ;
  assign n24664 = n179 | n4083 ;
  assign n24665 = n24663 & ~n24664 ;
  assign n24666 = n24665 ^ n7033 ^ 1'b0 ;
  assign n24667 = n24666 ^ n7369 ^ 1'b0 ;
  assign n24661 = n8334 | n10531 ;
  assign n24668 = n24667 ^ n24661 ^ 1'b0 ;
  assign n24669 = ~n129 & n10598 ;
  assign n24670 = n24669 ^ n8904 ^ 1'b0 ;
  assign n24671 = n24668 | n24670 ;
  assign n24672 = n14963 & ~n22022 ;
  assign n24673 = ~n3842 & n19912 ;
  assign n24674 = n11170 & ~n24673 ;
  assign n24675 = ~n8716 & n24674 ;
  assign n24676 = n10086 ^ n8362 ^ 1'b0 ;
  assign n24677 = ~n19931 & n24676 ;
  assign n24678 = ( n3428 & ~n14922 ) | ( n3428 & n22598 ) | ( ~n14922 & n22598 ) ;
  assign n24679 = n6157 & n24678 ;
  assign n24680 = ~n17901 & n24679 ;
  assign n24681 = n24680 ^ n13083 ^ 1'b0 ;
  assign n24682 = n10089 ^ n4401 ^ 1'b0 ;
  assign n24683 = n9249 | n10975 ;
  assign n24684 = n11613 | n24683 ;
  assign n24685 = n14489 | n24684 ;
  assign n24686 = n298 & n4357 ;
  assign n24687 = n24686 ^ n14525 ^ 1'b0 ;
  assign n24688 = n1943 & ~n2002 ;
  assign n24689 = ~n19535 & n24688 ;
  assign n24690 = ~n24687 & n24689 ;
  assign n24696 = n1138 & n22024 ;
  assign n24697 = n1517 | n24696 ;
  assign n24691 = n2754 & ~n8730 ;
  assign n24692 = n24691 ^ n3907 ^ 1'b0 ;
  assign n24693 = ~n5803 & n24692 ;
  assign n24694 = n24693 ^ n12035 ^ 1'b0 ;
  assign n24695 = n1304 & ~n24694 ;
  assign n24698 = n24697 ^ n24695 ^ 1'b0 ;
  assign n24699 = n19173 ^ n18485 ^ 1'b0 ;
  assign n24700 = n2940 | n12142 ;
  assign n24701 = n6027 ^ n4902 ^ 1'b0 ;
  assign n24702 = n24701 ^ n7257 ^ 1'b0 ;
  assign n24703 = n4039 | n24702 ;
  assign n24704 = n12299 ^ n4356 ^ 1'b0 ;
  assign n24705 = n24703 | n24704 ;
  assign n24706 = ( n19524 & ~n24700 ) | ( n19524 & n24705 ) | ( ~n24700 & n24705 ) ;
  assign n24707 = n21883 ^ n2532 ^ 1'b0 ;
  assign n24708 = n7451 & ~n24707 ;
  assign n24709 = ~n6085 & n8391 ;
  assign n24710 = n24709 ^ n9070 ^ 1'b0 ;
  assign n24711 = n24708 & n24710 ;
  assign n24712 = n11622 & n18708 ;
  assign n24713 = n15488 ^ n1548 ^ 1'b0 ;
  assign n24714 = n14606 ^ n881 ^ 1'b0 ;
  assign n24715 = n56 | n5416 ;
  assign n24716 = n24715 ^ n7856 ^ 1'b0 ;
  assign n24717 = n11440 ^ n2343 ^ 1'b0 ;
  assign n24718 = n11458 & n24717 ;
  assign n24719 = n24718 ^ n10112 ^ 1'b0 ;
  assign n24720 = n4365 | n10656 ;
  assign n24721 = n24719 | n24720 ;
  assign n24722 = n1553 & ~n24721 ;
  assign n24723 = n3927 ^ n2471 ^ 1'b0 ;
  assign n24729 = n6397 ^ n3343 ^ 1'b0 ;
  assign n24730 = n8239 & ~n24729 ;
  assign n24728 = n2794 & ~n5001 ;
  assign n24724 = n11435 ^ n6366 ^ 1'b0 ;
  assign n24725 = ~n4819 & n24724 ;
  assign n24726 = n24725 ^ n16052 ^ 1'b0 ;
  assign n24727 = n24726 ^ n6694 ^ 1'b0 ;
  assign n24731 = n24730 ^ n24728 ^ n24727 ;
  assign n24732 = n9335 ^ n5492 ^ 1'b0 ;
  assign n24733 = n24732 ^ n12559 ^ 1'b0 ;
  assign n24734 = n8717 & n24733 ;
  assign n24735 = n24734 ^ n3630 ^ n1392 ;
  assign n24736 = n24735 ^ n1570 ^ 1'b0 ;
  assign n24737 = n7918 ^ n3225 ^ 1'b0 ;
  assign n24738 = n19586 ^ n10805 ^ 1'b0 ;
  assign n24739 = ~n24737 & n24738 ;
  assign n24740 = n16920 ^ n15084 ^ 1'b0 ;
  assign n24741 = n23561 & n24740 ;
  assign n24742 = n20001 ^ n4290 ^ 1'b0 ;
  assign n24743 = n9354 | n14971 ;
  assign n24744 = n11861 ^ n466 ^ 1'b0 ;
  assign n24745 = n24744 ^ n13687 ^ 1'b0 ;
  assign n24746 = n13852 ^ n10086 ^ 1'b0 ;
  assign n24747 = n13011 & ~n24746 ;
  assign n24748 = n889 ^ n333 ^ 1'b0 ;
  assign n24749 = n13741 & n24748 ;
  assign n24750 = ~n9177 & n24749 ;
  assign n24751 = ~n1495 & n24750 ;
  assign n24752 = n1546 & n10634 ;
  assign n24753 = n2591 & n24752 ;
  assign n24754 = n24753 ^ n23630 ^ 1'b0 ;
  assign n24755 = ~n7873 & n24754 ;
  assign n24756 = n12777 ^ n6099 ^ n4946 ;
  assign n24757 = n3539 & ~n18359 ;
  assign n24758 = ~n8807 & n24757 ;
  assign n24759 = n24758 ^ n18046 ^ 1'b0 ;
  assign n24760 = ~n2562 & n22436 ;
  assign n24761 = n21187 & n22937 ;
  assign n24762 = ~n8490 & n24761 ;
  assign n24763 = n15906 ^ n3802 ^ 1'b0 ;
  assign n24764 = n24763 ^ n10855 ^ 1'b0 ;
  assign n24765 = n1467 ^ n56 ^ 1'b0 ;
  assign n24766 = n119 | n24765 ;
  assign n24770 = n12638 ^ n9707 ^ 1'b0 ;
  assign n24771 = n8302 & ~n24770 ;
  assign n24767 = n3186 ^ n503 ^ 1'b0 ;
  assign n24768 = n17335 & n24767 ;
  assign n24769 = n24768 ^ n7705 ^ 1'b0 ;
  assign n24772 = n24771 ^ n24769 ^ 1'b0 ;
  assign n24773 = ~n3968 & n24772 ;
  assign n24774 = n19298 ^ n9923 ^ 1'b0 ;
  assign n24775 = n4213 & n24774 ;
  assign n24776 = n24775 ^ n16382 ^ 1'b0 ;
  assign n24777 = n24776 ^ n565 ^ 1'b0 ;
  assign n24778 = n3545 & n24777 ;
  assign n24779 = n16106 ^ n1211 ^ 1'b0 ;
  assign n24780 = n1426 | n6640 ;
  assign n24781 = n24780 ^ n4639 ^ 1'b0 ;
  assign n24782 = n24781 ^ n18263 ^ 1'b0 ;
  assign n24783 = n4677 | n12088 ;
  assign n24784 = n24783 ^ n24380 ^ n12088 ;
  assign n24785 = ~n10738 & n17000 ;
  assign n24786 = ~n18864 & n24785 ;
  assign n24787 = n24786 ^ n11572 ^ 1'b0 ;
  assign n24789 = ~n5812 & n14802 ;
  assign n24790 = n3513 & n24789 ;
  assign n24788 = n3886 | n13324 ;
  assign n24791 = n24790 ^ n24788 ^ 1'b0 ;
  assign n24792 = n4853 ^ n216 ^ 1'b0 ;
  assign n24793 = n14775 & n24792 ;
  assign n24794 = n24791 & n24793 ;
  assign n24795 = n3320 & n5725 ;
  assign n24796 = n1179 & ~n6623 ;
  assign n24797 = n24796 ^ n4460 ^ 1'b0 ;
  assign n24798 = n24797 ^ n6844 ^ 1'b0 ;
  assign n24799 = n10403 ^ n3226 ^ 1'b0 ;
  assign n24800 = n6785 ^ n1109 ^ 1'b0 ;
  assign n24801 = n24800 ^ n21604 ^ 1'b0 ;
  assign n24802 = n24799 | n24801 ;
  assign n24803 = n6110 ^ n2826 ^ 1'b0 ;
  assign n24804 = n588 | n24803 ;
  assign n24805 = n3035 | n24804 ;
  assign n24806 = ~n65 & n5345 ;
  assign n24807 = n16872 & n24806 ;
  assign n24808 = n19237 ^ n18496 ^ 1'b0 ;
  assign n24809 = ( n1920 & ~n5664 ) | ( n1920 & n9905 ) | ( ~n5664 & n9905 ) ;
  assign n24810 = ~n2860 & n24809 ;
  assign n24811 = n5052 | n24810 ;
  assign n24812 = n5002 ^ n2211 ^ 1'b0 ;
  assign n24813 = n18099 & ~n24117 ;
  assign n24814 = n3471 ^ n3139 ^ 1'b0 ;
  assign n24815 = n24814 ^ n9337 ^ 1'b0 ;
  assign n24816 = n12343 ^ n136 ^ 1'b0 ;
  assign n24819 = n8330 ^ n4698 ^ n1891 ;
  assign n24817 = ~n1208 & n17762 ;
  assign n24818 = n24817 ^ n7401 ^ 1'b0 ;
  assign n24820 = n24819 ^ n24818 ^ 1'b0 ;
  assign n24821 = ~n9736 & n20249 ;
  assign n24822 = ~n6625 & n7136 ;
  assign n24823 = ~n5642 & n24822 ;
  assign n24824 = n1767 & n7589 ;
  assign n24825 = ~n20249 & n24824 ;
  assign n24826 = n24068 ^ n19186 ^ n15850 ;
  assign n24827 = n4547 ^ n23 ^ 1'b0 ;
  assign n24828 = n4838 & n24199 ;
  assign n24829 = ~n24827 & n24828 ;
  assign n24830 = n3052 | n3351 ;
  assign n24831 = n1277 & ~n5142 ;
  assign n24832 = n24831 ^ n1714 ^ 1'b0 ;
  assign n24833 = n19757 | n24832 ;
  assign n24834 = n24830 | n24833 ;
  assign n24835 = n15938 ^ n5215 ^ 1'b0 ;
  assign n24836 = n4809 & n11100 ;
  assign n24837 = n2571 | n7531 ;
  assign n24838 = n24837 ^ n12843 ^ 1'b0 ;
  assign n24839 = n24838 ^ n16485 ^ 1'b0 ;
  assign n24840 = n15872 & ~n24839 ;
  assign n24841 = ~n9203 & n24840 ;
  assign n24842 = n15393 & ~n16781 ;
  assign n24843 = n24841 & n24842 ;
  assign n24844 = ( ~n8903 & n9961 ) | ( ~n8903 & n24843 ) | ( n9961 & n24843 ) ;
  assign n24845 = n2612 | n22469 ;
  assign n24846 = n24845 ^ n7234 ^ 1'b0 ;
  assign n24847 = n696 & ~n13085 ;
  assign n24848 = n10716 & n24847 ;
  assign n24849 = n24848 ^ n2146 ^ 1'b0 ;
  assign n24850 = n19458 & ~n24849 ;
  assign n24851 = n9925 ^ n4525 ^ 1'b0 ;
  assign n24852 = n20543 ^ n4891 ^ 1'b0 ;
  assign n24853 = n9839 & n24852 ;
  assign n24854 = n6908 & n8078 ;
  assign n24855 = ~n5695 & n24854 ;
  assign n24856 = n24855 ^ n14934 ^ 1'b0 ;
  assign n24857 = n12322 ^ n11333 ^ 1'b0 ;
  assign n24858 = n9673 & ~n19129 ;
  assign n24860 = n2521 ^ n2322 ^ 1'b0 ;
  assign n24861 = n7554 & n24860 ;
  assign n24862 = n24861 ^ n16367 ^ n1187 ;
  assign n24859 = n14493 & n21121 ;
  assign n24863 = n24862 ^ n24859 ^ 1'b0 ;
  assign n24864 = n8111 | n13839 ;
  assign n24865 = n24864 ^ n16935 ^ 1'b0 ;
  assign n24866 = n6035 & ~n24865 ;
  assign n24867 = n18062 & n24866 ;
  assign n24868 = ~n12030 & n14710 ;
  assign n24869 = ~n12692 & n24868 ;
  assign n24870 = ( n5355 & n11873 ) | ( n5355 & ~n16221 ) | ( n11873 & ~n16221 ) ;
  assign n24871 = n867 | n24870 ;
  assign n24872 = n24869 & ~n24871 ;
  assign n24873 = n4741 & n8519 ;
  assign n24874 = ~n16069 & n24873 ;
  assign n24875 = n13726 ^ n5878 ^ 1'b0 ;
  assign n24876 = n8998 & n24875 ;
  assign n24877 = n481 | n5526 ;
  assign n24878 = n6982 & ~n24877 ;
  assign n24879 = n209 & ~n8677 ;
  assign n24880 = ~n716 & n24879 ;
  assign n24881 = n6945 & ~n24880 ;
  assign n24882 = n12451 ^ n10708 ^ n6314 ;
  assign n24883 = ( n4267 & ~n5150 ) | ( n4267 & n9201 ) | ( ~n5150 & n9201 ) ;
  assign n24884 = n5190 | n5425 ;
  assign n24885 = n19367 | n24884 ;
  assign n24886 = n2151 & n4493 ;
  assign n24887 = ~n22638 & n24886 ;
  assign n24888 = n12430 ^ n1808 ^ 1'b0 ;
  assign n24890 = n21452 & ~n21743 ;
  assign n24889 = n3408 ^ n2549 ^ 1'b0 ;
  assign n24891 = n24890 ^ n24889 ^ n21344 ;
  assign n24892 = n24708 ^ n23790 ^ 1'b0 ;
  assign n24893 = n6616 ^ n5548 ^ 1'b0 ;
  assign n24895 = n8304 ^ n5872 ^ n582 ;
  assign n24896 = n24895 ^ n1652 ^ 1'b0 ;
  assign n24897 = ~n1469 & n24896 ;
  assign n24894 = n11740 & n24514 ;
  assign n24898 = n24897 ^ n24894 ^ 1'b0 ;
  assign n24899 = n1469 | n4922 ;
  assign n24900 = n1469 & ~n24899 ;
  assign n24901 = n24900 ^ n6302 ^ 1'b0 ;
  assign n24902 = n24901 ^ n14360 ^ 1'b0 ;
  assign n24903 = n24898 | n24902 ;
  assign n24904 = n15602 ^ n8233 ^ n225 ;
  assign n24905 = n6645 | n24904 ;
  assign n24906 = n17482 ^ n2940 ^ n2682 ;
  assign n24907 = n24906 ^ n6203 ^ 1'b0 ;
  assign n24908 = ~n4218 & n24907 ;
  assign n24909 = n17900 ^ n15970 ^ 1'b0 ;
  assign n24910 = n7194 | n20340 ;
  assign n24911 = n3279 | n16367 ;
  assign n24912 = n9499 | n20670 ;
  assign n24913 = n16343 | n24912 ;
  assign n24914 = n918 & n24913 ;
  assign n24915 = n24911 & n24914 ;
  assign n24916 = n2103 | n18399 ;
  assign n24917 = n4440 | n24916 ;
  assign n24923 = n2905 & ~n19298 ;
  assign n24924 = n24923 ^ n23344 ^ 1'b0 ;
  assign n24925 = n9373 & ~n24924 ;
  assign n24926 = n24925 ^ n14429 ^ 1'b0 ;
  assign n24918 = n5950 & ~n9051 ;
  assign n24919 = n24918 ^ n5014 ^ 1'b0 ;
  assign n24920 = n8896 | n24919 ;
  assign n24921 = n24920 ^ n4074 ^ 1'b0 ;
  assign n24922 = n5758 & n24921 ;
  assign n24927 = n24926 ^ n24922 ^ 1'b0 ;
  assign n24928 = n16417 & n21849 ;
  assign n24929 = n24895 ^ n24182 ^ n15528 ;
  assign n24930 = ~n2330 & n22553 ;
  assign n24931 = ~n425 & n1347 ;
  assign n24932 = n11300 | n24839 ;
  assign n24933 = n24932 ^ n14757 ^ 1'b0 ;
  assign n24934 = n18803 & n23996 ;
  assign n24935 = n2481 & n24934 ;
  assign n24936 = n4657 & n10955 ;
  assign n24937 = ~n9796 & n24936 ;
  assign n24940 = n1080 & ~n16400 ;
  assign n24938 = n7167 ^ n6110 ^ 1'b0 ;
  assign n24939 = n24938 ^ n14038 ^ n7524 ;
  assign n24941 = n24940 ^ n24939 ^ 1'b0 ;
  assign n24942 = n24941 ^ n6719 ^ 1'b0 ;
  assign n24943 = n24937 | n24942 ;
  assign n24944 = ( n6979 & ~n13599 ) | ( n6979 & n24943 ) | ( ~n13599 & n24943 ) ;
  assign n24945 = n16891 ^ n5775 ^ 1'b0 ;
  assign n24946 = n18321 ^ n12456 ^ 1'b0 ;
  assign n24947 = n9676 & ~n24946 ;
  assign n24948 = n24947 ^ n18217 ^ 1'b0 ;
  assign n24949 = n16079 & n24948 ;
  assign n24950 = n17436 & n24949 ;
  assign n24951 = ~n18385 & n21855 ;
  assign n24952 = ~n5999 & n24951 ;
  assign n24953 = n832 & ~n18547 ;
  assign n24954 = n124 | n18514 ;
  assign n24955 = n3626 ^ n2869 ^ n755 ;
  assign n24956 = n3674 ^ n146 ^ 1'b0 ;
  assign n24957 = ( n23025 & n24955 ) | ( n23025 & ~n24956 ) | ( n24955 & ~n24956 ) ;
  assign n24958 = n3335 & ~n4361 ;
  assign n24959 = n5682 & ~n24078 ;
  assign n24961 = n253 & n6991 ;
  assign n24962 = n24961 ^ n11524 ^ 1'b0 ;
  assign n24960 = n9513 | n19305 ;
  assign n24963 = n24962 ^ n24960 ^ 1'b0 ;
  assign n24964 = n7114 | n8029 ;
  assign n24965 = n12376 ^ n459 ^ 1'b0 ;
  assign n24966 = ( n5366 & ~n7059 ) | ( n5366 & n23317 ) | ( ~n7059 & n23317 ) ;
  assign n24967 = ~n3080 & n24966 ;
  assign n24968 = x1 | n9087 ;
  assign n24969 = n24968 ^ n16942 ^ 1'b0 ;
  assign n24970 = n10491 | n24969 ;
  assign n24971 = n15142 | n24970 ;
  assign n24972 = n11880 ^ n7182 ^ n5714 ;
  assign n24973 = ~n3318 & n16975 ;
  assign n24975 = n11717 ^ n8834 ^ 1'b0 ;
  assign n24974 = n5028 | n15541 ;
  assign n24976 = n24975 ^ n24974 ^ 1'b0 ;
  assign n24977 = ( n261 & ~n10711 ) | ( n261 & n21579 ) | ( ~n10711 & n21579 ) ;
  assign n24978 = ~n22968 & n23240 ;
  assign n24979 = n17262 ^ n6360 ^ 1'b0 ;
  assign n24980 = n9832 & n24979 ;
  assign n24981 = n12974 & n24980 ;
  assign n24982 = n24981 ^ n8600 ^ 1'b0 ;
  assign n24983 = n3562 | n21581 ;
  assign n24984 = n641 | n7245 ;
  assign n24985 = n7153 & ~n24984 ;
  assign n24986 = n10752 | n24985 ;
  assign n24987 = n13874 ^ n806 ^ 1'b0 ;
  assign n24988 = n6024 & n24987 ;
  assign n24990 = n1635 & n15491 ;
  assign n24991 = n24990 ^ n13490 ^ 1'b0 ;
  assign n24989 = ( n6660 & n8550 ) | ( n6660 & ~n16460 ) | ( n8550 & ~n16460 ) ;
  assign n24992 = n24991 ^ n24989 ^ 1'b0 ;
  assign n24993 = n2335 & ~n8879 ;
  assign n24994 = n18831 & n24993 ;
  assign n24995 = n4704 & n7998 ;
  assign n24996 = n18962 & n24995 ;
  assign n24997 = ~n6883 & n10475 ;
  assign n24998 = n2730 & n9780 ;
  assign n24999 = ~n23369 & n24998 ;
  assign n25000 = ~n1159 & n7073 ;
  assign n25001 = n25000 ^ n17115 ^ 1'b0 ;
  assign n25002 = n8756 & n14371 ;
  assign n25003 = n25002 ^ n2242 ^ 1'b0 ;
  assign n25004 = n25003 ^ n20362 ^ n13505 ;
  assign n25005 = n22344 ^ n14284 ^ n13673 ;
  assign n25006 = n14297 & n25005 ;
  assign n25007 = x6 | n25006 ;
  assign n25008 = n1024 | n4685 ;
  assign n25009 = ~n13787 & n25008 ;
  assign n25010 = n25009 ^ n2829 ^ 1'b0 ;
  assign n25011 = n25010 ^ n6846 ^ 1'b0 ;
  assign n25012 = ~n20730 & n25011 ;
  assign n25013 = n4951 & ~n24895 ;
  assign n25014 = n25013 ^ n2327 ^ 1'b0 ;
  assign n25015 = n25014 ^ n6488 ^ 1'b0 ;
  assign n25016 = n2890 | n25015 ;
  assign n25017 = n20537 & n24669 ;
  assign n25018 = n23281 ^ n116 ^ 1'b0 ;
  assign n25019 = n2370 & ~n11407 ;
  assign n25020 = n5418 ^ n5344 ^ 1'b0 ;
  assign n25021 = n25020 ^ n3715 ^ 1'b0 ;
  assign n25022 = n23966 | n25021 ;
  assign n25023 = n25022 ^ n2401 ^ 1'b0 ;
  assign n25024 = n8244 ^ n6101 ^ n3777 ;
  assign n25025 = n15813 & ~n19173 ;
  assign n25026 = n22373 & n25025 ;
  assign n25027 = n25024 & n25026 ;
  assign n25028 = ~n17855 & n21187 ;
  assign n25029 = n7382 ^ n1684 ^ 1'b0 ;
  assign n25030 = n15493 ^ n5888 ^ 1'b0 ;
  assign n25031 = n83 | n25030 ;
  assign n25032 = n11498 & ~n19336 ;
  assign n25033 = ~n9032 & n18797 ;
  assign n25034 = ~n1280 & n3251 ;
  assign n25035 = n14034 | n25034 ;
  assign n25036 = n25035 ^ n1186 ^ 1'b0 ;
  assign n25037 = n18295 ^ n16343 ^ n6381 ;
  assign n25038 = n25037 ^ n15449 ^ 1'b0 ;
  assign n25039 = n23721 | n25038 ;
  assign n25040 = ( n1679 & n9417 ) | ( n1679 & n22007 ) | ( n9417 & n22007 ) ;
  assign n25041 = n25040 ^ n8536 ^ 1'b0 ;
  assign n25042 = n3849 & ~n15298 ;
  assign n25043 = n24015 ^ n10596 ^ 1'b0 ;
  assign n25044 = n21251 & ~n25043 ;
  assign n25045 = n25044 ^ n14276 ^ 1'b0 ;
  assign n25046 = ~n77 & n25045 ;
  assign n25047 = ( n4546 & n23190 ) | ( n4546 & ~n23619 ) | ( n23190 & ~n23619 ) ;
  assign n25048 = n16167 & ~n17369 ;
  assign n25049 = n5883 & n21457 ;
  assign n25050 = ~n2841 & n25049 ;
  assign n25051 = n482 & n14734 ;
  assign n25052 = n10624 & n25051 ;
  assign n25053 = n257 & ~n10220 ;
  assign n25054 = n25053 ^ n23362 ^ 1'b0 ;
  assign n25055 = x6 & n25054 ;
  assign n25056 = n18640 ^ n2284 ^ 1'b0 ;
  assign n25057 = n5909 & n25056 ;
  assign n25058 = n22283 & n25057 ;
  assign n25059 = ~n3958 & n19519 ;
  assign n25060 = ~n4094 & n25059 ;
  assign n25061 = n14081 ^ n5684 ^ n5352 ;
  assign n25062 = n19478 ^ n1438 ^ 1'b0 ;
  assign n25063 = n1853 & n8618 ;
  assign n25064 = n25063 ^ n9321 ^ 1'b0 ;
  assign n25065 = n24115 ^ n20201 ^ 1'b0 ;
  assign n25066 = n2967 | n3219 ;
  assign n25067 = n25066 ^ n7653 ^ 1'b0 ;
  assign n25068 = n14992 & n25067 ;
  assign n25069 = n2885 & n21707 ;
  assign n25070 = n9733 ^ n139 ^ 1'b0 ;
  assign n25071 = n25070 ^ n10653 ^ 1'b0 ;
  assign n25072 = n22150 & ~n25071 ;
  assign n25073 = n12996 ^ n3592 ^ 1'b0 ;
  assign n25074 = n2411 & ~n3017 ;
  assign n25075 = n25074 ^ n10473 ^ 1'b0 ;
  assign n25076 = n25075 ^ n4555 ^ 1'b0 ;
  assign n25077 = n6103 & ~n25076 ;
  assign n25078 = n19477 | n20163 ;
  assign n25079 = n14292 ^ n7567 ^ n3712 ;
  assign n25080 = n25079 ^ n3462 ^ 1'b0 ;
  assign n25081 = ~n14817 & n25080 ;
  assign n25082 = n25081 ^ n22436 ^ 1'b0 ;
  assign n25083 = n6527 & ~n18968 ;
  assign n25084 = n14087 ^ n700 ^ 1'b0 ;
  assign n25085 = n372 & ~n25084 ;
  assign n25086 = ~n1378 & n25085 ;
  assign n25087 = ~n7242 & n19402 ;
  assign n25088 = n16188 ^ n4038 ^ 1'b0 ;
  assign n25089 = n25088 ^ n18464 ^ n1293 ;
  assign n25090 = n8141 ^ n6016 ^ 1'b0 ;
  assign n25091 = n7727 | n25090 ;
  assign n25092 = ( n4977 & n5054 ) | ( n4977 & ~n9923 ) | ( n5054 & ~n9923 ) ;
  assign n25093 = ~n1985 & n3143 ;
  assign n25094 = n25093 ^ n8801 ^ 1'b0 ;
  assign n25095 = n841 & ~n7046 ;
  assign n25096 = ~n25094 & n25095 ;
  assign n25097 = n25096 ^ n20547 ^ 1'b0 ;
  assign n25098 = n4561 | n25097 ;
  assign n25099 = n1148 & ~n5413 ;
  assign n25100 = n21928 ^ n5839 ^ 1'b0 ;
  assign n25101 = n25099 | n25100 ;
  assign n25102 = n22274 | n25101 ;
  assign n25103 = n6156 & ~n6586 ;
  assign n25104 = n7623 & n25103 ;
  assign n25105 = n18672 ^ n17345 ^ n9539 ;
  assign n25106 = n25104 | n25105 ;
  assign n25107 = n25106 ^ n8843 ^ 1'b0 ;
  assign n25108 = n15605 ^ n7520 ^ 1'b0 ;
  assign n25109 = n25108 ^ n16085 ^ n15956 ;
  assign n25110 = n911 & ~n11849 ;
  assign n25111 = n2527 ^ n1073 ^ 1'b0 ;
  assign n25112 = ~n2076 & n25111 ;
  assign n25113 = ~n5929 & n25112 ;
  assign n25114 = ~n25110 & n25113 ;
  assign n25115 = n3691 & ~n25114 ;
  assign n25116 = n1947 & ~n13831 ;
  assign n25117 = ~n7725 & n25116 ;
  assign n25118 = n2227 & n18255 ;
  assign n25119 = n25118 ^ n2053 ^ 1'b0 ;
  assign n25120 = n25119 ^ n7160 ^ n6599 ;
  assign n25121 = n22888 ^ n15363 ^ n8194 ;
  assign n25122 = n6098 | n25121 ;
  assign n25123 = n12699 ^ n9324 ^ 1'b0 ;
  assign n25124 = n14871 & n25123 ;
  assign n25125 = n8771 | n14287 ;
  assign n25126 = n25125 ^ n2694 ^ 1'b0 ;
  assign n25127 = ( n484 & n9643 ) | ( n484 & ~n22427 ) | ( n9643 & ~n22427 ) ;
  assign n25128 = n24959 ^ n16414 ^ 1'b0 ;
  assign n25129 = n727 | n17024 ;
  assign n25130 = ~n339 & n6550 ;
  assign n25131 = ~n9748 & n25130 ;
  assign n25132 = n231 & n340 ;
  assign n25133 = ~n231 & n25132 ;
  assign n25134 = n340 & n782 ;
  assign n25135 = n25133 & n25134 ;
  assign n25136 = n25131 | n25135 ;
  assign n25137 = n25131 & ~n25136 ;
  assign n25138 = n8928 ^ n1905 ^ 1'b0 ;
  assign n25139 = ~n23160 & n25138 ;
  assign n25140 = n25139 ^ n7923 ^ 1'b0 ;
  assign n25141 = n22050 ^ n14047 ^ n5662 ;
  assign n25142 = n17507 | n23389 ;
  assign n25143 = n20128 | n25142 ;
  assign n25144 = n16213 & n25143 ;
  assign n25145 = n2927 | n7515 ;
  assign n25146 = n314 & ~n25145 ;
  assign n25147 = n25146 ^ n9597 ^ 1'b0 ;
  assign n25148 = n25147 ^ n3707 ^ 1'b0 ;
  assign n25149 = n18441 ^ n617 ^ 1'b0 ;
  assign n25150 = n1295 & ~n25149 ;
  assign n25151 = ~n8020 & n25150 ;
  assign n25152 = n24890 ^ n18393 ^ 1'b0 ;
  assign n25153 = ~n11628 & n20285 ;
  assign n25154 = n25153 ^ n5604 ^ 1'b0 ;
  assign n25155 = n6813 & n25154 ;
  assign n25156 = n18321 ^ n911 ^ 1'b0 ;
  assign n25157 = n6127 & n25156 ;
  assign n25158 = n4960 & n7734 ;
  assign n25159 = n20812 ^ n7087 ^ 1'b0 ;
  assign n25160 = n8215 & n25159 ;
  assign n25161 = n25160 ^ n15769 ^ 1'b0 ;
  assign n25162 = n11800 ^ n10439 ^ 1'b0 ;
  assign n25163 = n8635 & ~n25162 ;
  assign n25164 = n25163 ^ n21588 ^ 1'b0 ;
  assign n25165 = n8787 | n11913 ;
  assign n25166 = n25165 ^ n16777 ^ 1'b0 ;
  assign n25167 = ( n5592 & n9477 ) | ( n5592 & ~n16823 ) | ( n9477 & ~n16823 ) ;
  assign n25168 = n25167 ^ n19202 ^ 1'b0 ;
  assign n25169 = n511 | n8648 ;
  assign n25170 = n25169 ^ n3524 ^ 1'b0 ;
  assign n25171 = n3044 & ~n25170 ;
  assign n25172 = n7881 & ~n15109 ;
  assign n25173 = n25172 ^ n3917 ^ 1'b0 ;
  assign n25174 = n25173 ^ n867 ^ n35 ;
  assign n25175 = n13007 ^ n12547 ^ 1'b0 ;
  assign n25178 = n2424 & ~n6946 ;
  assign n25179 = ~n1845 & n25178 ;
  assign n25180 = n4268 & n25179 ;
  assign n25181 = n25180 ^ n12642 ^ 1'b0 ;
  assign n25176 = n5058 & ~n6923 ;
  assign n25177 = ~n287 & n25176 ;
  assign n25182 = n25181 ^ n25177 ^ 1'b0 ;
  assign n25183 = n983 | n1146 ;
  assign n25184 = n2363 & ~n25183 ;
  assign n25185 = ~n4273 & n13682 ;
  assign n25186 = n6650 | n25185 ;
  assign n25187 = n12666 ^ n1732 ^ 1'b0 ;
  assign n25188 = n22541 | n25187 ;
  assign n25189 = ( n1408 & n12025 ) | ( n1408 & n16313 ) | ( n12025 & n16313 ) ;
  assign n25190 = ~n13031 & n13462 ;
  assign n25191 = ~n6473 & n25190 ;
  assign n25192 = n25191 ^ n197 ^ 1'b0 ;
  assign n25193 = n4833 & ~n25192 ;
  assign n25194 = n20858 ^ n10760 ^ 1'b0 ;
  assign n25196 = n6871 ^ n6543 ^ 1'b0 ;
  assign n25195 = n1924 & ~n2634 ;
  assign n25197 = n25196 ^ n25195 ^ 1'b0 ;
  assign n25198 = ~n4593 & n25197 ;
  assign n25199 = ~n18307 & n25198 ;
  assign n25200 = n471 & ~n3777 ;
  assign n25201 = ~n11826 & n25200 ;
  assign n25202 = n5109 & ~n25201 ;
  assign n25203 = ~n5395 & n25202 ;
  assign n25204 = ~n8029 & n14366 ;
  assign n25205 = n25203 & n25204 ;
  assign n25206 = n17153 ^ n16900 ^ 1'b0 ;
  assign n25207 = n7730 | n25206 ;
  assign n25208 = n4187 & ~n8980 ;
  assign n25209 = n25208 ^ n2483 ^ 1'b0 ;
  assign n25210 = n7531 & ~n25209 ;
  assign n25211 = n4095 | n4442 ;
  assign n25212 = n12667 & ~n25211 ;
  assign n25213 = n8919 ^ n8308 ^ 1'b0 ;
  assign n25214 = n9210 & ~n25213 ;
  assign n25216 = n9727 ^ n6088 ^ 1'b0 ;
  assign n25217 = n5192 & ~n25216 ;
  assign n25215 = n21111 ^ n7180 ^ n6216 ;
  assign n25218 = n25217 ^ n25215 ^ 1'b0 ;
  assign n25221 = n25185 ^ n9467 ^ 1'b0 ;
  assign n25222 = n18416 & n25221 ;
  assign n25219 = n9117 ^ n2319 ^ 1'b0 ;
  assign n25220 = ~n5124 & n25219 ;
  assign n25223 = n25222 ^ n25220 ^ 1'b0 ;
  assign n25224 = n5871 | n17653 ;
  assign n25225 = ~n132 & n14441 ;
  assign n25226 = n25225 ^ n12475 ^ 1'b0 ;
  assign n25227 = n10153 | n12789 ;
  assign n25228 = n6777 & ~n25227 ;
  assign n25229 = n25228 ^ n15190 ^ 1'b0 ;
  assign n25230 = ( n23170 & ~n25226 ) | ( n23170 & n25229 ) | ( ~n25226 & n25229 ) ;
  assign n25231 = ~n2512 & n9112 ;
  assign n25232 = n13138 & n25210 ;
  assign n25233 = n7304 ^ n2082 ^ 1'b0 ;
  assign n25234 = n5155 & n25233 ;
  assign n25235 = n13983 ^ n12839 ^ 1'b0 ;
  assign n25236 = ~n3658 & n25235 ;
  assign n25237 = n7676 ^ n666 ^ 1'b0 ;
  assign n25238 = n5845 & n9048 ;
  assign n25239 = n20230 & n25238 ;
  assign n25240 = n25239 ^ n2843 ^ 1'b0 ;
  assign n25241 = ~n10517 & n25240 ;
  assign n25242 = n982 & ~n1211 ;
  assign n25243 = n10544 & n25242 ;
  assign n25244 = n11701 ^ n2262 ^ 1'b0 ;
  assign n25245 = n25243 | n25244 ;
  assign n25246 = n2626 & ~n25245 ;
  assign n25247 = n25246 ^ n1949 ^ 1'b0 ;
  assign n25248 = ~n15759 & n25247 ;
  assign n25249 = n25248 ^ n4547 ^ 1'b0 ;
  assign n25250 = ~n10143 & n13000 ;
  assign n25251 = ~n13612 & n25250 ;
  assign n25252 = ~n25249 & n25251 ;
  assign n25253 = n5510 & n16355 ;
  assign n25254 = ~n11860 & n25253 ;
  assign n25255 = n25254 ^ n16330 ^ 1'b0 ;
  assign n25256 = n20441 & n25255 ;
  assign n25257 = ~n25252 & n25256 ;
  assign n25258 = n11907 & ~n16690 ;
  assign n25259 = n4903 | n10387 ;
  assign n25260 = n3416 & ~n4381 ;
  assign n25261 = ~n10933 & n25260 ;
  assign n25262 = n25261 ^ n16464 ^ 1'b0 ;
  assign n25263 = n5348 | n25262 ;
  assign n25266 = n506 | n16184 ;
  assign n25267 = n25266 ^ n21444 ^ 1'b0 ;
  assign n25264 = n15213 ^ n4916 ^ 1'b0 ;
  assign n25265 = n5031 & ~n25264 ;
  assign n25268 = n25267 ^ n25265 ^ 1'b0 ;
  assign n25269 = ~n9896 & n25268 ;
  assign n25270 = n18315 ^ n10774 ^ 1'b0 ;
  assign n25271 = n7981 & n15324 ;
  assign n25272 = n1731 & n4287 ;
  assign n25273 = n25272 ^ n1724 ^ 1'b0 ;
  assign n25274 = n5099 & ~n5165 ;
  assign n25275 = n25274 ^ n2492 ^ 1'b0 ;
  assign n25276 = n7092 ^ n1771 ^ 1'b0 ;
  assign n25277 = ( n6154 & n25275 ) | ( n6154 & n25276 ) | ( n25275 & n25276 ) ;
  assign n25278 = n13231 | n25277 ;
  assign n25279 = n6036 | n25278 ;
  assign n25280 = n4903 & n14055 ;
  assign n25281 = n9212 & n25280 ;
  assign n25282 = n25281 ^ n11214 ^ n5309 ;
  assign n25283 = n8868 ^ n2498 ^ 1'b0 ;
  assign n25284 = n3970 & ~n25283 ;
  assign n25288 = n819 & ~n2700 ;
  assign n25289 = n4995 & n25288 ;
  assign n25290 = n9334 | n25289 ;
  assign n25285 = n24669 ^ n3987 ^ 1'b0 ;
  assign n25286 = n11680 & n25285 ;
  assign n25287 = n25286 ^ n1966 ^ 1'b0 ;
  assign n25291 = n25290 ^ n25287 ^ 1'b0 ;
  assign n25292 = ~n220 & n2644 ;
  assign n25293 = ~n10581 & n18101 ;
  assign n25294 = n860 | n3674 ;
  assign n25298 = n6446 ^ n755 ^ 1'b0 ;
  assign n25295 = n5940 | n15750 ;
  assign n25296 = n6435 & ~n25295 ;
  assign n25297 = n4608 & ~n25296 ;
  assign n25299 = n25298 ^ n25297 ^ 1'b0 ;
  assign n25300 = ~n5329 & n8405 ;
  assign n25301 = n1167 | n25300 ;
  assign n25302 = n659 | n4712 ;
  assign n25303 = n25302 ^ n6892 ^ 1'b0 ;
  assign n25304 = n25303 ^ n9380 ^ 1'b0 ;
  assign n25305 = n4092 & ~n25304 ;
  assign n25306 = n12696 & n14654 ;
  assign n25307 = ~n9848 & n25306 ;
  assign n25308 = n18073 | n25307 ;
  assign n25309 = n1745 & n25308 ;
  assign n25310 = n10844 ^ n671 ^ 1'b0 ;
  assign n25311 = n2046 | n25310 ;
  assign n25312 = n24304 & ~n25311 ;
  assign n25313 = ~n2352 & n5359 ;
  assign n25314 = n5531 & n25313 ;
  assign n25315 = n25314 ^ n12852 ^ 1'b0 ;
  assign n25316 = n12451 & n13471 ;
  assign n25317 = n18273 ^ n3137 ^ 1'b0 ;
  assign n25318 = n13593 & n25317 ;
  assign n25319 = n10874 ^ n2650 ^ 1'b0 ;
  assign n25320 = n25319 ^ n8705 ^ n3003 ;
  assign n25321 = n2763 & ~n4155 ;
  assign n25322 = ~n17878 & n25321 ;
  assign n25323 = n7292 & ~n11612 ;
  assign n25324 = ~n5199 & n18808 ;
  assign n25325 = ~n6011 & n25324 ;
  assign n25326 = n7940 | n14099 ;
  assign n25327 = n11064 & n13056 ;
  assign n25328 = ~n25326 & n25327 ;
  assign n25329 = ~n3116 & n3605 ;
  assign n25330 = n2598 & n25329 ;
  assign n25331 = n10917 | n25330 ;
  assign n25332 = n25331 ^ n10241 ^ 1'b0 ;
  assign n25333 = n1211 | n25332 ;
  assign n25334 = n18582 ^ n6218 ^ 1'b0 ;
  assign n25335 = n6296 & n25334 ;
  assign n25336 = ~n1946 & n25335 ;
  assign n25337 = n11394 | n17156 ;
  assign n25338 = n3488 ^ n2374 ^ 1'b0 ;
  assign n25339 = n17358 | n25338 ;
  assign n25340 = ( n21 & n2492 ) | ( n21 & n3864 ) | ( n2492 & n3864 ) ;
  assign n25341 = n24027 | n25340 ;
  assign n25342 = n25339 & ~n25341 ;
  assign n25343 = n647 & ~n11812 ;
  assign n25344 = n6060 & n25343 ;
  assign n25345 = n21218 & n25344 ;
  assign n25346 = n3565 | n10570 ;
  assign n25347 = n25346 ^ n3904 ^ 1'b0 ;
  assign n25348 = n4575 & n25347 ;
  assign n25349 = n25348 ^ n3906 ^ 1'b0 ;
  assign n25350 = n15096 | n24209 ;
  assign n25351 = n6154 & ~n25350 ;
  assign n25352 = n16167 ^ n10393 ^ 1'b0 ;
  assign n25353 = n8803 | n25352 ;
  assign n25354 = ~n19915 & n20533 ;
  assign n25355 = n25353 | n25354 ;
  assign n25356 = n8235 & ~n14667 ;
  assign n25358 = ~n7922 & n8885 ;
  assign n25359 = n25358 ^ n16874 ^ 1'b0 ;
  assign n25357 = n20522 | n21781 ;
  assign n25360 = n25359 ^ n25357 ^ 1'b0 ;
  assign n25363 = n14601 & ~n21108 ;
  assign n25361 = ~n1395 & n4315 ;
  assign n25362 = n11546 | n25361 ;
  assign n25364 = n25363 ^ n25362 ^ 1'b0 ;
  assign n25365 = n8211 ^ n1024 ^ 1'b0 ;
  assign n25366 = n3414 & n7020 ;
  assign n25367 = n6028 & n25366 ;
  assign n25369 = n12125 ^ n2080 ^ 1'b0 ;
  assign n25368 = n7396 | n20907 ;
  assign n25370 = n25369 ^ n25368 ^ 1'b0 ;
  assign n25371 = n11885 ^ n6387 ^ 1'b0 ;
  assign n25372 = n25371 ^ n25079 ^ 1'b0 ;
  assign n25373 = ~n7547 & n25372 ;
  assign n25374 = ~n25370 & n25373 ;
  assign n25375 = n269 & n19705 ;
  assign n25376 = ~n1366 & n11185 ;
  assign n25377 = n25376 ^ n8206 ^ 1'b0 ;
  assign n25378 = n25377 ^ n11489 ^ 1'b0 ;
  assign n25379 = n812 | n16513 ;
  assign n25380 = n25379 ^ n7986 ^ 1'b0 ;
  assign n25381 = n21049 & n25380 ;
  assign n25383 = n9854 & ~n10716 ;
  assign n25382 = ~n870 & n14951 ;
  assign n25384 = n25383 ^ n25382 ^ 1'b0 ;
  assign n25385 = n6256 ^ n5526 ^ 1'b0 ;
  assign n25386 = n8449 & ~n25385 ;
  assign n25387 = n25386 ^ n8876 ^ 1'b0 ;
  assign n25388 = n8399 | n10050 ;
  assign n25389 = n8039 & ~n25388 ;
  assign n25390 = ~n9775 & n25389 ;
  assign n25391 = ~n25387 & n25390 ;
  assign n25392 = n25391 ^ n1499 ^ 1'b0 ;
  assign n25393 = ~n25384 & n25392 ;
  assign n25394 = n929 & ~n20001 ;
  assign n25395 = n423 & ~n22107 ;
  assign n25396 = n13869 | n23244 ;
  assign n25397 = n25396 ^ n23427 ^ 1'b0 ;
  assign n25398 = n972 | n2773 ;
  assign n25399 = n25398 ^ n1430 ^ 1'b0 ;
  assign n25400 = ~n2730 & n25399 ;
  assign n25401 = n8869 & n25400 ;
  assign n25402 = n7966 | n14017 ;
  assign n25403 = n3811 & n25402 ;
  assign n25404 = n25403 ^ n14396 ^ n14240 ;
  assign n25405 = ( ~n695 & n2337 ) | ( ~n695 & n2460 ) | ( n2337 & n2460 ) ;
  assign n25406 = n15140 ^ n2634 ^ 1'b0 ;
  assign n25407 = ~n9919 & n25406 ;
  assign n25408 = ~n6229 & n25407 ;
  assign n25409 = n9085 ^ n2726 ^ 1'b0 ;
  assign n25410 = ~n25029 & n25409 ;
  assign n25411 = n7142 | n15163 ;
  assign n25412 = n22118 | n25411 ;
  assign n25413 = n495 & ~n21500 ;
  assign n25414 = n15680 ^ n12677 ^ 1'b0 ;
  assign n25415 = n7919 & n23705 ;
  assign n25416 = n737 & n6784 ;
  assign n25417 = n25416 ^ n21165 ^ 1'b0 ;
  assign n25418 = n8483 | n16756 ;
  assign n25419 = n9319 & ~n11141 ;
  assign n25420 = ~n7820 & n25419 ;
  assign n25421 = n334 & ~n7471 ;
  assign n25422 = n254 & ~n2131 ;
  assign n25423 = n25422 ^ n4868 ^ 1'b0 ;
  assign n25424 = n25423 ^ n16533 ^ 1'b0 ;
  assign n25425 = n5005 ^ n3906 ^ 1'b0 ;
  assign n25426 = n25425 ^ n14473 ^ 1'b0 ;
  assign n25427 = n10879 & ~n25426 ;
  assign n25428 = n10828 ^ n2008 ^ 1'b0 ;
  assign n25429 = ~n7510 & n14480 ;
  assign n25430 = ( ~n582 & n7076 ) | ( ~n582 & n10147 ) | ( n7076 & n10147 ) ;
  assign n25431 = n24583 ^ n11572 ^ 1'b0 ;
  assign n25432 = n25430 | n25431 ;
  assign n25433 = ( n25428 & ~n25429 ) | ( n25428 & n25432 ) | ( ~n25429 & n25432 ) ;
  assign n25435 = ~n4955 & n5145 ;
  assign n25436 = n25435 ^ n23318 ^ 1'b0 ;
  assign n25437 = n15964 & ~n25436 ;
  assign n25438 = ~n6839 & n25437 ;
  assign n25439 = n2574 & n22131 ;
  assign n25440 = n11758 ^ n9928 ^ 1'b0 ;
  assign n25441 = n25439 & ~n25440 ;
  assign n25442 = n25441 ^ n11945 ^ n8000 ;
  assign n25443 = ( n10330 & ~n25438 ) | ( n10330 & n25442 ) | ( ~n25438 & n25442 ) ;
  assign n25434 = n18379 ^ n13737 ^ 1'b0 ;
  assign n25444 = n25443 ^ n25434 ^ 1'b0 ;
  assign n25445 = n564 & n17731 ;
  assign n25446 = n25445 ^ n7729 ^ 1'b0 ;
  assign n25447 = n4990 | n6228 ;
  assign n25448 = ~n9153 & n25447 ;
  assign n25449 = n2427 & n25448 ;
  assign n25450 = n13082 ^ n10056 ^ 1'b0 ;
  assign n25451 = ~n25449 & n25450 ;
  assign n25453 = n3334 | n12576 ;
  assign n25452 = n5123 & ~n13147 ;
  assign n25454 = n25453 ^ n25452 ^ 1'b0 ;
  assign n25455 = n12016 ^ n2989 ^ n1306 ;
  assign n25456 = n25455 ^ n22391 ^ n5072 ;
  assign n25457 = n23495 ^ n20740 ^ n16162 ;
  assign n25458 = n24182 & n25457 ;
  assign n25459 = ~n14087 & n25458 ;
  assign n25460 = n750 | n1697 ;
  assign n25461 = n14360 | n25460 ;
  assign n25462 = n1336 & ~n8031 ;
  assign n25463 = n25462 ^ n3212 ^ 1'b0 ;
  assign n25464 = n7140 & ~n25463 ;
  assign n25465 = ~n907 & n17206 ;
  assign n25466 = n25465 ^ n18033 ^ 1'b0 ;
  assign n25467 = n15757 ^ n11152 ^ 1'b0 ;
  assign n25468 = n2118 | n25467 ;
  assign n25469 = ~n1366 & n5624 ;
  assign n25470 = n25469 ^ n3556 ^ n2973 ;
  assign n25471 = ~n17936 & n25470 ;
  assign n25472 = n5282 ^ n740 ^ 1'b0 ;
  assign n25473 = n14200 & n25472 ;
  assign n25474 = ~n10466 & n17792 ;
  assign n25475 = ~n1134 & n14121 ;
  assign n25476 = ~n11779 & n25475 ;
  assign n25477 = n7167 & n17405 ;
  assign n25478 = n25476 | n25477 ;
  assign n25479 = n5829 | n8024 ;
  assign n25480 = n3822 | n25479 ;
  assign n25481 = n9120 ^ n3254 ^ 1'b0 ;
  assign n25482 = n11524 | n25481 ;
  assign n25483 = n25482 ^ n3240 ^ 1'b0 ;
  assign n25484 = ~n9665 & n25483 ;
  assign n25485 = n24088 | n25484 ;
  assign n25486 = n8494 | n25485 ;
  assign n25487 = n12281 ^ n4328 ^ 1'b0 ;
  assign n25488 = ~n18950 & n25487 ;
  assign n25489 = n13463 & n25488 ;
  assign n25490 = n2336 | n16008 ;
  assign n25491 = n13520 & ~n16675 ;
  assign n25492 = ( n2284 & n20367 ) | ( n2284 & ~n24413 ) | ( n20367 & ~n24413 ) ;
  assign n25497 = n13663 & n17291 ;
  assign n25493 = n2154 | n8550 ;
  assign n25494 = n25493 ^ n5309 ^ 1'b0 ;
  assign n25495 = ( n2405 & n17061 ) | ( n2405 & ~n25494 ) | ( n17061 & ~n25494 ) ;
  assign n25496 = n25495 ^ n13123 ^ n5041 ;
  assign n25498 = n25497 ^ n25496 ^ 1'b0 ;
  assign n25499 = n165 & ~n1329 ;
  assign n25500 = n20254 & ~n25499 ;
  assign n25501 = n14087 ^ n6381 ^ n4280 ;
  assign n25502 = ~n25500 & n25501 ;
  assign n25503 = ~n1275 & n25502 ;
  assign n25504 = ~n1366 & n11068 ;
  assign n25505 = ~n2389 & n25504 ;
  assign n25506 = n12758 & ~n25505 ;
  assign n25507 = n25506 ^ n12013 ^ 1'b0 ;
  assign n25508 = n2796 & ~n12496 ;
  assign n25509 = n23634 ^ n2647 ^ 1'b0 ;
  assign n25510 = n3266 & ~n15415 ;
  assign n25511 = n25510 ^ n6781 ^ 1'b0 ;
  assign n25512 = n3056 | n25511 ;
  assign n25513 = n61 & n1117 ;
  assign n25514 = n25513 ^ n22924 ^ 1'b0 ;
  assign n25515 = ~n3915 & n13266 ;
  assign n25516 = ~n7668 & n25515 ;
  assign n25517 = n2967 | n25516 ;
  assign n25518 = n25517 ^ n23398 ^ 1'b0 ;
  assign n25519 = ~n2227 & n10131 ;
  assign n25520 = n25519 ^ n11452 ^ 1'b0 ;
  assign n25521 = ~n19818 & n25520 ;
  assign n25522 = n24585 | n25521 ;
  assign n25523 = n11512 ^ n9620 ^ 1'b0 ;
  assign n25524 = n1392 & ~n15850 ;
  assign n25525 = n20759 | n23905 ;
  assign n25526 = n25525 ^ n8662 ^ 1'b0 ;
  assign n25527 = n22114 ^ n8573 ^ 1'b0 ;
  assign n25528 = n25526 & ~n25527 ;
  assign n25529 = n13599 ^ n6584 ^ 1'b0 ;
  assign n25530 = ~n2185 & n25529 ;
  assign n25531 = n3349 & n24565 ;
  assign n25532 = n10782 & n11759 ;
  assign n25533 = n6236 & ~n22519 ;
  assign n25534 = n16874 & n25533 ;
  assign n25535 = n23272 ^ n6556 ^ n152 ;
  assign n25536 = n2108 | n25535 ;
  assign n25539 = n1471 | n7237 ;
  assign n25537 = n9940 ^ n8705 ^ 1'b0 ;
  assign n25538 = n24559 & n25537 ;
  assign n25540 = n25539 ^ n25538 ^ 1'b0 ;
  assign n25541 = ~n12025 & n22969 ;
  assign n25542 = ~n8129 & n25541 ;
  assign n25543 = n1081 | n25542 ;
  assign n25544 = n25543 ^ n314 ^ 1'b0 ;
  assign n25545 = n22313 | n25544 ;
  assign n25546 = n412 | n25545 ;
  assign n25547 = n2074 & n25546 ;
  assign n25548 = n10463 & n25547 ;
  assign n25549 = ( n7464 & ~n10475 ) | ( n7464 & n11608 ) | ( ~n10475 & n11608 ) ;
  assign n25550 = n9459 | n25549 ;
  assign n25551 = n16871 & n19007 ;
  assign n25552 = n25425 ^ n16607 ^ n7700 ;
  assign n25553 = n8338 ^ n4778 ^ 1'b0 ;
  assign n25555 = n15454 ^ n1079 ^ 1'b0 ;
  assign n25554 = n19729 ^ n19351 ^ 1'b0 ;
  assign n25556 = n25555 ^ n25554 ^ 1'b0 ;
  assign n25557 = ~n25553 & n25556 ;
  assign n25558 = n1200 | n23087 ;
  assign n25559 = n12150 ^ n9116 ^ n475 ;
  assign n25560 = n5549 | n25559 ;
  assign n25561 = ~n1207 & n16994 ;
  assign n25562 = n17632 ^ n1835 ^ 1'b0 ;
  assign n25563 = n5260 | n10399 ;
  assign n25564 = n25562 | n25563 ;
  assign n25565 = ( n582 & ~n675 ) | ( n582 & n1551 ) | ( ~n675 & n1551 ) ;
  assign n25566 = n3484 & ~n25565 ;
  assign n25567 = x5 & ~n25566 ;
  assign n25568 = n25567 ^ n14058 ^ 1'b0 ;
  assign n25569 = n23428 | n25568 ;
  assign n25570 = n19629 ^ n15587 ^ 1'b0 ;
  assign n25573 = n7813 ^ n712 ^ 1'b0 ;
  assign n25571 = ~n13212 & n24089 ;
  assign n25572 = n18578 & n25571 ;
  assign n25574 = n25573 ^ n25572 ^ 1'b0 ;
  assign n25575 = n3536 ^ n1744 ^ 1'b0 ;
  assign n25576 = n25575 ^ n9205 ^ 1'b0 ;
  assign n25577 = n5197 & ~n11227 ;
  assign n25594 = ~n16683 & n23351 ;
  assign n25595 = n25594 ^ n25112 ^ 1'b0 ;
  assign n25592 = n7589 ^ n65 ^ 1'b0 ;
  assign n25591 = n2201 & n7277 ;
  assign n25593 = n25592 ^ n25591 ^ 1'b0 ;
  assign n25578 = n1310 & n1826 ;
  assign n25579 = n25578 ^ n6045 ^ 1'b0 ;
  assign n25580 = ( n1516 & n11546 ) | ( n1516 & ~n25579 ) | ( n11546 & ~n25579 ) ;
  assign n25583 = n93 & n4350 ;
  assign n25584 = n25583 ^ n2469 ^ 1'b0 ;
  assign n25585 = n7042 ^ n423 ^ 1'b0 ;
  assign n25586 = n25584 & n25585 ;
  assign n25582 = n20032 ^ n9391 ^ n4434 ;
  assign n25587 = n25586 ^ n25582 ^ 1'b0 ;
  assign n25588 = n11232 | n25587 ;
  assign n25581 = n1944 & ~n10351 ;
  assign n25589 = n25588 ^ n25581 ^ n14559 ;
  assign n25590 = ( n7999 & n25580 ) | ( n7999 & n25589 ) | ( n25580 & n25589 ) ;
  assign n25596 = n25595 ^ n25593 ^ n25590 ;
  assign n25597 = ~n11212 & n17176 ;
  assign n25598 = ~n18431 & n25597 ;
  assign n25599 = n22538 ^ n3086 ^ 1'b0 ;
  assign n25600 = n4613 | n10537 ;
  assign n25601 = n10238 | n25600 ;
  assign n25604 = n1570 | n7493 ;
  assign n25605 = n1907 & ~n9495 ;
  assign n25606 = n4214 & n25605 ;
  assign n25607 = n25606 ^ n3442 ^ 1'b0 ;
  assign n25608 = n25604 & n25607 ;
  assign n25602 = n12849 & ~n14500 ;
  assign n25603 = n25602 ^ n18848 ^ 1'b0 ;
  assign n25609 = n25608 ^ n25603 ^ n2940 ;
  assign n25610 = ~n3992 & n24885 ;
  assign n25611 = n25610 ^ n20727 ^ 1'b0 ;
  assign n25612 = ( n1002 & ~n9455 ) | ( n1002 & n16290 ) | ( ~n9455 & n16290 ) ;
  assign n25613 = n10040 & ~n11797 ;
  assign n25614 = n18831 | n25613 ;
  assign n25615 = n1915 | n25614 ;
  assign n25616 = n8334 ^ n3221 ^ 1'b0 ;
  assign n25617 = n25616 ^ n4356 ^ 1'b0 ;
  assign n25618 = ~n25615 & n25617 ;
  assign n25619 = n3429 & n19949 ;
  assign n25620 = n21830 ^ n15095 ^ 1'b0 ;
  assign n25621 = n7578 & n25620 ;
  assign n25622 = n8145 ^ n3686 ^ 1'b0 ;
  assign n25623 = n2095 & ~n25622 ;
  assign n25624 = n12286 | n22252 ;
  assign n25625 = n5979 | n25624 ;
  assign n25626 = n19714 ^ n3347 ^ 1'b0 ;
  assign n25627 = n21218 | n25626 ;
  assign n25628 = n25627 ^ n7344 ^ 1'b0 ;
  assign n25630 = n8610 & n21814 ;
  assign n25631 = n25630 ^ n21535 ^ 1'b0 ;
  assign n25632 = n25631 ^ n13944 ^ n717 ;
  assign n25629 = n2415 | n13302 ;
  assign n25633 = n25632 ^ n25629 ^ 1'b0 ;
  assign n25634 = n11115 ^ n4036 ^ 1'b0 ;
  assign n25635 = n2486 & ~n5890 ;
  assign n25636 = n13186 & ~n14542 ;
  assign n25637 = ~n25635 & n25636 ;
  assign n25638 = n19705 | n25637 ;
  assign n25639 = n22148 | n25638 ;
  assign n25640 = n25639 ^ n9447 ^ 1'b0 ;
  assign n25644 = n12475 ^ n11308 ^ n5986 ;
  assign n25641 = n3726 & n9796 ;
  assign n25642 = n666 | n25641 ;
  assign n25643 = n8555 | n25642 ;
  assign n25645 = n25644 ^ n25643 ^ 1'b0 ;
  assign n25646 = n15102 ^ n13393 ^ 1'b0 ;
  assign n25647 = n25646 ^ n7545 ^ n4264 ;
  assign n25648 = n2856 ^ n233 ^ 1'b0 ;
  assign n25649 = n3052 | n9150 ;
  assign n25650 = n4366 & n15681 ;
  assign n25651 = ~n1157 & n25650 ;
  assign n25652 = n280 & ~n4974 ;
  assign n25653 = n24945 & n25652 ;
  assign n25654 = ~n6917 & n13671 ;
  assign n25655 = n6917 & n25654 ;
  assign n25656 = n468 | n10881 ;
  assign n25657 = n17108 | n25656 ;
  assign n25658 = n10451 & n25657 ;
  assign n25659 = ~n2033 & n25658 ;
  assign n25660 = n18330 | n25659 ;
  assign n25661 = ~n24130 & n25660 ;
  assign n25662 = n25655 & n25661 ;
  assign n25663 = n13343 ^ n13108 ^ 1'b0 ;
  assign n25664 = n16598 & n25663 ;
  assign n25665 = n10646 ^ n4732 ^ 1'b0 ;
  assign n25666 = n25664 & n25665 ;
  assign n25667 = n8332 & ~n24804 ;
  assign n25668 = n25667 ^ n15009 ^ 1'b0 ;
  assign n25669 = n14042 | n15657 ;
  assign n25670 = ( n3155 & n25668 ) | ( n3155 & ~n25669 ) | ( n25668 & ~n25669 ) ;
  assign n25674 = n8506 ^ n4946 ^ 1'b0 ;
  assign n25671 = n12180 ^ n5396 ^ 1'b0 ;
  assign n25672 = n25671 ^ n15136 ^ 1'b0 ;
  assign n25673 = ~n5344 & n25672 ;
  assign n25675 = n25674 ^ n25673 ^ 1'b0 ;
  assign n25676 = n17932 ^ n13545 ^ 1'b0 ;
  assign n25677 = ( n325 & ~n5632 ) | ( n325 & n16145 ) | ( ~n5632 & n16145 ) ;
  assign n25678 = n12740 ^ n1714 ^ 1'b0 ;
  assign n25679 = n181 | n25678 ;
  assign n25680 = n954 & ~n25679 ;
  assign n25681 = n25680 ^ n20136 ^ 1'b0 ;
  assign n25682 = n14345 | n25681 ;
  assign n25683 = n823 & n3568 ;
  assign n25684 = n4119 & n25683 ;
  assign n25685 = ( n1571 & n2121 ) | ( n1571 & n25684 ) | ( n2121 & n25684 ) ;
  assign n25686 = n25685 ^ n6655 ^ 1'b0 ;
  assign n25687 = ~n19918 & n25686 ;
  assign n25688 = n7824 | n11268 ;
  assign n25689 = n25688 ^ n1631 ^ 1'b0 ;
  assign n25690 = n25689 ^ n17370 ^ 1'b0 ;
  assign n25691 = ( ~n3147 & n7414 ) | ( ~n3147 & n11345 ) | ( n7414 & n11345 ) ;
  assign n25692 = n5206 & n13420 ;
  assign n25693 = n18893 ^ n3238 ^ 1'b0 ;
  assign n25694 = n25693 ^ n9694 ^ 1'b0 ;
  assign n25695 = n17079 & n25694 ;
  assign n25696 = n25692 & n25695 ;
  assign n25697 = n3113 | n13189 ;
  assign n25698 = n4141 & ~n25697 ;
  assign n25699 = ~n24911 & n25698 ;
  assign n25700 = n7963 & n12899 ;
  assign n25701 = n919 & n12821 ;
  assign n25702 = ~n11073 & n25701 ;
  assign n25703 = ~n1728 & n13406 ;
  assign n25704 = n14800 & ~n25703 ;
  assign n25705 = ~n14746 & n25704 ;
  assign n25706 = ~n8427 & n25705 ;
  assign n25707 = n13288 & ~n25706 ;
  assign n25708 = n16461 ^ n5484 ^ 1'b0 ;
  assign n25709 = n18950 ^ n4884 ^ 1'b0 ;
  assign n25710 = n700 | n16111 ;
  assign n25711 = n15751 & ~n25710 ;
  assign n25712 = n23397 | n25711 ;
  assign n25713 = n7649 & n15056 ;
  assign n25714 = n25713 ^ n6854 ^ 1'b0 ;
  assign n25715 = ( n614 & n9146 ) | ( n614 & ~n25714 ) | ( n9146 & ~n25714 ) ;
  assign n25716 = n14833 ^ n89 ^ 1'b0 ;
  assign n25717 = n1269 | n25716 ;
  assign n25718 = n13274 ^ n191 ^ 1'b0 ;
  assign n25719 = n11483 | n25718 ;
  assign n25720 = n25717 | n25719 ;
  assign n25721 = ~n14609 & n16640 ;
  assign n25722 = n15602 & n25721 ;
  assign n25724 = n2609 & n4214 ;
  assign n25725 = n3682 & n25724 ;
  assign n25726 = n25725 ^ n8448 ^ 1'b0 ;
  assign n25723 = ~n11616 & n15389 ;
  assign n25727 = n25726 ^ n25723 ^ 1'b0 ;
  assign n25728 = n3751 & n21402 ;
  assign n25732 = ~n6865 & n18803 ;
  assign n25733 = n5953 & n25732 ;
  assign n25729 = n12995 ^ n2427 ^ 1'b0 ;
  assign n25730 = n2845 & n7918 ;
  assign n25731 = n25729 & n25730 ;
  assign n25734 = n25733 ^ n25731 ^ 1'b0 ;
  assign n25735 = n25728 & ~n25734 ;
  assign n25736 = n8560 & ~n15684 ;
  assign n25737 = n25736 ^ n8299 ^ 1'b0 ;
  assign n25739 = n840 | n3444 ;
  assign n25738 = n2650 & ~n4990 ;
  assign n25740 = n25739 ^ n25738 ^ 1'b0 ;
  assign n25741 = n3671 & n18458 ;
  assign n25745 = n1109 ^ x1 ^ 1'b0 ;
  assign n25746 = n10793 | n25745 ;
  assign n25742 = ~n259 & n2593 ;
  assign n25743 = n25742 ^ n721 ^ 1'b0 ;
  assign n25744 = n3833 & ~n25743 ;
  assign n25747 = n25746 ^ n25744 ^ n25418 ;
  assign n25748 = n5306 | n10372 ;
  assign n25749 = ~n21484 & n25748 ;
  assign n25750 = n25749 ^ n24611 ^ n22833 ;
  assign n25751 = n23204 ^ n11244 ^ 1'b0 ;
  assign n25752 = n17156 & ~n25751 ;
  assign n25753 = n21217 | n22884 ;
  assign n25754 = n14960 & ~n25753 ;
  assign n25755 = n3903 & n22668 ;
  assign n25756 = n21949 & n25755 ;
  assign n25758 = n20016 ^ n5150 ^ 1'b0 ;
  assign n25759 = ~n4593 & n25758 ;
  assign n25757 = n13937 ^ n765 ^ 1'b0 ;
  assign n25760 = n25759 ^ n25757 ^ n22005 ;
  assign n25761 = n706 & n7466 ;
  assign n25762 = n7803 & ~n24658 ;
  assign n25763 = n4464 | n6553 ;
  assign n25764 = n6277 ^ n2772 ^ 1'b0 ;
  assign n25765 = n21818 ^ n9190 ^ n4423 ;
  assign n25766 = ~n25764 & n25765 ;
  assign n25767 = n8503 & ~n12045 ;
  assign n25768 = n25767 ^ n15893 ^ 1'b0 ;
  assign n25769 = n25768 ^ n14863 ^ 1'b0 ;
  assign n25770 = n17027 ^ n6184 ^ 1'b0 ;
  assign n25771 = ~n5444 & n25770 ;
  assign n25772 = n17322 ^ n10628 ^ n808 ;
  assign n25773 = n3414 & n22051 ;
  assign n25774 = n20426 ^ n12970 ^ n7722 ;
  assign n25775 = n7658 | n10961 ;
  assign n25776 = n25775 ^ n15681 ^ 1'b0 ;
  assign n25777 = n1743 | n25776 ;
  assign n25778 = ~n8459 & n25777 ;
  assign n25779 = n15511 & ~n25778 ;
  assign n25780 = n25774 & n25779 ;
  assign n25781 = n3331 & ~n3835 ;
  assign n25782 = n25781 ^ n9571 ^ 1'b0 ;
  assign n25783 = n25782 ^ n8776 ^ 1'b0 ;
  assign n25784 = ( n7497 & ~n8452 ) | ( n7497 & n25783 ) | ( ~n8452 & n25783 ) ;
  assign n25785 = n681 & ~n23922 ;
  assign n25786 = n5660 | n25785 ;
  assign n25787 = n7990 & ~n13805 ;
  assign n25788 = n23518 & n25787 ;
  assign n25789 = n25788 ^ n12694 ^ 1'b0 ;
  assign n25790 = n6070 ^ n903 ^ 1'b0 ;
  assign n25791 = n5979 & ~n25790 ;
  assign n25792 = ~n3425 & n6925 ;
  assign n25793 = ~n3140 & n25792 ;
  assign n25794 = n9410 & ~n25793 ;
  assign n25795 = n25794 ^ n9274 ^ 1'b0 ;
  assign n25796 = n25791 & ~n25795 ;
  assign n25798 = n5775 | n7100 ;
  assign n25797 = ( ~n1584 & n4276 ) | ( ~n1584 & n8230 ) | ( n4276 & n8230 ) ;
  assign n25799 = n25798 ^ n25797 ^ 1'b0 ;
  assign n25800 = n10194 | n19051 ;
  assign n25801 = ( ~n12693 & n20620 ) | ( ~n12693 & n25800 ) | ( n20620 & n25800 ) ;
  assign n25802 = ~n3601 & n6533 ;
  assign n25803 = n13559 & ~n25802 ;
  assign n25804 = ~n7148 & n25803 ;
  assign n25805 = n22603 & ~n25804 ;
  assign n25806 = n14964 ^ n4768 ^ n2861 ;
  assign n25807 = n25806 ^ n2091 ^ 1'b0 ;
  assign n25808 = n21681 | n25807 ;
  assign n25809 = ~n4635 & n14483 ;
  assign n25810 = n147 & ~n22086 ;
  assign n25811 = n5282 ^ n1266 ^ 1'b0 ;
  assign n25812 = n868 & ~n25811 ;
  assign n25813 = n12344 ^ n2996 ^ n1187 ;
  assign n25814 = n999 | n12248 ;
  assign n25815 = n25814 ^ n3181 ^ 1'b0 ;
  assign n25816 = n5697 | n25815 ;
  assign n25817 = n3003 | n25816 ;
  assign n25818 = n25817 ^ n8553 ^ 1'b0 ;
  assign n25819 = n25813 & ~n25818 ;
  assign n25820 = n18360 ^ n17300 ^ 1'b0 ;
  assign n25827 = ~n4215 & n4439 ;
  assign n25828 = n25827 ^ n10101 ^ 1'b0 ;
  assign n25821 = n4914 & ~n18544 ;
  assign n25822 = ~n6250 & n25821 ;
  assign n25823 = n7018 & ~n25822 ;
  assign n25824 = n13283 & n25823 ;
  assign n25825 = n25824 ^ n2991 ^ 1'b0 ;
  assign n25826 = n25825 ^ n18376 ^ 1'b0 ;
  assign n25829 = n25828 ^ n25826 ^ 1'b0 ;
  assign n25830 = n3179 & ~n11211 ;
  assign n25831 = n17694 & n25830 ;
  assign n25832 = ~n548 & n2871 ;
  assign n25833 = n548 & n25832 ;
  assign n25834 = ~n2380 & n6287 ;
  assign n25835 = n2380 & n25834 ;
  assign n25836 = n25833 | n25835 ;
  assign n25837 = n2652 | n5016 ;
  assign n25838 = n2652 & ~n25837 ;
  assign n25839 = n2193 | n25838 ;
  assign n25840 = n3150 & ~n4229 ;
  assign n25841 = ~n3150 & n25840 ;
  assign n25842 = n25839 & ~n25841 ;
  assign n25843 = ~n25839 & n25842 ;
  assign n25844 = n8983 | n25843 ;
  assign n25845 = n25843 & ~n25844 ;
  assign n25846 = n24009 | n25845 ;
  assign n25847 = n25846 ^ n25558 ^ 1'b0 ;
  assign n25848 = ~n25836 & n25847 ;
  assign n25849 = ~n6396 & n7349 ;
  assign n25850 = ~n205 & n1351 ;
  assign n25851 = n792 | n19365 ;
  assign n25852 = ~n8482 & n16319 ;
  assign n25853 = n25851 & n25852 ;
  assign n25855 = n9145 ^ n440 ^ 1'b0 ;
  assign n25854 = n1271 | n4698 ;
  assign n25856 = n25855 ^ n25854 ^ 1'b0 ;
  assign n25857 = ( n4103 & n19060 ) | ( n4103 & n25856 ) | ( n19060 & n25856 ) ;
  assign n25858 = ~n1172 & n23570 ;
  assign n25859 = n7042 & ~n9917 ;
  assign n25860 = n11369 ^ n9536 ^ n4926 ;
  assign n25861 = ~n5965 & n10812 ;
  assign n25862 = n16371 ^ n5126 ^ 1'b0 ;
  assign n25863 = ~n25861 & n25862 ;
  assign n25864 = n12449 & ~n25863 ;
  assign n25865 = ~n24638 & n25864 ;
  assign n25866 = n22427 ^ n9014 ^ 1'b0 ;
  assign n25867 = n21241 | n25866 ;
  assign n25868 = n4801 & ~n5166 ;
  assign n25871 = n3066 & n6331 ;
  assign n25872 = n1574 & n5802 ;
  assign n25873 = ~n25871 & n25872 ;
  assign n25874 = n25873 ^ n3671 ^ 1'b0 ;
  assign n25875 = n7873 & ~n25874 ;
  assign n25869 = n11740 ^ n8788 ^ 1'b0 ;
  assign n25870 = ~n16392 & n25869 ;
  assign n25876 = n25875 ^ n25870 ^ 1'b0 ;
  assign n25877 = n23803 ^ n3442 ^ 1'b0 ;
  assign n25878 = n36 | n16923 ;
  assign n25879 = n4727 & n25878 ;
  assign n25880 = n19563 | n22704 ;
  assign n25882 = ~n6543 & n7402 ;
  assign n25881 = n6573 & ~n25862 ;
  assign n25883 = n25882 ^ n25881 ^ 1'b0 ;
  assign n25884 = n25880 & n25883 ;
  assign n25885 = n16743 ^ n6829 ^ 1'b0 ;
  assign n25886 = n25885 ^ n13059 ^ 1'b0 ;
  assign n25887 = ~n14880 & n25886 ;
  assign n25888 = n19118 & ~n24700 ;
  assign n25889 = n2591 ^ n956 ^ 1'b0 ;
  assign n25890 = ~n1174 & n25889 ;
  assign n25891 = n10796 ^ n5150 ^ 1'b0 ;
  assign n25892 = n19113 | n25891 ;
  assign n25893 = ( n13097 & ~n25890 ) | ( n13097 & n25892 ) | ( ~n25890 & n25892 ) ;
  assign n25894 = n12015 & n24686 ;
  assign n25895 = n25894 ^ n15782 ^ 1'b0 ;
  assign n25896 = ( n5743 & n7402 ) | ( n5743 & ~n25895 ) | ( n7402 & ~n25895 ) ;
  assign n25897 = n633 & ~n1455 ;
  assign n25898 = n2855 | n25897 ;
  assign n25899 = n25898 ^ n10484 ^ 1'b0 ;
  assign n25900 = n19456 ^ n12000 ^ n1531 ;
  assign n25901 = n25900 ^ n1289 ^ 1'b0 ;
  assign n25902 = n21918 ^ n11081 ^ 1'b0 ;
  assign n25903 = n13425 & ~n14058 ;
  assign n25904 = ~n5282 & n23295 ;
  assign n25905 = n25760 ^ n7265 ^ 1'b0 ;
  assign n25906 = n745 & ~n6818 ;
  assign n25907 = n22994 ^ n8960 ^ 1'b0 ;
  assign n25908 = n6281 & n25907 ;
  assign n25909 = n10814 | n20175 ;
  assign n25910 = n972 & n5401 ;
  assign n25911 = n15130 & n17781 ;
  assign n25912 = n5864 & n24107 ;
  assign n25913 = n25912 ^ n4357 ^ 1'b0 ;
  assign n25914 = n25913 ^ n19934 ^ n18328 ;
  assign n25915 = n1538 | n10577 ;
  assign n25916 = n25915 ^ n787 ^ 1'b0 ;
  assign n25917 = n5999 | n25916 ;
  assign n25918 = n3763 & ~n25917 ;
  assign n25919 = n25918 ^ n1845 ^ 1'b0 ;
  assign n25920 = n11836 & n13422 ;
  assign n25921 = n25919 & n25920 ;
  assign n25922 = n8450 ^ n8313 ^ n4926 ;
  assign n25923 = n6669 & ~n9461 ;
  assign n25924 = n25923 ^ n17816 ^ 1'b0 ;
  assign n25925 = n1823 & ~n9779 ;
  assign n25926 = n4252 & n7076 ;
  assign n25927 = n23854 ^ n17874 ^ n10052 ;
  assign n25928 = ~n5084 & n25927 ;
  assign n25929 = n14958 & ~n25928 ;
  assign n25930 = ~n15547 & n25929 ;
  assign n25931 = n6551 & n25930 ;
  assign n25932 = n2120 & ~n7015 ;
  assign n25933 = n10452 & n25932 ;
  assign n25934 = n14873 | n25933 ;
  assign n25935 = n25934 ^ n2267 ^ 1'b0 ;
  assign n25936 = ~n12636 & n19799 ;
  assign n25937 = n25936 ^ n13174 ^ 1'b0 ;
  assign n25938 = n1273 & n24749 ;
  assign n25939 = n5779 ^ n5170 ^ 1'b0 ;
  assign n25940 = n302 & ~n25939 ;
  assign n25941 = ~n22158 & n25940 ;
  assign n25942 = ~n4082 & n4341 ;
  assign n25943 = ~n11934 & n25942 ;
  assign n25944 = n23456 ^ n5039 ^ 1'b0 ;
  assign n25945 = n6770 ^ n1802 ^ 1'b0 ;
  assign n25946 = n8832 ^ n2063 ^ 1'b0 ;
  assign n25947 = n2068 | n7627 ;
  assign n25948 = n25947 ^ n6062 ^ 1'b0 ;
  assign n25949 = n8033 ^ n3777 ^ 1'b0 ;
  assign n25950 = n25948 | n25949 ;
  assign n25951 = n1561 & n25950 ;
  assign n25952 = n5851 ^ n3848 ^ 1'b0 ;
  assign n25953 = n6181 & n25952 ;
  assign n25954 = n25953 ^ n24491 ^ 1'b0 ;
  assign n25955 = n511 & ~n25954 ;
  assign n25956 = ( n968 & n6626 ) | ( n968 & ~n16157 ) | ( n6626 & ~n16157 ) ;
  assign n25957 = ( n11737 & n18779 ) | ( n11737 & ~n25956 ) | ( n18779 & ~n25956 ) ;
  assign n25958 = n4545 ^ n2522 ^ 1'b0 ;
  assign n25959 = n15915 ^ n12280 ^ 1'b0 ;
  assign n25960 = ~n25958 & n25959 ;
  assign n25961 = n20410 ^ n2170 ^ 1'b0 ;
  assign n25962 = n8971 | n25961 ;
  assign n25963 = n20648 ^ n20355 ^ 1'b0 ;
  assign n25964 = n11717 ^ n205 ^ 1'b0 ;
  assign n25967 = ~n2030 & n2292 ;
  assign n25968 = n12307 & n25967 ;
  assign n25965 = n25579 ^ n20835 ^ 1'b0 ;
  assign n25966 = n20243 & n25965 ;
  assign n25969 = n25968 ^ n25966 ^ 1'b0 ;
  assign n25970 = ~n2036 & n12821 ;
  assign n25971 = n2097 & ~n2382 ;
  assign n25972 = ~n25970 & n25971 ;
  assign n25973 = ( n1123 & ~n2309 ) | ( n1123 & n11187 ) | ( ~n2309 & n11187 ) ;
  assign n25974 = n20974 & ~n25973 ;
  assign n25975 = ( n5977 & n11162 ) | ( n5977 & ~n25974 ) | ( n11162 & ~n25974 ) ;
  assign n25976 = n6045 & ~n6469 ;
  assign n25977 = n23253 ^ n12494 ^ 1'b0 ;
  assign n25978 = n451 & ~n12816 ;
  assign n25979 = n3026 | n20911 ;
  assign n25980 = n25978 | n25979 ;
  assign n25981 = ( ~n2641 & n6437 ) | ( ~n2641 & n19638 ) | ( n6437 & n19638 ) ;
  assign n25982 = n25981 ^ n31 ^ 1'b0 ;
  assign n25983 = ~n4411 & n25982 ;
  assign n25990 = n150 | n607 ;
  assign n25991 = n150 & ~n25990 ;
  assign n25992 = ~n2170 & n3600 ;
  assign n25993 = n25991 & n25992 ;
  assign n25994 = n10183 | n25993 ;
  assign n25988 = n11755 & n12077 ;
  assign n25989 = n16780 | n25988 ;
  assign n25984 = ~n10950 & n15984 ;
  assign n25985 = ~n15984 & n25984 ;
  assign n25986 = ~n16247 & n18917 ;
  assign n25987 = n25985 & n25986 ;
  assign n25995 = n25994 ^ n25989 ^ n25987 ;
  assign n25996 = n978 & ~n7375 ;
  assign n25997 = n25996 ^ n14720 ^ 1'b0 ;
  assign n25998 = n19382 ^ n2433 ^ 1'b0 ;
  assign n25999 = n25998 ^ n20604 ^ 1'b0 ;
  assign n26000 = ~n4147 & n25999 ;
  assign n26001 = n9375 ^ n4919 ^ 1'b0 ;
  assign n26002 = n25075 & n26001 ;
  assign n26003 = n3408 & n26002 ;
  assign n26004 = ~n23133 & n26003 ;
  assign n26005 = n10227 ^ n3386 ^ 1'b0 ;
  assign n26006 = ~n8156 & n26005 ;
  assign n26007 = n26006 ^ n9102 ^ 1'b0 ;
  assign n26008 = n16871 ^ n11908 ^ n6813 ;
  assign n26009 = n18838 ^ n2199 ^ 1'b0 ;
  assign n26010 = n27 & n14727 ;
  assign n26011 = n26010 ^ n3262 ^ 1'b0 ;
  assign n26012 = n10180 & n20013 ;
  assign n26013 = n620 ^ n440 ^ 1'b0 ;
  assign n26014 = n14484 ^ n11691 ^ 1'b0 ;
  assign n26015 = n26013 & n26014 ;
  assign n26016 = n733 & ~n1420 ;
  assign n26017 = ~n733 & n26016 ;
  assign n26018 = n12550 & ~n26017 ;
  assign n26019 = ~n12550 & n26018 ;
  assign n26020 = n1049 | n6595 ;
  assign n26021 = n2355 | n26020 ;
  assign n26022 = n26021 ^ n7624 ^ n7515 ;
  assign n26023 = n1747 & ~n13478 ;
  assign n26024 = ~n16059 & n26023 ;
  assign n26025 = n10489 ^ n3811 ^ 1'b0 ;
  assign n26026 = ~n26024 & n26025 ;
  assign n26027 = n22218 ^ n19726 ^ 1'b0 ;
  assign n26028 = n15308 ^ n13299 ^ 1'b0 ;
  assign n26029 = ~n4604 & n14612 ;
  assign n26030 = n26029 ^ n19714 ^ 1'b0 ;
  assign n26031 = n1024 & n20615 ;
  assign n26032 = n26031 ^ n24898 ^ 1'b0 ;
  assign n26033 = n13436 ^ n3809 ^ 1'b0 ;
  assign n26034 = n2524 & ~n26033 ;
  assign n26035 = ~n14904 & n26034 ;
  assign n26040 = ~n8847 & n9746 ;
  assign n26037 = n3775 & ~n16353 ;
  assign n26038 = ~n7388 & n26037 ;
  assign n26039 = n1369 & n26038 ;
  assign n26036 = ~n8292 & n14171 ;
  assign n26041 = n26040 ^ n26039 ^ n26036 ;
  assign n26042 = n22337 & ~n24632 ;
  assign n26043 = n1439 & ~n10220 ;
  assign n26044 = n26043 ^ n1460 ^ 1'b0 ;
  assign n26045 = n7759 ^ n7368 ^ 1'b0 ;
  assign n26046 = n4583 & n12468 ;
  assign n26047 = n20533 & ~n26046 ;
  assign n26048 = n12661 & n26047 ;
  assign n26049 = n26045 & ~n26048 ;
  assign n26050 = ~n25532 & n26049 ;
  assign n26051 = n1159 & n2033 ;
  assign n26052 = n4044 | n7413 ;
  assign n26053 = ~n428 & n5021 ;
  assign n26054 = n867 & n26053 ;
  assign n26055 = n26054 ^ n10411 ^ n1631 ;
  assign n26056 = n14672 | n26055 ;
  assign n26057 = n26052 & ~n26056 ;
  assign n26058 = n26057 ^ n10477 ^ 1'b0 ;
  assign n26059 = n13340 & n26058 ;
  assign n26060 = ~n5658 & n9143 ;
  assign n26061 = n16356 | n26060 ;
  assign n26062 = n26061 ^ n13096 ^ 1'b0 ;
  assign n26063 = n5747 ^ n4267 ^ 1'b0 ;
  assign n26066 = n1544 ^ n270 ^ 1'b0 ;
  assign n26067 = n2458 ^ n205 ^ 1'b0 ;
  assign n26068 = ~n26066 & n26067 ;
  assign n26069 = ~n2044 & n26068 ;
  assign n26064 = n231 | n5264 ;
  assign n26065 = n12133 & ~n26064 ;
  assign n26070 = n26069 ^ n26065 ^ 1'b0 ;
  assign n26071 = n3657 & n3893 ;
  assign n26072 = n7405 | n24804 ;
  assign n26073 = n26072 ^ n2796 ^ 1'b0 ;
  assign n26074 = n26071 & n26073 ;
  assign n26075 = n25466 ^ n9096 ^ 1'b0 ;
  assign n26076 = ( n112 & n7527 ) | ( n112 & ~n21806 ) | ( n7527 & ~n21806 ) ;
  assign n26077 = x1 & n54 ;
  assign n26078 = ~n54 & n26077 ;
  assign n26079 = n26078 ^ n11934 ^ 1'b0 ;
  assign n26081 = ~n7759 & n21212 ;
  assign n26082 = ~n21212 & n26081 ;
  assign n26080 = ~n2649 & n19776 ;
  assign n26083 = n26082 ^ n26080 ^ 1'b0 ;
  assign n26084 = n26079 & n26083 ;
  assign n26085 = ~n26079 & n26084 ;
  assign n26086 = n1912 & n4949 ;
  assign n26087 = ~n4949 & n26086 ;
  assign n26088 = n14864 & n26087 ;
  assign n26089 = n26088 ^ n12038 ^ 1'b0 ;
  assign n26090 = n20158 ^ n2060 ^ 1'b0 ;
  assign n26091 = n26090 ^ n12919 ^ 1'b0 ;
  assign n26092 = n24049 & n26091 ;
  assign n26093 = ~n26089 & n26092 ;
  assign n26094 = n7403 & ~n11967 ;
  assign n26095 = ~n18936 & n26094 ;
  assign n26096 = ~n2780 & n4564 ;
  assign n26097 = n19367 & n26096 ;
  assign n26098 = n12397 ^ n10603 ^ 1'b0 ;
  assign n26099 = n922 | n3182 ;
  assign n26100 = n6447 | n26099 ;
  assign n26101 = n1745 & n19427 ;
  assign n26102 = n26100 & ~n26101 ;
  assign n26103 = ~n26098 & n26102 ;
  assign n26104 = n16898 ^ n192 ^ 1'b0 ;
  assign n26105 = ~n1771 & n21255 ;
  assign n26106 = n11456 | n21307 ;
  assign n26107 = ~n6296 & n11741 ;
  assign n26108 = n16933 & n26107 ;
  assign n26109 = n16294 ^ n11312 ^ 1'b0 ;
  assign n26110 = n4747 ^ n2147 ^ 1'b0 ;
  assign n26111 = n13105 | n26110 ;
  assign n26112 = n6193 & n13023 ;
  assign n26113 = ( n2407 & n5001 ) | ( n2407 & ~n24492 ) | ( n5001 & ~n24492 ) ;
  assign n26114 = n18044 ^ n4754 ^ 1'b0 ;
  assign n26115 = n20340 & ~n26114 ;
  assign n26116 = n4745 ^ n852 ^ 1'b0 ;
  assign n26117 = n12640 & n20119 ;
  assign n26118 = n26117 ^ n14422 ^ 1'b0 ;
  assign n26119 = n15215 & n26118 ;
  assign n26120 = n26119 ^ n12604 ^ n9844 ;
  assign n26121 = ( n727 & ~n21200 ) | ( n727 & n26120 ) | ( ~n21200 & n26120 ) ;
  assign n26122 = ( ~n8740 & n9753 ) | ( ~n8740 & n12593 ) | ( n9753 & n12593 ) ;
  assign n26123 = ~n8625 & n12422 ;
  assign n26124 = n13454 & n26123 ;
  assign n26125 = n1513 & ~n1878 ;
  assign n26126 = ~n12970 & n26125 ;
  assign n26127 = n9943 & ~n26126 ;
  assign n26128 = ~n11283 & n23155 ;
  assign n26129 = ( n3437 & n8273 ) | ( n3437 & ~n26098 ) | ( n8273 & ~n26098 ) ;
  assign n26130 = n6434 & n6745 ;
  assign n26131 = ~n16931 & n26130 ;
  assign n26132 = n22985 ^ n11515 ^ 1'b0 ;
  assign n26133 = n1354 | n26132 ;
  assign n26134 = n10036 | n11697 ;
  assign n26135 = n7187 | n25668 ;
  assign n26136 = n26135 ^ n9962 ^ 1'b0 ;
  assign n26137 = n21516 ^ n13941 ^ n10500 ;
  assign n26138 = n15782 ^ n1023 ^ 1'b0 ;
  assign n26139 = n3584 & n16071 ;
  assign n26140 = n26138 & n26139 ;
  assign n26141 = n5064 ^ n4857 ^ 1'b0 ;
  assign n26142 = ~n8749 & n25272 ;
  assign n26143 = n7757 & ~n8274 ;
  assign n26144 = ~n901 & n3826 ;
  assign n26145 = ~n3826 & n26144 ;
  assign n26146 = n26145 ^ n22187 ^ 1'b0 ;
  assign n26147 = n1991 & n2900 ;
  assign n26148 = ~n2900 & n26147 ;
  assign n26149 = n15856 | n26148 ;
  assign n26150 = n26146 | n26149 ;
  assign n26151 = ( n2121 & ~n15220 ) | ( n2121 & n26150 ) | ( ~n15220 & n26150 ) ;
  assign n26152 = n24830 ^ n1416 ^ 1'b0 ;
  assign n26153 = n16804 ^ n14460 ^ 1'b0 ;
  assign n26154 = ~n8459 & n26153 ;
  assign n26155 = ~n12307 & n13607 ;
  assign n26156 = n4215 & n26155 ;
  assign n26157 = n717 ^ n105 ^ 1'b0 ;
  assign n26158 = n365 & ~n26157 ;
  assign n26159 = n11431 ^ n2715 ^ 1'b0 ;
  assign n26160 = ~n26158 & n26159 ;
  assign n26161 = n26160 ^ n1933 ^ 1'b0 ;
  assign n26162 = n15708 | n26161 ;
  assign n26163 = n13342 ^ n6576 ^ n2462 ;
  assign n26164 = n7877 ^ n2610 ^ 1'b0 ;
  assign n26165 = n14288 & n26164 ;
  assign n26166 = n26165 ^ n15966 ^ n2154 ;
  assign n26167 = n10882 | n12132 ;
  assign n26168 = n26167 ^ n352 ^ 1'b0 ;
  assign n26169 = n326 & ~n6931 ;
  assign n26170 = n3121 | n26169 ;
  assign n26171 = n26170 ^ n924 ^ 1'b0 ;
  assign n26172 = n11169 ^ n1264 ^ 1'b0 ;
  assign n26173 = n10021 | n12863 ;
  assign n26174 = n12578 | n26173 ;
  assign n26175 = n26174 ^ n12974 ^ 1'b0 ;
  assign n26176 = ~n8962 & n26175 ;
  assign n26177 = n528 & ~n3193 ;
  assign n26178 = ~n2987 & n26177 ;
  assign n26179 = n26178 ^ n6408 ^ 1'b0 ;
  assign n26180 = n2097 | n26179 ;
  assign n26181 = n2444 & ~n26180 ;
  assign n26182 = ~n1196 & n12228 ;
  assign n26183 = n26182 ^ n17421 ^ 1'b0 ;
  assign n26184 = n26183 ^ n8042 ^ 1'b0 ;
  assign n26185 = n8843 & n19163 ;
  assign n26186 = n21786 ^ n15166 ^ 1'b0 ;
  assign n26187 = n24162 & ~n26186 ;
  assign n26188 = n15499 & ~n17622 ;
  assign n26189 = ~n9645 & n26188 ;
  assign n26190 = n9178 & ~n26189 ;
  assign n26194 = ~n2656 & n22624 ;
  assign n26191 = ~n989 & n2176 ;
  assign n26192 = n26191 ^ n459 ^ 1'b0 ;
  assign n26193 = ~n152 & n26192 ;
  assign n26195 = n26194 ^ n26193 ^ 1'b0 ;
  assign n26196 = ( n4685 & n6838 ) | ( n4685 & n7927 ) | ( n6838 & n7927 ) ;
  assign n26197 = n26196 ^ n23065 ^ 1'b0 ;
  assign n26198 = n9601 | n26197 ;
  assign n26199 = n5765 & ~n6399 ;
  assign n26200 = n6625 & n22448 ;
  assign n26201 = n16508 | n26200 ;
  assign n26202 = ~n9222 & n16221 ;
  assign n26203 = n1346 & n26202 ;
  assign n26204 = n26203 ^ n2662 ^ 1'b0 ;
  assign n26205 = n21150 | n22522 ;
  assign n26206 = n23734 & ~n26205 ;
  assign n26207 = n2818 | n21573 ;
  assign n26208 = n26207 ^ n21432 ^ n13625 ;
  assign n26209 = n16085 & n26208 ;
  assign n26210 = n3576 | n14676 ;
  assign n26211 = n26210 ^ n18579 ^ 1'b0 ;
  assign n26212 = n6456 & n26211 ;
  assign n26213 = n14183 ^ n8901 ^ 1'b0 ;
  assign n26214 = n26212 & ~n26213 ;
  assign n26215 = n2562 & n23936 ;
  assign n26216 = ~n18885 & n26215 ;
  assign n26217 = n8411 ^ n2655 ^ 1'b0 ;
  assign n26218 = n26217 ^ n23556 ^ 1'b0 ;
  assign n26219 = n22857 & ~n26218 ;
  assign n26220 = ~n851 & n17496 ;
  assign n26221 = n26220 ^ n19529 ^ 1'b0 ;
  assign n26222 = n11425 ^ n10370 ^ 1'b0 ;
  assign n26223 = n4341 & ~n26222 ;
  assign n26224 = n26223 ^ n12551 ^ 1'b0 ;
  assign n26225 = ~n13488 & n26224 ;
  assign n26226 = n26225 ^ n10552 ^ n9334 ;
  assign n26227 = ~n22739 & n26226 ;
  assign n26228 = n1695 & ~n5579 ;
  assign n26229 = n26228 ^ n11637 ^ 1'b0 ;
  assign n26230 = n17108 ^ n6761 ^ 1'b0 ;
  assign n26231 = n3680 & n26230 ;
  assign n26232 = n26231 ^ n5810 ^ 1'b0 ;
  assign n26233 = n26229 & ~n26232 ;
  assign n26234 = n3730 ^ n574 ^ 1'b0 ;
  assign n26235 = n8948 & n26234 ;
  assign n26236 = ~n184 & n26235 ;
  assign n26237 = ~n26233 & n26236 ;
  assign n26238 = n6799 | n9680 ;
  assign n26239 = n26238 ^ n2954 ^ 1'b0 ;
  assign n26240 = n26239 ^ n19464 ^ 1'b0 ;
  assign n26241 = n250 | n26240 ;
  assign n26242 = n21664 ^ n13194 ^ 1'b0 ;
  assign n26243 = n18626 ^ n16056 ^ n8677 ;
  assign n26244 = n26243 ^ n9150 ^ 1'b0 ;
  assign n26245 = n23688 ^ n6182 ^ 1'b0 ;
  assign n26248 = n6979 | n12377 ;
  assign n26249 = n11776 & ~n26248 ;
  assign n26247 = n4788 & n12851 ;
  assign n26250 = n26249 ^ n26247 ^ 1'b0 ;
  assign n26246 = ~n7999 & n16910 ;
  assign n26251 = n26250 ^ n26246 ^ n19910 ;
  assign n26252 = n1580 & ~n20725 ;
  assign n26253 = n26252 ^ n25224 ^ 1'b0 ;
  assign n26255 = n2262 ^ n1811 ^ 1'b0 ;
  assign n26256 = n4561 | n26255 ;
  assign n26254 = ~n4097 & n15047 ;
  assign n26257 = n26256 ^ n26254 ^ 1'b0 ;
  assign n26258 = ~n10790 & n19283 ;
  assign n26259 = n26257 & ~n26258 ;
  assign n26260 = ~n3045 & n14785 ;
  assign n26261 = ~n14785 & n26260 ;
  assign n26262 = n119 | n26261 ;
  assign n26263 = n119 & ~n26262 ;
  assign n26264 = n7048 & ~n26263 ;
  assign n26265 = ~n7048 & n26264 ;
  assign n26266 = n2353 | n26265 ;
  assign n26267 = n83 & n574 ;
  assign n26268 = ~n83 & n26267 ;
  assign n26269 = n26266 | n26268 ;
  assign n26270 = n26266 & ~n26269 ;
  assign n26271 = n24050 & ~n26270 ;
  assign n26272 = ~n532 & n26271 ;
  assign n26273 = n4313 ^ n2821 ^ 1'b0 ;
  assign n26274 = ~n3044 & n26273 ;
  assign n26275 = ( n5249 & n14153 ) | ( n5249 & n26274 ) | ( n14153 & n26274 ) ;
  assign n26276 = n26275 ^ n11692 ^ 1'b0 ;
  assign n26277 = n14203 & n14998 ;
  assign n26278 = ~n14998 & n26277 ;
  assign n26279 = n9998 & ~n26278 ;
  assign n26280 = n19882 ^ n286 ^ 1'b0 ;
  assign n26281 = ( ~n3023 & n14500 ) | ( ~n3023 & n26280 ) | ( n14500 & n26280 ) ;
  assign n26282 = n1842 & ~n18964 ;
  assign n26283 = ~n4676 & n26282 ;
  assign n26284 = n18195 ^ n15807 ^ 1'b0 ;
  assign n26285 = n3713 | n26284 ;
  assign n26286 = n6159 & n9268 ;
  assign n26287 = n6741 | n26286 ;
  assign n26288 = n26287 ^ n7471 ^ 1'b0 ;
  assign n26289 = n3909 & ~n26288 ;
  assign n26290 = n26289 ^ n11714 ^ 1'b0 ;
  assign n26291 = ~n4019 & n17935 ;
  assign n26292 = n2078 & n7632 ;
  assign n26293 = n5482 & ~n26292 ;
  assign n26294 = n5249 & ~n11366 ;
  assign n26295 = ~n26293 & n26294 ;
  assign n26296 = n5154 | n24228 ;
  assign n26297 = n489 & n3558 ;
  assign n26298 = n6522 ^ n1154 ^ 1'b0 ;
  assign n26299 = ( n3971 & ~n4147 ) | ( n3971 & n26298 ) | ( ~n4147 & n26298 ) ;
  assign n26300 = n5268 & n26299 ;
  assign n26301 = n343 & n26300 ;
  assign n26302 = n26297 & ~n26301 ;
  assign n26303 = n24146 & n26302 ;
  assign n26304 = n21279 ^ n1216 ^ 1'b0 ;
  assign n26305 = n22540 | n24136 ;
  assign n26306 = n2872 & ~n26305 ;
  assign n26307 = n7256 & n25370 ;
  assign n26308 = ~n2517 & n8775 ;
  assign n26309 = n2517 & n26308 ;
  assign n26310 = n2428 & ~n26309 ;
  assign n26311 = n26310 ^ n13661 ^ 1'b0 ;
  assign n26312 = n13393 & ~n14343 ;
  assign n26313 = n4583 & n13152 ;
  assign n26314 = n26312 & n26313 ;
  assign n26315 = n3665 & ~n6919 ;
  assign n26316 = n26315 ^ n12906 ^ 1'b0 ;
  assign n26317 = n26314 & ~n26316 ;
  assign n26318 = n1700 | n3583 ;
  assign n26319 = n18142 & n26318 ;
  assign n26320 = n26319 ^ n533 ^ 1'b0 ;
  assign n26321 = ~n7998 & n26320 ;
  assign n26322 = n10085 ^ n192 ^ 1'b0 ;
  assign n26323 = ~n12118 & n26322 ;
  assign n26324 = ( n16430 & n17834 ) | ( n16430 & n26323 ) | ( n17834 & n26323 ) ;
  assign n26325 = n26324 ^ n7973 ^ 1'b0 ;
  assign n26326 = n8450 & n11532 ;
  assign n26327 = n26326 ^ n19362 ^ 1'b0 ;
  assign n26328 = n15603 ^ n4018 ^ 1'b0 ;
  assign n26329 = n398 & n15614 ;
  assign n26330 = n26329 ^ n8819 ^ 1'b0 ;
  assign n26331 = n1131 | n4931 ;
  assign n26332 = n26330 | n26331 ;
  assign n26333 = n8008 & ~n8915 ;
  assign n26334 = n6851 ^ n5179 ^ 1'b0 ;
  assign n26335 = n22601 & ~n26334 ;
  assign n26336 = ~n8958 & n10692 ;
  assign n26337 = n12922 & n26336 ;
  assign n26338 = n5363 | n18393 ;
  assign n26339 = ~n15010 & n22073 ;
  assign n26340 = n26339 ^ n1516 ^ 1'b0 ;
  assign n26341 = n26340 ^ n17100 ^ n6145 ;
  assign n26342 = ~n4087 & n12835 ;
  assign n26343 = n18831 ^ n8879 ^ 1'b0 ;
  assign n26344 = n2211 & ~n26343 ;
  assign n26345 = n16560 & n21081 ;
  assign n26346 = n26345 ^ n11727 ^ 1'b0 ;
  assign n26347 = n18167 | n26346 ;
  assign n26348 = n7494 & ~n26347 ;
  assign n26349 = n17038 ^ n10728 ^ n1293 ;
  assign n26350 = ( n4261 & n4698 ) | ( n4261 & n24732 ) | ( n4698 & n24732 ) ;
  assign n26351 = n26350 ^ n12832 ^ 1'b0 ;
  assign n26352 = ~n13204 & n23445 ;
  assign n26353 = n15404 | n16430 ;
  assign n26354 = n26353 ^ n12249 ^ 1'b0 ;
  assign n26355 = n22291 ^ n13011 ^ n431 ;
  assign n26356 = n712 & n1335 ;
  assign n26357 = n26356 ^ n919 ^ 1'b0 ;
  assign n26358 = n26357 ^ n423 ^ 1'b0 ;
  assign n26359 = n6922 | n26358 ;
  assign n26360 = ~n19911 & n21350 ;
  assign n26361 = n11980 & n26360 ;
  assign n26362 = n26359 & n26361 ;
  assign n26363 = ~n11489 & n26362 ;
  assign n26364 = ~n850 & n12988 ;
  assign n26365 = n1150 & n26364 ;
  assign n26366 = n26365 ^ n12483 ^ 1'b0 ;
  assign n26367 = ~n780 & n1513 ;
  assign n26368 = n26367 ^ n3726 ^ 1'b0 ;
  assign n26369 = ~n5206 & n26368 ;
  assign n26370 = n26369 ^ n13279 ^ 1'b0 ;
  assign n26371 = n10519 & ~n26370 ;
  assign n26372 = n8867 ^ n5507 ^ 1'b0 ;
  assign n26373 = n26372 ^ n14352 ^ n184 ;
  assign n26374 = ( n3428 & n5915 ) | ( n3428 & ~n13321 ) | ( n5915 & ~n13321 ) ;
  assign n26375 = n540 & n12735 ;
  assign n26376 = n4294 ^ n3430 ^ 1'b0 ;
  assign n26377 = ~n4809 & n26376 ;
  assign n26378 = n12393 ^ n9049 ^ 1'b0 ;
  assign n26379 = n26377 & ~n26378 ;
  assign n26380 = n10908 & n11652 ;
  assign n26381 = n3783 ^ n1352 ^ 1'b0 ;
  assign n26382 = n10168 ^ n8734 ^ 1'b0 ;
  assign n26383 = ~n26381 & n26382 ;
  assign n26384 = ~n12812 & n26383 ;
  assign n26385 = n26380 | n26384 ;
  assign n26386 = n8523 & n10027 ;
  assign n26387 = n26386 ^ n22951 ^ 1'b0 ;
  assign n26388 = n7259 ^ n5795 ^ n2568 ;
  assign n26389 = ~n5984 & n21463 ;
  assign n26390 = n8407 ^ n1800 ^ 1'b0 ;
  assign n26391 = n26390 ^ n2695 ^ 1'b0 ;
  assign n26392 = n3011 & n20547 ;
  assign n26393 = n317 & ~n17874 ;
  assign n26394 = n26393 ^ n3979 ^ 1'b0 ;
  assign n26395 = ~n26393 & n26394 ;
  assign n26396 = ~n26392 & n26395 ;
  assign n26397 = n26396 ^ n6694 ^ 1'b0 ;
  assign n26398 = n2408 | n8312 ;
  assign n26399 = n7943 | n26398 ;
  assign n26400 = n26399 ^ n4650 ^ 1'b0 ;
  assign n26401 = n26377 & ~n26400 ;
  assign n26402 = n26401 ^ n7869 ^ 1'b0 ;
  assign n26403 = ~n694 & n26402 ;
  assign n26404 = n13732 ^ n423 ^ 1'b0 ;
  assign n26405 = n26404 ^ n14270 ^ n4737 ;
  assign n26406 = n18676 & n21042 ;
  assign n26407 = n26406 ^ n5801 ^ 1'b0 ;
  assign n26408 = ( ~n26403 & n26405 ) | ( ~n26403 & n26407 ) | ( n26405 & n26407 ) ;
  assign n26409 = ( n17022 & ~n17658 ) | ( n17022 & n25980 ) | ( ~n17658 & n25980 ) ;
  assign n26410 = n3609 | n24199 ;
  assign n26412 = n6498 & n9623 ;
  assign n26413 = n1689 & ~n26412 ;
  assign n26414 = n26413 ^ n716 ^ 1'b0 ;
  assign n26411 = n18209 | n22440 ;
  assign n26415 = n26414 ^ n26411 ^ 1'b0 ;
  assign n26417 = n4545 | n16233 ;
  assign n26416 = n11416 & n18420 ;
  assign n26418 = n26417 ^ n26416 ^ 1'b0 ;
  assign n26419 = n22574 ^ n5222 ^ n2484 ;
  assign n26420 = n26419 ^ n16502 ^ 1'b0 ;
  assign n26421 = ~n11876 & n23927 ;
  assign n26422 = ~n968 & n4224 ;
  assign n26423 = n7929 & ~n15431 ;
  assign n26424 = n26423 ^ n15766 ^ 1'b0 ;
  assign n26425 = n10237 & n26424 ;
  assign n26426 = ~n26422 & n26425 ;
  assign n26432 = n11691 ^ n108 ^ 1'b0 ;
  assign n26427 = n7900 ^ n815 ^ n500 ;
  assign n26428 = n26427 ^ n25419 ^ 1'b0 ;
  assign n26429 = n17598 ^ n9835 ^ 1'b0 ;
  assign n26430 = n18389 & ~n26429 ;
  assign n26431 = n26428 & n26430 ;
  assign n26433 = n26432 ^ n26431 ^ 1'b0 ;
  assign n26434 = n21652 ^ n19473 ^ 1'b0 ;
  assign n26439 = ( n2283 & n3409 ) | ( n2283 & ~n6590 ) | ( n3409 & ~n6590 ) ;
  assign n26440 = ~n2510 & n3731 ;
  assign n26441 = ~n1329 & n26440 ;
  assign n26442 = n26441 ^ n25170 ^ 1'b0 ;
  assign n26443 = ~n1590 & n26442 ;
  assign n26444 = n15781 & n26443 ;
  assign n26445 = n26444 ^ n22242 ^ 1'b0 ;
  assign n26446 = ~n26439 & n26445 ;
  assign n26447 = n26446 ^ n4528 ^ 1'b0 ;
  assign n26435 = n1648 & n2683 ;
  assign n26436 = n2004 & n26435 ;
  assign n26437 = n19820 & ~n26436 ;
  assign n26438 = n26437 ^ n9304 ^ 1'b0 ;
  assign n26448 = n26447 ^ n26438 ^ n22854 ;
  assign n26449 = n2794 & ~n5953 ;
  assign n26454 = n12165 ^ n5329 ^ 1'b0 ;
  assign n26450 = ~n2879 & n14282 ;
  assign n26451 = n26450 ^ n5458 ^ 1'b0 ;
  assign n26452 = n5058 & n26451 ;
  assign n26453 = ~n5578 & n26452 ;
  assign n26455 = n26454 ^ n26453 ^ 1'b0 ;
  assign n26456 = n11431 & ~n16910 ;
  assign n26457 = n4711 | n12511 ;
  assign n26458 = ~n4338 & n23444 ;
  assign n26459 = n26458 ^ n15937 ^ 1'b0 ;
  assign n26460 = n3004 | n10286 ;
  assign n26461 = n26460 ^ n7458 ^ 1'b0 ;
  assign n26462 = ~n7621 & n26461 ;
  assign n26463 = n26462 ^ n8505 ^ 1'b0 ;
  assign n26464 = n13495 | n17857 ;
  assign n26465 = n15386 & ~n26464 ;
  assign n26466 = ( n12781 & n26463 ) | ( n12781 & n26465 ) | ( n26463 & n26465 ) ;
  assign n26467 = n22094 ^ n6937 ^ 1'b0 ;
  assign n26468 = n10874 & ~n26467 ;
  assign n26469 = n22703 | n25117 ;
  assign n26470 = n22436 & n25974 ;
  assign n26471 = n26470 ^ n23505 ^ 1'b0 ;
  assign n26472 = n13270 ^ n12943 ^ n8001 ;
  assign n26473 = n26472 ^ n23244 ^ 1'b0 ;
  assign n26474 = n3638 ^ n2244 ^ 1'b0 ;
  assign n26475 = ~n1700 & n26474 ;
  assign n26476 = n8403 & n15672 ;
  assign n26477 = n10093 | n26476 ;
  assign n26478 = n2216 & ~n26477 ;
  assign n26479 = ~n1819 & n16725 ;
  assign n26480 = ~n11124 & n26479 ;
  assign n26481 = n18888 | n26480 ;
  assign n26482 = n26481 ^ n10364 ^ 1'b0 ;
  assign n26483 = n1768 & n26482 ;
  assign n26484 = n26483 ^ n669 ^ 1'b0 ;
  assign n26485 = n15653 ^ n12924 ^ 1'b0 ;
  assign n26486 = ~n5267 & n18307 ;
  assign n26487 = n17931 ^ n3042 ^ 1'b0 ;
  assign n26488 = n4540 ^ n3892 ^ 1'b0 ;
  assign n26489 = n21083 | n26488 ;
  assign n26490 = n6426 | n9899 ;
  assign n26491 = n24875 ^ n9239 ^ 1'b0 ;
  assign n26492 = ~n13500 & n26491 ;
  assign n26493 = n12602 & n14545 ;
  assign n26494 = ( n1563 & n6867 ) | ( n1563 & ~n26393 ) | ( n6867 & ~n26393 ) ;
  assign n26495 = n6944 ^ n1525 ^ 1'b0 ;
  assign n26496 = ~n9984 & n26495 ;
  assign n26497 = n10259 & ~n12045 ;
  assign n26498 = n13413 & n26497 ;
  assign n26499 = n9670 ^ n8443 ^ 1'b0 ;
  assign n26500 = n8823 & ~n26499 ;
  assign n26501 = n26500 ^ n9525 ^ 1'b0 ;
  assign n26502 = n11283 & ~n26501 ;
  assign n26503 = n10761 & n24173 ;
  assign n26504 = n26503 ^ n5933 ^ 1'b0 ;
  assign n26505 = n10284 ^ n4712 ^ 1'b0 ;
  assign n26506 = n6922 | n13566 ;
  assign n26507 = n1809 & n13345 ;
  assign n26508 = n2134 & n26507 ;
  assign n26509 = n4799 & ~n18220 ;
  assign n26510 = n11182 & n26509 ;
  assign n26511 = n11423 ^ n10117 ^ 1'b0 ;
  assign n26512 = n12157 & ~n26511 ;
  assign n26513 = ( n4624 & n26510 ) | ( n4624 & ~n26512 ) | ( n26510 & ~n26512 ) ;
  assign n26514 = ( n25752 & n26508 ) | ( n25752 & ~n26513 ) | ( n26508 & ~n26513 ) ;
  assign n26515 = n1484 & n2085 ;
  assign n26516 = n26515 ^ n3211 ^ 1'b0 ;
  assign n26517 = n16391 ^ n5181 ^ 1'b0 ;
  assign n26518 = n10948 | n26517 ;
  assign n26519 = n8208 & n26518 ;
  assign n26520 = n22741 ^ n6534 ^ 1'b0 ;
  assign n26521 = n26520 ^ n6947 ^ 1'b0 ;
  assign n26522 = n7067 & ~n26521 ;
  assign n26523 = n10029 ^ n690 ^ 1'b0 ;
  assign n26524 = n26523 ^ n18244 ^ 1'b0 ;
  assign n26525 = n22217 ^ n14545 ^ 1'b0 ;
  assign n26526 = n11033 ^ n6885 ^ 1'b0 ;
  assign n26527 = n208 & ~n26526 ;
  assign n26528 = n11286 | n20510 ;
  assign n26529 = n26528 ^ n17156 ^ 1'b0 ;
  assign n26530 = ~n3521 & n19478 ;
  assign n26531 = n26530 ^ n2785 ^ 1'b0 ;
  assign n26532 = n8305 ^ n3611 ^ 1'b0 ;
  assign n26533 = n5443 ^ n827 ^ 1'b0 ;
  assign n26534 = n26533 ^ n3487 ^ 1'b0 ;
  assign n26535 = ( n16702 & n26532 ) | ( n16702 & ~n26534 ) | ( n26532 & ~n26534 ) ;
  assign n26536 = n2918 & ~n26535 ;
  assign n26537 = n26536 ^ n1574 ^ 1'b0 ;
  assign n26538 = n8942 ^ n8132 ^ 1'b0 ;
  assign n26539 = ~n1456 & n26538 ;
  assign n26540 = ~n22257 & n26539 ;
  assign n26541 = n4750 & n26540 ;
  assign n26543 = ( n2535 & n7254 ) | ( n2535 & ~n11977 ) | ( n7254 & ~n11977 ) ;
  assign n26542 = ( n592 & ~n4768 ) | ( n592 & n16640 ) | ( ~n4768 & n16640 ) ;
  assign n26544 = n26543 ^ n26542 ^ 1'b0 ;
  assign n26545 = ~n24256 & n26544 ;
  assign n26546 = n22501 ^ n11932 ^ n2572 ;
  assign n26548 = n3186 & ~n12317 ;
  assign n26547 = n4583 | n22231 ;
  assign n26549 = n26548 ^ n26547 ^ 1'b0 ;
  assign n26550 = n26549 ^ n13033 ^ 1'b0 ;
  assign n26551 = n7785 ^ n4865 ^ 1'b0 ;
  assign n26552 = n2150 & n26551 ;
  assign n26553 = n10073 ^ n513 ^ 1'b0 ;
  assign n26554 = n26552 & ~n26553 ;
  assign n26555 = n2501 & n26554 ;
  assign n26556 = n6762 | n26555 ;
  assign n26557 = n2593 & ~n12579 ;
  assign n26558 = n17294 ^ n3660 ^ 1'b0 ;
  assign n26559 = n26557 & n26558 ;
  assign n26560 = n14039 ^ n9141 ^ 1'b0 ;
  assign n26561 = ~n15363 & n26560 ;
  assign n26562 = ~n6054 & n26561 ;
  assign n26563 = n1327 & ~n7123 ;
  assign n26564 = ( n2468 & ~n2671 ) | ( n2468 & n26563 ) | ( ~n2671 & n26563 ) ;
  assign n26565 = n8486 ^ n6528 ^ 1'b0 ;
  assign n26566 = ( n1958 & n22782 ) | ( n1958 & n26565 ) | ( n22782 & n26565 ) ;
  assign n26569 = n23584 & ~n26104 ;
  assign n26570 = n26569 ^ n17285 ^ 1'b0 ;
  assign n26571 = n6140 & ~n26570 ;
  assign n26567 = n7427 & n13021 ;
  assign n26568 = n13747 | n26567 ;
  assign n26572 = n26571 ^ n26568 ^ 1'b0 ;
  assign n26573 = n21293 ^ n14401 ^ 1'b0 ;
  assign n26574 = n821 & ~n26573 ;
  assign n26575 = n130 & n13690 ;
  assign n26576 = n302 | n1967 ;
  assign n26577 = n26576 ^ n9233 ^ 1'b0 ;
  assign n26578 = n9975 & n26577 ;
  assign n26579 = ~n11863 & n26578 ;
  assign n26582 = n1194 ^ n1010 ^ 1'b0 ;
  assign n26580 = n13694 & ~n15459 ;
  assign n26581 = n26580 ^ n1674 ^ 1'b0 ;
  assign n26583 = n26582 ^ n26581 ^ 1'b0 ;
  assign n26584 = ~n26579 & n26583 ;
  assign n26585 = n10287 & n11673 ;
  assign n26586 = n20046 ^ n2453 ^ 1'b0 ;
  assign n26587 = n8156 | n11295 ;
  assign n26588 = n20489 ^ n10861 ^ n6254 ;
  assign n26589 = n8534 ^ n3477 ^ n2994 ;
  assign n26591 = n2960 & ~n3129 ;
  assign n26592 = n26591 ^ n6174 ^ 1'b0 ;
  assign n26590 = n4170 & n16399 ;
  assign n26593 = n26592 ^ n26590 ^ n12678 ;
  assign n26594 = n15783 ^ n9528 ^ 1'b0 ;
  assign n26595 = n23883 & ~n26594 ;
  assign n26596 = ~n18465 & n26595 ;
  assign n26597 = n26596 ^ n15016 ^ 1'b0 ;
  assign n26598 = ~n7697 & n22705 ;
  assign n26599 = n7917 & ~n10624 ;
  assign n26600 = n8845 & ~n15365 ;
  assign n26601 = n996 & n21765 ;
  assign n26602 = n26601 ^ n4679 ^ 1'b0 ;
  assign n26603 = n5805 & n9940 ;
  assign n26604 = ~n9768 & n12039 ;
  assign n26605 = n26604 ^ n133 ^ 1'b0 ;
  assign n26606 = n26603 | n26605 ;
  assign n26607 = n17214 ^ x6 ^ 1'b0 ;
  assign n26608 = ~n11312 & n18033 ;
  assign n26609 = ~n25003 & n26608 ;
  assign n26610 = n26609 ^ n988 ^ 1'b0 ;
  assign n26611 = n21466 ^ n627 ^ 1'b0 ;
  assign n26612 = n23427 & ~n26611 ;
  assign n26613 = n9084 ^ n2474 ^ 1'b0 ;
  assign n26614 = n15614 & ~n26613 ;
  assign n26615 = n1237 & ~n26614 ;
  assign n26616 = ~n3527 & n26615 ;
  assign n26617 = n24015 & n25189 ;
  assign n26618 = n26617 ^ n22024 ^ 1'b0 ;
  assign n26619 = n16810 & n21313 ;
  assign n26620 = n3638 & n5613 ;
  assign n26621 = n6389 & ~n14578 ;
  assign n26622 = n13896 ^ n7958 ^ 1'b0 ;
  assign n26623 = n20607 & ~n26622 ;
  assign n26624 = n26623 ^ n2922 ^ n1887 ;
  assign n26625 = n7398 ^ n2460 ^ 1'b0 ;
  assign n26626 = n10795 ^ n5890 ^ 1'b0 ;
  assign n26627 = ~n1353 & n26626 ;
  assign n26628 = n23962 ^ n10872 ^ 1'b0 ;
  assign n26629 = n20920 ^ n3480 ^ 1'b0 ;
  assign n26630 = n26628 | n26629 ;
  assign n26631 = n984 | n2529 ;
  assign n26632 = n26631 ^ n124 ^ 1'b0 ;
  assign n26637 = n1184 & n1800 ;
  assign n26638 = ~n1752 & n26637 ;
  assign n26633 = n3802 & ~n15487 ;
  assign n26634 = n26633 ^ n20302 ^ 1'b0 ;
  assign n26635 = n26634 ^ n13732 ^ 1'b0 ;
  assign n26636 = n3375 | n26635 ;
  assign n26639 = n26638 ^ n26636 ^ 1'b0 ;
  assign n26640 = n6235 | n24447 ;
  assign n26641 = n17869 & ~n26640 ;
  assign n26642 = ~n459 & n4525 ;
  assign n26643 = n26642 ^ n17084 ^ 1'b0 ;
  assign n26644 = ~n19972 & n26643 ;
  assign n26646 = ~n5107 & n5139 ;
  assign n26647 = n26646 ^ n5632 ^ 1'b0 ;
  assign n26645 = n3194 & n21371 ;
  assign n26648 = n26647 ^ n26645 ^ 1'b0 ;
  assign n26649 = n2338 & n2567 ;
  assign n26650 = n26649 ^ n2346 ^ 1'b0 ;
  assign n26651 = n26648 & ~n26650 ;
  assign n26652 = n4440 ^ n3308 ^ 1'b0 ;
  assign n26653 = n15741 & ~n26652 ;
  assign n26655 = n16175 ^ n8735 ^ 1'b0 ;
  assign n26656 = n7285 & ~n26655 ;
  assign n26654 = n560 | n5985 ;
  assign n26657 = n26656 ^ n26654 ^ 1'b0 ;
  assign n26658 = n3619 & n5052 ;
  assign n26659 = n19053 & ~n26658 ;
  assign n26660 = n26659 ^ n9296 ^ 1'b0 ;
  assign n26661 = n10888 | n22425 ;
  assign n26662 = n26661 ^ n3706 ^ 1'b0 ;
  assign n26663 = ( n2146 & n13357 ) | ( n2146 & ~n18069 ) | ( n13357 & ~n18069 ) ;
  assign n26664 = n26663 ^ n19367 ^ 1'b0 ;
  assign n26665 = ~n2560 & n9863 ;
  assign n26666 = n2042 | n16319 ;
  assign n26667 = n26665 & ~n26666 ;
  assign n26668 = ~n727 & n26667 ;
  assign n26669 = n7502 ^ n7137 ^ n6069 ;
  assign n26670 = n26669 ^ n7080 ^ 1'b0 ;
  assign n26671 = n5489 ^ n4714 ^ n3266 ;
  assign n26672 = n2671 & n14223 ;
  assign n26673 = n26671 & ~n26672 ;
  assign n26674 = n12823 | n21271 ;
  assign n26675 = ~n13911 & n26674 ;
  assign n26676 = ~n18960 & n26675 ;
  assign n26677 = n5592 & ~n15596 ;
  assign n26678 = n24334 ^ n12285 ^ 1'b0 ;
  assign n26679 = n8212 ^ n5957 ^ 1'b0 ;
  assign n26680 = n2554 ^ n493 ^ 1'b0 ;
  assign n26681 = n2324 & n10997 ;
  assign n26682 = ~n26680 & n26681 ;
  assign n26683 = n6995 & n10426 ;
  assign n26684 = n26682 & n26683 ;
  assign n26685 = n8281 ^ n2869 ^ 1'b0 ;
  assign n26686 = n12549 & ~n26685 ;
  assign n26687 = n6018 & ~n12340 ;
  assign n26688 = ~n16275 & n26687 ;
  assign n26689 = n10959 ^ n8599 ^ 1'b0 ;
  assign n26690 = n13498 | n26689 ;
  assign n26691 = n21261 | n26690 ;
  assign n26692 = n24814 | n26691 ;
  assign n26693 = n26692 ^ n615 ^ 1'b0 ;
  assign n26694 = n6868 & n12921 ;
  assign n26695 = n1308 & n26694 ;
  assign n26696 = n10511 ^ n7193 ^ 1'b0 ;
  assign n26697 = n10751 & n26696 ;
  assign n26698 = n26697 ^ n12119 ^ 1'b0 ;
  assign n26699 = x1 | n5311 ;
  assign n26700 = n2114 | n26699 ;
  assign n26701 = n9205 & ~n14304 ;
  assign n26702 = n26701 ^ n6254 ^ 1'b0 ;
  assign n26703 = n26700 | n26702 ;
  assign n26704 = n26703 ^ n7717 ^ 1'b0 ;
  assign n26705 = n4229 | n4789 ;
  assign n26706 = n26705 ^ n4340 ^ 1'b0 ;
  assign n26707 = n23643 | n26706 ;
  assign n26708 = n9459 ^ n1613 ^ 1'b0 ;
  assign n26709 = n26707 & n26708 ;
  assign n26710 = n6817 ^ n1734 ^ 1'b0 ;
  assign n26711 = n26710 ^ n4916 ^ n43 ;
  assign n26712 = n26709 | n26711 ;
  assign n26715 = n8500 & ~n9693 ;
  assign n26713 = n2917 ^ n124 ^ 1'b0 ;
  assign n26714 = n2101 & ~n26713 ;
  assign n26716 = n26715 ^ n26714 ^ n7119 ;
  assign n26718 = n19897 ^ n8287 ^ 1'b0 ;
  assign n26719 = n9717 & ~n26718 ;
  assign n26717 = ~n2217 & n17745 ;
  assign n26720 = n26719 ^ n26717 ^ 1'b0 ;
  assign n26721 = n10701 ^ n4068 ^ 1'b0 ;
  assign n26722 = n22593 & ~n26721 ;
  assign n26723 = n2812 ^ n1196 ^ 1'b0 ;
  assign n26724 = n21052 & ~n24487 ;
  assign n26725 = n20289 & n24329 ;
  assign n26726 = n13855 ^ n12589 ^ 1'b0 ;
  assign n26727 = n10298 & n26726 ;
  assign n26728 = n676 & n26727 ;
  assign n26729 = ~n6878 & n26728 ;
  assign n26730 = n503 | n4807 ;
  assign n26731 = ~n26729 & n26730 ;
  assign n26732 = n21935 ^ n4438 ^ 1'b0 ;
  assign n26733 = n412 & ~n19918 ;
  assign n26734 = n26733 ^ n9090 ^ 1'b0 ;
  assign n26735 = n22939 ^ n16926 ^ 1'b0 ;
  assign n26736 = ~n26734 & n26735 ;
  assign n26737 = n26736 ^ n1987 ^ 1'b0 ;
  assign n26738 = n5699 | n21474 ;
  assign n26739 = n15571 ^ n7398 ^ 1'b0 ;
  assign n26740 = n6093 | n18409 ;
  assign n26744 = n18797 ^ n11909 ^ 1'b0 ;
  assign n26741 = n6128 & ~n12583 ;
  assign n26742 = n26741 ^ n2549 ^ 1'b0 ;
  assign n26743 = n26742 ^ n20346 ^ 1'b0 ;
  assign n26745 = n26744 ^ n26743 ^ 1'b0 ;
  assign n26746 = n4070 & n11295 ;
  assign n26747 = n4644 | n7272 ;
  assign n26748 = n26747 ^ n18310 ^ n16002 ;
  assign n26749 = n26748 ^ n12716 ^ 1'b0 ;
  assign n26750 = ~n2214 & n26749 ;
  assign n26751 = n4644 ^ n2610 ^ 1'b0 ;
  assign n26752 = n8659 & n9661 ;
  assign n26753 = n16582 ^ n3751 ^ 1'b0 ;
  assign n26754 = n7788 & ~n26753 ;
  assign n26755 = n1099 ^ n740 ^ 1'b0 ;
  assign n26756 = n164 & ~n26755 ;
  assign n26757 = n2555 | n7529 ;
  assign n26758 = n26756 | n26757 ;
  assign n26759 = n9500 ^ n5727 ^ 1'b0 ;
  assign n26760 = n26758 & ~n26759 ;
  assign n26761 = n1843 & n9851 ;
  assign n26762 = n25296 ^ n20787 ^ 1'b0 ;
  assign n26763 = n26498 & n26762 ;
  assign n26767 = n10153 ^ n6742 ^ 1'b0 ;
  assign n26766 = n2370 ^ n725 ^ 1'b0 ;
  assign n26764 = n19808 ^ n17085 ^ 1'b0 ;
  assign n26765 = ~n6463 & n26764 ;
  assign n26768 = n26767 ^ n26766 ^ n26765 ;
  assign n26769 = n8107 ^ n7713 ^ 1'b0 ;
  assign n26770 = n26769 ^ n16495 ^ 1'b0 ;
  assign n26771 = n1772 & ~n8987 ;
  assign n26772 = n26771 ^ n3896 ^ 1'b0 ;
  assign n26773 = n26770 & n26772 ;
  assign n26774 = n1802 | n13876 ;
  assign n26775 = n12821 & ~n25122 ;
  assign n26776 = n2337 ^ n20 ^ 1'b0 ;
  assign n26777 = n237 & n26776 ;
  assign n26778 = n3174 & ~n26777 ;
  assign n26779 = n20392 ^ n9190 ^ n2317 ;
  assign n26780 = n15292 ^ n10978 ^ 1'b0 ;
  assign n26781 = ~n6744 & n26780 ;
  assign n26782 = n26781 ^ n4741 ^ 1'b0 ;
  assign n26783 = n7839 | n14505 ;
  assign n26784 = ( n772 & n1623 ) | ( n772 & n14975 ) | ( n1623 & n14975 ) ;
  assign n26785 = n8292 | n26784 ;
  assign n26786 = n26783 & ~n26785 ;
  assign n26787 = n26786 ^ n7482 ^ 1'b0 ;
  assign n26788 = n7199 & ~n26787 ;
  assign n26789 = n26788 ^ n4589 ^ 1'b0 ;
  assign n26790 = n25033 ^ n3279 ^ 1'b0 ;
  assign n26791 = n3724 | n9611 ;
  assign n26792 = n12426 & ~n26791 ;
  assign n26793 = n15127 | n22936 ;
  assign n26794 = n5139 & ~n26793 ;
  assign n26795 = n23886 & ~n26794 ;
  assign n26796 = n26795 ^ n1337 ^ 1'b0 ;
  assign n26797 = n26796 ^ n23011 ^ 1'b0 ;
  assign n26798 = ~n13085 & n26797 ;
  assign n26799 = n23331 ^ n331 ^ 1'b0 ;
  assign n26800 = ~n1943 & n26799 ;
  assign n26801 = n26800 ^ n19195 ^ 1'b0 ;
  assign n26802 = n8098 ^ n47 ^ 1'b0 ;
  assign n26803 = n6492 | n26802 ;
  assign n26804 = ~n7506 & n7989 ;
  assign n26805 = ~n22942 & n26804 ;
  assign n26806 = ~n317 & n26805 ;
  assign n26807 = n16057 & n26806 ;
  assign n26808 = n13041 ^ n5742 ^ 1'b0 ;
  assign n26809 = ~n3042 & n5136 ;
  assign n26810 = n26809 ^ n2108 ^ 1'b0 ;
  assign n26811 = n11423 & ~n26810 ;
  assign n26812 = ~n26808 & n26811 ;
  assign n26813 = n20007 ^ n12941 ^ 1'b0 ;
  assign n26814 = ~n26812 & n26813 ;
  assign n26815 = n2574 & n6274 ;
  assign n26816 = ~n6274 & n26815 ;
  assign n26817 = ~n3566 & n26816 ;
  assign n26818 = n3566 & n26817 ;
  assign n26819 = n11210 & ~n26818 ;
  assign n26820 = n26819 ^ n17409 ^ 1'b0 ;
  assign n26821 = n14354 ^ n1337 ^ 1'b0 ;
  assign n26822 = n4081 & ~n18209 ;
  assign n26823 = n23432 ^ n6444 ^ 1'b0 ;
  assign n26824 = ~n25897 & n26823 ;
  assign n26825 = ( ~n1187 & n15622 ) | ( ~n1187 & n19702 ) | ( n15622 & n19702 ) ;
  assign n26826 = n11668 ^ n4327 ^ 1'b0 ;
  assign n26827 = ~n6399 & n23318 ;
  assign n26828 = n26827 ^ n1213 ^ 1'b0 ;
  assign n26829 = n910 | n26828 ;
  assign n26830 = ~n3924 & n7397 ;
  assign n26831 = n4016 ^ n940 ^ 1'b0 ;
  assign n26832 = n26831 ^ n22046 ^ n9269 ;
  assign n26833 = ~n654 & n26832 ;
  assign n26834 = n18295 & ~n26833 ;
  assign n26835 = n16443 ^ n6981 ^ n4884 ;
  assign n26836 = n14413 | n21048 ;
  assign n26837 = ~n4496 & n25428 ;
  assign n26838 = n26837 ^ n10973 ^ 1'b0 ;
  assign n26839 = n26838 ^ n14828 ^ 1'b0 ;
  assign n26840 = ~n13490 & n22974 ;
  assign n26841 = n12576 & n26840 ;
  assign n26842 = n26841 ^ n13671 ^ 1'b0 ;
  assign n26843 = n26842 ^ n24926 ^ n23281 ;
  assign n26844 = n26843 ^ n8539 ^ 1'b0 ;
  assign n26845 = ~n7846 & n13314 ;
  assign n26846 = n3858 & n26845 ;
  assign n26847 = n3502 & ~n7835 ;
  assign n26848 = n10168 & n26847 ;
  assign n26849 = n16788 ^ n7112 ^ n6318 ;
  assign n26850 = ~n16727 & n26849 ;
  assign n26851 = ~n9232 & n26850 ;
  assign n26852 = n10405 | n15867 ;
  assign n26853 = ( n948 & ~n9198 ) | ( n948 & n9965 ) | ( ~n9198 & n9965 ) ;
  assign n26854 = ( n9360 & n26852 ) | ( n9360 & ~n26853 ) | ( n26852 & ~n26853 ) ;
  assign n26855 = n8254 ^ n4228 ^ 1'b0 ;
  assign n26856 = n9546 & n26855 ;
  assign n26857 = n17583 & n26856 ;
  assign n26858 = n26857 ^ n4461 ^ 1'b0 ;
  assign n26861 = n17362 ^ n7346 ^ 1'b0 ;
  assign n26862 = ~n2612 & n26861 ;
  assign n26859 = n12550 ^ n8704 ^ 1'b0 ;
  assign n26860 = n18721 & n26859 ;
  assign n26863 = n26862 ^ n26860 ^ 1'b0 ;
  assign n26864 = n1810 & ~n23523 ;
  assign n26865 = ~n1810 & n26864 ;
  assign n26870 = n2445 & n21245 ;
  assign n26871 = n26870 ^ n5420 ^ 1'b0 ;
  assign n26872 = n19051 & n26871 ;
  assign n26873 = n26872 ^ n9191 ^ 1'b0 ;
  assign n26866 = n1830 | n11711 ;
  assign n26867 = n7749 & ~n26866 ;
  assign n26868 = n26867 ^ n1157 ^ 1'b0 ;
  assign n26869 = n874 | n26868 ;
  assign n26874 = n26873 ^ n26869 ^ 1'b0 ;
  assign n26875 = n9254 ^ n1839 ^ 1'b0 ;
  assign n26876 = n11689 & ~n20257 ;
  assign n26877 = ~n800 & n5289 ;
  assign n26878 = n26877 ^ n23108 ^ n9401 ;
  assign n26879 = ~n5416 & n11849 ;
  assign n26880 = n13761 ^ n5477 ^ 1'b0 ;
  assign n26881 = ~n2640 & n26880 ;
  assign n26882 = n4827 & ~n12052 ;
  assign n26883 = n477 & ~n11688 ;
  assign n26884 = n26883 ^ n15842 ^ 1'b0 ;
  assign n26885 = n26884 ^ n12115 ^ 1'b0 ;
  assign n26887 = n4276 | n12501 ;
  assign n26888 = n26887 ^ n6766 ^ 1'b0 ;
  assign n26886 = n8515 & ~n12467 ;
  assign n26889 = n26888 ^ n26886 ^ 1'b0 ;
  assign n26890 = n12993 ^ n11427 ^ 1'b0 ;
  assign n26891 = n14639 & ~n15368 ;
  assign n26892 = n26891 ^ n14302 ^ 1'b0 ;
  assign n26893 = n12002 ^ n5765 ^ n3314 ;
  assign n26894 = n9024 & ~n26893 ;
  assign n26895 = n26894 ^ n2494 ^ 1'b0 ;
  assign n26896 = n11088 & n21245 ;
  assign n26897 = n26896 ^ n23087 ^ 1'b0 ;
  assign n26898 = n26897 ^ n6560 ^ n4616 ;
  assign n26899 = ~n8731 & n13119 ;
  assign n26900 = n2906 | n26566 ;
  assign n26901 = n26900 ^ n17833 ^ 1'b0 ;
  assign n26902 = ( ~n6635 & n7695 ) | ( ~n6635 & n10245 ) | ( n7695 & n10245 ) ;
  assign n26904 = n5558 | n15232 ;
  assign n26903 = n3083 | n7368 ;
  assign n26905 = n26904 ^ n26903 ^ 1'b0 ;
  assign n26906 = ( n9380 & n10740 ) | ( n9380 & n11274 ) | ( n10740 & n11274 ) ;
  assign n26907 = n7245 & n26906 ;
  assign n26908 = n3695 ^ n420 ^ 1'b0 ;
  assign n26909 = n10565 & n26908 ;
  assign n26910 = n12501 & n26909 ;
  assign n26911 = n22703 ^ n1269 ^ 1'b0 ;
  assign n26912 = n9714 & n26911 ;
  assign n26913 = n13130 ^ n6081 ^ n1961 ;
  assign n26914 = n19067 & n26913 ;
  assign n26915 = n26914 ^ n14983 ^ 1'b0 ;
  assign n26916 = n25955 ^ n12561 ^ 1'b0 ;
  assign n26917 = n14177 | n26916 ;
  assign n26918 = n14406 ^ n12133 ^ 1'b0 ;
  assign n26919 = n26918 ^ n24063 ^ n18742 ;
  assign n26920 = ~n3122 & n20469 ;
  assign n26921 = n26920 ^ n1853 ^ 1'b0 ;
  assign n26922 = n26921 ^ n24342 ^ 1'b0 ;
  assign n26923 = n7628 & ~n22740 ;
  assign n26924 = n292 | n19074 ;
  assign n26925 = n2539 & n14750 ;
  assign n26926 = n26925 ^ n4434 ^ 1'b0 ;
  assign n26927 = n26926 ^ n17927 ^ 1'b0 ;
  assign n26928 = ( n950 & ~n13809 ) | ( n950 & n23534 ) | ( ~n13809 & n23534 ) ;
  assign n26929 = n16028 ^ n8357 ^ 1'b0 ;
  assign n26930 = n26928 & ~n26929 ;
  assign n26931 = ~n18425 & n26201 ;
  assign n26933 = n8830 ^ n5130 ^ 1'b0 ;
  assign n26934 = n6740 & ~n26933 ;
  assign n26932 = ~n14385 & n20475 ;
  assign n26935 = n26934 ^ n26932 ^ 1'b0 ;
  assign n26936 = n11334 ^ n150 ^ 1'b0 ;
  assign n26937 = n15782 ^ n1786 ^ 1'b0 ;
  assign n26938 = n26936 | n26937 ;
  assign n26945 = n3901 ^ n2824 ^ 1'b0 ;
  assign n26940 = n1310 & n5308 ;
  assign n26939 = ~n6269 & n21402 ;
  assign n26941 = n26940 ^ n26939 ^ 1'b0 ;
  assign n26942 = n13240 ^ n8679 ^ 1'b0 ;
  assign n26943 = n19854 & n26942 ;
  assign n26944 = n26941 & n26943 ;
  assign n26946 = n26945 ^ n26944 ^ 1'b0 ;
  assign n26947 = ~n7964 & n17792 ;
  assign n26948 = n9851 & n26947 ;
  assign n26949 = n1932 | n26296 ;
  assign n26950 = n20829 ^ n1469 ^ 1'b0 ;
  assign n26951 = ~n21326 & n26950 ;
  assign n26952 = n1095 & ~n22683 ;
  assign n26957 = n61 & n2871 ;
  assign n26958 = n26957 ^ n2272 ^ 1'b0 ;
  assign n26953 = n9620 ^ n5675 ^ 1'b0 ;
  assign n26954 = ~n2728 & n26953 ;
  assign n26955 = ~n25377 & n26954 ;
  assign n26956 = n26955 ^ n4206 ^ 1'b0 ;
  assign n26959 = n26958 ^ n26956 ^ n6351 ;
  assign n26960 = n2996 | n4451 ;
  assign n26961 = n4632 ^ n2038 ^ 1'b0 ;
  assign n26962 = n26961 ^ n1699 ^ 1'b0 ;
  assign n26963 = n3547 ^ n1004 ^ 1'b0 ;
  assign n26964 = n10542 | n26963 ;
  assign n26965 = n26961 | n26964 ;
  assign n26966 = n7681 ^ n3017 ^ 1'b0 ;
  assign n26967 = ~n18096 & n26966 ;
  assign n26968 = n891 | n6825 ;
  assign n26969 = n26967 & ~n26968 ;
  assign n26970 = n26565 ^ n3027 ^ 1'b0 ;
  assign n26971 = ~n515 & n26970 ;
  assign n26972 = n26971 ^ n2873 ^ 1'b0 ;
  assign n26973 = n7112 ^ n4609 ^ n2796 ;
  assign n26974 = n26973 ^ n24271 ^ 1'b0 ;
  assign n26975 = n14804 & ~n22093 ;
  assign n26976 = ~n7757 & n9777 ;
  assign n26977 = n4965 & n26976 ;
  assign n26978 = ( ~n1929 & n4235 ) | ( ~n1929 & n8562 ) | ( n4235 & n8562 ) ;
  assign n26979 = n17560 | n26978 ;
  assign n26980 = n26977 & ~n26979 ;
  assign n26985 = n17829 ^ n267 ^ 1'b0 ;
  assign n26981 = n3564 & n5847 ;
  assign n26982 = ~n1525 & n26981 ;
  assign n26983 = n1190 & n1573 ;
  assign n26984 = ~n26982 & n26983 ;
  assign n26986 = n26985 ^ n26984 ^ 1'b0 ;
  assign n26987 = n15094 ^ n3558 ^ 1'b0 ;
  assign n26988 = ~n788 & n23048 ;
  assign n26989 = n10144 ^ n4284 ^ 1'b0 ;
  assign n26990 = n311 | n2356 ;
  assign n26991 = n26990 ^ n24861 ^ 1'b0 ;
  assign n26992 = n26991 ^ n12559 ^ 1'b0 ;
  assign n26993 = n8993 | n12659 ;
  assign n26994 = ~n20860 & n26993 ;
  assign n26995 = n26994 ^ n21555 ^ 1'b0 ;
  assign n26996 = n11358 ^ n2780 ^ 1'b0 ;
  assign n26997 = ~n8792 & n26996 ;
  assign n26998 = n11860 & ~n21309 ;
  assign n26999 = ~n6775 & n26998 ;
  assign n27000 = n26997 | n26999 ;
  assign n27001 = n6681 & n7385 ;
  assign n27002 = n18925 | n27001 ;
  assign n27003 = n9935 & n15748 ;
  assign n27004 = n1257 | n27003 ;
  assign n27005 = n11737 ^ n344 ^ 1'b0 ;
  assign n27006 = ~n1522 & n14624 ;
  assign n27007 = ~n17099 & n27006 ;
  assign n27008 = n19780 ^ n5451 ^ 1'b0 ;
  assign n27009 = ~n27007 & n27008 ;
  assign n27010 = n16501 ^ n582 ^ 1'b0 ;
  assign n27011 = n27009 & n27010 ;
  assign n27012 = n14999 ^ n12513 ^ 1'b0 ;
  assign n27013 = ~n23630 & n27012 ;
  assign n27014 = ~n1438 & n18685 ;
  assign n27015 = n27014 ^ n2206 ^ 1'b0 ;
  assign n27016 = n2912 ^ n1691 ^ 1'b0 ;
  assign n27017 = n27016 ^ n17257 ^ 1'b0 ;
  assign n27018 = n6949 & ~n15925 ;
  assign n27019 = ( n183 & n4016 ) | ( n183 & n10790 ) | ( n4016 & n10790 ) ;
  assign n27020 = n7061 & ~n8334 ;
  assign n27021 = n27019 | n27020 ;
  assign n27022 = ~n12649 & n18383 ;
  assign n27023 = n27022 ^ n15462 ^ 1'b0 ;
  assign n27024 = n13218 & ~n27023 ;
  assign n27025 = n27024 ^ n2853 ^ 1'b0 ;
  assign n27026 = ( n5401 & n12516 ) | ( n5401 & n19365 ) | ( n12516 & n19365 ) ;
  assign n27027 = n4526 | n11162 ;
  assign n27029 = ~n8506 & n9116 ;
  assign n27030 = ~n11920 & n27029 ;
  assign n27031 = n20296 & n27030 ;
  assign n27028 = n1429 ^ n1012 ^ 1'b0 ;
  assign n27032 = n27031 ^ n27028 ^ 1'b0 ;
  assign n27033 = n7145 ^ n5138 ^ 1'b0 ;
  assign n27034 = n27033 ^ n10294 ^ 1'b0 ;
  assign n27035 = n11721 | n12839 ;
  assign n27038 = n7171 & ~n8975 ;
  assign n27037 = n3218 & ~n8322 ;
  assign n27039 = n27038 ^ n27037 ^ 1'b0 ;
  assign n27036 = n521 & ~n24006 ;
  assign n27040 = n27039 ^ n27036 ^ 1'b0 ;
  assign n27041 = n9432 & ~n15287 ;
  assign n27042 = n11253 & n27041 ;
  assign n27043 = n1907 & n27042 ;
  assign n27044 = n27043 ^ n11909 ^ 1'b0 ;
  assign n27045 = n12275 & n27044 ;
  assign n27046 = n2907 & n3766 ;
  assign n27047 = n23948 ^ n5117 ^ 1'b0 ;
  assign n27048 = n27046 & n27047 ;
  assign n27049 = n3202 & ~n4621 ;
  assign n27050 = n27049 ^ n9063 ^ 1'b0 ;
  assign n27051 = n27050 ^ n3327 ^ 1'b0 ;
  assign n27053 = n6458 & ~n12541 ;
  assign n27054 = n27053 ^ n6100 ^ 1'b0 ;
  assign n27052 = n4707 | n12417 ;
  assign n27055 = n27054 ^ n27052 ^ 1'b0 ;
  assign n27056 = n13589 & n26100 ;
  assign n27057 = n22496 ^ n12713 ^ 1'b0 ;
  assign n27058 = n13126 & n27057 ;
  assign n27060 = n5570 ^ n1504 ^ 1'b0 ;
  assign n27059 = n8081 | n12637 ;
  assign n27061 = n27060 ^ n27059 ^ 1'b0 ;
  assign n27062 = n19770 & n27061 ;
  assign n27063 = n13550 ^ n10839 ^ 1'b0 ;
  assign n27064 = n17723 ^ n105 ^ 1'b0 ;
  assign n27065 = n8130 & ~n27064 ;
  assign n27067 = n9060 | n26201 ;
  assign n27066 = n725 | n16923 ;
  assign n27068 = n27067 ^ n27066 ^ 1'b0 ;
  assign n27069 = ~n503 & n2614 ;
  assign n27070 = n7604 & ~n27069 ;
  assign n27071 = n27070 ^ x7 ^ 1'b0 ;
  assign n27072 = n6025 & n27071 ;
  assign n27073 = n5576 & n5662 ;
  assign n27074 = ~n19207 & n27073 ;
  assign n27076 = ~n802 & n2917 ;
  assign n27075 = n14845 ^ n12105 ^ 1'b0 ;
  assign n27077 = n27076 ^ n27075 ^ n4024 ;
  assign n27078 = ~n3813 & n12046 ;
  assign n27079 = n3437 ^ n2441 ^ 1'b0 ;
  assign n27080 = n4205 | n27079 ;
  assign n27081 = n27080 ^ n5167 ^ 1'b0 ;
  assign n27082 = n13520 & ~n27081 ;
  assign n27083 = ( n12145 & n14997 ) | ( n12145 & ~n27082 ) | ( n14997 & ~n27082 ) ;
  assign n27084 = ( n774 & n9955 ) | ( n774 & ~n14728 ) | ( n9955 & ~n14728 ) ;
  assign n27085 = ~n481 & n27084 ;
  assign n27086 = n1933 & n18961 ;
  assign n27087 = n27086 ^ n7609 ^ 1'b0 ;
  assign n27088 = n16747 ^ n4738 ^ 1'b0 ;
  assign n27089 = ~n17183 & n27088 ;
  assign n27090 = n1267 & n27089 ;
  assign n27091 = n1542 & n7084 ;
  assign n27093 = ( n1266 & ~n5007 ) | ( n1266 & n5189 ) | ( ~n5007 & n5189 ) ;
  assign n27092 = n6283 | n11176 ;
  assign n27094 = n27093 ^ n27092 ^ 1'b0 ;
  assign n27095 = n27091 | n27094 ;
  assign n27096 = n27095 ^ n25403 ^ 1'b0 ;
  assign n27097 = n17781 ^ n11489 ^ 1'b0 ;
  assign n27098 = n24959 ^ n14950 ^ 1'b0 ;
  assign n27100 = n1941 | n2448 ;
  assign n27099 = n8058 & ~n16648 ;
  assign n27101 = n27100 ^ n27099 ^ 1'b0 ;
  assign n27105 = n1358 | n13509 ;
  assign n27106 = n27105 ^ n15819 ^ 1'b0 ;
  assign n27102 = ~n3887 & n8077 ;
  assign n27103 = n27102 ^ n19142 ^ 1'b0 ;
  assign n27104 = ( n1570 & n10367 ) | ( n1570 & ~n27103 ) | ( n10367 & ~n27103 ) ;
  assign n27107 = n27106 ^ n27104 ^ 1'b0 ;
  assign n27109 = n423 | n21087 ;
  assign n27108 = n2859 & n17579 ;
  assign n27110 = n27109 ^ n27108 ^ 1'b0 ;
  assign n27111 = n1987 | n27110 ;
  assign n27112 = n10919 & ~n12086 ;
  assign n27113 = n16147 & n27112 ;
  assign n27114 = n2946 & ~n15051 ;
  assign n27115 = n27114 ^ n11583 ^ 1'b0 ;
  assign n27116 = ( n4801 & n5044 ) | ( n4801 & n27115 ) | ( n5044 & n27115 ) ;
  assign n27117 = n1641 & ~n3003 ;
  assign n27118 = n8268 ^ n1843 ^ 1'b0 ;
  assign n27119 = n27117 & n27118 ;
  assign n27120 = n27119 ^ n12824 ^ 1'b0 ;
  assign n27121 = n10720 & ~n27120 ;
  assign n27122 = n13732 & ~n21066 ;
  assign n27123 = ~n983 & n27122 ;
  assign n27124 = n9923 ^ n540 ^ 1'b0 ;
  assign n27125 = ~n1413 & n27124 ;
  assign n27126 = n3298 ^ n2127 ^ 1'b0 ;
  assign n27127 = n9210 & ~n27126 ;
  assign n27128 = n25336 ^ n14286 ^ 1'b0 ;
  assign n27130 = n286 & n1832 ;
  assign n27129 = ~n4343 & n12996 ;
  assign n27131 = n27130 ^ n27129 ^ 1'b0 ;
  assign n27132 = ( n1726 & n2663 ) | ( n1726 & n8499 ) | ( n2663 & n8499 ) ;
  assign n27133 = n27132 ^ n3145 ^ 1'b0 ;
  assign n27134 = n18359 ^ n9215 ^ n5077 ;
  assign n27135 = n666 | n16231 ;
  assign n27136 = ~n208 & n25108 ;
  assign n27137 = n5883 & n10361 ;
  assign n27138 = n27137 ^ n4938 ^ 1'b0 ;
  assign n27139 = ( n459 & ~n2179 ) | ( n459 & n5688 ) | ( ~n2179 & n5688 ) ;
  assign n27140 = ( ~n21478 & n23920 ) | ( ~n21478 & n27139 ) | ( n23920 & n27139 ) ;
  assign n27141 = ~n7111 & n17671 ;
  assign n27142 = ~n16330 & n18347 ;
  assign n27143 = n27142 ^ n25759 ^ 1'b0 ;
  assign n27144 = n6911 ^ n1288 ^ 1'b0 ;
  assign n27145 = n5028 | n7513 ;
  assign n27146 = n27145 ^ n15175 ^ 1'b0 ;
  assign n27147 = n27144 & ~n27146 ;
  assign n27148 = n12718 & ~n27147 ;
  assign n27149 = n3569 ^ n3086 ^ 1'b0 ;
  assign n27150 = n5982 & ~n27149 ;
  assign n27151 = n27150 ^ n8596 ^ 1'b0 ;
  assign n27152 = n14343 | n27151 ;
  assign n27153 = n17300 & ~n27152 ;
  assign n27154 = n7785 | n27153 ;
  assign n27155 = n27148 | n27154 ;
  assign n27156 = ~n8227 & n27155 ;
  assign n27157 = n27156 ^ n22962 ^ 1'b0 ;
  assign n27158 = n20460 ^ n9974 ^ 1'b0 ;
  assign n27159 = n74 & ~n680 ;
  assign n27160 = ~n74 & n27159 ;
  assign n27161 = n27160 ^ n21863 ^ 1'b0 ;
  assign n27162 = n4402 | n27161 ;
  assign n27163 = n4468 & n15461 ;
  assign n27164 = n27163 ^ n7787 ^ 1'b0 ;
  assign n27165 = ~n27162 & n27164 ;
  assign n27166 = n11726 & n27165 ;
  assign n27167 = ~n4399 & n27166 ;
  assign n27168 = ~n20704 & n27167 ;
  assign n27169 = n21967 | n27168 ;
  assign n27170 = ~n224 & n25019 ;
  assign n27171 = n27170 ^ n22571 ^ 1'b0 ;
  assign n27172 = n231 & n15966 ;
  assign n27173 = n697 & n27172 ;
  assign n27174 = ( ~n24264 & n26229 ) | ( ~n24264 & n27173 ) | ( n26229 & n27173 ) ;
  assign n27175 = ~n12983 & n24728 ;
  assign n27176 = n27175 ^ n6522 ^ 1'b0 ;
  assign n27177 = n2478 & ~n21674 ;
  assign n27178 = n511 | n27177 ;
  assign n27179 = n27178 ^ n5076 ^ 1'b0 ;
  assign n27180 = n2634 ^ n425 ^ 1'b0 ;
  assign n27181 = ~n22708 & n27180 ;
  assign n27182 = n15531 & n27181 ;
  assign n27183 = n26761 ^ n14471 ^ 1'b0 ;
  assign n27184 = n24467 & n27183 ;
  assign n27186 = ~n3498 & n5189 ;
  assign n27187 = ~n211 & n27186 ;
  assign n27188 = n6367 & n27187 ;
  assign n27185 = n24919 ^ n7128 ^ 1'b0 ;
  assign n27189 = n27188 ^ n27185 ^ 1'b0 ;
  assign n27190 = n15824 | n27189 ;
  assign n27196 = n7810 ^ n6363 ^ 1'b0 ;
  assign n27191 = n22231 ^ n2803 ^ 1'b0 ;
  assign n27192 = ~n3050 & n27191 ;
  assign n27193 = n2474 & ~n17449 ;
  assign n27194 = n18770 & n27193 ;
  assign n27195 = n27192 & ~n27194 ;
  assign n27197 = n27196 ^ n27195 ^ 1'b0 ;
  assign n27198 = n9833 ^ n7377 ^ 1'b0 ;
  assign n27199 = ~n11047 & n27198 ;
  assign n27200 = n3725 & n27199 ;
  assign n27201 = n23363 ^ n16909 ^ 1'b0 ;
  assign n27202 = n25254 | n27201 ;
  assign n27203 = n3649 ^ n695 ^ 1'b0 ;
  assign n27204 = n6100 ^ n189 ^ 1'b0 ;
  assign n27205 = n1609 & ~n4519 ;
  assign n27206 = n7110 | n27205 ;
  assign n27207 = n3646 & ~n27206 ;
  assign n27208 = n24578 ^ n16726 ^ 1'b0 ;
  assign n27209 = n27207 | n27208 ;
  assign n27210 = n19767 ^ n14928 ^ 1'b0 ;
  assign n27211 = ~n27209 & n27210 ;
  assign n27212 = n2341 & ~n9049 ;
  assign n27213 = ~n11400 & n27212 ;
  assign n27214 = n16578 ^ n14324 ^ 1'b0 ;
  assign n27215 = ~n8452 & n27214 ;
  assign n27216 = n27213 & n27215 ;
  assign n27217 = n15885 ^ n7626 ^ 1'b0 ;
  assign n27218 = n23061 ^ n11251 ^ 1'b0 ;
  assign n27219 = n20682 & n27218 ;
  assign n27220 = n3967 & n16902 ;
  assign n27221 = n27220 ^ n5480 ^ 1'b0 ;
  assign n27222 = n27221 ^ n17080 ^ n6098 ;
  assign n27223 = ~n27219 & n27222 ;
  assign n27224 = n27217 & n27223 ;
  assign n27225 = n9751 & ~n16640 ;
  assign n27226 = n11523 | n13257 ;
  assign n27229 = n1152 | n2805 ;
  assign n27230 = n27229 ^ n3462 ^ 1'b0 ;
  assign n27231 = n27230 ^ n13094 ^ n7208 ;
  assign n27227 = n5541 ^ n4738 ^ 1'b0 ;
  assign n27228 = ~n6857 & n27227 ;
  assign n27232 = n27231 ^ n27228 ^ 1'b0 ;
  assign n27233 = n13553 | n18333 ;
  assign n27234 = n8868 ^ n417 ^ 1'b0 ;
  assign n27238 = n5971 | n7591 ;
  assign n27235 = n12673 ^ n8157 ^ 1'b0 ;
  assign n27236 = ( ~n195 & n7027 ) | ( ~n195 & n23552 ) | ( n7027 & n23552 ) ;
  assign n27237 = n27235 & n27236 ;
  assign n27239 = n27238 ^ n27237 ^ 1'b0 ;
  assign n27240 = n27239 ^ n16543 ^ 1'b0 ;
  assign n27241 = n863 & n3403 ;
  assign n27242 = n17403 & n27241 ;
  assign n27243 = n27242 ^ n19173 ^ n6027 ;
  assign n27244 = n27243 ^ n17693 ^ n15934 ;
  assign n27245 = ~n23038 & n27244 ;
  assign n27246 = ~n11006 & n27245 ;
  assign n27247 = ~n2967 & n7449 ;
  assign n27248 = ~n18119 & n27247 ;
  assign n27249 = n27248 ^ n14068 ^ n5806 ;
  assign n27250 = n386 & n443 ;
  assign n27251 = n19762 ^ n2914 ^ 1'b0 ;
  assign n27252 = n27251 ^ n2179 ^ 1'b0 ;
  assign n27253 = n12546 & n27252 ;
  assign n27254 = ( ~n6075 & n6593 ) | ( ~n6075 & n27253 ) | ( n6593 & n27253 ) ;
  assign n27256 = n1829 & ~n2682 ;
  assign n27255 = n3308 | n7576 ;
  assign n27257 = n27256 ^ n27255 ^ 1'b0 ;
  assign n27258 = n445 & ~n2697 ;
  assign n27259 = n7066 & ~n10177 ;
  assign n27260 = ~n4969 & n7528 ;
  assign n27261 = n27260 ^ n1961 ^ 1'b0 ;
  assign n27262 = n11644 ^ n6030 ^ 1'b0 ;
  assign n27263 = ~n9199 & n27262 ;
  assign n27264 = ~n5277 & n12513 ;
  assign n27265 = n11552 & n27264 ;
  assign n27266 = n896 | n27265 ;
  assign n27267 = n27263 | n27266 ;
  assign n27268 = n27267 ^ n18164 ^ 1'b0 ;
  assign n27269 = n1014 & n27268 ;
  assign n27270 = n14254 ^ n9594 ^ 1'b0 ;
  assign n27271 = n7298 & ~n9528 ;
  assign n27272 = n5856 & ~n14930 ;
  assign n27273 = ~n27271 & n27272 ;
  assign n27274 = n6350 & n17605 ;
  assign n27275 = n27274 ^ n25235 ^ 1'b0 ;
  assign n27278 = ( n2353 & n10370 ) | ( n2353 & ~n26723 ) | ( n10370 & ~n26723 ) ;
  assign n27276 = ( n4102 & n7343 ) | ( n4102 & ~n19509 ) | ( n7343 & ~n19509 ) ;
  assign n27277 = ~n2813 & n27276 ;
  assign n27279 = n27278 ^ n27277 ^ 1'b0 ;
  assign n27280 = n4914 & n23953 ;
  assign n27281 = n27280 ^ n959 ^ 1'b0 ;
  assign n27283 = ~n10018 & n24101 ;
  assign n27284 = ~n6074 & n27283 ;
  assign n27282 = n4121 & n5201 ;
  assign n27285 = n27284 ^ n27282 ^ n673 ;
  assign n27286 = n4716 | n6231 ;
  assign n27287 = n27286 ^ n12131 ^ 1'b0 ;
  assign n27288 = n27287 ^ n25346 ^ n10272 ;
  assign n27289 = n9550 & ~n27288 ;
  assign n27290 = n27289 ^ n14453 ^ 1'b0 ;
  assign n27291 = ~n6413 & n23812 ;
  assign n27292 = n27291 ^ n23698 ^ 1'b0 ;
  assign n27293 = n13125 | n17256 ;
  assign n27294 = n1556 | n5260 ;
  assign n27295 = n12309 ^ n2093 ^ 1'b0 ;
  assign n27296 = n3852 | n27295 ;
  assign n27297 = n27296 ^ n15825 ^ 1'b0 ;
  assign n27298 = ~n27294 & n27297 ;
  assign n27299 = n3042 & n27298 ;
  assign n27300 = n1771 & ~n18402 ;
  assign n27301 = ( ~n3382 & n5785 ) | ( ~n3382 & n6116 ) | ( n5785 & n6116 ) ;
  assign n27302 = ~n6082 & n27301 ;
  assign n27303 = n27302 ^ n2560 ^ 1'b0 ;
  assign n27304 = n1887 ^ n927 ^ 1'b0 ;
  assign n27305 = n27304 ^ n8924 ^ 1'b0 ;
  assign n27306 = ~n27303 & n27305 ;
  assign n27307 = n1884 & n5816 ;
  assign n27308 = n1749 | n23958 ;
  assign n27309 = ( n20641 & n27307 ) | ( n20641 & ~n27308 ) | ( n27307 & ~n27308 ) ;
  assign n27310 = n10618 ^ n10143 ^ 1'b0 ;
  assign n27311 = n27310 ^ n13758 ^ n7965 ;
  assign n27312 = n23053 ^ n5244 ^ 1'b0 ;
  assign n27313 = ~n7898 & n13108 ;
  assign n27314 = ~n25268 & n27313 ;
  assign n27315 = n24886 ^ n13085 ^ 1'b0 ;
  assign n27317 = n7735 & ~n17191 ;
  assign n27318 = n27317 ^ n6876 ^ 1'b0 ;
  assign n27316 = n2097 | n23917 ;
  assign n27319 = n27318 ^ n27316 ^ 1'b0 ;
  assign n27320 = n19110 ^ n2102 ^ 1'b0 ;
  assign n27321 = n5518 & ~n9755 ;
  assign n27322 = n26697 ^ n22870 ^ 1'b0 ;
  assign n27323 = n27321 & ~n27322 ;
  assign n27324 = n26983 ^ n2442 ^ 1'b0 ;
  assign n27326 = n14842 ^ n7842 ^ 1'b0 ;
  assign n27325 = ~n5095 & n14642 ;
  assign n27327 = n27326 ^ n27325 ^ 1'b0 ;
  assign n27328 = ~n2391 & n27327 ;
  assign n27329 = ~n14010 & n27328 ;
  assign n27330 = n22927 ^ n11383 ^ n7077 ;
  assign n27331 = n27330 ^ n23275 ^ n7001 ;
  assign n27332 = ~n7531 & n9790 ;
  assign n27333 = ( n780 & ~n8756 ) | ( n780 & n15151 ) | ( ~n8756 & n15151 ) ;
  assign n27334 = n4568 & n5141 ;
  assign n27335 = n12949 | n27334 ;
  assign n27336 = n15230 | n27335 ;
  assign n27337 = ~n8370 & n27336 ;
  assign n27338 = n2309 & ~n20236 ;
  assign n27339 = n18968 | n27144 ;
  assign n27340 = ( ~n15798 & n22181 ) | ( ~n15798 & n27339 ) | ( n22181 & n27339 ) ;
  assign n27341 = n788 | n13601 ;
  assign n27342 = n15119 ^ n9121 ^ 1'b0 ;
  assign n27343 = n24974 & ~n27342 ;
  assign n27344 = ~n685 & n2216 ;
  assign n27345 = n27344 ^ n2999 ^ 1'b0 ;
  assign n27346 = n16299 | n27345 ;
  assign n27347 = n654 | n754 ;
  assign n27348 = n11358 | n27347 ;
  assign n27349 = ~n40 & n27348 ;
  assign n27350 = n17054 & n23948 ;
  assign n27351 = n8547 & ~n17712 ;
  assign n27352 = n27351 ^ n7294 ^ 1'b0 ;
  assign n27356 = n5719 | n19516 ;
  assign n27357 = n16747 ^ n4537 ^ 1'b0 ;
  assign n27358 = n27356 & ~n27357 ;
  assign n27359 = n27358 ^ n8566 ^ 1'b0 ;
  assign n27353 = n1219 & ~n11786 ;
  assign n27354 = n4875 | n27353 ;
  assign n27355 = n3414 | n27354 ;
  assign n27360 = n27359 ^ n27355 ^ 1'b0 ;
  assign n27361 = n13218 | n17853 ;
  assign n27362 = n12788 | n27361 ;
  assign n27363 = n5206 ^ n4605 ^ 1'b0 ;
  assign n27364 = n3724 | n10173 ;
  assign n27365 = n27364 ^ n6254 ^ 1'b0 ;
  assign n27366 = n27365 ^ n2273 ^ n949 ;
  assign n27367 = n6110 | n27366 ;
  assign n27368 = n27367 ^ n18751 ^ 1'b0 ;
  assign n27369 = ( ~n5443 & n27363 ) | ( ~n5443 & n27368 ) | ( n27363 & n27368 ) ;
  assign n27370 = n2040 | n7597 ;
  assign n27371 = ( n7008 & n23066 ) | ( n7008 & n27370 ) | ( n23066 & n27370 ) ;
  assign n27372 = n27371 ^ n5636 ^ 1'b0 ;
  assign n27373 = n27321 & n27372 ;
  assign n27374 = n3211 | n9457 ;
  assign n27375 = n20207 & ~n27374 ;
  assign n27376 = ( n5244 & n6563 ) | ( n5244 & n27375 ) | ( n6563 & n27375 ) ;
  assign n27377 = ~n2661 & n27376 ;
  assign n27378 = n2661 & n27377 ;
  assign n27379 = n27373 & ~n27378 ;
  assign n27380 = ~n27373 & n27379 ;
  assign n27381 = n7459 ^ n4053 ^ 1'b0 ;
  assign n27382 = n7321 & n27381 ;
  assign n27383 = ~n1354 & n20226 ;
  assign n27384 = n3424 ^ n439 ^ 1'b0 ;
  assign n27385 = n2873 & n27384 ;
  assign n27386 = n5328 | n7066 ;
  assign n27387 = n12891 ^ n6273 ^ n5497 ;
  assign n27388 = n19062 & n23798 ;
  assign n27389 = ~n11126 & n27388 ;
  assign n27390 = n3444 | n10069 ;
  assign n27391 = n10069 & ~n27390 ;
  assign n27392 = n27391 ^ n1493 ^ 1'b0 ;
  assign n27393 = n10294 | n25684 ;
  assign n27394 = n243 | n27393 ;
  assign n27395 = ~n19889 & n20994 ;
  assign n27396 = n27395 ^ n22533 ^ n21433 ;
  assign n27397 = n22157 ^ n8573 ^ 1'b0 ;
  assign n27398 = n2112 | n3125 ;
  assign n27399 = n15699 ^ n3477 ^ 1'b0 ;
  assign n27400 = n27398 & ~n27399 ;
  assign n27401 = n189 | n1040 ;
  assign n27402 = n27400 | n27401 ;
  assign n27403 = n4180 ^ n525 ^ 1'b0 ;
  assign n27405 = n19018 ^ n8565 ^ 1'b0 ;
  assign n27404 = n17124 ^ n3314 ^ 1'b0 ;
  assign n27406 = n27405 ^ n27404 ^ n13384 ;
  assign n27407 = n22191 ^ n5638 ^ n1570 ;
  assign n27408 = n27407 ^ n12805 ^ 1'b0 ;
  assign n27409 = n8060 & n27408 ;
  assign n27410 = n18945 & n27409 ;
  assign n27411 = ~n1329 & n18534 ;
  assign n27412 = ~n16467 & n27411 ;
  assign n27413 = n27412 ^ n17461 ^ 1'b0 ;
  assign n27414 = ~n16935 & n27413 ;
  assign n27415 = n765 & ~n9056 ;
  assign n27416 = n27415 ^ n21800 ^ 1'b0 ;
  assign n27417 = n18435 ^ n13402 ^ 1'b0 ;
  assign n27418 = n6437 ^ n2082 ^ 1'b0 ;
  assign n27419 = n27418 ^ n1469 ^ 1'b0 ;
  assign n27420 = n1823 & n27419 ;
  assign n27421 = ~n27417 & n27420 ;
  assign n27422 = n3796 & ~n13582 ;
  assign n27423 = n27422 ^ n5423 ^ 1'b0 ;
  assign n27424 = n4819 & ~n25436 ;
  assign n27425 = ~n10945 & n27424 ;
  assign n27426 = n9522 | n26052 ;
  assign n27427 = n7045 & ~n27426 ;
  assign n27428 = n27427 ^ n4795 ^ 1'b0 ;
  assign n27429 = n19339 ^ n16026 ^ 1'b0 ;
  assign n27430 = ~n9797 & n27429 ;
  assign n27431 = n27430 ^ n15203 ^ 1'b0 ;
  assign n27432 = ~n9549 & n9663 ;
  assign n27433 = n340 & ~n5317 ;
  assign n27434 = ( n11445 & n27432 ) | ( n11445 & ~n27433 ) | ( n27432 & ~n27433 ) ;
  assign n27435 = n10319 ^ n7961 ^ 1'b0 ;
  assign n27436 = n27434 | n27435 ;
  assign n27437 = n16021 | n27436 ;
  assign n27438 = n7887 ^ n790 ^ 1'b0 ;
  assign n27439 = n1329 & ~n27438 ;
  assign n27440 = n827 & n27439 ;
  assign n27441 = ~n24543 & n27440 ;
  assign n27442 = n306 & ~n18295 ;
  assign n27443 = n27441 & n27442 ;
  assign n27445 = n2952 & n21029 ;
  assign n27446 = n27445 ^ n4333 ^ 1'b0 ;
  assign n27444 = ~n6475 & n9674 ;
  assign n27447 = n27446 ^ n27444 ^ 1'b0 ;
  assign n27448 = n5121 & ~n8258 ;
  assign n27449 = ~n10023 & n10958 ;
  assign n27450 = ~n10024 & n15084 ;
  assign n27451 = n27450 ^ n1941 ^ 1'b0 ;
  assign n27452 = n9147 ^ n3214 ^ 1'b0 ;
  assign n27453 = n1469 & ~n27452 ;
  assign n27454 = n10031 | n25152 ;
  assign n27455 = n17124 ^ n4095 ^ 1'b0 ;
  assign n27458 = ~n12368 & n14138 ;
  assign n27459 = ~n3835 & n27458 ;
  assign n27456 = n4386 & ~n5868 ;
  assign n27457 = ~n24442 & n27456 ;
  assign n27460 = n27459 ^ n27457 ^ 1'b0 ;
  assign n27461 = n4757 ^ n1804 ^ 1'b0 ;
  assign n27462 = n10356 ^ n2474 ^ 1'b0 ;
  assign n27463 = n1460 | n27462 ;
  assign n27464 = n16803 & ~n27463 ;
  assign n27466 = n4538 ^ n2604 ^ 1'b0 ;
  assign n27467 = n27466 ^ n15389 ^ 1'b0 ;
  assign n27468 = n6524 & n27467 ;
  assign n27469 = n27468 ^ n271 ^ 1'b0 ;
  assign n27470 = n27469 ^ n15009 ^ 1'b0 ;
  assign n27465 = n2352 | n25388 ;
  assign n27471 = n27470 ^ n27465 ^ 1'b0 ;
  assign n27472 = n27469 ^ n11870 ^ 1'b0 ;
  assign n27473 = n4241 & n15953 ;
  assign n27474 = ~n15953 & n27473 ;
  assign n27475 = n16847 | n27474 ;
  assign n27476 = n27475 ^ n4298 ^ 1'b0 ;
  assign n27477 = n7443 & n11712 ;
  assign n27478 = n2991 & n10166 ;
  assign n27479 = n15653 & n27478 ;
  assign n27480 = n3280 & n27479 ;
  assign n27481 = n415 | n14351 ;
  assign n27482 = n27481 ^ n1962 ^ 1'b0 ;
  assign n27483 = n4989 & ~n11292 ;
  assign n27484 = ~n13837 & n27483 ;
  assign n27485 = n27484 ^ n367 ^ 1'b0 ;
  assign n27486 = n22918 & n24510 ;
  assign n27487 = n551 | n6291 ;
  assign n27488 = n16923 & ~n27487 ;
  assign n27489 = n3409 & ~n27488 ;
  assign n27490 = n4207 & ~n17479 ;
  assign n27491 = n27490 ^ n23956 ^ 1'b0 ;
  assign n27492 = n17499 & n27491 ;
  assign n27493 = ~n10803 & n19931 ;
  assign n27494 = n21293 ^ n9194 ^ 1'b0 ;
  assign n27495 = ~n27493 & n27494 ;
  assign n27496 = n10315 & ~n25403 ;
  assign n27497 = n27496 ^ n13823 ^ 1'b0 ;
  assign n27498 = n2246 ^ n1701 ^ 1'b0 ;
  assign n27499 = n27498 ^ n2649 ^ 1'b0 ;
  assign n27500 = n5442 & ~n6726 ;
  assign n27501 = n9724 & n27500 ;
  assign n27502 = n27501 ^ n7140 ^ 1'b0 ;
  assign n27503 = ~n22224 & n27502 ;
  assign n27504 = n27499 & n27503 ;
  assign n27505 = n1883 ^ n1852 ^ 1'b0 ;
  assign n27506 = n7609 | n27505 ;
  assign n27507 = n3564 ^ n2808 ^ 1'b0 ;
  assign n27508 = n7067 ^ n6527 ^ 1'b0 ;
  assign n27509 = n88 | n10584 ;
  assign n27510 = ~n15147 & n27509 ;
  assign n27511 = n11320 & n27510 ;
  assign n27512 = n26730 ^ n7979 ^ n647 ;
  assign n27513 = n26357 & ~n27512 ;
  assign n27514 = ( n6394 & n14123 ) | ( n6394 & ~n27513 ) | ( n14123 & ~n27513 ) ;
  assign n27515 = ( n5143 & ~n6254 ) | ( n5143 & n23389 ) | ( ~n6254 & n23389 ) ;
  assign n27519 = n15468 ^ n2694 ^ 1'b0 ;
  assign n27516 = n12383 & n25005 ;
  assign n27517 = n4182 & ~n27516 ;
  assign n27518 = ~n21792 & n27517 ;
  assign n27520 = n27519 ^ n27518 ^ 1'b0 ;
  assign n27521 = ~n27515 & n27520 ;
  assign n27522 = n5005 | n26789 ;
  assign n27523 = n8119 & ~n26858 ;
  assign n27524 = n2373 & n4074 ;
  assign n27525 = n15769 | n27524 ;
  assign n27526 = ~n16010 & n16806 ;
  assign n27527 = n27526 ^ n2849 ^ 1'b0 ;
  assign n27528 = n18164 ^ n6124 ^ 1'b0 ;
  assign n27529 = n1347 & ~n27528 ;
  assign n27530 = n7588 & n27312 ;
  assign n27531 = n27530 ^ n6472 ^ 1'b0 ;
  assign n27533 = n3072 & ~n5188 ;
  assign n27532 = n9137 & n17337 ;
  assign n27534 = n27533 ^ n27532 ^ 1'b0 ;
  assign n27535 = n8230 ^ n4960 ^ 1'b0 ;
  assign n27536 = n25604 ^ n16062 ^ 1'b0 ;
  assign n27537 = n11274 & n15005 ;
  assign n27538 = ~n6060 & n27537 ;
  assign n27539 = n21402 ^ n93 ^ 1'b0 ;
  assign n27540 = n8970 | n27539 ;
  assign n27541 = n27540 ^ x1 ^ 1'b0 ;
  assign n27542 = n18934 ^ n5781 ^ 1'b0 ;
  assign n27543 = n27542 ^ n26541 ^ 1'b0 ;
  assign n27544 = n146 | n9850 ;
  assign n27545 = n17802 | n27544 ;
  assign n27546 = n2872 & n8732 ;
  assign n27547 = n27546 ^ n5708 ^ 1'b0 ;
  assign n27548 = ~n26405 & n27547 ;
  assign n27549 = n19060 & n21889 ;
  assign n27550 = ( n5371 & n6927 ) | ( n5371 & ~n26975 ) | ( n6927 & ~n26975 ) ;
  assign n27551 = n12291 & n18992 ;
  assign n27552 = ~n625 & n27551 ;
  assign n27553 = n9680 | n12344 ;
  assign n27558 = n5929 | n15584 ;
  assign n27554 = ( n690 & ~n3177 ) | ( n690 & n3586 ) | ( ~n3177 & n3586 ) ;
  assign n27555 = ~n12618 & n27554 ;
  assign n27556 = n27555 ^ n1809 ^ n1653 ;
  assign n27557 = n9316 & n27556 ;
  assign n27559 = n27558 ^ n27557 ^ 1'b0 ;
  assign n27560 = n15893 ^ n14844 ^ 1'b0 ;
  assign n27561 = n966 & ~n27560 ;
  assign n27562 = n4173 ^ n3813 ^ 1'b0 ;
  assign n27563 = n25557 & ~n27562 ;
  assign n27564 = n741 | n18418 ;
  assign n27565 = n27369 & ~n27564 ;
  assign n27566 = n5047 ^ n3255 ^ n2444 ;
  assign n27567 = n22757 & n27566 ;
  assign n27568 = n27567 ^ n6292 ^ 1'b0 ;
  assign n27569 = n16670 ^ n7303 ^ 1'b0 ;
  assign n27570 = n17115 ^ n7352 ^ 1'b0 ;
  assign n27571 = ~n23693 & n27570 ;
  assign n27572 = ~n7842 & n26550 ;
  assign n27573 = ~n27571 & n27572 ;
  assign n27574 = ~n4009 & n6757 ;
  assign n27575 = n27574 ^ n998 ^ 1'b0 ;
  assign n27576 = n25975 ^ n5974 ^ 1'b0 ;
  assign n27579 = n23997 ^ n21941 ^ 1'b0 ;
  assign n27577 = n5911 | n13990 ;
  assign n27578 = n14555 & ~n27577 ;
  assign n27580 = n27579 ^ n27578 ^ 1'b0 ;
  assign n27581 = n1439 & n9433 ;
  assign n27582 = n27581 ^ n2719 ^ 1'b0 ;
  assign n27583 = n27582 ^ n17704 ^ 1'b0 ;
  assign n27584 = ~n1590 & n27583 ;
  assign n27585 = ~n8012 & n20191 ;
  assign n27586 = n4114 | n27585 ;
  assign n27587 = ~n3039 & n4926 ;
  assign n27588 = n27586 & ~n27587 ;
  assign n27589 = n27588 ^ n15662 ^ 1'b0 ;
  assign n27590 = n2141 & n9369 ;
  assign n27591 = n27590 ^ n388 ^ 1'b0 ;
  assign n27592 = ~n16720 & n27591 ;
  assign n27593 = n5394 | n7808 ;
  assign n27594 = ~n5314 & n7359 ;
  assign n27595 = n27594 ^ n10790 ^ 1'b0 ;
  assign n27596 = n1932 | n12307 ;
  assign n27597 = n27596 ^ n5985 ^ 1'b0 ;
  assign n27599 = n6925 ^ n6271 ^ 1'b0 ;
  assign n27598 = n17683 & n25457 ;
  assign n27600 = n27599 ^ n27598 ^ n17605 ;
  assign n27601 = n27600 ^ n7366 ^ n3136 ;
  assign n27602 = n3384 ^ n1697 ^ 1'b0 ;
  assign n27603 = n18760 & n23331 ;
  assign n27604 = n27603 ^ n25732 ^ 1'b0 ;
  assign n27605 = n25307 ^ n13904 ^ 1'b0 ;
  assign n27606 = n781 & ~n13155 ;
  assign n27607 = n1157 & n11077 ;
  assign n27608 = n27606 & n27607 ;
  assign n27609 = n1382 & ~n27608 ;
  assign n27610 = n27609 ^ n19034 ^ 1'b0 ;
  assign n27611 = n18923 & n27610 ;
  assign n27612 = n6333 ^ n903 ^ 1'b0 ;
  assign n27613 = ( n16508 & n27312 ) | ( n16508 & n27612 ) | ( n27312 & n27612 ) ;
  assign n27614 = n1988 & ~n21186 ;
  assign n27615 = n4537 ^ n312 ^ 1'b0 ;
  assign n27616 = n4979 & n27615 ;
  assign n27617 = n3828 & n10209 ;
  assign n27618 = n27617 ^ n15948 ^ 1'b0 ;
  assign n27619 = n27616 & ~n27618 ;
  assign n27620 = ( n1301 & ~n6264 ) | ( n1301 & n9539 ) | ( ~n6264 & n9539 ) ;
  assign n27621 = n10470 ^ n9500 ^ 1'b0 ;
  assign n27622 = n24281 | n27621 ;
  assign n27623 = n27620 & ~n27622 ;
  assign n27624 = ~n4991 & n8441 ;
  assign n27625 = n13059 ^ n6051 ^ n1295 ;
  assign n27626 = n3530 ^ n1816 ^ 1'b0 ;
  assign n27627 = n12754 | n27626 ;
  assign n27628 = n69 & ~n27627 ;
  assign n27629 = ~n27625 & n27628 ;
  assign n27630 = n27624 & n27629 ;
  assign n27631 = n6643 & n27630 ;
  assign n27632 = n7277 ^ n4995 ^ 1'b0 ;
  assign n27633 = n2343 & ~n27632 ;
  assign n27638 = ~n3498 & n4859 ;
  assign n27639 = n27638 ^ n7536 ^ 1'b0 ;
  assign n27634 = ~n815 & n1832 ;
  assign n27635 = ~n4359 & n27634 ;
  assign n27636 = n27635 ^ n13412 ^ n4241 ;
  assign n27637 = ~n6774 & n27636 ;
  assign n27640 = n27639 ^ n27637 ^ 1'b0 ;
  assign n27641 = n2721 ^ n437 ^ 1'b0 ;
  assign n27642 = n27641 ^ n6860 ^ 1'b0 ;
  assign n27643 = n27642 ^ n13438 ^ 1'b0 ;
  assign n27644 = n25910 ^ n13585 ^ 1'b0 ;
  assign n27645 = ~n2262 & n16407 ;
  assign n27651 = n17287 & ~n26577 ;
  assign n27646 = n14277 ^ n5166 ^ 1'b0 ;
  assign n27647 = n7715 & ~n27646 ;
  assign n27648 = n8275 & ~n13596 ;
  assign n27649 = ~n15076 & n27648 ;
  assign n27650 = n27647 | n27649 ;
  assign n27652 = n27651 ^ n27650 ^ 1'b0 ;
  assign n27653 = n27645 | n27652 ;
  assign n27654 = n736 & n1596 ;
  assign n27655 = n27654 ^ n8763 ^ 1'b0 ;
  assign n27656 = n27655 ^ n25998 ^ 1'b0 ;
  assign n27657 = n1574 & ~n27656 ;
  assign n27658 = ~n14030 & n21950 ;
  assign n27659 = n27658 ^ n1714 ^ 1'b0 ;
  assign n27660 = n10465 & ~n11304 ;
  assign n27661 = n27660 ^ n2780 ^ 1'b0 ;
  assign n27662 = n20547 ^ n20260 ^ 1'b0 ;
  assign n27663 = n27661 & ~n27662 ;
  assign n27664 = n27663 ^ n14835 ^ 1'b0 ;
  assign n27665 = n4523 | n22445 ;
  assign n27666 = n9651 | n27665 ;
  assign n27667 = n3513 | n11273 ;
  assign n27668 = n5644 | n27667 ;
  assign n27669 = ~n115 & n27668 ;
  assign n27670 = n7927 & ~n27669 ;
  assign n27671 = n9639 & ~n20996 ;
  assign n27672 = n27671 ^ n20812 ^ 1'b0 ;
  assign n27673 = ~n12654 & n21320 ;
  assign n27674 = n25567 ^ n22448 ^ 1'b0 ;
  assign n27675 = n8869 ^ n6452 ^ 1'b0 ;
  assign n27676 = n27674 | n27675 ;
  assign n27677 = n27676 ^ n5300 ^ 1'b0 ;
  assign n27678 = n27673 & n27677 ;
  assign n27679 = n3052 | n11476 ;
  assign n27680 = n27679 ^ n23595 ^ 1'b0 ;
  assign n27681 = ~n11899 & n16062 ;
  assign n27682 = n4506 ^ n1405 ^ n459 ;
  assign n27683 = n27682 ^ n1337 ^ 1'b0 ;
  assign n27684 = x1 & n27683 ;
  assign n27685 = n26520 ^ n6885 ^ n3212 ;
  assign n27686 = ~n20131 & n22781 ;
  assign n27687 = n27686 ^ n16019 ^ 1'b0 ;
  assign n27688 = ~n26688 & n27687 ;
  assign n27690 = n488 & n14518 ;
  assign n27691 = n10319 & n27690 ;
  assign n27689 = n5034 & ~n26837 ;
  assign n27692 = n27691 ^ n27689 ^ 1'b0 ;
  assign n27693 = ~n6749 & n27692 ;
  assign n27694 = ~n26571 & n27693 ;
  assign n27695 = ~n16044 & n17128 ;
  assign n27696 = n27694 & n27695 ;
  assign n27697 = n11068 ^ n5190 ^ 1'b0 ;
  assign n27698 = n1726 | n27697 ;
  assign n27699 = n6409 ^ n4976 ^ 1'b0 ;
  assign n27700 = n2639 & n27699 ;
  assign n27701 = ~n27698 & n27700 ;
  assign n27702 = n27701 ^ n11905 ^ 1'b0 ;
  assign n27705 = ~n9145 & n15027 ;
  assign n27706 = n27705 ^ n24162 ^ 1'b0 ;
  assign n27703 = ( ~n10963 & n17499 ) | ( ~n10963 & n22218 ) | ( n17499 & n22218 ) ;
  assign n27704 = ~n11153 & n27703 ;
  assign n27707 = n27706 ^ n27704 ^ 1'b0 ;
  assign n27708 = ~n4560 & n5259 ;
  assign n27709 = n27708 ^ n4884 ^ 1'b0 ;
  assign n27710 = ~n2835 & n7632 ;
  assign n27711 = n27709 & n27710 ;
  assign n27712 = ~n3802 & n27711 ;
  assign n27713 = n14582 & ~n27712 ;
  assign n27714 = ~n14325 & n15596 ;
  assign n27715 = n27714 ^ n8136 ^ 1'b0 ;
  assign n27716 = n9331 ^ n2359 ^ 1'b0 ;
  assign n27717 = ( n2421 & n2754 ) | ( n2421 & n12763 ) | ( n2754 & n12763 ) ;
  assign n27718 = n1551 & ~n4833 ;
  assign n27719 = n2415 | n12485 ;
  assign n27720 = ~n304 & n27719 ;
  assign n27721 = ~n14728 & n21884 ;
  assign n27722 = n765 & n5630 ;
  assign n27723 = n27722 ^ n18359 ^ 1'b0 ;
  assign n27724 = n10958 ^ n3017 ^ 1'b0 ;
  assign n27725 = n27723 & ~n27724 ;
  assign n27726 = ( n290 & n17891 ) | ( n290 & ~n27725 ) | ( n17891 & ~n27725 ) ;
  assign n27727 = n4088 & n6998 ;
  assign n27728 = n27727 ^ n16714 ^ n15376 ;
  assign n27729 = n27728 ^ n6857 ^ 1'b0 ;
  assign n27730 = ~n2004 & n2847 ;
  assign n27731 = n3867 ^ n2753 ^ 1'b0 ;
  assign n27732 = n11169 ^ n1157 ^ 1'b0 ;
  assign n27733 = n16720 & n27732 ;
  assign n27734 = n9319 | n20505 ;
  assign n27735 = n22538 & ~n27734 ;
  assign n27736 = n3483 & ~n4937 ;
  assign n27737 = ~n3021 & n27736 ;
  assign n27738 = n703 & n5202 ;
  assign n27739 = ~n13704 & n15443 ;
  assign n27740 = n27739 ^ n18195 ^ 1'b0 ;
  assign n27741 = n10879 & n27740 ;
  assign n27742 = ~n27370 & n27741 ;
  assign n27743 = n27738 | n27742 ;
  assign n27744 = n27743 ^ n8822 ^ 1'b0 ;
  assign n27745 = n2628 ^ n184 ^ 1'b0 ;
  assign n27746 = n7251 & ~n27745 ;
  assign n27747 = n1186 | n8031 ;
  assign n27748 = n27747 ^ n4175 ^ 1'b0 ;
  assign n27749 = n12836 & ~n27748 ;
  assign n27750 = n27749 ^ n7198 ^ n255 ;
  assign n27751 = n16405 ^ n9325 ^ 1'b0 ;
  assign n27752 = n1933 | n2317 ;
  assign n27753 = n490 & ~n3760 ;
  assign n27760 = n25131 ^ n3726 ^ 1'b0 ;
  assign n27761 = n8145 & n27760 ;
  assign n27754 = n19494 ^ n14587 ^ 1'b0 ;
  assign n27755 = n13555 | n27754 ;
  assign n27756 = n22779 & ~n27755 ;
  assign n27757 = n27756 ^ n22057 ^ n14235 ;
  assign n27758 = n1969 & ~n5323 ;
  assign n27759 = ~n27757 & n27758 ;
  assign n27762 = n27761 ^ n27759 ^ 1'b0 ;
  assign n27763 = n5051 & n18255 ;
  assign n27764 = n27763 ^ n4479 ^ 1'b0 ;
  assign n27765 = n26468 & ~n27764 ;
  assign n27766 = ~n6663 & n20642 ;
  assign n27767 = n7835 | n9630 ;
  assign n27768 = n12901 ^ n1071 ^ 1'b0 ;
  assign n27769 = n502 & n27768 ;
  assign n27770 = n430 & n13487 ;
  assign n27771 = n10001 & n27770 ;
  assign n27772 = n591 ^ n287 ^ 1'b0 ;
  assign n27773 = n18260 & ~n27772 ;
  assign n27775 = ( n1267 & n9077 ) | ( n1267 & n10460 ) | ( n9077 & n10460 ) ;
  assign n27774 = n4931 & n11234 ;
  assign n27776 = n27775 ^ n27774 ^ 1'b0 ;
  assign n27777 = n23720 ^ n22744 ^ n15876 ;
  assign n27778 = n6927 | n17994 ;
  assign n27779 = n22629 ^ n1372 ^ n395 ;
  assign n27780 = ~n18124 & n27779 ;
  assign n27781 = n8505 ^ n30 ^ 1'b0 ;
  assign n27782 = n27781 ^ n946 ^ 1'b0 ;
  assign n27783 = ~n27780 & n27782 ;
  assign n27784 = n2895 & n18647 ;
  assign n27785 = n9091 & n27784 ;
  assign n27786 = ~n792 & n8824 ;
  assign n27787 = ~n17459 & n27786 ;
  assign n27788 = n6563 ^ n4805 ^ 1'b0 ;
  assign n27789 = n17788 ^ n4033 ^ 1'b0 ;
  assign n27790 = n27788 & ~n27789 ;
  assign n27791 = n27790 ^ n3909 ^ 1'b0 ;
  assign n27792 = ~n27787 & n27791 ;
  assign n27793 = ~n9564 & n26727 ;
  assign n27794 = n7881 & ~n17233 ;
  assign n27795 = n21916 & n27794 ;
  assign n27796 = n20440 | n27795 ;
  assign n27797 = n9662 & ~n19906 ;
  assign n27798 = n27797 ^ n2772 ^ 1'b0 ;
  assign n27799 = ~n15191 & n22406 ;
  assign n27800 = n11891 ^ n2373 ^ 1'b0 ;
  assign n27801 = n378 | n24667 ;
  assign n27802 = n27801 ^ n3571 ^ 1'b0 ;
  assign n27803 = n13730 ^ n12523 ^ 1'b0 ;
  assign n27804 = n10460 & n27803 ;
  assign n27805 = n1141 & n27804 ;
  assign n27806 = n17198 & n27805 ;
  assign n27807 = n8220 & ~n22983 ;
  assign n27809 = n12719 & n23233 ;
  assign n27810 = n9432 & n27809 ;
  assign n27808 = ~n6074 & n8959 ;
  assign n27811 = n27810 ^ n27808 ^ 1'b0 ;
  assign n27812 = ~n1226 & n22936 ;
  assign n27813 = n19639 ^ n6316 ^ 1'b0 ;
  assign n27814 = n4010 & n12361 ;
  assign n27815 = n3390 & ~n20362 ;
  assign n27816 = n8208 ^ n4581 ^ n4555 ;
  assign n27817 = n27816 ^ n11816 ^ n10209 ;
  assign n27818 = n12103 ^ n4009 ^ 1'b0 ;
  assign n27819 = ( n1987 & n8349 ) | ( n1987 & n27818 ) | ( n8349 & n27818 ) ;
  assign n27820 = n27819 ^ n519 ^ 1'b0 ;
  assign n27821 = n13041 & ~n27820 ;
  assign n27822 = n1173 & n19710 ;
  assign n27823 = n6869 | n27822 ;
  assign n27824 = n27823 ^ n14351 ^ 1'b0 ;
  assign n27825 = n6774 | n15000 ;
  assign n27826 = n10646 ^ n5869 ^ 1'b0 ;
  assign n27827 = n17767 | n27826 ;
  assign n27828 = ~n768 & n7513 ;
  assign n27829 = ~n4040 & n27828 ;
  assign n27830 = n17129 ^ n5226 ^ 1'b0 ;
  assign n27832 = n315 | n7270 ;
  assign n27831 = ~n13342 & n20350 ;
  assign n27833 = n27832 ^ n27831 ^ 1'b0 ;
  assign n27834 = n14739 ^ n14081 ^ 1'b0 ;
  assign n27835 = n8931 | n27834 ;
  assign n27836 = n774 & n27835 ;
  assign n27838 = n6961 & n9832 ;
  assign n27839 = n7067 & n27838 ;
  assign n27837 = n13381 | n24248 ;
  assign n27840 = n27839 ^ n27837 ^ 1'b0 ;
  assign n27841 = ~n3809 & n27840 ;
  assign n27842 = n15893 ^ n10212 ^ n2108 ;
  assign n27843 = n2764 & n27842 ;
  assign n27844 = n846 | n18510 ;
  assign n27845 = n22233 | n27844 ;
  assign n27846 = n27845 ^ n25447 ^ 1'b0 ;
  assign n27847 = ~n2703 & n15138 ;
  assign n27848 = n2335 & n2665 ;
  assign n27849 = n1385 & n27848 ;
  assign n27850 = ~n373 & n13212 ;
  assign n27851 = n27850 ^ n4058 ^ 1'b0 ;
  assign n27852 = n27849 | n27851 ;
  assign n27853 = n7500 & ~n27852 ;
  assign n27854 = n5485 & ~n21545 ;
  assign n27855 = n14938 & n27854 ;
  assign n27856 = n27855 ^ n3617 ^ 1'b0 ;
  assign n27857 = n7147 & n11276 ;
  assign n27858 = n6256 & ~n17358 ;
  assign n27859 = n9170 | n27858 ;
  assign n27860 = n21557 | n27859 ;
  assign n27861 = n7130 ^ n1488 ^ 1'b0 ;
  assign n27862 = n1542 & ~n27861 ;
  assign n27863 = n2140 & n27862 ;
  assign n27864 = n27863 ^ n3428 ^ 1'b0 ;
  assign n27865 = n23772 ^ n1466 ^ 1'b0 ;
  assign n27866 = n27864 | n27865 ;
  assign n27867 = n5136 & n7675 ;
  assign n27868 = n27867 ^ n13699 ^ 1'b0 ;
  assign n27869 = n7237 & ~n14092 ;
  assign n27870 = n254 & n675 ;
  assign n27871 = ~n9921 & n27870 ;
  assign n27872 = n27871 ^ n5880 ^ 1'b0 ;
  assign n27873 = n5546 & n23834 ;
  assign n27874 = ( ~n27869 & n27872 ) | ( ~n27869 & n27873 ) | ( n27872 & n27873 ) ;
  assign n27875 = n13841 ^ n3420 ^ 1'b0 ;
  assign n27876 = n14299 & n27875 ;
  assign n27877 = n5630 ^ n5235 ^ 1'b0 ;
  assign n27878 = n2098 & n27877 ;
  assign n27879 = n864 | n12062 ;
  assign n27880 = n27879 ^ n16580 ^ 1'b0 ;
  assign n27881 = n7207 | n27880 ;
  assign n27882 = n18909 & n25960 ;
  assign n27883 = n27882 ^ n13356 ^ 1'b0 ;
  assign n27884 = n8366 ^ n2741 ^ 1'b0 ;
  assign n27885 = n22923 ^ n6745 ^ n3213 ;
  assign n27886 = ( n23207 & n27884 ) | ( n23207 & n27885 ) | ( n27884 & n27885 ) ;
  assign n27887 = n10783 & n12239 ;
  assign n27888 = n27887 ^ n255 ^ 1'b0 ;
  assign n27889 = n27888 ^ n453 ^ 1'b0 ;
  assign n27893 = n13192 | n14994 ;
  assign n27894 = n924 | n27893 ;
  assign n27890 = n18191 ^ n571 ^ 1'b0 ;
  assign n27891 = n1211 & ~n27890 ;
  assign n27892 = n22205 | n27891 ;
  assign n27895 = n27894 ^ n27892 ^ 1'b0 ;
  assign n27896 = n12133 & n18222 ;
  assign n27897 = n4346 & n27896 ;
  assign n27898 = n3408 & ~n26296 ;
  assign n27899 = ~n27897 & n27898 ;
  assign n27900 = n6527 ^ n74 ^ 1'b0 ;
  assign n27901 = ~n6568 & n8177 ;
  assign n27902 = n27901 ^ n20796 ^ 1'b0 ;
  assign n27903 = n19714 | n27902 ;
  assign n27904 = n7749 & ~n27903 ;
  assign n27905 = n2108 ^ n772 ^ 1'b0 ;
  assign n27906 = n9959 | n27905 ;
  assign n27907 = ( n3169 & n9868 ) | ( n3169 & n22596 ) | ( n9868 & n22596 ) ;
  assign n27908 = ~n481 & n13999 ;
  assign n27909 = n27907 & n27908 ;
  assign n27910 = n16069 & ~n27909 ;
  assign n27911 = n27910 ^ n4615 ^ 1'b0 ;
  assign n27912 = ( n183 & ~n21608 ) | ( n183 & n27911 ) | ( ~n21608 & n27911 ) ;
  assign n27913 = ( ~n574 & n27906 ) | ( ~n574 & n27912 ) | ( n27906 & n27912 ) ;
  assign n27914 = n23156 & n23355 ;
  assign n27915 = ~n18167 & n23520 ;
  assign n27916 = ~n1887 & n27915 ;
  assign n27917 = n22558 & n24728 ;
  assign n27918 = n19262 & n24678 ;
  assign n27919 = ~n283 & n5815 ;
  assign n27920 = n3636 ^ n571 ^ 1'b0 ;
  assign n27921 = n27920 ^ n16909 ^ 1'b0 ;
  assign n27922 = ~n27919 & n27921 ;
  assign n27923 = n16744 | n25806 ;
  assign n27924 = n1111 & ~n2772 ;
  assign n27925 = n3990 & n27924 ;
  assign n27926 = n19995 ^ n5535 ^ 1'b0 ;
  assign n27927 = n633 | n27926 ;
  assign n27928 = n16612 ^ n374 ^ 1'b0 ;
  assign n27929 = n27927 | n27928 ;
  assign n27930 = n3257 | n19521 ;
  assign n27931 = n23292 & n27930 ;
  assign n27932 = ~n20279 & n27931 ;
  assign n27933 = n56 & n687 ;
  assign n27934 = n27932 & n27933 ;
  assign n27935 = ( n2568 & n12623 ) | ( n2568 & ~n25619 ) | ( n12623 & ~n25619 ) ;
  assign n27936 = ~n518 & n612 ;
  assign n27937 = ~n612 & n27936 ;
  assign n27938 = n5911 | n27937 ;
  assign n27939 = n27938 ^ n18573 ^ n6564 ;
  assign n27940 = ~n5811 & n26975 ;
  assign n27942 = n20679 ^ n14356 ^ 1'b0 ;
  assign n27943 = ~n11793 & n27942 ;
  assign n27941 = n12673 & ~n13730 ;
  assign n27944 = n27943 ^ n27941 ^ 1'b0 ;
  assign n27945 = n13028 & n27944 ;
  assign n27946 = n2469 ^ x1 ^ 1'b0 ;
  assign n27947 = n27946 ^ n7134 ^ 1'b0 ;
  assign n27948 = ~n17573 & n27947 ;
  assign n27949 = ~n20174 & n27525 ;
  assign n27950 = n4814 & n18307 ;
  assign n27951 = n27950 ^ n3652 ^ 1'b0 ;
  assign n27952 = n4379 ^ n3762 ^ 1'b0 ;
  assign n27953 = n5499 & n27952 ;
  assign n27954 = ~n8301 & n27953 ;
  assign n27955 = ~n2535 & n21111 ;
  assign n27956 = n24506 & n27955 ;
  assign n27957 = n9601 & n20308 ;
  assign n27958 = n15470 ^ n13258 ^ 1'b0 ;
  assign n27959 = ~n27957 & n27958 ;
  assign n27960 = n10345 ^ n4833 ^ 1'b0 ;
  assign n27961 = n9332 | n25041 ;
  assign n27962 = n6439 & ~n27961 ;
  assign n27963 = ~n2158 & n11682 ;
  assign n27964 = n27963 ^ n7159 ^ 1'b0 ;
  assign n27965 = n18665 ^ n445 ^ 1'b0 ;
  assign n27966 = n1933 & n7189 ;
  assign n27967 = n27966 ^ n2812 ^ 1'b0 ;
  assign n27968 = ~n13037 & n27967 ;
  assign n27969 = n27968 ^ n7656 ^ 1'b0 ;
  assign n27970 = n27965 & n27969 ;
  assign n27971 = n9536 ^ n7588 ^ 1'b0 ;
  assign n27972 = n21241 | n27971 ;
  assign n27973 = ~n4021 & n11023 ;
  assign n27974 = n15825 & ~n17610 ;
  assign n27975 = n27973 & n27974 ;
  assign n27976 = n26604 & n27975 ;
  assign n27977 = n8122 & ~n16423 ;
  assign n27979 = n4256 ^ n3349 ^ 1'b0 ;
  assign n27978 = n133 | n19409 ;
  assign n27980 = n27979 ^ n27978 ^ 1'b0 ;
  assign n27981 = n3683 & n27980 ;
  assign n27982 = ~n16132 & n27981 ;
  assign n27983 = n20403 ^ n9022 ^ 1'b0 ;
  assign n27984 = ~n1416 & n27983 ;
  assign n27985 = ( n540 & n1481 ) | ( n540 & n1771 ) | ( n1481 & n1771 ) ;
  assign n27986 = n27985 ^ n5647 ^ 1'b0 ;
  assign n27987 = ( n5005 & n10749 ) | ( n5005 & ~n27986 ) | ( n10749 & ~n27986 ) ;
  assign n27988 = ( n6330 & n7259 ) | ( n6330 & n7401 ) | ( n7259 & n7401 ) ;
  assign n27989 = n27988 ^ n49 ^ 1'b0 ;
  assign n27990 = n14686 | n15232 ;
  assign n27991 = n16627 & ~n27990 ;
  assign n27992 = n13355 & ~n18386 ;
  assign n27993 = n299 & n25022 ;
  assign n27994 = n19505 ^ n1495 ^ 1'b0 ;
  assign n27995 = n194 & n27994 ;
  assign n27998 = n1685 | n9478 ;
  assign n27999 = n27998 ^ n40 ^ 1'b0 ;
  assign n28000 = n22580 & n27999 ;
  assign n27996 = ( ~n1389 & n13826 ) | ( ~n1389 & n24680 ) | ( n13826 & n24680 ) ;
  assign n27997 = n9560 & ~n27996 ;
  assign n28001 = n28000 ^ n27997 ^ 1'b0 ;
  assign n28002 = n11527 & ~n19395 ;
  assign n28003 = n6355 & n28002 ;
  assign n28004 = n5756 & ~n28003 ;
  assign n28005 = n28004 ^ n14660 ^ 1'b0 ;
  assign n28017 = ( ~n522 & n2902 ) | ( ~n522 & n3544 ) | ( n2902 & n3544 ) ;
  assign n28014 = n864 | n7156 ;
  assign n28015 = n8086 | n28014 ;
  assign n28016 = n2974 & n28015 ;
  assign n28018 = n28017 ^ n28016 ^ 1'b0 ;
  assign n28010 = n4009 ^ n2549 ^ 1'b0 ;
  assign n28011 = n7552 & n28010 ;
  assign n28006 = n7368 | n7949 ;
  assign n28007 = n28006 ^ n7298 ^ 1'b0 ;
  assign n28008 = ~n13990 & n28007 ;
  assign n28009 = n28008 ^ n17294 ^ 1'b0 ;
  assign n28012 = n28011 ^ n28009 ^ 1'b0 ;
  assign n28013 = n7394 & ~n28012 ;
  assign n28019 = n28018 ^ n28013 ^ 1'b0 ;
  assign n28020 = n485 & ~n6971 ;
  assign n28021 = n6808 | n18068 ;
  assign n28022 = n18192 & ~n28021 ;
  assign n28023 = ~n12195 & n28022 ;
  assign n28024 = ~n8225 & n11176 ;
  assign n28025 = ~n5685 & n28024 ;
  assign n28026 = n14111 & n18711 ;
  assign n28027 = n5217 & ~n26835 ;
  assign n28028 = n6864 & n8978 ;
  assign n28029 = n28028 ^ n189 ^ 1'b0 ;
  assign n28030 = n28029 ^ n19645 ^ n1989 ;
  assign n28031 = n28030 ^ n10476 ^ 1'b0 ;
  assign n28032 = n1837 | n28031 ;
  assign n28034 = n1446 | n17737 ;
  assign n28033 = n588 | n19918 ;
  assign n28035 = n28034 ^ n28033 ^ 1'b0 ;
  assign n28036 = n12625 ^ n4291 ^ 1'b0 ;
  assign n28037 = n10505 | n28036 ;
  assign n28038 = ( n1884 & n2679 ) | ( n1884 & n6312 ) | ( n2679 & n6312 ) ;
  assign n28039 = n23286 | n28038 ;
  assign n28040 = n25264 ^ n21664 ^ 1'b0 ;
  assign n28041 = n15390 & ~n20142 ;
  assign n28042 = ~n135 & n5228 ;
  assign n28043 = n28042 ^ n17946 ^ 1'b0 ;
  assign n28044 = n22347 & n27485 ;
  assign n28045 = n28044 ^ n7836 ^ 1'b0 ;
  assign n28046 = n631 & n9224 ;
  assign n28047 = n28046 ^ n6179 ^ 1'b0 ;
  assign n28048 = n28047 ^ n105 ^ 1'b0 ;
  assign n28049 = ~n14190 & n19645 ;
  assign n28050 = n28049 ^ n18129 ^ 1'b0 ;
  assign n28051 = n22624 ^ n9958 ^ 1'b0 ;
  assign n28052 = n8208 ^ n493 ^ 1'b0 ;
  assign n28053 = ~n13299 & n28052 ;
  assign n28054 = n10858 & ~n28053 ;
  assign n28055 = n28051 & n28054 ;
  assign n28056 = n9270 ^ n7722 ^ 1'b0 ;
  assign n28057 = n2424 & ~n28056 ;
  assign n28058 = n9528 | n19062 ;
  assign n28059 = n28058 ^ n12380 ^ 1'b0 ;
  assign n28060 = n12219 & ~n19201 ;
  assign n28061 = ( n3300 & n14521 ) | ( n3300 & ~n28060 ) | ( n14521 & ~n28060 ) ;
  assign n28062 = ~n11451 & n26253 ;
  assign n28063 = ~n2989 & n6991 ;
  assign n28064 = n11683 ^ n9373 ^ 1'b0 ;
  assign n28065 = n9341 | n13946 ;
  assign n28066 = n12908 | n28065 ;
  assign n28067 = ~n7089 & n9309 ;
  assign n28068 = n28067 ^ n1955 ^ 1'b0 ;
  assign n28069 = n2423 | n16111 ;
  assign n28070 = n28069 ^ n1694 ^ 1'b0 ;
  assign n28071 = n28068 & ~n28070 ;
  assign n28072 = ~n19615 & n28071 ;
  assign n28073 = n2527 & n10166 ;
  assign n28074 = n6157 | n28073 ;
  assign n28075 = n28074 ^ n13618 ^ 1'b0 ;
  assign n28076 = n132 & ~n874 ;
  assign n28077 = n23154 & n28076 ;
  assign n28078 = n5085 | n11604 ;
  assign n28079 = n4665 | n28078 ;
  assign n28080 = n339 & ~n6119 ;
  assign n28081 = ~n28079 & n28080 ;
  assign n28082 = n2619 & ~n8474 ;
  assign n28083 = ~n5274 & n28082 ;
  assign n28084 = n28083 ^ n11052 ^ 1'b0 ;
  assign n28085 = n6238 & ~n28084 ;
  assign n28086 = n28085 ^ n13086 ^ 1'b0 ;
  assign n28087 = ~n7566 & n28086 ;
  assign n28088 = n28087 ^ n15582 ^ 1'b0 ;
  assign n28089 = n19421 ^ n9054 ^ 1'b0 ;
  assign n28090 = n3657 | n28089 ;
  assign n28091 = n28090 ^ n3880 ^ 1'b0 ;
  assign n28092 = n2146 & ~n28091 ;
  assign n28093 = ~n14289 & n28092 ;
  assign n28094 = n28093 ^ n9636 ^ 1'b0 ;
  assign n28095 = n9833 ^ n4250 ^ 1'b0 ;
  assign n28096 = n11211 | n28095 ;
  assign n28099 = ~n4297 & n5823 ;
  assign n28097 = n27398 ^ n8241 ^ 1'b0 ;
  assign n28098 = ( n16161 & ~n25434 ) | ( n16161 & n28097 ) | ( ~n25434 & n28097 ) ;
  assign n28100 = n28099 ^ n28098 ^ 1'b0 ;
  assign n28101 = n3521 | n4218 ;
  assign n28102 = n28101 ^ n10688 ^ 1'b0 ;
  assign n28103 = n12045 ^ n10841 ^ n10131 ;
  assign n28104 = n21904 & ~n28103 ;
  assign n28105 = n25615 ^ n17140 ^ 1'b0 ;
  assign n28106 = n28104 & n28105 ;
  assign n28107 = n4732 & n6907 ;
  assign n28108 = n28107 ^ n23632 ^ n12495 ;
  assign n28109 = n28108 ^ n18348 ^ 1'b0 ;
  assign n28110 = n7741 ^ n911 ^ 1'b0 ;
  assign n28111 = n1467 | n11359 ;
  assign n28112 = n28111 ^ n9049 ^ 1'b0 ;
  assign n28113 = n2451 | n26364 ;
  assign n28114 = n23356 ^ n6333 ^ 1'b0 ;
  assign n28115 = n21867 | n28114 ;
  assign n28116 = n5470 ^ n582 ^ 1'b0 ;
  assign n28117 = n2833 & ~n28116 ;
  assign n28118 = ( n8819 & n15850 ) | ( n8819 & ~n28117 ) | ( n15850 & ~n28117 ) ;
  assign n28119 = n28118 ^ n14997 ^ 1'b0 ;
  assign n28120 = n14559 ^ n1927 ^ 1'b0 ;
  assign n28121 = n28120 ^ n27515 ^ n13331 ;
  assign n28122 = n19040 ^ n17494 ^ 1'b0 ;
  assign n28123 = ~n23205 & n28122 ;
  assign n28124 = n28123 ^ n13386 ^ 1'b0 ;
  assign n28125 = n5228 & ~n10656 ;
  assign n28126 = n28125 ^ n26884 ^ n25160 ;
  assign n28127 = ~n1152 & n28126 ;
  assign n28128 = ~n15128 & n18706 ;
  assign n28129 = n4081 & ~n10311 ;
  assign n28130 = n28129 ^ n3349 ^ 1'b0 ;
  assign n28131 = n28130 ^ n20803 ^ n16604 ;
  assign n28132 = n16532 & ~n21769 ;
  assign n28133 = n2798 | n18456 ;
  assign n28134 = n28133 ^ n18549 ^ 1'b0 ;
  assign n28135 = n16455 | n22394 ;
  assign n28136 = n430 & ~n659 ;
  assign n28137 = n28136 ^ n208 ^ 1'b0 ;
  assign n28138 = n28137 ^ n15630 ^ n14563 ;
  assign n28139 = n7835 & ~n12575 ;
  assign n28140 = ~n21523 & n28139 ;
  assign n28141 = ~n28138 & n28140 ;
  assign n28142 = n19428 ^ n11710 ^ 1'b0 ;
  assign n28143 = ~n13304 & n28142 ;
  assign n28144 = n28003 | n28143 ;
  assign n28145 = n15283 ^ n6885 ^ 1'b0 ;
  assign n28146 = n11560 ^ n9564 ^ n5541 ;
  assign n28147 = n28146 ^ n13050 ^ 1'b0 ;
  assign n28148 = n25968 ^ n12695 ^ n3110 ;
  assign n28149 = n28147 & ~n28148 ;
  assign n28150 = n3828 & ~n28149 ;
  assign n28151 = n2094 & n10134 ;
  assign n28152 = n1202 | n21266 ;
  assign n28153 = n25665 & ~n28152 ;
  assign n28154 = n411 | n18382 ;
  assign n28155 = n4871 | n28154 ;
  assign n28156 = n8674 ^ n4326 ^ 1'b0 ;
  assign n28157 = n2513 | n28156 ;
  assign n28158 = n28155 & ~n28157 ;
  assign n28159 = n28158 ^ n7078 ^ 1'b0 ;
  assign n28160 = n6662 | n9358 ;
  assign n28163 = n8279 ^ n7935 ^ 1'b0 ;
  assign n28162 = n3301 | n7077 ;
  assign n28161 = n2981 | n24442 ;
  assign n28164 = n28163 ^ n28162 ^ n28161 ;
  assign n28165 = n3622 | n6294 ;
  assign n28166 = n28165 ^ n24214 ^ 1'b0 ;
  assign n28171 = n727 | n16144 ;
  assign n28167 = n11614 | n19534 ;
  assign n28168 = n4449 & ~n28167 ;
  assign n28169 = n12865 ^ n1796 ^ 1'b0 ;
  assign n28170 = n28168 | n28169 ;
  assign n28172 = n28171 ^ n28170 ^ 1'b0 ;
  assign n28173 = n22653 & n28172 ;
  assign n28174 = ~n11167 & n13179 ;
  assign n28175 = ( ~n3258 & n10277 ) | ( ~n3258 & n28174 ) | ( n10277 & n28174 ) ;
  assign n28176 = n13848 & ~n18830 ;
  assign n28177 = n28176 ^ n22029 ^ 1'b0 ;
  assign n28178 = n21485 & n21798 ;
  assign n28179 = n28178 ^ n14489 ^ 1'b0 ;
  assign n28181 = n7080 ^ n7019 ^ 1'b0 ;
  assign n28180 = n20305 | n25606 ;
  assign n28182 = n28181 ^ n28180 ^ 1'b0 ;
  assign n28183 = n103 | n3073 ;
  assign n28184 = n15863 & n28183 ;
  assign n28185 = n28184 ^ n26121 ^ 1'b0 ;
  assign n28186 = n12952 | n15975 ;
  assign n28187 = n28186 ^ n19338 ^ 1'b0 ;
  assign n28188 = ~n2871 & n18034 ;
  assign n28189 = n26425 ^ n1023 ^ 1'b0 ;
  assign n28190 = n7532 | n28189 ;
  assign n28191 = n19526 ^ n13306 ^ 1'b0 ;
  assign n28192 = n7140 | n28191 ;
  assign n28193 = n4213 & ~n27740 ;
  assign n28194 = ~n3428 & n13422 ;
  assign n28195 = n2648 | n9963 ;
  assign n28196 = n15341 & ~n28195 ;
  assign n28197 = n28196 ^ n19158 ^ 1'b0 ;
  assign n28198 = n28194 & ~n28197 ;
  assign n28199 = ~n593 & n3890 ;
  assign n28200 = ~n10836 & n28199 ;
  assign n28201 = n27469 ^ n5872 ^ n4401 ;
  assign n28202 = ~n6479 & n21404 ;
  assign n28203 = ~n11722 & n28202 ;
  assign n28204 = ( ~n6040 & n10357 ) | ( ~n6040 & n21889 ) | ( n10357 & n21889 ) ;
  assign n28205 = n23797 ^ n9151 ^ 1'b0 ;
  assign n28210 = n13557 ^ n5254 ^ 1'b0 ;
  assign n28206 = n770 | n16155 ;
  assign n28207 = n4976 & ~n28206 ;
  assign n28208 = ( n1464 & ~n7574 ) | ( n1464 & n28207 ) | ( ~n7574 & n28207 ) ;
  assign n28209 = n2172 | n28208 ;
  assign n28211 = n28210 ^ n28209 ^ 1'b0 ;
  assign n28212 = n1552 & n17115 ;
  assign n28213 = ~n17709 & n28212 ;
  assign n28214 = n21398 | n28213 ;
  assign n28215 = n28214 ^ n16415 ^ 1'b0 ;
  assign n28216 = n1897 | n21812 ;
  assign n28217 = n28215 & ~n28216 ;
  assign n28218 = ~n367 & n2128 ;
  assign n28219 = n22370 & n28218 ;
  assign n28220 = n135 & n12058 ;
  assign n28221 = ~n1419 & n9368 ;
  assign n28222 = n16734 & ~n28221 ;
  assign n28223 = n13012 & n22040 ;
  assign n28224 = ~n17 & n28223 ;
  assign n28225 = n2746 ^ n2030 ^ 1'b0 ;
  assign n28226 = n1277 | n28225 ;
  assign n28227 = n5467 | n28226 ;
  assign n28231 = ~n4282 & n14693 ;
  assign n28232 = n28231 ^ n8724 ^ 1'b0 ;
  assign n28228 = n16389 ^ n4643 ^ 1'b0 ;
  assign n28229 = n25208 & ~n28228 ;
  assign n28230 = n28229 ^ n7880 ^ 1'b0 ;
  assign n28233 = n28232 ^ n28230 ^ n26922 ;
  assign n28234 = n5999 & ~n21531 ;
  assign n28235 = n28234 ^ n65 ^ 1'b0 ;
  assign n28236 = n28235 ^ n5499 ^ 1'b0 ;
  assign n28237 = ~n318 & n24084 ;
  assign n28238 = n7254 | n10875 ;
  assign n28239 = n28237 & ~n28238 ;
  assign n28240 = n13331 ^ n12458 ^ 1'b0 ;
  assign n28241 = n7204 | n28240 ;
  assign n28242 = ~n1852 & n4701 ;
  assign n28243 = n28242 ^ n8186 ^ 1'b0 ;
  assign n28244 = n28241 | n28243 ;
  assign n28245 = n20158 ^ n14024 ^ n2060 ;
  assign n28246 = ~n28244 & n28245 ;
  assign n28247 = n4863 & n14977 ;
  assign n28248 = n28247 ^ n4364 ^ 1'b0 ;
  assign n28249 = n14388 & n28248 ;
  assign n28250 = n17704 & ~n26963 ;
  assign n28251 = n28250 ^ n17088 ^ 1'b0 ;
  assign n28252 = n28251 ^ n5172 ^ 1'b0 ;
  assign n28253 = ~n28249 & n28252 ;
  assign n28254 = n7023 & ~n18950 ;
  assign n28255 = n14958 ^ n3758 ^ 1'b0 ;
  assign n28256 = n23893 ^ n15992 ^ n712 ;
  assign n28257 = ~n28255 & n28256 ;
  assign n28258 = ~n28254 & n28257 ;
  assign n28260 = n202 & n16144 ;
  assign n28259 = ~n5865 & n6235 ;
  assign n28261 = n28260 ^ n28259 ^ n17418 ;
  assign n28262 = n28261 ^ n6596 ^ 1'b0 ;
  assign n28263 = ( n7062 & ~n15119 ) | ( n7062 & n25881 ) | ( ~n15119 & n25881 ) ;
  assign n28264 = n4637 & ~n28263 ;
  assign n28265 = n28264 ^ n7998 ^ 1'b0 ;
  assign n28266 = ~n7206 & n26622 ;
  assign n28267 = n28266 ^ n4690 ^ 1'b0 ;
  assign n28268 = n10719 & n20614 ;
  assign n28269 = n12671 | n18519 ;
  assign n28270 = n28269 ^ n20719 ^ 1'b0 ;
  assign n28271 = n67 | n18535 ;
  assign n28272 = n9831 & ~n28271 ;
  assign n28273 = n28272 ^ n12854 ^ n10789 ;
  assign n28274 = ~n7867 & n9955 ;
  assign n28275 = n28273 & n28274 ;
  assign n28276 = n28275 ^ n19438 ^ n2192 ;
  assign n28277 = n5059 & ~n7784 ;
  assign n28278 = n5525 & ~n8131 ;
  assign n28279 = n19695 ^ n14904 ^ 1'b0 ;
  assign n28280 = ~n28278 & n28279 ;
  assign n28281 = ~n7718 & n7756 ;
  assign n28282 = n10239 | n19750 ;
  assign n28283 = n28282 ^ n922 ^ 1'b0 ;
  assign n28284 = n3429 & ~n11675 ;
  assign n28285 = n28284 ^ n4005 ^ 1'b0 ;
  assign n28286 = n8367 & ~n27851 ;
  assign n28287 = ~n26533 & n28286 ;
  assign n28288 = n2577 | n21623 ;
  assign n28290 = n7792 & ~n9468 ;
  assign n28291 = n28290 ^ n22024 ^ 1'b0 ;
  assign n28289 = n7960 | n8889 ;
  assign n28292 = n28291 ^ n28289 ^ 1'b0 ;
  assign n28293 = n2701 | n4097 ;
  assign n28295 = n12202 ^ n10259 ^ 1'b0 ;
  assign n28294 = n4106 ^ n3797 ^ 1'b0 ;
  assign n28296 = n28295 ^ n28294 ^ n22622 ;
  assign n28297 = n28296 ^ n8950 ^ 1'b0 ;
  assign n28298 = ~n28293 & n28297 ;
  assign n28299 = n12504 ^ n9031 ^ 1'b0 ;
  assign n28300 = n17254 & n25586 ;
  assign n28301 = n28300 ^ n2417 ^ 1'b0 ;
  assign n28302 = n28301 ^ n3612 ^ 1'b0 ;
  assign n28303 = n13465 ^ n2004 ^ 1'b0 ;
  assign n28304 = n5136 & n28303 ;
  assign n28305 = ~n28302 & n28304 ;
  assign n28306 = ~n19965 & n25157 ;
  assign n28307 = ~n1430 & n28306 ;
  assign n28308 = ~n17629 & n28307 ;
  assign n28309 = n11778 ^ n2294 ^ 1'b0 ;
  assign n28310 = n14240 & n28309 ;
  assign n28311 = n28310 ^ n2941 ^ 1'b0 ;
  assign n28312 = ( n439 & n11759 ) | ( n439 & ~n15145 ) | ( n11759 & ~n15145 ) ;
  assign n28313 = ~n28311 & n28312 ;
  assign n28314 = ~n13321 & n28313 ;
  assign n28315 = n15313 & n19651 ;
  assign n28316 = n5686 | n18797 ;
  assign n28317 = n28315 | n28316 ;
  assign n28318 = n13699 ^ n1213 ^ 1'b0 ;
  assign n28319 = n27622 ^ n3731 ^ 1'b0 ;
  assign n28320 = n28318 | n28319 ;
  assign n28321 = ( n5535 & n8531 ) | ( n5535 & n21791 ) | ( n8531 & n21791 ) ;
  assign n28322 = ~n2452 & n15728 ;
  assign n28323 = n28322 ^ n15140 ^ 1'b0 ;
  assign n28324 = n28323 ^ n8980 ^ 1'b0 ;
  assign n28325 = ( n9050 & n10270 ) | ( n9050 & ~n22013 ) | ( n10270 & ~n22013 ) ;
  assign n28326 = n996 & n1688 ;
  assign n28327 = n28326 ^ n25449 ^ 1'b0 ;
  assign n28328 = ~n7825 & n10031 ;
  assign n28329 = n28328 ^ n6514 ^ 1'b0 ;
  assign n28330 = n14666 & ~n20310 ;
  assign n28331 = n8549 & n28330 ;
  assign n28332 = n21249 ^ n13355 ^ 1'b0 ;
  assign n28333 = ~n8939 & n16636 ;
  assign n28334 = n15887 & n28333 ;
  assign n28335 = ~n26137 & n28334 ;
  assign n28340 = n3058 & n8432 ;
  assign n28337 = n5958 | n19647 ;
  assign n28338 = n28337 ^ n8128 ^ 1'b0 ;
  assign n28336 = ~n6553 & n6756 ;
  assign n28339 = n28338 ^ n28336 ^ 1'b0 ;
  assign n28341 = n28340 ^ n28339 ^ n4131 ;
  assign n28343 = n3820 | n3996 ;
  assign n28344 = n10844 | n28343 ;
  assign n28345 = ( n4360 & ~n7679 ) | ( n4360 & n28344 ) | ( ~n7679 & n28344 ) ;
  assign n28342 = n5151 & ~n9670 ;
  assign n28346 = n28345 ^ n28342 ^ 1'b0 ;
  assign n28347 = n6305 & n28346 ;
  assign n28348 = ( n738 & n2176 ) | ( n738 & ~n8577 ) | ( n2176 & ~n8577 ) ;
  assign n28349 = n19014 ^ n2045 ^ 1'b0 ;
  assign n28350 = n28349 ^ n17229 ^ 1'b0 ;
  assign n28351 = ( n2093 & n28348 ) | ( n2093 & ~n28350 ) | ( n28348 & ~n28350 ) ;
  assign n28352 = n6201 ^ n1580 ^ 1'b0 ;
  assign n28353 = n3127 | n23335 ;
  assign n28354 = n28353 ^ n20262 ^ 1'b0 ;
  assign n28355 = ( ~n1182 & n28352 ) | ( ~n1182 & n28354 ) | ( n28352 & n28354 ) ;
  assign n28362 = n20281 ^ n17931 ^ 1'b0 ;
  assign n28356 = n7889 | n12673 ;
  assign n28357 = n4300 | n28356 ;
  assign n28358 = n28357 ^ n10904 ^ 1'b0 ;
  assign n28359 = n6464 ^ n6196 ^ 1'b0 ;
  assign n28360 = n22125 & n28359 ;
  assign n28361 = n28358 & n28360 ;
  assign n28363 = n28362 ^ n28361 ^ 1'b0 ;
  assign n28364 = n3749 & ~n8128 ;
  assign n28365 = n28364 ^ n21444 ^ 1'b0 ;
  assign n28366 = n28365 ^ n5796 ^ 1'b0 ;
  assign n28367 = n14586 | n20341 ;
  assign n28368 = n25919 ^ n1295 ^ 1'b0 ;
  assign n28369 = n28368 ^ n27196 ^ n2193 ;
  assign n28370 = ( n3298 & n4563 ) | ( n3298 & ~n5154 ) | ( n4563 & ~n5154 ) ;
  assign n28371 = ~n10112 & n11194 ;
  assign n28372 = n2726 & n28371 ;
  assign n28373 = n15000 & ~n28372 ;
  assign n28374 = n9238 ^ n8672 ^ 1'b0 ;
  assign n28375 = ~n11329 & n28374 ;
  assign n28376 = n9182 & n28375 ;
  assign n28377 = n28376 ^ n10145 ^ 1'b0 ;
  assign n28378 = n7182 & n8944 ;
  assign n28379 = n28378 ^ n26223 ^ 1'b0 ;
  assign n28380 = ~n873 & n4709 ;
  assign n28381 = ( n3282 & ~n6161 ) | ( n3282 & n28380 ) | ( ~n6161 & n28380 ) ;
  assign n28382 = n28381 ^ n6662 ^ 1'b0 ;
  assign n28383 = n17577 | n28382 ;
  assign n28384 = ~n3901 & n6613 ;
  assign n28385 = n16512 & n28384 ;
  assign n28386 = n28383 & n28385 ;
  assign n28387 = n26630 ^ n3489 ^ 1'b0 ;
  assign n28388 = n9598 ^ n5692 ^ 1'b0 ;
  assign n28389 = ~n9332 & n28388 ;
  assign n28390 = n1208 | n28389 ;
  assign n28391 = n27524 ^ n13797 ^ 1'b0 ;
  assign n28392 = n23761 & ~n28391 ;
  assign n28393 = n20657 ^ n11509 ^ 1'b0 ;
  assign n28394 = n3913 | n4328 ;
  assign n28395 = n28394 ^ n5054 ^ 1'b0 ;
  assign n28396 = ~n18956 & n28395 ;
  assign n28397 = n28396 ^ n23155 ^ 1'b0 ;
  assign n28398 = n2093 ^ n224 ^ 1'b0 ;
  assign n28399 = n25613 & n28398 ;
  assign n28400 = n28399 ^ n494 ^ 1'b0 ;
  assign n28401 = n21436 ^ n10480 ^ n4559 ;
  assign n28402 = n28401 ^ n12721 ^ 1'b0 ;
  assign n28403 = n28400 & n28402 ;
  assign n28404 = n28403 ^ n25373 ^ 1'b0 ;
  assign n28405 = n6563 & ~n28404 ;
  assign n28406 = ( ~n2588 & n6221 ) | ( ~n2588 & n10235 ) | ( n6221 & n10235 ) ;
  assign n28407 = n16040 & ~n28406 ;
  assign n28408 = ( n1770 & n7471 ) | ( n1770 & ~n28407 ) | ( n7471 & ~n28407 ) ;
  assign n28409 = n453 & ~n15641 ;
  assign n28410 = n28409 ^ n15952 ^ 1'b0 ;
  assign n28411 = n5206 | n15922 ;
  assign n28412 = n22360 | n28411 ;
  assign n28413 = n765 | n4709 ;
  assign n28414 = ~n2324 & n28413 ;
  assign n28415 = ( n7086 & n13891 ) | ( n7086 & ~n16356 ) | ( n13891 & ~n16356 ) ;
  assign n28416 = ~n9037 & n28415 ;
  assign n28417 = n5646 & n28416 ;
  assign n28418 = n28417 ^ n1439 ^ 1'b0 ;
  assign n28419 = ~n3037 & n18856 ;
  assign n28420 = n578 & n13169 ;
  assign n28421 = n11621 & n28420 ;
  assign n28422 = n9309 ^ n4888 ^ 1'b0 ;
  assign n28423 = ~n28421 & n28422 ;
  assign n28424 = n5364 ^ n1607 ^ 1'b0 ;
  assign n28425 = n751 | n10295 ;
  assign n28426 = ~n23566 & n27874 ;
  assign n28427 = n28426 ^ n16460 ^ 1'b0 ;
  assign n28428 = n14708 ^ n7633 ^ n1460 ;
  assign n28429 = ~n6610 & n28428 ;
  assign n28430 = n25047 ^ n4687 ^ 1'b0 ;
  assign n28431 = ~n657 & n28430 ;
  assign n28432 = n3464 | n4024 ;
  assign n28433 = n28432 ^ n10747 ^ 1'b0 ;
  assign n28434 = n6045 ^ n522 ^ 1'b0 ;
  assign n28435 = n8118 & n16015 ;
  assign n28436 = n4436 & n28435 ;
  assign n28437 = n12573 & n28436 ;
  assign n28438 = n28437 ^ n14248 ^ 1'b0 ;
  assign n28439 = ~n6099 & n28438 ;
  assign n28440 = ~n24438 & n28439 ;
  assign n28441 = n15548 ^ n6891 ^ 1'b0 ;
  assign n28442 = ~n20234 & n28441 ;
  assign n28443 = n22083 ^ n3030 ^ 1'b0 ;
  assign n28444 = ( n2815 & n11638 ) | ( n2815 & n19512 ) | ( n11638 & n19512 ) ;
  assign n28445 = n25218 ^ n10231 ^ 1'b0 ;
  assign n28446 = n23209 ^ n3761 ^ 1'b0 ;
  assign n28447 = n7299 & ~n28446 ;
  assign n28448 = n1251 & ~n2356 ;
  assign n28449 = n12430 & n28448 ;
  assign n28450 = ~n6069 & n28449 ;
  assign n28451 = n28450 ^ n16968 ^ 1'b0 ;
  assign n28452 = n4075 & ~n25565 ;
  assign n28453 = n28452 ^ n13117 ^ 1'b0 ;
  assign n28454 = ~n437 & n28453 ;
  assign n28455 = n17701 ^ n5535 ^ n3536 ;
  assign n28457 = n12265 | n23202 ;
  assign n28458 = n28457 ^ n4991 ^ 1'b0 ;
  assign n28459 = n16227 | n28458 ;
  assign n28456 = n9714 ^ n4685 ^ 1'b0 ;
  assign n28460 = n28459 ^ n28456 ^ 1'b0 ;
  assign n28461 = n21803 | n27281 ;
  assign n28462 = n2556 ^ n1400 ^ 1'b0 ;
  assign n28463 = n498 & ~n28462 ;
  assign n28464 = n1396 | n9753 ;
  assign n28465 = n9753 & ~n28464 ;
  assign n28466 = n9464 & ~n28465 ;
  assign n28467 = n28465 & n28466 ;
  assign n28468 = n28467 ^ n2933 ^ 1'b0 ;
  assign n28469 = n2240 | n28468 ;
  assign n28470 = n28463 | n28469 ;
  assign n28471 = ~n6179 & n10359 ;
  assign n28472 = n28471 ^ n10500 ^ 1'b0 ;
  assign n28473 = n14773 & n28472 ;
  assign n28474 = ( n3701 & n8230 ) | ( n3701 & n28473 ) | ( n8230 & n28473 ) ;
  assign n28475 = ~n22020 & n28342 ;
  assign n28476 = n3264 & n9106 ;
  assign n28477 = n28476 ^ n11754 ^ 1'b0 ;
  assign n28478 = n18766 & n28477 ;
  assign n28479 = n10839 ^ n1637 ^ 1'b0 ;
  assign n28480 = n9153 & ~n28479 ;
  assign n28481 = n4432 & ~n5866 ;
  assign n28482 = n13513 & ~n28481 ;
  assign n28483 = n14558 ^ n2330 ^ 1'b0 ;
  assign n28484 = n15671 & ~n28483 ;
  assign n28485 = ~n9292 & n19372 ;
  assign n28486 = n9546 ^ n6818 ^ 1'b0 ;
  assign n28487 = ~n12272 & n28486 ;
  assign n28488 = ~n809 & n10134 ;
  assign n28489 = n13843 | n23806 ;
  assign n28490 = n28489 ^ n19193 ^ 1'b0 ;
  assign n28491 = n28490 ^ n24500 ^ 1'b0 ;
  assign n28492 = n27555 ^ n22215 ^ n2876 ;
  assign n28493 = n12634 ^ n6122 ^ 1'b0 ;
  assign n28494 = n8068 & ~n14667 ;
  assign n28495 = n28494 ^ n2181 ^ 1'b0 ;
  assign n28496 = ~n28493 & n28495 ;
  assign n28497 = n10695 ^ n1740 ^ 1'b0 ;
  assign n28498 = n1987 | n28497 ;
  assign n28501 = n25938 ^ n16833 ^ n6927 ;
  assign n28499 = n368 & ~n6006 ;
  assign n28500 = n9319 | n28499 ;
  assign n28502 = n28501 ^ n28500 ^ 1'b0 ;
  assign n28503 = n5724 | n11486 ;
  assign n28504 = n12011 | n13130 ;
  assign n28505 = n28504 ^ n911 ^ n31 ;
  assign n28506 = ~n3566 & n8879 ;
  assign n28507 = n16401 & n20460 ;
  assign n28508 = n13771 & n28507 ;
  assign n28509 = n4084 & n16094 ;
  assign n28510 = n15454 ^ n15452 ^ n9692 ;
  assign n28511 = n9163 & ~n28510 ;
  assign n28512 = n9752 & n28511 ;
  assign n28513 = ~n8093 & n28512 ;
  assign n28514 = n209 & ~n28513 ;
  assign n28515 = ~n28509 & n28514 ;
  assign n28516 = n26348 ^ n4326 ^ 1'b0 ;
  assign n28518 = n241 & n2721 ;
  assign n28519 = n28518 ^ n18908 ^ 1'b0 ;
  assign n28520 = n28519 ^ n7506 ^ 1'b0 ;
  assign n28517 = n5244 & n11458 ;
  assign n28521 = n28520 ^ n28517 ^ 1'b0 ;
  assign n28522 = n7578 ^ n1570 ^ 1'b0 ;
  assign n28523 = n19218 ^ n1318 ^ 1'b0 ;
  assign n28524 = n28522 | n28523 ;
  assign n28525 = n28183 ^ n3226 ^ 1'b0 ;
  assign n28526 = n1984 & n9012 ;
  assign n28527 = n4707 ^ n466 ^ 1'b0 ;
  assign n28528 = n1460 & ~n16077 ;
  assign n28529 = n5005 | n26350 ;
  assign n28531 = n12062 ^ n2552 ^ 1'b0 ;
  assign n28532 = n439 & ~n28531 ;
  assign n28530 = n8684 | n17313 ;
  assign n28533 = n28532 ^ n28530 ^ 1'b0 ;
  assign n28534 = n25387 & ~n28533 ;
  assign n28535 = n3907 & n9258 ;
  assign n28536 = n19924 ^ n6387 ^ 1'b0 ;
  assign n28537 = ~n28535 & n28536 ;
  assign n28540 = n5806 ^ n541 ^ 1'b0 ;
  assign n28538 = n1123 & ~n5357 ;
  assign n28539 = ~n19609 & n28538 ;
  assign n28541 = n28540 ^ n28539 ^ 1'b0 ;
  assign n28542 = n21493 & n28541 ;
  assign n28543 = ~n9544 & n19062 ;
  assign n28544 = n28543 ^ n1806 ^ 1'b0 ;
  assign n28545 = n11489 ^ n8000 ^ 1'b0 ;
  assign n28546 = n28544 & n28545 ;
  assign n28547 = n14778 ^ n2435 ^ 1'b0 ;
  assign n28548 = n28547 ^ n21623 ^ 1'b0 ;
  assign n28549 = n7494 & n28548 ;
  assign n28550 = n3331 | n28549 ;
  assign n28551 = n682 | n15059 ;
  assign n28552 = n21883 | n28551 ;
  assign n28553 = n20335 ^ n1897 ^ 1'b0 ;
  assign n28554 = n1010 | n9548 ;
  assign n28555 = ~n6986 & n28554 ;
  assign n28556 = ~n10501 & n28555 ;
  assign n28557 = n20764 | n28556 ;
  assign n28558 = n421 & ~n10624 ;
  assign n28559 = n5113 & n22785 ;
  assign n28560 = ~n3366 & n5549 ;
  assign n28561 = n2700 & n25584 ;
  assign n28562 = n20406 & n28561 ;
  assign n28563 = ~n9526 & n10688 ;
  assign n28564 = n12993 ^ n9319 ^ 1'b0 ;
  assign n28565 = n20530 ^ n3359 ^ 1'b0 ;
  assign n28566 = n2688 & n22354 ;
  assign n28567 = n28566 ^ n2000 ^ 1'b0 ;
  assign n28568 = n6157 & ~n25717 ;
  assign n28569 = ~n6157 & n28568 ;
  assign n28570 = n637 & ~n11852 ;
  assign n28571 = n11852 & n28570 ;
  assign n28572 = n5558 & ~n28571 ;
  assign n28573 = n28571 & n28572 ;
  assign n28574 = n28569 | n28573 ;
  assign n28575 = n28574 ^ n13452 ^ n5800 ;
  assign n28576 = n7482 & n22826 ;
  assign n28577 = n3827 & n28576 ;
  assign n28578 = n23226 ^ n4750 ^ 1'b0 ;
  assign n28579 = ~n18984 & n28578 ;
  assign n28580 = n26837 ^ n3762 ^ 1'b0 ;
  assign n28581 = ~n28579 & n28580 ;
  assign n28582 = n8222 & ~n10845 ;
  assign n28583 = n2595 & n6099 ;
  assign n28584 = n3289 & n28583 ;
  assign n28585 = n5933 & n8154 ;
  assign n28586 = n3488 & ~n9806 ;
  assign n28587 = n28586 ^ n22292 ^ 1'b0 ;
  assign n28588 = n12578 ^ n3924 ^ 1'b0 ;
  assign n28589 = n8631 & ~n17492 ;
  assign n28590 = n18813 & ~n28589 ;
  assign n28591 = ~n28588 & n28590 ;
  assign n28592 = n11118 ^ n6176 ^ n2765 ;
  assign n28593 = n7500 | n28592 ;
  assign n28594 = ~n2427 & n6151 ;
  assign n28595 = n25275 ^ n17418 ^ 1'b0 ;
  assign n28596 = n28594 | n28595 ;
  assign n28597 = ~n10283 & n11295 ;
  assign n28598 = n470 & n28597 ;
  assign n28599 = n2101 & n28598 ;
  assign n28600 = n8952 & ~n15484 ;
  assign n28601 = ~n194 & n28600 ;
  assign n28602 = n28601 ^ n25028 ^ 1'b0 ;
  assign n28603 = ~n6155 & n21836 ;
  assign n28604 = n28603 ^ n8208 ^ 1'b0 ;
  assign n28606 = ~n2588 & n4105 ;
  assign n28605 = n9411 ^ n3853 ^ 1'b0 ;
  assign n28607 = n28606 ^ n28605 ^ 1'b0 ;
  assign n28608 = ~n3972 & n28607 ;
  assign n28609 = ~n1109 & n28608 ;
  assign n28610 = n2453 | n3508 ;
  assign n28611 = n9787 & ~n28610 ;
  assign n28612 = ~n8176 & n12123 ;
  assign n28613 = n2955 & n16603 ;
  assign n28614 = n8595 & n12894 ;
  assign n28615 = n14031 ^ n1464 ^ 1'b0 ;
  assign n28616 = n6099 & n28615 ;
  assign n28617 = n582 & n28616 ;
  assign n28618 = n28617 ^ n6099 ^ 1'b0 ;
  assign n28619 = n3687 | n28618 ;
  assign n28620 = n2660 & ~n24874 ;
  assign n28621 = n22306 ^ n864 ^ n612 ;
  assign n28622 = n15363 & ~n28621 ;
  assign n28623 = ~n9105 & n18383 ;
  assign n28624 = ~n13293 & n28623 ;
  assign n28625 = ~n5619 & n23560 ;
  assign n28626 = n28625 ^ n6119 ^ 1'b0 ;
  assign n28627 = n8354 & ~n8607 ;
  assign n28628 = ~n15680 & n28627 ;
  assign n28630 = n5911 | n9443 ;
  assign n28631 = n28630 ^ n13354 ^ 1'b0 ;
  assign n28629 = n16221 & ~n25114 ;
  assign n28632 = n28631 ^ n28629 ^ 1'b0 ;
  assign n28633 = ( n17399 & n21291 ) | ( n17399 & ~n26622 ) | ( n21291 & ~n26622 ) ;
  assign n28634 = n12705 & ~n21243 ;
  assign n28635 = ~n11217 & n17964 ;
  assign n28636 = n28635 ^ n13621 ^ 1'b0 ;
  assign n28637 = n5227 & ~n13298 ;
  assign n28638 = n18046 | n28637 ;
  assign n28639 = n28638 ^ n11694 ^ 1'b0 ;
  assign n28640 = n21961 | n26229 ;
  assign n28641 = n8154 ^ n4860 ^ n3004 ;
  assign n28642 = n823 & ~n3094 ;
  assign n28643 = n28642 ^ n12902 ^ 1'b0 ;
  assign n28644 = n28641 & n28643 ;
  assign n28645 = n3091 & ~n13390 ;
  assign n28646 = n3136 & n5646 ;
  assign n28647 = ~n3136 & n28646 ;
  assign n28648 = ~n5900 & n23274 ;
  assign n28649 = n2265 | n28648 ;
  assign n28650 = n28648 & ~n28649 ;
  assign n28651 = n28647 & ~n28650 ;
  assign n28652 = n1609 & ~n10652 ;
  assign n28653 = n15295 & ~n28652 ;
  assign n28654 = n28651 & n28653 ;
  assign n28655 = n10925 | n28654 ;
  assign n28656 = n10925 & ~n28655 ;
  assign n28657 = n233 & ~n1972 ;
  assign n28658 = ~n233 & n28657 ;
  assign n28659 = n4368 | n28658 ;
  assign n28660 = ~n127 & n14701 ;
  assign n28661 = n17008 ^ n10642 ^ 1'b0 ;
  assign n28662 = n28660 & n28661 ;
  assign n28663 = ~n21040 & n28662 ;
  assign n28664 = n28659 & n28663 ;
  assign n28665 = n28656 | n28664 ;
  assign n28666 = n249 | n28665 ;
  assign n28667 = n2048 | n20936 ;
  assign n28668 = n8341 ^ n5469 ^ 1'b0 ;
  assign n28669 = n2007 & ~n7808 ;
  assign n28670 = n28669 ^ n18906 ^ 1'b0 ;
  assign n28671 = n28670 ^ n13661 ^ 1'b0 ;
  assign n28672 = n28668 & n28671 ;
  assign n28673 = n6385 & n28672 ;
  assign n28674 = n28673 ^ n14888 ^ 1'b0 ;
  assign n28675 = n2147 & ~n5268 ;
  assign n28676 = n28675 ^ n25215 ^ n23649 ;
  assign n28677 = n6540 & ~n12156 ;
  assign n28678 = n28677 ^ n19463 ^ 1'b0 ;
  assign n28679 = n25104 ^ n20662 ^ 1'b0 ;
  assign n28680 = n28678 | n28679 ;
  assign n28681 = n13157 ^ n6669 ^ 1'b0 ;
  assign n28682 = n14691 & ~n23133 ;
  assign n28683 = n28682 ^ n5786 ^ 1'b0 ;
  assign n28684 = n28683 ^ n28610 ^ 1'b0 ;
  assign n28685 = n28681 & n28684 ;
  assign n28686 = n4785 ^ n170 ^ 1'b0 ;
  assign n28687 = n16719 | n28686 ;
  assign n28688 = n12449 ^ n1124 ^ 1'b0 ;
  assign n28689 = n15109 & n28688 ;
  assign n28690 = n28687 & n28689 ;
  assign n28691 = n1896 & n15600 ;
  assign n28692 = n4241 & n7763 ;
  assign n28693 = n12680 ^ n3193 ^ 1'b0 ;
  assign n28694 = ~n28692 & n28693 ;
  assign n28695 = n28691 | n28694 ;
  assign n28696 = ( n2919 & ~n9985 ) | ( n2919 & n28695 ) | ( ~n9985 & n28695 ) ;
  assign n28697 = ( ~n16725 & n21564 ) | ( ~n16725 & n28696 ) | ( n21564 & n28696 ) ;
  assign n28698 = ~n3716 & n14010 ;
  assign n28699 = n13809 | n28698 ;
  assign n28700 = n21635 ^ n11865 ^ 1'b0 ;
  assign n28701 = n11743 ^ n8277 ^ 1'b0 ;
  assign n28702 = n6026 & ~n28701 ;
  assign n28703 = n28702 ^ n10687 ^ 1'b0 ;
  assign n28704 = ~n19178 & n24181 ;
  assign n28705 = n4191 & ~n10463 ;
  assign n28706 = n28705 ^ n5748 ^ 1'b0 ;
  assign n28707 = n12400 ^ n1466 ^ 1'b0 ;
  assign n28708 = n18591 | n28707 ;
  assign n28712 = n25519 ^ n16600 ^ n105 ;
  assign n28709 = n14238 ^ n269 ^ 1'b0 ;
  assign n28710 = n28709 ^ n10545 ^ n8896 ;
  assign n28711 = n21668 & ~n28710 ;
  assign n28713 = n28712 ^ n28711 ^ 1'b0 ;
  assign n28714 = ~n4724 & n12125 ;
  assign n28715 = n9631 ^ n9538 ^ 1'b0 ;
  assign n28716 = ~n28714 & n28715 ;
  assign n28717 = n7965 & n26627 ;
  assign n28718 = ~n11918 & n28717 ;
  assign n28719 = n5707 & n6311 ;
  assign n28720 = n1372 | n1465 ;
  assign n28721 = n16156 ^ n11638 ^ 1'b0 ;
  assign n28722 = n28720 & n28721 ;
  assign n28723 = n28722 ^ n2112 ^ 1'b0 ;
  assign n28724 = n1379 & n11137 ;
  assign n28725 = n26297 & ~n28724 ;
  assign n28726 = n8324 ^ n2773 ^ 1'b0 ;
  assign n28727 = n20281 | n28726 ;
  assign n28728 = n28727 ^ n19118 ^ 1'b0 ;
  assign n28729 = n21944 ^ n16430 ^ 1'b0 ;
  assign n28730 = ~n2381 & n3285 ;
  assign n28731 = n28730 ^ n5916 ^ 1'b0 ;
  assign n28732 = n25408 | n28731 ;
  assign n28733 = n10096 & n10241 ;
  assign n28734 = n28733 ^ n2938 ^ 1'b0 ;
  assign n28735 = n14403 ^ n10929 ^ 1'b0 ;
  assign n28736 = n2225 & ~n28735 ;
  assign n28737 = ~n6574 & n26403 ;
  assign n28738 = n21114 ^ n3004 ^ 1'b0 ;
  assign n28739 = n26648 & n28738 ;
  assign n28740 = ~n146 & n28739 ;
  assign n28741 = n1018 & n28740 ;
  assign n28742 = n16518 ^ n4588 ^ 1'b0 ;
  assign n28743 = ~n7476 & n16010 ;
  assign n28744 = ~n23281 & n27933 ;
  assign n28745 = n28744 ^ n13954 ^ 1'b0 ;
  assign n28746 = n4753 & ~n10475 ;
  assign n28747 = n7111 & n28746 ;
  assign n28748 = n6641 ^ n1764 ^ 1'b0 ;
  assign n28749 = ~n6240 & n28748 ;
  assign n28750 = ( n2432 & ~n5109 ) | ( n2432 & n28749 ) | ( ~n5109 & n28749 ) ;
  assign n28751 = n18513 & n28750 ;
  assign n28752 = n10280 | n17439 ;
  assign n28753 = n28752 ^ n1718 ^ 1'b0 ;
  assign n28754 = ~n9588 & n28753 ;
  assign n28755 = n28754 ^ n17818 ^ n17598 ;
  assign n28756 = n5897 ^ n1588 ^ 1'b0 ;
  assign n28757 = ~n553 & n16788 ;
  assign n28758 = n28756 & n28757 ;
  assign n28759 = n938 | n10836 ;
  assign n28760 = n6945 & n28759 ;
  assign n28761 = n28760 ^ n19235 ^ 1'b0 ;
  assign n28762 = n536 & ~n9597 ;
  assign n28763 = n16971 & ~n28762 ;
  assign n28764 = n11355 ^ n3833 ^ 1'b0 ;
  assign n28765 = n26480 & ~n28764 ;
  assign n28766 = n492 & ~n5929 ;
  assign n28767 = n28766 ^ n875 ^ 1'b0 ;
  assign n28768 = n7929 ^ n4505 ^ 1'b0 ;
  assign n28769 = n28768 ^ n14955 ^ 1'b0 ;
  assign n28770 = n1592 & ~n28769 ;
  assign n28771 = n28767 & n28770 ;
  assign n28772 = ~n2721 & n22353 ;
  assign n28773 = n28771 | n28772 ;
  assign n28774 = n20667 | n28773 ;
  assign n28775 = ~n28765 & n28774 ;
  assign n28776 = ~n23951 & n28775 ;
  assign n28777 = n17907 ^ n1438 ^ 1'b0 ;
  assign n28778 = n5827 | n13413 ;
  assign n28779 = ~n2885 & n12786 ;
  assign n28780 = n28779 ^ n439 ^ 1'b0 ;
  assign n28781 = n28778 | n28780 ;
  assign n28782 = ~n6494 & n28781 ;
  assign n28783 = n1024 | n5447 ;
  assign n28784 = n28783 ^ n535 ^ 1'b0 ;
  assign n28785 = n18711 ^ n3833 ^ 1'b0 ;
  assign n28786 = n28784 & n28785 ;
  assign n28787 = n28786 ^ n3811 ^ 1'b0 ;
  assign n28788 = n1481 & n25455 ;
  assign n28789 = n28788 ^ n11406 ^ 1'b0 ;
  assign n28790 = n6088 ^ n2780 ^ 1'b0 ;
  assign n28791 = n15737 & n28790 ;
  assign n28792 = ~n7054 & n10432 ;
  assign n28793 = ~n28791 & n28792 ;
  assign n28794 = n18760 ^ n16809 ^ 1'b0 ;
  assign n28795 = ~n10553 & n17103 ;
  assign n28796 = n563 & n28795 ;
  assign n28797 = n28796 ^ n7342 ^ 1'b0 ;
  assign n28798 = ~n2747 & n28797 ;
  assign n28801 = n6988 & n17887 ;
  assign n28800 = n8357 & ~n9803 ;
  assign n28802 = n28801 ^ n28800 ^ 1'b0 ;
  assign n28803 = n28802 ^ n4434 ^ n2082 ;
  assign n28799 = n13891 & n25752 ;
  assign n28804 = n28803 ^ n28799 ^ n14206 ;
  assign n28805 = n14276 & n22884 ;
  assign n28806 = n4780 & n12596 ;
  assign n28807 = n16285 ^ n14081 ^ 1'b0 ;
  assign n28808 = ~n7109 & n28807 ;
  assign n28809 = ~n8998 & n17730 ;
  assign n28810 = n9583 & ~n28809 ;
  assign n28814 = n1340 & ~n3382 ;
  assign n28815 = n10253 & n28814 ;
  assign n28811 = n592 | n1865 ;
  assign n28812 = n28811 ^ n7657 ^ 1'b0 ;
  assign n28813 = n28812 ^ n18395 ^ 1'b0 ;
  assign n28816 = n28815 ^ n28813 ^ 1'b0 ;
  assign n28817 = n17170 | n18363 ;
  assign n28818 = n28816 | n28817 ;
  assign n28819 = n8010 ^ n3574 ^ 1'b0 ;
  assign n28820 = n13977 & ~n28819 ;
  assign n28823 = n17198 ^ n4082 ^ 1'b0 ;
  assign n28824 = n3372 | n28476 ;
  assign n28825 = n28823 & ~n28824 ;
  assign n28821 = n16303 ^ n14753 ^ 1'b0 ;
  assign n28822 = ~n11437 & n28821 ;
  assign n28826 = n28825 ^ n28822 ^ 1'b0 ;
  assign n28827 = n10452 ^ n3109 ^ n3040 ;
  assign n28828 = n11223 & ~n28406 ;
  assign n28829 = ~n6444 & n16425 ;
  assign n28830 = n18372 & ~n28829 ;
  assign n28831 = n28830 ^ n2356 ^ 1'b0 ;
  assign n28832 = n22235 ^ n16087 ^ 1'b0 ;
  assign n28833 = n414 | n28832 ;
  assign n28834 = n9895 & n11550 ;
  assign n28835 = ~n2940 & n16177 ;
  assign n28836 = n28835 ^ n5671 ^ 1'b0 ;
  assign n28837 = n2473 ^ n1738 ^ 1'b0 ;
  assign n28838 = n5106 & ~n24779 ;
  assign n28839 = n28838 ^ n17662 ^ 1'b0 ;
  assign n28840 = ( n10140 & n28837 ) | ( n10140 & ~n28839 ) | ( n28837 & ~n28839 ) ;
  assign n28841 = n22117 | n26543 ;
  assign n28842 = n3958 & ~n28841 ;
  assign n28843 = n10117 ^ n1779 ^ 1'b0 ;
  assign n28844 = ~n28842 & n28843 ;
  assign n28845 = ~n1392 & n28844 ;
  assign n28846 = n3113 | n5579 ;
  assign n28847 = n28846 ^ n24304 ^ 1'b0 ;
  assign n28848 = ~n17427 & n24889 ;
  assign n28849 = ~n4751 & n28848 ;
  assign n28851 = n91 & ~n2915 ;
  assign n28850 = n1770 & n2389 ;
  assign n28852 = n28851 ^ n28850 ^ 1'b0 ;
  assign n28853 = ~n5049 & n28852 ;
  assign n28854 = n3476 | n12126 ;
  assign n28855 = n28854 ^ n6020 ^ 1'b0 ;
  assign n28856 = ( n12551 & ~n26595 ) | ( n12551 & n28855 ) | ( ~n26595 & n28855 ) ;
  assign n28857 = n3257 & ~n21916 ;
  assign n28858 = n28857 ^ n28425 ^ 1'b0 ;
  assign n28861 = n11552 | n19317 ;
  assign n28859 = ~n5551 & n18765 ;
  assign n28860 = n1360 & n28859 ;
  assign n28862 = n28861 ^ n28860 ^ 1'b0 ;
  assign n28863 = n2909 ^ n1408 ^ 1'b0 ;
  assign n28864 = n1624 | n6308 ;
  assign n28865 = n28864 ^ n15588 ^ 1'b0 ;
  assign n28866 = ( ~n16117 & n28863 ) | ( ~n16117 & n28865 ) | ( n28863 & n28865 ) ;
  assign n28870 = n765 & n2645 ;
  assign n28871 = n2569 & ~n28870 ;
  assign n28872 = ~n1469 & n28871 ;
  assign n28868 = n6479 ^ n6397 ^ 1'b0 ;
  assign n28869 = n6032 & n28868 ;
  assign n28873 = n28872 ^ n28869 ^ 1'b0 ;
  assign n28867 = n23481 ^ n21182 ^ 1'b0 ;
  assign n28874 = n28873 ^ n28867 ^ 1'b0 ;
  assign n28875 = ~n28866 & n28874 ;
  assign n28877 = n12320 ^ n3766 ^ 1'b0 ;
  assign n28878 = n12368 & n28877 ;
  assign n28876 = n15467 | n17126 ;
  assign n28879 = n28878 ^ n28876 ^ 1'b0 ;
  assign n28880 = ~n755 & n14737 ;
  assign n28881 = n547 & n692 ;
  assign n28882 = ~n692 & n28881 ;
  assign n28883 = n24391 ^ n302 ^ 1'b0 ;
  assign n28884 = n10998 & n28883 ;
  assign n28885 = ~n10337 & n28884 ;
  assign n28886 = n28882 & n28885 ;
  assign n28887 = ( n13573 & n15403 ) | ( n13573 & ~n28886 ) | ( n15403 & ~n28886 ) ;
  assign n28888 = n1006 ^ n184 ^ 1'b0 ;
  assign n28889 = ~n8977 & n27970 ;
  assign n28890 = n28889 ^ n18986 ^ 1'b0 ;
  assign n28891 = ~n8373 & n21391 ;
  assign n28892 = n18068 & n28891 ;
  assign n28893 = ( ~n1182 & n1862 ) | ( ~n1182 & n8604 ) | ( n1862 & n8604 ) ;
  assign n28894 = n28893 ^ n27332 ^ n18628 ;
  assign n28895 = n21759 & ~n25010 ;
  assign n28896 = n28895 ^ n5618 ^ 1'b0 ;
  assign n28897 = n7541 ^ n3554 ^ 1'b0 ;
  assign n28898 = n1471 | n7660 ;
  assign n28899 = n19904 | n28898 ;
  assign n28900 = n710 & n17529 ;
  assign n28901 = n28900 ^ n20240 ^ 1'b0 ;
  assign n28902 = n10107 ^ n3226 ^ 1'b0 ;
  assign n28903 = n28902 ^ n19797 ^ 1'b0 ;
  assign n28904 = n7542 ^ n5518 ^ 1'b0 ;
  assign n28905 = n5803 | n15321 ;
  assign n28906 = n3041 | n28905 ;
  assign n28907 = n1217 | n13794 ;
  assign n28908 = n28907 ^ n17116 ^ 1'b0 ;
  assign n28909 = n28908 ^ n10507 ^ 1'b0 ;
  assign n28910 = n1944 | n28909 ;
  assign n28911 = ~n770 & n4419 ;
  assign n28917 = n12799 ^ n4833 ^ 1'b0 ;
  assign n28912 = ~n15447 & n21868 ;
  assign n28913 = n28912 ^ n2034 ^ 1'b0 ;
  assign n28914 = n4991 & n12077 ;
  assign n28915 = n28914 ^ n20969 ^ 1'b0 ;
  assign n28916 = n28913 & ~n28915 ;
  assign n28918 = n28917 ^ n28916 ^ 1'b0 ;
  assign n28919 = n27529 ^ n8235 ^ 1'b0 ;
  assign n28920 = n3361 | n28919 ;
  assign n28921 = n28920 ^ n17043 ^ n197 ;
  assign n28922 = n18048 ^ n3417 ^ 1'b0 ;
  assign n28923 = n7004 | n28922 ;
  assign n28924 = ( ~n614 & n1703 ) | ( ~n614 & n28923 ) | ( n1703 & n28923 ) ;
  assign n28925 = n15337 & n18817 ;
  assign n28926 = n23115 ^ n22852 ^ 1'b0 ;
  assign n28927 = ~n1912 & n4005 ;
  assign n28928 = n3687 & ~n5139 ;
  assign n28929 = n25521 ^ n4835 ^ 1'b0 ;
  assign n28930 = n9020 | n28929 ;
  assign n28931 = n6473 | n28930 ;
  assign n28932 = n10653 ^ n5700 ^ 1'b0 ;
  assign n28933 = n7414 & n28932 ;
  assign n28934 = n22893 ^ n18381 ^ 1'b0 ;
  assign n28935 = n1660 & ~n6473 ;
  assign n28936 = ~n695 & n28415 ;
  assign n28937 = n17352 ^ n17166 ^ 1'b0 ;
  assign n28938 = ~n13850 & n28937 ;
  assign n28939 = n28938 ^ n28817 ^ n12725 ;
  assign n28940 = n362 & ~n14820 ;
  assign n28941 = n17420 ^ n14431 ^ 1'b0 ;
  assign n28942 = n26004 ^ n25289 ^ 1'b0 ;
  assign n28943 = n28941 & n28942 ;
  assign n28944 = ~n3444 & n15481 ;
  assign n28945 = n28944 ^ n2173 ^ 1'b0 ;
  assign n28946 = n4860 ^ n2938 ^ 1'b0 ;
  assign n28947 = n1658 & ~n15028 ;
  assign n28948 = n25948 | n27498 ;
  assign n28949 = ~n4762 & n13352 ;
  assign n28950 = n28949 ^ n7685 ^ 1'b0 ;
  assign n28951 = n28950 ^ n13857 ^ n12392 ;
  assign n28952 = n16815 & ~n28951 ;
  assign n28953 = n9664 & ~n19050 ;
  assign n28954 = n4668 & n28953 ;
  assign n28955 = n5740 | n28954 ;
  assign n28956 = n2805 | n28955 ;
  assign n28957 = n10866 & ~n28956 ;
  assign n28958 = n24089 ^ n15203 ^ 1'b0 ;
  assign n28959 = n2876 & n28958 ;
  assign n28960 = ( n3647 & n6931 ) | ( n3647 & n9276 ) | ( n6931 & n9276 ) ;
  assign n28961 = n24007 | n28960 ;
  assign n28962 = n28961 ^ n23790 ^ 1'b0 ;
  assign n28963 = n4395 & ~n6316 ;
  assign n28964 = ~n28962 & n28963 ;
  assign n28965 = ( n14614 & ~n20512 ) | ( n14614 & n28520 ) | ( ~n20512 & n28520 ) ;
  assign n28966 = n11471 & n27843 ;
  assign n28967 = n14392 | n21772 ;
  assign n28972 = n1138 & ~n17880 ;
  assign n28973 = n28972 ^ n1900 ^ 1'b0 ;
  assign n28974 = ~n8258 & n28973 ;
  assign n28968 = n11300 ^ n6102 ^ 1'b0 ;
  assign n28969 = n14032 & ~n28968 ;
  assign n28970 = n14913 & n28969 ;
  assign n28971 = ( x8 & n19879 ) | ( x8 & n28970 ) | ( n19879 & n28970 ) ;
  assign n28975 = n28974 ^ n28971 ^ n16237 ;
  assign n28976 = n8174 ^ n3425 ^ 1'b0 ;
  assign n28977 = n19489 ^ n4744 ^ 1'b0 ;
  assign n28978 = ~n28976 & n28977 ;
  assign n28979 = ~n11333 & n26274 ;
  assign n28980 = n8667 & n28979 ;
  assign n28981 = n13743 ^ n8885 ^ 1'b0 ;
  assign n28982 = n15134 | n28981 ;
  assign n28983 = n26873 & ~n28982 ;
  assign n28984 = n1211 & n11179 ;
  assign n28985 = ~n7449 & n12516 ;
  assign n28986 = ~n13 & n6740 ;
  assign n28987 = n28986 ^ n2780 ^ 1'b0 ;
  assign n28988 = n21441 ^ n11286 ^ n10000 ;
  assign n28989 = n2614 | n28988 ;
  assign n28990 = n28989 ^ n11470 ^ 1'b0 ;
  assign n28991 = n8000 | n28335 ;
  assign n28992 = n2507 & ~n4781 ;
  assign n28996 = ~n13137 & n20521 ;
  assign n28997 = n28996 ^ n14384 ^ 1'b0 ;
  assign n28993 = n14511 ^ n6608 ^ 1'b0 ;
  assign n28994 = n8233 & n28993 ;
  assign n28995 = ~n2560 & n28994 ;
  assign n28998 = n28997 ^ n28995 ^ 1'b0 ;
  assign n28999 = ~n1334 & n9880 ;
  assign n29000 = n28999 ^ n12985 ^ n7156 ;
  assign n29001 = n29000 ^ n4080 ^ 1'b0 ;
  assign n29002 = ~n8697 & n29001 ;
  assign n29003 = n16758 ^ n6180 ^ 1'b0 ;
  assign n29004 = n2317 | n29003 ;
  assign n29005 = n29004 ^ n28258 ^ 1'b0 ;
  assign n29006 = n2488 & ~n29005 ;
  assign n29007 = n8974 ^ n4203 ^ 1'b0 ;
  assign n29008 = n29007 ^ n7267 ^ n6494 ;
  assign n29009 = n11122 ^ n11115 ^ 1'b0 ;
  assign n29010 = n7735 | n29009 ;
  assign n29011 = ~n8074 & n29010 ;
  assign n29012 = ~n2621 & n29011 ;
  assign n29013 = n11234 & ~n13884 ;
  assign n29014 = n29013 ^ n9294 ^ 1'b0 ;
  assign n29015 = ~n25757 & n29014 ;
  assign n29016 = n25379 ^ n5734 ^ 1'b0 ;
  assign n29017 = ~n13708 & n29016 ;
  assign n29018 = ( ~n7407 & n8486 ) | ( ~n7407 & n11717 ) | ( n8486 & n11717 ) ;
  assign n29019 = ( n2120 & ~n4793 ) | ( n2120 & n29018 ) | ( ~n4793 & n29018 ) ;
  assign n29020 = n10929 & ~n12976 ;
  assign n29021 = n6750 ^ n4741 ^ 1'b0 ;
  assign n29022 = n10598 & n29021 ;
  assign n29023 = n18162 & n29022 ;
  assign n29025 = n12819 ^ n8064 ^ 1'b0 ;
  assign n29026 = n10715 & n29025 ;
  assign n29024 = n3408 & n16933 ;
  assign n29027 = n29026 ^ n29024 ^ 1'b0 ;
  assign n29028 = n18772 ^ n6610 ^ n2258 ;
  assign n29029 = ( n12682 & n22308 ) | ( n12682 & ~n29028 ) | ( n22308 & ~n29028 ) ;
  assign n29030 = n14957 ^ n456 ^ 1'b0 ;
  assign n29031 = n2101 & ~n20598 ;
  assign n29034 = n4017 | n5791 ;
  assign n29035 = n2724 | n29034 ;
  assign n29032 = n19404 ^ n38 ^ 1'b0 ;
  assign n29033 = n29032 ^ n368 ^ 1'b0 ;
  assign n29036 = n29035 ^ n29033 ^ n24545 ;
  assign n29037 = n13668 ^ n8117 ^ 1'b0 ;
  assign n29038 = n2655 & ~n29037 ;
  assign n29039 = n20846 & n29038 ;
  assign n29040 = n10298 & n29039 ;
  assign n29041 = n229 & ~n4523 ;
  assign n29042 = n4523 & n29041 ;
  assign n29043 = n5320 | n29042 ;
  assign n29044 = n3349 | n29043 ;
  assign n29045 = n5226 ^ n3328 ^ 1'b0 ;
  assign n29046 = n6464 & n29045 ;
  assign n29047 = n17661 & n27618 ;
  assign n29048 = ~n29046 & n29047 ;
  assign n29049 = n136 | n29048 ;
  assign n29050 = n17932 & ~n29049 ;
  assign n29051 = n29044 | n29050 ;
  assign n29052 = ( n1853 & n3252 ) | ( n1853 & ~n11481 ) | ( n3252 & ~n11481 ) ;
  assign n29053 = n29052 ^ n15958 ^ 1'b0 ;
  assign n29054 = n16208 & n29053 ;
  assign n29055 = n18065 ^ n16257 ^ 1'b0 ;
  assign n29056 = ~n8024 & n29055 ;
  assign n29057 = n810 & n1771 ;
  assign n29058 = n1969 & n29057 ;
  assign n29059 = n3578 & ~n24256 ;
  assign n29060 = n29059 ^ n6472 ^ 1'b0 ;
  assign n29061 = ~n13138 & n18462 ;
  assign n29062 = ~n29060 & n29061 ;
  assign n29063 = n19680 & ~n26169 ;
  assign n29064 = n23649 ^ n8600 ^ 1'b0 ;
  assign n29065 = ~n379 & n27943 ;
  assign n29066 = ~n3359 & n13272 ;
  assign n29067 = n10145 & n29066 ;
  assign n29068 = n3909 & n14111 ;
  assign n29069 = n29068 ^ n16098 ^ 1'b0 ;
  assign n29070 = n21823 ^ n966 ^ n625 ;
  assign n29071 = n24886 ^ n12781 ^ 1'b0 ;
  assign n29072 = n3774 | n29071 ;
  assign n29074 = n8958 ^ n4180 ^ 1'b0 ;
  assign n29073 = n564 & ~n12916 ;
  assign n29075 = n29074 ^ n29073 ^ 1'b0 ;
  assign n29076 = n14516 | n17025 ;
  assign n29077 = n29076 ^ n1377 ^ 1'b0 ;
  assign n29078 = n22632 & ~n29077 ;
  assign n29079 = n29078 ^ n25504 ^ 1'b0 ;
  assign n29086 = n4374 & ~n9511 ;
  assign n29080 = n4317 & ~n8630 ;
  assign n29081 = n17404 & ~n29080 ;
  assign n29082 = ~n4789 & n29081 ;
  assign n29083 = n15796 & n29082 ;
  assign n29084 = n29083 ^ n360 ^ 1'b0 ;
  assign n29085 = n8689 & n29084 ;
  assign n29087 = n29086 ^ n29085 ^ n6269 ;
  assign n29088 = n23846 ^ n7400 ^ 1'b0 ;
  assign n29089 = n24311 ^ n4460 ^ 1'b0 ;
  assign n29091 = n14331 ^ n8887 ^ 1'b0 ;
  assign n29092 = n20628 & ~n29091 ;
  assign n29090 = n21496 ^ n5982 ^ 1'b0 ;
  assign n29093 = n29092 ^ n29090 ^ n4886 ;
  assign n29094 = n8724 & ~n19377 ;
  assign n29095 = n29094 ^ n12634 ^ 1'b0 ;
  assign n29096 = n2315 | n29095 ;
  assign n29097 = n273 & ~n4378 ;
  assign n29098 = n5810 & ~n14640 ;
  assign n29099 = n3428 & ~n18264 ;
  assign n29100 = n29099 ^ x5 ^ 1'b0 ;
  assign n29101 = n27277 ^ n24140 ^ n12258 ;
  assign n29106 = n12658 & ~n13723 ;
  assign n29107 = n29106 ^ n5968 ^ 1'b0 ;
  assign n29102 = n8969 & ~n13175 ;
  assign n29103 = ~n2656 & n29102 ;
  assign n29104 = n29103 ^ n23645 ^ 1'b0 ;
  assign n29105 = n6586 | n29104 ;
  assign n29108 = n29107 ^ n29105 ^ n7490 ;
  assign n29109 = ( n235 & n4004 ) | ( n235 & n29108 ) | ( n4004 & n29108 ) ;
  assign n29110 = x10 & ~n831 ;
  assign n29111 = ~x10 & n29110 ;
  assign n29112 = n5803 & ~n29111 ;
  assign n29113 = n1383 & n7968 ;
  assign n29114 = ~n7968 & n29113 ;
  assign n29115 = n1434 | n2094 ;
  assign n29116 = n2094 & ~n29115 ;
  assign n29117 = n29114 & ~n29116 ;
  assign n29118 = n1382 & ~n6065 ;
  assign n29119 = ~n1382 & n29118 ;
  assign n29120 = n29117 | n29119 ;
  assign n29121 = n29117 & ~n29120 ;
  assign n29122 = n8551 | n29121 ;
  assign n29123 = n29121 & ~n29122 ;
  assign n29124 = n29123 ^ n17763 ^ 1'b0 ;
  assign n29125 = ~n29112 & n29124 ;
  assign n29126 = n2656 & ~n24558 ;
  assign n29127 = n29126 ^ n6095 ^ 1'b0 ;
  assign n29128 = ~n7710 & n14992 ;
  assign n29129 = n10665 ^ n1157 ^ 1'b0 ;
  assign n29130 = n12015 ^ n6184 ^ 1'b0 ;
  assign n29131 = n17506 & ~n23055 ;
  assign n29132 = n9151 ^ n6431 ^ 1'b0 ;
  assign n29133 = n1484 & ~n29132 ;
  assign n29134 = n16190 ^ n11968 ^ 1'b0 ;
  assign n29135 = n29133 & ~n29134 ;
  assign n29136 = n6176 & ~n8596 ;
  assign n29137 = ~n3531 & n5492 ;
  assign n29138 = n29137 ^ n5380 ^ 1'b0 ;
  assign n29139 = n2435 | n25340 ;
  assign n29140 = n3955 | n29139 ;
  assign n29141 = n29140 ^ n7093 ^ 1'b0 ;
  assign n29142 = n29138 | n29141 ;
  assign n29143 = n29136 & ~n29142 ;
  assign n29144 = n29143 ^ n14374 ^ 1'b0 ;
  assign n29145 = n16305 & ~n29144 ;
  assign n29146 = n14563 & n29145 ;
  assign n29147 = n623 & ~n1944 ;
  assign n29148 = n15368 & ~n25909 ;
  assign n29149 = n20719 ^ n12965 ^ 1'b0 ;
  assign n29150 = ~n12594 & n17771 ;
  assign n29151 = n4395 ^ n243 ^ 1'b0 ;
  assign n29152 = n25926 ^ n2507 ^ 1'b0 ;
  assign n29153 = n16310 | n21618 ;
  assign n29154 = n24779 ^ n4344 ^ 1'b0 ;
  assign n29160 = n22235 ^ n10775 ^ 1'b0 ;
  assign n29155 = n25571 ^ n18114 ^ 1'b0 ;
  assign n29156 = n22984 & ~n29155 ;
  assign n29157 = ~n6040 & n29156 ;
  assign n29158 = ~n14735 & n14883 ;
  assign n29159 = n29157 & n29158 ;
  assign n29161 = n29160 ^ n29159 ^ 1'b0 ;
  assign n29162 = n7344 | n22286 ;
  assign n29163 = ( n4317 & n4885 ) | ( n4317 & ~n16055 ) | ( n4885 & ~n16055 ) ;
  assign n29164 = ( ~n26880 & n29162 ) | ( ~n26880 & n29163 ) | ( n29162 & n29163 ) ;
  assign n29165 = n20045 ^ n2715 ^ 1'b0 ;
  assign n29166 = n23309 ^ n7704 ^ 1'b0 ;
  assign n29167 = n12260 & ~n29166 ;
  assign n29168 = n29167 ^ n11383 ^ 1'b0 ;
  assign n29169 = n21381 ^ n14254 ^ 1'b0 ;
  assign n29170 = n29168 & n29169 ;
  assign n29172 = n1304 & n2656 ;
  assign n29171 = n18920 | n20685 ;
  assign n29173 = n29172 ^ n29171 ^ 1'b0 ;
  assign n29174 = n2489 & n9319 ;
  assign n29175 = n29174 ^ n3981 ^ 1'b0 ;
  assign n29176 = ~n3348 & n29175 ;
  assign n29177 = n7883 | n29176 ;
  assign n29178 = n19150 ^ n15185 ^ n12198 ;
  assign n29179 = n58 & ~n152 ;
  assign n29180 = ~n58 & n29179 ;
  assign n29181 = n3798 & ~n29180 ;
  assign n29182 = n29180 & n29181 ;
  assign n29183 = n365 & n479 ;
  assign n29184 = ~n365 & n29183 ;
  assign n29185 = ~n1212 & n1401 ;
  assign n29186 = n1212 & n29185 ;
  assign n29187 = n29184 & ~n29186 ;
  assign n29188 = n4949 & ~n5981 ;
  assign n29189 = n29187 & n29188 ;
  assign n29190 = n3277 | n29189 ;
  assign n29191 = n3277 & ~n29190 ;
  assign n29192 = n29191 ^ n2258 ^ 1'b0 ;
  assign n29193 = n29192 ^ n13493 ^ 1'b0 ;
  assign n29194 = ~n29182 & n29193 ;
  assign n29195 = n22660 ^ n12130 ^ 1'b0 ;
  assign n29196 = ~n8992 & n29195 ;
  assign n29197 = ( n29178 & n29194 ) | ( n29178 & ~n29196 ) | ( n29194 & ~n29196 ) ;
  assign n29198 = n6434 & ~n27787 ;
  assign n29199 = n10610 & n29198 ;
  assign n29200 = n7020 & ~n9416 ;
  assign n29201 = n29199 & n29200 ;
  assign n29202 = n3020 | n22611 ;
  assign n29203 = n13008 | n29202 ;
  assign n29204 = n1079 | n22496 ;
  assign n29205 = n29204 ^ n1936 ^ 1'b0 ;
  assign n29206 = ( n4526 & n13891 ) | ( n4526 & n23299 ) | ( n13891 & n23299 ) ;
  assign n29207 = ( n1542 & ~n6794 ) | ( n1542 & n29206 ) | ( ~n6794 & n29206 ) ;
  assign n29208 = n4754 | n8502 ;
  assign n29209 = n26853 & ~n29208 ;
  assign n29210 = n7643 | n18389 ;
  assign n29213 = n150 & ~n9775 ;
  assign n29214 = n6278 & ~n29213 ;
  assign n29211 = n15677 & n25308 ;
  assign n29212 = ~n8100 & n29211 ;
  assign n29215 = n29214 ^ n29212 ^ 1'b0 ;
  assign n29216 = ~n12868 & n29215 ;
  assign n29217 = n4952 ^ n4263 ^ 1'b0 ;
  assign n29218 = ~n9837 & n29217 ;
  assign n29219 = n24050 ^ n22221 ^ 1'b0 ;
  assign n29220 = n29218 & ~n29219 ;
  assign n29221 = n2355 & n12794 ;
  assign n29222 = ~n2141 & n29221 ;
  assign n29223 = ( n978 & n3106 ) | ( n978 & n21847 ) | ( n3106 & n21847 ) ;
  assign n29224 = n746 & n8834 ;
  assign n29225 = ~n29223 & n29224 ;
  assign n29226 = n10403 & ~n11600 ;
  assign n29227 = ( ~n4533 & n6506 ) | ( ~n4533 & n29226 ) | ( n6506 & n29226 ) ;
  assign n29228 = n7839 ^ n886 ^ 1'b0 ;
  assign n29229 = n11659 | n12081 ;
  assign n29230 = n29229 ^ n14687 ^ 1'b0 ;
  assign n29231 = n12985 ^ n5547 ^ 1'b0 ;
  assign n29232 = n551 & ~n1945 ;
  assign n29233 = n3886 & n29232 ;
  assign n29234 = n11576 & ~n12405 ;
  assign n29235 = n29234 ^ n1469 ^ 1'b0 ;
  assign n29236 = n29235 ^ n24969 ^ 1'b0 ;
  assign n29237 = ~n14953 & n29236 ;
  assign n29238 = n12513 & ~n16251 ;
  assign n29239 = n24669 ^ n2399 ^ 1'b0 ;
  assign n29240 = n4888 & ~n22221 ;
  assign n29241 = n9584 & n29240 ;
  assign n29242 = n2619 & n29241 ;
  assign n29243 = ~n4169 & n5886 ;
  assign n29244 = ~n5886 & n29243 ;
  assign n29245 = n6479 & ~n29244 ;
  assign n29246 = n372 | n29245 ;
  assign n29247 = n29246 ^ n11523 ^ 1'b0 ;
  assign n29248 = n16667 & ~n29247 ;
  assign n29249 = n9189 | n25027 ;
  assign n29250 = n29248 | n29249 ;
  assign n29251 = n1071 | n28257 ;
  assign n29252 = n11367 ^ n2635 ^ 1'b0 ;
  assign n29253 = n23274 & n29252 ;
  assign n29254 = ~n4267 & n5849 ;
  assign n29255 = ~n16772 & n29254 ;
  assign n29256 = n8789 | n29255 ;
  assign n29257 = n29256 ^ n16435 ^ 1'b0 ;
  assign n29258 = n29253 | n29257 ;
  assign n29259 = n184 | n645 ;
  assign n29260 = n645 & ~n29259 ;
  assign n29261 = n235 & n29260 ;
  assign n29262 = n277 | n29261 ;
  assign n29263 = n26 | n296 ;
  assign n29264 = n296 & ~n29263 ;
  assign n29265 = n29262 | n29264 ;
  assign n29266 = n29262 & ~n29265 ;
  assign n29267 = n305 & n509 ;
  assign n29268 = ~n509 & n29267 ;
  assign n29269 = n1142 & ~n29268 ;
  assign n29270 = n29266 & n29269 ;
  assign n29271 = n3580 & ~n29270 ;
  assign n29272 = n12924 ^ n2526 ^ 1'b0 ;
  assign n29273 = n29271 & n29272 ;
  assign n29274 = n27 & ~n4259 ;
  assign n29275 = n29274 ^ n12175 ^ 1'b0 ;
  assign n29276 = n1128 | n29275 ;
  assign n29277 = ( n17644 & n24123 ) | ( n17644 & ~n29276 ) | ( n24123 & ~n29276 ) ;
  assign n29280 = n2891 & n6149 ;
  assign n29278 = n9553 & ~n10755 ;
  assign n29279 = ~n5045 & n29278 ;
  assign n29281 = n29280 ^ n29279 ^ 1'b0 ;
  assign n29282 = n12007 ^ n3589 ^ 1'b0 ;
  assign n29283 = n21105 | n29282 ;
  assign n29284 = ( n5756 & n29281 ) | ( n5756 & ~n29283 ) | ( n29281 & ~n29283 ) ;
  assign n29285 = n16861 ^ n1902 ^ 1'b0 ;
  assign n29286 = n1650 | n29285 ;
  assign n29287 = n29286 ^ n21469 ^ 1'b0 ;
  assign n29288 = n26954 & ~n29287 ;
  assign n29289 = n15347 | n27519 ;
  assign n29290 = n29289 ^ n16092 ^ 1'b0 ;
  assign n29291 = n29290 ^ n15221 ^ 1'b0 ;
  assign n29292 = n10114 & n29291 ;
  assign n29293 = n11352 ^ n9198 ^ 1'b0 ;
  assign n29294 = n14937 & ~n29293 ;
  assign n29295 = n29294 ^ n7830 ^ n3565 ;
  assign n29296 = n4154 & n15086 ;
  assign n29297 = ~n27234 & n29296 ;
  assign n29298 = n17156 & n19158 ;
  assign n29299 = n28495 ^ n26187 ^ 1'b0 ;
  assign n29300 = n13593 ^ n4274 ^ 1'b0 ;
  assign n29301 = n20862 | n27299 ;
  assign n29302 = n4931 & ~n29301 ;
  assign n29303 = n2408 | n10177 ;
  assign n29304 = n29303 ^ n9326 ^ 1'b0 ;
  assign n29305 = n29304 ^ n9912 ^ 1'b0 ;
  assign n29306 = n20431 ^ n8001 ^ 1'b0 ;
  assign n29307 = n29305 & ~n29306 ;
  assign n29308 = ~n28400 & n29307 ;
  assign n29309 = n10211 ^ n1545 ^ 1'b0 ;
  assign n29310 = n20391 ^ n11308 ^ 1'b0 ;
  assign n29311 = n29309 | n29310 ;
  assign n29312 = ( ~n3030 & n10567 ) | ( ~n3030 & n21445 ) | ( n10567 & n21445 ) ;
  assign n29313 = ~n6581 & n10837 ;
  assign n29314 = n29313 ^ n7447 ^ 1'b0 ;
  assign n29315 = n18969 & ~n29314 ;
  assign n29316 = ~n1227 & n29315 ;
  assign n29317 = n25549 ^ n5893 ^ 1'b0 ;
  assign n29318 = n7753 | n11276 ;
  assign n29319 = n29318 ^ n9010 ^ 1'b0 ;
  assign n29320 = n29317 & n29319 ;
  assign n29321 = n29320 ^ n13454 ^ 1'b0 ;
  assign n29322 = ( n3060 & ~n9391 ) | ( n3060 & n10045 ) | ( ~n9391 & n10045 ) ;
  assign n29327 = n896 & n8887 ;
  assign n29323 = n8445 | n17404 ;
  assign n29324 = n4395 & ~n29323 ;
  assign n29325 = n8106 & n11547 ;
  assign n29326 = ( n1741 & n29324 ) | ( n1741 & ~n29325 ) | ( n29324 & ~n29325 ) ;
  assign n29328 = n29327 ^ n29326 ^ 1'b0 ;
  assign n29329 = n12393 | n22893 ;
  assign n29330 = n20724 & ~n29329 ;
  assign n29331 = n3157 ^ n1825 ^ 1'b0 ;
  assign n29332 = n23108 & ~n29331 ;
  assign n29333 = n27050 & ~n29332 ;
  assign n29334 = n3536 & ~n8419 ;
  assign n29335 = n12160 & n29334 ;
  assign n29336 = n8403 ^ n7665 ^ 1'b0 ;
  assign n29337 = n9324 & n29336 ;
  assign n29338 = n29337 ^ n4660 ^ 1'b0 ;
  assign n29339 = n11708 & ~n29338 ;
  assign n29340 = n8659 ^ n7588 ^ 1'b0 ;
  assign n29341 = n6666 | n29340 ;
  assign n29342 = n9642 ^ n6623 ^ 1'b0 ;
  assign n29343 = n4175 & n29342 ;
  assign n29344 = n16435 ^ n10377 ^ 1'b0 ;
  assign n29345 = n16673 ^ n4583 ^ 1'b0 ;
  assign n29346 = ~n3135 & n7971 ;
  assign n29347 = n29346 ^ n23936 ^ 1'b0 ;
  assign n29348 = n29347 ^ n16460 ^ 1'b0 ;
  assign n29349 = n23658 ^ n5580 ^ 1'b0 ;
  assign n29350 = n17415 & ~n29349 ;
  assign n29351 = n6224 ^ n1002 ^ 1'b0 ;
  assign n29352 = n29351 ^ n24141 ^ 1'b0 ;
  assign n29353 = ~n1994 & n29352 ;
  assign n29354 = n17364 ^ n1323 ^ 1'b0 ;
  assign n29355 = n18540 & ~n29354 ;
  assign n29356 = n18639 & n29355 ;
  assign n29357 = ~n25468 & n29356 ;
  assign n29358 = n514 & n2563 ;
  assign n29359 = n29358 ^ n8612 ^ 1'b0 ;
  assign n29360 = n19112 ^ n4629 ^ 1'b0 ;
  assign n29361 = n8281 & n29360 ;
  assign n29362 = ~n29359 & n29361 ;
  assign n29363 = n27624 ^ n2411 ^ 1'b0 ;
  assign n29364 = n14253 & n29363 ;
  assign n29365 = ( n16394 & ~n19144 ) | ( n16394 & n29364 ) | ( ~n19144 & n29364 ) ;
  assign n29366 = n12699 & ~n29365 ;
  assign n29367 = n4422 ^ n4405 ^ 1'b0 ;
  assign n29368 = n1761 & n27735 ;
  assign n29369 = n1938 & n2915 ;
  assign n29370 = n29369 ^ n1229 ^ 1'b0 ;
  assign n29372 = ( n1009 & n12317 ) | ( n1009 & ~n19088 ) | ( n12317 & ~n19088 ) ;
  assign n29371 = n22833 & n24776 ;
  assign n29373 = n29372 ^ n29371 ^ 1'b0 ;
  assign n29374 = n3240 | n28144 ;
  assign n29375 = n4787 & ~n23643 ;
  assign n29376 = n2085 & ~n29375 ;
  assign n29377 = n782 & n16813 ;
  assign n29378 = n18102 & ~n24599 ;
  assign n29381 = n17422 ^ n11749 ^ 1'b0 ;
  assign n29379 = ~n700 & n3818 ;
  assign n29380 = ~n23946 & n29379 ;
  assign n29382 = n29381 ^ n29380 ^ 1'b0 ;
  assign n29383 = n29382 ^ n18064 ^ 1'b0 ;
  assign n29384 = ~n5306 & n12373 ;
  assign n29385 = n997 & n29384 ;
  assign n29386 = n24653 ^ n11349 ^ 1'b0 ;
  assign n29387 = n29385 | n29386 ;
  assign n29388 = n5665 & ~n23216 ;
  assign n29389 = n4240 & ~n18973 ;
  assign n29390 = n5890 & n10027 ;
  assign n29391 = ~n867 & n3367 ;
  assign n29392 = ~n813 & n29391 ;
  assign n29393 = n13255 ^ n4147 ^ 1'b0 ;
  assign n29394 = ~n29392 & n29393 ;
  assign n29395 = n29394 ^ n25191 ^ 1'b0 ;
  assign n29396 = n8376 | n29395 ;
  assign n29397 = n12575 | n29396 ;
  assign n29398 = n29397 ^ n28927 ^ 1'b0 ;
  assign n29399 = n15691 ^ n5387 ^ 1'b0 ;
  assign n29400 = n8263 ^ n423 ^ 1'b0 ;
  assign n29401 = n29305 ^ n1993 ^ 1'b0 ;
  assign n29402 = ~n2849 & n29401 ;
  assign n29403 = ~n3370 & n29402 ;
  assign n29404 = n29403 ^ n5710 ^ 1'b0 ;
  assign n29405 = n8949 ^ n4545 ^ 1'b0 ;
  assign n29406 = n3568 & n24621 ;
  assign n29407 = n29406 ^ n16165 ^ 1'b0 ;
  assign n29408 = n74 & ~n25143 ;
  assign n29409 = ~n29407 & n29408 ;
  assign n29410 = n3195 & n29409 ;
  assign n29411 = n10809 ^ n7545 ^ 1'b0 ;
  assign n29412 = n10217 & ~n29411 ;
  assign n29413 = ~n8562 & n25138 ;
  assign n29414 = n7427 & ~n19074 ;
  assign n29415 = n26541 & n29414 ;
  assign n29418 = n7156 & n15858 ;
  assign n29416 = n5706 ^ n5126 ^ 1'b0 ;
  assign n29417 = n18312 | n29416 ;
  assign n29419 = n29418 ^ n29417 ^ 1'b0 ;
  assign n29420 = ~n1111 & n29419 ;
  assign n29421 = n22991 ^ n7936 ^ 1'b0 ;
  assign n29422 = n29421 ^ n27192 ^ n5697 ;
  assign n29423 = n19772 | n26323 ;
  assign n29424 = n29423 ^ n29000 ^ 1'b0 ;
  assign n29425 = n5497 & n11813 ;
  assign n29426 = n870 ^ n699 ^ 1'b0 ;
  assign n29427 = n2512 & n14338 ;
  assign n29428 = n29427 ^ n2066 ^ 1'b0 ;
  assign n29429 = n28759 ^ n27001 ^ n6551 ;
  assign n29430 = n7254 ^ n646 ^ 1'b0 ;
  assign n29431 = n18111 & n25319 ;
  assign n29432 = n29431 ^ n8855 ^ 1'b0 ;
  assign n29433 = n27717 ^ n9762 ^ 1'b0 ;
  assign n29434 = n5222 | n29433 ;
  assign n29435 = n12228 & ~n22275 ;
  assign n29436 = n29435 ^ n1506 ^ 1'b0 ;
  assign n29437 = n27698 ^ n2779 ^ 1'b0 ;
  assign n29438 = n2148 & n13272 ;
  assign n29439 = n29438 ^ n8662 ^ 1'b0 ;
  assign n29440 = n14827 ^ n1904 ^ 1'b0 ;
  assign n29441 = n15598 ^ n9588 ^ 1'b0 ;
  assign n29442 = n6353 & ~n29441 ;
  assign n29443 = n3423 | n3957 ;
  assign n29444 = ~n29442 & n29443 ;
  assign n29445 = n23088 ^ n10752 ^ n6383 ;
  assign n29446 = n29445 ^ n17086 ^ 1'b0 ;
  assign n29447 = n5561 | n11810 ;
  assign n29448 = ~n19718 & n29447 ;
  assign n29449 = n29448 ^ n1038 ^ 1'b0 ;
  assign n29450 = ~n2076 & n8163 ;
  assign n29451 = n1201 & n29450 ;
  assign n29452 = n29451 ^ n12444 ^ 1'b0 ;
  assign n29453 = n4808 ^ n753 ^ 1'b0 ;
  assign n29454 = ~n6099 & n21073 ;
  assign n29455 = n29454 ^ n7476 ^ 1'b0 ;
  assign n29456 = n5979 & ~n8001 ;
  assign n29457 = n3840 & n29456 ;
  assign n29458 = n29457 ^ n6035 ^ 1'b0 ;
  assign n29459 = n3716 & ~n29458 ;
  assign n29460 = n1534 & ~n1571 ;
  assign n29461 = ~n1534 & n29460 ;
  assign n29462 = n29461 ^ n9670 ^ 1'b0 ;
  assign n29463 = ( n3266 & ~n15659 ) | ( n3266 & n29462 ) | ( ~n15659 & n29462 ) ;
  assign n29464 = n20759 ^ n1915 ^ 1'b0 ;
  assign n29465 = n29464 ^ n15007 ^ 1'b0 ;
  assign n29467 = n12067 ^ n10689 ^ 1'b0 ;
  assign n29468 = n4142 & ~n29467 ;
  assign n29466 = n18961 ^ n14729 ^ n2347 ;
  assign n29469 = n29468 ^ n29466 ^ 1'b0 ;
  assign n29470 = n27192 & ~n29469 ;
  assign n29471 = ~n5076 & n14637 ;
  assign n29472 = n6761 & n29471 ;
  assign n29473 = ~n29470 & n29472 ;
  assign n29474 = n162 & ~n6705 ;
  assign n29475 = n29474 ^ n428 ^ 1'b0 ;
  assign n29476 = ( n1884 & n11568 ) | ( n1884 & ~n27906 ) | ( n11568 & ~n27906 ) ;
  assign n29477 = n23067 & ~n29476 ;
  assign n29478 = n29477 ^ n24846 ^ 1'b0 ;
  assign n29479 = n11294 & n26449 ;
  assign n29480 = n29479 ^ n3962 ^ 1'b0 ;
  assign n29481 = n9788 & n10552 ;
  assign n29482 = n29481 ^ n1650 ^ 1'b0 ;
  assign n29483 = n29482 ^ n4167 ^ 1'b0 ;
  assign n29484 = n29483 ^ n11697 ^ 1'b0 ;
  assign n29485 = ~n23341 & n29484 ;
  assign n29486 = n13520 ^ n1387 ^ 1'b0 ;
  assign n29487 = n20054 | n29486 ;
  assign n29488 = n29487 ^ n5073 ^ 1'b0 ;
  assign n29489 = ~n883 & n29488 ;
  assign n29490 = n1293 ^ n1095 ^ 1'b0 ;
  assign n29491 = n29490 ^ n2670 ^ 1'b0 ;
  assign n29492 = n439 & ~n959 ;
  assign n29493 = ~n4558 & n29492 ;
  assign n29494 = n29493 ^ n5856 ^ 1'b0 ;
  assign n29495 = n29491 & ~n29494 ;
  assign n29496 = n18122 | n29495 ;
  assign n29498 = n15773 ^ n1284 ^ 1'b0 ;
  assign n29499 = n17008 & ~n29498 ;
  assign n29500 = n17863 & ~n29499 ;
  assign n29497 = n9526 | n12518 ;
  assign n29501 = n29500 ^ n29497 ^ 1'b0 ;
  assign n29502 = n23307 ^ n1705 ^ 1'b0 ;
  assign n29503 = n29502 ^ n23292 ^ 1'b0 ;
  assign n29504 = n9775 ^ n799 ^ 1'b0 ;
  assign n29505 = n18801 ^ n5168 ^ 1'b0 ;
  assign n29506 = n20179 ^ n14642 ^ 1'b0 ;
  assign n29507 = n19461 ^ n10083 ^ 1'b0 ;
  assign n29508 = n24875 | n29507 ;
  assign n29509 = n29508 ^ n12331 ^ n2358 ;
  assign n29510 = n11121 ^ n4326 ^ 1'b0 ;
  assign n29511 = ~n2186 & n11509 ;
  assign n29512 = n29511 ^ n1786 ^ 1'b0 ;
  assign n29513 = n2356 | n3906 ;
  assign n29518 = n1122 ^ n833 ^ 1'b0 ;
  assign n29519 = n5646 & ~n29518 ;
  assign n29516 = n11951 ^ n11018 ^ 1'b0 ;
  assign n29514 = n13196 ^ n12994 ^ n9508 ;
  assign n29515 = n12154 | n29514 ;
  assign n29517 = n29516 ^ n29515 ^ 1'b0 ;
  assign n29520 = n29519 ^ n29517 ^ 1'b0 ;
  assign n29521 = n29513 & n29520 ;
  assign n29522 = n28043 ^ n23997 ^ n494 ;
  assign n29523 = ~n3162 & n20313 ;
  assign n29524 = n29523 ^ n8058 ^ 1'b0 ;
  assign n29525 = n5789 & ~n13897 ;
  assign n29526 = n12149 ^ n1267 ^ 1'b0 ;
  assign n29527 = n5936 ^ n2382 ^ 1'b0 ;
  assign n29528 = n985 & ~n7329 ;
  assign n29529 = ~n7881 & n10118 ;
  assign n29530 = n29529 ^ n24496 ^ 1'b0 ;
  assign n29531 = n19518 ^ n19377 ^ 1'b0 ;
  assign n29532 = n29530 & n29531 ;
  assign n29533 = n2698 & ~n12261 ;
  assign n29534 = ~n21663 & n29533 ;
  assign n29535 = n5837 & n13251 ;
  assign n29536 = n29535 ^ n8076 ^ 1'b0 ;
  assign n29537 = n6275 ^ n17 ^ 1'b0 ;
  assign n29538 = n27952 & n29537 ;
  assign n29539 = n29538 ^ n7695 ^ 1'b0 ;
  assign n29540 = n9773 | n29539 ;
  assign n29541 = n10388 & n18525 ;
  assign n29542 = n4060 & n29541 ;
  assign n29543 = n4113 & n29542 ;
  assign n29544 = ~n4293 & n9062 ;
  assign n29545 = n14134 ^ n8039 ^ n7724 ;
  assign n29546 = n3127 | n19931 ;
  assign n29547 = n1293 & ~n2639 ;
  assign n29548 = ~n49 & n22955 ;
  assign n29549 = n29548 ^ n9943 ^ 1'b0 ;
  assign n29550 = n7209 & n29549 ;
  assign n29551 = n29547 & n29550 ;
  assign n29552 = n3571 & n26730 ;
  assign n29553 = n24446 ^ n22917 ^ 1'b0 ;
  assign n29554 = ~n12181 & n29553 ;
  assign n29555 = n23467 ^ n8480 ^ 1'b0 ;
  assign n29556 = n17012 ^ n9023 ^ 1'b0 ;
  assign n29557 = n15282 & ~n15898 ;
  assign n29558 = n29557 ^ n24266 ^ 1'b0 ;
  assign n29559 = n14471 ^ n5589 ^ 1'b0 ;
  assign n29560 = n10248 ^ n292 ^ 1'b0 ;
  assign n29564 = n741 & n1047 ;
  assign n29562 = n4277 | n23786 ;
  assign n29561 = n2668 & ~n18798 ;
  assign n29563 = n29562 ^ n29561 ^ 1'b0 ;
  assign n29565 = n29564 ^ n29563 ^ 1'b0 ;
  assign n29566 = n15777 ^ n8944 ^ 1'b0 ;
  assign n29567 = ( n124 & n20030 ) | ( n124 & ~n29566 ) | ( n20030 & ~n29566 ) ;
  assign n29568 = n11194 & ~n22083 ;
  assign n29569 = ~n4264 & n29568 ;
  assign n29570 = n29567 | n29569 ;
  assign n29571 = n29570 ^ n22448 ^ 1'b0 ;
  assign n29572 = n29571 ^ n22905 ^ 1'b0 ;
  assign n29573 = n27868 & n29572 ;
  assign n29574 = n163 & n14303 ;
  assign n29575 = n29574 ^ n24075 ^ 1'b0 ;
  assign n29576 = n4396 ^ n682 ^ 1'b0 ;
  assign n29577 = ( n1921 & n2247 ) | ( n1921 & n5658 ) | ( n2247 & n5658 ) ;
  assign n29578 = n366 & n29577 ;
  assign n29579 = n29578 ^ n22467 ^ n11858 ;
  assign n29580 = n29579 ^ n8055 ^ 1'b0 ;
  assign n29581 = n9511 | n17648 ;
  assign n29582 = n6099 | n6607 ;
  assign n29583 = n4098 & n29582 ;
  assign n29584 = n14206 ^ n12091 ^ 1'b0 ;
  assign n29585 = n3430 | n8819 ;
  assign n29586 = n6436 & n22454 ;
  assign n29587 = ~n18372 & n29586 ;
  assign n29588 = ~n2815 & n29587 ;
  assign n29589 = n29588 ^ n654 ^ 1'b0 ;
  assign n29590 = n1438 & ~n7479 ;
  assign n29591 = ( n3492 & ~n6052 ) | ( n3492 & n25300 ) | ( ~n6052 & n25300 ) ;
  assign n29592 = n29590 & n29591 ;
  assign n29593 = n29592 ^ n20992 ^ n357 ;
  assign n29594 = n5320 ^ n1770 ^ 1'b0 ;
  assign n29595 = n3455 & ~n29594 ;
  assign n29596 = n17650 & n29595 ;
  assign n29597 = ( n7530 & n22382 ) | ( n7530 & n29596 ) | ( n22382 & n29596 ) ;
  assign n29598 = n13871 & ~n16421 ;
  assign n29599 = n23272 & ~n29598 ;
  assign n29600 = n12677 & ~n22736 ;
  assign n29601 = n6256 & n29600 ;
  assign n29602 = n16482 ^ n9170 ^ 1'b0 ;
  assign n29603 = n2698 & n29602 ;
  assign n29604 = n29603 ^ n231 ^ 1'b0 ;
  assign n29605 = ~n10412 & n29604 ;
  assign n29606 = n29491 & n29605 ;
  assign n29607 = n8183 | n9949 ;
  assign n29608 = n29607 ^ n13559 ^ 1'b0 ;
  assign n29609 = n25791 & ~n29608 ;
  assign n29610 = n870 | n29609 ;
  assign n29611 = n6238 & n25546 ;
  assign n29612 = n10814 & n29611 ;
  assign n29613 = n6898 ^ n1705 ^ 1'b0 ;
  assign n29614 = n400 & ~n1461 ;
  assign n29615 = ~n400 & n29614 ;
  assign n29616 = n29615 ^ n7860 ^ 1'b0 ;
  assign n29617 = ~n24266 & n29616 ;
  assign n29618 = n24266 & n29617 ;
  assign n29619 = n7308 & ~n13404 ;
  assign n29620 = n22204 ^ n9065 ^ 1'b0 ;
  assign n29621 = ~n29619 & n29620 ;
  assign n29622 = n26098 ^ n25399 ^ 1'b0 ;
  assign n29623 = n10644 & n18912 ;
  assign n29624 = n1389 & ~n9049 ;
  assign n29625 = ~n17209 & n29624 ;
  assign n29626 = n2131 & ~n7081 ;
  assign n29627 = n20959 ^ n8714 ^ 1'b0 ;
  assign n29628 = n29627 ^ n24969 ^ n8503 ;
  assign n29629 = n29628 ^ n17415 ^ 1'b0 ;
  assign n29630 = n934 | n9579 ;
  assign n29631 = n25402 | n29630 ;
  assign n29632 = n12665 | n29631 ;
  assign n29633 = ( n4855 & n29629 ) | ( n4855 & n29632 ) | ( n29629 & n29632 ) ;
  assign n29637 = n6702 ^ n6539 ^ 1'b0 ;
  assign n29634 = n11535 & ~n17080 ;
  assign n29635 = ~n4121 & n29634 ;
  assign n29636 = n17112 & ~n29635 ;
  assign n29638 = n29637 ^ n29636 ^ 1'b0 ;
  assign n29639 = n4690 ^ n2535 ^ 1'b0 ;
  assign n29640 = ~n14863 & n29639 ;
  assign n29641 = n29640 ^ n13587 ^ 1'b0 ;
  assign n29642 = ~n19206 & n29641 ;
  assign n29643 = n2045 & ~n3465 ;
  assign n29644 = n24140 ^ n5921 ^ 1'b0 ;
  assign n29645 = ~n1556 & n29644 ;
  assign n29646 = n1207 | n17353 ;
  assign n29648 = n14979 ^ n4347 ^ 1'b0 ;
  assign n29647 = n5151 & ~n9232 ;
  assign n29649 = n29648 ^ n29647 ^ 1'b0 ;
  assign n29650 = n20856 ^ n9703 ^ 1'b0 ;
  assign n29651 = n29649 | n29650 ;
  assign n29652 = n1109 ^ n165 ^ 1'b0 ;
  assign n29653 = n29652 ^ n1570 ^ 1'b0 ;
  assign n29654 = n3166 | n19226 ;
  assign n29655 = n29654 ^ n10075 ^ 1'b0 ;
  assign n29656 = n10374 & ~n29655 ;
  assign n29657 = n29653 & n29656 ;
  assign n29658 = ( n7823 & ~n29651 ) | ( n7823 & n29657 ) | ( ~n29651 & n29657 ) ;
  assign n29659 = n21116 ^ n13664 ^ 1'b0 ;
  assign n29660 = n6950 & n22203 ;
  assign n29661 = n3823 & n29660 ;
  assign n29662 = ~n158 & n12030 ;
  assign n29663 = ~n10749 & n29662 ;
  assign n29664 = n16931 ^ n4034 ^ 1'b0 ;
  assign n29665 = n29663 | n29664 ;
  assign n29666 = ( n9427 & n11088 ) | ( n9427 & ~n29665 ) | ( n11088 & ~n29665 ) ;
  assign n29667 = n23931 ^ n14561 ^ 1'b0 ;
  assign n29669 = ~n7344 & n12488 ;
  assign n29668 = n1847 & ~n26323 ;
  assign n29670 = n29669 ^ n29668 ^ 1'b0 ;
  assign n29671 = n6442 | n26923 ;
  assign n29672 = n4252 ^ n2671 ^ 1'b0 ;
  assign n29673 = n27217 | n29672 ;
  assign n29675 = n2074 & n2130 ;
  assign n29676 = ~n1318 & n29675 ;
  assign n29674 = ~n3726 & n4022 ;
  assign n29677 = n29676 ^ n29674 ^ 1'b0 ;
  assign n29679 = n11076 ^ n2328 ^ 1'b0 ;
  assign n29680 = ~n2317 & n29679 ;
  assign n29678 = n266 & ~n9585 ;
  assign n29681 = n29680 ^ n29678 ^ 1'b0 ;
  assign n29682 = n9762 | n29681 ;
  assign n29683 = n29677 & n29682 ;
  assign n29684 = ~n15062 & n29683 ;
  assign n29685 = n11176 & ~n19835 ;
  assign n29686 = n9461 & n16146 ;
  assign n29687 = n11489 | n26324 ;
  assign n29688 = n9010 & n28348 ;
  assign n29689 = n17630 & ~n29688 ;
  assign n29690 = n12107 & ~n29689 ;
  assign n29691 = n14135 & n29690 ;
  assign n29692 = ~n1542 & n27668 ;
  assign n29693 = n20785 ^ n3981 ^ 1'b0 ;
  assign n29694 = n3558 | n29693 ;
  assign n29695 = ( n698 & n16931 ) | ( n698 & ~n29694 ) | ( n16931 & ~n29694 ) ;
  assign n29696 = n11222 & ~n29695 ;
  assign n29697 = n29696 ^ n26395 ^ 1'b0 ;
  assign n29699 = ( n12740 & n16910 ) | ( n12740 & n21460 ) | ( n16910 & n21460 ) ;
  assign n29698 = ~n6316 & n18941 ;
  assign n29700 = n29699 ^ n29698 ^ 1'b0 ;
  assign n29701 = n24653 ^ n2974 ^ 1'b0 ;
  assign n29702 = n1138 | n5010 ;
  assign n29703 = n9245 | n14183 ;
  assign n29704 = n2092 & ~n29703 ;
  assign n29705 = n29704 ^ n4376 ^ 1'b0 ;
  assign n29706 = ~n29702 & n29705 ;
  assign n29707 = n7116 ^ n6991 ^ 1'b0 ;
  assign n29708 = n11230 & ~n29707 ;
  assign n29709 = ~n746 & n23317 ;
  assign n29710 = n29709 ^ n7556 ^ 1'b0 ;
  assign n29711 = n2268 | n29710 ;
  assign n29712 = n12580 & n20146 ;
  assign n29713 = ~n24768 & n29712 ;
  assign n29714 = n3599 & ~n29713 ;
  assign n29715 = n18621 & n29714 ;
  assign n29716 = n19310 ^ n3060 ^ 1'b0 ;
  assign n29717 = ~n7718 & n29716 ;
  assign n29720 = n17712 ^ n12588 ^ 1'b0 ;
  assign n29718 = n1392 | n18069 ;
  assign n29719 = n14564 | n29718 ;
  assign n29721 = n29720 ^ n29719 ^ 1'b0 ;
  assign n29722 = n29721 ^ n12324 ^ 1'b0 ;
  assign n29723 = n3672 | n29722 ;
  assign n29729 = n3548 & ~n4095 ;
  assign n29730 = n29729 ^ n4379 ^ 1'b0 ;
  assign n29724 = n19945 & n22757 ;
  assign n29725 = n604 & n11124 ;
  assign n29726 = n1994 & n29725 ;
  assign n29727 = n2429 & ~n29726 ;
  assign n29728 = n29724 & ~n29727 ;
  assign n29731 = n29730 ^ n29728 ^ 1'b0 ;
  assign n29732 = n24790 ^ n2432 ^ 1'b0 ;
  assign n29733 = n7078 ^ n6925 ^ 1'b0 ;
  assign n29734 = ( n7057 & n10935 ) | ( n7057 & n29733 ) | ( n10935 & n29733 ) ;
  assign n29735 = n12591 ^ n9522 ^ n1052 ;
  assign n29736 = n18582 | n29735 ;
  assign n29737 = n29736 ^ n14340 ^ 1'b0 ;
  assign n29738 = n21209 & n22952 ;
  assign n29739 = ~n29737 & n29738 ;
  assign n29740 = n5940 ^ n2235 ^ 1'b0 ;
  assign n29742 = n13830 ^ n9364 ^ 1'b0 ;
  assign n29741 = n7114 & ~n15529 ;
  assign n29743 = n29742 ^ n29741 ^ 1'b0 ;
  assign n29744 = n8239 & n29743 ;
  assign n29745 = n7781 & n29744 ;
  assign n29746 = n12906 | n19780 ;
  assign n29747 = ~n12079 & n26664 ;
  assign n29748 = n29747 ^ n372 ^ 1'b0 ;
  assign n29749 = n26314 ^ n3349 ^ 1'b0 ;
  assign n29750 = n14053 & ~n29749 ;
  assign n29751 = ~n3109 & n24692 ;
  assign n29752 = n29751 ^ n20600 ^ 1'b0 ;
  assign n29753 = n28053 ^ n4081 ^ 1'b0 ;
  assign n29754 = n1014 & n29753 ;
  assign n29755 = n11212 & ~n16651 ;
  assign n29756 = n23727 ^ n18305 ^ n17333 ;
  assign n29757 = n17144 & ~n29756 ;
  assign n29758 = n5091 & n12395 ;
  assign n29759 = n29758 ^ n15406 ^ 1'b0 ;
  assign n29760 = n22671 ^ n17436 ^ 1'b0 ;
  assign n29761 = n18449 & ~n29760 ;
  assign n29762 = ( ~n2775 & n14128 ) | ( ~n2775 & n21297 ) | ( n14128 & n21297 ) ;
  assign n29763 = n1962 & n9069 ;
  assign n29764 = n15523 & ~n29763 ;
  assign n29765 = n29764 ^ n8874 ^ 1'b0 ;
  assign n29766 = n11697 & ~n26609 ;
  assign n29767 = n4666 | n13252 ;
  assign n29768 = n465 & ~n29767 ;
  assign n29769 = n13500 | n18003 ;
  assign n29770 = n29769 ^ n25581 ^ 1'b0 ;
  assign n29771 = n4005 ^ n1769 ^ 1'b0 ;
  assign n29772 = n25383 & ~n28025 ;
  assign n29773 = n1164 ^ n1062 ^ 1'b0 ;
  assign n29774 = n29773 ^ n29449 ^ 1'b0 ;
  assign n29775 = n2494 & ~n29774 ;
  assign n29776 = n2004 ^ n1000 ^ 1'b0 ;
  assign n29777 = n2966 & ~n3529 ;
  assign n29778 = n11106 | n29777 ;
  assign n29779 = n1568 | n29778 ;
  assign n29780 = ~n11007 & n29779 ;
  assign n29781 = n29780 ^ n5401 ^ 1'b0 ;
  assign n29782 = n10452 | n29781 ;
  assign n29783 = n12474 ^ n5699 ^ 1'b0 ;
  assign n29784 = n11160 & ~n29783 ;
  assign n29785 = ~n4691 & n9773 ;
  assign n29786 = n6445 & n29785 ;
  assign n29787 = n29786 ^ n2158 ^ 1'b0 ;
  assign n29788 = n29519 & ~n29787 ;
  assign n29789 = n9963 & ~n29788 ;
  assign n29791 = ~n2518 & n18228 ;
  assign n29790 = n1891 | n5982 ;
  assign n29792 = n29791 ^ n29790 ^ 1'b0 ;
  assign n29793 = n221 & ~n577 ;
  assign n29794 = n577 & n29793 ;
  assign n29795 = n1988 & n29794 ;
  assign n29796 = ~n787 & n29795 ;
  assign n29797 = n787 & n29796 ;
  assign n29798 = n631 & n9405 ;
  assign n29799 = ~n9405 & n29798 ;
  assign n29800 = ~n218 & n29799 ;
  assign n29801 = ~n1131 & n29800 ;
  assign n29802 = n1131 & n29801 ;
  assign n29803 = n692 & ~n29802 ;
  assign n29804 = n29797 & n29803 ;
  assign n29805 = n5067 & ~n29804 ;
  assign n29806 = ~n5067 & n29805 ;
  assign n29807 = n675 & n29806 ;
  assign n29808 = ( ~n6564 & n8460 ) | ( ~n6564 & n29807 ) | ( n8460 & n29807 ) ;
  assign n29809 = n26298 ^ n18615 ^ 1'b0 ;
  assign n29810 = n29808 | n29809 ;
  assign n29811 = n12364 ^ n968 ^ 1'b0 ;
  assign n29812 = ~n29810 & n29811 ;
  assign n29813 = n29812 ^ n7919 ^ 1'b0 ;
  assign n29814 = n9542 & ~n21395 ;
  assign n29815 = ~n4916 & n23054 ;
  assign n29816 = n3518 & ~n4131 ;
  assign n29817 = n2438 & n29816 ;
  assign n29819 = n5246 & ~n9929 ;
  assign n29820 = n107 & n29819 ;
  assign n29818 = n3469 & n15424 ;
  assign n29821 = n29820 ^ n29818 ^ 1'b0 ;
  assign n29822 = n5016 | n5668 ;
  assign n29825 = n4700 & ~n11865 ;
  assign n29826 = ~n23 & n29825 ;
  assign n29823 = ( n482 & ~n13481 ) | ( n482 & n21221 ) | ( ~n13481 & n21221 ) ;
  assign n29824 = ~n14536 & n29823 ;
  assign n29827 = n29826 ^ n29824 ^ 1'b0 ;
  assign n29828 = n17201 | n29827 ;
  assign n29829 = n225 & n4544 ;
  assign n29830 = n29829 ^ n27929 ^ 1'b0 ;
  assign n29831 = ~n12217 & n26107 ;
  assign n29832 = n20304 ^ n4005 ^ n2902 ;
  assign n29833 = ~n22709 & n29832 ;
  assign n29834 = n8494 | n8961 ;
  assign n29835 = ~n16656 & n22895 ;
  assign n29836 = ~n29834 & n29835 ;
  assign n29837 = n14832 | n26715 ;
  assign n29838 = n13597 ^ n2864 ^ 1'b0 ;
  assign n29839 = n16136 & ~n17769 ;
  assign n29840 = n1534 & n29839 ;
  assign n29841 = n29840 ^ n22262 ^ 1'b0 ;
  assign n29842 = ~n2421 & n2883 ;
  assign n29843 = n15413 & n29842 ;
  assign n29844 = n466 & n1154 ;
  assign n29845 = ~n1958 & n27569 ;
  assign n29846 = ( n934 & n1900 ) | ( n934 & ~n9286 ) | ( n1900 & ~n9286 ) ;
  assign n29847 = n29846 ^ n774 ^ 1'b0 ;
  assign n29848 = ~n11047 & n16280 ;
  assign n29849 = n29847 | n29848 ;
  assign n29850 = n1741 & ~n29849 ;
  assign n29851 = n29823 ^ n6646 ^ 1'b0 ;
  assign n29853 = n2628 ^ n402 ^ 1'b0 ;
  assign n29854 = n3082 & n29853 ;
  assign n29852 = n5738 & n27959 ;
  assign n29855 = n29854 ^ n29852 ^ 1'b0 ;
  assign n29856 = n19399 ^ n13520 ^ 1'b0 ;
  assign n29857 = ~n12197 & n29856 ;
  assign n29858 = ~n796 & n29857 ;
  assign n29859 = n29858 ^ n7994 ^ 1'b0 ;
  assign n29860 = n1340 | n9929 ;
  assign n29861 = n29860 ^ n28960 ^ 1'b0 ;
  assign n29862 = n14905 ^ n5610 ^ n510 ;
  assign n29863 = n5357 & n6292 ;
  assign n29864 = n2900 & n29296 ;
  assign n29865 = ~n12786 & n29864 ;
  assign n29866 = n19831 & n29704 ;
  assign n29867 = n27834 ^ n5681 ^ 1'b0 ;
  assign n29868 = ( n1211 & n13939 ) | ( n1211 & ~n29867 ) | ( n13939 & ~n29867 ) ;
  assign n29869 = n6297 & ~n25101 ;
  assign n29870 = n15207 ^ n5616 ^ 1'b0 ;
  assign n29871 = n13388 | n29870 ;
  assign n29872 = n4313 & ~n6235 ;
  assign n29873 = n2586 | n20833 ;
  assign n29874 = n29873 ^ n26767 ^ 1'b0 ;
  assign n29875 = n152 & ~n6600 ;
  assign n29876 = n1523 & n29875 ;
  assign n29877 = n24208 ^ n8683 ^ 1'b0 ;
  assign n29879 = n20547 ^ n15206 ^ n7262 ;
  assign n29878 = n15697 | n18343 ;
  assign n29880 = n29879 ^ n29878 ^ 1'b0 ;
  assign n29881 = ~n133 & n2678 ;
  assign n29882 = n24953 & ~n27109 ;
  assign n29883 = n29882 ^ n3061 ^ 1'b0 ;
  assign n29884 = n12197 ^ n225 ^ 1'b0 ;
  assign n29885 = n12990 & n29884 ;
  assign n29886 = n29885 ^ n12479 ^ n892 ;
  assign n29887 = n2684 | n20230 ;
  assign n29888 = n24583 ^ n23767 ^ 1'b0 ;
  assign n29889 = n26647 ^ n11251 ^ 1'b0 ;
  assign n29890 = n27839 ^ n1439 ^ 1'b0 ;
  assign n29891 = n2769 ^ x5 ^ 1'b0 ;
  assign n29892 = n11305 ^ n6696 ^ 1'b0 ;
  assign n29893 = n29891 & ~n29892 ;
  assign n29894 = ~n16023 & n29893 ;
  assign n29895 = ~n5041 & n7091 ;
  assign n29896 = n29895 ^ n3359 ^ 1'b0 ;
  assign n29897 = n29896 ^ n6827 ^ 1'b0 ;
  assign n29898 = ~n25310 & n29897 ;
  assign n29899 = n22214 ^ n2545 ^ 1'b0 ;
  assign n29900 = n3983 | n5552 ;
  assign n29901 = n29900 ^ n403 ^ 1'b0 ;
  assign n29902 = n26825 ^ n25640 ^ 1'b0 ;
  assign n29903 = n4408 ^ n1426 ^ 1'b0 ;
  assign n29904 = n8760 & ~n29903 ;
  assign n29905 = n9085 ^ n61 ^ 1'b0 ;
  assign n29906 = n3003 & n29905 ;
  assign n29907 = n29906 ^ n4006 ^ 1'b0 ;
  assign n29908 = n27009 ^ n20048 ^ 1'b0 ;
  assign n29909 = n16527 | n29908 ;
  assign n29910 = n29907 & n29909 ;
  assign n29911 = ( ~n6935 & n29904 ) | ( ~n6935 & n29910 ) | ( n29904 & n29910 ) ;
  assign n29912 = n8163 ^ n3032 ^ 1'b0 ;
  assign n29913 = n9194 | n11846 ;
  assign n29914 = n29913 ^ n25241 ^ 1'b0 ;
  assign n29915 = n20457 ^ n5027 ^ 1'b0 ;
  assign n29916 = n1548 & n21264 ;
  assign n29917 = n29916 ^ n12125 ^ 1'b0 ;
  assign n29918 = n667 & n29917 ;
  assign n29919 = n19879 & ~n23770 ;
  assign n29920 = n5741 ^ n535 ^ 1'b0 ;
  assign n29921 = n4208 & n29920 ;
  assign n29922 = n20559 ^ n20268 ^ 1'b0 ;
  assign n29923 = n21228 ^ n17157 ^ 1'b0 ;
  assign n29924 = n3406 | n29923 ;
  assign n29925 = n2232 | n29924 ;
  assign n29926 = n11841 & n20362 ;
  assign n29927 = n16947 ^ n9203 ^ 1'b0 ;
  assign n29928 = n21868 & ~n29927 ;
  assign n29929 = n28605 & n29928 ;
  assign n29930 = ~n4056 & n19360 ;
  assign n29931 = n29930 ^ n3705 ^ 1'b0 ;
  assign n29932 = ~n223 & n4331 ;
  assign n29933 = ( ~n12179 & n13118 ) | ( ~n12179 & n29932 ) | ( n13118 & n29932 ) ;
  assign n29934 = n6645 & n29933 ;
  assign n29935 = n10368 & n29934 ;
  assign n29937 = n12579 ^ n1510 ^ 1'b0 ;
  assign n29936 = n17878 ^ n2337 ^ 1'b0 ;
  assign n29938 = n29937 ^ n29936 ^ n423 ;
  assign n29939 = n3102 | n12740 ;
  assign n29940 = n29939 ^ n18445 ^ n3080 ;
  assign n29941 = n25562 ^ n3082 ^ 1'b0 ;
  assign n29942 = n5036 & ~n26787 ;
  assign n29943 = n29942 ^ n16079 ^ n2399 ;
  assign n29944 = n4506 & ~n21545 ;
  assign n29945 = ~n20285 & n29944 ;
  assign n29946 = n4341 ^ n3279 ^ 1'b0 ;
  assign n29947 = n29945 | n29946 ;
  assign n29948 = n4525 & ~n5672 ;
  assign n29949 = n29948 ^ n1841 ^ 1'b0 ;
  assign n29950 = n4301 | n29949 ;
  assign n29951 = n10656 & n29950 ;
  assign n29953 = n56 & ~n10438 ;
  assign n29954 = n10438 & n29953 ;
  assign n29952 = n1929 & ~n7953 ;
  assign n29955 = n29954 ^ n29952 ^ 1'b0 ;
  assign n29956 = n29955 ^ n16252 ^ n704 ;
  assign n29957 = n12901 | n19173 ;
  assign n29958 = n29957 ^ n20617 ^ n13939 ;
  assign n29959 = n25047 ^ n1109 ^ 1'b0 ;
  assign n29960 = n19973 & ~n29959 ;
  assign n29961 = n8105 ^ n6498 ^ 1'b0 ;
  assign n29962 = n2284 & ~n4398 ;
  assign n29963 = n10403 & n29962 ;
  assign n29964 = n29963 ^ n16116 ^ 1'b0 ;
  assign n29965 = n18458 & n29964 ;
  assign n29967 = n14207 ^ n1407 ^ 1'b0 ;
  assign n29968 = n12144 & n29967 ;
  assign n29969 = n14123 & n29968 ;
  assign n29966 = n9857 & n19193 ;
  assign n29970 = n29969 ^ n29966 ^ 1'b0 ;
  assign n29971 = n7467 | n25763 ;
  assign n29972 = n8771 ^ n6633 ^ 1'b0 ;
  assign n29973 = n13557 & n29819 ;
  assign n29974 = n8874 & ~n9617 ;
  assign n29975 = n29974 ^ n1663 ^ 1'b0 ;
  assign n29976 = n29975 ^ n5897 ^ n4960 ;
  assign n29977 = n24415 ^ n2262 ^ 1'b0 ;
  assign n29978 = ~n18936 & n29977 ;
  assign n29979 = n29976 & n29978 ;
  assign n29980 = ~n2248 & n29645 ;
  assign n29981 = n5973 & ~n6370 ;
  assign n29982 = n16026 & ~n29981 ;
  assign n29983 = n2192 & ~n7360 ;
  assign n29984 = n29983 ^ n24664 ^ 1'b0 ;
  assign n29985 = n24973 ^ n4712 ^ 1'b0 ;
  assign n29986 = ~n12642 & n14937 ;
  assign n29987 = n16670 ^ n1276 ^ 1'b0 ;
  assign n29988 = n29987 ^ n23715 ^ 1'b0 ;
  assign n29989 = n29988 ^ n28060 ^ 1'b0 ;
  assign n29990 = n17314 ^ n11150 ^ 1'b0 ;
  assign n29991 = ~n16974 & n21235 ;
  assign n29992 = ~n27636 & n29991 ;
  assign n29993 = n14244 ^ n10345 ^ 1'b0 ;
  assign n29994 = n24380 ^ n220 ^ 1'b0 ;
  assign n29995 = n29993 | n29994 ;
  assign n29996 = n6878 ^ n5286 ^ 1'b0 ;
  assign n29997 = n15009 & ~n29996 ;
  assign n29998 = n29997 ^ n4180 ^ 1'b0 ;
  assign n29999 = ~n29995 & n29998 ;
  assign n30002 = n18031 ^ n9657 ^ 1'b0 ;
  assign n30003 = n18616 & n30002 ;
  assign n30000 = ( n10740 & ~n12046 ) | ( n10740 & n14667 ) | ( ~n12046 & n14667 ) ;
  assign n30001 = ~n10129 & n30000 ;
  assign n30004 = n30003 ^ n30001 ^ 1'b0 ;
  assign n30005 = n6804 | n30004 ;
  assign n30006 = n7463 & ~n30005 ;
  assign n30007 = n7916 & n8391 ;
  assign n30008 = ~n5823 & n30007 ;
  assign n30009 = n8860 & ~n30008 ;
  assign n30010 = ~n11164 & n30009 ;
  assign n30011 = n2923 & ~n18662 ;
  assign n30012 = n17702 ^ n5663 ^ 1'b0 ;
  assign n30013 = n14200 & ~n14577 ;
  assign n30014 = ~n26511 & n30013 ;
  assign n30015 = n15213 & n30014 ;
  assign n30016 = n12013 ^ n9148 ^ 1'b0 ;
  assign n30017 = n30016 ^ n23264 ^ 1'b0 ;
  assign n30018 = n30017 ^ n21868 ^ n17220 ;
  assign n30019 = ( ~n20927 & n28335 ) | ( ~n20927 & n30018 ) | ( n28335 & n30018 ) ;
  assign n30020 = ~n21811 & n29997 ;
  assign n30021 = n22671 ^ n5183 ^ 1'b0 ;
  assign n30022 = n14353 & ~n29935 ;
  assign n30023 = n263 & n12502 ;
  assign n30024 = n1726 & ~n21427 ;
  assign n30025 = n30024 ^ n19931 ^ 1'b0 ;
  assign n30026 = ~n14343 & n14802 ;
  assign n30027 = n30026 ^ n4832 ^ 1'b0 ;
  assign n30028 = n2991 & ~n7109 ;
  assign n30029 = n30028 ^ n20400 ^ 1'b0 ;
  assign n30030 = n6467 & n11583 ;
  assign n30031 = ~n2634 & n4143 ;
  assign n30032 = ~n30030 & n30031 ;
  assign n30033 = n20157 | n29101 ;
  assign n30036 = ~n213 & n5184 ;
  assign n30037 = n5294 & n30036 ;
  assign n30038 = n30037 ^ n20489 ^ 1'b0 ;
  assign n30034 = ( n9583 & n15822 ) | ( n9583 & ~n24848 ) | ( n15822 & ~n24848 ) ;
  assign n30035 = n28211 & n30034 ;
  assign n30039 = n30038 ^ n30035 ^ 1'b0 ;
  assign n30040 = ~n10463 & n27263 ;
  assign n30041 = ~n18051 & n30040 ;
  assign n30042 = n4419 & ~n9946 ;
  assign n30043 = n2719 & n30042 ;
  assign n30044 = n30043 ^ n2556 ^ 1'b0 ;
  assign n30045 = n9009 | n30044 ;
  assign n30046 = n30041 | n30045 ;
  assign n30047 = ( n7197 & n18944 ) | ( n7197 & n30046 ) | ( n18944 & n30046 ) ;
  assign n30048 = n7999 | n15561 ;
  assign n30049 = n30048 ^ n3126 ^ 1'b0 ;
  assign n30050 = n30049 ^ n982 ^ 1'b0 ;
  assign n30051 = n15803 | n16829 ;
  assign n30052 = n30051 ^ n19934 ^ 1'b0 ;
  assign n30053 = n28391 | n30052 ;
  assign n30054 = n269 | n792 ;
  assign n30055 = n2202 | n30054 ;
  assign n30056 = n23286 ^ n6556 ^ 1'b0 ;
  assign n30057 = ~n1985 & n30056 ;
  assign n30058 = n4508 & ~n5190 ;
  assign n30059 = ~n365 & n30058 ;
  assign n30060 = n14994 ^ n5514 ^ 1'b0 ;
  assign n30061 = n3392 & n30060 ;
  assign n30062 = n30061 ^ n2771 ^ 1'b0 ;
  assign n30063 = n30059 | n30062 ;
  assign n30064 = n10235 | n18821 ;
  assign n30065 = n30063 & ~n30064 ;
  assign n30066 = n315 & ~n2874 ;
  assign n30067 = ~n15299 & n30066 ;
  assign n30068 = n23915 ^ n4345 ^ 1'b0 ;
  assign n30069 = n10369 | n30068 ;
  assign n30070 = n8500 | n30069 ;
  assign n30071 = n30070 ^ n5867 ^ 1'b0 ;
  assign n30072 = ~n21031 & n30071 ;
  assign n30073 = ( ~n9555 & n30067 ) | ( ~n9555 & n30072 ) | ( n30067 & n30072 ) ;
  assign n30074 = n26740 | n26805 ;
  assign n30075 = n1721 & ~n8662 ;
  assign n30076 = n30075 ^ n2034 ^ 1'b0 ;
  assign n30077 = n2424 & n10069 ;
  assign n30078 = ~n7948 & n12980 ;
  assign n30079 = n30077 & n30078 ;
  assign n30080 = n625 & n6464 ;
  assign n30081 = n30080 ^ n10703 ^ 1'b0 ;
  assign n30082 = n6846 | n7947 ;
  assign n30083 = n26298 | n30082 ;
  assign n30084 = n8233 ^ n1978 ^ 1'b0 ;
  assign n30085 = n9033 & n12015 ;
  assign n30086 = n25208 & n30085 ;
  assign n30087 = ~n918 & n22389 ;
  assign n30088 = n30087 ^ n3584 ^ 1'b0 ;
  assign n30089 = n3949 ^ n3445 ^ 1'b0 ;
  assign n30090 = n9022 & n30089 ;
  assign n30091 = n26719 ^ n5385 ^ 1'b0 ;
  assign n30092 = n9312 & ~n30091 ;
  assign n30093 = n3235 & ~n7567 ;
  assign n30094 = n29702 & n30093 ;
  assign n30095 = n24743 & n30094 ;
  assign n30096 = n22545 ^ n13540 ^ 1'b0 ;
  assign n30097 = ~n28278 & n30096 ;
  assign n30098 = n7308 & ~n17025 ;
  assign n30099 = n30098 ^ n704 ^ 1'b0 ;
  assign n30100 = n9963 ^ n4683 ^ 1'b0 ;
  assign n30101 = n725 & n30100 ;
  assign n30102 = ~n11994 & n30101 ;
  assign n30103 = n6023 | n9983 ;
  assign n30104 = n30103 ^ n14253 ^ 1'b0 ;
  assign n30105 = n30102 & ~n30104 ;
  assign n30106 = n30105 ^ n14057 ^ n4328 ;
  assign n30107 = n11911 ^ n6978 ^ 1'b0 ;
  assign n30108 = n30107 ^ n12423 ^ 1'b0 ;
  assign n30109 = n5988 | n23176 ;
  assign n30110 = n24489 | n30109 ;
  assign n30111 = n806 & ~n3885 ;
  assign n30112 = ( n423 & ~n14305 ) | ( n423 & n30111 ) | ( ~n14305 & n30111 ) ;
  assign n30113 = n5262 & ~n17711 ;
  assign n30114 = ~n19129 & n29499 ;
  assign n30115 = ~n30113 & n30114 ;
  assign n30116 = n30115 ^ n22969 ^ 1'b0 ;
  assign n30117 = n9925 | n30116 ;
  assign n30118 = n6156 & ~n26556 ;
  assign n30122 = n6224 ^ n5728 ^ 1'b0 ;
  assign n30119 = n22697 ^ n1603 ^ 1'b0 ;
  assign n30120 = n23112 & n30119 ;
  assign n30121 = n30120 ^ n1312 ^ 1'b0 ;
  assign n30123 = n30122 ^ n30121 ^ 1'b0 ;
  assign n30124 = n1574 | n22128 ;
  assign n30125 = n26369 ^ n8730 ^ 1'b0 ;
  assign n30126 = n30125 ^ n6912 ^ 1'b0 ;
  assign n30127 = ( n8476 & ~n10828 ) | ( n8476 & n12860 ) | ( ~n10828 & n12860 ) ;
  assign n30128 = n21926 & ~n30127 ;
  assign n30129 = n14570 ^ n6479 ^ n2851 ;
  assign n30130 = n2038 | n30129 ;
  assign n30131 = n3449 | n7413 ;
  assign n30132 = ~n14558 & n28618 ;
  assign n30133 = n7893 ^ n2284 ^ 1'b0 ;
  assign n30134 = n9651 & ~n30133 ;
  assign n30135 = n19203 & n30134 ;
  assign n30136 = ~n5872 & n30135 ;
  assign n30137 = n12376 ^ n9332 ^ 1'b0 ;
  assign n30138 = n2953 & ~n23790 ;
  assign n30139 = n1157 & n8646 ;
  assign n30140 = n30139 ^ n22791 ^ 1'b0 ;
  assign n30141 = n600 & ~n11066 ;
  assign n30142 = n30140 & n30141 ;
  assign n30143 = ~n25785 & n30142 ;
  assign n30144 = n12187 & ~n30143 ;
  assign n30145 = ~n4976 & n11704 ;
  assign n30146 = n19658 & ~n30145 ;
  assign n30147 = n8099 ^ n863 ^ 1'b0 ;
  assign n30148 = n14665 & ~n30147 ;
  assign n30149 = n10256 & n22382 ;
  assign n30150 = ( n25629 & n30148 ) | ( n25629 & n30149 ) | ( n30148 & n30149 ) ;
  assign n30151 = ~n4593 & n5921 ;
  assign n30152 = n30151 ^ n26169 ^ 1'b0 ;
  assign n30153 = n23558 ^ n13238 ^ 1'b0 ;
  assign n30154 = ~n61 & n30153 ;
  assign n30155 = n30154 ^ n17829 ^ 1'b0 ;
  assign n30156 = n8557 | n15934 ;
  assign n30157 = n15426 & ~n30156 ;
  assign n30158 = n3955 & ~n5912 ;
  assign n30159 = n5422 ^ n4670 ^ 1'b0 ;
  assign n30160 = n30158 | n30159 ;
  assign n30161 = n11039 ^ n7386 ^ 1'b0 ;
  assign n30162 = ~n11964 & n30161 ;
  assign n30163 = n13018 ^ n6925 ^ 1'b0 ;
  assign n30164 = n30162 & ~n30163 ;
  assign n30165 = n30160 & n30164 ;
  assign n30166 = n7590 | n19595 ;
  assign n30167 = ~n4884 & n30166 ;
  assign n30168 = n24860 ^ n609 ^ 1'b0 ;
  assign n30169 = n13136 ^ n5974 ^ 1'b0 ;
  assign n30170 = ~n17420 & n19629 ;
  assign n30171 = n11068 ^ n3940 ^ 1'b0 ;
  assign n30172 = n7948 | n30171 ;
  assign n30173 = n7476 & n9036 ;
  assign n30174 = n30173 ^ n11978 ^ 1'b0 ;
  assign n30175 = n30172 | n30174 ;
  assign n30176 = n24543 ^ n2833 ^ 1'b0 ;
  assign n30177 = n2279 | n8070 ;
  assign n30178 = n7778 | n23354 ;
  assign n30179 = ~n21139 & n30178 ;
  assign n30180 = n14212 ^ n2623 ^ 1'b0 ;
  assign n30181 = ( n2632 & ~n8689 ) | ( n2632 & n17142 ) | ( ~n8689 & n17142 ) ;
  assign n30182 = ~n16701 & n30181 ;
  assign n30183 = ~n7124 & n29035 ;
  assign n30184 = n30183 ^ n23149 ^ 1'b0 ;
  assign n30185 = n16004 | n20455 ;
  assign n30186 = n17563 & ~n30185 ;
  assign n30189 = n6898 ^ n3917 ^ 1'b0 ;
  assign n30187 = n19537 ^ n2461 ^ 1'b0 ;
  assign n30188 = n14226 & ~n30187 ;
  assign n30190 = n30189 ^ n30188 ^ 1'b0 ;
  assign n30192 = n3006 & ~n4870 ;
  assign n30193 = n17604 & n30192 ;
  assign n30194 = n30193 ^ n5067 ^ 1'b0 ;
  assign n30191 = n362 & n2398 ;
  assign n30195 = n30194 ^ n30191 ^ 1'b0 ;
  assign n30196 = ~n6234 & n6272 ;
  assign n30197 = n30196 ^ n40 ^ 1'b0 ;
  assign n30198 = n3052 & ~n18382 ;
  assign n30199 = n14558 ^ n3013 ^ 1'b0 ;
  assign n30200 = n26 | n30199 ;
  assign n30201 = n11771 | n30200 ;
  assign n30202 = n9361 & ~n30201 ;
  assign n30203 = n19153 ^ n5491 ^ 1'b0 ;
  assign n30204 = ( n4951 & n15023 ) | ( n4951 & n24155 ) | ( n15023 & n24155 ) ;
  assign n30205 = ~n10171 & n13351 ;
  assign n30206 = n22986 ^ n11772 ^ 1'b0 ;
  assign n30207 = ~n536 & n30206 ;
  assign n30208 = ~n27209 & n30207 ;
  assign n30209 = n30205 & n30208 ;
  assign n30210 = n1196 & ~n8939 ;
  assign n30211 = n15054 & ~n30210 ;
  assign n30212 = n28968 & n30211 ;
  assign n30213 = n27668 & ~n30212 ;
  assign n30214 = n6690 ^ n5273 ^ 1'b0 ;
  assign n30215 = ~n7955 & n30214 ;
  assign n30216 = n30215 ^ n20433 ^ 1'b0 ;
  assign n30217 = n6128 & ~n30216 ;
  assign n30218 = n4174 ^ n2749 ^ 1'b0 ;
  assign n30219 = ~n13673 & n30218 ;
  assign n30220 = n30219 ^ n16909 ^ 1'b0 ;
  assign n30221 = n25794 ^ n18961 ^ n8712 ;
  assign n30222 = n22161 & n26530 ;
  assign n30223 = n10083 & n13699 ;
  assign n30224 = n19059 ^ n16325 ^ 1'b0 ;
  assign n30225 = n10462 & n30224 ;
  assign n30226 = n30225 ^ n15092 ^ 1'b0 ;
  assign n30227 = n18411 & ~n20552 ;
  assign n30228 = n11122 & n30227 ;
  assign n30229 = n12718 & n14489 ;
  assign n30230 = ~n14489 & n30229 ;
  assign n30231 = n659 | n22835 ;
  assign n30232 = n3207 & ~n16331 ;
  assign n30233 = n16331 & n30232 ;
  assign n30234 = ~n4834 & n16577 ;
  assign n30235 = n30233 & n30234 ;
  assign n30236 = n30235 ^ n428 ^ 1'b0 ;
  assign n30237 = n30231 & ~n30236 ;
  assign n30238 = n30237 ^ n30103 ^ 1'b0 ;
  assign n30239 = n3899 & ~n12932 ;
  assign n30240 = n588 ^ n248 ^ 1'b0 ;
  assign n30241 = n12299 & n30240 ;
  assign n30242 = n30239 | n30241 ;
  assign n30243 = n23556 ^ n7990 ^ 1'b0 ;
  assign n30244 = n957 & n11193 ;
  assign n30245 = n10424 & n11737 ;
  assign n30246 = n8390 ^ n2388 ^ 1'b0 ;
  assign n30247 = n30245 & n30246 ;
  assign n30248 = n14156 | n25307 ;
  assign n30249 = n30248 ^ n3147 ^ n522 ;
  assign n30250 = n16691 & ~n30249 ;
  assign n30251 = n30250 ^ n3790 ^ 1'b0 ;
  assign n30252 = n482 & n10756 ;
  assign n30253 = n8020 & n30252 ;
  assign n30254 = n30253 ^ n25732 ^ 1'b0 ;
  assign n30255 = n30254 ^ n18575 ^ n3817 ;
  assign n30256 = n28 & n1246 ;
  assign n30257 = n10497 ^ n229 ^ 1'b0 ;
  assign n30258 = n3760 | n30257 ;
  assign n30259 = n30256 & n30258 ;
  assign n30260 = n21251 | n30259 ;
  assign n30261 = n16762 & n21792 ;
  assign n30262 = ~n13061 & n30261 ;
  assign n30263 = n30262 ^ n10185 ^ 1'b0 ;
  assign n30264 = n7010 & n30263 ;
  assign n30265 = n23880 ^ n12320 ^ 1'b0 ;
  assign n30266 = ~n16613 & n22344 ;
  assign n30267 = n30266 ^ n22501 ^ 1'b0 ;
  assign n30269 = n18191 ^ n7735 ^ 1'b0 ;
  assign n30268 = n20904 | n24580 ;
  assign n30270 = n30269 ^ n30268 ^ 1'b0 ;
  assign n30271 = ~n5956 & n8906 ;
  assign n30272 = ~n9178 & n30271 ;
  assign n30273 = n30272 ^ n4681 ^ 1'b0 ;
  assign n30274 = n22496 ^ n9985 ^ 1'b0 ;
  assign n30275 = n7459 ^ n2872 ^ 1'b0 ;
  assign n30276 = n841 & n30275 ;
  assign n30277 = n4975 & n30276 ;
  assign n30278 = ~n133 & n30277 ;
  assign n30279 = n10041 ^ n4681 ^ 1'b0 ;
  assign n30280 = ~n15944 & n20034 ;
  assign n30281 = n30280 ^ n5979 ^ 1'b0 ;
  assign n30282 = n6358 | n11499 ;
  assign n30283 = ~n23593 & n26747 ;
  assign n30284 = ~n30282 & n30283 ;
  assign n30285 = n23142 ^ n5217 ^ 1'b0 ;
  assign n30286 = n19937 | n27758 ;
  assign n30287 = n30286 ^ n17162 ^ 1'b0 ;
  assign n30289 = n3798 | n10544 ;
  assign n30288 = n13826 ^ n10449 ^ 1'b0 ;
  assign n30290 = n30289 ^ n30288 ^ n25989 ;
  assign n30291 = n26712 ^ n3514 ^ 1'b0 ;
  assign n30292 = ~n9045 & n30291 ;
  assign n30293 = n27117 ^ n15742 ^ 1'b0 ;
  assign n30294 = n15299 | n27566 ;
  assign n30297 = ~n8032 & n23766 ;
  assign n30298 = ( n9542 & n15025 ) | ( n9542 & ~n30297 ) | ( n15025 & ~n30297 ) ;
  assign n30295 = n12757 & n13287 ;
  assign n30296 = ~n24317 & n30295 ;
  assign n30299 = n30298 ^ n30296 ^ 1'b0 ;
  assign n30300 = n6736 ^ n3670 ^ 1'b0 ;
  assign n30301 = ~n4024 & n30300 ;
  assign n30302 = ( n663 & ~n1385 ) | ( n663 & n4193 ) | ( ~n1385 & n4193 ) ;
  assign n30303 = n30302 ^ n3974 ^ 1'b0 ;
  assign n30304 = n20287 & n30303 ;
  assign n30305 = n6164 & ~n10119 ;
  assign n30306 = n30305 ^ n25747 ^ 1'b0 ;
  assign n30307 = n19772 | n30306 ;
  assign n30308 = n30307 ^ n85 ^ 1'b0 ;
  assign n30309 = ~n3044 & n9770 ;
  assign n30310 = ~n8573 & n30309 ;
  assign n30311 = ~n1688 & n30310 ;
  assign n30312 = n21439 ^ n9043 ^ 1'b0 ;
  assign n30313 = ~n30311 & n30312 ;
  assign n30314 = n30313 ^ n2085 ^ 1'b0 ;
  assign n30315 = n16972 ^ n13578 ^ 1'b0 ;
  assign n30316 = ~n714 & n1323 ;
  assign n30317 = n30316 ^ n14434 ^ 1'b0 ;
  assign n30318 = n15662 ^ n10083 ^ n9768 ;
  assign n30319 = ~n18062 & n30318 ;
  assign n30320 = n15211 ^ n5227 ^ n3280 ;
  assign n30321 = n3058 & n4007 ;
  assign n30322 = ~n579 & n30321 ;
  assign n30323 = n3414 & ~n30322 ;
  assign n30324 = n30320 & n30323 ;
  assign n30325 = ~n14301 & n27485 ;
  assign n30326 = n16245 & n30325 ;
  assign n30327 = n24667 ^ n5651 ^ 1'b0 ;
  assign n30328 = n8933 & n30327 ;
  assign n30329 = ( ~n1325 & n22791 ) | ( ~n1325 & n30328 ) | ( n22791 & n30328 ) ;
  assign n30330 = n5001 & ~n15155 ;
  assign n30331 = ~n366 & n19394 ;
  assign n30332 = ~n2014 & n30331 ;
  assign n30333 = n7744 & ~n19515 ;
  assign n30334 = n732 | n29283 ;
  assign n30335 = n22761 & ~n30334 ;
  assign n30336 = ( n1383 & ~n5520 ) | ( n1383 & n22959 ) | ( ~n5520 & n22959 ) ;
  assign n30337 = n30336 ^ n10724 ^ 1'b0 ;
  assign n30338 = n12433 & ~n30337 ;
  assign n30339 = n5217 & n10031 ;
  assign n30340 = n30339 ^ n290 ^ 1'b0 ;
  assign n30341 = n30340 ^ n2961 ^ 1'b0 ;
  assign n30342 = ( n2439 & ~n30338 ) | ( n2439 & n30341 ) | ( ~n30338 & n30341 ) ;
  assign n30343 = ~n1908 & n20496 ;
  assign n30344 = n1857 & ~n8731 ;
  assign n30345 = ~n545 & n30344 ;
  assign n30346 = n8381 | n30345 ;
  assign n30347 = n14687 ^ n1396 ^ n545 ;
  assign n30348 = n1688 | n9886 ;
  assign n30349 = n30348 ^ n6065 ^ 1'b0 ;
  assign n30350 = n30349 ^ n20037 ^ 1'b0 ;
  assign n30351 = ( n4267 & n30347 ) | ( n4267 & n30350 ) | ( n30347 & n30350 ) ;
  assign n30352 = ~n577 & n855 ;
  assign n30353 = n30352 ^ x8 ^ 1'b0 ;
  assign n30354 = ( n7832 & n11386 ) | ( n7832 & ~n21902 ) | ( n11386 & ~n21902 ) ;
  assign n30355 = n692 & ~n30354 ;
  assign n30356 = n30355 ^ n28122 ^ 1'b0 ;
  assign n30357 = n9216 & n16599 ;
  assign n30358 = n19281 ^ n11860 ^ 1'b0 ;
  assign n30359 = n30357 & n30358 ;
  assign n30360 = n30359 ^ n2327 ^ 1'b0 ;
  assign n30361 = n7930 ^ n485 ^ 1'b0 ;
  assign n30362 = n15479 | n30361 ;
  assign n30363 = n13547 & n18373 ;
  assign n30364 = ~n17044 & n30363 ;
  assign n30365 = n14431 ^ n7546 ^ 1'b0 ;
  assign n30366 = n11768 & n30365 ;
  assign n30367 = n3968 | n9542 ;
  assign n30368 = n19191 & n30367 ;
  assign n30369 = n21674 & n30368 ;
  assign n30370 = n26472 ^ n21515 ^ 1'b0 ;
  assign n30371 = n30370 ^ n17649 ^ 1'b0 ;
  assign n30372 = ( n12692 & n20669 ) | ( n12692 & ~n30371 ) | ( n20669 & ~n30371 ) ;
  assign n30373 = n7639 & n11146 ;
  assign n30374 = n9215 ^ n4218 ^ 1'b0 ;
  assign n30375 = n30373 & n30374 ;
  assign n30376 = n9072 | n19338 ;
  assign n30377 = n4395 | n30376 ;
  assign n30378 = n6126 ^ n4145 ^ 1'b0 ;
  assign n30379 = n7688 & n30378 ;
  assign n30380 = n30379 ^ n10463 ^ 1'b0 ;
  assign n30381 = n13086 ^ n1408 ^ 1'b0 ;
  assign n30382 = n30380 & ~n30381 ;
  assign n30383 = n12185 & ~n22040 ;
  assign n30384 = n17420 & n26589 ;
  assign n30385 = ( n6655 & ~n7490 ) | ( n6655 & n15792 ) | ( ~n7490 & n15792 ) ;
  assign n30387 = n4123 | n11858 ;
  assign n30388 = n3078 & ~n30387 ;
  assign n30389 = n1469 | n30388 ;
  assign n30386 = ~n10182 & n17887 ;
  assign n30390 = n30389 ^ n30386 ^ 1'b0 ;
  assign n30391 = n19808 & ~n24928 ;
  assign n30392 = n8073 | n16809 ;
  assign n30393 = n30391 & ~n30392 ;
  assign n30394 = n27018 ^ n3461 ^ 1'b0 ;
  assign n30395 = ~n27976 & n30394 ;
  assign n30396 = n19245 & ~n28687 ;
  assign n30397 = n17209 ^ n9177 ^ 1'b0 ;
  assign n30398 = n4622 | n26405 ;
  assign n30401 = ~n1095 & n5662 ;
  assign n30402 = n30401 ^ n6557 ^ 1'b0 ;
  assign n30399 = n10684 | n26543 ;
  assign n30400 = n30399 ^ n19262 ^ n855 ;
  assign n30403 = n30402 ^ n30400 ^ 1'b0 ;
  assign n30404 = ~n17539 & n30403 ;
  assign n30405 = n4986 & ~n16221 ;
  assign n30406 = n3114 & n30405 ;
  assign n30407 = n30406 ^ n9094 ^ 1'b0 ;
  assign n30408 = ~n12494 & n30407 ;
  assign n30409 = n2655 ^ n182 ^ 1'b0 ;
  assign n30410 = n9349 ^ n7408 ^ 1'b0 ;
  assign n30411 = n13875 | n19063 ;
  assign n30412 = n2154 & ~n30411 ;
  assign n30413 = n3422 & n5353 ;
  assign n30414 = n16493 ^ n6142 ^ 1'b0 ;
  assign n30415 = n7937 & ~n30414 ;
  assign n30416 = n7737 & ~n23092 ;
  assign n30417 = n30416 ^ n12867 ^ 1'b0 ;
  assign n30418 = ~n27748 & n30417 ;
  assign n30419 = ( n2653 & ~n12047 ) | ( n2653 & n19168 ) | ( ~n12047 & n19168 ) ;
  assign n30420 = n2682 & ~n24578 ;
  assign n30421 = ~n2682 & n30420 ;
  assign n30422 = n312 & ~n22325 ;
  assign n30423 = n22325 & n30422 ;
  assign n30424 = n30423 ^ n21087 ^ 1'b0 ;
  assign n30425 = n30424 ^ n30314 ^ 1'b0 ;
  assign n30426 = ~n30421 & n30425 ;
  assign n30427 = n10348 & n15406 ;
  assign n30428 = ( n910 & n6690 ) | ( n910 & ~n18772 ) | ( n6690 & ~n18772 ) ;
  assign n30429 = n18742 ^ n1838 ^ n1551 ;
  assign n30430 = n30428 & ~n30429 ;
  assign n30431 = n7119 ^ n3062 ^ 1'b0 ;
  assign n30432 = n2117 & ~n30431 ;
  assign n30433 = n22540 | n30432 ;
  assign n30434 = ~n17749 & n30433 ;
  assign n30435 = ~n30430 & n30434 ;
  assign n30436 = ~n1337 & n19271 ;
  assign n30437 = n30436 ^ n5909 ^ 1'b0 ;
  assign n30438 = n30437 ^ n15347 ^ 1'b0 ;
  assign n30439 = n4259 | n6307 ;
  assign n30440 = n19605 | n30439 ;
  assign n30441 = n14117 & n30440 ;
  assign n30442 = ~n1235 & n1700 ;
  assign n30443 = n30442 ^ n9772 ^ 1'b0 ;
  assign n30444 = n16295 ^ n13044 ^ 1'b0 ;
  assign n30445 = n1191 | n4159 ;
  assign n30446 = n27370 ^ n4657 ^ 1'b0 ;
  assign n30447 = n9224 & n30446 ;
  assign n30448 = n26275 & ~n30447 ;
  assign n30449 = ~n14472 & n29108 ;
  assign n30450 = n28101 ^ n23727 ^ 1'b0 ;
  assign n30451 = ~n81 & n24308 ;
  assign n30452 = n28009 ^ n25824 ^ n4405 ;
  assign n30453 = ~n18603 & n30452 ;
  assign n30454 = n6006 | n12339 ;
  assign n30455 = n30454 ^ n347 ^ 1'b0 ;
  assign n30456 = n1276 & ~n16089 ;
  assign n30457 = ~n30455 & n30456 ;
  assign n30458 = n30457 ^ n17883 ^ 1'b0 ;
  assign n30459 = n968 & ~n30458 ;
  assign n30460 = ~n6036 & n30459 ;
  assign n30461 = n28139 & n30460 ;
  assign n30462 = n10751 | n30461 ;
  assign n30465 = n9592 ^ n8572 ^ 1'b0 ;
  assign n30463 = n1148 & ~n3842 ;
  assign n30464 = ~n4508 & n30463 ;
  assign n30466 = n30465 ^ n30464 ^ n11406 ;
  assign n30467 = n2226 ^ n983 ^ 1'b0 ;
  assign n30468 = n2693 & ~n30467 ;
  assign n30469 = n379 | n29466 ;
  assign n30470 = n5188 | n8849 ;
  assign n30471 = n30470 ^ n5655 ^ 1'b0 ;
  assign n30472 = n30471 ^ n700 ^ 1'b0 ;
  assign n30473 = n28011 ^ n6808 ^ 1'b0 ;
  assign n30474 = n6773 | n13837 ;
  assign n30475 = n10723 & n12215 ;
  assign n30476 = ~n16560 & n30475 ;
  assign n30477 = n30476 ^ n27307 ^ 1'b0 ;
  assign n30478 = ~n26636 & n30477 ;
  assign n30479 = n13355 | n16423 ;
  assign n30480 = n30479 ^ n29619 ^ 1'b0 ;
  assign n30481 = ~n1207 & n1707 ;
  assign n30482 = n683 & n30481 ;
  assign n30483 = n1079 & ~n30482 ;
  assign n30484 = n2586 ^ n212 ^ 1'b0 ;
  assign n30485 = n30483 & ~n30484 ;
  assign n30486 = n3392 & ~n30485 ;
  assign n30487 = n4722 | n17214 ;
  assign n30488 = n910 | n24792 ;
  assign n30489 = ( n2032 & n25443 ) | ( n2032 & n30215 ) | ( n25443 & n30215 ) ;
  assign n30490 = n3961 & n30489 ;
  assign n30492 = n24255 ^ n2802 ^ n28 ;
  assign n30493 = n21 | n30492 ;
  assign n30494 = n30493 ^ n26897 ^ 1'b0 ;
  assign n30491 = n10448 | n14934 ;
  assign n30495 = n30494 ^ n30491 ^ 1'b0 ;
  assign n30497 = n5305 & ~n6365 ;
  assign n30498 = n13946 ^ n788 ^ 1'b0 ;
  assign n30499 = n30497 | n30498 ;
  assign n30496 = n21767 ^ n1562 ^ 1'b0 ;
  assign n30500 = n30499 ^ n30496 ^ 1'b0 ;
  assign n30501 = n1182 & ~n30500 ;
  assign n30502 = n12366 ^ n7105 ^ n1025 ;
  assign n30504 = n14347 ^ n1736 ^ 1'b0 ;
  assign n30505 = n4276 | n30504 ;
  assign n30503 = n3239 & ~n21741 ;
  assign n30506 = n30505 ^ n30503 ^ 1'b0 ;
  assign n30507 = ~n1703 & n8049 ;
  assign n30508 = n10459 & n30507 ;
  assign n30509 = n2029 | n8915 ;
  assign n30510 = n30508 | n30509 ;
  assign n30511 = n162 & ~n17410 ;
  assign n30512 = n30510 & n30511 ;
  assign n30513 = n6860 & ~n12449 ;
  assign n30514 = n22517 & ~n30513 ;
  assign n30515 = n6133 ^ n2754 ^ n582 ;
  assign n30516 = n7337 | n9418 ;
  assign n30517 = n2236 | n30516 ;
  assign n30518 = n16360 ^ n9060 ^ 1'b0 ;
  assign n30519 = n23365 ^ n11346 ^ 1'b0 ;
  assign n30520 = ~n30518 & n30519 ;
  assign n30521 = n4374 ^ n3284 ^ 1'b0 ;
  assign n30522 = n18894 | n30521 ;
  assign n30523 = n30522 ^ n4195 ^ 1'b0 ;
  assign n30524 = n17822 & n29023 ;
  assign n30525 = ~n2109 & n10081 ;
  assign n30526 = n30525 ^ n17744 ^ 1'b0 ;
  assign n30527 = n12618 ^ n3983 ^ 1'b0 ;
  assign n30528 = n9769 & ~n30527 ;
  assign n30529 = n30528 ^ n20996 ^ 1'b0 ;
  assign n30530 = n24937 | n30529 ;
  assign n30531 = n30530 ^ n5829 ^ 1'b0 ;
  assign n30532 = n20988 & n30531 ;
  assign n30533 = ~n30526 & n30532 ;
  assign n30534 = n14194 ^ n14059 ^ 1'b0 ;
  assign n30535 = n6796 | n30534 ;
  assign n30536 = n30535 ^ n18635 ^ 1'b0 ;
  assign n30537 = n12807 & n30536 ;
  assign n30538 = n17788 & n30537 ;
  assign n30539 = n9735 ^ n560 ^ 1'b0 ;
  assign n30540 = n19237 | n30539 ;
  assign n30541 = n9354 & n17366 ;
  assign n30542 = n8258 ^ n2073 ^ 1'b0 ;
  assign n30543 = n2444 | n16209 ;
  assign n30544 = n24529 & ~n30543 ;
  assign n30545 = n19980 & n30544 ;
  assign n30546 = n16117 ^ n188 ^ 1'b0 ;
  assign n30547 = n6149 & ~n30546 ;
  assign n30548 = ~n16906 & n30547 ;
  assign n30549 = n29756 ^ n15289 ^ 1'b0 ;
  assign n30550 = n957 & ~n11027 ;
  assign n30551 = ~n17506 & n30550 ;
  assign n30552 = n30551 ^ n26988 ^ 1'b0 ;
  assign n30553 = n18631 | n20611 ;
  assign n30554 = n26200 ^ n21030 ^ 1'b0 ;
  assign n30555 = n12906 ^ n11595 ^ x5 ;
  assign n30556 = n10081 ^ n2349 ^ 1'b0 ;
  assign n30557 = ~n854 & n30556 ;
  assign n30558 = n30557 ^ n26877 ^ 1'b0 ;
  assign n30560 = n7825 | n8101 ;
  assign n30559 = n995 | n15478 ;
  assign n30561 = n30560 ^ n30559 ^ 1'b0 ;
  assign n30562 = ~n1360 & n2478 ;
  assign n30563 = n9134 & ~n11356 ;
  assign n30564 = n30562 & n30563 ;
  assign n30565 = n7314 & n26657 ;
  assign n30566 = n4575 | n7940 ;
  assign n30567 = n1734 & ~n4510 ;
  assign n30568 = n30567 ^ n9837 ^ 1'b0 ;
  assign n30569 = n2480 & n14362 ;
  assign n30570 = n18307 & n27884 ;
  assign n30571 = n24421 & n30570 ;
  assign n30572 = ~n698 & n1304 ;
  assign n30573 = n30572 ^ n18875 ^ 1'b0 ;
  assign n30574 = n27674 ^ n14808 ^ 1'b0 ;
  assign n30575 = ~n2843 & n30574 ;
  assign n30576 = n18556 & n28257 ;
  assign n30577 = n6630 ^ n5304 ^ 1'b0 ;
  assign n30578 = n15328 & n30577 ;
  assign n30579 = ~n30576 & n30578 ;
  assign n30580 = n2405 & n11621 ;
  assign n30581 = n27417 ^ n22442 ^ 1'b0 ;
  assign n30582 = n6980 & ~n30581 ;
  assign n30583 = n4046 & n16667 ;
  assign n30584 = n30583 ^ n3611 ^ 1'b0 ;
  assign n30585 = ~n3465 & n7327 ;
  assign n30586 = n19548 ^ n16335 ^ 1'b0 ;
  assign n30587 = n30586 ^ n1893 ^ 1'b0 ;
  assign n30588 = n24132 & n30587 ;
  assign n30589 = n5727 | n23396 ;
  assign n30590 = n30589 ^ n5587 ^ 1'b0 ;
  assign n30591 = n27242 | n30590 ;
  assign n30592 = n4293 ^ n3423 ^ 1'b0 ;
  assign n30593 = n2845 & ~n30592 ;
  assign n30594 = ~n19090 & n23486 ;
  assign n30595 = n1863 & n28070 ;
  assign n30596 = n30595 ^ n18963 ^ n5245 ;
  assign n30607 = n3006 & ~n7808 ;
  assign n30598 = n17980 ^ n7482 ^ 1'b0 ;
  assign n30599 = n2492 ^ n367 ^ 1'b0 ;
  assign n30600 = n28 & ~n2657 ;
  assign n30601 = ~n30599 & n30600 ;
  assign n30602 = n12474 & ~n30601 ;
  assign n30603 = n1422 & ~n30602 ;
  assign n30604 = n30603 ^ n5310 ^ n1453 ;
  assign n30605 = n30598 & ~n30604 ;
  assign n30606 = ~n16367 & n30605 ;
  assign n30608 = n30607 ^ n30606 ^ 1'b0 ;
  assign n30597 = n533 | n6439 ;
  assign n30609 = n30608 ^ n30597 ^ 1'b0 ;
  assign n30610 = n1438 | n4637 ;
  assign n30615 = ~n682 & n19150 ;
  assign n30616 = n682 & n30615 ;
  assign n30612 = ( n790 & ~n5638 ) | ( n790 & n7469 ) | ( ~n5638 & n7469 ) ;
  assign n30611 = n362 & ~n10244 ;
  assign n30613 = n30612 ^ n30611 ^ 1'b0 ;
  assign n30614 = n30613 ^ n21586 ^ 1'b0 ;
  assign n30617 = n30616 ^ n30614 ^ 1'b0 ;
  assign n30618 = n9121 & n30617 ;
  assign n30619 = n12988 ^ n204 ^ 1'b0 ;
  assign n30620 = n20822 | n30619 ;
  assign n30621 = ~n722 & n1699 ;
  assign n30622 = ~n14456 & n30621 ;
  assign n30623 = n2677 & ~n16478 ;
  assign n30624 = n9260 | n30623 ;
  assign n30625 = n28695 | n30624 ;
  assign n30626 = n23256 & ~n26768 ;
  assign n30627 = ~n6468 & n25651 ;
  assign n30628 = n21323 & n30627 ;
  assign n30629 = n4195 ^ n1148 ^ 1'b0 ;
  assign n30630 = n18389 ^ n7545 ^ 1'b0 ;
  assign n30631 = n7599 & ~n30630 ;
  assign n30632 = n30631 ^ n9187 ^ 1'b0 ;
  assign n30633 = n12228 & n30632 ;
  assign n30634 = n13823 & ~n30633 ;
  assign n30635 = n3052 & n4912 ;
  assign n30636 = n22524 ^ n17503 ^ 1'b0 ;
  assign n30637 = n4452 & n30636 ;
  assign n30638 = ~n4510 & n7556 ;
  assign n30639 = n14347 & n30638 ;
  assign n30640 = n30102 ^ n12751 ^ 1'b0 ;
  assign n30641 = n4741 | n30640 ;
  assign n30642 = ~n23454 & n30641 ;
  assign n30643 = n14736 | n23327 ;
  assign n30644 = n21535 & ~n30643 ;
  assign n30646 = n485 | n1469 ;
  assign n30647 = n18888 | n30646 ;
  assign n30648 = n30647 ^ n14768 ^ 1'b0 ;
  assign n30649 = n15404 ^ n6669 ^ 1'b0 ;
  assign n30650 = ~n30648 & n30649 ;
  assign n30645 = n7538 & ~n29050 ;
  assign n30651 = n30650 ^ n30645 ^ 1'b0 ;
  assign n30652 = n2053 & n3668 ;
  assign n30653 = n30652 ^ n16259 ^ 1'b0 ;
  assign n30654 = n30653 ^ n18307 ^ 1'b0 ;
  assign n30655 = ~n30651 & n30654 ;
  assign n30656 = n30655 ^ n27694 ^ 1'b0 ;
  assign n30662 = n30402 ^ n10819 ^ 1'b0 ;
  assign n30663 = ~n177 & n30662 ;
  assign n30657 = n21459 ^ n19267 ^ 1'b0 ;
  assign n30658 = ~n11329 & n30657 ;
  assign n30659 = n30658 ^ n20579 ^ 1'b0 ;
  assign n30660 = n1353 & n30659 ;
  assign n30661 = n30660 ^ n5775 ^ 1'b0 ;
  assign n30664 = n30663 ^ n30661 ^ 1'b0 ;
  assign n30665 = n23125 ^ n4070 ^ 1'b0 ;
  assign n30666 = n27349 ^ n26098 ^ 1'b0 ;
  assign n30667 = n11439 ^ n5391 ^ 1'b0 ;
  assign n30668 = n551 & n30667 ;
  assign n30669 = n3852 | n20759 ;
  assign n30670 = n13717 & ~n30669 ;
  assign n30671 = n873 & ~n30670 ;
  assign n30672 = n30671 ^ n6180 ^ 1'b0 ;
  assign n30673 = n16788 & ~n19555 ;
  assign n30674 = ~n30672 & n30673 ;
  assign n30675 = n24465 ^ n3052 ^ 1'b0 ;
  assign n30676 = n3636 | n30675 ;
  assign n30677 = n18726 | n30676 ;
  assign n30678 = n30677 ^ n6568 ^ 1'b0 ;
  assign n30679 = n19949 ^ n3280 ^ 1'b0 ;
  assign n30680 = ~n13601 & n30679 ;
  assign n30681 = n30680 ^ n11316 ^ 1'b0 ;
  assign n30682 = n12562 | n21003 ;
  assign n30683 = n2258 & ~n12407 ;
  assign n30685 = n788 & n1004 ;
  assign n30684 = n27802 & n28283 ;
  assign n30686 = n30685 ^ n30684 ^ 1'b0 ;
  assign n30687 = n27920 ^ n14053 ^ 1'b0 ;
  assign n30688 = ~n29403 & n30687 ;
  assign n30689 = n16491 | n29817 ;
  assign n30690 = n30688 | n30689 ;
  assign n30691 = n29311 ^ n14066 ^ 1'b0 ;
  assign n30692 = n16603 & ~n30691 ;
  assign n30693 = n631 & n16482 ;
  assign n30694 = ~n5900 & n30693 ;
  assign n30695 = n8313 ^ n2560 ^ 1'b0 ;
  assign n30696 = n30694 | n30695 ;
  assign n30697 = n19647 | n21225 ;
  assign n30698 = n15692 & ~n30697 ;
  assign n30699 = n18473 & n25195 ;
  assign n30700 = n22022 & n27970 ;
  assign n30701 = n30700 ^ n19697 ^ 1'b0 ;
  assign n30702 = n17482 ^ n6145 ^ 1'b0 ;
  assign n30703 = n2680 | n30702 ;
  assign n30704 = n630 & ~n30703 ;
  assign n30705 = n20425 & ~n24431 ;
  assign n30706 = n19051 ^ n1025 ^ 1'b0 ;
  assign n30707 = n7116 | n30706 ;
  assign n30708 = n30707 ^ n5057 ^ 1'b0 ;
  assign n30709 = n30708 ^ n12790 ^ 1'b0 ;
  assign n30710 = ~n11439 & n30709 ;
  assign n30711 = n343 | n805 ;
  assign n30712 = n17253 ^ n8944 ^ n8495 ;
  assign n30713 = n28681 ^ n3985 ^ 1'b0 ;
  assign n30714 = n28867 & ~n30713 ;
  assign n30715 = n18706 ^ n16085 ^ 1'b0 ;
  assign n30716 = n379 & ~n30715 ;
  assign n30717 = n1653 & ~n3827 ;
  assign n30718 = ( ~n5606 & n11233 ) | ( ~n5606 & n30717 ) | ( n11233 & n30717 ) ;
  assign n30721 = n856 | n1455 ;
  assign n30722 = n30721 ^ n397 ^ 1'b0 ;
  assign n30719 = n12744 & n19629 ;
  assign n30720 = n30719 ^ n10063 ^ 1'b0 ;
  assign n30723 = n30722 ^ n30720 ^ 1'b0 ;
  assign n30724 = ~n30718 & n30723 ;
  assign n30725 = ~n30716 & n30724 ;
  assign n30726 = n8582 & ~n30725 ;
  assign n30727 = n14246 & n20769 ;
  assign n30728 = n1947 & n2468 ;
  assign n30729 = n30728 ^ n12193 ^ 1'b0 ;
  assign n30730 = n13369 & n18909 ;
  assign n30731 = n3333 & n30730 ;
  assign n30732 = n24093 ^ n466 ^ 1'b0 ;
  assign n30733 = n9928 ^ n3500 ^ 1'b0 ;
  assign n30734 = n30733 ^ n13675 ^ 1'b0 ;
  assign n30735 = n30732 | n30734 ;
  assign n30736 = n12966 & n19416 ;
  assign n30737 = n30736 ^ n17537 ^ 1'b0 ;
  assign n30738 = n8211 & ~n30737 ;
  assign n30739 = n21466 ^ n19881 ^ 1'b0 ;
  assign n30740 = ( n4722 & n5828 ) | ( n4722 & ~n30739 ) | ( n5828 & ~n30739 ) ;
  assign n30741 = ~n852 & n4738 ;
  assign n30742 = n30741 ^ n7746 ^ 1'b0 ;
  assign n30743 = ~n30740 & n30742 ;
  assign n30744 = n24478 ^ n2463 ^ 1'b0 ;
  assign n30745 = n4757 & n30744 ;
  assign n30746 = ~n2431 & n30745 ;
  assign n30747 = n13608 & n30746 ;
  assign n30748 = n30747 ^ n2389 ^ 1'b0 ;
  assign n30749 = n25176 ^ n12801 ^ 1'b0 ;
  assign n30750 = ( n625 & n30748 ) | ( n625 & n30749 ) | ( n30748 & n30749 ) ;
  assign n30751 = ~n3113 & n6366 ;
  assign n30752 = n5970 & ~n15293 ;
  assign n30753 = n29666 & ~n30752 ;
  assign n30754 = n30753 ^ n790 ^ 1'b0 ;
  assign n30755 = n522 | n11169 ;
  assign n30756 = n757 ^ n382 ^ 1'b0 ;
  assign n30757 = n9057 & ~n30756 ;
  assign n30758 = n23033 & n30757 ;
  assign n30759 = n24078 & n30758 ;
  assign n30760 = n30759 ^ n11193 ^ 1'b0 ;
  assign n30761 = n6128 & ~n30760 ;
  assign n30762 = n2893 & ~n3915 ;
  assign n30763 = n30762 ^ n27227 ^ 1'b0 ;
  assign n30764 = n4439 & ~n30763 ;
  assign n30765 = ~n18199 & n30764 ;
  assign n30766 = n20340 ^ n3578 ^ 1'b0 ;
  assign n30767 = ( ~n2390 & n22099 ) | ( ~n2390 & n30766 ) | ( n22099 & n30766 ) ;
  assign n30768 = n10603 ^ n7707 ^ 1'b0 ;
  assign n30769 = n2754 & ~n6475 ;
  assign n30770 = n19593 ^ n18563 ^ 1'b0 ;
  assign n30771 = ( n30768 & n30769 ) | ( n30768 & ~n30770 ) | ( n30769 & ~n30770 ) ;
  assign n30772 = n22660 ^ n9100 ^ n1591 ;
  assign n30773 = n26943 & n30772 ;
  assign n30774 = n3584 & ~n20971 ;
  assign n30775 = n12424 & n30774 ;
  assign n30776 = n9108 & n11909 ;
  assign n30777 = n30775 | n30776 ;
  assign n30778 = n6836 | n30777 ;
  assign n30779 = n30778 ^ n11770 ^ 1'b0 ;
  assign n30781 = n18276 ^ n10540 ^ 1'b0 ;
  assign n30782 = n14032 & ~n30781 ;
  assign n30780 = n6423 | n7972 ;
  assign n30783 = n30782 ^ n30780 ^ 1'b0 ;
  assign n30784 = n655 | n1845 ;
  assign n30785 = n4175 & ~n24078 ;
  assign n30786 = n6949 & ~n17973 ;
  assign n30787 = n30786 ^ n11925 ^ n7420 ;
  assign n30788 = ( n314 & ~n9570 ) | ( n314 & n30787 ) | ( ~n9570 & n30787 ) ;
  assign n30789 = n12829 ^ n6954 ^ 1'b0 ;
  assign n30790 = ~n8341 & n30789 ;
  assign n30791 = n21778 & ~n26317 ;
  assign n30792 = ~n8266 & n22846 ;
  assign n30793 = n447 & n18939 ;
  assign n30794 = n4473 | n30793 ;
  assign n30795 = ~n2137 & n23658 ;
  assign n30797 = n9713 ^ n2668 ^ 1'b0 ;
  assign n30798 = n10782 & ~n30797 ;
  assign n30799 = n9364 | n30798 ;
  assign n30796 = n7379 & ~n12423 ;
  assign n30800 = n30799 ^ n30796 ^ 1'b0 ;
  assign n30801 = n15997 | n30800 ;
  assign n30802 = n30801 ^ n6153 ^ 1'b0 ;
  assign n30803 = n25878 ^ n11429 ^ 1'b0 ;
  assign n30804 = n1576 & n28181 ;
  assign n30805 = n30804 ^ n3537 ^ 1'b0 ;
  assign n30806 = n28081 | n30805 ;
  assign n30807 = n14337 & ~n30806 ;
  assign n30808 = n7588 ^ n5157 ^ 1'b0 ;
  assign n30809 = n6196 | n30808 ;
  assign n30810 = n10711 & ~n13717 ;
  assign n30811 = ~n4264 & n30810 ;
  assign n30812 = n30809 | n30811 ;
  assign n30813 = n30812 ^ n28368 ^ 1'b0 ;
  assign n30815 = n12533 ^ n1189 ^ 1'b0 ;
  assign n30816 = ~n9686 & n30815 ;
  assign n30814 = n8989 ^ n8216 ^ 1'b0 ;
  assign n30817 = n30816 ^ n30814 ^ 1'b0 ;
  assign n30818 = n25929 & ~n30817 ;
  assign n30819 = n9539 & n30818 ;
  assign n30820 = n1670 & n5682 ;
  assign n30821 = n30820 ^ n28960 ^ 1'b0 ;
  assign n30822 = n924 & ~n5475 ;
  assign n30823 = ~n5809 & n18127 ;
  assign n30824 = n30823 ^ n11524 ^ 1'b0 ;
  assign n30825 = n4432 & ~n30824 ;
  assign n30826 = n19468 & n29933 ;
  assign n30827 = n4044 & n8532 ;
  assign n30828 = n30827 ^ n2796 ^ 1'b0 ;
  assign n30829 = n23396 ^ n13971 ^ n11847 ;
  assign n30830 = ~n2914 & n7403 ;
  assign n30831 = n30830 ^ n2919 ^ 1'b0 ;
  assign n30832 = n28762 | n30831 ;
  assign n30833 = n2313 & n24976 ;
  assign n30834 = n30833 ^ n26119 ^ 1'b0 ;
  assign n30835 = n11846 ^ n11286 ^ 1'b0 ;
  assign n30836 = n18256 ^ n11466 ^ 1'b0 ;
  assign n30837 = ~n9358 & n13524 ;
  assign n30838 = n16906 ^ n8206 ^ 1'b0 ;
  assign n30839 = n5390 & ~n5823 ;
  assign n30843 = ~n3039 & n10147 ;
  assign n30844 = n22691 | n30843 ;
  assign n30840 = n11554 ^ n3727 ^ 1'b0 ;
  assign n30841 = n27230 & ~n30840 ;
  assign n30842 = n15332 | n30841 ;
  assign n30845 = n30844 ^ n30842 ^ 1'b0 ;
  assign n30846 = ~n10425 & n12337 ;
  assign n30847 = ~n7287 & n13436 ;
  assign n30848 = n30847 ^ n5184 ^ 1'b0 ;
  assign n30849 = n7256 & n30848 ;
  assign n30850 = n5744 & n30849 ;
  assign n30851 = ~n27519 & n30850 ;
  assign n30852 = n1688 & n25053 ;
  assign n30853 = ( n16193 & n17788 ) | ( n16193 & n30805 ) | ( n17788 & n30805 ) ;
  assign n30854 = n10545 & ~n16127 ;
  assign n30855 = n5160 | n7443 ;
  assign n30856 = n30854 & ~n30855 ;
  assign n30857 = n30856 ^ n26888 ^ 1'b0 ;
  assign n30858 = n2405 & n30857 ;
  assign n30859 = n6511 ^ n1853 ^ n1392 ;
  assign n30860 = n30859 ^ n2513 ^ 1'b0 ;
  assign n30861 = n5915 & ~n30860 ;
  assign n30862 = n21333 ^ n8915 ^ 1'b0 ;
  assign n30863 = ~n18977 & n30862 ;
  assign n30864 = n30863 ^ n488 ^ 1'b0 ;
  assign n30865 = n5435 & n6809 ;
  assign n30866 = n30865 ^ n2114 ^ 1'b0 ;
  assign n30867 = n4276 | n30866 ;
  assign n30868 = n30867 ^ n21890 ^ 1'b0 ;
  assign n30869 = n2041 & n30868 ;
  assign n30870 = ~n12897 & n30869 ;
  assign n30871 = n17370 | n22901 ;
  assign n30872 = n30871 ^ n1648 ^ 1'b0 ;
  assign n30873 = n15196 & ~n30872 ;
  assign n30874 = n30256 ^ n22497 ^ 1'b0 ;
  assign n30875 = n30873 & n30874 ;
  assign n30876 = n14274 ^ n4622 ^ 1'b0 ;
  assign n30877 = n14999 & n30876 ;
  assign n30878 = n10614 | n13041 ;
  assign n30879 = n5621 | n30878 ;
  assign n30880 = ~n13912 & n30879 ;
  assign n30881 = n16463 & n30880 ;
  assign n30882 = n10998 & n14798 ;
  assign n30883 = ( ~n6950 & n17899 ) | ( ~n6950 & n28648 ) | ( n17899 & n28648 ) ;
  assign n30884 = n30883 ^ n3731 ^ 1'b0 ;
  assign n30885 = n4835 & ~n30884 ;
  assign n30886 = n30885 ^ n1186 ^ 1'b0 ;
  assign n30887 = n4401 & ~n30886 ;
  assign n30888 = ~n10405 & n30887 ;
  assign n30889 = n22029 ^ n16721 ^ 1'b0 ;
  assign n30890 = n30889 ^ n26231 ^ 1'b0 ;
  assign n30891 = n12765 ^ n9699 ^ 1'b0 ;
  assign n30892 = n15885 ^ n5284 ^ n4809 ;
  assign n30893 = n30892 ^ n13403 ^ 1'b0 ;
  assign n30894 = n12950 ^ n9074 ^ n5866 ;
  assign n30895 = ~n4667 & n30894 ;
  assign n30896 = n4365 & ~n9709 ;
  assign n30897 = ~n5587 & n30896 ;
  assign n30898 = n1969 & n26126 ;
  assign n30899 = n21767 & n30898 ;
  assign n30900 = n30899 ^ n15684 ^ 1'b0 ;
  assign n30901 = n27368 ^ n19274 ^ 1'b0 ;
  assign n30902 = n21090 ^ n11269 ^ 1'b0 ;
  assign n30903 = n3467 ^ n3050 ^ 1'b0 ;
  assign n30904 = n197 & ~n1969 ;
  assign n30905 = n6359 & n26287 ;
  assign n30906 = n219 & n30905 ;
  assign n30907 = n30904 & ~n30906 ;
  assign n30908 = ~n13578 & n30907 ;
  assign n30909 = n14080 & ~n25384 ;
  assign n30910 = ~n19993 & n30909 ;
  assign n30911 = n19210 & n30447 ;
  assign n30912 = n30911 ^ n6216 ^ 1'b0 ;
  assign n30913 = ~n1647 & n24797 ;
  assign n30914 = ~n30912 & n30913 ;
  assign n30915 = n23872 & ~n30914 ;
  assign n30916 = ( n12153 & n12169 ) | ( n12153 & ~n28463 ) | ( n12169 & ~n28463 ) ;
  assign n30917 = ( ~n5511 & n11784 ) | ( ~n5511 & n30916 ) | ( n11784 & n30916 ) ;
  assign n30918 = n754 | n16323 ;
  assign n30919 = n7086 & ~n30918 ;
  assign n30920 = n30919 ^ n21184 ^ 1'b0 ;
  assign n30921 = n14766 ^ n8688 ^ 1'b0 ;
  assign n30922 = n1385 | n30921 ;
  assign n30923 = n6934 & ~n30922 ;
  assign n30924 = n30923 ^ n3221 ^ 1'b0 ;
  assign n30925 = n9553 ^ n4804 ^ 1'b0 ;
  assign n30926 = n30924 & ~n30925 ;
  assign n30927 = ~n347 & n15614 ;
  assign n30928 = n24180 & n30927 ;
  assign n30929 = n13977 ^ n12327 ^ 1'b0 ;
  assign n30930 = ~n2510 & n30929 ;
  assign n30931 = n30930 ^ n3544 ^ 1'b0 ;
  assign n30932 = n1142 & ~n9202 ;
  assign n30933 = n30932 ^ n894 ^ 1'b0 ;
  assign n30934 = n30933 ^ n14066 ^ n8183 ;
  assign n30936 = n3119 & ~n7108 ;
  assign n30937 = n30936 ^ x0 ^ 1'b0 ;
  assign n30935 = n2798 ^ n1080 ^ n511 ;
  assign n30938 = n30937 ^ n30935 ^ 1'b0 ;
  assign n30939 = n9833 | n30938 ;
  assign n30940 = n30939 ^ n192 ^ 1'b0 ;
  assign n30941 = n1277 & n3671 ;
  assign n30942 = ~n20093 & n30941 ;
  assign n30943 = n30942 ^ n8283 ^ 1'b0 ;
  assign n30944 = ~n8896 & n13772 ;
  assign n30945 = n17593 ^ n7271 ^ 1'b0 ;
  assign n30946 = n1068 | n1582 ;
  assign n30947 = n1851 & n30946 ;
  assign n30948 = n28670 ^ n347 ^ 1'b0 ;
  assign n30949 = n11500 ^ n6660 ^ 1'b0 ;
  assign n30950 = n16387 & ~n24637 ;
  assign n30951 = ~n30949 & n30950 ;
  assign n30952 = n24645 | n30951 ;
  assign n30953 = n30952 ^ n1770 ^ 1'b0 ;
  assign n30954 = ~n7595 & n20158 ;
  assign n30955 = ~n12788 & n30954 ;
  assign n30956 = n30953 & ~n30955 ;
  assign n30957 = n3295 & n30956 ;
  assign n30958 = n10430 | n20577 ;
  assign n30959 = n3869 & ~n18873 ;
  assign n30960 = n30959 ^ n3366 ^ 1'b0 ;
  assign n30961 = n10158 & n30960 ;
  assign n30962 = n14675 ^ n4956 ^ 1'b0 ;
  assign n30963 = ( n248 & n1582 ) | ( n248 & ~n3550 ) | ( n1582 & ~n3550 ) ;
  assign n30964 = ( n528 & ~n30745 ) | ( n528 & n30963 ) | ( ~n30745 & n30963 ) ;
  assign n30965 = n30550 ^ n23806 ^ 1'b0 ;
  assign n30966 = n9952 ^ n7437 ^ 1'b0 ;
  assign n30967 = n22654 | n22862 ;
  assign n30968 = n16918 ^ n13500 ^ 1'b0 ;
  assign n30969 = n28068 & n30968 ;
  assign n30970 = n5054 & ~n13288 ;
  assign n30971 = n15923 & n24616 ;
  assign n30972 = n16286 ^ n5909 ^ n1592 ;
  assign n30973 = n23398 ^ n2216 ^ 1'b0 ;
  assign n30974 = n22349 & n30973 ;
  assign n30975 = n8308 & ~n13342 ;
  assign n30976 = n10415 | n30975 ;
  assign n30977 = n4571 & n8817 ;
  assign n30978 = n30977 ^ n983 ^ 1'b0 ;
  assign n30979 = n15257 & n30978 ;
  assign n30980 = n15078 & n28119 ;
  assign n30984 = n1327 | n2769 ;
  assign n30985 = n2327 & ~n30984 ;
  assign n30981 = n30354 ^ n8850 ^ 1'b0 ;
  assign n30982 = n12938 & ~n30981 ;
  assign n30983 = n14249 & n30982 ;
  assign n30986 = n30985 ^ n30983 ^ 1'b0 ;
  assign n30987 = n7655 & n9731 ;
  assign n30988 = n3143 | n27093 ;
  assign n30989 = n23433 ^ n15618 ^ n7188 ;
  assign n30990 = n5269 | n15265 ;
  assign n30991 = n30990 ^ n30737 ^ 1'b0 ;
  assign n30992 = n1743 & n30991 ;
  assign n30997 = ~n3574 & n11694 ;
  assign n30998 = n30997 ^ n20785 ^ n2141 ;
  assign n30999 = n30998 ^ n7397 ^ 1'b0 ;
  assign n30993 = n7399 ^ n472 ^ 1'b0 ;
  assign n30994 = n30993 ^ n1551 ^ 1'b0 ;
  assign n30995 = n16758 & n30994 ;
  assign n30996 = n30995 ^ n9957 ^ 1'b0 ;
  assign n31000 = n30999 ^ n30996 ^ 1'b0 ;
  assign n31001 = n30992 & ~n31000 ;
  assign n31002 = n7280 ^ n2550 ^ 1'b0 ;
  assign n31003 = n11146 & ~n27276 ;
  assign n31004 = ~n25014 & n31003 ;
  assign n31005 = n31002 & n31004 ;
  assign n31006 = n4891 & ~n12076 ;
  assign n31007 = ~n5865 & n18963 ;
  assign n31008 = n31006 & n31007 ;
  assign n31009 = n31008 ^ n1908 ^ 1'b0 ;
  assign n31010 = n12202 ^ n11088 ^ 1'b0 ;
  assign n31011 = n23185 & ~n31010 ;
  assign n31012 = n1878 | n17172 ;
  assign n31013 = n31012 ^ n26364 ^ 1'b0 ;
  assign n31014 = n2382 | n31013 ;
  assign n31015 = n27984 ^ n3367 ^ n564 ;
  assign n31016 = n31015 ^ n18986 ^ n6749 ;
  assign n31017 = n522 & ~n26455 ;
  assign n31018 = ~n21178 & n31017 ;
  assign n31019 = n25096 ^ n7816 ^ n5150 ;
  assign n31020 = n18981 ^ n8118 ^ 1'b0 ;
  assign n31021 = n17329 ^ n7523 ^ n5364 ;
  assign n31022 = n7867 & n9276 ;
  assign n31023 = n31022 ^ n10945 ^ 1'b0 ;
  assign n31024 = n31023 ^ n28902 ^ 1'b0 ;
  assign n31025 = n31021 & n31024 ;
  assign n31026 = n4732 ^ n1775 ^ 1'b0 ;
  assign n31027 = n31026 ^ n3521 ^ 1'b0 ;
  assign n31028 = n12228 & n31027 ;
  assign n31029 = n11515 & ~n31028 ;
  assign n31030 = n10245 & n25446 ;
  assign n31031 = n10998 & ~n26660 ;
  assign n31032 = n27045 & n31031 ;
  assign n31033 = ~n31030 & n31032 ;
  assign n31034 = n23222 ^ n22133 ^ 1'b0 ;
  assign n31035 = n5497 ^ n3979 ^ 1'b0 ;
  assign n31036 = n28520 & n30769 ;
  assign n31037 = n31036 ^ n14926 ^ 1'b0 ;
  assign n31038 = ( ~n2474 & n13957 ) | ( ~n2474 & n31037 ) | ( n13957 & n31037 ) ;
  assign n31040 = n13735 & n25185 ;
  assign n31039 = n11119 ^ n5122 ^ n1966 ;
  assign n31041 = n31040 ^ n31039 ^ 1'b0 ;
  assign n31042 = n4845 & ~n18310 ;
  assign n31043 = n21514 & n31042 ;
  assign n31044 = n1534 & ~n8246 ;
  assign n31045 = n31044 ^ n10778 ^ 1'b0 ;
  assign n31046 = n25813 | n31045 ;
  assign n31047 = n1546 & ~n12808 ;
  assign n31048 = n31047 ^ n19219 ^ 1'b0 ;
  assign n31049 = n2492 | n6241 ;
  assign n31050 = ( n13677 & ~n16512 ) | ( n13677 & n31049 ) | ( ~n16512 & n31049 ) ;
  assign n31051 = n20838 ^ n12496 ^ 1'b0 ;
  assign n31052 = n31051 ^ n19064 ^ n5209 ;
  assign n31053 = n27545 | n31052 ;
  assign n31054 = n13346 ^ n7403 ^ 1'b0 ;
  assign n31055 = n16538 & n31054 ;
  assign n31056 = ~n8310 & n19973 ;
  assign n31057 = ~n20030 & n31056 ;
  assign n31058 = ~n7206 & n8111 ;
  assign n31059 = n31058 ^ n4142 ^ 1'b0 ;
  assign n31060 = n18696 & ~n31059 ;
  assign n31061 = n31057 & n31060 ;
  assign n31062 = n21843 | n31061 ;
  assign n31063 = n2108 & ~n30830 ;
  assign n31064 = n15374 ^ n9608 ^ 1'b0 ;
  assign n31065 = n8438 ^ n1338 ^ 1'b0 ;
  assign n31066 = ~n18156 & n31065 ;
  assign n31067 = n9775 & ~n26697 ;
  assign n31068 = ~n5544 & n31067 ;
  assign n31069 = n4171 | n20136 ;
  assign n31070 = n31069 ^ n9287 ^ 1'b0 ;
  assign n31071 = n13876 ^ n4364 ^ 1'b0 ;
  assign n31072 = n233 & n31071 ;
  assign n31073 = ~n31070 & n31072 ;
  assign n31074 = n28387 & n31073 ;
  assign n31075 = n24137 & ~n24317 ;
  assign n31076 = n31075 ^ n26229 ^ 1'b0 ;
  assign n31077 = n1743 | n17417 ;
  assign n31078 = n15324 | n31077 ;
  assign n31079 = n7327 | n8588 ;
  assign n31080 = n25685 & ~n31079 ;
  assign n31081 = n31080 ^ n1134 ^ 1'b0 ;
  assign n31082 = n25731 | n31081 ;
  assign n31083 = n15374 | n30320 ;
  assign n31084 = n31083 ^ n2978 ^ 1'b0 ;
  assign n31085 = n26045 ^ n20498 ^ 1'b0 ;
  assign n31086 = n13469 & n31085 ;
  assign n31087 = n31086 ^ n5076 ^ 1'b0 ;
  assign n31088 = n9050 & ~n10277 ;
  assign n31089 = n7672 & ~n15420 ;
  assign n31090 = n29847 & n31089 ;
  assign n31092 = n4479 & ~n5353 ;
  assign n31093 = n3094 & n31092 ;
  assign n31091 = n6342 ^ n4394 ^ n2864 ;
  assign n31094 = n31093 ^ n31091 ^ 1'b0 ;
  assign n31095 = n9562 | n15287 ;
  assign n31096 = n9562 & ~n31095 ;
  assign n31097 = n6527 | n21170 ;
  assign n31098 = n31096 & ~n31097 ;
  assign n31099 = n17121 | n31098 ;
  assign n31100 = n17121 & ~n31099 ;
  assign n31101 = n26644 ^ n19984 ^ n6931 ;
  assign n31102 = n21954 ^ n15030 ^ 1'b0 ;
  assign n31103 = n7134 & ~n31102 ;
  assign n31104 = n31103 ^ n249 ^ 1'b0 ;
  assign n31105 = n26667 ^ n15114 ^ n7820 ;
  assign n31106 = ~n26054 & n31105 ;
  assign n31107 = n2155 ^ n387 ^ 1'b0 ;
  assign n31108 = n7523 & ~n16406 ;
  assign n31109 = n31108 ^ n23908 ^ n6063 ;
  assign n31110 = n25081 ^ n3050 ^ 1'b0 ;
  assign n31111 = n2953 ^ n93 ^ 1'b0 ;
  assign n31112 = n9305 & ~n31111 ;
  assign n31113 = n31112 ^ n623 ^ 1'b0 ;
  assign n31114 = ~n16543 & n19322 ;
  assign n31115 = n31114 ^ n9319 ^ 1'b0 ;
  assign n31116 = ~n9974 & n26949 ;
  assign n31117 = ~n5570 & n31116 ;
  assign n31118 = ~n183 & n3118 ;
  assign n31119 = n9253 ^ n4526 ^ 1'b0 ;
  assign n31120 = n16002 & n25579 ;
  assign n31121 = n25977 | n31120 ;
  assign n31122 = n30703 & ~n31121 ;
  assign n31123 = n14349 ^ n9419 ^ 1'b0 ;
  assign n31124 = n28490 & n31123 ;
  assign n31125 = n31124 ^ n3173 ^ 1'b0 ;
  assign n31126 = n31125 ^ n8870 ^ 1'b0 ;
  assign n31127 = ~n17280 & n31126 ;
  assign n31128 = n27188 ^ n13753 ^ 1'b0 ;
  assign n31129 = n11942 ^ n3248 ^ 1'b0 ;
  assign n31130 = n31128 & n31129 ;
  assign n31131 = n8815 ^ n7577 ^ n3705 ;
  assign n31132 = ~n4873 & n31131 ;
  assign n31133 = n24331 ^ n22590 ^ 1'b0 ;
  assign n31135 = ~n2900 & n3229 ;
  assign n31134 = n16004 & ~n27856 ;
  assign n31136 = n31135 ^ n31134 ^ 1'b0 ;
  assign n31137 = n7342 ^ n2783 ^ n810 ;
  assign n31138 = n15600 & ~n31137 ;
  assign n31139 = n31138 ^ n13462 ^ 1'b0 ;
  assign n31140 = n13879 | n31139 ;
  assign n31141 = n2445 | n31140 ;
  assign n31142 = n6488 & n14001 ;
  assign n31143 = n372 & n31142 ;
  assign n31144 = n13785 ^ n8879 ^ n551 ;
  assign n31145 = n31144 ^ n2356 ^ 1'b0 ;
  assign n31146 = n14884 ^ n3083 ^ 1'b0 ;
  assign n31147 = n13083 | n31146 ;
  assign n31152 = n273 & ~n1201 ;
  assign n31153 = n1201 & n31152 ;
  assign n31148 = ~n362 & n1570 ;
  assign n31149 = n362 & n31148 ;
  assign n31150 = ~n4116 & n31149 ;
  assign n31151 = n14652 & n31150 ;
  assign n31154 = n31153 ^ n31151 ^ 1'b0 ;
  assign n31155 = ~n5097 & n31154 ;
  assign n31156 = n5097 & n31155 ;
  assign n31157 = ~n1205 & n2607 ;
  assign n31158 = ~n2607 & n31157 ;
  assign n31159 = n31158 ^ n11257 ^ 1'b0 ;
  assign n31160 = ~n948 & n31159 ;
  assign n31161 = n31160 ^ n23030 ^ 1'b0 ;
  assign n31162 = ~n31156 & n31161 ;
  assign n31167 = ~n11196 & n11489 ;
  assign n31163 = n13682 ^ n2498 ^ 1'b0 ;
  assign n31164 = ~n16295 & n31163 ;
  assign n31165 = ~n7562 & n31164 ;
  assign n31166 = n7526 & n31165 ;
  assign n31168 = n31167 ^ n31166 ^ 1'b0 ;
  assign n31170 = n27235 ^ n6554 ^ 1'b0 ;
  assign n31171 = n5195 & ~n31170 ;
  assign n31169 = n7308 & n27363 ;
  assign n31172 = n31171 ^ n31169 ^ 1'b0 ;
  assign n31173 = n16101 | n31172 ;
  assign n31174 = n4082 & ~n15557 ;
  assign n31175 = ~n22073 & n31174 ;
  assign n31176 = n334 & ~n18958 ;
  assign n31177 = n31176 ^ n2361 ^ 1'b0 ;
  assign n31178 = n23716 & ~n31177 ;
  assign n31179 = n6318 & ~n11383 ;
  assign n31180 = n16596 & n31179 ;
  assign n31181 = n5736 ^ n2549 ^ 1'b0 ;
  assign n31182 = ~n24692 & n31181 ;
  assign n31183 = ( ~n1688 & n10227 ) | ( ~n1688 & n26511 ) | ( n10227 & n26511 ) ;
  assign n31184 = n31183 ^ n7534 ^ 1'b0 ;
  assign n31185 = ( n31180 & ~n31182 ) | ( n31180 & n31184 ) | ( ~n31182 & n31184 ) ;
  assign n31186 = ~n9624 & n12470 ;
  assign n31187 = n25402 ^ n6878 ^ 1'b0 ;
  assign n31188 = n31187 ^ n7509 ^ n5039 ;
  assign n31189 = n31186 & ~n31188 ;
  assign n31191 = n16298 ^ n3323 ^ 1'b0 ;
  assign n31192 = n1941 & ~n31191 ;
  assign n31193 = n14948 & ~n31192 ;
  assign n31190 = n5524 & ~n15184 ;
  assign n31194 = n31193 ^ n31190 ^ 1'b0 ;
  assign n31195 = n582 | n12647 ;
  assign n31199 = n8433 | n14136 ;
  assign n31198 = n25732 ^ n22829 ^ n2415 ;
  assign n31196 = n9596 ^ n2446 ^ 1'b0 ;
  assign n31197 = n22474 & n31196 ;
  assign n31200 = n31199 ^ n31198 ^ n31197 ;
  assign n31201 = n4160 | n30759 ;
  assign n31202 = n23811 | n31201 ;
  assign n31203 = n11876 ^ n7360 ^ 1'b0 ;
  assign n31204 = n13582 | n31203 ;
  assign n31205 = n3736 | n19805 ;
  assign n31206 = n31205 ^ n20168 ^ 1'b0 ;
  assign n31207 = n31206 ^ n8783 ^ n682 ;
  assign n31208 = n820 & n8779 ;
  assign n31209 = n5564 & n31208 ;
  assign n31210 = ~n31207 & n31209 ;
  assign n31211 = n5685 & ~n31210 ;
  assign n31212 = n25604 ^ n21046 ^ 1'b0 ;
  assign n31213 = n5010 & ~n21030 ;
  assign n31214 = n31213 ^ n13240 ^ 1'b0 ;
  assign n31215 = n31214 ^ n27668 ^ 1'b0 ;
  assign n31216 = n5151 & ~n10468 ;
  assign n31217 = ~n17927 & n31216 ;
  assign n31218 = n18899 ^ n15246 ^ 1'b0 ;
  assign n31219 = n31217 | n31218 ;
  assign n31220 = n2906 ^ n839 ^ 1'b0 ;
  assign n31221 = n2197 | n31220 ;
  assign n31222 = n418 & n26556 ;
  assign n31223 = n30315 ^ n16751 ^ n13449 ;
  assign n31224 = n2101 & ~n10050 ;
  assign n31225 = n16703 ^ n12453 ^ 1'b0 ;
  assign n31226 = n23550 | n31225 ;
  assign n31227 = n31226 ^ n18006 ^ 1'b0 ;
  assign n31228 = ~n26630 & n31227 ;
  assign n31229 = ~n13451 & n31228 ;
  assign n31230 = n16112 ^ n14780 ^ n4260 ;
  assign n31231 = n10481 & ~n31230 ;
  assign n31232 = n4357 & n31231 ;
  assign n31233 = n3000 & n12103 ;
  assign n31234 = ~n3500 & n31233 ;
  assign n31235 = n2548 | n31234 ;
  assign n31236 = n5468 & ~n31235 ;
  assign n31237 = x11 & n9036 ;
  assign n31238 = ~n9036 & n31237 ;
  assign n31239 = n701 & n3400 ;
  assign n31240 = ~n1697 & n31239 ;
  assign n31241 = n28357 ^ n11978 ^ 1'b0 ;
  assign n31242 = ~n17474 & n31241 ;
  assign n31243 = ~n31240 & n31242 ;
  assign n31244 = ~n19045 & n31243 ;
  assign n31245 = n31244 ^ n30247 ^ 1'b0 ;
  assign n31246 = n31238 | n31245 ;
  assign n31247 = n2549 | n6760 ;
  assign n31248 = n31247 ^ n6210 ^ 1'b0 ;
  assign n31249 = n4746 & ~n31248 ;
  assign n31250 = n30089 ^ n6876 ^ 1'b0 ;
  assign n31251 = n10656 & ~n31250 ;
  assign n31252 = n5562 & n31251 ;
  assign n31253 = n11331 & n11759 ;
  assign n31254 = n18907 ^ n9474 ^ 1'b0 ;
  assign n31255 = n1141 & ~n31254 ;
  assign n31256 = n1697 | n31255 ;
  assign n31257 = n5680 ^ n1099 ^ 1'b0 ;
  assign n31258 = n3240 & n19903 ;
  assign n31259 = n31257 & n31258 ;
  assign n31260 = n3027 & ~n6373 ;
  assign n31261 = n2784 & n6998 ;
  assign n31262 = n28056 & n31261 ;
  assign n31263 = n13475 & ~n30259 ;
  assign n31264 = n31262 & n31263 ;
  assign n31265 = n24805 | n31264 ;
  assign n31266 = n31265 ^ n7588 ^ 1'b0 ;
  assign n31267 = n21253 & ~n30803 ;
  assign n31268 = n9725 & n31267 ;
  assign n31269 = n21651 ^ n17934 ^ 1'b0 ;
  assign n31270 = n30752 & n31269 ;
  assign n31271 = ~n11251 & n30823 ;
  assign n31272 = n11383 ^ n2728 ^ 1'b0 ;
  assign n31273 = n9077 ^ n8387 ^ 1'b0 ;
  assign n31274 = n9884 & ~n31273 ;
  assign n31275 = n5558 & ~n12740 ;
  assign n31276 = n12317 ^ n1471 ^ 1'b0 ;
  assign n31277 = ~n2411 & n31276 ;
  assign n31278 = n31275 & n31277 ;
  assign n31279 = n15970 ^ n15470 ^ 1'b0 ;
  assign n31280 = n18219 ^ n1352 ^ 1'b0 ;
  assign n31281 = n29968 & n31280 ;
  assign n31287 = ( n6292 & ~n7681 ) | ( n6292 & n20067 ) | ( ~n7681 & n20067 ) ;
  assign n31288 = n3934 | n31287 ;
  assign n31289 = n31288 ^ n18898 ^ 1'b0 ;
  assign n31282 = n16998 ^ n1450 ^ 1'b0 ;
  assign n31283 = n20419 & ~n31282 ;
  assign n31284 = n31283 ^ n4977 ^ 1'b0 ;
  assign n31285 = n1050 & n31284 ;
  assign n31286 = n18169 & n31285 ;
  assign n31290 = n31289 ^ n31286 ^ 1'b0 ;
  assign n31291 = n23303 ^ n17511 ^ 1'b0 ;
  assign n31292 = n11409 & ~n31291 ;
  assign n31293 = ~n1181 & n21823 ;
  assign n31294 = n1413 | n31164 ;
  assign n31295 = ~n22477 & n24603 ;
  assign n31296 = n18228 & n25160 ;
  assign n31297 = ~n31295 & n31296 ;
  assign n31298 = n8525 & ~n13144 ;
  assign n31299 = n2270 & n31298 ;
  assign n31300 = n31297 & n31299 ;
  assign n31301 = n2132 | n8594 ;
  assign n31302 = n31301 ^ n7147 ^ 1'b0 ;
  assign n31303 = n1609 | n15902 ;
  assign n31304 = n886 | n31303 ;
  assign n31305 = ~n11524 & n13033 ;
  assign n31306 = n25370 & n31305 ;
  assign n31307 = n1315 | n12385 ;
  assign n31308 = n31307 ^ n3420 ^ 1'b0 ;
  assign n31309 = n15423 ^ n6764 ^ 1'b0 ;
  assign n31310 = n31309 ^ n3759 ^ 1'b0 ;
  assign n31311 = n1370 & n15995 ;
  assign n31312 = n11979 ^ n1918 ^ 1'b0 ;
  assign n31313 = n1216 & n31312 ;
  assign n31314 = ( n12899 & n31311 ) | ( n12899 & n31313 ) | ( n31311 & n31313 ) ;
  assign n31315 = n13108 ^ n7990 ^ 1'b0 ;
  assign n31317 = n15467 & n26135 ;
  assign n31318 = n31317 ^ n7589 ^ 1'b0 ;
  assign n31316 = ~n11446 & n16846 ;
  assign n31319 = n31318 ^ n31316 ^ 1'b0 ;
  assign n31320 = n10647 ^ n7493 ^ 1'b0 ;
  assign n31321 = n10593 & n31320 ;
  assign n31322 = ~n11500 & n31321 ;
  assign n31323 = n11462 & ~n31322 ;
  assign n31324 = n31323 ^ n3840 ^ 1'b0 ;
  assign n31325 = ~n28537 & n31324 ;
  assign n31326 = n24715 & n31325 ;
  assign n31327 = n29865 ^ n25189 ^ 1'b0 ;
  assign n31328 = n7463 | n31327 ;
  assign n31329 = n29324 ^ n15906 ^ n9831 ;
  assign n31330 = n21 & ~n31329 ;
  assign n31331 = n2066 & n7499 ;
  assign n31332 = n31330 & n31331 ;
  assign n31333 = n6893 ^ n3268 ^ 1'b0 ;
  assign n31334 = ~n13594 & n31333 ;
  assign n31335 = ~n1525 & n31334 ;
  assign n31336 = n31335 ^ n18934 ^ 1'b0 ;
  assign n31337 = n875 & ~n14670 ;
  assign n31338 = ~n4008 & n23856 ;
  assign n31339 = n1505 & n23214 ;
  assign n31340 = ~n24324 & n31339 ;
  assign n31341 = n31340 ^ n14111 ^ 1'b0 ;
  assign n31342 = n31338 | n31341 ;
  assign n31343 = n3268 & ~n31342 ;
  assign n31344 = n26015 & n31343 ;
  assign n31345 = ( ~n2005 & n6610 ) | ( ~n2005 & n11295 ) | ( n6610 & n11295 ) ;
  assign n31346 = n31345 ^ n11573 ^ 1'b0 ;
  assign n31347 = n24514 & n31346 ;
  assign n31348 = n21818 ^ n2594 ^ 1'b0 ;
  assign n31349 = n772 | n31348 ;
  assign n31350 = n29046 ^ n28857 ^ 1'b0 ;
  assign n31351 = n8688 | n10363 ;
  assign n31352 = n31351 ^ n3011 ^ 1'b0 ;
  assign n31353 = n6811 | n31352 ;
  assign n31354 = n5027 | n10883 ;
  assign n31355 = ~n456 & n7259 ;
  assign n31356 = n9598 ^ n5684 ^ 1'b0 ;
  assign n31357 = n5660 | n31356 ;
  assign n31358 = n31355 & ~n31357 ;
  assign n31359 = n31354 & ~n31358 ;
  assign n31360 = n10426 ^ n8054 ^ 1'b0 ;
  assign n31361 = n10003 | n31360 ;
  assign n31362 = ~n21021 & n27199 ;
  assign n31363 = n31362 ^ n18111 ^ 1'b0 ;
  assign n31364 = n10031 | n31363 ;
  assign n31365 = n6043 | n26066 ;
  assign n31366 = n31365 ^ n3214 ^ 1'b0 ;
  assign n31367 = n6393 | n12616 ;
  assign n31368 = n31367 ^ n10670 ^ 1'b0 ;
  assign n31369 = n4747 & n16682 ;
  assign n31370 = n12511 & n31369 ;
  assign n31371 = n31370 ^ n16941 ^ n7732 ;
  assign n31372 = n25584 ^ n22956 ^ 1'b0 ;
  assign n31373 = n26763 & ~n31244 ;
  assign n31374 = n16961 & n31373 ;
  assign n31375 = n25207 ^ n3818 ^ 1'b0 ;
  assign n31376 = n6524 & n16920 ;
  assign n31377 = ~n25154 & n31376 ;
  assign n31378 = n12585 & ~n31377 ;
  assign n31379 = ~n30380 & n31378 ;
  assign n31380 = ~n2049 & n26592 ;
  assign n31381 = n30593 & n31380 ;
  assign n31382 = n31381 ^ n21293 ^ 1'b0 ;
  assign n31383 = n898 & ~n10391 ;
  assign n31384 = n31383 ^ n8542 ^ 1'b0 ;
  assign n31385 = n1655 & ~n22321 ;
  assign n31386 = n12206 & ~n26711 ;
  assign n31387 = n11446 | n21293 ;
  assign n31388 = n23673 & ~n31387 ;
  assign n31389 = n7105 & ~n13042 ;
  assign n31390 = n798 & ~n31389 ;
  assign n31391 = n13397 ^ n5492 ^ 1'b0 ;
  assign n31392 = n8607 | n31391 ;
  assign n31393 = n31392 ^ n7562 ^ 1'b0 ;
  assign n31394 = n26821 ^ n3736 ^ 1'b0 ;
  assign n31395 = n7921 | n31394 ;
  assign n31396 = n631 & n2236 ;
  assign n31397 = n31396 ^ n11576 ^ 1'b0 ;
  assign n31398 = n31397 ^ n12393 ^ 1'b0 ;
  assign n31399 = n16361 & ~n21478 ;
  assign n31400 = n6771 & ~n31399 ;
  assign n31401 = n7965 ^ n6316 ^ n194 ;
  assign n31402 = n31401 ^ n13345 ^ 1'b0 ;
  assign n31403 = n31026 ^ n21217 ^ 1'b0 ;
  assign n31404 = n2303 & ~n31403 ;
  assign n31405 = n31404 ^ n14311 ^ 1'b0 ;
  assign n31406 = ~n3064 & n16084 ;
  assign n31407 = n15542 ^ n9258 ^ 1'b0 ;
  assign n31408 = n3756 & n31407 ;
  assign n31409 = ~n3742 & n12817 ;
  assign n31410 = n31409 ^ n3081 ^ 1'b0 ;
  assign n31411 = ~n3299 & n31410 ;
  assign n31412 = n31411 ^ n9057 ^ 1'b0 ;
  assign n31413 = ~n2175 & n17678 ;
  assign n31414 = n31412 & n31413 ;
  assign n31415 = ( n31406 & n31408 ) | ( n31406 & ~n31414 ) | ( n31408 & ~n31414 ) ;
  assign n31416 = n31415 ^ n14949 ^ 1'b0 ;
  assign n31417 = n8844 | n10963 ;
  assign n31418 = ( n5525 & ~n6556 ) | ( n5525 & n7083 ) | ( ~n6556 & n7083 ) ;
  assign n31419 = ~n12303 & n17745 ;
  assign n31420 = n31419 ^ n21038 ^ 1'b0 ;
  assign n31421 = n14963 ^ n4679 ^ 1'b0 ;
  assign n31422 = n14206 & ~n31421 ;
  assign n31426 = n31112 ^ n5589 ^ 1'b0 ;
  assign n31423 = n14038 & n22983 ;
  assign n31424 = n19997 & n31423 ;
  assign n31425 = n2346 & n31424 ;
  assign n31427 = n31426 ^ n31425 ^ n12312 ;
  assign n31428 = n12781 | n27507 ;
  assign n31429 = n1161 & n9760 ;
  assign n31430 = n31429 ^ n14106 ^ 1'b0 ;
  assign n31431 = n3472 & n24998 ;
  assign n31432 = n31431 ^ n30916 ^ 1'b0 ;
  assign n31433 = n23973 | n28772 ;
  assign n31434 = n4947 | n31433 ;
  assign n31435 = n16833 | n17113 ;
  assign n31436 = n24468 ^ n4328 ^ n390 ;
  assign n31437 = ( ~n25217 & n30074 ) | ( ~n25217 & n31436 ) | ( n30074 & n31436 ) ;
  assign n31439 = n4850 | n20191 ;
  assign n31440 = n31439 ^ n19163 ^ 1'b0 ;
  assign n31438 = n609 & ~n7953 ;
  assign n31441 = n31440 ^ n31438 ^ 1'b0 ;
  assign n31442 = n2313 | n8372 ;
  assign n31443 = n31442 ^ n13868 ^ 1'b0 ;
  assign n31444 = n6114 | n31443 ;
  assign n31445 = n3197 & ~n31444 ;
  assign n31446 = n31445 ^ n22789 ^ 1'b0 ;
  assign n31447 = n9090 & ~n23867 ;
  assign n31448 = n311 | n14305 ;
  assign n31449 = n31448 ^ n3609 ^ 1'b0 ;
  assign n31450 = n18417 & ~n31449 ;
  assign n31451 = ~n1297 & n31450 ;
  assign n31452 = n31451 ^ n9839 ^ 1'b0 ;
  assign n31453 = n7659 ^ n290 ^ 1'b0 ;
  assign n31454 = ~n5632 & n31453 ;
  assign n31458 = n19246 ^ n13855 ^ 1'b0 ;
  assign n31455 = n16568 ^ n12258 ^ 1'b0 ;
  assign n31456 = n29327 & n31455 ;
  assign n31457 = n31456 ^ n29564 ^ 1'b0 ;
  assign n31459 = n31458 ^ n31457 ^ n8124 ;
  assign n31460 = n17540 & ~n18039 ;
  assign n31461 = n31460 ^ n11954 ^ 1'b0 ;
  assign n31462 = n22691 ^ n44 ^ 1'b0 ;
  assign n31463 = n17632 & ~n31462 ;
  assign n31464 = n6145 ^ n5878 ^ 1'b0 ;
  assign n31465 = n12240 ^ n3080 ^ 1'b0 ;
  assign n31466 = n31464 & ~n31465 ;
  assign n31467 = n23905 ^ n14149 ^ 1'b0 ;
  assign n31468 = n31466 & ~n31467 ;
  assign n31469 = n19647 ^ n9049 ^ 1'b0 ;
  assign n31470 = n31468 & ~n31469 ;
  assign n31471 = ~n18496 & n31470 ;
  assign n31472 = n31471 ^ n7604 ^ 1'b0 ;
  assign n31473 = n7984 | n14395 ;
  assign n31474 = ( n24180 & n29590 ) | ( n24180 & ~n31473 ) | ( n29590 & ~n31473 ) ;
  assign n31475 = n31474 ^ n21389 ^ n10728 ;
  assign n31476 = n11014 ^ n5350 ^ 1'b0 ;
  assign n31477 = n19359 ^ n18650 ^ 1'b0 ;
  assign n31478 = ( ~n1545 & n31476 ) | ( ~n1545 & n31477 ) | ( n31476 & n31477 ) ;
  assign n31479 = ~n142 & n24553 ;
  assign n31480 = n31479 ^ n229 ^ 1'b0 ;
  assign n31481 = n30309 ^ n4395 ^ 1'b0 ;
  assign n31482 = n31480 & n31481 ;
  assign n31483 = n31482 ^ n4254 ^ 1'b0 ;
  assign n31484 = n22360 & n31483 ;
  assign n31485 = n31484 ^ n1636 ^ 1'b0 ;
  assign n31486 = n8565 | n12366 ;
  assign n31487 = n31486 ^ n16536 ^ 1'b0 ;
  assign n31488 = n31487 ^ n8757 ^ 1'b0 ;
  assign n31489 = n31488 ^ n17493 ^ 1'b0 ;
  assign n31490 = n31489 ^ n9192 ^ 1'b0 ;
  assign n31491 = n23647 & n24657 ;
  assign n31492 = n369 & n31491 ;
  assign n31493 = n482 & ~n7670 ;
  assign n31494 = n14480 & n31493 ;
  assign n31495 = n26671 & n31494 ;
  assign n31496 = n24545 ^ n24016 ^ 1'b0 ;
  assign n31497 = ~n13229 & n13279 ;
  assign n31498 = n31497 ^ n14311 ^ 1'b0 ;
  assign n31499 = n12553 & n31498 ;
  assign n31500 = n14426 & n31499 ;
  assign n31501 = n31500 ^ n22952 ^ 1'b0 ;
  assign n31502 = n3163 & n3992 ;
  assign n31503 = n31502 ^ n2159 ^ 1'b0 ;
  assign n31504 = n7499 & ~n31503 ;
  assign n31505 = n19931 ^ n19688 ^ n3939 ;
  assign n31506 = n5559 ^ n1816 ^ 1'b0 ;
  assign n31507 = ~n20458 & n31506 ;
  assign n31508 = n5598 & ~n31507 ;
  assign n31509 = n20500 & n21132 ;
  assign n31510 = n17741 ^ n13208 ^ n11997 ;
  assign n31511 = n4079 | n31510 ;
  assign n31512 = n3227 & ~n4691 ;
  assign n31513 = n1591 & n31512 ;
  assign n31514 = n7475 & n31513 ;
  assign n31515 = n31514 ^ n5045 ^ 1'b0 ;
  assign n31516 = n13342 & ~n31515 ;
  assign n31517 = ~n5334 & n31516 ;
  assign n31518 = n1880 | n27432 ;
  assign n31519 = n5277 & ~n31518 ;
  assign n31520 = n31519 ^ n17605 ^ 1'b0 ;
  assign n31521 = n20338 | n31520 ;
  assign n31522 = n31521 ^ n9088 ^ 1'b0 ;
  assign n31523 = n20138 & n31522 ;
  assign n31524 = n7397 & ~n19062 ;
  assign n31525 = n11900 ^ n9522 ^ 1'b0 ;
  assign n31526 = n609 & n31525 ;
  assign n31527 = n26542 & n31526 ;
  assign n31528 = n31527 ^ n12766 ^ 1'b0 ;
  assign n31531 = n6623 | n17841 ;
  assign n31529 = n8551 | n19402 ;
  assign n31530 = n31529 ^ n7876 ^ 1'b0 ;
  assign n31532 = n31531 ^ n31530 ^ 1'b0 ;
  assign n31533 = n21516 & n31532 ;
  assign n31534 = n23765 ^ n8737 ^ 1'b0 ;
  assign n31535 = n5091 & ~n31534 ;
  assign n31536 = n14523 | n17778 ;
  assign n31537 = n9258 & ~n31536 ;
  assign n31538 = ( n6489 & ~n25971 ) | ( n6489 & n31537 ) | ( ~n25971 & n31537 ) ;
  assign n31539 = n27137 ^ n606 ^ 1'b0 ;
  assign n31540 = n17477 | n31539 ;
  assign n31541 = n31538 & ~n31540 ;
  assign n31542 = ( n74 & n10479 ) | ( n74 & n26137 ) | ( n10479 & n26137 ) ;
  assign n31543 = n3488 & n13427 ;
  assign n31544 = ~n8344 & n10601 ;
  assign n31545 = ~n77 & n2053 ;
  assign n31546 = n31545 ^ n24079 ^ 1'b0 ;
  assign n31547 = n21981 & n22681 ;
  assign n31548 = n9916 & n11446 ;
  assign n31549 = n21748 ^ n8219 ^ 1'b0 ;
  assign n31550 = n31549 ^ n25070 ^ 1'b0 ;
  assign n31551 = n31548 & n31550 ;
  assign n31552 = ~n22819 & n27060 ;
  assign n31553 = n4800 ^ n294 ^ 1'b0 ;
  assign n31554 = ~n3047 & n31553 ;
  assign n31555 = ( n10449 & n12015 ) | ( n10449 & n31554 ) | ( n12015 & n31554 ) ;
  assign n31556 = n31552 & ~n31555 ;
  assign n31557 = n25784 ^ n14063 ^ 1'b0 ;
  assign n31558 = ~n20539 & n31557 ;
  assign n31559 = n19615 ^ n13480 ^ n2671 ;
  assign n31560 = n22776 ^ n6834 ^ 1'b0 ;
  assign n31561 = ~n10399 & n15571 ;
  assign n31562 = n15261 ^ n7303 ^ 1'b0 ;
  assign n31564 = ~n2781 & n5350 ;
  assign n31565 = n31564 ^ n294 ^ 1'b0 ;
  assign n31563 = n9069 & ~n16473 ;
  assign n31566 = n31565 ^ n31563 ^ 1'b0 ;
  assign n31567 = n13331 & ~n31566 ;
  assign n31568 = n29602 ^ n12198 ^ 1'b0 ;
  assign n31569 = ~n1079 & n31568 ;
  assign n31570 = n1003 | n28056 ;
  assign n31571 = n31570 ^ n5281 ^ 1'b0 ;
  assign n31572 = n3319 & n15719 ;
  assign n31573 = n4141 & n31572 ;
  assign n31574 = n31573 ^ n21775 ^ 1'b0 ;
  assign n31575 = n29399 & ~n31574 ;
  assign n31576 = n31571 & n31575 ;
  assign n31577 = n17554 ^ n8367 ^ 1'b0 ;
  assign n31578 = ~n31576 & n31577 ;
  assign n31579 = n13843 & n31578 ;
  assign n31580 = n22712 ^ n2202 ^ 1'b0 ;
  assign n31581 = n9643 & n31580 ;
  assign n31582 = ~n1631 & n31581 ;
  assign n31583 = ~n10115 & n22704 ;
  assign n31584 = n31583 ^ n27884 ^ 1'b0 ;
  assign n31585 = n1497 & n10761 ;
  assign n31586 = ( n22552 & ~n23226 ) | ( n22552 & n27591 ) | ( ~n23226 & n27591 ) ;
  assign n31587 = n12038 & n25119 ;
  assign n31588 = n8747 & ~n17155 ;
  assign n31589 = n31588 ^ n11318 ^ 1'b0 ;
  assign n31590 = n7816 ^ n493 ^ 1'b0 ;
  assign n31591 = n17449 | n31590 ;
  assign n31592 = n25044 | n31591 ;
  assign n31593 = n16170 & ~n31592 ;
  assign n31594 = n502 & n7889 ;
  assign n31595 = n31594 ^ n14268 ^ 1'b0 ;
  assign n31596 = n30355 ^ n24493 ^ 1'b0 ;
  assign n31597 = n3915 | n17228 ;
  assign n31598 = n31597 ^ n774 ^ 1'b0 ;
  assign n31599 = n31391 ^ n5541 ^ 1'b0 ;
  assign n31600 = n31598 & n31599 ;
  assign n31601 = n2812 & ~n5469 ;
  assign n31602 = n31601 ^ n7871 ^ 1'b0 ;
  assign n31603 = n26002 & ~n31602 ;
  assign n31604 = n16769 & n31603 ;
  assign n31605 = n13223 ^ n10882 ^ n61 ;
  assign n31606 = n1210 | n7480 ;
  assign n31607 = n31605 & ~n31606 ;
  assign n31610 = n4263 & n26951 ;
  assign n31608 = n15426 ^ n10883 ^ 1'b0 ;
  assign n31609 = n31143 & n31608 ;
  assign n31611 = n31610 ^ n31609 ^ 1'b0 ;
  assign n31612 = n25222 ^ n4263 ^ 1'b0 ;
  assign n31613 = n5348 ^ n2630 ^ 1'b0 ;
  assign n31614 = n15342 & ~n31613 ;
  assign n31615 = n6941 & n31614 ;
  assign n31616 = n23523 & ~n23583 ;
  assign n31617 = n6947 | n9251 ;
  assign n31618 = ( n9288 & n11074 ) | ( n9288 & n31617 ) | ( n11074 & n31617 ) ;
  assign n31619 = ~n21125 & n31466 ;
  assign n31620 = ~n5991 & n16361 ;
  assign n31621 = n23054 & n31620 ;
  assign n31622 = ~n18626 & n21941 ;
  assign n31623 = n2002 & n31622 ;
  assign n31624 = n29542 & n31623 ;
  assign n31625 = n13386 & ~n22432 ;
  assign n31626 = ( n7602 & n10544 ) | ( n7602 & ~n31625 ) | ( n10544 & ~n31625 ) ;
  assign n31627 = n30639 & n31626 ;
  assign n31628 = ~n8055 & n31627 ;
  assign n31629 = n4501 ^ n1987 ^ 1'b0 ;
  assign n31630 = ~n10272 & n31629 ;
  assign n31631 = n12379 & n31630 ;
  assign n31632 = n13451 ^ n4365 ^ n74 ;
  assign n31633 = n31476 ^ n5898 ^ 1'b0 ;
  assign n31634 = ~n16525 & n31633 ;
  assign n31635 = ~n2843 & n20294 ;
  assign n31636 = ~n16408 & n31635 ;
  assign n31637 = n14778 ^ n6738 ^ 1'b0 ;
  assign n31638 = ~n25385 & n25584 ;
  assign n31639 = n12832 & n31638 ;
  assign n31640 = n31639 ^ n16244 ^ 1'b0 ;
  assign n31641 = n22531 & ~n31640 ;
  assign n31642 = ~n16670 & n26858 ;
  assign n31643 = n1570 | n4657 ;
  assign n31644 = n31642 & n31643 ;
  assign n31647 = n20649 ^ n4947 ^ n1264 ;
  assign n31645 = n16580 ^ n3720 ^ n3369 ;
  assign n31646 = ( n25719 & n27418 ) | ( n25719 & n31645 ) | ( n27418 & n31645 ) ;
  assign n31648 = n31647 ^ n31646 ^ n18538 ;
  assign n31649 = ~n10094 & n17874 ;
  assign n31650 = n20976 ^ n11290 ^ 1'b0 ;
  assign n31651 = ~n5981 & n10716 ;
  assign n31652 = ~n6009 & n25300 ;
  assign n31653 = ~n22934 & n31652 ;
  assign n31654 = n6768 & n21347 ;
  assign n31655 = n31654 ^ n7583 ^ 1'b0 ;
  assign n31656 = n10762 & ~n23770 ;
  assign n31657 = n6384 ^ n2778 ^ 1'b0 ;
  assign n31658 = n28278 | n31657 ;
  assign n31659 = n31658 ^ n404 ^ 1'b0 ;
  assign n31660 = n3352 & ~n7455 ;
  assign n31661 = ~n3352 & n31660 ;
  assign n31662 = ~n732 & n31661 ;
  assign n31665 = n2275 ^ n2267 ^ 1'b0 ;
  assign n31666 = n5543 | n31665 ;
  assign n31667 = n5543 & ~n31666 ;
  assign n31668 = n31667 ^ n16004 ^ 1'b0 ;
  assign n31663 = n7208 | n8362 ;
  assign n31664 = n8362 & ~n31663 ;
  assign n31669 = n31668 ^ n31664 ^ 1'b0 ;
  assign n31670 = n31662 | n31669 ;
  assign n31672 = n4555 & n6919 ;
  assign n31673 = n31672 ^ n12442 ^ 1'b0 ;
  assign n31674 = n31673 ^ n15426 ^ n3315 ;
  assign n31671 = n4260 & n19416 ;
  assign n31675 = n31674 ^ n31671 ^ 1'b0 ;
  assign n31676 = ~n4681 & n13274 ;
  assign n31677 = ~n12860 & n23478 ;
  assign n31678 = n11636 & n31677 ;
  assign n31679 = ~n12126 & n28816 ;
  assign n31680 = ~n2425 & n31679 ;
  assign n31681 = n10654 & ~n14598 ;
  assign n31682 = ~n8304 & n31681 ;
  assign n31683 = ~n9886 & n20682 ;
  assign n31684 = n31682 & n31683 ;
  assign n31685 = n163 & n1897 ;
  assign n31686 = n21308 & ~n24179 ;
  assign n31697 = n3644 | n10473 ;
  assign n31698 = n3644 & ~n31697 ;
  assign n31699 = n6110 | n8243 ;
  assign n31700 = n31698 & ~n31699 ;
  assign n31701 = n4429 | n31700 ;
  assign n31702 = n4429 & ~n31701 ;
  assign n31694 = ~n5097 & n8127 ;
  assign n31695 = ~n8127 & n31694 ;
  assign n31696 = n13821 | n31695 ;
  assign n31703 = n31702 ^ n31696 ^ 1'b0 ;
  assign n31687 = n1660 & n2277 ;
  assign n31688 = n11719 & n31687 ;
  assign n31689 = ~n2735 & n25504 ;
  assign n31690 = ~n25504 & n31689 ;
  assign n31691 = n31690 ^ n10543 ^ 1'b0 ;
  assign n31692 = n21554 | n31691 ;
  assign n31693 = n31688 & ~n31692 ;
  assign n31704 = n31703 ^ n31693 ^ n31573 ;
  assign n31705 = n2019 | n3202 ;
  assign n31706 = n478 | n31705 ;
  assign n31707 = n23115 & ~n31706 ;
  assign n31708 = n12059 | n31451 ;
  assign n31709 = n1152 ^ n692 ^ 1'b0 ;
  assign n31710 = n11841 ^ n7703 ^ 1'b0 ;
  assign n31711 = n3619 & n15586 ;
  assign n31712 = n31711 ^ n19677 ^ 1'b0 ;
  assign n31713 = n11383 ^ n7704 ^ 1'b0 ;
  assign n31714 = n609 | n31713 ;
  assign n31715 = n27674 ^ n6436 ^ 1'b0 ;
  assign n31716 = ~n10330 & n31715 ;
  assign n31717 = n31716 ^ n8388 ^ 1'b0 ;
  assign n31718 = n5805 | n17642 ;
  assign n31719 = n31718 ^ n1588 ^ 1'b0 ;
  assign n31721 = ( n8399 & ~n8462 ) | ( n8399 & n28034 ) | ( ~n8462 & n28034 ) ;
  assign n31720 = n9584 | n22020 ;
  assign n31722 = n31721 ^ n31720 ^ 1'b0 ;
  assign n31723 = n5402 & ~n25725 ;
  assign n31724 = n31723 ^ n3902 ^ 1'b0 ;
  assign n31725 = ~n8758 & n31724 ;
  assign n31726 = n31725 ^ n23898 ^ 1'b0 ;
  assign n31727 = n1477 & n4261 ;
  assign n31728 = n31727 ^ n21249 ^ 1'b0 ;
  assign n31729 = ~n2703 & n31728 ;
  assign n31730 = n31729 ^ n1018 ^ 1'b0 ;
  assign n31731 = n31730 ^ n14134 ^ 1'b0 ;
  assign n31732 = n19645 & n31334 ;
  assign n31733 = n6927 & ~n19094 ;
  assign n31734 = n16389 & n31733 ;
  assign n31735 = n21035 ^ n5825 ^ 1'b0 ;
  assign n31736 = ~n6023 & n31735 ;
  assign n31737 = n31736 ^ n3671 ^ 1'b0 ;
  assign n31738 = n414 & ~n30012 ;
  assign n31739 = n7368 | n18498 ;
  assign n31740 = ~n3748 & n28363 ;
  assign n31741 = n4299 & n23517 ;
  assign n31742 = n31741 ^ n3030 ^ 1'b0 ;
  assign n31743 = n14456 ^ n3023 ^ 1'b0 ;
  assign n31744 = n10295 | n31743 ;
  assign n31745 = n31744 ^ n7367 ^ 1'b0 ;
  assign n31747 = ~n3367 & n30049 ;
  assign n31748 = n1823 & ~n31747 ;
  assign n31749 = n31748 ^ n8413 ^ 1'b0 ;
  assign n31746 = n24035 & n31404 ;
  assign n31750 = n31749 ^ n31746 ^ 1'b0 ;
  assign n31751 = n31750 ^ n29058 ^ 1'b0 ;
  assign n31752 = n12157 & n23555 ;
  assign n31753 = n14303 | n19725 ;
  assign n31754 = n3122 ^ n2282 ^ 1'b0 ;
  assign n31755 = ~n667 & n31754 ;
  assign n31756 = n25571 ^ n3047 ^ 1'b0 ;
  assign n31757 = n31756 ^ n16896 ^ 1'b0 ;
  assign n31758 = n31755 & ~n31757 ;
  assign n31759 = n31758 ^ n16204 ^ 1'b0 ;
  assign n31760 = n13545 ^ n5378 ^ 1'b0 ;
  assign n31761 = n31760 ^ n15388 ^ n6927 ;
  assign n31762 = n18519 | n31761 ;
  assign n31763 = n8404 & ~n31762 ;
  assign n31764 = n3071 | n21769 ;
  assign n31765 = n12202 & n23031 ;
  assign n31766 = n17193 & n22082 ;
  assign n31767 = ( n6337 & n9983 ) | ( n6337 & ~n21632 ) | ( n9983 & ~n21632 ) ;
  assign n31768 = n31767 ^ n21564 ^ 1'b0 ;
  assign n31769 = n31766 & n31768 ;
  assign n31770 = ~n10473 & n29893 ;
  assign n31771 = ( n3221 & ~n9282 ) | ( n3221 & n25793 ) | ( ~n9282 & n25793 ) ;
  assign n31772 = n2706 & ~n31771 ;
  assign n31773 = n2356 & n31772 ;
  assign n31774 = ~n770 & n2468 ;
  assign n31775 = n20662 ^ n1644 ^ 1'b0 ;
  assign n31776 = n14887 & ~n31775 ;
  assign n31777 = ~n21596 & n31776 ;
  assign n31778 = n31777 ^ n844 ^ 1'b0 ;
  assign n31779 = ~n8814 & n31778 ;
  assign n31780 = n31779 ^ n4750 ^ 1'b0 ;
  assign n31781 = n1511 & ~n3641 ;
  assign n31782 = ~n13569 & n31781 ;
  assign n31783 = n6954 & ~n31782 ;
  assign n31784 = n1377 & ~n5388 ;
  assign n31785 = ( n2048 & ~n10499 ) | ( n2048 & n11470 ) | ( ~n10499 & n11470 ) ;
  assign n31786 = n6610 | n26229 ;
  assign n31787 = n31785 & n31786 ;
  assign n31788 = ~n16395 & n26419 ;
  assign n31789 = n11803 ^ n1165 ^ 1'b0 ;
  assign n31790 = n31789 ^ n2103 ^ 1'b0 ;
  assign n31791 = n31788 & ~n31790 ;
  assign n31792 = ~n14259 & n22474 ;
  assign n31793 = n25170 ^ n15109 ^ 1'b0 ;
  assign n31794 = n31793 ^ n2832 ^ 1'b0 ;
  assign n31796 = n4077 & ~n11013 ;
  assign n31797 = n31796 ^ n28103 ^ 1'b0 ;
  assign n31795 = n687 & n4613 ;
  assign n31798 = n31797 ^ n31795 ^ 1'b0 ;
  assign n31799 = n31794 & n31798 ;
  assign n31800 = n9209 & ~n9884 ;
  assign n31801 = n31800 ^ n10281 ^ 1'b0 ;
  assign n31802 = ~n4748 & n29213 ;
  assign n31803 = n7544 & ~n17339 ;
  assign n31804 = n23619 & ~n31803 ;
  assign n31805 = n29146 ^ n785 ^ 1'b0 ;
  assign n31806 = n4301 | n31805 ;
  assign n31807 = n29730 ^ n11286 ^ 1'b0 ;
  assign n31808 = n9837 ^ n5439 ^ n1322 ;
  assign n31809 = n31808 ^ n16966 ^ 1'b0 ;
  assign n31810 = n8507 ^ n1116 ^ 1'b0 ;
  assign n31811 = ~n11121 & n31810 ;
  assign n31812 = n6380 ^ n1312 ^ 1'b0 ;
  assign n31813 = n10119 ^ n2674 ^ 1'b0 ;
  assign n31814 = ~n31812 & n31813 ;
  assign n31815 = n21339 ^ n4038 ^ 1'b0 ;
  assign n31816 = n31603 & ~n31815 ;
  assign n31817 = n657 & n31816 ;
  assign n31818 = n8534 & n31817 ;
  assign n31819 = n44 & ~n31193 ;
  assign n31820 = ~n31818 & n31819 ;
  assign n31821 = n1653 & ~n21127 ;
  assign n31822 = n31821 ^ n10634 ^ 1'b0 ;
  assign n31823 = n10965 | n13774 ;
  assign n31824 = n13393 | n31823 ;
  assign n31825 = ~n3713 & n7919 ;
  assign n31826 = ~n31824 & n31825 ;
  assign n31827 = n3884 & ~n4090 ;
  assign n31828 = n31827 ^ n13380 ^ 1'b0 ;
  assign n31829 = ~n2217 & n2769 ;
  assign n31830 = n31829 ^ n20005 ^ n16606 ;
  assign n31831 = ~n8688 & n20739 ;
  assign n31832 = n1391 | n31831 ;
  assign n31834 = n7466 | n9344 ;
  assign n31833 = n11791 & n24561 ;
  assign n31835 = n31834 ^ n31833 ^ 1'b0 ;
  assign n31836 = n17253 ^ n2124 ^ 1'b0 ;
  assign n31837 = n11529 | n31836 ;
  assign n31838 = ( n6762 & n9371 ) | ( n6762 & ~n26121 ) | ( n9371 & ~n26121 ) ;
  assign n31839 = n965 & ~n3738 ;
  assign n31840 = n6470 & ~n31839 ;
  assign n31841 = n5157 ^ n4214 ^ 1'b0 ;
  assign n31842 = n31015 ^ n18414 ^ 1'b0 ;
  assign n31843 = n31841 | n31842 ;
  assign n31844 = n12644 ^ n7317 ^ 1'b0 ;
  assign n31845 = n244 | n21229 ;
  assign n31846 = ( n466 & n10298 ) | ( n466 & n14396 ) | ( n10298 & n14396 ) ;
  assign n31847 = n7369 & ~n9851 ;
  assign n31851 = n326 & n3006 ;
  assign n31852 = n31851 ^ n4252 ^ 1'b0 ;
  assign n31853 = n31852 ^ n6716 ^ 1'b0 ;
  assign n31854 = n7876 & ~n31853 ;
  assign n31848 = n10956 ^ n3278 ^ n1816 ;
  assign n31849 = n31848 ^ n2137 ^ n1586 ;
  assign n31850 = ( ~n631 & n16874 ) | ( ~n631 & n31849 ) | ( n16874 & n31849 ) ;
  assign n31855 = n31854 ^ n31850 ^ 1'b0 ;
  assign n31856 = n22959 ^ n13026 ^ n5399 ;
  assign n31857 = n30417 ^ n20472 ^ n12309 ;
  assign n31858 = n6314 & n30725 ;
  assign n31859 = n31858 ^ n443 ^ 1'b0 ;
  assign n31860 = ~n2265 & n31859 ;
  assign n31861 = ~n8436 & n31860 ;
  assign n31862 = n1374 & ~n8630 ;
  assign n31863 = n31862 ^ n1010 ^ 1'b0 ;
  assign n31864 = n11193 | n31863 ;
  assign n31865 = n1816 | n22147 ;
  assign n31866 = n31865 ^ n22214 ^ 1'b0 ;
  assign n31867 = n28863 ^ n18664 ^ n3150 ;
  assign n31868 = n31867 ^ n26977 ^ 1'b0 ;
  assign n31869 = n21393 ^ n9557 ^ 1'b0 ;
  assign n31870 = n12514 | n29524 ;
  assign n31871 = n17014 & ~n31870 ;
  assign n31872 = n30457 ^ n20498 ^ n9156 ;
  assign n31873 = ( n3930 & n13193 ) | ( n3930 & ~n31872 ) | ( n13193 & ~n31872 ) ;
  assign n31874 = ( n4637 & n6809 ) | ( n4637 & ~n9192 ) | ( n6809 & ~n9192 ) ;
  assign n31875 = n9208 & n14968 ;
  assign n31876 = n31875 ^ n23827 ^ 1'b0 ;
  assign n31877 = n18273 | n27287 ;
  assign n31883 = n5367 & ~n7004 ;
  assign n31884 = n31883 ^ n20927 ^ 1'b0 ;
  assign n31885 = n31884 ^ n31105 ^ n7007 ;
  assign n31878 = n2796 ^ n2356 ^ 1'b0 ;
  assign n31879 = ~n9674 & n31878 ;
  assign n31880 = n2095 & n31879 ;
  assign n31881 = n31880 ^ n13785 ^ 1'b0 ;
  assign n31882 = ~n8814 & n31881 ;
  assign n31886 = n31885 ^ n31882 ^ 1'b0 ;
  assign n31887 = n19769 & n27973 ;
  assign n31888 = n31887 ^ n14351 ^ 1'b0 ;
  assign n31889 = n29772 & n31888 ;
  assign n31890 = ( n4738 & n5888 ) | ( n4738 & ~n18825 ) | ( n5888 & ~n18825 ) ;
  assign n31891 = n20816 | n23919 ;
  assign n31892 = n31890 | n31891 ;
  assign n31893 = ~n12067 & n15087 ;
  assign n31894 = n19173 | n31893 ;
  assign n31895 = n12395 ^ n7827 ^ 1'b0 ;
  assign n31896 = n28275 & ~n31895 ;
  assign n31898 = n16517 ^ n8728 ^ n3672 ;
  assign n31897 = ( n253 & n682 ) | ( n253 & n8303 ) | ( n682 & n8303 ) ;
  assign n31899 = n31898 ^ n31897 ^ n7556 ;
  assign n31900 = n7322 & ~n31899 ;
  assign n31901 = n14311 | n15272 ;
  assign n31902 = n31901 ^ n3955 ^ 1'b0 ;
  assign n31903 = ~n3115 & n31902 ;
  assign n31904 = n30409 | n31903 ;
  assign n31905 = n12525 | n13545 ;
  assign n31906 = n130 & n708 ;
  assign n31907 = ~n29632 & n31906 ;
  assign n31908 = ( ~n23966 & n26941 ) | ( ~n23966 & n31907 ) | ( n26941 & n31907 ) ;
  assign n31909 = n7676 & n21651 ;
  assign n31910 = ~n8972 & n26441 ;
  assign n31911 = ~n14378 & n31910 ;
  assign n31912 = n11813 & ~n12053 ;
  assign n31913 = n3726 & n31912 ;
  assign n31914 = n4914 & n15317 ;
  assign n31915 = ~n7265 & n31914 ;
  assign n31916 = ~n4586 & n20191 ;
  assign n31917 = n8122 ^ n4280 ^ 1'b0 ;
  assign n31918 = n2694 | n31917 ;
  assign n31919 = n22939 ^ n898 ^ 1'b0 ;
  assign n31920 = n31919 ^ n8057 ^ 1'b0 ;
  assign n31921 = n14338 & n31920 ;
  assign n31922 = ( n9321 & n31918 ) | ( n9321 & n31921 ) | ( n31918 & n31921 ) ;
  assign n31923 = n18286 ^ n3252 ^ 1'b0 ;
  assign n31924 = n6449 & ~n31923 ;
  assign n31925 = n26638 ^ n16290 ^ 1'b0 ;
  assign n31926 = n31925 ^ n1116 ^ n356 ;
  assign n31927 = n8860 & ~n24071 ;
  assign n31928 = n4114 & ~n31927 ;
  assign n31929 = n14208 & n18127 ;
  assign n31930 = n17320 & n31929 ;
  assign n31931 = ~n996 & n5452 ;
  assign n31932 = ~n3744 & n31931 ;
  assign n31933 = n18268 ^ n6844 ^ 1'b0 ;
  assign n31934 = n31932 & ~n31933 ;
  assign n31935 = n25608 ^ n14291 ^ 1'b0 ;
  assign n31936 = n2065 & n17461 ;
  assign n31937 = n31936 ^ n15246 ^ 1'b0 ;
  assign n31938 = ~n4937 & n14875 ;
  assign n31939 = n31938 ^ n14726 ^ 1'b0 ;
  assign n31940 = n31939 ^ n31643 ^ 1'b0 ;
  assign n31941 = ~n14468 & n31940 ;
  assign n31942 = n3725 | n9709 ;
  assign n31943 = n31942 ^ n12692 ^ 1'b0 ;
  assign n31944 = n31943 ^ n9600 ^ 1'b0 ;
  assign n31945 = ~n10510 & n31944 ;
  assign n31946 = n1539 & ~n16148 ;
  assign n31947 = ~n110 & n5058 ;
  assign n31948 = ~n17209 & n31947 ;
  assign n31949 = ~n14356 & n31948 ;
  assign n31950 = n18217 ^ n12729 ^ 1'b0 ;
  assign n31951 = n7357 & ~n27906 ;
  assign n31952 = n445 | n31951 ;
  assign n31953 = n31952 ^ n28678 ^ 1'b0 ;
  assign n31954 = n16325 ^ n2063 ^ 1'b0 ;
  assign n31955 = n31954 ^ n7707 ^ 1'b0 ;
  assign n31956 = n3163 & ~n6381 ;
  assign n31957 = n31956 ^ n2540 ^ 1'b0 ;
  assign n31958 = n31957 ^ n23490 ^ 1'b0 ;
  assign n31960 = n255 | n890 ;
  assign n31961 = n890 & ~n31960 ;
  assign n31959 = n11954 & n14632 ;
  assign n31962 = n31961 ^ n31959 ^ 1'b0 ;
  assign n31963 = ( n6750 & ~n9178 ) | ( n6750 & n31962 ) | ( ~n9178 & n31962 ) ;
  assign n31964 = n31963 ^ n27243 ^ 1'b0 ;
  assign n31965 = n4859 & ~n30158 ;
  assign n31966 = ( n21534 & ~n23312 ) | ( n21534 & n31965 ) | ( ~n23312 & n31965 ) ;
  assign n31967 = ( ~n8909 & n14851 ) | ( ~n8909 & n18951 ) | ( n14851 & n18951 ) ;
  assign n31968 = n26317 | n28685 ;
  assign n31969 = n13 | n17511 ;
  assign n31970 = n13951 | n31969 ;
  assign n31971 = n10106 | n31970 ;
  assign n31972 = n14861 ^ n6279 ^ 1'b0 ;
  assign n31973 = n27353 & n31972 ;
  assign n31974 = n31973 ^ n31856 ^ 1'b0 ;
  assign n31975 = n3455 ^ n1226 ^ 1'b0 ;
  assign n31976 = ( n6470 & ~n12856 ) | ( n6470 & n31975 ) | ( ~n12856 & n31975 ) ;
  assign n31977 = n9386 & ~n15387 ;
  assign n31978 = ~n9051 & n31977 ;
  assign n31979 = n31978 ^ n20574 ^ 1'b0 ;
  assign n31980 = n398 & n25025 ;
  assign n31981 = n31980 ^ n1207 ^ 1'b0 ;
  assign n31982 = n24328 ^ n23761 ^ 1'b0 ;
  assign n31983 = ~n1414 & n5493 ;
  assign n31984 = n7962 ^ n7071 ^ 1'b0 ;
  assign n31985 = ( n4962 & ~n14924 ) | ( n4962 & n19148 ) | ( ~n14924 & n19148 ) ;
  assign n31986 = n10713 & ~n12275 ;
  assign n31987 = n31986 ^ n115 ^ 1'b0 ;
  assign n31988 = n28 & n14213 ;
  assign n31989 = ~n3891 & n31988 ;
  assign n31990 = n17860 ^ n2101 ^ 1'b0 ;
  assign n31991 = n5005 | n28968 ;
  assign n31992 = n23093 & ~n31991 ;
  assign n31993 = n9894 & ~n29052 ;
  assign n31994 = n31993 ^ n25812 ^ 1'b0 ;
  assign n31995 = n10944 ^ n1182 ^ 1'b0 ;
  assign n31996 = ~n6472 & n11578 ;
  assign n31997 = n15844 ^ n741 ^ 1'b0 ;
  assign n32000 = n1485 | n24550 ;
  assign n31998 = n6396 & ~n11044 ;
  assign n31999 = ~n17201 & n31998 ;
  assign n32001 = n32000 ^ n31999 ^ 1'b0 ;
  assign n32002 = n3020 | n23295 ;
  assign n32003 = n25201 & ~n32002 ;
  assign n32004 = n8647 ^ n5860 ^ 1'b0 ;
  assign n32005 = n8454 & ~n32004 ;
  assign n32006 = n28878 ^ n2867 ^ 1'b0 ;
  assign n32007 = n4451 ^ n451 ^ 1'b0 ;
  assign n32008 = n7110 | n7914 ;
  assign n32010 = n11044 & ~n12024 ;
  assign n32009 = n26009 ^ n4746 ^ 1'b0 ;
  assign n32011 = n32010 ^ n32009 ^ 1'b0 ;
  assign n32012 = n9598 & ~n32011 ;
  assign n32013 = n8830 | n28205 ;
  assign n32014 = n8830 & ~n32013 ;
  assign n32015 = ~n13138 & n32014 ;
  assign n32016 = n1841 & n2799 ;
  assign n32017 = ~n2799 & n32016 ;
  assign n32018 = n27253 & ~n32017 ;
  assign n32019 = ~n27253 & n32018 ;
  assign n32020 = n24172 & ~n32019 ;
  assign n32021 = n32020 ^ n10411 ^ 1'b0 ;
  assign n32022 = n32015 & n32021 ;
  assign n32023 = n30555 ^ n9631 ^ 1'b0 ;
  assign n32024 = n2403 & n32023 ;
  assign n32025 = n9808 ^ n402 ^ 1'b0 ;
  assign n32026 = n5118 & ~n32025 ;
  assign n32027 = n20005 & n20113 ;
  assign n32028 = n22010 & n32027 ;
  assign n32029 = n7611 | n14748 ;
  assign n32030 = n32029 ^ n23 ^ 1'b0 ;
  assign n32031 = ~n10944 & n32030 ;
  assign n32032 = ~n2051 & n32031 ;
  assign n32033 = n2634 & n32032 ;
  assign n32034 = n21733 ^ n15698 ^ 1'b0 ;
  assign n32035 = n32033 & n32034 ;
  assign n32036 = n2273 & ~n10610 ;
  assign n32037 = n3111 & n11836 ;
  assign n32038 = n32037 ^ n18231 ^ 1'b0 ;
  assign n32039 = n17244 | n32038 ;
  assign n32040 = ( ~n14345 & n19966 ) | ( ~n14345 & n32039 ) | ( n19966 & n32039 ) ;
  assign n32041 = ( n1237 & ~n1603 ) | ( n1237 & n1832 ) | ( ~n1603 & n1832 ) ;
  assign n32042 = n18502 & ~n25420 ;
  assign n32043 = n150 & n29910 ;
  assign n32044 = n20002 ^ n5886 ^ 1'b0 ;
  assign n32045 = n32044 ^ n30414 ^ n16640 ;
  assign n32046 = n6088 ^ n2093 ^ n917 ;
  assign n32047 = n25593 ^ n8675 ^ 1'b0 ;
  assign n32048 = n32046 | n32047 ;
  assign n32049 = n32048 ^ n2080 ^ 1'b0 ;
  assign n32050 = n32049 ^ n31517 ^ 1'b0 ;
  assign n32051 = ~n3209 & n6630 ;
  assign n32052 = n6560 ^ n4780 ^ 1'b0 ;
  assign n32053 = ~n13259 & n32052 ;
  assign n32054 = n32051 & n32053 ;
  assign n32055 = n7624 ^ n582 ^ 1'b0 ;
  assign n32056 = n16580 | n32055 ;
  assign n32057 = n23552 | n32056 ;
  assign n32058 = n2989 | n17189 ;
  assign n32059 = n32058 ^ n5422 ^ 1'b0 ;
  assign n32060 = n7788 & ~n19413 ;
  assign n32061 = ( n1184 & n32059 ) | ( n1184 & n32060 ) | ( n32059 & n32060 ) ;
  assign n32062 = n1395 & ~n25720 ;
  assign n32063 = n887 & n32062 ;
  assign n32064 = n31524 ^ n11238 ^ 1'b0 ;
  assign n32065 = n20880 | n23160 ;
  assign n32066 = n12201 & n28249 ;
  assign n32067 = ( n15442 & n21331 ) | ( n15442 & n32066 ) | ( n21331 & n32066 ) ;
  assign n32068 = n12201 ^ n6953 ^ 1'b0 ;
  assign n32069 = n1035 & n13996 ;
  assign n32070 = n2570 & n32069 ;
  assign n32071 = n32070 ^ n828 ^ 1'b0 ;
  assign n32072 = n6917 & ~n32071 ;
  assign n32073 = n32072 ^ n12938 ^ 1'b0 ;
  assign n32074 = ~n16062 & n20419 ;
  assign n32075 = n4785 & n32074 ;
  assign n32076 = ( ~n14094 & n22501 ) | ( ~n14094 & n32075 ) | ( n22501 & n32075 ) ;
  assign n32077 = n7797 & n13901 ;
  assign n32080 = ( n454 & ~n14478 ) | ( n454 & n16835 ) | ( ~n14478 & n16835 ) ;
  assign n32081 = n28301 & ~n29311 ;
  assign n32082 = n32080 & n32081 ;
  assign n32078 = n19973 ^ n2798 ^ 1'b0 ;
  assign n32079 = ~n3741 & n32078 ;
  assign n32083 = n32082 ^ n32079 ^ 1'b0 ;
  assign n32084 = n2802 | n4348 ;
  assign n32085 = n1862 & n3027 ;
  assign n32086 = ~n32084 & n32085 ;
  assign n32087 = ~n6488 & n32086 ;
  assign n32088 = n31287 | n32087 ;
  assign n32089 = n12825 | n32088 ;
  assign n32090 = ~n817 & n18492 ;
  assign n32091 = n32090 ^ n28816 ^ n15972 ;
  assign n32092 = ( n7749 & n12105 ) | ( n7749 & ~n26543 ) | ( n12105 & ~n26543 ) ;
  assign n32093 = ( n11479 & n24172 ) | ( n11479 & ~n32092 ) | ( n24172 & ~n32092 ) ;
  assign n32094 = n21393 ^ n15614 ^ 1'b0 ;
  assign n32095 = ~n6108 & n32094 ;
  assign n32096 = n4346 & n14872 ;
  assign n32097 = n22217 & n32096 ;
  assign n32098 = n20382 & ~n32097 ;
  assign n32099 = n9377 & n32098 ;
  assign n32100 = ~n218 & n4899 ;
  assign n32101 = n32100 ^ n20545 ^ 1'b0 ;
  assign n32102 = n32101 ^ n5406 ^ 1'b0 ;
  assign n32103 = ~n17474 & n28030 ;
  assign n32104 = n7132 & n8169 ;
  assign n32105 = n11917 & n24156 ;
  assign n32106 = n32104 & n32105 ;
  assign n32107 = n8153 ^ n6959 ^ 1'b0 ;
  assign n32108 = ~n32106 & n32107 ;
  assign n32109 = ( n12354 & n16197 ) | ( n12354 & n23203 ) | ( n16197 & n23203 ) ;
  assign n32110 = n1216 & ~n8906 ;
  assign n32111 = n19334 ^ n15413 ^ n1571 ;
  assign n32112 = n7245 | n9883 ;
  assign n32113 = n20397 | n32112 ;
  assign n32114 = n1839 | n21505 ;
  assign n32115 = ( n1868 & n2438 ) | ( n1868 & ~n24439 ) | ( n2438 & ~n24439 ) ;
  assign n32116 = n22347 ^ n3384 ^ 1'b0 ;
  assign n32117 = n2254 | n32116 ;
  assign n32118 = n6437 & ~n32117 ;
  assign n32119 = n9660 ^ n472 ^ 1'b0 ;
  assign n32120 = ~n32118 & n32119 ;
  assign n32121 = n5765 & n32120 ;
  assign n32122 = n56 & n6933 ;
  assign n32123 = n32122 ^ n4676 ^ 1'b0 ;
  assign n32124 = ~n226 & n32123 ;
  assign n32125 = n12137 ^ n7404 ^ 1'b0 ;
  assign n32126 = n3034 & n7674 ;
  assign n32127 = ~n32125 & n32126 ;
  assign n32128 = ~n17831 & n32127 ;
  assign n32129 = n5012 & n6910 ;
  assign n32130 = n18950 ^ n5250 ^ 1'b0 ;
  assign n32131 = n32129 & n32130 ;
  assign n32132 = n22954 ^ n6360 ^ 1'b0 ;
  assign n32133 = n19513 & n32132 ;
  assign n32134 = ( ~n2199 & n31789 ) | ( ~n2199 & n32133 ) | ( n31789 & n32133 ) ;
  assign n32135 = n3915 ^ n2277 ^ 1'b0 ;
  assign n32136 = n18171 | n32135 ;
  assign n32137 = n8212 | n23027 ;
  assign n32138 = n25279 ^ n18113 ^ 1'b0 ;
  assign n32139 = n32137 & ~n32138 ;
  assign n32140 = n19046 | n25725 ;
  assign n32141 = n28109 | n32140 ;
  assign n32142 = n30612 ^ n30611 ^ n21586 ;
  assign n32143 = n26821 ^ n21192 ^ 1'b0 ;
  assign n32144 = ~n708 & n2864 ;
  assign n32145 = n6063 & ~n8542 ;
  assign n32146 = ~n9783 & n32145 ;
  assign n32147 = n19983 ^ n7599 ^ 1'b0 ;
  assign n32148 = n2656 & n32147 ;
  assign n32149 = n31565 ^ n9511 ^ 1'b0 ;
  assign n32150 = n19034 & n20799 ;
  assign n32151 = n3284 | n7448 ;
  assign n32152 = n29339 & ~n32151 ;
  assign n32153 = n9559 | n11951 ;
  assign n32154 = ( ~n2103 & n7719 ) | ( ~n2103 & n17855 ) | ( n7719 & n17855 ) ;
  assign n32155 = ( n6318 & n6794 ) | ( n6318 & n20184 ) | ( n6794 & n20184 ) ;
  assign n32156 = x1 | n7014 ;
  assign n32157 = n11038 & ~n11850 ;
  assign n32158 = n16987 & n32157 ;
  assign n32159 = n16213 ^ n2796 ^ 1'b0 ;
  assign n32160 = n7730 | n32159 ;
  assign n32161 = n1769 ^ n659 ^ 1'b0 ;
  assign n32162 = n16171 & n27820 ;
  assign n32167 = n3331 & n15633 ;
  assign n32168 = ( ~x1 & n15111 ) | ( ~x1 & n32167 ) | ( n15111 & n32167 ) ;
  assign n32169 = ~n19607 & n32168 ;
  assign n32163 = n4464 | n12368 ;
  assign n32164 = n3785 & ~n32163 ;
  assign n32165 = ~n8098 & n32164 ;
  assign n32166 = n15446 | n32165 ;
  assign n32170 = n32169 ^ n32166 ^ 1'b0 ;
  assign n32171 = ( n4002 & n5168 ) | ( n4002 & n7713 ) | ( n5168 & n7713 ) ;
  assign n32172 = n14848 ^ n13375 ^ 1'b0 ;
  assign n32173 = ~n7209 & n32172 ;
  assign n32174 = n32173 ^ n12559 ^ 1'b0 ;
  assign n32175 = n32171 & ~n32174 ;
  assign n32176 = n23291 ^ n16534 ^ 1'b0 ;
  assign n32177 = n32176 ^ n22783 ^ 1'b0 ;
  assign n32178 = n5799 & ~n14616 ;
  assign n32179 = n6621 & ~n12353 ;
  assign n32180 = n13594 & n32179 ;
  assign n32181 = n6551 | n32180 ;
  assign n32182 = n3798 & ~n6833 ;
  assign n32183 = n4335 & n32182 ;
  assign n32184 = ~n14582 & n17387 ;
  assign n32185 = n5480 ^ n165 ^ 1'b0 ;
  assign n32186 = n32185 ^ n1469 ^ 1'b0 ;
  assign n32187 = n17488 | n28170 ;
  assign n32188 = ~n5768 & n8917 ;
  assign n32189 = n19330 ^ n19189 ^ 1'b0 ;
  assign n32190 = ~n22898 & n32189 ;
  assign n32191 = n21666 ^ n7399 ^ 1'b0 ;
  assign n32192 = n5444 & n32191 ;
  assign n32193 = n32192 ^ n25144 ^ 1'b0 ;
  assign n32194 = n4298 & n11107 ;
  assign n32195 = n9688 | n18041 ;
  assign n32197 = n9153 ^ n6274 ^ 1'b0 ;
  assign n32196 = ~n5710 & n6296 ;
  assign n32198 = n32197 ^ n32196 ^ 1'b0 ;
  assign n32199 = n1329 & n32198 ;
  assign n32200 = n32199 ^ n24611 ^ 1'b0 ;
  assign n32201 = n1073 | n4794 ;
  assign n32202 = n15684 & ~n32201 ;
  assign n32203 = n29296 ^ n3405 ^ 1'b0 ;
  assign n32204 = n32202 & ~n32203 ;
  assign n32205 = ( n10027 & n11468 ) | ( n10027 & ~n15417 ) | ( n11468 & ~n15417 ) ;
  assign n32206 = n32205 ^ n4328 ^ 1'b0 ;
  assign n32207 = n12373 & n32206 ;
  assign n32208 = n77 | n11561 ;
  assign n32209 = n32208 ^ n189 ^ 1'b0 ;
  assign n32210 = n13883 & ~n32209 ;
  assign n32211 = n15174 ^ n6825 ^ 1'b0 ;
  assign n32212 = n16162 & ~n32211 ;
  assign n32213 = n32212 ^ n9731 ^ n7233 ;
  assign n32214 = n32210 | n32213 ;
  assign n32215 = n16251 ^ n10039 ^ 1'b0 ;
  assign n32216 = ~n7150 & n32215 ;
  assign n32217 = n26671 ^ n1878 ^ 1'b0 ;
  assign n32218 = n2671 & n32217 ;
  assign n32219 = ~n32216 & n32218 ;
  assign n32220 = ( n1501 & ~n2618 ) | ( n1501 & n20785 ) | ( ~n2618 & n20785 ) ;
  assign n32221 = n32220 ^ n8347 ^ 1'b0 ;
  assign n32222 = n28652 | n32221 ;
  assign n32223 = ( n19052 & n32219 ) | ( n19052 & n32222 ) | ( n32219 & n32222 ) ;
  assign n32224 = n32223 ^ n22915 ^ 1'b0 ;
  assign n32225 = ~n753 & n4369 ;
  assign n32226 = n32225 ^ n1510 ^ 1'b0 ;
  assign n32227 = n10322 | n32226 ;
  assign n32228 = n7052 ^ n335 ^ 1'b0 ;
  assign n32229 = n15757 | n32228 ;
  assign n32230 = n32229 ^ n25855 ^ 1'b0 ;
  assign n32231 = n32227 & ~n32230 ;
  assign n32232 = n13628 ^ n10603 ^ 1'b0 ;
  assign n32233 = ~n10173 & n32232 ;
  assign n32234 = n436 & n4579 ;
  assign n32235 = ~n4579 & n32234 ;
  assign n32236 = n79 & ~n857 ;
  assign n32237 = n857 & n32236 ;
  assign n32238 = ~n9363 & n21963 ;
  assign n32239 = n32237 & n32238 ;
  assign n32240 = n32239 ^ n26987 ^ 1'b0 ;
  assign n32241 = n32235 | n32240 ;
  assign n32242 = n32235 & ~n32241 ;
  assign n32243 = n16721 ^ n5684 ^ 1'b0 ;
  assign n32244 = n30782 ^ n25960 ^ n13462 ;
  assign n32245 = n12002 ^ n1202 ^ 1'b0 ;
  assign n32246 = ~n1016 & n14509 ;
  assign n32247 = n11817 & ~n20176 ;
  assign n32248 = n32246 & n32247 ;
  assign n32249 = n21948 ^ n4940 ^ 1'b0 ;
  assign n32250 = n2556 | n26670 ;
  assign n32251 = n1767 & n4960 ;
  assign n32252 = ~n28357 & n32251 ;
  assign n32253 = n25782 & ~n32252 ;
  assign n32254 = n32250 & n32253 ;
  assign n32255 = n2100 | n21302 ;
  assign n32256 = n8969 | n32255 ;
  assign n32257 = n32256 ^ n18583 ^ 1'b0 ;
  assign n32260 = n2926 & n11406 ;
  assign n32258 = n4693 | n8156 ;
  assign n32259 = n10443 & ~n32258 ;
  assign n32261 = n32260 ^ n32259 ^ 1'b0 ;
  assign n32262 = n2738 & n7659 ;
  assign n32263 = n6559 ^ n1551 ^ 1'b0 ;
  assign n32264 = ~n32262 & n32263 ;
  assign n32265 = n32264 ^ n25669 ^ 1'b0 ;
  assign n32266 = ~n7965 & n32265 ;
  assign n32268 = ~n15205 & n24280 ;
  assign n32267 = n9451 & ~n14772 ;
  assign n32269 = n32268 ^ n32267 ^ 1'b0 ;
  assign n32270 = n4037 & ~n21038 ;
  assign n32273 = n9962 ^ n2350 ^ 1'b0 ;
  assign n32271 = ~n3111 & n20169 ;
  assign n32272 = n32271 ^ n11285 ^ 1'b0 ;
  assign n32274 = n32273 ^ n32272 ^ 1'b0 ;
  assign n32275 = n12750 ^ n1267 ^ 1'b0 ;
  assign n32276 = ~n6817 & n32275 ;
  assign n32277 = n32276 ^ n27485 ^ n1868 ;
  assign n32278 = n5262 & n30169 ;
  assign n32279 = ~n32277 & n32278 ;
  assign n32280 = n22581 & ~n28692 ;
  assign n32281 = n32280 ^ n28509 ^ 1'b0 ;
  assign n32282 = n13096 & n14208 ;
  assign n32283 = n23099 & n32282 ;
  assign n32284 = n4264 & n24473 ;
  assign n32285 = n23880 | n32284 ;
  assign n32286 = n5510 & ~n32285 ;
  assign n32287 = n32286 ^ n16407 ^ 1'b0 ;
  assign n32288 = ( n1327 & ~n19893 ) | ( n1327 & n28118 ) | ( ~n19893 & n28118 ) ;
  assign n32289 = n22479 ^ n5001 ^ 1'b0 ;
  assign n32290 = n18817 & n32289 ;
  assign n32291 = ~n10171 & n14086 ;
  assign n32292 = ~n12338 & n32291 ;
  assign n32293 = n1937 & ~n16854 ;
  assign n32294 = n32293 ^ n1707 ^ 1'b0 ;
  assign n32295 = n14356 | n32294 ;
  assign n32296 = n30603 | n32295 ;
  assign n32297 = ~n9667 & n23352 ;
  assign n32298 = n8275 & n14925 ;
  assign n32299 = n6408 & n32298 ;
  assign n32300 = n2885 & ~n12303 ;
  assign n32301 = n32300 ^ n6999 ^ 1'b0 ;
  assign n32302 = n15712 ^ n6757 ^ 1'b0 ;
  assign n32304 = n22325 ^ n16021 ^ n15444 ;
  assign n32303 = ~n5064 & n9437 ;
  assign n32305 = n32304 ^ n32303 ^ 1'b0 ;
  assign n32306 = n10319 ^ n798 ^ 1'b0 ;
  assign n32307 = n9051 & ~n27332 ;
  assign n32308 = n1680 | n11630 ;
  assign n32309 = n32308 ^ n165 ^ 1'b0 ;
  assign n32310 = n9808 ^ n8152 ^ 1'b0 ;
  assign n32311 = n13954 & ~n32310 ;
  assign n32312 = n32309 & ~n32311 ;
  assign n32313 = n978 | n27756 ;
  assign n32314 = n32313 ^ n835 ^ 1'b0 ;
  assign n32315 = n17052 | n32314 ;
  assign n32316 = n19530 & n29332 ;
  assign n32317 = n11822 | n14697 ;
  assign n32318 = n32317 ^ n27797 ^ 1'b0 ;
  assign n32319 = n16716 ^ n5268 ^ 1'b0 ;
  assign n32320 = n2469 | n32319 ;
  assign n32321 = ~n1466 & n4432 ;
  assign n32322 = n32321 ^ n12502 ^ 1'b0 ;
  assign n32323 = n27586 ^ n26045 ^ n2747 ;
  assign n32324 = n32323 ^ n4641 ^ 1'b0 ;
  assign n32325 = n32322 & ~n32324 ;
  assign n32326 = ( n7086 & ~n9271 ) | ( n7086 & n15113 ) | ( ~n9271 & n15113 ) ;
  assign n32327 = n1758 | n32326 ;
  assign n32328 = ~n4240 & n6210 ;
  assign n32329 = n798 ^ n699 ^ 1'b0 ;
  assign n32330 = ~n19382 & n32329 ;
  assign n32333 = n23512 & ~n31059 ;
  assign n32331 = n19248 ^ n11300 ^ 1'b0 ;
  assign n32332 = n6581 | n32331 ;
  assign n32334 = n32333 ^ n32332 ^ 1'b0 ;
  assign n32335 = n32334 ^ n29251 ^ 1'b0 ;
  assign n32336 = n32330 & n32335 ;
  assign n32337 = n7297 & ~n13809 ;
  assign n32338 = n7889 & n32337 ;
  assign n32339 = ~n17320 & n32338 ;
  assign n32340 = ~n6348 & n9046 ;
  assign n32341 = n12860 ^ n2161 ^ 1'b0 ;
  assign n32342 = n6176 | n32341 ;
  assign n32343 = n2604 & ~n18441 ;
  assign n32345 = n508 | n18961 ;
  assign n32346 = n5769 | n32345 ;
  assign n32344 = n2634 | n3375 ;
  assign n32347 = n32346 ^ n32344 ^ 1'b0 ;
  assign n32348 = n17827 | n25477 ;
  assign n32349 = n18213 & ~n23558 ;
  assign n32350 = n18799 & n32349 ;
  assign n32351 = n492 & n4873 ;
  assign n32352 = n2170 & n32351 ;
  assign n32353 = n32352 ^ n493 ^ 1'b0 ;
  assign n32354 = n12816 & ~n32353 ;
  assign n32355 = n812 & n22044 ;
  assign n32356 = n19902 | n23171 ;
  assign n32357 = n8809 | n32356 ;
  assign n32358 = n32357 ^ n9534 ^ n1176 ;
  assign n32359 = n20533 | n21800 ;
  assign n32360 = n18199 & n32359 ;
  assign n32361 = ( n29485 & ~n32358 ) | ( n29485 & n32360 ) | ( ~n32358 & n32360 ) ;
  assign n32362 = n19534 ^ n11905 ^ 1'b0 ;
  assign n32363 = n17798 | n32362 ;
  assign n32364 = n6370 & ~n32363 ;
  assign n32365 = n32364 ^ n21769 ^ 1'b0 ;
  assign n32367 = n6299 ^ n3932 ^ 1'b0 ;
  assign n32368 = ~n10852 & n32367 ;
  assign n32369 = ~n3058 & n32368 ;
  assign n32366 = n12828 & n20475 ;
  assign n32370 = n32369 ^ n32366 ^ 1'b0 ;
  assign n32371 = ( n782 & n15292 ) | ( n782 & ~n27411 ) | ( n15292 & ~n27411 ) ;
  assign n32372 = ~n22308 & n24029 ;
  assign n32373 = ~n854 & n32372 ;
  assign n32375 = n29305 ^ n10753 ^ 1'b0 ;
  assign n32374 = ~n18458 & n19084 ;
  assign n32376 = n32375 ^ n32374 ^ 1'b0 ;
  assign n32377 = ~n291 & n32376 ;
  assign n32378 = n15618 | n20048 ;
  assign n32379 = n6278 & ~n15324 ;
  assign n32380 = ~n3891 & n32379 ;
  assign n32381 = n32380 ^ n10240 ^ 1'b0 ;
  assign n32382 = n9192 & ~n32381 ;
  assign n32383 = n32382 ^ n6797 ^ 1'b0 ;
  assign n32384 = n13942 & ~n32383 ;
  assign n32385 = n32384 ^ n25760 ^ 1'b0 ;
  assign n32386 = n3045 ^ n1530 ^ 1'b0 ;
  assign n32387 = n4021 & n11918 ;
  assign n32388 = n12701 ^ x6 ^ 1'b0 ;
  assign n32389 = ~n3939 & n9860 ;
  assign n32390 = n14795 & n32389 ;
  assign n32391 = n9098 | n11872 ;
  assign n32392 = n1627 & ~n27550 ;
  assign n32393 = n16033 & n23134 ;
  assign n32394 = n32393 ^ n24839 ^ 1'b0 ;
  assign n32395 = n18034 ^ n15750 ^ n7299 ;
  assign n32396 = ( ~n15413 & n32198 ) | ( ~n15413 & n32395 ) | ( n32198 & n32395 ) ;
  assign n32397 = n162 | n27213 ;
  assign n32398 = n21195 & n26808 ;
  assign n32399 = n15516 ^ n1955 ^ 1'b0 ;
  assign n32400 = n32261 ^ n1442 ^ 1'b0 ;
  assign n32401 = n31571 ^ n19087 ^ n2118 ;
  assign n32402 = n4835 & n8325 ;
  assign n32403 = n32402 ^ n7951 ^ n7324 ;
  assign n32404 = ( n5594 & n29927 ) | ( n5594 & ~n32403 ) | ( n29927 & ~n32403 ) ;
  assign n32405 = n29365 ^ n9037 ^ 1'b0 ;
  assign n32406 = n8975 | n32405 ;
  assign n32407 = n8591 & n17919 ;
  assign n32408 = n25571 ^ n20870 ^ 1'b0 ;
  assign n32409 = n24620 ^ n13413 ^ 1'b0 ;
  assign n32412 = n17151 ^ n2253 ^ 1'b0 ;
  assign n32410 = n1050 & n18111 ;
  assign n32411 = n8130 & ~n32410 ;
  assign n32413 = n32412 ^ n32411 ^ 1'b0 ;
  assign n32414 = ~n11870 & n24049 ;
  assign n32415 = n27331 & ~n32414 ;
  assign n32416 = ~n8710 & n9271 ;
  assign n32417 = n32416 ^ n16938 ^ n1791 ;
  assign n32418 = n7699 | n13557 ;
  assign n32419 = n32418 ^ n806 ^ 1'b0 ;
  assign n32420 = n22940 & ~n32419 ;
  assign n32421 = n12047 & ~n23558 ;
  assign n32422 = n4009 ^ n946 ^ 1'b0 ;
  assign n32423 = n26243 & ~n32422 ;
  assign n32424 = n13520 ^ n5552 ^ 1'b0 ;
  assign n32425 = n20662 | n32424 ;
  assign n32426 = n28706 | n32425 ;
  assign n32427 = n13675 ^ n404 ^ 1'b0 ;
  assign n32428 = n15400 ^ n12503 ^ 1'b0 ;
  assign n32429 = n839 & n25387 ;
  assign n32430 = ~n32428 & n32429 ;
  assign n32431 = n10828 ^ n1369 ^ 1'b0 ;
  assign n32432 = n14806 & ~n23636 ;
  assign n32442 = n149 | n5923 ;
  assign n32443 = n5923 & ~n32442 ;
  assign n32444 = n32443 ^ n13108 ^ 1'b0 ;
  assign n32437 = ~n150 & n1806 ;
  assign n32438 = n150 & n32437 ;
  assign n32439 = ~n1594 & n1863 ;
  assign n32440 = n32438 & n32439 ;
  assign n32441 = n548 & n32440 ;
  assign n32445 = n32444 ^ n32441 ^ 1'b0 ;
  assign n32446 = ~n2177 & n32445 ;
  assign n32433 = n3952 & ~n4976 ;
  assign n32434 = n4976 & n32433 ;
  assign n32435 = ~n659 & n32434 ;
  assign n32436 = ~n24996 & n32435 ;
  assign n32447 = n32446 ^ n32436 ^ 1'b0 ;
  assign n32448 = n16957 ^ n12690 ^ 1'b0 ;
  assign n32449 = n4113 & ~n23233 ;
  assign n32450 = n7299 | n7884 ;
  assign n32451 = n32449 | n32450 ;
  assign n32452 = n1767 & n32451 ;
  assign n32453 = n31091 ^ n22793 ^ 1'b0 ;
  assign n32454 = n6750 ^ n5880 ^ 1'b0 ;
  assign n32455 = n32454 ^ n15451 ^ 1'b0 ;
  assign n32456 = ~n7075 & n32455 ;
  assign n32457 = n7300 & ~n14356 ;
  assign n32458 = n32457 ^ n9701 ^ 1'b0 ;
  assign n32459 = n15953 ^ n7806 ^ 1'b0 ;
  assign n32460 = ~n32458 & n32459 ;
  assign n32461 = ~n7159 & n23875 ;
  assign n32462 = n13168 ^ n10904 ^ 1'b0 ;
  assign n32463 = ~n7149 & n32462 ;
  assign n32464 = n23481 ^ n7093 ^ 1'b0 ;
  assign n32465 = n5391 ^ n4019 ^ 1'b0 ;
  assign n32466 = n32465 ^ n20065 ^ 1'b0 ;
  assign n32467 = n6676 ^ n904 ^ 1'b0 ;
  assign n32468 = ~n32466 & n32467 ;
  assign n32469 = n7241 & ~n7685 ;
  assign n32470 = n24911 | n32469 ;
  assign n32471 = n32470 ^ n21323 ^ 1'b0 ;
  assign n32472 = n24697 ^ n813 ^ 1'b0 ;
  assign n32473 = n10434 ^ n8432 ^ 1'b0 ;
  assign n32474 = n7478 & n32473 ;
  assign n32475 = n32474 ^ n681 ^ 1'b0 ;
  assign n32476 = n7806 & ~n10259 ;
  assign n32477 = n205 & n32476 ;
  assign n32479 = n12514 ^ n4738 ^ 1'b0 ;
  assign n32480 = n15805 | n32479 ;
  assign n32478 = n5482 & ~n32391 ;
  assign n32481 = n32480 ^ n32478 ^ 1'b0 ;
  assign n32482 = n14542 | n30872 ;
  assign n32483 = n717 & ~n10194 ;
  assign n32484 = n3437 & n15515 ;
  assign n32485 = ~n9611 & n32484 ;
  assign n32486 = n6394 & n22704 ;
  assign n32488 = n4590 & ~n11778 ;
  assign n32487 = n11030 & ~n28112 ;
  assign n32489 = n32488 ^ n32487 ^ 1'b0 ;
  assign n32490 = n1212 ^ n253 ^ 1'b0 ;
  assign n32491 = n2389 & ~n21534 ;
  assign n32492 = n357 & n32491 ;
  assign n32493 = n9332 ^ n2179 ^ n1103 ;
  assign n32494 = n32493 ^ n30028 ^ 1'b0 ;
  assign n32497 = n2905 & n4208 ;
  assign n32498 = n32497 ^ n3602 ^ 1'b0 ;
  assign n32495 = n5982 ^ n2893 ^ 1'b0 ;
  assign n32496 = n24919 | n32495 ;
  assign n32499 = n32498 ^ n32496 ^ 1'b0 ;
  assign n32502 = n30345 ^ n4260 ^ 1'b0 ;
  assign n32503 = ( n800 & n23601 ) | ( n800 & n32502 ) | ( n23601 & n32502 ) ;
  assign n32504 = n31028 ^ n1533 ^ 1'b0 ;
  assign n32505 = n32503 & ~n32504 ;
  assign n32500 = n21883 ^ n4914 ^ 1'b0 ;
  assign n32501 = n17439 & n32500 ;
  assign n32506 = n32505 ^ n32501 ^ 1'b0 ;
  assign n32507 = n30766 ^ n23065 ^ 1'b0 ;
  assign n32508 = n23612 ^ n12854 ^ 1'b0 ;
  assign n32509 = n13436 | n17610 ;
  assign n32510 = n32509 ^ n8906 ^ 1'b0 ;
  assign n32511 = n32510 ^ n3292 ^ 1'b0 ;
  assign n32512 = n7403 & ~n32511 ;
  assign n32513 = n29502 ^ n28006 ^ 1'b0 ;
  assign n32514 = n10269 & ~n32513 ;
  assign n32515 = n32512 & n32514 ;
  assign n32516 = n32515 ^ n30777 ^ 1'b0 ;
  assign n32517 = n23112 ^ n14790 ^ 1'b0 ;
  assign n32518 = n32516 & n32517 ;
  assign n32519 = n8106 ^ n1617 ^ 1'b0 ;
  assign n32521 = ~n3745 & n9825 ;
  assign n32520 = n4104 & n9733 ;
  assign n32522 = n32521 ^ n32520 ^ 1'b0 ;
  assign n32523 = n3955 & ~n22675 ;
  assign n32524 = n32523 ^ n31361 ^ 1'b0 ;
  assign n32525 = n4189 & n4773 ;
  assign n32526 = n6256 | n32525 ;
  assign n32527 = n20199 & ~n28714 ;
  assign n32528 = n14868 | n32180 ;
  assign n32529 = n2883 & n3150 ;
  assign n32530 = ~n21714 & n21865 ;
  assign n32531 = ~n32529 & n32530 ;
  assign n32532 = n14885 ^ n10675 ^ 1'b0 ;
  assign n32533 = n5372 | n16361 ;
  assign n32534 = ~n6442 & n8541 ;
  assign n32535 = n27234 ^ n6121 ^ 1'b0 ;
  assign n32536 = n19704 ^ n4114 ^ 1'b0 ;
  assign n32537 = n27668 & n32536 ;
  assign n32538 = n14827 ^ n1392 ^ 1'b0 ;
  assign n32539 = n2438 | n32538 ;
  assign n32540 = ~n2146 & n26665 ;
  assign n32541 = n24637 | n32540 ;
  assign n32542 = n27173 & ~n32541 ;
  assign n32543 = n32539 | n32542 ;
  assign n32544 = n32537 | n32543 ;
  assign n32545 = n3017 & ~n30492 ;
  assign n32546 = n32545 ^ n29107 ^ 1'b0 ;
  assign n32548 = n4034 & n8177 ;
  assign n32549 = n32548 ^ n4229 ^ 1'b0 ;
  assign n32547 = n47 | n14371 ;
  assign n32550 = n32549 ^ n32547 ^ 1'b0 ;
  assign n32551 = n7765 | n32550 ;
  assign n32552 = n7996 | n16872 ;
  assign n32553 = n32551 & ~n32552 ;
  assign n32554 = n21287 ^ n4754 ^ 1'b0 ;
  assign n32555 = ( n2240 & n20105 ) | ( n2240 & n32173 ) | ( n20105 & n32173 ) ;
  assign n32556 = n9411 | n32555 ;
  assign n32557 = n25321 | n32556 ;
  assign n32558 = ~n15415 & n20075 ;
  assign n32559 = ~n12474 & n32558 ;
  assign n32560 = n27904 ^ n2661 ^ 1'b0 ;
  assign n32561 = n21807 & n32560 ;
  assign n32562 = n10903 & ~n22567 ;
  assign n32563 = n28816 ^ n10812 ^ 1'b0 ;
  assign n32564 = ~n3044 & n32563 ;
  assign n32565 = ~n7400 & n26298 ;
  assign n32566 = n31105 ^ n27323 ^ 1'b0 ;
  assign n32568 = n14248 ^ n3011 ^ 1'b0 ;
  assign n32567 = n20191 ^ n19235 ^ 1'b0 ;
  assign n32569 = n32568 ^ n32567 ^ 1'b0 ;
  assign n32570 = n32566 & ~n32569 ;
  assign n32571 = n2358 & n18416 ;
  assign n32572 = n32571 ^ n27583 ^ 1'b0 ;
  assign n32573 = n21670 ^ n1443 ^ 1'b0 ;
  assign n32574 = n25685 & ~n32573 ;
  assign n32575 = ~n6052 & n32574 ;
  assign n32576 = n4142 & n8130 ;
  assign n32577 = n12271 & n12584 ;
  assign n32578 = n32577 ^ n24797 ^ 1'b0 ;
  assign n32579 = n32578 ^ n13200 ^ 1'b0 ;
  assign n32580 = n1403 | n19737 ;
  assign n32581 = ~n8321 & n23075 ;
  assign n32582 = n110 & ~n5810 ;
  assign n32583 = n17605 & n19347 ;
  assign n32584 = n32582 & n32583 ;
  assign n32585 = n456 ^ n132 ^ 1'b0 ;
  assign n32586 = n1035 & n32585 ;
  assign n32587 = n25641 | n32586 ;
  assign n32588 = n32587 ^ n30192 ^ n15451 ;
  assign n32589 = n16263 ^ n10941 ^ 1'b0 ;
  assign n32590 = n30428 & ~n32589 ;
  assign n32591 = ~n32588 & n32590 ;
  assign n32593 = n6641 ^ n5724 ^ 1'b0 ;
  assign n32594 = ~n6004 & n32593 ;
  assign n32592 = n26973 ^ n2860 ^ 1'b0 ;
  assign n32595 = n32594 ^ n32592 ^ 1'b0 ;
  assign n32596 = n12651 ^ n10749 ^ 1'b0 ;
  assign n32597 = n3628 & n32596 ;
  assign n32598 = n24380 | n32597 ;
  assign n32599 = n5464 | n15678 ;
  assign n32600 = n32599 ^ n12260 ^ 1'b0 ;
  assign n32601 = n22538 | n32600 ;
  assign n32602 = n25849 ^ n14866 ^ n10092 ;
  assign n32603 = ~n1060 & n2784 ;
  assign n32604 = n32603 ^ n10481 ^ 1'b0 ;
  assign n32605 = n15956 & n32604 ;
  assign n32606 = n11070 & n32605 ;
  assign n32607 = n3744 & n8743 ;
  assign n32608 = n4463 | n5495 ;
  assign n32609 = ~n7800 & n13513 ;
  assign n32610 = n4075 ^ n1395 ^ 1'b0 ;
  assign n32611 = n32609 & n32610 ;
  assign n32612 = n32611 ^ n2784 ^ 1'b0 ;
  assign n32613 = n31113 ^ n7623 ^ 1'b0 ;
  assign n32614 = n16912 ^ n12154 ^ 1'b0 ;
  assign n32615 = n12902 & n32614 ;
  assign n32616 = ~n2515 & n3319 ;
  assign n32617 = n3761 | n6629 ;
  assign n32618 = n5235 | n32617 ;
  assign n32619 = n11670 ^ n11605 ^ 1'b0 ;
  assign n32620 = n32618 & n32619 ;
  assign n32621 = n30727 ^ n23683 ^ n3472 ;
  assign n32622 = n29255 ^ n28 ^ 1'b0 ;
  assign n32623 = n1284 & n11546 ;
  assign n32624 = n27670 & n32623 ;
  assign n32625 = n18582 & ~n32624 ;
  assign n32629 = n8058 & n25495 ;
  assign n32626 = n20522 ^ n5166 ^ 1'b0 ;
  assign n32627 = ~n1456 & n32626 ;
  assign n32628 = ~n3425 & n32627 ;
  assign n32630 = n32629 ^ n32628 ^ 1'b0 ;
  assign n32631 = n7893 | n8110 ;
  assign n32632 = n32631 ^ n9519 ^ 1'b0 ;
  assign n32633 = n20662 ^ n3315 ^ 1'b0 ;
  assign n32634 = ~n5704 & n32633 ;
  assign n32635 = ~n1363 & n8080 ;
  assign n32636 = n32635 ^ n12451 ^ n6573 ;
  assign n32637 = n261 | n4322 ;
  assign n32638 = n32637 ^ n30320 ^ 1'b0 ;
  assign n32639 = n5104 & ~n7162 ;
  assign n32640 = n10614 | n32639 ;
  assign n32641 = ( n4207 & n7344 ) | ( n4207 & ~n8095 ) | ( n7344 & ~n8095 ) ;
  assign n32642 = ~n16947 & n19151 ;
  assign n32643 = ( ~n24068 & n32641 ) | ( ~n24068 & n32642 ) | ( n32641 & n32642 ) ;
  assign n32644 = n183 & n26129 ;
  assign n32645 = ~n18460 & n19432 ;
  assign n32646 = n18327 & ~n21857 ;
  assign n32647 = n9630 ^ n5468 ^ 1'b0 ;
  assign n32648 = n8147 & ~n32647 ;
  assign n32649 = n12934 & n32648 ;
  assign n32650 = n32649 ^ n9639 ^ 1'b0 ;
  assign n32651 = n356 | n14108 ;
  assign n32652 = n32651 ^ n860 ^ 1'b0 ;
  assign n32653 = ~n3768 & n32652 ;
  assign n32654 = n7139 & n32408 ;
  assign n32655 = n10823 & ~n25117 ;
  assign n32656 = n32655 ^ n17729 ^ 1'b0 ;
  assign n32657 = n24804 & n32656 ;
  assign n32658 = n12673 ^ n4010 ^ 1'b0 ;
  assign n32659 = ~n16683 & n32658 ;
  assign n32660 = n30217 & n32659 ;
  assign n32661 = n32660 ^ n12744 ^ 1'b0 ;
  assign n32662 = n5524 & ~n31182 ;
  assign n32665 = n11717 & ~n24938 ;
  assign n32663 = n4952 & n14164 ;
  assign n32664 = n5179 & n32663 ;
  assign n32666 = n32665 ^ n32664 ^ 1'b0 ;
  assign n32667 = ~n2637 & n7352 ;
  assign n32668 = n10832 | n19774 ;
  assign n32669 = n32667 | n32668 ;
  assign n32670 = ( n390 & n21843 ) | ( n390 & ~n32669 ) | ( n21843 & ~n32669 ) ;
  assign n32671 = ~n11122 & n25581 ;
  assign n32672 = n32671 ^ n10364 ^ 1'b0 ;
  assign n32673 = n5809 | n32672 ;
  assign n32674 = n32673 ^ n24827 ^ 1'b0 ;
  assign n32675 = n31105 ^ n7488 ^ n1057 ;
  assign n32676 = n17051 | n32675 ;
  assign n32677 = n129 & n26852 ;
  assign n32678 = n32677 ^ n17677 ^ 1'b0 ;
  assign n32679 = n7873 & n32678 ;
  assign n32687 = n669 & ~n2483 ;
  assign n32688 = ~n669 & n32687 ;
  assign n32682 = n539 | n3389 ;
  assign n32683 = n539 & ~n32682 ;
  assign n32684 = n226 & n32683 ;
  assign n32685 = n117 | n32684 ;
  assign n32686 = n16340 & ~n32685 ;
  assign n32680 = n14551 & ~n19096 ;
  assign n32681 = n6299 & n32680 ;
  assign n32689 = n32688 ^ n32686 ^ n32681 ;
  assign n32690 = n7316 & n26660 ;
  assign n32691 = n9324 | n16486 ;
  assign n32692 = n32691 ^ n12294 ^ n6447 ;
  assign n32693 = n4432 & ~n5706 ;
  assign n32694 = ~n5897 & n32693 ;
  assign n32695 = n32694 ^ n2319 ^ 1'b0 ;
  assign n32696 = n3521 & ~n21003 ;
  assign n32697 = n6528 & n10933 ;
  assign n32698 = n2478 | n32697 ;
  assign n32699 = n667 ^ n631 ^ 1'b0 ;
  assign n32700 = n27668 & n32699 ;
  assign n32701 = n15896 & ~n23654 ;
  assign n32702 = n6245 ^ n5323 ^ 1'b0 ;
  assign n32703 = n2006 | n11552 ;
  assign n32704 = n9609 & ~n32703 ;
  assign n32705 = n30679 | n32704 ;
  assign n32706 = n11920 & ~n14636 ;
  assign n32707 = n224 & n32706 ;
  assign n32708 = n21857 ^ n1392 ^ 1'b0 ;
  assign n32709 = ~n32707 & n32708 ;
  assign n32710 = n32709 ^ n7798 ^ n6756 ;
  assign n32711 = n11377 & n22601 ;
  assign n32712 = n5933 & n28490 ;
  assign n32713 = n32712 ^ n11238 ^ 1'b0 ;
  assign n32714 = n6976 ^ n466 ^ 1'b0 ;
  assign n32715 = n642 & ~n8071 ;
  assign n32716 = n14544 ^ n9754 ^ 1'b0 ;
  assign n32717 = ~n13893 & n32716 ;
  assign n32718 = n21666 ^ n890 ^ 1'b0 ;
  assign n32719 = n32717 & ~n32718 ;
  assign n32720 = n1219 & n5945 ;
  assign n32721 = n12091 & n32720 ;
  assign n32722 = n875 & n7493 ;
  assign n32723 = ( ~n9386 & n25719 ) | ( ~n9386 & n32722 ) | ( n25719 & n32722 ) ;
  assign n32724 = n14724 | n32723 ;
  assign n32725 = n175 & ~n32724 ;
  assign n32726 = n11673 ^ n2190 ^ 1'b0 ;
  assign n32727 = n32726 ^ n6236 ^ 1'b0 ;
  assign n32728 = n11147 | n32727 ;
  assign n32729 = ~n302 & n1980 ;
  assign n32730 = n32729 ^ n8338 ^ 1'b0 ;
  assign n32731 = n10454 & ~n32730 ;
  assign n32732 = ~n19659 & n32731 ;
  assign n32733 = n32732 ^ n9145 ^ n3599 ;
  assign n32734 = n25330 | n32733 ;
  assign n32735 = n14247 ^ n738 ^ 1'b0 ;
  assign n32736 = ~n16925 & n32735 ;
  assign n32737 = n13695 & n14292 ;
  assign n32738 = n7984 ^ n7707 ^ 1'b0 ;
  assign n32739 = n29423 ^ n9913 ^ 1'b0 ;
  assign n32740 = n26750 & n32739 ;
  assign n32741 = n28710 ^ n12985 ^ n1256 ;
  assign n32742 = n15241 & ~n32741 ;
  assign n32743 = ( n7153 & n7403 ) | ( n7153 & ~n18647 ) | ( n7403 & ~n18647 ) ;
  assign n32744 = n12043 & ~n32743 ;
  assign n32745 = n21960 & n32744 ;
  assign n32746 = n6265 | n27343 ;
  assign n32747 = n8412 & ~n10354 ;
  assign n32748 = n32747 ^ n841 ^ 1'b0 ;
  assign n32749 = ( n16106 & ~n30368 ) | ( n16106 & n32748 ) | ( ~n30368 & n32748 ) ;
  assign n32750 = n13412 ^ n10098 ^ 1'b0 ;
  assign n32751 = n32750 ^ n29689 ^ n3095 ;
  assign n32752 = n20281 ^ n11383 ^ 1'b0 ;
  assign n32753 = n4245 & n32752 ;
  assign n32754 = n32753 ^ n23367 ^ 1'b0 ;
  assign n32755 = n12661 & n14667 ;
  assign n32756 = n12551 & n32755 ;
  assign n32757 = ~n2398 & n32756 ;
  assign n32758 = n9653 | n28771 ;
  assign n32759 = ~n21326 & n29382 ;
  assign n32760 = n32759 ^ n8176 ^ 1'b0 ;
  assign n32761 = n2108 & n5118 ;
  assign n32762 = n32761 ^ n1267 ^ 1'b0 ;
  assign n32763 = ~n12214 & n32762 ;
  assign n32764 = n13883 | n14390 ;
  assign n32765 = n2262 ^ n614 ^ 1'b0 ;
  assign n32766 = n20815 | n32765 ;
  assign n32767 = ~n20759 & n30220 ;
  assign n32771 = n4377 & n9121 ;
  assign n32768 = n13870 ^ n8321 ^ 1'b0 ;
  assign n32769 = n15506 & n32768 ;
  assign n32770 = n26101 & n32769 ;
  assign n32772 = n32771 ^ n32770 ^ 1'b0 ;
  assign n32773 = ~n1361 & n17746 ;
  assign n32776 = n3600 & ~n19918 ;
  assign n32777 = n32776 ^ n28893 ^ 1'b0 ;
  assign n32774 = n27278 ^ n22748 ^ 1'b0 ;
  assign n32775 = n28315 & n32774 ;
  assign n32778 = n32777 ^ n32775 ^ 1'b0 ;
  assign n32779 = ~n7289 & n10479 ;
  assign n32783 = n9760 & n22044 ;
  assign n32784 = ~n5071 & n32783 ;
  assign n32780 = n1217 & n4572 ;
  assign n32781 = ~n2498 & n32780 ;
  assign n32782 = ~n5165 & n32781 ;
  assign n32785 = n32784 ^ n32782 ^ 1'b0 ;
  assign n32786 = ~n21371 & n25530 ;
  assign n32787 = n1329 | n26508 ;
  assign n32788 = n32787 ^ n7107 ^ 1'b0 ;
  assign n32789 = n1701 & ~n12996 ;
  assign n32790 = n32789 ^ n22039 ^ 1'b0 ;
  assign n32791 = n7145 | n15198 ;
  assign n32792 = ~n4864 & n5664 ;
  assign n32793 = n14969 | n28590 ;
  assign n32794 = n20281 | n31968 ;
  assign n32795 = n32793 | n32794 ;
  assign n32796 = ~n9689 & n15004 ;
  assign n32797 = n15748 & ~n28812 ;
  assign n32798 = n32797 ^ n8244 ^ 1'b0 ;
  assign n32799 = ~n2753 & n5253 ;
  assign n32800 = ~n934 & n32799 ;
  assign n32801 = n5439 & n32800 ;
  assign n32802 = n32801 ^ n20423 ^ 1'b0 ;
  assign n32803 = n32798 & ~n32802 ;
  assign n32804 = n9491 ^ n2349 ^ 1'b0 ;
  assign n32805 = n9403 & n32804 ;
  assign n32806 = n7322 & n32805 ;
  assign n32807 = n32806 ^ n21782 ^ 1'b0 ;
  assign n32808 = n3632 & n26448 ;
  assign n32809 = ~n32807 & n32808 ;
  assign n32810 = n22871 ^ n521 ^ 1'b0 ;
  assign n32811 = n24028 ^ n4271 ^ 1'b0 ;
  assign n32812 = n32811 ^ n20 ^ 1'b0 ;
  assign n32813 = n32810 & n32812 ;
  assign n32814 = n15590 ^ n4762 ^ 1'b0 ;
  assign n32815 = n661 & ~n32814 ;
  assign n32816 = ~n32813 & n32815 ;
  assign n32817 = ( ~n1381 & n8101 ) | ( ~n1381 & n32816 ) | ( n8101 & n32816 ) ;
  assign n32818 = n1179 & n13900 ;
  assign n32819 = ~n1246 & n32818 ;
  assign n32820 = n13543 ^ n9180 ^ 1'b0 ;
  assign n32821 = n11848 & n32820 ;
  assign n32822 = ~n30353 & n32821 ;
  assign n32823 = n2953 | n15559 ;
  assign n32824 = ~n6311 & n25316 ;
  assign n32825 = ~n27980 & n32824 ;
  assign n32826 = n30134 ^ n27418 ^ 1'b0 ;
  assign n32827 = ~n8198 & n24885 ;
  assign n32828 = ~n4914 & n26770 ;
  assign n32829 = n7534 | n19226 ;
  assign n32830 = n25272 | n32829 ;
  assign n32831 = n2465 & n2954 ;
  assign n32832 = ( n729 & n32830 ) | ( n729 & ~n32831 ) | ( n32830 & ~n32831 ) ;
  assign n32833 = n24769 & n24832 ;
  assign n32834 = n26000 ^ n16847 ^ 1'b0 ;
  assign n32835 = ~n21509 & n32834 ;
  assign n32836 = n6100 ^ n2906 ^ 1'b0 ;
  assign n32837 = n9941 & n32836 ;
  assign n32838 = n32837 ^ n8525 ^ 1'b0 ;
  assign n32839 = n6149 ^ n1488 ^ 1'b0 ;
  assign n32840 = n14388 | n32839 ;
  assign n32841 = n32840 ^ n16415 ^ 1'b0 ;
  assign n32842 = n6290 & n32841 ;
  assign n32843 = n12489 & ~n13342 ;
  assign n32844 = n32843 ^ n26352 ^ 1'b0 ;
  assign n32845 = n16367 ^ n16270 ^ 1'b0 ;
  assign n32846 = n30026 & ~n32589 ;
  assign n32847 = n788 | n5249 ;
  assign n32848 = ~n8487 & n32847 ;
  assign n32849 = n453 | n32848 ;
  assign n32851 = ( n434 & n2238 ) | ( n434 & ~n10345 ) | ( n2238 & ~n10345 ) ;
  assign n32850 = n17183 | n29649 ;
  assign n32852 = n32851 ^ n32850 ^ 1'b0 ;
  assign n32853 = n32849 & n32852 ;
  assign n32854 = n32853 ^ n26099 ^ 1'b0 ;
  assign n32855 = n12122 ^ n1955 ^ n749 ;
  assign n32856 = n6116 | n32855 ;
  assign n32857 = n978 & ~n32856 ;
  assign n32858 = n32857 ^ n15390 ^ 1'b0 ;
  assign n32859 = n19821 ^ n7798 ^ 1'b0 ;
  assign n32860 = n20816 & ~n32859 ;
  assign n32861 = ( x1 & n25504 ) | ( x1 & ~n32860 ) | ( n25504 & ~n32860 ) ;
  assign n32862 = n6568 & ~n16470 ;
  assign n32863 = n32862 ^ n2283 ^ 1'b0 ;
  assign n32864 = ~n290 & n17130 ;
  assign n32865 = n401 & ~n32864 ;
  assign n32866 = n1434 & n32865 ;
  assign n32867 = ~n2852 & n7056 ;
  assign n32868 = ~n12899 & n32867 ;
  assign n32869 = n19611 | n32868 ;
  assign n32870 = n23861 ^ n22121 ^ 1'b0 ;
  assign n32871 = ~n20460 & n32870 ;
  assign n32872 = n1983 & n8084 ;
  assign n32873 = n28594 & n32872 ;
  assign n32874 = n11419 | n32873 ;
  assign n32875 = n23593 & ~n32874 ;
  assign n32876 = n8313 & ~n10485 ;
  assign n32877 = n32876 ^ n8972 ^ 1'b0 ;
  assign n32878 = ~n13737 & n19257 ;
  assign n32879 = ~n32877 & n32878 ;
  assign n32880 = n32879 ^ n6426 ^ 1'b0 ;
  assign n32881 = n32880 ^ n4070 ^ 1'b0 ;
  assign n32882 = n10452 | n32881 ;
  assign n32883 = n14997 ^ n1119 ^ 1'b0 ;
  assign n32884 = n32883 ^ n5379 ^ n2228 ;
  assign n32885 = n14249 ^ n668 ^ 1'b0 ;
  assign n32887 = n8867 ^ n86 ^ 1'b0 ;
  assign n32886 = n5183 | n15354 ;
  assign n32888 = n32887 ^ n32886 ^ 1'b0 ;
  assign n32889 = n1275 ^ n683 ^ 1'b0 ;
  assign n32890 = n32889 ^ n13322 ^ 1'b0 ;
  assign n32891 = ~n6588 & n32890 ;
  assign n32892 = n25964 & n32891 ;
  assign n32893 = n11951 & n32892 ;
  assign n32894 = n14285 & ~n18386 ;
  assign n32895 = n32893 & n32894 ;
  assign n32896 = n24114 ^ n9231 ^ 1'b0 ;
  assign n32897 = n3447 ^ n1052 ^ 1'b0 ;
  assign n32898 = n11103 | n32897 ;
  assign n32899 = n10188 | n11636 ;
  assign n32900 = n32899 ^ n7263 ^ 1'b0 ;
  assign n32901 = n32900 ^ n16604 ^ 1'b0 ;
  assign n32902 = n16463 & n32901 ;
  assign n32903 = n32902 ^ n2060 ^ 1'b0 ;
  assign n32904 = n31042 & n32903 ;
  assign n32905 = n32898 & n32904 ;
  assign n32907 = n19112 ^ n393 ^ 1'b0 ;
  assign n32908 = n32907 ^ n13283 ^ 1'b0 ;
  assign n32906 = n17822 ^ n12450 ^ 1'b0 ;
  assign n32909 = n32908 ^ n32906 ^ n4895 ;
  assign n32910 = n19485 ^ n11471 ^ n27 ;
  assign n32911 = ~n2217 & n12000 ;
  assign n32912 = n23953 ^ n1403 ^ 1'b0 ;
  assign n32913 = n228 | n32912 ;
  assign n32914 = n6043 | n32913 ;
  assign n32915 = n18808 & ~n23028 ;
  assign n32916 = n32915 ^ n15016 ^ 1'b0 ;
  assign n32917 = n6676 & n17542 ;
  assign n32918 = n32917 ^ n10497 ^ 1'b0 ;
  assign n32919 = ~n3324 & n5263 ;
  assign n32920 = ~n6605 & n12584 ;
  assign n32921 = n577 & n32920 ;
  assign n32922 = n32921 ^ n24955 ^ 1'b0 ;
  assign n32923 = ~n32919 & n32922 ;
  assign n32924 = ~n6989 & n18349 ;
  assign n32925 = n11551 & n32924 ;
  assign n32926 = n17417 | n32925 ;
  assign n32927 = n32926 ^ n13797 ^ 1'b0 ;
  assign n32928 = ~n2628 & n7237 ;
  assign n32929 = n11483 & ~n21788 ;
  assign n32930 = n9522 & ~n22386 ;
  assign n32931 = ~n13802 & n17945 ;
  assign n32932 = ~n8091 & n32931 ;
  assign n32934 = ~n2094 & n20672 ;
  assign n32935 = n26597 ^ n8223 ^ 1'b0 ;
  assign n32936 = n32934 & n32935 ;
  assign n32933 = ~n15898 & n21161 ;
  assign n32937 = n32936 ^ n32933 ^ 1'b0 ;
  assign n32938 = n28357 ^ n23318 ^ 1'b0 ;
  assign n32939 = n7298 & ~n19421 ;
  assign n32940 = n7832 & n32939 ;
  assign n32941 = ( n8494 & n18007 ) | ( n8494 & n32940 ) | ( n18007 & n32940 ) ;
  assign n32942 = n3918 | n32941 ;
  assign n32943 = n32942 ^ n29158 ^ n25592 ;
  assign n32945 = ~n162 & n10434 ;
  assign n32946 = n28018 & n32945 ;
  assign n32944 = n9624 & n25108 ;
  assign n32947 = n32946 ^ n32944 ^ 1'b0 ;
  assign n32948 = n15488 ^ n4962 ^ 1'b0 ;
  assign n32949 = n320 & ~n32948 ;
  assign n32950 = n14037 & ~n15650 ;
  assign n32951 = n25492 ^ n9864 ^ 1'b0 ;
  assign n32952 = n28511 & n32951 ;
  assign n32953 = n8505 | n17052 ;
  assign n32954 = n32953 ^ n30380 ^ 1'b0 ;
  assign n32955 = n10793 | n32954 ;
  assign n32956 = n32955 ^ n27829 ^ 1'b0 ;
  assign n32957 = n147 & ~n3698 ;
  assign n32958 = n11106 & n32957 ;
  assign n32959 = n32958 ^ n4061 ^ 1'b0 ;
  assign n32960 = n18981 | n32959 ;
  assign n32961 = n32960 ^ n18033 ^ 1'b0 ;
  assign n32962 = n22646 & ~n32961 ;
  assign n32963 = ( n1246 & n5606 ) | ( n1246 & ~n22473 ) | ( n5606 & ~n22473 ) ;
  assign n32964 = n16000 ^ n14249 ^ 1'b0 ;
  assign n32965 = n23197 & n32964 ;
  assign n32966 = n28762 ^ n13758 ^ 1'b0 ;
  assign n32967 = n8510 & ~n32966 ;
  assign n32968 = ~n1054 & n8305 ;
  assign n32969 = n32968 ^ n7110 ^ 1'b0 ;
  assign n32970 = n19664 | n32969 ;
  assign n32971 = n32970 ^ n14541 ^ 1'b0 ;
  assign n32972 = ~n8156 & n32971 ;
  assign n32973 = n32972 ^ n22126 ^ 1'b0 ;
  assign n32974 = n18424 ^ n16225 ^ 1'b0 ;
  assign n32975 = n19206 | n32974 ;
  assign n32976 = n32975 ^ n28547 ^ 1'b0 ;
  assign n32977 = ~n12004 & n13840 ;
  assign n32978 = ~n2610 & n24030 ;
  assign n32979 = n800 & n3599 ;
  assign n32980 = n32979 ^ n27862 ^ 1'b0 ;
  assign n32981 = n10837 & ~n13002 ;
  assign n32982 = ~n485 & n567 ;
  assign n32983 = n3023 & ~n11238 ;
  assign n32984 = n32983 ^ n22059 ^ 1'b0 ;
  assign n32985 = n7447 & ~n14539 ;
  assign n32986 = n32984 & n32985 ;
  assign n32987 = n10836 & n14345 ;
  assign n32990 = n16931 ^ n7717 ^ n892 ;
  assign n32989 = n18027 | n28958 ;
  assign n32991 = n32990 ^ n32989 ^ 1'b0 ;
  assign n32992 = n13110 | n32991 ;
  assign n32988 = n11428 & ~n30091 ;
  assign n32993 = n32992 ^ n32988 ^ 1'b0 ;
  assign n32994 = n20101 ^ n18919 ^ 1'b0 ;
  assign n32995 = n1413 & n32994 ;
  assign n32996 = n32995 ^ n21800 ^ 1'b0 ;
  assign n32997 = n32079 & ~n32996 ;
  assign n33004 = ( ~n2802 & n5267 ) | ( ~n2802 & n22020 ) | ( n5267 & n22020 ) ;
  assign n32998 = n1002 & n4768 ;
  assign n32999 = ~n1002 & n32998 ;
  assign n33000 = n6570 & ~n32999 ;
  assign n33001 = n32999 & n33000 ;
  assign n33002 = n24485 & ~n33001 ;
  assign n33003 = n16044 & n33002 ;
  assign n33005 = n33004 ^ n33003 ^ 1'b0 ;
  assign n33006 = n4340 & ~n17571 ;
  assign n33007 = n33006 ^ n5591 ^ 1'b0 ;
  assign n33010 = n17221 ^ n5866 ^ 1'b0 ;
  assign n33008 = ~n10610 & n13776 ;
  assign n33009 = n33008 ^ n6991 ^ 1'b0 ;
  assign n33011 = n33010 ^ n33009 ^ 1'b0 ;
  assign n33012 = n7600 & ~n29347 ;
  assign n33013 = n2313 & n8721 ;
  assign n33014 = n3330 & n17549 ;
  assign n33015 = n9012 & n33014 ;
  assign n33016 = n2118 ^ n85 ^ 1'b0 ;
  assign n33017 = n33016 ^ n23949 ^ 1'b0 ;
  assign n33018 = n23355 | n33017 ;
  assign n33019 = n22600 ^ n20881 ^ 1'b0 ;
  assign n33020 = n33019 ^ n29914 ^ 1'b0 ;
  assign n33021 = n16411 & ~n33020 ;
  assign n33022 = ~n3045 & n6842 ;
  assign n33023 = n33022 ^ n17221 ^ 1'b0 ;
  assign n33024 = n15388 ^ n10180 ^ 1'b0 ;
  assign n33025 = n31123 ^ n4668 ^ 1'b0 ;
  assign n33026 = ( n1810 & n33024 ) | ( n1810 & n33025 ) | ( n33024 & n33025 ) ;
  assign n33027 = ~n16442 & n24084 ;
  assign n33028 = n19767 ^ n9351 ^ 1'b0 ;
  assign n33029 = ( n1986 & n5340 ) | ( n1986 & n25521 ) | ( n5340 & n25521 ) ;
  assign n33030 = n33029 ^ n6874 ^ n3428 ;
  assign n33031 = n33030 ^ n16540 ^ 1'b0 ;
  assign n33032 = n30028 & ~n33031 ;
  assign n33033 = n4024 & ~n23922 ;
  assign n33034 = n33033 ^ n11757 ^ 1'b0 ;
  assign n33035 = n18602 | n33034 ;
  assign n33036 = n33035 ^ n5151 ^ 1'b0 ;
  assign n33037 = n7907 ^ n291 ^ 1'b0 ;
  assign n33038 = n33037 ^ n15207 ^ 1'b0 ;
  assign n33039 = n536 & n21619 ;
  assign n33040 = n30483 ^ n10154 ^ 1'b0 ;
  assign n33041 = n3118 & n18375 ;
  assign n33042 = n33041 ^ n4009 ^ 1'b0 ;
  assign n33043 = n30285 & n33042 ;
  assign n33044 = n2796 | n11861 ;
  assign n33045 = n33044 ^ n3308 ^ 1'b0 ;
  assign n33046 = n26379 | n33045 ;
  assign n33047 = n32165 ^ n15060 ^ 1'b0 ;
  assign n33048 = ~n12057 & n26189 ;
  assign n33049 = ( n5320 & n11704 ) | ( n5320 & ~n23456 ) | ( n11704 & ~n23456 ) ;
  assign n33050 = n3415 & ~n22386 ;
  assign n33051 = ~n2346 & n33050 ;
  assign n33052 = n29918 ^ n12651 ^ 1'b0 ;
  assign n33053 = n21383 & ~n33052 ;
  assign n33054 = n33051 & n33053 ;
  assign n33055 = n5274 & ~n19064 ;
  assign n33056 = ( n13909 & n23377 ) | ( n13909 & ~n33055 ) | ( n23377 & ~n33055 ) ;
  assign n33057 = n32483 ^ n23580 ^ 1'b0 ;
  assign n33058 = ~n33056 & n33057 ;
  assign n33059 = n15390 ^ n7924 ^ 1'b0 ;
  assign n33060 = ( n4977 & n11013 ) | ( n4977 & ~n11425 ) | ( n11013 & ~n11425 ) ;
  assign n33061 = ( n3042 & n9134 ) | ( n3042 & n12995 ) | ( n9134 & n12995 ) ;
  assign n33062 = n7109 ^ n403 ^ 1'b0 ;
  assign n33063 = n23207 & n33062 ;
  assign n33064 = ~n11798 & n33063 ;
  assign n33065 = n13605 | n32667 ;
  assign n33066 = ~n15 & n33065 ;
  assign n33067 = n33066 ^ n14520 ^ 1'b0 ;
  assign n33068 = n11273 ^ n7471 ^ 1'b0 ;
  assign n33069 = n33068 ^ n11151 ^ 1'b0 ;
  assign n33070 = n27115 ^ n20113 ^ 1'b0 ;
  assign n33071 = n6671 | n33070 ;
  assign n33072 = ( ~n6271 & n8787 ) | ( ~n6271 & n33071 ) | ( n8787 & n33071 ) ;
  assign n33077 = n3851 & n21240 ;
  assign n33074 = n18474 & ~n29514 ;
  assign n33075 = ~n96 & n33074 ;
  assign n33073 = n1542 & ~n14081 ;
  assign n33076 = n33075 ^ n33073 ^ n8805 ;
  assign n33078 = n33077 ^ n33076 ^ 1'b0 ;
  assign n33079 = n14360 & ~n33078 ;
  assign n33080 = n20820 ^ n17424 ^ 1'b0 ;
  assign n33081 = n167 & ~n33080 ;
  assign n33082 = ~n20484 & n33081 ;
  assign n33083 = ~n6714 & n33082 ;
  assign n33084 = n6441 | n9279 ;
  assign n33085 = n33084 ^ n10409 ^ 1'b0 ;
  assign n33086 = ~n5374 & n33085 ;
  assign n33087 = ~n6133 & n33086 ;
  assign n33088 = n33087 ^ n5088 ^ 1'b0 ;
  assign n33089 = n23022 | n33088 ;
  assign n33090 = n19235 ^ n3056 ^ 1'b0 ;
  assign n33094 = n65 | n25251 ;
  assign n33095 = n33094 ^ n21490 ^ 1'b0 ;
  assign n33091 = n9781 & ~n32666 ;
  assign n33092 = n33091 ^ n28207 ^ 1'b0 ;
  assign n33093 = ~n21071 & n33092 ;
  assign n33096 = n33095 ^ n33093 ^ 1'b0 ;
  assign n33097 = ~n14331 & n14997 ;
  assign n33098 = n9694 & ~n25251 ;
  assign n33099 = n33098 ^ n14911 ^ 1'b0 ;
  assign n33100 = n20207 ^ n12941 ^ 1'b0 ;
  assign n33101 = ~n33099 & n33100 ;
  assign n33102 = n16768 & n33101 ;
  assign n33103 = n18183 & n33102 ;
  assign n33104 = n33103 ^ n12831 ^ n404 ;
  assign n33105 = n2784 & n14142 ;
  assign n33106 = ~n11784 & n33105 ;
  assign n33107 = n1395 | n33106 ;
  assign n33109 = n4567 ^ n1251 ^ 1'b0 ;
  assign n33110 = ~n31442 & n33109 ;
  assign n33108 = n12301 | n23351 ;
  assign n33111 = n33110 ^ n33108 ^ 1'b0 ;
  assign n33112 = n1907 | n25468 ;
  assign n33113 = n28710 & ~n33112 ;
  assign n33114 = ~n6394 & n18889 ;
  assign n33115 = n25903 & n33114 ;
  assign n33116 = n33115 ^ n6082 ^ 1'b0 ;
  assign n33117 = ~n33113 & n33116 ;
  assign n33118 = n1975 | n25196 ;
  assign n33122 = n21417 ^ n7046 ^ 1'b0 ;
  assign n33119 = n31613 ^ n13266 ^ 1'b0 ;
  assign n33120 = n1980 & ~n33119 ;
  assign n33121 = n13366 & n33120 ;
  assign n33123 = n33122 ^ n33121 ^ 1'b0 ;
  assign n33124 = n14750 & n15863 ;
  assign n33125 = n16473 & n33124 ;
  assign n33126 = n33125 ^ n13258 ^ n7048 ;
  assign n33127 = ( n104 & n2648 ) | ( n104 & ~n3726 ) | ( n2648 & ~n3726 ) ;
  assign n33128 = n3715 & n15782 ;
  assign n33129 = n15516 & n33128 ;
  assign n33130 = n33129 ^ n31674 ^ 1'b0 ;
  assign n33131 = n33127 & ~n33130 ;
  assign n33132 = ~n14078 & n33131 ;
  assign n33133 = n18128 & n33132 ;
  assign n33134 = ( n205 & n2138 ) | ( n205 & ~n2462 ) | ( n2138 & ~n2462 ) ;
  assign n33135 = ~n14873 & n33134 ;
  assign n33136 = n33135 ^ n9726 ^ 1'b0 ;
  assign n33137 = n8573 & ~n22322 ;
  assign n33138 = n12024 ^ n8233 ^ 1'b0 ;
  assign n33139 = n9701 & ~n23287 ;
  assign n33140 = n33139 ^ n698 ^ 1'b0 ;
  assign n33141 = n33140 ^ n4486 ^ 1'b0 ;
  assign n33142 = n12781 ^ n445 ^ 1'b0 ;
  assign n33143 = n20962 & n33142 ;
  assign n33144 = n31819 & n33143 ;
  assign n33145 = n20137 ^ n1289 ^ 1'b0 ;
  assign n33146 = n1628 & n33145 ;
  assign n33147 = n3227 & n18411 ;
  assign n33148 = n29032 ^ n10603 ^ 1'b0 ;
  assign n33149 = n10501 & n23810 ;
  assign n33150 = n33149 ^ n4037 ^ 1'b0 ;
  assign n33151 = n727 | n32552 ;
  assign n33152 = n33151 ^ n729 ^ 1'b0 ;
  assign n33153 = n15775 & ~n33152 ;
  assign n33154 = n11445 & n28590 ;
  assign n33155 = n33153 & n33154 ;
  assign n33156 = n19293 | n26322 ;
  assign n33157 = n29817 ^ n24926 ^ 1'b0 ;
  assign n33158 = n8907 & n33157 ;
  assign n33159 = ~n26897 & n30513 ;
  assign n33160 = n18134 & ~n18952 ;
  assign n33161 = n33160 ^ n18821 ^ 1'b0 ;
  assign n33162 = ( n4263 & ~n6353 ) | ( n4263 & n8867 ) | ( ~n6353 & n8867 ) ;
  assign n33163 = ( n1159 & n16573 ) | ( n1159 & ~n33162 ) | ( n16573 & ~n33162 ) ;
  assign n33164 = n18648 ^ n16885 ^ 1'b0 ;
  assign n33165 = n33164 ^ n17087 ^ 1'b0 ;
  assign n33166 = n1014 & ~n22886 ;
  assign n33168 = n2127 & ~n22939 ;
  assign n33167 = ~n1932 & n4569 ;
  assign n33169 = n33168 ^ n33167 ^ n9391 ;
  assign n33170 = ~n33166 & n33169 ;
  assign n33171 = ~n6052 & n33170 ;
  assign n33172 = n33171 ^ n6041 ^ 1'b0 ;
  assign n33173 = n24297 ^ n4131 ^ 1'b0 ;
  assign n33174 = n10300 & ~n33173 ;
  assign n33175 = n19004 ^ n2129 ^ 1'b0 ;
  assign n33176 = ~n3724 & n7132 ;
  assign n33177 = ( n1835 & n31392 ) | ( n1835 & n32893 ) | ( n31392 & n32893 ) ;
  assign n33178 = n634 | n17493 ;
  assign n33179 = n33178 ^ n27294 ^ 1'b0 ;
  assign n33180 = n7916 & n29757 ;
  assign n33181 = n33180 ^ n13438 ^ 1'b0 ;
  assign n33182 = n22438 ^ n16565 ^ 1'b0 ;
  assign n33183 = n12375 & n33182 ;
  assign n33184 = n7793 & n33183 ;
  assign n33185 = n33184 ^ n17735 ^ 1'b0 ;
  assign n33186 = n15602 ^ n14586 ^ 1'b0 ;
  assign n33187 = n11189 ^ n10544 ^ 1'b0 ;
  assign n33188 = n33187 ^ n23749 ^ 1'b0 ;
  assign n33189 = ~n12053 & n25110 ;
  assign n33190 = n33189 ^ n24540 ^ 1'b0 ;
  assign n33191 = n33190 ^ n6969 ^ 1'b0 ;
  assign n33192 = n9222 | n33191 ;
  assign n33193 = ( n21772 & ~n33188 ) | ( n21772 & n33192 ) | ( ~n33188 & n33192 ) ;
  assign n33194 = n15089 & ~n19754 ;
  assign n33195 = n33194 ^ n8427 ^ 1'b0 ;
  assign n33196 = n6447 & n21090 ;
  assign n33197 = ~n14125 & n33196 ;
  assign n33198 = n33197 ^ n2129 ^ 1'b0 ;
  assign n33199 = n2835 & ~n31360 ;
  assign n33200 = n33199 ^ n16087 ^ 1'b0 ;
  assign n33201 = n30272 ^ n26869 ^ 1'b0 ;
  assign n33205 = n5915 ^ n822 ^ 1'b0 ;
  assign n33206 = n33205 ^ n8054 ^ 1'b0 ;
  assign n33202 = ~n4064 & n9532 ;
  assign n33203 = ~n12580 & n33202 ;
  assign n33204 = n33203 ^ n1964 ^ 1'b0 ;
  assign n33207 = n33206 ^ n33204 ^ 1'b0 ;
  assign n33208 = n8989 ^ n7014 ^ 1'b0 ;
  assign n33209 = n17640 | n33208 ;
  assign n33210 = n5634 & ~n19283 ;
  assign n33211 = n11371 ^ n10147 ^ 1'b0 ;
  assign n33212 = n6591 & ~n33211 ;
  assign n33213 = ( n2902 & n4335 ) | ( n2902 & n10465 ) | ( n4335 & n10465 ) ;
  assign n33214 = n33213 ^ n16523 ^ 1'b0 ;
  assign n33215 = n33212 & n33214 ;
  assign n33216 = n7124 ^ n4409 ^ 1'b0 ;
  assign n33217 = ~n1072 & n9518 ;
  assign n33218 = n33217 ^ n6535 ^ 1'b0 ;
  assign n33221 = ~n4675 & n17108 ;
  assign n33222 = n10070 | n33221 ;
  assign n33219 = ( n2584 & n4800 ) | ( n2584 & n5864 ) | ( n4800 & n5864 ) ;
  assign n33220 = n33219 ^ n10277 ^ 1'b0 ;
  assign n33223 = n33222 ^ n33220 ^ n26364 ;
  assign n33224 = n13311 & n25653 ;
  assign n33225 = n33224 ^ n9074 ^ 1'b0 ;
  assign n33226 = n9621 ^ n3462 ^ 1'b0 ;
  assign n33227 = n25917 & n33226 ;
  assign n33228 = n7251 ^ n1723 ^ 1'b0 ;
  assign n33229 = n10059 ^ n6128 ^ 1'b0 ;
  assign n33230 = n20031 ^ n10120 ^ n4925 ;
  assign n33231 = n33230 ^ n15415 ^ n5859 ;
  assign n33232 = ~n8062 & n12371 ;
  assign n33233 = n33232 ^ n13495 ^ 1'b0 ;
  assign n33234 = n17810 | n27582 ;
  assign n33235 = n33234 ^ n16124 ^ 1'b0 ;
  assign n33236 = n22683 & ~n33235 ;
  assign n33237 = n6566 ^ n447 ^ 1'b0 ;
  assign n33238 = n11098 ^ n10245 ^ 1'b0 ;
  assign n33239 = ( ~n2721 & n7081 ) | ( ~n2721 & n7143 ) | ( n7081 & n7143 ) ;
  assign n33240 = n11811 & ~n33239 ;
  assign n33241 = ~n5181 & n33240 ;
  assign n33242 = ( n1789 & n16861 ) | ( n1789 & ~n25554 ) | ( n16861 & ~n25554 ) ;
  assign n33243 = n9358 | n27512 ;
  assign n33244 = n33243 ^ n33161 ^ 1'b0 ;
  assign n33245 = n9928 | n16532 ;
  assign n33246 = n8230 & ~n33245 ;
  assign n33247 = n8716 & n25941 ;
  assign n33248 = n33247 ^ n31042 ^ 1'b0 ;
  assign n33249 = n8204 ^ n2930 ^ 1'b0 ;
  assign n33250 = n25968 | n33249 ;
  assign n33251 = n12400 & ~n26292 ;
  assign n33252 = n16673 ^ n11209 ^ n1202 ;
  assign n33253 = n11198 | n33252 ;
  assign n33254 = n20608 ^ n19601 ^ 1'b0 ;
  assign n33255 = n21907 | n33254 ;
  assign n33256 = n10217 & ~n23372 ;
  assign n33257 = n8478 & n33256 ;
  assign n33258 = ~n30178 & n33257 ;
  assign n33259 = n33258 ^ n31422 ^ 1'b0 ;
  assign n33260 = n4573 ^ n2999 ^ 1'b0 ;
  assign n33261 = ( ~n5595 & n12893 ) | ( ~n5595 & n22065 ) | ( n12893 & n22065 ) ;
  assign n33262 = n1416 | n2431 ;
  assign n33263 = n7292 | n33262 ;
  assign n33264 = n27458 ^ n10049 ^ 1'b0 ;
  assign n33265 = n4596 & ~n5747 ;
  assign n33266 = n33265 ^ n8229 ^ n415 ;
  assign n33267 = n10366 | n33266 ;
  assign n33268 = n33267 ^ n33068 ^ 1'b0 ;
  assign n33269 = n5517 ^ n3370 ^ 1'b0 ;
  assign n33270 = n428 | n6885 ;
  assign n33271 = n33270 ^ n16483 ^ 1'b0 ;
  assign n33272 = n33269 & n33271 ;
  assign n33273 = n5814 & ~n27204 ;
  assign n33274 = n229 | n2264 ;
  assign n33275 = n33274 ^ n14962 ^ 1'b0 ;
  assign n33276 = n2066 & n33275 ;
  assign n33277 = n33276 ^ n3763 ^ 1'b0 ;
  assign n33278 = n23010 | n33277 ;
  assign n33279 = n33278 ^ n7935 ^ 1'b0 ;
  assign n33284 = n7749 ^ n1929 ^ 1'b0 ;
  assign n33285 = n11146 & ~n33284 ;
  assign n33282 = n2588 ^ n331 ^ 1'b0 ;
  assign n33280 = n10614 ^ n8291 ^ 1'b0 ;
  assign n33281 = n24749 & n33280 ;
  assign n33283 = n33282 ^ n33281 ^ 1'b0 ;
  assign n33286 = n33285 ^ n33283 ^ n9372 ;
  assign n33287 = n4974 & ~n7293 ;
  assign n33288 = n16268 & ~n18209 ;
  assign n33289 = n33287 & n33288 ;
  assign n33290 = n6368 & ~n33289 ;
  assign n33291 = n33290 ^ n4701 ^ 1'b0 ;
  assign n33292 = n11360 ^ n7027 ^ 1'b0 ;
  assign n33293 = n3732 & ~n33292 ;
  assign n33294 = n18542 & ~n33293 ;
  assign n33295 = ~n11872 & n25532 ;
  assign n33296 = n17291 & n24493 ;
  assign n33297 = ~n471 & n33296 ;
  assign n33298 = n431 | n5354 ;
  assign n33299 = n33298 ^ n20785 ^ 1'b0 ;
  assign n33300 = n33299 ^ n163 ^ 1'b0 ;
  assign n33304 = n11498 | n30443 ;
  assign n33305 = n33304 ^ n22603 ^ 1'b0 ;
  assign n33301 = n9770 & ~n19720 ;
  assign n33302 = n1944 & ~n33301 ;
  assign n33303 = ~n15703 & n33302 ;
  assign n33306 = n33305 ^ n33303 ^ 1'b0 ;
  assign n33307 = n33306 ^ n14878 ^ n12013 ;
  assign n33308 = n9795 ^ n1590 ^ 1'b0 ;
  assign n33309 = ~n10275 & n10598 ;
  assign n33310 = n1845 & n5549 ;
  assign n33311 = n33310 ^ n18885 ^ 1'b0 ;
  assign n33312 = n18177 & ~n33311 ;
  assign n33313 = n16671 ^ n11274 ^ 1'b0 ;
  assign n33314 = n4338 | n9260 ;
  assign n33315 = n1590 & ~n33314 ;
  assign n33316 = ~n482 & n10103 ;
  assign n33317 = n23727 ^ n703 ^ 1'b0 ;
  assign n33318 = ~n33316 & n33317 ;
  assign n33319 = n31743 ^ n1688 ^ 1'b0 ;
  assign n33320 = n466 & ~n33319 ;
  assign n33321 = n26243 & ~n31136 ;
  assign n33322 = n7744 ^ n5374 ^ 1'b0 ;
  assign n33323 = n21928 & ~n33322 ;
  assign n33324 = n33323 ^ n6643 ^ 1'b0 ;
  assign n33325 = n9074 & n11081 ;
  assign n33326 = n222 & n33325 ;
  assign n33327 = ( ~n3171 & n6129 ) | ( ~n3171 & n27822 ) | ( n6129 & n27822 ) ;
  assign n33328 = n18393 & ~n22373 ;
  assign n33329 = n12393 | n20648 ;
  assign n33330 = n33329 ^ n436 ^ 1'b0 ;
  assign n33331 = ~n6070 & n33330 ;
  assign n33332 = n3802 & ~n15229 ;
  assign n33333 = n33332 ^ n12005 ^ 1'b0 ;
  assign n33334 = n27836 & n31728 ;
  assign n33335 = n33334 ^ n25896 ^ 1'b0 ;
  assign n33336 = n12837 | n16544 ;
  assign n33337 = n4007 | n33336 ;
  assign n33338 = n3293 & n9923 ;
  assign n33339 = n33338 ^ n2496 ^ 1'b0 ;
  assign n33340 = n8606 ^ n7208 ^ 1'b0 ;
  assign n33341 = n4180 & ~n16463 ;
  assign n33342 = n4329 & ~n13031 ;
  assign n33343 = n33341 & n33342 ;
  assign n33344 = n8599 | n15743 ;
  assign n33345 = n33344 ^ n13298 ^ n7909 ;
  assign n33346 = n18137 & ~n25328 ;
  assign n33347 = n33346 ^ n5152 ^ 1'b0 ;
  assign n33348 = n3409 & n22373 ;
  assign n33349 = n19809 & n25590 ;
  assign n33350 = ( ~n10696 & n22580 ) | ( ~n10696 & n31206 ) | ( n22580 & n31206 ) ;
  assign n33351 = n7095 & ~n10084 ;
  assign n33352 = n33351 ^ n9756 ^ 1'b0 ;
  assign n33353 = n5461 & ~n33352 ;
  assign n33354 = n33350 & n33353 ;
  assign n33355 = n33354 ^ n4211 ^ 1'b0 ;
  assign n33356 = ~n2723 & n8898 ;
  assign n33357 = n11256 ^ n7657 ^ 1'b0 ;
  assign n33358 = ~n22925 & n33357 ;
  assign n33359 = n33358 ^ n2409 ^ 1'b0 ;
  assign n33360 = n4776 & ~n18777 ;
  assign n33361 = n25741 & ~n33360 ;
  assign n33363 = n7407 ^ n5200 ^ 1'b0 ;
  assign n33364 = ~n3250 & n33363 ;
  assign n33365 = n1453 & ~n33364 ;
  assign n33362 = ~n11431 & n12994 ;
  assign n33366 = n33365 ^ n33362 ^ 1'b0 ;
  assign n33367 = ~n11729 & n33366 ;
  assign n33368 = ~n20799 & n33367 ;
  assign n33369 = n19339 ^ n758 ^ 1'b0 ;
  assign n33370 = ~n991 & n33369 ;
  assign n33371 = n23619 ^ n6933 ^ 1'b0 ;
  assign n33372 = n130 | n3185 ;
  assign n33373 = n11274 & ~n16106 ;
  assign n33374 = n33373 ^ n8850 ^ 1'b0 ;
  assign n33375 = n4216 & n33374 ;
  assign n33376 = n29893 ^ n10031 ^ 1'b0 ;
  assign n33377 = n11009 & n33376 ;
  assign n33378 = n620 & n2151 ;
  assign n33379 = n1306 & ~n16509 ;
  assign n33380 = n2163 & n33379 ;
  assign n33381 = n29815 ^ n13913 ^ 1'b0 ;
  assign n33382 = n2185 & n15916 ;
  assign n33383 = ~n18628 & n33382 ;
  assign n33384 = n24401 ^ n4444 ^ 1'b0 ;
  assign n33385 = n2732 ^ n2640 ^ 1'b0 ;
  assign n33386 = n12480 & n33385 ;
  assign n33387 = n26707 ^ n16673 ^ n12557 ;
  assign n33388 = n6814 | n10752 ;
  assign n33389 = n3992 ^ n1695 ^ 1'b0 ;
  assign n33390 = n33389 ^ n8830 ^ 1'b0 ;
  assign n33391 = n33388 | n33390 ;
  assign n33392 = n20410 | n30340 ;
  assign n33393 = n5234 & n8166 ;
  assign n33394 = n32495 ^ n20039 ^ 1'b0 ;
  assign n33395 = n33393 | n33394 ;
  assign n33396 = n11205 & n12433 ;
  assign n33397 = n33396 ^ n18046 ^ 1'b0 ;
  assign n33398 = ~n2541 & n33397 ;
  assign n33399 = n33398 ^ n3510 ^ 1'b0 ;
  assign n33400 = n12057 & ~n33399 ;
  assign n33401 = n33400 ^ n9046 ^ n8206 ;
  assign n33402 = n33401 ^ n33075 ^ n4718 ;
  assign n33403 = n5216 & ~n10412 ;
  assign n33404 = n33403 ^ n208 ^ 1'b0 ;
  assign n33405 = n15719 & ~n33404 ;
  assign n33406 = n4773 & n8468 ;
  assign n33407 = ~n2366 & n33406 ;
  assign n33409 = n22571 ^ n9049 ^ 1'b0 ;
  assign n33408 = n667 & ~n9592 ;
  assign n33410 = n33409 ^ n33408 ^ 1'b0 ;
  assign n33411 = n5890 ^ n971 ^ 1'b0 ;
  assign n33412 = ~n3264 & n11048 ;
  assign n33413 = n16654 ^ n13171 ^ 1'b0 ;
  assign n33414 = n25495 | n33413 ;
  assign n33415 = n2724 & ~n33414 ;
  assign n33416 = n22615 & n33415 ;
  assign n33417 = n2971 | n10177 ;
  assign n33418 = n3349 | n12106 ;
  assign n33419 = n27200 | n33418 ;
  assign n33420 = n8410 & ~n24645 ;
  assign n33421 = ~n18421 & n33420 ;
  assign n33422 = n10553 ^ n4338 ^ 1'b0 ;
  assign n33423 = n6166 | n22870 ;
  assign n33424 = n33423 ^ n18295 ^ n12515 ;
  assign n33425 = n1742 & n3721 ;
  assign n33426 = ~n16337 & n33425 ;
  assign n33427 = ~n758 & n33426 ;
  assign n33428 = n14500 | n20395 ;
  assign n33429 = n33428 ^ n10699 ^ 1'b0 ;
  assign n33430 = ~n33427 & n33429 ;
  assign n33431 = n33430 ^ n395 ^ 1'b0 ;
  assign n33432 = n22000 ^ n9062 ^ 1'b0 ;
  assign n33433 = ~n14200 & n23810 ;
  assign n33434 = n33433 ^ n12422 ^ 1'b0 ;
  assign n33435 = n11162 & ~n33434 ;
  assign n33436 = n18664 ^ n8989 ^ 1'b0 ;
  assign n33437 = ~n229 & n9193 ;
  assign n33438 = n23969 & n33437 ;
  assign n33439 = n19188 | n26873 ;
  assign n33440 = n10305 ^ n1207 ^ 1'b0 ;
  assign n33441 = ~n3405 & n33440 ;
  assign n33442 = n3219 | n19647 ;
  assign n33443 = n3274 & ~n33442 ;
  assign n33444 = n26869 & n33443 ;
  assign n33445 = n4088 ^ n411 ^ 1'b0 ;
  assign n33446 = n2754 & ~n9724 ;
  assign n33447 = n33445 | n33446 ;
  assign n33448 = ~n6643 & n16725 ;
  assign n33449 = n33448 ^ n9084 ^ 1'b0 ;
  assign n33450 = n6523 & ~n11162 ;
  assign n33451 = ~n1372 & n32422 ;
  assign n33452 = ~n33145 & n33451 ;
  assign n33453 = n13364 & n27508 ;
  assign n33454 = n15394 & n33453 ;
  assign n33455 = ( n5151 & n7396 ) | ( n5151 & ~n18511 ) | ( n7396 & ~n18511 ) ;
  assign n33456 = n2885 & ~n23817 ;
  assign n33457 = n6754 & n33456 ;
  assign n33458 = n11240 ^ n4746 ^ n4095 ;
  assign n33459 = n6383 & n33458 ;
  assign n33460 = n2070 & n33459 ;
  assign n33461 = n3802 & ~n33460 ;
  assign n33462 = ~n33457 & n33461 ;
  assign n33463 = n894 & ~n6754 ;
  assign n33464 = n282 & ~n22110 ;
  assign n33465 = n3758 ^ n3131 ^ 1'b0 ;
  assign n33466 = ~n13665 & n14007 ;
  assign n33467 = n10895 & n33466 ;
  assign n33468 = ~n26360 & n26714 ;
  assign n33469 = n33468 ^ n10634 ^ 1'b0 ;
  assign n33470 = n16439 ^ n13832 ^ 1'b0 ;
  assign n33471 = n33470 ^ n2552 ^ 1'b0 ;
  assign n33472 = n9770 & ~n27430 ;
  assign n33473 = n98 | n33472 ;
  assign n33474 = n19926 & ~n33473 ;
  assign n33475 = n33474 ^ n2000 ^ 1'b0 ;
  assign n33476 = n32097 ^ n4588 ^ 1'b0 ;
  assign n33477 = n25924 ^ n17193 ^ 1'b0 ;
  assign n33478 = n22902 & ~n33477 ;
  assign n33479 = n32202 ^ n13012 ^ 1'b0 ;
  assign n33480 = n28490 ^ n10621 ^ 1'b0 ;
  assign n33481 = ~n25958 & n33480 ;
  assign n33482 = ( ~n1543 & n18867 ) | ( ~n1543 & n33481 ) | ( n18867 & n33481 ) ;
  assign n33483 = n6764 & ~n25287 ;
  assign n33484 = n16410 & n25447 ;
  assign n33485 = n33249 & n33484 ;
  assign n33486 = n4081 ^ n3909 ^ 1'b0 ;
  assign n33487 = n13002 & n33486 ;
  assign n33488 = n33485 & n33487 ;
  assign n33489 = ( n1269 & ~n5258 ) | ( n1269 & n16580 ) | ( ~n5258 & n16580 ) ;
  assign n33490 = n33489 ^ n15015 ^ 1'b0 ;
  assign n33491 = ~n30239 & n33490 ;
  assign n33492 = n3582 & n13150 ;
  assign n33493 = n33491 | n33492 ;
  assign n33494 = n1868 & ~n4449 ;
  assign n33495 = ~n1786 & n33090 ;
  assign n33496 = n33495 ^ n31335 ^ 1'b0 ;
  assign n33497 = n22914 ^ n8712 ^ n963 ;
  assign n33500 = n96 & ~n5686 ;
  assign n33501 = n819 & n6719 ;
  assign n33502 = ~n33500 & n33501 ;
  assign n33503 = n22857 & ~n33502 ;
  assign n33498 = ~n4372 & n7968 ;
  assign n33499 = ~n13750 & n33498 ;
  assign n33504 = n33503 ^ n33499 ^ 1'b0 ;
  assign n33505 = n996 | n2421 ;
  assign n33506 = n33505 ^ n11704 ^ 1'b0 ;
  assign n33507 = n13277 | n33506 ;
  assign n33508 = n33507 ^ n4539 ^ 1'b0 ;
  assign n33509 = n33508 ^ n459 ^ 1'b0 ;
  assign n33510 = n2415 | n8042 ;
  assign n33511 = n33510 ^ n205 ^ 1'b0 ;
  assign n33512 = ~n649 & n8834 ;
  assign n33513 = n16083 ^ n11285 ^ n5690 ;
  assign n33514 = n33513 ^ n28820 ^ 1'b0 ;
  assign n33515 = n13437 ^ n5540 ^ n826 ;
  assign n33516 = n33515 ^ n28454 ^ 1'b0 ;
  assign n33517 = n1544 & n15213 ;
  assign n33518 = n26225 ^ n17417 ^ 1'b0 ;
  assign n33519 = n18828 ^ n8421 ^ 1'b0 ;
  assign n33520 = n27810 | n33519 ;
  assign n33521 = n7233 & n11827 ;
  assign n33522 = n33521 ^ n15562 ^ 1'b0 ;
  assign n33523 = n11627 | n18347 ;
  assign n33524 = n2813 ^ n159 ^ 1'b0 ;
  assign n33525 = n191 | n414 ;
  assign n33526 = n33525 ^ n36 ^ 1'b0 ;
  assign n33527 = ~n33524 & n33526 ;
  assign n33528 = n33524 & n33527 ;
  assign n33529 = n15195 | n32800 ;
  assign n33530 = n33529 ^ n15796 ^ 1'b0 ;
  assign n33531 = ( n1473 & n7146 ) | ( n1473 & n20149 ) | ( n7146 & n20149 ) ;
  assign n33532 = n33029 ^ n30852 ^ 1'b0 ;
  assign n33533 = n30438 & n33532 ;
  assign n33534 = n24398 ^ n10500 ^ 1'b0 ;
  assign n33535 = n20641 & ~n33269 ;
  assign n33536 = n7404 | n8478 ;
  assign n33537 = n33536 ^ n16042 ^ 1'b0 ;
  assign n33538 = n6586 | n9858 ;
  assign n33539 = n33538 ^ n7187 ^ 1'b0 ;
  assign n33540 = n30447 ^ n22065 ^ n61 ;
  assign n33541 = n430 & n17620 ;
  assign n33542 = n33541 ^ n221 ^ 1'b0 ;
  assign n33543 = ~n863 & n2895 ;
  assign n33544 = n33543 ^ n1781 ^ 1'b0 ;
  assign n33545 = ~n33542 & n33544 ;
  assign n33546 = ( ~n3331 & n23583 ) | ( ~n3331 & n33545 ) | ( n23583 & n33545 ) ;
  assign n33547 = n24199 ^ n3453 ^ 1'b0 ;
  assign n33549 = n6878 ^ n3867 ^ 1'b0 ;
  assign n33550 = n3193 | n33549 ;
  assign n33548 = n4173 & n9860 ;
  assign n33551 = n33550 ^ n33548 ^ 1'b0 ;
  assign n33552 = n20414 ^ n4451 ^ 1'b0 ;
  assign n33553 = n4754 | n33552 ;
  assign n33554 = n9958 ^ n3082 ^ 1'b0 ;
  assign n33555 = n21533 & n33554 ;
  assign n33556 = n33555 ^ n30482 ^ 1'b0 ;
  assign n33557 = n17416 & n32645 ;
  assign n33558 = n33557 ^ n22347 ^ 1'b0 ;
  assign n33559 = n12449 ^ n4674 ^ 1'b0 ;
  assign n33560 = ~n1217 & n5602 ;
  assign n33561 = n2996 & ~n33560 ;
  assign n33562 = n3035 & ~n33561 ;
  assign n33563 = n2871 & n33562 ;
  assign n33564 = n21187 ^ n5880 ^ 1'b0 ;
  assign n33565 = ( n7529 & ~n8778 ) | ( n7529 & n13117 ) | ( ~n8778 & n13117 ) ;
  assign n33566 = ( n3158 & n6959 ) | ( n3158 & ~n33565 ) | ( n6959 & ~n33565 ) ;
  assign n33567 = n33566 ^ n10670 ^ 1'b0 ;
  assign n33568 = n33564 | n33567 ;
  assign n33569 = n11306 ^ n8542 ^ 1'b0 ;
  assign n33570 = n33568 | n33569 ;
  assign n33571 = n5320 ^ n4087 ^ n3980 ;
  assign n33572 = n1055 & ~n9205 ;
  assign n33573 = n33572 ^ n4774 ^ 1'b0 ;
  assign n33574 = n33571 | n33573 ;
  assign n33575 = n29314 ^ n22872 ^ 1'b0 ;
  assign n33576 = ~n3135 & n5863 ;
  assign n33577 = n33576 ^ n7514 ^ 1'b0 ;
  assign n33578 = n31168 | n33518 ;
  assign n33579 = n33577 & ~n33578 ;
  assign n33580 = n1256 & ~n30435 ;
  assign n33581 = ~n403 & n1437 ;
  assign n33582 = n21952 ^ n18849 ^ 1'b0 ;
  assign n33583 = ~n10437 & n33582 ;
  assign n33584 = n19911 | n32583 ;
  assign n33585 = n8447 | n18525 ;
  assign n33586 = n14601 & ~n33585 ;
  assign n33587 = n6243 & n21101 ;
  assign n33588 = n10305 & n33587 ;
  assign n33589 = n33588 ^ n20533 ^ 1'b0 ;
  assign n33590 = n1574 & ~n22646 ;
  assign n33591 = n33589 & ~n33590 ;
  assign n33592 = n11124 ^ n4021 ^ 1'b0 ;
  assign n33593 = n24084 ^ n16164 ^ 1'b0 ;
  assign n33594 = n33593 ^ n2955 ^ 1'b0 ;
  assign n33595 = n33592 | n33594 ;
  assign n33596 = n854 & n18983 ;
  assign n33597 = n19588 & n33596 ;
  assign n33598 = n12365 ^ n1769 ^ 1'b0 ;
  assign n33599 = n33597 & ~n33598 ;
  assign n33600 = n1539 ^ n459 ^ 1'b0 ;
  assign n33601 = n18453 & ~n22052 ;
  assign n33602 = n8076 | n33601 ;
  assign n33603 = n33602 ^ n6041 ^ 1'b0 ;
  assign n33604 = n14566 ^ n6039 ^ 1'b0 ;
  assign n33605 = n9178 & n18678 ;
  assign n33606 = n23696 ^ n654 ^ 1'b0 ;
  assign n33609 = ~n6308 & n24531 ;
  assign n33607 = n28058 ^ n18786 ^ 1'b0 ;
  assign n33608 = n1025 & n33607 ;
  assign n33610 = n33609 ^ n33608 ^ 1'b0 ;
  assign n33611 = ~n22689 & n33610 ;
  assign n33612 = n19473 ^ n9886 ^ 1'b0 ;
  assign n33613 = n63 & ~n1615 ;
  assign n33614 = n16079 | n28701 ;
  assign n33615 = ( ~n1365 & n33613 ) | ( ~n1365 & n33614 ) | ( n33613 & n33614 ) ;
  assign n33616 = ( n19186 & n33170 ) | ( n19186 & ~n33615 ) | ( n33170 & ~n33615 ) ;
  assign n33617 = n1329 ^ n823 ^ 1'b0 ;
  assign n33618 = ~n9621 & n33617 ;
  assign n33619 = n5195 & ~n14672 ;
  assign n33620 = n25924 ^ n10822 ^ 1'b0 ;
  assign n33621 = ~n14767 & n33620 ;
  assign n33622 = ~n16790 & n33621 ;
  assign n33623 = n33622 ^ n4610 ^ 1'b0 ;
  assign n33624 = n19891 | n31070 ;
  assign n33625 = n2132 & n32261 ;
  assign n33626 = ~n28363 & n33625 ;
  assign n33628 = n15514 ^ n3738 ^ 1'b0 ;
  assign n33629 = n9419 | n33628 ;
  assign n33630 = n7842 ^ n105 ^ 1'b0 ;
  assign n33631 = ~n6630 & n33630 ;
  assign n33632 = n33629 & n33631 ;
  assign n33627 = n849 & n4587 ;
  assign n33633 = n33632 ^ n33627 ^ 1'b0 ;
  assign n33634 = n28360 ^ n4278 ^ 1'b0 ;
  assign n33635 = n23325 & ~n24573 ;
  assign n33636 = n33635 ^ n10893 ^ 1'b0 ;
  assign n33637 = n12147 | n22847 ;
  assign n33638 = n14160 ^ n4741 ^ 1'b0 ;
  assign n33639 = n33638 ^ n29030 ^ 1'b0 ;
  assign n33640 = n27304 ^ n20562 ^ 1'b0 ;
  assign n33641 = ( n24108 & n32285 ) | ( n24108 & ~n33640 ) | ( n32285 & ~n33640 ) ;
  assign n33642 = n33641 ^ n1819 ^ 1'b0 ;
  assign n33643 = n31280 & n33642 ;
  assign n33644 = n1276 ^ n74 ^ 1'b0 ;
  assign n33645 = n24326 | n33644 ;
  assign n33646 = n33645 ^ n3992 ^ 1'b0 ;
  assign n33647 = n16281 & ~n27130 ;
  assign n33648 = n1898 & ~n12611 ;
  assign n33649 = n21718 ^ n13728 ^ n6998 ;
  assign n33650 = n20933 ^ n5522 ^ 1'b0 ;
  assign n33651 = n33650 ^ n411 ^ 1'b0 ;
  assign n33652 = ~n5604 & n15206 ;
  assign n33653 = n33652 ^ n32484 ^ n12983 ;
  assign n33654 = n30612 ^ n13046 ^ 1'b0 ;
  assign n33655 = n347 | n10361 ;
  assign n33656 = ( n4347 & ~n6111 ) | ( n4347 & n7515 ) | ( ~n6111 & n7515 ) ;
  assign n33657 = n33656 ^ n10855 ^ 1'b0 ;
  assign n33658 = ~n2539 & n9873 ;
  assign n33659 = n2660 & n4780 ;
  assign n33660 = ~n4780 & n33659 ;
  assign n33661 = n3255 | n15467 ;
  assign n33662 = ( ~n4058 & n33660 ) | ( ~n4058 & n33661 ) | ( n33660 & n33661 ) ;
  assign n33663 = ~n3649 & n7696 ;
  assign n33664 = n33663 ^ n6151 ^ 1'b0 ;
  assign n33665 = ( n4357 & ~n20772 ) | ( n4357 & n33664 ) | ( ~n20772 & n33664 ) ;
  assign n33666 = n5567 | n33665 ;
  assign n33671 = n23532 ^ n10085 ^ 1'b0 ;
  assign n33672 = n10740 & n33671 ;
  assign n33669 = n7261 | n9539 ;
  assign n33670 = n33669 ^ n28375 ^ 1'b0 ;
  assign n33667 = ~n7530 & n10049 ;
  assign n33668 = n33667 ^ n24092 ^ n5886 ;
  assign n33673 = n33672 ^ n33670 ^ n33668 ;
  assign n33674 = ~n2304 & n4021 ;
  assign n33675 = n33674 ^ n33220 ^ 1'b0 ;
  assign n33677 = ~n892 & n14558 ;
  assign n33676 = n14299 & n22443 ;
  assign n33678 = n33677 ^ n33676 ^ 1'b0 ;
  assign n33679 = n17415 ^ n15095 ^ n724 ;
  assign n33680 = ( ~n6347 & n10105 ) | ( ~n6347 & n33679 ) | ( n10105 & n33679 ) ;
  assign n33681 = n33680 ^ n1035 ^ 1'b0 ;
  assign n33682 = n9762 & n24897 ;
  assign n33683 = n17749 & n33682 ;
  assign n33684 = n14266 ^ n8868 ^ 1'b0 ;
  assign n33685 = n33683 | n33684 ;
  assign n33690 = n12243 ^ n9020 ^ 1'b0 ;
  assign n33686 = n4870 & ~n18442 ;
  assign n33687 = ~n8675 & n33686 ;
  assign n33688 = n33687 ^ n19195 ^ n5107 ;
  assign n33689 = ( n3785 & n8616 ) | ( n3785 & ~n33688 ) | ( n8616 & ~n33688 ) ;
  assign n33691 = n33690 ^ n33689 ^ n13182 ;
  assign n33692 = n31648 & n33101 ;
  assign n33693 = n33692 ^ n2258 ^ 1'b0 ;
  assign n33694 = n28006 ^ n21350 ^ n9941 ;
  assign n33695 = n23078 & n33694 ;
  assign n33696 = n13013 & n33695 ;
  assign n33697 = n862 & ~n4048 ;
  assign n33698 = n33697 ^ n7376 ^ 1'b0 ;
  assign n33699 = n4597 & ~n15111 ;
  assign n33700 = n21461 | n33699 ;
  assign n33701 = n33700 ^ n32326 ^ 1'b0 ;
  assign n33702 = n493 & ~n29926 ;
  assign n33703 = n15624 ^ n10789 ^ 1'b0 ;
  assign n33704 = n6080 | n33703 ;
  assign n33705 = n33704 ^ n11460 ^ 1'b0 ;
  assign n33706 = ~n14724 & n28598 ;
  assign n33707 = n33706 ^ n7824 ^ 1'b0 ;
  assign n33708 = ~n6488 & n27423 ;
  assign n33710 = n18840 ^ n855 ^ 1'b0 ;
  assign n33709 = n8480 & n31477 ;
  assign n33711 = n33710 ^ n33709 ^ 1'b0 ;
  assign n33712 = ~n511 & n6226 ;
  assign n33713 = n4846 & n11523 ;
  assign n33714 = n19387 & n33713 ;
  assign n33715 = n33714 ^ n23619 ^ 1'b0 ;
  assign n33716 = n33311 | n33715 ;
  assign n33717 = ~n11805 & n33716 ;
  assign n33718 = n33665 ^ n2233 ^ 1'b0 ;
  assign n33719 = n23571 & ~n33718 ;
  assign n33720 = n4451 & n13999 ;
  assign n33721 = ~n13175 & n26223 ;
  assign n33722 = n33721 ^ n10672 ^ 1'b0 ;
  assign n33723 = n17580 & n33722 ;
  assign n33724 = n33723 ^ n27655 ^ n15024 ;
  assign n33725 = n33724 ^ n19008 ^ 1'b0 ;
  assign n33726 = n5480 | n33725 ;
  assign n33727 = ( n5309 & n7030 ) | ( n5309 & ~n7734 ) | ( n7030 & ~n7734 ) ;
  assign n33728 = ( ~n1989 & n4859 ) | ( ~n1989 & n33727 ) | ( n4859 & n33727 ) ;
  assign n33729 = n6175 & n10106 ;
  assign n33730 = n7342 & n33729 ;
  assign n33731 = ~n24027 & n32226 ;
  assign n33738 = n1983 | n4486 ;
  assign n33739 = n33738 ^ n376 ^ 1'b0 ;
  assign n33736 = n18597 | n29090 ;
  assign n33737 = ~n16399 & n33736 ;
  assign n33732 = n10436 | n16743 ;
  assign n33733 = n33732 ^ n328 ^ 1'b0 ;
  assign n33734 = n28856 & n33733 ;
  assign n33735 = n33734 ^ n21145 ^ 1'b0 ;
  assign n33740 = n33739 ^ n33737 ^ n33735 ;
  assign n33741 = n9118 ^ n1031 ^ 1'b0 ;
  assign n33742 = n9585 & n33741 ;
  assign n33743 = n106 | n19302 ;
  assign n33744 = n33743 ^ n25104 ^ 1'b0 ;
  assign n33745 = n6915 & n11192 ;
  assign n33746 = ~n19324 & n31435 ;
  assign n33747 = n20733 & ~n33746 ;
  assign n33748 = n16893 | n20453 ;
  assign n33749 = n17607 | n33748 ;
  assign n33750 = n33749 ^ n15529 ^ n14184 ;
  assign n33751 = n33750 ^ n7672 ^ 1'b0 ;
  assign n33752 = n26848 | n31051 ;
  assign n33753 = n13620 ^ n13110 ^ 1'b0 ;
  assign n33754 = n33753 ^ n12586 ^ n10048 ;
  assign n33755 = ~n2796 & n8472 ;
  assign n33756 = n16463 ^ n16165 ^ 1'b0 ;
  assign n33757 = n33755 & n33756 ;
  assign n33758 = n21335 ^ n749 ^ 1'b0 ;
  assign n33759 = n18754 | n33758 ;
  assign n33760 = n4714 & n33759 ;
  assign n33761 = ~n20998 & n32277 ;
  assign n33762 = n27610 ^ n21277 ^ n12736 ;
  assign n33763 = n6033 & ~n33762 ;
  assign n33764 = n1477 & ~n33763 ;
  assign n33765 = n2701 | n3811 ;
  assign n33766 = n403 & ~n21054 ;
  assign n33767 = n33766 ^ n162 ^ 1'b0 ;
  assign n33768 = n33765 | n33767 ;
  assign n33769 = ~n2429 & n5461 ;
  assign n33770 = ~n11751 & n13092 ;
  assign n33771 = n31480 ^ n7766 ^ 1'b0 ;
  assign n33772 = n11811 & n14302 ;
  assign n33773 = n33772 ^ n32314 ^ 1'b0 ;
  assign n33774 = n18032 & ~n33773 ;
  assign n33775 = n2136 & ~n7579 ;
  assign n33776 = n33775 ^ n17759 ^ 1'b0 ;
  assign n33782 = n11940 ^ n8675 ^ 1'b0 ;
  assign n33783 = ( n10864 & n11005 ) | ( n10864 & ~n33782 ) | ( n11005 & ~n33782 ) ;
  assign n33777 = n19984 ^ n12511 ^ 1'b0 ;
  assign n33778 = n9048 & ~n25298 ;
  assign n33779 = n33777 | n33778 ;
  assign n33780 = n1655 & ~n33779 ;
  assign n33781 = n32294 | n33780 ;
  assign n33784 = n33783 ^ n33781 ^ 1'b0 ;
  assign n33785 = n14963 ^ n5297 ^ 1'b0 ;
  assign n33786 = n23490 & n33785 ;
  assign n33787 = ~n5803 & n25012 ;
  assign n33788 = n33787 ^ n3887 ^ 1'b0 ;
  assign n33789 = n24921 ^ n22389 ^ 1'b0 ;
  assign n33790 = ( ~n5049 & n7520 ) | ( ~n5049 & n16458 ) | ( n7520 & n16458 ) ;
  assign n33791 = n28519 ^ n5046 ^ 1'b0 ;
  assign n33792 = n14923 ^ n9113 ^ n5490 ;
  assign n33793 = ~n20223 & n33792 ;
  assign n33794 = n11060 ^ n10593 ^ 1'b0 ;
  assign n33795 = n9621 & ~n21786 ;
  assign n33796 = n6978 & ~n33795 ;
  assign n33797 = n33796 ^ n18416 ^ 1'b0 ;
  assign n33798 = n33794 & n33797 ;
  assign n33799 = ~n6045 & n6488 ;
  assign n33800 = n572 & n8621 ;
  assign n33801 = n33800 ^ n24580 ^ n11107 ;
  assign n33802 = n8958 | n12789 ;
  assign n33803 = n20804 ^ n10600 ^ 1'b0 ;
  assign n33804 = ~n7442 & n28715 ;
  assign n33805 = n12159 | n20563 ;
  assign n33806 = n2754 | n33805 ;
  assign n33807 = ~n5821 & n30455 ;
  assign n33808 = n33807 ^ n7294 ^ 1'b0 ;
  assign n33809 = n33806 & n33808 ;
  assign n33810 = n13463 ^ n7933 ^ 1'b0 ;
  assign n33811 = n17417 | n33810 ;
  assign n33812 = n14680 ^ n12967 ^ 1'b0 ;
  assign n33813 = n33811 | n33812 ;
  assign n33814 = n33813 ^ n29500 ^ 1'b0 ;
  assign n33815 = n3220 & ~n5374 ;
  assign n33816 = ~n26908 & n33815 ;
  assign n33817 = n3262 & ~n9159 ;
  assign n33818 = n16243 ^ n8697 ^ 1'b0 ;
  assign n33819 = ( ~n13414 & n33817 ) | ( ~n13414 & n33818 ) | ( n33817 & n33818 ) ;
  assign n33820 = n33819 ^ n14417 ^ 1'b0 ;
  assign n33821 = n5547 | n33820 ;
  assign n33822 = n33821 ^ n4558 ^ 1'b0 ;
  assign n33823 = ~n3242 & n26792 ;
  assign n33824 = n32126 ^ n25588 ^ n15892 ;
  assign n33825 = n31006 ^ n20652 ^ 1'b0 ;
  assign n33826 = n12101 | n29407 ;
  assign n33827 = n18675 ^ n10367 ^ 1'b0 ;
  assign n33828 = n3343 & n10692 ;
  assign n33829 = n7001 | n33828 ;
  assign n33830 = n33829 ^ n16953 ^ 1'b0 ;
  assign n33831 = n3225 & ~n33830 ;
  assign n33832 = ~n11801 & n12337 ;
  assign n33833 = n5293 ^ n4066 ^ 1'b0 ;
  assign n33834 = n8872 | n33833 ;
  assign n33835 = n21859 | n33834 ;
  assign n33836 = n14196 & ~n18209 ;
  assign n33837 = n605 & n33836 ;
  assign n33838 = n33837 ^ n28820 ^ n7556 ;
  assign n33839 = n8729 ^ n4485 ^ n4279 ;
  assign n33840 = n6959 ^ n4356 ^ 1'b0 ;
  assign n33841 = n8080 & n11740 ;
  assign n33842 = ~n6498 & n33841 ;
  assign n33843 = n12047 & n22226 ;
  assign n33844 = n33843 ^ n15793 ^ 1'b0 ;
  assign n33845 = ( n9332 & n9404 ) | ( n9332 & ~n17428 ) | ( n9404 & ~n17428 ) ;
  assign n33846 = n17675 ^ n733 ^ 1'b0 ;
  assign n33847 = ~n13833 & n33846 ;
  assign n33848 = n1293 & ~n2601 ;
  assign n33849 = n12058 & n29957 ;
  assign n33850 = ~n725 & n33849 ;
  assign n33851 = n20142 | n33850 ;
  assign n33852 = n5437 & n12238 ;
  assign n33853 = ~n6056 & n33852 ;
  assign n33854 = n12158 | n33853 ;
  assign n33855 = n6481 | n33854 ;
  assign n33856 = n849 | n20987 ;
  assign n33857 = n5935 ^ n4082 ^ 1'b0 ;
  assign n33858 = n11588 | n33857 ;
  assign n33859 = n26630 ^ n25354 ^ n14748 ;
  assign n33860 = n33859 ^ n14865 ^ 1'b0 ;
  assign n33861 = n11378 & ~n24341 ;
  assign n33862 = ~n31673 & n33861 ;
  assign n33863 = n3982 & n6583 ;
  assign n33864 = n19095 & n33863 ;
  assign n33865 = n20429 ^ n14085 ^ 1'b0 ;
  assign n33866 = n33865 ^ n991 ^ 1'b0 ;
  assign n33867 = n4741 ^ n1200 ^ 1'b0 ;
  assign n33868 = n33867 ^ n2367 ^ n2202 ;
  assign n33869 = n11164 ^ n1972 ^ 1'b0 ;
  assign n33872 = n1657 ^ n1321 ^ 1'b0 ;
  assign n33870 = n23705 ^ n19900 ^ 1'b0 ;
  assign n33871 = n10191 & ~n33870 ;
  assign n33873 = n33872 ^ n33871 ^ 1'b0 ;
  assign n33874 = n320 | n29476 ;
  assign n33875 = n33874 ^ n17809 ^ 1'b0 ;
  assign n33876 = n16113 ^ n8494 ^ 1'b0 ;
  assign n33877 = ~n15088 & n33876 ;
  assign n33878 = n19248 & ~n31782 ;
  assign n33879 = n10955 & n17704 ;
  assign n33880 = ~n26767 & n33879 ;
  assign n33881 = n6899 & n7189 ;
  assign n33882 = n17599 | n33881 ;
  assign n33883 = n17876 ^ n15285 ^ n7877 ;
  assign n33884 = ~n1645 & n3131 ;
  assign n33885 = n33884 ^ n26393 ^ 1'b0 ;
  assign n33886 = n19164 ^ n4687 ^ 1'b0 ;
  assign n33887 = n33885 & n33886 ;
  assign n33888 = ( n10538 & ~n12283 ) | ( n10538 & n12877 ) | ( ~n12283 & n12877 ) ;
  assign n33889 = n33888 ^ n18803 ^ 1'b0 ;
  assign n33890 = n5042 | n33889 ;
  assign n33891 = ( n4226 & n28400 ) | ( n4226 & n33890 ) | ( n28400 & n33890 ) ;
  assign n33892 = n3591 & n33891 ;
  assign n33893 = n10787 ^ n10048 ^ 1'b0 ;
  assign n33894 = n4797 | n6166 ;
  assign n33895 = n6540 | n33894 ;
  assign n33896 = n7268 & ~n12323 ;
  assign n33897 = n15224 ^ n14505 ^ 1'b0 ;
  assign n33898 = n12938 & n33897 ;
  assign n33899 = ~n10430 & n33898 ;
  assign n33900 = n33899 ^ n3440 ^ 1'b0 ;
  assign n33901 = n31108 & ~n33900 ;
  assign n33902 = n17608 & ~n24167 ;
  assign n33903 = ~n12040 & n33902 ;
  assign n33904 = n12675 | n20561 ;
  assign n33905 = n33904 ^ n9372 ^ 1'b0 ;
  assign n33906 = n20140 ^ n5747 ^ n579 ;
  assign n33907 = n4349 & ~n33906 ;
  assign n33908 = ~n33905 & n33907 ;
  assign n33909 = n22594 & n26825 ;
  assign n33910 = n28756 & n33909 ;
  assign n33911 = n1941 | n24117 ;
  assign n33912 = n33911 ^ n32186 ^ 1'b0 ;
  assign n33913 = n15 | n19293 ;
  assign n33914 = n3628 | n33913 ;
  assign n33915 = n1841 | n5543 ;
  assign n33916 = ~n21440 & n22924 ;
  assign n33917 = n26115 ^ n19896 ^ 1'b0 ;
  assign n33918 = n8220 & n33917 ;
  assign n33919 = n33918 ^ n21251 ^ 1'b0 ;
  assign n33922 = n2735 | n33543 ;
  assign n33920 = ~n2125 & n11525 ;
  assign n33921 = ~n18742 & n33920 ;
  assign n33923 = n33922 ^ n33921 ^ n7313 ;
  assign n33924 = n2614 | n6533 ;
  assign n33925 = n30393 | n33924 ;
  assign n33926 = n33925 ^ n4639 ^ 1'b0 ;
  assign n33928 = n3953 | n16296 ;
  assign n33929 = n6766 & ~n33928 ;
  assign n33930 = ~n15134 & n16069 ;
  assign n33931 = n33929 & n33930 ;
  assign n33927 = n2668 | n7825 ;
  assign n33932 = n33931 ^ n33927 ^ 1'b0 ;
  assign n33933 = n3558 | n5803 ;
  assign n33934 = n25555 & ~n33933 ;
  assign n33935 = n8981 & ~n20970 ;
  assign n33936 = n22445 & n33935 ;
  assign n33937 = n1349 | n33936 ;
  assign n33938 = n3772 & ~n33937 ;
  assign n33939 = n33710 & n33938 ;
  assign n33940 = n2914 & n8759 ;
  assign n33941 = n1993 & ~n33940 ;
  assign n33942 = n5136 & n30834 ;
  assign n33943 = n33942 ^ n12622 ^ 1'b0 ;
  assign n33944 = ~n12927 & n14429 ;
  assign n33945 = ~n16236 & n33944 ;
  assign n33946 = n14551 & n33945 ;
  assign n33947 = n4085 & ~n10489 ;
  assign n33948 = n26469 & ~n33947 ;
  assign n33949 = ~n32522 & n33948 ;
  assign n33950 = n16974 ^ n9104 ^ 1'b0 ;
  assign n33951 = n12317 & n16512 ;
  assign n33952 = ~n3686 & n33951 ;
  assign n33953 = n1522 & n33952 ;
  assign n33955 = n6727 ^ n3003 ^ 1'b0 ;
  assign n33954 = n15481 & n22683 ;
  assign n33956 = n33955 ^ n33954 ^ n15226 ;
  assign n33957 = n11738 & n12803 ;
  assign n33958 = ~n9324 & n33957 ;
  assign n33959 = n33958 ^ n15024 ^ 1'b0 ;
  assign n33960 = n12525 | n33959 ;
  assign n33961 = ~n2728 & n3367 ;
  assign n33962 = ~n4588 & n33961 ;
  assign n33963 = n33962 ^ n13254 ^ 1'b0 ;
  assign n33964 = n33963 ^ n22962 ^ 1'b0 ;
  assign n33965 = n1199 | n17677 ;
  assign n33966 = n22274 ^ n16747 ^ 1'b0 ;
  assign n33967 = n31144 ^ n12475 ^ 1'b0 ;
  assign n33968 = n30631 & ~n33967 ;
  assign n33969 = n33968 ^ n25161 ^ 1'b0 ;
  assign n33972 = n827 & n15416 ;
  assign n33970 = ~n5809 & n31797 ;
  assign n33971 = n33970 ^ n17737 ^ 1'b0 ;
  assign n33973 = n33972 ^ n33971 ^ n17293 ;
  assign n33974 = n29451 ^ n12937 ^ 1'b0 ;
  assign n33975 = ( ~n10300 & n16004 ) | ( ~n10300 & n24580 ) | ( n16004 & n24580 ) ;
  assign n33976 = n33975 ^ n12665 ^ n1085 ;
  assign n33977 = n17358 ^ n16563 ^ n3025 ;
  assign n33978 = ~n2920 & n12404 ;
  assign n33979 = n33978 ^ n31422 ^ 1'b0 ;
  assign n33980 = ( n7038 & n21059 ) | ( n7038 & ~n26159 ) | ( n21059 & ~n26159 ) ;
  assign n33981 = n28375 & ~n33980 ;
  assign n33982 = n33981 ^ n765 ^ 1'b0 ;
  assign n33983 = n13942 & n33982 ;
  assign n33984 = n33983 ^ n26666 ^ 1'b0 ;
  assign n33985 = n17841 & ~n33637 ;
  assign n33986 = n19665 ^ n9530 ^ 1'b0 ;
  assign n33987 = n17369 | n33986 ;
  assign n33988 = ~n10142 & n27263 ;
  assign n33989 = n33988 ^ n5219 ^ 1'b0 ;
  assign n33990 = n33989 ^ n10008 ^ 1'b0 ;
  assign n33991 = n2197 | n16923 ;
  assign n33993 = n13106 ^ n9736 ^ 1'b0 ;
  assign n33992 = n12889 & n14403 ;
  assign n33994 = n33993 ^ n33992 ^ n805 ;
  assign n33995 = n33991 | n33994 ;
  assign n33997 = n3054 ^ n1215 ^ 1'b0 ;
  assign n33996 = ~n6261 & n24164 ;
  assign n33998 = n33997 ^ n33996 ^ 1'b0 ;
  assign n33999 = n28208 ^ n26296 ^ 1'b0 ;
  assign n34000 = n17590 & n30748 ;
  assign n34001 = n2626 & n3611 ;
  assign n34002 = ~n3312 & n34001 ;
  assign n34003 = n16983 & n34002 ;
  assign n34004 = n1544 & n2225 ;
  assign n34005 = n1267 & n34004 ;
  assign n34006 = n9002 ^ n7007 ^ 1'b0 ;
  assign n34007 = n34006 ^ n31164 ^ 1'b0 ;
  assign n34008 = n408 & n9672 ;
  assign n34009 = ~n10816 & n29779 ;
  assign n34010 = n34009 ^ n1024 ^ 1'b0 ;
  assign n34011 = n21148 & n34010 ;
  assign n34012 = n8910 | n34011 ;
  assign n34013 = n16987 ^ n1445 ^ 1'b0 ;
  assign n34014 = n13404 | n34013 ;
  assign n34015 = n34014 ^ n10395 ^ 1'b0 ;
  assign n34016 = n34015 ^ n13327 ^ n3111 ;
  assign n34017 = n3597 & n6275 ;
  assign n34018 = n34017 ^ n23286 ^ 1'b0 ;
  assign n34019 = n25210 ^ n1377 ^ 1'b0 ;
  assign n34020 = n27003 | n34019 ;
  assign n34021 = n18041 ^ n17005 ^ 1'b0 ;
  assign n34022 = n4954 & ~n11885 ;
  assign n34023 = n13904 & n34022 ;
  assign n34024 = n2157 | n8922 ;
  assign n34025 = n34024 ^ n30599 ^ 1'b0 ;
  assign n34026 = ( n7614 & n20548 ) | ( n7614 & n31292 ) | ( n20548 & n31292 ) ;
  assign n34027 = ~n12479 & n29218 ;
  assign n34028 = n27268 ^ n25193 ^ 1'b0 ;
  assign n34032 = n14667 ^ n8159 ^ 1'b0 ;
  assign n34033 = n34032 ^ n10437 ^ 1'b0 ;
  assign n34034 = n34033 ^ n1659 ^ 1'b0 ;
  assign n34035 = n13393 & ~n34034 ;
  assign n34029 = n3466 ^ n1662 ^ 1'b0 ;
  assign n34030 = ~n7865 & n34029 ;
  assign n34031 = ( n6881 & n32469 ) | ( n6881 & n34030 ) | ( n32469 & n34030 ) ;
  assign n34036 = n34035 ^ n34031 ^ 1'b0 ;
  assign n34037 = n750 | n5880 ;
  assign n34038 = n34036 | n34037 ;
  assign n34039 = ( ~n2682 & n4962 ) | ( ~n2682 & n14173 ) | ( n4962 & n14173 ) ;
  assign n34040 = n26243 & ~n34039 ;
  assign n34041 = n34040 ^ n15649 ^ 1'b0 ;
  assign n34042 = ~n7040 & n34041 ;
  assign n34043 = n25067 | n27571 ;
  assign n34044 = n22115 ^ n19831 ^ n17079 ;
  assign n34045 = n16388 & ~n34044 ;
  assign n34046 = n13252 & n27093 ;
  assign n34047 = n7897 & ~n13230 ;
  assign n34048 = ( n9328 & ~n23749 ) | ( n9328 & n33834 ) | ( ~n23749 & n33834 ) ;
  assign n34049 = n17070 & n23547 ;
  assign n34050 = n34048 & n34049 ;
  assign n34051 = n1791 & ~n2525 ;
  assign n34052 = ~n107 & n34051 ;
  assign n34053 = n3238 & n34052 ;
  assign n34054 = n6903 ^ n6200 ^ 1'b0 ;
  assign n34055 = n26034 & n34054 ;
  assign n34056 = n6601 | n14373 ;
  assign n34057 = n1513 | n34056 ;
  assign n34058 = n8608 & n34057 ;
  assign n34059 = n33458 ^ n8716 ^ n3791 ;
  assign n34060 = ~n6906 & n34059 ;
  assign n34061 = n171 & ~n3221 ;
  assign n34062 = ~n34060 & n34061 ;
  assign n34063 = n23644 ^ n248 ^ 1'b0 ;
  assign n34064 = n21496 ^ n10022 ^ 1'b0 ;
  assign n34065 = n16469 | n24380 ;
  assign n34066 = n28745 ^ n25207 ^ n12935 ;
  assign n34067 = n10711 ^ n592 ^ 1'b0 ;
  assign n34068 = ~n8827 & n34067 ;
  assign n34069 = n34068 ^ n10651 ^ 1'b0 ;
  assign n34070 = n13290 ^ n7308 ^ 1'b0 ;
  assign n34071 = ~n16106 & n34070 ;
  assign n34072 = ( n5686 & ~n12773 ) | ( n5686 & n34071 ) | ( ~n12773 & n34071 ) ;
  assign n34073 = n23124 ^ n10372 ^ 1'b0 ;
  assign n34074 = n34072 & n34073 ;
  assign n34076 = n2929 ^ n1811 ^ 1'b0 ;
  assign n34077 = ~n4097 & n34076 ;
  assign n34078 = n1749 & ~n27787 ;
  assign n34079 = n18303 & n34078 ;
  assign n34080 = n24653 | n34079 ;
  assign n34081 = n34080 ^ n15909 ^ 1'b0 ;
  assign n34082 = ( n18371 & ~n34077 ) | ( n18371 & n34081 ) | ( ~n34077 & n34081 ) ;
  assign n34075 = n7568 ^ n228 ^ n105 ;
  assign n34083 = n34082 ^ n34075 ^ 1'b0 ;
  assign n34084 = n22584 ^ n11956 ^ 1'b0 ;
  assign n34085 = n3284 | n34084 ;
  assign n34086 = n13037 ^ n12585 ^ 1'b0 ;
  assign n34087 = ( n1985 & n6869 ) | ( n1985 & n20045 ) | ( n6869 & n20045 ) ;
  assign n34088 = n18511 ^ n12198 ^ 1'b0 ;
  assign n34089 = n10287 & n34088 ;
  assign n34090 = n34089 ^ n18360 ^ 1'b0 ;
  assign n34091 = ~n19400 & n34090 ;
  assign n34092 = ( n9139 & ~n9326 ) | ( n9139 & n11515 ) | ( ~n9326 & n11515 ) ;
  assign n34093 = n34092 ^ n11095 ^ 1'b0 ;
  assign n34094 = n17747 & ~n23254 ;
  assign n34095 = ~n11113 & n34094 ;
  assign n34096 = n5473 & n34095 ;
  assign n34097 = n4357 | n13359 ;
  assign n34098 = n34097 ^ n9896 ^ 1'b0 ;
  assign n34099 = n223 & n34098 ;
  assign n34100 = n34099 ^ n7454 ^ n5413 ;
  assign n34101 = n8147 & ~n28598 ;
  assign n34102 = n19529 ^ n1551 ^ 1'b0 ;
  assign n34103 = ~n7312 & n34102 ;
  assign n34104 = n488 & ~n34103 ;
  assign n34106 = n33929 ^ n1360 ^ 1'b0 ;
  assign n34107 = n34106 ^ n22572 ^ 1'b0 ;
  assign n34108 = n16828 & ~n34107 ;
  assign n34105 = n3163 & ~n7972 ;
  assign n34109 = n34108 ^ n34105 ^ 1'b0 ;
  assign n34110 = n5381 ^ n249 ^ 1'b0 ;
  assign n34111 = ~n15129 & n34110 ;
  assign n34112 = n6122 | n28172 ;
  assign n34113 = n8340 | n34112 ;
  assign n34114 = n14324 & n24162 ;
  assign n34115 = ( ~n15262 & n22075 ) | ( ~n15262 & n34114 ) | ( n22075 & n34114 ) ;
  assign n34116 = n34115 ^ n17499 ^ 1'b0 ;
  assign n34117 = n4947 & n10893 ;
  assign n34118 = ~n32566 & n34117 ;
  assign n34119 = n1377 | n1653 ;
  assign n34120 = n8978 | n34119 ;
  assign n34121 = n18494 ^ n9674 ^ 1'b0 ;
  assign n34122 = n4454 & ~n34121 ;
  assign n34123 = n34122 ^ n22888 ^ 1'b0 ;
  assign n34124 = ~n7257 & n34123 ;
  assign n34125 = n6442 & n34124 ;
  assign n34126 = n15071 & ~n34125 ;
  assign n34127 = n34120 & ~n34126 ;
  assign n34128 = ( ~n465 & n3574 ) | ( ~n465 & n4659 ) | ( n3574 & n4659 ) ;
  assign n34129 = ~n2423 & n32929 ;
  assign n34130 = n27832 ^ n9369 ^ 1'b0 ;
  assign n34131 = n3588 & ~n34130 ;
  assign n34132 = n26350 ^ n20759 ^ 1'b0 ;
  assign n34133 = n89 & n15598 ;
  assign n34134 = n25391 & ~n30651 ;
  assign n34135 = n5118 & ~n27738 ;
  assign n34136 = n34135 ^ n6048 ^ n2184 ;
  assign n34137 = n34136 ^ n25927 ^ 1'b0 ;
  assign n34138 = n7273 | n13486 ;
  assign n34139 = n5935 | n13623 ;
  assign n34140 = ~n20 & n5734 ;
  assign n34141 = ~n2921 & n34140 ;
  assign n34142 = n34141 ^ n3980 ^ 1'b0 ;
  assign n34144 = n26020 ^ n14894 ^ 1'b0 ;
  assign n34143 = n9193 & ~n27177 ;
  assign n34145 = n34144 ^ n34143 ^ 1'b0 ;
  assign n34146 = n5613 ^ n3302 ^ 1'b0 ;
  assign n34147 = ~n29464 & n34146 ;
  assign n34154 = n8433 & ~n8942 ;
  assign n34155 = n34154 ^ n19725 ^ 1'b0 ;
  assign n34152 = n15527 | n15752 ;
  assign n34151 = n11165 | n16889 ;
  assign n34153 = n34152 ^ n34151 ^ 1'b0 ;
  assign n34156 = n34155 ^ n34153 ^ 1'b0 ;
  assign n34148 = n30583 ^ n13797 ^ 1'b0 ;
  assign n34149 = ~n25276 & n34148 ;
  assign n34150 = ~n9588 & n34149 ;
  assign n34157 = n34156 ^ n34150 ^ 1'b0 ;
  assign n34158 = ~n34147 & n34157 ;
  assign n34159 = n25077 & n28642 ;
  assign n34160 = ~n34077 & n34159 ;
  assign n34161 = n2626 & n24309 ;
  assign n34162 = n23395 ^ n20826 ^ 1'b0 ;
  assign n34163 = n2045 & n34162 ;
  assign n34164 = n7546 ^ n6198 ^ 1'b0 ;
  assign n34165 = n34163 & ~n34164 ;
  assign n34166 = n7004 ^ n2137 ^ 1'b0 ;
  assign n34167 = n34166 ^ n6387 ^ 1'b0 ;
  assign n34168 = n1174 | n31380 ;
  assign n34169 = n24250 ^ n12862 ^ 1'b0 ;
  assign n34170 = n1522 | n13861 ;
  assign n34171 = n34170 ^ n32038 ^ 1'b0 ;
  assign n34172 = n34171 ^ n26324 ^ n14136 ;
  assign n34173 = n30239 ^ n14356 ^ 1'b0 ;
  assign n34174 = n4250 & ~n26573 ;
  assign n34175 = n34174 ^ n20172 ^ 1'b0 ;
  assign n34179 = n15430 ^ n7585 ^ 1'b0 ;
  assign n34176 = n13676 & n17620 ;
  assign n34177 = n34176 ^ n5562 ^ 1'b0 ;
  assign n34178 = n14885 & ~n34177 ;
  assign n34180 = n34179 ^ n34178 ^ n16400 ;
  assign n34181 = ~n26359 & n34180 ;
  assign n34182 = n32207 ^ n16769 ^ 1'b0 ;
  assign n34183 = n8728 | n21593 ;
  assign n34184 = ~n28499 & n33027 ;
  assign n34185 = ~n513 & n34184 ;
  assign n34186 = n3068 | n12428 ;
  assign n34187 = n34186 ^ n22443 ^ n9233 ;
  assign n34188 = n13422 & n27650 ;
  assign n34189 = n20318 ^ n12618 ^ 1'b0 ;
  assign n34190 = n5215 | n7971 ;
  assign n34191 = n34190 ^ n1590 ^ 1'b0 ;
  assign n34192 = n3413 & ~n16056 ;
  assign n34193 = n21714 ^ n738 ^ 1'b0 ;
  assign n34194 = n34192 | n34193 ;
  assign n34195 = n33813 ^ n26768 ^ 1'b0 ;
  assign n34196 = n28248 ^ n24653 ^ 1'b0 ;
  assign n34197 = n19146 | n34196 ;
  assign n34198 = n34197 ^ n7965 ^ 1'b0 ;
  assign n34199 = ~n6228 & n34198 ;
  assign n34200 = n18525 ^ n10706 ^ 1'b0 ;
  assign n34201 = n29963 ^ n18329 ^ n2101 ;
  assign n34202 = n7180 & n14448 ;
  assign n34203 = n1141 & n12589 ;
  assign n34204 = ~n5143 & n14773 ;
  assign n34205 = n22577 ^ n10970 ^ 1'b0 ;
  assign n34206 = n5257 | n34205 ;
  assign n34207 = ~n946 & n8091 ;
  assign n34208 = n19101 ^ n6946 ^ 1'b0 ;
  assign n34209 = ~n4442 & n14011 ;
  assign n34210 = n1141 & n34209 ;
  assign n34211 = ~n10795 & n34210 ;
  assign n34212 = n1143 & n34211 ;
  assign n34213 = n2137 ^ n2000 ^ 1'b0 ;
  assign n34214 = n14369 | n34213 ;
  assign n34215 = n24065 & ~n34214 ;
  assign n34216 = n23888 ^ n14525 ^ 1'b0 ;
  assign n34217 = ~n34215 & n34216 ;
  assign n34218 = n7455 ^ n7252 ^ 1'b0 ;
  assign n34219 = n17795 & n34218 ;
  assign n34220 = ( n2600 & n6206 ) | ( n2600 & ~n14635 ) | ( n6206 & ~n14635 ) ;
  assign n34221 = n10702 | n23307 ;
  assign n34222 = n34221 ^ n11077 ^ 1'b0 ;
  assign n34223 = n34222 ^ n24381 ^ 1'b0 ;
  assign n34224 = n13966 ^ n5965 ^ 1'b0 ;
  assign n34225 = n2236 & n22636 ;
  assign n34226 = n34225 ^ n15757 ^ 1'b0 ;
  assign n34227 = n23919 ^ n22917 ^ 1'b0 ;
  assign n34228 = n18871 & n34227 ;
  assign n34229 = n25651 ^ n16458 ^ 1'b0 ;
  assign n34230 = ~n21791 & n34229 ;
  assign n34231 = n3225 & n17608 ;
  assign n34232 = ~n27834 & n34231 ;
  assign n34233 = n28043 ^ n1114 ^ 1'b0 ;
  assign n34234 = n18549 & ~n25500 ;
  assign n34235 = n34234 ^ n23891 ^ 1'b0 ;
  assign n34236 = n34235 ^ n27523 ^ 1'b0 ;
  assign n34238 = n11642 ^ n7789 ^ 1'b0 ;
  assign n34239 = n127 | n25516 ;
  assign n34240 = n34238 | n34239 ;
  assign n34237 = n27340 ^ n25114 ^ 1'b0 ;
  assign n34241 = n34240 ^ n34237 ^ 1'b0 ;
  assign n34242 = ~n2635 & n7566 ;
  assign n34243 = n297 & ~n1442 ;
  assign n34244 = n32551 ^ n14439 ^ 1'b0 ;
  assign n34245 = ~n2203 & n27877 ;
  assign n34246 = n5036 & n5513 ;
  assign n34247 = n34246 ^ n2655 ^ n2244 ;
  assign n34248 = ~n11891 & n23402 ;
  assign n34249 = ~n19595 & n34248 ;
  assign n34250 = n2404 & ~n34249 ;
  assign n34251 = n34250 ^ n12664 ^ 1'b0 ;
  assign n34252 = n4962 & n19072 ;
  assign n34253 = ( n43 & n724 ) | ( n43 & ~n2728 ) | ( n724 & ~n2728 ) ;
  assign n34254 = ~n7369 & n34253 ;
  assign n34255 = n34254 ^ n5369 ^ n1821 ;
  assign n34256 = n17387 ^ n8987 ^ 1'b0 ;
  assign n34257 = n34256 ^ n33249 ^ 1'b0 ;
  assign n34258 = n3584 & ~n28751 ;
  assign n34259 = n7568 | n16252 ;
  assign n34260 = ~n16923 & n34259 ;
  assign n34261 = n34260 ^ n15915 ^ 1'b0 ;
  assign n34262 = n6934 ^ n695 ^ 1'b0 ;
  assign n34263 = ~n13454 & n22990 ;
  assign n34264 = n1670 & n14080 ;
  assign n34265 = ~n21938 & n34264 ;
  assign n34266 = n34263 & n34265 ;
  assign n34267 = ~n2671 & n11918 ;
  assign n34268 = n34267 ^ n5700 ^ 1'b0 ;
  assign n34269 = n10775 & ~n11692 ;
  assign n34270 = n8659 & n15231 ;
  assign n34271 = n7990 & ~n34270 ;
  assign n34272 = n34271 ^ n6166 ^ 1'b0 ;
  assign n34273 = n34272 ^ n2552 ^ 1'b0 ;
  assign n34274 = n34273 ^ n10263 ^ 1'b0 ;
  assign n34275 = n34274 ^ n13833 ^ 1'b0 ;
  assign n34276 = n3688 & n20785 ;
  assign n34277 = n34276 ^ n6102 ^ 1'b0 ;
  assign n34278 = ~n30641 & n34277 ;
  assign n34279 = n34278 ^ n18772 ^ 1'b0 ;
  assign n34280 = n10277 & ~n29060 ;
  assign n34281 = n34280 ^ n27916 ^ 1'b0 ;
  assign n34282 = ~n7949 & n34281 ;
  assign n34283 = ~n2338 & n20015 ;
  assign n34284 = n11055 ^ n4479 ^ 1'b0 ;
  assign n34285 = n12421 | n13376 ;
  assign n34286 = n11577 ^ n8287 ^ 1'b0 ;
  assign n34287 = n31566 ^ n28306 ^ 1'b0 ;
  assign n34288 = n7233 ^ n5237 ^ 1'b0 ;
  assign n34289 = n15915 | n28155 ;
  assign n34290 = n30539 ^ n29325 ^ n7792 ;
  assign n34291 = n34290 ^ n4949 ^ 1'b0 ;
  assign n34292 = n34289 & n34291 ;
  assign n34293 = n34292 ^ n16040 ^ 1'b0 ;
  assign n34294 = n2885 | n8936 ;
  assign n34295 = n29452 | n34294 ;
  assign n34296 = ~n1851 & n11065 ;
  assign n34297 = ~n34295 & n34296 ;
  assign n34298 = ~n1711 & n14348 ;
  assign n34299 = n34298 ^ n22737 ^ 1'b0 ;
  assign n34300 = n16497 & n34299 ;
  assign n34301 = n17677 & n34300 ;
  assign n34302 = n1783 & n4651 ;
  assign n34303 = n34302 ^ n21386 ^ n11392 ;
  assign n34304 = ~n26240 & n27368 ;
  assign n34305 = ~n34303 & n34304 ;
  assign n34306 = n32697 ^ n291 ^ 1'b0 ;
  assign n34307 = ~n34305 & n34306 ;
  assign n34308 = n1337 & n20999 ;
  assign n34311 = n4280 & ~n8110 ;
  assign n34312 = n34311 ^ n10207 ^ 1'b0 ;
  assign n34313 = ~n323 & n34312 ;
  assign n34309 = n635 & n23318 ;
  assign n34310 = n34309 ^ n2930 ^ 1'b0 ;
  assign n34314 = n34313 ^ n34310 ^ n15452 ;
  assign n34315 = n29280 ^ n15078 ^ 1'b0 ;
  assign n34316 = n5991 | n10315 ;
  assign n34317 = n27980 | n34316 ;
  assign n34318 = n13015 ^ n1933 ^ 1'b0 ;
  assign n34319 = n26511 & ~n30262 ;
  assign n34320 = n17993 ^ n592 ^ 1'b0 ;
  assign n34321 = n9205 & n32377 ;
  assign n34322 = n34321 ^ n26441 ^ 1'b0 ;
  assign n34323 = n2767 | n5103 ;
  assign n34324 = n14680 & ~n34323 ;
  assign n34325 = n34324 ^ n11162 ^ 1'b0 ;
  assign n34326 = n7952 & n19360 ;
  assign n34327 = ( n21748 & ~n34325 ) | ( n21748 & n34326 ) | ( ~n34325 & n34326 ) ;
  assign n34328 = n15236 & ~n26892 ;
  assign n34329 = n34327 | n34328 ;
  assign n34330 = n3822 | n34329 ;
  assign n34331 = n26282 ^ n17470 ^ 1'b0 ;
  assign n34332 = n22173 | n34331 ;
  assign n34333 = n31176 ^ n18022 ^ 1'b0 ;
  assign n34334 = n2941 & ~n34333 ;
  assign n34335 = n34334 ^ n26967 ^ 1'b0 ;
  assign n34336 = ~n2811 & n5991 ;
  assign n34337 = n7437 & ~n10223 ;
  assign n34338 = n27326 & n34337 ;
  assign n34339 = n28395 ^ n26359 ^ n10205 ;
  assign n34340 = n24776 ^ n2671 ^ 1'b0 ;
  assign n34341 = n8663 & n34340 ;
  assign n34342 = n2835 & n34341 ;
  assign n34343 = ~n6282 & n34342 ;
  assign n34344 = n23203 ^ n7550 ^ 1'b0 ;
  assign n34345 = n13024 ^ n12673 ^ 1'b0 ;
  assign n34346 = n29606 ^ n6616 ^ 1'b0 ;
  assign n34347 = n23375 & n26176 ;
  assign n34348 = ~n5906 & n17527 ;
  assign n34349 = n34348 ^ n1422 ^ 1'b0 ;
  assign n34350 = n12617 & n34349 ;
  assign n34351 = n13900 & ~n34350 ;
  assign n34352 = n1987 & ~n5138 ;
  assign n34353 = n6898 & ~n14602 ;
  assign n34354 = n1534 & ~n26743 ;
  assign n34355 = ~n2376 & n32870 ;
  assign n34356 = ~n3524 & n13482 ;
  assign n34357 = n7294 & ~n34356 ;
  assign n34358 = n30868 ^ n15270 ^ 1'b0 ;
  assign n34359 = n3748 & n34358 ;
  assign n34360 = n11198 ^ n2555 ^ 1'b0 ;
  assign n34361 = n26322 | n34360 ;
  assign n34362 = ~n14304 & n18955 ;
  assign n34363 = ~n7238 & n34362 ;
  assign n34364 = ~n8126 & n18328 ;
  assign n34365 = n34364 ^ n20245 ^ 1'b0 ;
  assign n34366 = ~n34363 & n34365 ;
  assign n34367 = n9794 | n21436 ;
  assign n34368 = n34367 ^ n29022 ^ 1'b0 ;
  assign n34369 = n116 | n2583 ;
  assign n34370 = n2583 & ~n34369 ;
  assign n34371 = n509 & ~n856 ;
  assign n34372 = n34370 & n34371 ;
  assign n34373 = n34372 ^ n2927 ^ 1'b0 ;
  assign n34374 = n12570 | n34373 ;
  assign n34375 = n34373 & ~n34374 ;
  assign n34376 = n1251 & n4263 ;
  assign n34377 = n34375 & n34376 ;
  assign n34378 = n2473 | n34377 ;
  assign n34379 = n34377 & ~n34378 ;
  assign n34383 = n2492 & ~n9277 ;
  assign n34384 = ( n11249 & n14380 ) | ( n11249 & n34383 ) | ( n14380 & n34383 ) ;
  assign n34382 = n7391 & n8611 ;
  assign n34385 = n34384 ^ n34382 ^ 1'b0 ;
  assign n34380 = n29983 ^ n13477 ^ 1'b0 ;
  assign n34381 = n22628 | n34380 ;
  assign n34386 = n34385 ^ n34381 ^ 1'b0 ;
  assign n34387 = n34379 | n34386 ;
  assign n34388 = n34387 ^ n4701 ^ 1'b0 ;
  assign n34389 = ~n2467 & n25201 ;
  assign n34390 = n26152 | n34389 ;
  assign n34391 = n17434 & ~n34390 ;
  assign n34392 = n27080 ^ n5151 ^ 1'b0 ;
  assign n34393 = n5538 | n34392 ;
  assign n34394 = n11277 ^ n5638 ^ 1'b0 ;
  assign n34395 = n13559 & ~n21514 ;
  assign n34396 = n13059 ^ n9949 ^ 1'b0 ;
  assign n34397 = n34041 | n34396 ;
  assign n34398 = ( ~n5773 & n9497 ) | ( ~n5773 & n23025 ) | ( n9497 & n23025 ) ;
  assign n34399 = n14228 ^ n5810 ^ 1'b0 ;
  assign n34400 = n10248 & n34399 ;
  assign n34401 = n12776 | n18064 ;
  assign n34402 = ~n14500 & n34401 ;
  assign n34403 = n9468 & n31856 ;
  assign n34404 = n18779 ^ n2689 ^ 1'b0 ;
  assign n34405 = ~n20943 & n34404 ;
  assign n34406 = n33393 ^ n19070 ^ 1'b0 ;
  assign n34407 = n9770 & n34406 ;
  assign n34408 = ~n34405 & n34407 ;
  assign n34409 = n14082 & ~n34408 ;
  assign n34410 = n34409 ^ n16174 ^ 1'b0 ;
  assign n34412 = n10022 ^ n9975 ^ n2961 ;
  assign n34413 = n1880 | n34412 ;
  assign n34411 = n5765 ^ n395 ^ 1'b0 ;
  assign n34414 = n34413 ^ n34411 ^ n9264 ;
  assign n34415 = n2411 & ~n7025 ;
  assign n34418 = n12828 ^ n8119 ^ n5728 ;
  assign n34419 = n2109 | n34418 ;
  assign n34420 = n34419 ^ n10866 ^ 1'b0 ;
  assign n34421 = n7949 ^ n6714 ^ 1'b0 ;
  assign n34422 = n34420 | n34421 ;
  assign n34416 = ~n6557 & n11300 ;
  assign n34417 = n25911 & n34416 ;
  assign n34423 = n34422 ^ n34417 ^ 1'b0 ;
  assign n34424 = n17427 & ~n30922 ;
  assign n34425 = n31785 ^ n1298 ^ 1'b0 ;
  assign n34426 = ~n4331 & n34425 ;
  assign n34427 = ~n774 & n14384 ;
  assign n34429 = n1497 & ~n9719 ;
  assign n34430 = ~n8174 & n34429 ;
  assign n34431 = n15170 & ~n34430 ;
  assign n34432 = n4140 & n34431 ;
  assign n34428 = n8124 | n33218 ;
  assign n34433 = n34432 ^ n34428 ^ 1'b0 ;
  assign n34434 = n34433 ^ n25104 ^ 1'b0 ;
  assign n34435 = ~n34427 & n34434 ;
  assign n34436 = ~n20844 & n34435 ;
  assign n34437 = n34436 ^ n28872 ^ 1'b0 ;
  assign n34438 = n7080 ^ n4264 ^ 1'b0 ;
  assign n34439 = n14472 ^ n4056 ^ 1'b0 ;
  assign n34440 = n24945 & ~n34439 ;
  assign n34441 = n13183 & ~n24310 ;
  assign n34442 = n29276 ^ n20980 ^ 1'b0 ;
  assign n34443 = n27957 | n34442 ;
  assign n34444 = n12050 ^ n9612 ^ n7241 ;
  assign n34445 = n12563 ^ n9810 ^ 1'b0 ;
  assign n34446 = ( ~n4409 & n22796 ) | ( ~n4409 & n34445 ) | ( n22796 & n34445 ) ;
  assign n34447 = n34446 ^ n30309 ^ 1'b0 ;
  assign n34448 = ~n16453 & n27459 ;
  assign n34449 = n34448 ^ n4444 ^ 1'b0 ;
  assign n34450 = n6366 ^ n5632 ^ n3383 ;
  assign n34451 = n34449 | n34450 ;
  assign n34452 = n29354 ^ n13597 ^ 1'b0 ;
  assign n34453 = n6370 | n34452 ;
  assign n34455 = ~n188 & n4570 ;
  assign n34454 = n8366 & ~n10673 ;
  assign n34456 = n34455 ^ n34454 ^ 1'b0 ;
  assign n34457 = n17182 ^ n3359 ^ 1'b0 ;
  assign n34459 = n7932 & ~n9983 ;
  assign n34460 = n11659 & n34459 ;
  assign n34461 = n13 | n34460 ;
  assign n34462 = n34461 ^ n15776 ^ 1'b0 ;
  assign n34458 = n1834 | n19978 ;
  assign n34463 = n34462 ^ n34458 ^ 1'b0 ;
  assign n34464 = n18218 & n32852 ;
  assign n34465 = n607 | n22425 ;
  assign n34466 = n34465 ^ n23402 ^ 1'b0 ;
  assign n34467 = n9629 ^ n9190 ^ 1'b0 ;
  assign n34468 = n18348 | n34467 ;
  assign n34469 = n34468 ^ n11435 ^ 1'b0 ;
  assign n34470 = n11552 | n17634 ;
  assign n34471 = n34470 ^ n7965 ^ 1'b0 ;
  assign n34472 = ~n34469 & n34471 ;
  assign n34473 = n2395 & n34472 ;
  assign n34474 = n10156 ^ n8327 ^ 1'b0 ;
  assign n34475 = n34474 ^ n8519 ^ n3917 ;
  assign n34476 = n14261 | n15495 ;
  assign n34477 = n34476 ^ n248 ^ 1'b0 ;
  assign n34478 = n28928 | n34477 ;
  assign n34479 = n2895 & ~n13831 ;
  assign n34480 = ~n10729 & n34479 ;
  assign n34481 = n34480 ^ n16337 ^ 1'b0 ;
  assign n34482 = n2387 & n34481 ;
  assign n34483 = ~n13180 & n34482 ;
  assign n34484 = n16119 & ~n20755 ;
  assign n34485 = n34484 ^ n22648 ^ 1'b0 ;
  assign n34486 = n21383 & ~n34485 ;
  assign n34487 = ~n27459 & n34486 ;
  assign n34488 = n9725 | n19688 ;
  assign n34489 = n5001 & ~n34488 ;
  assign n34490 = n34487 & n34489 ;
  assign n34491 = n13302 ^ n627 ^ 1'b0 ;
  assign n34492 = x1 & n8916 ;
  assign n34493 = n7011 & n34492 ;
  assign n34494 = n1550 & ~n34493 ;
  assign n34495 = n34494 ^ n26038 ^ 1'b0 ;
  assign n34496 = n33572 ^ n11977 ^ n6984 ;
  assign n34497 = n34496 ^ n12176 ^ 1'b0 ;
  assign n34498 = n9720 & ~n34497 ;
  assign n34499 = n34495 & ~n34498 ;
  assign n34500 = n15586 ^ n8672 ^ n2867 ;
  assign n34501 = ~n33209 & n34500 ;
  assign n34502 = n7767 & n34501 ;
  assign n34503 = n11708 & ~n26216 ;
  assign n34504 = n34503 ^ n15622 ^ 1'b0 ;
  assign n34505 = ~n3524 & n25319 ;
  assign n34506 = n34505 ^ n12585 ^ 1'b0 ;
  assign n34507 = n15542 ^ n15508 ^ 1'b0 ;
  assign n34508 = n34506 & ~n34507 ;
  assign n34509 = n22633 & n34508 ;
  assign n34510 = n34509 ^ n24094 ^ 1'b0 ;
  assign n34511 = n17243 | n27849 ;
  assign n34512 = n34511 ^ n31005 ^ 1'b0 ;
  assign n34513 = n727 & ~n5465 ;
  assign n34514 = n34512 & n34513 ;
  assign n34515 = n14759 ^ n2478 ^ 1'b0 ;
  assign n34516 = n2526 & n21506 ;
  assign n34517 = n4328 & n34516 ;
  assign n34518 = n1161 & ~n10530 ;
  assign n34519 = n765 & ~n34518 ;
  assign n34520 = n848 | n5571 ;
  assign n34521 = n34520 ^ n1275 ^ 1'b0 ;
  assign n34522 = n7507 | n32248 ;
  assign n34523 = n18553 | n34522 ;
  assign n34524 = n29090 ^ n22661 ^ 1'b0 ;
  assign n34525 = ~n19563 & n34475 ;
  assign n34526 = n551 | n559 ;
  assign n34527 = n34526 ^ n13519 ^ 1'b0 ;
  assign n34528 = n34527 ^ n4639 ^ 1'b0 ;
  assign n34529 = n10877 & n34528 ;
  assign n34530 = n26625 & n34529 ;
  assign n34531 = ~n16849 & n34530 ;
  assign n34532 = ( n522 & n15165 ) | ( n522 & ~n23506 ) | ( n15165 & ~n23506 ) ;
  assign n34533 = n8906 | n9703 ;
  assign n34534 = n17938 & n27804 ;
  assign n34535 = n34534 ^ n3486 ^ 1'b0 ;
  assign n34536 = n725 & n27214 ;
  assign n34537 = ~n30404 & n34536 ;
  assign n34538 = n30637 ^ n25691 ^ n9090 ;
  assign n34539 = n8195 ^ n3671 ^ 1'b0 ;
  assign n34540 = n6200 & ~n32946 ;
  assign n34541 = ~n15760 & n31766 ;
  assign n34542 = n3849 & n29098 ;
  assign n34543 = n16399 & n29500 ;
  assign n34544 = n6238 & ~n9802 ;
  assign n34545 = n34544 ^ n4960 ^ 1'b0 ;
  assign n34546 = n34545 ^ n6545 ^ n1845 ;
  assign n34547 = n8675 ^ n1394 ^ 1'b0 ;
  assign n34548 = ~n15390 & n34547 ;
  assign n34549 = n6122 & ~n20002 ;
  assign n34550 = n13520 & ~n34549 ;
  assign n34551 = ~n14587 & n16016 ;
  assign n34552 = n12400 & ~n16504 ;
  assign n34553 = n34552 ^ n2747 ^ 1'b0 ;
  assign n34554 = ~n9693 & n34553 ;
  assign n34555 = n34554 ^ n3221 ^ 1'b0 ;
  assign n34556 = n17707 ^ n4819 ^ 1'b0 ;
  assign n34558 = n6714 & ~n22884 ;
  assign n34557 = ~n5584 & n23049 ;
  assign n34559 = n34558 ^ n34557 ^ 1'b0 ;
  assign n34560 = n34559 ^ n8136 ^ 1'b0 ;
  assign n34561 = ~n4547 & n34560 ;
  assign n34562 = n27651 ^ n22802 ^ 1'b0 ;
  assign n34563 = n15800 ^ n11012 ^ 1'b0 ;
  assign n34564 = ~n33593 & n34563 ;
  assign n34565 = n220 & n9760 ;
  assign n34566 = n10851 ^ n8987 ^ 1'b0 ;
  assign n34567 = n2638 ^ n1072 ^ 1'b0 ;
  assign n34568 = n17601 | n34567 ;
  assign n34569 = n5350 & ~n10394 ;
  assign n34570 = ~n9508 & n11111 ;
  assign n34573 = ~n1985 & n26384 ;
  assign n34574 = n34573 ^ n14080 ^ 1'b0 ;
  assign n34571 = n492 | n20226 ;
  assign n34572 = n10391 & n34571 ;
  assign n34575 = n34574 ^ n34572 ^ 1'b0 ;
  assign n34576 = ( ~n6796 & n10486 ) | ( ~n6796 & n11123 ) | ( n10486 & n11123 ) ;
  assign n34577 = ~n27727 & n34576 ;
  assign n34578 = ~n1434 & n18858 ;
  assign n34579 = n34578 ^ n3093 ^ 1'b0 ;
  assign n34580 = ~n13675 & n34579 ;
  assign n34581 = ~n11055 & n34580 ;
  assign n34582 = n6787 | n13884 ;
  assign n34583 = n298 | n10852 ;
  assign n34584 = n10681 | n34583 ;
  assign n34585 = n9253 ^ n5073 ^ 1'b0 ;
  assign n34586 = n34584 & ~n34585 ;
  assign n34587 = n2164 | n22126 ;
  assign n34588 = n34586 | n34587 ;
  assign n34589 = ~n16126 & n34588 ;
  assign n34590 = ~n34582 & n34589 ;
  assign n34591 = n8091 ^ n6428 ^ 1'b0 ;
  assign n34592 = n25273 | n34591 ;
  assign n34593 = n34592 ^ n6834 ^ 1'b0 ;
  assign n34594 = n3050 & ~n8262 ;
  assign n34595 = n8209 | n33257 ;
  assign n34596 = n34594 & ~n34595 ;
  assign n34597 = ~n30661 & n30670 ;
  assign n34599 = ( ~n2458 & n12698 ) | ( ~n2458 & n20330 ) | ( n12698 & n20330 ) ;
  assign n34598 = n5936 & ~n24108 ;
  assign n34600 = n34599 ^ n34598 ^ 1'b0 ;
  assign n34601 = n12947 ^ n10235 ^ 1'b0 ;
  assign n34602 = n13422 ^ n1545 ^ 1'b0 ;
  assign n34603 = n34601 & n34602 ;
  assign n34604 = n22293 & ~n26068 ;
  assign n34605 = ~n3531 & n22135 ;
  assign n34606 = n34605 ^ n23595 ^ 1'b0 ;
  assign n34607 = n9375 & ~n10468 ;
  assign n34608 = ~n34606 & n34607 ;
  assign n34609 = n20172 | n31290 ;
  assign n34610 = n34609 ^ n23133 ^ 1'b0 ;
  assign n34611 = n13763 & ~n24531 ;
  assign n34612 = n17324 ^ n9570 ^ 1'b0 ;
  assign n34613 = n23936 ^ n4164 ^ 1'b0 ;
  assign n34614 = n22454 & ~n34613 ;
  assign n34615 = n2917 | n9287 ;
  assign n34616 = n21611 ^ n21291 ^ 1'b0 ;
  assign n34617 = n34171 ^ n2051 ^ 1'b0 ;
  assign n34618 = n4613 | n10056 ;
  assign n34619 = n5751 | n12302 ;
  assign n34620 = n3225 | n5418 ;
  assign n34621 = n3187 | n3292 ;
  assign n34622 = n34620 | n34621 ;
  assign n34624 = n8482 & n12338 ;
  assign n34625 = n34624 ^ n1174 ^ 1'b0 ;
  assign n34626 = n34625 ^ n20520 ^ 1'b0 ;
  assign n34623 = n9433 & ~n21719 ;
  assign n34627 = n34626 ^ n34623 ^ 1'b0 ;
  assign n34628 = ( n3330 & ~n19146 ) | ( n3330 & n34627 ) | ( ~n19146 & n34627 ) ;
  assign n34629 = ~n14738 & n23506 ;
  assign n34630 = n34629 ^ n22709 ^ 1'b0 ;
  assign n34631 = n13264 ^ n8263 ^ 1'b0 ;
  assign n34632 = ( ~n8973 & n9416 ) | ( ~n8973 & n34631 ) | ( n9416 & n34631 ) ;
  assign n34633 = n9611 & n34632 ;
  assign n34634 = ( n7287 & n17172 ) | ( n7287 & ~n18275 ) | ( n17172 & ~n18275 ) ;
  assign n34635 = n20573 ^ n9923 ^ 1'b0 ;
  assign n34636 = n16455 & n34635 ;
  assign n34637 = ~n5423 & n34636 ;
  assign n34638 = ~n10550 & n34637 ;
  assign n34639 = n3706 & ~n21239 ;
  assign n34640 = n1435 | n34639 ;
  assign n34641 = n34640 ^ n4180 ^ 1'b0 ;
  assign n34642 = ~n5005 & n34641 ;
  assign n34643 = n31262 & n34642 ;
  assign n34644 = ~n11818 & n22017 ;
  assign n34645 = n34644 ^ n23395 ^ 1'b0 ;
  assign n34646 = n13520 ^ n9792 ^ 1'b0 ;
  assign n34647 = n1055 & ~n22243 ;
  assign n34648 = n423 | n25675 ;
  assign n34649 = n34648 ^ n29486 ^ 1'b0 ;
  assign n34650 = n33632 & ~n34649 ;
  assign n34651 = n16395 ^ n11688 ^ 1'b0 ;
  assign n34652 = n26991 | n34651 ;
  assign n34653 = n2634 | n4810 ;
  assign n34654 = n34652 & ~n34653 ;
  assign n34655 = ( n1962 & ~n26352 ) | ( n1962 & n27761 ) | ( ~n26352 & n27761 ) ;
  assign n34656 = ( n6028 & ~n7469 ) | ( n6028 & n16536 ) | ( ~n7469 & n16536 ) ;
  assign n34657 = n26625 ^ n372 ^ 1'b0 ;
  assign n34658 = n20460 | n34657 ;
  assign n34659 = n23794 ^ n18871 ^ 1'b0 ;
  assign n34660 = n13792 & ~n34659 ;
  assign n34661 = n6662 & ~n28278 ;
  assign n34662 = n277 & n34661 ;
  assign n34663 = n22974 ^ n14156 ^ 1'b0 ;
  assign n34664 = n34662 | n34663 ;
  assign n34665 = n1244 & n7418 ;
  assign n34666 = n10196 & ~n34665 ;
  assign n34667 = ~n6871 & n34666 ;
  assign n34668 = n9785 | n11852 ;
  assign n34669 = n2671 | n34668 ;
  assign n34670 = n10582 | n18121 ;
  assign n34671 = n28012 ^ n1966 ^ 1'b0 ;
  assign n34676 = ~n1141 & n3166 ;
  assign n34677 = n34676 ^ n9880 ^ 1'b0 ;
  assign n34678 = n4962 & ~n34677 ;
  assign n34673 = ~n489 & n8778 ;
  assign n34674 = ~n1211 & n34673 ;
  assign n34675 = n12985 & n34674 ;
  assign n34672 = ( ~n4636 & n5697 ) | ( ~n4636 & n9821 ) | ( n5697 & n9821 ) ;
  assign n34679 = n34678 ^ n34675 ^ n34672 ;
  assign n34680 = ( ~n8309 & n10312 ) | ( ~n8309 & n34679 ) | ( n10312 & n34679 ) ;
  assign n34681 = n7160 & n34122 ;
  assign n34682 = n5095 & n34681 ;
  assign n34683 = n27674 | n34682 ;
  assign n34684 = n11878 & ~n34683 ;
  assign n34685 = ~n74 & n24081 ;
  assign n34686 = n832 | n34685 ;
  assign n34687 = n262 & ~n34686 ;
  assign n34688 = n12549 ^ n8430 ^ n2735 ;
  assign n34689 = n34688 ^ n26286 ^ n15523 ;
  assign n34690 = n9203 & n19821 ;
  assign n34691 = n34690 ^ n25614 ^ 1'b0 ;
  assign n34692 = ~n11273 & n31608 ;
  assign n34693 = n34692 ^ n10598 ^ 1'b0 ;
  assign n34699 = n3409 | n14818 ;
  assign n34694 = n33962 ^ n26369 ^ 1'b0 ;
  assign n34695 = n9053 & ~n34694 ;
  assign n34696 = n34695 ^ n26099 ^ 1'b0 ;
  assign n34697 = n34696 ^ n26304 ^ 1'b0 ;
  assign n34698 = n7919 & n34697 ;
  assign n34700 = n34699 ^ n34698 ^ 1'b0 ;
  assign n34701 = n6419 & ~n7340 ;
  assign n34702 = ~n3233 & n34701 ;
  assign n34703 = n19442 ^ n7837 ^ 1'b0 ;
  assign n34704 = ~n2683 & n34703 ;
  assign n34705 = n34702 | n34704 ;
  assign n34706 = n11456 & n34705 ;
  assign n34707 = n1210 & n34706 ;
  assign n34708 = n5789 & n23223 ;
  assign n34709 = n3544 & n34708 ;
  assign n34710 = n34709 ^ n20201 ^ n6039 ;
  assign n34711 = ~n8503 & n17924 ;
  assign n34712 = n34710 & n34711 ;
  assign n34714 = ~n2195 & n5499 ;
  assign n34713 = n7050 | n32106 ;
  assign n34715 = n34714 ^ n34713 ^ 1'b0 ;
  assign n34716 = n21080 & ~n27219 ;
  assign n34717 = n28803 ^ n28295 ^ n6943 ;
  assign n34718 = n25407 & n25565 ;
  assign n34719 = n7975 | n11681 ;
  assign n34720 = n11046 & ~n13230 ;
  assign n34721 = ~n34719 & n34720 ;
  assign n34722 = n27269 ^ n765 ^ 1'b0 ;
  assign n34723 = n2576 & n11747 ;
  assign n34724 = n860 | n34723 ;
  assign n34725 = n34724 ^ n31429 ^ 1'b0 ;
  assign n34726 = n5940 & n34325 ;
  assign n34727 = n6869 | n11102 ;
  assign n34728 = n34726 | n34727 ;
  assign n34729 = n19716 ^ n6797 ^ 1'b0 ;
  assign n34730 = n34729 ^ n7538 ^ 1'b0 ;
  assign n34731 = n148 | n13603 ;
  assign n34732 = n11315 | n34731 ;
  assign n34733 = n28537 ^ n4852 ^ 1'b0 ;
  assign n34734 = n14184 ^ n3315 ^ 1'b0 ;
  assign n34735 = n5866 & ~n13383 ;
  assign n34736 = ( n1902 & n15660 ) | ( n1902 & ~n22354 ) | ( n15660 & ~n22354 ) ;
  assign n34737 = ~n2853 & n28999 ;
  assign n34738 = n34737 ^ n27466 ^ 1'b0 ;
  assign n34739 = n14351 & n21814 ;
  assign n34740 = n30704 & ~n34739 ;
  assign n34741 = n34740 ^ n1116 ^ 1'b0 ;
  assign n34742 = ~n2852 & n11466 ;
  assign n34743 = n34742 ^ n3861 ^ 1'b0 ;
  assign n34744 = n3556 & n34743 ;
  assign n34745 = n34744 ^ n30175 ^ 1'b0 ;
  assign n34746 = n20044 ^ n17903 ^ n15841 ;
  assign n34747 = n20367 ^ n2728 ^ 1'b0 ;
  assign n34748 = n10120 & n13342 ;
  assign n34749 = ( ~n1568 & n3338 ) | ( ~n1568 & n22226 ) | ( n3338 & n22226 ) ;
  assign n34750 = ~n9354 & n20946 ;
  assign n34751 = ~n9213 & n34750 ;
  assign n34752 = n34749 | n34751 ;
  assign n34753 = n620 & ~n10702 ;
  assign n34754 = n7075 | n34753 ;
  assign n34755 = n33689 | n34754 ;
  assign n34756 = ~n11314 & n17427 ;
  assign n34757 = n5380 ^ n1237 ^ 1'b0 ;
  assign n34758 = ( n5425 & n24895 ) | ( n5425 & ~n25085 ) | ( n24895 & ~n25085 ) ;
  assign n34759 = n564 | n15193 ;
  assign n34760 = n571 | n34759 ;
  assign n34761 = ~n12363 & n34760 ;
  assign n34762 = n22314 & n34761 ;
  assign n34763 = n559 & ~n19888 ;
  assign n34764 = n1172 & ~n2855 ;
  assign n34765 = n1467 | n34764 ;
  assign n34766 = n592 ^ n552 ^ 1'b0 ;
  assign n34767 = n6974 & ~n9385 ;
  assign n34768 = n34766 & n34767 ;
  assign n34769 = n14694 & n25566 ;
  assign n34770 = n34769 ^ n8425 ^ 1'b0 ;
  assign n34771 = ~n5380 & n34770 ;
  assign n34772 = ~n699 & n2474 ;
  assign n34773 = n34772 ^ n10040 ^ 1'b0 ;
  assign n34774 = n14369 ^ n13477 ^ 1'b0 ;
  assign n34775 = ~n10527 & n13432 ;
  assign n34776 = n6615 | n32921 ;
  assign n34777 = n34776 ^ n386 ^ 1'b0 ;
  assign n34778 = ( n3961 & n13322 ) | ( n3961 & n34777 ) | ( n13322 & n34777 ) ;
  assign n34780 = n2856 | n9058 ;
  assign n34781 = n34780 ^ n3044 ^ 1'b0 ;
  assign n34779 = n286 & ~n31087 ;
  assign n34782 = n34781 ^ n34779 ^ 1'b0 ;
  assign n34783 = ( n8492 & ~n18421 ) | ( n8492 & n34782 ) | ( ~n18421 & n34782 ) ;
  assign n34784 = ~n25604 & n34783 ;
  assign n34785 = n1889 | n34282 ;
  assign n34786 = n5269 | n9047 ;
  assign n34787 = n13868 ^ n11876 ^ 1'b0 ;
  assign n34788 = n32990 | n34787 ;
  assign n34789 = n23641 & ~n34788 ;
  assign n34790 = n1269 & n34789 ;
  assign n34791 = n4365 | n28372 ;
  assign n34792 = n34791 ^ n31398 ^ 1'b0 ;
  assign n34793 = n34790 | n34792 ;
  assign n34794 = ( n1276 & n6885 ) | ( n1276 & ~n7616 ) | ( n6885 & ~n7616 ) ;
  assign n34795 = n34794 ^ n10819 ^ 1'b0 ;
  assign n34796 = ~n1186 & n34795 ;
  assign n34797 = n9208 ^ n3600 ^ 1'b0 ;
  assign n34798 = n23619 ^ n15527 ^ n1029 ;
  assign n34799 = n34798 ^ n19900 ^ 1'b0 ;
  assign n34800 = n3325 & n15467 ;
  assign n34801 = n26627 ^ n15578 ^ 1'b0 ;
  assign n34802 = n363 & n30898 ;
  assign n34803 = n34802 ^ n13841 ^ 1'b0 ;
  assign n34804 = n6326 | n11882 ;
  assign n34805 = n34803 | n34804 ;
  assign n34806 = n25252 ^ n3388 ^ n2451 ;
  assign n34807 = n2489 & ~n9812 ;
  assign n34808 = ( n6416 & n32925 ) | ( n6416 & ~n34807 ) | ( n32925 & ~n34807 ) ;
  assign n34809 = n28395 ^ n24870 ^ 1'b0 ;
  assign n34810 = n20 & n31043 ;
  assign n34811 = n34810 ^ n4837 ^ 1'b0 ;
  assign n34812 = n14087 & ~n27790 ;
  assign n34814 = n13274 | n14229 ;
  assign n34815 = n13196 & ~n34814 ;
  assign n34816 = n19008 | n34815 ;
  assign n34813 = ~n2060 & n12228 ;
  assign n34817 = n34816 ^ n34813 ^ 1'b0 ;
  assign n34818 = ~n195 & n23797 ;
  assign n34819 = n4271 & ~n4670 ;
  assign n34820 = n798 | n34819 ;
  assign n34821 = n34818 | n34820 ;
  assign n34822 = ~n18999 & n34821 ;
  assign n34823 = ~n34821 & n34822 ;
  assign n34824 = n3580 & ~n19248 ;
  assign n34825 = ~n19924 & n28121 ;
  assign n34826 = n34825 ^ n924 ^ 1'b0 ;
  assign n34828 = n24311 ^ n8620 ^ 1'b0 ;
  assign n34827 = n13723 | n25316 ;
  assign n34829 = n34828 ^ n34827 ^ 1'b0 ;
  assign n34833 = n6475 & n17298 ;
  assign n34834 = n667 | n1201 ;
  assign n34835 = n1201 & ~n34834 ;
  assign n34836 = n765 & n34835 ;
  assign n34837 = n29140 & ~n34836 ;
  assign n34838 = ~n34833 & n34837 ;
  assign n34830 = n11724 | n19014 ;
  assign n34831 = n19014 & ~n34830 ;
  assign n34832 = n20535 | n34831 ;
  assign n34839 = n34838 ^ n34832 ^ 1'b0 ;
  assign n34840 = n23393 & n33969 ;
  assign n34841 = n34313 ^ n6966 ^ 1'b0 ;
  assign n34842 = n20577 | n34841 ;
  assign n34843 = n33076 ^ n26099 ^ n1995 ;
  assign n34844 = n5604 ^ n2856 ^ 1'b0 ;
  assign n34845 = n34844 ^ n2662 ^ n1758 ;
  assign n34846 = n8608 ^ n6056 ^ n5535 ;
  assign n34847 = n20442 & n31038 ;
  assign n34848 = ~n34846 & n34847 ;
  assign n34849 = n7609 & ~n25029 ;
  assign n34850 = ~n11556 & n34849 ;
  assign n34851 = ~n31943 & n34850 ;
  assign n34852 = n19741 ^ n18271 ^ n1257 ;
  assign n34853 = n34852 ^ n19094 ^ 1'b0 ;
  assign n34854 = n26436 ^ n17136 ^ 1'b0 ;
  assign n34855 = n17577 & n22710 ;
  assign n34856 = n34855 ^ n25385 ^ n7466 ;
  assign n34857 = n6600 | n32862 ;
  assign n34858 = n14593 | n15032 ;
  assign n34859 = n34858 ^ n17366 ^ 1'b0 ;
  assign n34860 = n3333 ^ n2918 ^ 1'b0 ;
  assign n34861 = ~n10638 & n34860 ;
  assign n34862 = n7379 & ~n18010 ;
  assign n34863 = n28714 & n34862 ;
  assign n34864 = n32798 ^ n22203 ^ n5270 ;
  assign n34865 = n14728 & ~n28230 ;
  assign n34866 = n22629 & n34865 ;
  assign n34868 = n942 | n4056 ;
  assign n34869 = n34868 ^ n6472 ^ 1'b0 ;
  assign n34867 = ~n11390 & n19961 ;
  assign n34870 = n34869 ^ n34867 ^ 1'b0 ;
  assign n34871 = ~n116 & n19603 ;
  assign n34872 = n34871 ^ n18675 ^ 1'b0 ;
  assign n34873 = n2318 & n34872 ;
  assign n34875 = n1307 & ~n4921 ;
  assign n34876 = n1658 & n34875 ;
  assign n34874 = n3797 | n3833 ;
  assign n34877 = n34876 ^ n34874 ^ 1'b0 ;
  assign n34878 = n14555 | n22099 ;
  assign n34879 = n30733 & n34878 ;
  assign n34880 = n25179 ^ n4770 ^ 1'b0 ;
  assign n34881 = n10886 & ~n34880 ;
  assign n34882 = n2515 & ~n25958 ;
  assign n34883 = n16145 ^ n11046 ^ 1'b0 ;
  assign n34884 = n1469 & ~n34883 ;
  assign n34885 = ~n13767 & n34884 ;
  assign n34886 = n15099 ^ n14371 ^ 1'b0 ;
  assign n34887 = n28866 | n34886 ;
  assign n34888 = n20801 ^ n12927 ^ 1'b0 ;
  assign n34889 = ~n4731 & n34888 ;
  assign n34890 = ( n11218 & n34099 ) | ( n11218 & n34889 ) | ( n34099 & n34889 ) ;
  assign n34891 = n34166 ^ n16990 ^ 1'b0 ;
  assign n34892 = ( ~n1207 & n4365 ) | ( ~n1207 & n32125 ) | ( n4365 & n32125 ) ;
  assign n34893 = ~n20266 & n34892 ;
  assign n34894 = n8401 & n9104 ;
  assign n34895 = ( n749 & n11021 ) | ( n749 & n34894 ) | ( n11021 & n34894 ) ;
  assign n34896 = n34895 ^ n19339 ^ 1'b0 ;
  assign n34897 = n40 & n1712 ;
  assign n34898 = ~n14221 & n34897 ;
  assign n34899 = n961 | n34898 ;
  assign n34900 = n5487 | n34899 ;
  assign n34901 = n12116 & ~n34900 ;
  assign n34902 = ~n1042 & n14673 ;
  assign n34903 = n34901 | n34902 ;
  assign n34904 = n5231 & ~n34903 ;
  assign n34905 = n6719 & ~n14327 ;
  assign n34906 = ~n2547 & n34905 ;
  assign n34907 = n3004 & n16208 ;
  assign n34908 = n34907 ^ n9546 ^ 1'b0 ;
  assign n34909 = ~n7369 & n19343 ;
  assign n34910 = ( n4429 & n7030 ) | ( n4429 & ~n34909 ) | ( n7030 & ~n34909 ) ;
  assign n34911 = n9077 & n12470 ;
  assign n34912 = n34911 ^ n6271 ^ 1'b0 ;
  assign n34913 = n25101 & n34912 ;
  assign n34914 = n34913 ^ n14485 ^ 1'b0 ;
  assign n34915 = n419 ^ n259 ^ 1'b0 ;
  assign n34916 = ~n3176 & n34915 ;
  assign n34917 = n12988 & n34916 ;
  assign n34918 = n34917 ^ n23805 ^ 1'b0 ;
  assign n34920 = n5025 & ~n20840 ;
  assign n34921 = n34920 ^ n32216 ^ 1'b0 ;
  assign n34919 = n2478 & ~n5667 ;
  assign n34922 = n34921 ^ n34919 ^ 1'b0 ;
  assign n34923 = n1150 & ~n15302 ;
  assign n34924 = n34923 ^ n1456 ^ 1'b0 ;
  assign n34925 = n34924 ^ n20726 ^ 1'b0 ;
  assign n34926 = n3687 | n14642 ;
  assign n34927 = n34925 & ~n34926 ;
  assign n34928 = n34927 ^ n1205 ^ 1'b0 ;
  assign n34929 = ~n3135 & n34928 ;
  assign n34930 = ~n22477 & n25608 ;
  assign n34931 = n372 & n34930 ;
  assign n34932 = n13002 | n34931 ;
  assign n34933 = n17760 ^ n5581 ^ 1'b0 ;
  assign n34934 = ~n9084 & n34933 ;
  assign n34935 = n24548 & n28054 ;
  assign n34936 = n4931 & ~n14381 ;
  assign n34937 = n34936 ^ n661 ^ 1'b0 ;
  assign n34938 = n14474 & ~n34937 ;
  assign n34939 = n34938 ^ n9768 ^ 1'b0 ;
  assign n34940 = n7865 & ~n14894 ;
  assign n34941 = n16920 ^ n7630 ^ 1'b0 ;
  assign n34942 = ~n34940 & n34941 ;
  assign n34943 = n532 & n1589 ;
  assign n34944 = ~n532 & n34943 ;
  assign n34945 = ~n10678 & n34944 ;
  assign n34946 = n34945 ^ n20641 ^ 1'b0 ;
  assign n34947 = n5163 | n7079 ;
  assign n34948 = n27756 | n34947 ;
  assign n34949 = n8607 & ~n34948 ;
  assign n34950 = n34946 | n34949 ;
  assign n34951 = n25546 | n34950 ;
  assign n34952 = n11225 ^ n474 ^ 1'b0 ;
  assign n34953 = ( n5393 & ~n10140 ) | ( n5393 & n34952 ) | ( ~n10140 & n34952 ) ;
  assign n34954 = n34953 ^ n33940 ^ n16621 ;
  assign n34955 = ~n15215 & n34954 ;
  assign n34956 = ~n9819 & n34955 ;
  assign n34957 = n944 | n7448 ;
  assign n34958 = n34957 ^ n4765 ^ 1'b0 ;
  assign n34959 = ( n968 & n2635 ) | ( n968 & n9046 ) | ( n2635 & n9046 ) ;
  assign n34960 = n14656 ^ n11189 ^ 1'b0 ;
  assign n34961 = n450 & n22094 ;
  assign n34962 = n13922 ^ n5149 ^ 1'b0 ;
  assign n34963 = ~n16218 & n34962 ;
  assign n34964 = n12849 & n34963 ;
  assign n34965 = n34961 & ~n34964 ;
  assign n34966 = n8331 & ~n16599 ;
  assign n34967 = n33911 & n34966 ;
  assign n34968 = ( n13083 & ~n13480 ) | ( n13083 & n34714 ) | ( ~n13480 & n34714 ) ;
  assign n34969 = n1231 & ~n5634 ;
  assign n34970 = ~n8338 & n32213 ;
  assign n34971 = ~n3805 & n34970 ;
  assign n34972 = n1631 & n5137 ;
  assign n34973 = n15646 ^ n11550 ^ 1'b0 ;
  assign n34974 = n15276 & ~n34973 ;
  assign n34975 = n14927 & n34974 ;
  assign n34976 = ~n2127 & n7656 ;
  assign n34977 = n9571 | n34976 ;
  assign n34978 = n1591 | n34977 ;
  assign n34979 = n5071 | n8850 ;
  assign n34980 = n34979 ^ n45 ^ 1'b0 ;
  assign n34981 = n527 & ~n13747 ;
  assign n34982 = ( ~n23066 & n25128 ) | ( ~n23066 & n34981 ) | ( n25128 & n34981 ) ;
  assign n34983 = n3261 ^ n2317 ^ n1409 ;
  assign n34984 = n7062 ^ n6081 ^ 1'b0 ;
  assign n34985 = n34983 | n34984 ;
  assign n34986 = n34985 ^ n29402 ^ 1'b0 ;
  assign n34987 = n27878 ^ n5528 ^ 1'b0 ;
  assign n34988 = n18040 ^ n1192 ^ 1'b0 ;
  assign n34989 = n21100 ^ n892 ^ 1'b0 ;
  assign n34990 = ~n14401 & n22110 ;
  assign n34991 = n3255 | n17760 ;
  assign n34992 = ~n373 & n8204 ;
  assign n34993 = n29716 & n34992 ;
  assign n34994 = n34993 ^ n15101 ^ 1'b0 ;
  assign n34995 = ( n5340 & n20662 ) | ( n5340 & n34952 ) | ( n20662 & n34952 ) ;
  assign n34996 = n9065 & ~n14963 ;
  assign n34997 = n10249 & n34996 ;
  assign n34998 = n28360 & n34997 ;
  assign n34999 = n34995 & n34998 ;
  assign n35000 = n15472 ^ n4436 ^ 1'b0 ;
  assign n35001 = ~n2900 & n35000 ;
  assign n35002 = n20657 ^ n14097 ^ n3818 ;
  assign n35003 = ~n35001 & n35002 ;
  assign n35004 = n6435 & n33382 ;
  assign n35005 = n15110 & n26987 ;
  assign n35006 = n35005 ^ n12826 ^ 1'b0 ;
  assign n35007 = ~n4313 & n35006 ;
  assign n35008 = n3995 ^ n878 ^ 1'b0 ;
  assign n35009 = n31412 | n34664 ;
  assign n35010 = n35009 ^ n2092 ^ 1'b0 ;
  assign n35013 = n17172 | n29385 ;
  assign n35011 = n1918 | n33262 ;
  assign n35012 = n6605 | n35011 ;
  assign n35014 = n35013 ^ n35012 ^ 1'b0 ;
  assign n35015 = n6084 | n14558 ;
  assign n35016 = ~n9631 & n13033 ;
  assign n35017 = n35016 ^ n30303 ^ n23817 ;
  assign n35018 = n27568 & ~n35013 ;
  assign n35019 = n4644 ^ n4095 ^ 1'b0 ;
  assign n35020 = n8898 & ~n35019 ;
  assign n35021 = n12800 ^ n1939 ^ 1'b0 ;
  assign n35022 = ~n16373 & n35021 ;
  assign n35023 = n12098 & n35022 ;
  assign n35024 = n15682 ^ n533 ^ 1'b0 ;
  assign n35025 = ~n10545 & n35024 ;
  assign n35026 = ~n35023 & n35025 ;
  assign n35027 = ~n26502 & n35026 ;
  assign n35028 = ~n2818 & n23256 ;
  assign n35029 = n35028 ^ n12204 ^ 1'b0 ;
  assign n35030 = n16346 ^ n8249 ^ n4583 ;
  assign n35031 = n28120 ^ n8145 ^ 1'b0 ;
  assign n35032 = n9274 & ~n28260 ;
  assign n35033 = n34786 ^ n509 ^ 1'b0 ;
  assign n35034 = n29925 ^ n9386 ^ 1'b0 ;
  assign n35035 = n16695 & n29497 ;
  assign n35036 = ~n2056 & n21271 ;
  assign n35037 = n1596 & ~n6919 ;
  assign n35038 = ~n30494 & n35037 ;
  assign n35039 = n5809 & ~n9360 ;
  assign n35040 = n35039 ^ n18073 ^ 1'b0 ;
  assign n35041 = ( n1726 & n4389 ) | ( n1726 & n35040 ) | ( n4389 & n35040 ) ;
  assign n35042 = n3875 ^ n1528 ^ 1'b0 ;
  assign n35043 = ~n12649 & n15433 ;
  assign n35044 = n590 & n35043 ;
  assign n35045 = n32811 ^ n11208 ^ 1'b0 ;
  assign n35046 = n7541 & n30105 ;
  assign n35047 = n10823 | n18654 ;
  assign n35048 = n35047 ^ n26130 ^ n3545 ;
  assign n35049 = n14303 & n28229 ;
  assign n35050 = n35049 ^ n19173 ^ 1'b0 ;
  assign n35051 = n7972 ^ n2637 ^ 1'b0 ;
  assign n35052 = n19189 & ~n35051 ;
  assign n35053 = ~n35050 & n35052 ;
  assign n35054 = n20940 & n25937 ;
  assign n35055 = ~n4425 & n6272 ;
  assign n35056 = n35055 ^ n27408 ^ 1'b0 ;
  assign n35059 = n4780 & ~n5893 ;
  assign n35060 = n11242 & n35059 ;
  assign n35057 = n16829 ^ n10157 ^ 1'b0 ;
  assign n35058 = n12740 & ~n35057 ;
  assign n35061 = n35060 ^ n35058 ^ 1'b0 ;
  assign n35062 = ( ~n8430 & n8809 ) | ( ~n8430 & n25201 ) | ( n8809 & n25201 ) ;
  assign n35063 = ~n325 & n35062 ;
  assign n35064 = n18572 & n35063 ;
  assign n35065 = ( n24157 & n26512 ) | ( n24157 & n35064 ) | ( n26512 & n35064 ) ;
  assign n35066 = n7918 ^ n7841 ^ 1'b0 ;
  assign n35067 = ~n5375 & n35066 ;
  assign n35068 = n24415 & ~n28295 ;
  assign n35069 = n28501 ^ n13687 ^ 1'b0 ;
  assign n35070 = n35068 | n35069 ;
  assign n35071 = n27147 ^ n25028 ^ 1'b0 ;
  assign n35072 = n9785 & ~n19283 ;
  assign n35073 = ~n3712 & n35072 ;
  assign n35074 = n35073 ^ n14428 ^ 1'b0 ;
  assign n35075 = ~n12860 & n35074 ;
  assign n35076 = n33239 ^ n12595 ^ 1'b0 ;
  assign n35077 = ~n431 & n35076 ;
  assign n35078 = n3647 | n35077 ;
  assign n35079 = ~n8992 & n12007 ;
  assign n35080 = ( ~n27150 & n32502 ) | ( ~n27150 & n35079 ) | ( n32502 & n35079 ) ;
  assign n35081 = n12950 | n29352 ;
  assign n35082 = n12548 ^ n11509 ^ n1701 ;
  assign n35085 = n25759 ^ n362 ^ 1'b0 ;
  assign n35083 = ( n317 & ~n4522 ) | ( n317 & n20453 ) | ( ~n4522 & n20453 ) ;
  assign n35084 = n19801 & n35083 ;
  assign n35086 = n35085 ^ n35084 ^ 1'b0 ;
  assign n35087 = n35082 & ~n35086 ;
  assign n35088 = n22257 & n35087 ;
  assign n35089 = ~n31879 & n33302 ;
  assign n35090 = n28725 ^ n3429 ^ 1'b0 ;
  assign n35091 = n33863 ^ n6560 ^ 1'b0 ;
  assign n35092 = n18009 & n35091 ;
  assign n35093 = n17407 ^ n7933 ^ 1'b0 ;
  assign n35094 = n16986 | n20573 ;
  assign n35095 = ~n15691 & n30916 ;
  assign n35097 = n27583 ^ n15103 ^ 1'b0 ;
  assign n35098 = ~n9837 & n35097 ;
  assign n35096 = n3392 & ~n6367 ;
  assign n35099 = n35098 ^ n35096 ^ 1'b0 ;
  assign n35100 = ~n22353 & n25370 ;
  assign n35102 = n936 & n4474 ;
  assign n35103 = n1933 & n35102 ;
  assign n35101 = n11234 & n11719 ;
  assign n35104 = n35103 ^ n35101 ^ 1'b0 ;
  assign n35105 = ~n11556 & n24543 ;
  assign n35106 = n26667 | n35105 ;
  assign n35107 = n10211 | n30539 ;
  assign n35108 = n21582 ^ n16405 ^ 1'b0 ;
  assign n35109 = n5510 & ~n35108 ;
  assign n35110 = ( ~n5309 & n21023 ) | ( ~n5309 & n35109 ) | ( n21023 & n35109 ) ;
  assign n35111 = n12665 ^ n9143 ^ n132 ;
  assign n35112 = n8201 ^ n3578 ^ n2429 ;
  assign n35113 = n35111 & ~n35112 ;
  assign n35114 = n35113 ^ n5916 ^ 1'b0 ;
  assign n35115 = ~n21559 & n35114 ;
  assign n35116 = n23124 & ~n27632 ;
  assign n35117 = ~n3939 & n11787 ;
  assign n35118 = n19380 ^ n1441 ^ 1'b0 ;
  assign n35119 = n13108 & ~n35118 ;
  assign n35120 = n35117 | n35119 ;
  assign n35121 = n20479 & n35120 ;
  assign n35122 = n6671 & n35121 ;
  assign n35123 = n747 | n2322 ;
  assign n35124 = n3685 & ~n35123 ;
  assign n35125 = n2056 ^ n2034 ^ 1'b0 ;
  assign n35126 = ~n35124 & n35125 ;
  assign n35127 = n13698 ^ n968 ^ 1'b0 ;
  assign n35128 = n765 & n35127 ;
  assign n35129 = n35128 ^ n25881 ^ 1'b0 ;
  assign n35130 = n35129 ^ n22187 ^ 1'b0 ;
  assign n35131 = n536 | n24044 ;
  assign n35132 = ~n18288 & n33097 ;
  assign n35133 = n35132 ^ n9215 ^ 1'b0 ;
  assign n35135 = n985 & n9673 ;
  assign n35136 = ~n21405 & n35135 ;
  assign n35134 = n13871 & ~n34253 ;
  assign n35137 = n35136 ^ n35134 ^ 1'b0 ;
  assign n35138 = ( n2130 & n2694 ) | ( n2130 & ~n4480 ) | ( n2694 & ~n4480 ) ;
  assign n35139 = n23767 ^ n58 ^ 1'b0 ;
  assign n35140 = n10642 & ~n35139 ;
  assign n35141 = n13613 & n35140 ;
  assign n35142 = n9483 & n35141 ;
  assign n35143 = n35142 ^ n31863 ^ n16004 ;
  assign n35144 = n10421 & n34259 ;
  assign n35145 = n9697 & n35144 ;
  assign n35146 = n15351 & n18845 ;
  assign n35147 = n23398 ^ n5651 ^ 1'b0 ;
  assign n35148 = n13618 | n35147 ;
  assign n35149 = n428 & n3374 ;
  assign n35150 = n35148 & n35149 ;
  assign n35151 = n35150 ^ n20255 ^ 1'b0 ;
  assign n35152 = n21586 ^ n14123 ^ 1'b0 ;
  assign n35153 = n30358 & n35152 ;
  assign n35154 = n35153 ^ n7361 ^ 1'b0 ;
  assign n35155 = n25671 ^ n23 ^ 1'b0 ;
  assign n35156 = n4430 & ~n35155 ;
  assign n35157 = n35156 ^ n8584 ^ 1'b0 ;
  assign n35158 = n32549 ^ n4479 ^ 1'b0 ;
  assign n35159 = n633 | n11147 ;
  assign n35160 = n35159 ^ n32922 ^ 1'b0 ;
  assign n35161 = ~n1714 & n12076 ;
  assign n35162 = n5719 ^ n1530 ^ 1'b0 ;
  assign n35163 = n13077 | n35162 ;
  assign n35164 = n35163 ^ n2732 ^ 1'b0 ;
  assign n35165 = ~n18167 & n35164 ;
  assign n35166 = n18621 ^ n7591 ^ 1'b0 ;
  assign n35167 = n9543 ^ n606 ^ 1'b0 ;
  assign n35168 = n2079 & ~n35167 ;
  assign n35169 = n35168 ^ n14227 ^ 1'b0 ;
  assign n35170 = n33750 ^ n14578 ^ 1'b0 ;
  assign n35171 = n9207 & ~n13436 ;
  assign n35172 = n16523 & n35171 ;
  assign n35173 = ~n6527 & n14474 ;
  assign n35174 = n24283 ^ n3774 ^ 1'b0 ;
  assign n35175 = n29582 ^ n18534 ^ 1'b0 ;
  assign n35176 = n31519 | n35175 ;
  assign n35177 = n15157 ^ n2217 ^ 1'b0 ;
  assign n35178 = n9630 | n12680 ;
  assign n35179 = n6539 & ~n35178 ;
  assign n35180 = n31489 ^ n30521 ^ 1'b0 ;
  assign n35181 = n16550 ^ n7948 ^ n1566 ;
  assign n35182 = n1745 & n12988 ;
  assign n35183 = n13370 & ~n35182 ;
  assign n35184 = n18717 ^ n17709 ^ 1'b0 ;
  assign n35185 = n4913 & ~n35184 ;
  assign n35191 = n9983 & n30113 ;
  assign n35192 = n35191 ^ n25143 ^ 1'b0 ;
  assign n35193 = ~n540 & n3833 ;
  assign n35194 = n35193 ^ n6271 ^ 1'b0 ;
  assign n35195 = ~n23203 & n35194 ;
  assign n35196 = n35192 & n35195 ;
  assign n35186 = n8977 | n28101 ;
  assign n35187 = ~n12211 & n19339 ;
  assign n35188 = n35187 ^ n14419 ^ 1'b0 ;
  assign n35189 = n19602 & ~n35188 ;
  assign n35190 = ~n35186 & n35189 ;
  assign n35197 = n35196 ^ n35190 ^ 1'b0 ;
  assign n35198 = n17056 & ~n23437 ;
  assign n35199 = ~n11425 & n35198 ;
  assign n35200 = n35199 ^ n15282 ^ n12453 ;
  assign n35201 = n16747 & n24906 ;
  assign n35202 = ~n20332 & n25929 ;
  assign n35203 = n28407 ^ n19542 ^ 1'b0 ;
  assign n35204 = n243 & n35203 ;
  assign n35205 = n270 | n30066 ;
  assign n35206 = n35205 ^ n22135 ^ 1'b0 ;
  assign n35207 = n12299 & n35206 ;
  assign n35209 = n33828 ^ n21676 ^ 1'b0 ;
  assign n35210 = n22575 & n35209 ;
  assign n35208 = n1525 & ~n13573 ;
  assign n35211 = n35210 ^ n35208 ^ 1'b0 ;
  assign n35212 = n5007 & n25501 ;
  assign n35213 = n17411 ^ n2978 ^ 1'b0 ;
  assign n35214 = n11914 | n35213 ;
  assign n35215 = n9775 | n15372 ;
  assign n35216 = ~n14542 & n16464 ;
  assign n35217 = n17901 & n35216 ;
  assign n35218 = n4236 & n20344 ;
  assign n35219 = n848 & n35218 ;
  assign n35220 = n1624 & ~n4442 ;
  assign n35221 = n7478 & ~n35220 ;
  assign n35222 = n32042 ^ n1355 ^ 1'b0 ;
  assign n35223 = ~n13526 & n35222 ;
  assign n35224 = n1501 | n16138 ;
  assign n35225 = n4034 & n12188 ;
  assign n35226 = n35225 ^ n10703 ^ 1'b0 ;
  assign n35227 = n5332 & ~n35226 ;
  assign n35228 = n35227 ^ n2602 ^ 1'b0 ;
  assign n35229 = n12123 ^ n9047 ^ 1'b0 ;
  assign n35230 = n25498 & n35229 ;
  assign n35231 = n35230 ^ n18293 ^ 1'b0 ;
  assign n35232 = n34959 ^ n924 ^ 1'b0 ;
  assign n35233 = n1718 & ~n35232 ;
  assign n35234 = n27225 ^ n12549 ^ 1'b0 ;
  assign n35235 = n30960 ^ n493 ^ 1'b0 ;
  assign n35236 = ~n9684 & n35235 ;
  assign n35237 = n5510 & n35236 ;
  assign n35238 = n3972 | n13393 ;
  assign n35239 = ( n2384 & n20379 ) | ( n2384 & ~n33024 ) | ( n20379 & ~n33024 ) ;
  assign n35240 = ~n2010 & n28785 ;
  assign n35241 = ~n34384 & n35240 ;
  assign n35242 = ~n6969 & n20092 ;
  assign n35243 = n35242 ^ n2443 ^ 1'b0 ;
  assign n35244 = n19050 | n29929 ;
  assign n35245 = n1016 & ~n1029 ;
  assign n35246 = n10857 & ~n35245 ;
  assign n35247 = n35246 ^ n3896 ^ 1'b0 ;
  assign n35248 = n14390 & ~n35247 ;
  assign n35249 = n17427 | n26794 ;
  assign n35250 = n16263 & ~n35249 ;
  assign n35251 = n35250 ^ n16312 ^ 1'b0 ;
  assign n35256 = n7245 | n12142 ;
  assign n35257 = n35256 ^ n667 ^ 1'b0 ;
  assign n35258 = n35257 ^ n10269 ^ 1'b0 ;
  assign n35252 = ~n5166 & n26318 ;
  assign n35253 = n35252 ^ n7842 ^ 1'b0 ;
  assign n35254 = n15239 & n35253 ;
  assign n35255 = n35254 ^ n29860 ^ 1'b0 ;
  assign n35259 = n35258 ^ n35255 ^ 1'b0 ;
  assign n35260 = n11485 ^ n11353 ^ 1'b0 ;
  assign n35261 = n28227 & ~n35260 ;
  assign n35262 = n35261 ^ n18621 ^ 1'b0 ;
  assign n35263 = n5311 ^ n342 ^ 1'b0 ;
  assign n35264 = ~n19423 & n35263 ;
  assign n35265 = n16478 ^ n6452 ^ 1'b0 ;
  assign n35266 = n3209 | n35265 ;
  assign n35267 = n35266 ^ n21042 ^ 1'b0 ;
  assign n35268 = ~n901 & n17528 ;
  assign n35269 = ~n15413 & n35268 ;
  assign n35270 = n6216 | n35269 ;
  assign n35271 = n25446 ^ n14871 ^ 1'b0 ;
  assign n35272 = ~n1580 & n13139 ;
  assign n35273 = n14603 ^ n13363 ^ 1'b0 ;
  assign n35274 = n4168 & ~n35273 ;
  assign n35275 = n18740 ^ n14677 ^ 1'b0 ;
  assign n35276 = n7494 & n35275 ;
  assign n35277 = ~n24580 & n35276 ;
  assign n35279 = n13947 & n25399 ;
  assign n35280 = n35279 ^ n11900 ^ 1'b0 ;
  assign n35281 = n9931 & n35280 ;
  assign n35282 = n35281 ^ n12758 ^ 1'b0 ;
  assign n35278 = n30041 ^ n10024 ^ 1'b0 ;
  assign n35283 = n35282 ^ n35278 ^ 1'b0 ;
  assign n35284 = n312 & ~n11147 ;
  assign n35285 = n35284 ^ n9639 ^ 1'b0 ;
  assign n35286 = n2912 & n35285 ;
  assign n35287 = ( n2125 & ~n25143 ) | ( n2125 & n35286 ) | ( ~n25143 & n35286 ) ;
  assign n35288 = n12264 ^ n10952 ^ 1'b0 ;
  assign n35289 = ~n8331 & n22105 ;
  assign n35290 = ~n4913 & n35289 ;
  assign n35291 = n10152 & ~n35290 ;
  assign n35292 = n35291 ^ n14498 ^ 1'b0 ;
  assign n35293 = n10239 & ~n10979 ;
  assign n35294 = n18046 | n35293 ;
  assign n35295 = n4070 & ~n9419 ;
  assign n35296 = n2522 | n27412 ;
  assign n35297 = n35295 | n35296 ;
  assign n35298 = n23219 & n35297 ;
  assign n35299 = n8387 ^ n1858 ^ 1'b0 ;
  assign n35300 = n13809 | n35299 ;
  assign n35301 = n7541 ^ n3745 ^ 1'b0 ;
  assign n35302 = ~n11232 & n35301 ;
  assign n35303 = n35300 | n35302 ;
  assign n35304 = n26697 ^ n25704 ^ n6304 ;
  assign n35305 = n11676 & n13934 ;
  assign n35306 = n35305 ^ n7948 ^ 1'b0 ;
  assign n35307 = ~n19247 & n35306 ;
  assign n35308 = n35307 ^ n16600 ^ 1'b0 ;
  assign n35309 = n530 & n12090 ;
  assign n35310 = n625 & n35309 ;
  assign n35311 = n35310 ^ n2489 ^ 1'b0 ;
  assign n35312 = n35311 ^ n4857 ^ 1'b0 ;
  assign n35313 = n35308 | n35312 ;
  assign n35314 = n7871 & n10656 ;
  assign n35315 = n18958 & n35314 ;
  assign n35316 = n6236 ^ n1734 ^ 1'b0 ;
  assign n35317 = n35316 ^ n10121 ^ 1'b0 ;
  assign n35318 = n35315 | n35317 ;
  assign n35319 = n323 & ~n5113 ;
  assign n35320 = n7430 ^ n3663 ^ 1'b0 ;
  assign n35321 = n35320 ^ n22068 ^ 1'b0 ;
  assign n35322 = n35032 ^ n9050 ^ n4910 ;
  assign n35323 = ( n12375 & n12432 ) | ( n12375 & n17964 ) | ( n12432 & n17964 ) ;
  assign n35324 = n27929 ^ n26052 ^ 1'b0 ;
  assign n35325 = ~n4021 & n35324 ;
  assign n35326 = n13996 | n18571 ;
  assign n35328 = n3319 | n29325 ;
  assign n35329 = n35328 ^ n11697 ^ 1'b0 ;
  assign n35327 = n780 | n16517 ;
  assign n35330 = n35329 ^ n35327 ^ 1'b0 ;
  assign n35331 = n25933 & ~n33572 ;
  assign n35334 = ~n2421 & n12040 ;
  assign n35332 = n7033 | n7550 ;
  assign n35333 = n35332 ^ n33577 ^ 1'b0 ;
  assign n35335 = n35334 ^ n35333 ^ n6091 ;
  assign n35336 = n7189 & ~n35335 ;
  assign n35337 = n35336 ^ n5458 ^ 1'b0 ;
  assign n35338 = ~n1864 & n4666 ;
  assign n35339 = n35338 ^ n9721 ^ 1'b0 ;
  assign n35340 = n4233 | n10073 ;
  assign n35341 = ~n35339 & n35340 ;
  assign n35342 = n5999 ^ n2754 ^ 1'b0 ;
  assign n35343 = n18169 & n35342 ;
  assign n35344 = ~n35341 & n35343 ;
  assign n35345 = n20869 ^ n6252 ^ 1'b0 ;
  assign n35346 = ( n11340 & n16988 ) | ( n11340 & ~n31925 ) | ( n16988 & ~n31925 ) ;
  assign n35347 = n11391 & n35346 ;
  assign n35348 = n17561 | n20255 ;
  assign n35349 = n35348 ^ n5935 ^ 1'b0 ;
  assign n35352 = n20272 ^ n11710 ^ n8315 ;
  assign n35353 = n3259 & ~n35352 ;
  assign n35350 = n28017 ^ n9049 ^ n1613 ;
  assign n35351 = n35350 ^ n16719 ^ n6626 ;
  assign n35354 = n35353 ^ n35351 ^ n25262 ;
  assign n35355 = n3233 & ~n31153 ;
  assign n35356 = n4555 & n31961 ;
  assign n35357 = ~n14821 & n35356 ;
  assign n35358 = n35355 & ~n35357 ;
  assign n35359 = n35358 ^ n10536 ^ 1'b0 ;
  assign n35360 = ( n6758 & ~n27732 ) | ( n6758 & n35359 ) | ( ~n27732 & n35359 ) ;
  assign n35361 = n6124 | n15071 ;
  assign n35362 = n35361 ^ n7437 ^ 1'b0 ;
  assign n35363 = n18412 ^ n14558 ^ 1'b0 ;
  assign n35364 = ~n184 & n35363 ;
  assign n35365 = n10796 | n24131 ;
  assign n35366 = ~n6100 & n11334 ;
  assign n35367 = n4333 & n35366 ;
  assign n35368 = ~n25626 & n35367 ;
  assign n35369 = n17881 ^ n7699 ^ 1'b0 ;
  assign n35370 = n35369 ^ n21256 ^ 1'b0 ;
  assign n35371 = n11346 & n35370 ;
  assign n35372 = n11458 ^ n7254 ^ 1'b0 ;
  assign n35373 = n35371 & ~n35372 ;
  assign n35374 = n3962 ^ n379 ^ 1'b0 ;
  assign n35375 = ~n163 & n7390 ;
  assign n35376 = n21253 ^ n16156 ^ 1'b0 ;
  assign n35377 = ~n35375 & n35376 ;
  assign n35378 = ~n1312 & n35377 ;
  assign n35379 = ~n16790 & n35378 ;
  assign n35380 = ~n12523 & n33365 ;
  assign n35381 = n23203 | n35380 ;
  assign n35382 = n30178 & ~n35381 ;
  assign n35383 = ~n3280 & n10970 ;
  assign n35384 = n33891 | n35383 ;
  assign n35385 = n35384 ^ n29689 ^ 1'b0 ;
  assign n35388 = n1416 & n1969 ;
  assign n35389 = n35388 ^ n28138 ^ 1'b0 ;
  assign n35386 = n10324 | n23061 ;
  assign n35387 = n468 & ~n35386 ;
  assign n35390 = n35389 ^ n35387 ^ 1'b0 ;
  assign n35391 = n2336 & ~n13444 ;
  assign n35392 = ~n11404 & n35391 ;
  assign n35393 = ~n1392 & n32408 ;
  assign n35394 = ~n9002 & n35393 ;
  assign n35395 = n26390 | n30210 ;
  assign n35396 = n35395 ^ n8462 ^ 1'b0 ;
  assign n35397 = n9207 ^ n5623 ^ 1'b0 ;
  assign n35398 = ( n9949 & n14937 ) | ( n9949 & ~n35397 ) | ( n14937 & ~n35397 ) ;
  assign n35399 = ( n1845 & n13893 ) | ( n1845 & ~n16683 ) | ( n13893 & ~n16683 ) ;
  assign n35400 = n35399 ^ n1157 ^ 1'b0 ;
  assign n35401 = n4622 | n35400 ;
  assign n35402 = n17760 | n18385 ;
  assign n35403 = n13124 & ~n35402 ;
  assign n35404 = ~n26137 & n30210 ;
  assign n35405 = n23363 & n35404 ;
  assign n35406 = n4782 | n5052 ;
  assign n35407 = n20997 & ~n35406 ;
  assign n35408 = n35405 | n35407 ;
  assign n35409 = n1191 & ~n28154 ;
  assign n35410 = ~n9192 & n35409 ;
  assign n35411 = ~n24799 & n35410 ;
  assign n35412 = n2103 ^ n1816 ^ n124 ;
  assign n35413 = n439 & n35412 ;
  assign n35414 = n35413 ^ n25537 ^ 1'b0 ;
  assign n35415 = n32823 ^ n16057 ^ 1'b0 ;
  assign n35416 = n35414 | n35415 ;
  assign n35417 = n34599 ^ n33740 ^ 1'b0 ;
  assign n35418 = n8355 | n35417 ;
  assign n35419 = n1918 ^ n1044 ^ 1'b0 ;
  assign n35420 = ( n676 & n14460 ) | ( n676 & ~n35419 ) | ( n14460 & ~n35419 ) ;
  assign n35421 = n17259 ^ n11498 ^ 1'b0 ;
  assign n35422 = n35420 & ~n35421 ;
  assign n35423 = ~n32540 & n34694 ;
  assign n35424 = ~n3045 & n25261 ;
  assign n35425 = n7483 ^ n3437 ^ 1'b0 ;
  assign n35426 = n1161 & n35425 ;
  assign n35427 = n35426 ^ n28070 ^ 1'b0 ;
  assign n35428 = n35427 ^ n16777 ^ 1'b0 ;
  assign n35429 = n8000 ^ n3111 ^ 1'b0 ;
  assign n35430 = n4729 & n9772 ;
  assign n35431 = n35430 ^ n8005 ^ 1'b0 ;
  assign n35432 = n35429 | n35431 ;
  assign n35433 = ~n20341 & n35432 ;
  assign n35434 = n13380 ^ n152 ^ 1'b0 ;
  assign n35435 = n2440 & n35434 ;
  assign n35436 = n9917 & ~n12474 ;
  assign n35437 = ~n22634 & n32154 ;
  assign n35438 = n11872 ^ n6372 ^ 1'b0 ;
  assign n35439 = n1569 & n35438 ;
  assign n35440 = n18929 ^ n17441 ^ 1'b0 ;
  assign n35441 = n27727 ^ n1023 ^ 1'b0 ;
  assign n35442 = n18616 & ~n35441 ;
  assign n35443 = n35442 ^ n2711 ^ 1'b0 ;
  assign n35444 = n5431 | n31832 ;
  assign n35445 = n15527 & ~n35444 ;
  assign n35446 = n26473 ^ n4301 ^ 1'b0 ;
  assign n35447 = n7518 ^ n4960 ^ 1'b0 ;
  assign n35449 = n5350 ^ n4182 ^ n56 ;
  assign n35448 = n10195 | n30838 ;
  assign n35450 = n35449 ^ n35448 ^ 1'b0 ;
  assign n35451 = n29353 ^ n4707 ^ 1'b0 ;
  assign n35452 = n7862 ^ n1829 ^ 1'b0 ;
  assign n35453 = ~n13287 & n35452 ;
  assign n35454 = n8173 & n35453 ;
  assign n35455 = ( ~n1479 & n2045 ) | ( ~n1479 & n2859 ) | ( n2045 & n2859 ) ;
  assign n35456 = n35455 ^ n4451 ^ 1'b0 ;
  assign n35457 = ( n17492 & n35454 ) | ( n17492 & n35456 ) | ( n35454 & n35456 ) ;
  assign n35458 = n16669 ^ n12007 ^ 1'b0 ;
  assign n35459 = n13283 | n35458 ;
  assign n35460 = n35459 ^ n9534 ^ 1'b0 ;
  assign n35461 = ~n21131 & n35460 ;
  assign n35462 = n35461 ^ n6988 ^ 1'b0 ;
  assign n35463 = n13218 | n34386 ;
  assign n35464 = n35463 ^ n18605 ^ 1'b0 ;
  assign n35465 = n12692 & ~n23817 ;
  assign n35466 = n35465 ^ n5188 ^ 1'b0 ;
  assign n35469 = n2829 & n23065 ;
  assign n35467 = ~n13920 & n14052 ;
  assign n35468 = n35467 ^ n8829 ^ 1'b0 ;
  assign n35470 = n35469 ^ n35468 ^ n10831 ;
  assign n35471 = n35470 ^ n25188 ^ 1'b0 ;
  assign n35472 = n23810 & ~n35471 ;
  assign n35473 = ( n6854 & ~n9372 ) | ( n6854 & n12271 ) | ( ~n9372 & n12271 ) ;
  assign n35474 = n11409 ^ n1653 ^ 1'b0 ;
  assign n35475 = n35473 | n35474 ;
  assign n35476 = n2697 | n8089 ;
  assign n35477 = n35475 | n35476 ;
  assign n35478 = n28762 ^ n7298 ^ 1'b0 ;
  assign n35479 = ~n262 & n35478 ;
  assign n35480 = n9940 | n17974 ;
  assign n35481 = ~n23555 & n30036 ;
  assign n35482 = ~n11839 & n35481 ;
  assign n35483 = n7257 ^ n3295 ^ n1157 ;
  assign n35484 = n17383 & n35483 ;
  assign n35485 = n35484 ^ n7884 ^ 1'b0 ;
  assign n35486 = n16745 & ~n26126 ;
  assign n35487 = n33016 ^ n30725 ^ 1'b0 ;
  assign n35488 = ~n5493 & n19710 ;
  assign n35489 = n11068 & ~n35488 ;
  assign n35490 = n35489 ^ n318 ^ 1'b0 ;
  assign n35491 = n18941 | n22558 ;
  assign n35492 = n8267 | n23093 ;
  assign n35493 = n11837 ^ n4087 ^ 1'b0 ;
  assign n35494 = n3520 | n35493 ;
  assign n35495 = n35494 ^ n4848 ^ 1'b0 ;
  assign n35496 = n14601 ^ n8144 ^ 1'b0 ;
  assign n35497 = ~n6694 & n35496 ;
  assign n35498 = ( n1329 & ~n21473 ) | ( n1329 & n35497 ) | ( ~n21473 & n35497 ) ;
  assign n35499 = n9437 & n20521 ;
  assign n35500 = n35499 ^ n22720 ^ 1'b0 ;
  assign n35503 = n17350 ^ n6041 ^ 1'b0 ;
  assign n35504 = n4083 & ~n35503 ;
  assign n35505 = n35504 ^ n13891 ^ 1'b0 ;
  assign n35506 = n35483 & ~n35505 ;
  assign n35507 = ~n8495 & n35506 ;
  assign n35501 = ~n14458 & n16236 ;
  assign n35502 = n4367 & n35501 ;
  assign n35508 = n35507 ^ n35502 ^ 1'b0 ;
  assign n35509 = n7473 ^ n5282 ^ 1'b0 ;
  assign n35510 = n1768 ^ n1142 ^ 1'b0 ;
  assign n35511 = n10620 & ~n20207 ;
  assign n35512 = ~n35510 & n35511 ;
  assign n35513 = n30433 ^ n20294 ^ 1'b0 ;
  assign n35514 = ~n12655 & n35513 ;
  assign n35515 = n31301 ^ n21176 ^ 1'b0 ;
  assign n35516 = n9386 & n35515 ;
  assign n35517 = n35516 ^ n18573 ^ 1'b0 ;
  assign n35518 = n257 | n10953 ;
  assign n35519 = n22112 | n35518 ;
  assign n35520 = n17887 ^ n1422 ^ 1'b0 ;
  assign n35521 = n8014 & n35520 ;
  assign n35522 = ~n11409 & n22520 ;
  assign n35523 = ~n32510 & n35522 ;
  assign n35524 = ~n6304 & n14031 ;
  assign n35525 = n5936 & n35524 ;
  assign n35526 = n35525 ^ n33087 ^ n12422 ;
  assign n35528 = n5809 | n27698 ;
  assign n35527 = n2300 & n3995 ;
  assign n35529 = n35528 ^ n35527 ^ 1'b0 ;
  assign n35530 = ~n33940 & n35529 ;
  assign n35531 = n35530 ^ n17153 ^ 1'b0 ;
  assign n35532 = n3500 & n21463 ;
  assign n35536 = n5490 & ~n35389 ;
  assign n35533 = ~n9684 & n25008 ;
  assign n35534 = n18292 & n35533 ;
  assign n35535 = n27 | n35534 ;
  assign n35537 = n35536 ^ n35535 ^ 1'b0 ;
  assign n35538 = n13523 | n35537 ;
  assign n35539 = n35538 ^ n17120 ^ 1'b0 ;
  assign n35540 = n1863 & n24454 ;
  assign n35541 = n35540 ^ n11018 ^ 1'b0 ;
  assign n35542 = n31048 | n35541 ;
  assign n35543 = n35542 ^ n14340 ^ 1'b0 ;
  assign n35544 = ~n15935 & n35543 ;
  assign n35545 = n8553 ^ n5915 ^ 1'b0 ;
  assign n35546 = ~n17142 & n35545 ;
  assign n35547 = n16940 ^ n8042 ^ 1'b0 ;
  assign n35548 = n4369 & n35547 ;
  assign n35549 = n14251 ^ n5349 ^ 1'b0 ;
  assign n35550 = n3188 & ~n8445 ;
  assign n35551 = n13352 & n35550 ;
  assign n35552 = n35551 ^ n30899 ^ n10361 ;
  assign n35553 = n7487 ^ n1003 ^ 1'b0 ;
  assign n35554 = n4477 | n35553 ;
  assign n35555 = n35554 ^ n7918 ^ 1'b0 ;
  assign n35556 = ~n9507 & n16896 ;
  assign n35557 = n18828 & n35556 ;
  assign n35558 = n593 | n3414 ;
  assign n35559 = n7399 | n35558 ;
  assign n35560 = n35559 ^ n25439 ^ 1'b0 ;
  assign n35561 = n21512 & n35560 ;
  assign n35564 = n349 & ~n28605 ;
  assign n35565 = n35564 ^ n21880 ^ 1'b0 ;
  assign n35562 = n11800 ^ n9264 ^ n8194 ;
  assign n35563 = ~n4094 & n35562 ;
  assign n35566 = n35565 ^ n35563 ^ 1'b0 ;
  assign n35567 = n35566 ^ n9296 ^ n2971 ;
  assign n35568 = n11374 & n35567 ;
  assign n35569 = n15421 & ~n35568 ;
  assign n35570 = n11421 | n30349 ;
  assign n35571 = n9216 | n35570 ;
  assign n35572 = n30292 ^ n9941 ^ 1'b0 ;
  assign n35573 = n35571 & n35572 ;
  assign n35574 = n35573 ^ n34821 ^ 1'b0 ;
  assign n35575 = n16857 | n29387 ;
  assign n35576 = ~n3116 & n3897 ;
  assign n35577 = ~n3802 & n35576 ;
  assign n35578 = n7086 ^ n3877 ^ 1'b0 ;
  assign n35579 = n2723 & ~n35578 ;
  assign n35580 = n15923 ^ n144 ^ 1'b0 ;
  assign n35581 = n6647 | n35580 ;
  assign n35582 = n8267 & ~n35581 ;
  assign n35583 = ~n35579 & n35582 ;
  assign n35584 = ~n2460 & n5974 ;
  assign n35585 = n697 & n35584 ;
  assign n35586 = n35585 ^ n663 ^ 1'b0 ;
  assign n35587 = ~n10935 & n35586 ;
  assign n35588 = ( n2079 & n7893 ) | ( n2079 & n8081 ) | ( n7893 & n8081 ) ;
  assign n35589 = n35588 ^ n10352 ^ 1'b0 ;
  assign n35590 = ( n15333 & n24853 ) | ( n15333 & n35589 ) | ( n24853 & n35589 ) ;
  assign n35591 = n18017 & n35590 ;
  assign n35597 = n14624 ^ n9048 ^ 1'b0 ;
  assign n35594 = ( ~n14580 & n21130 ) | ( ~n14580 & n24492 ) | ( n21130 & n24492 ) ;
  assign n35595 = n35594 ^ n1291 ^ 1'b0 ;
  assign n35593 = n16994 ^ n12314 ^ 1'b0 ;
  assign n35596 = n35595 ^ n35593 ^ 1'b0 ;
  assign n35598 = n35597 ^ n35596 ^ 1'b0 ;
  assign n35599 = ~n25529 & n35598 ;
  assign n35592 = n30368 & n31459 ;
  assign n35600 = n35599 ^ n35592 ^ 1'b0 ;
  assign n35601 = n18964 & n35194 ;
  assign n35602 = n14471 & ~n16781 ;
  assign n35603 = n35602 ^ n18635 ^ 1'b0 ;
  assign n35604 = n28397 & ~n35603 ;
  assign n35605 = n16513 ^ n14942 ^ 1'b0 ;
  assign n35606 = n11547 & ~n13544 ;
  assign n35607 = n35606 ^ n12597 ^ 1'b0 ;
  assign n35608 = n27117 | n35607 ;
  assign n35609 = n18142 | n35608 ;
  assign n35610 = n35609 ^ n23270 ^ 1'b0 ;
  assign n35611 = ~n35605 & n35610 ;
  assign n35612 = n9797 ^ n3009 ^ 1'b0 ;
  assign n35614 = ~n2645 & n32665 ;
  assign n35613 = n1814 & ~n30569 ;
  assign n35615 = n35614 ^ n35613 ^ 1'b0 ;
  assign n35616 = n31898 ^ n11668 ^ 1'b0 ;
  assign n35617 = n17637 & ~n35616 ;
  assign n35618 = ~n9277 & n9611 ;
  assign n35619 = n5525 & ~n35618 ;
  assign n35620 = ~n35617 & n35619 ;
  assign n35621 = n1372 | n13564 ;
  assign n35622 = n14750 | n35621 ;
  assign n35623 = ~n4070 & n8529 ;
  assign n35624 = n18603 | n35623 ;
  assign n35625 = n33951 | n35624 ;
  assign n35626 = n14978 & n35625 ;
  assign n35627 = ~n33127 & n35626 ;
  assign n35628 = n5727 | n6923 ;
  assign n35630 = n2749 & n20168 ;
  assign n35629 = n13324 | n15261 ;
  assign n35631 = n35630 ^ n35629 ^ 1'b0 ;
  assign n35632 = n18641 ^ n9832 ^ 1'b0 ;
  assign n35633 = n1617 & n35632 ;
  assign n35634 = n35633 ^ n3505 ^ 1'b0 ;
  assign n35635 = n35631 | n35634 ;
  assign n35636 = n35635 ^ n33391 ^ 1'b0 ;
  assign n35637 = n9850 ^ n5467 ^ 1'b0 ;
  assign n35638 = n13855 | n35637 ;
  assign n35639 = n10477 & ~n35638 ;
  assign n35640 = n10438 ^ n737 ^ 1'b0 ;
  assign n35641 = ( ~n13919 & n22793 ) | ( ~n13919 & n35640 ) | ( n22793 & n35640 ) ;
  assign n35642 = n5364 ^ n2940 ^ 1'b0 ;
  assign n35643 = n26299 | n35642 ;
  assign n35644 = n4624 & n29250 ;
  assign n35645 = ~n1939 & n7164 ;
  assign n35646 = n28241 & n35645 ;
  assign n35647 = n6257 & n8012 ;
  assign n35648 = n12214 ^ n2970 ^ 1'b0 ;
  assign n35649 = n9104 & ~n10056 ;
  assign n35650 = n7202 & n35649 ;
  assign n35651 = ( ~n3165 & n35648 ) | ( ~n3165 & n35650 ) | ( n35648 & n35650 ) ;
  assign n35652 = n7699 & ~n22272 ;
  assign n35653 = n18186 | n35652 ;
  assign n35654 = ~n16042 & n34153 ;
  assign n35655 = ~n35653 & n35654 ;
  assign n35656 = n2460 | n24875 ;
  assign n35657 = n8187 | n30107 ;
  assign n35658 = n35656 & ~n35657 ;
  assign n35659 = ~n9912 & n22153 ;
  assign n35660 = ~n27591 & n35659 ;
  assign n35661 = n10929 ^ n8212 ^ 1'b0 ;
  assign n35662 = n24543 & ~n35661 ;
  assign n35664 = n17700 ^ n1971 ^ 1'b0 ;
  assign n35665 = n18898 & n35664 ;
  assign n35663 = n13926 & ~n17239 ;
  assign n35666 = n35665 ^ n35663 ^ 1'b0 ;
  assign n35667 = n10919 | n35666 ;
  assign n35668 = n17781 ^ n5126 ^ 1'b0 ;
  assign n35669 = n19408 ^ n16721 ^ 1'b0 ;
  assign n35670 = n9749 & n35669 ;
  assign n35671 = n34236 ^ n24102 ^ 1'b0 ;
  assign n35672 = n19210 ^ n11292 ^ 1'b0 ;
  assign n35673 = n12199 & ~n14466 ;
  assign n35674 = ( n2639 & n16940 ) | ( n2639 & n27524 ) | ( n16940 & n27524 ) ;
  assign n35675 = n35674 ^ n15557 ^ 1'b0 ;
  assign n35676 = n1286 & n17136 ;
  assign n35677 = n10967 ^ n6658 ^ 1'b0 ;
  assign n35678 = n35676 & n35677 ;
  assign n35679 = n16497 & ~n27459 ;
  assign n35680 = n20809 ^ n6751 ^ 1'b0 ;
  assign n35681 = n22579 & n35680 ;
  assign n35682 = n12863 ^ n777 ^ 1'b0 ;
  assign n35683 = ( n4065 & n14564 ) | ( n4065 & n28171 ) | ( n14564 & n28171 ) ;
  assign n35684 = n22854 & ~n35683 ;
  assign n35685 = ~n7877 & n35684 ;
  assign n35686 = n14341 | n26967 ;
  assign n35687 = n19588 ^ n15075 ^ 1'b0 ;
  assign n35688 = n15252 | n21059 ;
  assign n35689 = n35687 & ~n35688 ;
  assign n35690 = n1781 | n3592 ;
  assign n35691 = ~n378 & n35690 ;
  assign n35692 = n3428 | n24491 ;
  assign n35693 = n35691 | n35692 ;
  assign n35694 = n30661 ^ n3139 ^ 1'b0 ;
  assign n35695 = n530 & ~n35694 ;
  assign n35696 = ~n6719 & n35695 ;
  assign n35697 = n28482 ^ n6228 ^ n3374 ;
  assign n35698 = n4276 | n35697 ;
  assign n35699 = n6578 ^ n5089 ^ 1'b0 ;
  assign n35700 = n35699 ^ n26995 ^ 1'b0 ;
  assign n35701 = n6366 & ~n35700 ;
  assign n35702 = n33712 ^ n9858 ^ 1'b0 ;
  assign n35703 = n16986 & n35702 ;
  assign n35704 = ~n11942 & n16770 ;
  assign n35705 = n35704 ^ n33019 ^ 1'b0 ;
  assign n35706 = ~n6832 & n8491 ;
  assign n35707 = n35706 ^ n30904 ^ 1'b0 ;
  assign n35708 = n12776 | n35707 ;
  assign n35709 = n7722 & ~n27019 ;
  assign n35710 = n35709 ^ n32642 ^ 1'b0 ;
  assign n35711 = n7963 ^ n1686 ^ 1'b0 ;
  assign n35712 = n2146 | n35711 ;
  assign n35713 = n6250 & ~n35712 ;
  assign n35714 = ~n35710 & n35713 ;
  assign n35715 = n5459 | n15122 ;
  assign n35716 = n35715 ^ n21743 ^ 1'b0 ;
  assign n35717 = n10298 & n14295 ;
  assign n35718 = ~n25759 & n35717 ;
  assign n35719 = ~n6818 & n10115 ;
  assign n35720 = n4307 ^ n3193 ^ 1'b0 ;
  assign n35721 = n1761 & ~n35720 ;
  assign n35722 = n35721 ^ n4273 ^ 1'b0 ;
  assign n35723 = n35722 ^ n1210 ^ 1'b0 ;
  assign n35724 = n5741 ^ n2923 ^ 1'b0 ;
  assign n35725 = n2517 & ~n12877 ;
  assign n35726 = n35725 ^ n33924 ^ 1'b0 ;
  assign n35727 = n1617 & n26561 ;
  assign n35728 = n11202 | n27849 ;
  assign n35729 = n35728 ^ n29721 ^ 1'b0 ;
  assign n35730 = n8154 | n18856 ;
  assign n35731 = n35730 ^ n3037 ^ 1'b0 ;
  assign n35732 = n15795 & n26805 ;
  assign n35733 = n35732 ^ n30200 ^ 1'b0 ;
  assign n35734 = n35731 & n35733 ;
  assign n35735 = n35734 ^ n30732 ^ 1'b0 ;
  assign n35736 = n35735 ^ n16872 ^ 1'b0 ;
  assign n35737 = n18641 & ~n35736 ;
  assign n35738 = ~n25 & n345 ;
  assign n35739 = n3017 | n11167 ;
  assign n35740 = n25732 ^ n21061 ^ 1'b0 ;
  assign n35741 = ~n35739 & n35740 ;
  assign n35742 = n11897 & ~n21005 ;
  assign n35743 = ~n35741 & n35742 ;
  assign n35744 = n98 | n25075 ;
  assign n35745 = ( n7873 & n28183 ) | ( n7873 & ~n35744 ) | ( n28183 & ~n35744 ) ;
  assign n35746 = ~n29142 & n29842 ;
  assign n35747 = n35745 & n35746 ;
  assign n35748 = n24118 ^ n23324 ^ 1'b0 ;
  assign n35749 = n2306 & ~n35748 ;
  assign n35750 = n12763 & ~n21379 ;
  assign n35751 = n35750 ^ n1743 ^ 1'b0 ;
  assign n35752 = n35751 ^ n9244 ^ 1'b0 ;
  assign n35753 = n9133 | n17940 ;
  assign n35754 = n9507 & ~n35753 ;
  assign n35755 = n14445 | n35754 ;
  assign n35757 = n19784 & n35297 ;
  assign n35756 = n4609 & n5851 ;
  assign n35758 = n35757 ^ n35756 ^ 1'b0 ;
  assign n35759 = n12580 & ~n24565 ;
  assign n35762 = n14270 | n14878 ;
  assign n35760 = n5451 ^ n3993 ^ 1'b0 ;
  assign n35761 = n27078 & ~n35760 ;
  assign n35763 = n35762 ^ n35761 ^ 1'b0 ;
  assign n35764 = n10370 ^ n4519 ^ 1'b0 ;
  assign n35765 = n35764 ^ n8545 ^ 1'b0 ;
  assign n35766 = n28777 ^ n12690 ^ 1'b0 ;
  assign n35767 = n35 & n536 ;
  assign n35768 = ~n35 & n35767 ;
  assign n35769 = n509 & ~n35768 ;
  assign n35770 = n35768 & n35769 ;
  assign n35771 = n260 | n35770 ;
  assign n35772 = n14701 & ~n35771 ;
  assign n35773 = ~n106 & n2087 ;
  assign n35774 = n106 & n35773 ;
  assign n35775 = n10533 | n35774 ;
  assign n35776 = n35772 & ~n35775 ;
  assign n35777 = n874 & ~n35776 ;
  assign n35778 = n3647 | n4240 ;
  assign n35779 = n3647 & ~n35778 ;
  assign n35780 = n931 & ~n31153 ;
  assign n35781 = ~n931 & n35780 ;
  assign n35782 = n2005 & ~n4178 ;
  assign n35783 = n35781 & n35782 ;
  assign n35784 = n35779 | n35783 ;
  assign n35785 = n35777 & ~n35784 ;
  assign n35786 = ~n6271 & n28928 ;
  assign n35787 = ~n35083 & n35786 ;
  assign n35788 = n13232 | n35787 ;
  assign n35789 = ~n5152 & n35788 ;
  assign n35790 = n28338 & n35789 ;
  assign n35791 = ~n3101 & n4566 ;
  assign n35792 = n27263 & n35791 ;
  assign n35793 = n5505 & n12137 ;
  assign n35794 = n20298 | n35793 ;
  assign n35796 = n1981 | n27606 ;
  assign n35797 = n35796 ^ n6678 ^ 1'b0 ;
  assign n35798 = n27276 | n35797 ;
  assign n35795 = ~n12356 & n26799 ;
  assign n35799 = n35798 ^ n35795 ^ 1'b0 ;
  assign n35800 = n33650 ^ n33622 ^ 1'b0 ;
  assign n35801 = n27946 | n35800 ;
  assign n35802 = n3583 & ~n10839 ;
  assign n35803 = n20101 | n35802 ;
  assign n35804 = n35801 & ~n35803 ;
  assign n35805 = n3259 & n12575 ;
  assign n35806 = ~n2749 & n35805 ;
  assign n35807 = n34639 ^ n19528 ^ 1'b0 ;
  assign n35808 = n19645 & n35807 ;
  assign n35809 = n28428 ^ n515 ^ 1'b0 ;
  assign n35810 = n20352 ^ n9017 ^ 1'b0 ;
  assign n35811 = n67 | n35810 ;
  assign n35812 = n3054 & n4888 ;
  assign n35816 = n10329 | n11831 ;
  assign n35817 = n4768 | n35816 ;
  assign n35813 = n11630 ^ n10610 ^ 1'b0 ;
  assign n35814 = n5142 | n10215 ;
  assign n35815 = n35813 | n35814 ;
  assign n35818 = n35817 ^ n35815 ^ 1'b0 ;
  assign n35823 = n13144 ^ n8879 ^ 1'b0 ;
  assign n35824 = n3152 & ~n35823 ;
  assign n35819 = n11820 ^ n11576 ^ n6262 ;
  assign n35820 = n14538 ^ n2745 ^ 1'b0 ;
  assign n35821 = ~n35819 & n35820 ;
  assign n35822 = n35821 ^ n16833 ^ 1'b0 ;
  assign n35825 = n35824 ^ n35822 ^ n23335 ;
  assign n35826 = n18143 & ~n33092 ;
  assign n35827 = n18978 & n26249 ;
  assign n35828 = n15541 ^ n3556 ^ 1'b0 ;
  assign n35829 = n31730 & n35828 ;
  assign n35830 = n1542 & ~n25637 ;
  assign n35831 = n35830 ^ n32276 ^ 1'b0 ;
  assign n35832 = n27916 ^ n9912 ^ 1'b0 ;
  assign n35833 = ~n5416 & n35832 ;
  assign n35834 = ~n10900 & n25888 ;
  assign n35835 = ~n13373 & n35834 ;
  assign n35836 = n13792 & n21473 ;
  assign n35837 = n35835 & n35836 ;
  assign n35839 = ~n11099 & n31192 ;
  assign n35840 = n35839 ^ n3276 ^ 1'b0 ;
  assign n35841 = n5470 & n35840 ;
  assign n35842 = n24548 & n35841 ;
  assign n35838 = n12357 & n25716 ;
  assign n35843 = n35842 ^ n35838 ^ n18327 ;
  assign n35844 = n6035 ^ n1657 ^ 1'b0 ;
  assign n35845 = ~n9443 & n35844 ;
  assign n35846 = n35845 ^ n29995 ^ 1'b0 ;
  assign n35847 = n30935 | n35846 ;
  assign n35848 = n4550 & n20467 ;
  assign n35849 = n10121 | n35848 ;
  assign n35850 = n15066 & n23031 ;
  assign n35851 = n24657 ^ n16619 ^ 1'b0 ;
  assign n35852 = ~n1023 & n35851 ;
  assign n35853 = ( n911 & n9716 ) | ( n911 & n19165 ) | ( n9716 & n19165 ) ;
  assign n35854 = n35853 ^ n21386 ^ 1'b0 ;
  assign n35855 = n13480 & ~n35854 ;
  assign n35860 = n5908 & ~n8200 ;
  assign n35861 = n35860 ^ n15905 ^ 1'b0 ;
  assign n35859 = n2641 & n33818 ;
  assign n35862 = n35861 ^ n35859 ^ 1'b0 ;
  assign n35856 = n1073 | n13564 ;
  assign n35857 = n35856 ^ n27106 ^ 1'b0 ;
  assign n35858 = ~n23329 & n35857 ;
  assign n35863 = n35862 ^ n35858 ^ 1'b0 ;
  assign n35864 = n3529 | n7635 ;
  assign n35865 = n35864 ^ n1984 ^ 1'b0 ;
  assign n35866 = n35865 ^ n16905 ^ 1'b0 ;
  assign n35867 = n17434 | n28724 ;
  assign n35868 = n667 & ~n35867 ;
  assign n35869 = n7986 ^ n5497 ^ 1'b0 ;
  assign n35870 = n4555 | n20101 ;
  assign n35871 = n20101 & ~n35870 ;
  assign n35872 = ( ~n9899 & n31579 ) | ( ~n9899 & n35871 ) | ( n31579 & n35871 ) ;
  assign n35874 = ~n2950 & n11154 ;
  assign n35875 = n35874 ^ n15159 ^ 1'b0 ;
  assign n35873 = ~n654 & n7732 ;
  assign n35876 = n35875 ^ n35873 ^ 1'b0 ;
  assign n35877 = n9049 | n35876 ;
  assign n35878 = n30465 ^ n25668 ^ 1'b0 ;
  assign n35879 = n31995 & ~n35878 ;
  assign n35880 = ~n3912 & n20001 ;
  assign n35881 = n35880 ^ n18573 ^ 1'b0 ;
  assign n35882 = n1981 ^ n1502 ^ 1'b0 ;
  assign n35883 = n31072 ^ n27912 ^ 1'b0 ;
  assign n35884 = ~n11657 & n33872 ;
  assign n35885 = n35884 ^ n30521 ^ 1'b0 ;
  assign n35888 = n1276 ^ n578 ^ 1'b0 ;
  assign n35889 = n7208 & n35888 ;
  assign n35886 = n25010 & n29046 ;
  assign n35887 = ~n7193 & n35886 ;
  assign n35890 = n35889 ^ n35887 ^ 1'b0 ;
  assign n35891 = n28828 | n35890 ;
  assign n35892 = n35891 ^ n5946 ^ 1'b0 ;
  assign n35893 = ( n10149 & ~n35885 ) | ( n10149 & n35892 ) | ( ~n35885 & n35892 ) ;
  assign n35898 = n5241 ^ n1851 ^ 1'b0 ;
  assign n35899 = n6213 & n35898 ;
  assign n35900 = n25559 & n35899 ;
  assign n35894 = n7670 ^ n3268 ^ 1'b0 ;
  assign n35895 = n14459 | n29458 ;
  assign n35896 = n35894 | n35895 ;
  assign n35897 = n19983 & n35896 ;
  assign n35901 = n35900 ^ n35897 ^ 1'b0 ;
  assign n35902 = n4891 ^ n4433 ^ 1'b0 ;
  assign n35903 = n28311 ^ n17431 ^ 1'b0 ;
  assign n35904 = n9891 | n17917 ;
  assign n35905 = n13475 & ~n18566 ;
  assign n35906 = n35904 & n35905 ;
  assign n35910 = n25283 ^ n2634 ^ 1'b0 ;
  assign n35911 = ~n4593 & n35910 ;
  assign n35907 = n20949 ^ n9941 ^ 1'b0 ;
  assign n35908 = n8782 & n35907 ;
  assign n35909 = n12528 | n35908 ;
  assign n35912 = n35911 ^ n35909 ^ 1'b0 ;
  assign n35913 = ~n2670 & n35912 ;
  assign n35914 = n3584 & n35913 ;
  assign n35915 = n6618 & ~n13082 ;
  assign n35916 = n12195 & n35915 ;
  assign n35917 = n12759 ^ n5637 ^ 1'b0 ;
  assign n35918 = ( n14815 & ~n16442 ) | ( n14815 & n35917 ) | ( ~n16442 & n35917 ) ;
  assign n35919 = n35918 ^ n31867 ^ 1'b0 ;
  assign n35920 = n3111 & ~n3295 ;
  assign n35921 = n14248 & n35920 ;
  assign n35922 = n35921 ^ n25637 ^ 1'b0 ;
  assign n35923 = ~n5157 & n35922 ;
  assign n35924 = ~n33016 & n35923 ;
  assign n35925 = n2653 & n3437 ;
  assign n35926 = ~n21921 & n35925 ;
  assign n35927 = n1837 & n35926 ;
  assign n35928 = n136 | n15746 ;
  assign n35929 = n35928 ^ n15213 ^ 1'b0 ;
  assign n35930 = ( n997 & n2366 ) | ( n997 & n19534 ) | ( n2366 & n19534 ) ;
  assign n35931 = n28117 & n35930 ;
  assign n35932 = n22492 & ~n35931 ;
  assign n35933 = n20169 | n35932 ;
  assign n35934 = n16925 ^ n11000 ^ 1'b0 ;
  assign n35939 = n7016 | n20093 ;
  assign n35935 = n20232 ^ n4600 ^ 1'b0 ;
  assign n35936 = n25110 & ~n35935 ;
  assign n35937 = n12854 & ~n35936 ;
  assign n35938 = ~n4632 & n35937 ;
  assign n35940 = n35939 ^ n35938 ^ 1'b0 ;
  assign n35941 = ~n10670 & n35940 ;
  assign n35942 = n27785 ^ n25829 ^ 1'b0 ;
  assign n35943 = ~n9286 & n16896 ;
  assign n35944 = ~n35316 & n35943 ;
  assign n35945 = n14085 ^ n12656 ^ 1'b0 ;
  assign n35946 = ~n35944 & n35945 ;
  assign n35947 = n35946 ^ n27722 ^ 1'b0 ;
  assign n35948 = n33765 ^ n17005 ^ 1'b0 ;
  assign n35949 = ~n3522 & n6644 ;
  assign n35950 = ~n12471 & n35949 ;
  assign n35951 = n942 | n20367 ;
  assign n35952 = n11675 ^ n1609 ^ 1'b0 ;
  assign n35953 = n10728 ^ n10235 ^ 1'b0 ;
  assign n35954 = ~n35952 & n35953 ;
  assign n35955 = n3667 | n6293 ;
  assign n35956 = n35955 ^ n19946 ^ 1'b0 ;
  assign n35957 = n15783 & n35956 ;
  assign n35959 = n2173 & ~n11095 ;
  assign n35958 = n1969 & n2816 ;
  assign n35960 = n35959 ^ n35958 ^ 1'b0 ;
  assign n35961 = ~n961 & n35960 ;
  assign n35962 = n22600 ^ n12643 ^ 1'b0 ;
  assign n35963 = n30716 & ~n35962 ;
  assign n35964 = n35963 ^ n34432 ^ 1'b0 ;
  assign n35965 = n16915 | n20702 ;
  assign n35966 = n16528 ^ n13687 ^ 1'b0 ;
  assign n35967 = n13251 ^ n2491 ^ 1'b0 ;
  assign n35968 = ~n18927 & n35967 ;
  assign n35969 = n6741 & n35968 ;
  assign n35970 = n27980 & ~n35969 ;
  assign n35971 = n35966 & n35970 ;
  assign n35972 = ( ~n22153 & n27342 ) | ( ~n22153 & n35064 ) | ( n27342 & n35064 ) ;
  assign n35973 = ( n6856 & n35971 ) | ( n6856 & ~n35972 ) | ( n35971 & ~n35972 ) ;
  assign n35974 = n23327 ^ n14817 ^ n14038 ;
  assign n35975 = n11201 & n35974 ;
  assign n35976 = n11159 & n27224 ;
  assign n35977 = n24563 ^ n12433 ^ 1'b0 ;
  assign n35978 = n27781 & n35977 ;
  assign n35979 = n11758 | n20451 ;
  assign n35980 = n35978 | n35979 ;
  assign n35981 = ( n3040 & ~n8545 ) | ( n3040 & n21573 ) | ( ~n8545 & n21573 ) ;
  assign n35982 = n2346 & n7516 ;
  assign n35983 = n2176 & ~n35982 ;
  assign n35984 = n35983 ^ n12246 ^ 1'b0 ;
  assign n35985 = ( n11423 & n19975 ) | ( n11423 & ~n35984 ) | ( n19975 & ~n35984 ) ;
  assign n35986 = ~n15028 & n18547 ;
  assign n35987 = ~n35985 & n35986 ;
  assign n35988 = n5052 & ~n6452 ;
  assign n35989 = n35988 ^ n6095 ^ 1'b0 ;
  assign n35990 = ~n3951 & n35989 ;
  assign n35991 = ~n21189 & n35990 ;
  assign n35992 = n10901 & n35991 ;
  assign n35993 = n634 | n5984 ;
  assign n35994 = n18031 & n35993 ;
  assign n35995 = ~n8911 & n19428 ;
  assign n35996 = n4813 | n5742 ;
  assign n35997 = n11059 | n35996 ;
  assign n35998 = n7234 & ~n35997 ;
  assign n36000 = n3227 & ~n5626 ;
  assign n35999 = n799 & n8613 ;
  assign n36001 = n36000 ^ n35999 ^ 1'b0 ;
  assign n36002 = ~n2260 & n26176 ;
  assign n36003 = n36001 & n36002 ;
  assign n36004 = ( n9931 & n26322 ) | ( n9931 & n36003 ) | ( n26322 & n36003 ) ;
  assign n36005 = ~n14736 & n35129 ;
  assign n36006 = n14561 | n29541 ;
  assign n36007 = n18946 ^ n8951 ^ 1'b0 ;
  assign n36008 = n13157 | n13481 ;
  assign n36009 = n7916 | n36008 ;
  assign n36010 = n9882 ^ n2042 ^ 1'b0 ;
  assign n36011 = n6200 | n36010 ;
  assign n36015 = n1080 & n14798 ;
  assign n36012 = n1244 & ~n7802 ;
  assign n36013 = n36012 ^ n5057 ^ 1'b0 ;
  assign n36014 = n36013 ^ n9384 ^ 1'b0 ;
  assign n36016 = n36015 ^ n36014 ^ n14297 ;
  assign n36017 = ( n135 & ~n3780 ) | ( n135 & n17031 ) | ( ~n3780 & n17031 ) ;
  assign n36018 = n2719 ^ n1908 ^ 1'b0 ;
  assign n36019 = n36017 & n36018 ;
  assign n36020 = n19163 & n31109 ;
  assign n36021 = n36020 ^ n30169 ^ 1'b0 ;
  assign n36022 = ~n6831 & n8712 ;
  assign n36023 = n36022 ^ n1014 ^ 1'b0 ;
  assign n36024 = ~n21769 & n36023 ;
  assign n36029 = ( ~n1884 & n18540 ) | ( ~n1884 & n21390 ) | ( n18540 & n21390 ) ;
  assign n36025 = n12666 ^ n8717 ^ 1'b0 ;
  assign n36026 = ~n5260 & n36025 ;
  assign n36027 = ~n9133 & n35593 ;
  assign n36028 = n36026 & ~n36027 ;
  assign n36030 = n36029 ^ n36028 ^ 1'b0 ;
  assign n36031 = n36024 | n36030 ;
  assign n36032 = ~n18553 & n36031 ;
  assign n36033 = n14652 ^ n7266 ^ n6839 ;
  assign n36034 = n14597 | n36033 ;
  assign n36035 = n16221 & ~n32171 ;
  assign n36036 = ~n36034 & n36035 ;
  assign n36037 = n36036 ^ n32839 ^ 1'b0 ;
  assign n36038 = n36037 ^ n2108 ^ 1'b0 ;
  assign n36039 = n12651 & ~n17388 ;
  assign n36040 = n4804 ^ n365 ^ 1'b0 ;
  assign n36041 = n4402 ^ n1660 ^ n536 ;
  assign n36042 = ~n36040 & n36041 ;
  assign n36043 = n7569 | n36042 ;
  assign n36044 = n2719 & ~n24461 ;
  assign n36045 = n489 & n5371 ;
  assign n36046 = n6236 & n7138 ;
  assign n36047 = ~n8894 & n17092 ;
  assign n36048 = ~n36046 & n36047 ;
  assign n36049 = n4607 & ~n10056 ;
  assign n36050 = n8249 & n36049 ;
  assign n36051 = n21404 & n33491 ;
  assign n36052 = ~n11009 & n36051 ;
  assign n36053 = n36052 ^ n35072 ^ n4170 ;
  assign n36054 = n8197 ^ n1134 ^ 1'b0 ;
  assign n36055 = n1023 | n36054 ;
  assign n36056 = n1517 & ~n36055 ;
  assign n36057 = n1165 & ~n3609 ;
  assign n36058 = ~n1165 & n36057 ;
  assign n36059 = ~n7270 & n9401 ;
  assign n36060 = n7270 & n36059 ;
  assign n36061 = n36058 | n36060 ;
  assign n36062 = n36061 ^ n5796 ^ 1'b0 ;
  assign n36063 = n36062 ^ n29237 ^ 1'b0 ;
  assign n36064 = n19509 ^ n11794 ^ 1'b0 ;
  assign n36065 = n5404 & n36064 ;
  assign n36066 = n29935 & n36065 ;
  assign n36067 = n20281 | n22891 ;
  assign n36068 = n36067 ^ n23766 ^ 1'b0 ;
  assign n36069 = ~n21418 & n21438 ;
  assign n36070 = n8449 ^ n220 ^ 1'b0 ;
  assign n36071 = n36069 & ~n36070 ;
  assign n36072 = n31480 ^ n27923 ^ n7536 ;
  assign n36073 = n36072 ^ n18072 ^ n11523 ;
  assign n36074 = n36037 ^ n23496 ^ 1'b0 ;
  assign n36075 = n10720 ^ n10183 ^ 1'b0 ;
  assign n36076 = n33819 ^ n18856 ^ 1'b0 ;
  assign n36077 = n28509 & n36076 ;
  assign n36078 = n31645 ^ n11162 ^ n4551 ;
  assign n36079 = n8217 | n35706 ;
  assign n36080 = n36078 & ~n36079 ;
  assign n36081 = ~n19019 & n23252 ;
  assign n36082 = n36081 ^ n813 ^ 1'b0 ;
  assign n36083 = n18635 & ~n28903 ;
  assign n36084 = n7798 & ~n24130 ;
  assign n36085 = n7194 ^ n3274 ^ 1'b0 ;
  assign n36086 = n8281 & n36085 ;
  assign n36087 = n36086 ^ n4819 ^ 1'b0 ;
  assign n36088 = n4895 & ~n19180 ;
  assign n36089 = n182 & ~n25314 ;
  assign n36090 = n36089 ^ n1455 ^ 1'b0 ;
  assign n36091 = ( n2238 & ~n2628 ) | ( n2238 & n36090 ) | ( ~n2628 & n36090 ) ;
  assign n36092 = n36091 ^ n7369 ^ 1'b0 ;
  assign n36093 = ~n36088 & n36092 ;
  assign n36094 = ~n14589 & n23695 ;
  assign n36095 = n34974 & n36094 ;
  assign n36098 = n3644 ^ n527 ^ 1'b0 ;
  assign n36097 = n2600 & n15635 ;
  assign n36099 = n36098 ^ n36097 ^ 1'b0 ;
  assign n36096 = n12726 & ~n29866 ;
  assign n36100 = n36099 ^ n36096 ^ 1'b0 ;
  assign n36101 = ~n511 & n22859 ;
  assign n36102 = n1814 | n30134 ;
  assign n36103 = n1329 & n20279 ;
  assign n36104 = n27470 ^ n2854 ^ 1'b0 ;
  assign n36105 = n4083 & n21863 ;
  assign n36106 = ~n11258 & n36105 ;
  assign n36107 = n12833 | n30562 ;
  assign n36108 = n20959 ^ n8525 ^ 1'b0 ;
  assign n36109 = ~n19170 & n35857 ;
  assign n36110 = ~n36108 & n36109 ;
  assign n36111 = n18138 ^ n1116 ^ 1'b0 ;
  assign n36112 = ~n22177 & n36111 ;
  assign n36113 = n36112 ^ n15588 ^ 1'b0 ;
  assign n36114 = ( n578 & n15699 ) | ( n578 & n22056 ) | ( n15699 & n22056 ) ;
  assign n36115 = n31967 & n36114 ;
  assign n36116 = n36115 ^ n9478 ^ 1'b0 ;
  assign n36117 = n31587 & ~n36116 ;
  assign n36118 = n3939 & n36117 ;
  assign n36119 = ~n310 & n5353 ;
  assign n36120 = ~n9151 & n36119 ;
  assign n36122 = n6768 & n19945 ;
  assign n36123 = n36122 ^ n26156 ^ 1'b0 ;
  assign n36121 = ~n3674 & n25373 ;
  assign n36124 = n36123 ^ n36121 ^ 1'b0 ;
  assign n36125 = ~n22901 & n30599 ;
  assign n36126 = ~n10816 & n36125 ;
  assign n36127 = n8324 | n36126 ;
  assign n36128 = n36127 ^ n11599 ^ 1'b0 ;
  assign n36129 = n15017 ^ n85 ^ 1'b0 ;
  assign n36130 = n36129 ^ n29156 ^ 1'b0 ;
  assign n36131 = ~n13136 & n36130 ;
  assign n36132 = n4757 & n25565 ;
  assign n36133 = n36132 ^ n2137 ^ 1'b0 ;
  assign n36134 = ~n13657 & n36133 ;
  assign n36135 = n36134 ^ n5483 ^ 1'b0 ;
  assign n36136 = ( ~n2390 & n9653 ) | ( ~n2390 & n36135 ) | ( n9653 & n36135 ) ;
  assign n36137 = ~n22313 & n28815 ;
  assign n36138 = ~n22321 & n36137 ;
  assign n36139 = n36138 ^ n4301 ^ 1'b0 ;
  assign n36140 = n2379 | n8553 ;
  assign n36141 = n31248 & ~n36140 ;
  assign n36142 = n23821 ^ n7822 ^ 1'b0 ;
  assign n36143 = n21902 ^ n302 ^ 1'b0 ;
  assign n36144 = n459 | n13707 ;
  assign n36145 = n36144 ^ n9401 ^ 1'b0 ;
  assign n36146 = ( n15878 & ~n26874 ) | ( n15878 & n36145 ) | ( ~n26874 & n36145 ) ;
  assign n36147 = n20702 | n36146 ;
  assign n36148 = n30438 ^ n83 ^ 1'b0 ;
  assign n36149 = n5714 & n36148 ;
  assign n36150 = n1690 & ~n11523 ;
  assign n36151 = n12104 & n32198 ;
  assign n36152 = ( ~n8529 & n36150 ) | ( ~n8529 & n36151 ) | ( n36150 & n36151 ) ;
  assign n36153 = n13557 ^ n3745 ^ 1'b0 ;
  assign n36154 = n11274 | n36153 ;
  assign n36155 = n36154 ^ n7690 ^ 1'b0 ;
  assign n36156 = n138 & ~n10783 ;
  assign n36157 = n11751 & n36156 ;
  assign n36158 = n27682 & ~n30935 ;
  assign n36159 = n36158 ^ n2066 ^ 1'b0 ;
  assign n36160 = ~n11198 & n12438 ;
  assign n36161 = n36160 ^ n11253 ^ 1'b0 ;
  assign n36162 = n36159 & ~n36161 ;
  assign n36163 = n36162 ^ n4267 ^ 1'b0 ;
  assign n36164 = n36157 & n36163 ;
  assign n36165 = ~n6647 & n32532 ;
  assign n36166 = n27075 & n36165 ;
  assign n36167 = n27152 ^ n890 ^ 1'b0 ;
  assign n36169 = ~n31713 & n34110 ;
  assign n36168 = n25469 ^ n8480 ^ 1'b0 ;
  assign n36170 = n36169 ^ n36168 ^ 1'b0 ;
  assign n36177 = n22005 ^ n7335 ^ 1'b0 ;
  assign n36178 = n1286 | n36177 ;
  assign n36175 = n13139 ^ n13122 ^ n8099 ;
  assign n36173 = ~n6388 & n20702 ;
  assign n36174 = ~n5501 & n36173 ;
  assign n36176 = n36175 ^ n36174 ^ 1'b0 ;
  assign n36171 = ~n682 & n2079 ;
  assign n36172 = n36171 ^ n379 ^ 1'b0 ;
  assign n36179 = n36178 ^ n36176 ^ n36172 ;
  assign n36180 = n36179 ^ n1843 ^ 1'b0 ;
  assign n36181 = n19851 & ~n25588 ;
  assign n36184 = n22835 & n33037 ;
  assign n36182 = n43 & n5472 ;
  assign n36183 = n36182 ^ n20169 ^ 1'b0 ;
  assign n36185 = n36184 ^ n36183 ^ 1'b0 ;
  assign n36186 = n611 | n9281 ;
  assign n36187 = ( n7137 & n33491 ) | ( n7137 & n36186 ) | ( n33491 & n36186 ) ;
  assign n36188 = n26258 ^ n7924 ^ 1'b0 ;
  assign n36189 = n17929 | n36188 ;
  assign n36190 = n4958 & n5181 ;
  assign n36191 = n34694 & n36190 ;
  assign n36192 = n16084 & n24986 ;
  assign n36193 = n1069 & n36192 ;
  assign n36194 = ~n24758 & n36193 ;
  assign n36195 = n9427 & n25429 ;
  assign n36196 = ( ~n1973 & n4780 ) | ( ~n1973 & n36195 ) | ( n4780 & n36195 ) ;
  assign n36197 = n12996 & ~n22464 ;
  assign n36198 = n1434 | n36197 ;
  assign n36199 = n5938 & n36198 ;
  assign n36200 = n36199 ^ n15 ^ 1'b0 ;
  assign n36201 = ~n49 & n17017 ;
  assign n36202 = n24633 ^ n13184 ^ 1'b0 ;
  assign n36203 = ~n36201 & n36202 ;
  assign n36204 = n6057 & n9848 ;
  assign n36205 = ~n33993 & n36204 ;
  assign n36206 = n20506 | n30364 ;
  assign n36207 = n220 & ~n36206 ;
  assign n36208 = n3124 & ~n10220 ;
  assign n36209 = n36208 ^ n17682 ^ 1'b0 ;
  assign n36210 = n20346 & n36209 ;
  assign n36211 = n1918 | n24719 ;
  assign n36212 = n36211 ^ n5350 ^ 1'b0 ;
  assign n36213 = n5136 & ~n25462 ;
  assign n36214 = n13855 | n23824 ;
  assign n36215 = ~n13167 & n14221 ;
  assign n36216 = n36215 ^ n11194 ^ 1'b0 ;
  assign n36217 = n1978 & ~n36216 ;
  assign n36218 = n36217 ^ n31674 ^ 1'b0 ;
  assign n36220 = n18981 ^ n18074 ^ n1834 ;
  assign n36219 = ~n4276 & n13091 ;
  assign n36221 = n36220 ^ n36219 ^ 1'b0 ;
  assign n36222 = n2236 & n5016 ;
  assign n36223 = n36222 ^ n13899 ^ 1'b0 ;
  assign n36224 = n29584 ^ n11437 ^ 1'b0 ;
  assign n36225 = n36223 & n36224 ;
  assign n36226 = n21848 & ~n35708 ;
  assign n36227 = n36226 ^ n19443 ^ 1'b0 ;
  assign n36228 = n4121 ^ n2044 ^ 1'b0 ;
  assign n36229 = ~n4305 & n25681 ;
  assign n36230 = ~n9916 & n36229 ;
  assign n36231 = n3193 ^ n57 ^ 1'b0 ;
  assign n36232 = n8150 ^ n3894 ^ 1'b0 ;
  assign n36233 = ~n16111 & n36232 ;
  assign n36234 = n13393 ^ n12211 ^ 1'b0 ;
  assign n36235 = ~n8708 & n17718 ;
  assign n36236 = n3449 & n36235 ;
  assign n36237 = n2983 | n26743 ;
  assign n36238 = n36236 & ~n36237 ;
  assign n36239 = n25598 & n32361 ;
  assign n36240 = n10761 & n36239 ;
  assign n36241 = n1264 & n16650 ;
  assign n36242 = n36241 ^ n19520 ^ 1'b0 ;
  assign n36243 = n12994 & n23884 ;
  assign n36245 = n9180 ^ n6312 ^ 1'b0 ;
  assign n36244 = n400 | n12043 ;
  assign n36246 = n36245 ^ n36244 ^ 1'b0 ;
  assign n36247 = ~n2826 & n11289 ;
  assign n36248 = n36247 ^ n13821 ^ 1'b0 ;
  assign n36249 = n13117 | n31576 ;
  assign n36250 = n36249 ^ n18099 ^ 1'b0 ;
  assign n36251 = n36250 ^ n24256 ^ 1'b0 ;
  assign n36252 = n764 & ~n3315 ;
  assign n36253 = ~n764 & n36252 ;
  assign n36254 = n3280 & ~n36253 ;
  assign n36255 = ~n3280 & n36254 ;
  assign n36256 = n36255 ^ n16669 ^ 1'b0 ;
  assign n36265 = ~n31 & n849 ;
  assign n36266 = n31 & n36265 ;
  assign n36257 = ~n588 & n2355 ;
  assign n36258 = n588 & n36257 ;
  assign n36259 = n27 & n552 ;
  assign n36260 = ~n27 & n36259 ;
  assign n36261 = n4895 & n36260 ;
  assign n36262 = ~n2824 & n36261 ;
  assign n36263 = n36258 & n36262 ;
  assign n36264 = n2282 | n36263 ;
  assign n36267 = n36266 ^ n36264 ^ 1'b0 ;
  assign n36268 = n36256 & ~n36267 ;
  assign n36269 = ~n36256 & n36268 ;
  assign n36270 = n23490 & ~n25824 ;
  assign n36271 = n36270 ^ n14351 ^ 1'b0 ;
  assign n36272 = n12226 | n18706 ;
  assign n36273 = n36271 | n36272 ;
  assign n36274 = ~n3388 & n36273 ;
  assign n36275 = n36269 & n36274 ;
  assign n36276 = ( n6219 & n13285 ) | ( n6219 & ~n13306 ) | ( n13285 & ~n13306 ) ;
  assign n36277 = n36276 ^ n23767 ^ 1'b0 ;
  assign n36278 = ~n1901 & n8346 ;
  assign n36279 = n3139 | n36278 ;
  assign n36280 = n36279 ^ n11927 ^ 1'b0 ;
  assign n36281 = n28588 | n36280 ;
  assign n36282 = n20801 ^ n5901 ^ 1'b0 ;
  assign n36283 = n2883 & n36282 ;
  assign n36284 = n17129 & n32934 ;
  assign n36285 = n1975 ^ n1422 ^ 1'b0 ;
  assign n36286 = n34147 ^ n251 ^ 1'b0 ;
  assign n36287 = n598 & n36286 ;
  assign n36288 = n9151 ^ n1323 ^ 1'b0 ;
  assign n36289 = n7476 & ~n36288 ;
  assign n36290 = n10171 & n10323 ;
  assign n36291 = n36290 ^ n34893 ^ n11477 ;
  assign n36292 = ~n1020 & n13707 ;
  assign n36293 = n36292 ^ n36245 ^ 1'b0 ;
  assign n36294 = ( n12799 & n17189 ) | ( n12799 & n36293 ) | ( n17189 & n36293 ) ;
  assign n36295 = n11637 ^ n9536 ^ 1'b0 ;
  assign n36296 = n1771 | n36295 ;
  assign n36297 = n11553 & ~n25466 ;
  assign n36298 = n36296 & n36297 ;
  assign n36299 = n24094 | n36298 ;
  assign n36300 = n26400 ^ n19566 ^ n10537 ;
  assign n36301 = n5563 & n36300 ;
  assign n36302 = n15468 ^ x6 ^ 1'b0 ;
  assign n36303 = n36302 ^ n6805 ^ 1'b0 ;
  assign n36304 = n36301 & n36303 ;
  assign n36305 = n9261 & n30548 ;
  assign n36306 = n1337 & n36305 ;
  assign n36307 = ~n8058 & n11501 ;
  assign n36308 = ~n3361 & n36307 ;
  assign n36309 = n6176 ^ n3305 ^ 1'b0 ;
  assign n36310 = n32555 ^ n24664 ^ n15185 ;
  assign n36311 = n26602 ^ n8224 ^ 1'b0 ;
  assign n36312 = n14598 ^ n1743 ^ 1'b0 ;
  assign n36313 = n15038 & ~n36312 ;
  assign n36314 = n2258 ^ n2158 ^ 1'b0 ;
  assign n36315 = n16811 | n36314 ;
  assign n36316 = n36315 ^ n19182 ^ 1'b0 ;
  assign n36317 = n18587 ^ n3574 ^ 1'b0 ;
  assign n36318 = n36317 ^ n13091 ^ n12513 ;
  assign n36319 = ~n371 & n16391 ;
  assign n36320 = n36319 ^ n1372 ^ n1003 ;
  assign n36321 = n36320 ^ n31773 ^ 1'b0 ;
  assign n36322 = n996 & n23997 ;
  assign n36323 = n16705 & ~n22558 ;
  assign n36324 = n35312 ^ n30653 ^ n5867 ;
  assign n36325 = n36324 ^ n6326 ^ n40 ;
  assign n36326 = n5518 & n11336 ;
  assign n36327 = n36326 ^ n3124 ^ 1'b0 ;
  assign n36328 = ~n7918 & n36327 ;
  assign n36329 = n7893 & ~n36328 ;
  assign n36330 = n1347 & n4328 ;
  assign n36331 = n36330 ^ n12183 ^ 1'b0 ;
  assign n36332 = n27080 | n34325 ;
  assign n36333 = n23188 ^ n8784 ^ 1'b0 ;
  assign n36334 = n2735 & n36333 ;
  assign n36335 = ~n16020 & n17221 ;
  assign n36336 = ~n36334 & n36335 ;
  assign n36337 = n23243 & n36129 ;
  assign n36338 = n36337 ^ n19774 ^ 1'b0 ;
  assign n36339 = n15254 & n26783 ;
  assign n36340 = ~n18473 & n36339 ;
  assign n36341 = n9758 ^ n908 ^ 1'b0 ;
  assign n36342 = n11391 & n36341 ;
  assign n36343 = n36342 ^ n17823 ^ n11215 ;
  assign n36344 = ~n15622 & n23573 ;
  assign n36345 = n2521 | n4137 ;
  assign n36346 = n36345 ^ n36207 ^ 1'b0 ;
  assign n36347 = n25269 | n28267 ;
  assign n36348 = n36347 ^ n4789 ^ 1'b0 ;
  assign n36349 = n26196 & n29997 ;
  assign n36350 = n36349 ^ n11338 ^ 1'b0 ;
  assign n36351 = n1662 | n10391 ;
  assign n36352 = n4856 & ~n36351 ;
  assign n36353 = n16659 ^ n3718 ^ 1'b0 ;
  assign n36354 = n36352 | n36353 ;
  assign n36355 = n26680 & n33929 ;
  assign n36356 = n3277 | n13413 ;
  assign n36357 = n6442 & ~n36356 ;
  assign n36358 = n17099 & n17364 ;
  assign n36359 = n36357 & n36358 ;
  assign n36360 = ~n1445 & n2940 ;
  assign n36361 = ( n1398 & ~n14428 ) | ( n1398 & n32382 ) | ( ~n14428 & n32382 ) ;
  assign n36362 = n2460 & ~n36361 ;
  assign n36363 = n9908 | n36362 ;
  assign n36364 = n4222 & ~n36363 ;
  assign n36365 = n81 & ~n10495 ;
  assign n36366 = n2222 & n12718 ;
  assign n36367 = n13825 & n14484 ;
  assign n36368 = n36367 ^ n7293 ^ 1'b0 ;
  assign n36369 = n11438 & n28352 ;
  assign n36370 = ( n1363 & ~n12831 ) | ( n1363 & n19356 ) | ( ~n12831 & n19356 ) ;
  assign n36371 = n5743 & ~n12592 ;
  assign n36372 = n684 & n5933 ;
  assign n36373 = n36372 ^ n5144 ^ 1'b0 ;
  assign n36374 = n4279 & n12576 ;
  assign n36375 = n3633 & n36374 ;
  assign n36376 = n6001 & n14845 ;
  assign n36377 = n29491 ^ n21651 ^ 1'b0 ;
  assign n36378 = ~n12829 & n36377 ;
  assign n36379 = ~n29723 & n36378 ;
  assign n36380 = n17467 & n36379 ;
  assign n36381 = n28750 | n36380 ;
  assign n36382 = ~n11951 & n24137 ;
  assign n36383 = n9810 & n36382 ;
  assign n36384 = n16536 | n25639 ;
  assign n36385 = ~n5478 & n19526 ;
  assign n36386 = n29486 | n36385 ;
  assign n36387 = n36384 & ~n36386 ;
  assign n36388 = n18550 ^ n1939 ^ 1'b0 ;
  assign n36389 = n36388 ^ n23375 ^ 1'b0 ;
  assign n36390 = n13934 & n36389 ;
  assign n36391 = ~n200 & n14159 ;
  assign n36392 = ~n10396 & n36391 ;
  assign n36393 = n14652 ^ n2580 ^ 1'b0 ;
  assign n36394 = ~n8714 & n36393 ;
  assign n36395 = n12390 & n36394 ;
  assign n36396 = n12507 ^ n8582 ^ n2338 ;
  assign n36397 = ~n6574 & n36396 ;
  assign n36398 = n36397 ^ n1834 ^ 1'b0 ;
  assign n36399 = n36398 ^ n23160 ^ n10675 ;
  assign n36400 = ( ~n304 & n9029 ) | ( ~n304 & n36399 ) | ( n9029 & n36399 ) ;
  assign n36401 = ~n12055 & n35467 ;
  assign n36407 = n9071 | n27616 ;
  assign n36403 = n18866 & ~n22834 ;
  assign n36402 = n16801 | n16887 ;
  assign n36404 = n36403 ^ n36402 ^ 1'b0 ;
  assign n36405 = n9693 ^ n5592 ^ 1'b0 ;
  assign n36406 = ~n36404 & n36405 ;
  assign n36408 = n36407 ^ n36406 ^ 1'b0 ;
  assign n36409 = n36401 & ~n36408 ;
  assign n36410 = n4332 | n13526 ;
  assign n36411 = n5362 & ~n36410 ;
  assign n36412 = n8120 & n11567 ;
  assign n36413 = n36412 ^ n33895 ^ n28750 ;
  assign n36414 = n15992 & n36413 ;
  assign n36415 = ~n29879 & n36414 ;
  assign n36416 = n22145 ^ n17592 ^ 1'b0 ;
  assign n36417 = ( n2946 & n20263 ) | ( n2946 & ~n36416 ) | ( n20263 & ~n36416 ) ;
  assign n36418 = n1697 & ~n20037 ;
  assign n36419 = n36418 ^ n5739 ^ 1'b0 ;
  assign n36420 = n17017 ^ n4346 ^ 1'b0 ;
  assign n36421 = n11697 & n36420 ;
  assign n36422 = n9260 & n36421 ;
  assign n36423 = n13587 & n15246 ;
  assign n36424 = n27849 & n36423 ;
  assign n36425 = n7243 & n10892 ;
  assign n36426 = n4841 ^ n1908 ^ 1'b0 ;
  assign n36427 = n36426 ^ n34576 ^ n20769 ;
  assign n36428 = n18007 ^ n9596 ^ 1'b0 ;
  assign n36429 = n1542 & ~n35169 ;
  assign n36430 = n13136 | n21435 ;
  assign n36431 = n36430 ^ n8021 ^ 1'b0 ;
  assign n36432 = n12573 & n36431 ;
  assign n36433 = n6898 & n7357 ;
  assign n36434 = n36433 ^ n11701 ^ 1'b0 ;
  assign n36437 = n3613 & ~n6556 ;
  assign n36438 = n6051 & n36437 ;
  assign n36435 = n23208 ^ n10183 ^ 1'b0 ;
  assign n36436 = n35494 | n36435 ;
  assign n36439 = n36438 ^ n36436 ^ 1'b0 ;
  assign n36440 = n3587 & n36439 ;
  assign n36441 = n36440 ^ n26359 ^ 1'b0 ;
  assign n36442 = n36441 ^ n25550 ^ 1'b0 ;
  assign n36443 = ~n33203 & n36442 ;
  assign n36444 = ( n15159 & ~n36434 ) | ( n15159 & n36443 ) | ( ~n36434 & n36443 ) ;
  assign n36445 = n36444 ^ n1712 ^ 1'b0 ;
  assign n36446 = ( n9000 & n22140 ) | ( n9000 & n23571 ) | ( n22140 & n23571 ) ;
  assign n36447 = n2067 | n15646 ;
  assign n36448 = n14404 & ~n31451 ;
  assign n36449 = n36448 ^ n802 ^ 1'b0 ;
  assign n36450 = n19153 ^ n10740 ^ 1'b0 ;
  assign n36451 = n6707 & ~n36450 ;
  assign n36452 = n14067 & ~n23491 ;
  assign n36453 = n11404 | n17989 ;
  assign n36454 = n12984 & ~n36453 ;
  assign n36455 = n36454 ^ n4428 ^ 1'b0 ;
  assign n36456 = n36455 ^ n12941 ^ 1'b0 ;
  assign n36457 = n19511 & n36456 ;
  assign n36458 = n4121 | n34446 ;
  assign n36459 = n36458 ^ n318 ^ 1'b0 ;
  assign n36460 = ~n16696 & n24197 ;
  assign n36461 = n36460 ^ n7242 ^ 1'b0 ;
  assign n36462 = n27002 & ~n36461 ;
  assign n36463 = ~n9772 & n23067 ;
  assign n36464 = n36463 ^ n33130 ^ n1392 ;
  assign n36465 = ~n33220 & n36464 ;
  assign n36466 = n24931 & n36465 ;
  assign n36467 = n15069 ^ n9887 ^ 1'b0 ;
  assign n36468 = ~n24550 & n28592 ;
  assign n36469 = n36467 & n36468 ;
  assign n36470 = ~n121 & n36469 ;
  assign n36471 = n36470 ^ n3500 ^ 1'b0 ;
  assign n36472 = n899 | n22107 ;
  assign n36473 = n36472 ^ n20354 ^ n20001 ;
  assign n36474 = n3071 | n14165 ;
  assign n36475 = n16294 | n36474 ;
  assign n36476 = n13529 & ~n36475 ;
  assign n36477 = n36476 ^ n32943 ^ 1'b0 ;
  assign n36478 = n4506 & n36477 ;
  assign n36479 = ~n1182 & n3391 ;
  assign n36480 = n5458 & n36479 ;
  assign n36481 = n1933 & n36480 ;
  assign n36482 = n4570 | n5510 ;
  assign n36483 = ~n795 & n3512 ;
  assign n36484 = n36483 ^ n1590 ^ 1'b0 ;
  assign n36488 = n25096 ^ n71 ^ 1'b0 ;
  assign n36489 = n7735 & n36488 ;
  assign n36485 = ~n7484 & n10345 ;
  assign n36486 = n16393 | n36485 ;
  assign n36487 = n22379 & ~n36486 ;
  assign n36490 = n36489 ^ n36487 ^ n7668 ;
  assign n36491 = n459 & ~n35393 ;
  assign n36492 = n914 & n14087 ;
  assign n36493 = ~n32514 & n36492 ;
  assign n36494 = ~n13562 & n36493 ;
  assign n36495 = n23467 ^ n12690 ^ 1'b0 ;
  assign n36496 = ~n3042 & n32041 ;
  assign n36497 = n3610 | n4501 ;
  assign n36498 = n33481 ^ n6704 ^ 1'b0 ;
  assign n36499 = n8289 & ~n36083 ;
  assign n36500 = n1851 & ~n8297 ;
  assign n36501 = ~n36364 & n36500 ;
  assign n36502 = ~n19997 & n36501 ;
  assign n36505 = n2128 & ~n3698 ;
  assign n36503 = n488 & ~n4119 ;
  assign n36504 = n10231 & ~n36503 ;
  assign n36506 = n36505 ^ n36504 ^ 1'b0 ;
  assign n36507 = n6814 ^ n1327 ^ 1'b0 ;
  assign n36508 = n16167 | n36507 ;
  assign n36509 = n36508 ^ n21091 ^ n12466 ;
  assign n36510 = n29980 ^ n9089 ^ 1'b0 ;
  assign n36511 = n10646 & ~n36510 ;
  assign n36512 = n14402 ^ n8621 ^ 1'b0 ;
  assign n36513 = n27186 ^ n7847 ^ n1918 ;
  assign n36514 = n7792 | n36513 ;
  assign n36515 = n9687 ^ n1431 ^ 1'b0 ;
  assign n36516 = n36515 ^ n9525 ^ n1199 ;
  assign n36517 = ~n4422 & n20913 ;
  assign n36518 = n3444 & n36517 ;
  assign n36519 = n24658 | n36518 ;
  assign n36520 = n31002 ^ n21967 ^ 1'b0 ;
  assign n36521 = n3550 ^ n2093 ^ 1'b0 ;
  assign n36522 = ~n31808 & n34219 ;
  assign n36523 = n6618 & ~n14897 ;
  assign n36524 = n25743 ^ n7887 ^ 1'b0 ;
  assign n36525 = ( n29483 & ~n36523 ) | ( n29483 & n36524 ) | ( ~n36523 & n36524 ) ;
  assign n36526 = n470 & ~n3584 ;
  assign n36527 = n36526 ^ n7038 ^ 1'b0 ;
  assign n36528 = n12144 | n36527 ;
  assign n36529 = n33699 & ~n36528 ;
  assign n36530 = n1360 & ~n12342 ;
  assign n36531 = n36530 ^ n13048 ^ 1'b0 ;
  assign n36532 = ~n463 & n34066 ;
  assign n36533 = ~n36531 & n36532 ;
  assign n36534 = ( ~n10166 & n16453 ) | ( ~n10166 & n34760 ) | ( n16453 & n34760 ) ;
  assign n36535 = n36534 ^ n1191 ^ 1'b0 ;
  assign n36536 = ~n23540 & n36535 ;
  assign n36537 = n34073 ^ n33031 ^ 1'b0 ;
  assign n36538 = n5076 | n9748 ;
  assign n36539 = n3080 | n31777 ;
  assign n36540 = n33059 ^ n17876 ^ 1'b0 ;
  assign n36541 = n5001 & n36540 ;
  assign n36542 = n14848 & n15851 ;
  assign n36543 = n36542 ^ n13905 ^ 1'b0 ;
  assign n36544 = n1422 & n36543 ;
  assign n36545 = ~n3674 & n36544 ;
  assign n36546 = n18051 & n36545 ;
  assign n36547 = n30358 ^ n23395 ^ 1'b0 ;
  assign n36548 = n18858 ^ n2683 ^ 1'b0 ;
  assign n36549 = n32612 ^ n5648 ^ 1'b0 ;
  assign n36550 = n36548 & ~n36549 ;
  assign n36551 = n16777 ^ n3758 ^ 1'b0 ;
  assign n36552 = n16843 & n36551 ;
  assign n36553 = n11065 ^ n2287 ^ 1'b0 ;
  assign n36554 = n36553 ^ n15406 ^ 1'b0 ;
  assign n36555 = ( n489 & ~n24325 ) | ( n489 & n36554 ) | ( ~n24325 & n36554 ) ;
  assign n36556 = n15828 & ~n24014 ;
  assign n36557 = n25363 ^ n17369 ^ 1'b0 ;
  assign n36558 = n8763 & ~n9850 ;
  assign n36559 = n36558 ^ n7630 ^ 1'b0 ;
  assign n36560 = n27033 & ~n36559 ;
  assign n36561 = n36560 ^ n6140 ^ 1'b0 ;
  assign n36562 = ~n4013 & n36561 ;
  assign n36563 = n28203 ^ n20685 ^ 1'b0 ;
  assign n36564 = ~n16062 & n36563 ;
  assign n36566 = n6231 | n18905 ;
  assign n36565 = n4613 | n22086 ;
  assign n36567 = n36566 ^ n36565 ^ 1'b0 ;
  assign n36568 = n7921 ^ n453 ^ 1'b0 ;
  assign n36569 = n32982 & ~n36568 ;
  assign n36570 = n36569 ^ n3449 ^ 1'b0 ;
  assign n36571 = n36570 ^ n8287 ^ 1'b0 ;
  assign n36572 = n25351 ^ n20108 ^ 1'b0 ;
  assign n36573 = n94 & ~n714 ;
  assign n36574 = ~n14244 & n36573 ;
  assign n36575 = n36574 ^ n11211 ^ 1'b0 ;
  assign n36576 = n9163 & n36575 ;
  assign n36577 = n3257 & ~n32667 ;
  assign n36578 = n19395 ^ n4956 ^ 1'b0 ;
  assign n36579 = n22314 | n36578 ;
  assign n36580 = n25289 ^ n15347 ^ n2317 ;
  assign n36581 = n16268 & ~n26734 ;
  assign n36582 = ~n7285 & n28958 ;
  assign n36583 = ~n10033 & n12111 ;
  assign n36584 = n27644 & n35306 ;
  assign n36585 = ~n445 & n36584 ;
  assign n36586 = n27336 ^ n13975 ^ 1'b0 ;
  assign n36587 = n36586 ^ n18264 ^ 1'b0 ;
  assign n36588 = n4659 | n36587 ;
  assign n36589 = n17314 & ~n27634 ;
  assign n36590 = n24384 & ~n36589 ;
  assign n36591 = ( ~n6995 & n34924 ) | ( ~n6995 & n36590 ) | ( n34924 & n36590 ) ;
  assign n36592 = n8124 & n13712 ;
  assign n36593 = n28968 & n36592 ;
  assign n36594 = n36593 ^ n11175 ^ 1'b0 ;
  assign n36595 = n7034 & n16384 ;
  assign n36596 = ~n18191 & n36595 ;
  assign n36597 = ~n5580 & n8256 ;
  assign n36598 = n4970 | n34303 ;
  assign n36599 = n1740 & ~n17411 ;
  assign n36600 = n20 & ~n10268 ;
  assign n36601 = n4036 & ~n6765 ;
  assign n36602 = ~n5018 & n36601 ;
  assign n36603 = n6280 ^ n3881 ^ 1'b0 ;
  assign n36604 = ~n36602 & n36603 ;
  assign n36605 = n35083 & ~n36604 ;
  assign n36606 = n6794 & n10230 ;
  assign n36607 = ~n36041 & n36606 ;
  assign n36608 = n9343 & n28554 ;
  assign n36609 = n36608 ^ n18685 ^ 1'b0 ;
  assign n36610 = n8958 | n36609 ;
  assign n36611 = n31968 ^ n28387 ^ 1'b0 ;
  assign n36612 = n33794 & n36611 ;
  assign n36613 = ( n22051 & ~n34310 ) | ( n22051 & n36612 ) | ( ~n34310 & n36612 ) ;
  assign n36614 = n1430 | n8963 ;
  assign n36615 = n36614 ^ n13281 ^ 1'b0 ;
  assign n36616 = n367 & n15928 ;
  assign n36617 = n7080 & n36616 ;
  assign n36618 = ~n16726 & n17643 ;
  assign n36619 = n16268 ^ n15406 ^ 1'b0 ;
  assign n36620 = n36618 & n36619 ;
  assign n36621 = ~n36617 & n36620 ;
  assign n36622 = ~n33226 & n36621 ;
  assign n36623 = n4937 | n22470 ;
  assign n36624 = n9555 ^ n8285 ^ 1'b0 ;
  assign n36625 = n13568 | n36624 ;
  assign n36626 = n36625 ^ n19088 ^ 1'b0 ;
  assign n36627 = n15690 & n36626 ;
  assign n36628 = n32246 ^ n16421 ^ n489 ;
  assign n36629 = n1636 & n4256 ;
  assign n36630 = ~n4346 & n36629 ;
  assign n36633 = n4997 ^ n345 ^ 1'b0 ;
  assign n36634 = n27980 & n36633 ;
  assign n36631 = n6858 & ~n7007 ;
  assign n36632 = ( n9002 & n14087 ) | ( n9002 & ~n36631 ) | ( n14087 & ~n36631 ) ;
  assign n36635 = n36634 ^ n36632 ^ n13550 ;
  assign n36636 = n8685 ^ n4741 ^ n896 ;
  assign n36637 = n36636 ^ n6017 ^ 1'b0 ;
  assign n36638 = n1848 ^ n1356 ^ 1'b0 ;
  assign n36639 = n36637 & n36638 ;
  assign n36640 = n36639 ^ n31422 ^ n23893 ;
  assign n36641 = n14061 ^ n837 ^ 1'b0 ;
  assign n36642 = n32859 ^ n17858 ^ 1'b0 ;
  assign n36643 = n2028 | n36642 ;
  assign n36644 = n36643 ^ n8283 ^ 1'b0 ;
  assign n36645 = n36641 | n36644 ;
  assign n36646 = ~n21998 & n24527 ;
  assign n36647 = ( n2502 & n17369 ) | ( n2502 & n22718 ) | ( n17369 & n22718 ) ;
  assign n36648 = ~n6836 & n36647 ;
  assign n36651 = ~n9790 & n17234 ;
  assign n36649 = n29457 ^ n9943 ^ 1'b0 ;
  assign n36650 = n25069 & n36649 ;
  assign n36652 = n36651 ^ n36650 ^ 1'b0 ;
  assign n36653 = n20410 & n36652 ;
  assign n36654 = n9193 & n25391 ;
  assign n36655 = ~n6647 & n17936 ;
  assign n36656 = n15906 & n36655 ;
  assign n36659 = n6834 ^ n899 ^ 1'b0 ;
  assign n36657 = n11070 ^ n6058 ^ 1'b0 ;
  assign n36658 = n15440 & ~n36657 ;
  assign n36660 = n36659 ^ n36658 ^ n3158 ;
  assign n36661 = ( n7467 & n36472 ) | ( n7467 & n36660 ) | ( n36472 & n36660 ) ;
  assign n36662 = n7953 | n16446 ;
  assign n36663 = n124 & ~n36662 ;
  assign n36664 = ( n20740 & n28066 ) | ( n20740 & ~n36663 ) | ( n28066 & ~n36663 ) ;
  assign n36666 = n15782 | n23389 ;
  assign n36667 = n21872 & ~n36666 ;
  assign n36665 = n6455 & n12718 ;
  assign n36668 = n36667 ^ n36665 ^ 1'b0 ;
  assign n36670 = ( ~n1877 & n5394 ) | ( ~n1877 & n19853 ) | ( n5394 & n19853 ) ;
  assign n36669 = n12642 ^ n7234 ^ 1'b0 ;
  assign n36671 = n36670 ^ n36669 ^ 1'b0 ;
  assign n36672 = n23115 ^ n12576 ^ 1'b0 ;
  assign n36673 = n28273 & n36672 ;
  assign n36674 = ~n4111 & n6164 ;
  assign n36675 = n7784 ^ n2183 ^ 1'b0 ;
  assign n36676 = n16559 & ~n36675 ;
  assign n36677 = n5091 & n18063 ;
  assign n36678 = ~n36676 & n36677 ;
  assign n36679 = n7248 & n25089 ;
  assign n36680 = ~n14785 & n36679 ;
  assign n36681 = n15407 ^ n3519 ^ n1539 ;
  assign n36682 = n12950 & ~n30611 ;
  assign n36683 = n26787 & n36682 ;
  assign n36684 = n36681 & n36683 ;
  assign n36685 = n34749 ^ n5591 ^ 1'b0 ;
  assign n36686 = n4461 | n10852 ;
  assign n36687 = n1697 & ~n36686 ;
  assign n36688 = n25195 & ~n36687 ;
  assign n36689 = n5721 & n36688 ;
  assign n36690 = n30943 | n32226 ;
  assign n36691 = n15198 ^ n1014 ^ 1'b0 ;
  assign n36692 = n26983 ^ n10149 ^ n3307 ;
  assign n36693 = n5308 | n36692 ;
  assign n36694 = n36693 ^ n17319 ^ 1'b0 ;
  assign n36695 = ~n27071 & n36694 ;
  assign n36696 = n8419 ^ n3333 ^ 1'b0 ;
  assign n36697 = n21239 & n36696 ;
  assign n36698 = n27775 ^ n13304 ^ 1'b0 ;
  assign n36699 = n10296 | n36698 ;
  assign n36702 = ~n9017 & n23546 ;
  assign n36703 = n30508 & n36702 ;
  assign n36700 = n23958 & ~n27407 ;
  assign n36701 = n29671 & n36700 ;
  assign n36704 = n36703 ^ n36701 ^ 1'b0 ;
  assign n36705 = n8604 | n12038 ;
  assign n36706 = n36705 ^ n35005 ^ 1'b0 ;
  assign n36707 = n7399 ^ n782 ^ 1'b0 ;
  assign n36708 = n12338 & n26697 ;
  assign n36709 = n36707 & n36708 ;
  assign n36710 = n10288 & ~n36709 ;
  assign n36711 = ~n36706 & n36710 ;
  assign n36712 = n10497 & ~n18270 ;
  assign n36713 = ~n18328 & n36712 ;
  assign n36714 = n11682 & n36713 ;
  assign n36715 = n3904 & n5151 ;
  assign n36716 = n14343 & n36715 ;
  assign n36717 = n20798 ^ n10620 ^ 1'b0 ;
  assign n36718 = n19182 & n36717 ;
  assign n36719 = n3535 ^ n1862 ^ n481 ;
  assign n36720 = n36719 ^ n2218 ^ 1'b0 ;
  assign n36721 = n36361 | n36720 ;
  assign n36722 = n19881 & ~n36721 ;
  assign n36723 = n36722 ^ n12541 ^ n372 ;
  assign n36725 = ( n11287 & n17759 ) | ( n11287 & n26340 ) | ( n17759 & n26340 ) ;
  assign n36724 = n13389 | n34627 ;
  assign n36726 = n36725 ^ n36724 ^ 1'b0 ;
  assign n36727 = n27832 ^ n7947 ^ 1'b0 ;
  assign n36728 = n11295 & ~n36727 ;
  assign n36729 = ~n2826 & n27545 ;
  assign n36730 = n32233 ^ n23944 ^ 1'b0 ;
  assign n36731 = ~n1889 & n25101 ;
  assign n36732 = n6559 & n13451 ;
  assign n36733 = n36732 ^ n7586 ^ 1'b0 ;
  assign n36734 = n36731 & n36733 ;
  assign n36736 = n12049 & ~n23778 ;
  assign n36735 = n25138 | n35312 ;
  assign n36737 = n36736 ^ n36735 ^ 1'b0 ;
  assign n36738 = n8312 & n31493 ;
  assign n36739 = ~n8420 & n30097 ;
  assign n36740 = ~n36738 & n36739 ;
  assign n36741 = ~n12930 & n16627 ;
  assign n36742 = ~n2346 & n17881 ;
  assign n36743 = n18031 | n27923 ;
  assign n36744 = n9090 | n36743 ;
  assign n36745 = n25852 ^ n3358 ^ 1'b0 ;
  assign n36746 = n3665 & ~n23150 ;
  assign n36747 = n9522 | n9544 ;
  assign n36748 = n36747 ^ n35267 ^ n26298 ;
  assign n36749 = ( n4356 & n4525 ) | ( n4356 & ~n28764 ) | ( n4525 & ~n28764 ) ;
  assign n36750 = n36026 ^ n14891 ^ 1'b0 ;
  assign n36751 = n36749 & n36750 ;
  assign n36752 = n6277 | n36518 ;
  assign n36753 = n6870 & ~n36752 ;
  assign n36754 = n17939 ^ n14673 ^ x6 ;
  assign n36755 = ( n2152 & n12587 ) | ( n2152 & ~n36754 ) | ( n12587 & ~n36754 ) ;
  assign n36756 = n24208 ^ n4809 ^ 1'b0 ;
  assign n36757 = n12812 & ~n20689 ;
  assign n36758 = n11666 & ~n36757 ;
  assign n36759 = n36758 ^ n3794 ^ 1'b0 ;
  assign n36760 = n6833 | n17412 ;
  assign n36761 = n7197 & ~n7749 ;
  assign n36762 = n36761 ^ n21350 ^ n16727 ;
  assign n36763 = n36762 ^ n13755 ^ 1'b0 ;
  assign n36764 = n9700 & ~n36763 ;
  assign n36765 = n29007 ^ n16714 ^ 1'b0 ;
  assign n36766 = ~n17327 & n25441 ;
  assign n36767 = n12616 & n36766 ;
  assign n36768 = n34295 ^ n588 ^ 1'b0 ;
  assign n36769 = ~n20248 & n27721 ;
  assign n36770 = n36768 & n36769 ;
  assign n36771 = n23550 ^ n439 ^ 1'b0 ;
  assign n36772 = n3293 & ~n36771 ;
  assign n36773 = n7554 & ~n36772 ;
  assign n36774 = ~n1880 & n18888 ;
  assign n36775 = n36774 ^ n17549 ^ 1'b0 ;
  assign n36776 = n30404 & n36775 ;
  assign n36777 = n34575 ^ n33411 ^ 1'b0 ;
  assign n36778 = n19105 & n36777 ;
  assign n36779 = ~n4547 & n22833 ;
  assign n36780 = ~n1895 & n36779 ;
  assign n36781 = n949 & n32618 ;
  assign n36782 = n36781 ^ n373 ^ 1'b0 ;
  assign n36783 = n10071 & n28938 ;
  assign n36784 = n36782 & n36783 ;
  assign n36785 = ~n11331 & n12719 ;
  assign n36786 = ( n5580 & n6431 ) | ( n5580 & n29595 ) | ( n6431 & n29595 ) ;
  assign n36787 = ~n4025 & n14580 ;
  assign n36788 = n13850 | n24334 ;
  assign n36789 = n200 & ~n26511 ;
  assign n36791 = ~n51 & n2065 ;
  assign n36792 = n36791 ^ n10595 ^ 1'b0 ;
  assign n36790 = n26743 & ~n35605 ;
  assign n36793 = n36792 ^ n36790 ^ 1'b0 ;
  assign n36794 = ~n13302 & n20234 ;
  assign n36795 = n36794 ^ n12414 ^ 1'b0 ;
  assign n36796 = n18672 ^ n219 ^ 1'b0 ;
  assign n36797 = n1701 & n36796 ;
  assign n36798 = n5144 & ~n36797 ;
  assign n36799 = n19 & n17231 ;
  assign n36800 = n21715 | n27346 ;
  assign n36801 = n36800 ^ n9428 ^ 1'b0 ;
  assign n36802 = ( ~n4346 & n36799 ) | ( ~n4346 & n36801 ) | ( n36799 & n36801 ) ;
  assign n36803 = n4048 | n19440 ;
  assign n36804 = ~n220 & n3214 ;
  assign n36805 = ~n36075 & n36804 ;
  assign n36806 = n6021 & n36805 ;
  assign n36807 = n20959 ^ n4267 ^ 1'b0 ;
  assign n36808 = n16728 | n17187 ;
  assign n36809 = n36807 | n36808 ;
  assign n36810 = n6161 & ~n14894 ;
  assign n36811 = n231 & ~n12286 ;
  assign n36812 = n2621 & n36811 ;
  assign n36813 = ( ~n17611 & n31363 ) | ( ~n17611 & n36812 ) | ( n31363 & n36812 ) ;
  assign n36814 = n36813 ^ n1141 ^ 1'b0 ;
  assign n36815 = n36810 & ~n36814 ;
  assign n36816 = n16847 ^ n15377 ^ 1'b0 ;
  assign n36817 = n20719 & n36816 ;
  assign n36818 = n302 & ~n6769 ;
  assign n36819 = n2601 & n11826 ;
  assign n36820 = n36819 ^ n25175 ^ 1'b0 ;
  assign n36821 = n13877 & ~n36820 ;
  assign n36822 = ~n2802 & n9163 ;
  assign n36823 = n36822 ^ n17193 ^ 1'b0 ;
  assign n36824 = n2555 & ~n3298 ;
  assign n36825 = ( n4095 & ~n14253 ) | ( n4095 & n36824 ) | ( ~n14253 & n36824 ) ;
  assign n36827 = ~n2334 & n5644 ;
  assign n36828 = n36827 ^ n5111 ^ 1'b0 ;
  assign n36829 = n35862 & ~n36828 ;
  assign n36826 = ~n9204 & n20381 ;
  assign n36830 = n36829 ^ n36826 ^ 1'b0 ;
  assign n36831 = n347 & n13205 ;
  assign n36832 = n717 & n36831 ;
  assign n36833 = ( n14343 & n34099 ) | ( n14343 & ~n36832 ) | ( n34099 & ~n36832 ) ;
  assign n36834 = n8603 & n36833 ;
  assign n36835 = n15008 ^ n1005 ^ 1'b0 ;
  assign n36836 = n996 & n36835 ;
  assign n36837 = n2193 & n32643 ;
  assign n36838 = ~n16046 & n36837 ;
  assign n36839 = n8448 & ~n30461 ;
  assign n36840 = ~n24219 & n27732 ;
  assign n36841 = n23481 & ~n24898 ;
  assign n36842 = n36841 ^ n16328 ^ 1'b0 ;
  assign n36843 = n7681 & n17035 ;
  assign n36844 = n36843 ^ n3618 ^ 1'b0 ;
  assign n36845 = n1381 | n27173 ;
  assign n36846 = n36845 ^ n2379 ^ 1'b0 ;
  assign n36847 = n23283 ^ n9000 ^ 1'b0 ;
  assign n36848 = n1641 & ~n36847 ;
  assign n36849 = n15800 | n34975 ;
  assign n36850 = n17613 ^ n5799 ^ 1'b0 ;
  assign n36851 = n13566 | n36850 ;
  assign n36852 = ( n5821 & ~n6615 ) | ( n5821 & n21892 ) | ( ~n6615 & n21892 ) ;
  assign n36853 = n6338 | n6375 ;
  assign n36854 = n36852 & ~n36853 ;
  assign n36855 = n31503 ^ n20155 ^ 1'b0 ;
  assign n36856 = n26769 & ~n36855 ;
  assign n36857 = ~n298 & n6372 ;
  assign n36858 = ~n12294 & n36857 ;
  assign n36859 = ~n14248 & n29621 ;
  assign n36860 = ~n31676 & n36859 ;
  assign n36861 = ~n36858 & n36860 ;
  assign n36863 = n18881 ^ n7693 ^ 1'b0 ;
  assign n36862 = n6427 & n20163 ;
  assign n36864 = n36863 ^ n36862 ^ n28 ;
  assign n36865 = n13503 ^ n1570 ^ 1'b0 ;
  assign n36866 = ~n2353 & n36865 ;
  assign n36867 = n14135 ^ n8939 ^ 1'b0 ;
  assign n36868 = n3228 & n36867 ;
  assign n36869 = n21323 ^ n1539 ^ 1'b0 ;
  assign n36870 = ~n7327 & n36869 ;
  assign n36871 = n15360 ^ n2535 ^ 1'b0 ;
  assign n36872 = ~n12937 & n21239 ;
  assign n36873 = n36872 ^ n12302 ^ 1'b0 ;
  assign n36874 = ~n36871 & n36873 ;
  assign n36875 = n8582 & n14796 ;
  assign n36876 = n29583 ^ n9282 ^ 1'b0 ;
  assign n36877 = ~n28851 & n36876 ;
  assign n36878 = ~n15230 & n29918 ;
  assign n36879 = ~n29918 & n36878 ;
  assign n36880 = ~n18414 & n36879 ;
  assign n36881 = n3058 & n13885 ;
  assign n36883 = n27155 & n27723 ;
  assign n36882 = n1609 | n3305 ;
  assign n36884 = n36883 ^ n36882 ^ 1'b0 ;
  assign n36885 = n4039 | n36884 ;
  assign n36886 = n36881 & ~n36885 ;
  assign n36887 = n14828 & n27303 ;
  assign n36888 = n33813 ^ n19612 ^ 1'b0 ;
  assign n36889 = n17971 | n36888 ;
  assign n36890 = n36889 ^ n23817 ^ 1'b0 ;
  assign n36891 = n9584 & n36890 ;
  assign n36892 = n30072 ^ n19035 ^ 1'b0 ;
  assign n36893 = n9069 ^ n4089 ^ 1'b0 ;
  assign n36894 = n21064 & ~n36893 ;
  assign n36895 = n36894 ^ n13342 ^ 1'b0 ;
  assign n36896 = n6069 ^ n4750 ^ 1'b0 ;
  assign n36897 = ~n6008 & n36896 ;
  assign n36898 = ~n4183 & n36897 ;
  assign n36899 = n36898 ^ n8229 ^ 1'b0 ;
  assign n36900 = n21682 ^ n6566 ^ 1'b0 ;
  assign n36901 = ~n3533 & n36900 ;
  assign n36904 = n22865 ^ n5474 ^ 1'b0 ;
  assign n36905 = n18347 & n36904 ;
  assign n36902 = ( ~n8453 & n14994 ) | ( ~n8453 & n15479 ) | ( n14994 & n15479 ) ;
  assign n36903 = ~n17908 & n36902 ;
  assign n36906 = n36905 ^ n36903 ^ n21865 ;
  assign n36907 = n4298 & ~n7307 ;
  assign n36908 = n36907 ^ n3066 ^ 1'b0 ;
  assign n36909 = n1812 | n36908 ;
  assign n36910 = n13569 | n36909 ;
  assign n36911 = n36910 ^ n695 ^ 1'b0 ;
  assign n36912 = n22556 ^ n15885 ^ n15559 ;
  assign n36913 = n36911 & n36912 ;
  assign n36914 = n6790 ^ n2605 ^ 1'b0 ;
  assign n36915 = ~n13792 & n36914 ;
  assign n36916 = n11786 & n36915 ;
  assign n36917 = ~n3613 & n36916 ;
  assign n36918 = n8101 & ~n36917 ;
  assign n36919 = n10736 ^ n2802 ^ n356 ;
  assign n36920 = n15492 & n36919 ;
  assign n36921 = n36920 ^ n22860 ^ 1'b0 ;
  assign n36922 = n7046 ^ n6435 ^ 1'b0 ;
  assign n36923 = n11218 & ~n33542 ;
  assign n36924 = n36923 ^ n11120 ^ 1'b0 ;
  assign n36925 = n36924 ^ n28428 ^ 1'b0 ;
  assign n36927 = n10003 & n17964 ;
  assign n36928 = n36927 ^ n25567 ^ 1'b0 ;
  assign n36926 = n7464 & n23390 ;
  assign n36929 = n36928 ^ n36926 ^ 1'b0 ;
  assign n36930 = n13666 ^ n3122 ^ 1'b0 ;
  assign n36931 = n28098 & ~n36930 ;
  assign n36932 = ( n11497 & n27341 ) | ( n11497 & n28981 ) | ( n27341 & n28981 ) ;
  assign n36933 = n4086 & ~n24680 ;
  assign n36934 = n36933 ^ n22777 ^ 1'b0 ;
  assign n36935 = n28526 & n36934 ;
  assign n36936 = n8869 & n28591 ;
  assign n36937 = n6210 & n26716 ;
  assign n36938 = n27470 ^ n16003 ^ 1'b0 ;
  assign n36939 = n36937 & n36938 ;
  assign n36940 = n12513 & n34499 ;
  assign n36941 = n11187 & ~n35845 ;
  assign n36942 = n19799 ^ n4983 ^ n627 ;
  assign n36943 = ~n5721 & n5803 ;
  assign n36944 = n22469 & n36943 ;
  assign n36945 = n36944 ^ n26788 ^ n1900 ;
  assign n36955 = n12103 & n26194 ;
  assign n36956 = n12149 & n36955 ;
  assign n36957 = n18914 & ~n36956 ;
  assign n36958 = ~n15600 & n36957 ;
  assign n36959 = n11805 | n36958 ;
  assign n36960 = n20646 & ~n36959 ;
  assign n36961 = ( n1845 & n16786 ) | ( n1845 & n36960 ) | ( n16786 & n36960 ) ;
  assign n36948 = n27375 ^ n1627 ^ 1'b0 ;
  assign n36949 = n13699 ^ n2048 ^ 1'b0 ;
  assign n36950 = n25791 & n36949 ;
  assign n36951 = ~n8997 & n36950 ;
  assign n36952 = n36948 & n36951 ;
  assign n36953 = n9538 | n36952 ;
  assign n36954 = n3341 | n36953 ;
  assign n36962 = n36961 ^ n36954 ^ n9983 ;
  assign n36946 = n6769 & n12656 ;
  assign n36947 = n16548 | n36946 ;
  assign n36963 = n36962 ^ n36947 ^ 1'b0 ;
  assign n36964 = n36963 ^ n2605 ^ 1'b0 ;
  assign n36965 = n17627 & n36964 ;
  assign n36966 = ( n3466 & n9906 ) | ( n3466 & n21614 ) | ( n9906 & n21614 ) ;
  assign n36967 = n12850 | n36966 ;
  assign n36968 = ( n12288 & n14987 ) | ( n12288 & n36967 ) | ( n14987 & n36967 ) ;
  assign n36969 = n3246 & n36968 ;
  assign n36970 = n28725 & n36969 ;
  assign n36971 = n5598 | n24835 ;
  assign n36972 = n21074 ^ n1944 ^ 1'b0 ;
  assign n36973 = n23490 | n36972 ;
  assign n36974 = n36973 ^ n21636 ^ 1'b0 ;
  assign n36975 = n8608 & ~n19224 ;
  assign n36976 = n36975 ^ n720 ^ 1'b0 ;
  assign n36977 = ~n31503 & n36976 ;
  assign n36978 = ~n26211 & n36977 ;
  assign n36979 = n3082 & ~n36978 ;
  assign n36980 = n35608 ^ n5763 ^ n1119 ;
  assign n36981 = ~n12664 & n21283 ;
  assign n36982 = ~n15459 & n28634 ;
  assign n36983 = n36982 ^ n34308 ^ 1'b0 ;
  assign n36984 = n27321 | n31118 ;
  assign n36985 = n8633 & ~n36984 ;
  assign n36986 = ~n32971 & n36985 ;
  assign n36987 = ~n2282 & n2845 ;
  assign n36988 = n36987 ^ n13364 ^ 1'b0 ;
  assign n36989 = n14338 ^ n5821 ^ 1'b0 ;
  assign n36990 = n36988 | n36989 ;
  assign n36991 = n2212 ^ n657 ^ 1'b0 ;
  assign n36992 = ~n36990 & n36991 ;
  assign n36993 = n36992 ^ n8083 ^ 1'b0 ;
  assign n36994 = ~n36986 & n36993 ;
  assign n36995 = n20845 & ~n30322 ;
  assign n36996 = n2603 & n36995 ;
  assign n36997 = n36996 ^ n27638 ^ 1'b0 ;
  assign n36998 = n27705 | n36997 ;
  assign n37001 = n6492 ^ n4551 ^ 1'b0 ;
  assign n36999 = n17167 | n20095 ;
  assign n37000 = n36999 ^ n3075 ^ 1'b0 ;
  assign n37002 = n37001 ^ n37000 ^ n26441 ;
  assign n37003 = ( n5453 & ~n11414 ) | ( n5453 & n28476 ) | ( ~n11414 & n28476 ) ;
  assign n37004 = n23677 ^ n12030 ^ 1'b0 ;
  assign n37005 = n3665 & ~n37004 ;
  assign n37006 = ~n7921 & n14386 ;
  assign n37007 = n37006 ^ n17409 ^ 1'b0 ;
  assign n37008 = n13625 & n13897 ;
  assign n37009 = n37007 & ~n37008 ;
  assign n37010 = ~n37005 & n37009 ;
  assign n37011 = n8577 & n24926 ;
  assign n37012 = n37011 ^ n551 ^ 1'b0 ;
  assign n37013 = n6583 | n12125 ;
  assign n37014 = ~n14177 & n37013 ;
  assign n37015 = ~n1012 & n37014 ;
  assign n37016 = ~n3826 & n27629 ;
  assign n37017 = n37016 ^ n11060 ^ 1'b0 ;
  assign n37018 = n11193 & ~n27967 ;
  assign n37019 = n1000 & ~n2498 ;
  assign n37020 = ~n37018 & n37019 ;
  assign n37021 = n23146 ^ n13710 ^ 1'b0 ;
  assign n37022 = ~n37020 & n37021 ;
  assign n37023 = n7271 & ~n28505 ;
  assign n37024 = n1080 & n37023 ;
  assign n37025 = ~n25389 & n32798 ;
  assign n37026 = ( n2940 & n10840 ) | ( n2940 & n11572 ) | ( n10840 & n11572 ) ;
  assign n37027 = n13427 & n37026 ;
  assign n37028 = n24304 & n37027 ;
  assign n37029 = n34014 ^ n20430 ^ 1'b0 ;
  assign n37030 = ~n1085 & n11378 ;
  assign n37031 = n11552 & n37030 ;
  assign n37032 = n37031 ^ n11073 ^ n146 ;
  assign n37033 = ~n14184 & n31365 ;
  assign n37034 = n5819 | n6578 ;
  assign n37035 = n37034 ^ n26379 ^ 1'b0 ;
  assign n37036 = n4909 ^ n668 ^ 1'b0 ;
  assign n37037 = ~n2317 & n37036 ;
  assign n37038 = n11331 & n23242 ;
  assign n37039 = ~n37037 & n37038 ;
  assign n37040 = ~n23746 & n37039 ;
  assign n37041 = n4903 & n25960 ;
  assign n37042 = ~n31765 & n37041 ;
  assign n37043 = ~n22634 & n27733 ;
  assign n37044 = ~n3833 & n21635 ;
  assign n37045 = n25974 & n37044 ;
  assign n37046 = n6618 ^ n3298 ^ 1'b0 ;
  assign n37047 = n14462 | n37046 ;
  assign n37048 = n37047 ^ n12254 ^ 1'b0 ;
  assign n37049 = n37048 ^ n17326 ^ n11266 ;
  assign n37050 = n37049 ^ n19942 ^ 1'b0 ;
  assign n37051 = n23488 & ~n37050 ;
  assign n37052 = n30949 ^ n9413 ^ 1'b0 ;
  assign n37053 = n1584 | n28513 ;
  assign n37054 = n37052 | n37053 ;
  assign n37055 = ~n5747 & n28038 ;
  assign n37056 = ( n21816 & n31365 ) | ( n21816 & n37055 ) | ( n31365 & n37055 ) ;
  assign n37057 = n19131 | n22353 ;
  assign n37058 = ~n22784 & n24407 ;
  assign n37059 = n19680 & ~n26669 ;
  assign n37060 = n37059 ^ n772 ^ 1'b0 ;
  assign n37061 = n37060 ^ n34245 ^ 1'b0 ;
  assign n37062 = ~n28863 & n37061 ;
  assign n37063 = n23203 ^ n5242 ^ 1'b0 ;
  assign n37064 = n11644 & ~n35460 ;
  assign n37065 = n2359 & n37064 ;
  assign n37066 = ~n8027 & n27830 ;
  assign n37067 = n37066 ^ n7895 ^ 1'b0 ;
  assign n37068 = n17346 ^ n10945 ^ 1'b0 ;
  assign n37069 = ~n27 & n37068 ;
  assign n37070 = n27078 & n37069 ;
  assign n37071 = n22918 ^ n20917 ^ 1'b0 ;
  assign n37072 = n10387 | n37071 ;
  assign n37074 = ~n11897 & n24489 ;
  assign n37073 = n5350 & ~n6252 ;
  assign n37075 = n37074 ^ n37073 ^ 1'b0 ;
  assign n37076 = n37075 ^ n27493 ^ 1'b0 ;
  assign n37077 = n27467 ^ n3455 ^ 1'b0 ;
  assign n37078 = ~n6111 & n17479 ;
  assign n37079 = ~n905 & n37078 ;
  assign n37080 = n37079 ^ n8421 ^ 1'b0 ;
  assign n37081 = n5798 & ~n11504 ;
  assign n37082 = n37081 ^ n8728 ^ 1'b0 ;
  assign n37083 = ~n16010 & n32798 ;
  assign n37084 = n37083 ^ n2548 ^ 1'b0 ;
  assign n37085 = n37084 ^ n14520 ^ 1'b0 ;
  assign n37086 = n9719 | n15516 ;
  assign n37087 = n492 & ~n37086 ;
  assign n37088 = n20458 ^ n4946 ^ 1'b0 ;
  assign n37089 = ~n11235 & n37088 ;
  assign n37090 = ~n12746 & n37089 ;
  assign n37091 = n28931 ^ n10868 ^ n443 ;
  assign n37092 = n37091 ^ n16164 ^ n2022 ;
  assign n37093 = n20423 ^ n15 ^ 1'b0 ;
  assign n37094 = n20525 & n20988 ;
  assign n37095 = n8735 | n23880 ;
  assign n37096 = n6307 | n37095 ;
  assign n37097 = n1884 | n7889 ;
  assign n37098 = n9088 & ~n37097 ;
  assign n37099 = n4164 & ~n37098 ;
  assign n37100 = n11697 ^ n8703 ^ 1'b0 ;
  assign n37101 = n1079 | n33206 ;
  assign n37102 = n37100 & ~n37101 ;
  assign n37103 = ( n5219 & n37099 ) | ( n5219 & n37102 ) | ( n37099 & n37102 ) ;
  assign n37104 = n12036 | n14969 ;
  assign n37105 = n10726 | n12909 ;
  assign n37106 = n37105 ^ n24720 ^ 1'b0 ;
  assign n37107 = n8825 & ~n22969 ;
  assign n37108 = n37107 ^ n21226 ^ 1'b0 ;
  assign n37109 = n1929 & n18084 ;
  assign n37110 = n37109 ^ n16327 ^ 1'b0 ;
  assign n37111 = ( ~n17742 & n33389 ) | ( ~n17742 & n37110 ) | ( n33389 & n37110 ) ;
  assign n37112 = n23315 & ~n27550 ;
  assign n37113 = n14603 & ~n19769 ;
  assign n37114 = n813 & ~n1035 ;
  assign n37115 = n37114 ^ n2321 ^ 1'b0 ;
  assign n37116 = n7397 & ~n37115 ;
  assign n37117 = ~n7259 & n37116 ;
  assign n37118 = n459 | n3405 ;
  assign n37119 = n37118 ^ n11783 ^ 1'b0 ;
  assign n37120 = n7665 & n37119 ;
  assign n37121 = ~n11220 & n37120 ;
  assign n37122 = n37121 ^ n33792 ^ 1'b0 ;
  assign n37123 = n2122 & ~n37122 ;
  assign n37124 = n37123 ^ n2922 ^ 1'b0 ;
  assign n37125 = ~n18004 & n37124 ;
  assign n37126 = n19280 & ~n37125 ;
  assign n37128 = n27407 & ~n27470 ;
  assign n37127 = ~n18202 & n31577 ;
  assign n37129 = n37128 ^ n37127 ^ 1'b0 ;
  assign n37130 = n725 & ~n3665 ;
  assign n37131 = n37130 ^ n10978 ^ 1'b0 ;
  assign n37132 = n25075 ^ n21830 ^ 1'b0 ;
  assign n37133 = n17084 & ~n37132 ;
  assign n37134 = ( n1329 & n21259 ) | ( n1329 & ~n24182 ) | ( n21259 & ~n24182 ) ;
  assign n37135 = n17584 ^ n600 ^ 1'b0 ;
  assign n37136 = n37135 ^ n14022 ^ n10886 ;
  assign n37137 = n6492 & n12082 ;
  assign n37138 = n37137 ^ n16188 ^ 1'b0 ;
  assign n37139 = n27998 ^ n10232 ^ 1'b0 ;
  assign n37140 = n315 & ~n37139 ;
  assign n37141 = n11550 ^ n8903 ^ 1'b0 ;
  assign n37142 = n37140 & ~n37141 ;
  assign n37143 = ~n15290 & n37142 ;
  assign n37144 = n37143 ^ n4254 ^ 1'b0 ;
  assign n37145 = n8681 & ~n9266 ;
  assign n37146 = n2283 & n37145 ;
  assign n37147 = n11369 & ~n33482 ;
  assign n37148 = ( n5328 & n10094 ) | ( n5328 & n28113 ) | ( n10094 & n28113 ) ;
  assign n37150 = n12059 ^ n2114 ^ 1'b0 ;
  assign n37149 = n2055 & ~n2773 ;
  assign n37151 = n37150 ^ n37149 ^ 1'b0 ;
  assign n37152 = n3201 & ~n13963 ;
  assign n37153 = n31623 & ~n37152 ;
  assign n37154 = ( n17284 & n17625 ) | ( n17284 & ~n27030 ) | ( n17625 & ~n27030 ) ;
  assign n37155 = ~n11959 & n20157 ;
  assign n37156 = n8652 ^ n1517 ^ 1'b0 ;
  assign n37157 = ~n36304 & n37156 ;
  assign n37158 = n2273 | n8787 ;
  assign n37159 = n23762 ^ n23395 ^ 1'b0 ;
  assign n37160 = n7368 ^ n4973 ^ n4106 ;
  assign n37161 = n37160 ^ n12595 ^ 1'b0 ;
  assign n37162 = n21468 | n37161 ;
  assign n37163 = ( n1247 & n11123 ) | ( n1247 & ~n22524 ) | ( n11123 & ~n22524 ) ;
  assign n37164 = n2133 & ~n5448 ;
  assign n37165 = n8459 & n37164 ;
  assign n37166 = n7808 | n37165 ;
  assign n37167 = n37166 ^ n6749 ^ 1'b0 ;
  assign n37168 = n368 | n16010 ;
  assign n37169 = n317 & ~n13371 ;
  assign n37170 = n26474 & n37169 ;
  assign n37171 = n37170 ^ n7739 ^ 1'b0 ;
  assign n37172 = ~n2967 & n12713 ;
  assign n37173 = n37172 ^ n5474 ^ 1'b0 ;
  assign n37174 = n4007 | n29317 ;
  assign n37175 = n24594 & n37174 ;
  assign n37176 = n2747 | n28612 ;
  assign n37177 = n14825 ^ n546 ^ 1'b0 ;
  assign n37178 = ~n13129 & n37177 ;
  assign n37179 = n5948 | n12513 ;
  assign n37180 = ~n18199 & n28199 ;
  assign n37181 = n37179 | n37180 ;
  assign n37182 = n4159 & ~n35587 ;
  assign n37183 = n1150 | n21569 ;
  assign n37184 = n37183 ^ n4420 ^ 1'b0 ;
  assign n37185 = ~n1069 & n17366 ;
  assign n37186 = n14107 & n36011 ;
  assign n37187 = ~n8295 & n37186 ;
  assign n37188 = n6191 | n7909 ;
  assign n37189 = ( n186 & n25196 ) | ( n186 & ~n37188 ) | ( n25196 & ~n37188 ) ;
  assign n37190 = n28348 ^ n6040 ^ 1'b0 ;
  assign n37191 = n24861 & ~n37190 ;
  assign n37192 = ~n1229 & n37191 ;
  assign n37193 = n17309 | n37192 ;
  assign n37194 = n35048 | n37193 ;
  assign n37195 = n4164 & ~n37194 ;
  assign n37198 = n27498 ^ n12115 ^ 1'b0 ;
  assign n37199 = n6271 | n37198 ;
  assign n37196 = n3280 & ~n32051 ;
  assign n37197 = n37196 ^ n17773 ^ 1'b0 ;
  assign n37200 = n37199 ^ n37197 ^ n23373 ;
  assign n37201 = n26850 & ~n37200 ;
  assign n37202 = n20163 & ~n32004 ;
  assign n37203 = n423 & n28047 ;
  assign n37204 = n26435 | n26983 ;
  assign n37205 = n21277 ^ n13308 ^ n2382 ;
  assign n37206 = n5372 & n13126 ;
  assign n37207 = n2350 | n9500 ;
  assign n37208 = n3428 & n4034 ;
  assign n37209 = n37208 ^ n5871 ^ 1'b0 ;
  assign n37210 = n16630 & ~n35744 ;
  assign n37211 = n18152 & ~n37210 ;
  assign n37212 = n3477 | n9613 ;
  assign n37213 = n37212 ^ n19 ^ 1'b0 ;
  assign n37214 = n37213 ^ n10436 ^ 1'b0 ;
  assign n37215 = n9577 & n23553 ;
  assign n37216 = n37215 ^ n17353 ^ 1'b0 ;
  assign n37217 = ~n588 & n5288 ;
  assign n37218 = ~n5288 & n37217 ;
  assign n37219 = n37216 & ~n37218 ;
  assign n37220 = ~n37216 & n37219 ;
  assign n37221 = n20014 ^ n19685 ^ 1'b0 ;
  assign n37222 = n1360 & ~n6082 ;
  assign n37223 = n37222 ^ n4380 ^ 1'b0 ;
  assign n37224 = n18359 | n37223 ;
  assign n37225 = n22418 ^ n10066 ^ 1'b0 ;
  assign n37226 = n23287 | n37225 ;
  assign n37227 = ~n17427 & n19172 ;
  assign n37228 = ~n1469 & n37227 ;
  assign n37229 = ( n34344 & n37226 ) | ( n34344 & ~n37228 ) | ( n37226 & ~n37228 ) ;
  assign n37230 = n1176 ^ n421 ^ 1'b0 ;
  assign n37231 = n16837 | n37230 ;
  assign n37232 = n37231 ^ n33262 ^ 1'b0 ;
  assign n37233 = n37232 ^ n14087 ^ n3035 ;
  assign n37234 = n3893 & ~n24305 ;
  assign n37235 = n37234 ^ n11095 ^ 1'b0 ;
  assign n37236 = n26052 ^ n21924 ^ 1'b0 ;
  assign n37237 = n6860 & ~n11954 ;
  assign n37238 = n37237 ^ n35648 ^ 1'b0 ;
  assign n37239 = n23426 & n25501 ;
  assign n37240 = n37239 ^ n14057 ^ 1'b0 ;
  assign n37241 = n3114 & ~n37240 ;
  assign n37242 = n13055 & ~n33470 ;
  assign n37243 = n37242 ^ n17124 ^ 1'b0 ;
  assign n37244 = n36099 ^ n2934 ^ 1'b0 ;
  assign n37245 = ~n17169 & n17176 ;
  assign n37246 = n5974 & n37245 ;
  assign n37247 = n17548 & ~n37246 ;
  assign n37248 = n14082 & n29854 ;
  assign n37249 = n37248 ^ n1267 ^ 1'b0 ;
  assign n37250 = ( n465 & n29598 ) | ( n465 & n37249 ) | ( n29598 & n37249 ) ;
  assign n37251 = n2802 | n16740 ;
  assign n37252 = n6257 & ~n37251 ;
  assign n37253 = n15680 ^ n5438 ^ 1'b0 ;
  assign n37254 = n29490 & ~n37253 ;
  assign n37255 = n37254 ^ n3574 ^ 1'b0 ;
  assign n37256 = ~n13238 & n23075 ;
  assign n37257 = n37255 & n37256 ;
  assign n37258 = n31834 ^ n3355 ^ 1'b0 ;
  assign n37259 = n24930 | n37258 ;
  assign n37260 = n21905 & ~n37259 ;
  assign n37261 = n6322 & n35124 ;
  assign n37262 = n24313 & ~n37261 ;
  assign n37263 = ~n2609 & n37262 ;
  assign n37264 = ( n27687 & n35505 ) | ( n27687 & n36639 ) | ( n35505 & n36639 ) ;
  assign n37265 = n18563 ^ n7509 ^ 1'b0 ;
  assign n37266 = n37264 | n37265 ;
  assign n37267 = n7987 ^ n1010 ^ 1'b0 ;
  assign n37268 = n23619 & ~n37267 ;
  assign n37269 = n2340 & n37268 ;
  assign n37270 = n15999 & ~n37269 ;
  assign n37271 = n21461 & n37270 ;
  assign n37272 = n37271 ^ n9892 ^ 1'b0 ;
  assign n37273 = n1625 & n21353 ;
  assign n37274 = n37273 ^ n32848 ^ 1'b0 ;
  assign n37275 = n695 | n5874 ;
  assign n37276 = n5538 | n15867 ;
  assign n37277 = n1273 & ~n37276 ;
  assign n37278 = n37275 & ~n37277 ;
  assign n37279 = ~n20144 & n37278 ;
  assign n37280 = n37279 ^ n34179 ^ 1'b0 ;
  assign n37281 = ~n20510 & n35743 ;
  assign n37282 = n18146 ^ n11973 ^ 1'b0 ;
  assign n37283 = n5957 & ~n37282 ;
  assign n37284 = n23040 & ~n37283 ;
  assign n37285 = ~n12640 & n24587 ;
  assign n37286 = n9632 ^ n3958 ^ 1'b0 ;
  assign n37287 = n31397 | n37286 ;
  assign n37288 = n37287 ^ n25399 ^ 1'b0 ;
  assign n37289 = n28260 & n37288 ;
  assign n37290 = ~n192 & n18232 ;
  assign n37291 = ~n10352 & n37290 ;
  assign n37292 = n37291 ^ n22984 ^ 1'b0 ;
  assign n37293 = n15876 | n37292 ;
  assign n37294 = ~n12935 & n15659 ;
  assign n37295 = n37294 ^ n33239 ^ 1'b0 ;
  assign n37296 = ( n31061 & ~n37293 ) | ( n31061 & n37295 ) | ( ~n37293 & n37295 ) ;
  assign n37297 = n26321 & n34166 ;
  assign n37298 = n29730 ^ n17079 ^ 1'b0 ;
  assign n37299 = ~n6312 & n25451 ;
  assign n37300 = ~n30744 & n37299 ;
  assign n37301 = n14498 ^ n6182 ^ 1'b0 ;
  assign n37302 = n26550 & n37301 ;
  assign n37303 = n32958 ^ n12969 ^ 1'b0 ;
  assign n37304 = n37303 ^ n25972 ^ n7429 ;
  assign n37306 = n4231 & n29332 ;
  assign n37305 = ~n10877 & n16968 ;
  assign n37307 = n37306 ^ n37305 ^ 1'b0 ;
  assign n37308 = n12050 & ~n37307 ;
  assign n37309 = n19675 ^ n12502 ^ 1'b0 ;
  assign n37310 = n8738 & ~n15822 ;
  assign n37311 = n37310 ^ n14612 ^ 1'b0 ;
  assign n37312 = n11251 | n32432 ;
  assign n37313 = n37312 ^ n6878 ^ 1'b0 ;
  assign n37314 = n9465 | n37313 ;
  assign n37315 = n37314 ^ n13540 ^ 1'b0 ;
  assign n37316 = n1307 & ~n6948 ;
  assign n37317 = ~n10715 & n37316 ;
  assign n37318 = n18836 & ~n26258 ;
  assign n37319 = n11689 & n37318 ;
  assign n37320 = n14950 & ~n19411 ;
  assign n37321 = ~n11908 & n37320 ;
  assign n37322 = n19834 ^ n610 ^ 1'b0 ;
  assign n37323 = n7046 | n37322 ;
  assign n37324 = n20046 & n32755 ;
  assign n37325 = n31324 ^ n12224 ^ 1'b0 ;
  assign n37326 = n19166 | n22526 ;
  assign n37327 = n4347 & n13139 ;
  assign n37328 = ~n4006 & n37327 ;
  assign n37329 = n16297 & n23488 ;
  assign n37330 = n43 & n15839 ;
  assign n37331 = n37330 ^ n2547 ^ 1'b0 ;
  assign n37332 = ~n12052 & n37331 ;
  assign n37333 = n1501 | n3315 ;
  assign n37334 = n37333 ^ n14144 ^ 1'b0 ;
  assign n37335 = n21883 & n24047 ;
  assign n37336 = n3272 | n37335 ;
  assign n37337 = n14583 & n18582 ;
  assign n37338 = n16184 & n23912 ;
  assign n37339 = n2602 & ~n13356 ;
  assign n37340 = ( n9133 & n16558 ) | ( n9133 & ~n28779 ) | ( n16558 & ~n28779 ) ;
  assign n37341 = n6588 | n8460 ;
  assign n37342 = n37341 ^ n6378 ^ 1'b0 ;
  assign n37343 = n37342 ^ n30560 ^ 1'b0 ;
  assign n37344 = ~n8030 & n11813 ;
  assign n37346 = n26314 ^ n1395 ^ 1'b0 ;
  assign n37345 = n725 | n33432 ;
  assign n37347 = n37346 ^ n37345 ^ 1'b0 ;
  assign n37348 = n3135 | n10425 ;
  assign n37349 = n37348 ^ n7041 ^ 1'b0 ;
  assign n37350 = n20029 & n37349 ;
  assign n37351 = n34881 ^ n682 ^ 1'b0 ;
  assign n37352 = n15437 ^ n11196 ^ 1'b0 ;
  assign n37353 = ~n1198 & n14730 ;
  assign n37354 = n37353 ^ n6838 ^ 1'b0 ;
  assign n37355 = ~n9874 & n34003 ;
  assign n37356 = ( n6980 & n28610 ) | ( n6980 & ~n34350 ) | ( n28610 & ~n34350 ) ;
  assign n37357 = n13103 & n32929 ;
  assign n37358 = ~n2989 & n37357 ;
  assign n37359 = n8068 ^ n1951 ^ 1'b0 ;
  assign n37360 = n17714 ^ n15188 ^ 1'b0 ;
  assign n37361 = ~n14487 & n37360 ;
  assign n37362 = ~n3386 & n10218 ;
  assign n37363 = n474 & n37362 ;
  assign n37364 = ~n2547 & n16165 ;
  assign n37369 = n3693 | n4590 ;
  assign n37365 = ~n17195 & n29281 ;
  assign n37366 = n37365 ^ n695 ^ 1'b0 ;
  assign n37367 = n37366 ^ n20822 ^ 1'b0 ;
  assign n37368 = n8331 & n37367 ;
  assign n37370 = n37369 ^ n37368 ^ n36838 ;
  assign n37371 = n11117 & n29485 ;
  assign n37372 = n11959 & ~n37371 ;
  assign n37373 = n26604 ^ n914 ^ 1'b0 ;
  assign n37374 = n1252 & n16000 ;
  assign n37375 = n23633 & n37374 ;
  assign n37376 = ( ~n1207 & n3165 ) | ( ~n1207 & n9850 ) | ( n3165 & n9850 ) ;
  assign n37377 = n37376 ^ n17325 ^ 1'b0 ;
  assign n37378 = ~n37375 & n37377 ;
  assign n37379 = n19195 ^ n5475 ^ 1'b0 ;
  assign n37380 = n33125 ^ n23828 ^ 1'b0 ;
  assign n37381 = ~n9756 & n37380 ;
  assign n37382 = n35901 & ~n37381 ;
  assign n37383 = ~n18040 & n36098 ;
  assign n37384 = n4053 | n29031 ;
  assign n37385 = n37384 ^ n12072 ^ 1'b0 ;
  assign n37386 = n4390 | n20796 ;
  assign n37387 = n37386 ^ n2425 ^ 1'b0 ;
  assign n37388 = n5104 & ~n6535 ;
  assign n37389 = n17038 & n19980 ;
  assign n37390 = n4006 & ~n37389 ;
  assign n37391 = ~n996 & n37390 ;
  assign n37392 = n8338 & n10052 ;
  assign n37393 = n3295 & n12752 ;
  assign n37394 = ~n27565 & n34108 ;
  assign n37395 = n37393 & n37394 ;
  assign n37396 = ~n5264 & n35997 ;
  assign n37397 = n37396 ^ n808 ^ 1'b0 ;
  assign n37398 = ( ~n25708 & n32697 ) | ( ~n25708 & n37397 ) | ( n32697 & n37397 ) ;
  assign n37399 = n18714 ^ n160 ^ 1'b0 ;
  assign n37400 = n7270 ^ n5410 ^ 1'b0 ;
  assign n37401 = n565 & ~n37400 ;
  assign n37402 = n13462 ^ n708 ^ 1'b0 ;
  assign n37403 = ~n15174 & n37402 ;
  assign n37404 = n27923 | n31925 ;
  assign n37405 = n4615 & ~n37404 ;
  assign n37406 = n6672 ^ n3197 ^ 1'b0 ;
  assign n37407 = n6103 & n37406 ;
  assign n37408 = n14053 | n37407 ;
  assign n37409 = n37408 ^ n19904 ^ 1'b0 ;
  assign n37410 = n35932 | n37409 ;
  assign n37411 = ~n5562 & n32656 ;
  assign n37412 = n37411 ^ n25571 ^ 1'b0 ;
  assign n37413 = n1016 & n19921 ;
  assign n37414 = n22449 & n31787 ;
  assign n37415 = n10543 & n37414 ;
  assign n37416 = n4733 & ~n15449 ;
  assign n37417 = n37416 ^ n15817 ^ 1'b0 ;
  assign n37418 = n11164 & ~n26987 ;
  assign n37419 = n28154 & n37418 ;
  assign n37420 = n8723 & ~n37419 ;
  assign n37421 = n4946 ^ n4345 ^ 1'b0 ;
  assign n37422 = n1479 & n37421 ;
  assign n37423 = ( n3740 & n36835 ) | ( n3740 & n37422 ) | ( n36835 & n37422 ) ;
  assign n37424 = n21386 ^ n3740 ^ 1'b0 ;
  assign n37425 = n23688 & n37424 ;
  assign n37426 = n16156 & ~n25544 ;
  assign n37427 = n14238 & n37426 ;
  assign n37428 = n11683 & n30433 ;
  assign n37429 = n37427 & n37428 ;
  assign n37436 = ( n8232 & n11467 ) | ( n8232 & n28122 ) | ( n11467 & n28122 ) ;
  assign n37430 = n16533 | n27200 ;
  assign n37431 = n29052 ^ n1650 ^ 1'b0 ;
  assign n37432 = ~n37430 & n37431 ;
  assign n37433 = n10546 | n14899 ;
  assign n37434 = n28863 & ~n37433 ;
  assign n37435 = n37432 & ~n37434 ;
  assign n37437 = n37436 ^ n37435 ^ 1'b0 ;
  assign n37438 = n29058 | n37437 ;
  assign n37439 = n1207 & ~n37438 ;
  assign n37444 = n11885 & ~n22068 ;
  assign n37440 = n22017 ^ n6430 ^ n6347 ;
  assign n37441 = n12432 | n37440 ;
  assign n37442 = n16463 & ~n37441 ;
  assign n37443 = n7590 & n37442 ;
  assign n37445 = n37444 ^ n37443 ^ 1'b0 ;
  assign n37446 = n7986 & ~n10717 ;
  assign n37447 = n37446 ^ n33357 ^ 1'b0 ;
  assign n37448 = n8225 | n24454 ;
  assign n37449 = n29326 ^ n15240 ^ n1385 ;
  assign n37450 = n37448 | n37449 ;
  assign n37451 = n29907 ^ n14667 ^ n5518 ;
  assign n37452 = ~n7369 & n9979 ;
  assign n37453 = n14504 | n14610 ;
  assign n37454 = n6566 & n37453 ;
  assign n37455 = n37454 ^ n28211 ^ 1'b0 ;
  assign n37458 = n19178 ^ n961 ^ 1'b0 ;
  assign n37459 = ~n18602 & n37458 ;
  assign n37456 = n7765 & n30602 ;
  assign n37457 = n1528 & n37456 ;
  assign n37460 = n37459 ^ n37457 ^ 1'b0 ;
  assign n37461 = n28157 & n35990 ;
  assign n37462 = ~n737 & n2522 ;
  assign n37463 = n12588 & n37462 ;
  assign n37464 = n37463 ^ n30641 ^ 1'b0 ;
  assign n37465 = n19993 & n28424 ;
  assign n37466 = ~n16495 & n16867 ;
  assign n37467 = n7400 & ~n20964 ;
  assign n37468 = n37467 ^ n28208 ^ 1'b0 ;
  assign n37469 = n1099 & ~n11533 ;
  assign n37470 = n37469 ^ n17615 ^ 1'b0 ;
  assign n37471 = n37468 & n37470 ;
  assign n37472 = n1320 | n21619 ;
  assign n37473 = n37472 ^ n7721 ^ 1'b0 ;
  assign n37474 = n30346 ^ n5188 ^ 1'b0 ;
  assign n37475 = ~n592 & n37474 ;
  assign n37476 = ~n8793 & n17015 ;
  assign n37477 = n6589 & ~n9798 ;
  assign n37478 = n1886 & n18678 ;
  assign n37479 = ~n17209 & n37478 ;
  assign n37480 = n13505 ^ n7971 ^ n2134 ;
  assign n37481 = n37480 ^ n10737 ^ 1'b0 ;
  assign n37482 = n37481 ^ n33332 ^ 1'b0 ;
  assign n37483 = n22541 & n37216 ;
  assign n37484 = n5346 & n28490 ;
  assign n37485 = n11741 & n37484 ;
  assign n37486 = n37485 ^ n10311 ^ n961 ;
  assign n37487 = ( n4095 & ~n37483 ) | ( n4095 & n37486 ) | ( ~n37483 & n37486 ) ;
  assign n37488 = ( ~n10903 & n14391 ) | ( ~n10903 & n15276 ) | ( n14391 & n15276 ) ;
  assign n37489 = n31400 & ~n37488 ;
  assign n37490 = ~n18426 & n37489 ;
  assign n37491 = n24713 ^ n4275 ^ 1'b0 ;
  assign n37492 = n2389 & n37491 ;
  assign n37493 = n28999 & n34052 ;
  assign n37494 = n35168 ^ n32375 ^ n14246 ;
  assign n37495 = n19188 ^ n630 ^ 1'b0 ;
  assign n37496 = n320 & ~n37495 ;
  assign n37497 = n23516 ^ n14536 ^ 1'b0 ;
  assign n37498 = n37496 & ~n37497 ;
  assign n37499 = ~n15239 & n37498 ;
  assign n37500 = n10101 | n14503 ;
  assign n37501 = n37500 ^ n22728 ^ 1'b0 ;
  assign n37503 = n14106 & n35597 ;
  assign n37504 = n37503 ^ n14541 ^ 1'b0 ;
  assign n37502 = n1771 | n7311 ;
  assign n37505 = n37504 ^ n37502 ^ 1'b0 ;
  assign n37506 = n7499 & n12735 ;
  assign n37507 = n27080 ^ n6394 ^ n192 ;
  assign n37508 = n21420 ^ n10092 ^ 1'b0 ;
  assign n37510 = n22828 ^ n9356 ^ 1'b0 ;
  assign n37511 = ~n29445 & n37510 ;
  assign n37509 = n8344 & n21132 ;
  assign n37512 = n37511 ^ n37509 ^ 1'b0 ;
  assign n37513 = ~n1643 & n13096 ;
  assign n37514 = n25861 ^ n13069 ^ 1'b0 ;
  assign n37515 = n21998 | n37514 ;
  assign n37516 = n11378 | n37515 ;
  assign n37517 = n35152 ^ n2796 ^ 1'b0 ;
  assign n37518 = n5007 | n10347 ;
  assign n37519 = n37518 ^ n7493 ^ 1'b0 ;
  assign n37520 = n13893 | n37519 ;
  assign n37522 = n3891 & n4546 ;
  assign n37523 = n37522 ^ n30766 ^ 1'b0 ;
  assign n37521 = n13607 & ~n24253 ;
  assign n37524 = n37523 ^ n37521 ^ 1'b0 ;
  assign n37525 = n29744 ^ n5563 ^ 1'b0 ;
  assign n37526 = n567 & ~n18036 ;
  assign n37527 = n37526 ^ n17275 ^ 1'b0 ;
  assign n37528 = n37527 ^ n1049 ^ 1'b0 ;
  assign n37529 = n7067 | n23293 ;
  assign n37530 = n2101 & ~n37529 ;
  assign n37531 = ~n10656 & n29977 ;
  assign n37532 = ~n27057 & n37531 ;
  assign n37533 = n13068 ^ n6891 ^ 1'b0 ;
  assign n37534 = n22164 | n37471 ;
  assign n37535 = ~n5933 & n22881 ;
  assign n37536 = n13449 ^ n659 ^ 1'b0 ;
  assign n37537 = n14580 | n16136 ;
  assign n37538 = n14907 ^ n6711 ^ 1'b0 ;
  assign n37539 = n37537 & n37538 ;
  assign n37540 = ~n8405 & n37539 ;
  assign n37541 = ~n2092 & n2319 ;
  assign n37542 = n2092 & n37541 ;
  assign n37543 = n666 | n37542 ;
  assign n37544 = n37543 ^ n23067 ^ 1'b0 ;
  assign n37545 = ( n571 & ~n7715 ) | ( n571 & n26439 ) | ( ~n7715 & n26439 ) ;
  assign n37546 = n27093 ^ n11452 ^ 1'b0 ;
  assign n37547 = ( n9577 & ~n37545 ) | ( n9577 & n37546 ) | ( ~n37545 & n37546 ) ;
  assign n37548 = n3602 ^ n1808 ^ 1'b0 ;
  assign n37549 = ( n4346 & ~n8401 ) | ( n4346 & n37548 ) | ( ~n8401 & n37548 ) ;
  assign n37550 = n28958 ^ n8037 ^ 1'b0 ;
  assign n37551 = n28652 | n37550 ;
  assign n37552 = n29504 ^ n25704 ^ 1'b0 ;
  assign n37553 = n1191 & ~n3177 ;
  assign n37554 = n37552 & n37553 ;
  assign n37555 = n37554 ^ n27421 ^ 1'b0 ;
  assign n37556 = n26814 ^ n5223 ^ 1'b0 ;
  assign n37557 = n1896 & ~n9437 ;
  assign n37559 = ( ~n5583 & n23271 ) | ( ~n5583 & n30412 ) | ( n23271 & n30412 ) ;
  assign n37558 = n541 & n6170 ;
  assign n37560 = n37559 ^ n37558 ^ 1'b0 ;
  assign n37561 = ~n22050 & n23898 ;
  assign n37562 = n37561 ^ n3672 ^ 1'b0 ;
  assign n37563 = ~n3037 & n37562 ;
  assign n37564 = n2897 | n28421 ;
  assign n37565 = n37564 ^ n5116 ^ 1'b0 ;
  assign n37566 = n2044 & n5414 ;
  assign n37567 = n9674 & ~n37566 ;
  assign n37568 = n37565 | n37567 ;
  assign n37569 = n28168 & ~n37568 ;
  assign n37570 = ~n8608 & n12823 ;
  assign n37571 = ( n19440 & ~n29160 ) | ( n19440 & n35749 ) | ( ~n29160 & n35749 ) ;
  assign n37572 = n37570 | n37571 ;
  assign n37573 = n26667 ^ n11800 ^ 1'b0 ;
  assign n37574 = ~n5396 & n37573 ;
  assign n37575 = ( n1014 & n6705 ) | ( n1014 & n16453 ) | ( n6705 & n16453 ) ;
  assign n37576 = n15279 ^ n12234 ^ 1'b0 ;
  assign n37577 = n23092 | n37576 ;
  assign n37578 = n13573 | n37577 ;
  assign n37579 = n37575 | n37578 ;
  assign n37580 = ~n30696 & n37357 ;
  assign n37581 = n37580 ^ n30977 ^ 1'b0 ;
  assign n37582 = n11923 & n33196 ;
  assign n37583 = n37582 ^ n31466 ^ 1'b0 ;
  assign n37584 = n3036 & n16328 ;
  assign n37585 = ~n13204 & n28865 ;
  assign n37586 = n37584 & n37585 ;
  assign n37587 = n26480 ^ n2136 ^ 1'b0 ;
  assign n37588 = n13849 ^ n1724 ^ 1'b0 ;
  assign n37589 = n37588 ^ n20 ^ 1'b0 ;
  assign n37590 = n37587 & ~n37589 ;
  assign n37591 = n27651 ^ n194 ^ 1'b0 ;
  assign n37592 = n2743 & n17366 ;
  assign n37593 = n28368 & n37592 ;
  assign n37594 = n20080 ^ n16461 ^ 1'b0 ;
  assign n37595 = n4813 & ~n37594 ;
  assign n37596 = n19450 ^ n10022 ^ 1'b0 ;
  assign n37597 = n27456 ^ n14201 ^ 1'b0 ;
  assign n37598 = ( n3037 & ~n10665 ) | ( n3037 & n37597 ) | ( ~n10665 & n37597 ) ;
  assign n37599 = n20414 ^ n3271 ^ 1'b0 ;
  assign n37600 = n2139 & ~n8798 ;
  assign n37601 = n18177 ^ n12865 ^ 1'b0 ;
  assign n37602 = n25147 ^ n1192 ^ 1'b0 ;
  assign n37603 = n37601 & ~n37602 ;
  assign n37604 = n813 & n17115 ;
  assign n37605 = ~n6024 & n37604 ;
  assign n37606 = n11698 ^ n975 ^ 1'b0 ;
  assign n37607 = n37605 | n37606 ;
  assign n37608 = n16707 & n24405 ;
  assign n37609 = n37608 ^ n20386 ^ 1'b0 ;
  assign n37610 = n37609 ^ n10138 ^ 1'b0 ;
  assign n37611 = n37074 ^ n8776 ^ 1'b0 ;
  assign n37612 = n13410 & n37611 ;
  assign n37613 = n4017 & ~n14525 ;
  assign n37614 = n20808 & n37613 ;
  assign n37615 = n15792 & n37614 ;
  assign n37616 = n6136 ^ n3139 ^ 1'b0 ;
  assign n37617 = n8161 | n37616 ;
  assign n37618 = n33612 ^ n5803 ^ 1'b0 ;
  assign n37619 = n9627 | n37618 ;
  assign n37620 = n28537 ^ n18754 ^ 1'b0 ;
  assign n37625 = n760 & ~n2541 ;
  assign n37626 = ~n8076 & n26631 ;
  assign n37627 = ( n18154 & n37625 ) | ( n18154 & ~n37626 ) | ( n37625 & ~n37626 ) ;
  assign n37621 = n5453 & ~n24455 ;
  assign n37622 = n37621 ^ n4218 ^ 1'b0 ;
  assign n37623 = n37622 ^ n31315 ^ n29720 ;
  assign n37624 = n4857 & n37623 ;
  assign n37628 = n37627 ^ n37624 ^ 1'b0 ;
  assign n37629 = n21964 ^ n3171 ^ 1'b0 ;
  assign n37630 = ( n148 & n16906 ) | ( n148 & n37629 ) | ( n16906 & n37629 ) ;
  assign n37631 = n25791 ^ n4581 ^ 1'b0 ;
  assign n37632 = n16408 ^ n10297 ^ 1'b0 ;
  assign n37633 = n26665 & n37632 ;
  assign n37634 = n37633 ^ n18856 ^ 1'b0 ;
  assign n37635 = n557 | n6233 ;
  assign n37636 = n11458 & n13255 ;
  assign n37637 = ~n31166 & n37636 ;
  assign n37638 = n37637 ^ n9684 ^ 1'b0 ;
  assign n37639 = n3060 & n37638 ;
  assign n37640 = n14020 & ~n37639 ;
  assign n37641 = n23016 ^ n8301 ^ 1'b0 ;
  assign n37642 = n17083 | n37641 ;
  assign n37643 = ( n2074 & n35221 ) | ( n2074 & ~n37642 ) | ( n35221 & ~n37642 ) ;
  assign n37644 = n20443 ^ n4348 ^ 1'b0 ;
  assign n37645 = n36484 & ~n37644 ;
  assign n37646 = n911 | n13695 ;
  assign n37647 = n37646 ^ n13216 ^ 1'b0 ;
  assign n37648 = n7316 & n21326 ;
  assign n37649 = n24931 & ~n34109 ;
  assign n37650 = n28479 | n35554 ;
  assign n37651 = n5513 & n17845 ;
  assign n37652 = n37651 ^ n18834 ^ 1'b0 ;
  assign n37653 = n37652 ^ n4082 ^ 1'b0 ;
  assign n37654 = ~n37650 & n37653 ;
  assign n37655 = n3572 & ~n6989 ;
  assign n37656 = n37655 ^ n27192 ^ 1'b0 ;
  assign n37657 = n15876 | n37656 ;
  assign n37658 = ~n9663 & n33727 ;
  assign n37659 = n37658 ^ n15263 ^ n8368 ;
  assign n37660 = ( n10502 & n11520 ) | ( n10502 & ~n12507 ) | ( n11520 & ~n12507 ) ;
  assign n37661 = n37660 ^ n36368 ^ 1'b0 ;
  assign n37662 = n17749 | n37661 ;
  assign n37663 = n773 | n1469 ;
  assign n37664 = n37663 ^ n1680 ^ 1'b0 ;
  assign n37665 = n2574 & n37664 ;
  assign n37666 = n22668 & n37665 ;
  assign n37667 = ~n3541 & n37666 ;
  assign n37668 = n19680 | n37667 ;
  assign n37669 = ~n23018 & n37668 ;
  assign n37670 = n15210 & ~n16508 ;
  assign n37671 = n2023 & n5192 ;
  assign n37672 = n37671 ^ n3894 ^ 1'b0 ;
  assign n37673 = ~n34694 & n37672 ;
  assign n37674 = ~n5870 & n37673 ;
  assign n37675 = ( ~n4914 & n5968 ) | ( ~n4914 & n27271 ) | ( n5968 & n27271 ) ;
  assign n37676 = n20801 ^ n16083 ^ 1'b0 ;
  assign n37677 = n37675 & n37676 ;
  assign n37678 = ~n12426 & n14379 ;
  assign n37679 = n37678 ^ n29833 ^ 1'b0 ;
  assign n37684 = ~n299 & n21157 ;
  assign n37685 = n14351 | n37684 ;
  assign n37686 = n8971 & ~n37685 ;
  assign n37680 = n896 | n35051 ;
  assign n37681 = n30061 | n37680 ;
  assign n37682 = n14614 | n37681 ;
  assign n37683 = ( ~n480 & n22171 ) | ( ~n480 & n37682 ) | ( n22171 & n37682 ) ;
  assign n37687 = n37686 ^ n37683 ^ 1'b0 ;
  assign n37688 = ( n6578 & n18215 ) | ( n6578 & n19115 ) | ( n18215 & n19115 ) ;
  assign n37689 = ( n2491 & n2915 ) | ( n2491 & ~n37688 ) | ( n2915 & ~n37688 ) ;
  assign n37690 = n358 & ~n9970 ;
  assign n37691 = n34194 ^ n28533 ^ 1'b0 ;
  assign n37692 = n15478 | n37691 ;
  assign n37693 = n17065 | n17492 ;
  assign n37694 = n37693 ^ n15226 ^ 1'b0 ;
  assign n37695 = n37694 ^ n36285 ^ 1'b0 ;
  assign n37696 = ~n37692 & n37695 ;
  assign n37697 = n2950 | n3917 ;
  assign n37698 = n2219 | n37697 ;
  assign n37699 = n6762 ^ n4357 ^ 1'b0 ;
  assign n37700 = n37698 & n37699 ;
  assign n37701 = n35238 ^ n22046 ^ 1'b0 ;
  assign n37702 = n37700 & ~n37701 ;
  assign n37703 = n37702 ^ n2373 ^ 1'b0 ;
  assign n37704 = ~n6185 & n10345 ;
  assign n37705 = n4302 | n28195 ;
  assign n37706 = n1379 | n4612 ;
  assign n37707 = ~n798 & n37706 ;
  assign n37708 = n32723 ^ n19056 ^ 1'b0 ;
  assign n37709 = ~n1416 & n37708 ;
  assign n37710 = ~n4224 & n31455 ;
  assign n37711 = ~n25978 & n37710 ;
  assign n37712 = n35224 ^ n9085 ^ 1'b0 ;
  assign n37715 = ( n1918 & ~n9249 ) | ( n1918 & n15094 ) | ( ~n9249 & n15094 ) ;
  assign n37714 = n488 & n844 ;
  assign n37716 = n37715 ^ n37714 ^ 1'b0 ;
  assign n37717 = n37716 ^ n30521 ^ 1'b0 ;
  assign n37713 = n27599 ^ n582 ^ 1'b0 ;
  assign n37718 = n37717 ^ n37713 ^ 1'b0 ;
  assign n37719 = n6638 & n21457 ;
  assign n37720 = n30324 | n32948 ;
  assign n37721 = n13809 & ~n37720 ;
  assign n37722 = n32101 ^ n24518 ^ 1'b0 ;
  assign n37723 = ~n37721 & n37722 ;
  assign n37726 = n21333 ^ n3535 ^ 1'b0 ;
  assign n37724 = n12593 & n24271 ;
  assign n37725 = n37724 ^ n21150 ^ 1'b0 ;
  assign n37727 = n37726 ^ n37725 ^ n21627 ;
  assign n37728 = n1814 & ~n12784 ;
  assign n37729 = ~n37727 & n37728 ;
  assign n37730 = n37729 ^ n34009 ^ n15578 ;
  assign n37731 = ( n16779 & ~n23741 ) | ( n16779 & n35253 ) | ( ~n23741 & n35253 ) ;
  assign n37732 = n18628 ^ n12315 ^ n1758 ;
  assign n37733 = n630 | n37732 ;
  assign n37734 = n155 & n34846 ;
  assign n37735 = n25968 & n37734 ;
  assign n37736 = n19453 | n37735 ;
  assign n37737 = n1202 & n19319 ;
  assign n37738 = n11044 | n27303 ;
  assign n37740 = ~n1851 & n4871 ;
  assign n37741 = n37740 ^ n21155 ^ 1'b0 ;
  assign n37739 = n9245 & n15034 ;
  assign n37742 = n37741 ^ n37739 ^ 1'b0 ;
  assign n37743 = n13905 ^ n6273 ^ 1'b0 ;
  assign n37744 = n28199 & n37743 ;
  assign n37745 = n8952 ^ n767 ^ 1'b0 ;
  assign n37746 = ( n2688 & n8454 ) | ( n2688 & n14365 ) | ( n8454 & n14365 ) ;
  assign n37747 = n37746 ^ n425 ^ 1'b0 ;
  assign n37748 = n23152 | n37747 ;
  assign n37749 = n37748 ^ n8010 ^ 1'b0 ;
  assign n37750 = n24937 ^ n8973 ^ 1'b0 ;
  assign n37751 = n4315 & ~n37750 ;
  assign n37752 = n16844 & ~n29142 ;
  assign n37753 = n11484 & n32172 ;
  assign n37754 = n18135 & n37753 ;
  assign n37755 = n33710 & n37754 ;
  assign n37756 = n8702 ^ n7546 ^ 1'b0 ;
  assign n37757 = n37756 ^ n19999 ^ 1'b0 ;
  assign n37758 = ~n9970 & n37757 ;
  assign n37759 = n17015 ^ n14117 ^ 1'b0 ;
  assign n37760 = n37758 & ~n37759 ;
  assign n37761 = n14837 ^ n7929 ^ 1'b0 ;
  assign n37762 = n37760 & ~n37761 ;
  assign n37763 = n4022 & n26822 ;
  assign n37764 = n37763 ^ n4997 ^ 1'b0 ;
  assign n37765 = n37764 ^ n5467 ^ 1'b0 ;
  assign n37766 = ( n260 & n3243 ) | ( n260 & n7526 ) | ( n3243 & n7526 ) ;
  assign n37767 = n22874 ^ n10736 ^ 1'b0 ;
  assign n37768 = n26765 ^ n24500 ^ 1'b0 ;
  assign n37769 = ~n37767 & n37768 ;
  assign n37770 = n37766 & ~n37769 ;
  assign n37771 = ( n15430 & n23905 ) | ( n15430 & ~n37770 ) | ( n23905 & ~n37770 ) ;
  assign n37772 = n20580 ^ n2114 ^ 1'b0 ;
  assign n37773 = n3374 & n37772 ;
  assign n37774 = n6080 ^ n4917 ^ 1'b0 ;
  assign n37775 = n37773 & n37774 ;
  assign n37776 = n1469 & ~n23587 ;
  assign n37777 = n37776 ^ n34561 ^ 1'b0 ;
  assign n37778 = n11244 ^ n4483 ^ 1'b0 ;
  assign n37779 = n37778 ^ n9523 ^ 1'b0 ;
  assign n37780 = n33162 & n37779 ;
  assign n37781 = ( n3479 & ~n3811 ) | ( n3479 & n8815 ) | ( ~n3811 & n8815 ) ;
  assign n37782 = n37781 ^ n13134 ^ 1'b0 ;
  assign n37783 = n37782 ^ n4857 ^ n593 ;
  assign n37784 = n37783 ^ n14951 ^ 1'b0 ;
  assign n37785 = ~n6216 & n37784 ;
  assign n37786 = ~n2277 & n37785 ;
  assign n37787 = ( n5151 & n8040 ) | ( n5151 & n16654 ) | ( n8040 & n16654 ) ;
  assign n37788 = n2403 & n29579 ;
  assign n37789 = n37788 ^ n34782 ^ 1'b0 ;
  assign n37791 = n12983 ^ n11973 ^ 1'b0 ;
  assign n37792 = ~n21302 & n37791 ;
  assign n37790 = ~n1089 & n12690 ;
  assign n37793 = n37792 ^ n37790 ^ 1'b0 ;
  assign n37794 = ~n17564 & n37793 ;
  assign n37795 = n11857 ^ n1600 ^ 1'b0 ;
  assign n37796 = n36389 & ~n37795 ;
  assign n37797 = n1668 & ~n3328 ;
  assign n37798 = ~n74 & n8570 ;
  assign n37799 = n19923 & n20035 ;
  assign n37800 = n22048 ^ n14810 ^ 1'b0 ;
  assign n37801 = n37799 & ~n37800 ;
  assign n37802 = ~n991 & n28672 ;
  assign n37803 = ~n996 & n37802 ;
  assign n37804 = n37803 ^ n34755 ^ 1'b0 ;
  assign n37805 = n8247 | n37804 ;
  assign n37806 = n34412 ^ n2097 ^ 1'b0 ;
  assign n37807 = n19393 | n37806 ;
  assign n37808 = n1887 & n9336 ;
  assign n37809 = n37808 ^ n9224 ^ n7697 ;
  assign n37810 = n24507 & n37809 ;
  assign n37811 = n37063 ^ n9970 ^ 1'b0 ;
  assign n37812 = n870 | n37811 ;
  assign n37813 = n1608 & ~n11312 ;
  assign n37814 = n37813 ^ n425 ^ 1'b0 ;
  assign n37815 = n14829 & n24913 ;
  assign n37816 = n37815 ^ n11849 ^ 1'b0 ;
  assign n37818 = ( n6704 & n10609 ) | ( n6704 & n36747 ) | ( n10609 & n36747 ) ;
  assign n37819 = n6084 | n37818 ;
  assign n37820 = n877 & ~n37819 ;
  assign n37817 = n511 & n37712 ;
  assign n37821 = n37820 ^ n37817 ^ 1'b0 ;
  assign n37822 = n2940 | n32227 ;
  assign n37824 = ( ~n401 & n1865 ) | ( ~n401 & n4059 ) | ( n1865 & n4059 ) ;
  assign n37823 = n227 | n10656 ;
  assign n37825 = n37824 ^ n37823 ^ 1'b0 ;
  assign n37826 = n37825 ^ n16729 ^ 1'b0 ;
  assign n37827 = n4970 & n20625 ;
  assign n37828 = n8122 & ~n23039 ;
  assign n37829 = ~n20191 & n30848 ;
  assign n37830 = ~n37828 & n37829 ;
  assign n37831 = ~n7917 & n21675 ;
  assign n37832 = n17797 & n37831 ;
  assign n37833 = n5760 | n7804 ;
  assign n37834 = n34591 & ~n37833 ;
  assign n37835 = n19202 ^ n10085 ^ n7356 ;
  assign n37836 = n12612 ^ n333 ^ 1'b0 ;
  assign n37837 = ~n10232 & n37836 ;
  assign n37838 = n37837 ^ n6813 ^ 1'b0 ;
  assign n37839 = n37838 ^ n24686 ^ n21798 ;
  assign n37840 = ~n18770 & n25974 ;
  assign n37841 = n20202 & ~n22603 ;
  assign n37842 = n31 | n18392 ;
  assign n37843 = n37842 ^ n3292 ^ 1'b0 ;
  assign n37844 = n25960 ^ n1109 ^ 1'b0 ;
  assign n37845 = n34641 & ~n37844 ;
  assign n37846 = n9109 ^ n8693 ^ 1'b0 ;
  assign n37847 = ~n5174 & n17237 ;
  assign n37848 = ~n20257 & n32641 ;
  assign n37849 = n37847 & n37848 ;
  assign n37850 = n25902 | n29058 ;
  assign n37851 = n37850 ^ n23822 ^ 1'b0 ;
  assign n37852 = ( n4814 & ~n37849 ) | ( n4814 & n37851 ) | ( ~n37849 & n37851 ) ;
  assign n37853 = n28348 ^ n12836 ^ 1'b0 ;
  assign n37854 = n4366 & n37853 ;
  assign n37855 = n37854 ^ n4905 ^ 1'b0 ;
  assign n37856 = n6506 & ~n12930 ;
  assign n37857 = n24048 & ~n32227 ;
  assign n37858 = n14135 ^ n820 ^ 1'b0 ;
  assign n37859 = n9166 | n37858 ;
  assign n37860 = n37859 ^ n34995 ^ n2155 ;
  assign n37861 = n31119 & ~n37860 ;
  assign n37862 = n1485 & n37861 ;
  assign n37863 = ~n37857 & n37862 ;
  assign n37864 = n3584 ^ n3486 ^ 1'b0 ;
  assign n37865 = n37303 ^ n24790 ^ 1'b0 ;
  assign n37866 = ~n25553 & n37865 ;
  assign n37867 = ~n3498 & n20577 ;
  assign n37868 = n34826 | n36017 ;
  assign n37869 = n7685 ^ n2140 ^ 1'b0 ;
  assign n37870 = n37869 ^ n36967 ^ 1'b0 ;
  assign n37871 = n12322 ^ n8286 ^ 1'b0 ;
  assign n37872 = ~n37870 & n37871 ;
  assign n37873 = n31477 ^ n27180 ^ 1'b0 ;
  assign n37874 = n37872 & n37873 ;
  assign n37875 = n26010 ^ n9267 ^ 1'b0 ;
  assign n37876 = n27940 & ~n37875 ;
  assign n37877 = n4104 & ~n4650 ;
  assign n37878 = ~n9586 & n37877 ;
  assign n37879 = n23798 | n37878 ;
  assign n37880 = n18236 | n33936 ;
  assign n37881 = n29840 | n37880 ;
  assign n37882 = n4290 | n8917 ;
  assign n37883 = ( n5708 & ~n14019 ) | ( n5708 & n37882 ) | ( ~n14019 & n37882 ) ;
  assign n37884 = n835 | n37883 ;
  assign n37885 = ~n22432 & n26745 ;
  assign n37886 = n959 | n3372 ;
  assign n37887 = n37886 ^ n3012 ^ 1'b0 ;
  assign n37888 = n17763 | n32879 ;
  assign n37889 = n37888 ^ n20095 ^ 1'b0 ;
  assign n37890 = n37889 ^ n29819 ^ n1920 ;
  assign n37891 = ~n475 & n17258 ;
  assign n37892 = ~n7655 & n37891 ;
  assign n37893 = n931 & n37892 ;
  assign n37894 = n36582 & ~n37893 ;
  assign n37895 = n3740 | n33269 ;
  assign n37896 = n24548 | n37895 ;
  assign n37897 = n37896 ^ n502 ^ 1'b0 ;
  assign n37898 = n4470 & n6610 ;
  assign n37899 = n33739 | n36713 ;
  assign n37900 = n24325 ^ n140 ^ 1'b0 ;
  assign n37901 = n21488 ^ n2539 ^ 1'b0 ;
  assign n37902 = n642 & ~n8664 ;
  assign n37903 = n23266 & n37902 ;
  assign n37904 = n9289 & n37903 ;
  assign n37905 = n37904 ^ n31269 ^ 1'b0 ;
  assign n37906 = n400 & ~n37905 ;
  assign n37907 = n16933 & n37906 ;
  assign n37908 = n37907 ^ n36082 ^ 1'b0 ;
  assign n37909 = ~n10809 & n21857 ;
  assign n37910 = n37909 ^ n502 ^ 1'b0 ;
  assign n37911 = ( n8927 & n14305 ) | ( n8927 & n27435 ) | ( n14305 & n27435 ) ;
  assign n37912 = n37911 ^ n14749 ^ 1'b0 ;
  assign n37913 = n13959 ^ n2776 ^ 1'b0 ;
  assign n37914 = n560 & n19038 ;
  assign n37916 = n4401 & ~n15200 ;
  assign n37915 = n6867 & n12322 ;
  assign n37917 = n37916 ^ n37915 ^ 1'b0 ;
  assign n37918 = n409 & n28365 ;
  assign n37919 = n860 & n37918 ;
  assign n37920 = n14798 & n16404 ;
  assign n37921 = ( n15872 & ~n19291 ) | ( n15872 & n24148 ) | ( ~n19291 & n24148 ) ;
  assign n37922 = n646 & n37921 ;
  assign n37923 = n23861 | n28381 ;
  assign n37924 = ~n2273 & n14374 ;
  assign n37925 = n37924 ^ n26744 ^ 1'b0 ;
  assign n37926 = ~n7640 & n23120 ;
  assign n37927 = n37926 ^ n26997 ^ 1'b0 ;
  assign n37928 = n12628 | n37927 ;
  assign n37929 = n5191 ^ n3173 ^ 1'b0 ;
  assign n37930 = n6020 & n36425 ;
  assign n37931 = n37930 ^ n4519 ^ 1'b0 ;
  assign n37932 = n1356 | n14614 ;
  assign n37933 = n37932 ^ n3118 ^ 1'b0 ;
  assign n37934 = n1493 | n5289 ;
  assign n37935 = n37933 | n37934 ;
  assign n37936 = ( n10015 & ~n10895 ) | ( n10015 & n37935 ) | ( ~n10895 & n37935 ) ;
  assign n37937 = n26926 ^ n3588 ^ 1'b0 ;
  assign n37938 = n8805 | n37937 ;
  assign n37939 = n29992 ^ n20509 ^ 1'b0 ;
  assign n37940 = n31856 & n37939 ;
  assign n37941 = n22341 & ~n29402 ;
  assign n37942 = n8321 ^ n4327 ^ 1'b0 ;
  assign n37943 = ~n18037 & n37942 ;
  assign n37944 = n10477 | n19903 ;
  assign n37945 = ~n5206 & n30848 ;
  assign n37946 = n37945 ^ n7193 ^ n4095 ;
  assign n37947 = n3530 ^ n896 ^ 1'b0 ;
  assign n37948 = ~n14439 & n32352 ;
  assign n37949 = n8001 | n37948 ;
  assign n37950 = n791 & ~n37949 ;
  assign n37951 = ~n934 & n5534 ;
  assign n37952 = ~n24228 & n26223 ;
  assign n37953 = n37952 ^ n18507 ^ 1'b0 ;
  assign n37954 = ~n37951 & n37953 ;
  assign n37955 = n5988 & ~n23395 ;
  assign n37956 = ~n11435 & n33508 ;
  assign n37957 = x10 & n3112 ;
  assign n37958 = n37957 ^ n22550 ^ 1'b0 ;
  assign n37959 = n23864 & n37958 ;
  assign n37960 = ~n2132 & n37959 ;
  assign n37961 = n37960 ^ n12116 ^ 1'b0 ;
  assign n37962 = ~n28698 & n37961 ;
  assign n37963 = n16860 ^ n12777 ^ 1'b0 ;
  assign n37964 = n445 ^ n342 ^ 1'b0 ;
  assign n37965 = ~n3595 & n37964 ;
  assign n37966 = n12450 & n37965 ;
  assign n37967 = ~n19902 & n37966 ;
  assign n37968 = n37967 ^ n16889 ^ 1'b0 ;
  assign n37969 = n15331 ^ n12990 ^ 1'b0 ;
  assign n37970 = n37969 ^ n10778 ^ 1'b0 ;
  assign n37971 = n23240 & n37970 ;
  assign n37972 = n870 & ~n37971 ;
  assign n37973 = ~n6750 & n6933 ;
  assign n37974 = ~n8490 & n12740 ;
  assign n37975 = ~n6378 & n37974 ;
  assign n37976 = n37975 ^ n18619 ^ n15616 ;
  assign n37977 = n3547 | n16010 ;
  assign n37978 = n7238 | n37977 ;
  assign n37979 = n37978 ^ n7388 ^ 1'b0 ;
  assign n37980 = n4718 | n16588 ;
  assign n37981 = n37980 ^ n3513 ^ 1'b0 ;
  assign n37982 = n20447 & n21114 ;
  assign n37983 = n4846 ^ n4641 ^ n2211 ;
  assign n37984 = n37983 ^ n25637 ^ n5872 ;
  assign n37985 = n15699 | n20242 ;
  assign n37986 = ~n2574 & n37985 ;
  assign n37987 = n37986 ^ n11559 ^ 1'b0 ;
  assign n37988 = n510 & n19201 ;
  assign n37989 = n37988 ^ n2389 ^ 1'b0 ;
  assign n37990 = n753 | n37989 ;
  assign n37991 = n5077 & ~n14384 ;
  assign n37992 = n11541 & n33630 ;
  assign n37993 = n37991 & n37992 ;
  assign n37994 = n165 & ~n16431 ;
  assign n37995 = n37994 ^ n423 ^ 1'b0 ;
  assign n37996 = n20001 & ~n37995 ;
  assign n37997 = n3643 & n27599 ;
  assign n37998 = n37997 ^ n10852 ^ 1'b0 ;
  assign n37999 = ~n10950 & n37998 ;
  assign n38000 = ~n24112 & n37999 ;
  assign n38001 = n4551 | n10538 ;
  assign n38002 = n36635 | n38001 ;
  assign n38003 = n27653 ^ n3112 ^ 1'b0 ;
  assign n38004 = n24326 ^ n5001 ^ 1'b0 ;
  assign n38005 = n38004 ^ n24587 ^ 1'b0 ;
  assign n38006 = n2408 & n38005 ;
  assign n38007 = ( n3331 & n38003 ) | ( n3331 & n38006 ) | ( n38003 & n38006 ) ;
  assign n38008 = n7134 & n25798 ;
  assign n38009 = n38008 ^ n28121 ^ n212 ;
  assign n38010 = ~n606 & n5849 ;
  assign n38011 = ~n14566 & n38010 ;
  assign n38012 = ~n5623 & n38011 ;
  assign n38013 = n4370 & ~n38012 ;
  assign n38014 = n38013 ^ n21969 ^ 1'b0 ;
  assign n38015 = n3992 ^ n1636 ^ 1'b0 ;
  assign n38016 = ~n13173 & n16117 ;
  assign n38017 = ~n38015 & n38016 ;
  assign n38018 = n13393 & ~n15607 ;
  assign n38019 = ~n7616 & n38018 ;
  assign n38020 = n7825 ^ n3954 ^ 1'b0 ;
  assign n38021 = n38020 ^ n1736 ^ 1'b0 ;
  assign n38022 = ( ~n3526 & n23962 ) | ( ~n3526 & n38021 ) | ( n23962 & n38021 ) ;
  assign n38023 = n3695 & ~n4095 ;
  assign n38024 = n21467 ^ n15087 ^ 1'b0 ;
  assign n38025 = ~n5355 & n38024 ;
  assign n38026 = n38025 ^ n35622 ^ n13929 ;
  assign n38027 = n34046 ^ n23104 ^ 1'b0 ;
  assign n38028 = n18679 | n38027 ;
  assign n38029 = n10803 & ~n15552 ;
  assign n38030 = ~n3762 & n27765 ;
  assign n38031 = n34628 ^ n9083 ^ 1'b0 ;
  assign n38032 = ( n565 & n6613 ) | ( n565 & ~n10475 ) | ( n6613 & ~n10475 ) ;
  assign n38033 = ~n17220 & n17774 ;
  assign n38034 = n10508 & n38033 ;
  assign n38035 = n2128 & n24524 ;
  assign n38036 = n38034 & n38035 ;
  assign n38039 = n2816 & n22379 ;
  assign n38038 = n8705 & n12322 ;
  assign n38040 = n38039 ^ n38038 ^ 1'b0 ;
  assign n38037 = ~n6590 & n37292 ;
  assign n38041 = n38040 ^ n38037 ^ 1'b0 ;
  assign n38042 = n16976 | n31365 ;
  assign n38043 = n38042 ^ n1852 ^ 1'b0 ;
  assign n38044 = n30917 & ~n38043 ;
  assign n38045 = n38041 & n38044 ;
  assign n38046 = n1119 & n16007 ;
  assign n38047 = n38046 ^ n15963 ^ 1'b0 ;
  assign n38048 = ( n1100 & n2288 ) | ( n1100 & n18703 ) | ( n2288 & n18703 ) ;
  assign n38049 = n4636 & n38048 ;
  assign n38050 = n38047 & n38049 ;
  assign n38051 = n10968 | n17341 ;
  assign n38052 = n13937 & ~n38051 ;
  assign n38053 = n3592 & n7565 ;
  assign n38054 = n3068 & ~n4447 ;
  assign n38055 = n38054 ^ n26837 ^ 1'b0 ;
  assign n38056 = ( ~n3488 & n12103 ) | ( ~n3488 & n38055 ) | ( n12103 & n38055 ) ;
  assign n38057 = n38053 & ~n38056 ;
  assign n38058 = n6351 ^ n4928 ^ 1'b0 ;
  assign n38059 = ~n10628 & n32399 ;
  assign n38060 = n7360 & n38059 ;
  assign n38061 = n22833 & n31656 ;
  assign n38063 = n11348 ^ n2199 ^ 1'b0 ;
  assign n38064 = n15607 ^ n14511 ^ 1'b0 ;
  assign n38065 = n38063 & n38064 ;
  assign n38062 = n4341 & n33647 ;
  assign n38066 = n38065 ^ n38062 ^ 1'b0 ;
  assign n38067 = n33485 ^ n1700 ^ n1327 ;
  assign n38068 = ~n5044 & n22357 ;
  assign n38069 = ~n24208 & n38068 ;
  assign n38070 = n38069 ^ n8457 ^ 1'b0 ;
  assign n38071 = n15463 | n35565 ;
  assign n38072 = n13454 ^ n5751 ^ 1'b0 ;
  assign n38073 = n22262 ^ n9792 ^ 1'b0 ;
  assign n38074 = n13414 & ~n38073 ;
  assign n38075 = n16621 ^ n11000 ^ 1'b0 ;
  assign n38076 = n18179 & n38075 ;
  assign n38077 = n11453 ^ n7369 ^ 1'b0 ;
  assign n38078 = n38077 ^ n9078 ^ n372 ;
  assign n38079 = n4859 ^ n1662 ^ 1'b0 ;
  assign n38081 = n28341 ^ n1381 ^ 1'b0 ;
  assign n38080 = n6274 & n31766 ;
  assign n38082 = n38081 ^ n38080 ^ 1'b0 ;
  assign n38083 = ~n15948 & n21171 ;
  assign n38084 = n21518 ^ n13998 ^ 1'b0 ;
  assign n38085 = ~n14598 & n38084 ;
  assign n38086 = ~n11597 & n38085 ;
  assign n38087 = n38086 ^ n14962 ^ 1'b0 ;
  assign n38088 = n38087 ^ n10389 ^ 1'b0 ;
  assign n38089 = n37885 ^ n22658 ^ 1'b0 ;
  assign n38090 = ~n38088 & n38089 ;
  assign n38091 = n3361 | n7486 ;
  assign n38092 = n38091 ^ n2141 ^ 1'b0 ;
  assign n38093 = n9117 & n38092 ;
  assign n38094 = n35247 & n38093 ;
  assign n38095 = ~n23573 & n31780 ;
  assign n38098 = n22601 ^ n11175 ^ 1'b0 ;
  assign n38099 = ~n9792 & n38098 ;
  assign n38096 = ~n2429 & n22284 ;
  assign n38097 = n968 & n38096 ;
  assign n38100 = n38099 ^ n38097 ^ n9693 ;
  assign n38101 = ~n3334 & n11044 ;
  assign n38102 = n14259 & n17206 ;
  assign n38103 = n38102 ^ n12561 ^ 1'b0 ;
  assign n38104 = ( n13603 & n22345 ) | ( n13603 & ~n24117 ) | ( n22345 & ~n24117 ) ;
  assign n38105 = n8235 | n20643 ;
  assign n38106 = n25419 | n38105 ;
  assign n38107 = n4510 ^ n1976 ^ 1'b0 ;
  assign n38108 = n21242 & ~n38107 ;
  assign n38109 = ~n6591 & n38108 ;
  assign n38110 = n18930 ^ n4897 ^ 1'b0 ;
  assign n38111 = n6526 & ~n27880 ;
  assign n38112 = n38111 ^ n5390 ^ 1'b0 ;
  assign n38113 = ( n729 & n3880 ) | ( n729 & ~n10215 ) | ( n3880 & ~n10215 ) ;
  assign n38114 = n1539 | n38113 ;
  assign n38115 = n681 & n4990 ;
  assign n38116 = n8424 & ~n13840 ;
  assign n38117 = n38116 ^ n4870 ^ 1'b0 ;
  assign n38118 = ~n5034 & n5563 ;
  assign n38119 = n18137 | n38118 ;
  assign n38120 = n11168 ^ n1014 ^ 1'b0 ;
  assign n38121 = n13875 & ~n38120 ;
  assign n38122 = n8971 ^ n342 ^ 1'b0 ;
  assign n38123 = n38122 ^ n12682 ^ 1'b0 ;
  assign n38124 = n10302 ^ n6534 ^ 1'b0 ;
  assign n38125 = ~n17065 & n38124 ;
  assign n38126 = n5149 | n28015 ;
  assign n38127 = n6764 & n7031 ;
  assign n38128 = n38127 ^ n2197 ^ 1'b0 ;
  assign n38129 = ~n5507 & n38128 ;
  assign n38130 = n11956 & n38129 ;
  assign n38131 = n3974 ^ n1424 ^ 1'b0 ;
  assign n38132 = n38131 ^ n24284 ^ 1'b0 ;
  assign n38133 = n12346 | n38132 ;
  assign n38136 = n19416 & n28415 ;
  assign n38137 = n38136 ^ n3636 ^ 1'b0 ;
  assign n38134 = n1863 & ~n17491 ;
  assign n38135 = n38134 ^ n7873 ^ 1'b0 ;
  assign n38138 = n38137 ^ n38135 ^ n3406 ;
  assign n38139 = n9043 & ~n10232 ;
  assign n38140 = n38139 ^ n24170 ^ 1'b0 ;
  assign n38141 = n38138 & ~n38140 ;
  assign n38142 = n2973 | n7839 ;
  assign n38143 = n11007 | n14350 ;
  assign n38144 = n38143 ^ n17627 ^ 1'b0 ;
  assign n38145 = n8698 & ~n38144 ;
  assign n38146 = n38145 ^ n14262 ^ 1'b0 ;
  assign n38147 = n24448 & n31415 ;
  assign n38148 = ~n5499 & n32922 ;
  assign n38149 = n4335 | n6827 ;
  assign n38150 = n3446 & ~n38149 ;
  assign n38151 = ( n916 & n5244 ) | ( n916 & n8246 ) | ( n5244 & n8246 ) ;
  assign n38152 = ~n3489 & n38151 ;
  assign n38153 = n38152 ^ n28318 ^ 1'b0 ;
  assign n38154 = n38153 ^ n24895 ^ n21843 ;
  assign n38155 = n5664 & n29713 ;
  assign n38156 = n38155 ^ n35641 ^ n7282 ;
  assign n38157 = n9773 & ~n11486 ;
  assign n38158 = n38157 ^ n6813 ^ 1'b0 ;
  assign n38159 = n21418 ^ n11837 ^ 1'b0 ;
  assign n38160 = n16204 ^ n11359 ^ 1'b0 ;
  assign n38161 = n8070 & ~n38160 ;
  assign n38162 = n8508 & n28181 ;
  assign n38163 = ~n38161 & n38162 ;
  assign n38164 = n30697 ^ n339 ^ 1'b0 ;
  assign n38165 = n19369 ^ n11949 ^ 1'b0 ;
  assign n38166 = n37292 & ~n38165 ;
  assign n38168 = n8456 | n14560 ;
  assign n38167 = n13343 | n26010 ;
  assign n38169 = n38168 ^ n38167 ^ 1'b0 ;
  assign n38170 = ~n269 & n1690 ;
  assign n38171 = ~n38169 & n38170 ;
  assign n38172 = n20724 & ~n26473 ;
  assign n38173 = n4914 & n5689 ;
  assign n38174 = ~n5689 & n38173 ;
  assign n38175 = n26627 | n38174 ;
  assign n38176 = ~n38172 & n38175 ;
  assign n38177 = n38172 & n38176 ;
  assign n38180 = ~n1598 & n9840 ;
  assign n38181 = n38180 ^ n1812 ^ 1'b0 ;
  assign n38182 = n15775 & n38181 ;
  assign n38178 = n17275 | n30289 ;
  assign n38179 = n15319 | n38178 ;
  assign n38183 = n38182 ^ n38179 ^ 1'b0 ;
  assign n38184 = n1355 & n9373 ;
  assign n38185 = n38120 & n38184 ;
  assign n38186 = n33503 & n38185 ;
  assign n38187 = n7700 ^ n7520 ^ 1'b0 ;
  assign n38188 = n34098 | n38187 ;
  assign n38189 = n38188 ^ n26383 ^ 1'b0 ;
  assign n38190 = n23919 ^ n17503 ^ 1'b0 ;
  assign n38191 = n20367 | n38190 ;
  assign n38192 = n38191 ^ n12057 ^ 1'b0 ;
  assign n38193 = n31897 ^ n21881 ^ n19808 ;
  assign n38194 = ~n1701 & n38193 ;
  assign n38195 = n16410 & n38194 ;
  assign n38196 = n22743 & n38195 ;
  assign n38197 = n4407 ^ n611 ^ 1'b0 ;
  assign n38198 = n38197 ^ n13925 ^ 1'b0 ;
  assign n38199 = ~n1688 & n38198 ;
  assign n38200 = n6176 & n26743 ;
  assign n38201 = n38200 ^ n18858 ^ 1'b0 ;
  assign n38202 = n17600 & n32977 ;
  assign n38203 = n7844 & n28113 ;
  assign n38204 = n14008 & n38203 ;
  assign n38205 = n3473 ^ n2376 ^ 1'b0 ;
  assign n38206 = n782 & n2738 ;
  assign n38207 = ~n782 & n38206 ;
  assign n38208 = n290 & n38207 ;
  assign n38209 = n38208 ^ n19924 ^ 1'b0 ;
  assign n38210 = n81 & ~n110 ;
  assign n38211 = n110 & n38210 ;
  assign n38212 = n1075 & n1132 ;
  assign n38213 = ~n1132 & n38212 ;
  assign n38214 = n29260 | n38213 ;
  assign n38215 = ~n38211 & n38214 ;
  assign n38216 = n38209 & n38215 ;
  assign n38217 = n12529 | n38216 ;
  assign n38218 = n38216 & ~n38217 ;
  assign n38219 = ( ~n1050 & n20467 ) | ( ~n1050 & n38218 ) | ( n20467 & n38218 ) ;
  assign n38220 = ~n38205 & n38219 ;
  assign n38221 = n2626 & n7408 ;
  assign n38222 = n38221 ^ n1814 ^ 1'b0 ;
  assign n38223 = n7891 & n38222 ;
  assign n38224 = n38223 ^ n24014 ^ 1'b0 ;
  assign n38225 = ~n2848 & n38224 ;
  assign n38226 = n38225 ^ n18483 ^ 1'b0 ;
  assign n38227 = n10327 ^ n188 ^ 1'b0 ;
  assign n38228 = n26563 ^ n22633 ^ 1'b0 ;
  assign n38229 = ~n33980 & n38228 ;
  assign n38230 = n2563 ^ n1050 ^ 1'b0 ;
  assign n38232 = ~n2310 & n6847 ;
  assign n38233 = n38232 ^ n8663 ^ 1'b0 ;
  assign n38231 = n17416 & ~n22679 ;
  assign n38234 = n38233 ^ n38231 ^ 1'b0 ;
  assign n38235 = ~n33739 & n38234 ;
  assign n38236 = n38235 ^ n37597 ^ 1'b0 ;
  assign n38237 = n38236 ^ n12856 ^ n11360 ;
  assign n38238 = ~n38230 & n38237 ;
  assign n38239 = n1615 & ~n18106 ;
  assign n38240 = ~n12496 & n35066 ;
  assign n38241 = ~n2662 & n38240 ;
  assign n38242 = n28110 ^ n7621 ^ 1'b0 ;
  assign n38243 = n28590 & ~n38242 ;
  assign n38244 = n33019 ^ n5982 ^ 1'b0 ;
  assign n38245 = n33989 ^ n5545 ^ n1530 ;
  assign n38246 = ( n1987 & n23760 ) | ( n1987 & n32498 ) | ( n23760 & n32498 ) ;
  assign n38247 = n29290 ^ n27668 ^ 1'b0 ;
  assign n38248 = n31217 ^ n2125 ^ 1'b0 ;
  assign n38249 = ~n2989 & n23621 ;
  assign n38250 = n38249 ^ n13863 ^ 1'b0 ;
  assign n38251 = n788 & ~n38250 ;
  assign n38252 = n33694 ^ n2154 ^ 1'b0 ;
  assign n38253 = ( n767 & n3531 ) | ( n767 & ~n14785 ) | ( n3531 & ~n14785 ) ;
  assign n38254 = ~n17 & n38253 ;
  assign n38255 = ( n13986 & n26692 ) | ( n13986 & n28796 ) | ( n26692 & n28796 ) ;
  assign n38256 = n4177 & ~n16720 ;
  assign n38257 = ~n1675 & n19449 ;
  assign n38258 = n12294 & ~n38257 ;
  assign n38259 = n5775 & n7300 ;
  assign n38260 = n38259 ^ n13852 ^ 1'b0 ;
  assign n38261 = n38260 ^ n86 ^ 1'b0 ;
  assign n38262 = n27972 | n38261 ;
  assign n38263 = n38262 ^ n5399 ^ 1'b0 ;
  assign n38267 = n18909 ^ n1574 ^ 1'b0 ;
  assign n38268 = ~n9687 & n38267 ;
  assign n38269 = n20168 & n38268 ;
  assign n38264 = n27152 ^ n6727 ^ 1'b0 ;
  assign n38265 = ~n1901 & n38264 ;
  assign n38266 = n3837 & n38265 ;
  assign n38270 = n38269 ^ n38266 ^ 1'b0 ;
  assign n38271 = n9048 ^ n4479 ^ 1'b0 ;
  assign n38275 = n15792 | n28947 ;
  assign n38272 = n3567 | n4098 ;
  assign n38273 = n1021 & ~n32710 ;
  assign n38274 = n38272 & n38273 ;
  assign n38276 = n38275 ^ n38274 ^ n2460 ;
  assign n38277 = n4824 | n38276 ;
  assign n38278 = n15086 & n22646 ;
  assign n38279 = n38278 ^ n4660 ^ 1'b0 ;
  assign n38280 = ~n5529 & n38279 ;
  assign n38281 = ( n2743 & ~n7620 ) | ( n2743 & n38280 ) | ( ~n7620 & n38280 ) ;
  assign n38282 = n1877 & ~n10459 ;
  assign n38286 = n24117 ^ n14650 ^ 1'b0 ;
  assign n38283 = n3212 | n11133 ;
  assign n38284 = n38283 ^ n12575 ^ 1'b0 ;
  assign n38285 = n38284 ^ n26843 ^ 1'b0 ;
  assign n38287 = n38286 ^ n38285 ^ n15944 ;
  assign n38288 = n7488 & n16684 ;
  assign n38289 = n38288 ^ n2317 ^ 1'b0 ;
  assign n38290 = n21714 | n33382 ;
  assign n38291 = n13007 & ~n22941 ;
  assign n38292 = ( ~n10055 & n16714 ) | ( ~n10055 & n33865 ) | ( n16714 & n33865 ) ;
  assign n38293 = n11717 & n32048 ;
  assign n38294 = ~n38292 & n38293 ;
  assign n38295 = n6093 & n38294 ;
  assign n38296 = n7802 ^ n3930 ^ 1'b0 ;
  assign n38297 = n13843 | n38296 ;
  assign n38298 = n38297 ^ n16795 ^ 1'b0 ;
  assign n38299 = n7623 | n23727 ;
  assign n38300 = n28547 ^ n27230 ^ n24832 ;
  assign n38301 = n38300 ^ n6542 ^ 1'b0 ;
  assign n38302 = n30637 ^ n8256 ^ 1'b0 ;
  assign n38303 = n6129 & ~n19456 ;
  assign n38304 = n19926 & n38303 ;
  assign n38305 = n15230 & ~n23146 ;
  assign n38306 = n38305 ^ n19586 ^ 1'b0 ;
  assign n38307 = n13079 & ~n24848 ;
  assign n38308 = n38307 ^ n6756 ^ 1'b0 ;
  assign n38309 = n21612 | n24380 ;
  assign n38310 = n10212 & ~n21588 ;
  assign n38311 = ~n15471 & n19365 ;
  assign n38312 = n7702 & ~n38311 ;
  assign n38313 = n38312 ^ n27366 ^ n1562 ;
  assign n38314 = n1580 & ~n2078 ;
  assign n38315 = n38314 ^ n4685 ^ 1'b0 ;
  assign n38316 = n38315 ^ n14494 ^ 1'b0 ;
  assign n38317 = n7744 & n8098 ;
  assign n38318 = n2349 | n37228 ;
  assign n38319 = n38318 ^ n21009 ^ 1'b0 ;
  assign n38320 = ~n1944 & n17839 ;
  assign n38321 = n1230 & n38320 ;
  assign n38322 = n38321 ^ n26068 ^ 1'b0 ;
  assign n38323 = n5818 | n24326 ;
  assign n38324 = ~n5439 & n5628 ;
  assign n38325 = n22504 & ~n38324 ;
  assign n38326 = n38325 ^ n17717 ^ 1'b0 ;
  assign n38327 = n864 ^ n290 ^ 1'b0 ;
  assign n38329 = n2151 & n2648 ;
  assign n38330 = n38329 ^ n8421 ^ 1'b0 ;
  assign n38328 = n13588 & n25601 ;
  assign n38331 = n38330 ^ n38328 ^ 1'b0 ;
  assign n38332 = ~n35136 & n38331 ;
  assign n38333 = n15781 ^ n10432 ^ 1'b0 ;
  assign n38334 = n10785 ^ n846 ^ 1'b0 ;
  assign n38336 = n10274 & n29635 ;
  assign n38335 = ~n4147 & n16971 ;
  assign n38337 = n38336 ^ n38335 ^ 1'b0 ;
  assign n38338 = n7030 | n10443 ;
  assign n38339 = n5046 | n38338 ;
  assign n38340 = n38339 ^ n6348 ^ 1'b0 ;
  assign n38341 = n18534 | n33571 ;
  assign n38342 = n38341 ^ n6982 ^ 1'b0 ;
  assign n38343 = n38342 ^ n1667 ^ 1'b0 ;
  assign n38344 = n19777 & ~n38343 ;
  assign n38345 = n1460 & n38344 ;
  assign n38346 = ( n15367 & n23081 ) | ( n15367 & n38345 ) | ( n23081 & n38345 ) ;
  assign n38347 = n36398 ^ n11194 ^ 1'b0 ;
  assign n38348 = n6362 & ~n36348 ;
  assign n38350 = n5883 ^ n2330 ^ 1'b0 ;
  assign n38351 = n18374 & n38350 ;
  assign n38352 = n38351 ^ n7951 ^ 1'b0 ;
  assign n38353 = n23792 | n38352 ;
  assign n38349 = n32787 ^ n19369 ^ 1'b0 ;
  assign n38354 = n38353 ^ n38349 ^ 1'b0 ;
  assign n38355 = n30 & ~n142 ;
  assign n38356 = n38355 ^ n74 ^ 1'b0 ;
  assign n38357 = n38356 ^ n13251 ^ 1'b0 ;
  assign n38358 = n5030 & n15996 ;
  assign n38359 = n927 | n2791 ;
  assign n38360 = n13422 | n38359 ;
  assign n38361 = n38358 & ~n38360 ;
  assign n38362 = ~n17437 & n38361 ;
  assign n38363 = n23746 & n38362 ;
  assign n38364 = n36198 & ~n36678 ;
  assign n38365 = n13342 | n34976 ;
  assign n38366 = n22492 & n38365 ;
  assign n38367 = n27477 ^ n5929 ^ 1'b0 ;
  assign n38368 = n22519 | n38367 ;
  assign n38369 = n35079 & ~n38368 ;
  assign n38370 = n31795 ^ n22010 ^ n6836 ;
  assign n38371 = ~n7324 & n9288 ;
  assign n38372 = n1229 | n38371 ;
  assign n38373 = ( n3726 & n24230 ) | ( n3726 & ~n38372 ) | ( n24230 & ~n38372 ) ;
  assign n38374 = ~n5662 & n14460 ;
  assign n38375 = n38374 ^ n2192 ^ 1'b0 ;
  assign n38376 = n3610 | n8860 ;
  assign n38380 = ( ~n6157 & n7685 ) | ( ~n6157 & n22042 ) | ( n7685 & n22042 ) ;
  assign n38378 = n7749 | n14680 ;
  assign n38377 = n563 & n12582 ;
  assign n38379 = n38378 ^ n38377 ^ 1'b0 ;
  assign n38381 = n38380 ^ n38379 ^ 1'b0 ;
  assign n38382 = n38376 & ~n38381 ;
  assign n38383 = n8679 | n14134 ;
  assign n38384 = n38383 ^ n18784 ^ 1'b0 ;
  assign n38385 = n13582 ^ n8951 ^ 1'b0 ;
  assign n38386 = n35371 & ~n38385 ;
  assign n38387 = n38384 & n38386 ;
  assign n38388 = ( n3766 & n25553 ) | ( n3766 & ~n38387 ) | ( n25553 & ~n38387 ) ;
  assign n38389 = n34277 ^ n27488 ^ n16871 ;
  assign n38390 = n6321 & ~n26000 ;
  assign n38391 = n2150 & n29756 ;
  assign n38392 = n38391 ^ n3572 ^ 1'b0 ;
  assign n38393 = ~n38390 & n38392 ;
  assign n38394 = ~n3721 & n19265 ;
  assign n38395 = ~n4448 & n38394 ;
  assign n38396 = n11605 & ~n38395 ;
  assign n38397 = n1038 & ~n4054 ;
  assign n38398 = ~n10825 & n12258 ;
  assign n38399 = n23093 | n38398 ;
  assign n38400 = n1771 & ~n38399 ;
  assign n38401 = n25569 & n32259 ;
  assign n38402 = ~n4487 & n9899 ;
  assign n38403 = n4538 & ~n17113 ;
  assign n38404 = ( n27509 & n31187 ) | ( n27509 & n38403 ) | ( n31187 & n38403 ) ;
  assign n38405 = n5600 & n19045 ;
  assign n38406 = n11409 & ~n37855 ;
  assign n38407 = n5192 | n18281 ;
  assign n38408 = ~n5093 & n38407 ;
  assign n38409 = ~n3486 & n38408 ;
  assign n38410 = n38409 ^ n6575 ^ 1'b0 ;
  assign n38411 = ( n214 & n522 ) | ( n214 & n1327 ) | ( n522 & n1327 ) ;
  assign n38412 = n38411 ^ n2131 ^ 1'b0 ;
  assign n38413 = n26893 & n35683 ;
  assign n38414 = n38413 ^ n14244 ^ 1'b0 ;
  assign n38415 = n12516 | n38414 ;
  assign n38416 = n8896 | n37236 ;
  assign n38417 = n17170 & ~n38416 ;
  assign n38418 = ~n18908 & n35017 ;
  assign n38419 = ~n6198 & n38418 ;
  assign n38420 = n30723 & n31028 ;
  assign n38421 = n30217 ^ n20962 ^ 1'b0 ;
  assign n38422 = ~n7369 & n38421 ;
  assign n38423 = n22094 ^ n17507 ^ n2954 ;
  assign n38424 = n3341 & ~n4948 ;
  assign n38425 = n38424 ^ n3330 ^ 1'b0 ;
  assign n38426 = n12326 | n17048 ;
  assign n38427 = n38426 ^ n23790 ^ 1'b0 ;
  assign n38428 = ~n13358 & n23100 ;
  assign n38429 = n7677 & n18813 ;
  assign n38430 = n38429 ^ n9322 ^ 1'b0 ;
  assign n38431 = n10205 & ~n38430 ;
  assign n38432 = n38431 ^ n6330 ^ 1'b0 ;
  assign n38433 = ( n511 & ~n2177 ) | ( n511 & n5809 ) | ( ~n2177 & n5809 ) ;
  assign n38434 = n17692 ^ n4357 ^ 1'b0 ;
  assign n38435 = n6175 & n38434 ;
  assign n38436 = n13896 & n38435 ;
  assign n38437 = n22547 & n35295 ;
  assign n38438 = ~n6804 & n38437 ;
  assign n38439 = n38436 & n38438 ;
  assign n38440 = n25693 ^ n798 ^ 1'b0 ;
  assign n38441 = n19274 ^ n1110 ^ 1'b0 ;
  assign n38442 = n4356 | n38441 ;
  assign n38443 = n25008 ^ n19937 ^ 1'b0 ;
  assign n38444 = n10705 ^ n8901 ^ 1'b0 ;
  assign n38445 = n38443 | n38444 ;
  assign n38446 = n38445 ^ n28348 ^ n12740 ;
  assign n38447 = n2841 ^ n270 ^ 1'b0 ;
  assign n38448 = ( n30924 & n38056 ) | ( n30924 & ~n38447 ) | ( n38056 & ~n38447 ) ;
  assign n38449 = n5352 | n9319 ;
  assign n38450 = n1550 | n38449 ;
  assign n38451 = n5872 & ~n18899 ;
  assign n38452 = n15068 & n38451 ;
  assign n38453 = n32790 ^ n27840 ^ 1'b0 ;
  assign n38454 = n38452 | n38453 ;
  assign n38459 = n6885 ^ n2732 ^ 1'b0 ;
  assign n38455 = n14536 & ~n33221 ;
  assign n38456 = n23361 ^ n3162 ^ 1'b0 ;
  assign n38457 = ~n35226 & n38456 ;
  assign n38458 = ~n38455 & n38457 ;
  assign n38460 = n38459 ^ n38458 ^ 1'b0 ;
  assign n38461 = n8799 ^ n4618 ^ 1'b0 ;
  assign n38462 = n6542 | n38461 ;
  assign n38463 = n24827 & ~n38462 ;
  assign n38464 = n38460 & n38463 ;
  assign n38465 = ( n13 & ~n880 ) | ( n13 & n14405 ) | ( ~n880 & n14405 ) ;
  assign n38466 = ~n6065 & n14604 ;
  assign n38467 = n38466 ^ n24188 ^ 1'b0 ;
  assign n38468 = ~n16523 & n38467 ;
  assign n38469 = n5881 ^ n2393 ^ 1'b0 ;
  assign n38470 = n17059 | n38469 ;
  assign n38471 = n6291 & ~n20860 ;
  assign n38472 = n23792 & n28218 ;
  assign n38473 = n625 & ~n10387 ;
  assign n38474 = n25307 & n38473 ;
  assign n38475 = n9698 ^ n7615 ^ 1'b0 ;
  assign n38476 = n8452 & n13794 ;
  assign n38477 = n22963 ^ n14137 ^ 1'b0 ;
  assign n38478 = n5946 & n37845 ;
  assign n38479 = n38478 ^ n15825 ^ 1'b0 ;
  assign n38481 = n919 & n5727 ;
  assign n38480 = ~n466 & n3547 ;
  assign n38482 = n38481 ^ n38480 ^ n7149 ;
  assign n38483 = n34103 ^ n22626 ^ 1'b0 ;
  assign n38484 = n38482 | n38483 ;
  assign n38485 = n3246 & n15438 ;
  assign n38486 = n13311 & ~n38485 ;
  assign n38487 = n38484 & n38486 ;
  assign n38489 = n6868 & ~n36082 ;
  assign n38490 = ~n12214 & n38489 ;
  assign n38488 = n14091 & n29107 ;
  assign n38491 = n38490 ^ n38488 ^ 1'b0 ;
  assign n38492 = n38491 ^ n5188 ^ 1'b0 ;
  assign n38493 = n14149 & n38492 ;
  assign n38494 = ~n14295 & n38493 ;
  assign n38495 = n22927 & n37182 ;
  assign n38496 = n17135 & n17583 ;
  assign n38497 = n9076 & n38496 ;
  assign n38498 = n11552 & n38497 ;
  assign n38499 = n14497 & n38498 ;
  assign n38500 = n34961 ^ n845 ^ 1'b0 ;
  assign n38501 = n25468 | n38500 ;
  assign n38502 = n38501 ^ n15667 ^ 1'b0 ;
  assign n38503 = n6472 | n10248 ;
  assign n38504 = n38503 ^ n4712 ^ 1'b0 ;
  assign n38505 = n4380 & ~n18067 ;
  assign n38506 = n120 & ~n15351 ;
  assign n38507 = n17629 & ~n38506 ;
  assign n38508 = n38505 & ~n38507 ;
  assign n38509 = n15076 ^ n889 ^ 1'b0 ;
  assign n38510 = n3634 & ~n4143 ;
  assign n38511 = n38510 ^ n10388 ^ 1'b0 ;
  assign n38512 = n13052 | n38511 ;
  assign n38513 = ~n34899 & n38512 ;
  assign n38514 = n38513 ^ n1554 ^ 1'b0 ;
  assign n38515 = n14920 ^ n4997 ^ 1'b0 ;
  assign n38516 = ~n791 & n38515 ;
  assign n38517 = n38516 ^ n34909 ^ 1'b0 ;
  assign n38518 = n2829 & ~n11140 ;
  assign n38519 = ~n19759 & n38518 ;
  assign n38520 = n22884 | n32403 ;
  assign n38521 = n3990 & ~n38520 ;
  assign n38522 = n38521 ^ n34560 ^ n2820 ;
  assign n38523 = n20500 ^ n6149 ^ 1'b0 ;
  assign n38524 = n30748 & ~n33869 ;
  assign n38525 = n5776 & ~n34145 ;
  assign n38526 = n6127 ^ n4914 ^ 1'b0 ;
  assign n38527 = n16642 ^ n1907 ^ 1'b0 ;
  assign n38528 = n38526 | n38527 ;
  assign n38529 = n6406 | n38528 ;
  assign n38530 = n6456 & n38529 ;
  assign n38531 = n762 | n15182 ;
  assign n38532 = n18072 ^ n2864 ^ 1'b0 ;
  assign n38533 = ~n5097 & n38532 ;
  assign n38534 = n38531 & ~n38533 ;
  assign n38535 = n25657 ^ n7898 ^ 1'b0 ;
  assign n38536 = n453 & ~n16236 ;
  assign n38537 = ~n38535 & n38536 ;
  assign n38538 = n16319 ^ n5760 ^ 1'b0 ;
  assign n38539 = n10238 & ~n18046 ;
  assign n38540 = n12361 ^ n7589 ^ 1'b0 ;
  assign n38541 = n4529 | n7626 ;
  assign n38542 = n7626 & ~n38541 ;
  assign n38543 = n3732 & ~n38542 ;
  assign n38544 = n38543 ^ n3395 ^ 1'b0 ;
  assign n38546 = n18239 ^ n10322 ^ 1'b0 ;
  assign n38545 = n798 | n5352 ;
  assign n38547 = n38546 ^ n38545 ^ n20533 ;
  assign n38548 = ( ~n16854 & n38544 ) | ( ~n16854 & n38547 ) | ( n38544 & n38547 ) ;
  assign n38549 = n829 & ~n1717 ;
  assign n38550 = ~n27998 & n38549 ;
  assign n38551 = n18844 & ~n38550 ;
  assign n38552 = ~n9748 & n15579 ;
  assign n38553 = n38552 ^ n18494 ^ 1'b0 ;
  assign n38554 = n38553 ^ n34940 ^ n4570 ;
  assign n38555 = n2028 ^ n1065 ^ 1'b0 ;
  assign n38556 = n1510 | n38555 ;
  assign n38557 = n38556 ^ n17320 ^ 1'b0 ;
  assign n38558 = n1853 & n30231 ;
  assign n38559 = n38557 & n38558 ;
  assign n38560 = n26217 & ~n34059 ;
  assign n38561 = n12224 ^ n5802 ^ 1'b0 ;
  assign n38562 = n34277 ^ n10749 ^ n640 ;
  assign n38564 = n8518 & n12073 ;
  assign n38565 = n17611 & n38564 ;
  assign n38563 = n214 & n1705 ;
  assign n38566 = n38565 ^ n38563 ^ 1'b0 ;
  assign n38567 = n4863 & n10222 ;
  assign n38572 = n17131 ^ n11316 ^ 1'b0 ;
  assign n38568 = ~n8073 & n16832 ;
  assign n38569 = n19577 | n28870 ;
  assign n38570 = n8204 | n38569 ;
  assign n38571 = n38568 & n38570 ;
  assign n38573 = n38572 ^ n38571 ^ 1'b0 ;
  assign n38574 = n30141 ^ n1703 ^ 1'b0 ;
  assign n38576 = n15796 & ~n27092 ;
  assign n38577 = n29379 & ~n38576 ;
  assign n38578 = n71 & n38577 ;
  assign n38579 = n38578 ^ n24669 ^ 1'b0 ;
  assign n38575 = ( n3665 & ~n18351 ) | ( n3665 & n24389 ) | ( ~n18351 & n24389 ) ;
  assign n38580 = n38579 ^ n38575 ^ n11458 ;
  assign n38581 = n6037 & n6089 ;
  assign n38582 = n13988 ^ n1829 ^ 1'b0 ;
  assign n38583 = n38581 | n38582 ;
  assign n38584 = ~n17976 & n30155 ;
  assign n38585 = n3280 | n7007 ;
  assign n38586 = n38585 ^ n9385 ^ 1'b0 ;
  assign n38587 = n38586 ^ n36357 ^ 1'b0 ;
  assign n38588 = n5528 & ~n38587 ;
  assign n38589 = n4171 | n23043 ;
  assign n38590 = n38589 ^ n35369 ^ 1'b0 ;
  assign n38591 = n32454 ^ n21963 ^ n4221 ;
  assign n38592 = n606 & n13212 ;
  assign n38593 = ( n38590 & ~n38591 ) | ( n38590 & n38592 ) | ( ~n38591 & n38592 ) ;
  assign n38594 = n28454 & ~n32855 ;
  assign n38595 = n38594 ^ n8376 ^ n4776 ;
  assign n38596 = n8357 & n24439 ;
  assign n38597 = n4135 & ~n5213 ;
  assign n38598 = n6472 | n8087 ;
  assign n38599 = n38598 ^ n2565 ^ 1'b0 ;
  assign n38600 = n2519 & n38599 ;
  assign n38601 = n38600 ^ n38151 ^ 1'b0 ;
  assign n38602 = n20475 & ~n21466 ;
  assign n38603 = n1023 & ~n38602 ;
  assign n38604 = n37957 ^ n9560 ^ 1'b0 ;
  assign n38605 = n38604 ^ n6461 ^ n1816 ;
  assign n38606 = n25668 ^ n17329 ^ 1'b0 ;
  assign n38607 = n22646 & n31353 ;
  assign n38608 = n38606 & n38607 ;
  assign n38609 = n14203 ^ n13673 ^ 1'b0 ;
  assign n38610 = ~n26156 & n26913 ;
  assign n38611 = n777 | n6765 ;
  assign n38612 = n14285 | n38611 ;
  assign n38613 = n2958 | n8598 ;
  assign n38614 = n38613 ^ n34801 ^ 1'b0 ;
  assign n38615 = ~n38613 & n38614 ;
  assign n38616 = n651 & ~n798 ;
  assign n38617 = n3979 & n38616 ;
  assign n38618 = n30935 | n34709 ;
  assign n38619 = n38617 & ~n38618 ;
  assign n38620 = n38619 ^ n22373 ^ 1'b0 ;
  assign n38621 = n4366 & n8995 ;
  assign n38622 = n4619 & n27968 ;
  assign n38623 = n38622 ^ n8023 ^ 1'b0 ;
  assign n38625 = n25615 ^ n957 ^ 1'b0 ;
  assign n38626 = n38625 ^ n21612 ^ n6157 ;
  assign n38624 = n5168 & ~n32400 ;
  assign n38627 = n38626 ^ n38624 ^ 1'b0 ;
  assign n38628 = n38627 ^ n33241 ^ 1'b0 ;
  assign n38629 = n15677 & n38628 ;
  assign n38630 = n24252 ^ n22068 ^ 1'b0 ;
  assign n38631 = ~n3923 & n25581 ;
  assign n38632 = ( ~n8799 & n28784 ) | ( ~n8799 & n30518 ) | ( n28784 & n30518 ) ;
  assign n38633 = n1918 & ~n16607 ;
  assign n38634 = n38633 ^ n4639 ^ 1'b0 ;
  assign n38635 = n17584 ^ n1826 ^ 1'b0 ;
  assign n38636 = n20846 ^ n4275 ^ 1'b0 ;
  assign n38637 = n12573 & ~n38636 ;
  assign n38638 = n24601 | n38637 ;
  assign n38639 = n19575 ^ n16327 ^ 1'b0 ;
  assign n38640 = ~n8566 & n38639 ;
  assign n38641 = n38640 ^ n24541 ^ 1'b0 ;
  assign n38642 = n10775 | n18573 ;
  assign n38643 = n18310 ^ n4856 ^ 1'b0 ;
  assign n38644 = n37462 & n38643 ;
  assign n38645 = n20 & n38644 ;
  assign n38646 = n11474 & n38645 ;
  assign n38647 = n38646 ^ n7382 ^ 1'b0 ;
  assign n38648 = n253 & ~n22131 ;
  assign n38649 = ~n1347 & n38648 ;
  assign n38650 = n38649 ^ x7 ^ 1'b0 ;
  assign n38651 = n13632 | n38650 ;
  assign n38652 = n35567 ^ n17293 ^ 1'b0 ;
  assign n38653 = n13922 | n38652 ;
  assign n38654 = ~n20785 & n23908 ;
  assign n38655 = n1235 | n21685 ;
  assign n38656 = n13884 | n38655 ;
  assign n38657 = ( n8223 & ~n17924 ) | ( n8223 & n37269 ) | ( ~n17924 & n37269 ) ;
  assign n38658 = n7766 ^ n7219 ^ 1'b0 ;
  assign n38659 = n7696 & ~n9304 ;
  assign n38660 = n21644 ^ n4399 ^ 1'b0 ;
  assign n38661 = n38659 & ~n38660 ;
  assign n38662 = n38661 ^ n3178 ^ 1'b0 ;
  assign n38663 = n16257 & ~n25006 ;
  assign n38664 = n38662 & n38663 ;
  assign n38665 = n1306 & ~n3783 ;
  assign n38667 = ~n1205 & n13541 ;
  assign n38666 = n3696 | n18921 ;
  assign n38668 = n38667 ^ n38666 ^ 1'b0 ;
  assign n38669 = n38668 ^ n13225 ^ 1'b0 ;
  assign n38670 = n8254 | n23879 ;
  assign n38671 = n38669 | n38670 ;
  assign n38672 = ~n774 & n17999 ;
  assign n38673 = n10935 | n24252 ;
  assign n38674 = n9218 & n20657 ;
  assign n38675 = n38674 ^ n1701 ^ 1'b0 ;
  assign n38676 = n15915 & ~n20621 ;
  assign n38677 = n36503 ^ n32097 ^ 1'b0 ;
  assign n38678 = n15086 & n38677 ;
  assign n38679 = n26701 ^ n20291 ^ 1'b0 ;
  assign n38680 = ( n20313 & n38678 ) | ( n20313 & ~n38679 ) | ( n38678 & ~n38679 ) ;
  assign n38681 = n21947 ^ n17011 ^ n1256 ;
  assign n38682 = n23013 & ~n35754 ;
  assign n38683 = n38682 ^ n14269 ^ 1'b0 ;
  assign n38686 = n4976 ^ n3949 ^ 1'b0 ;
  assign n38684 = n23633 ^ n6576 ^ 1'b0 ;
  assign n38685 = n31240 | n38684 ;
  assign n38687 = n38686 ^ n38685 ^ 1'b0 ;
  assign n38688 = n8310 & ~n38687 ;
  assign n38689 = n8750 | n23230 ;
  assign n38690 = n11812 | n38689 ;
  assign n38691 = n24897 ^ n5152 ^ 1'b0 ;
  assign n38692 = n1170 | n13311 ;
  assign n38693 = n38692 ^ n35260 ^ 1'b0 ;
  assign n38694 = ~n4468 & n38693 ;
  assign n38696 = n4037 & ~n11577 ;
  assign n38697 = ~n354 & n38696 ;
  assign n38695 = n2426 & ~n6833 ;
  assign n38698 = n38697 ^ n38695 ^ 1'b0 ;
  assign n38699 = n513 & n7185 ;
  assign n38700 = n38699 ^ n1636 ^ 1'b0 ;
  assign n38701 = n38700 ^ n17594 ^ 1'b0 ;
  assign n38702 = ~n4367 & n5872 ;
  assign n38703 = ~n38701 & n38702 ;
  assign n38704 = n4381 & n38703 ;
  assign n38705 = n38704 ^ n12769 ^ 1'b0 ;
  assign n38706 = n3193 & n38705 ;
  assign n38707 = n4201 & ~n11119 ;
  assign n38708 = n38707 ^ n29020 ^ 1'b0 ;
  assign n38709 = n25231 ^ n15892 ^ 1'b0 ;
  assign n38710 = n1363 & ~n38709 ;
  assign n38711 = n17778 ^ n16135 ^ 1'b0 ;
  assign n38712 = n12038 | n38711 ;
  assign n38713 = n27489 | n38712 ;
  assign n38714 = n3110 & ~n38713 ;
  assign n38715 = n14368 ^ n2406 ^ 1'b0 ;
  assign n38716 = n3349 & ~n11605 ;
  assign n38717 = ~n3764 & n38716 ;
  assign n38718 = n11703 & ~n24162 ;
  assign n38719 = n38718 ^ n12165 ^ 1'b0 ;
  assign n38720 = n23715 & ~n38719 ;
  assign n38721 = ~n6116 & n6291 ;
  assign n38722 = n38721 ^ n9022 ^ 1'b0 ;
  assign n38723 = n12867 | n38722 ;
  assign n38724 = n38723 ^ n38286 ^ 1'b0 ;
  assign n38725 = n9511 & ~n20928 ;
  assign n38732 = n15856 | n16613 ;
  assign n38733 = n38732 ^ n14530 ^ 1'b0 ;
  assign n38726 = n24791 ^ n8072 ^ 1'b0 ;
  assign n38727 = n7400 & n17114 ;
  assign n38728 = n38726 & n38727 ;
  assign n38729 = n38728 ^ n18100 ^ 1'b0 ;
  assign n38730 = ~n4547 & n38729 ;
  assign n38731 = ~n35904 & n38730 ;
  assign n38734 = n38733 ^ n38731 ^ 1'b0 ;
  assign n38735 = ~n4438 & n13444 ;
  assign n38736 = n2993 & n38735 ;
  assign n38737 = n17404 | n38736 ;
  assign n38738 = n465 & ~n38737 ;
  assign n38739 = ~n13693 & n24304 ;
  assign n38740 = n3488 & n18662 ;
  assign n38741 = n21229 & ~n38740 ;
  assign n38742 = n38741 ^ n38724 ^ 1'b0 ;
  assign n38743 = ~n38739 & n38742 ;
  assign n38744 = n18900 & n19846 ;
  assign n38745 = n10391 | n38744 ;
  assign n38748 = ( n4423 & n5562 ) | ( n4423 & ~n30059 ) | ( n5562 & ~n30059 ) ;
  assign n38749 = n38748 ^ n519 ^ 1'b0 ;
  assign n38746 = n5584 | n17802 ;
  assign n38747 = n3896 & n38746 ;
  assign n38750 = n38749 ^ n38747 ^ 1'b0 ;
  assign n38751 = n20521 ^ n3088 ^ 1'b0 ;
  assign n38752 = n11005 | n38751 ;
  assign n38753 = n19150 ^ n4593 ^ 1'b0 ;
  assign n38754 = x6 & n12836 ;
  assign n38755 = n36049 & n38754 ;
  assign n38756 = n11907 & ~n38755 ;
  assign n38757 = ~n15446 & n21061 ;
  assign n38758 = n2391 & ~n38757 ;
  assign n38760 = n18104 ^ n3766 ^ 1'b0 ;
  assign n38759 = n10764 & n24905 ;
  assign n38761 = n38760 ^ n38759 ^ 1'b0 ;
  assign n38762 = n6664 & n13354 ;
  assign n38763 = n15714 & n38762 ;
  assign n38764 = n38020 | n38763 ;
  assign n38765 = n38764 ^ n19409 ^ 1'b0 ;
  assign n38766 = n158 | n8246 ;
  assign n38767 = n38766 ^ n13600 ^ n2508 ;
  assign n38768 = n22341 ^ n16823 ^ 1'b0 ;
  assign n38769 = n23403 | n38768 ;
  assign n38770 = n38769 ^ n25296 ^ 1'b0 ;
  assign n38771 = n5898 | n9823 ;
  assign n38772 = n19305 & ~n38771 ;
  assign n38773 = n1944 | n28837 ;
  assign n38774 = n38772 & ~n38773 ;
  assign n38775 = ~n12158 & n21473 ;
  assign n38776 = n38775 ^ n17407 ^ 1'b0 ;
  assign n38777 = n38776 ^ n22743 ^ 1'b0 ;
  assign n38778 = n1383 & n38777 ;
  assign n38779 = n340 & n32574 ;
  assign n38780 = n19657 & n38779 ;
  assign n38781 = n12594 ^ n5130 ^ 1'b0 ;
  assign n38782 = n22286 & ~n38781 ;
  assign n38783 = n31657 & n38782 ;
  assign n38784 = n3632 & ~n13328 ;
  assign n38785 = n12361 ^ n4461 ^ 1'b0 ;
  assign n38786 = n21836 ^ n10154 ^ 1'b0 ;
  assign n38787 = ~n23020 & n38786 ;
  assign n38788 = ( n508 & n2881 ) | ( n508 & n13685 ) | ( n2881 & n13685 ) ;
  assign n38789 = n38788 ^ n19206 ^ 1'b0 ;
  assign n38790 = ~n38787 & n38789 ;
  assign n38791 = n38790 ^ n5444 ^ n1759 ;
  assign n38792 = ~n38785 & n38791 ;
  assign n38793 = n37413 & ~n38792 ;
  assign n38794 = n13601 | n36851 ;
  assign n38795 = n38794 ^ n25717 ^ 1'b0 ;
  assign n38796 = n5067 & ~n23405 ;
  assign n38797 = n27031 ^ n20203 ^ 1'b0 ;
  assign n38798 = n33019 & ~n38797 ;
  assign n38799 = n38798 ^ n26803 ^ 1'b0 ;
  assign n38800 = n30814 ^ n26312 ^ 1'b0 ;
  assign n38801 = n23065 | n37712 ;
  assign n38802 = n1174 & ~n7862 ;
  assign n38803 = n21547 & n38802 ;
  assign n38804 = n38803 ^ n8233 ^ 1'b0 ;
  assign n38805 = n15153 & ~n38804 ;
  assign n38806 = n5138 ^ n4191 ^ 1'b0 ;
  assign n38807 = n38805 & ~n38806 ;
  assign n38808 = n5618 | n7369 ;
  assign n38809 = n38808 ^ n810 ^ 1'b0 ;
  assign n38810 = n20693 & n38809 ;
  assign n38811 = n12598 & n38810 ;
  assign n38814 = n8840 & ~n19336 ;
  assign n38815 = ~n14054 & n38814 ;
  assign n38812 = ~n2127 & n6029 ;
  assign n38813 = ~n4091 & n38812 ;
  assign n38816 = n38815 ^ n38813 ^ 1'b0 ;
  assign n38817 = n286 & ~n988 ;
  assign n38818 = ~n286 & n38817 ;
  assign n38819 = ~n1611 & n38818 ;
  assign n38820 = ~n38818 & n38819 ;
  assign n38821 = n2227 & n21753 ;
  assign n38822 = n38821 ^ n7108 ^ 1'b0 ;
  assign n38823 = ~n38820 & n38822 ;
  assign n38824 = n38823 ^ n22059 ^ n5518 ;
  assign n38825 = n37065 ^ n8975 ^ 1'b0 ;
  assign n38826 = n38824 | n38825 ;
  assign n38827 = n1031 | n28254 ;
  assign n38828 = n10002 | n38827 ;
  assign n38829 = n10452 ^ n710 ^ 1'b0 ;
  assign n38830 = n14057 & ~n38829 ;
  assign n38831 = n3954 & ~n9719 ;
  assign n38832 = ~n8016 & n38831 ;
  assign n38833 = ( ~n32425 & n38830 ) | ( ~n32425 & n38832 ) | ( n38830 & n38832 ) ;
  assign n38834 = n24219 & ~n30120 ;
  assign n38835 = ~n10728 & n38834 ;
  assign n38836 = n9179 & n15262 ;
  assign n38837 = ~n14112 & n14838 ;
  assign n38838 = ~n6762 & n33783 ;
  assign n38839 = n29595 ^ n10372 ^ 1'b0 ;
  assign n38840 = n38839 ^ n30960 ^ n5115 ;
  assign n38841 = n20499 ^ n15436 ^ 1'b0 ;
  assign n38847 = n996 | n13037 ;
  assign n38848 = n996 & ~n38847 ;
  assign n38842 = n446 & ~n6923 ;
  assign n38843 = ~n446 & n38842 ;
  assign n38844 = ~n12135 & n36312 ;
  assign n38845 = n12135 & n38844 ;
  assign n38846 = n38843 | n38845 ;
  assign n38849 = n38848 ^ n38846 ^ 1'b0 ;
  assign n38850 = ~n8312 & n20257 ;
  assign n38851 = n25349 ^ n7093 ^ 1'b0 ;
  assign n38852 = n21399 | n38851 ;
  assign n38853 = n18455 & ~n38852 ;
  assign n38854 = n25404 ^ n1554 ^ 1'b0 ;
  assign n38855 = n7319 ^ n6760 ^ n2940 ;
  assign n38856 = n8010 & n8840 ;
  assign n38857 = n35825 & n38856 ;
  assign n38858 = n35595 & n36577 ;
  assign n38859 = n304 & n38858 ;
  assign n38860 = n1254 & ~n13706 ;
  assign n38861 = n31166 & n38860 ;
  assign n38862 = n17284 ^ n8823 ^ 1'b0 ;
  assign n38863 = n874 | n38862 ;
  assign n38864 = n86 & ~n38863 ;
  assign n38865 = n38864 ^ n14454 ^ 1'b0 ;
  assign n38866 = n10657 ^ n7243 ^ n1369 ;
  assign n38867 = ~n25010 & n38866 ;
  assign n38868 = ~n19271 & n38867 ;
  assign n38869 = ~n466 & n23214 ;
  assign n38870 = n169 & n38869 ;
  assign n38871 = n32176 | n38870 ;
  assign n38872 = n38871 ^ n19821 ^ 1'b0 ;
  assign n38873 = n38872 ^ n19240 ^ n5323 ;
  assign n38874 = n14560 & n31718 ;
  assign n38875 = n28267 | n38874 ;
  assign n38876 = n38875 ^ n24669 ^ 1'b0 ;
  assign n38877 = n6257 & n11274 ;
  assign n38878 = n38877 ^ n4224 ^ 1'b0 ;
  assign n38879 = ( n438 & n20080 ) | ( n438 & ~n38878 ) | ( n20080 & ~n38878 ) ;
  assign n38880 = n7952 ^ n5242 ^ n2845 ;
  assign n38881 = ~n37778 & n38880 ;
  assign n38882 = n38879 & ~n38881 ;
  assign n38883 = n16161 | n18010 ;
  assign n38884 = n34997 ^ n15750 ^ 1'b0 ;
  assign n38885 = n2649 ^ n470 ^ 1'b0 ;
  assign n38886 = n1918 & ~n38885 ;
  assign n38887 = n5076 & n38886 ;
  assign n38888 = n19680 & n38887 ;
  assign n38889 = ~n1853 & n38888 ;
  assign n38890 = n2815 & n9934 ;
  assign n38892 = n158 | n23221 ;
  assign n38891 = n11474 | n14863 ;
  assign n38893 = n38892 ^ n38891 ^ 1'b0 ;
  assign n38894 = n30508 ^ n15763 ^ 1'b0 ;
  assign n38895 = n27606 ^ n4085 ^ n586 ;
  assign n38896 = n3475 & n19368 ;
  assign n38897 = n25584 & n31117 ;
  assign n38898 = n32811 ^ n13068 ^ 1'b0 ;
  assign n38899 = ~n19153 & n38898 ;
  assign n38900 = n2478 ^ n1260 ^ 1'b0 ;
  assign n38901 = n2711 ^ n1870 ^ 1'b0 ;
  assign n38902 = n38900 & n38901 ;
  assign n38903 = ( n26906 & n38899 ) | ( n26906 & n38902 ) | ( n38899 & n38902 ) ;
  assign n38904 = n823 & ~n4400 ;
  assign n38905 = ~n8248 & n11635 ;
  assign n38906 = n38905 ^ n2448 ^ 1'b0 ;
  assign n38907 = ~n2213 & n6698 ;
  assign n38908 = n38907 ^ n417 ^ 1'b0 ;
  assign n38909 = ~n23875 & n38908 ;
  assign n38910 = n38906 & n38909 ;
  assign n38911 = ~n20946 & n38155 ;
  assign n38912 = ~n2859 & n13015 ;
  assign n38913 = n21867 ^ n18486 ^ n5866 ;
  assign n38914 = ~n3101 & n8885 ;
  assign n38915 = n5419 & n38914 ;
  assign n38916 = n38915 ^ n16050 ^ 1'b0 ;
  assign n38917 = n33993 ^ n3774 ^ 1'b0 ;
  assign n38918 = ~n38916 & n38917 ;
  assign n38919 = n38918 ^ n28381 ^ 1'b0 ;
  assign n38920 = ~n2379 & n11471 ;
  assign n38921 = n23269 | n38920 ;
  assign n38922 = ~n25508 & n27321 ;
  assign n38923 = n277 & n38922 ;
  assign n38924 = n5396 & n8729 ;
  assign n38925 = n38924 ^ n6923 ^ 1'b0 ;
  assign n38928 = n21008 & ~n28771 ;
  assign n38926 = ~n18744 & n28359 ;
  assign n38927 = n6866 & ~n38926 ;
  assign n38929 = n38928 ^ n38927 ^ 1'b0 ;
  assign n38930 = ~n1819 & n19436 ;
  assign n38931 = n38930 ^ n5885 ^ 1'b0 ;
  assign n38932 = n22338 & ~n37408 ;
  assign n38933 = n17935 ^ n4993 ^ 1'b0 ;
  assign n38935 = n835 & ~n22248 ;
  assign n38934 = n2443 & ~n16463 ;
  assign n38936 = n38935 ^ n38934 ^ 1'b0 ;
  assign n38937 = n7153 | n29149 ;
  assign n38938 = n38937 ^ n11061 ^ 1'b0 ;
  assign n38939 = n30834 & ~n31488 ;
  assign n38940 = ~n439 & n38939 ;
  assign n38941 = ~n16897 & n22338 ;
  assign n38942 = n26941 ^ n2164 ^ 1'b0 ;
  assign n38943 = n4576 & ~n38942 ;
  assign n38944 = ~n29399 & n38943 ;
  assign n38945 = n18274 ^ n14156 ^ 1'b0 ;
  assign n38946 = n14126 ^ n12659 ^ n2324 ;
  assign n38947 = n38945 & ~n38946 ;
  assign n38948 = n22651 ^ n17737 ^ 1'b0 ;
  assign n38949 = n20732 ^ n6764 ^ 1'b0 ;
  assign n38950 = n15923 | n38949 ;
  assign n38951 = ~n9667 & n32522 ;
  assign n38952 = n34567 & n38951 ;
  assign n38953 = n5470 & n28771 ;
  assign n38954 = n38566 ^ n10094 ^ 1'b0 ;
  assign n38955 = n35467 & n38954 ;
  assign n38956 = n5628 & ~n13555 ;
  assign n38957 = n2811 & n38956 ;
  assign n38958 = n38957 ^ n31767 ^ 1'b0 ;
  assign n38959 = ( n1763 & n16559 ) | ( n1763 & ~n36561 ) | ( n16559 & ~n36561 ) ;
  assign n38960 = n15200 & ~n38023 ;
  assign n38961 = n2917 | n12754 ;
  assign n38962 = n14301 ^ n7665 ^ 1'b0 ;
  assign n38963 = n19636 ^ n18031 ^ 1'b0 ;
  assign n38964 = n7089 ^ n2824 ^ 1'b0 ;
  assign n38965 = ~n10337 & n38964 ;
  assign n38966 = ( n1434 & n15690 ) | ( n1434 & n38965 ) | ( n15690 & n38965 ) ;
  assign n38967 = n22173 ^ n12990 ^ n6156 ;
  assign n38968 = n28540 & n38967 ;
  assign n38969 = n38968 ^ n3211 ^ 1'b0 ;
  assign n38970 = n24074 ^ n21849 ^ 1'b0 ;
  assign n38971 = n38969 & n38970 ;
  assign n38972 = n2256 & n7277 ;
  assign n38973 = n38972 ^ n4738 ^ 1'b0 ;
  assign n38974 = n8944 & ~n38973 ;
  assign n38975 = n38974 ^ n27312 ^ 1'b0 ;
  assign n38976 = n18049 & ~n30084 ;
  assign n38977 = n38976 ^ n37754 ^ 1'b0 ;
  assign n38978 = n10092 | n10909 ;
  assign n38979 = n4367 | n38978 ;
  assign n38980 = n12902 ^ n11572 ^ 1'b0 ;
  assign n38981 = ~n15624 & n38980 ;
  assign n38982 = n18732 & n23654 ;
  assign n38983 = ~n38981 & n38982 ;
  assign n38984 = ~n167 & n10342 ;
  assign n38985 = ~n4381 & n11803 ;
  assign n38986 = n2837 | n38985 ;
  assign n38987 = n6035 & n11624 ;
  assign n38988 = n38987 ^ n6240 ^ 1'b0 ;
  assign n38989 = n10303 & n12060 ;
  assign n38990 = ~n3626 & n38989 ;
  assign n38991 = ( n10529 & n11402 ) | ( n10529 & ~n14960 ) | ( n11402 & ~n14960 ) ;
  assign n38992 = n6398 & n38991 ;
  assign n38993 = n1434 | n31594 ;
  assign n38994 = n21765 & n23133 ;
  assign n38995 = n4942 | n13346 ;
  assign n38996 = ~n2051 & n3995 ;
  assign n38997 = ~n21834 & n35101 ;
  assign n38998 = ~n6834 & n33661 ;
  assign n38999 = n15117 & n38998 ;
  assign n39000 = n9224 & ~n23309 ;
  assign n39001 = n39000 ^ n1786 ^ 1'b0 ;
  assign n39002 = n39001 ^ n8878 ^ 1'b0 ;
  assign n39003 = n3393 & ~n39002 ;
  assign n39004 = n2954 | n6392 ;
  assign n39005 = n13194 & n39004 ;
  assign n39006 = n17689 ^ n5493 ^ 1'b0 ;
  assign n39007 = n5861 | n39006 ;
  assign n39008 = ~n11942 & n39007 ;
  assign n39009 = n6347 ^ n2837 ^ 1'b0 ;
  assign n39010 = ~n39008 & n39009 ;
  assign n39011 = ~n11535 & n11869 ;
  assign n39012 = n39010 | n39011 ;
  assign n39013 = n790 | n1732 ;
  assign n39014 = ( n3210 & n8570 ) | ( n3210 & ~n18232 ) | ( n8570 & ~n18232 ) ;
  assign n39015 = n8082 & ~n24126 ;
  assign n39016 = n4683 & ~n18277 ;
  assign n39017 = n13852 | n29683 ;
  assign n39018 = n2433 | n24372 ;
  assign n39019 = n24621 | n39018 ;
  assign n39020 = n1968 & ~n2326 ;
  assign n39021 = n39020 ^ n1286 ^ 1'b0 ;
  assign n39022 = n17319 & ~n39021 ;
  assign n39023 = n2433 | n16851 ;
  assign n39024 = n2433 & ~n39023 ;
  assign n39025 = n23290 ^ n16295 ^ 1'b0 ;
  assign n39026 = n39024 | n39025 ;
  assign n39027 = n39026 ^ n21165 ^ 1'b0 ;
  assign n39028 = n39022 & n39027 ;
  assign n39029 = n35057 ^ n5474 ^ 1'b0 ;
  assign n39030 = ~n17087 & n39029 ;
  assign n39031 = n24107 | n27166 ;
  assign n39032 = ~n9247 & n10191 ;
  assign n39033 = n39032 ^ n6126 ^ 1'b0 ;
  assign n39034 = ~n29845 & n39033 ;
  assign n39035 = ~n25580 & n39034 ;
  assign n39036 = n197 & n4849 ;
  assign n39037 = n39036 ^ n2746 ^ 1'b0 ;
  assign n39038 = n6256 & ~n39037 ;
  assign n39039 = n38063 & ~n39038 ;
  assign n39040 = n24799 | n39039 ;
  assign n39041 = n24667 & ~n39040 ;
  assign n39042 = n15009 & ~n20842 ;
  assign n39043 = n39042 ^ n37107 ^ 1'b0 ;
  assign n39044 = n1430 | n2732 ;
  assign n39045 = ( ~n2017 & n17935 ) | ( ~n2017 & n39044 ) | ( n17935 & n39044 ) ;
  assign n39046 = ( ~n1080 & n3790 ) | ( ~n1080 & n5522 ) | ( n3790 & n5522 ) ;
  assign n39047 = n39046 ^ n27816 ^ n9459 ;
  assign n39048 = n5549 & ~n26493 ;
  assign n39049 = ~n2252 & n7570 ;
  assign n39050 = n39049 ^ n34710 ^ 1'b0 ;
  assign n39051 = ~n10242 & n11423 ;
  assign n39052 = n14863 & n39051 ;
  assign n39053 = ~n18355 & n32567 ;
  assign n39054 = n8101 ^ n7891 ^ 1'b0 ;
  assign n39055 = n14716 ^ n9198 ^ n7471 ;
  assign n39056 = n13429 & ~n39055 ;
  assign n39057 = ~n3646 & n39056 ;
  assign n39058 = n39057 ^ n4213 ^ 1'b0 ;
  assign n39059 = n4229 ^ n2735 ^ 1'b0 ;
  assign n39060 = n944 | n39059 ;
  assign n39061 = ( n2755 & n10944 ) | ( n2755 & ~n13776 ) | ( n10944 & ~n13776 ) ;
  assign n39062 = ~n39060 & n39061 ;
  assign n39063 = n4693 | n19835 ;
  assign n39064 = n39063 ^ n13665 ^ 1'b0 ;
  assign n39065 = n39064 ^ n17155 ^ n848 ;
  assign n39066 = n25539 ^ n225 ^ 1'b0 ;
  assign n39067 = n16508 & n24229 ;
  assign n39068 = n39067 ^ n8408 ^ 1'b0 ;
  assign n39069 = n3221 | n39068 ;
  assign n39070 = n5085 & ~n11300 ;
  assign n39071 = n39070 ^ n12867 ^ 1'b0 ;
  assign n39072 = n9952 & ~n39071 ;
  assign n39073 = ~n18961 & n39072 ;
  assign n39074 = n18179 | n34988 ;
  assign n39075 = n6937 & n28959 ;
  assign n39076 = n1853 & n38603 ;
  assign n39077 = n39076 ^ n11481 ^ 1'b0 ;
  assign n39078 = n11898 | n30509 ;
  assign n39079 = n2377 | n39078 ;
  assign n39080 = n11133 & ~n14580 ;
  assign n39081 = ~n39079 & n39080 ;
  assign n39082 = ~n6534 & n7798 ;
  assign n39083 = n7280 | n18192 ;
  assign n39084 = n39083 ^ n3370 ^ 1'b0 ;
  assign n39085 = n39084 ^ n20242 ^ 1'b0 ;
  assign n39086 = n39082 & ~n39085 ;
  assign n39087 = n12131 & n21369 ;
  assign n39088 = ~n14848 & n39087 ;
  assign n39089 = n26871 ^ n15488 ^ 1'b0 ;
  assign n39090 = n6070 & n10656 ;
  assign n39091 = n39090 ^ n9082 ^ 1'b0 ;
  assign n39092 = n22425 ^ n10897 ^ 1'b0 ;
  assign n39093 = n18312 ^ n3310 ^ 1'b0 ;
  assign n39094 = n39092 & n39093 ;
  assign n39095 = n7803 & n39094 ;
  assign n39096 = n24904 ^ n15122 ^ 1'b0 ;
  assign n39097 = ~n14334 & n20128 ;
  assign n39098 = ~n19903 & n39097 ;
  assign n39099 = n9933 & ~n10154 ;
  assign n39100 = n19479 & ~n39099 ;
  assign n39101 = n4886 ^ n4774 ^ 1'b0 ;
  assign n39102 = n11982 & ~n39101 ;
  assign n39103 = ~n18542 & n39102 ;
  assign n39104 = n4856 & n38495 ;
  assign n39105 = ~n2134 & n29938 ;
  assign n39106 = n39105 ^ n28146 ^ 1'b0 ;
  assign n39107 = ( n28865 & ~n35653 ) | ( n28865 & n39106 ) | ( ~n35653 & n39106 ) ;
  assign n39108 = n302 & n6760 ;
  assign n39109 = n3488 & ~n19110 ;
  assign n39110 = n33016 ^ n27873 ^ 1'b0 ;
  assign n39111 = n4857 & ~n39110 ;
  assign n39112 = n13192 ^ n8383 ^ 1'b0 ;
  assign n39113 = n18832 | n39112 ;
  assign n39114 = n39113 ^ n21065 ^ 1'b0 ;
  assign n39115 = n14577 | n19409 ;
  assign n39116 = n4922 | n6583 ;
  assign n39117 = n9906 | n39116 ;
  assign n39118 = ~n13172 & n29421 ;
  assign n39119 = ~n39117 & n39118 ;
  assign n39120 = n3030 & n18696 ;
  assign n39124 = n9606 & n23898 ;
  assign n39121 = n12535 ^ n4741 ^ 1'b0 ;
  assign n39122 = n2721 & ~n39121 ;
  assign n39123 = n16346 & n39122 ;
  assign n39125 = n39124 ^ n39123 ^ 1'b0 ;
  assign n39126 = ~n11959 & n24703 ;
  assign n39128 = n20119 ^ n4234 ^ 1'b0 ;
  assign n39129 = ~n9129 & n39128 ;
  assign n39127 = n14221 & ~n33179 ;
  assign n39130 = n39129 ^ n39127 ^ n25698 ;
  assign n39131 = n2452 & n10333 ;
  assign n39132 = ~n28853 & n39131 ;
  assign n39133 = ( ~n11605 & n30770 ) | ( ~n11605 & n39132 ) | ( n30770 & n39132 ) ;
  assign n39136 = ~n2137 & n24573 ;
  assign n39134 = n2886 & n37357 ;
  assign n39135 = ~n15579 & n39134 ;
  assign n39137 = n39136 ^ n39135 ^ 1'b0 ;
  assign n39138 = ~n5998 & n39137 ;
  assign n39139 = n35595 | n35676 ;
  assign n39140 = n31672 & ~n39139 ;
  assign n39142 = n2504 | n16637 ;
  assign n39141 = n18515 & n27629 ;
  assign n39143 = n39142 ^ n39141 ^ 1'b0 ;
  assign n39144 = n19544 | n33349 ;
  assign n39145 = n15087 ^ n7565 ^ 1'b0 ;
  assign n39146 = n24835 ^ n16414 ^ 1'b0 ;
  assign n39147 = n39145 & n39146 ;
  assign n39148 = n11729 & ~n13320 ;
  assign n39149 = n39148 ^ n22638 ^ 1'b0 ;
  assign n39151 = n8725 ^ n2185 ^ 1'b0 ;
  assign n39152 = n29502 ^ n7031 ^ 1'b0 ;
  assign n39153 = n39151 & n39152 ;
  assign n39154 = n16736 ^ x0 ^ 1'b0 ;
  assign n39155 = ~n39153 & n39154 ;
  assign n39150 = n4033 | n16155 ;
  assign n39156 = n39155 ^ n39150 ^ 1'b0 ;
  assign n39157 = n12980 & n15544 ;
  assign n39158 = n39157 ^ n420 ^ 1'b0 ;
  assign n39159 = n12927 ^ n3243 ^ 1'b0 ;
  assign n39160 = n23048 & n39159 ;
  assign n39161 = n13061 & ~n28119 ;
  assign n39162 = n39161 ^ n27354 ^ 1'b0 ;
  assign n39163 = n2755 & n8986 ;
  assign n39164 = n7923 & n14997 ;
  assign n39165 = n13442 & ~n39164 ;
  assign n39166 = n39165 ^ n23516 ^ 1'b0 ;
  assign n39167 = ( ~n4137 & n12458 ) | ( ~n4137 & n39166 ) | ( n12458 & n39166 ) ;
  assign n39168 = n18351 | n36505 ;
  assign n39169 = ~n93 & n39168 ;
  assign n39170 = n4460 & n24224 ;
  assign n39171 = n241 & ~n8758 ;
  assign n39172 = n39171 ^ n25369 ^ 1'b0 ;
  assign n39173 = n10950 | n37663 ;
  assign n39174 = n24810 & ~n39173 ;
  assign n39175 = n39174 ^ n17737 ^ 1'b0 ;
  assign n39176 = ~n39172 & n39175 ;
  assign n39177 = ~n559 & n5150 ;
  assign n39178 = ~n6716 & n39177 ;
  assign n39179 = n9106 ^ n6164 ^ 1'b0 ;
  assign n39180 = n17422 & ~n39179 ;
  assign n39181 = ~n26582 & n29750 ;
  assign n39182 = n7008 | n13580 ;
  assign n39183 = n32388 & ~n39182 ;
  assign n39184 = ( n5501 & ~n23443 ) | ( n5501 & n31489 ) | ( ~n23443 & n31489 ) ;
  assign n39185 = n2444 | n8906 ;
  assign n39186 = n15130 | n39185 ;
  assign n39187 = n1083 & n24734 ;
  assign n39188 = n19636 ^ n7516 ^ n6441 ;
  assign n39189 = n38021 ^ n27906 ^ n7109 ;
  assign n39190 = n18665 ^ n2467 ^ 1'b0 ;
  assign n39191 = n10689 & ~n39190 ;
  assign n39192 = n22613 | n31256 ;
  assign n39193 = n39192 ^ n22524 ^ 1'b0 ;
  assign n39194 = n30242 ^ n3047 ^ 1'b0 ;
  assign n39195 = n26130 & n39194 ;
  assign n39196 = n5417 & ~n35559 ;
  assign n39197 = n10167 | n29599 ;
  assign n39198 = n21111 & n39197 ;
  assign n39199 = n2784 & ~n16084 ;
  assign n39200 = n18885 ^ n10822 ^ 1'b0 ;
  assign n39201 = n28211 & ~n39200 ;
  assign n39202 = ( n10083 & n10092 ) | ( n10083 & ~n35302 ) | ( n10092 & ~n35302 ) ;
  assign n39203 = n34807 & ~n35992 ;
  assign n39204 = ~n4483 & n39203 ;
  assign n39205 = ~n2353 & n8037 ;
  assign n39206 = n14926 ^ n4722 ^ 1'b0 ;
  assign n39207 = n3229 & n39206 ;
  assign n39208 = n24428 ^ n9875 ^ 1'b0 ;
  assign n39209 = n25761 | n39208 ;
  assign n39210 = n39209 ^ n11635 ^ 1'b0 ;
  assign n39211 = n39210 ^ n19482 ^ n1994 ;
  assign n39212 = n3725 & n3762 ;
  assign n39213 = n39212 ^ n10595 ^ n2758 ;
  assign n39214 = n28601 ^ n12091 ^ 1'b0 ;
  assign n39215 = n2399 & n39214 ;
  assign n39216 = n9765 | n39215 ;
  assign n39217 = n39216 ^ n774 ^ 1'b0 ;
  assign n39218 = ( n846 & ~n1313 ) | ( n846 & n26987 ) | ( ~n1313 & n26987 ) ;
  assign n39219 = n39218 ^ n14651 ^ 1'b0 ;
  assign n39220 = n39219 ^ n20641 ^ 1'b0 ;
  assign n39221 = n22781 ^ n15953 ^ n86 ;
  assign n39222 = n39220 & ~n39221 ;
  assign n39223 = n39222 ^ n682 ^ 1'b0 ;
  assign n39224 = n841 | n7804 ;
  assign n39225 = n39224 ^ n34452 ^ 1'b0 ;
  assign n39226 = n30471 ^ n19638 ^ n18080 ;
  assign n39227 = n7883 & n16508 ;
  assign n39228 = n17001 ^ n7875 ^ 1'b0 ;
  assign n39229 = ( n8695 & n13083 ) | ( n8695 & ~n18784 ) | ( n13083 & ~n18784 ) ;
  assign n39230 = n11805 | n39229 ;
  assign n39231 = n3871 | n39230 ;
  assign n39232 = n17701 & ~n39231 ;
  assign n39233 = n27728 ^ n16321 ^ 1'b0 ;
  assign n39234 = n23606 & ~n39233 ;
  assign n39235 = n37988 ^ n15594 ^ n3694 ;
  assign n39236 = ~n39234 & n39235 ;
  assign n39237 = n7206 & n15659 ;
  assign n39238 = n11458 & n22625 ;
  assign n39239 = n39238 ^ n21125 ^ 1'b0 ;
  assign n39240 = ~n7167 & n7476 ;
  assign n39241 = n39240 ^ n5273 ^ 1'b0 ;
  assign n39242 = n22073 ^ n21346 ^ 1'b0 ;
  assign n39243 = n7204 | n39242 ;
  assign n39244 = n27944 & ~n35825 ;
  assign n39245 = n38621 ^ n38353 ^ 1'b0 ;
  assign n39246 = ~n36352 & n39245 ;
  assign n39247 = n4063 & n16823 ;
  assign n39248 = n36586 ^ n2442 ^ 1'b0 ;
  assign n39249 = n39247 & n39248 ;
  assign n39250 = n25340 ^ n7321 ^ 1'b0 ;
  assign n39251 = n6945 & ~n39250 ;
  assign n39252 = n14544 ^ n10582 ^ 1'b0 ;
  assign n39253 = n1216 & n39252 ;
  assign n39254 = n10640 & n39253 ;
  assign n39255 = n39254 ^ n2309 ^ 1'b0 ;
  assign n39256 = n2376 | n39255 ;
  assign n39257 = n39251 | n39256 ;
  assign n39258 = n14600 & ~n33434 ;
  assign n39259 = n39258 ^ n3708 ^ 1'b0 ;
  assign n39260 = n34893 ^ n25691 ^ 1'b0 ;
  assign n39261 = ~n30404 & n39260 ;
  assign n39262 = n11486 & ~n19173 ;
  assign n39263 = n19173 & n39262 ;
  assign n39264 = n14949 & ~n15817 ;
  assign n39265 = ~n26005 & n39264 ;
  assign n39266 = ~n1973 & n29237 ;
  assign n39267 = n18842 ^ n14758 ^ 1'b0 ;
  assign n39268 = n36007 ^ n24196 ^ 1'b0 ;
  assign n39269 = n19409 | n39268 ;
  assign n39270 = n3755 | n8435 ;
  assign n39271 = n8435 & ~n39270 ;
  assign n39272 = ~n3792 & n39271 ;
  assign n39273 = n30343 | n39272 ;
  assign n39274 = n19702 & n35993 ;
  assign n39275 = ~n28101 & n39274 ;
  assign n39276 = ~n37099 & n39275 ;
  assign n39277 = n7806 & ~n9048 ;
  assign n39278 = n39277 ^ n31884 ^ 1'b0 ;
  assign n39279 = n6282 ^ n1832 ^ 1'b0 ;
  assign n39280 = n39279 ^ n8550 ^ 1'b0 ;
  assign n39281 = ~n39278 & n39280 ;
  assign n39282 = n12544 & n15907 ;
  assign n39283 = n34561 & n39282 ;
  assign n39284 = n21243 | n37646 ;
  assign n39285 = ~n23635 & n28865 ;
  assign n39286 = n1663 & n12576 ;
  assign n39287 = n2853 & n39286 ;
  assign n39288 = n17268 & ~n39287 ;
  assign n39289 = ( ~n18190 & n35824 ) | ( ~n18190 & n39288 ) | ( n35824 & n39288 ) ;
  assign n39290 = ( n7876 & ~n39285 ) | ( n7876 & n39289 ) | ( ~n39285 & n39289 ) ;
  assign n39291 = n6975 | n19182 ;
  assign n39292 = n15406 | n39291 ;
  assign n39293 = n25791 & ~n39292 ;
  assign n39294 = n39293 ^ n15129 ^ 1'b0 ;
  assign n39295 = n30718 ^ n2689 ^ 1'b0 ;
  assign n39296 = n2909 & n39295 ;
  assign n39297 = n27970 & ~n39296 ;
  assign n39298 = n7259 & n10237 ;
  assign n39299 = n26523 & n39298 ;
  assign n39300 = n39299 ^ n11931 ^ 1'b0 ;
  assign n39301 = n2668 & n5147 ;
  assign n39302 = n39301 ^ n11187 ^ 1'b0 ;
  assign n39303 = n31172 ^ n17407 ^ 1'b0 ;
  assign n39304 = x1 & ~n39303 ;
  assign n39305 = n10948 & ~n19933 ;
  assign n39306 = n1853 & n17387 ;
  assign n39307 = n22930 & n39306 ;
  assign n39308 = n34894 ^ n34401 ^ 1'b0 ;
  assign n39309 = n24144 ^ n7744 ^ 1'b0 ;
  assign n39310 = n5986 | n26542 ;
  assign n39311 = n28424 & ~n39310 ;
  assign n39312 = n39311 ^ n30459 ^ 1'b0 ;
  assign n39313 = n9390 & ~n16463 ;
  assign n39314 = ~n24311 & n39313 ;
  assign n39315 = n12230 ^ n4583 ^ 1'b0 ;
  assign n39316 = n24211 ^ n9314 ^ 1'b0 ;
  assign n39317 = n11476 | n39316 ;
  assign n39318 = ( n19455 & n20112 ) | ( n19455 & n21880 ) | ( n20112 & n21880 ) ;
  assign n39319 = n11913 ^ n9542 ^ 1'b0 ;
  assign n39320 = ~n179 & n4823 ;
  assign n39321 = n3985 | n39320 ;
  assign n39322 = n5234 & n24140 ;
  assign n39323 = n22192 & n39322 ;
  assign n39324 = n4733 & n20303 ;
  assign n39325 = n2081 & n39324 ;
  assign n39326 = n2353 | n39325 ;
  assign n39327 = n9153 | n15515 ;
  assign n39328 = n39326 | n39327 ;
  assign n39329 = ( n1821 & n15856 ) | ( n1821 & ~n20233 ) | ( n15856 & ~n20233 ) ;
  assign n39330 = n5132 & n14126 ;
  assign n39331 = n18561 | n26167 ;
  assign n39332 = n39330 | n39331 ;
  assign n39333 = n39332 ^ n12058 ^ 1'b0 ;
  assign n39334 = ~n12921 & n39333 ;
  assign n39336 = n28205 ^ n21981 ^ 1'b0 ;
  assign n39335 = n4976 | n12520 ;
  assign n39337 = n39336 ^ n39335 ^ 1'b0 ;
  assign n39338 = n263 | n39337 ;
  assign n39339 = n1551 & n30277 ;
  assign n39340 = n39339 ^ n29642 ^ 1'b0 ;
  assign n39341 = n39340 ^ n15597 ^ n9518 ;
  assign n39342 = n1023 | n39341 ;
  assign n39343 = n14246 | n39342 ;
  assign n39344 = n32768 ^ n21818 ^ 1'b0 ;
  assign n39346 = n33055 ^ n21509 ^ 1'b0 ;
  assign n39345 = n31380 ^ n31342 ^ 1'b0 ;
  assign n39347 = n39346 ^ n39345 ^ 1'b0 ;
  assign n39348 = n33890 ^ n15928 ^ 1'b0 ;
  assign n39349 = n28634 & n35315 ;
  assign n39350 = n5367 & n39349 ;
  assign n39351 = n29129 ^ n6811 ^ 1'b0 ;
  assign n39352 = n22885 & n39351 ;
  assign n39353 = ~n6885 & n33560 ;
  assign n39354 = n2346 & ~n3818 ;
  assign n39355 = n11929 ^ n2184 ^ 1'b0 ;
  assign n39356 = n1187 & n31806 ;
  assign n39357 = n11570 & ~n34044 ;
  assign n39358 = ~n22983 & n39357 ;
  assign n39359 = n1369 | n2806 ;
  assign n39360 = n2806 & ~n39359 ;
  assign n39361 = n28513 ^ n20864 ^ 1'b0 ;
  assign n39362 = n39361 ^ n18731 ^ 1'b0 ;
  assign n39363 = n39360 | n39362 ;
  assign n39365 = n8230 & n20393 ;
  assign n39364 = n11234 & n15217 ;
  assign n39366 = n39365 ^ n39364 ^ 1'b0 ;
  assign n39367 = n39366 ^ n23675 ^ n4081 ;
  assign n39368 = n39367 ^ n270 ^ 1'b0 ;
  assign n39369 = n3636 ^ n1724 ^ 1'b0 ;
  assign n39370 = ~n19664 & n39369 ;
  assign n39371 = n5385 ^ n1167 ^ 1'b0 ;
  assign n39372 = n35822 ^ n33059 ^ 1'b0 ;
  assign n39373 = n16010 & ~n39372 ;
  assign n39374 = ~n39371 & n39373 ;
  assign n39375 = n15423 ^ n8827 ^ 1'b0 ;
  assign n39376 = n4405 ^ n1574 ^ 1'b0 ;
  assign n39377 = n15267 ^ n11292 ^ 1'b0 ;
  assign n39378 = n7003 | n39377 ;
  assign n39379 = n4355 & ~n39378 ;
  assign n39380 = n39379 ^ n13491 ^ 1'b0 ;
  assign n39381 = n26384 & ~n39380 ;
  assign n39383 = ~n800 & n5417 ;
  assign n39384 = n39383 ^ n885 ^ 1'b0 ;
  assign n39385 = n39384 ^ n19780 ^ 1'b0 ;
  assign n39386 = n12862 | n39385 ;
  assign n39387 = n39386 ^ n25707 ^ 1'b0 ;
  assign n39382 = ~n2486 & n37985 ;
  assign n39388 = n39387 ^ n39382 ^ 1'b0 ;
  assign n39389 = n35559 ^ n4256 ^ 1'b0 ;
  assign n39390 = n3647 & ~n26288 ;
  assign n39391 = n2853 | n31223 ;
  assign n39392 = n39391 ^ n4359 ^ 1'b0 ;
  assign n39393 = n14208 ^ n2630 ^ 1'b0 ;
  assign n39396 = n19114 ^ n12472 ^ 1'b0 ;
  assign n39397 = n6714 & n39396 ;
  assign n39394 = n2980 & n28616 ;
  assign n39395 = n39394 ^ n4250 ^ 1'b0 ;
  assign n39398 = n39397 ^ n39395 ^ 1'b0 ;
  assign n39399 = ( ~n2094 & n6213 ) | ( ~n2094 & n16423 ) | ( n6213 & n16423 ) ;
  assign n39400 = n1961 | n39399 ;
  assign n39401 = n23363 & ~n39400 ;
  assign n39402 = ~n14153 & n39401 ;
  assign n39403 = n39402 ^ n35972 ^ 1'b0 ;
  assign n39404 = n39398 | n39403 ;
  assign n39405 = n16881 | n21623 ;
  assign n39406 = n25685 ^ n15541 ^ 1'b0 ;
  assign n39407 = ~n39405 & n39406 ;
  assign n39408 = n5813 & n22613 ;
  assign n39409 = ( n3442 & n11597 ) | ( n3442 & ~n17116 ) | ( n11597 & ~n17116 ) ;
  assign n39410 = n9715 & n27407 ;
  assign n39411 = n9183 ^ n892 ^ 1'b0 ;
  assign n39412 = ( ~n4483 & n14670 ) | ( ~n4483 & n39411 ) | ( n14670 & n39411 ) ;
  assign n39413 = n39412 ^ n4991 ^ 1'b0 ;
  assign n39414 = ~n17162 & n39413 ;
  assign n39415 = n3696 & ~n7682 ;
  assign n39416 = n27709 & ~n39415 ;
  assign n39417 = n12008 & n17206 ;
  assign n39418 = n39416 & n39417 ;
  assign n39419 = n11276 ^ n3968 ^ 1'b0 ;
  assign n39420 = ( n271 & ~n22340 ) | ( n271 & n39419 ) | ( ~n22340 & n39419 ) ;
  assign n39421 = n14284 & ~n15099 ;
  assign n39422 = n39421 ^ n5365 ^ 1'b0 ;
  assign n39423 = n31519 ^ n25757 ^ 1'b0 ;
  assign n39424 = n39422 | n39423 ;
  assign n39425 = n4888 & n7495 ;
  assign n39426 = n39425 ^ n18781 ^ 1'b0 ;
  assign n39427 = n1374 & n28544 ;
  assign n39428 = n2206 & n6714 ;
  assign n39429 = n2258 | n28911 ;
  assign n39430 = n13131 ^ n2008 ^ 1'b0 ;
  assign n39431 = n16795 & ~n39430 ;
  assign n39432 = n14614 & ~n29526 ;
  assign n39433 = ~n9023 & n39432 ;
  assign n39434 = n4519 | n6943 ;
  assign n39436 = n16681 ^ n10728 ^ 1'b0 ;
  assign n39437 = n13318 & n34210 ;
  assign n39438 = n39436 | n39437 ;
  assign n39435 = n10306 | n25215 ;
  assign n39439 = n39438 ^ n39435 ^ 1'b0 ;
  assign n39440 = ~n29387 & n39439 ;
  assign n39441 = ( ~n1071 & n3646 ) | ( ~n1071 & n11024 ) | ( n3646 & n11024 ) ;
  assign n39442 = n29842 & ~n39441 ;
  assign n39443 = n39442 ^ n5150 ^ 1'b0 ;
  assign n39444 = n39443 ^ n3384 ^ 1'b0 ;
  assign n39445 = n14372 & n21209 ;
  assign n39446 = n39445 ^ n9116 ^ 1'b0 ;
  assign n39447 = n15394 ^ n10612 ^ 1'b0 ;
  assign n39448 = ~n37756 & n39447 ;
  assign n39449 = n23136 & n33109 ;
  assign n39450 = ~n12972 & n39449 ;
  assign n39451 = ( n4170 & ~n39448 ) | ( n4170 & n39450 ) | ( ~n39448 & n39450 ) ;
  assign n39452 = n39451 ^ n27060 ^ 1'b0 ;
  assign n39453 = n1285 & ~n24211 ;
  assign n39454 = ~n17099 & n39453 ;
  assign n39456 = ~n6878 & n12899 ;
  assign n39457 = n39456 ^ n2183 ^ 1'b0 ;
  assign n39458 = ~n12008 & n39457 ;
  assign n39455 = n9589 & n27082 ;
  assign n39459 = n39458 ^ n39455 ^ 1'b0 ;
  assign n39460 = n3403 & ~n23167 ;
  assign n39461 = n29909 ^ n13687 ^ 1'b0 ;
  assign n39462 = n8616 | n39461 ;
  assign n39463 = n39462 ^ n559 ^ 1'b0 ;
  assign n39464 = ~n39460 & n39463 ;
  assign n39465 = n277 | n2755 ;
  assign n39466 = n39465 ^ n31967 ^ 1'b0 ;
  assign n39467 = n32807 ^ n1308 ^ 1'b0 ;
  assign n39468 = n9261 & n39467 ;
  assign n39469 = n38638 ^ n21260 ^ 1'b0 ;
  assign n39470 = n18585 & n39469 ;
  assign n39471 = n13445 | n21993 ;
  assign n39472 = n39471 ^ n343 ^ 1'b0 ;
  assign n39473 = n11338 ^ n528 ^ 1'b0 ;
  assign n39474 = n39473 ^ n4644 ^ 1'b0 ;
  assign n39475 = ( ~n7462 & n18450 ) | ( ~n7462 & n39474 ) | ( n18450 & n39474 ) ;
  assign n39476 = n6302 & ~n9899 ;
  assign n39477 = n39476 ^ n13878 ^ 1'b0 ;
  assign n39478 = n10720 ^ n2872 ^ 1'b0 ;
  assign n39479 = n1976 & n32322 ;
  assign n39480 = n39479 ^ n26849 ^ n13884 ;
  assign n39481 = ( n21059 & n39478 ) | ( n21059 & n39480 ) | ( n39478 & n39480 ) ;
  assign n39482 = n6185 | n8735 ;
  assign n39483 = n39481 & ~n39482 ;
  assign n39484 = n2632 & n3556 ;
  assign n39485 = n39484 ^ n11727 ^ 1'b0 ;
  assign n39486 = n2791 | n39485 ;
  assign n39487 = n2583 | n4526 ;
  assign n39488 = n39487 ^ n20936 ^ 1'b0 ;
  assign n39489 = n17902 & n23243 ;
  assign n39490 = ~n12825 & n39489 ;
  assign n39491 = n9865 | n26312 ;
  assign n39492 = n39490 & ~n39491 ;
  assign n39493 = ~n10321 & n16969 ;
  assign n39494 = n6716 & n39493 ;
  assign n39495 = n39492 & n39494 ;
  assign n39496 = n35695 ^ n22862 ^ 1'b0 ;
  assign n39497 = n25112 & ~n39496 ;
  assign n39498 = ~n8312 & n8368 ;
  assign n39499 = n37105 ^ n22825 ^ 1'b0 ;
  assign n39500 = n39498 | n39499 ;
  assign n39501 = n39500 ^ n33162 ^ 1'b0 ;
  assign n39502 = ( n608 & ~n4408 ) | ( n608 & n18812 ) | ( ~n4408 & n18812 ) ;
  assign n39503 = n16847 ^ n2173 ^ 1'b0 ;
  assign n39504 = n20251 & n39503 ;
  assign n39505 = n14469 ^ n3572 ^ 1'b0 ;
  assign n39506 = n10628 | n39505 ;
  assign n39507 = n13279 ^ n8602 ^ 1'b0 ;
  assign n39508 = n780 | n798 ;
  assign n39509 = n11371 | n39508 ;
  assign n39510 = ~n37282 & n39509 ;
  assign n39511 = n37230 ^ n27641 ^ n22148 ;
  assign n39512 = n32410 ^ n17903 ^ n4478 ;
  assign n39513 = n27238 ^ n24217 ^ 1'b0 ;
  assign n39514 = ( n4106 & n14677 ) | ( n4106 & ~n21324 ) | ( n14677 & ~n21324 ) ;
  assign n39515 = n175 | n25671 ;
  assign n39516 = n9231 & ~n39515 ;
  assign n39517 = ~n39514 & n39516 ;
  assign n39518 = n8053 ^ n609 ^ 1'b0 ;
  assign n39519 = n3105 & n39518 ;
  assign n39520 = n7703 & ~n27224 ;
  assign n39521 = n27130 ^ n24692 ^ 1'b0 ;
  assign n39522 = ~n19202 & n39521 ;
  assign n39523 = n39522 ^ n33818 ^ 1'b0 ;
  assign n39527 = n7437 ^ n3437 ^ 1'b0 ;
  assign n39524 = ( n8104 & n9156 ) | ( n8104 & n19921 ) | ( n9156 & n19921 ) ;
  assign n39525 = n39524 ^ n3445 ^ 1'b0 ;
  assign n39526 = n24150 | n39525 ;
  assign n39528 = n39527 ^ n39526 ^ 1'b0 ;
  assign n39529 = ~n4344 & n12438 ;
  assign n39530 = n39529 ^ n21934 ^ 1'b0 ;
  assign n39531 = n26276 ^ n601 ^ 1'b0 ;
  assign n39532 = ( ~n2347 & n2754 ) | ( ~n2347 & n4006 ) | ( n2754 & n4006 ) ;
  assign n39533 = n12023 & ~n37087 ;
  assign n39534 = ~n34334 & n39533 ;
  assign n39535 = n13493 ^ n11137 ^ 1'b0 ;
  assign n39536 = n4802 ^ n4593 ^ 1'b0 ;
  assign n39537 = n16364 & n39536 ;
  assign n39538 = n2563 & ~n28779 ;
  assign n39539 = n39537 & n39538 ;
  assign n39540 = n39539 ^ n3626 ^ 1'b0 ;
  assign n39541 = ~n750 & n17582 ;
  assign n39542 = ~n2587 & n39541 ;
  assign n39543 = n16617 | n22154 ;
  assign n39544 = n5057 ^ n4088 ^ 1'b0 ;
  assign n39545 = n6305 & n25104 ;
  assign n39546 = n11826 | n15415 ;
  assign n39547 = n39546 ^ n181 ^ 1'b0 ;
  assign n39548 = n14748 ^ n7348 ^ 1'b0 ;
  assign n39549 = n20739 & ~n39548 ;
  assign n39550 = n28159 ^ n9177 ^ 1'b0 ;
  assign n39551 = n574 | n39550 ;
  assign n39552 = n13311 ^ n12487 ^ 1'b0 ;
  assign n39553 = ~n581 & n25874 ;
  assign n39554 = ~n39552 & n39553 ;
  assign n39555 = n867 & ~n39554 ;
  assign n39556 = n7966 & n17497 ;
  assign n39557 = n13266 ^ n6176 ^ 1'b0 ;
  assign n39558 = n21054 | n39557 ;
  assign n39559 = n38403 ^ n34468 ^ n11655 ;
  assign n39560 = n37978 ^ n2657 ^ 1'b0 ;
  assign n39561 = ~n8792 & n32135 ;
  assign n39562 = n39561 ^ n805 ^ 1'b0 ;
  assign n39563 = n20002 | n39562 ;
  assign n39564 = n39563 ^ n15424 ^ n11726 ;
  assign n39565 = ~n243 & n4914 ;
  assign n39566 = ( n7100 & n11313 ) | ( n7100 & n39565 ) | ( n11313 & n39565 ) ;
  assign n39568 = n9222 ^ n1921 ^ 1'b0 ;
  assign n39569 = n26613 | n39568 ;
  assign n39567 = n1517 | n17477 ;
  assign n39570 = n39569 ^ n39567 ^ 1'b0 ;
  assign n39571 = n33683 ^ n33136 ^ 1'b0 ;
  assign n39572 = n19707 & n39571 ;
  assign n39573 = n8436 & ~n16511 ;
  assign n39574 = n39573 ^ n344 ^ 1'b0 ;
  assign n39575 = n8465 ^ n8366 ^ 1'b0 ;
  assign n39576 = n39574 & ~n39575 ;
  assign n39577 = n15492 & ~n16340 ;
  assign n39578 = n39577 ^ n11648 ^ 1'b0 ;
  assign n39579 = n4059 & ~n16404 ;
  assign n39580 = ~n39578 & n39579 ;
  assign n39581 = n3345 | n6184 ;
  assign n39582 = n39581 ^ n1196 ^ 1'b0 ;
  assign n39583 = ~n39580 & n39582 ;
  assign n39584 = n980 ^ n614 ^ n536 ;
  assign n39585 = n17493 & n21506 ;
  assign n39586 = ~n263 & n39585 ;
  assign n39587 = n9667 ^ n2022 ^ 1'b0 ;
  assign n39588 = ~n31623 & n39587 ;
  assign n39589 = n590 | n1208 ;
  assign n39590 = n39589 ^ n8604 ^ 1'b0 ;
  assign n39591 = n25034 & ~n39590 ;
  assign n39592 = n39591 ^ n30367 ^ 1'b0 ;
  assign n39593 = n39592 ^ n30272 ^ 1'b0 ;
  assign n39594 = n21650 & ~n39593 ;
  assign n39595 = n39594 ^ n25824 ^ 1'b0 ;
  assign n39596 = n19013 & n21277 ;
  assign n39597 = ~n14351 & n20611 ;
  assign n39598 = n39597 ^ n21293 ^ 1'b0 ;
  assign n39599 = n470 | n37156 ;
  assign n39600 = ~n938 & n38981 ;
  assign n39601 = n39600 ^ n22776 ^ 1'b0 ;
  assign n39602 = n2954 & ~n10428 ;
  assign n39603 = n15940 ^ n286 ^ 1'b0 ;
  assign n39604 = n32346 ^ n27757 ^ n13376 ;
  assign n39605 = n39604 ^ n17891 ^ 1'b0 ;
  assign n39606 = ~n14249 & n17245 ;
  assign n39607 = n6972 | n39606 ;
  assign n39608 = n14343 ^ n3034 ^ 1'b0 ;
  assign n39609 = n39608 ^ n10913 ^ 1'b0 ;
  assign n39610 = ~n21772 & n39609 ;
  assign n39611 = ( n33446 & n39607 ) | ( n33446 & n39610 ) | ( n39607 & n39610 ) ;
  assign n39612 = ~n6410 & n33110 ;
  assign n39613 = ~n25956 & n39612 ;
  assign n39614 = n1528 | n22177 ;
  assign n39615 = n37342 ^ n22888 ^ 1'b0 ;
  assign n39616 = n28538 & ~n39615 ;
  assign n39617 = n39614 & n39616 ;
  assign n39618 = n10025 ^ n47 ^ 1'b0 ;
  assign n39619 = ~n1694 & n19060 ;
  assign n39620 = n39619 ^ n14429 ^ 1'b0 ;
  assign n39621 = n25252 ^ n6470 ^ 1'b0 ;
  assign n39622 = ( n2290 & n19027 ) | ( n2290 & n28341 ) | ( n19027 & n28341 ) ;
  assign n39623 = ~n32301 & n33533 ;
  assign n39624 = n37714 & n39623 ;
  assign n39625 = n6151 | n10003 ;
  assign n39626 = n39625 ^ n3315 ^ 1'b0 ;
  assign n39627 = ~n14378 & n39626 ;
  assign n39628 = n31102 & ~n39627 ;
  assign n39630 = n3301 ^ n199 ^ 1'b0 ;
  assign n39629 = n22556 & n30551 ;
  assign n39631 = n39630 ^ n39629 ^ 1'b0 ;
  assign n39632 = n9503 ^ n8898 ^ 1'b0 ;
  assign n39633 = ~n24722 & n39632 ;
  assign n39634 = n15230 & n39633 ;
  assign n39635 = n6609 & n38455 ;
  assign n39636 = n19008 | n33872 ;
  assign n39637 = n1742 ^ n982 ^ 1'b0 ;
  assign n39638 = ~n5689 & n39637 ;
  assign n39639 = n39638 ^ n2428 ^ 1'b0 ;
  assign n39640 = ~n2649 & n39639 ;
  assign n39641 = n21427 & ~n39479 ;
  assign n39642 = n18019 | n36017 ;
  assign n39643 = ~n1186 & n30432 ;
  assign n39644 = n29057 & n39643 ;
  assign n39645 = n39644 ^ n22289 ^ 1'b0 ;
  assign n39646 = n6435 | n31916 ;
  assign n39647 = n12750 | n39646 ;
  assign n39648 = n37303 ^ n8459 ^ 1'b0 ;
  assign n39649 = ~n7007 & n14276 ;
  assign n39650 = n26926 & n39649 ;
  assign n39651 = n8201 ^ n4610 ^ 1'b0 ;
  assign n39652 = n39651 ^ n22158 ^ 1'b0 ;
  assign n39653 = n4757 & n39652 ;
  assign n39654 = n39653 ^ n19215 ^ 1'b0 ;
  assign n39655 = n26658 ^ n4926 ^ 1'b0 ;
  assign n39656 = n7952 & ~n19225 ;
  assign n39657 = n23555 & n39656 ;
  assign n39660 = n13318 ^ n4863 ^ n2980 ;
  assign n39658 = ( n5268 & ~n7342 ) | ( n5268 & n12656 ) | ( ~n7342 & n12656 ) ;
  assign n39659 = ~n13162 & n39658 ;
  assign n39661 = n39660 ^ n39659 ^ 1'b0 ;
  assign n39662 = ~n14735 & n24955 ;
  assign n39663 = ~n105 & n39662 ;
  assign n39664 = n39663 ^ n29893 ^ n11664 ;
  assign n39665 = n32810 & ~n39664 ;
  assign n39666 = n2257 ^ n1050 ^ 1'b0 ;
  assign n39667 = ~n4039 & n39666 ;
  assign n39668 = n39667 ^ n451 ^ 1'b0 ;
  assign n39669 = n20540 | n39668 ;
  assign n39670 = ( n18660 & ~n20325 ) | ( n18660 & n39669 ) | ( ~n20325 & n39669 ) ;
  assign n39671 = n578 & n9760 ;
  assign n39672 = n39671 ^ n5938 ^ 1'b0 ;
  assign n39673 = n16052 & ~n39672 ;
  assign n39674 = ~n205 & n39673 ;
  assign n39675 = n4260 ^ n1445 ^ 1'b0 ;
  assign n39676 = n12090 & ~n39675 ;
  assign n39677 = n35293 ^ n19810 ^ 1'b0 ;
  assign n39678 = n4004 | n39677 ;
  assign n39679 = n39678 ^ n4741 ^ 1'b0 ;
  assign n39680 = n36000 ^ n5789 ^ 1'b0 ;
  assign n39681 = ~n25909 & n39680 ;
  assign n39682 = n28879 ^ n13772 ^ 1'b0 ;
  assign n39683 = n39681 & n39682 ;
  assign n39684 = n15997 | n39174 ;
  assign n39685 = n13183 ^ n3981 ^ 1'b0 ;
  assign n39686 = n13267 & n39685 ;
  assign n39687 = n39686 ^ n29827 ^ 1'b0 ;
  assign n39688 = n2193 & n39687 ;
  assign n39689 = ~n15061 & n39688 ;
  assign n39690 = n13292 ^ n299 ^ 1'b0 ;
  assign n39691 = n39690 ^ n6385 ^ 1'b0 ;
  assign n39692 = n37320 & n39691 ;
  assign n39693 = n18607 ^ n1694 ^ 1'b0 ;
  assign n39694 = n22634 & n39693 ;
  assign n39695 = n25289 ^ n2326 ^ 1'b0 ;
  assign n39696 = n4053 | n39695 ;
  assign n39697 = n1227 & n25217 ;
  assign n39698 = n39697 ^ n10189 ^ 1'b0 ;
  assign n39699 = n10246 ^ n2087 ^ 1'b0 ;
  assign n39700 = ( n6013 & n10879 ) | ( n6013 & n36352 ) | ( n10879 & n36352 ) ;
  assign n39701 = n4241 & n5734 ;
  assign n39702 = n39701 ^ n1783 ^ 1'b0 ;
  assign n39703 = n12890 | n14863 ;
  assign n39704 = n39703 ^ n22646 ^ 1'b0 ;
  assign n39705 = n6898 & n21324 ;
  assign n39706 = n39705 ^ n38342 ^ 1'b0 ;
  assign n39707 = n619 & ~n15876 ;
  assign n39708 = n12283 & n39707 ;
  assign n39709 = ~n13879 & n39708 ;
  assign n39710 = n39709 ^ n24305 ^ n3438 ;
  assign n39711 = n492 | n9419 ;
  assign n39712 = n4555 & ~n17370 ;
  assign n39713 = n39712 ^ n20475 ^ 1'b0 ;
  assign n39714 = n12269 & n39713 ;
  assign n39715 = n5021 & ~n26212 ;
  assign n39716 = n17190 & ~n24523 ;
  assign n39717 = n13557 ^ n423 ^ 1'b0 ;
  assign n39718 = n11815 ^ n7292 ^ 1'b0 ;
  assign n39719 = ~n14523 & n39718 ;
  assign n39720 = ~n12283 & n19144 ;
  assign n39721 = n39720 ^ n4019 ^ 1'b0 ;
  assign n39722 = n25196 ^ n9912 ^ 1'b0 ;
  assign n39723 = n39721 & ~n39722 ;
  assign n39724 = n6527 & n39723 ;
  assign n39725 = n39724 ^ n22418 ^ 1'b0 ;
  assign n39726 = n13844 ^ n8070 ^ 1'b0 ;
  assign n39729 = n363 & n2322 ;
  assign n39727 = n1363 & n5393 ;
  assign n39728 = ~n8523 & n39727 ;
  assign n39730 = n39729 ^ n39728 ^ 1'b0 ;
  assign n39731 = n20614 ^ n1991 ^ 1'b0 ;
  assign n39732 = ~n39730 & n39731 ;
  assign n39733 = n39341 ^ n22943 ^ 1'b0 ;
  assign n39734 = n5547 & n39733 ;
  assign n39735 = ~n11235 & n21596 ;
  assign n39736 = n39735 ^ n12628 ^ 1'b0 ;
  assign n39737 = ~n38363 & n39736 ;
  assign n39738 = ~n39734 & n39737 ;
  assign n39739 = n1023 | n36136 ;
  assign n39740 = n7425 & ~n39739 ;
  assign n39741 = ( ~n3264 & n15578 ) | ( ~n3264 & n28259 ) | ( n15578 & n28259 ) ;
  assign n39742 = ~n11266 & n13323 ;
  assign n39743 = n39742 ^ n11008 ^ 1'b0 ;
  assign n39744 = n12972 & n20270 ;
  assign n39745 = n39744 ^ n27403 ^ 1'b0 ;
  assign n39746 = n29742 ^ n14765 ^ 1'b0 ;
  assign n39747 = n25796 & ~n39746 ;
  assign n39748 = n20659 & ~n29208 ;
  assign n39749 = n21200 ^ n8060 ^ 1'b0 ;
  assign n39750 = n33380 ^ n5473 ^ 1'b0 ;
  assign n39751 = n24890 ^ n2531 ^ 1'b0 ;
  assign n39752 = n16596 | n27705 ;
  assign n39753 = n24540 ^ n10117 ^ n1204 ;
  assign n39754 = n8871 ^ n7287 ^ 1'b0 ;
  assign n39755 = n33593 | n39754 ;
  assign n39756 = n22277 ^ n8880 ^ 1'b0 ;
  assign n39757 = n18037 ^ n611 ^ 1'b0 ;
  assign n39758 = n26335 ^ n5439 ^ 1'b0 ;
  assign n39759 = n12758 & n39758 ;
  assign n39760 = ~n8482 & n11876 ;
  assign n39761 = ~n6524 & n28785 ;
  assign n39762 = ~n6233 & n17584 ;
  assign n39763 = n39762 ^ n10883 ^ 1'b0 ;
  assign n39764 = n6258 | n14563 ;
  assign n39765 = ~n39763 & n39764 ;
  assign n39766 = n32840 & n39765 ;
  assign n39767 = ( n1047 & n5612 ) | ( n1047 & ~n13488 ) | ( n5612 & ~n13488 ) ;
  assign n39768 = n28352 & n39767 ;
  assign n39769 = n163 | n5893 ;
  assign n39770 = ( n6954 & ~n11757 ) | ( n6954 & n39769 ) | ( ~n11757 & n39769 ) ;
  assign n39771 = n8037 ^ n831 ^ 1'b0 ;
  assign n39772 = n39771 ^ n15491 ^ 1'b0 ;
  assign n39773 = ~n3323 & n39772 ;
  assign n39774 = n18319 ^ n12425 ^ 1'b0 ;
  assign n39775 = ~n10581 & n12593 ;
  assign n39776 = n39775 ^ n30997 ^ 1'b0 ;
  assign n39777 = n39776 ^ n373 ^ 1'b0 ;
  assign n39778 = ~n16613 & n28913 ;
  assign n39779 = n18083 & n39778 ;
  assign n39780 = ~n16206 & n18393 ;
  assign n39781 = n39780 ^ n5704 ^ 1'b0 ;
  assign n39782 = n39781 ^ n5289 ^ n4148 ;
  assign n39783 = n24051 ^ n132 ^ 1'b0 ;
  assign n39784 = ~n30350 & n39783 ;
  assign n39785 = n5172 | n10264 ;
  assign n39786 = n7137 & ~n39785 ;
  assign n39787 = n17640 ^ n1563 ^ 1'b0 ;
  assign n39788 = n39787 ^ n10721 ^ n1122 ;
  assign n39789 = ~n6623 & n7095 ;
  assign n39790 = ~n5475 & n39789 ;
  assign n39791 = n16847 ^ n14213 ^ 1'b0 ;
  assign n39792 = ~n323 & n39791 ;
  assign n39793 = ~n39790 & n39792 ;
  assign n39795 = n22556 ^ n15268 ^ 1'b0 ;
  assign n39796 = n23580 & n39795 ;
  assign n39794 = n1337 | n7617 ;
  assign n39797 = n39796 ^ n39794 ^ 1'b0 ;
  assign n39798 = n37224 ^ n18572 ^ 1'b0 ;
  assign n39799 = n39797 & n39798 ;
  assign n39800 = n4012 & n8295 ;
  assign n39801 = n14259 & n39800 ;
  assign n39803 = n2732 & ~n2980 ;
  assign n39802 = n5893 | n8461 ;
  assign n39804 = n39803 ^ n39802 ^ 1'b0 ;
  assign n39805 = n38155 ^ n4838 ^ 1'b0 ;
  assign n39806 = n17081 & ~n18092 ;
  assign n39808 = n754 | n1398 ;
  assign n39807 = ~n597 & n29038 ;
  assign n39809 = n39808 ^ n39807 ^ 1'b0 ;
  assign n39810 = n15406 ^ n6600 ^ 1'b0 ;
  assign n39811 = n5237 & ~n39810 ;
  assign n39812 = n20102 | n35594 ;
  assign n39813 = n2790 | n33226 ;
  assign n39814 = n39813 ^ n20322 ^ 1'b0 ;
  assign n39815 = n5656 & n6297 ;
  assign n39816 = ~n1700 & n8717 ;
  assign n39817 = n29466 & n39816 ;
  assign n39818 = n23468 ^ n22080 ^ 1'b0 ;
  assign n39819 = ~n39817 & n39818 ;
  assign n39820 = n11819 ^ n7744 ^ 1'b0 ;
  assign n39821 = n16299 & n18809 ;
  assign n39822 = ~n39820 & n39821 ;
  assign n39823 = n11175 & n11503 ;
  assign n39824 = n39823 ^ n34468 ^ n11356 ;
  assign n39825 = n18585 ^ n9854 ^ 1'b0 ;
  assign n39826 = n1054 | n39825 ;
  assign n39827 = n34039 | n39826 ;
  assign n39828 = ( n5395 & ~n21348 ) | ( n5395 & n28851 ) | ( ~n21348 & n28851 ) ;
  assign n39829 = n1763 | n39828 ;
  assign n39830 = n2272 ^ n831 ^ 1'b0 ;
  assign n39831 = n14295 & ~n39830 ;
  assign n39832 = n39831 ^ n19710 ^ 1'b0 ;
  assign n39833 = ~n1306 & n39832 ;
  assign n39834 = n36577 ^ n21240 ^ n10729 ;
  assign n39835 = n39834 ^ n3194 ^ 1'b0 ;
  assign n39836 = n12039 ^ n11273 ^ 1'b0 ;
  assign n39837 = n18020 | n39836 ;
  assign n39838 = n39837 ^ n5449 ^ 1'b0 ;
  assign n39839 = n32280 ^ n25498 ^ 1'b0 ;
  assign n39840 = n9423 & ~n39839 ;
  assign n39841 = n1843 & n7494 ;
  assign n39842 = n23220 ^ n14420 ^ 1'b0 ;
  assign n39843 = n5547 | n39842 ;
  assign n39844 = ( n16096 & n31192 ) | ( n16096 & n39843 ) | ( n31192 & n39843 ) ;
  assign n39845 = n39841 | n39844 ;
  assign n39846 = n7876 & ~n19264 ;
  assign n39847 = n14959 & ~n19094 ;
  assign n39848 = n39847 ^ n3665 ^ 1'b0 ;
  assign n39849 = n39848 ^ n27443 ^ 1'b0 ;
  assign n39850 = n33879 & n39849 ;
  assign n39852 = n8787 & n15424 ;
  assign n39851 = n17566 ^ n15198 ^ 1'b0 ;
  assign n39853 = n39852 ^ n39851 ^ n8098 ;
  assign n39854 = n16197 | n25429 ;
  assign n39855 = ( n10345 & ~n24007 ) | ( n10345 & n39854 ) | ( ~n24007 & n39854 ) ;
  assign n39856 = n4448 & n28870 ;
  assign n39857 = n39856 ^ n18059 ^ 1'b0 ;
  assign n39858 = n39061 | n39857 ;
  assign n39859 = n32629 ^ n23905 ^ n22577 ;
  assign n39860 = n16556 & ~n39859 ;
  assign n39861 = n223 & ~n10023 ;
  assign n39862 = ~n6035 & n39861 ;
  assign n39863 = n39862 ^ n22888 ^ 1'b0 ;
  assign n39864 = n23546 ^ n21682 ^ 1'b0 ;
  assign n39865 = n6121 & ~n39864 ;
  assign n39866 = n39863 & n39865 ;
  assign n39873 = ( ~n1010 & n1199 ) | ( ~n1010 & n7560 ) | ( n1199 & n7560 ) ;
  assign n39874 = n21520 & n39873 ;
  assign n39875 = n21501 & n39874 ;
  assign n39867 = n22714 ^ n8427 ^ 1'b0 ;
  assign n39868 = n21498 & n27136 ;
  assign n39869 = n39867 & n39868 ;
  assign n39870 = n14491 | n39869 ;
  assign n39871 = n39870 ^ n1703 ^ 1'b0 ;
  assign n39872 = n30582 & ~n39871 ;
  assign n39876 = n39875 ^ n39872 ^ 1'b0 ;
  assign n39877 = n29208 ^ n21582 ^ 1'b0 ;
  assign n39878 = ( n27117 & ~n38568 ) | ( n27117 & n39877 ) | ( ~n38568 & n39877 ) ;
  assign n39879 = n535 & ~n9907 ;
  assign n39880 = n33759 & ~n39879 ;
  assign n39881 = n4085 & n6542 ;
  assign n39882 = ~n7722 & n18783 ;
  assign n39884 = ~n10886 & n26461 ;
  assign n39883 = n26229 & n27497 ;
  assign n39885 = n39884 ^ n39883 ^ 1'b0 ;
  assign n39886 = n38693 ^ n33265 ^ n17490 ;
  assign n39887 = ~n3663 & n39886 ;
  assign n39888 = n39887 ^ n37013 ^ 1'b0 ;
  assign n39889 = n10913 ^ n7948 ^ 1'b0 ;
  assign n39890 = n1471 & ~n29975 ;
  assign n39891 = n39889 & n39890 ;
  assign n39892 = n451 & ~n3723 ;
  assign n39893 = ~n18983 & n31865 ;
  assign n39894 = n20903 ^ n11789 ^ 1'b0 ;
  assign n39895 = n7951 & ~n39894 ;
  assign n39896 = n17513 & ~n39895 ;
  assign n39897 = n29544 ^ n27164 ^ n16217 ;
  assign n39898 = n39897 ^ n31744 ^ n19675 ;
  assign n39899 = n2328 & ~n25239 ;
  assign n39900 = ~n19941 & n39899 ;
  assign n39901 = n39900 ^ n26249 ^ 1'b0 ;
  assign n39902 = n9086 & n20724 ;
  assign n39903 = n39902 ^ n6345 ^ 1'b0 ;
  assign n39904 = n15698 ^ n5697 ^ 1'b0 ;
  assign n39905 = n3896 | n9102 ;
  assign n39906 = n37278 ^ n15690 ^ 1'b0 ;
  assign n39907 = n13173 ^ n5630 ^ 1'b0 ;
  assign n39908 = n2835 & n26829 ;
  assign n39910 = n20875 ^ n12658 ^ n8515 ;
  assign n39909 = n782 & n4319 ;
  assign n39911 = n39910 ^ n39909 ^ 1'b0 ;
  assign n39912 = n1455 & ~n2340 ;
  assign n39913 = n39912 ^ n15834 ^ 1'b0 ;
  assign n39914 = n34006 | n39913 ;
  assign n39915 = n8199 & ~n10691 ;
  assign n39916 = ~n13233 & n39915 ;
  assign n39917 = n16482 ^ n13470 ^ 1'b0 ;
  assign n39918 = n24694 | n34961 ;
  assign n39919 = ~n13750 & n39638 ;
  assign n39920 = ~n37110 & n39919 ;
  assign n39921 = n8662 & ~n39920 ;
  assign n39922 = n1204 & n23273 ;
  assign n39923 = n16633 ^ n14823 ^ 1'b0 ;
  assign n39924 = n21678 ^ n16998 ^ 1'b0 ;
  assign n39925 = n39923 | n39924 ;
  assign n39926 = n34852 & ~n39925 ;
  assign n39927 = n13228 & n39926 ;
  assign n39928 = n17081 ^ n654 ^ 1'b0 ;
  assign n39929 = n39928 ^ n24164 ^ n15283 ;
  assign n39930 = n16597 | n35077 ;
  assign n39931 = n14385 ^ n8774 ^ 1'b0 ;
  assign n39932 = n39399 | n39931 ;
  assign n39933 = n11820 ^ n11142 ^ 1'b0 ;
  assign n39934 = n428 & n1289 ;
  assign n39935 = ~n428 & n39934 ;
  assign n39936 = n445 | n1966 ;
  assign n39937 = n39935 & ~n39936 ;
  assign n39938 = n39933 | n39937 ;
  assign n39939 = n39933 & ~n39938 ;
  assign n39940 = n24986 | n39939 ;
  assign n39941 = n27878 ^ n2016 ^ 1'b0 ;
  assign n39942 = n39940 & n39941 ;
  assign n39943 = n28513 ^ n24518 ^ 1'b0 ;
  assign n39944 = ~n3579 & n39943 ;
  assign n39945 = n39944 ^ n10769 ^ n318 ;
  assign n39946 = n39945 ^ n7294 ^ 1'b0 ;
  assign n39947 = n21385 & ~n39061 ;
  assign n39948 = n38803 ^ n3166 ^ 1'b0 ;
  assign n39949 = n4044 & ~n21320 ;
  assign n39950 = n39948 & ~n39949 ;
  assign n39951 = n10114 & n25646 ;
  assign n39952 = n39951 ^ n15138 ^ n11680 ;
  assign n39953 = n3366 | n8266 ;
  assign n39954 = n32367 | n39953 ;
  assign n39955 = n39954 ^ n7360 ^ 1'b0 ;
  assign n39956 = n6271 | n39955 ;
  assign n39957 = ~n20002 & n39921 ;
  assign n39958 = n39957 ^ n9701 ^ 1'b0 ;
  assign n39959 = n14998 & n21411 ;
  assign n39960 = n620 & n36979 ;
  assign n39961 = n7655 | n23067 ;
  assign n39962 = n249 | n26787 ;
  assign n39963 = ~n20317 & n25882 ;
  assign n39964 = n39963 ^ n32768 ^ 1'b0 ;
  assign n39965 = n15754 ^ n11906 ^ 1'b0 ;
  assign n39966 = ~n10231 & n39965 ;
  assign n39967 = n33397 ^ n12284 ^ 1'b0 ;
  assign n39968 = n19466 | n39967 ;
  assign n39969 = n25619 & ~n39968 ;
  assign n39970 = n4241 | n13821 ;
  assign n39971 = ( n6195 & n12884 ) | ( n6195 & ~n13687 ) | ( n12884 & ~n13687 ) ;
  assign n39972 = n39971 ^ n30861 ^ 1'b0 ;
  assign n39973 = ~n39970 & n39972 ;
  assign n39974 = ~n5992 & n27881 ;
  assign n39975 = n39974 ^ n5517 ^ 1'b0 ;
  assign n39976 = n35997 ^ n7087 ^ 1'b0 ;
  assign n39977 = n15719 & n20621 ;
  assign n39978 = ~n34075 & n39977 ;
  assign n39979 = n2986 & n36418 ;
  assign n39980 = n10900 & n39979 ;
  assign n39981 = n1235 | n22581 ;
  assign n39982 = n6408 & ~n39981 ;
  assign n39983 = n23383 | n39982 ;
  assign n39984 = ( n14226 & ~n20010 ) | ( n14226 & n30185 ) | ( ~n20010 & n30185 ) ;
  assign n39985 = n39984 ^ n4139 ^ 1'b0 ;
  assign n39986 = n6196 | n39985 ;
  assign n39987 = n23133 ^ n3700 ^ 1'b0 ;
  assign n39988 = n33828 & n39987 ;
  assign n39989 = ~n19622 & n39988 ;
  assign n39990 = n3096 | n5839 ;
  assign n39991 = n14349 | n16790 ;
  assign n39992 = n33701 & n39991 ;
  assign n39993 = n14948 & ~n25919 ;
  assign n39994 = n14198 & n31442 ;
  assign n39995 = n39994 ^ n7358 ^ 1'b0 ;
  assign n39996 = n36946 ^ n25917 ^ 1'b0 ;
  assign n39997 = n31357 ^ n12587 ^ 1'b0 ;
  assign n39998 = n3934 | n39997 ;
  assign n39999 = n39998 ^ n14164 ^ 1'b0 ;
  assign n40000 = n11701 ^ n7941 ^ 1'b0 ;
  assign n40001 = n25234 | n40000 ;
  assign n40002 = n14039 ^ n13285 ^ 1'b0 ;
  assign n40003 = n14235 | n40002 ;
  assign n40004 = n11759 & n38639 ;
  assign n40005 = n6893 & n40004 ;
  assign n40006 = ( n19617 & ~n40003 ) | ( n19617 & n40005 ) | ( ~n40003 & n40005 ) ;
  assign n40007 = n2349 & n29443 ;
  assign n40008 = n40007 ^ n11688 ^ 1'b0 ;
  assign n40009 = ~n2806 & n22143 ;
  assign n40010 = n10150 ^ n74 ^ 1'b0 ;
  assign n40011 = n37307 ^ n14555 ^ 1'b0 ;
  assign n40012 = n14330 ^ n14112 ^ 1'b0 ;
  assign n40013 = n24188 | n40012 ;
  assign n40014 = n2572 & n8340 ;
  assign n40015 = n40014 ^ n34586 ^ 1'b0 ;
  assign n40016 = ~n1031 & n1548 ;
  assign n40017 = n40015 & n40016 ;
  assign n40018 = n39488 ^ n2708 ^ 1'b0 ;
  assign n40019 = n19446 ^ n12715 ^ 1'b0 ;
  assign n40020 = n26095 & ~n40019 ;
  assign n40021 = ~n19163 & n40020 ;
  assign n40022 = n13612 & n28274 ;
  assign n40023 = n17123 ^ n8712 ^ 1'b0 ;
  assign n40024 = ~n2491 & n16028 ;
  assign n40025 = n5825 | n20177 ;
  assign n40026 = n4478 & ~n16047 ;
  assign n40027 = ~n33648 & n40026 ;
  assign n40028 = n40027 ^ n27779 ^ 1'b0 ;
  assign n40029 = n31549 ^ n10389 ^ 1'b0 ;
  assign n40030 = n15130 ^ n9931 ^ n9704 ;
  assign n40031 = ( n26711 & ~n40029 ) | ( n26711 & n40030 ) | ( ~n40029 & n40030 ) ;
  assign n40032 = n1615 | n26958 ;
  assign n40033 = n13304 ^ n9704 ^ 1'b0 ;
  assign n40034 = ~n881 & n40033 ;
  assign n40035 = n21967 ^ n21337 ^ 1'b0 ;
  assign n40036 = n9901 & ~n27516 ;
  assign n40037 = n8939 & n40036 ;
  assign n40038 = n8862 ^ n3454 ^ 1'b0 ;
  assign n40039 = n1567 | n5154 ;
  assign n40040 = n835 & ~n40039 ;
  assign n40041 = n2143 ^ n1703 ^ 1'b0 ;
  assign n40042 = n890 & n11932 ;
  assign n40043 = ( n40040 & n40041 ) | ( n40040 & ~n40042 ) | ( n40041 & ~n40042 ) ;
  assign n40044 = n13712 & n20313 ;
  assign n40045 = ~n14388 & n40044 ;
  assign n40046 = n40045 ^ n39067 ^ n8225 ;
  assign n40047 = n16473 | n32384 ;
  assign n40048 = n32857 & ~n40047 ;
  assign n40049 = n30085 ^ n21916 ^ n14785 ;
  assign n40050 = n21325 ^ n3039 ^ 1'b0 ;
  assign n40051 = n5217 | n40050 ;
  assign n40052 = n15509 & ~n40051 ;
  assign n40053 = ~n40049 & n40052 ;
  assign n40054 = n19728 | n40053 ;
  assign n40055 = n17852 ^ n17409 ^ 1'b0 ;
  assign n40056 = n7405 & ~n40055 ;
  assign n40057 = n11781 ^ n2763 ^ 1'b0 ;
  assign n40058 = ~n4583 & n33958 ;
  assign n40059 = n788 & n22017 ;
  assign n40060 = n5333 & n40059 ;
  assign n40061 = n40060 ^ n20406 ^ n16756 ;
  assign n40062 = ~n25191 & n27995 ;
  assign n40063 = ~n1435 & n40062 ;
  assign n40064 = n14827 ^ n10119 ^ 1'b0 ;
  assign n40065 = n40064 ^ n8282 ^ 1'b0 ;
  assign n40066 = ~n32702 & n40065 ;
  assign n40067 = ~n9553 & n40066 ;
  assign n40069 = n466 ^ n367 ^ 1'b0 ;
  assign n40070 = n40069 ^ n3760 ^ 1'b0 ;
  assign n40068 = n12588 & ~n22630 ;
  assign n40071 = n40070 ^ n40068 ^ 1'b0 ;
  assign n40072 = n11682 | n12625 ;
  assign n40073 = n2292 & ~n5866 ;
  assign n40074 = n6271 & n40073 ;
  assign n40075 = n33554 & ~n40074 ;
  assign n40076 = ~n12264 & n40075 ;
  assign n40077 = n40076 ^ n16795 ^ 1'b0 ;
  assign n40078 = n12390 ^ n9846 ^ n3579 ;
  assign n40079 = ~n30534 & n40078 ;
  assign n40080 = n40077 | n40079 ;
  assign n40081 = ~n27540 & n40080 ;
  assign n40082 = ~n13385 & n13934 ;
  assign n40083 = n582 & n40082 ;
  assign n40084 = n40083 ^ n8190 ^ 1'b0 ;
  assign n40085 = x11 & ~n19967 ;
  assign n40086 = n40085 ^ n25955 ^ 1'b0 ;
  assign n40087 = n35316 ^ n15196 ^ n9356 ;
  assign n40089 = n2588 & ~n14559 ;
  assign n40088 = n6809 & ~n13192 ;
  assign n40090 = n40089 ^ n40088 ^ n21461 ;
  assign n40091 = n40090 ^ n4837 ^ 1'b0 ;
  assign n40093 = n29929 ^ n9270 ^ 1'b0 ;
  assign n40094 = ~n25336 & n40093 ;
  assign n40092 = n9404 & ~n14236 ;
  assign n40095 = n40094 ^ n40092 ^ 1'b0 ;
  assign n40096 = n33806 & ~n40095 ;
  assign n40097 = ~n11759 & n40096 ;
  assign n40098 = n25254 ^ n20492 ^ 1'b0 ;
  assign n40099 = n18062 | n40098 ;
  assign n40101 = n9922 ^ n9290 ^ 1'b0 ;
  assign n40100 = ( n6722 & n10175 ) | ( n6722 & ~n32618 ) | ( n10175 & ~n32618 ) ;
  assign n40102 = n40101 ^ n40100 ^ n30069 ;
  assign n40103 = n11525 & ~n22929 ;
  assign n40104 = n10484 | n14034 ;
  assign n40105 = n40104 ^ n18510 ^ 1'b0 ;
  assign n40106 = n11296 | n40105 ;
  assign n40107 = ~n8016 & n40106 ;
  assign n40108 = n14235 ^ n9746 ^ 1'b0 ;
  assign n40109 = ~n17511 & n40108 ;
  assign n40110 = n25017 ^ n2377 ^ 1'b0 ;
  assign n40111 = n30701 | n40110 ;
  assign n40112 = n39395 ^ n36876 ^ 1'b0 ;
  assign n40113 = n10167 & ~n40112 ;
  assign n40114 = n13594 & n27174 ;
  assign n40115 = n11470 & ~n15531 ;
  assign n40116 = n40115 ^ n2202 ^ 1'b0 ;
  assign n40117 = n13010 | n13980 ;
  assign n40118 = n17054 ^ n8584 ^ n6447 ;
  assign n40119 = n40118 ^ n4856 ^ 1'b0 ;
  assign n40120 = ~n6849 & n10456 ;
  assign n40121 = n40120 ^ n3539 ^ 1'b0 ;
  assign n40122 = ~n2039 & n40121 ;
  assign n40123 = n40122 ^ n6997 ^ 1'b0 ;
  assign n40124 = n40119 & n40123 ;
  assign n40125 = n6081 ^ n3442 ^ 1'b0 ;
  assign n40126 = n40125 ^ n27017 ^ n3270 ;
  assign n40127 = n14682 & n18060 ;
  assign n40128 = ( n17439 & n37914 ) | ( n17439 & n40127 ) | ( n37914 & n40127 ) ;
  assign n40129 = n4499 | n33219 ;
  assign n40130 = n40129 ^ n9453 ^ 1'b0 ;
  assign n40131 = n296 & ~n2791 ;
  assign n40132 = ~n12404 & n40131 ;
  assign n40133 = n10472 ^ n461 ^ 1'b0 ;
  assign n40134 = n35342 ^ n14804 ^ 1'b0 ;
  assign n40135 = n40133 | n40134 ;
  assign n40136 = n4537 & ~n31493 ;
  assign n40137 = n1542 & ~n12116 ;
  assign n40138 = ~n16335 & n40137 ;
  assign n40139 = ( ~n9264 & n11527 ) | ( ~n9264 & n40138 ) | ( n11527 & n40138 ) ;
  assign n40140 = n31301 | n37714 ;
  assign n40141 = n20721 ^ n3504 ^ 1'b0 ;
  assign n40142 = n3484 & n40141 ;
  assign n40143 = n2691 & ~n24009 ;
  assign n40144 = n3838 & n27174 ;
  assign n40145 = n40144 ^ n16241 ^ 1'b0 ;
  assign n40146 = ( ~n738 & n15897 ) | ( ~n738 & n24666 ) | ( n15897 & n24666 ) ;
  assign n40147 = ( n4512 & n27814 ) | ( n4512 & ~n40146 ) | ( n27814 & ~n40146 ) ;
  assign n40148 = ( n7631 & n23570 ) | ( n7631 & n29871 ) | ( n23570 & n29871 ) ;
  assign n40149 = ( n11664 & n16103 ) | ( n11664 & ~n40148 ) | ( n16103 & ~n40148 ) ;
  assign n40150 = n30853 & n34217 ;
  assign n40151 = n7042 | n8229 ;
  assign n40152 = n21170 & ~n31180 ;
  assign n40153 = n1351 & n34327 ;
  assign n40154 = n40153 ^ n23854 ^ 1'b0 ;
  assign n40156 = n14559 ^ n11020 ^ n7814 ;
  assign n40155 = n37527 ^ n34983 ^ n19418 ;
  assign n40157 = n40156 ^ n40155 ^ n30914 ;
  assign n40158 = n35082 ^ n27454 ^ n15680 ;
  assign n40159 = n8811 | n16062 ;
  assign n40160 = n40159 ^ n5566 ^ 1'b0 ;
  assign n40161 = n2038 & ~n40160 ;
  assign n40162 = n30187 ^ n8457 ^ 1'b0 ;
  assign n40163 = n1441 ^ n571 ^ 1'b0 ;
  assign n40164 = n28355 ^ n1269 ^ 1'b0 ;
  assign n40165 = ~n1794 & n37891 ;
  assign n40166 = ~n18664 & n40165 ;
  assign n40167 = n6037 & n11934 ;
  assign n40168 = n40166 & n40167 ;
  assign n40169 = n1075 & n40168 ;
  assign n40170 = n15515 & n17314 ;
  assign n40171 = n40170 ^ n1980 ^ 1'b0 ;
  assign n40172 = ~n3831 & n20518 ;
  assign n40173 = n39873 ^ n36634 ^ 1'b0 ;
  assign n40174 = ~n7004 & n22676 ;
  assign n40175 = n40174 ^ n9124 ^ 1'b0 ;
  assign n40176 = n17074 & n40175 ;
  assign n40177 = ~n35516 & n40176 ;
  assign n40178 = n21715 | n40177 ;
  assign n40179 = n11020 ^ n9969 ^ 1'b0 ;
  assign n40180 = n15273 & ~n40179 ;
  assign n40181 = n40180 ^ n24496 ^ 1'b0 ;
  assign n40182 = n5319 ^ n1566 ^ 1'b0 ;
  assign n40183 = n40182 ^ n25802 ^ n20315 ;
  assign n40184 = n9611 ^ n5276 ^ 1'b0 ;
  assign n40185 = n26301 & ~n40184 ;
  assign n40186 = n18402 & n34124 ;
  assign n40187 = ~n9953 & n40186 ;
  assign n40188 = n28413 & n40187 ;
  assign n40189 = n3781 & n40188 ;
  assign n40190 = n19690 ^ n3730 ^ 1'b0 ;
  assign n40191 = n9468 | n40190 ;
  assign n40192 = n22541 ^ n7340 ^ 1'b0 ;
  assign n40193 = ( n1915 & n9289 ) | ( n1915 & ~n15000 ) | ( n9289 & ~n15000 ) ;
  assign n40194 = n22923 ^ n8803 ^ 1'b0 ;
  assign n40195 = n21201 ^ n1603 ^ 1'b0 ;
  assign n40196 = ~n25793 & n40195 ;
  assign n40197 = n40009 ^ n12773 ^ 1'b0 ;
  assign n40198 = n21434 | n40197 ;
  assign n40199 = ( n22022 & ~n28481 ) | ( n22022 & n33316 ) | ( ~n28481 & n33316 ) ;
  assign n40200 = n40199 ^ n23738 ^ 1'b0 ;
  assign n40201 = n1657 | n9803 ;
  assign n40202 = n3231 & ~n40201 ;
  assign n40203 = n40202 ^ n24897 ^ 1'b0 ;
  assign n40204 = n3212 | n29017 ;
  assign n40205 = n659 | n39457 ;
  assign n40206 = n19842 & ~n36387 ;
  assign n40207 = n38498 & n40206 ;
  assign n40208 = n6702 | n12470 ;
  assign n40209 = ~n8136 & n40208 ;
  assign n40210 = n12405 | n40209 ;
  assign n40211 = n15546 ^ n14961 ^ 1'b0 ;
  assign n40212 = n4301 | n5749 ;
  assign n40213 = n23040 & ~n40212 ;
  assign n40214 = n40213 ^ n481 ^ 1'b0 ;
  assign n40215 = n37625 ^ n24179 ^ n11512 ;
  assign n40216 = n21223 & n40215 ;
  assign n40217 = n40216 ^ n33632 ^ 1'b0 ;
  assign n40218 = n2941 & ~n29214 ;
  assign n40219 = ~n24597 & n32468 ;
  assign n40220 = n5395 & ~n27858 ;
  assign n40225 = n18375 ^ n8926 ^ 1'b0 ;
  assign n40221 = n2840 & ~n8750 ;
  assign n40222 = ~n11086 & n40221 ;
  assign n40223 = n1072 & n40222 ;
  assign n40224 = n18723 & ~n40223 ;
  assign n40226 = n40225 ^ n40224 ^ 1'b0 ;
  assign n40227 = n40190 ^ n14385 ^ 1'b0 ;
  assign n40228 = n27369 ^ n14192 ^ 1'b0 ;
  assign n40229 = n40227 | n40228 ;
  assign n40230 = n9518 ^ n4754 ^ n3636 ;
  assign n40231 = n12929 & n40230 ;
  assign n40232 = ~n11524 & n14059 ;
  assign n40233 = n40232 ^ n4074 ^ 1'b0 ;
  assign n40234 = n9226 | n14537 ;
  assign n40235 = n19473 & ~n40234 ;
  assign n40236 = n40235 ^ n23020 ^ 1'b0 ;
  assign n40237 = n9825 | n40236 ;
  assign n40238 = n6753 & n7806 ;
  assign n40239 = n20045 ^ n16774 ^ 1'b0 ;
  assign n40240 = n4242 & ~n16358 ;
  assign n40241 = ~n4944 & n38395 ;
  assign n40242 = n3049 & n16536 ;
  assign n40243 = ~n8302 & n40242 ;
  assign n40244 = n40243 ^ n16394 ^ 1'b0 ;
  assign n40245 = n29255 | n40244 ;
  assign n40246 = n3312 | n40245 ;
  assign n40247 = n15787 | n24230 ;
  assign n40248 = ~n9102 & n11505 ;
  assign n40249 = n40248 ^ n13994 ^ 1'b0 ;
  assign n40250 = ~n9253 & n40123 ;
  assign n40252 = n2085 ^ n612 ^ 1'b0 ;
  assign n40251 = n1045 & ~n33299 ;
  assign n40253 = n40252 ^ n40251 ^ 1'b0 ;
  assign n40254 = ~n24931 & n40253 ;
  assign n40256 = ~n7961 & n17584 ;
  assign n40257 = n22986 & n40256 ;
  assign n40255 = n4984 & ~n19881 ;
  assign n40258 = n40257 ^ n40255 ^ 1'b0 ;
  assign n40259 = ( ~n582 & n5237 ) | ( ~n582 & n5646 ) | ( n5237 & n5646 ) ;
  assign n40260 = n40259 ^ n38639 ^ 1'b0 ;
  assign n40261 = ~n38260 & n40260 ;
  assign n40262 = n24115 ^ n16462 ^ 1'b0 ;
  assign n40263 = n10418 & n40262 ;
  assign n40264 = n40263 ^ n2287 ^ 1'b0 ;
  assign n40265 = n27729 & ~n40264 ;
  assign n40266 = n6376 & n13915 ;
  assign n40267 = n40266 ^ n14164 ^ 1'b0 ;
  assign n40268 = n25643 ^ n19941 ^ n7798 ;
  assign n40269 = n16147 ^ n13101 ^ 1'b0 ;
  assign n40270 = ( ~n2352 & n7149 ) | ( ~n2352 & n40269 ) | ( n7149 & n40269 ) ;
  assign n40271 = n25163 ^ n9700 ^ 1'b0 ;
  assign n40272 = n40270 & n40271 ;
  assign n40273 = n2571 & ~n25544 ;
  assign n40274 = n34460 & n40273 ;
  assign n40275 = n11073 & n11765 ;
  assign n40276 = ~n6164 & n40275 ;
  assign n40277 = ( n7360 & n40257 ) | ( n7360 & ~n40276 ) | ( n40257 & ~n40276 ) ;
  assign n40278 = n16941 ^ n3699 ^ 1'b0 ;
  assign n40279 = n11632 & n40278 ;
  assign n40280 = n40279 ^ n39875 ^ n5697 ;
  assign n40281 = ~n28421 & n39626 ;
  assign n40282 = n6016 & ~n21593 ;
  assign n40283 = n40282 ^ n19336 ^ 1'b0 ;
  assign n40284 = n25597 ^ n17739 ^ 1'b0 ;
  assign n40285 = ~n8715 & n40284 ;
  assign n40286 = ~n16275 & n27888 ;
  assign n40287 = n40286 ^ n22174 ^ 1'b0 ;
  assign n40288 = n40285 & ~n40287 ;
  assign n40289 = n20527 ^ n3616 ^ 1'b0 ;
  assign n40290 = ~n24038 & n29910 ;
  assign n40291 = ( n2080 & ~n8323 ) | ( n2080 & n15822 ) | ( ~n8323 & n15822 ) ;
  assign n40292 = n11994 ^ n5531 ^ 1'b0 ;
  assign n40293 = ~n5388 & n35869 ;
  assign n40294 = n40293 ^ n2596 ^ 1'b0 ;
  assign n40295 = n40292 | n40294 ;
  assign n40296 = n40291 & ~n40295 ;
  assign n40297 = n32639 ^ n425 ^ 1'b0 ;
  assign n40298 = n25580 ^ n11153 ^ 1'b0 ;
  assign n40299 = n387 | n40298 ;
  assign n40300 = n1331 | n24632 ;
  assign n40301 = n24336 ^ n20862 ^ 1'b0 ;
  assign n40302 = n12109 & ~n40301 ;
  assign n40303 = ~n2781 & n8370 ;
  assign n40304 = n3214 & n40303 ;
  assign n40305 = n3558 | n40304 ;
  assign n40306 = n13275 | n40305 ;
  assign n40307 = n14500 & n23230 ;
  assign n40308 = ~n15631 & n40307 ;
  assign n40309 = n17572 & n24541 ;
  assign n40310 = n40309 ^ n625 ^ 1'b0 ;
  assign n40311 = n229 | n20405 ;
  assign n40312 = n40311 ^ n15651 ^ 1'b0 ;
  assign n40313 = ~n19240 & n40312 ;
  assign n40314 = n24838 & n40313 ;
  assign n40315 = ~n20455 & n36525 ;
  assign n40316 = ~n1961 & n40315 ;
  assign n40317 = n22779 | n33708 ;
  assign n40318 = n34400 ^ n2401 ^ 1'b0 ;
  assign n40319 = ~n16028 & n31777 ;
  assign n40320 = ~n6941 & n10197 ;
  assign n40321 = n40320 ^ n25384 ^ 1'b0 ;
  assign n40322 = n35186 ^ n69 ^ 1'b0 ;
  assign n40323 = n3802 & ~n5783 ;
  assign n40325 = n12644 ^ n108 ^ 1'b0 ;
  assign n40324 = n15605 & n20628 ;
  assign n40326 = n40325 ^ n40324 ^ 1'b0 ;
  assign n40327 = ~n712 & n4829 ;
  assign n40328 = n40326 | n40327 ;
  assign n40329 = n9208 & ~n40328 ;
  assign n40330 = n23707 & n40329 ;
  assign n40331 = n29475 ^ n23637 ^ 1'b0 ;
  assign n40332 = n26288 ^ n9049 ^ 1'b0 ;
  assign n40333 = n25826 ^ n16292 ^ 1'b0 ;
  assign n40334 = ~n17893 & n31315 ;
  assign n40335 = ~n40333 & n40334 ;
  assign n40336 = n10048 ^ n5994 ^ 1'b0 ;
  assign n40337 = ~n40018 & n40336 ;
  assign n40338 = n17128 & ~n36650 ;
  assign n40340 = n4780 & n17849 ;
  assign n40341 = n1724 & n40340 ;
  assign n40339 = n12042 | n24196 ;
  assign n40342 = n40341 ^ n40339 ^ 1'b0 ;
  assign n40343 = n3383 | n30402 ;
  assign n40344 = n10601 & n40343 ;
  assign n40345 = n10196 & n40344 ;
  assign n40346 = n40345 ^ n5161 ^ 1'b0 ;
  assign n40347 = n10603 & n17072 ;
  assign n40349 = n9715 ^ n6827 ^ 1'b0 ;
  assign n40348 = ~n4493 & n28323 ;
  assign n40350 = n40349 ^ n40348 ^ 1'b0 ;
  assign n40351 = ~n6299 & n40350 ;
  assign n40352 = ~n40347 & n40351 ;
  assign n40354 = n10245 & ~n21213 ;
  assign n40355 = ( n1211 & ~n10875 ) | ( n1211 & n40354 ) | ( ~n10875 & n40354 ) ;
  assign n40353 = ~n4025 & n19759 ;
  assign n40356 = n40355 ^ n40353 ^ 1'b0 ;
  assign n40357 = n2885 ^ n1234 ^ 1'b0 ;
  assign n40358 = n4545 | n40357 ;
  assign n40359 = n4823 | n40358 ;
  assign n40360 = n11371 ^ n325 ^ 1'b0 ;
  assign n40361 = ~n13207 & n40360 ;
  assign n40362 = n5158 & n23433 ;
  assign n40363 = n8604 | n16647 ;
  assign n40364 = n40363 ^ n14123 ^ 1'b0 ;
  assign n40365 = n40364 ^ n37422 ^ 1'b0 ;
  assign n40366 = n20165 & n40365 ;
  assign n40368 = n5182 | n34807 ;
  assign n40367 = n3768 | n22501 ;
  assign n40369 = n40368 ^ n40367 ^ 1'b0 ;
  assign n40370 = n39422 ^ n26922 ^ 1'b0 ;
  assign n40371 = n2343 & ~n35107 ;
  assign n40372 = ~n40370 & n40371 ;
  assign n40373 = ~n6015 & n6216 ;
  assign n40374 = n8406 & ~n40373 ;
  assign n40375 = ~n3090 & n3628 ;
  assign n40376 = n2012 | n40375 ;
  assign n40377 = n40376 ^ n34717 ^ 1'b0 ;
  assign n40378 = n40377 ^ n20472 ^ 1'b0 ;
  assign n40379 = n5992 & n40378 ;
  assign n40380 = n24701 & ~n39003 ;
  assign n40381 = ~n5731 & n40380 ;
  assign n40382 = n3335 & n40381 ;
  assign n40383 = n40382 ^ n38768 ^ n24642 ;
  assign n40384 = n376 & ~n2476 ;
  assign n40385 = ~n376 & n40384 ;
  assign n40386 = ( n29451 & n30256 ) | ( n29451 & ~n40385 ) | ( n30256 & ~n40385 ) ;
  assign n40387 = ( n15588 & n21326 ) | ( n15588 & ~n27454 ) | ( n21326 & ~n27454 ) ;
  assign n40388 = ( n5333 & ~n40386 ) | ( n5333 & n40387 ) | ( ~n40386 & n40387 ) ;
  assign n40389 = n1178 & n21457 ;
  assign n40390 = n5836 & n40389 ;
  assign n40391 = n2876 & ~n19186 ;
  assign n40392 = n10378 & n40391 ;
  assign n40393 = n6114 | n16889 ;
  assign n40394 = n746 | n40393 ;
  assign n40395 = n13186 & n30648 ;
  assign n40396 = n1867 ^ n1853 ^ 1'b0 ;
  assign n40397 = ~n2673 & n6272 ;
  assign n40398 = n40397 ^ n23569 ^ 1'b0 ;
  assign n40399 = n6663 | n11743 ;
  assign n40400 = n6766 & ~n40399 ;
  assign n40401 = n10565 | n33507 ;
  assign n40402 = ~n40400 & n40401 ;
  assign n40403 = ~n3547 & n9848 ;
  assign n40404 = n40403 ^ n26794 ^ 1'b0 ;
  assign n40405 = n39319 ^ n38674 ^ 1'b0 ;
  assign n40406 = n5321 | n5704 ;
  assign n40407 = n5584 & ~n40406 ;
  assign n40408 = ( ~n1994 & n25643 ) | ( ~n1994 & n40407 ) | ( n25643 & n40407 ) ;
  assign n40409 = n12125 ^ n528 ^ 1'b0 ;
  assign n40410 = n33554 ^ n19458 ^ 1'b0 ;
  assign n40411 = n12747 & n33187 ;
  assign n40412 = n12646 & ~n28237 ;
  assign n40413 = ~n31565 & n40412 ;
  assign n40414 = n20042 ^ n443 ^ 1'b0 ;
  assign n40415 = n1513 & ~n7940 ;
  assign n40416 = n40415 ^ n991 ^ 1'b0 ;
  assign n40417 = n25616 ^ n4066 ^ 1'b0 ;
  assign n40418 = n40416 & ~n40417 ;
  assign n40419 = ( n33365 & n37622 ) | ( n33365 & n40418 ) | ( n37622 & n40418 ) ;
  assign n40420 = n7067 ^ n3240 ^ 1'b0 ;
  assign n40421 = n8681 | n40420 ;
  assign n40422 = ~n3992 & n32069 ;
  assign n40423 = n40422 ^ n29512 ^ 1'b0 ;
  assign n40424 = n3349 | n39663 ;
  assign n40425 = n6265 ^ n4163 ^ 1'b0 ;
  assign n40426 = n4757 & n24926 ;
  assign n40427 = n40425 & n40426 ;
  assign n40428 = n872 ^ n88 ^ 1'b0 ;
  assign n40429 = n1044 | n40428 ;
  assign n40430 = n31495 | n34014 ;
  assign n40431 = n40429 & ~n40430 ;
  assign n40432 = ~n7374 & n38491 ;
  assign n40433 = n15023 & n40432 ;
  assign n40434 = n40433 ^ n23778 ^ 1'b0 ;
  assign n40435 = ~n36290 & n40434 ;
  assign n40436 = n17142 & n40435 ;
  assign n40437 = n21606 | n34064 ;
  assign n40439 = n3917 | n24768 ;
  assign n40438 = n515 & ~n13165 ;
  assign n40440 = n40439 ^ n40438 ^ 1'b0 ;
  assign n40441 = n22071 ^ n6599 ^ 1'b0 ;
  assign n40442 = ~n25340 & n40441 ;
  assign n40443 = n40442 ^ n139 ^ 1'b0 ;
  assign n40444 = n3430 | n40443 ;
  assign n40445 = n7528 & ~n40444 ;
  assign n40446 = n40445 ^ n27740 ^ 1'b0 ;
  assign n40447 = n15206 & n40446 ;
  assign n40448 = ( n18363 & ~n31197 ) | ( n18363 & n40447 ) | ( ~n31197 & n40447 ) ;
  assign n40449 = n1685 & ~n9701 ;
  assign n40450 = n29697 ^ n77 ^ 1'b0 ;
  assign n40451 = n40449 & n40450 ;
  assign n40452 = n4930 & n12078 ;
  assign n40453 = n40452 ^ n37770 ^ 1'b0 ;
  assign n40454 = n3763 & n4077 ;
  assign n40455 = n31370 & n40454 ;
  assign n40456 = n5897 & n40455 ;
  assign n40457 = n10048 & ~n40456 ;
  assign n40458 = n33436 ^ n12773 ^ 1'b0 ;
  assign n40459 = n25708 ^ n13352 ^ 1'b0 ;
  assign n40460 = n32181 ^ n17345 ^ n5492 ;
  assign n40461 = n8390 ^ n3522 ^ 1'b0 ;
  assign n40462 = n40461 ^ n12528 ^ 1'b0 ;
  assign n40463 = n35559 & ~n40462 ;
  assign n40464 = ~n5900 & n40463 ;
  assign n40465 = n3738 & n24217 ;
  assign n40466 = n14312 | n24983 ;
  assign n40467 = n40466 ^ n18080 ^ 1'b0 ;
  assign n40468 = n318 & ~n40467 ;
  assign n40469 = n29707 ^ n15488 ^ n2645 ;
  assign n40470 = n16943 ^ n3145 ^ 1'b0 ;
  assign n40471 = n315 & ~n9837 ;
  assign n40472 = ~n27082 & n40471 ;
  assign n40473 = n37249 ^ n23547 ^ 1'b0 ;
  assign n40474 = n23751 ^ n8273 ^ 1'b0 ;
  assign n40475 = n10804 ^ n4843 ^ 1'b0 ;
  assign n40476 = n21791 & n40475 ;
  assign n40477 = n40476 ^ n11439 ^ n694 ;
  assign n40478 = ~n40474 & n40477 ;
  assign n40479 = n12271 ^ n7816 ^ 1'b0 ;
  assign n40480 = n24197 & n35196 ;
  assign n40481 = n40480 ^ n24041 ^ 1'b0 ;
  assign n40482 = n40479 & n40481 ;
  assign n40483 = n6282 & n26604 ;
  assign n40484 = n40483 ^ n16111 ^ 1'b0 ;
  assign n40485 = n38536 ^ n2140 ^ 1'b0 ;
  assign n40486 = n4910 ^ n2996 ^ 1'b0 ;
  assign n40487 = n2348 & n40486 ;
  assign n40488 = n40487 ^ n3426 ^ 1'b0 ;
  assign n40489 = n10782 ^ n387 ^ 1'b0 ;
  assign n40490 = n8054 ^ n1079 ^ 1'b0 ;
  assign n40491 = n11553 ^ n6314 ^ 1'b0 ;
  assign n40492 = n11353 | n40491 ;
  assign n40493 = n40492 ^ n24974 ^ 1'b0 ;
  assign n40494 = n21952 | n26075 ;
  assign n40495 = n10300 ^ n277 ^ 1'b0 ;
  assign n40496 = n32681 | n40495 ;
  assign n40497 = n40496 ^ n12525 ^ 1'b0 ;
  assign n40498 = n38973 | n40497 ;
  assign n40499 = n13794 ^ n3455 ^ 1'b0 ;
  assign n40500 = n5501 | n40499 ;
  assign n40501 = n40500 ^ n38452 ^ 1'b0 ;
  assign n40502 = n5758 & n40501 ;
  assign n40503 = n11741 ^ n4353 ^ 1'b0 ;
  assign n40504 = ~n4347 & n40503 ;
  assign n40505 = ~n40502 & n40504 ;
  assign n40506 = n27031 ^ n15429 ^ 1'b0 ;
  assign n40507 = ~n39867 & n40506 ;
  assign n40508 = n1414 & n4981 ;
  assign n40509 = n446 & ~n16493 ;
  assign n40510 = n5935 & n40509 ;
  assign n40511 = n20505 | n40510 ;
  assign n40512 = n2872 & ~n40511 ;
  assign n40513 = n32514 | n40512 ;
  assign n40514 = ~n5490 & n10592 ;
  assign n40515 = ( ~n2481 & n5529 ) | ( ~n2481 & n40514 ) | ( n5529 & n40514 ) ;
  assign n40516 = n40515 ^ n5742 ^ 1'b0 ;
  assign n40517 = n11242 ^ n322 ^ 1'b0 ;
  assign n40518 = ~n24671 & n40517 ;
  assign n40519 = n40518 ^ n28378 ^ 1'b0 ;
  assign n40520 = n33333 & ~n40519 ;
  assign n40521 = n4302 & n40520 ;
  assign n40522 = n16464 & n31051 ;
  assign n40523 = n140 & n40522 ;
  assign n40524 = n40523 ^ n29669 ^ 1'b0 ;
  assign n40525 = n315 & ~n26253 ;
  assign n40526 = n32301 ^ n3388 ^ 1'b0 ;
  assign n40527 = n28641 ^ n18158 ^ n4128 ;
  assign n40528 = n13147 ^ n4478 ^ n3726 ;
  assign n40529 = n2146 & n7877 ;
  assign n40530 = n9131 & n40529 ;
  assign n40531 = n23913 ^ n4119 ^ 1'b0 ;
  assign n40532 = n19840 | n40531 ;
  assign n40533 = n4732 | n40532 ;
  assign n40534 = n8663 | n40533 ;
  assign n40535 = n21344 ^ n2907 ^ 1'b0 ;
  assign n40536 = n17155 & n20573 ;
  assign n40537 = n40536 ^ n7008 ^ n1603 ;
  assign n40538 = ( n2203 & n3188 ) | ( n2203 & ~n4236 ) | ( n3188 & ~n4236 ) ;
  assign n40539 = n40538 ^ n2455 ^ 1'b0 ;
  assign n40540 = n575 | n4296 ;
  assign n40541 = n40540 ^ n8553 ^ 1'b0 ;
  assign n40542 = n25775 ^ n9279 ^ n6811 ;
  assign n40543 = n21982 ^ n7927 ^ 1'b0 ;
  assign n40544 = n40542 & n40543 ;
  assign n40545 = n7520 & n10128 ;
  assign n40546 = n22271 | n40545 ;
  assign n40547 = n40546 ^ n23855 ^ 1'b0 ;
  assign n40548 = n16203 | n30534 ;
  assign n40549 = n6995 | n40548 ;
  assign n40550 = n29961 & n40549 ;
  assign n40551 = n40550 ^ n15541 ^ 1'b0 ;
  assign n40552 = n14194 ^ n11182 ^ 1'b0 ;
  assign n40553 = ( n23283 & n23541 ) | ( n23283 & n40552 ) | ( n23541 & n40552 ) ;
  assign n40554 = ( n24478 & n28490 ) | ( n24478 & n40553 ) | ( n28490 & n40553 ) ;
  assign n40555 = n12606 ^ n3760 ^ 1'b0 ;
  assign n40556 = ~n7455 & n40555 ;
  assign n40557 = ~n466 & n40556 ;
  assign n40558 = n37213 ^ n4480 ^ 1'b0 ;
  assign n40559 = n4600 | n6599 ;
  assign n40560 = n7116 | n40559 ;
  assign n40561 = ~n6598 & n8477 ;
  assign n40562 = n40561 ^ n2914 ^ 1'b0 ;
  assign n40563 = n7271 | n9887 ;
  assign n40564 = n40563 ^ n23627 ^ n13373 ;
  assign n40565 = n2596 ^ n1093 ^ 1'b0 ;
  assign n40566 = n2859 & n32795 ;
  assign n40567 = n34258 & n40566 ;
  assign n40568 = n10281 & ~n40567 ;
  assign n40569 = n40565 & n40568 ;
  assign n40570 = n12485 ^ n135 ^ 1'b0 ;
  assign n40571 = n5093 | n40570 ;
  assign n40572 = n14525 & ~n40571 ;
  assign n40573 = n6216 ^ n3646 ^ 1'b0 ;
  assign n40574 = n9356 & n40573 ;
  assign n40578 = ~n2856 & n5067 ;
  assign n40576 = n29504 ^ n9311 ^ 1'b0 ;
  assign n40577 = n15128 | n40576 ;
  assign n40575 = n1845 ^ n58 ^ 1'b0 ;
  assign n40579 = n40578 ^ n40577 ^ n40575 ;
  assign n40580 = n9267 ^ n6184 ^ 1'b0 ;
  assign n40581 = n40579 | n40580 ;
  assign n40582 = n2164 & ~n14928 ;
  assign n40583 = n12049 & n28719 ;
  assign n40584 = n9193 ^ n6542 ^ n821 ;
  assign n40588 = ( n2816 & n3915 ) | ( n2816 & ~n18177 ) | ( n3915 & ~n18177 ) ;
  assign n40585 = n5360 & ~n5487 ;
  assign n40586 = n40585 ^ n39320 ^ 1'b0 ;
  assign n40587 = ~n420 & n40586 ;
  assign n40589 = n40588 ^ n40587 ^ 1'b0 ;
  assign n40590 = n40584 & ~n40589 ;
  assign n40591 = n27979 ^ n14092 ^ 1'b0 ;
  assign n40592 = ~n20159 & n40591 ;
  assign n40593 = n263 & n20558 ;
  assign n40594 = n40593 ^ n387 ^ 1'b0 ;
  assign n40595 = ~n712 & n25349 ;
  assign n40596 = ~n11876 & n40595 ;
  assign n40598 = n1843 | n18689 ;
  assign n40599 = n1843 & ~n40598 ;
  assign n40600 = n311 & ~n347 ;
  assign n40601 = n347 & n40600 ;
  assign n40602 = n40599 | n40601 ;
  assign n40603 = n40599 & ~n40602 ;
  assign n40604 = n1229 | n40603 ;
  assign n40605 = n40603 & ~n40604 ;
  assign n40606 = n12689 | n40605 ;
  assign n40607 = n40606 ^ n7652 ^ 1'b0 ;
  assign n40608 = n31206 | n40607 ;
  assign n40597 = ~n9823 & n26130 ;
  assign n40609 = n40608 ^ n40597 ^ 1'b0 ;
  assign n40611 = n2033 | n16164 ;
  assign n40610 = n7069 & ~n9515 ;
  assign n40612 = n40611 ^ n40610 ^ 1'b0 ;
  assign n40613 = n13321 ^ n8872 ^ n2455 ;
  assign n40614 = n13182 ^ n2086 ^ 1'b0 ;
  assign n40615 = n11794 & ~n40614 ;
  assign n40616 = n24800 ^ n6294 ^ 1'b0 ;
  assign n40617 = n3616 & ~n40616 ;
  assign n40618 = n40617 ^ n36670 ^ n21081 ;
  assign n40619 = n38287 | n40618 ;
  assign n40620 = n40619 ^ n8963 ^ 1'b0 ;
  assign n40621 = n3924 & ~n30593 ;
  assign n40622 = n1590 & n28435 ;
  assign n40623 = n21926 & n40622 ;
  assign n40624 = n15596 ^ n2481 ^ 1'b0 ;
  assign n40625 = n26744 ^ n2451 ^ 1'b0 ;
  assign n40626 = n6048 | n40625 ;
  assign n40627 = n40626 ^ n31957 ^ 1'b0 ;
  assign n40628 = n14244 ^ n6042 ^ 1'b0 ;
  assign n40629 = n12688 & ~n40628 ;
  assign n40630 = ~n37422 & n40629 ;
  assign n40631 = n16657 ^ n6063 ^ 1'b0 ;
  assign n40632 = n6865 | n40631 ;
  assign n40633 = n10657 | n12921 ;
  assign n40634 = n40632 & ~n40633 ;
  assign n40635 = n7059 & ~n40634 ;
  assign n40636 = n5028 & n40635 ;
  assign n40637 = ~n26348 & n40636 ;
  assign n40638 = ~n5511 & n20545 ;
  assign n40639 = n16042 & n40638 ;
  assign n40640 = n16615 ^ n2818 ^ 1'b0 ;
  assign n40641 = n34629 & ~n40640 ;
  assign n40642 = n22517 ^ n3748 ^ 1'b0 ;
  assign n40643 = n3397 | n9785 ;
  assign n40644 = n7804 | n11790 ;
  assign n40645 = n39554 ^ n30532 ^ 1'b0 ;
  assign n40646 = n5520 | n40645 ;
  assign n40647 = ( n31335 & ~n40644 ) | ( n31335 & n40646 ) | ( ~n40644 & n40646 ) ;
  assign n40648 = n19069 ^ n266 ^ 1'b0 ;
  assign n40649 = n20846 ^ n18879 ^ 1'b0 ;
  assign n40650 = n30432 & n40649 ;
  assign n40651 = n40650 ^ n4369 ^ 1'b0 ;
  assign n40652 = ~n32666 & n40651 ;
  assign n40653 = n20962 ^ n13247 ^ 1'b0 ;
  assign n40654 = n25209 & n40653 ;
  assign n40655 = n14959 ^ n1893 ^ 1'b0 ;
  assign n40656 = n7457 & ~n40655 ;
  assign n40657 = n28018 & n40656 ;
  assign n40658 = n39366 ^ n32539 ^ n13515 ;
  assign n40659 = ~n14452 & n24620 ;
  assign n40660 = n2971 & ~n26465 ;
  assign n40661 = n20571 & n40660 ;
  assign n40662 = n40661 ^ n4401 ^ 1'b0 ;
  assign n40663 = n8487 | n40662 ;
  assign n40664 = ( n382 & n2595 ) | ( n382 & ~n3194 ) | ( n2595 & ~n3194 ) ;
  assign n40665 = n24093 & n40664 ;
  assign n40666 = ~n24093 & n40665 ;
  assign n40674 = n21631 ^ n20268 ^ 1'b0 ;
  assign n40675 = n40674 ^ n3402 ^ 1'b0 ;
  assign n40667 = n737 & n1312 ;
  assign n40668 = ~n1312 & n40667 ;
  assign n40669 = n25504 & n40668 ;
  assign n40670 = n23770 ^ n8727 ^ 1'b0 ;
  assign n40671 = n5781 | n40670 ;
  assign n40672 = n40669 | n40671 ;
  assign n40673 = n40669 & ~n40672 ;
  assign n40676 = n40675 ^ n40673 ^ 1'b0 ;
  assign n40677 = n3828 & ~n40676 ;
  assign n40678 = n40666 & n40677 ;
  assign n40679 = n4044 | n24283 ;
  assign n40680 = n15641 & n17325 ;
  assign n40681 = ~n1755 & n5328 ;
  assign n40682 = n40681 ^ n13677 ^ 1'b0 ;
  assign n40683 = n9940 | n13010 ;
  assign n40684 = n40683 ^ n20458 ^ 1'b0 ;
  assign n40685 = n40684 ^ n38702 ^ n6993 ;
  assign n40686 = ~n40346 & n40685 ;
  assign n40687 = n40686 ^ n28701 ^ 1'b0 ;
  assign n40688 = ( n3877 & n29317 ) | ( n3877 & ~n29642 ) | ( n29317 & ~n29642 ) ;
  assign n40689 = n8513 & n9873 ;
  assign n40690 = n40689 ^ n7620 ^ 1'b0 ;
  assign n40691 = n4468 & n21201 ;
  assign n40692 = ~n9874 & n18939 ;
  assign n40693 = n3153 | n36670 ;
  assign n40694 = n24703 ^ n3708 ^ 1'b0 ;
  assign n40695 = n5952 & n14825 ;
  assign n40696 = n40695 ^ n29327 ^ 1'b0 ;
  assign n40697 = n18727 ^ n7614 ^ 1'b0 ;
  assign n40698 = n40696 & ~n40697 ;
  assign n40699 = n1928 | n5522 ;
  assign n40700 = n40699 ^ n1249 ^ 1'b0 ;
  assign n40701 = n40700 ^ n10211 ^ 1'b0 ;
  assign n40702 = ~n6436 & n40701 ;
  assign n40703 = n8534 & ~n40702 ;
  assign n40704 = n1071 & n2567 ;
  assign n40705 = n15111 & n40704 ;
  assign n40706 = n12599 ^ n9680 ^ 1'b0 ;
  assign n40707 = n23793 & ~n40706 ;
  assign n40708 = n11763 | n40707 ;
  assign n40709 = n25611 ^ n1083 ^ 1'b0 ;
  assign n40710 = n33982 & n40709 ;
  assign n40711 = n4074 & n11176 ;
  assign n40712 = n40711 ^ n8456 ^ 1'b0 ;
  assign n40713 = ( n2273 & ~n33109 ) | ( n2273 & n40712 ) | ( ~n33109 & n40712 ) ;
  assign n40714 = n36055 ^ n5306 ^ 1'b0 ;
  assign n40715 = n4007 & n40714 ;
  assign n40716 = ~n3242 & n40715 ;
  assign n40717 = n40716 ^ n12190 ^ 1'b0 ;
  assign n40718 = ( n12100 & n33980 ) | ( n12100 & n40717 ) | ( n33980 & n40717 ) ;
  assign n40720 = n17792 & ~n28181 ;
  assign n40719 = n10315 & n37609 ;
  assign n40721 = n40720 ^ n40719 ^ 1'b0 ;
  assign n40722 = n934 | n35053 ;
  assign n40723 = n5593 & ~n14184 ;
  assign n40724 = n23897 ^ n13062 ^ 1'b0 ;
  assign n40725 = n40724 ^ n8036 ^ 1'b0 ;
  assign n40726 = ~n19042 & n40725 ;
  assign n40727 = n21845 & n40726 ;
  assign n40728 = n40727 ^ n167 ^ 1'b0 ;
  assign n40729 = n2649 | n22873 ;
  assign n40730 = n8210 | n40729 ;
  assign n40733 = ~n3671 & n13267 ;
  assign n40734 = n13844 | n40733 ;
  assign n40731 = ~n12541 & n30741 ;
  assign n40732 = n7510 & n40731 ;
  assign n40735 = n40734 ^ n40732 ^ 1'b0 ;
  assign n40737 = n17644 & n23736 ;
  assign n40736 = n448 | n11016 ;
  assign n40738 = n40737 ^ n40736 ^ n19978 ;
  assign n40739 = n11153 ^ n2401 ^ 1'b0 ;
  assign n40740 = n38928 ^ n7891 ^ 1'b0 ;
  assign n40741 = n26759 & n40740 ;
  assign n40742 = n13456 & n40741 ;
  assign n40743 = n2403 ^ n453 ^ 1'b0 ;
  assign n40744 = n20946 & ~n27973 ;
  assign n40745 = ~n40743 & n40744 ;
  assign n40746 = n17535 | n40512 ;
  assign n40747 = n4522 ^ n4014 ^ 1'b0 ;
  assign n40748 = n18900 & n40747 ;
  assign n40749 = n13059 & ~n40748 ;
  assign n40750 = n5390 ^ n682 ^ 1'b0 ;
  assign n40751 = ~n24985 & n40750 ;
  assign n40752 = n40751 ^ n28211 ^ 1'b0 ;
  assign n40753 = ~n122 & n9248 ;
  assign n40754 = n40753 ^ n35745 ^ n4775 ;
  assign n40755 = n7570 | n40754 ;
  assign n40756 = n15697 & ~n40755 ;
  assign n40757 = n16935 & ~n26038 ;
  assign n40758 = n2723 & n40757 ;
  assign n40759 = n32125 ^ n8411 ^ 1'b0 ;
  assign n40760 = ~n3687 & n40759 ;
  assign n40761 = n18960 | n40760 ;
  assign n40762 = n2315 & ~n6006 ;
  assign n40763 = n40762 ^ n695 ^ 1'b0 ;
  assign n40764 = n100 | n25267 ;
  assign n40765 = n10962 ^ n461 ^ 1'b0 ;
  assign n40766 = ~n40764 & n40765 ;
  assign n40767 = n28643 ^ n18252 ^ 1'b0 ;
  assign n40768 = ~n2109 & n14750 ;
  assign n40769 = n40768 ^ n17361 ^ 1'b0 ;
  assign n40770 = n10500 ^ n9159 ^ 1'b0 ;
  assign n40771 = n7233 & n40770 ;
  assign n40772 = n8324 | n8410 ;
  assign n40773 = n14396 & ~n33123 ;
  assign n40774 = n8909 | n23039 ;
  assign n40775 = n30763 ^ n24041 ^ n15641 ;
  assign n40776 = ~n466 & n2032 ;
  assign n40777 = ~n8168 & n40776 ;
  assign n40778 = n6225 ^ n4894 ^ 1'b0 ;
  assign n40779 = n26913 & n40778 ;
  assign n40780 = n315 & ~n4254 ;
  assign n40781 = n40780 ^ n7130 ^ 1'b0 ;
  assign n40782 = n20260 | n40781 ;
  assign n40783 = n40782 ^ n26130 ^ 1'b0 ;
  assign n40784 = n5675 & n40783 ;
  assign n40785 = n1344 & n16554 ;
  assign n40786 = n40785 ^ n1469 ^ 1'b0 ;
  assign n40787 = ~n10124 & n21239 ;
  assign n40788 = n27383 & n40787 ;
  assign n40789 = n16408 & ~n18603 ;
  assign n40790 = n40788 & n40789 ;
  assign n40791 = n165 & ~n28837 ;
  assign n40792 = n20697 & n40791 ;
  assign n40793 = n1718 & ~n19004 ;
  assign n40794 = n40793 ^ n3211 ^ 1'b0 ;
  assign n40795 = n24368 & ~n40794 ;
  assign n40796 = n7647 ^ n3522 ^ n1707 ;
  assign n40797 = n12809 ^ n1853 ^ 1'b0 ;
  assign n40798 = ~n6829 & n40797 ;
  assign n40799 = ~n40796 & n40798 ;
  assign n40800 = n35071 ^ n20155 ^ 1'b0 ;
  assign n40801 = n40799 | n40800 ;
  assign n40802 = n7632 ^ n360 ^ 1'b0 ;
  assign n40803 = n1895 & n16995 ;
  assign n40804 = ~n4724 & n40803 ;
  assign n40805 = n40802 & n40804 ;
  assign n40806 = n37451 ^ n36471 ^ 1'b0 ;
  assign n40807 = n2321 & ~n35293 ;
  assign n40808 = n22858 & n40807 ;
  assign n40809 = n8161 | n17679 ;
  assign n40810 = n280 & ~n14094 ;
  assign n40811 = n40809 & n40810 ;
  assign n40812 = n40811 ^ n21308 ^ 1'b0 ;
  assign n40813 = n40812 ^ n29707 ^ 1'b0 ;
  assign n40814 = n700 | n25973 ;
  assign n40815 = n13547 | n40814 ;
  assign n40816 = ~n40813 & n40815 ;
  assign n40817 = ~n40733 & n40816 ;
  assign n40818 = n31890 | n32184 ;
  assign n40819 = n13599 & n20919 ;
  assign n40820 = n29649 & n40819 ;
  assign n40821 = ~n17416 & n40820 ;
  assign n40822 = n4780 ^ n1864 ^ 1'b0 ;
  assign n40823 = n40822 ^ n24637 ^ 1'b0 ;
  assign n40824 = ~n49 & n3859 ;
  assign n40825 = n40824 ^ n31674 ^ 1'b0 ;
  assign n40826 = n32167 ^ n16254 ^ 1'b0 ;
  assign n40827 = n19918 ^ n4634 ^ 1'b0 ;
  assign n40828 = n459 & ~n30768 ;
  assign n40829 = n40828 ^ n29176 ^ 1'b0 ;
  assign n40830 = n56 & ~n3612 ;
  assign n40831 = ~n56 & n40830 ;
  assign n40832 = ~n356 & n1943 ;
  assign n40833 = n356 & n40832 ;
  assign n40834 = n40833 ^ n16388 ^ 1'b0 ;
  assign n40835 = n14337 | n40834 ;
  assign n40836 = n40835 ^ n1551 ^ 1'b0 ;
  assign n40837 = n40831 | n40836 ;
  assign n40838 = n5734 & n17771 ;
  assign n40839 = n40837 & n40838 ;
  assign n40840 = n19967 ^ n146 ^ 1'b0 ;
  assign n40841 = n411 & ~n9048 ;
  assign n40842 = n36908 & n40841 ;
  assign n40843 = n40842 ^ n12535 ^ 1'b0 ;
  assign n40844 = n9940 | n38935 ;
  assign n40845 = ( n14885 & n34528 ) | ( n14885 & ~n39970 ) | ( n34528 & ~n39970 ) ;
  assign n40846 = n4476 & n26131 ;
  assign n40847 = n439 & n40846 ;
  assign n40848 = n12576 | n40847 ;
  assign n40849 = n40848 ^ n11876 ^ 1'b0 ;
  assign n40850 = ( n438 & ~n5599 ) | ( n438 & n17189 ) | ( ~n5599 & n17189 ) ;
  assign n40851 = n40850 ^ n20318 ^ 1'b0 ;
  assign n40852 = n5801 | n40851 ;
  assign n40853 = n39604 & ~n40852 ;
  assign n40854 = n40853 ^ n2346 ^ 1'b0 ;
  assign n40855 = n23632 ^ n23291 ^ 1'b0 ;
  assign n40856 = n21539 ^ n6573 ^ 1'b0 ;
  assign n40857 = n13101 ^ n12529 ^ 1'b0 ;
  assign n40858 = ~n17615 & n39521 ;
  assign n40859 = n40858 ^ n38928 ^ 1'b0 ;
  assign n40860 = n22974 & n32891 ;
  assign n40861 = n12725 ^ n10844 ^ 1'b0 ;
  assign n40862 = ~n34190 & n40861 ;
  assign n40863 = ~n15344 & n40862 ;
  assign n40864 = ~n40860 & n40863 ;
  assign n40865 = ~n20653 & n35875 ;
  assign n40866 = ( n13159 & n15068 ) | ( n13159 & n40865 ) | ( n15068 & n40865 ) ;
  assign n40868 = n20700 & ~n34924 ;
  assign n40867 = ~n13150 & n13218 ;
  assign n40869 = n40868 ^ n40867 ^ 1'b0 ;
  assign n40870 = n40869 ^ n36213 ^ 1'b0 ;
  assign n40871 = n33281 & ~n40870 ;
  assign n40872 = n31832 ^ n31463 ^ 1'b0 ;
  assign n40873 = ~n11701 & n40872 ;
  assign n40874 = n20533 ^ n15594 ^ 1'b0 ;
  assign n40875 = n27788 ^ n19473 ^ 1'b0 ;
  assign n40879 = n17631 ^ n8263 ^ 1'b0 ;
  assign n40880 = n24509 | n40879 ;
  assign n40876 = n35665 ^ n30428 ^ n29248 ;
  assign n40877 = n181 & ~n40876 ;
  assign n40878 = ~n8485 & n40877 ;
  assign n40881 = n40880 ^ n40878 ^ n16016 ;
  assign n40882 = n31798 & ~n34079 ;
  assign n40883 = n40679 ^ n14242 ^ 1'b0 ;
  assign n40885 = n14327 ^ n13481 ^ 1'b0 ;
  assign n40886 = ~n20838 & n40885 ;
  assign n40884 = n731 & ~n12968 ;
  assign n40887 = n40886 ^ n40884 ^ 1'b0 ;
  assign n40888 = n20813 ^ n3259 ^ 1'b0 ;
  assign n40889 = n7128 & n22859 ;
  assign n40890 = n15789 & n40889 ;
  assign n40891 = n40890 ^ n33447 ^ 1'b0 ;
  assign n40892 = n9339 & n36317 ;
  assign n40893 = n5973 & n40892 ;
  assign n40894 = n34798 ^ n12793 ^ 1'b0 ;
  assign n40895 = n8995 | n9996 ;
  assign n40896 = n40895 ^ n11969 ^ 1'b0 ;
  assign n40897 = ~n21042 & n21383 ;
  assign n40898 = n29026 & n40897 ;
  assign n40899 = n5247 | n7261 ;
  assign n40900 = ~n188 & n40899 ;
  assign n40901 = n21487 & n35092 ;
  assign n40902 = n25593 & n40901 ;
  assign n40903 = ~n918 & n16745 ;
  assign n40904 = n3445 | n5229 ;
  assign n40905 = n40904 ^ n1157 ^ 1'b0 ;
  assign n40906 = n27723 ^ n16994 ^ 1'b0 ;
  assign n40907 = n4870 & ~n40906 ;
  assign n40908 = n29562 ^ n15068 ^ 1'b0 ;
  assign n40909 = n23361 ^ n4051 ^ 1'b0 ;
  assign n40910 = n31881 ^ n9710 ^ n7673 ;
  assign n40911 = n8906 ^ n3811 ^ 1'b0 ;
  assign n40912 = ~n13326 & n36064 ;
  assign n40913 = n40912 ^ n30889 ^ 1'b0 ;
  assign n40914 = n7936 & ~n21905 ;
  assign n40915 = n19226 & n40914 ;
  assign n40916 = ~n34672 & n39220 ;
  assign n40917 = n11133 ^ n2112 ^ 1'b0 ;
  assign n40918 = ( n22231 & n34153 ) | ( n22231 & n40917 ) | ( n34153 & n40917 ) ;
  assign n40919 = n40532 ^ n22833 ^ 1'b0 ;
  assign n40920 = n21407 | n40919 ;
  assign n40921 = n21490 & n22637 ;
  assign n40922 = n28157 & n40921 ;
  assign n40923 = ~n6213 & n40922 ;
  assign n40924 = n1312 & n9171 ;
  assign n40925 = n21192 & n23276 ;
  assign n40926 = n32412 & n40925 ;
  assign n40927 = ~n39771 & n40926 ;
  assign n40928 = n18871 ^ n3971 ^ 1'b0 ;
  assign n40929 = n11273 | n15829 ;
  assign n40930 = n6353 & n12705 ;
  assign n40931 = n21087 | n38985 ;
  assign n40932 = n12597 | n40931 ;
  assign n40933 = n33875 & n40932 ;
  assign n40934 = ( ~n8945 & n13389 ) | ( ~n8945 & n21859 ) | ( n13389 & n21859 ) ;
  assign n40935 = n40934 ^ n13035 ^ 1'b0 ;
  assign n40936 = ~n21410 & n34277 ;
  assign n40937 = n40936 ^ n33694 ^ n33289 ;
  assign n40938 = ~n3025 & n21944 ;
  assign n40939 = n40938 ^ n40065 ^ 1'b0 ;
  assign n40940 = n12843 & n23577 ;
  assign n40941 = n40940 ^ n17880 ^ 1'b0 ;
  assign n40942 = n5982 & ~n26425 ;
  assign n40943 = n40942 ^ n23179 ^ 1'b0 ;
  assign n40944 = ~n12614 & n17876 ;
  assign n40945 = ~n2550 & n30653 ;
  assign n40946 = n14751 ^ n11955 ^ n2008 ;
  assign n40947 = n40945 & ~n40946 ;
  assign n40948 = n25339 ^ n7889 ^ 1'b0 ;
  assign n40949 = n28458 & n40948 ;
  assign n40950 = n40011 ^ n11546 ^ 1'b0 ;
  assign n40951 = n15969 & n27655 ;
  assign n40952 = n37660 ^ n18219 ^ 1'b0 ;
  assign n40953 = n7624 ^ n875 ^ 1'b0 ;
  assign n40954 = n6637 | n40953 ;
  assign n40955 = n6428 & ~n40954 ;
  assign n40956 = n10498 | n23556 ;
  assign n40957 = n21037 | n40956 ;
  assign n40958 = n2764 & n7705 ;
  assign n40959 = n40958 ^ n27398 ^ 1'b0 ;
  assign n40960 = n40957 & n40959 ;
  assign n40962 = n5755 & ~n7836 ;
  assign n40963 = n40962 ^ n1138 ^ 1'b0 ;
  assign n40961 = n18854 | n22545 ;
  assign n40964 = n40963 ^ n40961 ^ 1'b0 ;
  assign n40965 = n1714 & ~n32789 ;
  assign n40966 = n2815 & n35886 ;
  assign n40967 = n11760 & n40966 ;
  assign n40968 = n21395 ^ n7940 ^ 1'b0 ;
  assign n40969 = n40967 & ~n40968 ;
  assign n40970 = n12939 | n35236 ;
  assign n40971 = ( ~n29827 & n35929 ) | ( ~n29827 & n40970 ) | ( n35929 & n40970 ) ;
  assign n40972 = n5154 & n31078 ;
  assign n40973 = n40972 ^ n280 ^ 1'b0 ;
  assign n40974 = n29030 ^ n2044 ^ 1'b0 ;
  assign n40975 = ~n16470 & n28928 ;
  assign n40976 = n40975 ^ n27087 ^ 1'b0 ;
  assign n40977 = n18190 & n40976 ;
  assign n40980 = n1808 | n37726 ;
  assign n40981 = n1967 & ~n40980 ;
  assign n40978 = n9606 ^ n7156 ^ 1'b0 ;
  assign n40979 = n3576 | n40978 ;
  assign n40982 = n40981 ^ n40979 ^ 1'b0 ;
  assign n40983 = n2594 & ~n40982 ;
  assign n40984 = n18175 & ~n25081 ;
  assign n40985 = ( n7632 & ~n10787 ) | ( n7632 & n15527 ) | ( ~n10787 & n15527 ) ;
  assign n40986 = n36198 ^ n61 ^ 1'b0 ;
  assign n40987 = n24940 & ~n40986 ;
  assign n40988 = n35186 ^ n2262 ^ 1'b0 ;
  assign n40989 = n40988 ^ n15784 ^ 1'b0 ;
  assign n40990 = ~n8648 & n40989 ;
  assign n40991 = n5413 & n31314 ;
  assign n40992 = n2796 & n40991 ;
  assign n40993 = n18379 ^ n12625 ^ 1'b0 ;
  assign n40994 = ~n27425 & n39395 ;
  assign n40995 = n26792 ^ n3213 ^ 1'b0 ;
  assign n40996 = n19207 & ~n40995 ;
  assign n40997 = n3410 & ~n16872 ;
  assign n40998 = n2172 & n40997 ;
  assign n40999 = n40998 ^ n5700 ^ 1'b0 ;
  assign n41000 = n2139 | n34413 ;
  assign n41001 = ( n15877 & n33169 ) | ( n15877 & n41000 ) | ( n33169 & n41000 ) ;
  assign n41002 = n641 | n1174 ;
  assign n41003 = n27629 ^ n7681 ^ 1'b0 ;
  assign n41004 = n1720 | n9153 ;
  assign n41005 = n41004 ^ n15413 ^ 1'b0 ;
  assign n41006 = n6043 & n28066 ;
  assign n41007 = n17219 & n41006 ;
  assign n41008 = n31444 ^ n13823 ^ 1'b0 ;
  assign n41009 = n41007 | n41008 ;
  assign n41010 = n19368 & n40223 ;
  assign n41011 = ~n10612 & n12700 ;
  assign n41012 = n27496 & n41011 ;
  assign n41013 = n11931 ^ n4775 ^ 1'b0 ;
  assign n41014 = n3669 & n8107 ;
  assign n41015 = n41013 & n41014 ;
  assign n41016 = ( n3763 & ~n8001 ) | ( n3763 & n41015 ) | ( ~n8001 & n41015 ) ;
  assign n41017 = ~n13228 & n17045 ;
  assign n41018 = ~n16136 & n41017 ;
  assign n41019 = n1613 | n9063 ;
  assign n41020 = n37157 & ~n41019 ;
  assign n41021 = n14109 & n14839 ;
  assign n41022 = n7391 & n41021 ;
  assign n41023 = n41022 ^ n7152 ^ 1'b0 ;
  assign n41024 = n3574 & n13389 ;
  assign n41025 = n13535 & n37401 ;
  assign n41026 = n41025 ^ n8131 ^ 1'b0 ;
  assign n41027 = n3721 & ~n16359 ;
  assign n41028 = n15360 | n41027 ;
  assign n41029 = n41028 ^ n18236 ^ 1'b0 ;
  assign n41030 = n16223 ^ n4327 ^ 1'b0 ;
  assign n41031 = n35374 & ~n41030 ;
  assign n41032 = n27414 & n30140 ;
  assign n41033 = n13266 & ~n31014 ;
  assign n41034 = n41033 ^ n28642 ^ 1'b0 ;
  assign n41035 = n17744 ^ n1212 ^ n790 ;
  assign n41036 = n37098 & n41035 ;
  assign n41037 = n39703 ^ n14962 ^ n14833 ;
  assign n41038 = ~n6809 & n12868 ;
  assign n41039 = n14009 ^ n4289 ^ 1'b0 ;
  assign n41040 = ~n20559 & n41039 ;
  assign n41041 = n40796 ^ n27466 ^ n8549 ;
  assign n41042 = ~n8376 & n41041 ;
  assign n41043 = ~n21379 & n41042 ;
  assign n41044 = n41043 ^ n22436 ^ 1'b0 ;
  assign n41045 = n3111 & ~n33259 ;
  assign n41046 = ~n15319 & n41045 ;
  assign n41047 = n1247 | n6267 ;
  assign n41048 = n41047 ^ n12840 ^ 1'b0 ;
  assign n41049 = ~n13254 & n17855 ;
  assign n41050 = n7443 & n16690 ;
  assign n41051 = n41050 ^ n15916 ^ 1'b0 ;
  assign n41052 = ~n41049 & n41051 ;
  assign n41053 = n38200 ^ n32977 ^ n14413 ;
  assign n41054 = n35754 ^ n29486 ^ n3766 ;
  assign n41055 = ~n6338 & n14248 ;
  assign n41056 = n26758 ^ n8633 ^ 1'b0 ;
  assign n41057 = n261 | n29227 ;
  assign n41058 = n41056 & ~n41057 ;
  assign n41059 = n32941 ^ n7538 ^ 1'b0 ;
  assign n41060 = ~n33188 & n41059 ;
  assign n41061 = n9821 & ~n41060 ;
  assign n41062 = n17309 ^ n7248 ^ n20 ;
  assign n41063 = n5787 | n26627 ;
  assign n41064 = n41063 ^ n2327 ^ 1'b0 ;
  assign n41065 = n8724 & n24755 ;
  assign n41066 = n5584 & n10223 ;
  assign n41067 = n4916 & n41066 ;
  assign n41068 = n6785 & ~n21315 ;
  assign n41069 = n20039 ^ n18773 ^ 1'b0 ;
  assign n41070 = ~n32751 & n41069 ;
  assign n41071 = ( ~n31264 & n41068 ) | ( ~n31264 & n41070 ) | ( n41068 & n41070 ) ;
  assign n41072 = ~n10645 & n18388 ;
  assign n41073 = n7473 | n27707 ;
  assign n41074 = n26972 & n41073 ;
  assign n41075 = n12013 | n41074 ;
  assign n41076 = ~n25752 & n41075 ;
  assign n41077 = n1134 | n8233 ;
  assign n41078 = n14896 & n24725 ;
  assign n41079 = n14824 & ~n41078 ;
  assign n41080 = n10760 ^ n6969 ^ 1'b0 ;
  assign n41081 = n30997 ^ n8961 ^ 1'b0 ;
  assign n41082 = n25191 | n41081 ;
  assign n41083 = n26249 & n41082 ;
  assign n41084 = n6651 | n41083 ;
  assign n41085 = n37442 ^ n15634 ^ 1'b0 ;
  assign n41086 = n666 & n13798 ;
  assign n41087 = n862 ^ n445 ^ 1'b0 ;
  assign n41088 = n2784 | n41087 ;
  assign n41089 = ~n12967 & n30120 ;
  assign n41090 = n41089 ^ n26700 ^ 1'b0 ;
  assign n41091 = n4690 | n41090 ;
  assign n41092 = n17639 | n40781 ;
  assign n41093 = n41092 ^ n25163 ^ 1'b0 ;
  assign n41094 = n86 & ~n1186 ;
  assign n41095 = n41094 ^ n2940 ^ 1'b0 ;
  assign n41096 = ~n32180 & n34901 ;
  assign n41097 = n9754 ^ n6852 ^ 1'b0 ;
  assign n41098 = n19019 | n41097 ;
  assign n41099 = n3206 & n23927 ;
  assign n41100 = n41099 ^ n25571 ^ 1'b0 ;
  assign n41101 = n29140 ^ n23397 ^ 1'b0 ;
  assign n41102 = n27907 | n41101 ;
  assign n41103 = n17210 | n35387 ;
  assign n41104 = ~n8761 & n9264 ;
  assign n41105 = n27080 & n41104 ;
  assign n41106 = n41105 ^ n22470 ^ 1'b0 ;
  assign n41107 = n41106 ^ n267 ^ 1'b0 ;
  assign n41108 = n30032 ^ n11218 ^ 1'b0 ;
  assign n41109 = ~n30088 & n31442 ;
  assign n41110 = n41109 ^ n28791 ^ 1'b0 ;
  assign n41111 = n5734 & ~n9043 ;
  assign n41112 = n41111 ^ n40548 ^ 1'b0 ;
  assign n41113 = ~n23327 & n41112 ;
  assign n41114 = n2824 | n35608 ;
  assign n41115 = ~n6781 & n16236 ;
  assign n41116 = n2527 & n10158 ;
  assign n41117 = n8147 & n14088 ;
  assign n41118 = ~n41116 & n41117 ;
  assign n41120 = n25488 ^ n15906 ^ n901 ;
  assign n41119 = ~n11559 & n34384 ;
  assign n41121 = n41120 ^ n41119 ^ 1'b0 ;
  assign n41122 = ~n8628 & n11074 ;
  assign n41123 = n41122 ^ n188 ^ 1'b0 ;
  assign n41124 = n6608 | n8346 ;
  assign n41125 = n41124 ^ n3455 ^ 1'b0 ;
  assign n41126 = n41125 ^ n5497 ^ 1'b0 ;
  assign n41127 = n14371 ^ n5022 ^ 1'b0 ;
  assign n41128 = n4949 & ~n41127 ;
  assign n41129 = ( n8725 & ~n36129 ) | ( n8725 & n41128 ) | ( ~n36129 & n41128 ) ;
  assign n41130 = n7413 & ~n21034 ;
  assign n41131 = n29686 ^ n1031 ^ 1'b0 ;
  assign n41132 = n41130 | n41131 ;
  assign n41135 = n14817 ^ n8594 ^ 1'b0 ;
  assign n41136 = n23786 | n41135 ;
  assign n41137 = n17503 & ~n41136 ;
  assign n41133 = n1337 & ~n1743 ;
  assign n41134 = ~n33814 & n41133 ;
  assign n41138 = n41137 ^ n41134 ^ 1'b0 ;
  assign n41140 = n1265 & ~n5145 ;
  assign n41139 = n9348 & n15404 ;
  assign n41141 = n41140 ^ n41139 ^ 1'b0 ;
  assign n41142 = n1656 & ~n41141 ;
  assign n41143 = n22243 ^ n14941 ^ 1'b0 ;
  assign n41144 = n41142 & n41143 ;
  assign n41145 = n37639 ^ n22563 ^ 1'b0 ;
  assign n41146 = n1984 | n11216 ;
  assign n41147 = n7033 ^ n3820 ^ n2370 ;
  assign n41148 = ~n1267 & n37174 ;
  assign n41149 = ~n14499 & n41148 ;
  assign n41150 = ~n5562 & n17321 ;
  assign n41151 = n13933 & ~n16478 ;
  assign n41152 = n41151 ^ n33409 ^ 1'b0 ;
  assign n41153 = n28203 ^ n21892 ^ 1'b0 ;
  assign n41154 = ~n41152 & n41153 ;
  assign n41155 = n41154 ^ n3853 ^ 1'b0 ;
  assign n41156 = n41150 & n41155 ;
  assign n41157 = n25646 ^ n9004 ^ 1'b0 ;
  assign n41158 = n21461 ^ n5952 ^ 1'b0 ;
  assign n41159 = n2018 ^ n1566 ^ 1'b0 ;
  assign n41160 = n12736 & ~n27554 ;
  assign n41161 = n41159 & n41160 ;
  assign n41162 = n13131 | n41161 ;
  assign n41163 = ~n8176 & n10500 ;
  assign n41164 = ~n1235 & n8285 ;
  assign n41165 = ~n27661 & n41164 ;
  assign n41166 = n36673 & n41165 ;
  assign n41167 = n31280 ^ n15101 ^ 1'b0 ;
  assign n41168 = n41167 ^ n26945 ^ n23633 ;
  assign n41169 = n25356 ^ n2118 ^ 1'b0 ;
  assign n41170 = n29442 & n41169 ;
  assign n41171 = n745 & ~n13903 ;
  assign n41172 = ~n12986 & n41171 ;
  assign n41173 = n5995 & n23824 ;
  assign n41174 = n11902 ^ n7784 ^ n4848 ;
  assign n41175 = n8879 & n28667 ;
  assign n41176 = n19770 & ~n34811 ;
  assign n41177 = n1381 | n14594 ;
  assign n41178 = n27312 ^ n8237 ^ 1'b0 ;
  assign n41179 = n41177 | n41178 ;
  assign n41180 = n9923 & n12084 ;
  assign n41181 = n41180 ^ n11055 ^ 1'b0 ;
  assign n41182 = ( ~n19475 & n27515 ) | ( ~n19475 & n41181 ) | ( n27515 & n41181 ) ;
  assign n41183 = n5551 | n6228 ;
  assign n41184 = n24854 | n41183 ;
  assign n41185 = n2980 | n10282 ;
  assign n41186 = ~n12897 & n35528 ;
  assign n41187 = n41186 ^ n1441 ^ 1'b0 ;
  assign n41188 = n26439 ^ n20531 ^ 1'b0 ;
  assign n41189 = n41188 ^ n38329 ^ n8270 ;
  assign n41190 = ~n8009 & n11181 ;
  assign n41191 = ( ~n3695 & n12413 ) | ( ~n3695 & n41190 ) | ( n12413 & n41190 ) ;
  assign n41192 = n6277 | n41191 ;
  assign n41193 = n31207 & ~n41192 ;
  assign n41194 = ( n25890 & n38398 ) | ( n25890 & ~n41193 ) | ( n38398 & ~n41193 ) ;
  assign n41195 = n6128 & ~n34323 ;
  assign n41196 = n700 | n11498 ;
  assign n41197 = n22633 | n41196 ;
  assign n41198 = n20332 & n26727 ;
  assign n41199 = n41198 ^ n16470 ^ 1'b0 ;
  assign n41200 = n15261 ^ n11402 ^ 1'b0 ;
  assign n41201 = n5609 & n19485 ;
  assign n41202 = n41201 ^ n9981 ^ 1'b0 ;
  assign n41203 = n41202 ^ n10616 ^ 1'b0 ;
  assign n41204 = n35539 ^ n8960 ^ 1'b0 ;
  assign n41205 = n5086 | n13620 ;
  assign n41206 = n41205 ^ n22130 ^ 1'b0 ;
  assign n41207 = n41206 ^ n5187 ^ 1'b0 ;
  assign n41208 = ~n19010 & n41207 ;
  assign n41209 = n122 & n4017 ;
  assign n41210 = n29666 ^ n14969 ^ 1'b0 ;
  assign n41211 = n41209 | n41210 ;
  assign n41212 = ( ~n680 & n8009 ) | ( ~n680 & n34673 ) | ( n8009 & n34673 ) ;
  assign n41213 = n41212 ^ n31808 ^ n23324 ;
  assign n41214 = n16439 & ~n36017 ;
  assign n41215 = n8555 & n17661 ;
  assign n41216 = n17465 & n41215 ;
  assign n41217 = ~n15359 & n41216 ;
  assign n41218 = n23677 ^ n10320 ^ 1'b0 ;
  assign n41219 = ~n12475 & n41218 ;
  assign n41220 = ~n2451 & n41219 ;
  assign n41221 = n41220 ^ n15380 ^ 1'b0 ;
  assign n41222 = ~n6101 & n10147 ;
  assign n41223 = ~n5394 & n41222 ;
  assign n41224 = n37070 & n41223 ;
  assign n41225 = n19160 ^ n1941 ^ 1'b0 ;
  assign n41226 = n8970 ^ n7159 ^ 1'b0 ;
  assign n41227 = n10162 & ~n15096 ;
  assign n41228 = n41227 ^ n19193 ^ 1'b0 ;
  assign n41229 = n13578 ^ n717 ^ 1'b0 ;
  assign n41230 = n30731 | n41229 ;
  assign n41231 = n41230 ^ n21259 ^ 1'b0 ;
  assign n41233 = n3143 & ~n5260 ;
  assign n41232 = n41087 ^ n30108 ^ 1'b0 ;
  assign n41234 = n41233 ^ n41232 ^ n35886 ;
  assign n41235 = n10901 ^ n9062 ^ 1'b0 ;
  assign n41236 = ~n41234 & n41235 ;
  assign n41237 = n9940 & ~n10126 ;
  assign n41238 = n9754 ^ n7208 ^ 1'b0 ;
  assign n41245 = n3519 | n33817 ;
  assign n41246 = n896 ^ n35 ^ 1'b0 ;
  assign n41247 = n41245 & n41246 ;
  assign n41239 = n22436 ^ n8334 ^ 1'b0 ;
  assign n41240 = n7162 & ~n41239 ;
  assign n41241 = n41240 ^ n10156 ^ 1'b0 ;
  assign n41242 = n21031 & ~n40577 ;
  assign n41243 = ~n41241 & n41242 ;
  assign n41244 = n14529 | n41243 ;
  assign n41248 = n41247 ^ n41244 ^ 1'b0 ;
  assign n41249 = n7713 | n9043 ;
  assign n41250 = n38269 | n41249 ;
  assign n41251 = n40294 ^ n14325 ^ 1'b0 ;
  assign n41252 = n34970 ^ n4063 ^ 1'b0 ;
  assign n41253 = ~n25091 & n41252 ;
  assign n41254 = ~n366 & n33665 ;
  assign n41255 = n17697 | n25896 ;
  assign n41256 = n13578 | n41255 ;
  assign n41257 = n1177 | n1973 ;
  assign n41258 = n22030 | n41257 ;
  assign n41259 = n16770 & n38387 ;
  assign n41260 = n2202 & ~n4229 ;
  assign n41261 = ~n10486 & n41260 ;
  assign n41262 = n12575 & n41261 ;
  assign n41263 = ( n10562 & n11637 ) | ( n10562 & n41262 ) | ( n11637 & n41262 ) ;
  assign n41264 = n13473 & n17880 ;
  assign n41265 = ~n10908 & n41264 ;
  assign n41266 = ~n27834 & n41265 ;
  assign n41267 = ( n15562 & n17790 ) | ( n15562 & ~n41266 ) | ( n17790 & ~n41266 ) ;
  assign n41268 = n4463 & ~n41267 ;
  assign n41269 = ~n29240 & n40463 ;
  assign n41270 = n26595 ^ n484 ^ 1'b0 ;
  assign n41271 = n24926 ^ n592 ^ 1'b0 ;
  assign n41272 = ~n11552 & n16598 ;
  assign n41273 = n37375 ^ n27045 ^ 1'b0 ;
  assign n41274 = n41272 & ~n41273 ;
  assign n41275 = n911 | n41274 ;
  assign n41277 = n9173 | n23546 ;
  assign n41276 = ~n2492 & n34719 ;
  assign n41278 = n41277 ^ n41276 ^ 1'b0 ;
  assign n41279 = n12448 ^ n1422 ^ 1'b0 ;
  assign n41280 = ~n36528 & n41279 ;
  assign n41281 = ( ~n27703 & n41278 ) | ( ~n27703 & n41280 ) | ( n41278 & n41280 ) ;
  assign n41282 = n7921 | n10598 ;
  assign n41283 = n39417 ^ n32391 ^ n1685 ;
  assign n41284 = n282 & n1701 ;
  assign n41285 = n22545 & n41284 ;
  assign n41286 = n15546 & n36085 ;
  assign n41287 = ~n12488 & n27110 ;
  assign n41288 = n41287 ^ n19535 ^ 1'b0 ;
  assign n41289 = n1530 & ~n8896 ;
  assign n41290 = n4180 & ~n15099 ;
  assign n41291 = ~n41289 & n41290 ;
  assign n41292 = n29914 ^ n12327 ^ 1'b0 ;
  assign n41293 = n2067 | n3449 ;
  assign n41294 = n19135 ^ n3361 ^ 1'b0 ;
  assign n41295 = ~n41293 & n41294 ;
  assign n41296 = n20469 & ~n41295 ;
  assign n41297 = n23814 ^ n14352 ^ 1'b0 ;
  assign n41298 = ( n1615 & n6323 ) | ( n1615 & n41297 ) | ( n6323 & n41297 ) ;
  assign n41299 = ~n3768 & n16084 ;
  assign n41300 = ~n14337 & n26009 ;
  assign n41301 = n41300 ^ n12209 ^ 1'b0 ;
  assign n41302 = x1 & n41301 ;
  assign n41303 = n39022 ^ n448 ^ 1'b0 ;
  assign n41304 = n4947 & ~n33075 ;
  assign n41305 = ~n4624 & n41304 ;
  assign n41306 = ~n3243 & n34833 ;
  assign n41307 = n41306 ^ n14066 ^ 1'b0 ;
  assign n41308 = n7623 | n10998 ;
  assign n41309 = n12187 ^ n8635 ^ 1'b0 ;
  assign n41310 = ~n7697 & n41309 ;
  assign n41311 = n10038 & n10159 ;
  assign n41312 = n6472 & n41311 ;
  assign n41313 = n6704 | n40100 ;
  assign n41314 = n41312 | n41313 ;
  assign n41316 = n3777 & n31482 ;
  assign n41317 = n2643 & n41316 ;
  assign n41318 = ~n49 & n41317 ;
  assign n41315 = ~n2217 & n37436 ;
  assign n41319 = n41318 ^ n41315 ^ 1'b0 ;
  assign n41320 = n5387 | n21152 ;
  assign n41321 = n41320 ^ n5935 ^ 1'b0 ;
  assign n41322 = n8879 ^ n7293 ^ 1'b0 ;
  assign n41323 = ~n27754 & n41322 ;
  assign n41324 = ~n15270 & n41323 ;
  assign n41325 = n20980 ^ n1563 ^ 1'b0 ;
  assign n41326 = n41324 | n41325 ;
  assign n41327 = n11238 & ~n41326 ;
  assign n41328 = n41327 ^ n20446 ^ 1'b0 ;
  assign n41329 = n41019 ^ n26838 ^ n26748 ;
  assign n41330 = n16876 ^ n7907 ^ 1'b0 ;
  assign n41331 = n835 | n13314 ;
  assign n41332 = n2662 & ~n32787 ;
  assign n41333 = ~n20252 & n34673 ;
  assign n41334 = n41333 ^ n19413 ^ 1'b0 ;
  assign n41335 = n8342 & n20397 ;
  assign n41336 = ~n17284 & n34412 ;
  assign n41337 = n41336 ^ n22024 ^ 1'b0 ;
  assign n41338 = ( n1767 & ~n38235 ) | ( n1767 & n41337 ) | ( ~n38235 & n41337 ) ;
  assign n41339 = n9797 | n41338 ;
  assign n41340 = n14184 ^ n7624 ^ 1'b0 ;
  assign n41341 = ~n3736 & n36673 ;
  assign n41342 = n36484 ^ n15760 ^ 1'b0 ;
  assign n41343 = n29129 ^ n1213 ^ 1'b0 ;
  assign n41344 = n17277 ^ n9829 ^ 1'b0 ;
  assign n41345 = n3930 | n8542 ;
  assign n41346 = n41345 ^ n24563 ^ 1'b0 ;
  assign n41347 = n41344 & n41346 ;
  assign n41348 = n41347 ^ n28959 ^ n22153 ;
  assign n41349 = n11070 | n28406 ;
  assign n41350 = n41349 ^ n34849 ^ 1'b0 ;
  assign n41351 = n10480 & n12994 ;
  assign n41352 = n20533 & n41351 ;
  assign n41353 = n20419 & n41352 ;
  assign n41354 = n7368 & ~n19377 ;
  assign n41355 = ~n41353 & n41354 ;
  assign n41356 = n17735 & n26922 ;
  assign n41357 = n41356 ^ n30406 ^ 1'b0 ;
  assign n41358 = n23200 ^ n1853 ^ 1'b0 ;
  assign n41359 = n37496 & n41358 ;
  assign n41360 = n13413 | n31503 ;
  assign n41361 = n34060 | n41360 ;
  assign n41362 = n31996 | n36271 ;
  assign n41363 = n20479 & n41362 ;
  assign n41364 = n41363 ^ n17177 ^ 1'b0 ;
  assign n41365 = n13716 ^ n5998 ^ 1'b0 ;
  assign n41366 = n26156 ^ n5490 ^ 1'b0 ;
  assign n41367 = n35916 ^ n14793 ^ 1'b0 ;
  assign n41368 = ~n1186 & n21135 ;
  assign n41369 = n10864 | n22041 ;
  assign n41370 = n41369 ^ n21447 ^ 1'b0 ;
  assign n41371 = ~n3720 & n5328 ;
  assign n41372 = ( n7497 & n41370 ) | ( n7497 & ~n41371 ) | ( n41370 & ~n41371 ) ;
  assign n41373 = n4087 & n33040 ;
  assign n41374 = n17372 ^ n3691 ^ 1'b0 ;
  assign n41375 = n41373 & n41374 ;
  assign n41376 = n12950 & ~n36318 ;
  assign n41377 = n41376 ^ n23571 ^ 1'b0 ;
  assign n41378 = ~n1956 & n2102 ;
  assign n41379 = n9173 ^ n7887 ^ 1'b0 ;
  assign n41380 = n4814 | n41379 ;
  assign n41382 = n1980 & n28870 ;
  assign n41381 = n10558 & ~n23637 ;
  assign n41383 = n41382 ^ n41381 ^ 1'b0 ;
  assign n41384 = n4993 ^ n738 ^ 1'b0 ;
  assign n41385 = n2336 & ~n17800 ;
  assign n41386 = ~n12293 & n41385 ;
  assign n41387 = ( n5316 & ~n41384 ) | ( n5316 & n41386 ) | ( ~n41384 & n41386 ) ;
  assign n41388 = n5480 & n17316 ;
  assign n41389 = ~n16517 & n41388 ;
  assign n41390 = n13308 ^ n2247 ^ 1'b0 ;
  assign n41391 = n41389 & ~n41390 ;
  assign n41392 = n8801 & n11588 ;
  assign n41393 = n41392 ^ n11515 ^ 1'b0 ;
  assign n41394 = n41393 ^ n17799 ^ 1'b0 ;
  assign n41395 = ~n6833 & n41394 ;
  assign n41396 = n41395 ^ n12576 ^ 1'b0 ;
  assign n41397 = n448 | n41396 ;
  assign n41398 = n16788 & ~n31010 ;
  assign n41399 = n41398 ^ n20844 ^ 1'b0 ;
  assign n41400 = n41399 ^ n30838 ^ 1'b0 ;
  assign n41401 = n10866 | n41400 ;
  assign n41403 = n2185 | n34635 ;
  assign n41402 = n5104 & ~n20063 ;
  assign n41404 = n41403 ^ n41402 ^ 1'b0 ;
  assign n41405 = n3770 & ~n38935 ;
  assign n41406 = n41405 ^ n5814 ^ 1'b0 ;
  assign n41407 = n41406 ^ n37986 ^ 1'b0 ;
  assign n41408 = n6989 | n22783 ;
  assign n41409 = n41408 ^ n26235 ^ 1'b0 ;
  assign n41410 = n26064 ^ n3985 ^ 1'b0 ;
  assign n41411 = n26901 & n41410 ;
  assign n41412 = n38125 ^ n1434 ^ 1'b0 ;
  assign n41413 = n18616 & ~n41412 ;
  assign n41414 = n5886 & ~n32940 ;
  assign n41415 = n4079 ^ n2876 ^ 1'b0 ;
  assign n41416 = n9598 & n41415 ;
  assign n41417 = n9827 ^ n3802 ^ 1'b0 ;
  assign n41418 = n41416 & ~n41417 ;
  assign n41419 = ( ~n6374 & n8478 ) | ( ~n6374 & n41418 ) | ( n8478 & n41418 ) ;
  assign n41420 = n9319 ^ n8451 ^ n3429 ;
  assign n41421 = n41420 ^ n25657 ^ 1'b0 ;
  assign n41422 = n21514 & ~n22445 ;
  assign n41423 = n41421 & n41422 ;
  assign n41425 = n8547 ^ n3350 ^ n1534 ;
  assign n41426 = n7830 & n41425 ;
  assign n41427 = ~n9732 & n41426 ;
  assign n41424 = ~n4442 & n38441 ;
  assign n41428 = n41427 ^ n41424 ^ 1'b0 ;
  assign n41429 = n15413 ^ n5589 ^ 1'b0 ;
  assign n41430 = n3049 & ~n41429 ;
  assign n41431 = n12911 & n41430 ;
  assign n41436 = n2219 & ~n3729 ;
  assign n41437 = n41436 ^ n7586 ^ 1'b0 ;
  assign n41432 = n18273 | n19351 ;
  assign n41433 = n8074 | n36692 ;
  assign n41434 = n41433 ^ n3335 ^ 1'b0 ;
  assign n41435 = ( n18784 & n41432 ) | ( n18784 & ~n41434 ) | ( n41432 & ~n41434 ) ;
  assign n41438 = n41437 ^ n41435 ^ n4964 ;
  assign n41439 = n6259 & ~n25298 ;
  assign n41440 = n9795 & n41439 ;
  assign n41441 = n6326 & ~n41440 ;
  assign n41442 = n41441 ^ n1138 ^ 1'b0 ;
  assign n41443 = ( n12185 & n17971 ) | ( n12185 & ~n41442 ) | ( n17971 & ~n41442 ) ;
  assign n41444 = n4486 & n18084 ;
  assign n41445 = n25296 ^ n3039 ^ 1'b0 ;
  assign n41446 = ~n30509 & n41445 ;
  assign n41447 = ~n26500 & n26756 ;
  assign n41448 = n8435 ^ n1419 ^ 1'b0 ;
  assign n41449 = n8593 & n11520 ;
  assign n41450 = n31338 & n41449 ;
  assign n41451 = ~n12897 & n15819 ;
  assign n41452 = n41451 ^ n16695 ^ 1'b0 ;
  assign n41453 = n40911 & n41452 ;
  assign n41454 = n41450 & n41453 ;
  assign n41455 = ~n999 & n39917 ;
  assign n41456 = n41455 ^ n17806 ^ 1'b0 ;
  assign n41457 = n15206 ^ n12323 ^ 1'b0 ;
  assign n41458 = n33962 ^ n1971 ^ 1'b0 ;
  assign n41459 = ~n11291 & n41458 ;
  assign n41460 = ~n4038 & n41459 ;
  assign n41461 = n30708 ^ n1653 ^ 1'b0 ;
  assign n41462 = n22636 & n41461 ;
  assign n41463 = n6690 & n32629 ;
  assign n41464 = n18108 & ~n35814 ;
  assign n41465 = n7984 | n12153 ;
  assign n41466 = ~n5821 & n32883 ;
  assign n41467 = n16381 | n41466 ;
  assign n41468 = n41467 ^ n4318 ^ 1'b0 ;
  assign n41469 = n8621 ^ n3066 ^ 1'b0 ;
  assign n41470 = n3906 & n5215 ;
  assign n41471 = ~n737 & n41470 ;
  assign n41472 = n41471 ^ n4832 ^ 1'b0 ;
  assign n41473 = n9067 & ~n41472 ;
  assign n41474 = n41473 ^ n6533 ^ 1'b0 ;
  assign n41475 = n41469 & ~n41474 ;
  assign n41476 = n2356 ^ n1235 ^ 1'b0 ;
  assign n41477 = ~n40545 & n41476 ;
  assign n41478 = n41477 ^ n40542 ^ n8376 ;
  assign n41479 = n21725 ^ n20393 ^ n3162 ;
  assign n41480 = n2448 & n6954 ;
  assign n41481 = n17973 & n41480 ;
  assign n41487 = n4164 & n16193 ;
  assign n41488 = n7624 & ~n41487 ;
  assign n41482 = n34753 ^ n11238 ^ 1'b0 ;
  assign n41483 = ~n6437 & n41482 ;
  assign n41484 = ~n10910 & n26113 ;
  assign n41485 = ~n41483 & n41484 ;
  assign n41486 = n13885 & ~n41485 ;
  assign n41489 = n41488 ^ n41486 ^ 1'b0 ;
  assign n41490 = n20114 ^ n11210 ^ 1'b0 ;
  assign n41491 = n33131 & n41490 ;
  assign n41492 = n9341 | n26347 ;
  assign n41494 = ~n6729 & n14092 ;
  assign n41493 = n19762 ^ n1884 ^ 1'b0 ;
  assign n41495 = n41494 ^ n41493 ^ n38371 ;
  assign n41496 = n1297 & n41495 ;
  assign n41497 = n9156 & n25144 ;
  assign n41498 = ~n41496 & n41497 ;
  assign n41499 = ~n5961 & n7908 ;
  assign n41500 = n41499 ^ n560 ^ 1'b0 ;
  assign n41501 = n21546 ^ n21111 ^ 1'b0 ;
  assign n41502 = n3078 | n41501 ;
  assign n41503 = n41502 ^ n29048 ^ 1'b0 ;
  assign n41504 = n17760 | n29788 ;
  assign n41505 = n8949 & n37845 ;
  assign n41506 = n20969 ^ n10624 ^ 1'b0 ;
  assign n41507 = ~n33016 & n41506 ;
  assign n41508 = ~n8906 & n41507 ;
  assign n41509 = n41508 ^ n20695 ^ 1'b0 ;
  assign n41510 = n8003 ^ n5562 ^ 1'b0 ;
  assign n41511 = ( ~n3417 & n18305 ) | ( ~n3417 & n41510 ) | ( n18305 & n41510 ) ;
  assign n41512 = n12188 & ~n24256 ;
  assign n41513 = ~n4363 & n41512 ;
  assign n41514 = ( n3783 & ~n9351 ) | ( n3783 & n41513 ) | ( ~n9351 & n41513 ) ;
  assign n41515 = n35863 ^ n6468 ^ 1'b0 ;
  assign n41516 = ~n4092 & n27373 ;
  assign n41517 = n23762 & n41516 ;
  assign n41518 = n3668 & ~n8771 ;
  assign n41519 = ~n30581 & n41518 ;
  assign n41520 = n22340 | n33349 ;
  assign n41521 = n41520 ^ n32672 ^ 1'b0 ;
  assign n41522 = n31918 ^ n27078 ^ 1'b0 ;
  assign n41523 = n6114 | n41522 ;
  assign n41524 = ( n7825 & n22857 ) | ( n7825 & n41352 ) | ( n22857 & n41352 ) ;
  assign n41525 = n41524 ^ n19595 ^ 1'b0 ;
  assign n41526 = n1401 & ~n41525 ;
  assign n41527 = n38356 ^ n20166 ^ 1'b0 ;
  assign n41529 = n3919 ^ n3571 ^ 1'b0 ;
  assign n41530 = n31728 & ~n41529 ;
  assign n41528 = n8596 | n28096 ;
  assign n41531 = n41530 ^ n41528 ^ 1'b0 ;
  assign n41532 = ~n2812 & n5086 ;
  assign n41533 = n41532 ^ n15403 ^ 1'b0 ;
  assign n41534 = ~n28872 & n41533 ;
  assign n41535 = ~n8435 & n32659 ;
  assign n41536 = n38003 ^ n26780 ^ 1'b0 ;
  assign n41537 = n12193 | n24886 ;
  assign n41538 = n41537 ^ n11905 ^ 1'b0 ;
  assign n41539 = ~n10033 & n41538 ;
  assign n41540 = n41539 ^ n40586 ^ 1'b0 ;
  assign n41541 = n15058 ^ n3001 ^ n1930 ;
  assign n41542 = ( ~n1267 & n2899 ) | ( ~n1267 & n6409 ) | ( n2899 & n6409 ) ;
  assign n41543 = n1450 & n41542 ;
  assign n41544 = n8216 & ~n41543 ;
  assign n41545 = n41544 ^ n14400 ^ 1'b0 ;
  assign n41546 = n41541 & ~n41545 ;
  assign n41547 = n8521 & n41546 ;
  assign n41548 = n23913 ^ n774 ^ 1'b0 ;
  assign n41549 = ~n25438 & n41548 ;
  assign n41550 = n5501 & ~n33221 ;
  assign n41551 = n35173 & ~n41550 ;
  assign n41552 = n6978 & ~n18582 ;
  assign n41553 = n41552 ^ n16549 ^ 1'b0 ;
  assign n41554 = n41553 ^ n15879 ^ 1'b0 ;
  assign n41555 = n15533 ^ n14207 ^ 1'b0 ;
  assign n41556 = n40064 & n41555 ;
  assign n41558 = n24054 & n35749 ;
  assign n41557 = n7528 & n23156 ;
  assign n41559 = n41558 ^ n41557 ^ 1'b0 ;
  assign n41560 = n16596 ^ n10146 ^ 1'b0 ;
  assign n41561 = n4479 | n41560 ;
  assign n41562 = n5982 ^ n311 ^ 1'b0 ;
  assign n41563 = n41562 ^ n24458 ^ 1'b0 ;
  assign n41564 = n24084 ^ n21045 ^ n14614 ;
  assign n41565 = n2373 & n41564 ;
  assign n41566 = ~n126 & n19702 ;
  assign n41567 = n1435 & ~n25937 ;
  assign n41568 = n3896 & n12379 ;
  assign n41569 = n24772 ^ n6457 ^ 1'b0 ;
  assign n41570 = n30302 ^ n331 ^ 1'b0 ;
  assign n41571 = n41570 ^ n36313 ^ 1'b0 ;
  assign n41572 = n41569 & n41571 ;
  assign n41573 = n18869 ^ n7697 ^ 1'b0 ;
  assign n41574 = ( ~n1983 & n7076 ) | ( ~n1983 & n20102 ) | ( n7076 & n20102 ) ;
  assign n41575 = ( ~n18516 & n41573 ) | ( ~n18516 & n41574 ) | ( n41573 & n41574 ) ;
  assign n41576 = n13346 & n36367 ;
  assign n41577 = n41576 ^ n21264 ^ 1'b0 ;
  assign n41578 = n14132 | n24703 ;
  assign n41579 = n41578 ^ n17204 ^ 1'b0 ;
  assign n41580 = ( n26549 & n29590 ) | ( n26549 & n41579 ) | ( n29590 & n41579 ) ;
  assign n41581 = n646 & ~n41580 ;
  assign n41582 = n3882 | n41581 ;
  assign n41583 = n41582 ^ n15279 ^ 1'b0 ;
  assign n41584 = n13541 ^ n7430 ^ 1'b0 ;
  assign n41585 = n41584 ^ n39686 ^ n17231 ;
  assign n41586 = n9364 | n15347 ;
  assign n41587 = n20530 ^ n11543 ^ 1'b0 ;
  assign n41588 = n11661 | n41587 ;
  assign n41589 = n28338 ^ n3962 ^ 1'b0 ;
  assign n41590 = n41588 | n41589 ;
  assign n41591 = n4679 & ~n41590 ;
  assign n41592 = ~n51 & n15656 ;
  assign n41593 = ~n18909 & n41592 ;
  assign n41594 = ( n515 & n6766 ) | ( n515 & ~n41593 ) | ( n6766 & ~n41593 ) ;
  assign n41595 = n24576 ^ n18980 ^ n3529 ;
  assign n41596 = n14658 & n41595 ;
  assign n41597 = n13327 | n16718 ;
  assign n41598 = n39218 & ~n41597 ;
  assign n41599 = n738 | n5901 ;
  assign n41600 = n7816 ^ n2678 ^ 1'b0 ;
  assign n41601 = n41599 & ~n41600 ;
  assign n41602 = ~n41371 & n41601 ;
  assign n41603 = n8008 | n41602 ;
  assign n41604 = ~n22929 & n33287 ;
  assign n41605 = n8012 | n23699 ;
  assign n41606 = n41605 ^ n5369 ^ 1'b0 ;
  assign n41607 = n41606 ^ n13134 ^ n3891 ;
  assign n41608 = n13270 ^ n10917 ^ 1'b0 ;
  assign n41609 = ~n12413 & n41608 ;
  assign n41610 = ~n17696 & n41609 ;
  assign n41611 = n21924 ^ n6127 ^ 1'b0 ;
  assign n41612 = n21843 | n41611 ;
  assign n41613 = n798 & ~n801 ;
  assign n41614 = n28061 & ~n41613 ;
  assign n41615 = n4933 & n41614 ;
  assign n41621 = ~n7100 & n7726 ;
  assign n41622 = n41621 ^ n2163 ^ 1'b0 ;
  assign n41616 = n3674 & ~n12592 ;
  assign n41617 = n3858 & n41616 ;
  assign n41618 = n5216 & ~n6898 ;
  assign n41619 = n41617 & n41618 ;
  assign n41620 = n5279 | n41619 ;
  assign n41623 = n41622 ^ n41620 ^ 1'b0 ;
  assign n41624 = n30499 ^ n9325 ^ 1'b0 ;
  assign n41625 = n7416 & ~n40792 ;
  assign n41626 = ~n5757 & n9114 ;
  assign n41627 = n41626 ^ n13616 ^ 1'b0 ;
  assign n41628 = n41627 ^ n28844 ^ n1907 ;
  assign n41629 = ~n39008 & n41628 ;
  assign n41630 = n35857 ^ n28583 ^ n1558 ;
  assign n41631 = n17773 | n41630 ;
  assign n41632 = ~n39683 & n41631 ;
  assign n41633 = n12375 | n33365 ;
  assign n41634 = n4665 & ~n5497 ;
  assign n41635 = n41634 ^ n8491 ^ 1'b0 ;
  assign n41636 = n12249 ^ n1024 ^ n339 ;
  assign n41637 = n41635 & ~n41636 ;
  assign n41638 = n41633 & n41637 ;
  assign n41639 = n5748 & n16364 ;
  assign n41640 = n41639 ^ n25233 ^ 1'b0 ;
  assign n41641 = n37694 ^ n22694 ^ 1'b0 ;
  assign n41642 = n356 & n23856 ;
  assign n41643 = n31315 ^ n2136 ^ 1'b0 ;
  assign n41644 = n5018 & ~n5610 ;
  assign n41645 = n41644 ^ n30374 ^ 1'b0 ;
  assign n41646 = n35861 ^ n14173 ^ 1'b0 ;
  assign n41647 = n17281 & n41646 ;
  assign n41648 = n13605 ^ n8243 ^ 1'b0 ;
  assign n41649 = n1967 & ~n5724 ;
  assign n41650 = n7270 & n41649 ;
  assign n41651 = n744 & ~n5508 ;
  assign n41652 = n41651 ^ n6273 ^ 1'b0 ;
  assign n41653 = ~n510 & n41652 ;
  assign n41654 = n41653 ^ n36669 ^ 1'b0 ;
  assign n41655 = n20772 | n28707 ;
  assign n41656 = n22863 & ~n41655 ;
  assign n41657 = n41656 ^ n41167 ^ 1'b0 ;
  assign n41658 = n26879 & n41657 ;
  assign n41659 = ~n5329 & n41658 ;
  assign n41660 = n26383 ^ n4413 ^ 1'b0 ;
  assign n41661 = ~n858 & n12354 ;
  assign n41662 = n41661 ^ n24493 ^ 1'b0 ;
  assign n41663 = n3331 & ~n7254 ;
  assign n41664 = ~n4975 & n35801 ;
  assign n41665 = n34913 ^ n16880 ^ n6350 ;
  assign n41666 = n2751 | n41665 ;
  assign n41667 = n2780 & n21784 ;
  assign n41668 = n3205 & ~n8012 ;
  assign n41669 = n10923 ^ n10893 ^ 1'b0 ;
  assign n41670 = n8195 ^ n2095 ^ 1'b0 ;
  assign n41671 = n14750 | n25385 ;
  assign n41672 = n25063 ^ n23621 ^ n21125 ;
  assign n41673 = n5906 ^ n2048 ^ 1'b0 ;
  assign n41674 = n11485 & ~n41673 ;
  assign n41675 = n22494 ^ n18665 ^ 1'b0 ;
  assign n41677 = n22218 ^ n1517 ^ 1'b0 ;
  assign n41676 = ~n4853 & n30783 ;
  assign n41678 = n41677 ^ n41676 ^ 1'b0 ;
  assign n41679 = n27692 ^ n26746 ^ 1'b0 ;
  assign n41680 = n20930 & n41679 ;
  assign n41681 = ~n36996 & n37085 ;
  assign n41682 = n10778 & ~n19664 ;
  assign n41685 = n8308 & n12026 ;
  assign n41686 = ~n24006 & n41685 ;
  assign n41687 = n41686 ^ n16007 ^ 1'b0 ;
  assign n41683 = n6100 | n29088 ;
  assign n41684 = n29060 | n41683 ;
  assign n41688 = n41687 ^ n41684 ^ 1'b0 ;
  assign n41689 = n38142 ^ n35625 ^ n33647 ;
  assign n41690 = n10886 ^ n1187 ^ 1'b0 ;
  assign n41691 = ~n630 & n19437 ;
  assign n41692 = n22885 ^ n7696 ^ 1'b0 ;
  assign n41693 = n18838 & n41692 ;
  assign n41694 = n3564 & n10245 ;
  assign n41695 = n12658 & ~n41694 ;
  assign n41696 = n5360 & n16130 ;
  assign n41697 = n37407 & n41696 ;
  assign n41699 = ( ~n19945 & n22871 ) | ( ~n19945 & n31085 ) | ( n22871 & n31085 ) ;
  assign n41698 = n1785 & n30382 ;
  assign n41700 = n41699 ^ n41698 ^ 1'b0 ;
  assign n41701 = ~n9535 & n15195 ;
  assign n41702 = n41701 ^ n9715 ^ 1'b0 ;
  assign n41703 = n41702 ^ n14750 ^ 1'b0 ;
  assign n41704 = n4473 | n16563 ;
  assign n41705 = ( n4772 & ~n6741 ) | ( n4772 & n41704 ) | ( ~n6741 & n41704 ) ;
  assign n41706 = n19681 ^ n11711 ^ 1'b0 ;
  assign n41707 = ~n9204 & n41706 ;
  assign n41708 = n23379 & n41707 ;
  assign n41709 = n2421 ^ n1946 ^ 1'b0 ;
  assign n41710 = n35401 & ~n41709 ;
  assign n41711 = n34567 ^ n27723 ^ 1'b0 ;
  assign n41712 = n37306 & ~n41711 ;
  assign n41713 = n41712 ^ n8989 ^ 1'b0 ;
  assign n41714 = n9155 & ~n19254 ;
  assign n41715 = n3533 & n15657 ;
  assign n41716 = n41715 ^ n18077 ^ 1'b0 ;
  assign n41717 = ~n10706 & n29879 ;
  assign n41718 = ( n2124 & ~n22445 ) | ( n2124 & n37075 ) | ( ~n22445 & n37075 ) ;
  assign n41719 = ( ~n304 & n2261 ) | ( ~n304 & n10552 ) | ( n2261 & n10552 ) ;
  assign n41720 = n7861 ^ n6203 ^ 1'b0 ;
  assign n41721 = n41720 ^ n2014 ^ 1'b0 ;
  assign n41722 = ~n11610 & n41721 ;
  assign n41723 = n21597 ^ n14904 ^ 1'b0 ;
  assign n41724 = n12842 | n41723 ;
  assign n41725 = n5629 ^ n3571 ^ 1'b0 ;
  assign n41726 = n18755 ^ n11813 ^ 1'b0 ;
  assign n41727 = n41726 ^ n21748 ^ 1'b0 ;
  assign n41728 = ~n18044 & n38349 ;
  assign n41729 = n1693 & ~n20840 ;
  assign n41730 = ~n3386 & n36151 ;
  assign n41731 = n41730 ^ n5420 ^ 1'b0 ;
  assign n41732 = ( n2242 & ~n16888 ) | ( n2242 & n36883 ) | ( ~n16888 & n36883 ) ;
  assign n41733 = n17601 & n26214 ;
  assign n41734 = n12534 & n21527 ;
  assign n41735 = n41734 ^ n2164 ^ 1'b0 ;
  assign n41736 = n24391 ^ n20969 ^ 1'b0 ;
  assign n41737 = ~n21562 & n41736 ;
  assign n41738 = ~n28101 & n41737 ;
  assign n41739 = n38047 ^ n5627 ^ 1'b0 ;
  assign n41740 = n34238 & ~n41739 ;
  assign n41741 = ~n12113 & n17050 ;
  assign n41742 = n16456 ^ n3174 ^ 1'b0 ;
  assign n41743 = n1876 & n41742 ;
  assign n41744 = n11358 & n41743 ;
  assign n41745 = ~n6032 & n41744 ;
  assign n41746 = n2773 | n3272 ;
  assign n41747 = n8352 & ~n41746 ;
  assign n41748 = n41745 & n41747 ;
  assign n41749 = n36835 & n41737 ;
  assign n41750 = n14264 & n41749 ;
  assign n41751 = n41750 ^ n1481 ^ 1'b0 ;
  assign n41752 = n31322 | n41751 ;
  assign n41753 = n17423 | n23961 ;
  assign n41754 = n33425 | n41753 ;
  assign n41755 = ( n1293 & n8512 ) | ( n1293 & ~n13986 ) | ( n8512 & ~n13986 ) ;
  assign n41756 = n19146 ^ n5514 ^ 1'b0 ;
  assign n41757 = ~n41755 & n41756 ;
  assign n41758 = n26838 ^ n3924 ^ 1'b0 ;
  assign n41759 = n41757 & ~n41758 ;
  assign n41760 = n26013 ^ n493 ^ n195 ;
  assign n41761 = ~n4422 & n12412 ;
  assign n41762 = ~n3764 & n41761 ;
  assign n41763 = n41762 ^ n22332 ^ n796 ;
  assign n41765 = ~n559 & n29648 ;
  assign n41766 = n2996 & n41765 ;
  assign n41764 = n8904 ^ n7057 ^ n673 ;
  assign n41767 = n41766 ^ n41764 ^ n25671 ;
  assign n41768 = n41763 & n41767 ;
  assign n41769 = n2389 ^ n368 ^ 1'b0 ;
  assign n41770 = n4390 | n41769 ;
  assign n41771 = n20868 ^ n12177 ^ 1'b0 ;
  assign n41772 = ~n5055 & n41771 ;
  assign n41773 = n41772 ^ n13299 ^ 1'b0 ;
  assign n41774 = n19982 | n41773 ;
  assign n41775 = n41770 & ~n41774 ;
  assign n41776 = ~n1664 & n3565 ;
  assign n41777 = n41776 ^ n2403 ^ 1'b0 ;
  assign n41778 = n41777 ^ n17378 ^ 1'b0 ;
  assign n41779 = n13287 ^ n160 ^ 1'b0 ;
  assign n41780 = n698 | n3932 ;
  assign n41781 = n41780 ^ n19975 ^ n7966 ;
  assign n41783 = n32597 ^ n32539 ^ 1'b0 ;
  assign n41782 = ~n22751 & n28007 ;
  assign n41784 = n41783 ^ n41782 ^ 1'b0 ;
  assign n41785 = n17220 ^ n13717 ^ 1'b0 ;
  assign n41786 = ~n41784 & n41785 ;
  assign n41787 = n40510 ^ n28003 ^ 1'b0 ;
  assign n41788 = n1337 & ~n12156 ;
  assign n41789 = ~n4770 & n41788 ;
  assign n41790 = n4142 & ~n41789 ;
  assign n41791 = n3032 & n41790 ;
  assign n41792 = n2358 | n16753 ;
  assign n41793 = n31625 ^ n24326 ^ 1'b0 ;
  assign n41794 = n4386 & n7375 ;
  assign n41795 = n16163 & n29025 ;
  assign n41796 = n41795 ^ n32694 ^ 1'b0 ;
  assign n41797 = n2532 & n20472 ;
  assign n41798 = n10300 & ~n21504 ;
  assign n41799 = n10245 & n10587 ;
  assign n41800 = n12715 & n41799 ;
  assign n41801 = n7520 ^ n568 ^ 1'b0 ;
  assign n41802 = n4347 & n34947 ;
  assign n41803 = ~n15252 & n22859 ;
  assign n41804 = n41803 ^ n4097 ^ 1'b0 ;
  assign n41805 = ~n17635 & n22029 ;
  assign n41806 = n41805 ^ n27349 ^ n15861 ;
  assign n41807 = n8983 | n27717 ;
  assign n41808 = n24678 | n41807 ;
  assign n41809 = n41808 ^ n33670 ^ 1'b0 ;
  assign n41810 = n5346 & n23077 ;
  assign n41811 = n9129 ^ n5692 ^ 1'b0 ;
  assign n41812 = n22359 & ~n41811 ;
  assign n41813 = n5258 | n6363 ;
  assign n41814 = n41813 ^ n36461 ^ 1'b0 ;
  assign n41815 = n21146 ^ n5827 ^ 1'b0 ;
  assign n41816 = n727 & n14637 ;
  assign n41817 = n33993 ^ n12731 ^ 1'b0 ;
  assign n41818 = n41816 & n41817 ;
  assign n41819 = n41818 ^ n2671 ^ 1'b0 ;
  assign n41820 = n25786 & n41819 ;
  assign n41821 = n41820 ^ n133 ^ 1'b0 ;
  assign n41822 = n5888 & ~n11133 ;
  assign n41823 = n271 & n41822 ;
  assign n41824 = n32201 & n41823 ;
  assign n41826 = n8519 ^ n1366 ^ 1'b0 ;
  assign n41827 = n8656 & ~n41826 ;
  assign n41825 = ~n135 & n4545 ;
  assign n41828 = n41827 ^ n41825 ^ 1'b0 ;
  assign n41829 = ~n2048 & n7797 ;
  assign n41830 = n41829 ^ n33349 ^ 1'b0 ;
  assign n41831 = ~n30249 & n41830 ;
  assign n41832 = n21730 ^ n2292 ^ 1'b0 ;
  assign n41833 = n21042 & n41832 ;
  assign n41834 = n16209 & ~n16343 ;
  assign n41835 = ~n29294 & n41834 ;
  assign n41836 = n41835 ^ n40988 ^ 1'b0 ;
  assign n41837 = n35708 ^ n17927 ^ 1'b0 ;
  assign n41844 = n2864 & n13690 ;
  assign n41838 = n10227 ^ n3108 ^ 1'b0 ;
  assign n41839 = ~n8720 & n41838 ;
  assign n41840 = n7601 | n18893 ;
  assign n41841 = n1723 & n41840 ;
  assign n41842 = ~n34493 & n41841 ;
  assign n41843 = ~n41839 & n41842 ;
  assign n41845 = n41844 ^ n41843 ^ 1'b0 ;
  assign n41846 = n16405 ^ n4461 ^ 1'b0 ;
  assign n41847 = ~n20457 & n41846 ;
  assign n41848 = n41847 ^ n14027 ^ 1'b0 ;
  assign n41849 = n7590 & n40899 ;
  assign n41850 = n41849 ^ n28762 ^ 1'b0 ;
  assign n41851 = n10361 & ~n41850 ;
  assign n41852 = ~n41848 & n41851 ;
  assign n41853 = n23715 ^ n302 ^ 1'b0 ;
  assign n41854 = n14385 ^ n1561 ^ 1'b0 ;
  assign n41855 = n1025 & ~n41854 ;
  assign n41856 = n41855 ^ n996 ^ 1'b0 ;
  assign n41857 = ~n22582 & n41856 ;
  assign n41858 = n7449 & ~n41857 ;
  assign n41859 = n23049 ^ n1469 ^ 1'b0 ;
  assign n41860 = n10915 & n41859 ;
  assign n41861 = n41860 ^ n1365 ^ 1'b0 ;
  assign n41862 = n41861 ^ n21447 ^ 1'b0 ;
  assign n41863 = n40234 ^ n7207 ^ 1'b0 ;
  assign n41864 = n14612 & ~n41863 ;
  assign n41865 = ~n10075 & n32172 ;
  assign n41866 = n41865 ^ n4216 ^ 1'b0 ;
  assign n41867 = n4313 & ~n41866 ;
  assign n41868 = ~n41864 & n41867 ;
  assign n41869 = n17881 ^ n3001 ^ 1'b0 ;
  assign n41870 = n27723 ^ n26701 ^ n12950 ;
  assign n41871 = ~n10558 & n22794 ;
  assign n41872 = n41871 ^ n16988 ^ 1'b0 ;
  assign n41873 = n11196 & n37322 ;
  assign n41874 = n18009 ^ n11099 ^ n2324 ;
  assign n41875 = ( ~n18301 & n41873 ) | ( ~n18301 & n41874 ) | ( n41873 & n41874 ) ;
  assign n41876 = n27802 & n41875 ;
  assign n41877 = n41876 ^ n6037 ^ 1'b0 ;
  assign n41878 = n41877 ^ n29772 ^ 1'b0 ;
  assign n41879 = n1226 & ~n25659 ;
  assign n41880 = n12558 & n41879 ;
  assign n41881 = n12490 ^ n6522 ^ 1'b0 ;
  assign n41882 = n15940 | n20233 ;
  assign n41883 = n41882 ^ n34186 ^ 1'b0 ;
  assign n41884 = n2283 | n24180 ;
  assign n41885 = n28675 ^ n3181 ^ 1'b0 ;
  assign n41886 = n41885 ^ n20662 ^ n4583 ;
  assign n41887 = n41886 ^ n25822 ^ 1'b0 ;
  assign n41888 = n41884 | n41887 ;
  assign n41889 = n26069 ^ n18664 ^ 1'b0 ;
  assign n41890 = ( ~n10234 & n17116 ) | ( ~n10234 & n20631 ) | ( n17116 & n20631 ) ;
  assign n41891 = n16455 & ~n41890 ;
  assign n41892 = n37453 ^ n36357 ^ 1'b0 ;
  assign n41893 = ~n2943 & n17981 ;
  assign n41894 = n41893 ^ n1476 ^ 1'b0 ;
  assign n41895 = n41894 ^ n26360 ^ n7482 ;
  assign n41896 = n31143 & ~n41895 ;
  assign n41897 = n1601 | n25340 ;
  assign n41898 = n18556 & ~n41897 ;
  assign n41899 = n7641 & n41898 ;
  assign n41900 = n448 & n41899 ;
  assign n41901 = n2288 | n16320 ;
  assign n41902 = n1865 & ~n41901 ;
  assign n41903 = n41902 ^ n27785 ^ 1'b0 ;
  assign n41904 = n22898 ^ n16356 ^ 1'b0 ;
  assign n41905 = n443 & n41904 ;
  assign n41908 = n2426 & ~n21168 ;
  assign n41906 = n11294 ^ n7518 ^ 1'b0 ;
  assign n41907 = n725 & ~n41906 ;
  assign n41909 = n41908 ^ n41907 ^ n2996 ;
  assign n41910 = n1811 & n2437 ;
  assign n41911 = n10828 | n17827 ;
  assign n41912 = n41910 | n41911 ;
  assign n41913 = n41912 ^ n24720 ^ n1029 ;
  assign n41914 = n13406 ^ n13272 ^ 1'b0 ;
  assign n41915 = n38102 & n41914 ;
  assign n41916 = ~n9232 & n12985 ;
  assign n41917 = ~n2469 & n12666 ;
  assign n41918 = n41916 & n41917 ;
  assign n41919 = n41918 ^ n10217 ^ 1'b0 ;
  assign n41920 = n3554 | n41919 ;
  assign n41921 = ( ~n746 & n2248 ) | ( ~n746 & n4688 ) | ( n2248 & n4688 ) ;
  assign n41922 = n41921 ^ n24860 ^ 1'b0 ;
  assign n41923 = x11 & n41922 ;
  assign n41924 = n41923 ^ n35452 ^ 1'b0 ;
  assign n41925 = n41924 ^ n36471 ^ 1'b0 ;
  assign n41926 = n35119 ^ n23601 ^ n16853 ;
  assign n41927 = ~n10996 & n41909 ;
  assign n41928 = n12335 | n38838 ;
  assign n41929 = n41928 ^ n40407 ^ 1'b0 ;
  assign n41930 = n5005 | n39223 ;
  assign n41931 = n386 & ~n41930 ;
  assign n41932 = ( n9433 & n39971 ) | ( n9433 & n41931 ) | ( n39971 & n41931 ) ;
  assign n41933 = n37507 ^ n23208 ^ n209 ;
  assign n41934 = ~n2539 & n26693 ;
  assign n41935 = n20781 ^ n18185 ^ 1'b0 ;
  assign n41936 = n23678 & n39253 ;
  assign n41937 = n5431 & n6527 ;
  assign n41938 = n41937 ^ n1469 ^ 1'b0 ;
  assign n41939 = n41936 & ~n41938 ;
  assign n41940 = n914 & ~n6832 ;
  assign n41941 = ~n16578 & n41940 ;
  assign n41942 = n19786 ^ n17491 ^ 1'b0 ;
  assign n41943 = ~n15120 & n41942 ;
  assign n41944 = n20460 ^ n963 ^ 1'b0 ;
  assign n41945 = n41943 & n41944 ;
  assign n41946 = n23243 & n41945 ;
  assign n41947 = ~n24313 & n41946 ;
  assign n41948 = n17812 ^ n13458 ^ 1'b0 ;
  assign n41949 = n4077 & n41948 ;
  assign n41950 = n23946 ^ n11364 ^ 1'b0 ;
  assign n41951 = n23891 & n41950 ;
  assign n41952 = ( n5992 & ~n10907 ) | ( n5992 & n18545 ) | ( ~n10907 & n18545 ) ;
  assign n41953 = ~n11014 & n22834 ;
  assign n41954 = ( n39884 & ~n41219 ) | ( n39884 & n41953 ) | ( ~n41219 & n41953 ) ;
  assign n41955 = n5103 & ~n6765 ;
  assign n41956 = n30532 & n40942 ;
  assign n41957 = n26472 ^ n21515 ^ n17649 ;
  assign n41958 = ( ~n17775 & n41956 ) | ( ~n17775 & n41957 ) | ( n41956 & n41957 ) ;
  assign n41959 = n18124 | n38371 ;
  assign n41960 = n2724 | n5684 ;
  assign n41961 = n41960 ^ n20056 ^ 1'b0 ;
  assign n41962 = n6293 | n9950 ;
  assign n41963 = n6024 | n37742 ;
  assign n41964 = n41963 ^ n3479 ^ 1'b0 ;
  assign n41965 = n582 & n8886 ;
  assign n41966 = n41965 ^ n13465 ^ n11689 ;
  assign n41967 = n1912 & ~n41966 ;
  assign n41968 = n6498 & ~n13488 ;
  assign n41969 = ~n41967 & n41968 ;
  assign n41970 = n3704 & ~n41969 ;
  assign n41971 = n6429 & n41970 ;
  assign n41972 = n18773 ^ n12040 ^ 1'b0 ;
  assign n41973 = ~n35628 & n41972 ;
  assign n41974 = n26858 | n41973 ;
  assign n41975 = n451 & ~n3741 ;
  assign n41976 = n39315 & n41975 ;
  assign n41977 = ( n379 & n13794 ) | ( n379 & n19702 ) | ( n13794 & n19702 ) ;
  assign n41978 = n22166 ^ n16387 ^ 1'b0 ;
  assign n41979 = n41978 ^ n40480 ^ n37650 ;
  assign n41980 = n18392 ^ n12608 ^ 1'b0 ;
  assign n41981 = n14503 ^ n7609 ^ 1'b0 ;
  assign n41982 = n41980 & ~n41981 ;
  assign n41983 = n36764 ^ n9270 ^ 1'b0 ;
  assign n41984 = n205 ^ n150 ^ 1'b0 ;
  assign n41985 = n5786 & ~n41984 ;
  assign n41986 = n12337 & ~n31511 ;
  assign n41987 = n10721 & ~n23287 ;
  assign n41988 = n41987 ^ n12757 ^ 1'b0 ;
  assign n41989 = n41988 ^ n35050 ^ 1'b0 ;
  assign n41991 = n10520 & ~n15117 ;
  assign n41992 = n20153 & n41991 ;
  assign n41993 = n41992 ^ n12131 ^ 1'b0 ;
  assign n41994 = n25215 | n41993 ;
  assign n41990 = n2925 & n24137 ;
  assign n41995 = n41994 ^ n41990 ^ 1'b0 ;
  assign n41996 = ~n85 & n4837 ;
  assign n41997 = n41996 ^ n23325 ^ 1'b0 ;
  assign n41998 = ( n2128 & ~n8070 ) | ( n2128 & n11105 ) | ( ~n8070 & n11105 ) ;
  assign n41999 = n41998 ^ n35116 ^ 1'b0 ;
  assign n42000 = n8105 & n32408 ;
  assign n42001 = n42000 ^ n40742 ^ 1'b0 ;
  assign n42002 = n18844 ^ n15816 ^ 1'b0 ;
  assign n42003 = n12450 ^ n667 ^ 1'b0 ;
  assign n42004 = n31290 | n42003 ;
  assign n42005 = n37001 ^ n32641 ^ n6844 ;
  assign n42006 = n42004 | n42005 ;
  assign n42007 = n38190 ^ n22597 ^ 1'b0 ;
  assign n42008 = n14152 | n42007 ;
  assign n42009 = n10552 | n12541 ;
  assign n42010 = n42009 ^ n30902 ^ 1'b0 ;
  assign n42011 = ( n4558 & ~n22101 ) | ( n4558 & n34039 ) | ( ~n22101 & n34039 ) ;
  assign n42013 = n6179 ^ n4048 ^ n2438 ;
  assign n42014 = ~n25902 & n42013 ;
  assign n42012 = n1016 & ~n23170 ;
  assign n42015 = n42014 ^ n42012 ^ 1'b0 ;
  assign n42017 = n11295 ^ n4767 ^ 1'b0 ;
  assign n42016 = n17866 ^ n2899 ^ 1'b0 ;
  assign n42018 = n42017 ^ n42016 ^ 1'b0 ;
  assign n42019 = n32709 & n42018 ;
  assign n42020 = n4028 ^ n776 ^ 1'b0 ;
  assign n42021 = n10048 | n10211 ;
  assign n42022 = n33153 ^ n7391 ^ 1'b0 ;
  assign n42023 = n42021 & ~n42022 ;
  assign n42024 = n32715 ^ n32525 ^ 1'b0 ;
  assign n42025 = n24273 & ~n42024 ;
  assign n42026 = n36550 & n42025 ;
  assign n42027 = ~n23541 & n42026 ;
  assign n42028 = n5224 & ~n9121 ;
  assign n42029 = n42028 ^ n21636 ^ n14823 ;
  assign n42034 = ~n2483 & n28752 ;
  assign n42035 = n42034 ^ n498 ^ 1'b0 ;
  assign n42036 = n26628 ^ n584 ^ 1'b0 ;
  assign n42037 = ~n42035 & n42036 ;
  assign n42030 = n18996 & ~n19005 ;
  assign n42031 = n42030 ^ n14787 ^ 1'b0 ;
  assign n42032 = n42031 ^ n2623 ^ 1'b0 ;
  assign n42033 = ~n4931 & n42032 ;
  assign n42038 = n42037 ^ n42033 ^ n132 ;
  assign n42039 = n737 | n9696 ;
  assign n42040 = n4651 | n42039 ;
  assign n42041 = n3062 & n12377 ;
  assign n42042 = ~n12377 & n19047 ;
  assign n42043 = n34924 ^ n612 ^ 1'b0 ;
  assign n42044 = n42042 & n42043 ;
  assign n42045 = n3674 ^ n3524 ^ 1'b0 ;
  assign n42046 = n42044 & n42045 ;
  assign n42047 = n846 | n23953 ;
  assign n42048 = ~n36436 & n42047 ;
  assign n42049 = n16699 ^ n16480 ^ 1'b0 ;
  assign n42050 = n42049 ^ n38993 ^ n21653 ;
  assign n42051 = n14376 & ~n32846 ;
  assign n42052 = n21965 & n42047 ;
  assign n42053 = ~n857 & n27236 ;
  assign n42054 = ~n27236 & n42053 ;
  assign n42055 = n4104 & ~n7188 ;
  assign n42056 = ~n4104 & n42055 ;
  assign n42057 = n42056 ^ n34630 ^ 1'b0 ;
  assign n42058 = n42057 ^ n38208 ^ 1'b0 ;
  assign n42059 = n42054 | n42058 ;
  assign n42060 = n4146 & n8281 ;
  assign n42061 = n10939 & n42060 ;
  assign n42062 = n42061 ^ n2258 ^ 1'b0 ;
  assign n42063 = n11961 ^ n3284 ^ 1'b0 ;
  assign n42064 = n23733 ^ n12009 ^ n5581 ;
  assign n42065 = ~n42063 & n42064 ;
  assign n42066 = n8230 ^ n6927 ^ 1'b0 ;
  assign n42067 = n15792 & n42066 ;
  assign n42068 = n214 & ~n846 ;
  assign n42069 = ~n723 & n42068 ;
  assign n42070 = n37922 & ~n42069 ;
  assign n42071 = n42070 ^ n23008 ^ 1'b0 ;
  assign n42072 = n7609 | n40232 ;
  assign n42073 = n42072 ^ n3835 ^ 1'b0 ;
  assign n42074 = ( n1466 & ~n10544 ) | ( n1466 & n42073 ) | ( ~n10544 & n42073 ) ;
  assign n42075 = ~n10814 & n22027 ;
  assign n42076 = n16768 ^ n10094 ^ 1'b0 ;
  assign n42077 = n19749 & ~n36030 ;
  assign n42078 = n42077 ^ n33357 ^ 1'b0 ;
  assign n42079 = n11532 & ~n42078 ;
  assign n42080 = ~n23015 & n42079 ;
  assign n42081 = n3455 & ~n11722 ;
  assign n42082 = n14594 & n28040 ;
  assign n42083 = n42082 ^ n10107 ^ 1'b0 ;
  assign n42085 = n3361 & ~n29877 ;
  assign n42084 = n12599 & ~n25764 ;
  assign n42086 = n42085 ^ n42084 ^ 1'b0 ;
  assign n42087 = n42086 ^ n2605 ^ 1'b0 ;
  assign n42088 = n39534 ^ n1513 ^ 1'b0 ;
  assign n42089 = n6299 & n16398 ;
  assign n42090 = ~n1563 & n42089 ;
  assign n42091 = n1138 & n42090 ;
  assign n42092 = ( n2980 & n13706 ) | ( n2980 & ~n16396 ) | ( n13706 & ~n16396 ) ;
  assign n42093 = n7188 | n8176 ;
  assign n42094 = ~n1353 & n14442 ;
  assign n42095 = n32173 ^ n11353 ^ 1'b0 ;
  assign n42096 = n42095 ^ n5612 ^ 1'b0 ;
  assign n42097 = n29972 | n42096 ;
  assign n42098 = n11727 & ~n42097 ;
  assign n42099 = n22563 ^ n5438 ^ 1'b0 ;
  assign n42100 = ~n26055 & n42099 ;
  assign n42101 = n24537 ^ n19192 ^ n6910 ;
  assign n42102 = n29296 & n42101 ;
  assign n42103 = ~n42100 & n42102 ;
  assign n42104 = n42103 ^ n36761 ^ 1'b0 ;
  assign n42105 = n29103 ^ n15484 ^ 1'b0 ;
  assign n42106 = ~n38377 & n42105 ;
  assign n42107 = n22558 & n42106 ;
  assign n42108 = ~n3977 & n16745 ;
  assign n42109 = n6472 & n42108 ;
  assign n42110 = n35909 ^ n29387 ^ 1'b0 ;
  assign n42111 = n14909 ^ n5892 ^ 1'b0 ;
  assign n42112 = n376 & n42111 ;
  assign n42113 = ~n42110 & n42112 ;
  assign n42114 = n2358 & n30272 ;
  assign n42115 = ~n13854 & n32279 ;
  assign n42116 = n2632 & ~n3182 ;
  assign n42117 = n8754 & n42116 ;
  assign n42118 = n42117 ^ n3770 ^ 1'b0 ;
  assign n42119 = n8281 & n12647 ;
  assign n42120 = n17927 ^ n3818 ^ 1'b0 ;
  assign n42121 = n33435 ^ n6088 ^ 1'b0 ;
  assign n42122 = ~n22756 & n36285 ;
  assign n42123 = ~n37322 & n42122 ;
  assign n42124 = n24664 ^ n23768 ^ 1'b0 ;
  assign n42125 = n10542 | n42124 ;
  assign n42126 = n2956 | n8279 ;
  assign n42127 = n33065 | n42126 ;
  assign n42128 = ~n1978 & n42127 ;
  assign n42129 = ~n14750 & n24807 ;
  assign n42130 = ( ~n19528 & n21105 ) | ( ~n19528 & n34334 ) | ( n21105 & n34334 ) ;
  assign n42131 = n8684 | n10526 ;
  assign n42132 = n42131 ^ n22799 ^ 1'b0 ;
  assign n42133 = ( n6267 & n31285 ) | ( n6267 & n42132 ) | ( n31285 & n42132 ) ;
  assign n42134 = n1943 & n32503 ;
  assign n42135 = n42134 ^ n13083 ^ 1'b0 ;
  assign n42136 = n12159 & n42135 ;
  assign n42137 = n14364 & n20616 ;
  assign n42138 = n19942 ^ n49 ^ 1'b0 ;
  assign n42139 = n42137 | n42138 ;
  assign n42140 = n7344 | n10944 ;
  assign n42141 = ( ~n1939 & n26663 ) | ( ~n1939 & n35224 ) | ( n26663 & n35224 ) ;
  assign n42142 = n13055 ^ n10841 ^ 1'b0 ;
  assign n42143 = ~n25232 & n38455 ;
  assign n42144 = n5600 | n42143 ;
  assign n42145 = n8156 ^ n5076 ^ 1'b0 ;
  assign n42146 = n22297 ^ n3235 ^ 1'b0 ;
  assign n42147 = n42146 ^ n2394 ^ 1'b0 ;
  assign n42148 = n3361 & ~n42147 ;
  assign n42149 = n42145 & n42148 ;
  assign n42150 = n42149 ^ n6120 ^ 1'b0 ;
  assign n42151 = n3279 ^ n1369 ^ 1'b0 ;
  assign n42152 = ~n24642 & n42151 ;
  assign n42153 = n3240 & n22341 ;
  assign n42154 = n7585 & n42153 ;
  assign n42155 = n42154 ^ n458 ^ 1'b0 ;
  assign n42156 = n38342 ^ n18946 ^ n14212 ;
  assign n42157 = n23938 ^ n10769 ^ n9751 ;
  assign n42158 = n32743 ^ n21533 ^ 1'b0 ;
  assign n42159 = ~n23714 & n38553 ;
  assign n42160 = n32921 & n42159 ;
  assign n42161 = n5905 | n30253 ;
  assign n42162 = n42161 ^ n3830 ^ 1'b0 ;
  assign n42163 = ~n7961 & n42162 ;
  assign n42164 = n42163 ^ n33863 ^ 1'b0 ;
  assign n42165 = ~n5154 & n25530 ;
  assign n42166 = ~n37369 & n42165 ;
  assign n42169 = n433 & ~n39763 ;
  assign n42167 = n17908 ^ n6662 ^ 1'b0 ;
  assign n42168 = n6742 | n42167 ;
  assign n42170 = n42169 ^ n42168 ^ 1'b0 ;
  assign n42171 = n15091 ^ n13897 ^ n4302 ;
  assign n42172 = n32399 ^ n22206 ^ 1'b0 ;
  assign n42173 = ~n23270 & n42172 ;
  assign n42174 = n42171 & n42173 ;
  assign n42175 = n25073 ^ n14215 ^ 1'b0 ;
  assign n42176 = n8507 & n42175 ;
  assign n42177 = ~n36954 & n42176 ;
  assign n42178 = ( ~n4034 & n7865 ) | ( ~n4034 & n14380 ) | ( n7865 & n14380 ) ;
  assign n42179 = n42178 ^ n13561 ^ 1'b0 ;
  assign n42180 = n2615 & n42179 ;
  assign n42181 = n16068 ^ n11118 ^ 1'b0 ;
  assign n42182 = n42180 | n42181 ;
  assign n42183 = ~n6553 & n9772 ;
  assign n42184 = n42183 ^ n8815 ^ 1'b0 ;
  assign n42185 = n9682 & n32662 ;
  assign n42186 = ~n42184 & n42185 ;
  assign n42187 = n13367 ^ n7268 ^ 1'b0 ;
  assign n42188 = n17714 ^ n11965 ^ 1'b0 ;
  assign n42189 = n27185 & n42188 ;
  assign n42190 = n31919 ^ n11764 ^ 1'b0 ;
  assign n42191 = ( ~n21296 & n23931 ) | ( ~n21296 & n37278 ) | ( n23931 & n37278 ) ;
  assign n42192 = n34425 ^ n8219 ^ 1'b0 ;
  assign n42193 = n283 & n42192 ;
  assign n42194 = n1907 & n41322 ;
  assign n42195 = n18175 & ~n29718 ;
  assign n42196 = ~n7696 & n42195 ;
  assign n42197 = n42196 ^ n39538 ^ 1'b0 ;
  assign n42198 = n15966 & ~n42197 ;
  assign n42199 = n32113 ^ n9934 ^ 1'b0 ;
  assign n42200 = ~n12303 & n39718 ;
  assign n42201 = ( n4729 & ~n4864 ) | ( n4729 & n8447 ) | ( ~n4864 & n8447 ) ;
  assign n42202 = n10720 & ~n42201 ;
  assign n42203 = ~n1080 & n42202 ;
  assign n42204 = n42203 ^ n38963 ^ 1'b0 ;
  assign n42205 = n24043 ^ n7185 ^ 1'b0 ;
  assign n42206 = n8814 ^ n5704 ^ 1'b0 ;
  assign n42207 = n42205 & n42206 ;
  assign n42208 = n42207 ^ n41874 ^ 1'b0 ;
  assign n42209 = n3303 ^ n1814 ^ 1'b0 ;
  assign n42210 = n19959 & ~n21213 ;
  assign n42211 = n9832 & n42210 ;
  assign n42212 = ( n4667 & n29791 ) | ( n4667 & n42211 ) | ( n29791 & n42211 ) ;
  assign n42213 = n4790 & ~n42212 ;
  assign n42214 = n42213 ^ n19726 ^ 1'b0 ;
  assign n42215 = n2568 & n7668 ;
  assign n42216 = n2854 & n10609 ;
  assign n42217 = n17917 & n42216 ;
  assign n42218 = n40081 ^ n5535 ^ 1'b0 ;
  assign n42219 = ( n7488 & n16744 ) | ( n7488 & ~n32839 ) | ( n16744 & ~n32839 ) ;
  assign n42220 = n10751 & n13331 ;
  assign n42221 = ~n42219 & n42220 ;
  assign n42224 = n20101 & n30517 ;
  assign n42225 = n5860 ^ n5325 ^ 1'b0 ;
  assign n42226 = ~n42224 & n42225 ;
  assign n42223 = n12640 & n35016 ;
  assign n42227 = n42226 ^ n42223 ^ n28403 ;
  assign n42222 = n4506 & ~n27628 ;
  assign n42228 = n42227 ^ n42222 ^ 1'b0 ;
  assign n42229 = n19558 ^ n10735 ^ 1'b0 ;
  assign n42230 = ~n9546 & n42229 ;
  assign n42231 = ~n436 & n32800 ;
  assign n42232 = ( n7713 & n20372 ) | ( n7713 & ~n32873 ) | ( n20372 & ~n32873 ) ;
  assign n42233 = n7972 | n21681 ;
  assign n42234 = n42232 & ~n42233 ;
  assign n42235 = n5444 & ~n12300 ;
  assign n42236 = n42235 ^ n24749 ^ 1'b0 ;
  assign n42237 = n28143 ^ n22474 ^ n9959 ;
  assign n42238 = n21077 ^ n9368 ^ 1'b0 ;
  assign n42239 = n42238 ^ n32328 ^ 1'b0 ;
  assign n42240 = n944 | n4512 ;
  assign n42241 = n15051 | n18324 ;
  assign n42242 = n42241 ^ n15843 ^ 1'b0 ;
  assign n42243 = n17123 & n42242 ;
  assign n42244 = ~n12825 & n42243 ;
  assign n42245 = n42244 ^ n6189 ^ 1'b0 ;
  assign n42246 = ~n2296 & n17686 ;
  assign n42247 = n9453 & n42246 ;
  assign n42248 = n11763 | n42247 ;
  assign n42249 = n26787 & ~n42248 ;
  assign n42250 = ~n5321 & n15760 ;
  assign n42251 = ~n7876 & n42250 ;
  assign n42252 = n18211 ^ n1961 ^ 1'b0 ;
  assign n42253 = n2440 & ~n19466 ;
  assign n42254 = n42253 ^ n1915 ^ 1'b0 ;
  assign n42255 = ( ~n39505 & n42252 ) | ( ~n39505 & n42254 ) | ( n42252 & n42254 ) ;
  assign n42256 = n4347 & ~n42255 ;
  assign n42257 = n42256 ^ n872 ^ 1'b0 ;
  assign n42258 = n3034 | n42257 ;
  assign n42259 = n32755 | n42258 ;
  assign n42260 = ( n10401 & ~n16751 ) | ( n10401 & n20333 ) | ( ~n16751 & n20333 ) ;
  assign n42261 = ( n1096 & n31372 ) | ( n1096 & ~n42260 ) | ( n31372 & ~n42260 ) ;
  assign n42262 = n21632 ^ n5001 ^ n269 ;
  assign n42263 = ~n3742 & n7307 ;
  assign n42264 = n29339 ^ n28119 ^ 1'b0 ;
  assign n42265 = n17906 & n42264 ;
  assign n42266 = ~n10143 & n42265 ;
  assign n42267 = ~n21765 & n42266 ;
  assign n42268 = n8525 | n42267 ;
  assign n42269 = n6185 & ~n6989 ;
  assign n42270 = n42269 ^ n27606 ^ 1'b0 ;
  assign n42271 = n4428 | n38834 ;
  assign n42272 = n6322 & n13002 ;
  assign n42273 = ~n5946 & n42272 ;
  assign n42274 = n35160 & ~n41784 ;
  assign n42275 = n42274 ^ n15719 ^ 1'b0 ;
  assign n42279 = n5829 ^ n4200 ^ 1'b0 ;
  assign n42276 = n37389 ^ n25469 ^ 1'b0 ;
  assign n42277 = n12018 & ~n42276 ;
  assign n42278 = n12760 & n42277 ;
  assign n42280 = n42279 ^ n42278 ^ 1'b0 ;
  assign n42281 = n34086 & ~n42280 ;
  assign n42282 = n11232 & n42281 ;
  assign n42283 = n42282 ^ n11315 ^ n7358 ;
  assign n42284 = ~n5757 & n10245 ;
  assign n42285 = ~n31967 & n42284 ;
  assign n42286 = n8981 ^ n7368 ^ 1'b0 ;
  assign n42287 = n33388 | n42286 ;
  assign n42288 = n11144 & n42287 ;
  assign n42289 = n37782 ^ n11573 ^ 1'b0 ;
  assign n42290 = ~n16696 & n26989 ;
  assign n42291 = n8608 | n29500 ;
  assign n42292 = ( ~n7067 & n19889 ) | ( ~n7067 & n42291 ) | ( n19889 & n42291 ) ;
  assign n42293 = ~n42257 & n42292 ;
  assign n42294 = ( n23555 & n27278 ) | ( n23555 & n28359 ) | ( n27278 & n28359 ) ;
  assign n42298 = ~n22915 & n33571 ;
  assign n42295 = n3446 | n28144 ;
  assign n42296 = n30032 | n42295 ;
  assign n42297 = n37399 & n42296 ;
  assign n42299 = n42298 ^ n42297 ^ 1'b0 ;
  assign n42300 = n8945 ^ n8057 ^ 1'b0 ;
  assign n42301 = n42299 & ~n42300 ;
  assign n42302 = n12433 & ~n25371 ;
  assign n42303 = n42302 ^ n3097 ^ 1'b0 ;
  assign n42304 = ~n4484 & n5847 ;
  assign n42305 = n42304 ^ n19032 ^ 1'b0 ;
  assign n42306 = n17281 & ~n19879 ;
  assign n42307 = n15120 | n15316 ;
  assign n42308 = n194 | n42307 ;
  assign n42309 = n13691 & ~n18303 ;
  assign n42310 = n42309 ^ n16234 ^ 1'b0 ;
  assign n42311 = n42310 ^ n23633 ^ 1'b0 ;
  assign n42312 = ~n12139 & n21086 ;
  assign n42313 = n1293 & n42312 ;
  assign n42314 = ( n13351 & n30437 ) | ( n13351 & n42313 ) | ( n30437 & n42313 ) ;
  assign n42315 = ~n2833 & n3070 ;
  assign n42316 = n9664 & ~n42315 ;
  assign n42317 = n42316 ^ n36293 ^ 1'b0 ;
  assign n42318 = n5719 | n27815 ;
  assign n42319 = n42318 ^ n9304 ^ 1'b0 ;
  assign n42320 = n22131 & n42319 ;
  assign n42321 = n25783 ^ n10137 ^ 1'b0 ;
  assign n42322 = ~n1897 & n13489 ;
  assign n42323 = ~n5682 & n42322 ;
  assign n42324 = n36974 ^ n29704 ^ 1'b0 ;
  assign n42325 = ~n21436 & n42324 ;
  assign n42327 = ~n6114 & n28120 ;
  assign n42328 = n5336 & n42327 ;
  assign n42329 = n42328 ^ n30941 ^ 1'b0 ;
  assign n42326 = ~n9383 & n26072 ;
  assign n42330 = n42329 ^ n42326 ^ 1'b0 ;
  assign n42331 = n15431 | n29545 ;
  assign n42332 = n5788 | n15542 ;
  assign n42333 = n24406 | n42332 ;
  assign n42334 = n6274 & n42333 ;
  assign n42335 = n1774 ^ n1715 ^ 1'b0 ;
  assign n42336 = n4519 | n42335 ;
  assign n42337 = n42336 ^ n262 ^ 1'b0 ;
  assign n42339 = ~n2865 & n5354 ;
  assign n42340 = ~n30276 & n42339 ;
  assign n42338 = n4754 | n12782 ;
  assign n42341 = n42340 ^ n42338 ^ 1'b0 ;
  assign n42342 = n7759 & ~n17648 ;
  assign n42343 = n13909 | n39753 ;
  assign n42344 = n6100 | n19884 ;
  assign n42345 = n42344 ^ n4474 ^ 1'b0 ;
  assign n42346 = n2543 & ~n14009 ;
  assign n42347 = n28421 & n42346 ;
  assign n42348 = n2802 | n7077 ;
  assign n42350 = n7322 & n22050 ;
  assign n42351 = n3279 & n42350 ;
  assign n42349 = n18509 & ~n32184 ;
  assign n42352 = n42351 ^ n42349 ^ n21555 ;
  assign n42353 = n42352 ^ n15727 ^ 1'b0 ;
  assign n42354 = n11675 & ~n40724 ;
  assign n42355 = ~n7765 & n9058 ;
  assign n42356 = n42355 ^ n6093 ^ 1'b0 ;
  assign n42357 = ~n1370 & n42356 ;
  assign n42358 = n42357 ^ n32940 ^ 1'b0 ;
  assign n42359 = ( n1323 & ~n6278 ) | ( n1323 & n14123 ) | ( ~n6278 & n14123 ) ;
  assign n42360 = n18526 | n42359 ;
  assign n42361 = n29491 ^ n3926 ^ 1'b0 ;
  assign n42362 = n10391 ^ n4634 ^ 1'b0 ;
  assign n42363 = n32422 & ~n42362 ;
  assign n42364 = n31524 ^ n825 ^ 1'b0 ;
  assign n42365 = n2138 & n2343 ;
  assign n42366 = n42365 ^ n32831 ^ 1'b0 ;
  assign n42367 = n2389 & n42151 ;
  assign n42368 = n1584 & n19274 ;
  assign n42369 = n983 & n42368 ;
  assign n42370 = ~n38261 & n42369 ;
  assign n42373 = n8495 & ~n28205 ;
  assign n42374 = n42373 ^ n3649 ^ 1'b0 ;
  assign n42375 = n4407 & ~n42374 ;
  assign n42376 = n13176 & n42375 ;
  assign n42371 = n430 & n2223 ;
  assign n42372 = ~n7412 & n42371 ;
  assign n42377 = n42376 ^ n42372 ^ 1'b0 ;
  assign n42378 = ~n6888 & n16106 ;
  assign n42379 = n14208 ^ n4914 ^ 1'b0 ;
  assign n42380 = n42378 & ~n42379 ;
  assign n42381 = n31221 ^ n3399 ^ 1'b0 ;
  assign n42382 = n40213 ^ n17221 ^ 1'b0 ;
  assign n42383 = n8200 | n11616 ;
  assign n42384 = n42383 ^ n8103 ^ 1'b0 ;
  assign n42385 = n42384 ^ n37515 ^ 1'b0 ;
  assign n42386 = n42162 & ~n42385 ;
  assign n42387 = n42386 ^ n12343 ^ 1'b0 ;
  assign n42388 = n13618 & n16286 ;
  assign n42389 = n42388 ^ n29987 ^ n26249 ;
  assign n42390 = n106 & n42389 ;
  assign n42391 = n1182 & n31617 ;
  assign n42392 = n37927 | n42391 ;
  assign n42393 = n3611 & ~n42392 ;
  assign n42394 = n8879 & ~n22982 ;
  assign n42395 = ~n27358 & n42394 ;
  assign n42396 = n42395 ^ n24038 ^ 1'b0 ;
  assign n42397 = ~n2900 & n42396 ;
  assign n42398 = n13777 ^ n8246 ^ 1'b0 ;
  assign n42399 = n16047 ^ n2313 ^ 1'b0 ;
  assign n42400 = n42398 & ~n42399 ;
  assign n42401 = ( n4357 & n20556 ) | ( n4357 & n42400 ) | ( n20556 & n42400 ) ;
  assign n42402 = ~n5814 & n42401 ;
  assign n42403 = n25325 ^ n7191 ^ 1'b0 ;
  assign n42404 = n15850 & n34360 ;
  assign n42405 = n11235 ^ n11135 ^ 1'b0 ;
  assign n42406 = n15193 & ~n22630 ;
  assign n42407 = n2956 | n35297 ;
  assign n42408 = ( n25929 & n42406 ) | ( n25929 & ~n42407 ) | ( n42406 & ~n42407 ) ;
  assign n42409 = n18616 ^ n1014 ^ 1'b0 ;
  assign n42410 = n16188 & n31657 ;
  assign n42411 = ~n10411 & n23505 ;
  assign n42412 = n42411 ^ n9827 ^ 1'b0 ;
  assign n42413 = n162 | n23285 ;
  assign n42414 = n780 & ~n42413 ;
  assign n42415 = ( n17416 & ~n22333 ) | ( n17416 & n42414 ) | ( ~n22333 & n42414 ) ;
  assign n42416 = n10575 ^ n6124 ^ 1'b0 ;
  assign n42417 = n21404 & n42416 ;
  assign n42418 = n37593 ^ n27471 ^ 1'b0 ;
  assign n42419 = n42417 & ~n42418 ;
  assign n42420 = ~n26569 & n42419 ;
  assign n42421 = n38342 ^ n10425 ^ 1'b0 ;
  assign n42422 = n3661 | n42421 ;
  assign n42423 = ~n14248 & n16791 ;
  assign n42424 = n42423 ^ n419 ^ 1'b0 ;
  assign n42425 = n3025 | n42424 ;
  assign n42426 = n14306 & ~n42425 ;
  assign n42427 = n17150 & ~n20724 ;
  assign n42428 = n13806 ^ n2917 ^ 1'b0 ;
  assign n42429 = n10885 ^ n10121 ^ 1'b0 ;
  assign n42430 = n42429 ^ n18816 ^ 1'b0 ;
  assign n42431 = n27732 ^ n23891 ^ 1'b0 ;
  assign n42432 = n33947 ^ n23762 ^ n4341 ;
  assign n42433 = n28288 ^ n3158 ^ 1'b0 ;
  assign n42434 = ~n26842 & n42433 ;
  assign n42435 = ~n2539 & n15140 ;
  assign n42436 = ( ~n6583 & n14160 ) | ( ~n6583 & n20303 ) | ( n14160 & n20303 ) ;
  assign n42437 = n42436 ^ n42085 ^ 1'b0 ;
  assign n42438 = n6612 | n8489 ;
  assign n42439 = n42438 ^ n19577 ^ 1'b0 ;
  assign n42440 = ( n2918 & n28414 ) | ( n2918 & ~n42439 ) | ( n28414 & ~n42439 ) ;
  assign n42441 = n74 & ~n2155 ;
  assign n42442 = n4451 | n40081 ;
  assign n42443 = n3698 | n9067 ;
  assign n42444 = ~n229 & n2366 ;
  assign n42445 = n42443 & n42444 ;
  assign n42446 = n2754 & ~n21101 ;
  assign n42447 = n19281 ^ n17981 ^ 1'b0 ;
  assign n42448 = n13272 & n42447 ;
  assign n42449 = n13131 & n42448 ;
  assign n42450 = n42449 ^ n22030 ^ 1'b0 ;
  assign n42451 = ~n22025 & n29788 ;
  assign n42452 = ~n3446 & n34926 ;
  assign n42453 = n30194 & ~n39160 ;
  assign n42454 = n5204 | n6754 ;
  assign n42455 = n42454 ^ n14798 ^ 1'b0 ;
  assign n42456 = n42455 ^ n6397 ^ 1'b0 ;
  assign n42457 = n2350 | n42456 ;
  assign n42458 = n12851 | n18027 ;
  assign n42459 = n29867 ^ n20561 ^ n8911 ;
  assign n42460 = n17836 | n24420 ;
  assign n42461 = n42459 & ~n42460 ;
  assign n42462 = n17378 & ~n24320 ;
  assign n42463 = n37244 | n42462 ;
  assign n42464 = n13996 ^ n8645 ^ 1'b0 ;
  assign n42465 = n41680 & n42464 ;
  assign n42466 = n42465 ^ n33971 ^ 1'b0 ;
  assign n42467 = ~n1635 & n16629 ;
  assign n42468 = ~n2799 & n12845 ;
  assign n42469 = n30856 & ~n42468 ;
  assign n42470 = n5016 & ~n15792 ;
  assign n42471 = n42470 ^ n17778 ^ 1'b0 ;
  assign n42472 = ~n39267 & n42471 ;
  assign n42473 = n11836 & n27622 ;
  assign n42474 = n30471 ^ n9191 ^ 1'b0 ;
  assign n42475 = ~n34156 & n42474 ;
  assign n42476 = n42475 ^ n36992 ^ 1'b0 ;
  assign n42480 = n4559 & ~n6304 ;
  assign n42481 = n7702 | n42480 ;
  assign n42477 = n16067 ^ n7416 ^ 1'b0 ;
  assign n42478 = ~n25706 & n42477 ;
  assign n42479 = n42478 ^ n15710 ^ 1'b0 ;
  assign n42482 = n42481 ^ n42479 ^ n1785 ;
  assign n42483 = n25277 ^ n23749 ^ n2609 ;
  assign n42484 = n14668 ^ n2292 ^ 1'b0 ;
  assign n42485 = n4328 | n42484 ;
  assign n42486 = n42485 ^ n7040 ^ 1'b0 ;
  assign n42487 = ~n32732 & n42486 ;
  assign n42488 = n42487 ^ n34252 ^ 1'b0 ;
  assign n42489 = n42483 | n42488 ;
  assign n42490 = ~n1095 & n18885 ;
  assign n42491 = n42490 ^ n8732 ^ 1'b0 ;
  assign n42492 = ~n13857 & n20543 ;
  assign n42493 = ~n6172 & n13592 ;
  assign n42494 = n31080 & n42493 ;
  assign n42495 = n11975 | n42494 ;
  assign n42496 = n2520 & ~n42495 ;
  assign n42498 = n3411 & n9586 ;
  assign n42499 = ~n3411 & n42498 ;
  assign n42500 = n42499 ^ n4559 ^ 1'b0 ;
  assign n42497 = n2987 | n6467 ;
  assign n42501 = n42500 ^ n42497 ^ 1'b0 ;
  assign n42502 = n10221 & ~n42501 ;
  assign n42503 = n26346 | n31777 ;
  assign n42504 = n41495 & ~n42503 ;
  assign n42505 = ~n23786 & n39848 ;
  assign n42506 = n31747 ^ n23838 ^ 1'b0 ;
  assign n42507 = n11811 & ~n15224 ;
  assign n42508 = ~n10630 & n42507 ;
  assign n42509 = n42048 | n42508 ;
  assign n42510 = n42509 ^ n32900 ^ 1'b0 ;
  assign n42511 = ~n3032 & n20225 ;
  assign n42512 = n6083 & n19933 ;
  assign n42513 = n7512 & ~n42512 ;
  assign n42514 = ~n42511 & n42513 ;
  assign n42515 = n20359 & n24663 ;
  assign n42516 = n7186 & n33950 ;
  assign n42517 = n14279 ^ n5724 ^ 1'b0 ;
  assign n42518 = n26348 & n42517 ;
  assign n42519 = n34422 ^ n18683 ^ 1'b0 ;
  assign n42520 = n21269 & ~n27235 ;
  assign n42521 = n1409 & ~n17717 ;
  assign n42522 = n41425 & n42521 ;
  assign n42523 = ~n10059 & n42522 ;
  assign n42524 = ~n26905 & n42523 ;
  assign n42526 = ~n395 & n6979 ;
  assign n42527 = n42526 ^ n2417 ^ 1'b0 ;
  assign n42528 = n5812 | n42527 ;
  assign n42529 = n42528 ^ n19644 ^ 1'b0 ;
  assign n42525 = n10147 | n25659 ;
  assign n42530 = n42529 ^ n42525 ^ 1'b0 ;
  assign n42531 = n18674 & n36862 ;
  assign n42532 = n7979 & n42531 ;
  assign n42533 = ( n35006 & ~n40655 ) | ( n35006 & n42532 ) | ( ~n40655 & n42532 ) ;
  assign n42534 = n23374 | n30955 ;
  assign n42535 = n19241 & ~n29886 ;
  assign n42537 = n439 & n34412 ;
  assign n42536 = ~n13283 & n24688 ;
  assign n42538 = n42537 ^ n42536 ^ 1'b0 ;
  assign n42541 = n5027 | n30322 ;
  assign n42539 = n1837 & n12937 ;
  assign n42540 = n17692 | n42539 ;
  assign n42542 = n42541 ^ n42540 ^ 1'b0 ;
  assign n42543 = n17 | n42542 ;
  assign n42545 = n1419 | n3250 ;
  assign n42544 = n12337 & n26552 ;
  assign n42546 = n42545 ^ n42544 ^ 1'b0 ;
  assign n42547 = n25660 & ~n42546 ;
  assign n42548 = n30440 ^ n10790 ^ 1'b0 ;
  assign n42549 = n6805 ^ n351 ^ 1'b0 ;
  assign n42550 = n195 | n42549 ;
  assign n42551 = n3105 & ~n31933 ;
  assign n42552 = n42550 & n42551 ;
  assign n42553 = n1219 & n17115 ;
  assign n42554 = n5100 & n42553 ;
  assign n42555 = ~n5953 & n42554 ;
  assign n42556 = ( ~n17737 & n23318 ) | ( ~n17737 & n42555 ) | ( n23318 & n42555 ) ;
  assign n42557 = ~n5677 & n16303 ;
  assign n42558 = ~n11875 & n42557 ;
  assign n42559 = n42558 ^ n5331 ^ n881 ;
  assign n42560 = n11564 ^ n4174 ^ 1'b0 ;
  assign n42561 = n30604 | n42560 ;
  assign n42562 = ~n7917 & n22603 ;
  assign n42563 = ~n8150 & n16359 ;
  assign n42564 = ~n3333 & n33401 ;
  assign n42565 = ~n5116 & n5501 ;
  assign n42566 = n42565 ^ n25316 ^ 1'b0 ;
  assign n42567 = n40343 ^ n27057 ^ 1'b0 ;
  assign n42568 = ~n42566 & n42567 ;
  assign n42569 = ( ~n7792 & n21838 ) | ( ~n7792 & n26961 ) | ( n21838 & n26961 ) ;
  assign n42570 = n27009 ^ n22080 ^ n3502 ;
  assign n42571 = n5569 & n18674 ;
  assign n42577 = n1650 | n7865 ;
  assign n42576 = n1271 | n26317 ;
  assign n42578 = n42577 ^ n42576 ^ 1'b0 ;
  assign n42572 = n3584 & ~n6302 ;
  assign n42573 = ~n10199 & n42572 ;
  assign n42574 = ( n27634 & ~n36757 ) | ( n27634 & n42573 ) | ( ~n36757 & n42573 ) ;
  assign n42575 = n29512 & ~n42574 ;
  assign n42579 = n42578 ^ n42575 ^ 1'b0 ;
  assign n42580 = n15322 & n16249 ;
  assign n42581 = n26828 ^ n1285 ^ 1'b0 ;
  assign n42582 = n365 & n6742 ;
  assign n42583 = ( n2550 & n5084 ) | ( n2550 & n12656 ) | ( n5084 & n12656 ) ;
  assign n42584 = n4632 | n20505 ;
  assign n42585 = n42584 ^ n10716 ^ 1'b0 ;
  assign n42586 = n12576 ^ n1505 ^ 1'b0 ;
  assign n42587 = n42585 | n42586 ;
  assign n42589 = ~n3901 & n6120 ;
  assign n42590 = n12717 & n42589 ;
  assign n42588 = n6589 | n25628 ;
  assign n42591 = n42590 ^ n42588 ^ 1'b0 ;
  assign n42592 = n17683 ^ n2785 ^ 1'b0 ;
  assign n42593 = n1914 & ~n42592 ;
  assign n42594 = n23238 & ~n38172 ;
  assign n42595 = n42594 ^ n11318 ^ 1'b0 ;
  assign n42596 = n6045 & ~n18110 ;
  assign n42597 = ~n3587 & n42596 ;
  assign n42598 = n25101 ^ n6299 ^ 1'b0 ;
  assign n42599 = n42597 | n42598 ;
  assign n42600 = n42599 ^ n19973 ^ n192 ;
  assign n42601 = n15454 ^ n13229 ^ 1'b0 ;
  assign n42602 = n2017 | n42601 ;
  assign n42603 = ~n4626 & n5624 ;
  assign n42604 = n5040 & n42603 ;
  assign n42605 = n29997 & n32977 ;
  assign n42606 = n26727 ^ n6496 ^ 1'b0 ;
  assign n42607 = n2847 & ~n4676 ;
  assign n42608 = n42607 ^ n13122 ^ 1'b0 ;
  assign n42609 = n2885 & n40785 ;
  assign n42610 = n42609 ^ n4741 ^ 1'b0 ;
  assign n42611 = ~n11651 & n12586 ;
  assign n42612 = n42610 & n42611 ;
  assign n42613 = n3909 & ~n29599 ;
  assign n42614 = n42613 ^ n27148 ^ 1'b0 ;
  assign n42615 = n8435 | n9763 ;
  assign n42616 = n42615 ^ n2909 ^ 1'b0 ;
  assign n42617 = n18347 ^ n15078 ^ 1'b0 ;
  assign n42618 = n42616 & n42617 ;
  assign n42619 = n42614 | n42618 ;
  assign n42620 = n5499 & ~n39010 ;
  assign n42621 = n42620 ^ n20810 ^ n11500 ;
  assign n42622 = n2609 & ~n35759 ;
  assign n42623 = ( ~n7599 & n32117 ) | ( ~n7599 & n41399 ) | ( n32117 & n41399 ) ;
  assign n42624 = n3017 | n42623 ;
  assign n42625 = n42624 ^ n2857 ^ 1'b0 ;
  assign n42626 = n1791 & ~n31280 ;
  assign n42627 = n32552 & n42626 ;
  assign n42628 = n6790 ^ n5981 ^ 1'b0 ;
  assign n42629 = n12495 ^ n568 ^ 1'b0 ;
  assign n42630 = n42628 & n42629 ;
  assign n42631 = n301 & n42630 ;
  assign n42632 = n42631 ^ n14152 ^ 1'b0 ;
  assign n42633 = n33898 & n41857 ;
  assign n42634 = ~n40534 & n42633 ;
  assign n42635 = n24407 | n28950 ;
  assign n42636 = ~n11032 & n32730 ;
  assign n42637 = n5058 & ~n17640 ;
  assign n42638 = n18161 | n19072 ;
  assign n42639 = n9560 | n42539 ;
  assign n42640 = n19610 ^ n19153 ^ 1'b0 ;
  assign n42641 = n21649 & ~n42640 ;
  assign n42642 = ~n6297 & n42641 ;
  assign n42643 = n7252 & ~n24694 ;
  assign n42644 = n27894 ^ n21786 ^ 1'b0 ;
  assign n42645 = n4977 & ~n17864 ;
  assign n42646 = ~n42644 & n42645 ;
  assign n42647 = n28399 ^ n20974 ^ 1'b0 ;
  assign n42648 = n91 & n42647 ;
  assign n42649 = n3446 ^ n2891 ^ 1'b0 ;
  assign n42650 = n42648 & n42649 ;
  assign n42651 = n593 & n3279 ;
  assign n42652 = n6526 & ~n11511 ;
  assign n42653 = n42652 ^ n31042 ^ 1'b0 ;
  assign n42654 = n18879 | n42653 ;
  assign n42655 = n9571 & n32226 ;
  assign n42657 = ( n9076 & n15523 ) | ( n9076 & ~n26274 ) | ( n15523 & ~n26274 ) ;
  assign n42656 = ~n261 & n14478 ;
  assign n42658 = n42657 ^ n42656 ^ 1'b0 ;
  assign n42659 = n8363 & n31206 ;
  assign n42660 = n1450 & n42659 ;
  assign n42661 = n25509 ^ n23131 ^ 1'b0 ;
  assign n42662 = ~n13092 & n41818 ;
  assign n42663 = n183 & n42662 ;
  assign n42664 = n5484 | n42663 ;
  assign n42665 = ( n7407 & n8706 ) | ( n7407 & n42664 ) | ( n8706 & n42664 ) ;
  assign n42666 = n42665 ^ n37017 ^ 1'b0 ;
  assign n42667 = n24407 & n42666 ;
  assign n42668 = n543 & ~n5759 ;
  assign n42669 = n42668 ^ n28018 ^ n11945 ;
  assign n42670 = n31214 ^ n4545 ^ 1'b0 ;
  assign n42671 = ~n2455 & n22757 ;
  assign n42672 = ~n9923 & n42671 ;
  assign n42673 = n42672 ^ n30989 ^ 1'b0 ;
  assign n42674 = n8827 & n18900 ;
  assign n42675 = ~n9277 & n13061 ;
  assign n42676 = ~n6280 & n42675 ;
  assign n42677 = ~n17621 & n42676 ;
  assign n42678 = n6006 ^ n3323 ^ n305 ;
  assign n42679 = n22598 ^ n1050 ^ 1'b0 ;
  assign n42680 = n25033 ^ n11714 ^ 1'b0 ;
  assign n42681 = n1083 & ~n1570 ;
  assign n42682 = ( n8683 & ~n14085 ) | ( n8683 & n18151 ) | ( ~n14085 & n18151 ) ;
  assign n42683 = ~n749 & n42682 ;
  assign n42684 = n16313 ^ n9153 ^ 1'b0 ;
  assign n42685 = n6850 & n42684 ;
  assign n42686 = n5637 ^ n1528 ^ 1'b0 ;
  assign n42687 = n42686 ^ n37177 ^ n155 ;
  assign n42688 = ( n6108 & n12082 ) | ( n6108 & ~n17383 ) | ( n12082 & ~n17383 ) ;
  assign n42689 = ( n17105 & ~n21611 ) | ( n17105 & n42688 ) | ( ~n21611 & n42688 ) ;
  assign n42690 = n28902 & ~n36503 ;
  assign n42691 = n7133 & n42690 ;
  assign n42692 = n18040 & n42691 ;
  assign n42693 = ~n42689 & n42692 ;
  assign n42694 = ( ~n12284 & n21786 ) | ( ~n12284 & n42693 ) | ( n21786 & n42693 ) ;
  assign n42695 = n42694 ^ n14830 ^ 1'b0 ;
  assign n42696 = ~n4679 & n13868 ;
  assign n42697 = n42696 ^ n28260 ^ 1'b0 ;
  assign n42698 = ~n8872 & n19983 ;
  assign n42699 = n42698 ^ n27654 ^ 1'b0 ;
  assign n42700 = n5264 | n42699 ;
  assign n42701 = n42700 ^ n30134 ^ 1'b0 ;
  assign n42702 = ~n3252 & n19771 ;
  assign n42703 = n12287 | n18442 ;
  assign n42704 = n42703 ^ n32255 ^ 1'b0 ;
  assign n42705 = n28513 & ~n42704 ;
  assign n42706 = n35186 ^ n1361 ^ 1'b0 ;
  assign n42707 = n42705 & n42706 ;
  assign n42708 = n21775 ^ n4282 ^ 1'b0 ;
  assign n42709 = n4813 | n7856 ;
  assign n42710 = ( n21271 & n42708 ) | ( n21271 & n42709 ) | ( n42708 & n42709 ) ;
  assign n42711 = n9560 & ~n30349 ;
  assign n42712 = n9511 & ~n33009 ;
  assign n42713 = n3319 & n30803 ;
  assign n42714 = n8574 ^ n7804 ^ 1'b0 ;
  assign n42715 = n22342 | n42714 ;
  assign n42716 = n42715 ^ n2940 ^ 1'b0 ;
  assign n42717 = n35248 ^ n29015 ^ 1'b0 ;
  assign n42718 = n2835 | n11636 ;
  assign n42719 = n39763 & ~n42718 ;
  assign n42720 = n26694 ^ n14736 ^ 1'b0 ;
  assign n42721 = n16236 ^ n1235 ^ 1'b0 ;
  assign n42722 = n22789 ^ n8254 ^ 1'b0 ;
  assign n42724 = n7971 ^ n4926 ^ 1'b0 ;
  assign n42725 = n19842 | n42724 ;
  assign n42723 = ~n7576 & n27226 ;
  assign n42726 = n42725 ^ n42723 ^ 1'b0 ;
  assign n42727 = n24516 & ~n34562 ;
  assign n42728 = ~n39402 & n42727 ;
  assign n42729 = n26322 ^ n8639 ^ 1'b0 ;
  assign n42730 = ~n30089 & n42729 ;
  assign n42731 = n901 & ~n42730 ;
  assign n42732 = ~n19170 & n42731 ;
  assign n42733 = n41910 ^ n32948 ^ n6799 ;
  assign n42734 = n12551 ^ n10177 ^ n2588 ;
  assign n42735 = n26987 ^ n16225 ^ 1'b0 ;
  assign n42736 = n3088 & n42735 ;
  assign n42737 = n29975 ^ n25537 ^ n181 ;
  assign n42738 = n37828 ^ n10530 ^ 1'b0 ;
  assign n42739 = n42737 | n42738 ;
  assign n42740 = n6124 | n23230 ;
  assign n42741 = n395 & n39135 ;
  assign n42742 = n15267 & ~n25094 ;
  assign n42744 = x10 & n6498 ;
  assign n42745 = n8928 | n13806 ;
  assign n42746 = ( n8036 & ~n42744 ) | ( n8036 & n42745 ) | ( ~n42744 & n42745 ) ;
  assign n42743 = n16355 | n40917 ;
  assign n42747 = n42746 ^ n42743 ^ 1'b0 ;
  assign n42748 = n34880 ^ n32451 ^ 1'b0 ;
  assign n42749 = n7053 & ~n40433 ;
  assign n42750 = n20374 & n42749 ;
  assign n42751 = n24211 ^ n8287 ^ 1'b0 ;
  assign n42752 = n19709 & n22463 ;
  assign n42755 = ~n11978 & n20127 ;
  assign n42756 = n42755 ^ n35247 ^ 1'b0 ;
  assign n42754 = n6353 ^ n6017 ^ 1'b0 ;
  assign n42753 = ~n1434 & n9290 ;
  assign n42757 = n42756 ^ n42754 ^ n42753 ;
  assign n42758 = n32089 & n32357 ;
  assign n42759 = n3923 | n42758 ;
  assign n42760 = n7948 | n14506 ;
  assign n42761 = ~n2900 & n42760 ;
  assign n42762 = n42439 ^ n26627 ^ 1'b0 ;
  assign n42763 = n28029 & ~n42762 ;
  assign n42764 = n42763 ^ n11971 ^ 1'b0 ;
  assign n42765 = ~n22220 & n42764 ;
  assign n42766 = n8908 & ~n20500 ;
  assign n42767 = n29981 ^ n4470 ^ 1'b0 ;
  assign n42768 = ~n796 & n42767 ;
  assign n42769 = n1325 | n42768 ;
  assign n42770 = n42769 ^ n24998 ^ n14063 ;
  assign n42771 = n1636 & ~n17766 ;
  assign n42772 = n25704 ^ n12575 ^ 1'b0 ;
  assign n42773 = n901 & ~n10178 ;
  assign n42774 = n42773 ^ n7842 ^ 1'b0 ;
  assign n42775 = ( n3817 & n36943 ) | ( n3817 & ~n41011 ) | ( n36943 & ~n41011 ) ;
  assign n42776 = n13021 | n28478 ;
  assign n42777 = n10962 ^ n522 ^ 1'b0 ;
  assign n42778 = n5756 ^ n2577 ^ 1'b0 ;
  assign n42779 = n29827 | n42778 ;
  assign n42780 = n33586 ^ n9163 ^ 1'b0 ;
  assign n42781 = ~n40100 & n42780 ;
  assign n42782 = n1217 & n12201 ;
  assign n42783 = ( n14545 & n14564 ) | ( n14545 & ~n26482 ) | ( n14564 & ~n26482 ) ;
  assign n42784 = n32346 ^ n11324 ^ n1157 ;
  assign n42785 = n42784 ^ n24693 ^ n1714 ;
  assign n42786 = n24007 ^ n6586 ^ 1'b0 ;
  assign n42787 = n18451 ^ n12483 ^ 1'b0 ;
  assign n42788 = ( ~n8084 & n9094 ) | ( ~n8084 & n35936 ) | ( n9094 & n35936 ) ;
  assign n42789 = ~n42787 & n42788 ;
  assign n42790 = n17130 ^ n11599 ^ n3425 ;
  assign n42791 = n31645 ^ n9907 ^ 1'b0 ;
  assign n42792 = n42790 & n42791 ;
  assign n42793 = n29365 ^ n17855 ^ 1'b0 ;
  assign n42794 = n42793 ^ n38 ^ 1'b0 ;
  assign n42795 = n1962 | n42794 ;
  assign n42796 = n42795 ^ n1329 ^ 1'b0 ;
  assign n42797 = n14796 ^ n4097 ^ n2151 ;
  assign n42798 = n42797 ^ n41890 ^ 1'b0 ;
  assign n42799 = n874 ^ n701 ^ 1'b0 ;
  assign n42800 = n28278 | n42799 ;
  assign n42801 = n42800 ^ n18191 ^ 1'b0 ;
  assign n42802 = ~n42798 & n42801 ;
  assign n42803 = n42802 ^ n6514 ^ 1'b0 ;
  assign n42804 = n489 & ~n18486 ;
  assign n42805 = n253 & ~n7921 ;
  assign n42806 = n42805 ^ n1584 ^ 1'b0 ;
  assign n42807 = ~n15773 & n42806 ;
  assign n42808 = n4343 & n42807 ;
  assign n42809 = n42804 | n42808 ;
  assign n42810 = n12145 & ~n26323 ;
  assign n42811 = n2941 & ~n12358 ;
  assign n42812 = n1454 | n29635 ;
  assign n42813 = n42812 ^ n4125 ^ 1'b0 ;
  assign n42814 = n41720 & ~n42813 ;
  assign n42815 = n11324 & n11586 ;
  assign n42816 = n42815 ^ n6429 ^ 1'b0 ;
  assign n42817 = n27488 ^ n24088 ^ n18980 ;
  assign n42818 = n19430 ^ n1769 ^ 1'b0 ;
  assign n42819 = n10183 | n42818 ;
  assign n42820 = n20175 | n42819 ;
  assign n42821 = n10797 ^ n8881 ^ 1'b0 ;
  assign n42822 = n15215 & ~n42821 ;
  assign n42823 = ( n8562 & ~n42820 ) | ( n8562 & n42822 ) | ( ~n42820 & n42822 ) ;
  assign n42824 = n35124 ^ n4993 ^ 1'b0 ;
  assign n42825 = ~n3042 & n42824 ;
  assign n42826 = n7965 | n21440 ;
  assign n42827 = n1363 & ~n2423 ;
  assign n42828 = n28012 & n42827 ;
  assign n42829 = n27923 ^ n13393 ^ 1'b0 ;
  assign n42830 = n16707 | n42829 ;
  assign n42832 = ~n2039 & n6867 ;
  assign n42833 = ~n27620 & n42832 ;
  assign n42831 = ~n17805 & n41154 ;
  assign n42834 = n42833 ^ n42831 ^ 1'b0 ;
  assign n42835 = n155 | n13594 ;
  assign n42836 = ( n9941 & ~n37605 ) | ( n9941 & n42835 ) | ( ~n37605 & n42835 ) ;
  assign n42837 = n11242 & ~n13179 ;
  assign n42838 = ~n9059 & n42837 ;
  assign n42839 = n42838 ^ n2564 ^ 1'b0 ;
  assign n42840 = n2031 | n42839 ;
  assign n42841 = n4372 & ~n42840 ;
  assign n42842 = ~n18307 & n42841 ;
  assign n42843 = n25865 | n35293 ;
  assign n42844 = n42843 ^ n10107 ^ 1'b0 ;
  assign n42845 = ~n16057 & n21981 ;
  assign n42846 = n42845 ^ n9685 ^ 1'b0 ;
  assign n42847 = n565 | n1095 ;
  assign n42848 = n1095 & ~n42847 ;
  assign n42861 = n354 & ~n2835 ;
  assign n42862 = n2835 & n42861 ;
  assign n42849 = n2199 & ~n2730 ;
  assign n42850 = ~n2199 & n42849 ;
  assign n42851 = n2883 & ~n42850 ;
  assign n42852 = n24360 & n42851 ;
  assign n42853 = ~n1750 & n42852 ;
  assign n42854 = n3437 & n42853 ;
  assign n42855 = n10403 & ~n42854 ;
  assign n42856 = ~n10403 & n42855 ;
  assign n42857 = n9096 & ~n42856 ;
  assign n42858 = n42856 & n42857 ;
  assign n42859 = n3097 | n42858 ;
  assign n42860 = n3097 & ~n42859 ;
  assign n42863 = n42862 ^ n42860 ^ 1'b0 ;
  assign n42864 = n7779 | n42863 ;
  assign n42865 = n42848 & ~n42864 ;
  assign n42866 = n848 & ~n1514 ;
  assign n42867 = ~n848 & n42866 ;
  assign n42868 = n23202 | n42867 ;
  assign n42869 = n23202 & ~n42868 ;
  assign n42870 = n42869 ^ n3710 ^ 1'b0 ;
  assign n42871 = n42870 ^ n3121 ^ 1'b0 ;
  assign n42872 = ~n42865 & n42871 ;
  assign n42873 = n9896 | n26987 ;
  assign n42874 = n42873 ^ n2090 ^ 1'b0 ;
  assign n42875 = n14375 & n42874 ;
  assign n42876 = ~n42872 & n42875 ;
  assign n42877 = n2177 | n34857 ;
  assign n42878 = n42876 & ~n42877 ;
  assign n42879 = n10150 & n32328 ;
  assign n42880 = n1230 & n4724 ;
  assign n42881 = n42880 ^ n30497 ^ n2594 ;
  assign n42882 = ( n208 & n3519 ) | ( n208 & n3939 ) | ( n3519 & n3939 ) ;
  assign n42883 = n42882 ^ n34432 ^ n11827 ;
  assign n42884 = n42883 ^ n33632 ^ 1'b0 ;
  assign n42885 = n5031 & n6988 ;
  assign n42886 = n42885 ^ n27222 ^ 1'b0 ;
  assign n42887 = n14246 & n31650 ;
  assign n42888 = ~n3555 & n5811 ;
  assign n42889 = n11268 ^ n8225 ^ 1'b0 ;
  assign n42890 = ~n28501 & n42889 ;
  assign n42891 = n7757 & n23252 ;
  assign n42892 = ( n9321 & ~n22907 ) | ( n9321 & n42891 ) | ( ~n22907 & n42891 ) ;
  assign n42893 = n32177 ^ n6685 ^ 1'b0 ;
  assign n42894 = ~n12211 & n29627 ;
  assign n42895 = n22847 & ~n36961 ;
  assign n42896 = n42894 & n42895 ;
  assign n42897 = n15356 ^ n9118 ^ 1'b0 ;
  assign n42898 = n26496 ^ n12784 ^ 1'b0 ;
  assign n42899 = ~n34803 & n42898 ;
  assign n42900 = n42897 | n42899 ;
  assign n42901 = n8208 & ~n31601 ;
  assign n42902 = ~n33145 & n42901 ;
  assign n42903 = n18037 | n38236 ;
  assign n42904 = n6375 & n9701 ;
  assign n42905 = n30271 ^ n8181 ^ 1'b0 ;
  assign n42906 = n1514 | n42905 ;
  assign n42907 = ~n2353 & n42906 ;
  assign n42908 = n2074 & ~n3052 ;
  assign n42909 = n42908 ^ n13850 ^ 1'b0 ;
  assign n42910 = ( n39001 & n42907 ) | ( n39001 & n42909 ) | ( n42907 & n42909 ) ;
  assign n42911 = n42904 & ~n42910 ;
  assign n42912 = ( n3866 & n17979 ) | ( n3866 & n21836 ) | ( n17979 & n21836 ) ;
  assign n42913 = n19524 ^ n15776 ^ 1'b0 ;
  assign n42914 = n16397 ^ n14896 ^ 1'b0 ;
  assign n42915 = n18303 & n21447 ;
  assign n42916 = n7830 & n8433 ;
  assign n42917 = n18005 & n42916 ;
  assign n42918 = n3715 | n16677 ;
  assign n42919 = n42918 ^ n17178 ^ 1'b0 ;
  assign n42920 = n31721 ^ n11524 ^ 1'b0 ;
  assign n42921 = n21632 ^ n1887 ^ 1'b0 ;
  assign n42922 = n4201 & ~n42921 ;
  assign n42923 = ~n14897 & n42922 ;
  assign n42924 = n5767 & n42923 ;
  assign n42925 = n2723 ^ n517 ^ 1'b0 ;
  assign n42926 = ~n5758 & n23048 ;
  assign n42927 = n42925 & n42926 ;
  assign n42928 = n19647 | n42927 ;
  assign n42929 = n42928 ^ n2930 ^ 1'b0 ;
  assign n42930 = ~n5379 & n7487 ;
  assign n42931 = n42930 ^ n5444 ^ 1'b0 ;
  assign n42932 = n14347 ^ n4180 ^ 1'b0 ;
  assign n42933 = n27238 & n42932 ;
  assign n42934 = n7155 | n10443 ;
  assign n42935 = n42934 ^ n16400 ^ 1'b0 ;
  assign n42936 = n23726 ^ n4201 ^ 1'b0 ;
  assign n42937 = n17319 & ~n42936 ;
  assign n42938 = n1672 | n17330 ;
  assign n42939 = n12932 | n42938 ;
  assign n42940 = n42939 ^ n31050 ^ 1'b0 ;
  assign n42941 = n36927 | n42940 ;
  assign n42942 = n9336 ^ n983 ^ 1'b0 ;
  assign n42943 = ~n2387 & n17481 ;
  assign n42944 = ~n42942 & n42943 ;
  assign n42945 = n20174 | n34937 ;
  assign n42946 = n21929 & ~n42945 ;
  assign n42947 = ~n6325 & n42590 ;
  assign n42948 = n42947 ^ n30107 ^ 1'b0 ;
  assign n42949 = n22394 & n31549 ;
  assign n42951 = n11954 ^ n3081 ^ 1'b0 ;
  assign n42952 = n16920 & ~n29457 ;
  assign n42953 = n42951 & n42952 ;
  assign n42954 = n25849 & n42953 ;
  assign n42955 = n42954 ^ n12058 ^ 1'b0 ;
  assign n42956 = n1995 & ~n42955 ;
  assign n42950 = n11520 | n18989 ;
  assign n42957 = n42956 ^ n42950 ^ n5002 ;
  assign n42958 = n612 & ~n33188 ;
  assign n42959 = ~n30677 & n42958 ;
  assign n42960 = n42959 ^ n33454 ^ 1'b0 ;
  assign n42961 = n42959 & n42960 ;
  assign n42962 = n42961 ^ n11170 ^ 1'b0 ;
  assign n42963 = ~n10890 & n31320 ;
  assign n42964 = n4702 & ~n11589 ;
  assign n42965 = n42964 ^ n3618 ^ 1'b0 ;
  assign n42966 = n42965 ^ n2061 ^ 1'b0 ;
  assign n42967 = ~n450 & n31429 ;
  assign n42968 = n1853 & n22865 ;
  assign n42969 = n273 & ~n20648 ;
  assign n42970 = ~n14031 & n42969 ;
  assign n42971 = n24279 & n42970 ;
  assign n42972 = n42968 & n42971 ;
  assign n42973 = ~n19 & n38371 ;
  assign n42974 = n23491 | n32117 ;
  assign n42975 = n42974 ^ n16164 ^ 1'b0 ;
  assign n42976 = n20015 & n42975 ;
  assign n42977 = n4116 & n42976 ;
  assign n42978 = n42315 ^ n5256 ^ 1'b0 ;
  assign n42979 = n4145 ^ n1327 ^ 1'b0 ;
  assign n42980 = n30543 ^ n11349 ^ 1'b0 ;
  assign n42981 = n42979 | n42980 ;
  assign n42982 = n7690 ^ n4521 ^ 1'b0 ;
  assign n42983 = n42981 & n42982 ;
  assign n42984 = n14716 & n20475 ;
  assign n42985 = n4114 & ~n41965 ;
  assign n42986 = n28610 ^ n3891 ^ 1'b0 ;
  assign n42987 = n19775 & ~n42986 ;
  assign n42988 = n2244 | n17027 ;
  assign n42989 = n4331 & n9336 ;
  assign n42990 = n26647 & n42989 ;
  assign n42991 = ~n30137 & n37613 ;
  assign n42992 = n2643 | n7443 ;
  assign n42993 = ( n13490 & ~n19436 ) | ( n13490 & n33287 ) | ( ~n19436 & n33287 ) ;
  assign n42994 = n42993 ^ n20383 ^ n2902 ;
  assign n42995 = n23790 & n24865 ;
  assign n42996 = n42995 ^ n6941 ^ 1'b0 ;
  assign n42997 = n21324 & n42996 ;
  assign n42998 = ~n905 & n30397 ;
  assign n42999 = n42998 ^ n32210 ^ 1'b0 ;
  assign n43000 = ~n16811 & n42999 ;
  assign n43001 = ~n31242 & n43000 ;
  assign n43002 = n8885 & ~n18544 ;
  assign n43003 = n43002 ^ n9476 ^ 1'b0 ;
  assign n43004 = n43001 | n43003 ;
  assign n43005 = n100 | n23287 ;
  assign n43006 = n43005 ^ n22442 ^ 1'b0 ;
  assign n43007 = n35253 & ~n43006 ;
  assign n43008 = n32121 & ~n39415 ;
  assign n43009 = n147 & n24116 ;
  assign n43010 = n43009 ^ n21714 ^ 1'b0 ;
  assign n43011 = n16929 | n26710 ;
  assign n43012 = n20279 ^ n19900 ^ n423 ;
  assign n43013 = n15206 & ~n19059 ;
  assign n43014 = n21249 & n43013 ;
  assign n43015 = ~n29286 & n37904 ;
  assign n43016 = n1816 ^ n1179 ^ 1'b0 ;
  assign n43017 = n20510 ^ n4095 ^ 1'b0 ;
  assign n43018 = ~n1247 & n28625 ;
  assign n43019 = n43018 ^ n7522 ^ 1'b0 ;
  assign n43020 = ( n11372 & ~n16008 ) | ( n11372 & n43019 ) | ( ~n16008 & n43019 ) ;
  assign n43021 = ( n1865 & n29608 ) | ( n1865 & ~n43020 ) | ( n29608 & ~n43020 ) ;
  assign n43022 = n6619 & ~n13127 ;
  assign n43023 = ~n11742 & n13500 ;
  assign n43024 = n31788 & n37044 ;
  assign n43025 = ~n43023 & n43024 ;
  assign n43026 = ~n15231 & n19942 ;
  assign n43027 = n18790 | n43026 ;
  assign n43028 = n6656 ^ n6570 ^ n2732 ;
  assign n43029 = n43028 ^ n18299 ^ 1'b0 ;
  assign n43030 = n34876 ^ n23705 ^ n11795 ;
  assign n43032 = n12070 & n14276 ;
  assign n43031 = n3518 & ~n9688 ;
  assign n43033 = n43032 ^ n43031 ^ 1'b0 ;
  assign n43034 = n24781 ^ n5443 ^ 1'b0 ;
  assign n43035 = n17391 & n37827 ;
  assign n43036 = ( n4590 & ~n13877 ) | ( n4590 & n20232 ) | ( ~n13877 & n20232 ) ;
  assign n43037 = ~n18883 & n43036 ;
  assign n43038 = n43037 ^ n3334 ^ 1'b0 ;
  assign n43039 = n12813 & ~n28132 ;
  assign n43040 = n43039 ^ n32509 ^ 1'b0 ;
  assign n43041 = n34302 ^ n23150 ^ 1'b0 ;
  assign n43042 = n21 | n43041 ;
  assign n43043 = n17729 & ~n43042 ;
  assign n43044 = ( n18587 & n23318 ) | ( n18587 & ~n27732 ) | ( n23318 & ~n27732 ) ;
  assign n43045 = n6827 & ~n11474 ;
  assign n43046 = n43044 & n43045 ;
  assign n43047 = n37656 ^ n1786 ^ 1'b0 ;
  assign n43048 = n24539 & ~n25081 ;
  assign n43049 = n19216 ^ n5610 ^ 1'b0 ;
  assign n43050 = n43049 ^ n9832 ^ 1'b0 ;
  assign n43051 = n36285 & n38513 ;
  assign n43052 = n43051 ^ n1517 ^ 1'b0 ;
  assign n43053 = n14405 & ~n22215 ;
  assign n43054 = n43053 ^ n34790 ^ 1'b0 ;
  assign n43055 = n40161 & n43054 ;
  assign n43056 = n14750 ^ n3011 ^ 1'b0 ;
  assign n43057 = n15381 | n43056 ;
  assign n43058 = n35596 ^ n23770 ^ n5602 ;
  assign n43059 = n9227 ^ n822 ^ 1'b0 ;
  assign n43060 = n27851 | n43059 ;
  assign n43061 = n43058 | n43060 ;
  assign n43062 = ~n4698 & n17050 ;
  assign n43063 = n43062 ^ n5052 ^ 1'b0 ;
  assign n43064 = ~n30518 & n43063 ;
  assign n43065 = ~n21739 & n43064 ;
  assign n43066 = ~n5963 & n43065 ;
  assign n43067 = n43061 | n43066 ;
  assign n43068 = n18719 & n34253 ;
  assign n43069 = n43068 ^ n38055 ^ 1'b0 ;
  assign n43070 = n13404 & n24313 ;
  assign n43071 = n16513 ^ n1605 ^ 1'b0 ;
  assign n43072 = n3195 ^ n1460 ^ 1'b0 ;
  assign n43073 = ~n33113 & n43072 ;
  assign n43075 = n21418 | n21518 ;
  assign n43076 = n5516 & ~n43075 ;
  assign n43074 = n20153 | n27866 ;
  assign n43077 = n43076 ^ n43074 ^ 1'b0 ;
  assign n43078 = n368 | n1312 ;
  assign n43079 = n43078 ^ n39983 ^ 1'b0 ;
  assign n43080 = ~n182 & n470 ;
  assign n43081 = n43080 ^ n18313 ^ n11619 ;
  assign n43082 = n32940 ^ n17050 ^ n4563 ;
  assign n43084 = ( n2151 & n4901 ) | ( n2151 & n13798 ) | ( n4901 & n13798 ) ;
  assign n43085 = n43084 ^ n17647 ^ 1'b0 ;
  assign n43086 = n2549 & ~n43085 ;
  assign n43087 = n43086 ^ n18516 ^ 1'b0 ;
  assign n43083 = n4216 & ~n27670 ;
  assign n43088 = n43087 ^ n43083 ^ 1'b0 ;
  assign n43089 = n14909 & n29988 ;
  assign n43090 = ~n7174 & n43089 ;
  assign n43091 = n43090 ^ n35710 ^ 1'b0 ;
  assign n43092 = n3598 & n12899 ;
  assign n43093 = n8276 | n13033 ;
  assign n43094 = n43093 ^ n2365 ^ 1'b0 ;
  assign n43095 = n20401 ^ n5636 ^ 1'b0 ;
  assign n43101 = ~n4765 & n21666 ;
  assign n43102 = ~n8408 & n43101 ;
  assign n43096 = n3667 | n6080 ;
  assign n43097 = n43096 ^ n22694 ^ 1'b0 ;
  assign n43098 = n17749 | n43097 ;
  assign n43099 = n43098 ^ n24694 ^ 1'b0 ;
  assign n43100 = ( n8685 & ~n20089 ) | ( n8685 & n43099 ) | ( ~n20089 & n43099 ) ;
  assign n43103 = n43102 ^ n43100 ^ 1'b0 ;
  assign n43104 = n23619 ^ n13879 ^ 1'b0 ;
  assign n43105 = n2309 & n4034 ;
  assign n43106 = ~n31328 & n43105 ;
  assign n43107 = n43106 ^ n26135 ^ 1'b0 ;
  assign n43108 = n37395 ^ n14478 ^ 1'b0 ;
  assign n43113 = n12107 & n14963 ;
  assign n43114 = n43113 ^ n12145 ^ 1'b0 ;
  assign n43115 = ~n12219 & n18389 ;
  assign n43116 = n43114 & n43115 ;
  assign n43109 = n58 & n8773 ;
  assign n43110 = ~n5136 & n43109 ;
  assign n43111 = n2675 | n43110 ;
  assign n43112 = n3445 & ~n43111 ;
  assign n43117 = n43116 ^ n43112 ^ 1'b0 ;
  assign n43120 = ~n1546 & n7735 ;
  assign n43121 = ( ~n14477 & n37627 ) | ( ~n14477 & n43120 ) | ( n37627 & n43120 ) ;
  assign n43118 = n10147 ^ n5080 ^ 1'b0 ;
  assign n43119 = n43118 ^ n4741 ^ n2056 ;
  assign n43122 = n43121 ^ n43119 ^ n910 ;
  assign n43123 = n8445 ^ n983 ^ 1'b0 ;
  assign n43124 = n33632 ^ n24945 ^ 1'b0 ;
  assign n43125 = n43123 & n43124 ;
  assign n43126 = n3573 | n9468 ;
  assign n43127 = n914 & n3172 ;
  assign n43128 = ~n914 & n43127 ;
  assign n43129 = ~n961 & n43128 ;
  assign n43130 = n540 | n3517 ;
  assign n43131 = n540 & ~n43130 ;
  assign n43132 = n1660 & ~n43131 ;
  assign n43133 = n43129 & n43132 ;
  assign n43134 = n4008 & n5155 ;
  assign n43135 = ~n4008 & n43134 ;
  assign n43136 = n36327 & ~n43135 ;
  assign n43137 = ~n36327 & n43136 ;
  assign n43138 = n5028 | n13650 ;
  assign n43139 = n13650 & ~n43138 ;
  assign n43140 = ~n10872 & n43139 ;
  assign n43141 = n43140 ^ n10345 ^ 1'b0 ;
  assign n43142 = n43137 | n43141 ;
  assign n43143 = n43133 | n43142 ;
  assign n43144 = n43126 & ~n43143 ;
  assign n43145 = n43144 ^ n36296 ^ 1'b0 ;
  assign n43147 = n6878 ^ n6011 ^ 1'b0 ;
  assign n43146 = n18392 | n25452 ;
  assign n43148 = n43147 ^ n43146 ^ 1'b0 ;
  assign n43149 = ~n11054 & n13551 ;
  assign n43150 = n43149 ^ n9738 ^ 1'b0 ;
  assign n43151 = ~n4893 & n26360 ;
  assign n43152 = ~n27952 & n43151 ;
  assign n43153 = n5883 ^ n2835 ^ 1'b0 ;
  assign n43154 = n2455 & n43153 ;
  assign n43155 = n43154 ^ n12193 ^ 1'b0 ;
  assign n43156 = n43155 ^ n11827 ^ n6229 ;
  assign n43157 = n21432 & ~n37246 ;
  assign n43158 = ( n12567 & n12641 ) | ( n12567 & n43157 ) | ( n12641 & n43157 ) ;
  assign n43159 = n19397 ^ n7883 ^ n1208 ;
  assign n43160 = n18580 ^ n13 ^ 1'b0 ;
  assign n43161 = n43159 | n43160 ;
  assign n43162 = n12236 | n41006 ;
  assign n43163 = n43162 ^ n4368 ^ 1'b0 ;
  assign n43164 = ~n18380 & n43163 ;
  assign n43165 = n11295 ^ n7138 ^ 1'b0 ;
  assign n43166 = n35738 | n43165 ;
  assign n43167 = n43166 ^ n13668 ^ 1'b0 ;
  assign n43168 = n35839 ^ n7731 ^ 1'b0 ;
  assign n43169 = ~n3820 & n43168 ;
  assign n43170 = n11443 & n14653 ;
  assign n43171 = ~n20923 & n31314 ;
  assign n43172 = n43171 ^ n20143 ^ 1'b0 ;
  assign n43173 = ~n6065 & n43172 ;
  assign n43174 = ~n2041 & n27248 ;
  assign n43175 = n43174 ^ n2833 ^ 1'b0 ;
  assign n43176 = n43175 ^ n3366 ^ 1'b0 ;
  assign n43178 = ~n33802 & n33829 ;
  assign n43179 = n43178 ^ n25484 ^ 1'b0 ;
  assign n43177 = n8555 | n39212 ;
  assign n43180 = n43179 ^ n43177 ^ 1'b0 ;
  assign n43181 = ~n35251 & n43084 ;
  assign n43182 = n8126 & n18324 ;
  assign n43183 = ~n33270 & n43182 ;
  assign n43184 = n6092 | n20730 ;
  assign n43185 = n11296 & n11491 ;
  assign n43186 = n12733 & n39473 ;
  assign n43187 = n11774 | n28157 ;
  assign n43188 = n43187 ^ n31827 ^ 1'b0 ;
  assign n43189 = n42011 ^ n40671 ^ 1'b0 ;
  assign n43190 = n2440 & ~n15390 ;
  assign n43191 = ( ~n3674 & n40064 ) | ( ~n3674 & n43190 ) | ( n40064 & n43190 ) ;
  assign n43192 = ~n20376 & n43191 ;
  assign n43193 = n26711 & n43192 ;
  assign n43194 = n18142 | n21100 ;
  assign n43195 = n11996 & n32327 ;
  assign n43196 = n6498 & ~n16940 ;
  assign n43197 = n13404 & n43196 ;
  assign n43198 = ~n33203 & n43197 ;
  assign n43199 = n5740 | n14901 ;
  assign n43200 = n43198 & ~n43199 ;
  assign n43201 = n24886 ^ n16135 ^ 1'b0 ;
  assign n43202 = n4177 & n43201 ;
  assign n43203 = ( n7694 & n43200 ) | ( n7694 & n43202 ) | ( n43200 & n43202 ) ;
  assign n43204 = n30586 ^ n750 ^ 1'b0 ;
  assign n43205 = ~n23372 & n43204 ;
  assign n43206 = ( n10846 & ~n36380 ) | ( n10846 & n43205 ) | ( ~n36380 & n43205 ) ;
  assign n43207 = n33597 ^ n6511 ^ 1'b0 ;
  assign n43208 = ~n4679 & n25494 ;
  assign n43209 = ~n11515 & n43208 ;
  assign n43210 = n5652 & n18134 ;
  assign n43211 = n43209 & n43210 ;
  assign n43212 = n27593 ^ n9031 ^ 1'b0 ;
  assign n43213 = n37324 & n43212 ;
  assign n43214 = n43213 ^ n3947 ^ 1'b0 ;
  assign n43215 = ~n11827 & n17319 ;
  assign n43216 = n33939 | n43215 ;
  assign n43217 = ~n3061 & n40327 ;
  assign n43218 = n41802 ^ n11356 ^ 1'b0 ;
  assign n43219 = n27527 ^ n26287 ^ n12435 ;
  assign n43220 = ~n489 & n6880 ;
  assign n43221 = ~n1843 & n43220 ;
  assign n43222 = n4687 & ~n18882 ;
  assign n43223 = n7814 | n12436 ;
  assign n43224 = n11006 & n19720 ;
  assign n43225 = n6198 & ~n43224 ;
  assign n43226 = n11295 | n33588 ;
  assign n43227 = n30242 ^ n13891 ^ 1'b0 ;
  assign n43228 = n39183 ^ n35842 ^ 1'b0 ;
  assign n43229 = n17422 & n23325 ;
  assign n43230 = n43229 ^ n12985 ^ 1'b0 ;
  assign n43231 = n4504 & ~n29325 ;
  assign n43232 = n10277 ^ n5606 ^ 1'b0 ;
  assign n43233 = n1182 & ~n43232 ;
  assign n43234 = n9945 ^ n6228 ^ 1'b0 ;
  assign n43235 = n43233 & ~n43234 ;
  assign n43236 = n11819 ^ n10023 ^ 1'b0 ;
  assign n43237 = n42511 ^ n36901 ^ 1'b0 ;
  assign n43238 = ~n10060 & n14672 ;
  assign n43239 = n43238 ^ n40461 ^ n21610 ;
  assign n43240 = n30402 ^ n13181 ^ 1'b0 ;
  assign n43241 = ~n21127 & n43240 ;
  assign n43242 = n13744 ^ n8896 ^ 1'b0 ;
  assign n43243 = n234 & ~n22591 ;
  assign n43244 = n12167 & ~n38760 ;
  assign n43245 = n2771 ^ n1207 ^ 1'b0 ;
  assign n43246 = ( ~n4722 & n31340 ) | ( ~n4722 & n43245 ) | ( n31340 & n43245 ) ;
  assign n43247 = n31793 & ~n43246 ;
  assign n43248 = n42407 ^ n22519 ^ 1'b0 ;
  assign n43249 = n1345 & n18969 ;
  assign n43250 = n28526 ^ n18731 ^ 1'b0 ;
  assign n43251 = n31839 | n32226 ;
  assign n43252 = n13668 & ~n43251 ;
  assign n43253 = n43252 ^ n23348 ^ 1'b0 ;
  assign n43254 = n43250 & ~n43253 ;
  assign n43255 = n11530 ^ n9067 ^ 1'b0 ;
  assign n43256 = n40664 ^ n22866 ^ 1'b0 ;
  assign n43257 = n33468 | n43256 ;
  assign n43258 = n9457 ^ n2042 ^ 1'b0 ;
  assign n43259 = ~n39022 & n43258 ;
  assign n43260 = n41762 ^ n20298 ^ 1'b0 ;
  assign n43261 = n17532 | n27432 ;
  assign n43262 = n43261 ^ n4085 ^ 1'b0 ;
  assign n43263 = n26756 ^ n4784 ^ 1'b0 ;
  assign n43264 = n24624 & n43263 ;
  assign n43265 = n14911 & n20467 ;
  assign n43266 = n3783 & n43265 ;
  assign n43267 = n43266 ^ n3272 ^ 1'b0 ;
  assign n43270 = ( ~n11523 & n17582 ) | ( ~n11523 & n22082 ) | ( n17582 & n22082 ) ;
  assign n43268 = ~n448 & n3292 ;
  assign n43269 = n43268 ^ n24419 ^ 1'b0 ;
  assign n43271 = n43270 ^ n43269 ^ n6749 ;
  assign n43272 = n8930 & n9961 ;
  assign n43273 = n43272 ^ n11170 ^ 1'b0 ;
  assign n43274 = ~n15013 & n43273 ;
  assign n43275 = ~n10015 & n43274 ;
  assign n43276 = n12713 | n17929 ;
  assign n43277 = ~n6748 & n36782 ;
  assign n43278 = n4782 ^ n261 ^ 1'b0 ;
  assign n43279 = ( ~n11668 & n19584 ) | ( ~n11668 & n43278 ) | ( n19584 & n43278 ) ;
  assign n43280 = ~n7696 & n40327 ;
  assign n43281 = ~n21798 & n35240 ;
  assign n43282 = n16693 ^ n1252 ^ 1'b0 ;
  assign n43283 = n688 & n43282 ;
  assign n43284 = n31945 & ~n32898 ;
  assign n43285 = n43284 ^ n7632 ^ 1'b0 ;
  assign n43286 = n7451 & ~n43285 ;
  assign n43287 = ~n2563 & n24217 ;
  assign n43294 = n32582 ^ n1252 ^ 1'b0 ;
  assign n43295 = n58 & ~n43294 ;
  assign n43296 = n43295 ^ n5397 ^ 1'b0 ;
  assign n43288 = ~n1432 & n7358 ;
  assign n43289 = n43288 ^ n5893 ^ 1'b0 ;
  assign n43291 = n9567 & ~n14378 ;
  assign n43290 = ~n6442 & n18413 ;
  assign n43292 = n43291 ^ n43290 ^ 1'b0 ;
  assign n43293 = n43289 & ~n43292 ;
  assign n43297 = n43296 ^ n43293 ^ 1'b0 ;
  assign n43298 = n38913 ^ n707 ^ 1'b0 ;
  assign n43299 = n9924 & ~n43298 ;
  assign n43300 = n24694 | n30803 ;
  assign n43301 = n7314 & ~n42255 ;
  assign n43302 = n19228 ^ n19203 ^ 1'b0 ;
  assign n43303 = n14460 & ~n43302 ;
  assign n43304 = n31272 ^ n22243 ^ 1'b0 ;
  assign n43305 = n39652 | n43304 ;
  assign n43306 = ~n1420 & n32468 ;
  assign n43307 = n20577 & n24264 ;
  assign n43308 = n29748 ^ n13258 ^ 1'b0 ;
  assign n43309 = n492 & ~n43308 ;
  assign n43310 = n43307 | n43309 ;
  assign n43311 = n7943 ^ n2118 ^ 1'b0 ;
  assign n43312 = ~n1622 & n43311 ;
  assign n43313 = n29176 & n43312 ;
  assign n43314 = n43313 ^ n4748 ^ 1'b0 ;
  assign n43315 = n6787 & ~n43314 ;
  assign n43316 = n8817 & n43224 ;
  assign n43317 = n43316 ^ n14481 ^ 1'b0 ;
  assign n43318 = ~n17025 & n43111 ;
  assign n43319 = n43318 ^ n28813 ^ n4547 ;
  assign n43320 = n29136 ^ n11230 ^ 1'b0 ;
  assign n43321 = n7152 | n16888 ;
  assign n43322 = n760 | n43321 ;
  assign n43323 = n30121 | n43322 ;
  assign n43324 = n14448 ^ n13583 ^ 1'b0 ;
  assign n43325 = n17256 ^ n8011 ^ 1'b0 ;
  assign n43326 = n27294 | n43325 ;
  assign n43327 = n10320 & ~n43326 ;
  assign n43328 = n2914 | n30125 ;
  assign n43329 = n43328 ^ n38741 ^ 1'b0 ;
  assign n43330 = n43329 ^ n38095 ^ n29107 ;
  assign n43331 = n6362 | n27447 ;
  assign n43332 = n43331 ^ n11837 ^ 1'b0 ;
  assign n43333 = n1285 & n25389 ;
  assign n43334 = n667 | n10945 ;
  assign n43335 = n34499 & n38268 ;
  assign n43336 = ~n24749 & n43335 ;
  assign n43337 = n19446 ^ x1 ^ 1'b0 ;
  assign n43338 = n43337 ^ n5936 ^ n3946 ;
  assign n43339 = n24809 ^ n6308 ^ 1'b0 ;
  assign n43340 = ~n7285 & n43339 ;
  assign n43341 = n5646 & n10872 ;
  assign n43342 = n43341 ^ n27670 ^ n17936 ;
  assign n43343 = n677 | n2902 ;
  assign n43344 = n30688 & ~n43343 ;
  assign n43345 = n6198 & ~n22164 ;
  assign n43346 = n12219 | n20148 ;
  assign n43347 = n514 & n25233 ;
  assign n43348 = n43347 ^ n10309 ^ 1'b0 ;
  assign n43349 = n13523 ^ n7569 ^ 1'b0 ;
  assign n43350 = n22537 & ~n31199 ;
  assign n43351 = ~n39458 & n43350 ;
  assign n43352 = ~n1173 & n7900 ;
  assign n43353 = n43352 ^ n10723 ^ 1'b0 ;
  assign n43354 = n25467 & ~n43353 ;
  assign n43355 = n21473 ^ n15062 ^ 1'b0 ;
  assign n43356 = n4503 ^ n2848 ^ 1'b0 ;
  assign n43357 = n27782 & ~n33704 ;
  assign n43358 = n11290 & n32594 ;
  assign n43359 = ~n19228 & n43358 ;
  assign n43360 = n8843 | n17695 ;
  assign n43361 = n2179 & ~n43360 ;
  assign n43362 = n34018 ^ n32855 ^ n24065 ;
  assign n43363 = n8499 & n14173 ;
  assign n43364 = n39047 ^ n4838 ^ 1'b0 ;
  assign n43365 = n43363 & ~n43364 ;
  assign n43366 = n6881 ^ n5581 ^ 1'b0 ;
  assign n43367 = ~n36416 & n43366 ;
  assign n43368 = ~n30914 & n43367 ;
  assign n43369 = n11747 & ~n34074 ;
  assign n43370 = ~n22847 & n43369 ;
  assign n43371 = n9311 & ~n22217 ;
  assign n43372 = n23963 ^ n15972 ^ n5872 ;
  assign n43373 = n8807 & n24401 ;
  assign n43374 = n22268 ^ n742 ^ 1'b0 ;
  assign n43375 = n26500 & n31761 ;
  assign n43376 = n3698 | n6651 ;
  assign n43377 = ~n218 & n22587 ;
  assign n43378 = ~n30207 & n43377 ;
  assign n43379 = n452 | n2647 ;
  assign n43380 = n3066 & n3314 ;
  assign n43381 = ~n43379 & n43380 ;
  assign n43382 = n43381 ^ n2562 ^ 1'b0 ;
  assign n43383 = n30711 & n43382 ;
  assign n43384 = n32741 ^ n18333 ^ n16438 ;
  assign n43385 = n6285 | n43384 ;
  assign n43387 = n8823 & ~n18062 ;
  assign n43388 = n43387 ^ n8537 ^ 1'b0 ;
  assign n43386 = n26288 | n43266 ;
  assign n43389 = n43388 ^ n43386 ^ 1'b0 ;
  assign n43390 = ~n479 & n27629 ;
  assign n43391 = n23100 & ~n23889 ;
  assign n43392 = ~n4327 & n22029 ;
  assign n43393 = n1111 | n8785 ;
  assign n43394 = ( n10719 & n16832 ) | ( n10719 & ~n21499 ) | ( n16832 & ~n21499 ) ;
  assign n43395 = n43394 ^ n19677 ^ 1'b0 ;
  assign n43396 = n43062 & ~n43395 ;
  assign n43397 = n14915 ^ n5432 ^ 1'b0 ;
  assign n43398 = ~n31821 & n43397 ;
  assign n43399 = ( ~n5099 & n8227 ) | ( ~n5099 & n43398 ) | ( n8227 & n43398 ) ;
  assign n43400 = n4740 & n18856 ;
  assign n43401 = n43400 ^ n30121 ^ 1'b0 ;
  assign n43402 = n20035 ^ n19367 ^ 1'b0 ;
  assign n43403 = n1723 & n43402 ;
  assign n43404 = n30465 ^ n25783 ^ n1080 ;
  assign n43405 = n22340 & n31472 ;
  assign n43406 = n11791 & n27485 ;
  assign n43407 = n43406 ^ n36302 ^ 1'b0 ;
  assign n43408 = ~n28359 & n35839 ;
  assign n43409 = n43408 ^ n4428 ^ 1'b0 ;
  assign n43410 = n43409 ^ n42670 ^ 1'b0 ;
  assign n43411 = n23273 & ~n43053 ;
  assign n43412 = n43411 ^ n26552 ^ 1'b0 ;
  assign n43413 = ~n16451 & n24720 ;
  assign n43414 = n8258 & n20048 ;
  assign n43415 = n27968 & n38880 ;
  assign n43416 = n33282 ^ n8183 ^ 1'b0 ;
  assign n43417 = n6492 | n25933 ;
  assign n43418 = n12704 & n19995 ;
  assign n43419 = n35889 ^ n8978 ^ n6548 ;
  assign n43420 = n7087 & ~n19914 ;
  assign n43421 = ( n221 & ~n7343 ) | ( n221 & n14649 ) | ( ~n7343 & n14649 ) ;
  assign n43423 = n1004 & n24819 ;
  assign n43424 = n43423 ^ n16150 ^ 1'b0 ;
  assign n43422 = n1918 & ~n20603 ;
  assign n43425 = n43424 ^ n43422 ^ n24220 ;
  assign n43426 = n19321 ^ n1141 ^ 1'b0 ;
  assign n43427 = n6660 | n39428 ;
  assign n43428 = n30030 ^ n2922 ^ 1'b0 ;
  assign n43429 = n38293 & ~n43428 ;
  assign n43430 = n14264 ^ n545 ^ 1'b0 ;
  assign n43431 = n1204 | n43430 ;
  assign n43432 = n16204 ^ n623 ^ 1'b0 ;
  assign n43433 = ~n43431 & n43432 ;
  assign n43434 = n727 | n40802 ;
  assign n43435 = n16726 & ~n30127 ;
  assign n43436 = n43435 ^ n18324 ^ 1'b0 ;
  assign n43437 = n17059 ^ n9886 ^ n5001 ;
  assign n43438 = ~n2615 & n15957 ;
  assign n43439 = n20770 | n41746 ;
  assign n43440 = n20230 & ~n43439 ;
  assign n43442 = n3444 & n8163 ;
  assign n43443 = ~n8163 & n43442 ;
  assign n43444 = ~n5853 & n12401 ;
  assign n43445 = n43443 & n43444 ;
  assign n43446 = n1573 | n42850 ;
  assign n43447 = n1573 & ~n43446 ;
  assign n43448 = n2920 | n7066 ;
  assign n43449 = n43447 & ~n43448 ;
  assign n43450 = n43445 | n43449 ;
  assign n43451 = n43445 & ~n43450 ;
  assign n43441 = n16077 & ~n21496 ;
  assign n43452 = n43451 ^ n43441 ^ 1'b0 ;
  assign n43453 = n1306 & n24800 ;
  assign n43454 = ~n17169 & n43453 ;
  assign n43455 = n43452 & n43454 ;
  assign n43456 = n43455 ^ n765 ^ 1'b0 ;
  assign n43457 = n26200 ^ n5581 ^ n1132 ;
  assign n43458 = ~n16106 & n43457 ;
  assign n43459 = ~n29397 & n43458 ;
  assign n43460 = n3448 | n43459 ;
  assign n43461 = n43460 ^ n18383 ^ 1'b0 ;
  assign n43462 = ~n8600 & n14566 ;
  assign n43463 = n43462 ^ n3229 ^ 1'b0 ;
  assign n43464 = ~n19514 & n43463 ;
  assign n43465 = n24545 | n33880 ;
  assign n43466 = n2924 | n6647 ;
  assign n43467 = n43466 ^ n28148 ^ n13526 ;
  assign n43468 = n20923 ^ n8806 ^ 1'b0 ;
  assign n43469 = n38681 ^ n4097 ^ 1'b0 ;
  assign n43470 = n43468 & n43469 ;
  assign n43471 = ( ~n3649 & n13004 ) | ( ~n3649 & n26612 ) | ( n13004 & n26612 ) ;
  assign n43472 = n43471 ^ n28208 ^ 1'b0 ;
  assign n43473 = n14484 | n18837 ;
  assign n43474 = n17330 & ~n43473 ;
  assign n43475 = n34949 ^ n11137 ^ 1'b0 ;
  assign n43476 = ~n43474 & n43475 ;
  assign n43477 = n973 & n31276 ;
  assign n43478 = ~n20864 & n41652 ;
  assign n43479 = n43478 ^ n15960 ^ 1'b0 ;
  assign n43482 = n43087 ^ n7531 ^ 1'b0 ;
  assign n43483 = n34420 | n43482 ;
  assign n43480 = ( n20157 & n22802 ) | ( n20157 & n32362 ) | ( n22802 & n32362 ) ;
  assign n43481 = n8663 & ~n43480 ;
  assign n43484 = n43483 ^ n43481 ^ 1'b0 ;
  assign n43485 = n43479 & n43484 ;
  assign n43486 = n14651 | n27975 ;
  assign n43487 = n43486 ^ n11770 ^ 1'b0 ;
  assign n43488 = n3637 | n8704 ;
  assign n43489 = n43487 | n43488 ;
  assign n43490 = n37698 ^ n5815 ^ n395 ;
  assign n43491 = n25399 ^ n6020 ^ 1'b0 ;
  assign n43492 = n2781 | n31953 ;
  assign n43493 = n43492 ^ n20600 ^ 1'b0 ;
  assign n43495 = n3418 & ~n9324 ;
  assign n43494 = n120 & ~n459 ;
  assign n43496 = n43495 ^ n43494 ^ 1'b0 ;
  assign n43497 = ~n16807 & n17398 ;
  assign n43498 = n43497 ^ n35323 ^ n25286 ;
  assign n43499 = n2789 ^ n2094 ^ 1'b0 ;
  assign n43500 = ( ~n766 & n15527 ) | ( ~n766 & n43499 ) | ( n15527 & n43499 ) ;
  assign n43501 = n26906 & ~n40696 ;
  assign n43502 = n6876 & n15206 ;
  assign n43503 = n511 & n36311 ;
  assign n43504 = ~n43502 & n43503 ;
  assign n43505 = n18329 & ~n19198 ;
  assign n43506 = ~n34916 & n43505 ;
  assign n43507 = ~n8542 & n38533 ;
  assign n43508 = n2807 | n9546 ;
  assign n43509 = n17294 & ~n43508 ;
  assign n43510 = ~n43312 & n43509 ;
  assign n43511 = n30768 ^ n7147 ^ 1'b0 ;
  assign n43512 = n13520 | n39672 ;
  assign n43513 = n14749 & ~n43512 ;
  assign n43514 = n15532 & ~n36017 ;
  assign n43515 = ( n436 & n2918 ) | ( n436 & n17795 ) | ( n2918 & n17795 ) ;
  assign n43516 = n19443 ^ n10818 ^ 1'b0 ;
  assign n43517 = ~n28244 & n43516 ;
  assign n43518 = n3185 | n16431 ;
  assign n43519 = n43517 | n43518 ;
  assign n43520 = n43515 & n43519 ;
  assign n43521 = ~n43514 & n43520 ;
  assign n43522 = n38181 ^ n19081 ^ n14364 ;
  assign n43523 = n23958 & n39365 ;
  assign n43524 = ~n34643 & n35529 ;
  assign n43525 = ~n11138 & n41635 ;
  assign n43526 = n24973 ^ n23146 ^ 1'b0 ;
  assign n43527 = n7913 & ~n43526 ;
  assign n43528 = ~n3917 & n30072 ;
  assign n43529 = n43528 ^ n13326 ^ 1'b0 ;
  assign n43530 = ~n2565 & n16671 ;
  assign n43531 = ( n21279 & ~n38973 ) | ( n21279 & n43530 ) | ( ~n38973 & n43530 ) ;
  assign n43532 = ( n2784 & ~n9163 ) | ( n2784 & n24565 ) | ( ~n9163 & n24565 ) ;
  assign n43533 = ~n24259 & n43532 ;
  assign n43534 = n19160 ^ n2462 ^ 1'b0 ;
  assign n43535 = n3118 & n43534 ;
  assign n43536 = n11727 ^ n2286 ^ 1'b0 ;
  assign n43537 = n21618 | n43536 ;
  assign n43538 = n21607 | n41023 ;
  assign n43539 = n43537 & ~n43538 ;
  assign n43540 = ~n8580 & n40040 ;
  assign n43541 = n8154 | n43540 ;
  assign n43542 = n874 | n43541 ;
  assign n43543 = n41755 ^ n29138 ^ n6282 ;
  assign n43544 = ~n5020 & n8060 ;
  assign n43545 = n438 & n1265 ;
  assign n43546 = n22135 | n25874 ;
  assign n43547 = n1486 & ~n43546 ;
  assign n43548 = n15578 ^ n2108 ^ 1'b0 ;
  assign n43549 = n29751 ^ n20600 ^ n11102 ;
  assign n43551 = n6081 & n36197 ;
  assign n43550 = n18191 | n36504 ;
  assign n43552 = n43551 ^ n43550 ^ 1'b0 ;
  assign n43553 = ~n1488 & n11812 ;
  assign n43554 = ~n30263 & n43553 ;
  assign n43555 = n1389 & ~n39814 ;
  assign n43556 = ~n3660 & n43555 ;
  assign n43557 = n6205 ^ n2159 ^ 1'b0 ;
  assign n43558 = n11092 | n43557 ;
  assign n43559 = n37237 ^ n16204 ^ 1'b0 ;
  assign n43560 = ~n4833 & n7473 ;
  assign n43561 = n23167 & n43560 ;
  assign n43562 = n1350 | n2798 ;
  assign n43563 = n1208 & n4931 ;
  assign n43564 = n43563 ^ n16947 ^ 1'b0 ;
  assign n43565 = n2505 & n43564 ;
  assign n43566 = n4573 & n10703 ;
  assign n43567 = ~n43565 & n43566 ;
  assign n43568 = n9441 | n18716 ;
  assign n43569 = n43568 ^ n18540 ^ 1'b0 ;
  assign n43570 = n24220 ^ n22041 ^ 1'b0 ;
  assign n43571 = n24372 ^ n1237 ^ 1'b0 ;
  assign n43572 = ~n43570 & n43571 ;
  assign n43573 = n26441 ^ n19489 ^ n5579 ;
  assign n43574 = n42628 ^ n5510 ^ 1'b0 ;
  assign n43575 = n4660 | n10674 ;
  assign n43576 = n43575 ^ n36586 ^ 1'b0 ;
  assign n43577 = n379 & ~n12836 ;
  assign n43578 = n38029 ^ n6029 ^ 1'b0 ;
  assign n43579 = n37335 & n43578 ;
  assign n43580 = n25269 & ~n41019 ;
  assign n43581 = n9294 & n30754 ;
  assign n43582 = ~n4671 & n43581 ;
  assign n43583 = n9795 & n30433 ;
  assign n43584 = n23529 & ~n43583 ;
  assign n43585 = n33853 & n43584 ;
  assign n43586 = n3830 | n8725 ;
  assign n43587 = n43586 ^ n38329 ^ 1'b0 ;
  assign n43588 = ( n7948 & n11144 ) | ( n7948 & n43587 ) | ( n11144 & n43587 ) ;
  assign n43589 = n43059 ^ n11407 ^ 1'b0 ;
  assign n43590 = n6527 & ~n23725 ;
  assign n43591 = ~n5058 & n43590 ;
  assign n43592 = n2338 ^ n344 ^ 1'b0 ;
  assign n43593 = n43591 | n43592 ;
  assign n43594 = n43593 ^ n25926 ^ 1'b0 ;
  assign n43595 = n14530 ^ n4461 ^ 1'b0 ;
  assign n43596 = n35442 ^ n17218 ^ 1'b0 ;
  assign n43597 = n2929 ^ n266 ^ 1'b0 ;
  assign n43598 = n41818 & ~n43597 ;
  assign n43599 = n27113 & ~n38701 ;
  assign n43600 = n26137 & n33746 ;
  assign n43601 = n43600 ^ n31827 ^ n29834 ;
  assign n43602 = n7972 ^ n470 ^ 1'b0 ;
  assign n43603 = ( n16533 & n20909 ) | ( n16533 & n43602 ) | ( n20909 & n43602 ) ;
  assign n43604 = n33033 & n43603 ;
  assign n43605 = n4222 & ~n43604 ;
  assign n43606 = n1469 | n3740 ;
  assign n43607 = n1904 | n43606 ;
  assign n43608 = n1237 & ~n1247 ;
  assign n43609 = n43608 ^ n5630 ^ 1'b0 ;
  assign n43610 = n1237 & ~n25249 ;
  assign n43611 = n43610 ^ n40060 ^ 1'b0 ;
  assign n43612 = n30885 ^ n6832 ^ n1884 ;
  assign n43613 = n8289 & ~n43612 ;
  assign n43614 = n4948 & n43613 ;
  assign n43615 = n3193 | n31389 ;
  assign n43616 = n4137 | n11735 ;
  assign n43617 = n23280 & ~n43616 ;
  assign n43618 = n12107 | n43617 ;
  assign n43619 = n306 & n43618 ;
  assign n43620 = n43619 ^ n18888 ^ 1'b0 ;
  assign n43621 = n16786 | n28311 ;
  assign n43622 = n43621 ^ n2971 ^ n77 ;
  assign n43623 = n14142 & ~n33106 ;
  assign n43624 = n11968 & n43623 ;
  assign n43626 = n8717 & ~n11238 ;
  assign n43627 = n43626 ^ n43126 ^ 1'b0 ;
  assign n43628 = n8610 & ~n43627 ;
  assign n43625 = n38782 ^ n2306 ^ 1'b0 ;
  assign n43629 = n43628 ^ n43625 ^ 1'b0 ;
  assign n43630 = ~n43624 & n43629 ;
  assign n43631 = n32448 ^ n19338 ^ 1'b0 ;
  assign n43632 = n1234 & n12111 ;
  assign n43633 = n43632 ^ n38376 ^ 1'b0 ;
  assign n43634 = n15034 & ~n17927 ;
  assign n43635 = ~n12011 & n43634 ;
  assign n43636 = n43635 ^ n11169 ^ 1'b0 ;
  assign n43637 = n43633 | n43636 ;
  assign n43638 = n7137 | n13111 ;
  assign n43639 = n5938 & ~n16313 ;
  assign n43640 = ~n20223 & n43639 ;
  assign n43641 = ~n1816 & n14963 ;
  assign n43642 = n13934 ^ n13328 ^ 1'b0 ;
  assign n43643 = ~n17172 & n25010 ;
  assign n43644 = ~n20831 & n21109 ;
  assign n43645 = n37540 ^ n36459 ^ 1'b0 ;
  assign n43646 = n181 & ~n39631 ;
  assign n43647 = ~n1978 & n43646 ;
  assign n43648 = n17855 & n38342 ;
  assign n43649 = n43648 ^ n1471 ^ 1'b0 ;
  assign n43650 = n1191 | n43649 ;
  assign n43651 = n32730 ^ n24054 ^ n20299 ;
  assign n43652 = n35248 ^ n7908 ^ n1534 ;
  assign n43653 = n8853 | n27207 ;
  assign n43654 = n6232 | n30464 ;
  assign n43655 = n11685 ^ n10288 ^ n1726 ;
  assign n43656 = n31493 & ~n43655 ;
  assign n43657 = n34405 ^ n270 ^ 1'b0 ;
  assign n43658 = ~n43656 & n43657 ;
  assign n43659 = n22988 & ~n25893 ;
  assign n43660 = n8312 & n14083 ;
  assign n43661 = n7123 ^ n492 ^ 1'b0 ;
  assign n43662 = n17335 & ~n43661 ;
  assign n43663 = ~n16285 & n33169 ;
  assign n43664 = n8107 | n13844 ;
  assign n43665 = n1157 & n10368 ;
  assign n43668 = n6235 ^ n1802 ^ 1'b0 ;
  assign n43669 = n26643 | n43668 ;
  assign n43666 = n11266 ^ n9055 ^ 1'b0 ;
  assign n43667 = n8782 & ~n43666 ;
  assign n43670 = n43669 ^ n43667 ^ 1'b0 ;
  assign n43672 = n5459 & ~n28764 ;
  assign n43673 = n43672 ^ n21207 ^ 1'b0 ;
  assign n43671 = n20249 & n38513 ;
  assign n43674 = n43673 ^ n43671 ^ 1'b0 ;
  assign n43675 = n2587 & ~n2638 ;
  assign n43676 = ~n12972 & n43675 ;
  assign n43677 = n25896 | n43676 ;
  assign n43678 = n3637 & ~n43677 ;
  assign n43679 = n14372 & ~n43678 ;
  assign n43680 = n43679 ^ n13087 ^ 1'b0 ;
  assign n43681 = n11406 & n17195 ;
  assign n43682 = n20010 & ~n43681 ;
  assign n43686 = n2005 | n36958 ;
  assign n43683 = n12189 & ~n14981 ;
  assign n43684 = ( n1546 & n13255 ) | ( n1546 & ~n43683 ) | ( n13255 & ~n43683 ) ;
  assign n43685 = n15250 & n43684 ;
  assign n43687 = n43686 ^ n43685 ^ 1'b0 ;
  assign n43688 = n10277 ^ n2349 ^ 1'b0 ;
  assign n43689 = ~n18867 & n21769 ;
  assign n43690 = n9783 & n16048 ;
  assign n43691 = n10121 & n43690 ;
  assign n43692 = n10580 ^ n2359 ^ 1'b0 ;
  assign n43693 = n8350 & n15087 ;
  assign n43694 = n21091 | n25022 ;
  assign n43695 = n6687 | n43694 ;
  assign n43696 = n32377 & n43695 ;
  assign n43697 = n43696 ^ n35912 ^ 1'b0 ;
  assign n43698 = n1617 & ~n10040 ;
  assign n43699 = n631 & ~n20148 ;
  assign n43700 = n14288 & n43699 ;
  assign n43701 = n34456 | n43700 ;
  assign n43702 = n37485 ^ n10441 ^ n4175 ;
  assign n43703 = ~n7669 & n10327 ;
  assign n43704 = n4191 | n43703 ;
  assign n43705 = n822 | n9029 ;
  assign n43706 = n43705 ^ n2104 ^ 1'b0 ;
  assign n43707 = n8908 & n10476 ;
  assign n43708 = n43707 ^ n8485 ^ 1'b0 ;
  assign n43709 = ~n36559 & n43708 ;
  assign n43710 = n43709 ^ n32451 ^ 1'b0 ;
  assign n43711 = n34901 ^ n15938 ^ 1'b0 ;
  assign n43712 = n8309 | n43711 ;
  assign n43714 = n2376 & n23798 ;
  assign n43713 = n26109 & n29812 ;
  assign n43715 = n43714 ^ n43713 ^ 1'b0 ;
  assign n43716 = n2185 | n30415 ;
  assign n43717 = ~n10481 & n28732 ;
  assign n43718 = n7968 & n8812 ;
  assign n43719 = n43718 ^ n11056 ^ 1'b0 ;
  assign n43720 = n27296 & n43719 ;
  assign n43721 = n24819 | n43720 ;
  assign n43722 = n3896 & ~n15451 ;
  assign n43723 = ~n19116 & n43722 ;
  assign n43724 = n33380 | n43723 ;
  assign n43725 = n4104 | n43724 ;
  assign n43726 = n17490 & ~n17594 ;
  assign n43727 = ~n1078 & n43726 ;
  assign n43729 = ~n4017 & n10298 ;
  assign n43728 = n27579 & ~n31457 ;
  assign n43730 = n43729 ^ n43728 ^ 1'b0 ;
  assign n43731 = n43727 | n43730 ;
  assign n43732 = n16590 ^ n8174 ^ 1'b0 ;
  assign n43733 = ~n20163 & n43732 ;
  assign n43734 = n13692 | n14387 ;
  assign n43735 = n15556 & ~n43734 ;
  assign n43736 = n13529 & ~n43735 ;
  assign n43737 = n23039 ^ n8243 ^ 1'b0 ;
  assign n43738 = ~n40051 & n43737 ;
  assign n43739 = ~n20804 & n31811 ;
  assign n43740 = ~n31733 & n43739 ;
  assign n43742 = n28764 ^ n10131 ^ n8080 ;
  assign n43741 = n6098 & n16734 ;
  assign n43743 = n43742 ^ n43741 ^ 1'b0 ;
  assign n43744 = n11216 ^ n4411 ^ 1'b0 ;
  assign n43745 = n15279 & ~n23125 ;
  assign n43746 = n40639 ^ n30094 ^ 1'b0 ;
  assign n43747 = n8338 & n43746 ;
  assign n43748 = n29276 ^ n20819 ^ 1'b0 ;
  assign n43749 = n2288 & n43748 ;
  assign n43750 = n3216 | n8697 ;
  assign n43751 = n41875 & n43750 ;
  assign n43752 = n9147 | n13639 ;
  assign n43753 = n43752 ^ n31127 ^ 1'b0 ;
  assign n43754 = ~n29148 & n29957 ;
  assign n43755 = n16083 & n43754 ;
  assign n43756 = ( n24454 & n29680 ) | ( n24454 & n43755 ) | ( n29680 & n43755 ) ;
  assign n43757 = n722 & ~n38736 ;
  assign n43758 = n17138 & n17370 ;
  assign n43759 = n22960 ^ n9629 ^ n1469 ;
  assign n43760 = n43759 ^ n35483 ^ 1'b0 ;
  assign n43761 = n43758 & ~n43760 ;
  assign n43762 = n37437 ^ n27174 ^ 1'b0 ;
  assign n43763 = n17491 | n43762 ;
  assign n43764 = ( n5165 & n29100 ) | ( n5165 & ~n40225 ) | ( n29100 & ~n40225 ) ;
  assign n43765 = n22075 & ~n31322 ;
  assign n43766 = n43765 ^ n1033 ^ 1'b0 ;
  assign n43767 = ~n1267 & n6333 ;
  assign n43768 = n43766 & n43767 ;
  assign n43769 = n2914 & ~n8602 ;
  assign n43770 = n43769 ^ n2399 ^ 1'b0 ;
  assign n43771 = n43770 ^ n19330 ^ 1'b0 ;
  assign n43772 = n31648 & n43771 ;
  assign n43773 = n43772 ^ n8308 ^ 1'b0 ;
  assign n43774 = ~n22749 & n23108 ;
  assign n43775 = n43774 ^ n8841 ^ 1'b0 ;
  assign n43776 = n18428 & ~n20842 ;
  assign n43777 = ~n25804 & n35839 ;
  assign n43778 = n43777 ^ n32080 ^ 1'b0 ;
  assign n43779 = ~n216 & n15152 ;
  assign n43780 = ( ~n7570 & n12466 ) | ( ~n7570 & n43779 ) | ( n12466 & n43779 ) ;
  assign n43781 = ( n6734 & n11402 ) | ( n6734 & n43780 ) | ( n11402 & n43780 ) ;
  assign n43782 = n9887 ^ n9372 ^ 1'b0 ;
  assign n43783 = n5093 | n43782 ;
  assign n43784 = n43783 ^ n36309 ^ 1'b0 ;
  assign n43785 = n19172 & n43784 ;
  assign n43786 = n43785 ^ n11164 ^ 1'b0 ;
  assign n43787 = n3088 & ~n13904 ;
  assign n43788 = n10863 ^ n305 ^ 1'b0 ;
  assign n43789 = n21948 | n43788 ;
  assign n43790 = n31590 ^ n3054 ^ 1'b0 ;
  assign n43791 = n6168 | n11076 ;
  assign n43792 = ( ~n11079 & n20242 ) | ( ~n11079 & n42196 ) | ( n20242 & n42196 ) ;
  assign n43793 = ~n5811 & n9253 ;
  assign n43794 = n43793 ^ n26004 ^ 1'b0 ;
  assign n43795 = ~n38505 & n42356 ;
  assign n43796 = ~n3944 & n43795 ;
  assign n43797 = n15112 & ~n43796 ;
  assign n43798 = n4167 & n43797 ;
  assign n43799 = n30922 ^ n19770 ^ 1'b0 ;
  assign n43800 = ~n19548 & n26688 ;
  assign n43801 = n35035 ^ n18598 ^ 1'b0 ;
  assign n43802 = ~n43800 & n43801 ;
  assign n43803 = n15602 ^ n10281 ^ 1'b0 ;
  assign n43804 = n3119 & ~n43803 ;
  assign n43805 = ~n19586 & n35258 ;
  assign n43806 = ~n43804 & n43805 ;
  assign n43807 = n27104 & n40308 ;
  assign n43808 = n30927 & ~n33784 ;
  assign n43809 = ~n13331 & n43808 ;
  assign n43810 = n9087 ^ n8549 ^ n273 ;
  assign n43811 = n14939 ^ n2885 ^ 1'b0 ;
  assign n43812 = n41385 ^ n18958 ^ 1'b0 ;
  assign n43813 = ~n12497 & n43812 ;
  assign n43814 = n43813 ^ n29825 ^ 1'b0 ;
  assign n43815 = n20069 ^ n9899 ^ 1'b0 ;
  assign n43816 = ~n43814 & n43815 ;
  assign n43817 = n43816 ^ n19767 ^ 1'b0 ;
  assign n43818 = n14896 & ~n43817 ;
  assign n43819 = n3564 & ~n4962 ;
  assign n43820 = n43819 ^ n2527 ^ 1'b0 ;
  assign n43821 = ~n36747 & n43462 ;
  assign n43822 = n43821 ^ n27767 ^ 1'b0 ;
  assign n43823 = n29385 | n43822 ;
  assign n43824 = n23179 ^ n15672 ^ 1'b0 ;
  assign n43825 = n30145 & ~n43824 ;
  assign n43826 = n12893 | n20959 ;
  assign n43827 = ~n2576 & n4914 ;
  assign n43828 = n1539 | n35189 ;
  assign n43829 = n34405 ^ n22024 ^ 1'b0 ;
  assign n43830 = n3710 | n30122 ;
  assign n43831 = n15413 & ~n43830 ;
  assign n43832 = n14494 & n31526 ;
  assign n43833 = n30982 ^ n19034 ^ 1'b0 ;
  assign n43834 = n7362 | n7597 ;
  assign n43835 = n43834 ^ n7550 ^ 1'b0 ;
  assign n43836 = n43835 ^ n19182 ^ 1'b0 ;
  assign n43837 = n19359 | n43836 ;
  assign n43838 = n8697 & ~n27334 ;
  assign n43839 = ~n17746 & n43838 ;
  assign n43840 = n36293 & n40019 ;
  assign n43841 = n18757 ^ n18526 ^ 1'b0 ;
  assign n43842 = n438 & ~n2605 ;
  assign n43843 = n2605 & n43842 ;
  assign n43844 = ~n9304 & n15397 ;
  assign n43845 = n43843 & n43844 ;
  assign n43851 = n298 & n500 ;
  assign n43852 = ~n298 & n43851 ;
  assign n43853 = n29854 & ~n43852 ;
  assign n43854 = n43852 & n43853 ;
  assign n43846 = n398 & ~n1337 ;
  assign n43847 = ~n398 & n43846 ;
  assign n43848 = n40 & ~n6035 ;
  assign n43849 = ~n40 & n43848 ;
  assign n43850 = n43847 | n43849 ;
  assign n43855 = n43854 ^ n43850 ^ 1'b0 ;
  assign n43856 = ~n7526 & n43634 ;
  assign n43857 = ~n43634 & n43856 ;
  assign n43858 = n43857 ^ n40603 ^ 1'b0 ;
  assign n43859 = ~n30482 & n43858 ;
  assign n43860 = ( ~n43845 & n43855 ) | ( ~n43845 & n43859 ) | ( n43855 & n43859 ) ;
  assign n43861 = ~n16287 & n16726 ;
  assign n43862 = n17329 | n21318 ;
  assign n43863 = n13205 ^ n2048 ^ 1'b0 ;
  assign n43864 = n8176 | n43863 ;
  assign n43865 = n1216 & n14382 ;
  assign n43866 = n43865 ^ n7597 ^ 1'b0 ;
  assign n43867 = ~n15067 & n29833 ;
  assign n43868 = ~n42684 & n43867 ;
  assign n43869 = n22454 ^ n7532 ^ n4547 ;
  assign n43870 = n2753 | n24423 ;
  assign n43871 = n23845 ^ n16796 ^ 1'b0 ;
  assign n43872 = n31812 ^ n11550 ^ 1'b0 ;
  assign n43873 = n26350 & ~n41792 ;
  assign n43874 = ~n9871 & n43873 ;
  assign n43875 = n8927 & n29652 ;
  assign n43876 = n43875 ^ n24797 ^ 1'b0 ;
  assign n43877 = n35589 ^ n6632 ^ 1'b0 ;
  assign n43878 = n43876 | n43877 ;
  assign n43879 = ~n883 & n32466 ;
  assign n43880 = n15102 | n16142 ;
  assign n43881 = n16142 & ~n43880 ;
  assign n43882 = n43881 ^ n10366 ^ 1'b0 ;
  assign n43883 = n2570 & ~n43882 ;
  assign n43884 = n30775 & n43883 ;
  assign n43885 = n33783 ^ n6330 ^ 1'b0 ;
  assign n43886 = n24180 ^ n593 ^ 1'b0 ;
  assign n43887 = ~n43885 & n43886 ;
  assign n43888 = n1686 | n43887 ;
  assign n43889 = n10430 & ~n32311 ;
  assign n43890 = n1961 | n43889 ;
  assign n43891 = n3257 & ~n26731 ;
  assign n43896 = n31948 ^ n1534 ^ 1'b0 ;
  assign n43895 = n7685 & ~n24326 ;
  assign n43897 = n43896 ^ n43895 ^ 1'b0 ;
  assign n43894 = n21965 ^ n17631 ^ 1'b0 ;
  assign n43892 = n23705 ^ n12047 ^ 1'b0 ;
  assign n43893 = n43892 ^ n28958 ^ n13850 ;
  assign n43898 = n43897 ^ n43894 ^ n43893 ;
  assign n43900 = n1841 & n3539 ;
  assign n43901 = ~n7024 & n43900 ;
  assign n43902 = ~n7030 & n18509 ;
  assign n43903 = n17849 & n43902 ;
  assign n43904 = n43901 | n43903 ;
  assign n43905 = n26604 | n43904 ;
  assign n43906 = n5940 ^ n5332 ^ 1'b0 ;
  assign n43907 = n43905 & ~n43906 ;
  assign n43899 = n10729 & n22186 ;
  assign n43908 = n43907 ^ n43899 ^ 1'b0 ;
  assign n43909 = n368 & n40587 ;
  assign n43910 = n28920 | n42010 ;
  assign n43911 = n1828 | n43910 ;
  assign n43912 = n4590 & n7913 ;
  assign n43913 = n43912 ^ n10610 ^ 1'b0 ;
  assign n43914 = ~n10946 & n43913 ;
  assign n43915 = n12771 ^ n1534 ^ 1'b0 ;
  assign n43916 = n14810 | n31527 ;
  assign n43917 = n43915 | n43916 ;
  assign n43918 = ~n5139 & n17040 ;
  assign n43919 = n20763 ^ n8451 ^ 1'b0 ;
  assign n43920 = ~n43918 & n43919 ;
  assign n43921 = n243 & ~n25623 ;
  assign n43922 = n4461 & n11535 ;
  assign n43923 = n43921 & n43922 ;
  assign n43924 = n18848 ^ n6398 ^ n5215 ;
  assign n43925 = n29980 & n43924 ;
  assign n43926 = n26511 & n43925 ;
  assign n43928 = ~n18945 & n39001 ;
  assign n43929 = ~n24409 & n43928 ;
  assign n43927 = n5569 | n9584 ;
  assign n43930 = n43929 ^ n43927 ^ 1'b0 ;
  assign n43931 = ( n7953 & n15442 ) | ( n7953 & ~n23846 ) | ( n15442 & ~n23846 ) ;
  assign n43932 = n23451 & n24969 ;
  assign n43933 = n13801 & ~n43932 ;
  assign n43934 = n37583 ^ n6387 ^ 1'b0 ;
  assign n43935 = n7312 | n21066 ;
  assign n43936 = n19072 | n43935 ;
  assign n43937 = n14456 & n17816 ;
  assign n43938 = n8404 & n43937 ;
  assign n43939 = n31391 ^ n6417 ^ 1'b0 ;
  assign n43940 = n29635 | n43939 ;
  assign n43942 = n11077 ^ n10403 ^ 1'b0 ;
  assign n43943 = ~n11613 & n43942 ;
  assign n43941 = n11256 ^ n1853 ^ 1'b0 ;
  assign n43944 = n43943 ^ n43941 ^ n22888 ;
  assign n43945 = n9213 & n43944 ;
  assign n43946 = n31515 | n43945 ;
  assign n43947 = n2240 | n7672 ;
  assign n43948 = ~n4767 & n43947 ;
  assign n43949 = n43948 ^ n8879 ^ 1'b0 ;
  assign n43950 = n159 & ~n34931 ;
  assign n43953 = ~n5224 & n6128 ;
  assign n43951 = n8506 | n17227 ;
  assign n43952 = ~n12807 & n43951 ;
  assign n43954 = n43953 ^ n43952 ^ 1'b0 ;
  assign n43955 = n2921 & n22531 ;
  assign n43956 = n43955 ^ n7268 ^ 1'b0 ;
  assign n43957 = n26912 ^ n18540 ^ n8253 ;
  assign n43958 = ~n31068 & n43957 ;
  assign n43959 = n43956 & n43958 ;
  assign n43960 = n15775 & n25231 ;
  assign n43961 = n7176 & ~n7208 ;
  assign n43962 = n5719 & n9284 ;
  assign n43963 = n43962 ^ n4986 ^ 1'b0 ;
  assign n43964 = n23339 & ~n43963 ;
  assign n43965 = n663 & ~n38707 ;
  assign n43966 = n16319 ^ n13393 ^ 1'b0 ;
  assign n43967 = n13702 | n43966 ;
  assign n43968 = n15275 & ~n31905 ;
  assign n43969 = n43968 ^ n21474 ^ 1'b0 ;
  assign n43970 = ( n4928 & ~n15636 ) | ( n4928 & n16237 ) | ( ~n15636 & n16237 ) ;
  assign n43971 = n27819 | n33866 ;
  assign n43972 = n24124 & n43971 ;
  assign n43973 = n43970 & n43972 ;
  assign n43974 = n7384 & ~n7675 ;
  assign n43975 = n43974 ^ n1915 ^ 1'b0 ;
  assign n43976 = n43975 ^ n16768 ^ 1'b0 ;
  assign n43977 = n24875 & n40945 ;
  assign n43978 = n9934 | n43977 ;
  assign n43979 = n8474 ^ n4158 ^ 1'b0 ;
  assign n43980 = ~n2474 & n43979 ;
  assign n43981 = n468 & n43980 ;
  assign n43982 = n11849 & n43981 ;
  assign n43983 = n15508 & ~n20302 ;
  assign n43984 = ( ~n5903 & n16675 ) | ( ~n5903 & n18929 ) | ( n16675 & n18929 ) ;
  assign n43985 = n15171 | n17622 ;
  assign n43986 = n43984 | n43985 ;
  assign n43987 = n10505 ^ n52 ^ 1'b0 ;
  assign n43988 = ~n20835 & n43987 ;
  assign n43989 = ~n38824 & n43988 ;
  assign n43991 = n15966 ^ n4088 ^ 1'b0 ;
  assign n43990 = ~n6883 & n24774 ;
  assign n43992 = n43991 ^ n43990 ^ 1'b0 ;
  assign n43993 = ( n22513 & ~n28043 ) | ( n22513 & n43992 ) | ( ~n28043 & n43992 ) ;
  assign n43994 = n6142 | n23484 ;
  assign n43995 = n43994 ^ n7936 ^ 1'b0 ;
  assign n43996 = n18648 & ~n31187 ;
  assign n43997 = n22051 ^ n12242 ^ n3347 ;
  assign n43998 = ~n19668 & n43997 ;
  assign n43999 = n326 | n17935 ;
  assign n44000 = n43999 ^ n11220 ^ n1806 ;
  assign n44001 = ~n19466 & n44000 ;
  assign n44002 = n41767 & n44001 ;
  assign n44004 = ~n14368 & n18426 ;
  assign n44003 = n11046 & ~n29831 ;
  assign n44005 = n44004 ^ n44003 ^ 1'b0 ;
  assign n44006 = ~n1098 & n10038 ;
  assign n44007 = n873 & ~n5438 ;
  assign n44008 = ~n12563 & n44007 ;
  assign n44012 = n9072 & ~n9287 ;
  assign n44013 = ~n7067 & n44012 ;
  assign n44014 = n8308 & ~n21496 ;
  assign n44015 = n44013 & n44014 ;
  assign n44009 = ~n7531 & n32498 ;
  assign n44010 = n24957 | n44009 ;
  assign n44011 = n22206 | n44010 ;
  assign n44016 = n44015 ^ n44011 ^ 1'b0 ;
  assign n44017 = n29727 ^ n16527 ^ 1'b0 ;
  assign n44018 = n682 | n30215 ;
  assign n44019 = n15804 & ~n16880 ;
  assign n44020 = n44019 ^ n10338 ^ 1'b0 ;
  assign n44021 = n44020 ^ n21675 ^ 1'b0 ;
  assign n44022 = ~n30908 & n33206 ;
  assign n44023 = n7036 & ~n10519 ;
  assign n44024 = ~n6444 & n44023 ;
  assign n44025 = n23621 ^ n3980 ^ 1'b0 ;
  assign n44026 = ~n6674 & n44025 ;
  assign n44027 = n19006 ^ n7859 ^ 1'b0 ;
  assign n44028 = ~n31309 & n44027 ;
  assign n44029 = n2040 & n6999 ;
  assign n44030 = n4627 & n44029 ;
  assign n44031 = ( n36357 & n42162 ) | ( n36357 & ~n44030 ) | ( n42162 & ~n44030 ) ;
  assign n44032 = n39247 ^ n8752 ^ 1'b0 ;
  assign n44033 = n14959 & ~n27498 ;
  assign n44034 = ~n27966 & n44033 ;
  assign n44035 = n34788 | n42686 ;
  assign n44036 = n10760 & ~n13971 ;
  assign n44037 = n44035 & n44036 ;
  assign n44038 = n3353 ^ n2796 ^ 1'b0 ;
  assign n44039 = n44038 ^ n30029 ^ 1'b0 ;
  assign n44040 = n28589 & ~n44039 ;
  assign n44041 = ~n1083 & n19249 ;
  assign n44042 = ~n16552 & n17099 ;
  assign n44043 = n44042 ^ n366 ^ 1'b0 ;
  assign n44044 = ~n1398 & n44043 ;
  assign n44045 = ~n32216 & n44044 ;
  assign n44046 = n44045 ^ n40457 ^ 1'b0 ;
  assign n44047 = ( n12994 & n18053 ) | ( n12994 & n32384 ) | ( n18053 & n32384 ) ;
  assign n44048 = n2940 ^ n1462 ^ 1'b0 ;
  assign n44049 = n44047 | n44048 ;
  assign n44050 = n813 & n10767 ;
  assign n44051 = n44050 ^ n12373 ^ 1'b0 ;
  assign n44052 = n1182 | n14916 ;
  assign n44053 = n37142 ^ n2619 ^ 1'b0 ;
  assign n44054 = n12815 & ~n27400 ;
  assign n44055 = ~n1596 & n16004 ;
  assign n44056 = n22566 & n44055 ;
  assign n44057 = n44056 ^ n2306 ^ n820 ;
  assign n44058 = ~n18277 & n24986 ;
  assign n44059 = ~n3512 & n15385 ;
  assign n44060 = n8512 & n44059 ;
  assign n44061 = n22044 | n44060 ;
  assign n44062 = n29397 ^ n22451 ^ 1'b0 ;
  assign n44063 = n44061 & ~n44062 ;
  assign n44064 = n19218 & ~n32968 ;
  assign n44065 = n19821 ^ n3725 ^ 1'b0 ;
  assign n44066 = n23504 | n44065 ;
  assign n44067 = n44066 ^ n27148 ^ 1'b0 ;
  assign n44068 = ( n7556 & n8436 ) | ( n7556 & n11013 ) | ( n8436 & n11013 ) ;
  assign n44069 = n44068 ^ n27498 ^ 1'b0 ;
  assign n44070 = n37135 & n44069 ;
  assign n44071 = n15105 ^ n10092 ^ 1'b0 ;
  assign n44072 = ~n9928 & n44071 ;
  assign n44073 = n5235 & n21432 ;
  assign n44074 = n2857 & n44073 ;
  assign n44075 = n13124 | n44074 ;
  assign n44076 = n44075 ^ n3564 ^ 1'b0 ;
  assign n44077 = n44076 ^ n608 ^ 1'b0 ;
  assign n44078 = n6322 & n27843 ;
  assign n44079 = n1570 & n44078 ;
  assign n44080 = n6617 ^ n5007 ^ 1'b0 ;
  assign n44081 = n744 & ~n44080 ;
  assign n44082 = ~n11098 & n37001 ;
  assign n44083 = n1271 | n44082 ;
  assign n44084 = n44083 ^ n1971 ^ 1'b0 ;
  assign n44085 = n37222 ^ n13557 ^ 1'b0 ;
  assign n44087 = ~n6852 & n21952 ;
  assign n44086 = ~n2401 & n41322 ;
  assign n44088 = n44087 ^ n44086 ^ 1'b0 ;
  assign n44089 = n13335 & n33885 ;
  assign n44090 = n5811 ^ n1346 ^ 1'b0 ;
  assign n44091 = ~n4103 & n24324 ;
  assign n44092 = n33755 ^ n23099 ^ n14676 ;
  assign n44093 = ~n23981 & n30897 ;
  assign n44094 = n2850 & ~n29279 ;
  assign n44095 = n5316 | n5417 ;
  assign n44096 = ~n5458 & n24543 ;
  assign n44097 = n42788 ^ n16810 ^ 1'b0 ;
  assign n44098 = n11940 & n44097 ;
  assign n44099 = n2481 ^ n2282 ^ 1'b0 ;
  assign n44100 = n6573 & n44099 ;
  assign n44101 = n26123 ^ n23367 ^ 1'b0 ;
  assign n44102 = n30605 & ~n44101 ;
  assign n44103 = ~n17189 & n44102 ;
  assign n44104 = n5758 ^ n1191 ^ 1'b0 ;
  assign n44105 = n23566 ^ n23084 ^ 1'b0 ;
  assign n44106 = ~n38276 & n44105 ;
  assign n44107 = n13223 ^ n11969 ^ 1'b0 ;
  assign n44108 = n41791 | n44107 ;
  assign n44109 = n10194 | n32864 ;
  assign n44110 = x6 | n15049 ;
  assign n44111 = n7596 | n36155 ;
  assign n44112 = n44111 ^ n33829 ^ 1'b0 ;
  assign n44113 = n27411 ^ n25892 ^ n12213 ;
  assign n44114 = ( n24897 & n25731 ) | ( n24897 & ~n38766 ) | ( n25731 & ~n38766 ) ;
  assign n44115 = n697 | n9287 ;
  assign n44116 = n44115 ^ n8884 ^ 1'b0 ;
  assign n44117 = n18042 & ~n18919 ;
  assign n44118 = n5958 | n9572 ;
  assign n44119 = n9572 & ~n44118 ;
  assign n44120 = n7430 & n44119 ;
  assign n44121 = n15906 | n44120 ;
  assign n44122 = n15906 & ~n44121 ;
  assign n44139 = ~n11025 & n26816 ;
  assign n44140 = ~n13238 & n44139 ;
  assign n44141 = n13238 & n44140 ;
  assign n44123 = n938 | n1040 ;
  assign n44124 = n938 & ~n44123 ;
  assign n44125 = n1927 & ~n44124 ;
  assign n44126 = n44124 & n44125 ;
  assign n44127 = n47 | n700 ;
  assign n44128 = n700 & ~n44127 ;
  assign n44129 = n44128 ^ n1912 ^ 1'b0 ;
  assign n44130 = n44129 ^ n1912 ^ 1'b0 ;
  assign n44131 = ~n1164 & n44130 ;
  assign n44132 = n723 & n1351 ;
  assign n44133 = ~n1351 & n44132 ;
  assign n44134 = n44133 ^ n2061 ^ 1'b0 ;
  assign n44135 = n44131 & ~n44134 ;
  assign n44136 = ~n44126 & n44135 ;
  assign n44137 = n44126 & n44136 ;
  assign n44138 = ~n1167 & n44137 ;
  assign n44142 = n44141 ^ n44138 ^ 1'b0 ;
  assign n44143 = ~n44122 & n44142 ;
  assign n44153 = ~n11230 & n18595 ;
  assign n44154 = ~n18595 & n44153 ;
  assign n44155 = ~n1240 & n3367 ;
  assign n44156 = n1240 & n44155 ;
  assign n44157 = n44154 | n44156 ;
  assign n44158 = n44154 & ~n44157 ;
  assign n44159 = n32025 & ~n44158 ;
  assign n44144 = n253 & n1978 ;
  assign n44145 = ~n253 & n44144 ;
  assign n44146 = n149 | n44145 ;
  assign n44147 = n44145 & ~n44146 ;
  assign n44148 = n13612 & ~n44147 ;
  assign n44149 = n1132 & ~n42848 ;
  assign n44150 = n42848 & n44149 ;
  assign n44151 = n15616 | n44150 ;
  assign n44152 = ( ~n1939 & n44148 ) | ( ~n1939 & n44151 ) | ( n44148 & n44151 ) ;
  assign n44160 = n44159 ^ n44152 ^ 1'b0 ;
  assign n44161 = n44143 & n44160 ;
  assign n44162 = ~n4648 & n44161 ;
  assign n44163 = n8122 | n12444 ;
  assign n44164 = n44162 | n44163 ;
  assign n44165 = n27751 | n38889 ;
  assign n44166 = n6216 & ~n44165 ;
  assign n44167 = n3619 & n23451 ;
  assign n44168 = n9821 ^ n4372 ^ 1'b0 ;
  assign n44169 = n2728 | n44168 ;
  assign n44170 = ~n31510 & n36056 ;
  assign n44171 = n3543 & n19463 ;
  assign n44172 = n21048 ^ n19356 ^ 1'b0 ;
  assign n44173 = n16825 | n44172 ;
  assign n44174 = n44171 | n44173 ;
  assign n44175 = n14913 & n44174 ;
  assign n44176 = n14240 ^ n7531 ^ 1'b0 ;
  assign n44177 = n5901 & ~n6637 ;
  assign n44178 = n44176 & n44177 ;
  assign n44179 = n23948 ^ n4137 ^ 1'b0 ;
  assign n44180 = n11411 & n17353 ;
  assign n44181 = ~n8440 & n21649 ;
  assign n44182 = n44181 ^ n19792 ^ 1'b0 ;
  assign n44183 = n39237 | n44182 ;
  assign n44184 = n44183 ^ n12831 ^ 1'b0 ;
  assign n44185 = n19363 & ~n40230 ;
  assign n44186 = n26212 ^ n11046 ^ 1'b0 ;
  assign n44187 = ~n44185 & n44186 ;
  assign n44188 = n27585 | n44187 ;
  assign n44189 = n13979 ^ n2843 ^ 1'b0 ;
  assign n44190 = n5967 | n44189 ;
  assign n44191 = n25719 ^ n23670 ^ 1'b0 ;
  assign n44192 = n3221 | n44191 ;
  assign n44193 = n2655 & ~n44192 ;
  assign n44194 = n10976 & n44193 ;
  assign n44195 = n44194 ^ n1337 ^ 1'b0 ;
  assign n44196 = n21303 ^ n20919 ^ n12788 ;
  assign n44198 = n16744 ^ n3471 ^ n3186 ;
  assign n44197 = n25972 ^ n14691 ^ 1'b0 ;
  assign n44199 = n44198 ^ n44197 ^ 1'b0 ;
  assign n44200 = ~n13875 & n23812 ;
  assign n44201 = n1688 | n20828 ;
  assign n44202 = n44201 ^ n7087 ^ 1'b0 ;
  assign n44203 = n2134 & ~n44202 ;
  assign n44204 = n16795 & ~n44203 ;
  assign n44205 = n18853 & n44204 ;
  assign n44206 = n510 ^ n235 ^ 1'b0 ;
  assign n44207 = n10603 & ~n29763 ;
  assign n44208 = n44207 ^ n14793 ^ 1'b0 ;
  assign n44210 = n11640 & n18348 ;
  assign n44211 = n44210 ^ n11772 ^ 1'b0 ;
  assign n44209 = n11032 | n12897 ;
  assign n44212 = n44211 ^ n44209 ^ 1'b0 ;
  assign n44213 = n44212 ^ n14555 ^ 1'b0 ;
  assign n44214 = n44213 ^ n19514 ^ 1'b0 ;
  assign n44215 = n22095 ^ n7963 ^ 1'b0 ;
  assign n44216 = n6813 & ~n44215 ;
  assign n44217 = ~n29447 & n44216 ;
  assign n44219 = n14038 & n41816 ;
  assign n44218 = n11118 ^ n4313 ^ 1'b0 ;
  assign n44220 = n44219 ^ n44218 ^ 1'b0 ;
  assign n44221 = n19978 ^ n19304 ^ 1'b0 ;
  assign n44222 = n25701 & n44221 ;
  assign n44223 = n22781 ^ n17177 ^ 1'b0 ;
  assign n44224 = n4455 & n12082 ;
  assign n44225 = n44224 ^ n35642 ^ 1'b0 ;
  assign n44226 = ~n11552 & n38447 ;
  assign n44227 = ~n44225 & n44226 ;
  assign n44228 = n27435 | n44227 ;
  assign n44229 = n5420 & n28867 ;
  assign n44230 = n44229 ^ n16582 ^ 1'b0 ;
  assign n44231 = n43617 ^ n16414 ^ n4731 ;
  assign n44232 = n38692 & ~n44231 ;
  assign n44233 = n8012 & n44232 ;
  assign n44234 = n44233 ^ n27218 ^ n3548 ;
  assign n44235 = ~n3919 & n41630 ;
  assign n44236 = n3531 | n44235 ;
  assign n44240 = n19561 & n32208 ;
  assign n44241 = n44240 ^ n9926 ^ 1'b0 ;
  assign n44237 = n18740 | n23699 ;
  assign n44238 = n11190 & n44237 ;
  assign n44239 = n18963 & n44238 ;
  assign n44242 = n44241 ^ n44239 ^ n21597 ;
  assign n44243 = n35589 ^ n32039 ^ n31234 ;
  assign n44244 = n19498 ^ n17113 ^ 1'b0 ;
  assign n44245 = n25540 & ~n44227 ;
  assign n44246 = n1700 & n27310 ;
  assign n44247 = n7482 & n44246 ;
  assign n44248 = n3541 & n44247 ;
  assign n44249 = n32260 ^ n17070 ^ n4531 ;
  assign n44250 = ~n9585 & n44249 ;
  assign n44251 = n44248 & n44250 ;
  assign n44252 = n4917 & n14317 ;
  assign n44253 = n44252 ^ n38181 ^ 1'b0 ;
  assign n44254 = n14160 ^ n3390 ^ 1'b0 ;
  assign n44255 = n7350 & ~n27366 ;
  assign n44256 = n44255 ^ n33763 ^ 1'b0 ;
  assign n44257 = n173 | n6485 ;
  assign n44258 = n11162 | n44257 ;
  assign n44259 = ~n8278 & n44258 ;
  assign n44261 = n11964 ^ n2101 ^ 1'b0 ;
  assign n44260 = n2478 | n12775 ;
  assign n44262 = n44261 ^ n44260 ^ 1'b0 ;
  assign n44263 = n44262 ^ n13252 ^ 1'b0 ;
  assign n44264 = n3235 & ~n29328 ;
  assign n44265 = n26958 ^ n4486 ^ 1'b0 ;
  assign n44266 = ( n14274 & n39912 ) | ( n14274 & n44265 ) | ( n39912 & n44265 ) ;
  assign n44267 = n44266 ^ n2094 ^ 1'b0 ;
  assign n44268 = n9660 & n26522 ;
  assign n44269 = n44268 ^ n43644 ^ 1'b0 ;
  assign n44271 = n8190 | n28764 ;
  assign n44270 = n3611 & ~n10601 ;
  assign n44272 = n44271 ^ n44270 ^ 1'b0 ;
  assign n44273 = n44272 ^ n27 ^ 1'b0 ;
  assign n44274 = n15018 & n20924 ;
  assign n44275 = n3152 & ~n4505 ;
  assign n44276 = n2256 & n44275 ;
  assign n44277 = n44276 ^ n19915 ^ 1'b0 ;
  assign n44278 = n35699 ^ n5793 ^ 1'b0 ;
  assign n44279 = ~n1261 & n44278 ;
  assign n44280 = n1176 & n44279 ;
  assign n44281 = n28749 ^ n26291 ^ n2185 ;
  assign n44282 = n6898 & n44281 ;
  assign n44283 = n31125 & n31958 ;
  assign n44284 = ~n28742 & n44283 ;
  assign n44285 = n40797 ^ n11498 ^ n7325 ;
  assign n44286 = ( n2145 & ~n26690 ) | ( n2145 & n35505 ) | ( ~n26690 & n35505 ) ;
  assign n44287 = ~n5311 & n44286 ;
  assign n44288 = ~n9210 & n44287 ;
  assign n44289 = n8138 ^ n5501 ^ 1'b0 ;
  assign n44290 = n16549 & ~n44289 ;
  assign n44291 = n31777 | n44290 ;
  assign n44295 = n7023 ^ n3003 ^ 1'b0 ;
  assign n44292 = n4559 | n16912 ;
  assign n44293 = n23714 & ~n44292 ;
  assign n44294 = n8147 & ~n44293 ;
  assign n44296 = n44295 ^ n44294 ^ 1'b0 ;
  assign n44297 = n24146 ^ n4040 ^ 1'b0 ;
  assign n44298 = n7463 & ~n9992 ;
  assign n44299 = n1538 | n2856 ;
  assign n44300 = n44299 ^ n1771 ^ 1'b0 ;
  assign n44301 = n34730 ^ n19821 ^ 1'b0 ;
  assign n44302 = ~n44300 & n44301 ;
  assign n44303 = n5041 | n17295 ;
  assign n44304 = n4593 | n23028 ;
  assign n44305 = n9405 | n44304 ;
  assign n44306 = n44305 ^ n37054 ^ 1'b0 ;
  assign n44307 = n19671 | n35894 ;
  assign n44308 = ~n14808 & n40074 ;
  assign n44309 = n5708 & ~n33322 ;
  assign n44310 = n44309 ^ n6526 ^ 1'b0 ;
  assign n44311 = ( n2193 & ~n30374 ) | ( n2193 & n44310 ) | ( ~n30374 & n44310 ) ;
  assign n44312 = n27219 ^ n18234 ^ 1'b0 ;
  assign n44313 = n31141 ^ n18393 ^ 1'b0 ;
  assign n44314 = n3794 & n31289 ;
  assign n44315 = n44314 ^ n6719 ^ 1'b0 ;
  assign n44316 = n553 | n7159 ;
  assign n44317 = n44316 ^ n35825 ^ 1'b0 ;
  assign n44318 = n38279 ^ n14546 ^ n13855 ;
  assign n44319 = n15826 & n37115 ;
  assign n44320 = n6997 | n13179 ;
  assign n44321 = n7616 & ~n40908 ;
  assign n44322 = ~n43531 & n44321 ;
  assign n44323 = n2131 ^ n961 ^ 1'b0 ;
  assign n44327 = n2666 | n22941 ;
  assign n44324 = n505 & ~n11390 ;
  assign n44325 = ~n2225 & n44324 ;
  assign n44326 = n21594 | n44325 ;
  assign n44328 = n44327 ^ n44326 ^ n36876 ;
  assign n44329 = n2313 & n5797 ;
  assign n44330 = n44329 ^ n20021 ^ 1'b0 ;
  assign n44331 = n11099 & n18111 ;
  assign n44332 = n1081 & n37625 ;
  assign n44333 = ~n6350 & n44332 ;
  assign n44334 = n19564 & ~n44333 ;
  assign n44335 = n11691 ^ n1700 ^ 1'b0 ;
  assign n44336 = n18624 & ~n37010 ;
  assign n44337 = n1539 & n44336 ;
  assign n44338 = n8868 & ~n20000 ;
  assign n44339 = n33389 ^ n10324 ^ n7966 ;
  assign n44340 = n1929 & n11296 ;
  assign n44341 = n13723 & n44340 ;
  assign n44342 = n9282 | n44341 ;
  assign n44343 = n44342 ^ n5431 ^ 1'b0 ;
  assign n44344 = n14484 & n43686 ;
  assign n44345 = ~n8700 & n21843 ;
  assign n44346 = ~n41393 & n44345 ;
  assign n44347 = n5450 & n44346 ;
  assign n44348 = n11423 ^ n8803 ^ n6042 ;
  assign n44349 = ~n14563 & n44348 ;
  assign n44350 = n19245 & n44349 ;
  assign n44351 = n29642 & n44350 ;
  assign n44352 = ~n5866 & n8154 ;
  assign n44353 = n4085 & n29562 ;
  assign n44354 = n23738 & n44353 ;
  assign n44355 = n5431 & ~n17682 ;
  assign n44356 = n44355 ^ n44181 ^ 1'b0 ;
  assign n44357 = n44356 ^ n28255 ^ n26786 ;
  assign n44358 = n28137 ^ n6825 ^ n828 ;
  assign n44359 = n44358 ^ n38901 ^ n18945 ;
  assign n44360 = n21315 & n29655 ;
  assign n44361 = n5471 & ~n7836 ;
  assign n44365 = n194 & ~n3363 ;
  assign n44362 = n21080 ^ n7759 ^ 1'b0 ;
  assign n44363 = n30258 | n44362 ;
  assign n44364 = n19160 & ~n44363 ;
  assign n44366 = n44365 ^ n44364 ^ 1'b0 ;
  assign n44367 = n23854 & ~n36357 ;
  assign n44368 = n33285 ^ n16900 ^ n4621 ;
  assign n44369 = n40970 ^ n25599 ^ 1'b0 ;
  assign n44370 = n600 & ~n6494 ;
  assign n44371 = n6494 & n44370 ;
  assign n44372 = n4065 & ~n8247 ;
  assign n44373 = n44371 & n44372 ;
  assign n44374 = n91 & ~n44373 ;
  assign n44375 = ~n91 & n44374 ;
  assign n44376 = ~n33 & n2905 ;
  assign n44377 = n33 & n44376 ;
  assign n44378 = x6 & ~n44377 ;
  assign n44379 = n44375 & n44378 ;
  assign n44380 = ~n9513 & n15147 ;
  assign n44381 = n27635 ^ n4952 ^ 1'b0 ;
  assign n44382 = n44380 | n44381 ;
  assign n44383 = n18781 | n44382 ;
  assign n44384 = n44382 & ~n44383 ;
  assign n44385 = n27205 | n44384 ;
  assign n44386 = n44379 & ~n44385 ;
  assign n44387 = n29544 | n44386 ;
  assign n44388 = n5182 | n44387 ;
  assign n44389 = n44387 & ~n44388 ;
  assign n44390 = n13343 | n19544 ;
  assign n44391 = n3885 | n44390 ;
  assign n44392 = ~n18807 & n44391 ;
  assign n44393 = n44389 & n44392 ;
  assign n44394 = n3470 & n31311 ;
  assign n44395 = ~n2864 & n40080 ;
  assign n44396 = n22891 | n44395 ;
  assign n44397 = n263 & n29583 ;
  assign n44398 = n12821 & ~n28043 ;
  assign n44399 = n44398 ^ n13957 ^ 1'b0 ;
  assign n44400 = n9427 & ~n23698 ;
  assign n44401 = n43804 ^ n12060 ^ 1'b0 ;
  assign n44402 = n704 & ~n12649 ;
  assign n44403 = ~n3930 & n44402 ;
  assign n44404 = n2406 | n24566 ;
  assign n44405 = n34389 ^ n328 ^ n253 ;
  assign n44406 = n31182 ^ n4163 ^ 1'b0 ;
  assign n44407 = ~n2062 & n44406 ;
  assign n44408 = n44407 ^ n22785 ^ 1'b0 ;
  assign n44409 = n44408 ^ n25787 ^ n1917 ;
  assign n44410 = n14032 & ~n28648 ;
  assign n44411 = n44410 ^ n33641 ^ 1'b0 ;
  assign n44413 = n12873 ^ n3791 ^ 1'b0 ;
  assign n44412 = n4780 & n7554 ;
  assign n44414 = n44413 ^ n44412 ^ 1'b0 ;
  assign n44415 = ~n1877 & n7739 ;
  assign n44416 = ( n8342 & n11292 ) | ( n8342 & n11977 ) | ( n11292 & n11977 ) ;
  assign n44417 = n44416 ^ n27909 ^ n11286 ;
  assign n44418 = n44417 ^ n23254 ^ 1'b0 ;
  assign n44419 = ~n44415 & n44418 ;
  assign n44420 = n564 & n12456 ;
  assign n44421 = ~n31939 & n44420 ;
  assign n44422 = n28086 | n31596 ;
  assign n44423 = n1276 & ~n25571 ;
  assign n44424 = n40171 | n44423 ;
  assign n44425 = n2314 & n5898 ;
  assign n44426 = n44425 ^ n10935 ^ 1'b0 ;
  assign n44427 = n6410 ^ n758 ^ 1'b0 ;
  assign n44428 = n25268 & ~n44427 ;
  assign n44429 = n5969 | n8650 ;
  assign n44430 = n11098 ^ n1576 ^ 1'b0 ;
  assign n44431 = n18031 | n44430 ;
  assign n44432 = n44431 ^ n16167 ^ n13071 ;
  assign n44433 = n1534 | n18220 ;
  assign n44434 = n2554 | n44433 ;
  assign n44435 = n44432 & ~n44434 ;
  assign n44436 = ~n2101 & n8795 ;
  assign n44437 = ~n31756 & n44436 ;
  assign n44438 = n44435 & n44437 ;
  assign n44439 = n32864 ^ n24726 ^ n24208 ;
  assign n44440 = n38265 ^ n12167 ^ 1'b0 ;
  assign n44441 = n298 & ~n44440 ;
  assign n44442 = n19910 ^ n104 ^ 1'b0 ;
  assign n44443 = n10797 | n44442 ;
  assign n44444 = n10425 & n16211 ;
  assign n44445 = n44443 & n44444 ;
  assign n44446 = n16448 & ~n22499 ;
  assign n44447 = n44445 & n44446 ;
  assign n44448 = n28443 & ~n44447 ;
  assign n44449 = n2283 & n44448 ;
  assign n44450 = n30843 ^ n18386 ^ n2568 ;
  assign n44451 = n28946 & n44450 ;
  assign n44452 = n21026 & ~n34885 ;
  assign n44453 = n44452 ^ n16876 ^ 1'b0 ;
  assign n44454 = n2303 & ~n32120 ;
  assign n44455 = ~n11911 & n44454 ;
  assign n44456 = n30873 & ~n39686 ;
  assign n44457 = ~n20004 & n44456 ;
  assign n44458 = n15499 & ~n30003 ;
  assign n44459 = n34041 ^ n17070 ^ 1'b0 ;
  assign n44460 = n11468 & ~n44459 ;
  assign n44461 = n24384 | n24753 ;
  assign n44462 = n32778 & ~n37948 ;
  assign n44463 = ~n135 & n44462 ;
  assign n44464 = n11111 ^ n1635 ^ 1'b0 ;
  assign n44465 = n12421 | n44464 ;
  assign n44466 = n16538 & n27886 ;
  assign n44467 = ~n27221 & n44466 ;
  assign n44468 = n5187 & n15436 ;
  assign n44469 = n34179 & n44468 ;
  assign n44470 = n12295 ^ n1411 ^ 1'b0 ;
  assign n44471 = ~n2161 & n13836 ;
  assign n44477 = n4347 ^ n3731 ^ 1'b0 ;
  assign n44474 = n10942 | n21867 ;
  assign n44475 = n35253 | n44474 ;
  assign n44476 = n44475 ^ n12393 ^ 1'b0 ;
  assign n44472 = ~n1109 & n13376 ;
  assign n44473 = ~n18900 & n44472 ;
  assign n44478 = n44477 ^ n44476 ^ n44473 ;
  assign n44479 = n796 | n25346 ;
  assign n44480 = n7759 & ~n44479 ;
  assign n44481 = n36742 & ~n44480 ;
  assign n44482 = ~n27353 & n44481 ;
  assign n44483 = n19980 ^ n15145 ^ 1'b0 ;
  assign n44484 = n18390 ^ n1631 ^ 1'b0 ;
  assign n44485 = n4377 ^ n4267 ^ 1'b0 ;
  assign n44486 = ~n21004 & n44485 ;
  assign n44487 = n44486 ^ n42196 ^ 1'b0 ;
  assign n44488 = n13700 ^ n13169 ^ n12686 ;
  assign n44489 = n16924 & ~n44488 ;
  assign n44490 = n44489 ^ n11779 ^ 1'b0 ;
  assign n44491 = n997 | n8555 ;
  assign n44492 = n12654 | n44491 ;
  assign n44493 = n17193 & n44492 ;
  assign n44495 = ~n9570 & n24126 ;
  assign n44496 = n16312 & n44495 ;
  assign n44494 = n9553 & n38757 ;
  assign n44497 = n44496 ^ n44494 ^ n5710 ;
  assign n44498 = n40851 ^ n15641 ^ 1'b0 ;
  assign n44499 = n12544 | n31035 ;
  assign n44500 = n15565 | n44499 ;
  assign n44501 = n11323 | n20927 ;
  assign n44502 = n28935 ^ n5010 ^ 1'b0 ;
  assign n44503 = n4903 | n44502 ;
  assign n44504 = ( ~n1981 & n3727 ) | ( ~n1981 & n4367 ) | ( n3727 & n4367 ) ;
  assign n44505 = n13172 | n44504 ;
  assign n44506 = ~n1431 & n10262 ;
  assign n44507 = ( n2480 & n18126 ) | ( n2480 & ~n34155 ) | ( n18126 & ~n34155 ) ;
  assign n44508 = n14727 | n35243 ;
  assign n44509 = n44507 | n44508 ;
  assign n44510 = n44509 ^ n4416 ^ 1'b0 ;
  assign n44511 = n16496 & ~n32223 ;
  assign n44512 = n36754 & n44511 ;
  assign n44513 = n21819 & ~n36485 ;
  assign n44514 = ~n5214 & n44513 ;
  assign n44515 = n14409 | n19831 ;
  assign n44516 = n840 & n7652 ;
  assign n44517 = n35339 | n44516 ;
  assign n44518 = n36919 ^ n17239 ^ n1237 ;
  assign n44519 = n5914 | n13293 ;
  assign n44520 = n3880 | n44519 ;
  assign n44521 = ~n1771 & n14676 ;
  assign n44522 = ~n11530 & n12588 ;
  assign n44523 = n44522 ^ n1513 ^ 1'b0 ;
  assign n44524 = n8273 | n16294 ;
  assign n44526 = n14471 & ~n23637 ;
  assign n44525 = n2403 & ~n35475 ;
  assign n44527 = n44526 ^ n44525 ^ 1'b0 ;
  assign n44528 = ( n2114 & n21657 ) | ( n2114 & n44527 ) | ( n21657 & n44527 ) ;
  assign n44530 = n27897 ^ n26465 ^ 1'b0 ;
  assign n44531 = ~n18004 & n44530 ;
  assign n44529 = n468 | n562 ;
  assign n44532 = n44531 ^ n44529 ^ 1'b0 ;
  assign n44533 = ( n625 & n5052 ) | ( n625 & n8536 ) | ( n5052 & n8536 ) ;
  assign n44534 = ( n10952 & n27635 ) | ( n10952 & n44533 ) | ( n27635 & n44533 ) ;
  assign n44535 = n41599 & n44534 ;
  assign n44536 = n44535 ^ n25796 ^ 1'b0 ;
  assign n44537 = n736 & n8578 ;
  assign n44538 = n7792 & n23944 ;
  assign n44539 = ~n28999 & n44538 ;
  assign n44540 = n32322 & ~n44539 ;
  assign n44541 = ~n44537 & n44540 ;
  assign n44542 = n11683 ^ n7844 ^ 1'b0 ;
  assign n44543 = ( ~n10083 & n12320 ) | ( ~n10083 & n21073 ) | ( n12320 & n21073 ) ;
  assign n44547 = n36628 ^ n2802 ^ 1'b0 ;
  assign n44544 = n2727 ^ n2381 ^ 1'b0 ;
  assign n44545 = n2828 | n44544 ;
  assign n44546 = n5455 & ~n44545 ;
  assign n44548 = n44547 ^ n44546 ^ 1'b0 ;
  assign n44549 = n3240 & ~n11899 ;
  assign n44550 = n44549 ^ n25255 ^ 1'b0 ;
  assign n44551 = n12679 & n14107 ;
  assign n44554 = n6861 & n17346 ;
  assign n44555 = ~n11258 & n44554 ;
  assign n44556 = n44555 ^ n9227 ^ 1'b0 ;
  assign n44552 = n31045 ^ n6663 ^ 1'b0 ;
  assign n44553 = ~n12195 & n44552 ;
  assign n44557 = n44556 ^ n44553 ^ 1'b0 ;
  assign n44558 = n30031 ^ n18317 ^ 1'b0 ;
  assign n44559 = ~n16941 & n44231 ;
  assign n44562 = n13230 | n31186 ;
  assign n44563 = n31186 & ~n44562 ;
  assign n44564 = n44563 ^ n2491 ^ 1'b0 ;
  assign n44560 = n14983 | n29395 ;
  assign n44561 = n14983 & ~n44560 ;
  assign n44565 = n44564 ^ n44561 ^ 1'b0 ;
  assign n44566 = n6161 ^ n3970 ^ 1'b0 ;
  assign n44567 = n11433 & n17084 ;
  assign n44568 = n8725 & n44567 ;
  assign n44569 = n24643 | n44568 ;
  assign n44570 = n44569 ^ n16236 ^ 1'b0 ;
  assign n44571 = n2355 | n34073 ;
  assign n44572 = ~n2554 & n3620 ;
  assign n44573 = ~n17855 & n44572 ;
  assign n44574 = n19347 ^ n493 ^ 1'b0 ;
  assign n44575 = n18773 & ~n44574 ;
  assign n44576 = n8030 & n44575 ;
  assign n44577 = n26643 ^ n14269 ^ 1'b0 ;
  assign n44578 = ~n5305 & n40763 ;
  assign n44579 = n14559 ^ n3118 ^ 1'b0 ;
  assign n44580 = ~n4497 & n44579 ;
  assign n44581 = ~n7975 & n14918 ;
  assign n44582 = n2306 | n44581 ;
  assign n44583 = ~n4159 & n44582 ;
  assign n44584 = n5247 ^ n3451 ^ n3412 ;
  assign n44585 = ( ~n14243 & n43367 ) | ( ~n14243 & n44584 ) | ( n43367 & n44584 ) ;
  assign n44586 = n3161 & n39531 ;
  assign n44587 = n13860 & n36681 ;
  assign n44588 = n6231 & ~n25191 ;
  assign n44589 = n44588 ^ n22050 ^ n4299 ;
  assign n44590 = n19281 & ~n44589 ;
  assign n44591 = ~n33995 & n44590 ;
  assign n44592 = ~n630 & n3242 ;
  assign n44594 = n2303 & n4984 ;
  assign n44595 = n44594 ^ n2885 ^ 1'b0 ;
  assign n44593 = ~n131 & n20706 ;
  assign n44596 = n44595 ^ n44593 ^ 1'b0 ;
  assign n44597 = n44596 ^ n1062 ^ 1'b0 ;
  assign n44598 = ~n1922 & n4007 ;
  assign n44599 = n484 & n27331 ;
  assign n44600 = n30258 & n44599 ;
  assign n44601 = ~n5397 & n40548 ;
  assign n44602 = n7000 & n26420 ;
  assign n44603 = ~n28126 & n44602 ;
  assign n44608 = n593 | n1499 ;
  assign n44609 = n1499 & ~n44608 ;
  assign n44604 = n344 | n10724 ;
  assign n44605 = n10724 & ~n44604 ;
  assign n44606 = n2924 | n44605 ;
  assign n44607 = n44605 & ~n44606 ;
  assign n44610 = n44609 ^ n44607 ^ n28815 ;
  assign n44611 = n7271 ^ n4593 ^ 1'b0 ;
  assign n44612 = n21921 | n44611 ;
  assign n44613 = n160 & ~n15365 ;
  assign n44614 = ~n44612 & n44613 ;
  assign n44615 = n44614 ^ n3081 ^ 1'b0 ;
  assign n44616 = n7926 | n35554 ;
  assign n44617 = n44616 ^ n30899 ^ 1'b0 ;
  assign n44618 = n31078 & n44617 ;
  assign n44619 = n44618 ^ n21640 ^ 1'b0 ;
  assign n44620 = n17044 & n22262 ;
  assign n44621 = n19201 ^ n4294 ^ 1'b0 ;
  assign n44622 = n24022 | n44621 ;
  assign n44626 = n6753 ^ n918 ^ 1'b0 ;
  assign n44623 = n7427 & n15953 ;
  assign n44624 = n44623 ^ n4336 ^ 1'b0 ;
  assign n44625 = n44624 ^ n40737 ^ n11032 ;
  assign n44627 = n44626 ^ n44625 ^ n31788 ;
  assign n44628 = n38963 ^ n24339 ^ 1'b0 ;
  assign n44629 = n21470 ^ n17341 ^ 1'b0 ;
  assign n44643 = n12599 ^ n188 ^ 1'b0 ;
  assign n44633 = n152 | n490 ;
  assign n44634 = n490 & ~n44633 ;
  assign n44635 = ~n192 & n1546 ;
  assign n44636 = n192 & n44635 ;
  assign n44637 = n44634 | n44636 ;
  assign n44638 = n44634 & ~n44637 ;
  assign n44630 = ~n305 & n3182 ;
  assign n44631 = ~n3182 & n44630 ;
  assign n44632 = n367 & n44631 ;
  assign n44639 = n44638 ^ n44632 ^ 1'b0 ;
  assign n44640 = ~n13797 & n27263 ;
  assign n44641 = ~n44639 & n44640 ;
  assign n44642 = n25865 | n44641 ;
  assign n44644 = n44643 ^ n44642 ^ 1'b0 ;
  assign n44645 = n1480 | n20077 ;
  assign n44646 = n44645 ^ n39344 ^ 1'b0 ;
  assign n44647 = n19220 ^ n16183 ^ 1'b0 ;
  assign n44648 = n3527 | n14538 ;
  assign n44649 = n41700 | n44648 ;
  assign n44650 = ~n60 & n40046 ;
  assign n44651 = n44650 ^ n25544 ^ 1'b0 ;
  assign n44652 = n21743 ^ n6179 ^ 1'b0 ;
  assign n44653 = n7800 ^ n4173 ^ 1'b0 ;
  assign n44654 = n44653 ^ n19886 ^ 1'b0 ;
  assign n44655 = n44652 | n44654 ;
  assign n44656 = n19899 ^ n5441 ^ 1'b0 ;
  assign n44657 = ( ~n279 & n8962 ) | ( ~n279 & n9735 ) | ( n8962 & n9735 ) ;
  assign n44658 = n44657 ^ n23785 ^ n676 ;
  assign n44659 = n37758 ^ n13488 ^ n667 ;
  assign n44660 = n2494 & n43995 ;
  assign n44661 = ~n23470 & n44660 ;
  assign n44662 = n31657 ^ n28581 ^ 1'b0 ;
  assign n44663 = n29103 ^ n20653 ^ 1'b0 ;
  assign n44664 = n44662 & ~n44663 ;
  assign n44665 = n1083 & n5217 ;
  assign n44666 = n32359 & n44665 ;
  assign n44667 = n6032 & n15657 ;
  assign n44668 = n15315 & n44667 ;
  assign n44669 = n44668 ^ n13314 ^ 1'b0 ;
  assign n44670 = n2131 & ~n44669 ;
  assign n44672 = n9848 ^ n5481 ^ 1'b0 ;
  assign n44673 = n27781 & ~n44672 ;
  assign n44671 = n34635 ^ n13609 ^ 1'b0 ;
  assign n44674 = n44673 ^ n44671 ^ 1'b0 ;
  assign n44675 = n4440 & ~n5526 ;
  assign n44676 = n33150 | n44675 ;
  assign n44677 = n20957 ^ n13130 ^ 1'b0 ;
  assign n44678 = ( n40377 & ~n44676 ) | ( n40377 & n44677 ) | ( ~n44676 & n44677 ) ;
  assign n44679 = n4700 & ~n13664 ;
  assign n44680 = n39094 ^ n38429 ^ 1'b0 ;
  assign n44681 = ( n38763 & n44679 ) | ( n38763 & n44680 ) | ( n44679 & n44680 ) ;
  assign n44682 = n1542 & n40421 ;
  assign n44683 = ~n5249 & n44682 ;
  assign n44684 = n14870 ^ n12593 ^ 1'b0 ;
  assign n44685 = n5266 & n44684 ;
  assign n44686 = n36736 ^ n2248 ^ 1'b0 ;
  assign n44687 = n30723 & n40236 ;
  assign n44688 = n33819 ^ n29972 ^ 1'b0 ;
  assign n44689 = n44687 & n44688 ;
  assign n44690 = n30728 ^ n667 ^ 1'b0 ;
  assign n44691 = n972 & n44690 ;
  assign n44692 = ~n15321 & n44691 ;
  assign n44693 = n14055 ^ n1645 ^ 1'b0 ;
  assign n44694 = n44693 ^ n22601 ^ n7087 ;
  assign n44696 = n3651 | n32069 ;
  assign n44697 = n709 | n44696 ;
  assign n44698 = n44697 ^ n19625 ^ 1'b0 ;
  assign n44695 = n5001 & ~n10888 ;
  assign n44699 = n44698 ^ n44695 ^ 1'b0 ;
  assign n44700 = ~n3564 & n6655 ;
  assign n44701 = n6009 & n14670 ;
  assign n44702 = n44701 ^ n15937 ^ 1'b0 ;
  assign n44703 = n44247 ^ n12762 ^ n12297 ;
  assign n44704 = n44702 & n44703 ;
  assign n44705 = n44700 | n44704 ;
  assign n44706 = n12985 & n44705 ;
  assign n44707 = n14161 ^ n8729 ^ 1'b0 ;
  assign n44708 = ~n2317 & n44707 ;
  assign n44709 = n2247 | n5930 ;
  assign n44710 = n44709 ^ n443 ^ 1'b0 ;
  assign n44711 = n44708 & ~n44710 ;
  assign n44712 = ~n17449 & n28785 ;
  assign n44713 = ~n13801 & n25549 ;
  assign n44714 = n44713 ^ n5991 ^ n5736 ;
  assign n44715 = n2308 & n44714 ;
  assign n44716 = ~n44712 & n44715 ;
  assign n44717 = ~n7803 & n13044 ;
  assign n44718 = ~n30 & n44717 ;
  assign n44719 = n35625 & ~n44718 ;
  assign n44721 = n14844 ^ n6749 ^ 1'b0 ;
  assign n44722 = n44721 ^ n13248 ^ n10812 ;
  assign n44720 = n6758 | n8904 ;
  assign n44723 = n44722 ^ n44720 ^ 1'b0 ;
  assign n44724 = ~n9522 & n13340 ;
  assign n44725 = n15896 ^ n5338 ^ 1'b0 ;
  assign n44726 = n4555 & ~n44725 ;
  assign n44727 = ~n26688 & n44726 ;
  assign n44728 = n36504 ^ n23896 ^ 1'b0 ;
  assign n44729 = ~n34739 & n44728 ;
  assign n44730 = n42127 ^ n2252 ^ 1'b0 ;
  assign n44731 = ~n6401 & n15769 ;
  assign n44732 = n17777 & n44731 ;
  assign n44733 = n39086 ^ n15406 ^ 1'b0 ;
  assign n44734 = ~n4916 & n13436 ;
  assign n44735 = n17167 & n44734 ;
  assign n44736 = n36083 | n44735 ;
  assign n44737 = n15898 & ~n44736 ;
  assign n44738 = ~n10378 & n15832 ;
  assign n44739 = n44738 ^ n5706 ^ 1'b0 ;
  assign n44740 = ~n6550 & n44739 ;
  assign n44741 = n6237 & ~n8475 ;
  assign n44742 = n16379 | n27565 ;
  assign n44743 = n44742 ^ n30985 ^ 1'b0 ;
  assign n44744 = n13182 ^ n7961 ^ n6065 ;
  assign n44745 = n7108 & n44744 ;
  assign n44746 = ~n13755 & n44745 ;
  assign n44747 = n44746 ^ n38943 ^ n37498 ;
  assign n44748 = n21366 & ~n43417 ;
  assign n44749 = n44748 ^ n24862 ^ 1'b0 ;
  assign n44750 = ~n18853 & n29474 ;
  assign n44751 = ( n22147 & n34147 ) | ( n22147 & n42111 ) | ( n34147 & n42111 ) ;
  assign n44752 = n18830 ^ n14358 ^ 1'b0 ;
  assign n44753 = ~n23571 & n44752 ;
  assign n44754 = n2845 & ~n41442 ;
  assign n44755 = n9193 & ~n31273 ;
  assign n44756 = n44755 ^ n8729 ^ 1'b0 ;
  assign n44757 = n12105 & n44756 ;
  assign n44758 = ~n25079 & n30181 ;
  assign n44759 = ( n15358 & ~n27625 ) | ( n15358 & n42219 ) | ( ~n27625 & n42219 ) ;
  assign n44760 = n33368 | n37855 ;
  assign n44761 = n31166 & ~n44760 ;
  assign n44762 = n25215 | n27751 ;
  assign n44763 = n22469 & ~n44762 ;
  assign n44764 = ~n2435 & n11400 ;
  assign n44765 = ~n9988 & n44764 ;
  assign n44766 = n29395 ^ n2137 ^ 1'b0 ;
  assign n44767 = n44766 ^ n34649 ^ 1'b0 ;
  assign n44768 = n12190 ^ n6383 ^ 1'b0 ;
  assign n44769 = ~n5179 & n44768 ;
  assign n44770 = n44769 ^ n38510 ^ 1'b0 ;
  assign n44771 = n44770 ^ n43682 ^ 1'b0 ;
  assign n44772 = n25418 & n39561 ;
  assign n44773 = ~n27227 & n44772 ;
  assign n44774 = n18227 ^ n7770 ^ n4028 ;
  assign n44775 = n9222 | n21215 ;
  assign n44776 = n44775 ^ n1044 ^ 1'b0 ;
  assign n44777 = n10247 & ~n44776 ;
  assign n44778 = n17075 ^ n5623 ^ 1'b0 ;
  assign n44779 = n11283 & n44778 ;
  assign n44780 = n18519 ^ n3985 ^ 1'b0 ;
  assign n44781 = ~n3004 & n9324 ;
  assign n44782 = n44781 ^ n315 ^ 1'b0 ;
  assign n44783 = n44782 ^ n470 ^ 1'b0 ;
  assign n44784 = n6919 & ~n14538 ;
  assign n44785 = n44784 ^ n35904 ^ 1'b0 ;
  assign n44786 = n1392 & n41416 ;
  assign n44787 = n5303 & n44786 ;
  assign n44788 = n34295 ^ n32627 ^ 1'b0 ;
  assign n44789 = n44476 ^ n6522 ^ 1'b0 ;
  assign n44790 = n18480 ^ n8857 ^ 1'b0 ;
  assign n44791 = ~n28985 & n44790 ;
  assign n44792 = ~n44789 & n44791 ;
  assign n44793 = n8233 & ~n10809 ;
  assign n44794 = ~n16639 & n25691 ;
  assign n44795 = n8443 | n21707 ;
  assign n44796 = n28490 | n44795 ;
  assign n44797 = ~n4626 & n6512 ;
  assign n44798 = n12754 & n44797 ;
  assign n44799 = n7864 & n23871 ;
  assign n44800 = n44798 & n44799 ;
  assign n44801 = n2018 ^ n885 ^ 1'b0 ;
  assign n44802 = n44801 ^ n29676 ^ 1'b0 ;
  assign n44803 = n21286 ^ n21026 ^ n12943 ;
  assign n44804 = n12279 ^ n6230 ^ 1'b0 ;
  assign n44805 = n16028 ^ n535 ^ 1'b0 ;
  assign n44806 = n17678 & ~n19295 ;
  assign n44807 = ~n44805 & n44806 ;
  assign n44808 = ( ~n18505 & n44804 ) | ( ~n18505 & n44807 ) | ( n44804 & n44807 ) ;
  assign n44809 = n4741 | n16820 ;
  assign n44810 = n17150 & ~n44809 ;
  assign n44811 = n44810 ^ n23200 ^ 1'b0 ;
  assign n44812 = ~n18191 & n44811 ;
  assign n44813 = n21892 & ~n31297 ;
  assign n44814 = n44813 ^ n6649 ^ 1'b0 ;
  assign n44815 = ~n5936 & n39983 ;
  assign n44816 = n9917 & n23573 ;
  assign n44817 = ~n27836 & n44816 ;
  assign n44818 = n13129 ^ n12450 ^ 1'b0 ;
  assign n44819 = n44818 ^ n42487 ^ 1'b0 ;
  assign n44820 = ( n2226 & n18347 ) | ( n2226 & ~n19050 ) | ( n18347 & ~n19050 ) ;
  assign n44821 = n3871 & n44820 ;
  assign n44822 = n39982 & ~n44821 ;
  assign n44823 = n302 & n5769 ;
  assign n44824 = n44823 ^ n15273 ^ n1428 ;
  assign n44825 = n44824 ^ n4997 ^ n576 ;
  assign n44826 = n15326 & ~n44825 ;
  assign n44827 = ~n21256 & n27239 ;
  assign n44828 = ~n28354 & n38337 ;
  assign n44829 = n18930 ^ n12007 ^ 1'b0 ;
  assign n44830 = ~n698 & n1658 ;
  assign n44831 = n13843 & n44830 ;
  assign n44832 = n20604 ^ n1528 ^ 1'b0 ;
  assign n44833 = n44831 | n44832 ;
  assign n44834 = n35345 & n44833 ;
  assign n44835 = n4060 & n35350 ;
  assign n44836 = n37346 ^ n18363 ^ 1'b0 ;
  assign n44837 = n44836 ^ n26631 ^ n18893 ;
  assign n44838 = n17197 ^ n7054 ^ 1'b0 ;
  assign n44839 = ( n13566 & ~n19198 ) | ( n13566 & n44838 ) | ( ~n19198 & n44838 ) ;
  assign n44841 = ~n6776 & n11657 ;
  assign n44840 = ~n8529 & n17873 ;
  assign n44842 = n44841 ^ n44840 ^ 1'b0 ;
  assign n44843 = n20606 ^ n1428 ^ 1'b0 ;
  assign n44844 = n7534 & n8697 ;
  assign n44845 = n44844 ^ n25017 ^ 1'b0 ;
  assign n44846 = n4082 | n44845 ;
  assign n44847 = n1215 & ~n8894 ;
  assign n44848 = ~n32815 & n44847 ;
  assign n44849 = n15370 | n44848 ;
  assign n44850 = n15920 | n44358 ;
  assign n44851 = ~n16671 & n24428 ;
  assign n44852 = ~n9177 & n33674 ;
  assign n44853 = ~n40712 & n44852 ;
  assign n44854 = ( n10124 & n21915 ) | ( n10124 & n42417 ) | ( n21915 & n42417 ) ;
  assign n44855 = n4560 | n9995 ;
  assign n44856 = n36151 | n44855 ;
  assign n44857 = n12520 ^ n4946 ^ n3554 ;
  assign n44858 = n2368 & n37274 ;
  assign n44859 = n3088 | n5685 ;
  assign n44860 = n2361 & ~n44859 ;
  assign n44861 = n8118 & n11562 ;
  assign n44862 = n8689 & ~n44861 ;
  assign n44863 = n20810 | n35802 ;
  assign n44864 = n4823 | n40578 ;
  assign n44865 = n6660 & ~n44864 ;
  assign n44866 = n5131 & ~n43770 ;
  assign n44867 = ~n23650 & n44866 ;
  assign n44868 = n4366 | n26702 ;
  assign n44869 = ~n2381 & n44868 ;
  assign n44870 = n41223 ^ n15105 ^ 1'b0 ;
  assign n44871 = ~n44869 & n44870 ;
  assign n44872 = n19548 & n44871 ;
  assign n44873 = ~n24773 & n29038 ;
  assign n44874 = n5270 & n17210 ;
  assign n44875 = ~n35861 & n44874 ;
  assign n44876 = ~n4139 & n11331 ;
  assign n44877 = n44876 ^ n4653 ^ 1'b0 ;
  assign n44878 = n44877 ^ n15416 ^ 1'b0 ;
  assign n44879 = n44878 ^ n26774 ^ 1'b0 ;
  assign n44880 = n11058 | n44879 ;
  assign n44881 = ( ~n17588 & n21052 ) | ( ~n17588 & n27586 ) | ( n21052 & n27586 ) ;
  assign n44882 = n640 & n44881 ;
  assign n44885 = n2298 | n4539 ;
  assign n44886 = n44885 ^ n8156 ^ 1'b0 ;
  assign n44887 = n27628 ^ n18963 ^ 1'b0 ;
  assign n44888 = ( n5364 & n44886 ) | ( n5364 & n44887 ) | ( n44886 & n44887 ) ;
  assign n44883 = ~n11846 & n18948 ;
  assign n44884 = n44883 ^ n21256 ^ 1'b0 ;
  assign n44889 = n44888 ^ n44884 ^ 1'b0 ;
  assign n44890 = n28133 ^ n23273 ^ 1'b0 ;
  assign n44891 = n15101 & n18559 ;
  assign n44892 = ~n44890 & n44891 ;
  assign n44893 = n38596 | n44892 ;
  assign n44894 = n6282 | n44893 ;
  assign n44895 = n11597 ^ n6874 ^ 1'b0 ;
  assign n44896 = n41806 | n44895 ;
  assign n44897 = n36906 | n44896 ;
  assign n44898 = n23120 ^ n19164 ^ 1'b0 ;
  assign n44899 = ~n8406 & n44898 ;
  assign n44900 = n26838 ^ n8659 ^ 1'b0 ;
  assign n44901 = ~n23202 & n44900 ;
  assign n44902 = n39655 & n44901 ;
  assign n44903 = n44902 ^ n28360 ^ 1'b0 ;
  assign n44904 = n9751 ^ n8815 ^ 1'b0 ;
  assign n44905 = n42880 ^ n39818 ^ n548 ;
  assign n44906 = n14076 ^ n1743 ^ 1'b0 ;
  assign n44907 = ~n19437 & n38892 ;
  assign n44908 = ~n18016 & n27972 ;
  assign n44909 = n15331 ^ n2498 ^ 1'b0 ;
  assign n44910 = ~n4211 & n44909 ;
  assign n44911 = n44910 ^ n32940 ^ 1'b0 ;
  assign n44912 = n31425 ^ n10968 ^ 1'b0 ;
  assign n44913 = ~n27042 & n44912 ;
  assign n44914 = n27009 ^ n7338 ^ 1'b0 ;
  assign n44915 = n16819 & n22436 ;
  assign n44916 = n5336 & ~n25933 ;
  assign n44917 = n481 & n9643 ;
  assign n44918 = n44917 ^ n4707 ^ 1'b0 ;
  assign n44919 = n44918 ^ n28784 ^ 1'b0 ;
  assign n44920 = n44916 & ~n44919 ;
  assign n44921 = ( n3823 & n41916 ) | ( n3823 & n44920 ) | ( n41916 & n44920 ) ;
  assign n44922 = n20295 & ~n20653 ;
  assign n44923 = n30839 ^ n584 ^ 1'b0 ;
  assign n44924 = n44923 ^ n34956 ^ 1'b0 ;
  assign n44925 = n2046 | n44924 ;
  assign n44926 = n11279 ^ n10359 ^ 1'b0 ;
  assign n44927 = n15834 & n15844 ;
  assign n44928 = ~n44926 & n44927 ;
  assign n44929 = ~n10556 & n43648 ;
  assign n44930 = n41770 ^ n24568 ^ 1'b0 ;
  assign n44931 = n6785 & ~n32704 ;
  assign n44932 = n18312 & n44931 ;
  assign n44933 = n44932 ^ n30204 ^ n7827 ;
  assign n44934 = n7579 | n8073 ;
  assign n44935 = n7579 & ~n44934 ;
  assign n44936 = n7722 & ~n44935 ;
  assign n44937 = n44935 & n44936 ;
  assign n44938 = n44937 ^ n16546 ^ 1'b0 ;
  assign n44939 = n6820 & ~n11951 ;
  assign n44940 = n36851 ^ n54 ^ 1'b0 ;
  assign n44941 = n10054 & n31554 ;
  assign n44942 = n44941 ^ n11899 ^ 1'b0 ;
  assign n44943 = n19655 & n44942 ;
  assign n44944 = n44943 ^ n9113 ^ 1'b0 ;
  assign n44945 = n20189 ^ n12393 ^ 1'b0 ;
  assign n44946 = n489 | n44945 ;
  assign n44947 = n13620 | n21588 ;
  assign n44948 = n44947 ^ n5851 ^ 1'b0 ;
  assign n44949 = n22679 & n44948 ;
  assign n44950 = n9220 | n44949 ;
  assign n44951 = n27441 ^ n24481 ^ 1'b0 ;
  assign n44952 = n21178 & n38460 ;
  assign n44953 = n25804 | n37098 ;
  assign n44954 = n6789 & ~n44953 ;
  assign n44955 = ( n2238 & ~n44952 ) | ( n2238 & n44954 ) | ( ~n44952 & n44954 ) ;
  assign n44956 = n4321 & ~n44955 ;
  assign n44957 = n34921 ^ n13053 ^ 1'b0 ;
  assign n44958 = ~n12837 & n21449 ;
  assign n44959 = ~n19182 & n44958 ;
  assign n44960 = n2802 | n44959 ;
  assign n44961 = n44957 | n44960 ;
  assign n44965 = ~n49 & n16342 ;
  assign n44966 = n16893 & n44965 ;
  assign n44967 = n5540 & ~n44966 ;
  assign n44968 = n44967 ^ n26407 ^ 1'b0 ;
  assign n44969 = n2944 & ~n22991 ;
  assign n44970 = n44968 & n44969 ;
  assign n44962 = n14011 ^ n2306 ^ 1'b0 ;
  assign n44963 = n15435 & ~n44962 ;
  assign n44964 = n12328 & n44963 ;
  assign n44971 = n44970 ^ n44964 ^ 1'b0 ;
  assign n44973 = n3934 | n9133 ;
  assign n44974 = n44973 ^ n41818 ^ 1'b0 ;
  assign n44972 = n4463 & n42004 ;
  assign n44975 = n44974 ^ n44972 ^ 1'b0 ;
  assign n44977 = n14219 | n16962 ;
  assign n44978 = n44977 ^ n16455 ^ 1'b0 ;
  assign n44979 = n44978 ^ n9852 ^ 1'b0 ;
  assign n44980 = ~n7948 & n44979 ;
  assign n44976 = n11064 | n33896 ;
  assign n44981 = n44980 ^ n44976 ^ 1'b0 ;
  assign n44984 = n3920 & n12126 ;
  assign n44982 = ~n15105 & n16425 ;
  assign n44983 = n7031 & n44982 ;
  assign n44985 = n44984 ^ n44983 ^ 1'b0 ;
  assign n44986 = n2448 & ~n10280 ;
  assign n44987 = n30520 & ~n44986 ;
  assign n44988 = n26744 ^ n4925 ^ 1'b0 ;
  assign n44989 = n30997 ^ n5854 ^ n1313 ;
  assign n44990 = n646 & n12271 ;
  assign n44991 = n35536 ^ n4226 ^ 1'b0 ;
  assign n44992 = n17887 & n18096 ;
  assign n44993 = n44992 ^ n29457 ^ 1'b0 ;
  assign n44994 = n20254 ^ n4667 ^ 1'b0 ;
  assign n44995 = n43541 & n44994 ;
  assign n44996 = n1989 & ~n5016 ;
  assign n44997 = n25998 & ~n44996 ;
  assign n44998 = ~n3044 & n7401 ;
  assign n44999 = n44998 ^ n18881 ^ n2432 ;
  assign n45000 = ( ~n6048 & n8857 ) | ( ~n6048 & n32512 ) | ( n8857 & n32512 ) ;
  assign n45001 = n40263 ^ n32384 ^ 1'b0 ;
  assign n45002 = n31603 ^ n13907 ^ 1'b0 ;
  assign n45003 = n34368 ^ n9247 ^ 1'b0 ;
  assign n45004 = n9952 & n45003 ;
  assign n45005 = n1000 & n28546 ;
  assign n45006 = n4589 & n45005 ;
  assign n45008 = n7146 & n11162 ;
  assign n45007 = n4408 & n5410 ;
  assign n45009 = n45008 ^ n45007 ^ 1'b0 ;
  assign n45010 = n8660 ^ n4600 ^ 1'b0 ;
  assign n45011 = ~n9687 & n45010 ;
  assign n45012 = ~n9577 & n45011 ;
  assign n45013 = ( n4007 & n34694 ) | ( n4007 & n45012 ) | ( n34694 & n45012 ) ;
  assign n45014 = n7268 & ~n8036 ;
  assign n45015 = n27144 ^ n8960 ^ 1'b0 ;
  assign n45016 = n11300 ^ n10939 ^ 1'b0 ;
  assign n45017 = n4631 & n45016 ;
  assign n45018 = n45017 ^ n37018 ^ 1'b0 ;
  assign n45019 = n5236 & ~n13379 ;
  assign n45020 = n408 & ~n24874 ;
  assign n45021 = ( n20 & n17325 ) | ( n20 & n45020 ) | ( n17325 & n45020 ) ;
  assign n45022 = n2173 & ~n17673 ;
  assign n45023 = ~n27881 & n39397 ;
  assign n45024 = n45023 ^ n17038 ^ 1'b0 ;
  assign n45025 = n16946 & ~n22744 ;
  assign n45026 = n1877 & ~n4745 ;
  assign n45027 = ~n25597 & n45026 ;
  assign n45028 = ( n25968 & ~n32056 ) | ( n25968 & n32706 ) | ( ~n32056 & n32706 ) ;
  assign n45029 = n23609 ^ n3740 ^ 1'b0 ;
  assign n45030 = ( ~n3231 & n44235 ) | ( ~n3231 & n45029 ) | ( n44235 & n45029 ) ;
  assign n45031 = n1613 | n26250 ;
  assign n45032 = n1613 & ~n45031 ;
  assign n45033 = n14471 & ~n45032 ;
  assign n45034 = n45033 ^ n22951 ^ 1'b0 ;
  assign n45035 = n7030 | n45034 ;
  assign n45036 = n12271 & ~n45035 ;
  assign n45037 = ~n1459 & n24638 ;
  assign n45038 = n45037 ^ n31108 ^ 1'b0 ;
  assign n45039 = n35133 & n36024 ;
  assign n45040 = n7443 & n40751 ;
  assign n45041 = n19265 ^ n3235 ^ 1'b0 ;
  assign n45042 = n22741 & ~n45041 ;
  assign n45043 = n45042 ^ n9083 ^ 1'b0 ;
  assign n45044 = ~n9017 & n45043 ;
  assign n45045 = ~n7484 & n30868 ;
  assign n45046 = n3274 & n13345 ;
  assign n45047 = ~n283 & n45046 ;
  assign n45048 = n12109 | n25243 ;
  assign n45049 = n27369 | n45048 ;
  assign n45050 = n45047 & ~n45049 ;
  assign n45051 = n27979 & n29846 ;
  assign n45052 = ~n37951 & n45051 ;
  assign n45053 = n4149 | n45052 ;
  assign n45054 = n7430 | n45053 ;
  assign n45055 = ~n1426 & n38718 ;
  assign n45056 = n45055 ^ n3582 ^ 1'b0 ;
  assign n45057 = ~n22305 & n37710 ;
  assign n45058 = n14500 & ~n23129 ;
  assign n45059 = ~n17167 & n17789 ;
  assign n45060 = n45058 & n45059 ;
  assign n45061 = n4131 ^ n3592 ^ 1'b0 ;
  assign n45062 = n15086 ^ n9049 ^ 1'b0 ;
  assign n45063 = ~n45061 & n45062 ;
  assign n45064 = ( n1993 & n20819 ) | ( n1993 & n44962 ) | ( n20819 & n44962 ) ;
  assign n45065 = ~n33575 & n45064 ;
  assign n45066 = n19905 | n20912 ;
  assign n45067 = n14452 & ~n45066 ;
  assign n45068 = ~n3009 & n37173 ;
  assign n45069 = n24864 ^ n8831 ^ 1'b0 ;
  assign n45070 = n8820 | n16442 ;
  assign n45071 = n45070 ^ n13566 ^ 1'b0 ;
  assign n45072 = n36098 & ~n45071 ;
  assign n45073 = n24263 & ~n29789 ;
  assign n45074 = n15207 ^ n5763 ^ 1'b0 ;
  assign n45075 = n39030 & ~n45074 ;
  assign n45076 = ~n45073 & n45075 ;
  assign n45077 = n25170 ^ n23063 ^ 1'b0 ;
  assign n45078 = n10915 & n45077 ;
  assign n45079 = n14251 ^ n4632 ^ 1'b0 ;
  assign n45080 = n729 | n7893 ;
  assign n45081 = n40307 ^ n1141 ^ 1'b0 ;
  assign n45082 = n7843 & ~n15561 ;
  assign n45083 = n17497 & n45082 ;
  assign n45084 = n11240 & n17637 ;
  assign n45085 = n6722 & n45084 ;
  assign n45086 = n45085 ^ n11772 ^ 1'b0 ;
  assign n45087 = ( n11717 & ~n45083 ) | ( n11717 & n45086 ) | ( ~n45083 & n45086 ) ;
  assign n45088 = n37199 ^ n9583 ^ 1'b0 ;
  assign n45089 = n1410 & ~n2361 ;
  assign n45090 = n45089 ^ n11875 ^ 1'b0 ;
  assign n45091 = n12483 ^ n205 ^ 1'b0 ;
  assign n45092 = n45090 | n45091 ;
  assign n45093 = ~n6590 & n18442 ;
  assign n45094 = ~n38493 & n45093 ;
  assign n45095 = n12489 ^ n6151 ^ n1464 ;
  assign n45096 = n3174 & ~n6880 ;
  assign n45097 = n45096 ^ n26906 ^ 1'b0 ;
  assign n45098 = n45095 & ~n45097 ;
  assign n45099 = ~n8293 & n33441 ;
  assign n45100 = ~n38692 & n45099 ;
  assign n45101 = n12483 ^ n10834 ^ 1'b0 ;
  assign n45102 = n7651 & ~n45101 ;
  assign n45103 = n26 & n45102 ;
  assign n45104 = n27067 & n45103 ;
  assign n45105 = n25496 ^ n9882 ^ 1'b0 ;
  assign n45106 = n34631 ^ n34620 ^ 1'b0 ;
  assign n45107 = n34235 ^ n30844 ^ 1'b0 ;
  assign n45108 = n32521 ^ n4496 ^ 1'b0 ;
  assign n45109 = ~n1845 & n45108 ;
  assign n45110 = n4546 & ~n14073 ;
  assign n45111 = ~n45109 & n45110 ;
  assign n45112 = n7451 & n36996 ;
  assign n45113 = n2330 & n14396 ;
  assign n45114 = n45113 ^ n33992 ^ 1'b0 ;
  assign n45115 = n45114 ^ n9428 ^ 1'b0 ;
  assign n45116 = ( n2266 & n3484 ) | ( n2266 & ~n27411 ) | ( n3484 & ~n27411 ) ;
  assign n45117 = n9970 ^ n7927 ^ n1707 ;
  assign n45118 = n9046 ^ n6650 ^ 1'b0 ;
  assign n45119 = n5885 & n6664 ;
  assign n45120 = n13193 & n21296 ;
  assign n45121 = ~n13735 & n45120 ;
  assign n45122 = n774 & n19610 ;
  assign n45123 = n45122 ^ n16435 ^ 1'b0 ;
  assign n45124 = ~n7721 & n19680 ;
  assign n45125 = ~n45123 & n45124 ;
  assign n45126 = n24536 | n25146 ;
  assign n45127 = n8190 & ~n45126 ;
  assign n45128 = n29744 | n45127 ;
  assign n45129 = ( n3310 & n14080 ) | ( n3310 & n30933 ) | ( n14080 & n30933 ) ;
  assign n45130 = n340 | n2798 ;
  assign n45131 = n19602 & ~n45130 ;
  assign n45132 = n45131 ^ n4747 ^ 1'b0 ;
  assign n45133 = ~n4807 & n33300 ;
  assign n45134 = n11043 & n45133 ;
  assign n45135 = n18899 | n27011 ;
  assign n45136 = n6456 & n23045 ;
  assign n45137 = n45135 & n45136 ;
  assign n45138 = n2813 | n10539 ;
  assign n45139 = n45138 ^ n22939 ^ 1'b0 ;
  assign n45140 = n45139 ^ n14303 ^ 1'b0 ;
  assign n45141 = n17789 | n22985 ;
  assign n45142 = ( n16091 & n45140 ) | ( n16091 & n45141 ) | ( n45140 & n45141 ) ;
  assign n45143 = n6997 & n15527 ;
  assign n45144 = n45143 ^ n5465 ^ 1'b0 ;
  assign n45145 = n34579 & ~n35221 ;
  assign n45146 = n45145 ^ n36518 ^ 1'b0 ;
  assign n45147 = n6008 | n23541 ;
  assign n45148 = n45147 ^ n37091 ^ 1'b0 ;
  assign n45149 = n20177 & n28229 ;
  assign n45150 = n2388 & n45149 ;
  assign n45151 = n20452 ^ n10545 ^ 1'b0 ;
  assign n45152 = n41063 & n45151 ;
  assign n45153 = n45152 ^ n23908 ^ 1'b0 ;
  assign n45154 = n11318 ^ n9058 ^ 1'b0 ;
  assign n45155 = n2588 & n45154 ;
  assign n45156 = n45155 ^ n23793 ^ n5800 ;
  assign n45157 = n2207 | n6808 ;
  assign n45158 = n22558 & n45157 ;
  assign n45159 = n10470 & ~n12625 ;
  assign n45160 = ~n903 & n45159 ;
  assign n45161 = n45160 ^ n16634 ^ n4074 ;
  assign n45162 = n42475 & n45161 ;
  assign n45163 = n45162 ^ n5636 ^ 1'b0 ;
  assign n45164 = n8874 & ~n19970 ;
  assign n45165 = n45164 ^ n2813 ^ 1'b0 ;
  assign n45166 = n45165 ^ n19716 ^ 1'b0 ;
  assign n45167 = ~n646 & n22870 ;
  assign n45168 = n45166 & n45167 ;
  assign n45169 = n39274 | n45168 ;
  assign n45170 = n7839 & ~n21062 ;
  assign n45171 = n22568 ^ n9584 ^ n5976 ;
  assign n45172 = ~n2922 & n36891 ;
  assign n45173 = ( n7100 & n9536 ) | ( n7100 & n19113 ) | ( n9536 & n19113 ) ;
  assign n45174 = n36534 ^ n3443 ^ 1'b0 ;
  assign n45175 = n45174 ^ n23482 ^ n20298 ;
  assign n45176 = ~n700 & n2721 ;
  assign n45177 = n22857 ^ n14550 ^ 1'b0 ;
  assign n45178 = n45176 & ~n45177 ;
  assign n45179 = n11704 & n24346 ;
  assign n45180 = n5672 & n45010 ;
  assign n45181 = ~n45179 & n45180 ;
  assign n45182 = n38715 ^ n7099 ^ 1'b0 ;
  assign n45183 = n19151 | n30733 ;
  assign n45184 = n1576 & ~n12328 ;
  assign n45185 = n45184 ^ n20370 ^ 1'b0 ;
  assign n45186 = n9148 | n45185 ;
  assign n45187 = ~n8144 & n24263 ;
  assign n45188 = n45186 & n45187 ;
  assign n45189 = n11535 | n20268 ;
  assign n45190 = n45189 ^ n21418 ^ n12225 ;
  assign n45191 = n45188 | n45190 ;
  assign n45192 = n45183 | n45191 ;
  assign n45193 = n19515 ^ n15301 ^ n1956 ;
  assign n45194 = n6504 & n6766 ;
  assign n45195 = n10758 | n39336 ;
  assign n45196 = n12906 & ~n45195 ;
  assign n45197 = n27302 & n45196 ;
  assign n45198 = n1987 | n2491 ;
  assign n45199 = n45198 ^ n1887 ^ 1'b0 ;
  assign n45201 = n34818 ^ n9391 ^ 1'b0 ;
  assign n45200 = ( ~n1099 & n1469 ) | ( ~n1099 & n40155 ) | ( n1469 & n40155 ) ;
  assign n45202 = n45201 ^ n45200 ^ n38617 ;
  assign n45203 = n3259 & n12189 ;
  assign n45204 = n45203 ^ n1069 ^ n220 ;
  assign n45205 = n29399 ^ n3825 ^ 1'b0 ;
  assign n45207 = n3377 & ~n6494 ;
  assign n45206 = n20333 ^ n15091 ^ n1491 ;
  assign n45208 = n45207 ^ n45206 ^ 1'b0 ;
  assign n45209 = ~n8368 & n30433 ;
  assign n45210 = ~n6296 & n45209 ;
  assign n45211 = n17812 & ~n40840 ;
  assign n45212 = n19305 | n22073 ;
  assign n45214 = n32185 ^ n19888 ^ 1'b0 ;
  assign n45213 = n14152 | n41510 ;
  assign n45215 = n45214 ^ n45213 ^ n6927 ;
  assign n45216 = n33851 ^ n24624 ^ 1'b0 ;
  assign n45217 = n24094 & n45216 ;
  assign n45218 = n11453 | n17402 ;
  assign n45219 = n45218 ^ n9477 ^ 1'b0 ;
  assign n45220 = n45219 ^ n33482 ^ 1'b0 ;
  assign n45221 = n19 & n7034 ;
  assign n45222 = n45221 ^ n13863 ^ 1'b0 ;
  assign n45223 = n5297 | n21710 ;
  assign n45224 = n2991 & ~n6834 ;
  assign n45225 = n45224 ^ n552 ^ 1'b0 ;
  assign n45226 = n108 & n10290 ;
  assign n45227 = n10967 & n25867 ;
  assign n45228 = ( n28070 & n31004 ) | ( n28070 & n45227 ) | ( n31004 & n45227 ) ;
  assign n45229 = n35128 ^ n10159 ^ n4707 ;
  assign n45230 = n45228 | n45229 ;
  assign n45231 = n45226 & ~n45230 ;
  assign n45235 = n10066 ^ n2074 ^ 1'b0 ;
  assign n45236 = n4203 & n45235 ;
  assign n45232 = n874 | n12125 ;
  assign n45233 = n27676 & ~n45232 ;
  assign n45234 = ( n5528 & n32227 ) | ( n5528 & n45233 ) | ( n32227 & n45233 ) ;
  assign n45237 = n45236 ^ n45234 ^ n43636 ;
  assign n45238 = n7617 & n28347 ;
  assign n45239 = n38987 ^ n3224 ^ n1566 ;
  assign n45240 = ~n9600 & n41702 ;
  assign n45241 = n29525 ^ n18962 ^ 1'b0 ;
  assign n45242 = n11383 & n27959 ;
  assign n45243 = n45242 ^ n1407 ^ 1'b0 ;
  assign n45244 = n45243 ^ n10851 ^ 1'b0 ;
  assign n45245 = ~n45241 & n45244 ;
  assign n45246 = n40771 ^ n32454 ^ n2164 ;
  assign n45247 = ( n18486 & ~n33127 ) | ( n18486 & n45246 ) | ( ~n33127 & n45246 ) ;
  assign n45248 = ~n642 & n10635 ;
  assign n45249 = ~n45247 & n45248 ;
  assign n45250 = n45249 ^ n38327 ^ 1'b0 ;
  assign n45251 = n29604 & ~n45250 ;
  assign n45253 = ~n12436 & n28927 ;
  assign n45254 = ~n9031 & n45253 ;
  assign n45252 = n2663 & n19903 ;
  assign n45255 = n45254 ^ n45252 ^ 1'b0 ;
  assign n45256 = n2022 | n18099 ;
  assign n45257 = n45256 ^ n17439 ^ 1'b0 ;
  assign n45258 = n45257 ^ n41209 ^ 1'b0 ;
  assign n45259 = ( ~n10709 & n33543 ) | ( ~n10709 & n43532 ) | ( n33543 & n43532 ) ;
  assign n45260 = n45259 ^ n32857 ^ 1'b0 ;
  assign n45261 = n37045 ^ n6030 ^ 1'b0 ;
  assign n45262 = n3583 & n45261 ;
  assign n45263 = ~n5660 & n41083 ;
  assign n45264 = ~n1667 & n35597 ;
  assign n45265 = n36114 ^ n20833 ^ 1'b0 ;
  assign n45266 = n4367 & ~n29076 ;
  assign n45267 = ( n25793 & ~n34883 ) | ( n25793 & n45266 ) | ( ~n34883 & n45266 ) ;
  assign n45268 = n17632 ^ n5497 ^ 1'b0 ;
  assign n45269 = n6762 | n18414 ;
  assign n45270 = n25234 ^ n11967 ^ 1'b0 ;
  assign n45271 = ~n19633 & n45270 ;
  assign n45272 = ( n22214 & n26071 ) | ( n22214 & ~n32038 ) | ( n26071 & ~n32038 ) ;
  assign n45273 = n43755 ^ n2946 ^ 1'b0 ;
  assign n45274 = n957 & n45273 ;
  assign n45275 = n45274 ^ n25913 ^ n10511 ;
  assign n45276 = n4432 & n30471 ;
  assign n45277 = n12261 & ~n45276 ;
  assign n45278 = n39336 ^ n13758 ^ 1'b0 ;
  assign n45279 = n1300 & ~n45278 ;
  assign n45281 = n7902 & ~n8487 ;
  assign n45282 = ~n31973 & n45281 ;
  assign n45283 = n45282 ^ n6975 ^ 1'b0 ;
  assign n45280 = ~n6454 & n35875 ;
  assign n45284 = n45283 ^ n45280 ^ 1'b0 ;
  assign n45285 = ~n17775 & n32780 ;
  assign n45286 = n45285 ^ n10299 ^ 1'b0 ;
  assign n45287 = n12974 & n38521 ;
  assign n45288 = n19581 & ~n21470 ;
  assign n45289 = n25146 & n45288 ;
  assign n45290 = n31965 ^ n10298 ^ 1'b0 ;
  assign n45291 = n45289 | n45290 ;
  assign n45292 = ~n17840 & n19834 ;
  assign n45293 = n45292 ^ n21391 ^ n56 ;
  assign n45294 = n6057 | n27296 ;
  assign n45295 = n43110 ^ n24480 ^ n17427 ;
  assign n45296 = n45295 ^ n5449 ^ 1'b0 ;
  assign n45297 = n27282 & n45296 ;
  assign n45298 = ~n38929 & n45297 ;
  assign n45299 = n45298 ^ n12337 ^ 1'b0 ;
  assign n45300 = ~n2361 & n7585 ;
  assign n45301 = n21575 & n45300 ;
  assign n45302 = n35862 ^ n13751 ^ 1'b0 ;
  assign n45303 = n28827 | n45302 ;
  assign n45304 = n44587 & ~n45303 ;
  assign n45305 = n16079 ^ n1381 ^ 1'b0 ;
  assign n45306 = n11772 | n45305 ;
  assign n45307 = ~n21733 & n45306 ;
  assign n45308 = n4971 & ~n8640 ;
  assign n45309 = n45308 ^ n21163 ^ 1'b0 ;
  assign n45310 = ~n1493 & n14024 ;
  assign n45311 = n45310 ^ n20971 ^ 1'b0 ;
  assign n45312 = ( n124 & ~n13708 ) | ( n124 & n45311 ) | ( ~n13708 & n45311 ) ;
  assign n45313 = n1387 & ~n45312 ;
  assign n45314 = n1211 | n7156 ;
  assign n45315 = n42145 ^ n11429 ^ 1'b0 ;
  assign n45316 = n45314 & ~n45315 ;
  assign n45317 = n11030 & n19062 ;
  assign n45318 = n28104 ^ n20408 ^ n6296 ;
  assign n45319 = ( n11613 & ~n13303 ) | ( n11613 & n31755 ) | ( ~n13303 & n31755 ) ;
  assign n45320 = n45319 ^ n13474 ^ n344 ;
  assign n45321 = ~n36573 & n45320 ;
  assign n45322 = n12208 & n45321 ;
  assign n45323 = n16590 ^ n2662 ^ 1'b0 ;
  assign n45324 = n25370 & ~n45323 ;
  assign n45325 = n11811 & ~n29339 ;
  assign n45326 = n45325 ^ n10740 ^ 1'b0 ;
  assign n45327 = n8985 & n20148 ;
  assign n45328 = n36776 ^ n22499 ^ 1'b0 ;
  assign n45329 = n14450 & ~n34766 ;
  assign n45330 = n45329 ^ n20106 ^ 1'b0 ;
  assign n45331 = n33134 & ~n33888 ;
  assign n45332 = n8798 | n14200 ;
  assign n45333 = n6200 & n45332 ;
  assign n45334 = n23695 & ~n30809 ;
  assign n45335 = ~n45333 & n45334 ;
  assign n45336 = ( n9941 & ~n16007 ) | ( n9941 & n44582 ) | ( ~n16007 & n44582 ) ;
  assign n45337 = n41831 ^ n10065 ^ 1'b0 ;
  assign n45338 = n8507 & ~n45337 ;
  assign n45339 = n8650 & ~n44643 ;
  assign n45340 = n45339 ^ n28154 ^ 1'b0 ;
  assign n45341 = ~n11223 & n16285 ;
  assign n45342 = n2930 | n28781 ;
  assign n45343 = n3940 & ~n45342 ;
  assign n45344 = ~n45341 & n45343 ;
  assign n45345 = n25108 ^ n19360 ^ 1'b0 ;
  assign n45346 = n33752 ^ n26711 ^ 1'b0 ;
  assign n45347 = ~n5801 & n7832 ;
  assign n45348 = n12943 ^ n6275 ^ 1'b0 ;
  assign n45349 = n35057 | n45348 ;
  assign n45350 = ( n12472 & n34011 ) | ( n12472 & n45349 ) | ( n34011 & n45349 ) ;
  assign n45351 = n2693 & n27890 ;
  assign n45352 = n45351 ^ n3292 ^ 1'b0 ;
  assign n45353 = ~n1161 & n5247 ;
  assign n45354 = n41266 ^ n9083 ^ 1'b0 ;
  assign n45355 = ( n3766 & n5903 ) | ( n3766 & ~n44258 ) | ( n5903 & ~n44258 ) ;
  assign n45356 = ~n5511 & n44435 ;
  assign n45357 = n18485 ^ n17112 ^ 1'b0 ;
  assign n45358 = ~n9800 & n31977 ;
  assign n45359 = n24336 & n45358 ;
  assign n45360 = ~n31728 & n45359 ;
  assign n45361 = n1545 & ~n35929 ;
  assign n45364 = n3867 ^ n488 ^ 1'b0 ;
  assign n45362 = n12849 ^ n4423 ^ n3428 ;
  assign n45363 = n45362 ^ n12016 ^ 1'b0 ;
  assign n45365 = n45364 ^ n45363 ^ 1'b0 ;
  assign n45366 = n1734 & n1958 ;
  assign n45367 = n45366 ^ n13069 ^ 1'b0 ;
  assign n45368 = n17206 & ~n45367 ;
  assign n45369 = n12585 & n34981 ;
  assign n45370 = n400 & n758 ;
  assign n45371 = ~n45369 & n45370 ;
  assign n45372 = n25887 ^ n4834 ^ 1'b0 ;
  assign n45373 = n45372 ^ n32485 ^ 1'b0 ;
  assign n45374 = n17256 & n45373 ;
  assign n45375 = n38379 | n45374 ;
  assign n45376 = n7941 ^ n2298 ^ 1'b0 ;
  assign n45377 = ( n1927 & n3299 ) | ( n1927 & ~n45376 ) | ( n3299 & ~n45376 ) ;
  assign n45378 = ~n5539 & n25773 ;
  assign n45379 = n12868 & n45378 ;
  assign n45380 = n708 & ~n45379 ;
  assign n45381 = ~n7664 & n45380 ;
  assign n45382 = n3513 | n45381 ;
  assign n45383 = n36891 ^ n1863 ^ 1'b0 ;
  assign n45384 = n2886 & n45383 ;
  assign n45385 = n13690 & n45214 ;
  assign n45386 = n19195 ^ n734 ^ 1'b0 ;
  assign n45387 = ~n45385 & n45386 ;
  assign n45388 = n11652 ^ n2877 ^ 1'b0 ;
  assign n45389 = ~n19772 & n45388 ;
  assign n45390 = n36034 ^ n6512 ^ 1'b0 ;
  assign n45391 = n16587 & ~n45390 ;
  assign n45392 = n45391 ^ n22041 ^ 1'b0 ;
  assign n45393 = n45392 ^ n24664 ^ 1'b0 ;
  assign n45397 = n19619 ^ n19372 ^ 1'b0 ;
  assign n45398 = ~n4841 & n45397 ;
  assign n45395 = n34060 ^ n17968 ^ 1'b0 ;
  assign n45396 = n19891 & ~n45395 ;
  assign n45394 = ~n1167 & n4088 ;
  assign n45399 = n45398 ^ n45396 ^ n45394 ;
  assign n45400 = n33293 ^ n23683 ^ 1'b0 ;
  assign n45401 = n13376 & n45400 ;
  assign n45402 = ~n10749 & n24621 ;
  assign n45403 = n39219 ^ n36852 ^ 1'b0 ;
  assign n45404 = n12368 & n45403 ;
  assign n45405 = n16829 | n24838 ;
  assign n45406 = n34916 | n45405 ;
  assign n45407 = n9940 | n18665 ;
  assign n45408 = n20785 | n45407 ;
  assign n45409 = n3972 | n29915 ;
  assign n45410 = n45409 ^ n8729 ^ 1'b0 ;
  assign n45411 = ( n34222 & ~n34625 ) | ( n34222 & n45410 ) | ( ~n34625 & n45410 ) ;
  assign n45412 = n539 | n5747 ;
  assign n45413 = n11049 & ~n45412 ;
  assign n45414 = n13481 & ~n23039 ;
  assign n45416 = n33409 ^ n17482 ^ n712 ;
  assign n45417 = ~n846 & n45416 ;
  assign n45415 = n5345 & n35559 ;
  assign n45418 = n45417 ^ n45415 ^ 1'b0 ;
  assign n45419 = ( n6153 & n13109 ) | ( n6153 & ~n21679 ) | ( n13109 & ~n21679 ) ;
  assign n45420 = ~n33140 & n45419 ;
  assign n45421 = n41024 & ~n45420 ;
  assign n45422 = ~n10002 & n31401 ;
  assign n45423 = n35924 & n45422 ;
  assign n45424 = ~n4546 & n17227 ;
  assign n45425 = n45424 ^ n23541 ^ 1'b0 ;
  assign n45426 = ~n2961 & n45425 ;
  assign n45427 = ( n19329 & ~n40587 ) | ( n19329 & n45426 ) | ( ~n40587 & n45426 ) ;
  assign n45428 = ~n6430 & n13480 ;
  assign n45429 = n790 & ~n40286 ;
  assign n45430 = n45428 & n45429 ;
  assign n45431 = n31 & n45430 ;
  assign n45432 = ~n35554 & n44996 ;
  assign n45433 = n15940 ^ n8284 ^ n749 ;
  assign n45434 = n14299 | n45433 ;
  assign n45435 = n35267 & n37773 ;
  assign n45436 = ~n15748 & n45435 ;
  assign n45437 = n3382 & ~n39057 ;
  assign n45438 = n2356 | n12159 ;
  assign n45439 = n2356 & ~n45438 ;
  assign n45440 = n45439 ^ n22147 ^ 1'b0 ;
  assign n45441 = n32165 ^ n25911 ^ 1'b0 ;
  assign n45442 = n45440 & ~n45441 ;
  assign n45443 = n12484 | n23541 ;
  assign n45444 = n19463 | n45443 ;
  assign n45445 = n2053 & n6280 ;
  assign n45446 = n45445 ^ n243 ^ 1'b0 ;
  assign n45447 = ~n20907 & n40094 ;
  assign n45448 = n15413 & n45447 ;
  assign n45449 = n14380 ^ n9819 ^ 1'b0 ;
  assign n45450 = n45448 | n45449 ;
  assign n45451 = n33971 ^ n30026 ^ 1'b0 ;
  assign n45452 = n34220 & n45451 ;
  assign n45453 = n18336 & n45452 ;
  assign n45454 = n40565 ^ n24853 ^ n5411 ;
  assign n45455 = n45454 ^ n22825 ^ 1'b0 ;
  assign n45456 = n6083 & ~n45455 ;
  assign n45457 = ~n21834 & n45456 ;
  assign n45458 = n24962 & n27884 ;
  assign n45459 = n41182 ^ n1055 ^ 1'b0 ;
  assign n45460 = n45458 | n45459 ;
  assign n45461 = n37846 ^ n31636 ^ 1'b0 ;
  assign n45462 = n15487 ^ n14228 ^ 1'b0 ;
  assign n45463 = n27235 & ~n45462 ;
  assign n45464 = n33345 ^ n26346 ^ 1'b0 ;
  assign n45465 = n18824 ^ n6371 ^ 1'b0 ;
  assign n45466 = n22231 & n45465 ;
  assign n45467 = n31975 ^ n2358 ^ 1'b0 ;
  assign n45468 = n765 & n12489 ;
  assign n45469 = n43042 & n45468 ;
  assign n45470 = n4085 & ~n34446 ;
  assign n45471 = n45470 ^ n4702 ^ 1'b0 ;
  assign n45472 = n21934 ^ n5362 ^ 1'b0 ;
  assign n45473 = ~n7949 & n45472 ;
  assign n45474 = n13789 ^ n6081 ^ 1'b0 ;
  assign n45475 = ~n6556 & n45474 ;
  assign n45476 = ~n29544 & n45475 ;
  assign n45477 = n45476 ^ n21366 ^ 1'b0 ;
  assign n45478 = n42770 & ~n45477 ;
  assign n45479 = ~n45473 & n45478 ;
  assign n45480 = n13561 ^ n7994 ^ 1'b0 ;
  assign n45481 = ~n2017 & n17551 ;
  assign n45482 = n45481 ^ n34569 ^ 1'b0 ;
  assign n45483 = n45480 & ~n45482 ;
  assign n45485 = n10003 ^ n7893 ^ n1994 ;
  assign n45486 = n3917 | n10150 ;
  assign n45487 = ( ~n4336 & n45485 ) | ( ~n4336 & n45486 ) | ( n45485 & n45486 ) ;
  assign n45484 = n12547 & ~n14694 ;
  assign n45488 = n45487 ^ n45484 ^ 1'b0 ;
  assign n45489 = n10185 ^ n4569 ^ 1'b0 ;
  assign n45490 = n24732 ^ n1741 ^ 1'b0 ;
  assign n45491 = n14092 & ~n27247 ;
  assign n45492 = n12432 ^ n11238 ^ 1'b0 ;
  assign n45493 = ~n34668 & n45492 ;
  assign n45494 = n20335 | n45493 ;
  assign n45495 = n23625 & ~n36396 ;
  assign n45496 = n45495 ^ n7936 ^ 1'b0 ;
  assign n45497 = n23081 | n33550 ;
  assign n45498 = n45497 ^ n10434 ^ 1'b0 ;
  assign n45499 = ~n4724 & n45498 ;
  assign n45500 = n45499 ^ n12137 ^ 1'b0 ;
  assign n45501 = n26921 ^ n17112 ^ n4092 ;
  assign n45502 = n4653 | n31006 ;
  assign n45503 = n45502 ^ n35300 ^ 1'b0 ;
  assign n45504 = n3694 & n4575 ;
  assign n45505 = n12565 & n45504 ;
  assign n45506 = n28431 & n45505 ;
  assign n45507 = n3991 | n9004 ;
  assign n45508 = n45507 ^ n6413 ^ 1'b0 ;
  assign n45509 = ~n4772 & n45508 ;
  assign n45510 = n24461 ^ n21859 ^ 1'b0 ;
  assign n45511 = n45509 & ~n45510 ;
  assign n45512 = n2172 & n45511 ;
  assign n45513 = n7448 & ~n8867 ;
  assign n45514 = n91 & n7791 ;
  assign n45515 = ~n45513 & n45514 ;
  assign n45516 = n41350 & ~n45515 ;
  assign n45517 = n43894 & n45516 ;
  assign n45518 = n9193 | n26348 ;
  assign n45519 = n45518 ^ n40763 ^ 1'b0 ;
  assign n45520 = n3442 & ~n9823 ;
  assign n45521 = ~n5671 & n16177 ;
  assign n45522 = n45520 & n45521 ;
  assign n45523 = n5872 ^ n4359 ^ 1'b0 ;
  assign n45524 = ( ~n1768 & n3583 ) | ( ~n1768 & n45523 ) | ( n3583 & n45523 ) ;
  assign n45525 = n13474 & n35425 ;
  assign n45526 = n4005 & n45525 ;
  assign n45527 = n9689 | n20906 ;
  assign n45528 = n45527 ^ n1194 ^ 1'b0 ;
  assign n45529 = n296 | n40177 ;
  assign n45530 = n8313 | n45529 ;
  assign n45531 = ~n6959 & n22298 ;
  assign n45532 = n45531 ^ n24310 ^ 1'b0 ;
  assign n45533 = n10319 ^ n8282 ^ 1'b0 ;
  assign n45534 = ~n8486 & n45533 ;
  assign n45539 = n14978 & ~n22379 ;
  assign n45536 = n4326 | n19433 ;
  assign n45535 = n220 & n7536 ;
  assign n45537 = n45536 ^ n45535 ^ 1'b0 ;
  assign n45538 = ~n16820 & n45537 ;
  assign n45540 = n45539 ^ n45538 ^ 1'b0 ;
  assign n45541 = n24982 & ~n45540 ;
  assign n45542 = n45541 ^ n6132 ^ 1'b0 ;
  assign n45543 = n7793 ^ n3146 ^ 1'b0 ;
  assign n45544 = n38787 ^ n12511 ^ n11817 ;
  assign n45545 = n20577 ^ n13981 ^ 1'b0 ;
  assign n45546 = n9421 ^ n3143 ^ 1'b0 ;
  assign n45547 = ~n19716 & n45546 ;
  assign n45548 = ~n26745 & n40896 ;
  assign n45549 = n1210 & n33483 ;
  assign n45550 = n45549 ^ n7143 ^ 1'b0 ;
  assign n45551 = n8712 & n10118 ;
  assign n45552 = n2367 | n12428 ;
  assign n45553 = n45552 ^ n1355 ^ 1'b0 ;
  assign n45554 = n45553 ^ n13393 ^ 1'b0 ;
  assign n45555 = n19784 & n45554 ;
  assign n45556 = ( n18675 & n27661 ) | ( n18675 & n27940 ) | ( n27661 & n27940 ) ;
  assign n45557 = n1329 & n29399 ;
  assign n45558 = n9559 | n39197 ;
  assign n45559 = n4238 | n10890 ;
  assign n45560 = n41846 ^ n23609 ^ n5438 ;
  assign n45561 = n45560 ^ n1450 ^ 1'b0 ;
  assign n45562 = ~n16275 & n39966 ;
  assign n45563 = n43023 ^ n9377 ^ 1'b0 ;
  assign n45564 = ~n20569 & n33162 ;
  assign n45565 = ~n12357 & n45564 ;
  assign n45566 = ( n7427 & n8281 ) | ( n7427 & n13618 ) | ( n8281 & n13618 ) ;
  assign n45568 = n6106 | n21135 ;
  assign n45569 = n45568 ^ n33187 ^ 1'b0 ;
  assign n45567 = n12082 & ~n43026 ;
  assign n45570 = n45569 ^ n45567 ^ 1'b0 ;
  assign n45571 = n340 & ~n5401 ;
  assign n45572 = n620 | n40679 ;
  assign n45573 = ~n11763 & n12592 ;
  assign n45574 = n13094 & n45573 ;
  assign n45575 = ~n2688 & n45574 ;
  assign n45576 = n40077 & ~n44355 ;
  assign n45577 = n28254 ^ n5805 ^ 1'b0 ;
  assign n45578 = n11659 & n30102 ;
  assign n45579 = n40166 ^ n25447 ^ 1'b0 ;
  assign n45580 = n6930 | n35053 ;
  assign n45581 = n45580 ^ n34044 ^ 1'b0 ;
  assign n45582 = ~n275 & n16063 ;
  assign n45583 = n9212 ^ n593 ^ 1'b0 ;
  assign n45584 = ~n5986 & n45583 ;
  assign n45585 = n45584 ^ n42508 ^ 1'b0 ;
  assign n45586 = n45582 & n45585 ;
  assign n45587 = ~n38620 & n45586 ;
  assign n45588 = n22801 & n45587 ;
  assign n45589 = n30053 ^ n21885 ^ 1'b0 ;
  assign n45590 = ~n13042 & n26971 ;
  assign n45592 = n9140 ^ n3909 ^ 1'b0 ;
  assign n45591 = n4863 & n16968 ;
  assign n45593 = n45592 ^ n45591 ^ 1'b0 ;
  assign n45594 = n26835 & n42567 ;
  assign n45595 = n15068 & n45594 ;
  assign n45596 = ~n2247 & n19669 ;
  assign n45597 = n45596 ^ n1387 ^ 1'b0 ;
  assign n45598 = n25369 & ~n32348 ;
  assign n45599 = ( n179 & n6011 ) | ( n179 & ~n26292 ) | ( n6011 & ~n26292 ) ;
  assign n45600 = n237 & n19307 ;
  assign n45601 = n45600 ^ n16230 ^ 1'b0 ;
  assign n45602 = n4148 & n5277 ;
  assign n45603 = n45602 ^ n4348 ^ 1'b0 ;
  assign n45604 = n45603 ^ n2772 ^ 1'b0 ;
  assign n45605 = n45601 & ~n45604 ;
  assign n45606 = n24862 | n40076 ;
  assign n45607 = n39706 ^ n6397 ^ 1'b0 ;
  assign n45608 = n45606 & ~n45607 ;
  assign n45613 = n24527 ^ n19076 ^ 1'b0 ;
  assign n45614 = ~n34449 & n45613 ;
  assign n45609 = n1653 & n3802 ;
  assign n45610 = n8725 & n45609 ;
  assign n45611 = n28365 & n45610 ;
  assign n45612 = n16983 & ~n45611 ;
  assign n45615 = n45614 ^ n45612 ^ 1'b0 ;
  assign n45616 = ~n6000 & n35827 ;
  assign n45617 = n1230 & ~n2902 ;
  assign n45618 = ~n14922 & n45617 ;
  assign n45619 = ~n11334 & n45618 ;
  assign n45620 = n45619 ^ n901 ^ 1'b0 ;
  assign n45621 = n18773 ^ n2604 ^ 1'b0 ;
  assign n45622 = n2389 & ~n19440 ;
  assign n45623 = n45621 & n45622 ;
  assign n45624 = n734 & n6095 ;
  assign n45625 = n45624 ^ n36179 ^ 1'b0 ;
  assign n45626 = n2835 ^ n170 ^ 1'b0 ;
  assign n45627 = n45626 ^ n26239 ^ 1'b0 ;
  assign n45628 = n11880 & n45627 ;
  assign n45629 = n11372 ^ n372 ^ 1'b0 ;
  assign n45630 = n3736 | n45629 ;
  assign n45631 = n45630 ^ n546 ^ 1'b0 ;
  assign n45632 = n5979 & n45631 ;
  assign n45633 = n16244 & n26963 ;
  assign n45634 = n700 & n45633 ;
  assign n45635 = n12022 | n45634 ;
  assign n45636 = n32736 & n45635 ;
  assign n45637 = ( ~n492 & n16669 ) | ( ~n492 & n18556 ) | ( n16669 & n18556 ) ;
  assign n45638 = ~n25138 & n45637 ;
  assign n45641 = n44568 ^ n11005 ^ 1'b0 ;
  assign n45639 = n18151 ^ n15220 ^ 1'b0 ;
  assign n45640 = ~n25619 & n45639 ;
  assign n45642 = n45641 ^ n45640 ^ n31782 ;
  assign n45643 = n20128 | n26983 ;
  assign n45644 = n30750 & n40945 ;
  assign n45645 = n10805 ^ n727 ^ 1'b0 ;
  assign n45646 = ~n1271 & n45645 ;
  assign n45647 = n7797 ^ n182 ^ 1'b0 ;
  assign n45648 = ( n9846 & n23403 ) | ( n9846 & ~n45647 ) | ( n23403 & ~n45647 ) ;
  assign n45649 = n20406 & ~n38668 ;
  assign n45650 = n45649 ^ n1714 ^ 1'b0 ;
  assign n45652 = n34639 ^ n16920 ^ n3867 ;
  assign n45651 = n7458 & ~n24283 ;
  assign n45653 = n45652 ^ n45651 ^ 1'b0 ;
  assign n45654 = n15934 ^ n9748 ^ 1'b0 ;
  assign n45655 = ~n19301 & n45654 ;
  assign n45656 = n15882 ^ n12323 ^ n6518 ;
  assign n45657 = n44776 & ~n45656 ;
  assign n45658 = n24937 ^ n13909 ^ n7729 ;
  assign n45660 = n15799 ^ n12664 ^ 1'b0 ;
  assign n45659 = n33995 & n41494 ;
  assign n45661 = n45660 ^ n45659 ^ 1'b0 ;
  assign n45662 = n19319 ^ n10883 ^ 1'b0 ;
  assign n45663 = n6290 ^ n6016 ^ 1'b0 ;
  assign n45664 = ~n5916 & n45663 ;
  assign n45665 = n7058 ^ n2803 ^ 1'b0 ;
  assign n45666 = n18106 | n45665 ;
  assign n45667 = n45666 ^ n16723 ^ 1'b0 ;
  assign n45668 = n45664 & n45667 ;
  assign n45669 = n24672 & n45668 ;
  assign n45670 = ~n19769 & n45669 ;
  assign n45671 = ( n8775 & n21373 ) | ( n8775 & n45166 ) | ( n21373 & n45166 ) ;
  assign n45672 = n7400 & n19629 ;
  assign n45673 = n45671 & n45672 ;
  assign n45674 = ~n4841 & n6866 ;
  assign n45675 = n45674 ^ n1812 ^ 1'b0 ;
  assign n45676 = ( ~n6552 & n17300 ) | ( ~n6552 & n18451 ) | ( n17300 & n18451 ) ;
  assign n45677 = n20835 ^ n16966 ^ 1'b0 ;
  assign n45678 = n21499 & ~n45677 ;
  assign n45679 = n45678 ^ n12507 ^ n1618 ;
  assign n45680 = n9268 & ~n43617 ;
  assign n45681 = n12935 & n45680 ;
  assign n45682 = n6415 | n45681 ;
  assign n45683 = n45682 ^ n35195 ^ 1'b0 ;
  assign n45684 = n19851 & n21031 ;
  assign n45685 = n5727 ^ n792 ^ 1'b0 ;
  assign n45686 = n22107 & n45685 ;
  assign n45687 = n10497 ^ n551 ^ 1'b0 ;
  assign n45688 = n26362 & ~n40813 ;
  assign n45689 = n43154 ^ n1716 ^ 1'b0 ;
  assign n45690 = n21418 | n45689 ;
  assign n45691 = n24111 & ~n40808 ;
  assign n45692 = ~n15707 & n45691 ;
  assign n45693 = n406 | n45692 ;
  assign n45694 = ~n17998 & n25635 ;
  assign n45695 = n45694 ^ n5948 ^ 1'b0 ;
  assign n45696 = n12553 & ~n40906 ;
  assign n45697 = ~n45695 & n45696 ;
  assign n45698 = n38726 ^ n15112 ^ n3181 ;
  assign n45699 = ~n16387 & n45698 ;
  assign n45700 = ~n10272 & n14402 ;
  assign n45701 = n45700 ^ n44921 ^ 1'b0 ;
  assign n45702 = n37652 & ~n45701 ;
  assign n45703 = n8283 & n17876 ;
  assign n45704 = n45703 ^ n10950 ^ 1'b0 ;
  assign n45705 = n11790 & ~n45704 ;
  assign n45706 = n7407 & ~n43111 ;
  assign n45707 = n10180 ^ n6507 ^ 1'b0 ;
  assign n45708 = ~n40946 & n45707 ;
  assign n45709 = n14360 ^ n9680 ^ n1269 ;
  assign n45710 = n39666 ^ n8989 ^ 1'b0 ;
  assign n45711 = n25156 ^ n16361 ^ n2170 ;
  assign n45712 = n4604 | n20347 ;
  assign n45713 = n532 & n1574 ;
  assign n45714 = n31559 & n45713 ;
  assign n45715 = n45714 ^ n18297 ^ 1'b0 ;
  assign n45716 = n34171 ^ n269 ^ 1'b0 ;
  assign n45717 = n1124 & n45716 ;
  assign n45718 = n43420 & n45717 ;
  assign n45719 = ~n38265 & n45718 ;
  assign n45720 = n12338 & n33572 ;
  assign n45721 = n45720 ^ n4446 ^ 1'b0 ;
  assign n45722 = n376 & n6574 ;
  assign n45723 = n37579 & n45722 ;
  assign n45724 = n45723 ^ n3034 ^ 1'b0 ;
  assign n45726 = n35468 | n40429 ;
  assign n45725 = n861 & ~n3587 ;
  assign n45727 = n45726 ^ n45725 ^ n20252 ;
  assign n45728 = n5725 & ~n24599 ;
  assign n45729 = n1459 & n45728 ;
  assign n45730 = n4666 & ~n8180 ;
  assign n45731 = ~n15822 & n45730 ;
  assign n45732 = n24290 & n45731 ;
  assign n45733 = ( ~n4962 & n40398 ) | ( ~n4962 & n41789 ) | ( n40398 & n41789 ) ;
  assign n45734 = ( n7076 & ~n13765 ) | ( n7076 & n35105 ) | ( ~n13765 & n35105 ) ;
  assign n45735 = n1077 | n3764 ;
  assign n45736 = ~n13056 & n28495 ;
  assign n45738 = ~n5893 & n11095 ;
  assign n45739 = n6949 & n45738 ;
  assign n45737 = n14350 | n16327 ;
  assign n45740 = n45739 ^ n45737 ^ 1'b0 ;
  assign n45741 = n22621 & n45740 ;
  assign n45742 = n3489 & n43215 ;
  assign n45743 = ~n91 & n2045 ;
  assign n45744 = n35311 ^ n11230 ^ 1'b0 ;
  assign n45745 = n45743 & n45744 ;
  assign n45746 = ( ~n30744 & n34852 ) | ( ~n30744 & n43591 ) | ( n34852 & n43591 ) ;
  assign n45751 = n61 | n6367 ;
  assign n45748 = ~n15694 & n28221 ;
  assign n45749 = ~n27884 & n45748 ;
  assign n45747 = ( ~n18156 & n24215 ) | ( ~n18156 & n44782 ) | ( n24215 & n44782 ) ;
  assign n45750 = n45749 ^ n45747 ^ 1'b0 ;
  assign n45752 = n45751 ^ n45750 ^ n3259 ;
  assign n45753 = ~n1385 & n25272 ;
  assign n45754 = n45753 ^ n43200 ^ 1'b0 ;
  assign n45755 = n40407 ^ n35 ^ 1'b0 ;
  assign n45756 = n6084 | n43554 ;
  assign n45757 = ~n8503 & n13708 ;
  assign n45758 = ( ~n17124 & n24518 ) | ( ~n17124 & n30637 ) | ( n24518 & n30637 ) ;
  assign n45759 = ( n25582 & n37660 ) | ( n25582 & n45758 ) | ( n37660 & n45758 ) ;
  assign n45760 = n2097 ^ n262 ^ 1'b0 ;
  assign n45761 = n12113 & n45760 ;
  assign n45762 = n15531 & n45761 ;
  assign n45763 = n13023 ^ n3121 ^ 1'b0 ;
  assign n45764 = n12881 & n37591 ;
  assign n45765 = n10146 | n32968 ;
  assign n45766 = n21042 ^ n12883 ^ 1'b0 ;
  assign n45767 = ~n45765 & n45766 ;
  assign n45769 = n27265 ^ n8230 ^ 1'b0 ;
  assign n45768 = ~n6043 & n29645 ;
  assign n45770 = n45769 ^ n45768 ^ 1'b0 ;
  assign n45771 = n6966 ^ n6468 ^ 1'b0 ;
  assign n45772 = ( ~n1189 & n1434 ) | ( ~n1189 & n7715 ) | ( n1434 & n7715 ) ;
  assign n45773 = n10069 | n45772 ;
  assign n45774 = n45771 & ~n45773 ;
  assign n45775 = ( n4302 & n4357 ) | ( n4302 & ~n45774 ) | ( n4357 & ~n45774 ) ;
  assign n45776 = n18409 ^ n2726 ^ 1'b0 ;
  assign n45777 = n17605 ^ n2796 ^ 1'b0 ;
  assign n45778 = ~n162 & n32862 ;
  assign n45779 = n45778 ^ n1050 ^ 1'b0 ;
  assign n45780 = n428 | n12050 ;
  assign n45781 = n24132 ^ n9795 ^ 1'b0 ;
  assign n45782 = ~n2048 & n43974 ;
  assign n45783 = n19323 & n45782 ;
  assign n45784 = n40783 & ~n45783 ;
  assign n45785 = n23786 & n45784 ;
  assign n45786 = n37941 | n45785 ;
  assign n45787 = n45786 ^ n24813 ^ 1'b0 ;
  assign n45788 = n12337 ^ n2361 ^ 1'b0 ;
  assign n45789 = n4336 ^ n2865 ^ 1'b0 ;
  assign n45790 = n412 & n1445 ;
  assign n45791 = ~n4244 & n45790 ;
  assign n45792 = ~n21811 & n40180 ;
  assign n45793 = n45792 ^ n30430 ^ n23302 ;
  assign n45794 = n45793 ^ n6093 ^ n4910 ;
  assign n45801 = n4969 ^ n1020 ^ 1'b0 ;
  assign n45795 = n7583 & n24454 ;
  assign n45796 = n45795 ^ n24678 ^ 1'b0 ;
  assign n45797 = ~n2367 & n45796 ;
  assign n45798 = n5375 & ~n18183 ;
  assign n45799 = ~n10970 & n45798 ;
  assign n45800 = ( n26694 & n45797 ) | ( n26694 & n45799 ) | ( n45797 & n45799 ) ;
  assign n45802 = n45801 ^ n45800 ^ 1'b0 ;
  assign n45803 = n39852 | n42006 ;
  assign n45804 = n5526 & ~n45803 ;
  assign n45805 = n37960 ^ n27623 ^ 1'b0 ;
  assign n45806 = n5867 & ~n45805 ;
  assign n45807 = n13330 ^ n12599 ^ 1'b0 ;
  assign n45808 = n14583 & n45807 ;
  assign n45809 = ~n12160 & n45808 ;
  assign n45810 = n45809 ^ n37769 ^ 1'b0 ;
  assign n45811 = n39279 ^ n7151 ^ 1'b0 ;
  assign n45812 = n3335 & n45811 ;
  assign n45813 = n19394 & ~n19792 ;
  assign n45814 = n38692 & n45813 ;
  assign n45815 = n45814 ^ n20744 ^ 1'b0 ;
  assign n45816 = n40274 | n45815 ;
  assign n45817 = n11908 & ~n20803 ;
  assign n45818 = n41260 & ~n45817 ;
  assign n45819 = n29733 ^ n3724 ^ 1'b0 ;
  assign n45820 = ( ~n15297 & n19064 ) | ( ~n15297 & n25036 ) | ( n19064 & n25036 ) ;
  assign n45821 = n3314 | n15273 ;
  assign n45822 = n7722 & ~n8190 ;
  assign n45823 = n45821 & n45822 ;
  assign n45824 = n45823 ^ n1361 ^ 1'b0 ;
  assign n45825 = n45537 & n45824 ;
  assign n45826 = n15550 & n45825 ;
  assign n45827 = ~n45820 & n45826 ;
  assign n45828 = ~n29052 & n45827 ;
  assign n45829 = n14883 ^ n3235 ^ 1'b0 ;
  assign n45830 = ~n13470 & n45829 ;
  assign n45831 = n45830 ^ n15491 ^ 1'b0 ;
  assign n45832 = n4891 | n45831 ;
  assign n45833 = n22386 | n45188 ;
  assign n45834 = n19837 ^ n6632 ^ n1396 ;
  assign n45835 = n45834 ^ n25532 ^ 1'b0 ;
  assign n45836 = n22159 & n45835 ;
  assign n45837 = n21919 & ~n23658 ;
  assign n45838 = n11759 & ~n20569 ;
  assign n45839 = n41725 | n45838 ;
  assign n45840 = n45837 & ~n45839 ;
  assign n45841 = n874 & n2368 ;
  assign n45842 = ~n19231 & n45841 ;
  assign n45843 = n9580 & ~n14320 ;
  assign n45844 = n45843 ^ n38139 ^ 1'b0 ;
  assign n45845 = n45844 ^ n18084 ^ 1'b0 ;
  assign n45846 = n6181 & ~n45845 ;
  assign n45847 = n28771 ^ n6976 ^ 1'b0 ;
  assign n45848 = n13024 | n26792 ;
  assign n45849 = n45848 ^ n3284 ^ 1'b0 ;
  assign n45850 = ( n31002 & n45847 ) | ( n31002 & ~n45849 ) | ( n45847 & ~n45849 ) ;
  assign n45851 = n43026 ^ n17723 ^ n6998 ;
  assign n45852 = n20287 ^ n15922 ^ 1'b0 ;
  assign n45853 = n15544 & ~n36156 ;
  assign n45855 = n38863 ^ n140 ^ 1'b0 ;
  assign n45856 = ~n13355 & n45855 ;
  assign n45857 = n14999 & n45856 ;
  assign n45854 = n17723 ^ n8650 ^ n7105 ;
  assign n45858 = n45857 ^ n45854 ^ 1'b0 ;
  assign n45859 = ~n2235 & n25936 ;
  assign n45860 = ~n1592 & n28138 ;
  assign n45861 = n45860 ^ n40909 ^ 1'b0 ;
  assign n45862 = n45859 & ~n45861 ;
  assign n45863 = n24391 ^ n21062 ^ 1'b0 ;
  assign n45864 = ~n21784 & n45863 ;
  assign n45865 = n17439 | n21965 ;
  assign n45866 = n31045 ^ n8559 ^ 1'b0 ;
  assign n45867 = n8815 & ~n35311 ;
  assign n45868 = n28272 ^ n7319 ^ 1'b0 ;
  assign n45869 = n30844 ^ n5080 ^ 1'b0 ;
  assign n45870 = n27723 ^ n3558 ^ 1'b0 ;
  assign n45871 = n16754 & n44436 ;
  assign n45872 = n45871 ^ n5731 ^ 1'b0 ;
  assign n45873 = n220 & ~n21302 ;
  assign n45874 = ~n45872 & n45873 ;
  assign n45875 = n45695 ^ n6949 ^ 1'b0 ;
  assign n45876 = n15198 | n45875 ;
  assign n45877 = n14460 & n20453 ;
  assign n45878 = n45877 ^ n8183 ^ 1'b0 ;
  assign n45879 = n45878 ^ n6472 ^ 1'b0 ;
  assign n45880 = n13369 & n45879 ;
  assign n45881 = n10976 & n41345 ;
  assign n45882 = n3867 & n18417 ;
  assign n45883 = n37646 & n45882 ;
  assign n45884 = n3194 ^ n2225 ^ 1'b0 ;
  assign n45885 = ~n3598 & n11194 ;
  assign n45886 = n825 & n45885 ;
  assign n45887 = n45886 ^ n17778 ^ 1'b0 ;
  assign n45888 = ( ~n22371 & n45884 ) | ( ~n22371 & n45887 ) | ( n45884 & n45887 ) ;
  assign n45889 = ( n11295 & n12677 ) | ( n11295 & n29699 ) | ( n12677 & n29699 ) ;
  assign n45890 = n105 & n160 ;
  assign n45891 = n5667 & n45890 ;
  assign n45892 = n1872 | n45891 ;
  assign n45893 = n4986 | n45892 ;
  assign n45894 = n1927 ^ n982 ^ 1'b0 ;
  assign n45895 = n25041 | n34235 ;
  assign n45896 = n45894 | n45895 ;
  assign n45897 = ( ~n45889 & n45893 ) | ( ~n45889 & n45896 ) | ( n45893 & n45896 ) ;
  assign n45898 = n38870 ^ n12405 ^ 1'b0 ;
  assign n45899 = n45897 & n45898 ;
  assign n45900 = ~n24381 & n35744 ;
  assign n45901 = n21824 ^ n3897 ^ 1'b0 ;
  assign n45902 = ( n154 & ~n423 ) | ( n154 & n2322 ) | ( ~n423 & n2322 ) ;
  assign n45903 = ~n27542 & n36480 ;
  assign n45904 = n19096 & n45903 ;
  assign n45905 = n45904 ^ n29020 ^ n2197 ;
  assign n45906 = n10354 | n18319 ;
  assign n45907 = n45906 ^ n9140 ^ 1'b0 ;
  assign n45908 = n45907 ^ n7897 ^ 1'b0 ;
  assign n45909 = n7524 & n45908 ;
  assign n45910 = n45909 ^ n12598 ^ 1'b0 ;
  assign n45911 = n2045 & ~n8743 ;
  assign n45912 = n45911 ^ n4838 ^ 1'b0 ;
  assign n45913 = n635 & ~n45912 ;
  assign n45914 = n45913 ^ n25806 ^ 1'b0 ;
  assign n45915 = n8040 & n13026 ;
  assign n45916 = n10073 | n33931 ;
  assign n45917 = n1491 & ~n45916 ;
  assign n45918 = ( n3185 & n3459 ) | ( n3185 & ~n45614 ) | ( n3459 & ~n45614 ) ;
  assign n45919 = ( n2403 & n16057 ) | ( n2403 & ~n16716 ) | ( n16057 & ~n16716 ) ;
  assign n45920 = n4694 ^ n1495 ^ 1'b0 ;
  assign n45921 = n42950 | n45920 ;
  assign n45922 = n33142 ^ n9437 ^ 1'b0 ;
  assign n45923 = n16926 & n45922 ;
  assign n45924 = ~n39229 & n45923 ;
  assign n45925 = n539 & n45924 ;
  assign n45926 = n11723 | n31897 ;
  assign n45927 = n45926 ^ n2185 ^ 1'b0 ;
  assign n45928 = n45927 ^ n36154 ^ n4234 ;
  assign n45929 = n45928 ^ n7175 ^ 1'b0 ;
  assign n45930 = n36720 | n45929 ;
  assign n45931 = n4975 | n8188 ;
  assign n45932 = n45930 & ~n45931 ;
  assign n45934 = n30443 ^ n6774 ^ n6615 ;
  assign n45935 = ( n16039 & n17408 ) | ( n16039 & ~n45934 ) | ( n17408 & ~n45934 ) ;
  assign n45933 = ~n948 & n9611 ;
  assign n45936 = n45935 ^ n45933 ^ 1'b0 ;
  assign n45937 = ~n20305 & n45936 ;
  assign n45938 = n21294 ^ n19996 ^ 1'b0 ;
  assign n45939 = n3391 & ~n45938 ;
  assign n45940 = n16562 & n26884 ;
  assign n45941 = ~n45939 & n45940 ;
  assign n45942 = ~n2101 & n28146 ;
  assign n45943 = n40503 & n45942 ;
  assign n45944 = n34751 ^ n23025 ^ 1'b0 ;
  assign n45945 = ~n26710 & n45944 ;
  assign n45946 = n32918 ^ n1542 ^ 1'b0 ;
  assign n45947 = ~n38872 & n45946 ;
  assign n45948 = n4291 ^ n2163 ^ 1'b0 ;
  assign n45949 = n4095 & n45948 ;
  assign n45950 = n38172 | n45949 ;
  assign n45951 = n23381 ^ n21514 ^ 1'b0 ;
  assign n45952 = n18964 | n27498 ;
  assign n45953 = n45952 ^ n592 ^ 1'b0 ;
  assign n45954 = n7238 & ~n45953 ;
  assign n45955 = n35367 ^ n5269 ^ 1'b0 ;
  assign n45956 = n45954 & n45955 ;
  assign n45957 = ( ~n2921 & n14106 ) | ( ~n2921 & n45956 ) | ( n14106 & n45956 ) ;
  assign n45958 = ( n26461 & n27303 ) | ( n26461 & ~n44494 ) | ( n27303 & ~n44494 ) ;
  assign n45960 = n746 & ~n3160 ;
  assign n45961 = n45960 ^ n1269 ^ 1'b0 ;
  assign n45962 = ~n32104 & n45961 ;
  assign n45959 = ~n3320 & n9232 ;
  assign n45963 = n45962 ^ n45959 ^ 1'b0 ;
  assign n45964 = n8934 & ~n14492 ;
  assign n45965 = n45964 ^ n17298 ^ 1'b0 ;
  assign n45966 = n13257 | n45965 ;
  assign n45967 = n17696 & n19769 ;
  assign n45968 = ~n41701 & n45967 ;
  assign n45969 = n2658 | n6312 ;
  assign n45970 = n1987 | n45969 ;
  assign n45971 = ~n1299 & n13484 ;
  assign n45972 = ( n3939 & n45970 ) | ( n3939 & n45971 ) | ( n45970 & n45971 ) ;
  assign n45974 = ~n6552 & n25871 ;
  assign n45973 = n1511 & n4583 ;
  assign n45975 = n45974 ^ n45973 ^ 1'b0 ;
  assign n45976 = n3147 & ~n45975 ;
  assign n45977 = n45976 ^ n39039 ^ 1'b0 ;
  assign n45978 = n24505 ^ n12009 ^ 1'b0 ;
  assign n45979 = n10051 | n45978 ;
  assign n45980 = n11741 | n45979 ;
  assign n45981 = n45980 ^ n36309 ^ 1'b0 ;
  assign n45982 = n4772 | n20155 ;
  assign n45983 = n13315 ^ n1276 ^ 1'b0 ;
  assign n45984 = n30414 ^ n2966 ^ 1'b0 ;
  assign n45985 = ~n14720 & n26205 ;
  assign n45986 = n41301 & n45985 ;
  assign n45987 = n1680 | n33543 ;
  assign n45988 = n45 & ~n45987 ;
  assign n45989 = n40718 & ~n45988 ;
  assign n45990 = n2871 & n45989 ;
  assign n45991 = n45990 ^ n22201 ^ 1'b0 ;
  assign n45992 = ~n927 & n7272 ;
  assign n45993 = n45992 ^ n11965 ^ n9360 ;
  assign n45994 = ~n3811 & n16568 ;
  assign n45995 = n22971 ^ n1656 ^ 1'b0 ;
  assign n45996 = n45994 & ~n45995 ;
  assign n45997 = n16257 & ~n22935 ;
  assign n45998 = ~n12187 & n45997 ;
  assign n45999 = n43003 ^ n15161 ^ n11295 ;
  assign n46000 = n45998 & ~n45999 ;
  assign n46001 = ~n768 & n4938 ;
  assign n46002 = n10711 & n46001 ;
  assign n46003 = n18672 ^ n2602 ^ 1'b0 ;
  assign n46004 = n25195 & ~n46003 ;
  assign n46005 = ~n7078 & n46004 ;
  assign n46006 = n46002 & n46005 ;
  assign n46007 = n9063 & ~n14057 ;
  assign n46008 = ~n21926 & n46007 ;
  assign n46009 = n46006 & n46008 ;
  assign n46010 = ~n7482 & n28978 ;
  assign n46011 = n46010 ^ n21877 ^ 1'b0 ;
  assign n46012 = n11318 & ~n12248 ;
  assign n46013 = n46012 ^ n44247 ^ 1'b0 ;
  assign n46014 = ~n8491 & n9325 ;
  assign n46015 = n30725 & n46014 ;
  assign n46016 = n15511 & n46015 ;
  assign n46017 = n14464 | n15487 ;
  assign n46018 = n46017 ^ n33329 ^ 1'b0 ;
  assign n46019 = n46018 ^ n12916 ^ 1'b0 ;
  assign n46021 = n8847 & n9464 ;
  assign n46020 = n19770 & ~n19846 ;
  assign n46022 = n46021 ^ n46020 ^ 1'b0 ;
  assign n46023 = n6584 | n16568 ;
  assign n46024 = n39684 ^ n2816 ^ 1'b0 ;
  assign n46025 = n6198 & ~n18743 ;
  assign n46026 = n10111 & n46025 ;
  assign n46027 = n9196 ^ n9129 ^ 1'b0 ;
  assign n46028 = n15275 | n23274 ;
  assign n46029 = ~n37376 & n38755 ;
  assign n46030 = n11481 ^ n1128 ^ 1'b0 ;
  assign n46031 = ~n13762 & n46030 ;
  assign n46032 = n46031 ^ n27871 ^ 1'b0 ;
  assign n46033 = n13406 | n25094 ;
  assign n46034 = n3268 | n9264 ;
  assign n46035 = n46034 ^ n41233 ^ 1'b0 ;
  assign n46036 = ~n12224 & n30912 ;
  assign n46037 = n46036 ^ n32167 ^ 1'b0 ;
  assign n46038 = n19931 & n46037 ;
  assign n46039 = n46038 ^ n45928 ^ n33572 ;
  assign n46040 = n2080 & n15343 ;
  assign n46041 = n33609 ^ n26992 ^ 1'b0 ;
  assign n46042 = n46040 | n46041 ;
  assign n46043 = ~n1395 & n5183 ;
  assign n46044 = n2317 & ~n45801 ;
  assign n46045 = n46044 ^ n6074 ^ 1'b0 ;
  assign n46046 = n7457 & ~n46045 ;
  assign n46047 = ~n3216 & n46046 ;
  assign n46048 = n11439 ^ n9124 ^ 1'b0 ;
  assign n46049 = n37983 ^ n17774 ^ 1'b0 ;
  assign n46050 = n46048 & ~n46049 ;
  assign n46051 = n43579 & ~n45520 ;
  assign n46052 = n46051 ^ n14939 ^ 1'b0 ;
  assign n46053 = ( n2239 & n12185 ) | ( n2239 & ~n30723 ) | ( n12185 & ~n30723 ) ;
  assign n46054 = n46053 ^ n8150 ^ 1'b0 ;
  assign n46055 = ~n3736 & n5765 ;
  assign n46056 = n46055 ^ n10558 ^ 1'b0 ;
  assign n46057 = n35853 ^ n18064 ^ n1811 ;
  assign n46058 = n14937 ^ n12322 ^ 1'b0 ;
  assign n46059 = n38917 & n46058 ;
  assign n46060 = n15699 | n34106 ;
  assign n46061 = n14456 & ~n46060 ;
  assign n46062 = n11958 ^ n4930 ^ 1'b0 ;
  assign n46063 = n21631 & n46062 ;
  assign n46064 = n3265 ^ n1403 ^ 1'b0 ;
  assign n46065 = ~n2311 & n46064 ;
  assign n46066 = n2311 & n46065 ;
  assign n46067 = ~n3155 & n46066 ;
  assign n46068 = n46067 ^ n33705 ^ 1'b0 ;
  assign n46069 = n45071 & ~n46068 ;
  assign n46070 = n23742 ^ n2173 ^ 1'b0 ;
  assign n46071 = ~n12784 & n46070 ;
  assign n46072 = n46071 ^ n7414 ^ 1'b0 ;
  assign n46074 = n39417 ^ n26454 ^ n2649 ;
  assign n46073 = n18625 | n38356 ;
  assign n46075 = n46074 ^ n46073 ^ 1'b0 ;
  assign n46076 = n34237 ^ n28772 ^ n3545 ;
  assign n46077 = ~n7313 & n9067 ;
  assign n46078 = n5149 & n46077 ;
  assign n46079 = ~n4531 & n12456 ;
  assign n46080 = n21735 ^ n17853 ^ 1'b0 ;
  assign n46081 = n11805 ^ n3351 ^ 1'b0 ;
  assign n46082 = n46081 ^ n45542 ^ 1'b0 ;
  assign n46083 = n25595 & n28592 ;
  assign n46084 = n46083 ^ n12727 ^ 1'b0 ;
  assign n46085 = n27966 ^ n8931 ^ 1'b0 ;
  assign n46086 = n46085 ^ n35302 ^ n27330 ;
  assign n46087 = ~n13458 & n39555 ;
  assign n46088 = ~n31030 & n46087 ;
  assign n46089 = ( n6675 & ~n13251 ) | ( n6675 & n31013 ) | ( ~n13251 & n31013 ) ;
  assign n46090 = n28719 | n46089 ;
  assign n46091 = n26045 & ~n36371 ;
  assign n46092 = n29279 & n46091 ;
  assign n46093 = ~n21068 & n27454 ;
  assign n46094 = n7127 ^ n1745 ^ 1'b0 ;
  assign n46095 = n46094 ^ n38701 ^ 1'b0 ;
  assign n46096 = ( n3384 & n7651 ) | ( n3384 & n14334 ) | ( n7651 & n14334 ) ;
  assign n46097 = n45212 & ~n46096 ;
  assign n46098 = n15394 & ~n28058 ;
  assign n46099 = ~n11049 & n14315 ;
  assign n46100 = ~n1471 & n15598 ;
  assign n46101 = n46100 ^ n12673 ^ 1'b0 ;
  assign n46102 = n2223 ^ n2151 ^ 1'b0 ;
  assign n46103 = n20366 ^ n15538 ^ 1'b0 ;
  assign n46104 = n17532 ^ n1800 ^ 1'b0 ;
  assign n46105 = n46104 ^ n15707 ^ n14835 ;
  assign n46106 = n18741 ^ n16851 ^ 1'b0 ;
  assign n46107 = n46106 ^ n35906 ^ 1'b0 ;
  assign n46108 = n17986 & ~n37741 ;
  assign n46109 = n46108 ^ n19659 ^ 1'b0 ;
  assign n46110 = n21023 ^ n1644 ^ 1'b0 ;
  assign n46111 = n25871 & ~n39873 ;
  assign n46112 = n24492 & n44739 ;
  assign n46113 = n9336 & ~n14586 ;
  assign n46114 = n46113 ^ n606 ^ 1'b0 ;
  assign n46115 = n12321 & n46114 ;
  assign n46116 = ~n5655 & n46115 ;
  assign n46117 = ( ~n7663 & n14751 ) | ( ~n7663 & n46116 ) | ( n14751 & n46116 ) ;
  assign n46118 = n17432 & n38048 ;
  assign n46119 = n11644 ^ n1999 ^ 1'b0 ;
  assign n46120 = n21533 ^ n16170 ^ 1'b0 ;
  assign n46121 = ~n46119 & n46120 ;
  assign n46122 = n8761 | n12671 ;
  assign n46123 = n19691 & ~n46122 ;
  assign n46124 = ~n29146 & n44657 ;
  assign n46125 = n88 | n26066 ;
  assign n46126 = n26317 & ~n35929 ;
  assign n46127 = ~n21736 & n46126 ;
  assign n46128 = n138 & n46127 ;
  assign n46129 = n8474 & n46128 ;
  assign n46130 = n15997 & n16983 ;
  assign n46131 = n46130 ^ n37902 ^ 1'b0 ;
  assign n46132 = n46131 ^ n10315 ^ 1'b0 ;
  assign n46133 = n10825 ^ n9779 ^ 1'b0 ;
  assign n46134 = n46132 & n46133 ;
  assign n46135 = n13091 ^ n2591 ^ 1'b0 ;
  assign n46136 = n2560 | n46135 ;
  assign n46137 = n20781 ^ n5648 ^ 1'b0 ;
  assign n46138 = n46136 | n46137 ;
  assign n46139 = n26134 ^ n22626 ^ 1'b0 ;
  assign n46140 = n35427 & n46139 ;
  assign n46141 = n36302 | n42146 ;
  assign n46142 = n46141 ^ n12870 ^ 1'b0 ;
  assign n46143 = n15699 & ~n16469 ;
  assign n46144 = n46143 ^ n23693 ^ 1'b0 ;
  assign n46145 = n30770 ^ n267 ^ 1'b0 ;
  assign n46146 = n9660 ^ n6040 ^ 1'b0 ;
  assign n46147 = n46145 & ~n46146 ;
  assign n46148 = ~n8104 & n39099 ;
  assign n46149 = n1943 & ~n19797 ;
  assign n46150 = n26906 ^ n22801 ^ 1'b0 ;
  assign n46151 = n2563 & n18906 ;
  assign n46152 = n46150 & ~n46151 ;
  assign n46153 = n13623 | n15897 ;
  assign n46154 = n22002 | n46153 ;
  assign n46155 = n17249 ^ n4687 ^ 1'b0 ;
  assign n46156 = n13840 & ~n14716 ;
  assign n46157 = n1989 & n15739 ;
  assign n46158 = n46157 ^ n22178 ^ 1'b0 ;
  assign n46159 = n113 & n5290 ;
  assign n46160 = ~n1395 & n46159 ;
  assign n46161 = n46160 ^ n11813 ^ 1'b0 ;
  assign n46162 = n20492 & n46161 ;
  assign n46163 = n20740 & ~n27960 ;
  assign n46164 = ~n23677 & n46163 ;
  assign n46165 = ( n8249 & n15641 ) | ( n8249 & ~n46164 ) | ( n15641 & ~n46164 ) ;
  assign n46166 = n2934 & n5853 ;
  assign n46167 = n46166 ^ n608 ^ 1'b0 ;
  assign n46168 = ~n17560 & n46167 ;
  assign n46169 = n19972 & n46168 ;
  assign n46170 = n46169 ^ n43102 ^ n5293 ;
  assign n46171 = n11890 ^ n5246 ^ 1'b0 ;
  assign n46172 = n17745 & ~n46171 ;
  assign n46173 = n46172 ^ n38796 ^ 1'b0 ;
  assign n46174 = n2040 & n13862 ;
  assign n46175 = n46173 & n46174 ;
  assign n46176 = n13254 ^ n7969 ^ 1'b0 ;
  assign n46177 = n709 | n46176 ;
  assign n46178 = n17206 ^ n7827 ^ 1'b0 ;
  assign n46179 = n46177 | n46178 ;
  assign n46180 = n31290 ^ n8031 ^ 1'b0 ;
  assign n46181 = n9650 & n10598 ;
  assign n46182 = n40769 & n46181 ;
  assign n46183 = n12998 & n46182 ;
  assign n46184 = n35628 & ~n46183 ;
  assign n46185 = n34824 ^ n29654 ^ 1'b0 ;
  assign n46186 = n46184 & ~n46185 ;
  assign n46187 = n14357 & n14670 ;
  assign n46188 = n23822 & n46187 ;
  assign n46189 = n22173 | n46188 ;
  assign n46190 = n46189 ^ n17935 ^ 1'b0 ;
  assign n46191 = n11479 ^ n135 ^ 1'b0 ;
  assign n46192 = n4324 & n46191 ;
  assign n46193 = n46192 ^ n16106 ^ 1'b0 ;
  assign n46194 = n924 & ~n7469 ;
  assign n46195 = n227 & n46194 ;
  assign n46196 = n46195 ^ n9261 ^ 1'b0 ;
  assign n46197 = n42951 ^ n22313 ^ 1'b0 ;
  assign n46198 = ~n22577 & n46197 ;
  assign n46199 = ( n7349 & n16145 ) | ( n7349 & n18462 ) | ( n16145 & n18462 ) ;
  assign n46200 = n35449 & n46199 ;
  assign n46201 = n46200 ^ n44750 ^ 1'b0 ;
  assign n46202 = n46198 & n46201 ;
  assign n46203 = n7342 ^ n1335 ^ 1'b0 ;
  assign n46204 = n18914 | n30053 ;
  assign n46205 = n1845 | n41897 ;
  assign n46206 = n46205 ^ n8522 ^ 1'b0 ;
  assign n46207 = n46206 ^ n43272 ^ 1'b0 ;
  assign n46208 = ~n4072 & n5416 ;
  assign n46209 = n12123 & n46208 ;
  assign n46210 = n18185 ^ n4143 ^ 1'b0 ;
  assign n46211 = n39183 ^ n848 ^ 1'b0 ;
  assign n46212 = ~n17277 & n46211 ;
  assign n46213 = ~n17607 & n18788 ;
  assign n46214 = ( n39274 & n42287 ) | ( n39274 & n46213 ) | ( n42287 & n46213 ) ;
  assign n46215 = n2155 & ~n2543 ;
  assign n46216 = ( n2252 & n13863 ) | ( n2252 & ~n46215 ) | ( n13863 & ~n46215 ) ;
  assign n46217 = n37642 ^ n23018 ^ 1'b0 ;
  assign n46218 = n2022 & ~n20740 ;
  assign n46219 = n5833 & n6594 ;
  assign n46220 = ~n23963 & n46219 ;
  assign n46221 = n21791 & ~n46220 ;
  assign n46222 = n46221 ^ n31049 ^ 1'b0 ;
  assign n46227 = n1973 | n27608 ;
  assign n46228 = n46227 ^ n13470 ^ 1'b0 ;
  assign n46229 = n31496 & ~n46228 ;
  assign n46230 = n46229 ^ n17662 ^ 1'b0 ;
  assign n46223 = n3334 & ~n9904 ;
  assign n46224 = n46223 ^ n5150 ^ 1'b0 ;
  assign n46225 = n27218 | n46224 ;
  assign n46226 = ~n4289 & n46225 ;
  assign n46231 = n46230 ^ n46226 ^ 1'b0 ;
  assign n46232 = n4503 ^ n4277 ^ 1'b0 ;
  assign n46233 = ~n17087 & n46232 ;
  assign n46234 = ~n4251 & n46233 ;
  assign n46235 = n46234 ^ n39417 ^ n10378 ;
  assign n46236 = ~n261 & n27830 ;
  assign n46237 = ~n17742 & n46236 ;
  assign n46238 = n4895 & n27722 ;
  assign n46239 = ~n13600 & n46238 ;
  assign n46240 = n19756 & n26159 ;
  assign n46241 = n46239 & n46240 ;
  assign n46242 = n36147 & ~n37849 ;
  assign n46243 = n18867 ^ n716 ^ 1'b0 ;
  assign n46244 = n11165 ^ n6922 ^ 1'b0 ;
  assign n46245 = ~n11968 & n46244 ;
  assign n46246 = ( n26474 & ~n28592 ) | ( n26474 & n37567 ) | ( ~n28592 & n37567 ) ;
  assign n46247 = n4116 ^ n1941 ^ 1'b0 ;
  assign n46248 = ~n13122 & n46247 ;
  assign n46249 = n46248 ^ n23650 ^ 1'b0 ;
  assign n46250 = ~n9056 & n46249 ;
  assign n46251 = n7875 & ~n8197 ;
  assign n46252 = n3114 & ~n24389 ;
  assign n46253 = n46252 ^ n40771 ^ 1'b0 ;
  assign n46254 = n26930 | n40697 ;
  assign n46255 = n16576 ^ n5007 ^ 1'b0 ;
  assign n46256 = n19319 | n46255 ;
  assign n46257 = n1947 & n6856 ;
  assign n46258 = n13125 ^ n5854 ^ n5385 ;
  assign n46259 = n15087 & ~n46258 ;
  assign n46260 = n7923 & ~n38041 ;
  assign n46261 = n35796 ^ n13845 ^ 1'b0 ;
  assign n46262 = n22642 & ~n24616 ;
  assign n46263 = n7344 | n23521 ;
  assign n46264 = n16562 | n20923 ;
  assign n46265 = n56 & n7277 ;
  assign n46266 = n46265 ^ n26697 ^ 1'b0 ;
  assign n46267 = n3412 | n46266 ;
  assign n46268 = ~n15051 & n39784 ;
  assign n46269 = n45055 & n46268 ;
  assign n46270 = n22395 ^ n11323 ^ 1'b0 ;
  assign n46271 = ( ~n4103 & n45525 ) | ( ~n4103 & n46270 ) | ( n45525 & n46270 ) ;
  assign n46272 = n6527 & n7806 ;
  assign n46273 = ~n46271 & n46272 ;
  assign n46274 = n43896 ^ n39038 ^ 1'b0 ;
  assign n46275 = n29751 | n46274 ;
  assign n46276 = ( ~n6297 & n26990 ) | ( ~n6297 & n37973 ) | ( n26990 & n37973 ) ;
  assign n46277 = n4879 & ~n40173 ;
  assign n46278 = n7427 | n8197 ;
  assign n46279 = n18961 ^ n12725 ^ 1'b0 ;
  assign n46282 = n4090 & n17099 ;
  assign n46283 = n18918 & n46282 ;
  assign n46284 = n1047 & n46283 ;
  assign n46280 = n18548 ^ n5417 ^ n4117 ;
  assign n46281 = n14274 & ~n46280 ;
  assign n46285 = n46284 ^ n46281 ^ 1'b0 ;
  assign n46286 = ( ~n21935 & n37588 ) | ( ~n21935 & n46285 ) | ( n37588 & n46285 ) ;
  assign n46287 = n40802 ^ n17876 ^ 1'b0 ;
  assign n46288 = n10048 ^ n3034 ^ 1'b0 ;
  assign n46289 = n19911 | n46288 ;
  assign n46290 = n12551 & ~n32539 ;
  assign n46291 = n17846 & n46290 ;
  assign n46292 = n40829 ^ n1769 ^ 1'b0 ;
  assign n46293 = n35857 | n46292 ;
  assign n46295 = n15766 ^ n11521 ^ 1'b0 ;
  assign n46294 = n6320 ^ n5104 ^ 1'b0 ;
  assign n46296 = n46295 ^ n46294 ^ n16627 ;
  assign n46297 = n7568 ^ n4242 ^ 1'b0 ;
  assign n46298 = n12053 & ~n46297 ;
  assign n46299 = n46298 ^ n2671 ^ 1'b0 ;
  assign n46300 = ( n20364 & ~n35280 ) | ( n20364 & n46299 ) | ( ~n35280 & n46299 ) ;
  assign n46301 = n43689 ^ n35802 ^ 1'b0 ;
  assign n46302 = n10403 & ~n39476 ;
  assign n46303 = n11243 & ~n39216 ;
  assign n46304 = ~n46302 & n46303 ;
  assign n46305 = n6658 & n12271 ;
  assign n46306 = ~n3226 & n46305 ;
  assign n46307 = n11460 | n46306 ;
  assign n46308 = n30670 | n45590 ;
  assign n46309 = n8230 & ~n9032 ;
  assign n46310 = n13174 & ~n23018 ;
  assign n46311 = ~n25436 & n41483 ;
  assign n46312 = n18723 & n18765 ;
  assign n46313 = n43970 ^ n24494 ^ 1'b0 ;
  assign n46314 = ~n36459 & n46313 ;
  assign n46315 = n4364 | n46314 ;
  assign n46316 = n18678 & n26904 ;
  assign n46317 = n13626 & n46316 ;
  assign n46318 = n20608 ^ n10391 ^ 1'b0 ;
  assign n46319 = ~n9453 & n15557 ;
  assign n46320 = n11619 & n46319 ;
  assign n46321 = n46320 ^ n15478 ^ 1'b0 ;
  assign n46322 = ~n2583 & n12484 ;
  assign n46323 = ~n15929 & n22927 ;
  assign n46324 = n46323 ^ n20119 ^ 1'b0 ;
  assign n46325 = n30379 ^ n7458 ^ 1'b0 ;
  assign n46326 = ~n7847 & n16627 ;
  assign n46327 = n15114 ^ n10728 ^ 1'b0 ;
  assign n46328 = ( n27775 & ~n46326 ) | ( n27775 & n46327 ) | ( ~n46326 & n46327 ) ;
  assign n46329 = ( n11406 & n12516 ) | ( n11406 & ~n29035 ) | ( n12516 & ~n29035 ) ;
  assign n46330 = ( ~n19319 & n21718 ) | ( ~n19319 & n35559 ) | ( n21718 & n35559 ) ;
  assign n46331 = n9670 | n18784 ;
  assign n46332 = n1943 | n46331 ;
  assign n46333 = n28785 & ~n46332 ;
  assign n46334 = n46330 | n46333 ;
  assign n46335 = n468 & ~n46334 ;
  assign n46336 = n19293 | n24280 ;
  assign n46337 = n46336 ^ n28084 ^ 1'b0 ;
  assign n46338 = n46337 ^ n20548 ^ 1'b0 ;
  assign n46339 = ~n21509 & n46338 ;
  assign n46340 = n725 | n19456 ;
  assign n46344 = n5796 ^ n4461 ^ 1'b0 ;
  assign n46341 = n15997 ^ n1109 ^ 1'b0 ;
  assign n46342 = n32830 & ~n46341 ;
  assign n46343 = n14749 & n46342 ;
  assign n46345 = n46344 ^ n46343 ^ 1'b0 ;
  assign n46346 = n33716 ^ n14888 ^ 1'b0 ;
  assign n46347 = n21767 & ~n40015 ;
  assign n46348 = n15524 | n39199 ;
  assign n46351 = n34962 ^ n1231 ^ 1'b0 ;
  assign n46349 = n1182 | n14351 ;
  assign n46350 = n16650 | n46349 ;
  assign n46352 = n46351 ^ n46350 ^ 1'b0 ;
  assign n46353 = n34925 ^ n360 ^ 1'b0 ;
  assign n46354 = n15600 & ~n46353 ;
  assign n46355 = ~n27244 & n46354 ;
  assign n46356 = n2512 & ~n19949 ;
  assign n46357 = n37933 & n46356 ;
  assign n46358 = n23155 & ~n46357 ;
  assign n46359 = n10872 ^ n58 ^ 1'b0 ;
  assign n46360 = n45161 ^ n5864 ^ 1'b0 ;
  assign n46361 = n8570 & ~n31176 ;
  assign n46362 = ~n4224 & n19601 ;
  assign n46363 = ( ~n13695 & n14538 ) | ( ~n13695 & n46362 ) | ( n14538 & n46362 ) ;
  assign n46364 = n16180 & ~n31897 ;
  assign n46365 = n46364 ^ n12261 ^ 1'b0 ;
  assign n46366 = n20580 & ~n46365 ;
  assign n46367 = n9553 | n19038 ;
  assign n46368 = n30238 & ~n33187 ;
  assign n46369 = n1023 & n46368 ;
  assign n46372 = n39651 & ~n42554 ;
  assign n46373 = ~n30000 & n46372 ;
  assign n46370 = ~n37017 & n44407 ;
  assign n46371 = n46370 ^ n11655 ^ 1'b0 ;
  assign n46374 = n46373 ^ n46371 ^ 1'b0 ;
  assign n46376 = n10365 & ~n42035 ;
  assign n46377 = n1598 | n46376 ;
  assign n46375 = ~n9891 & n14566 ;
  assign n46378 = n46377 ^ n46375 ^ 1'b0 ;
  assign n46379 = n41534 ^ n861 ^ 1'b0 ;
  assign n46380 = ( n2621 & n5662 ) | ( n2621 & n17181 ) | ( n5662 & n17181 ) ;
  assign n46381 = n41636 ^ n20390 ^ 1'b0 ;
  assign n46382 = n4081 | n25780 ;
  assign n46383 = n7010 & ~n46382 ;
  assign n46384 = n4940 & n21636 ;
  assign n46386 = n1066 | n2306 ;
  assign n46385 = n42585 ^ n17325 ^ n3335 ;
  assign n46387 = n46386 ^ n46385 ^ n15508 ;
  assign n46391 = n25254 ^ n3441 ^ 1'b0 ;
  assign n46392 = n4857 & ~n46391 ;
  assign n46388 = n16495 ^ n16218 ^ 1'b0 ;
  assign n46389 = n5388 | n46388 ;
  assign n46390 = n35255 & ~n46389 ;
  assign n46393 = n46392 ^ n46390 ^ n22520 ;
  assign n46394 = ( ~n12781 & n19473 ) | ( ~n12781 & n20769 ) | ( n19473 & n20769 ) ;
  assign n46395 = n46394 ^ n43330 ^ 1'b0 ;
  assign n46396 = ~n3763 & n19166 ;
  assign n46397 = n12239 & n46396 ;
  assign n46398 = n1307 & ~n20140 ;
  assign n46399 = ( n886 & n8401 ) | ( n886 & ~n10799 ) | ( n8401 & ~n10799 ) ;
  assign n46400 = n1428 & ~n46399 ;
  assign n46401 = n46400 ^ n8901 ^ 1'b0 ;
  assign n46402 = ~n4612 & n35320 ;
  assign n46403 = n6937 | n46402 ;
  assign n46404 = n46403 ^ n30121 ^ 1'b0 ;
  assign n46406 = n1779 | n26712 ;
  assign n46407 = n4116 & ~n46406 ;
  assign n46408 = n9371 & n13881 ;
  assign n46409 = n46407 & n46408 ;
  assign n46410 = ( n820 & ~n16485 ) | ( n820 & n46409 ) | ( ~n16485 & n46409 ) ;
  assign n46405 = ~n25449 & n36910 ;
  assign n46411 = n46410 ^ n46405 ^ 1'b0 ;
  assign n46412 = n2552 & n39714 ;
  assign n46413 = n16223 & n46412 ;
  assign n46414 = n16068 ^ n1891 ^ 1'b0 ;
  assign n46415 = ~n16933 & n46414 ;
  assign n46416 = n17257 ^ n119 ^ 1'b0 ;
  assign n46417 = n46416 ^ n25685 ^ n23207 ;
  assign n46418 = n1724 & ~n16216 ;
  assign n46419 = ~n27979 & n46418 ;
  assign n46420 = n11176 & ~n21514 ;
  assign n46421 = n2120 & n46420 ;
  assign n46427 = n15922 & ~n25281 ;
  assign n46423 = n6474 & ~n35311 ;
  assign n46424 = n17191 & n46423 ;
  assign n46425 = n46424 ^ n18854 ^ 1'b0 ;
  assign n46426 = n22822 & n46425 ;
  assign n46422 = n13254 ^ n31 ^ 1'b0 ;
  assign n46428 = n46427 ^ n46426 ^ n46422 ;
  assign n46429 = n1060 & n3041 ;
  assign n46430 = n1251 | n25008 ;
  assign n46431 = ~n13789 & n46430 ;
  assign n46432 = n37927 ^ n3552 ^ 1'b0 ;
  assign n46434 = n33560 ^ n3333 ^ 1'b0 ;
  assign n46435 = ~n4499 & n46434 ;
  assign n46433 = n22115 & ~n41617 ;
  assign n46436 = n46435 ^ n46433 ^ 1'b0 ;
  assign n46437 = n11323 ^ n10742 ^ 1'b0 ;
  assign n46438 = ~n26991 & n46437 ;
  assign n46439 = n46438 ^ n2236 ^ 1'b0 ;
  assign n46440 = n42368 & ~n46439 ;
  assign n46441 = ~n2213 & n26099 ;
  assign n46442 = n36906 ^ n27084 ^ 1'b0 ;
  assign n46443 = n46441 & n46442 ;
  assign n46444 = n38063 ^ n23949 ^ 1'b0 ;
  assign n46445 = ~n8620 & n46444 ;
  assign n46446 = n11242 | n11616 ;
  assign n46447 = ( ~n3949 & n13270 ) | ( ~n3949 & n16548 ) | ( n13270 & n16548 ) ;
  assign n46448 = n3358 | n16342 ;
  assign n46449 = n1140 & ~n46448 ;
  assign n46450 = ~n21663 & n25708 ;
  assign n46451 = n7731 ^ n3839 ^ 1'b0 ;
  assign n46452 = n20419 & n46451 ;
  assign n46453 = ~n11636 & n21818 ;
  assign n46454 = n46453 ^ n18479 ^ 1'b0 ;
  assign n46455 = n46452 & n46454 ;
  assign n46456 = n14054 | n16336 ;
  assign n46457 = n8332 & ~n46456 ;
  assign n46458 = ( n404 & n3672 ) | ( n404 & n9783 ) | ( n3672 & n9783 ) ;
  assign n46459 = n41705 | n46458 ;
  assign n46460 = n46459 ^ n18020 ^ 1'b0 ;
  assign n46461 = ~n1893 & n21135 ;
  assign n46462 = n23969 & n43655 ;
  assign n46463 = n6758 & n42508 ;
  assign n46464 = n46463 ^ n5108 ^ 1'b0 ;
  assign n46465 = n6911 ^ n2650 ^ 1'b0 ;
  assign n46469 = ~n30752 & n32917 ;
  assign n46470 = n46469 ^ n42795 ^ 1'b0 ;
  assign n46466 = n23225 ^ n17481 ^ 1'b0 ;
  assign n46467 = n33328 & n46466 ;
  assign n46468 = n14311 & n46467 ;
  assign n46471 = n46470 ^ n46468 ^ n6445 ;
  assign n46472 = ~n6589 & n12147 ;
  assign n46473 = n6060 ^ n4142 ^ 1'b0 ;
  assign n46474 = ~n13739 & n46473 ;
  assign n46475 = n3028 & ~n4312 ;
  assign n46476 = ( ~n22389 & n30897 ) | ( ~n22389 & n46475 ) | ( n30897 & n46475 ) ;
  assign n46477 = ( n46472 & n46474 ) | ( n46472 & ~n46476 ) | ( n46474 & ~n46476 ) ;
  assign n46478 = n1014 & n8494 ;
  assign n46479 = n46478 ^ n130 ^ 1'b0 ;
  assign n46480 = n362 & ~n46479 ;
  assign n46481 = n4214 & ~n37473 ;
  assign n46482 = n46481 ^ n3012 ^ 1'b0 ;
  assign n46483 = n23775 ^ n3574 ^ 1'b0 ;
  assign n46484 = n29471 & ~n46483 ;
  assign n46485 = n40503 ^ n26902 ^ 1'b0 ;
  assign n46486 = n46484 & ~n46485 ;
  assign n46487 = n24725 ^ n13101 ^ 1'b0 ;
  assign n46488 = n21069 | n36373 ;
  assign n46489 = n12884 & n22201 ;
  assign n46490 = ~n9383 & n46489 ;
  assign n46491 = ~n325 & n11852 ;
  assign n46492 = ~n46490 & n46491 ;
  assign n46493 = n4108 | n46492 ;
  assign n46494 = n12038 | n46493 ;
  assign n46495 = n44035 ^ n11483 ^ 1'b0 ;
  assign n46496 = ~n6377 & n46495 ;
  assign n46497 = n3442 | n21548 ;
  assign n46498 = n46497 ^ n26137 ^ 1'b0 ;
  assign n46499 = n2526 & ~n46498 ;
  assign n46500 = ~n12634 & n42351 ;
  assign n46501 = ~n17140 & n46500 ;
  assign n46502 = n46501 ^ n18111 ^ 1'b0 ;
  assign n46503 = n9235 | n16619 ;
  assign n46504 = n33190 ^ n24032 ^ n6468 ;
  assign n46505 = n23879 ^ n8131 ^ 1'b0 ;
  assign n46506 = n16677 & n27353 ;
  assign n46507 = n2185 & ~n46506 ;
  assign n46508 = n46507 ^ n776 ^ 1'b0 ;
  assign n46509 = n46508 ^ n45660 ^ n24996 ;
  assign n46510 = ~n1261 & n46509 ;
  assign n46511 = n15636 ^ x7 ^ 1'b0 ;
  assign n46512 = n37781 & n46511 ;
  assign n46513 = n36519 & n39085 ;
  assign n46514 = n10948 & n46513 ;
  assign n46515 = n20620 ^ n17634 ^ 1'b0 ;
  assign n46516 = n21493 & n46515 ;
  assign n46517 = n611 | n12479 ;
  assign n46518 = n9525 & n46517 ;
  assign n46519 = n46518 ^ n8011 ^ 1'b0 ;
  assign n46520 = ~n20690 & n46519 ;
  assign n46521 = n13274 ^ n6749 ^ 1'b0 ;
  assign n46522 = ~n4399 & n46521 ;
  assign n46523 = ( ~n7162 & n15007 ) | ( ~n7162 & n46522 ) | ( n15007 & n46522 ) ;
  assign n46524 = ~n1908 & n42827 ;
  assign n46525 = n46524 ^ n31280 ^ 1'b0 ;
  assign n46526 = n7702 | n8200 ;
  assign n46527 = n39001 | n46526 ;
  assign n46528 = n14371 | n46527 ;
  assign n46529 = n34313 ^ n2202 ^ 1'b0 ;
  assign n46530 = n4570 ^ n1219 ^ 1'b0 ;
  assign n46531 = n38021 ^ n3996 ^ 1'b0 ;
  assign n46532 = n13262 & ~n46531 ;
  assign n46533 = n46532 ^ n23541 ^ 1'b0 ;
  assign n46534 = ~n1141 & n3802 ;
  assign n46537 = n16218 ^ n3082 ^ 1'b0 ;
  assign n46538 = ~n518 & n19725 ;
  assign n46539 = n46537 & n46538 ;
  assign n46535 = n1878 & n36276 ;
  assign n46536 = n21804 | n46535 ;
  assign n46540 = n46539 ^ n46536 ^ 1'b0 ;
  assign n46541 = n46540 ^ n41194 ^ 1'b0 ;
  assign n46542 = n21928 & ~n46541 ;
  assign n46543 = n26958 ^ n4321 ^ 1'b0 ;
  assign n46544 = n25588 ^ n11384 ^ n5667 ;
  assign n46545 = n23290 ^ n10437 ^ 1'b0 ;
  assign n46546 = n34384 & n46545 ;
  assign n46547 = ( n9941 & n29547 ) | ( n9941 & n46546 ) | ( n29547 & n46546 ) ;
  assign n46548 = n4267 & n10476 ;
  assign n46549 = n10556 | n38332 ;
  assign n46550 = n39498 & ~n46549 ;
  assign n46551 = n2455 & ~n3936 ;
  assign n46552 = n46551 ^ n96 ^ 1'b0 ;
  assign n46553 = n18812 | n29280 ;
  assign n46554 = n46552 & ~n46553 ;
  assign n46555 = n475 ^ n376 ^ 1'b0 ;
  assign n46556 = n9182 & ~n46555 ;
  assign n46557 = n36891 & n46556 ;
  assign n46558 = n46557 ^ n46410 ^ 1'b0 ;
  assign n46559 = ~n13162 & n16087 ;
  assign n46560 = n18277 ^ n12947 ^ 1'b0 ;
  assign n46561 = n5284 | n46560 ;
  assign n46562 = ( n1542 & ~n11714 ) | ( n1542 & n31234 ) | ( ~n11714 & n31234 ) ;
  assign n46563 = ~n3111 & n37423 ;
  assign n46564 = n983 & ~n38881 ;
  assign n46565 = n14796 & ~n46564 ;
  assign n46566 = n7257 & ~n28070 ;
  assign n46567 = n3508 & ~n20460 ;
  assign n46568 = n5263 & n10892 ;
  assign n46569 = n46567 & n46568 ;
  assign n46570 = n13670 | n30876 ;
  assign n46571 = n46569 & ~n46570 ;
  assign n46572 = n24969 ^ n15448 ^ 1'b0 ;
  assign n46573 = n37782 & n46572 ;
  assign n46574 = n39011 ^ n10372 ^ 1'b0 ;
  assign n46575 = ( n19005 & ~n46573 ) | ( n19005 & n46574 ) | ( ~n46573 & n46574 ) ;
  assign n46576 = n39873 ^ n12244 ^ 1'b0 ;
  assign n46577 = n6230 & n46576 ;
  assign n46578 = ( ~n7285 & n7534 ) | ( ~n7285 & n12654 ) | ( n7534 & n12654 ) ;
  assign n46579 = ( n30539 & n46577 ) | ( n30539 & ~n46578 ) | ( n46577 & ~n46578 ) ;
  assign n46580 = ( n4410 & n5982 ) | ( n4410 & n7948 ) | ( n5982 & n7948 ) ;
  assign n46581 = n46580 ^ n39183 ^ 1'b0 ;
  assign n46582 = n188 & ~n3985 ;
  assign n46583 = n2888 & n46582 ;
  assign n46584 = n12157 | n15261 ;
  assign n46585 = n16418 & ~n37572 ;
  assign n46586 = ~n46584 & n46585 ;
  assign n46587 = n1631 & n37213 ;
  assign n46588 = n46587 ^ n23505 ^ 1'b0 ;
  assign n46589 = n26839 & ~n33097 ;
  assign n46590 = n5001 & ~n46589 ;
  assign n46591 = n27844 ^ n1273 ^ 1'b0 ;
  assign n46592 = n12344 & n13931 ;
  assign n46599 = n10311 & ~n21744 ;
  assign n46600 = n3224 & n46599 ;
  assign n46598 = n25140 ^ n5458 ^ 1'b0 ;
  assign n46594 = n3592 & n11923 ;
  assign n46595 = n46594 ^ n35997 ^ 1'b0 ;
  assign n46596 = n12408 & ~n46595 ;
  assign n46597 = ~n39797 & n46596 ;
  assign n46601 = n46600 ^ n46598 ^ n46597 ;
  assign n46593 = n8785 | n9808 ;
  assign n46602 = n46601 ^ n46593 ^ 1'b0 ;
  assign n46603 = n13063 ^ n5785 ^ 1'b0 ;
  assign n46604 = n46603 ^ n21293 ^ n411 ;
  assign n46605 = n46604 ^ n6377 ^ 1'b0 ;
  assign n46606 = n28938 ^ n21921 ^ 1'b0 ;
  assign n46607 = n28458 & n46563 ;
  assign n46608 = n37587 & n46607 ;
  assign n46609 = n3662 & n35652 ;
  assign n46610 = n25771 & ~n46609 ;
  assign n46611 = n6551 & ~n46610 ;
  assign n46612 = n34354 ^ n25079 ^ 1'b0 ;
  assign n46613 = n19769 & ~n46612 ;
  assign n46614 = n46613 ^ n40630 ^ 1'b0 ;
  assign n46615 = n10212 ^ n6156 ^ 1'b0 ;
  assign n46616 = n5821 & ~n46615 ;
  assign n46617 = n1689 & n33441 ;
  assign n46618 = n46617 ^ n4746 ^ 1'b0 ;
  assign n46619 = n46618 ^ n19290 ^ 1'b0 ;
  assign n46620 = n2653 & ~n46619 ;
  assign n46621 = n46620 ^ n32276 ^ 1'b0 ;
  assign n46622 = n36198 ^ n6474 ^ 1'b0 ;
  assign n46623 = n229 & ~n17555 ;
  assign n46624 = n17642 | n36280 ;
  assign n46625 = ~n9055 & n19651 ;
  assign n46626 = n8031 ^ n7816 ^ 1'b0 ;
  assign n46627 = ~n46625 & n46626 ;
  assign n46628 = n11949 & ~n46627 ;
  assign n46629 = n10044 | n40820 ;
  assign n46630 = n37537 ^ n24119 ^ 1'b0 ;
  assign n46631 = n41848 ^ n6381 ^ 1'b0 ;
  assign n46632 = n17051 | n46631 ;
  assign n46633 = ~n11052 & n14863 ;
  assign n46634 = ( ~n29010 & n41056 ) | ( ~n29010 & n46633 ) | ( n41056 & n46633 ) ;
  assign n46635 = ~n8062 & n15462 ;
  assign n46636 = n46635 ^ n14658 ^ 1'b0 ;
  assign n46637 = n11563 ^ n6712 ^ 1'b0 ;
  assign n46638 = ~n11283 & n46637 ;
  assign n46639 = ~n10720 & n26750 ;
  assign n46640 = n1205 & ~n43466 ;
  assign n46641 = n46640 ^ n21317 ^ 1'b0 ;
  assign n46642 = n14315 & n20498 ;
  assign n46643 = n46642 ^ n39686 ^ 1'b0 ;
  assign n46644 = n812 | n46643 ;
  assign n46645 = n46644 ^ n43531 ^ 1'b0 ;
  assign n46646 = n6333 & n46645 ;
  assign n46647 = n18438 ^ n17243 ^ 1'b0 ;
  assign n46648 = n3006 & ~n11002 ;
  assign n46649 = n46648 ^ n12797 ^ n11556 ;
  assign n46652 = n609 & n5417 ;
  assign n46650 = n22087 ^ n982 ^ 1'b0 ;
  assign n46651 = ~n45200 & n46650 ;
  assign n46653 = n46652 ^ n46651 ^ 1'b0 ;
  assign n46654 = x11 & n11884 ;
  assign n46655 = n46654 ^ n10460 ^ 1'b0 ;
  assign n46656 = n25966 ^ n12327 ^ n2480 ;
  assign n46657 = n996 | n12976 ;
  assign n46658 = n14837 | n32069 ;
  assign n46659 = n17888 & n46658 ;
  assign n46660 = n46659 ^ n40101 ^ 1'b0 ;
  assign n46661 = n6774 ^ n6271 ^ 1'b0 ;
  assign n46662 = ~n33687 & n46661 ;
  assign n46663 = n304 | n8026 ;
  assign n46664 = n5742 & ~n46663 ;
  assign n46665 = n36544 ^ n3576 ^ n225 ;
  assign n46666 = n8926 & n9237 ;
  assign n46667 = n44777 ^ n28293 ^ n7702 ;
  assign n46668 = n1644 & n46667 ;
  assign n46669 = n3470 & n26381 ;
  assign n46670 = n46669 ^ n11249 ^ 1'b0 ;
  assign n46671 = n31476 & ~n46670 ;
  assign n46673 = n7768 & ~n8099 ;
  assign n46674 = n17982 & n46673 ;
  assign n46675 = n46674 ^ n19938 ^ 1'b0 ;
  assign n46676 = ~n3800 & n46675 ;
  assign n46677 = n46676 ^ n29950 ^ n14571 ;
  assign n46672 = ~n8166 & n40796 ;
  assign n46678 = n46677 ^ n46672 ^ 1'b0 ;
  assign n46679 = n38265 ^ n1511 ^ 1'b0 ;
  assign n46680 = n466 & n46679 ;
  assign n46681 = n269 ^ n260 ^ 1'b0 ;
  assign n46682 = n46681 ^ n45362 ^ 1'b0 ;
  assign n46683 = n9059 & ~n15230 ;
  assign n46684 = n46683 ^ n4960 ^ 1'b0 ;
  assign n46685 = n46684 ^ n8483 ^ 1'b0 ;
  assign n46686 = ~n22638 & n46685 ;
  assign n46687 = ~n30876 & n46686 ;
  assign n46689 = n12813 ^ n7454 ^ 1'b0 ;
  assign n46688 = n4737 & n8014 ;
  assign n46690 = n46689 ^ n46688 ^ 1'b0 ;
  assign n46691 = n32921 ^ n2014 ^ 1'b0 ;
  assign n46692 = n7121 & ~n46691 ;
  assign n46693 = n46692 ^ n42047 ^ 1'b0 ;
  assign n46694 = n3107 & ~n44116 ;
  assign n46695 = n10834 & ~n16088 ;
  assign n46696 = n528 & n7693 ;
  assign n46697 = ~n875 & n46696 ;
  assign n46698 = n10217 & ~n46697 ;
  assign n46699 = ~n46695 & n46698 ;
  assign n46700 = n23805 & ~n44541 ;
  assign n46701 = n367 & n46700 ;
  assign n46702 = n13015 ^ n6074 ^ 1'b0 ;
  assign n46703 = n15660 & n32475 ;
  assign n46704 = n10550 & ~n23040 ;
  assign n46705 = n10616 & ~n38724 ;
  assign n46706 = n46705 ^ n33571 ^ 1'b0 ;
  assign n46708 = ~n1050 & n12575 ;
  assign n46707 = n7814 | n24044 ;
  assign n46709 = n46708 ^ n46707 ^ 1'b0 ;
  assign n46710 = n7973 & ~n27993 ;
  assign n46711 = n46710 ^ n32702 ^ 1'b0 ;
  assign n46712 = n29496 ^ n16363 ^ 1'b0 ;
  assign n46713 = n8567 | n46712 ;
  assign n46714 = n28170 | n46713 ;
  assign n46715 = n41095 ^ n18653 ^ 1'b0 ;
  assign n46716 = n20763 ^ n13760 ^ 1'b0 ;
  assign n46717 = ~n24447 & n46716 ;
  assign n46718 = n19659 & ~n43181 ;
  assign n46719 = n46718 ^ n34125 ^ 1'b0 ;
  assign n46720 = n25917 ^ n5183 ^ 1'b0 ;
  assign n46721 = ~n39199 & n46720 ;
  assign n46722 = n19093 | n31392 ;
  assign n46723 = n20472 & ~n23042 ;
  assign n46725 = ~n6554 & n16144 ;
  assign n46726 = n3124 & n46725 ;
  assign n46727 = ~n1949 & n3848 ;
  assign n46728 = n631 & n46727 ;
  assign n46729 = n19395 & n46728 ;
  assign n46730 = ( n23806 & ~n46726 ) | ( n23806 & n46729 ) | ( ~n46726 & n46729 ) ;
  assign n46731 = n46730 ^ n592 ^ 1'b0 ;
  assign n46724 = n6428 & ~n32388 ;
  assign n46732 = n46731 ^ n46724 ^ 1'b0 ;
  assign n46733 = n31219 ^ n4411 ^ 1'b0 ;
  assign n46734 = n46552 ^ n18563 ^ n9424 ;
  assign n46735 = ( n3775 & ~n14162 ) | ( n3775 & n32071 ) | ( ~n14162 & n32071 ) ;
  assign n46736 = n31401 ^ n2853 ^ 1'b0 ;
  assign n46737 = n39194 & ~n46736 ;
  assign n46739 = n8505 & ~n27594 ;
  assign n46740 = n46739 ^ n23013 ^ 1'b0 ;
  assign n46738 = ~n3031 & n13053 ;
  assign n46741 = n46740 ^ n46738 ^ 1'b0 ;
  assign n46742 = n20338 | n43198 ;
  assign n46743 = n2779 | n46742 ;
  assign n46744 = n29327 & ~n46743 ;
  assign n46745 = n19241 & ~n46744 ;
  assign n46746 = n11650 & n19991 ;
  assign n46747 = n150 & n46746 ;
  assign n46748 = n14102 ^ n4797 ^ 1'b0 ;
  assign n46749 = ( ~n3686 & n4350 ) | ( ~n3686 & n6697 ) | ( n4350 & n6697 ) ;
  assign n46750 = n2242 | n46749 ;
  assign n46751 = n46748 & n46750 ;
  assign n46752 = n4434 & n15367 ;
  assign n46753 = n46751 & n46752 ;
  assign n46754 = n19512 ^ n15632 ^ 1'b0 ;
  assign n46755 = n21107 ^ n1497 ^ 1'b0 ;
  assign n46756 = n541 & ~n4962 ;
  assign n46757 = ~n20016 & n46756 ;
  assign n46758 = n2129 | n10572 ;
  assign n46759 = n8844 & ~n46758 ;
  assign n46760 = n46757 & n46759 ;
  assign n46761 = n10238 & n31617 ;
  assign n46762 = n25154 & ~n39630 ;
  assign n46763 = n46762 ^ n2517 ^ 1'b0 ;
  assign n46764 = n46761 | n46763 ;
  assign n46765 = n23653 & n25956 ;
  assign n46766 = n44726 ^ n27598 ^ n18676 ;
  assign n46768 = n5755 & n9276 ;
  assign n46767 = n9043 ^ n3314 ^ 1'b0 ;
  assign n46769 = n46768 ^ n46767 ^ 1'b0 ;
  assign n46770 = ~n3690 & n13929 ;
  assign n46771 = n46770 ^ n8507 ^ 1'b0 ;
  assign n46772 = n12291 & n18685 ;
  assign n46773 = ~n25604 & n46772 ;
  assign n46774 = n8945 & n26096 ;
  assign n46775 = n46774 ^ n5459 ^ 1'b0 ;
  assign n46776 = n8208 & n46775 ;
  assign n46777 = n46773 & n46776 ;
  assign n46778 = n11691 ^ n845 ^ 1'b0 ;
  assign n46779 = n7507 & ~n46778 ;
  assign n46780 = n451 | n43084 ;
  assign n46781 = n6836 | n7369 ;
  assign n46782 = n46781 ^ n26877 ^ 1'b0 ;
  assign n46783 = ~n1956 & n46782 ;
  assign n46784 = n26604 ^ n22012 ^ 1'b0 ;
  assign n46785 = n22051 ^ n11981 ^ 1'b0 ;
  assign n46786 = n20740 & n46785 ;
  assign n46787 = n7427 ^ n311 ^ 1'b0 ;
  assign n46788 = n5751 & ~n8588 ;
  assign n46789 = ~n17232 & n43729 ;
  assign n46790 = n46789 ^ n17480 ^ 1'b0 ;
  assign n46791 = n30085 ^ n5482 ^ 1'b0 ;
  assign n46792 = n17482 | n43537 ;
  assign n46797 = n3954 & ~n30517 ;
  assign n46793 = n5165 & ~n11225 ;
  assign n46794 = n7617 & n46793 ;
  assign n46795 = n46794 ^ n11359 ^ 1'b0 ;
  assign n46796 = n21386 | n46795 ;
  assign n46798 = n46797 ^ n46796 ^ n45560 ;
  assign n46799 = n26729 & ~n46798 ;
  assign n46800 = n27057 ^ n24905 ^ 1'b0 ;
  assign n46801 = n34136 ^ n9251 ^ 1'b0 ;
  assign n46802 = n14240 & ~n46801 ;
  assign n46803 = n46802 ^ n13968 ^ 1'b0 ;
  assign n46804 = n46800 & ~n46803 ;
  assign n46805 = n23948 ^ n17216 ^ 1'b0 ;
  assign n46806 = n40064 & ~n46805 ;
  assign n46807 = n7369 | n34984 ;
  assign n46808 = n46806 | n46807 ;
  assign n46809 = n5158 ^ n4805 ^ 1'b0 ;
  assign n46810 = n6996 & n46809 ;
  assign n46811 = n46810 ^ n22101 ^ 1'b0 ;
  assign n46812 = n5218 | n26890 ;
  assign n46813 = n46812 ^ n1210 ^ 1'b0 ;
  assign n46814 = n14123 ^ n11055 ^ 1'b0 ;
  assign n46815 = n1499 | n8674 ;
  assign n46816 = n8674 & ~n46815 ;
  assign n46817 = ~n19423 & n27998 ;
  assign n46818 = ~n27998 & n46817 ;
  assign n46819 = n46816 | n46818 ;
  assign n46820 = n46816 & ~n46819 ;
  assign n46821 = n5395 & n46820 ;
  assign n46822 = n7393 | n9231 ;
  assign n46823 = n7393 & ~n46822 ;
  assign n46824 = n45225 & n46823 ;
  assign n46825 = n2986 & ~n46824 ;
  assign n46826 = ~n2986 & n46825 ;
  assign n46827 = n46821 | n46826 ;
  assign n46828 = n46821 & ~n46827 ;
  assign n46829 = n28709 & n46828 ;
  assign n46830 = n42052 & ~n46829 ;
  assign n46831 = n46829 & n46830 ;
  assign n46832 = n20107 ^ n11299 ^ 1'b0 ;
  assign n46833 = ~n4313 & n46832 ;
  assign n46834 = n11689 ^ n7326 ^ n423 ;
  assign n46835 = ~n46833 & n46834 ;
  assign n46836 = n31824 ^ n704 ^ 1'b0 ;
  assign n46837 = n11055 & n46836 ;
  assign n46838 = n37801 & n46837 ;
  assign n46839 = ( ~n7369 & n24381 ) | ( ~n7369 & n31785 ) | ( n24381 & n31785 ) ;
  assign n46840 = n19172 & n23715 ;
  assign n46841 = ~n1020 & n46840 ;
  assign n46842 = n46841 ^ n36851 ^ 1'b0 ;
  assign n46843 = n37107 & n46842 ;
  assign n46844 = n3233 & n11263 ;
  assign n46845 = ~n3443 & n46844 ;
  assign n46846 = n35247 & n46845 ;
  assign n46847 = n17638 & ~n46846 ;
  assign n46848 = n46847 ^ n12243 ^ 1'b0 ;
  assign n46849 = n23451 & n45540 ;
  assign n46850 = n29156 & ~n34074 ;
  assign n46851 = ~n14360 & n46850 ;
  assign n46852 = n27463 ^ n25144 ^ 1'b0 ;
  assign n46853 = n26408 | n46852 ;
  assign n46854 = n42657 ^ n22386 ^ 1'b0 ;
  assign n46855 = n32974 & ~n46854 ;
  assign n46856 = n10630 & ~n35342 ;
  assign n46857 = n15370 & ~n34781 ;
  assign n46858 = n46857 ^ n5071 ^ 1'b0 ;
  assign n46859 = n46856 & n46858 ;
  assign n46860 = ~n16627 & n18848 ;
  assign n46861 = n46860 ^ n13385 ^ 1'b0 ;
  assign n46862 = n5541 & ~n46861 ;
  assign n46863 = n15185 | n31328 ;
  assign n46864 = n266 & ~n4634 ;
  assign n46865 = ~n17145 & n46864 ;
  assign n46866 = ( ~n3504 & n29750 ) | ( ~n3504 & n38704 ) | ( n29750 & n38704 ) ;
  assign n46867 = n46866 ^ n12623 ^ 1'b0 ;
  assign n46868 = n46865 & ~n46867 ;
  assign n46869 = n16653 ^ n10094 ^ 1'b0 ;
  assign n46870 = n45751 ^ n26949 ^ n13776 ;
  assign n46871 = n7620 | n11334 ;
  assign n46872 = n24040 & n26859 ;
  assign n46873 = n25590 ^ n1219 ^ 1'b0 ;
  assign n46874 = n38546 & ~n46873 ;
  assign n46875 = n41243 ^ n16392 ^ 1'b0 ;
  assign n46876 = n27049 & n46875 ;
  assign n46877 = n2381 ^ n700 ^ 1'b0 ;
  assign n46878 = n46877 ^ n17010 ^ 1'b0 ;
  assign n46879 = ~n9046 & n46878 ;
  assign n46881 = ( ~n3135 & n4214 ) | ( ~n3135 & n27326 ) | ( n4214 & n27326 ) ;
  assign n46880 = n630 | n11939 ;
  assign n46882 = n46881 ^ n46880 ^ 1'b0 ;
  assign n46883 = n7657 ^ n7272 ^ 1'b0 ;
  assign n46884 = n19423 ^ n14676 ^ 1'b0 ;
  assign n46885 = n21759 & n46884 ;
  assign n46886 = ( n5564 & n46883 ) | ( n5564 & n46885 ) | ( n46883 & n46885 ) ;
  assign n46887 = n20330 & ~n21306 ;
  assign n46888 = n16576 ^ n302 ^ 1'b0 ;
  assign n46889 = n15184 ^ n7579 ^ 1'b0 ;
  assign n46890 = n46888 & n46889 ;
  assign n46891 = n33677 ^ n8971 ^ 1'b0 ;
  assign n46892 = n2317 | n10107 ;
  assign n46893 = n46892 ^ n9974 ^ 1'b0 ;
  assign n46894 = ~n971 & n13691 ;
  assign n46895 = n46894 ^ n18175 ^ 1'b0 ;
  assign n46896 = n1212 & n7735 ;
  assign n46899 = ( n4572 & n12450 ) | ( n4572 & n26912 ) | ( n12450 & n26912 ) ;
  assign n46897 = n12673 | n16853 ;
  assign n46898 = n11238 | n46897 ;
  assign n46900 = n46899 ^ n46898 ^ 1'b0 ;
  assign n46901 = n28096 | n46900 ;
  assign n46902 = n46901 ^ n44445 ^ 1'b0 ;
  assign n46903 = n9319 ^ n1073 ^ 1'b0 ;
  assign n46904 = ~n5408 & n46903 ;
  assign n46905 = n2854 & ~n46904 ;
  assign n46906 = n22382 | n43071 ;
  assign n46907 = n28119 ^ n18458 ^ 1'b0 ;
  assign n46908 = n14948 | n30210 ;
  assign n46909 = ~n3417 & n3967 ;
  assign n46910 = ~n4702 & n46909 ;
  assign n46911 = n26009 & ~n46910 ;
  assign n46912 = n46908 | n46911 ;
  assign n46913 = n34163 ^ n23948 ^ 1'b0 ;
  assign n46914 = ~n9840 & n12700 ;
  assign n46915 = n46914 ^ n35444 ^ 1'b0 ;
  assign n46916 = ( n11179 & ~n26152 ) | ( n11179 & n38578 ) | ( ~n26152 & n38578 ) ;
  assign n46917 = n2424 & n27353 ;
  assign n46918 = n46917 ^ n17219 ^ 1'b0 ;
  assign n46919 = n46918 ^ n787 ^ 1'b0 ;
  assign n46920 = n46916 & ~n46919 ;
  assign n46921 = n480 | n2902 ;
  assign n46922 = n46921 ^ n42081 ^ 1'b0 ;
  assign n46923 = n16163 ^ n11795 ^ 1'b0 ;
  assign n46924 = n45102 & n46923 ;
  assign n46925 = n33778 & n46924 ;
  assign n46926 = n36803 ^ n25423 ^ 1'b0 ;
  assign n46927 = ~n46925 & n46926 ;
  assign n46929 = ~n3723 & n4556 ;
  assign n46930 = n46929 ^ n1385 ^ 1'b0 ;
  assign n46928 = n378 & ~n19201 ;
  assign n46931 = n46930 ^ n46928 ^ 1'b0 ;
  assign n46932 = n37979 ^ n37607 ^ 1'b0 ;
  assign n46933 = n6940 & ~n11908 ;
  assign n46934 = n4461 & n46933 ;
  assign n46935 = ~n5453 & n46934 ;
  assign n46936 = n43672 ^ n14210 ^ 1'b0 ;
  assign n46937 = n29909 ^ n7167 ^ 1'b0 ;
  assign n46938 = n12740 ^ n3807 ^ 1'b0 ;
  assign n46939 = n4635 & n37376 ;
  assign n46943 = ~n7149 & n9022 ;
  assign n46944 = n46943 ^ n18984 ^ 1'b0 ;
  assign n46942 = ~n4056 & n6650 ;
  assign n46940 = n9994 & ~n15262 ;
  assign n46941 = n22580 & ~n46940 ;
  assign n46945 = n46944 ^ n46942 ^ n46941 ;
  assign n46946 = n28254 ^ n1741 ^ 1'b0 ;
  assign n46947 = n28948 | n29300 ;
  assign n46948 = n46947 ^ n18909 ^ 1'b0 ;
  assign n46949 = n5722 & n46948 ;
  assign n46950 = ~n8144 & n18514 ;
  assign n46951 = n46950 ^ n16094 ^ 1'b0 ;
  assign n46952 = n7317 ^ n5418 ^ 1'b0 ;
  assign n46953 = n2854 & n46952 ;
  assign n46954 = n46953 ^ n1914 ^ 1'b0 ;
  assign n46955 = n46951 | n46954 ;
  assign n46956 = n46636 ^ n7562 ^ 1'b0 ;
  assign n46957 = n2502 & n15741 ;
  assign n46958 = n46957 ^ n19881 ^ n16301 ;
  assign n46959 = n31415 & n46958 ;
  assign n46960 = n8738 ^ n2569 ^ 1'b0 ;
  assign n46961 = n6161 & n46960 ;
  assign n46962 = n46737 & n46961 ;
  assign n46963 = ~n46959 & n46962 ;
  assign n46964 = n12192 & ~n20944 ;
  assign n46965 = n14614 ^ n13186 ^ 1'b0 ;
  assign n46966 = n6783 & ~n46965 ;
  assign n46967 = n31085 ^ n4612 ^ 1'b0 ;
  assign n46968 = n46407 ^ n17333 ^ 1'b0 ;
  assign n46969 = n32201 | n46968 ;
  assign n46970 = n12534 ^ n8055 ^ 1'b0 ;
  assign n46971 = ~n46969 & n46970 ;
  assign n46973 = n7265 ^ n7237 ^ 1'b0 ;
  assign n46972 = ~n2653 & n7546 ;
  assign n46974 = n46973 ^ n46972 ^ n18063 ;
  assign n46975 = n664 | n1269 ;
  assign n46976 = n46975 ^ n10284 ^ 1'b0 ;
  assign n46977 = ( n5176 & ~n14227 ) | ( n5176 & n18926 ) | ( ~n14227 & n18926 ) ;
  assign n46978 = ( ~n25252 & n46976 ) | ( ~n25252 & n46977 ) | ( n46976 & n46977 ) ;
  assign n46979 = ~n11411 & n41848 ;
  assign n46980 = ~n21460 & n46636 ;
  assign n46981 = n4575 ^ n774 ^ 1'b0 ;
  assign n46982 = ~n1269 & n46981 ;
  assign n46983 = n7377 | n33368 ;
  assign n46984 = n46982 | n46983 ;
  assign n46985 = n9636 | n27668 ;
  assign n46986 = n857 | n18393 ;
  assign n46987 = n2170 | n17778 ;
  assign n46988 = n311 & ~n46987 ;
  assign n46989 = n2346 & ~n46988 ;
  assign n46990 = n40795 ^ n3647 ^ 1'b0 ;
  assign n46991 = n2371 & ~n37546 ;
  assign n46992 = n46991 ^ n27050 ^ 1'b0 ;
  assign n46993 = n1814 & ~n10129 ;
  assign n46994 = ~n29686 & n46993 ;
  assign n46995 = n886 & ~n46994 ;
  assign n46996 = ~n11443 & n46995 ;
  assign n46997 = n14750 ^ n13004 ^ 1'b0 ;
  assign n46998 = n25892 ^ n564 ^ 1'b0 ;
  assign n46999 = ~n6384 & n6662 ;
  assign n47000 = n46999 ^ n25989 ^ 1'b0 ;
  assign n47001 = n19360 ^ n10828 ^ 1'b0 ;
  assign n47002 = n18261 & ~n19555 ;
  assign n47003 = ~n47001 & n47002 ;
  assign n47004 = n23614 | n47003 ;
  assign n47005 = n13852 & ~n47004 ;
  assign n47006 = ( n817 & ~n29682 ) | ( n817 & n41861 ) | ( ~n29682 & n41861 ) ;
  assign n47007 = n16215 & ~n20630 ;
  assign n47008 = n47007 ^ n2476 ^ 1'b0 ;
  assign n47009 = n15904 & ~n23281 ;
  assign n47010 = n5561 & n47009 ;
  assign n47011 = n47010 ^ n16215 ^ 1'b0 ;
  assign n47012 = n47008 & ~n47011 ;
  assign n47013 = n8776 ^ n8370 ^ x1 ;
  assign n47014 = n1109 | n2094 ;
  assign n47015 = n47013 & ~n47014 ;
  assign n47016 = n17162 ^ n3071 ^ 1'b0 ;
  assign n47018 = n21679 ^ n14651 ^ 1'b0 ;
  assign n47017 = n21183 | n29841 ;
  assign n47019 = n47018 ^ n47017 ^ 1'b0 ;
  assign n47023 = ~n1666 & n13850 ;
  assign n47020 = n171 & ~n5571 ;
  assign n47021 = n23483 & n47020 ;
  assign n47022 = n8789 | n47021 ;
  assign n47024 = n47023 ^ n47022 ^ 1'b0 ;
  assign n47025 = n20143 ^ n16047 ^ 1'b0 ;
  assign n47026 = n11954 | n47025 ;
  assign n47027 = n47026 ^ n8390 ^ 1'b0 ;
  assign n47028 = n41599 ^ n7170 ^ n6245 ;
  assign n47029 = n15058 & ~n47028 ;
  assign n47030 = n8966 | n47029 ;
  assign n47031 = n12285 ^ n6298 ^ 1'b0 ;
  assign n47032 = n47031 ^ n42429 ^ n13821 ;
  assign n47033 = n8102 ^ n6622 ^ 1'b0 ;
  assign n47034 = ~n25903 & n32038 ;
  assign n47035 = ~n47033 & n47034 ;
  assign n47036 = n16556 ^ n2163 ^ 1'b0 ;
  assign n47037 = n8944 | n14558 ;
  assign n47038 = n1907 & n9724 ;
  assign n47039 = n2771 & n47038 ;
  assign n47040 = ( n8500 & n47037 ) | ( n8500 & ~n47039 ) | ( n47037 & ~n47039 ) ;
  assign n47041 = n18469 | n47040 ;
  assign n47042 = ~n9553 & n28802 ;
  assign n47043 = n23167 ^ n13030 ^ 1'b0 ;
  assign n47044 = n4636 & ~n38930 ;
  assign n47045 = n32551 & n47044 ;
  assign n47046 = n47045 ^ n1445 ^ 1'b0 ;
  assign n47047 = n34869 ^ n13979 ^ n4629 ;
  assign n47048 = ( n7600 & ~n10322 ) | ( n7600 & n12875 ) | ( ~n10322 & n12875 ) ;
  assign n47049 = n47048 ^ n44611 ^ 1'b0 ;
  assign n47050 = ~n409 & n17809 ;
  assign n47051 = n46162 | n47050 ;
  assign n47052 = n5514 ^ n668 ^ 1'b0 ;
  assign n47053 = n23790 & n47052 ;
  assign n47054 = n5867 & n47053 ;
  assign n47055 = n47054 ^ n15332 ^ 1'b0 ;
  assign n47056 = n9925 | n33122 ;
  assign n47057 = n15909 & n47056 ;
  assign n47058 = ~n2441 & n16291 ;
  assign n47059 = n47058 ^ n44415 ^ n7953 ;
  assign n47060 = n21717 & ~n26246 ;
  assign n47061 = n47060 ^ n30102 ^ 1'b0 ;
  assign n47062 = n6234 | n44065 ;
  assign n47063 = n47062 ^ n709 ^ 1'b0 ;
  assign n47064 = n24061 ^ n9319 ^ 1'b0 ;
  assign n47065 = ~n14353 & n35339 ;
  assign n47066 = n41060 ^ n2857 ^ n749 ;
  assign n47067 = ~n1109 & n45872 ;
  assign n47068 = n47067 ^ n2532 ^ 1'b0 ;
  assign n47069 = n47068 ^ n41226 ^ 1'b0 ;
  assign n47070 = n47066 & ~n47069 ;
  assign n47071 = n21675 ^ n17352 ^ 1'b0 ;
  assign n47072 = n17213 & n47071 ;
  assign n47073 = n15024 & n43876 ;
  assign n47074 = n6479 | n14564 ;
  assign n47076 = n27754 ^ n11608 ^ 1'b0 ;
  assign n47075 = n637 & ~n39609 ;
  assign n47077 = n47076 ^ n47075 ^ 1'b0 ;
  assign n47078 = ( n47073 & ~n47074 ) | ( n47073 & n47077 ) | ( ~n47074 & n47077 ) ;
  assign n47079 = n2098 & n3105 ;
  assign n47080 = n47079 ^ n2753 ^ 1'b0 ;
  assign n47081 = n25321 ^ n8233 ^ 1'b0 ;
  assign n47082 = n20789 ^ n7284 ^ 1'b0 ;
  assign n47083 = ~n11489 & n47082 ;
  assign n47084 = n1705 & ~n47083 ;
  assign n47085 = n2981 | n47084 ;
  assign n47086 = n47081 | n47085 ;
  assign n47087 = ( n12528 & n47080 ) | ( n12528 & n47086 ) | ( n47080 & n47086 ) ;
  assign n47088 = n4376 ^ n4224 ^ 1'b0 ;
  assign n47089 = n4629 ^ n3777 ^ 1'b0 ;
  assign n47090 = n2282 | n4581 ;
  assign n47091 = n4581 & ~n47090 ;
  assign n47105 = n1182 & n4877 ;
  assign n47106 = ~n4877 & n47105 ;
  assign n47107 = n7902 & n47106 ;
  assign n47108 = n9721 & n47107 ;
  assign n47092 = ~n1205 & n1278 ;
  assign n47093 = ~n1278 & n47092 ;
  assign n47094 = n1347 & ~n47093 ;
  assign n47095 = ~n1347 & n47094 ;
  assign n47096 = n12397 | n47095 ;
  assign n47097 = n12397 & ~n47096 ;
  assign n47098 = n47097 ^ n24940 ^ 1'b0 ;
  assign n47099 = n1400 & n2051 ;
  assign n47100 = ~n7325 & n47099 ;
  assign n47101 = n5071 | n47100 ;
  assign n47102 = n47100 & ~n47101 ;
  assign n47103 = n21360 & ~n47102 ;
  assign n47104 = ~n47098 & n47103 ;
  assign n47109 = n47108 ^ n47104 ^ n20654 ;
  assign n47110 = n47091 | n47109 ;
  assign n47111 = ( ~n13580 & n33859 ) | ( ~n13580 & n36586 ) | ( n33859 & n36586 ) ;
  assign n47112 = n16846 & n22255 ;
  assign n47113 = n2478 & ~n9363 ;
  assign n47114 = ~n16291 & n47113 ;
  assign n47115 = ~n21009 & n47114 ;
  assign n47116 = n33668 ^ n6201 ^ 1'b0 ;
  assign n47117 = n8516 & ~n10403 ;
  assign n47118 = ~n3383 & n47117 ;
  assign n47119 = n24830 ^ n11434 ^ 1'b0 ;
  assign n47120 = n47118 | n47119 ;
  assign n47121 = ~n3831 & n12082 ;
  assign n47122 = ~n1935 & n2230 ;
  assign n47123 = n47122 ^ n12726 ^ 1'b0 ;
  assign n47124 = n47123 ^ n43076 ^ n14416 ;
  assign n47125 = n47124 ^ n2560 ^ 1'b0 ;
  assign n47126 = ~n6111 & n8016 ;
  assign n47127 = n6102 | n8040 ;
  assign n47128 = n47127 ^ n34702 ^ 1'b0 ;
  assign n47129 = n47128 ^ n45052 ^ n42942 ;
  assign n47130 = ~n3347 & n15275 ;
  assign n47131 = ~n404 & n1403 ;
  assign n47132 = n47131 ^ n47037 ^ 1'b0 ;
  assign n47133 = n10403 | n47132 ;
  assign n47134 = n2248 | n47133 ;
  assign n47135 = n3314 ^ n553 ^ 1'b0 ;
  assign n47136 = ~n3369 & n47135 ;
  assign n47137 = n37412 | n47136 ;
  assign n47138 = n6628 & n20393 ;
  assign n47139 = n47138 ^ n45559 ^ 1'b0 ;
  assign n47140 = ~n3039 & n11551 ;
  assign n47141 = n34138 ^ n16596 ^ 1'b0 ;
  assign n47142 = ~n47140 & n47141 ;
  assign n47143 = n19196 ^ n7904 ^ 1'b0 ;
  assign n47144 = ( ~n3781 & n45487 ) | ( ~n3781 & n47143 ) | ( n45487 & n47143 ) ;
  assign n47145 = n42833 ^ n13753 ^ 1'b0 ;
  assign n47146 = ~n11723 & n16012 ;
  assign n47147 = ~n7704 & n47146 ;
  assign n47148 = n3583 & ~n47147 ;
  assign n47149 = n42186 | n47148 ;
  assign n47150 = n3989 & ~n7542 ;
  assign n47151 = n47150 ^ n9772 ^ 1'b0 ;
  assign n47152 = ~n1066 & n28117 ;
  assign n47153 = n5604 & n47152 ;
  assign n47154 = n4634 ^ n1233 ^ 1'b0 ;
  assign n47155 = ~n47153 & n47154 ;
  assign n47156 = n18677 ^ n13363 ^ 1'b0 ;
  assign n47157 = n44082 | n47156 ;
  assign n47158 = n19362 & n34416 ;
  assign n47159 = n20577 ^ n14153 ^ 1'b0 ;
  assign n47160 = n8265 ^ n7547 ^ n4169 ;
  assign n47161 = ~n11469 & n47160 ;
  assign n47162 = n9291 ^ n1605 ^ 1'b0 ;
  assign n47163 = n47162 ^ n44662 ^ n1812 ;
  assign n47164 = n10753 & ~n23013 ;
  assign n47165 = n3445 | n20523 ;
  assign n47166 = n47165 ^ n39022 ^ n13346 ;
  assign n47167 = n5458 & ~n30202 ;
  assign n47168 = ~n47166 & n47167 ;
  assign n47169 = n39706 ^ n4273 ^ 1'b0 ;
  assign n47170 = n13055 | n47169 ;
  assign n47174 = n25321 ^ n14805 ^ 1'b0 ;
  assign n47173 = ~n3397 & n15578 ;
  assign n47175 = n47174 ^ n47173 ^ 1'b0 ;
  assign n47171 = n11839 | n40908 ;
  assign n47172 = n17463 & n47171 ;
  assign n47176 = n47175 ^ n47172 ^ 1'b0 ;
  assign n47177 = n6023 | n7802 ;
  assign n47178 = n7963 | n47177 ;
  assign n47179 = n23272 ^ n14027 ^ 1'b0 ;
  assign n47180 = ( n7312 & n27099 ) | ( n7312 & ~n30353 ) | ( n27099 & ~n30353 ) ;
  assign n47181 = n3003 & ~n31026 ;
  assign n47182 = n47181 ^ n32833 ^ 1'b0 ;
  assign n47183 = n21857 & n47182 ;
  assign n47184 = ~n21152 & n45751 ;
  assign n47185 = n47184 ^ n33205 ^ 1'b0 ;
  assign n47186 = n47185 ^ n3058 ^ 1'b0 ;
  assign n47187 = n25704 & n47186 ;
  assign n47188 = n42010 & n47187 ;
  assign n47189 = n15781 & n30389 ;
  assign n47190 = n47189 ^ n20050 ^ 1'b0 ;
  assign n47191 = n12786 & ~n16087 ;
  assign n47192 = ~n47190 & n47191 ;
  assign n47193 = n17871 ^ n4636 ^ 1'b0 ;
  assign n47194 = n16308 | n47193 ;
  assign n47195 = ~n16359 & n25207 ;
  assign n47196 = n44804 ^ n2658 ^ 1'b0 ;
  assign n47197 = n29452 & ~n47196 ;
  assign n47198 = n3517 & n47197 ;
  assign n47199 = ( n7604 & ~n15088 ) | ( n7604 & n15571 ) | ( ~n15088 & n15571 ) ;
  assign n47200 = n47199 ^ n6084 ^ 1'b0 ;
  assign n47201 = n16683 ^ n12696 ^ 1'b0 ;
  assign n47202 = n11059 & ~n42408 ;
  assign n47203 = n47202 ^ n14948 ^ 1'b0 ;
  assign n47204 = n17364 ^ n6447 ^ 1'b0 ;
  assign n47205 = ~n36082 & n41843 ;
  assign n47206 = ~n19245 & n32805 ;
  assign n47207 = ~n22209 & n47206 ;
  assign n47208 = n47207 ^ n6943 ^ 1'b0 ;
  assign n47209 = n47208 ^ n33145 ^ 1'b0 ;
  assign n47210 = n3753 ^ n3554 ^ 1'b0 ;
  assign n47211 = n7485 & ~n47210 ;
  assign n47212 = n7816 & ~n47211 ;
  assign n47213 = n6048 & n47212 ;
  assign n47214 = n47213 ^ n29834 ^ n10681 ;
  assign n47215 = ~n10225 & n37769 ;
  assign n47216 = n47215 ^ n4267 ^ n1736 ;
  assign n47217 = n33483 & ~n47216 ;
  assign n47218 = ~n26906 & n47217 ;
  assign n47219 = ~n29709 & n40876 ;
  assign n47220 = n6751 | n33783 ;
  assign n47221 = n4461 | n47220 ;
  assign n47222 = n14675 & n17294 ;
  assign n47223 = n28157 & n47222 ;
  assign n47224 = n3576 | n26890 ;
  assign n47225 = n3331 | n47224 ;
  assign n47226 = n135 & n39484 ;
  assign n47227 = n24489 | n47226 ;
  assign n47228 = n10129 ^ n6145 ^ 1'b0 ;
  assign n47229 = ( n6748 & n26730 ) | ( n6748 & n47228 ) | ( n26730 & n47228 ) ;
  assign n47230 = n47227 & n47229 ;
  assign n47235 = n934 | n1962 ;
  assign n47234 = n500 & ~n44074 ;
  assign n47236 = n47235 ^ n47234 ^ 1'b0 ;
  assign n47237 = n18445 & n47236 ;
  assign n47232 = ~n1550 & n37625 ;
  assign n47231 = n12139 & n30786 ;
  assign n47233 = n47232 ^ n47231 ^ n32262 ;
  assign n47238 = n47237 ^ n47233 ^ 1'b0 ;
  assign n47239 = n35459 ^ n7628 ^ 1'b0 ;
  assign n47240 = n14242 & n47239 ;
  assign n47241 = ~n33350 & n47240 ;
  assign n47242 = n28767 ^ n27527 ^ 1'b0 ;
  assign n47243 = n5995 ^ n647 ^ 1'b0 ;
  assign n47244 = ~n433 & n47243 ;
  assign n47245 = n11233 & n47244 ;
  assign n47247 = n1588 & n37089 ;
  assign n47248 = n47247 ^ n2849 ^ 1'b0 ;
  assign n47246 = n6524 & n23606 ;
  assign n47249 = n47248 ^ n47246 ^ 1'b0 ;
  assign n47250 = ~n10743 & n17608 ;
  assign n47251 = ~n45116 & n47250 ;
  assign n47252 = n30414 ^ n733 ^ 1'b0 ;
  assign n47253 = n15432 & n18135 ;
  assign n47254 = n2322 ^ n1491 ^ 1'b0 ;
  assign n47255 = ~n39246 & n44722 ;
  assign n47256 = ~n9765 & n11849 ;
  assign n47257 = ~n20289 & n26859 ;
  assign n47258 = ~n47256 & n47257 ;
  assign n47259 = n40375 ^ n1902 ^ 1'b0 ;
  assign n47260 = n45589 ^ n2885 ^ 1'b0 ;
  assign n47261 = n14343 ^ n158 ^ 1'b0 ;
  assign n47262 = n37882 ^ n31422 ^ n10147 ;
  assign n47263 = n47262 ^ n14378 ^ n8761 ;
  assign n47264 = n31345 ^ n20665 ^ 1'b0 ;
  assign n47265 = ~n11564 & n19647 ;
  assign n47266 = ~n44472 & n47265 ;
  assign n47267 = n39193 ^ n3772 ^ 1'b0 ;
  assign n47268 = n44353 & ~n47267 ;
  assign n47269 = n3777 & n18920 ;
  assign n47270 = n47269 ^ n18918 ^ 1'b0 ;
  assign n47271 = n835 & n11377 ;
  assign n47272 = ~n30459 & n47271 ;
  assign n47273 = ( n2515 & ~n7185 ) | ( n2515 & n12740 ) | ( ~n7185 & n12740 ) ;
  assign n47274 = n10855 | n18305 ;
  assign n47275 = n47274 ^ n11834 ^ 1'b0 ;
  assign n47276 = n29744 ^ n8715 ^ 1'b0 ;
  assign n47277 = n7818 | n47276 ;
  assign n47278 = n14242 ^ n588 ^ 1'b0 ;
  assign n47279 = n44955 | n47278 ;
  assign n47280 = n3600 | n21795 ;
  assign n47281 = n31777 ^ n11264 ^ 1'b0 ;
  assign n47282 = ( n9964 & ~n27222 ) | ( n9964 & n46625 ) | ( ~n27222 & n46625 ) ;
  assign n47283 = n47282 ^ n41746 ^ 1'b0 ;
  assign n47284 = n9787 & ~n25646 ;
  assign n47285 = n5010 | n6431 ;
  assign n47286 = n24139 ^ n8664 ^ 1'b0 ;
  assign n47287 = n14342 | n23620 ;
  assign n47288 = n39045 ^ n22751 ^ 1'b0 ;
  assign n47289 = n17256 & ~n47288 ;
  assign n47290 = ( n3449 & n13743 ) | ( n3449 & n46930 ) | ( n13743 & n46930 ) ;
  assign n47291 = n30993 ^ n24581 ^ n22181 ;
  assign n47292 = n20236 ^ n15076 ^ 1'b0 ;
  assign n47293 = n11855 ^ n1538 ^ 1'b0 ;
  assign n47294 = n47292 | n47293 ;
  assign n47295 = n12817 & ~n34412 ;
  assign n47296 = n16406 ^ n13605 ^ n1407 ;
  assign n47297 = ~n685 & n18059 ;
  assign n47298 = n47296 & n47297 ;
  assign n47299 = n1295 & ~n47298 ;
  assign n47300 = ~n17036 & n32923 ;
  assign n47301 = ~n29997 & n47300 ;
  assign n47302 = n4746 & ~n5541 ;
  assign n47303 = ~n3573 & n36694 ;
  assign n47304 = n2828 & n47303 ;
  assign n47305 = n12636 | n36225 ;
  assign n47306 = n29964 & n33761 ;
  assign n47307 = n47306 ^ n16751 ^ 1'b0 ;
  assign n47308 = n2822 & ~n34567 ;
  assign n47309 = n47308 ^ n9330 ^ n49 ;
  assign n47310 = ~n8997 & n19060 ;
  assign n47311 = n47310 ^ n31404 ^ 1'b0 ;
  assign n47312 = ( ~n4438 & n16673 ) | ( ~n4438 & n41764 ) | ( n16673 & n41764 ) ;
  assign n47313 = n2421 | n31487 ;
  assign n47314 = n3198 & ~n47313 ;
  assign n47315 = ~n23484 & n26906 ;
  assign n47316 = n47314 & n47315 ;
  assign n47317 = n10103 & ~n47316 ;
  assign n47318 = n12402 & n47317 ;
  assign n47320 = n17639 ^ n3324 ^ 1'b0 ;
  assign n47319 = n36516 | n44477 ;
  assign n47321 = n47320 ^ n47319 ^ 1'b0 ;
  assign n47322 = n9403 ^ n1645 ^ n1152 ;
  assign n47323 = ~n22574 & n47322 ;
  assign n47324 = n4805 & ~n47323 ;
  assign n47325 = n3334 & ~n9542 ;
  assign n47326 = ~n10477 & n47325 ;
  assign n47327 = ~n47324 & n47326 ;
  assign n47328 = ~n546 & n1104 ;
  assign n47329 = n47328 ^ n45534 ^ 1'b0 ;
  assign n47330 = n43716 ^ n23767 ^ 1'b0 ;
  assign n47331 = n47329 | n47330 ;
  assign n47332 = n37960 | n40571 ;
  assign n47333 = n3818 & ~n7632 ;
  assign n47334 = n15263 & n23483 ;
  assign n47335 = n8918 & n20872 ;
  assign n47336 = ~n37444 & n37640 ;
  assign n47337 = n19669 & n36866 ;
  assign n47338 = n47337 ^ n44350 ^ 1'b0 ;
  assign n47339 = n5151 & ~n11485 ;
  assign n47340 = n4636 & ~n20737 ;
  assign n47341 = n6628 & ~n47340 ;
  assign n47342 = ~n684 & n47341 ;
  assign n47343 = n22477 ^ n10888 ^ n9913 ;
  assign n47344 = n21266 | n47343 ;
  assign n47345 = n40325 ^ n4433 ^ n488 ;
  assign n47346 = n47345 ^ n8603 ^ 1'b0 ;
  assign n47347 = ~n3181 & n47346 ;
  assign n47348 = n47347 ^ n34081 ^ 1'b0 ;
  assign n47349 = n7623 | n15036 ;
  assign n47350 = n47349 ^ n30361 ^ 1'b0 ;
  assign n47351 = n47350 ^ n9787 ^ n251 ;
  assign n47352 = n34280 ^ n22073 ^ 1'b0 ;
  assign n47353 = n31915 | n47352 ;
  assign n47354 = n25511 & ~n47353 ;
  assign n47355 = ~n35790 & n38329 ;
  assign n47356 = n47355 ^ n45272 ^ 1'b0 ;
  assign n47358 = n47040 ^ n5071 ^ n1313 ;
  assign n47357 = n10967 & ~n33414 ;
  assign n47359 = n47358 ^ n47357 ^ 1'b0 ;
  assign n47360 = n33025 ^ n15086 ^ 1'b0 ;
  assign n47361 = n40175 | n47360 ;
  assign n47362 = n20988 ^ n6869 ^ 1'b0 ;
  assign n47363 = ~n47361 & n47362 ;
  assign n47364 = n47153 ^ n21456 ^ 1'b0 ;
  assign n47365 = n17836 | n47364 ;
  assign n47366 = n1157 & ~n47365 ;
  assign n47367 = n30008 ^ n12589 ^ 1'b0 ;
  assign n47368 = n47367 ^ n25885 ^ 1'b0 ;
  assign n47369 = n2405 | n6981 ;
  assign n47370 = n2991 & n41219 ;
  assign n47371 = ~n21490 & n47370 ;
  assign n47372 = n19281 & ~n47371 ;
  assign n47373 = n47372 ^ n3527 ^ 1'b0 ;
  assign n47374 = n13234 | n47373 ;
  assign n47375 = n47369 | n47374 ;
  assign n47376 = n1778 & n41797 ;
  assign n47377 = n13388 & n47376 ;
  assign n47378 = ~n2713 & n4913 ;
  assign n47379 = n47378 ^ n8547 ^ 1'b0 ;
  assign n47380 = n7695 | n47379 ;
  assign n47381 = ( n18429 & ~n43935 ) | ( n18429 & n47380 ) | ( ~n43935 & n47380 ) ;
  assign n47382 = n724 | n32883 ;
  assign n47383 = n47382 ^ n10979 ^ 1'b0 ;
  assign n47384 = n20971 ^ n6464 ^ 1'b0 ;
  assign n47385 = n47383 & ~n47384 ;
  assign n47386 = n9117 ^ n1542 ^ 1'b0 ;
  assign n47387 = n20359 | n47386 ;
  assign n47388 = ~n2643 & n4559 ;
  assign n47389 = ~n4559 & n47388 ;
  assign n47390 = n14182 & ~n47389 ;
  assign n47391 = n3023 & n42769 ;
  assign n47392 = ~n47390 & n47391 ;
  assign n47393 = ~n7475 & n47392 ;
  assign n47394 = n3272 | n6290 ;
  assign n47395 = n29353 ^ n11666 ^ 1'b0 ;
  assign n47396 = n24553 & n47395 ;
  assign n47397 = n1546 & n41393 ;
  assign n47398 = ~n4538 & n5184 ;
  assign n47399 = n47398 ^ n5728 ^ 1'b0 ;
  assign n47400 = n12725 & ~n15760 ;
  assign n47401 = ( n35504 & n47399 ) | ( n35504 & n47400 ) | ( n47399 & n47400 ) ;
  assign n47402 = n14937 & n35485 ;
  assign n47403 = n11407 & n47402 ;
  assign n47404 = ~n20724 & n23692 ;
  assign n47405 = n47404 ^ n22689 ^ 1'b0 ;
  assign n47406 = n9404 & n47405 ;
  assign n47407 = n47406 ^ n34311 ^ 1'b0 ;
  assign n47408 = ~n28491 & n35562 ;
  assign n47409 = n47408 ^ n33948 ^ 1'b0 ;
  assign n47410 = n5864 & ~n10499 ;
  assign n47411 = n47410 ^ n31092 ^ 1'b0 ;
  assign n47412 = n13008 ^ n7804 ^ 1'b0 ;
  assign n47413 = n12233 ^ n671 ^ 1'b0 ;
  assign n47414 = n2029 & n47413 ;
  assign n47415 = n47414 ^ n9984 ^ 1'b0 ;
  assign n47416 = n47415 ^ n8355 ^ 1'b0 ;
  assign n47417 = ~n2363 & n47416 ;
  assign n47418 = n47417 ^ n17281 ^ 1'b0 ;
  assign n47419 = n6500 & n16689 ;
  assign n47420 = n39219 & n47419 ;
  assign n47427 = ~n18626 & n19182 ;
  assign n47428 = n47427 ^ n16142 ^ 1'b0 ;
  assign n47424 = n1525 | n20965 ;
  assign n47423 = n16039 | n28137 ;
  assign n47425 = n47424 ^ n47423 ^ 1'b0 ;
  assign n47421 = n10076 & ~n20341 ;
  assign n47422 = n1385 | n47421 ;
  assign n47426 = n47425 ^ n47422 ^ 1'b0 ;
  assign n47429 = n47428 ^ n47426 ^ 1'b0 ;
  assign n47430 = n19400 ^ n12638 ^ 1'b0 ;
  assign n47431 = n47429 | n47430 ;
  assign n47432 = n18255 & ~n22837 ;
  assign n47433 = ~n16777 & n22963 ;
  assign n47434 = n3703 & ~n4070 ;
  assign n47435 = n38524 & n47434 ;
  assign n47436 = n47435 ^ n35637 ^ 1'b0 ;
  assign n47437 = n4948 & n43924 ;
  assign n47438 = n33384 ^ n15544 ^ 1'b0 ;
  assign n47439 = n24167 ^ n14419 ^ 1'b0 ;
  assign n47440 = n3390 & n13146 ;
  assign n47441 = n47440 ^ n38495 ^ 1'b0 ;
  assign n47442 = ~n1677 & n4665 ;
  assign n47443 = n1677 & n47442 ;
  assign n47444 = n492 & ~n523 ;
  assign n47445 = n523 & n47444 ;
  assign n47446 = n2749 & ~n47445 ;
  assign n47447 = n47445 & n47446 ;
  assign n47448 = n47443 | n47447 ;
  assign n47449 = n35853 & ~n47448 ;
  assign n47450 = n47448 & n47449 ;
  assign n47451 = n23023 & ~n30694 ;
  assign n47452 = n1229 & n47451 ;
  assign n47453 = ~n47451 & n47452 ;
  assign n47454 = n47453 ^ n6794 ^ 1'b0 ;
  assign n47455 = ~n3386 & n47454 ;
  assign n47456 = n47450 & n47455 ;
  assign n47457 = n47456 ^ n20556 ^ n17428 ;
  assign n47458 = n4038 & ~n30004 ;
  assign n47459 = n47458 ^ n12805 ^ 1'b0 ;
  assign n47460 = ( n892 & n6149 ) | ( n892 & n47459 ) | ( n6149 & n47459 ) ;
  assign n47461 = n6088 | n10454 ;
  assign n47462 = n5753 & n47461 ;
  assign n47463 = ~n6149 & n47462 ;
  assign n47464 = n39654 ^ n34445 ^ 1'b0 ;
  assign n47465 = n4081 & ~n47464 ;
  assign n47466 = n32789 ^ n12986 ^ n6854 ;
  assign n47467 = n47465 & ~n47466 ;
  assign n47468 = n4947 & ~n10958 ;
  assign n47472 = ~n12746 & n12850 ;
  assign n47473 = ~n13053 & n47472 ;
  assign n47469 = n1002 & ~n4307 ;
  assign n47470 = n47469 ^ n6868 ^ 1'b0 ;
  assign n47471 = n3970 & ~n47470 ;
  assign n47474 = n47473 ^ n47471 ^ 1'b0 ;
  assign n47475 = n47474 ^ n3729 ^ 1'b0 ;
  assign n47476 = n20996 | n22806 ;
  assign n47478 = n13309 ^ n4932 ^ 1'b0 ;
  assign n47477 = n21341 ^ n15561 ^ 1'b0 ;
  assign n47479 = n47478 ^ n47477 ^ n36799 ;
  assign n47480 = n8274 | n9481 ;
  assign n47481 = ( n44248 & n45557 ) | ( n44248 & n47480 ) | ( n45557 & n47480 ) ;
  assign n47482 = n20320 & ~n40286 ;
  assign n47483 = ~n25069 & n47482 ;
  assign n47484 = n9580 | n47483 ;
  assign n47485 = ~n19702 & n37174 ;
  assign n47486 = n264 & ~n36401 ;
  assign n47487 = n456 & n40042 ;
  assign n47488 = ~n24191 & n47487 ;
  assign n47489 = ~n47486 & n47488 ;
  assign n47490 = n15752 & ~n41234 ;
  assign n47491 = n31297 ^ n23641 ^ 1'b0 ;
  assign n47492 = n2397 | n47491 ;
  assign n47493 = n20265 & ~n47492 ;
  assign n47494 = n5733 ^ n4332 ^ 1'b0 ;
  assign n47495 = ~n10155 & n47494 ;
  assign n47496 = n29474 ^ n7953 ^ 1'b0 ;
  assign n47497 = ~n34815 & n47496 ;
  assign n47498 = n7177 & n10348 ;
  assign n47499 = n47498 ^ n13208 ^ 1'b0 ;
  assign n47500 = n26284 ^ n12698 ^ 1'b0 ;
  assign n47501 = n12665 & ~n18385 ;
  assign n47502 = n47501 ^ n26563 ^ 1'b0 ;
  assign n47503 = n6037 & ~n41170 ;
  assign n47504 = ( n25862 & ~n28616 ) | ( n25862 & n47503 ) | ( ~n28616 & n47503 ) ;
  assign n47505 = n44266 ^ n12470 ^ 1'b0 ;
  assign n47506 = n46484 & ~n47505 ;
  assign n47507 = n3060 & ~n14541 ;
  assign n47508 = n13992 ^ n12713 ^ 1'b0 ;
  assign n47509 = n27267 & n47508 ;
  assign n47510 = n5025 & n47509 ;
  assign n47511 = ~n4340 & n47510 ;
  assign n47512 = n20379 | n46852 ;
  assign n47513 = n47512 ^ n5813 ^ 1'b0 ;
  assign n47514 = ~n11423 & n20068 ;
  assign n47515 = ~n7620 & n47514 ;
  assign n47516 = n10449 | n28006 ;
  assign n47517 = n9771 | n47516 ;
  assign n47518 = n6898 ^ n934 ^ 1'b0 ;
  assign n47519 = ~n654 & n47518 ;
  assign n47520 = ~n11608 & n47519 ;
  assign n47521 = ~n1055 & n47520 ;
  assign n47522 = n11383 ^ n4054 ^ 1'b0 ;
  assign n47523 = n30341 | n47522 ;
  assign n47524 = n11431 | n47523 ;
  assign n47525 = n47521 & ~n47524 ;
  assign n47526 = n1853 & n37986 ;
  assign n47527 = n26671 | n37784 ;
  assign n47528 = n47527 ^ n45907 ^ n1337 ;
  assign n47529 = n9515 | n9597 ;
  assign n47530 = n673 ^ n575 ^ 1'b0 ;
  assign n47531 = n36706 | n47530 ;
  assign n47532 = ( n3181 & ~n47529 ) | ( n3181 & n47531 ) | ( ~n47529 & n47531 ) ;
  assign n47533 = n21948 ^ n10962 ^ 1'b0 ;
  assign n47534 = n34152 ^ n8330 ^ 1'b0 ;
  assign n47535 = n9511 | n14486 ;
  assign n47536 = n22203 | n47535 ;
  assign n47537 = n46416 ^ n1237 ^ 1'b0 ;
  assign n47538 = n11164 ^ n4808 ^ 1'b0 ;
  assign n47539 = n16313 ^ n9673 ^ 1'b0 ;
  assign n47540 = n47539 ^ n16699 ^ n1229 ;
  assign n47541 = ~n3716 & n17781 ;
  assign n47542 = n2152 & n47541 ;
  assign n47543 = n40560 ^ n27700 ^ 1'b0 ;
  assign n47544 = n10500 ^ n7875 ^ 1'b0 ;
  assign n47545 = ~n11798 & n38637 ;
  assign n47546 = n3891 & n20031 ;
  assign n47547 = n2145 & n45878 ;
  assign n47548 = ~n47546 & n47547 ;
  assign n47549 = n47548 ^ n11813 ^ 1'b0 ;
  assign n47550 = n14349 ^ n1445 ^ 1'b0 ;
  assign n47551 = n8728 ^ n1385 ^ 1'b0 ;
  assign n47552 = n47551 ^ n22242 ^ 1'b0 ;
  assign n47553 = ~n47550 & n47552 ;
  assign n47554 = ~n13526 & n32542 ;
  assign n47555 = ~n4133 & n43676 ;
  assign n47556 = n47555 ^ n3591 ^ n563 ;
  assign n47557 = n47556 ^ n36810 ^ 1'b0 ;
  assign n47558 = n8303 ^ n6613 ^ 1'b0 ;
  assign n47559 = ~n47557 & n47558 ;
  assign n47560 = n47559 ^ n41407 ^ 1'b0 ;
  assign n47561 = n41278 & n47560 ;
  assign n47562 = n9585 ^ n9368 ^ n9163 ;
  assign n47563 = n35743 ^ n2926 ^ 1'b0 ;
  assign n47564 = n47562 & ~n47563 ;
  assign n47567 = n17630 ^ n8148 ^ 1'b0 ;
  assign n47568 = n5454 & ~n47567 ;
  assign n47569 = n47568 ^ n34981 ^ 1'b0 ;
  assign n47565 = n14564 | n35494 ;
  assign n47566 = n10002 & ~n47565 ;
  assign n47570 = n47569 ^ n47566 ^ 1'b0 ;
  assign n47571 = n6514 & ~n31765 ;
  assign n47572 = n3315 | n5178 ;
  assign n47573 = n47572 ^ n29304 ^ 1'b0 ;
  assign n47574 = n9860 & ~n12561 ;
  assign n47575 = ~n47573 & n47574 ;
  assign n47576 = ( n10211 & n39122 ) | ( n10211 & n47575 ) | ( n39122 & n47575 ) ;
  assign n47577 = ( n6285 & ~n9353 ) | ( n6285 & n29854 ) | ( ~n9353 & n29854 ) ;
  assign n47578 = n16846 & n47577 ;
  assign n47579 = n30215 ^ n12790 ^ 1'b0 ;
  assign n47580 = ~n326 & n23708 ;
  assign n47581 = n47580 ^ n33533 ^ 1'b0 ;
  assign n47582 = n47579 & ~n47581 ;
  assign n47583 = ~n6465 & n47582 ;
  assign n47584 = ( n26312 & n38586 ) | ( n26312 & ~n40375 ) | ( n38586 & ~n40375 ) ;
  assign n47585 = n10909 & ~n23572 ;
  assign n47586 = ~n47584 & n47585 ;
  assign n47587 = n47586 ^ n2955 ^ 1'b0 ;
  assign n47588 = ~n35163 & n47587 ;
  assign n47589 = n5689 & n8000 ;
  assign n47590 = n47589 ^ n6164 ^ 1'b0 ;
  assign n47591 = n1338 & n47590 ;
  assign n47592 = n47591 ^ n38391 ^ n18393 ;
  assign n47593 = n36826 ^ n11797 ^ 1'b0 ;
  assign n47594 = n4411 ^ n2677 ^ n1798 ;
  assign n47595 = n47594 ^ n4276 ^ 1'b0 ;
  assign n47596 = n21547 | n47595 ;
  assign n47597 = n47334 & n47596 ;
  assign n47598 = n19231 & ~n34786 ;
  assign n47599 = n47597 & n47598 ;
  assign n47600 = n9192 & ~n18963 ;
  assign n47601 = n17692 & n47600 ;
  assign n47602 = n33916 ^ n30650 ^ 1'b0 ;
  assign n47603 = n38993 ^ n7515 ^ 1'b0 ;
  assign n47604 = n8986 & n20187 ;
  assign n47605 = ~n3558 & n14160 ;
  assign n47606 = n10486 & n47605 ;
  assign n47607 = n5402 & ~n47606 ;
  assign n47608 = ( ~n2164 & n5008 ) | ( ~n2164 & n32454 ) | ( n5008 & n32454 ) ;
  assign n47609 = n16525 ^ n2028 ^ 1'b0 ;
  assign n47610 = ~n20457 & n47609 ;
  assign n47611 = n6656 & n38638 ;
  assign n47612 = n47611 ^ n4971 ^ 1'b0 ;
  assign n47613 = n8478 ^ n2594 ^ 1'b0 ;
  assign n47614 = ~n33727 & n47613 ;
  assign n47615 = n38462 ^ n21101 ^ 1'b0 ;
  assign n47616 = n19164 & ~n47615 ;
  assign n47617 = ~n16328 & n47616 ;
  assign n47618 = ( n325 & n28362 ) | ( n325 & ~n47617 ) | ( n28362 & ~n47617 ) ;
  assign n47619 = n34753 ^ n2326 ^ 1'b0 ;
  assign n47620 = ( n4103 & n27288 ) | ( n4103 & n30271 ) | ( n27288 & n30271 ) ;
  assign n47621 = ~n2397 & n34071 ;
  assign n47622 = n47621 ^ n42061 ^ 1'b0 ;
  assign n47623 = n47622 ^ n560 ^ 1'b0 ;
  assign n47624 = ~n47620 & n47623 ;
  assign n47625 = ( ~n65 & n7108 ) | ( ~n65 & n18712 ) | ( n7108 & n18712 ) ;
  assign n47626 = ~n2070 & n5866 ;
  assign n47627 = ~n5839 & n47626 ;
  assign n47628 = n33016 ^ n32509 ^ 1'b0 ;
  assign n47629 = n3633 | n47628 ;
  assign n47630 = n47629 ^ n43760 ^ n7539 ;
  assign n47631 = n1670 & ~n10189 ;
  assign n47632 = n47631 ^ n39085 ^ 1'b0 ;
  assign n47633 = n1025 & n16788 ;
  assign n47634 = n47633 ^ n29938 ^ 1'b0 ;
  assign n47635 = ~n39708 & n47634 ;
  assign n47637 = n96 & n33204 ;
  assign n47636 = ~n14735 & n37595 ;
  assign n47638 = n47637 ^ n47636 ^ 1'b0 ;
  assign n47639 = ~n47635 & n47638 ;
  assign n47640 = ~n27219 & n32654 ;
  assign n47641 = n17124 & n18371 ;
  assign n47642 = n47641 ^ n18859 ^ 1'b0 ;
  assign n47643 = ~n4924 & n47256 ;
  assign n47644 = n21480 ^ n5821 ^ n4341 ;
  assign n47645 = n28262 & n47644 ;
  assign n47646 = n47645 ^ n4879 ^ 1'b0 ;
  assign n47647 = n10568 ^ n5023 ^ 1'b0 ;
  assign n47648 = n13891 | n46376 ;
  assign n47649 = n34215 ^ n18371 ^ n14746 ;
  assign n47650 = ~n14877 & n17052 ;
  assign n47651 = n47649 & n47650 ;
  assign n47652 = n7191 | n17251 ;
  assign n47653 = n45909 ^ n2277 ^ n2256 ;
  assign n47654 = n29750 ^ n21586 ^ 1'b0 ;
  assign n47655 = n47653 & ~n47654 ;
  assign n47656 = n39336 ^ n8421 ^ 1'b0 ;
  assign n47657 = ~n6709 & n47656 ;
  assign n47660 = n2552 ^ n1745 ^ n1675 ;
  assign n47658 = n45077 ^ n37980 ^ 1'b0 ;
  assign n47659 = n41442 & n47658 ;
  assign n47661 = n47660 ^ n47659 ^ 1'b0 ;
  assign n47662 = n17414 & n24516 ;
  assign n47663 = n12596 ^ n343 ^ 1'b0 ;
  assign n47664 = n47663 ^ n26002 ^ 1'b0 ;
  assign n47665 = n12167 | n21241 ;
  assign n47666 = n47664 & ~n47665 ;
  assign n47667 = n15957 & n47666 ;
  assign n47668 = n16211 & n42786 ;
  assign n47669 = n6479 & n47668 ;
  assign n47670 = n3439 | n10019 ;
  assign n47671 = n26837 & ~n47670 ;
  assign n47672 = n47671 ^ n33216 ^ 1'b0 ;
  assign n47673 = n20393 ^ n4195 ^ 1'b0 ;
  assign n47674 = n39102 & ~n47673 ;
  assign n47675 = n47674 ^ n22173 ^ 1'b0 ;
  assign n47676 = n10059 ^ n8492 ^ 1'b0 ;
  assign n47678 = n19830 ^ n14099 ^ 1'b0 ;
  assign n47677 = n20168 | n33452 ;
  assign n47679 = n47678 ^ n47677 ^ 1'b0 ;
  assign n47680 = n24342 ^ n13179 ^ 1'b0 ;
  assign n47681 = n18129 | n47680 ;
  assign n47682 = n47681 ^ n21952 ^ 1'b0 ;
  assign n47683 = n18933 & n25955 ;
  assign n47684 = n298 & n7061 ;
  assign n47685 = n47684 ^ n2379 ^ 1'b0 ;
  assign n47686 = n23521 ^ n20906 ^ 1'b0 ;
  assign n47687 = n11884 & n14540 ;
  assign n47688 = n47687 ^ n2772 ^ 1'b0 ;
  assign n47689 = ( n9753 & n21919 ) | ( n9753 & n47688 ) | ( n21919 & n47688 ) ;
  assign n47690 = n47689 ^ n1439 ^ 1'b0 ;
  assign n47691 = ~n18704 & n26735 ;
  assign n47692 = n3282 | n7609 ;
  assign n47693 = n28154 | n47692 ;
  assign n47694 = n30154 & n33306 ;
  assign n47695 = n1897 | n47694 ;
  assign n47696 = n47693 | n47695 ;
  assign n47697 = ~n32345 & n37302 ;
  assign n47698 = n47697 ^ n13592 ^ 1'b0 ;
  assign n47699 = ( n5001 & ~n46748 ) | ( n5001 & n47698 ) | ( ~n46748 & n47698 ) ;
  assign n47700 = ~n4032 & n11276 ;
  assign n47701 = ( n7759 & ~n18333 ) | ( n7759 & n47700 ) | ( ~n18333 & n47700 ) ;
  assign n47702 = n27180 ^ n10935 ^ 1'b0 ;
  assign n47703 = n2446 | n47702 ;
  assign n47704 = n13073 & ~n47703 ;
  assign n47705 = n47704 ^ n2420 ^ 1'b0 ;
  assign n47706 = ( n5328 & n27288 ) | ( n5328 & ~n47519 ) | ( n27288 & ~n47519 ) ;
  assign n47707 = n34252 | n47706 ;
  assign n47708 = n36317 ^ n23790 ^ 1'b0 ;
  assign n47709 = n2693 & ~n34955 ;
  assign n47710 = n31918 & n47709 ;
  assign n47711 = n27897 ^ n25428 ^ n3080 ;
  assign n47712 = n8016 & ~n18075 ;
  assign n47713 = n2498 | n4213 ;
  assign n47714 = n47713 ^ n8385 ^ 1'b0 ;
  assign n47715 = n16596 ^ n7342 ^ 1'b0 ;
  assign n47716 = n20268 | n47715 ;
  assign n47717 = n24769 ^ n11008 ^ 1'b0 ;
  assign n47718 = ~n4485 & n7839 ;
  assign n47719 = n47718 ^ n668 ^ 1'b0 ;
  assign n47720 = ~n13452 & n45155 ;
  assign n47721 = n47720 ^ n10675 ^ 1'b0 ;
  assign n47722 = n3674 | n47721 ;
  assign n47723 = n47722 ^ n36844 ^ 1'b0 ;
  assign n47724 = ( ~n1662 & n2567 ) | ( ~n1662 & n47723 ) | ( n2567 & n47723 ) ;
  assign n47725 = ~n3393 & n15359 ;
  assign n47726 = n11946 ^ n3325 ^ 1'b0 ;
  assign n47727 = n10886 | n33647 ;
  assign n47731 = n44625 ^ n4455 ^ 1'b0 ;
  assign n47732 = n33515 | n47731 ;
  assign n47728 = ~n4707 & n29730 ;
  assign n47729 = n12047 & n47728 ;
  assign n47730 = n17477 & ~n47729 ;
  assign n47733 = n47732 ^ n47730 ^ 1'b0 ;
  assign n47734 = n14082 & n42939 ;
  assign n47735 = n47734 ^ n20191 ^ 1'b0 ;
  assign n47736 = n37281 ^ n32707 ^ 1'b0 ;
  assign n47737 = n22593 & n25319 ;
  assign n47738 = n47737 ^ n11664 ^ 1'b0 ;
  assign n47739 = ( n11824 & n12028 ) | ( n11824 & n47738 ) | ( n12028 & n47738 ) ;
  assign n47740 = ~n3827 & n16305 ;
  assign n47741 = n47740 ^ n1360 ^ 1'b0 ;
  assign n47742 = n26130 | n47741 ;
  assign n47743 = n9171 | n14362 ;
  assign n47744 = n19942 & ~n31756 ;
  assign n47745 = n47744 ^ n1306 ^ 1'b0 ;
  assign n47746 = n22596 ^ n18186 ^ 1'b0 ;
  assign n47747 = ~n47228 & n47746 ;
  assign n47748 = ~n4626 & n5576 ;
  assign n47749 = n7691 | n10504 ;
  assign n47750 = n47749 ^ n1109 ^ 1'b0 ;
  assign n47751 = n4448 & n32525 ;
  assign n47752 = n9865 & n47751 ;
  assign n47753 = n10007 ^ n1327 ^ 1'b0 ;
  assign n47754 = n47753 ^ n42301 ^ 1'b0 ;
  assign n47755 = n9892 | n31139 ;
  assign n47756 = n38104 & ~n47755 ;
  assign n47757 = n24864 ^ n22633 ^ n11276 ;
  assign n47758 = n6274 & ~n16902 ;
  assign n47759 = ~n42663 & n47758 ;
  assign n47760 = n12403 | n29030 ;
  assign n47761 = n1644 | n47760 ;
  assign n47762 = ~n9867 & n47761 ;
  assign n47763 = n5385 & n47762 ;
  assign n47764 = n47575 ^ n42155 ^ 1'b0 ;
  assign n47765 = n1312 | n18900 ;
  assign n47766 = n2367 ^ n1688 ^ 1'b0 ;
  assign n47767 = n2894 & ~n47766 ;
  assign n47768 = ~n495 & n24331 ;
  assign n47769 = n47768 ^ n16623 ^ 1'b0 ;
  assign n47770 = n43479 ^ n32157 ^ 1'b0 ;
  assign n47771 = n471 & ~n7606 ;
  assign n47772 = ~n3926 & n47771 ;
  assign n47773 = n5789 & n47772 ;
  assign n47774 = n9923 ^ n8350 ^ 1'b0 ;
  assign n47775 = ~n47773 & n47774 ;
  assign n47776 = ~n11717 & n47775 ;
  assign n47777 = n1000 & n12835 ;
  assign n47778 = n30551 ^ n27171 ^ 1'b0 ;
  assign n47779 = n22207 & ~n47778 ;
  assign n47780 = n11049 & n19515 ;
  assign n47781 = n34712 & n47780 ;
  assign n47782 = n35892 & ~n37342 ;
  assign n47783 = ~n28460 & n44909 ;
  assign n47784 = ~n649 & n47783 ;
  assign n47785 = n17309 ^ n4366 ^ 1'b0 ;
  assign n47786 = n22218 & ~n47785 ;
  assign n47787 = n34987 & n47786 ;
  assign n47788 = ~n7082 & n47787 ;
  assign n47789 = n20667 & ~n31408 ;
  assign n47790 = n47789 ^ n8920 ^ 1'b0 ;
  assign n47791 = n20032 | n47790 ;
  assign n47792 = n11816 ^ n4650 ^ 1'b0 ;
  assign n47793 = ~n3118 & n47792 ;
  assign n47797 = n19821 ^ n12055 ^ n1546 ;
  assign n47795 = n15388 ^ n849 ^ 1'b0 ;
  assign n47796 = n21083 | n47795 ;
  assign n47794 = n12086 ^ n4677 ^ 1'b0 ;
  assign n47798 = n47797 ^ n47796 ^ n47794 ;
  assign n47799 = n47798 ^ n14787 ^ 1'b0 ;
  assign n47800 = n47793 & ~n47799 ;
  assign n47801 = n17559 ^ n592 ^ 1'b0 ;
  assign n47802 = n32158 ^ n21217 ^ 1'b0 ;
  assign n47803 = n31015 & n47802 ;
  assign n47804 = n15826 ^ n5717 ^ 1'b0 ;
  assign n47805 = n5221 & ~n47804 ;
  assign n47806 = ~n32594 & n47805 ;
  assign n47807 = ( n4546 & n8949 ) | ( n4546 & n47806 ) | ( n8949 & n47806 ) ;
  assign n47808 = n47807 ^ n14200 ^ n3166 ;
  assign n47809 = n3504 | n6447 ;
  assign n47810 = n606 & ~n47809 ;
  assign n47811 = n15795 ^ n4297 ^ 1'b0 ;
  assign n47812 = n43557 & n47811 ;
  assign n47813 = n34986 & n47812 ;
  assign n47814 = ~n9183 & n47813 ;
  assign n47815 = n11221 ^ n3944 ^ 1'b0 ;
  assign n47816 = n15413 & n47815 ;
  assign n47817 = n40336 ^ n18108 ^ 1'b0 ;
  assign n47819 = n4545 | n33492 ;
  assign n47818 = n22489 & ~n26723 ;
  assign n47820 = n47819 ^ n47818 ^ 1'b0 ;
  assign n47821 = n19984 & ~n43728 ;
  assign n47822 = ~n47820 & n47821 ;
  assign n47824 = n12990 | n20812 ;
  assign n47823 = ~n6601 & n29310 ;
  assign n47825 = n47824 ^ n47823 ^ 1'b0 ;
  assign n47826 = n47825 ^ n9488 ^ 1'b0 ;
  assign n47827 = ( n41325 & ~n45969 ) | ( n41325 & n47826 ) | ( ~n45969 & n47826 ) ;
  assign n47828 = ~x5 & n29070 ;
  assign n47829 = n47828 ^ n8881 ^ 1'b0 ;
  assign n47830 = n11908 & ~n20457 ;
  assign n47831 = n24726 ^ n9523 ^ 1'b0 ;
  assign n47832 = n27336 & ~n47831 ;
  assign n47833 = n12829 | n47832 ;
  assign n47834 = ~n30397 & n31005 ;
  assign n47835 = n8811 ^ n519 ^ 1'b0 ;
  assign n47836 = ~n11543 & n47835 ;
  assign n47837 = n47836 ^ n25553 ^ 1'b0 ;
  assign n47838 = n18615 ^ n16978 ^ n16047 ;
  assign n47839 = n2038 ^ n615 ^ 1'b0 ;
  assign n47840 = ( ~n8150 & n42545 ) | ( ~n8150 & n47839 ) | ( n42545 & n47839 ) ;
  assign n47841 = n11852 ^ n1999 ^ n1419 ;
  assign n47842 = n27303 | n47841 ;
  assign n47843 = ~n27331 & n33215 ;
  assign n47844 = n1930 & ~n18958 ;
  assign n47845 = n9966 & n31793 ;
  assign n47846 = n10897 & ~n29020 ;
  assign n47847 = n10797 & n47846 ;
  assign n47848 = ~n2820 & n4019 ;
  assign n47849 = n4597 & n28171 ;
  assign n47850 = n47849 ^ n33249 ^ n24927 ;
  assign n47851 = n209 | n4916 ;
  assign n47852 = n1484 & n6174 ;
  assign n47853 = ( n14571 & ~n47851 ) | ( n14571 & n47852 ) | ( ~n47851 & n47852 ) ;
  assign n47854 = n2771 | n46351 ;
  assign n47855 = n2175 | n43381 ;
  assign n47856 = n3060 | n47855 ;
  assign n47857 = n31857 & n38598 ;
  assign n47858 = n47857 ^ n38828 ^ 1'b0 ;
  assign n47859 = n14569 & n41848 ;
  assign n47860 = ~n12251 & n28798 ;
  assign n47861 = n47859 & n47860 ;
  assign n47862 = ~n26796 & n47861 ;
  assign n47863 = ~n8940 & n11111 ;
  assign n47864 = n38297 & ~n41450 ;
  assign n47865 = n9848 & n47864 ;
  assign n47866 = ~n29107 & n47646 ;
  assign n47867 = n31272 ^ n3891 ^ 1'b0 ;
  assign n47868 = n12950 & n47867 ;
  assign n47869 = n571 & n9267 ;
  assign n47870 = n47869 ^ n11160 ^ 1'b0 ;
  assign n47874 = n1507 & n3258 ;
  assign n47871 = n20499 & n35704 ;
  assign n47872 = n47871 ^ n13053 ^ 1'b0 ;
  assign n47873 = n11504 | n47872 ;
  assign n47875 = n47874 ^ n47873 ^ 1'b0 ;
  assign n47876 = n19085 & n30723 ;
  assign n47877 = n2317 & n7782 ;
  assign n47878 = n7167 | n47877 ;
  assign n47879 = n3429 & ~n31424 ;
  assign n47880 = n47878 & n47879 ;
  assign n47881 = n8396 & n26744 ;
  assign n47882 = ~n30003 & n47881 ;
  assign n47883 = n47882 ^ n2890 ^ 1'b0 ;
  assign n47884 = n47880 & ~n47883 ;
  assign n47885 = n4775 ^ n3685 ^ 1'b0 ;
  assign n47886 = n8650 & ~n47885 ;
  assign n47887 = n10119 & n43274 ;
  assign n47888 = n22776 ^ n9808 ^ 1'b0 ;
  assign n47889 = ~n18888 & n47888 ;
  assign n47890 = ~n24875 & n47889 ;
  assign n47891 = n29921 ^ n11276 ^ 1'b0 ;
  assign n47892 = n47890 | n47891 ;
  assign n47893 = n8670 & ~n27092 ;
  assign n47894 = n47893 ^ n16725 ^ 1'b0 ;
  assign n47895 = n30521 | n41245 ;
  assign n47896 = ~n10894 & n33608 ;
  assign n47897 = n42072 ^ n13988 ^ 1'b0 ;
  assign n47898 = n16179 & ~n16743 ;
  assign n47899 = n47897 & n47898 ;
  assign n47900 = n27874 & ~n47899 ;
  assign n47901 = n4429 & n47900 ;
  assign n47902 = n22204 & ~n47901 ;
  assign n47903 = n47902 ^ n23253 ^ 1'b0 ;
  assign n47904 = n10797 & n14727 ;
  assign n47905 = n17210 & ~n27804 ;
  assign n47906 = ~n16555 & n23264 ;
  assign n47907 = n41682 & n47906 ;
  assign n47908 = n42468 ^ n23833 ^ n1697 ;
  assign n47909 = n8487 ^ n3800 ^ n2399 ;
  assign n47910 = n47874 & ~n47909 ;
  assign n47911 = n39759 ^ n9356 ^ 1'b0 ;
  assign n47912 = n9843 ^ n2309 ^ 1'b0 ;
  assign n47913 = n47912 ^ n35912 ^ n23865 ;
  assign n47914 = ~n4113 & n28631 ;
  assign n47915 = ~n42917 & n47914 ;
  assign n47916 = n47915 ^ n1623 ^ 1'b0 ;
  assign n47917 = n11116 & ~n32539 ;
  assign n47919 = n4329 & ~n12179 ;
  assign n47918 = n5285 | n23945 ;
  assign n47920 = n47919 ^ n47918 ^ 1'b0 ;
  assign n47921 = n47920 ^ n37793 ^ n7623 ;
  assign n47922 = n38746 ^ n5002 ^ 1'b0 ;
  assign n47923 = n36193 ^ n19200 ^ 1'b0 ;
  assign n47924 = n25214 & ~n47923 ;
  assign n47925 = n47924 ^ n26112 ^ 1'b0 ;
  assign n47926 = n26770 ^ n14940 ^ 1'b0 ;
  assign n47927 = n2980 | n47926 ;
  assign n47928 = n1466 & ~n28372 ;
  assign n47929 = ~n225 & n20021 ;
  assign n47930 = n19825 & n47929 ;
  assign n47931 = n47930 ^ n9495 ^ 1'b0 ;
  assign n47932 = ~n47928 & n47931 ;
  assign n47933 = n38385 ^ n16018 ^ 1'b0 ;
  assign n47934 = n2789 | n4305 ;
  assign n47935 = ~n14400 & n17399 ;
  assign n47936 = n16888 & n47935 ;
  assign n47937 = n47936 ^ n3108 ^ 1'b0 ;
  assign n47938 = n28354 ^ n23449 ^ n22235 ;
  assign n47939 = n47938 ^ n21958 ^ 1'b0 ;
  assign n47940 = n16059 & ~n21509 ;
  assign n47941 = n47940 ^ n31511 ^ 1'b0 ;
  assign n47942 = n27132 & n47941 ;
  assign n47943 = n17424 | n30534 ;
  assign n47944 = n35182 ^ n19995 ^ n1545 ;
  assign n47945 = n45777 & n47944 ;
  assign n47946 = n47945 ^ n32133 ^ 1'b0 ;
  assign n47948 = n20457 ^ n7389 ^ 1'b0 ;
  assign n47947 = ~n12494 & n13690 ;
  assign n47949 = n47948 ^ n47947 ^ 1'b0 ;
  assign n47950 = n5946 | n11546 ;
  assign n47951 = n3423 & ~n12204 ;
  assign n47952 = ~n2745 & n44172 ;
  assign n47953 = ~n21100 & n25777 ;
  assign n47954 = n17578 | n18568 ;
  assign n47955 = ~n34712 & n47954 ;
  assign n47956 = n47955 ^ n34072 ^ 1'b0 ;
  assign n47957 = n4947 & ~n18936 ;
  assign n47958 = n21490 ^ n16367 ^ 1'b0 ;
  assign n47959 = n16350 | n47958 ;
  assign n47960 = n22646 ^ n13311 ^ 1'b0 ;
  assign n47961 = n18565 & ~n47960 ;
  assign n47962 = n13505 & ~n14177 ;
  assign n47963 = n47962 ^ n11703 ^ 1'b0 ;
  assign n47964 = n36176 ^ n1075 ^ 1'b0 ;
  assign n47965 = ( n2382 & ~n45930 ) | ( n2382 & n47964 ) | ( ~n45930 & n47964 ) ;
  assign n47966 = n47830 ^ n20520 ^ 1'b0 ;
  assign n47967 = n14085 | n47966 ;
  assign n47968 = n619 & ~n24983 ;
  assign n47969 = n27585 ^ n4356 ^ 1'b0 ;
  assign n47970 = n13314 & n47969 ;
  assign n47971 = ~n14175 & n47970 ;
  assign n47972 = n31832 ^ n19400 ^ 1'b0 ;
  assign n47973 = n47971 & ~n47972 ;
  assign n47980 = n11159 ^ n6972 ^ n510 ;
  assign n47974 = ~n1441 & n7308 ;
  assign n47975 = n47974 ^ n5235 ^ 1'b0 ;
  assign n47976 = ~n9725 & n47975 ;
  assign n47977 = n821 & n47976 ;
  assign n47978 = n47977 ^ n1747 ^ 1'b0 ;
  assign n47979 = n47978 ^ n4497 ^ 1'b0 ;
  assign n47981 = n47980 ^ n47979 ^ n1069 ;
  assign n47982 = n7442 & ~n32418 ;
  assign n47983 = n47982 ^ n47477 ^ 1'b0 ;
  assign n47984 = ~n21170 & n47983 ;
  assign n47985 = ~n5264 & n11770 ;
  assign n47986 = n47985 ^ n27247 ^ 1'b0 ;
  assign n47987 = n47678 & ~n47986 ;
  assign n47988 = n35071 | n47987 ;
  assign n47989 = n23927 | n47988 ;
  assign n47990 = n1165 & ~n19747 ;
  assign n47991 = n296 & n47990 ;
  assign n47992 = n47991 ^ n22983 ^ 1'b0 ;
  assign n47993 = n14994 & ~n47992 ;
  assign n47994 = n6622 & ~n23520 ;
  assign n47995 = ~n24483 & n40578 ;
  assign n47996 = n845 & n11180 ;
  assign n47997 = n47996 ^ n8505 ^ 1'b0 ;
  assign n47998 = n41382 ^ n32816 ^ 1'b0 ;
  assign n47999 = n47998 ^ n15117 ^ 1'b0 ;
  assign n48000 = n38097 & ~n47999 ;
  assign n48001 = ~n11167 & n29493 ;
  assign n48002 = n12171 | n33203 ;
  assign n48003 = n48002 ^ n21245 ^ 1'b0 ;
  assign n48004 = ( n28342 & n41202 ) | ( n28342 & ~n48003 ) | ( n41202 & ~n48003 ) ;
  assign n48005 = n29286 ^ n12600 ^ 1'b0 ;
  assign n48006 = n4041 & ~n31758 ;
  assign n48007 = n25703 ^ n23518 ^ 1'b0 ;
  assign n48008 = ~n48006 & n48007 ;
  assign n48009 = n29279 ^ n860 ^ 1'b0 ;
  assign n48010 = n25546 & n48009 ;
  assign n48011 = n48010 ^ n33387 ^ 1'b0 ;
  assign n48012 = n24687 & ~n40304 ;
  assign n48013 = n48012 ^ n3930 ^ 1'b0 ;
  assign n48014 = n13863 & ~n48013 ;
  assign n48015 = n8405 & n48014 ;
  assign n48017 = ~n780 & n37991 ;
  assign n48016 = ~n4881 & n25370 ;
  assign n48018 = n48017 ^ n48016 ^ 1'b0 ;
  assign n48019 = n47335 & n48018 ;
  assign n48020 = ~n12817 & n48019 ;
  assign n48021 = n20472 & n37169 ;
  assign n48022 = ( n30044 & ~n45188 ) | ( n30044 & n48021 ) | ( ~n45188 & n48021 ) ;
  assign n48023 = ~n4903 & n14775 ;
  assign n48024 = n588 & n48023 ;
  assign n48025 = n30302 & n48024 ;
  assign n48026 = ~n291 & n954 ;
  assign n48027 = ~n12606 & n48026 ;
  assign n48028 = ~n3031 & n28389 ;
  assign n48029 = n48027 & n48028 ;
  assign n48030 = n468 | n48029 ;
  assign n48031 = n48030 ^ n31287 ^ 1'b0 ;
  assign n48032 = n14890 ^ n3951 ^ 1'b0 ;
  assign n48033 = n28280 & n48032 ;
  assign n48034 = ~n14439 & n33077 ;
  assign n48035 = ~n22893 & n46933 ;
  assign n48036 = ~n48034 & n48035 ;
  assign n48037 = n9288 & ~n11400 ;
  assign n48038 = n48037 ^ n6099 ^ 1'b0 ;
  assign n48039 = n10647 & n48038 ;
  assign n48040 = ( n28375 & ~n42156 ) | ( n28375 & n43292 ) | ( ~n42156 & n43292 ) ;
  assign n48045 = n1915 & n4146 ;
  assign n48043 = n21812 | n44365 ;
  assign n48044 = n48043 ^ n46392 ^ 1'b0 ;
  assign n48046 = n48045 ^ n48044 ^ 1'b0 ;
  assign n48041 = ~n14200 & n42711 ;
  assign n48042 = n48041 ^ n41855 ^ 1'b0 ;
  assign n48047 = n48046 ^ n48042 ^ 1'b0 ;
  assign n48048 = n9857 ^ n2772 ^ 1'b0 ;
  assign n48049 = ~n39948 & n48048 ;
  assign n48051 = n27728 ^ n9489 ^ 1'b0 ;
  assign n48050 = ~n35086 & n36983 ;
  assign n48052 = n48051 ^ n48050 ^ 1'b0 ;
  assign n48053 = n7492 & n33705 ;
  assign n48054 = n48053 ^ n28 ^ 1'b0 ;
  assign n48055 = ( n2735 & ~n42643 ) | ( n2735 & n45889 ) | ( ~n42643 & n45889 ) ;
  assign n48056 = ~n9463 & n12665 ;
  assign n48057 = n535 & n15159 ;
  assign n48058 = ( n5712 & n31517 ) | ( n5712 & ~n40936 ) | ( n31517 & ~n40936 ) ;
  assign n48059 = n48058 ^ n33060 ^ 1'b0 ;
  assign n48060 = n14887 & ~n48059 ;
  assign n48061 = n5030 | n20902 ;
  assign n48062 = n10144 & n41910 ;
  assign n48063 = ~n9055 & n11005 ;
  assign n48064 = n48063 ^ n1217 ^ 1'b0 ;
  assign n48065 = n7209 & ~n48064 ;
  assign n48066 = n18760 & n21344 ;
  assign n48067 = n39663 & n48066 ;
  assign n48068 = n40312 ^ n15705 ^ 1'b0 ;
  assign n48069 = n48067 | n48068 ;
  assign n48070 = n1382 & n19770 ;
  assign n48071 = ( ~n2076 & n10753 ) | ( ~n2076 & n30651 ) | ( n10753 & n30651 ) ;
  assign n48072 = n48071 ^ n14007 ^ 1'b0 ;
  assign n48073 = n439 & n48072 ;
  assign n48074 = ~n25277 & n39479 ;
  assign n48075 = n48074 ^ n10628 ^ 1'b0 ;
  assign n48076 = ~n27857 & n48075 ;
  assign n48077 = ~n26798 & n48076 ;
  assign n48078 = n4074 ^ n2031 ^ 1'b0 ;
  assign n48079 = n905 & ~n45363 ;
  assign n48080 = n48079 ^ n19698 ^ 1'b0 ;
  assign n48081 = n38190 ^ n33113 ^ 1'b0 ;
  assign n48082 = n48081 ^ n14208 ^ n8685 ;
  assign n48083 = n8980 | n29726 ;
  assign n48084 = n8980 & ~n48083 ;
  assign n48085 = x5 & n44145 ;
  assign n48086 = n15475 & ~n48085 ;
  assign n48087 = n48085 & n48086 ;
  assign n48088 = n5270 & ~n48087 ;
  assign n48089 = n4729 & ~n20895 ;
  assign n48090 = n20895 & n48089 ;
  assign n48091 = n1050 | n10428 ;
  assign n48092 = n10428 & ~n48091 ;
  assign n48093 = n11827 & ~n48092 ;
  assign n48094 = n1092 & n3080 ;
  assign n48095 = ~n1092 & n48094 ;
  assign n48096 = n48093 & ~n48095 ;
  assign n48097 = ~n48093 & n48096 ;
  assign n48098 = n48097 ^ n21366 ^ 1'b0 ;
  assign n48099 = n1159 | n48098 ;
  assign n48100 = n48090 & ~n48099 ;
  assign n48101 = n48088 & n48100 ;
  assign n48102 = n48084 & n48101 ;
  assign n48103 = n39200 ^ n7771 ^ 1'b0 ;
  assign n48104 = n22239 & ~n36529 ;
  assign n48105 = n48104 ^ n8664 ^ 1'b0 ;
  assign n48106 = ( n948 & n19489 ) | ( n948 & n42804 ) | ( n19489 & n42804 ) ;
  assign n48107 = ~n362 & n36590 ;
  assign n48108 = n5685 ^ n3270 ^ 1'b0 ;
  assign n48109 = n48107 & n48108 ;
  assign n48110 = n48109 ^ n4493 ^ 1'b0 ;
  assign n48111 = n9751 & ~n11824 ;
  assign n48112 = n19918 ^ n2791 ^ 1'b0 ;
  assign n48113 = ~n17578 & n48112 ;
  assign n48114 = n48113 ^ n5377 ^ 1'b0 ;
  assign n48115 = n21967 | n48114 ;
  assign n48116 = n13808 ^ n8801 ^ n3262 ;
  assign n48117 = n10979 | n48116 ;
  assign n48119 = n5555 | n23633 ;
  assign n48120 = n48119 ^ n505 ^ 1'b0 ;
  assign n48118 = n5364 | n46580 ;
  assign n48121 = n48120 ^ n48118 ^ 1'b0 ;
  assign n48122 = n5432 & ~n15166 ;
  assign n48123 = n30993 ^ n22034 ^ n15224 ;
  assign n48124 = n4056 | n48123 ;
  assign n48126 = n29653 ^ n5906 ^ 1'b0 ;
  assign n48125 = n33538 | n47179 ;
  assign n48127 = n48126 ^ n48125 ^ 1'b0 ;
  assign n48128 = n22276 ^ n21488 ^ n19228 ;
  assign n48129 = n19 & ~n24496 ;
  assign n48130 = n47018 & n48129 ;
  assign n48131 = n15514 | n48130 ;
  assign n48132 = n535 & ~n3325 ;
  assign n48133 = ~n30650 & n48132 ;
  assign n48134 = n7285 | n22046 ;
  assign n48135 = n48134 ^ n18425 ^ n1223 ;
  assign n48137 = n3112 & n9602 ;
  assign n48136 = ~n8979 & n16282 ;
  assign n48138 = n48137 ^ n48136 ^ 1'b0 ;
  assign n48139 = n48138 ^ n13389 ^ 1'b0 ;
  assign n48140 = n37148 & n48139 ;
  assign n48141 = n11035 | n48140 ;
  assign n48142 = n48135 | n48141 ;
  assign n48143 = n12104 & n19824 ;
  assign n48144 = ~n4651 & n48143 ;
  assign n48145 = n48144 ^ n44980 ^ n18066 ;
  assign n48146 = n16756 ^ n7990 ^ 1'b0 ;
  assign n48147 = n33214 | n48146 ;
  assign n48148 = n2637 ^ n316 ^ 1'b0 ;
  assign n48149 = ~n3833 & n12219 ;
  assign n48150 = ~n48148 & n48149 ;
  assign n48151 = n48150 ^ n41500 ^ 1'b0 ;
  assign n48152 = n21081 & ~n48151 ;
  assign n48155 = n9662 & n21074 ;
  assign n48156 = n5503 & n48155 ;
  assign n48153 = ~n667 & n19548 ;
  assign n48154 = n18049 & n48153 ;
  assign n48157 = n48156 ^ n48154 ^ 1'b0 ;
  assign n48158 = n38190 ^ n15193 ^ 1'b0 ;
  assign n48159 = n10225 & ~n39862 ;
  assign n48160 = ~n33667 & n48159 ;
  assign n48161 = ~n9418 & n10005 ;
  assign n48162 = n34215 & n48161 ;
  assign n48163 = n36046 & n39968 ;
  assign n48164 = ~n14793 & n42155 ;
  assign n48165 = ~n38861 & n48164 ;
  assign n48166 = n8388 & n48165 ;
  assign n48167 = n34463 ^ n30593 ^ 1'b0 ;
  assign n48168 = n39503 & n48167 ;
  assign n48169 = n48168 ^ n42234 ^ 1'b0 ;
  assign n48170 = n44603 ^ n4662 ^ 1'b0 ;
  assign n48171 = n16435 ^ n1426 ^ 1'b0 ;
  assign n48172 = n46618 & n48171 ;
  assign n48173 = n48172 ^ n40259 ^ n12862 ;
  assign n48174 = n25966 ^ n18562 ^ 1'b0 ;
  assign n48175 = n18215 | n19984 ;
  assign n48176 = n1454 | n5916 ;
  assign n48177 = n31771 | n38006 ;
  assign n48178 = n21217 | n38327 ;
  assign n48179 = ~n6416 & n39154 ;
  assign n48180 = n2049 | n30441 ;
  assign n48181 = n3056 & ~n48180 ;
  assign n48182 = n32925 ^ n19202 ^ 1'b0 ;
  assign n48183 = n19619 ^ n11458 ^ 1'b0 ;
  assign n48184 = n22228 ^ n18200 ^ 1'b0 ;
  assign n48185 = n18122 | n48184 ;
  assign n48186 = ~n17573 & n31007 ;
  assign n48187 = n48186 ^ n16172 ^ 1'b0 ;
  assign n48188 = n682 & n29326 ;
  assign n48189 = n26302 | n48188 ;
  assign n48190 = n48187 | n48189 ;
  assign n48191 = ( n2616 & n8901 ) | ( n2616 & n15315 ) | ( n8901 & n15315 ) ;
  assign n48192 = n29530 & n35467 ;
  assign n48193 = ~n8144 & n17326 ;
  assign n48194 = n48193 ^ n12579 ^ 1'b0 ;
  assign n48195 = n44415 & n48194 ;
  assign n48196 = ~n21021 & n32397 ;
  assign n48197 = ~n2971 & n35818 ;
  assign n48198 = n48197 ^ n44094 ^ 1'b0 ;
  assign n48199 = ~n20544 & n48198 ;
  assign n48200 = n47343 ^ n37213 ^ 1'b0 ;
  assign n48201 = ~n7836 & n48200 ;
  assign n48202 = n48201 ^ n19680 ^ 1'b0 ;
  assign n48203 = n16144 | n20755 ;
  assign n48204 = n7627 ^ n3858 ^ n1327 ;
  assign n48205 = n20067 | n48204 ;
  assign n48206 = n48205 ^ n27534 ^ 1'b0 ;
  assign n48207 = ~n48203 & n48206 ;
  assign n48208 = ~n23869 & n27395 ;
  assign n48209 = ~n35387 & n43291 ;
  assign n48210 = n14829 & n35339 ;
  assign n48211 = n16040 & n40803 ;
  assign n48212 = ~n3363 & n48211 ;
  assign n48213 = n83 | n43779 ;
  assign n48214 = n48213 ^ n21660 ^ 1'b0 ;
  assign n48215 = n22128 | n40264 ;
  assign n48216 = n8665 ^ n929 ^ 1'b0 ;
  assign n48217 = n2397 | n48216 ;
  assign n48218 = n44355 | n48217 ;
  assign n48219 = n48218 ^ n5082 ^ 1'b0 ;
  assign n48220 = n21735 & n48219 ;
  assign n48221 = ~n7130 & n48220 ;
  assign n48222 = n508 | n10298 ;
  assign n48223 = ~n29865 & n32104 ;
  assign n48224 = n12324 & ~n48223 ;
  assign n48225 = ~n48222 & n48224 ;
  assign n48228 = n5008 | n26525 ;
  assign n48229 = n5008 & ~n48228 ;
  assign n48226 = n17013 | n45569 ;
  assign n48227 = n48226 ^ n12979 ^ 1'b0 ;
  assign n48230 = n48229 ^ n48227 ^ n39637 ;
  assign n48231 = n37523 ^ n11374 ^ 1'b0 ;
  assign n48232 = n6802 & ~n43015 ;
  assign n48233 = n40138 ^ n2845 ^ 1'b0 ;
  assign n48234 = ( n2876 & n25977 ) | ( n2876 & n48233 ) | ( n25977 & n48233 ) ;
  assign n48235 = n44807 ^ n5911 ^ 1'b0 ;
  assign n48236 = n48234 & n48235 ;
  assign n48237 = n48236 ^ n12343 ^ n7140 ;
  assign n48238 = n47080 ^ n37729 ^ n16934 ;
  assign n48240 = ~n11752 & n40702 ;
  assign n48241 = n48240 ^ n870 ^ 1'b0 ;
  assign n48239 = n4267 | n39037 ;
  assign n48242 = n48241 ^ n48239 ^ 1'b0 ;
  assign n48243 = n48242 ^ n4891 ^ 1'b0 ;
  assign n48244 = ~n9823 & n16119 ;
  assign n48245 = n35382 ^ n24346 ^ 1'b0 ;
  assign n48246 = ~n5660 & n48245 ;
  assign n48247 = n29961 & n48246 ;
  assign n48248 = n11887 | n28482 ;
  assign n48249 = n8559 & ~n11829 ;
  assign n48250 = ( ~n7659 & n18908 ) | ( ~n7659 & n48249 ) | ( n18908 & n48249 ) ;
  assign n48251 = ( ~n8217 & n45458 ) | ( ~n8217 & n48250 ) | ( n45458 & n48250 ) ;
  assign n48252 = n8468 & ~n26453 ;
  assign n48253 = ~n19428 & n48252 ;
  assign n48254 = n4732 ^ n2426 ^ 1'b0 ;
  assign n48255 = n2326 | n31579 ;
  assign n48256 = n48254 & ~n48255 ;
  assign n48257 = n18041 ^ n10711 ^ 1'b0 ;
  assign n48258 = ~n28263 & n48257 ;
  assign n48259 = n48258 ^ n42795 ^ n17855 ;
  assign n48260 = ~n5452 & n48259 ;
  assign n48261 = n45308 ^ n21 ^ 1'b0 ;
  assign n48262 = n34890 ^ n7864 ^ 1'b0 ;
  assign n48263 = n17189 | n48262 ;
  assign n48264 = n7736 ^ n7497 ^ 1'b0 ;
  assign n48265 = n10055 | n48264 ;
  assign n48266 = ( n13 & ~n3315 ) | ( n13 & n48265 ) | ( ~n3315 & n48265 ) ;
  assign n48267 = n1376 & ~n7730 ;
  assign n48268 = n1663 & ~n3382 ;
  assign n48269 = n48268 ^ n16651 ^ n14329 ;
  assign n48270 = n36762 ^ n3724 ^ 1'b0 ;
  assign n48271 = ~n8785 & n48270 ;
  assign n48272 = n43603 ^ n9854 ^ 1'b0 ;
  assign n48273 = n26130 & n26729 ;
  assign n48274 = ~n39146 & n48273 ;
  assign n48275 = n466 & n14109 ;
  assign n48276 = n48275 ^ n20467 ^ 1'b0 ;
  assign n48277 = n10845 | n11605 ;
  assign n48278 = n48277 ^ n3730 ^ 1'b0 ;
  assign n48279 = n17339 & n48278 ;
  assign n48280 = n48279 ^ n34098 ^ 1'b0 ;
  assign n48281 = n48280 ^ n1763 ^ 1'b0 ;
  assign n48282 = n7734 | n48281 ;
  assign n48283 = ~n3139 & n6908 ;
  assign n48284 = n18395 & ~n32042 ;
  assign n48285 = ~n1083 & n9594 ;
  assign n48286 = n48285 ^ n10780 ^ 1'b0 ;
  assign n48287 = n48286 ^ n2478 ^ 1'b0 ;
  assign n48288 = n681 | n48287 ;
  assign n48289 = n48288 ^ n23544 ^ 1'b0 ;
  assign n48290 = n28955 & n42975 ;
  assign n48291 = n8497 & ~n14728 ;
  assign n48292 = n48291 ^ n24096 ^ 1'b0 ;
  assign n48293 = n6760 | n31322 ;
  assign n48294 = n48293 ^ n26057 ^ 1'b0 ;
  assign n48295 = n7185 & n14474 ;
  assign n48296 = ~n54 & n48295 ;
  assign n48297 = n34383 | n48296 ;
  assign n48298 = n13956 ^ n8331 ^ 1'b0 ;
  assign n48299 = n38566 ^ n23085 ^ 1'b0 ;
  assign n48300 = n42388 ^ n475 ^ 1'b0 ;
  assign n48301 = n1254 & ~n48300 ;
  assign n48302 = ~n32269 & n48301 ;
  assign n48303 = ~n29756 & n48302 ;
  assign n48304 = n16849 & ~n36958 ;
  assign n48305 = n48304 ^ n753 ^ 1'b0 ;
  assign n48306 = n15275 | n20904 ;
  assign n48307 = n13806 | n25565 ;
  assign n48308 = n10942 & ~n48307 ;
  assign n48309 = n47228 ^ n2838 ^ 1'b0 ;
  assign n48310 = ( n1618 & n26370 ) | ( n1618 & ~n48309 ) | ( n26370 & ~n48309 ) ;
  assign n48311 = n7973 & n48310 ;
  assign n48312 = n478 & ~n10858 ;
  assign n48313 = n29826 & ~n48312 ;
  assign n48314 = ~n927 & n31241 ;
  assign n48315 = ~n12158 & n13663 ;
  assign n48316 = n44312 ^ n6179 ^ 1'b0 ;
  assign n48317 = n48315 & n48316 ;
  assign n48319 = n12516 & n32928 ;
  assign n48320 = n48319 ^ n12679 ^ 1'b0 ;
  assign n48321 = n2377 | n48320 ;
  assign n48322 = n48321 ^ n28714 ^ 1'b0 ;
  assign n48318 = n1688 | n8891 ;
  assign n48323 = n48322 ^ n48318 ^ 1'b0 ;
  assign n48324 = n104 & ~n23720 ;
  assign n48325 = n3933 & n20308 ;
  assign n48326 = ~n48324 & n48325 ;
  assign n48327 = n8105 ^ n4250 ^ 1'b0 ;
  assign n48328 = ~n19854 & n30231 ;
  assign n48329 = n26789 ^ n6203 ^ 1'b0 ;
  assign n48330 = n3315 | n48329 ;
  assign n48332 = ( ~n15760 & n18900 ) | ( ~n15760 & n22740 ) | ( n18900 & n22740 ) ;
  assign n48331 = n664 | n4975 ;
  assign n48333 = n48332 ^ n48331 ^ 1'b0 ;
  assign n48334 = n35931 & n39067 ;
  assign n48335 = n942 & ~n8942 ;
  assign n48336 = n48335 ^ n15262 ^ 1'b0 ;
  assign n48337 = n1938 & n48336 ;
  assign n48338 = ~n667 & n21651 ;
  assign n48339 = n48338 ^ n38855 ^ n9889 ;
  assign n48340 = ~n23043 & n48339 ;
  assign n48341 = n47581 ^ n6857 ^ 1'b0 ;
  assign n48342 = n249 ^ n182 ^ 1'b0 ;
  assign n48343 = n27145 | n36524 ;
  assign n48344 = ( ~n493 & n16170 ) | ( ~n493 & n47140 ) | ( n16170 & n47140 ) ;
  assign n48345 = n48344 ^ n20419 ^ 1'b0 ;
  assign n48346 = n32771 & ~n48345 ;
  assign n48347 = ~n18817 & n48346 ;
  assign n48348 = n2817 & n15289 ;
  assign n48349 = n48348 ^ n2747 ^ 1'b0 ;
  assign n48350 = n12397 | n23327 ;
  assign n48351 = n48350 ^ n459 ^ 1'b0 ;
  assign n48352 = n12947 ^ n8901 ^ 1'b0 ;
  assign n48353 = n28694 ^ n959 ^ 1'b0 ;
  assign n48354 = n3732 & ~n48353 ;
  assign n48355 = n2760 & ~n17707 ;
  assign n48356 = ~n40622 & n48355 ;
  assign n48357 = n28360 ^ n302 ^ 1'b0 ;
  assign n48358 = n13519 & ~n48357 ;
  assign n48359 = n8408 & n48358 ;
  assign n48360 = n48356 & n48359 ;
  assign n48361 = n2211 & n47793 ;
  assign n48362 = n48361 ^ n47970 ^ 1'b0 ;
  assign n48363 = n6498 ^ n2051 ^ n1984 ;
  assign n48364 = n48363 ^ n29958 ^ 1'b0 ;
  assign n48365 = n19466 & n48364 ;
  assign n48366 = ~n24055 & n29700 ;
  assign n48367 = n14551 ^ n3669 ^ 1'b0 ;
  assign n48368 = ~n4121 & n48367 ;
  assign n48369 = n21021 ^ n15690 ^ 1'b0 ;
  assign n48370 = n354 & ~n24790 ;
  assign n48371 = n26302 ^ n22133 ^ 1'b0 ;
  assign n48372 = n22051 & n39688 ;
  assign n48373 = ~n11913 & n48372 ;
  assign n48374 = n39538 ^ n5443 ^ 1'b0 ;
  assign n48375 = ~n15380 & n25978 ;
  assign n48376 = n48375 ^ n37511 ^ n12902 ;
  assign n48377 = ( n4264 & ~n23520 ) | ( n4264 & n28767 ) | ( ~n23520 & n28767 ) ;
  assign n48378 = n27573 ^ n7766 ^ 1'b0 ;
  assign n48379 = ~n48377 & n48378 ;
  assign n48380 = n48379 ^ n34942 ^ 1'b0 ;
  assign n48381 = n9023 & n48380 ;
  assign n48382 = n48381 ^ n6955 ^ 1'b0 ;
  assign n48385 = ~n1908 & n44193 ;
  assign n48386 = n27016 & n48385 ;
  assign n48383 = n36388 ^ n26200 ^ 1'b0 ;
  assign n48384 = n19514 | n48383 ;
  assign n48387 = n48386 ^ n48384 ^ 1'b0 ;
  assign n48388 = n46740 ^ n32509 ^ n5111 ;
  assign n48389 = n48388 ^ n2719 ^ 1'b0 ;
  assign n48390 = n20030 ^ n12315 ^ 1'b0 ;
  assign n48391 = n14612 & n48390 ;
  assign n48392 = n17759 ^ n1202 ^ 1'b0 ;
  assign n48393 = n48391 & n48392 ;
  assign n48394 = n39879 ^ n23110 ^ 1'b0 ;
  assign n48395 = n3132 | n48394 ;
  assign n48396 = ( n3370 & n3425 ) | ( n3370 & n13031 ) | ( n3425 & n13031 ) ;
  assign n48397 = n21963 | n48396 ;
  assign n48398 = n6229 & n41923 ;
  assign n48399 = n46892 ^ n19300 ^ 1'b0 ;
  assign n48400 = n14460 ^ n12537 ^ 1'b0 ;
  assign n48401 = ~n2388 & n48400 ;
  assign n48402 = n11194 & n40404 ;
  assign n48403 = n8448 | n15877 ;
  assign n48404 = n48403 ^ n34644 ^ 1'b0 ;
  assign n48405 = n14939 | n15867 ;
  assign n48406 = n1829 | n48405 ;
  assign n48407 = n48406 ^ n9503 ^ 1'b0 ;
  assign n48408 = n5887 | n47367 ;
  assign n48409 = n48408 ^ n12414 ^ 1'b0 ;
  assign n48410 = n48409 ^ n18360 ^ 1'b0 ;
  assign n48411 = ~n25555 & n48410 ;
  assign n48412 = n14961 & n22714 ;
  assign n48413 = n21008 ^ n19967 ^ 1'b0 ;
  assign n48414 = n5553 & n15115 ;
  assign n48415 = n24518 & n48414 ;
  assign n48416 = n22209 & ~n32331 ;
  assign n48417 = n48416 ^ n12449 ^ 1'b0 ;
  assign n48418 = n12988 & n33898 ;
  assign n48419 = n29695 & n47244 ;
  assign n48424 = n1469 & n44698 ;
  assign n48421 = n5319 & n13848 ;
  assign n48422 = n14772 & n48421 ;
  assign n48420 = ~n19277 & n40270 ;
  assign n48423 = n48422 ^ n48420 ^ 1'b0 ;
  assign n48425 = n48424 ^ n48423 ^ 1'b0 ;
  assign n48427 = n623 & n8249 ;
  assign n48428 = n18062 & n48427 ;
  assign n48426 = n2670 & ~n24683 ;
  assign n48429 = n48428 ^ n48426 ^ 1'b0 ;
  assign n48430 = n8853 | n12916 ;
  assign n48431 = n9201 & ~n25231 ;
  assign n48432 = n48431 ^ n3246 ^ 1'b0 ;
  assign n48433 = ~n30914 & n33482 ;
  assign n48434 = n39497 ^ n35596 ^ 1'b0 ;
  assign n48435 = n42478 & n48434 ;
  assign n48436 = n48435 ^ n7953 ^ 1'b0 ;
  assign n48437 = n37432 ^ n26804 ^ 1'b0 ;
  assign n48438 = n1246 & n48437 ;
  assign n48439 = n5268 & n48438 ;
  assign n48440 = n224 & n48439 ;
  assign n48441 = ( ~n19324 & n44971 ) | ( ~n19324 & n48440 ) | ( n44971 & n48440 ) ;
  assign n48442 = ( ~n408 & n6776 ) | ( ~n408 & n8219 ) | ( n6776 & n8219 ) ;
  assign n48443 = n28064 & n48442 ;
  assign n48444 = n5893 & n48443 ;
  assign n48445 = n31626 ^ n2151 ^ 1'b0 ;
  assign n48446 = n10189 & n19766 ;
  assign n48447 = n48446 ^ n31426 ^ 1'b0 ;
  assign n48448 = n27878 ^ n8467 ^ 1'b0 ;
  assign n48449 = n45130 ^ n36480 ^ 1'b0 ;
  assign n48450 = ~n17449 & n37832 ;
  assign n48451 = ~n13941 & n48450 ;
  assign n48452 = n34229 ^ n8948 ^ 1'b0 ;
  assign n48453 = n2885 & ~n48452 ;
  assign n48454 = n28449 ^ n11458 ^ 1'b0 ;
  assign n48455 = n48454 ^ n26714 ^ n7325 ;
  assign n48456 = n5902 | n44015 ;
  assign n48457 = n48456 ^ n22695 ^ 1'b0 ;
  assign n48458 = n25452 & ~n48457 ;
  assign n48459 = n27509 ^ n18307 ^ 1'b0 ;
  assign n48460 = ~n20505 & n48459 ;
  assign n48461 = ~n3009 & n5344 ;
  assign n48462 = n2802 ^ n205 ^ 1'b0 ;
  assign n48463 = n9165 & n48462 ;
  assign n48464 = n48463 ^ n20041 ^ 1'b0 ;
  assign n48465 = n7507 ^ n4121 ^ 1'b0 ;
  assign n48466 = n23816 | n48465 ;
  assign n48467 = n43205 ^ n8296 ^ 1'b0 ;
  assign n48468 = n48466 & n48467 ;
  assign n48469 = n3044 | n19789 ;
  assign n48470 = n8414 & ~n48469 ;
  assign n48471 = n3284 | n12938 ;
  assign n48472 = ( n725 & ~n24169 ) | ( n725 & n48471 ) | ( ~n24169 & n48471 ) ;
  assign n48473 = n4034 & ~n13568 ;
  assign n48474 = ~n6035 & n48473 ;
  assign n48475 = ( ~n20559 & n24688 ) | ( ~n20559 & n48474 ) | ( n24688 & n48474 ) ;
  assign n48476 = n44520 ^ n27214 ^ 1'b0 ;
  assign n48477 = n16692 & n48476 ;
  assign n48478 = n16824 & ~n25022 ;
  assign n48479 = n26875 & n48478 ;
  assign n48480 = n7568 & n44082 ;
  assign n48481 = ~n23483 & n27092 ;
  assign n48485 = ~n13707 & n32811 ;
  assign n48486 = n20858 & n48485 ;
  assign n48482 = n16364 & ~n45226 ;
  assign n48483 = n48482 ^ n22796 ^ 1'b0 ;
  assign n48484 = n48483 ^ n15828 ^ 1'b0 ;
  assign n48487 = n48486 ^ n48484 ^ 1'b0 ;
  assign n48488 = n24911 ^ n20791 ^ 1'b0 ;
  assign n48489 = ~n18777 & n48488 ;
  assign n48490 = n25691 ^ n3962 ^ 1'b0 ;
  assign n48491 = n19759 & n27039 ;
  assign n48492 = ~n21488 & n48491 ;
  assign n48493 = n23627 ^ n19297 ^ 1'b0 ;
  assign n48494 = n7001 | n48493 ;
  assign n48495 = n48494 ^ n46535 ^ 1'b0 ;
  assign n48496 = n19980 | n25919 ;
  assign n48497 = n48496 ^ n2072 ^ 1'b0 ;
  assign n48498 = n35470 ^ n17343 ^ 1'b0 ;
  assign n48499 = n27516 ^ n3445 ^ 1'b0 ;
  assign n48500 = n48498 & n48499 ;
  assign n48501 = n30115 ^ n24624 ^ 1'b0 ;
  assign n48502 = ~n2486 & n48501 ;
  assign n48503 = n8173 ^ n6769 ^ 1'b0 ;
  assign n48504 = ( n2883 & ~n14896 ) | ( n2883 & n48503 ) | ( ~n14896 & n48503 ) ;
  assign n48505 = n43215 ^ n14474 ^ 1'b0 ;
  assign n48506 = ~n26414 & n31732 ;
  assign n48507 = n48505 & n48506 ;
  assign n48508 = n12634 ^ n10616 ^ n983 ;
  assign n48509 = n26602 | n48508 ;
  assign n48510 = n19300 & ~n48509 ;
  assign n48511 = n48510 ^ n26430 ^ 1'b0 ;
  assign n48512 = n23754 ^ n1186 ^ 1'b0 ;
  assign n48513 = n22242 | n48512 ;
  assign n48514 = ~n7933 & n18154 ;
  assign n48515 = n12018 & ~n29297 ;
  assign n48516 = n42298 ^ n41024 ^ 1'b0 ;
  assign n48517 = ~n42797 & n48516 ;
  assign n48518 = n1980 & n18990 ;
  assign n48519 = n48518 ^ n9282 ^ 1'b0 ;
  assign n48520 = n11855 & ~n48519 ;
  assign n48521 = n21569 ^ n13509 ^ 1'b0 ;
  assign n48522 = n949 & ~n11309 ;
  assign n48523 = n48522 ^ n40972 ^ 1'b0 ;
  assign n48524 = ~n1933 & n10033 ;
  assign n48525 = n4788 ^ n3218 ^ 1'b0 ;
  assign n48526 = ~n33962 & n48525 ;
  assign n48527 = n4881 | n48526 ;
  assign n48528 = n5276 & n41170 ;
  assign n48529 = n48528 ^ n12740 ^ 1'b0 ;
  assign n48530 = n36559 ^ n11701 ^ 1'b0 ;
  assign n48531 = n5084 & ~n10159 ;
  assign n48532 = ~n2838 & n18111 ;
  assign n48533 = n48531 & n48532 ;
  assign n48534 = n4521 & n48533 ;
  assign n48535 = n23645 ^ n1743 ^ 1'b0 ;
  assign n48536 = n12516 | n48535 ;
  assign n48537 = n48536 ^ n8326 ^ 1'b0 ;
  assign n48538 = n26667 ^ n8529 ^ 1'b0 ;
  assign n48539 = n5805 & ~n48538 ;
  assign n48540 = n48539 ^ n23544 ^ 1'b0 ;
  assign n48541 = n26732 & ~n30262 ;
  assign n48542 = n38881 & n48541 ;
  assign n48543 = n28985 ^ n18027 ^ 1'b0 ;
  assign n48544 = n14933 | n48543 ;
  assign n48545 = n36312 ^ n6195 ^ 1'b0 ;
  assign n48546 = n33205 ^ n26009 ^ 1'b0 ;
  assign n48547 = n5458 & n48546 ;
  assign n48548 = n8915 & n13694 ;
  assign n48549 = n47474 ^ n24328 ^ 1'b0 ;
  assign n48550 = ( ~n1157 & n3349 ) | ( ~n1157 & n19039 ) | ( n3349 & n19039 ) ;
  assign n48551 = ( n1517 & n4390 ) | ( n1517 & n48550 ) | ( n4390 & n48550 ) ;
  assign n48552 = n36154 ^ n10603 ^ n4525 ;
  assign n48553 = n4044 & ~n48552 ;
  assign n48554 = ~n41516 & n44296 ;
  assign n48555 = ~n29007 & n48554 ;
  assign n48556 = ~n3464 & n5655 ;
  assign n48557 = ~n6815 & n9532 ;
  assign n48558 = ~n23936 & n48557 ;
  assign n48559 = n3462 ^ n753 ^ 1'b0 ;
  assign n48560 = n791 | n15180 ;
  assign n48561 = n22135 & ~n48560 ;
  assign n48562 = n6488 ^ n1981 ^ 1'b0 ;
  assign n48563 = ~n18485 & n18674 ;
  assign n48564 = n48563 ^ x7 ^ 1'b0 ;
  assign n48565 = n8265 & n48564 ;
  assign n48567 = n2108 & n11430 ;
  assign n48566 = n920 & n2085 ;
  assign n48568 = n48567 ^ n48566 ^ 1'b0 ;
  assign n48569 = n30332 & ~n48568 ;
  assign n48570 = n6655 | n28170 ;
  assign n48571 = ( ~n13245 & n14957 ) | ( ~n13245 & n48570 ) | ( n14957 & n48570 ) ;
  assign n48572 = n26738 ^ n26541 ^ 1'b0 ;
  assign n48573 = n26549 ^ n14616 ^ 1'b0 ;
  assign n48574 = n12405 | n28476 ;
  assign n48575 = n48574 ^ n41634 ^ 1'b0 ;
  assign n48576 = n48575 ^ n8738 ^ 1'b0 ;
  assign n48577 = n48573 & n48576 ;
  assign n48578 = n1794 & n48577 ;
  assign n48579 = n1237 | n46346 ;
  assign n48580 = n3792 & ~n48579 ;
  assign n48581 = n15246 ^ n3772 ^ 1'b0 ;
  assign n48582 = n18232 & n48581 ;
  assign n48583 = n45525 ^ n34427 ^ n30447 ;
  assign n48584 = n5151 ^ n519 ^ 1'b0 ;
  assign n48585 = ~n6623 & n48584 ;
  assign n48586 = n10530 & ~n14642 ;
  assign n48587 = n34326 & n48586 ;
  assign n48588 = n48585 | n48587 ;
  assign n48589 = ~n6289 & n48588 ;
  assign n48590 = ~n13685 & n29846 ;
  assign n48591 = n12611 | n48590 ;
  assign n48592 = n46503 ^ n8246 ^ 1'b0 ;
  assign n48593 = n20709 ^ n15824 ^ n2986 ;
  assign n48594 = n11476 ^ n5425 ^ 1'b0 ;
  assign n48595 = n18185 ^ n2550 ^ 1'b0 ;
  assign n48596 = n8299 & ~n26436 ;
  assign n48597 = ~n19784 & n48596 ;
  assign n48598 = n48597 ^ n27940 ^ 1'b0 ;
  assign n48599 = n6488 & ~n48598 ;
  assign n48600 = ~n7624 & n17015 ;
  assign n48601 = ~n11501 & n48600 ;
  assign n48602 = n48601 ^ n20816 ^ 1'b0 ;
  assign n48603 = n10893 & n36334 ;
  assign n48604 = n729 & ~n7001 ;
  assign n48605 = n48604 ^ n3114 ^ 1'b0 ;
  assign n48606 = n4845 & n26975 ;
  assign n48607 = n48606 ^ n7360 ^ 1'b0 ;
  assign n48608 = n29965 & n47793 ;
  assign n48609 = n48608 ^ n6179 ^ 1'b0 ;
  assign n48610 = n3562 & ~n12248 ;
  assign n48611 = n48610 ^ n15594 ^ 1'b0 ;
  assign n48612 = n14785 & ~n48611 ;
  assign n48613 = n40404 ^ n26200 ^ 1'b0 ;
  assign n48614 = ~n42844 & n48613 ;
  assign n48615 = n5073 | n29294 ;
  assign n48616 = n48615 ^ n2382 ^ 1'b0 ;
  assign n48617 = ~n3096 & n12368 ;
  assign n48618 = ~n48616 & n48617 ;
  assign n48619 = n492 & ~n18435 ;
  assign n48620 = n48619 ^ n11583 ^ 1'b0 ;
  assign n48621 = n3858 | n41074 ;
  assign n48622 = ~n5334 & n27466 ;
  assign n48623 = ( n148 & ~n10488 ) | ( n148 & n42356 ) | ( ~n10488 & n42356 ) ;
  assign n48624 = n48623 ^ n2649 ^ 1'b0 ;
  assign n48625 = n34446 & n48624 ;
  assign n48626 = n27407 ^ n23772 ^ n11692 ;
  assign n48627 = n944 & n24316 ;
  assign n48628 = n21501 | n48627 ;
  assign n48629 = n48628 ^ n1568 ^ 1'b0 ;
  assign n48630 = n24709 | n25020 ;
  assign n48631 = n47416 ^ n6291 ^ n1975 ;
  assign n48632 = n48631 ^ n4199 ^ 1'b0 ;
  assign n48633 = n20157 ^ n551 ^ 1'b0 ;
  assign n48634 = n571 & ~n18042 ;
  assign n48635 = n48634 ^ n26 ^ 1'b0 ;
  assign n48636 = n13130 | n42351 ;
  assign n48637 = n48636 ^ n14071 ^ 1'b0 ;
  assign n48638 = n48637 ^ n19277 ^ n2146 ;
  assign n48639 = n22382 ^ n8126 ^ 1'b0 ;
  assign n48640 = n8019 & n48639 ;
  assign n48641 = ~n46392 & n48640 ;
  assign n48642 = ~n892 & n48641 ;
  assign n48643 = ~n4416 & n15581 ;
  assign n48644 = n25379 ^ n2093 ^ 1'b0 ;
  assign n48645 = n24120 | n48644 ;
  assign n48646 = n42792 ^ n362 ^ 1'b0 ;
  assign n48647 = ~n1842 & n3510 ;
  assign n48648 = n48647 ^ n21903 ^ 1'b0 ;
  assign n48649 = ~n6528 & n48648 ;
  assign n48650 = n16724 | n43036 ;
  assign n48651 = ~n7498 & n17781 ;
  assign n48652 = n22903 & n48651 ;
  assign n48653 = n48652 ^ n423 ^ 1'b0 ;
  assign n48654 = n7739 & n48653 ;
  assign n48655 = n436 & ~n16083 ;
  assign n48656 = n10653 ^ n5342 ^ n780 ;
  assign n48657 = n35488 ^ n4367 ^ 1'b0 ;
  assign n48658 = n8879 & n22968 ;
  assign n48659 = n33164 ^ n13309 ^ 1'b0 ;
  assign n48660 = n21514 | n39378 ;
  assign n48661 = n48659 | n48660 ;
  assign n48662 = n4040 | n19097 ;
  assign n48663 = n48662 ^ n9271 ^ 1'b0 ;
  assign n48664 = n48663 ^ n18635 ^ 1'b0 ;
  assign n48665 = n3228 & ~n12142 ;
  assign n48666 = n28225 & n48665 ;
  assign n48667 = n20798 | n46330 ;
  assign n48668 = n30026 ^ n6716 ^ 1'b0 ;
  assign n48669 = n1742 & ~n48668 ;
  assign n48670 = ~n1212 & n18199 ;
  assign n48671 = n7507 & ~n22541 ;
  assign n48672 = n7645 & ~n48671 ;
  assign n48673 = n12030 | n41023 ;
  assign n48674 = n8391 & ~n22044 ;
  assign n48675 = n6413 | n48674 ;
  assign n48676 = ~n15919 & n24886 ;
  assign n48677 = n16308 | n17488 ;
  assign n48678 = n48677 ^ n16795 ^ n9823 ;
  assign n48679 = n9564 & n23600 ;
  assign n48680 = n28764 & ~n48679 ;
  assign n48681 = ~n25388 & n48680 ;
  assign n48682 = n18165 ^ n16394 ^ 1'b0 ;
  assign n48683 = n901 | n29553 ;
  assign n48684 = n38505 ^ n11390 ^ 1'b0 ;
  assign n48685 = n10031 ^ n4419 ^ 1'b0 ;
  assign n48686 = ~n30259 & n35539 ;
  assign n48687 = ( n16898 & n18458 ) | ( n16898 & n33702 ) | ( n18458 & n33702 ) ;
  assign n48688 = ( n16846 & ~n17436 ) | ( n16846 & n48687 ) | ( ~n17436 & n48687 ) ;
  assign n48689 = ~n2504 & n3139 ;
  assign n48690 = ~n3139 & n48689 ;
  assign n48691 = n10498 | n48690 ;
  assign n48692 = n48690 & ~n48691 ;
  assign n48693 = n48692 ^ n9491 ^ n3041 ;
  assign n48694 = n4794 & ~n13042 ;
  assign n48695 = n41006 ^ n34046 ^ 1'b0 ;
  assign n48696 = ~n8136 & n8413 ;
  assign n48697 = n14832 & n25470 ;
  assign n48698 = n21632 | n36352 ;
  assign n48699 = n48698 ^ n601 ^ 1'b0 ;
  assign n48700 = n43949 ^ n11650 ^ n7926 ;
  assign n48701 = n9014 | n9860 ;
  assign n48702 = n23741 ^ n3744 ^ 1'b0 ;
  assign n48703 = n1724 | n40476 ;
  assign n48704 = n8252 | n28672 ;
  assign n48705 = n340 & ~n38164 ;
  assign n48706 = n9455 ^ n3071 ^ 1'b0 ;
  assign n48707 = n48706 ^ n36524 ^ n565 ;
  assign n48708 = n34500 ^ n12793 ^ n6507 ;
  assign n48709 = n24131 ^ n3003 ^ 1'b0 ;
  assign n48710 = n21816 & ~n48709 ;
  assign n48711 = n1430 | n48710 ;
  assign n48713 = n14066 ^ n9557 ^ 1'b0 ;
  assign n48712 = ( n5719 & n7478 ) | ( n5719 & n17189 ) | ( n7478 & n17189 ) ;
  assign n48714 = n48713 ^ n48712 ^ 1'b0 ;
  assign n48715 = ~n6216 & n38466 ;
  assign n48716 = n30322 ^ n13893 ^ n8973 ;
  assign n48717 = n6237 & ~n29580 ;
  assign n48718 = n8608 & ~n9687 ;
  assign n48719 = n48718 ^ n17439 ^ 1'b0 ;
  assign n48720 = n42254 ^ n22469 ^ n1007 ;
  assign n48721 = n3917 | n48720 ;
  assign n48722 = n48721 ^ n13304 ^ 1'b0 ;
  assign n48723 = n47434 ^ n46260 ^ 1'b0 ;
  assign n48724 = n11909 & n26966 ;
  assign n48725 = ~n21411 & n48724 ;
  assign n48726 = n48725 ^ n34277 ^ 1'b0 ;
  assign n48727 = n5155 & n48726 ;
  assign n48728 = ~n26678 & n48727 ;
  assign n48729 = ~n10944 & n48728 ;
  assign n48730 = n45801 ^ n16453 ^ 1'b0 ;
  assign n48731 = ~n36822 & n48730 ;
  assign n48732 = n20840 ^ n7626 ^ 1'b0 ;
  assign n48733 = n29579 & ~n48732 ;
  assign n48734 = n48733 ^ n15865 ^ 1'b0 ;
  assign n48735 = n18092 ^ n14976 ^ 1'b0 ;
  assign n48736 = n277 | n1647 ;
  assign n48737 = ~n11691 & n14805 ;
  assign n48738 = ( n13232 & n30101 ) | ( n13232 & ~n48737 ) | ( n30101 & ~n48737 ) ;
  assign n48739 = n16597 | n19069 ;
  assign n48740 = n9405 | n48739 ;
  assign n48741 = ~n1075 & n48740 ;
  assign n48742 = ~n48738 & n48741 ;
  assign n48743 = n38557 ^ n6838 ^ 1'b0 ;
  assign n48744 = ~n1786 & n10312 ;
  assign n48745 = ~n7963 & n48744 ;
  assign n48746 = n26488 ^ n7238 ^ 1'b0 ;
  assign n48747 = n34030 & n48746 ;
  assign n48748 = n16894 ^ n8513 ^ 1'b0 ;
  assign n48749 = ( n48745 & n48747 ) | ( n48745 & n48748 ) | ( n48747 & n48748 ) ;
  assign n48750 = ~n4688 & n6575 ;
  assign n48751 = ~n9795 & n13097 ;
  assign n48752 = n48750 & n48751 ;
  assign n48753 = n11468 & n48752 ;
  assign n48754 = n46517 ^ n7508 ^ 1'b0 ;
  assign n48755 = n4092 & ~n7766 ;
  assign n48756 = n48754 & n48755 ;
  assign n48757 = n2413 | n6966 ;
  assign n48758 = ( ~n10107 & n46371 ) | ( ~n10107 & n48757 ) | ( n46371 & n48757 ) ;
  assign n48759 = ~n13167 & n27638 ;
  assign n48760 = n48759 ^ n8363 ^ 1'b0 ;
  assign n48762 = n24517 ^ n226 ^ 1'b0 ;
  assign n48763 = n10306 | n48762 ;
  assign n48761 = ~n6833 & n7989 ;
  assign n48764 = n48763 ^ n48761 ^ 1'b0 ;
  assign n48765 = n34559 | n34873 ;
  assign n48766 = n48764 | n48765 ;
  assign n48767 = n35652 ^ n19151 ^ 1'b0 ;
  assign n48768 = n25024 ^ n12049 ^ 1'b0 ;
  assign n48769 = n2068 | n48768 ;
  assign n48770 = n14976 & n48769 ;
  assign n48771 = n48767 & n48770 ;
  assign n48772 = n4444 & ~n8946 ;
  assign n48773 = n15278 & n48772 ;
  assign n48774 = n48773 ^ n26618 ^ 1'b0 ;
  assign n48775 = ~n14787 & n45022 ;
  assign n48776 = ~n48774 & n48775 ;
  assign n48777 = ~n16490 & n36625 ;
  assign n48778 = ( n3060 & ~n6095 ) | ( n3060 & n48777 ) | ( ~n6095 & n48777 ) ;
  assign n48779 = n14378 | n17563 ;
  assign n48780 = n26480 & ~n48779 ;
  assign n48781 = n6741 | n45400 ;
  assign n48782 = n432 & ~n17596 ;
  assign n48783 = n48781 & n48782 ;
  assign n48784 = ~n10885 & n37878 ;
  assign n48785 = n45186 ^ n13460 ^ 1'b0 ;
  assign n48786 = n48784 | n48785 ;
  assign n48787 = n29590 ^ n12565 ^ n12451 ;
  assign n48788 = n16157 ^ n8506 ^ 1'b0 ;
  assign n48789 = n13896 ^ n11852 ^ 1'b0 ;
  assign n48790 = ~n30464 & n48789 ;
  assign n48791 = n22779 ^ n2304 ^ 1'b0 ;
  assign n48792 = n10728 & n48791 ;
  assign n48793 = n48792 ^ n19821 ^ 1'b0 ;
  assign n48794 = ( n11439 & ~n37882 ) | ( n11439 & n42554 ) | ( ~n37882 & n42554 ) ;
  assign n48795 = n802 & n12494 ;
  assign n48796 = n159 | n48795 ;
  assign n48797 = ( n22959 & ~n48794 ) | ( n22959 & n48796 ) | ( ~n48794 & n48796 ) ;
  assign n48798 = n10603 & ~n19220 ;
  assign n48799 = n9606 ^ n3788 ^ 1'b0 ;
  assign n48800 = n2310 | n48799 ;
  assign n48801 = n30557 & ~n48425 ;
  assign n48802 = n48801 ^ n23108 ^ 1'b0 ;
  assign n48803 = n9343 & ~n23509 ;
  assign n48804 = n34157 & ~n48803 ;
  assign n48805 = ( ~n7739 & n17133 ) | ( ~n7739 & n19225 ) | ( n17133 & n19225 ) ;
  assign n48806 = n48805 ^ n17962 ^ 1'b0 ;
  assign n48807 = n48804 & ~n48806 ;
  assign n48808 = n1342 | n14085 ;
  assign n48809 = n14085 & ~n48808 ;
  assign n48810 = n21672 | n48809 ;
  assign n48811 = n48810 ^ n23593 ^ 1'b0 ;
  assign n48812 = n12609 ^ n2086 ^ 1'b0 ;
  assign n48813 = n48811 | n48812 ;
  assign n48814 = n48813 ^ n11692 ^ 1'b0 ;
  assign n48815 = n9927 ^ n4351 ^ 1'b0 ;
  assign n48816 = n35930 | n48815 ;
  assign n48817 = n38496 & ~n42095 ;
  assign n48818 = n9478 & n20133 ;
  assign n48819 = n4814 & n9196 ;
  assign n48820 = n7713 | n48819 ;
  assign n48821 = n48820 ^ n37515 ^ 1'b0 ;
  assign n48822 = n875 & n27251 ;
  assign n48823 = n17714 & n41787 ;
  assign n48824 = n48823 ^ n12503 ^ 1'b0 ;
  assign n48825 = n14546 ^ n924 ^ 1'b0 ;
  assign n48826 = n15457 & n39756 ;
  assign n48827 = n42838 | n46606 ;
  assign n48828 = n48827 ^ n2872 ^ 1'b0 ;
  assign n48829 = n19675 ^ n5942 ^ 1'b0 ;
  assign n48830 = ( n283 & ~n4977 ) | ( n283 & n36527 ) | ( ~n4977 & n36527 ) ;
  assign n48831 = n15324 & ~n36819 ;
  assign n48832 = n35204 | n48831 ;
  assign n48833 = n13 | n17191 ;
  assign n48834 = n13044 | n48833 ;
  assign n48835 = n25046 ^ n10975 ^ 1'b0 ;
  assign n48836 = n25553 & ~n48835 ;
  assign n48837 = n18416 | n18878 ;
  assign n48838 = n12977 & n13285 ;
  assign n48839 = n42421 & n48838 ;
  assign n48840 = n25452 & n32172 ;
  assign n48841 = n7399 & n48840 ;
  assign n48842 = n48841 ^ n7921 ^ 1'b0 ;
  assign n48843 = n2520 | n24438 ;
  assign n48844 = n15707 & n37650 ;
  assign n48845 = n48844 ^ n42721 ^ 1'b0 ;
  assign n48846 = n34401 & ~n35764 ;
  assign n48847 = n16301 ^ n11927 ^ 1'b0 ;
  assign n48848 = n4170 & n42407 ;
  assign n48849 = ~n41956 & n48848 ;
  assign n48850 = n9158 ^ n6013 ^ 1'b0 ;
  assign n48851 = ~n15446 & n48850 ;
  assign n48852 = n48851 ^ n1395 ^ 1'b0 ;
  assign n48853 = n14343 | n48852 ;
  assign n48854 = n18493 & n19627 ;
  assign n48855 = n4399 ^ n806 ^ 1'b0 ;
  assign n48856 = ( n7516 & n12732 ) | ( n7516 & n48855 ) | ( n12732 & n48855 ) ;
  assign n48857 = n47852 ^ n30324 ^ 1'b0 ;
  assign n48858 = ~n33973 & n48857 ;
  assign n48859 = n21668 & n35602 ;
  assign n48860 = n48859 ^ n31275 ^ 1'b0 ;
  assign n48861 = n620 & n28726 ;
  assign n48862 = n27269 & n48861 ;
  assign n48863 = ~n48860 & n48862 ;
  assign n48864 = ( n12324 & n15175 ) | ( n12324 & n40523 ) | ( n15175 & n40523 ) ;
  assign n48865 = n44423 ^ n20740 ^ 1'b0 ;
  assign n48866 = n24071 & n48865 ;
  assign n48867 = n24597 ^ n17470 ^ 1'b0 ;
  assign n48868 = n7624 | n18544 ;
  assign n48869 = n12320 | n48868 ;
  assign n48870 = n23775 ^ n4434 ^ 1'b0 ;
  assign n48871 = n4146 & ~n48870 ;
  assign n48872 = n48871 ^ n38455 ^ 1'b0 ;
  assign n48873 = n10668 | n23142 ;
  assign n48874 = n48873 ^ n44901 ^ 1'b0 ;
  assign n48875 = n125 & ~n21878 ;
  assign n48876 = n32665 ^ n6307 ^ 1'b0 ;
  assign n48877 = n25283 | n48876 ;
  assign n48878 = n3556 ^ n188 ^ 1'b0 ;
  assign n48879 = n31301 & ~n48878 ;
  assign n48880 = n35726 & n48879 ;
  assign n48881 = n48877 & n48880 ;
  assign n48882 = n14080 ^ n8057 ^ 1'b0 ;
  assign n48883 = ~n21339 & n40349 ;
  assign n48884 = ~n548 & n16268 ;
  assign n48885 = n47679 | n48884 ;
  assign n48886 = n13114 ^ n11355 ^ n115 ;
  assign n48887 = ( ~n4914 & n20213 ) | ( ~n4914 & n48886 ) | ( n20213 & n48886 ) ;
  assign n48888 = n8387 & ~n29160 ;
  assign n48889 = ~n23785 & n25771 ;
  assign n48890 = n16400 & n48889 ;
  assign n48891 = n30204 & ~n34302 ;
  assign n48892 = n48891 ^ n4005 ^ 1'b0 ;
  assign n48896 = n40957 ^ n20577 ^ n16067 ;
  assign n48897 = n30217 & n48896 ;
  assign n48893 = n1574 & n39092 ;
  assign n48894 = n1389 & n48893 ;
  assign n48895 = n9148 | n48894 ;
  assign n48898 = n48897 ^ n48895 ^ 1'b0 ;
  assign n48899 = ~n30065 & n48898 ;
  assign n48900 = n27717 ^ n17849 ^ 1'b0 ;
  assign n48901 = n11383 & ~n29514 ;
  assign n48902 = n48901 ^ n43499 ^ n30751 ;
  assign n48903 = n9624 & n32781 ;
  assign n48904 = n13251 & ~n34645 ;
  assign n48905 = ~n40664 & n48904 ;
  assign n48907 = n7977 ^ n7539 ^ 1'b0 ;
  assign n48908 = ~n13582 & n48907 ;
  assign n48909 = n42106 ^ n493 ^ 1'b0 ;
  assign n48910 = n48908 & n48909 ;
  assign n48906 = n667 | n31372 ;
  assign n48911 = n48910 ^ n48906 ^ 1'b0 ;
  assign n48912 = n14890 | n15694 ;
  assign n48913 = ~n12651 & n47227 ;
  assign n48914 = n30405 & n48913 ;
  assign n48915 = n6264 | n39321 ;
  assign n48916 = n1783 | n48915 ;
  assign n48917 = n48916 ^ n10320 ^ 1'b0 ;
  assign n48919 = n44535 ^ n8478 ^ 1'b0 ;
  assign n48918 = n43876 ^ n19844 ^ 1'b0 ;
  assign n48920 = n48919 ^ n48918 ^ n31230 ;
  assign n48921 = ~n1172 & n20725 ;
  assign n48922 = ~n1122 & n12559 ;
  assign n48923 = ~n40630 & n42097 ;
  assign n48924 = ~n48922 & n48923 ;
  assign n48925 = ~n7307 & n9479 ;
  assign n48926 = ( n1460 & ~n2551 ) | ( n1460 & n6099 ) | ( ~n2551 & n6099 ) ;
  assign n48927 = n2050 | n6059 ;
  assign n48928 = n253 | n48927 ;
  assign n48929 = ~n39038 & n48928 ;
  assign n48930 = n48929 ^ n22633 ^ 1'b0 ;
  assign n48931 = n11860 & n48930 ;
  assign n48932 = n48926 | n48931 ;
  assign n48933 = n782 | n48932 ;
  assign n48934 = n31343 ^ n8265 ^ 1'b0 ;
  assign n48935 = n48933 & ~n48934 ;
  assign n48936 = n183 | n3209 ;
  assign n48937 = n33458 | n48936 ;
  assign n48938 = n48937 ^ n16305 ^ 1'b0 ;
  assign n48939 = n18412 ^ n1609 ^ 1'b0 ;
  assign n48940 = n6833 | n27578 ;
  assign n48941 = n10158 | n48940 ;
  assign n48942 = ( n22313 & n23142 ) | ( n22313 & n48941 ) | ( n23142 & n48941 ) ;
  assign n48943 = n8705 ^ n4226 ^ 1'b0 ;
  assign n48944 = n7524 ^ n5812 ^ 1'b0 ;
  assign n48945 = ~n6598 & n6813 ;
  assign n48946 = n22937 | n48945 ;
  assign n48950 = n484 & ~n8567 ;
  assign n48951 = n2494 & ~n48950 ;
  assign n48947 = n2910 & ~n10073 ;
  assign n48948 = n48947 ^ n23351 ^ 1'b0 ;
  assign n48949 = n12458 | n48948 ;
  assign n48952 = n48951 ^ n48949 ^ 1'b0 ;
  assign n48953 = n5473 | n22332 ;
  assign n48954 = n6297 & ~n15695 ;
  assign n48955 = n48954 ^ n8721 ^ 1'b0 ;
  assign n48956 = ~n10443 & n48955 ;
  assign n48957 = n48956 ^ n13219 ^ 1'b0 ;
  assign n48958 = n9769 | n48957 ;
  assign n48959 = n12678 ^ n12119 ^ 1'b0 ;
  assign n48960 = n7803 & ~n10780 ;
  assign n48961 = n48960 ^ n2478 ^ 1'b0 ;
  assign n48962 = ~n33106 & n48961 ;
  assign n48963 = n4581 | n16650 ;
  assign n48964 = n32925 ^ n16707 ^ 1'b0 ;
  assign n48965 = ~n8138 & n48964 ;
  assign n48966 = n48965 ^ n12812 ^ 1'b0 ;
  assign n48967 = n17421 & ~n48966 ;
  assign n48968 = ( n2738 & n32880 ) | ( n2738 & n48967 ) | ( n32880 & n48967 ) ;
  assign n48969 = n36401 ^ n13108 ^ 1'b0 ;
  assign n48970 = n731 & ~n48969 ;
  assign n48971 = n48970 ^ n2314 ^ 1'b0 ;
  assign n48972 = n13553 | n32604 ;
  assign n48973 = n48972 ^ n12119 ^ 1'b0 ;
  assign n48974 = n48973 ^ n582 ^ 1'b0 ;
  assign n48975 = ~n27871 & n48974 ;
  assign n48976 = n18662 ^ n8131 ^ 1'b0 ;
  assign n48977 = n44744 ^ n216 ^ 1'b0 ;
  assign n48978 = ~n48976 & n48977 ;
  assign n48981 = n4590 & n22448 ;
  assign n48982 = n48981 ^ n27625 ^ 1'b0 ;
  assign n48980 = ~n2566 & n13303 ;
  assign n48983 = n48982 ^ n48980 ^ 1'b0 ;
  assign n48979 = n10620 & ~n10758 ;
  assign n48984 = n48983 ^ n48979 ^ 1'b0 ;
  assign n48985 = ~n5161 & n27729 ;
  assign n48986 = n48985 ^ n31391 ^ 1'b0 ;
  assign n48987 = n3510 & ~n43939 ;
  assign n48988 = ~n19984 & n32505 ;
  assign n48989 = n21834 ^ n7953 ^ 1'b0 ;
  assign n48991 = n14905 ^ n14670 ^ 1'b0 ;
  assign n48992 = ~n42485 & n48991 ;
  assign n48990 = n4366 & n11144 ;
  assign n48993 = n48992 ^ n48990 ^ 1'b0 ;
  assign n48994 = n212 & ~n37663 ;
  assign n48995 = n37663 & n48994 ;
  assign n48996 = n14068 & ~n48995 ;
  assign n48997 = ~n14068 & n48996 ;
  assign n48998 = n46399 | n48997 ;
  assign n48999 = n48997 & ~n48998 ;
  assign n49000 = n2252 & ~n7645 ;
  assign n49001 = ( n16969 & n48999 ) | ( n16969 & n49000 ) | ( n48999 & n49000 ) ;
  assign n49002 = n3601 & n11170 ;
  assign n49003 = ~n42566 & n49002 ;
  assign n49004 = n16627 | n23003 ;
  assign n49005 = n6764 & ~n12053 ;
  assign n49006 = ~n2550 & n49005 ;
  assign n49007 = n14001 & n49006 ;
  assign n49011 = ~n12555 & n24075 ;
  assign n49012 = n49011 ^ n2202 ^ 1'b0 ;
  assign n49008 = n5755 | n15579 ;
  assign n49009 = ( ~n9351 & n14420 ) | ( ~n9351 & n49008 ) | ( n14420 & n49008 ) ;
  assign n49010 = n27534 & n49009 ;
  assign n49013 = n49012 ^ n49010 ^ 1'b0 ;
  assign n49014 = n1804 & n43084 ;
  assign n49015 = n32165 & n49014 ;
  assign n49016 = n11442 & ~n12126 ;
  assign n49017 = n49015 & n49016 ;
  assign n49018 = n49017 ^ n33637 ^ 1'b0 ;
  assign n49019 = n1745 & n49018 ;
  assign n49020 = n3447 ^ n2639 ^ 1'b0 ;
  assign n49021 = n15865 & n49020 ;
  assign n49022 = ~n22384 & n49021 ;
  assign n49023 = n2665 | n12591 ;
  assign n49024 = n8806 & n49023 ;
  assign n49025 = ~n2267 & n3580 ;
  assign n49026 = n49024 & n49025 ;
  assign n49027 = n2884 & ~n7338 ;
  assign n49028 = ~n8865 & n49027 ;
  assign n49029 = ( n2222 & ~n29078 ) | ( n2222 & n42086 ) | ( ~n29078 & n42086 ) ;
  assign n49030 = n43835 ^ n4533 ^ n3106 ;
  assign n49031 = n45127 | n49030 ;
  assign n49032 = n1851 | n34109 ;
  assign n49033 = n23722 ^ n431 ^ 1'b0 ;
  assign n49034 = n49033 ^ n22288 ^ n914 ;
  assign n49035 = n49034 ^ n24156 ^ 1'b0 ;
  assign n49036 = ( n6799 & ~n39611 ) | ( n6799 & n49035 ) | ( ~n39611 & n49035 ) ;
  assign n49037 = ~n48564 & n49036 ;
  assign n49038 = n30158 & n49037 ;
  assign n49039 = n49038 ^ n12132 ^ 1'b0 ;
  assign n49040 = n19581 ^ n5497 ^ 1'b0 ;
  assign n49041 = n7050 | n49040 ;
  assign n49042 = n17931 & n20093 ;
  assign n49043 = n22365 & n49042 ;
  assign n49044 = n30309 & n48509 ;
  assign n49045 = n16935 & n19941 ;
  assign n49046 = ~n6891 & n47229 ;
  assign n49047 = n28859 ^ n16225 ^ n6122 ;
  assign n49048 = n31172 ^ n2981 ^ 1'b0 ;
  assign n49049 = ~n12126 & n49048 ;
  assign n49050 = ~n1047 & n2336 ;
  assign n49051 = n29630 & ~n40521 ;
  assign n49052 = n8391 & ~n30877 ;
  assign n49053 = n13503 ^ n2185 ^ 1'b0 ;
  assign n49054 = n34238 & ~n49053 ;
  assign n49055 = n22857 ^ n22834 ^ 1'b0 ;
  assign n49056 = ~n15016 & n49055 ;
  assign n49057 = n49056 ^ n4007 ^ 1'b0 ;
  assign n49058 = ~n1999 & n42512 ;
  assign n49059 = n45965 & n49058 ;
  assign n49060 = n106 & n7031 ;
  assign n49061 = n28687 ^ n8254 ^ 1'b0 ;
  assign n49062 = ~n8243 & n49061 ;
  assign n49063 = ( ~n2080 & n9631 ) | ( ~n2080 & n49062 ) | ( n9631 & n49062 ) ;
  assign n49064 = n49063 ^ n21894 ^ 1'b0 ;
  assign n49065 = n7617 | n49064 ;
  assign n49066 = n20299 | n32191 ;
  assign n49067 = n18941 & ~n26438 ;
  assign n49068 = n12081 ^ n4301 ^ 1'b0 ;
  assign n49069 = ~n49067 & n49068 ;
  assign n49070 = n35199 & ~n35383 ;
  assign n49071 = n14366 & ~n39997 ;
  assign n49072 = ~n3731 & n49071 ;
  assign n49073 = n19831 & n24386 ;
  assign n49074 = n49072 & n49073 ;
  assign n49075 = n21638 & ~n44082 ;
  assign n49076 = n8076 ^ n7649 ^ 1'b0 ;
  assign n49077 = n32848 | n49076 ;
  assign n49078 = n10302 & n15342 ;
  assign n49079 = ~n24035 & n49078 ;
  assign n49080 = n10201 | n15319 ;
  assign n49081 = n4254 | n15618 ;
  assign n49082 = n13007 | n24723 ;
  assign n49083 = n49082 ^ n33399 ^ 1'b0 ;
  assign n49084 = n16675 | n24032 ;
  assign n49085 = ~n56 & n15819 ;
  assign n49086 = n31747 & n49085 ;
  assign n49088 = n46975 ^ n9390 ^ 1'b0 ;
  assign n49087 = n5358 & ~n27925 ;
  assign n49089 = n49088 ^ n49087 ^ 1'b0 ;
  assign n49090 = n12055 | n41724 ;
  assign n49091 = n49090 ^ n8534 ^ 1'b0 ;
  assign n49092 = n17243 ^ n13911 ^ 1'b0 ;
  assign n49093 = n1576 | n10090 ;
  assign n49094 = n235 | n49093 ;
  assign n49095 = n3987 | n28513 ;
  assign n49096 = n19136 ^ n15091 ^ 1'b0 ;
  assign n49097 = n3214 & ~n49096 ;
  assign n49098 = ~n15634 & n17326 ;
  assign n49099 = n49098 ^ n14063 ^ 1'b0 ;
  assign n49100 = n36436 ^ n31642 ^ 1'b0 ;
  assign n49101 = ~n720 & n49100 ;
  assign n49102 = n49101 ^ n37923 ^ 1'b0 ;
  assign n49103 = n49099 & ~n49102 ;
  assign n49104 = n20147 ^ n774 ^ 1'b0 ;
  assign n49105 = n7240 & ~n21054 ;
  assign n49106 = n49104 & n49105 ;
  assign n49107 = n8761 & ~n13939 ;
  assign n49108 = n13848 & ~n29567 ;
  assign n49109 = ~n738 & n49108 ;
  assign n49110 = n30219 & ~n48805 ;
  assign n49112 = n7694 ^ n2492 ^ 1'b0 ;
  assign n49111 = ~n17563 & n18011 ;
  assign n49113 = n49112 ^ n49111 ^ 1'b0 ;
  assign n49114 = n884 & n23035 ;
  assign n49115 = n49114 ^ n19177 ^ 1'b0 ;
  assign n49116 = n42390 | n49115 ;
  assign n49117 = n9063 & ~n24275 ;
  assign n49118 = n49117 ^ n6325 ^ 1'b0 ;
  assign n49119 = n15007 | n37572 ;
  assign n49120 = n14503 & ~n49119 ;
  assign n49123 = n19297 ^ n17065 ^ 1'b0 ;
  assign n49124 = n2519 & ~n49123 ;
  assign n49122 = n17745 ^ n5842 ^ 1'b0 ;
  assign n49125 = n49124 ^ n49122 ^ n5014 ;
  assign n49121 = n4862 | n5916 ;
  assign n49126 = n49125 ^ n49121 ^ 1'b0 ;
  assign n49127 = n9039 & ~n41201 ;
  assign n49128 = ( n6142 & n10364 ) | ( n6142 & n12525 ) | ( n10364 & n12525 ) ;
  assign n49129 = n49128 ^ n445 ^ 1'b0 ;
  assign n49130 = ~n19423 & n49129 ;
  assign n49131 = ~n38908 & n49130 ;
  assign n49132 = ~n11561 & n23167 ;
  assign n49133 = n38997 ^ n14796 ^ 1'b0 ;
  assign n49134 = n14798 & n49133 ;
  assign n49135 = ( n1269 & ~n3649 ) | ( n1269 & n13508 ) | ( ~n3649 & n13508 ) ;
  assign n49136 = n823 | n49135 ;
  assign n49137 = n49136 ^ n37271 ^ 1'b0 ;
  assign n49138 = n1337 & ~n1803 ;
  assign n49139 = n24897 ^ n19356 ^ 1'b0 ;
  assign n49140 = n49138 | n49139 ;
  assign n49141 = ~n2917 & n33867 ;
  assign n49142 = ( n3280 & n35848 ) | ( n3280 & n36145 ) | ( n35848 & n36145 ) ;
  assign n49143 = n13868 | n49142 ;
  assign n49144 = ~n5880 & n12812 ;
  assign n49145 = ( n10822 & n49143 ) | ( n10822 & n49144 ) | ( n49143 & n49144 ) ;
  assign n49146 = ~n48296 & n49145 ;
  assign n49147 = n17411 & ~n19482 ;
  assign n49148 = ~n6730 & n49147 ;
  assign n49149 = n9762 & n21886 ;
  assign n49150 = n24666 ^ n3233 ^ 1'b0 ;
  assign n49151 = ~n40223 & n49150 ;
  assign n49152 = ~n49149 & n49151 ;
  assign n49153 = n1182 & n10855 ;
  assign n49154 = n3333 & ~n49153 ;
  assign n49155 = n2537 & ~n18441 ;
  assign n49156 = ~n2537 & n49155 ;
  assign n49157 = n1591 & n49156 ;
  assign n49158 = ( n8710 & n26532 ) | ( n8710 & n49157 ) | ( n26532 & n49157 ) ;
  assign n49159 = n49158 ^ n40443 ^ 1'b0 ;
  assign n49160 = n28858 & ~n49159 ;
  assign n49161 = n49160 ^ n14981 ^ 1'b0 ;
  assign n49162 = n20346 | n35072 ;
  assign n49163 = n41895 ^ n7893 ^ n7717 ;
  assign n49165 = n47872 ^ n46200 ^ n8858 ;
  assign n49164 = n4919 & ~n31760 ;
  assign n49166 = n49165 ^ n49164 ^ 1'b0 ;
  assign n49167 = n11551 | n33834 ;
  assign n49168 = n8326 | n12915 ;
  assign n49169 = ( ~n18102 & n20250 ) | ( ~n18102 & n28278 ) | ( n20250 & n28278 ) ;
  assign n49170 = n15686 & ~n21618 ;
  assign n49171 = n49170 ^ n23280 ^ n15997 ;
  assign n49172 = ~n3009 & n32483 ;
  assign n49173 = n49172 ^ n8867 ^ 1'b0 ;
  assign n49174 = n451 | n26987 ;
  assign n49175 = n5041 | n8476 ;
  assign n49176 = n11194 & ~n35086 ;
  assign n49178 = n10616 & ~n12262 ;
  assign n49179 = n5165 & n49178 ;
  assign n49177 = n5379 | n11122 ;
  assign n49180 = n49179 ^ n49177 ^ 1'b0 ;
  assign n49181 = n6258 ^ n2208 ^ 1'b0 ;
  assign n49182 = n26214 & ~n49181 ;
  assign n49183 = n2336 | n27203 ;
  assign n49184 = n49183 ^ n1050 ^ 1'b0 ;
  assign n49185 = n13389 ^ n9667 ^ 1'b0 ;
  assign n49186 = n49185 ^ n35346 ^ n13364 ;
  assign n49187 = n5256 & n6166 ;
  assign n49188 = n43238 & ~n49187 ;
  assign n49189 = n36927 ^ n162 ^ 1'b0 ;
  assign n49190 = n11150 | n49189 ;
  assign n49191 = n365 & ~n11255 ;
  assign n49192 = n44676 ^ n14102 ^ n4438 ;
  assign n49193 = n6215 & n49192 ;
  assign n49194 = n49193 ^ n35247 ^ 1'b0 ;
  assign n49195 = n30074 & n40968 ;
  assign n49196 = n32868 | n33932 ;
  assign n49197 = n49196 ^ n12576 ^ 1'b0 ;
  assign n49198 = ~n366 & n12020 ;
  assign n49199 = n49198 ^ n41662 ^ 1'b0 ;
  assign n49200 = n4942 | n49199 ;
  assign n49201 = n6429 | n6641 ;
  assign n49202 = n10785 | n26302 ;
  assign n49203 = n9578 ^ n3660 ^ 1'b0 ;
  assign n49204 = n21675 | n35787 ;
  assign n49205 = n6524 & ~n7570 ;
  assign n49206 = n22572 & ~n49205 ;
  assign n49207 = n49206 ^ n9549 ^ 1'b0 ;
  assign n49208 = n155 & n6489 ;
  assign n49209 = n11043 ^ n10357 ^ n5598 ;
  assign n49210 = n49209 ^ n23932 ^ n21836 ;
  assign n49211 = n38604 ^ n12244 ^ n8279 ;
  assign n49212 = ~n447 & n49211 ;
  assign n49213 = n547 & ~n49212 ;
  assign n49214 = n571 & ~n49213 ;
  assign n49215 = n5108 & ~n27332 ;
  assign n49217 = n5727 ^ n4731 ^ 1'b0 ;
  assign n49216 = n8299 & ~n28137 ;
  assign n49218 = n49217 ^ n49216 ^ 1'b0 ;
  assign n49219 = ~n12025 & n19079 ;
  assign n49220 = n31943 ^ n29784 ^ 1'b0 ;
  assign n49221 = ( n7262 & n10692 ) | ( n7262 & n46206 ) | ( n10692 & n46206 ) ;
  assign n49222 = n9784 ^ n8602 ^ 1'b0 ;
  assign n49223 = n6095 & n40650 ;
  assign n49224 = ~n49222 & n49223 ;
  assign n49225 = n15616 & n28631 ;
  assign n49226 = n7768 & ~n43921 ;
  assign n49227 = n49226 ^ n37123 ^ 1'b0 ;
  assign n49228 = n3357 & n12050 ;
  assign n49229 = n15704 & n49228 ;
  assign n49230 = n9151 & n13850 ;
  assign n49231 = n1119 & ~n8445 ;
  assign n49232 = ~n4359 & n12825 ;
  assign n49233 = ~n49231 & n49232 ;
  assign n49234 = n3012 & ~n12447 ;
  assign n49235 = n49234 ^ n23101 ^ 1'b0 ;
  assign n49236 = n49235 ^ n6180 ^ 1'b0 ;
  assign n49237 = n49186 ^ n8263 ^ 1'b0 ;
  assign n49238 = n44791 & n49237 ;
  assign n49239 = n1925 | n36527 ;
  assign n49240 = ~n44848 & n49239 ;
  assign n49241 = n41543 ^ n23561 ^ 1'b0 ;
  assign n49242 = n3339 & n29918 ;
  assign n49243 = n49242 ^ n21839 ^ 1'b0 ;
  assign n49244 = ~n26803 & n43889 ;
  assign n49245 = n19136 ^ n3126 ^ 1'b0 ;
  assign n49246 = ~n481 & n49245 ;
  assign n49247 = n23292 ^ n3017 ^ 1'b0 ;
  assign n49248 = ~n27113 & n49247 ;
  assign n49249 = ~n6332 & n49248 ;
  assign n49250 = n49249 ^ n25917 ^ 1'b0 ;
  assign n49251 = n36099 & ~n46213 ;
  assign n49252 = n20605 ^ n8728 ^ 1'b0 ;
  assign n49253 = n12028 & n20002 ;
  assign n49254 = n49253 ^ n40118 ^ n16336 ;
  assign n49255 = n30277 & n49254 ;
  assign n49256 = n9208 ^ n2320 ^ n1455 ;
  assign n49257 = n47636 ^ n20621 ^ 1'b0 ;
  assign n49258 = n34527 ^ n7579 ^ 1'b0 ;
  assign n49259 = ( ~n167 & n15477 ) | ( ~n167 & n17265 ) | ( n15477 & n17265 ) ;
  assign n49260 = n49259 ^ n1229 ^ 1'b0 ;
  assign n49261 = n3822 ^ n885 ^ 1'b0 ;
  assign n49262 = n1590 & n49261 ;
  assign n49263 = n49262 ^ n7370 ^ 1'b0 ;
  assign n49264 = n22073 & ~n49263 ;
  assign n49265 = n36197 & ~n49264 ;
  assign n49266 = n49265 ^ n18010 ^ 1'b0 ;
  assign n49267 = n29736 | n49266 ;
  assign n49268 = n33016 ^ n9261 ^ 1'b0 ;
  assign n49269 = n49268 ^ n16670 ^ 1'b0 ;
  assign n49270 = n34668 | n49269 ;
  assign n49271 = n2239 | n49270 ;
  assign n49272 = n19967 & ~n49271 ;
  assign n49273 = n49272 ^ n32157 ^ n14357 ;
  assign n49274 = n45643 ^ n14778 ^ 1'b0 ;
  assign n49275 = ~n22386 & n22942 ;
  assign n49276 = ( n2029 & ~n49274 ) | ( n2029 & n49275 ) | ( ~n49274 & n49275 ) ;
  assign n49277 = n37231 | n43689 ;
  assign n49278 = n16280 & ~n49277 ;
  assign n49279 = n38502 ^ n11827 ^ 1'b0 ;
  assign n49280 = n32322 & n49279 ;
  assign n49284 = n17084 & n44076 ;
  assign n49285 = n33393 & n49284 ;
  assign n49286 = n6631 | n49285 ;
  assign n49287 = n12126 & ~n49286 ;
  assign n49281 = n24620 | n36434 ;
  assign n49282 = n37998 | n49281 ;
  assign n49283 = n48033 & n49282 ;
  assign n49288 = n49287 ^ n49283 ^ 1'b0 ;
  assign n49289 = n6949 ^ n4384 ^ 1'b0 ;
  assign n49290 = n25181 ^ n11546 ^ 1'b0 ;
  assign n49291 = n4932 & n49290 ;
  assign n49292 = n45954 ^ n40017 ^ 1'b0 ;
  assign n49293 = n46021 ^ n12159 ^ n1853 ;
  assign n49294 = ~n3738 & n4347 ;
  assign n49295 = n6174 & n49294 ;
  assign n49296 = n49295 ^ n22566 ^ 1'b0 ;
  assign n49297 = n10711 & ~n31583 ;
  assign n49298 = ~n7148 & n49297 ;
  assign n49299 = n20233 ^ n3940 ^ 1'b0 ;
  assign n49300 = n25598 & n49299 ;
  assign n49301 = n37188 ^ n14897 ^ 1'b0 ;
  assign n49302 = ~n33203 & n35317 ;
  assign n49303 = ~n3064 & n35974 ;
  assign n49304 = ~n225 & n49303 ;
  assign n49305 = n26640 & n49304 ;
  assign n49306 = n24446 ^ n1121 ^ 1'b0 ;
  assign n49307 = n11546 & ~n49306 ;
  assign n49308 = ~n5763 & n16846 ;
  assign n49309 = n8815 & n49308 ;
  assign n49310 = ( n150 & n2343 ) | ( n150 & ~n4439 ) | ( n2343 & ~n4439 ) ;
  assign n49311 = n11100 | n13172 ;
  assign n49312 = ~n12808 & n49311 ;
  assign n49313 = n9124 ^ n144 ^ 1'b0 ;
  assign n49314 = n40813 & ~n49313 ;
  assign n49315 = ~n7156 & n27613 ;
  assign n49316 = ~n19513 & n49315 ;
  assign n49317 = n340 | n20768 ;
  assign n49318 = n35013 & n49317 ;
  assign n49319 = n28772 | n34781 ;
  assign n49320 = n10016 & ~n23375 ;
  assign n49321 = n49320 ^ n21839 ^ 1'b0 ;
  assign n49322 = ~n29297 & n40717 ;
  assign n49323 = n49322 ^ n23258 ^ n6790 ;
  assign n49324 = ~n7724 & n28884 ;
  assign n49325 = n49324 ^ n31457 ^ 1'b0 ;
  assign n49326 = n2812 | n4151 ;
  assign n49327 = n16055 & n49326 ;
  assign n49328 = n49327 ^ n37330 ^ 1'b0 ;
  assign n49329 = n46713 ^ n135 ^ 1'b0 ;
  assign n49330 = n11917 & n49329 ;
  assign n49331 = n8109 & n49330 ;
  assign n49332 = ~n8889 & n49331 ;
  assign n49333 = n2024 & n13190 ;
  assign n49334 = n6489 & n49333 ;
  assign n49335 = n1896 & ~n15926 ;
  assign n49336 = n2604 & n49335 ;
  assign n49337 = n402 & n14227 ;
  assign n49338 = n49337 ^ n18740 ^ 1'b0 ;
  assign n49339 = n1843 & ~n13407 ;
  assign n49340 = ~n1177 & n24088 ;
  assign n49341 = ( n46224 & ~n49339 ) | ( n46224 & n49340 ) | ( ~n49339 & n49340 ) ;
  assign n49343 = n3349 & ~n9190 ;
  assign n49342 = ~n81 & n11000 ;
  assign n49344 = n49343 ^ n49342 ^ 1'b0 ;
  assign n49345 = ~n35204 & n49344 ;
  assign n49346 = n25806 ^ n9369 ^ 1'b0 ;
  assign n49347 = n16190 & ~n49346 ;
  assign n49348 = n19418 ^ n7712 ^ n4091 ;
  assign n49349 = n16587 ^ n7128 ^ 1'b0 ;
  assign n49350 = n49348 & ~n49349 ;
  assign n49351 = n18790 | n39020 ;
  assign n49352 = ~n16888 & n37278 ;
  assign n49353 = n7299 ^ n6645 ^ 1'b0 ;
  assign n49354 = n49352 | n49353 ;
  assign n49355 = n49354 ^ n6893 ^ 1'b0 ;
  assign n49356 = n6092 & n35101 ;
  assign n49357 = n32038 ^ n10670 ^ 1'b0 ;
  assign n49358 = ~n3226 & n49357 ;
  assign n49359 = n44074 & n49358 ;
  assign n49360 = n41474 | n49359 ;
  assign n49361 = n4357 | n43337 ;
  assign n49362 = n47529 ^ n8068 ^ 1'b0 ;
  assign n49363 = n27356 ^ n11034 ^ 1'b0 ;
  assign n49364 = n22654 & ~n49363 ;
  assign n49365 = n3996 & n9191 ;
  assign n49366 = n4554 | n49365 ;
  assign n49367 = n35371 | n49366 ;
  assign n49368 = n21142 ^ n11205 ^ 1'b0 ;
  assign n49369 = n39509 & n49368 ;
  assign n49370 = n19408 & n35597 ;
  assign n49373 = n1853 & ~n5032 ;
  assign n49374 = n7933 & ~n10177 ;
  assign n49375 = ~n29490 & n49374 ;
  assign n49376 = ( n25430 & n49373 ) | ( n25430 & ~n49375 ) | ( n49373 & ~n49375 ) ;
  assign n49371 = n5027 ^ n3197 ^ 1'b0 ;
  assign n49372 = n21 | n49371 ;
  assign n49377 = n49376 ^ n49372 ^ 1'b0 ;
  assign n49378 = n3813 | n7460 ;
  assign n49379 = n49377 | n49378 ;
  assign n49380 = n36278 ^ n32974 ^ n17701 ;
  assign n49381 = n49380 ^ n35749 ^ n428 ;
  assign n49382 = n19595 ^ n17103 ^ 1'b0 ;
  assign n49383 = n36455 | n49382 ;
  assign n49384 = n36862 ^ n304 ^ 1'b0 ;
  assign n49385 = n6296 & ~n49384 ;
  assign n49386 = n49385 ^ n40534 ^ 1'b0 ;
  assign n49387 = n1002 & n49386 ;
  assign n49388 = n7889 | n45621 ;
  assign n49389 = n14155 & ~n49388 ;
  assign n49390 = n49389 ^ n19949 ^ 1'b0 ;
  assign n49391 = ~n1083 & n13615 ;
  assign n49392 = n49391 ^ n10897 ^ 1'b0 ;
  assign n49393 = n14237 & ~n49392 ;
  assign n49394 = ~n49390 & n49393 ;
  assign n49395 = n17627 ^ n1473 ^ 1'b0 ;
  assign n49396 = n12970 | n49395 ;
  assign n49398 = ~n3477 & n15042 ;
  assign n49399 = n47470 & n49398 ;
  assign n49397 = n6749 ^ n5209 ^ 1'b0 ;
  assign n49400 = n49399 ^ n49397 ^ n8365 ;
  assign n49401 = n49400 ^ n6764 ^ 1'b0 ;
  assign n49403 = n4349 | n8594 ;
  assign n49402 = n4634 & ~n6666 ;
  assign n49404 = n49403 ^ n49402 ^ 1'b0 ;
  assign n49405 = n20902 & ~n49404 ;
  assign n49406 = ~n15018 & n49405 ;
  assign n49407 = n49406 ^ n13557 ^ 1'b0 ;
  assign n49408 = n35409 | n44625 ;
  assign n49409 = ( ~n942 & n6479 ) | ( ~n942 & n46441 ) | ( n6479 & n46441 ) ;
  assign n49410 = n609 | n48377 ;
  assign n49411 = n37625 | n49410 ;
  assign n49412 = n49411 ^ n30989 ^ n6176 ;
  assign n49413 = n25233 ^ n3992 ^ 1'b0 ;
  assign n49414 = n2222 & ~n49413 ;
  assign n49415 = n9365 | n29546 ;
  assign n49416 = ~n9322 & n31325 ;
  assign n49417 = n328 & n21091 ;
  assign n49418 = n15367 ^ n152 ^ 1'b0 ;
  assign n49419 = n25436 ^ n18927 ^ 1'b0 ;
  assign n49420 = n45 | n24727 ;
  assign n49421 = n12760 | n49420 ;
  assign n49422 = n25334 & ~n30013 ;
  assign n49423 = n49422 ^ n32154 ^ 1'b0 ;
  assign n49424 = n21679 ^ n8133 ^ 1'b0 ;
  assign n49425 = n10143 | n49424 ;
  assign n49426 = n49425 ^ n5332 ^ n1157 ;
  assign n49427 = n33568 | n38281 ;
  assign n49428 = n29368 ^ n15413 ^ 1'b0 ;
  assign n49429 = ~n5976 & n49428 ;
  assign n49430 = n28072 | n41835 ;
  assign n49431 = n49429 | n49430 ;
  assign n49432 = n26808 ^ n10792 ^ 1'b0 ;
  assign n49433 = n31993 & ~n49432 ;
  assign n49434 = n11733 | n44626 ;
  assign n49435 = n15888 | n49434 ;
  assign n49436 = n6281 | n49435 ;
  assign n49437 = n49436 ^ n40779 ^ 1'b0 ;
  assign n49438 = n18723 & n49437 ;
  assign n49439 = ~n13567 & n20799 ;
  assign n49440 = n12700 ^ n8552 ^ 1'b0 ;
  assign n49441 = n49439 & ~n49440 ;
  assign n49442 = n49441 ^ n29587 ^ n1263 ;
  assign n49443 = n4014 & n49442 ;
  assign n49444 = n24089 & ~n28448 ;
  assign n49445 = n1481 & ~n18832 ;
  assign n49446 = ~n29652 & n49445 ;
  assign n49447 = n29368 | n49446 ;
  assign n49448 = n21591 ^ n4409 ^ 1'b0 ;
  assign n49449 = n49448 ^ n19105 ^ 1'b0 ;
  assign n49450 = ~n12751 & n49449 ;
  assign n49451 = n4808 | n29677 ;
  assign n49452 = n3068 & ~n16285 ;
  assign n49453 = n49452 ^ n13173 ^ 1'b0 ;
  assign n49454 = ~n1367 & n27464 ;
  assign n49455 = n8281 & ~n22326 ;
  assign n49456 = ~n30069 & n49455 ;
  assign n49457 = n24673 & n49456 ;
  assign n49458 = n20577 ^ n5121 ^ 1'b0 ;
  assign n49459 = n2346 & n4170 ;
  assign n49460 = ~n49458 & n49459 ;
  assign n49461 = n10267 & n49460 ;
  assign n49462 = ~n1570 & n49461 ;
  assign n49463 = n49457 & n49462 ;
  assign n49464 = n38034 ^ n6714 ^ 1'b0 ;
  assign n49465 = n4604 | n24829 ;
  assign n49466 = n5396 & n47261 ;
  assign n49467 = n49466 ^ n14235 ^ 1'b0 ;
  assign n49468 = n17480 ^ n13640 ^ 1'b0 ;
  assign n49471 = ~n5116 & n15616 ;
  assign n49469 = n41544 ^ n13190 ^ 1'b0 ;
  assign n49470 = n49469 ^ n8430 ^ n7927 ;
  assign n49472 = n49471 ^ n49470 ^ 1'b0 ;
  assign n49473 = n19062 & n29028 ;
  assign n49474 = ~n18565 & n49473 ;
  assign n49475 = n216 & ~n38736 ;
  assign n49476 = n49474 | n49475 ;
  assign n49477 = n36406 ^ n25708 ^ 1'b0 ;
  assign n49478 = ~n49476 & n49477 ;
  assign n49479 = n14007 ^ n2381 ^ 1'b0 ;
  assign n49480 = n24023 | n49479 ;
  assign n49481 = n18429 & ~n36503 ;
  assign n49482 = n49481 ^ n42016 ^ 1'b0 ;
  assign n49483 = n3720 | n19795 ;
  assign n49484 = n49483 ^ n25316 ^ 1'b0 ;
  assign n49485 = n22854 | n47688 ;
  assign n49486 = n31118 ^ n8457 ^ 1'b0 ;
  assign n49487 = n17283 & ~n49486 ;
  assign n49488 = n38158 ^ n7462 ^ 1'b0 ;
  assign n49489 = ( ~n30811 & n49487 ) | ( ~n30811 & n49488 ) | ( n49487 & n49488 ) ;
  assign n49490 = n2118 | n3331 ;
  assign n49491 = n49490 ^ n30993 ^ 1'b0 ;
  assign n49492 = n19912 & ~n49491 ;
  assign n49493 = n22990 ^ n6181 ^ 1'b0 ;
  assign n49494 = ~n10486 & n49493 ;
  assign n49495 = n30249 ^ n28954 ^ n16275 ;
  assign n49496 = n7913 | n49495 ;
  assign n49497 = ~n3314 & n21049 ;
  assign n49498 = ~n5767 & n49497 ;
  assign n49499 = n822 & n27880 ;
  assign n49500 = n17866 & ~n49499 ;
  assign n49501 = n49500 ^ n6748 ^ 1'b0 ;
  assign n49502 = ~n49498 & n49501 ;
  assign n49503 = ~n20669 & n49502 ;
  assign n49504 = n19551 ^ n2519 ^ 1'b0 ;
  assign n49505 = n16885 & ~n49504 ;
  assign n49506 = n35432 ^ n4263 ^ 1'b0 ;
  assign n49507 = ( n302 & ~n13163 ) | ( n302 & n48864 ) | ( ~n13163 & n48864 ) ;
  assign n49508 = n8578 & ~n28894 ;
  assign n49509 = n33010 ^ n48 ^ 1'b0 ;
  assign n49510 = n49508 & ~n49509 ;
  assign n49511 = n10298 ^ n4751 ^ 1'b0 ;
  assign n49512 = ~n45023 & n49511 ;
  assign n49513 = n49512 ^ n41487 ^ n11374 ;
  assign n49514 = n42331 ^ n18783 ^ 1'b0 ;
  assign n49515 = n1403 & ~n49514 ;
  assign n49517 = ~n16507 & n34432 ;
  assign n49516 = ~n27207 & n32791 ;
  assign n49518 = n49517 ^ n49516 ^ 1'b0 ;
  assign n49519 = n3601 & n6526 ;
  assign n49520 = ~n16308 & n49519 ;
  assign n49521 = n17420 & ~n49520 ;
  assign n49522 = n22467 | n27758 ;
  assign n49523 = n42833 | n49522 ;
  assign n49524 = ~n1422 & n49523 ;
  assign n49525 = n4015 | n49524 ;
  assign n49526 = n48894 ^ n6640 ^ n1434 ;
  assign n49527 = n3639 & ~n11208 ;
  assign n49528 = ~n3639 & n49527 ;
  assign n49529 = n1141 | n49528 ;
  assign n49530 = n49529 ^ n26048 ^ 1'b0 ;
  assign n49531 = n1254 & ~n49530 ;
  assign n49532 = n17689 & n49531 ;
  assign n49533 = n29096 & n32787 ;
  assign n49534 = n49533 ^ n514 ^ 1'b0 ;
  assign n49535 = n34422 ^ n4976 ^ 1'b0 ;
  assign n49536 = n9288 | n49017 ;
  assign n49537 = n11536 ^ n10935 ^ n7254 ;
  assign n49538 = n30894 & ~n49537 ;
  assign n49543 = ~n1574 & n5262 ;
  assign n49544 = n11252 & n49543 ;
  assign n49542 = n4182 & n47546 ;
  assign n49545 = n49544 ^ n49542 ^ 1'b0 ;
  assign n49539 = n28561 ^ n4990 ^ 1'b0 ;
  assign n49540 = n1360 & n49539 ;
  assign n49541 = n3758 & n49540 ;
  assign n49546 = n49545 ^ n49541 ^ n31867 ;
  assign n49547 = n23600 ^ n12996 ^ 1'b0 ;
  assign n49548 = ~n31 & n5346 ;
  assign n49549 = n1808 | n13809 ;
  assign n49550 = n49549 ^ n8454 ^ 1'b0 ;
  assign n49551 = n49548 | n49550 ;
  assign n49552 = n22580 & ~n30031 ;
  assign n49553 = n49552 ^ n39614 ^ 1'b0 ;
  assign n49554 = n12544 & ~n31818 ;
  assign n49555 = n18177 ^ n11550 ^ 1'b0 ;
  assign n49556 = ~n23393 & n49555 ;
  assign n49557 = n49556 ^ n8181 ^ 1'b0 ;
  assign n49558 = n28199 ^ n3218 ^ 1'b0 ;
  assign n49559 = n48042 ^ n29950 ^ 1'b0 ;
  assign n49560 = n8453 & n12740 ;
  assign n49561 = ~n44581 & n47530 ;
  assign n49562 = n26116 ^ n12195 ^ 1'b0 ;
  assign n49563 = ~n10860 & n49562 ;
  assign n49564 = n38498 ^ n13456 ^ 1'b0 ;
  assign n49565 = n15792 & ~n27943 ;
  assign n49566 = n45226 ^ n17005 ^ 1'b0 ;
  assign n49567 = n7031 | n20819 ;
  assign n49568 = n49567 ^ n11899 ^ 1'b0 ;
  assign n49569 = n49566 & n49568 ;
  assign n49570 = n1570 & ~n2803 ;
  assign n49571 = ~n48278 & n49570 ;
  assign n49572 = n20864 | n49571 ;
  assign n49573 = n27871 & ~n49572 ;
  assign n49574 = n28294 & ~n49573 ;
  assign n49575 = ~n16313 & n49574 ;
  assign n49576 = n26104 | n49575 ;
  assign n49577 = n43921 & ~n49576 ;
  assign n49578 = n4976 | n44888 ;
  assign n49579 = n8643 & ~n49578 ;
  assign n49580 = n25953 ^ n17979 ^ 1'b0 ;
  assign n49581 = n9798 | n24263 ;
  assign n49582 = n49581 ^ n24727 ^ 1'b0 ;
  assign n49583 = ~n6040 & n14946 ;
  assign n49584 = n49583 ^ n28637 ^ 1'b0 ;
  assign n49585 = n257 | n17775 ;
  assign n49586 = n16239 & n20831 ;
  assign n49587 = n49586 ^ n5857 ^ 1'b0 ;
  assign n49588 = n16926 ^ n4425 ^ 1'b0 ;
  assign n49589 = n49587 | n49588 ;
  assign n49590 = n5270 & n31971 ;
  assign n49591 = n49590 ^ n48315 ^ 1'b0 ;
  assign n49592 = n4553 & ~n27463 ;
  assign n49593 = ~n47344 & n49592 ;
  assign n49594 = ~n24263 & n49593 ;
  assign n49595 = n26235 ^ n9494 ^ 1'b0 ;
  assign n49596 = n1385 | n16721 ;
  assign n49597 = n49596 ^ n5400 ^ 1'b0 ;
  assign n49598 = n49597 ^ n7010 ^ 1'b0 ;
  assign n49599 = n19642 & n49598 ;
  assign n49600 = n44939 ^ n5194 ^ 1'b0 ;
  assign n49601 = n37395 | n49600 ;
  assign n49602 = n47917 ^ n12150 ^ 1'b0 ;
  assign n49603 = ( n3408 & n8449 ) | ( n3408 & n40785 ) | ( n8449 & n40785 ) ;
  assign n49604 = n13544 ^ n9636 ^ 1'b0 ;
  assign n49605 = n11954 ^ n4408 ^ 1'b0 ;
  assign n49606 = n7082 ^ n52 ^ 1'b0 ;
  assign n49607 = n17566 & ~n49606 ;
  assign n49612 = n6250 & ~n19159 ;
  assign n49608 = n181 & n4002 ;
  assign n49609 = n49608 ^ n7125 ^ 1'b0 ;
  assign n49610 = n1845 | n49609 ;
  assign n49611 = n11312 & ~n49610 ;
  assign n49613 = n49612 ^ n49611 ^ 1'b0 ;
  assign n49614 = ~n13059 & n19300 ;
  assign n49615 = ~n9051 & n22948 ;
  assign n49616 = n5387 ^ n991 ^ 1'b0 ;
  assign n49617 = ( n7833 & n48586 ) | ( n7833 & n49616 ) | ( n48586 & n49616 ) ;
  assign n49618 = ~n18374 & n28490 ;
  assign n49619 = n5872 & n7897 ;
  assign n49620 = n32113 & ~n49619 ;
  assign n49621 = n49620 ^ n16295 ^ 1'b0 ;
  assign n49622 = n35186 ^ n2838 ^ 1'b0 ;
  assign n49623 = n904 & n49622 ;
  assign n49624 = n49623 ^ n1700 ^ 1'b0 ;
  assign n49625 = n49621 & ~n49624 ;
  assign n49626 = ( n16600 & n49618 ) | ( n16600 & n49625 ) | ( n49618 & n49625 ) ;
  assign n49627 = n2658 & n34959 ;
  assign n49628 = n165 & ~n21029 ;
  assign n49629 = n49628 ^ n31225 ^ n11927 ;
  assign n49630 = n49629 ^ n21990 ^ 1'b0 ;
  assign n49631 = n14382 & n49630 ;
  assign n49632 = ~n41726 & n49631 ;
  assign n49633 = n43005 ^ n12678 ^ 1'b0 ;
  assign n49634 = n22099 & n44509 ;
  assign n49635 = n1413 & n49634 ;
  assign n49636 = n6545 & n22380 ;
  assign n49637 = n19100 ^ n15684 ^ 1'b0 ;
  assign n49638 = n24096 & n49637 ;
  assign n49639 = ( n2046 & n2390 ) | ( n2046 & ~n31457 ) | ( n2390 & ~n31457 ) ;
  assign n49640 = n34598 ^ n3113 ^ 1'b0 ;
  assign n49641 = n40401 | n49640 ;
  assign n49642 = n8879 & n36940 ;
  assign n49643 = n11345 ^ n3574 ^ 1'b0 ;
  assign n49644 = n6615 | n49643 ;
  assign n49645 = n48950 | n49644 ;
  assign n49646 = n12215 & ~n36573 ;
  assign n49647 = n19888 & ~n49646 ;
  assign n49648 = n27169 ^ n11291 ^ 1'b0 ;
  assign n49649 = n29240 ^ n4712 ^ 1'b0 ;
  assign n49650 = n43080 ^ n1038 ^ 1'b0 ;
  assign n49651 = n2324 & n49650 ;
  assign n49652 = n49651 ^ n41246 ^ n6380 ;
  assign n49653 = n1242 ^ n317 ^ 1'b0 ;
  assign n49654 = n28884 & n40941 ;
  assign n49655 = n49654 ^ n11291 ^ 1'b0 ;
  assign n49656 = ~n5885 & n49655 ;
  assign n49657 = n2361 | n44065 ;
  assign n49658 = n49657 ^ n28344 ^ 1'b0 ;
  assign n49659 = n49658 ^ n4586 ^ 1'b0 ;
  assign n49660 = n1905 & ~n49659 ;
  assign n49661 = n5106 & n47529 ;
  assign n49662 = n49661 ^ n19912 ^ 1'b0 ;
  assign n49663 = n8500 | n36218 ;
  assign n49664 = n27661 | n49663 ;
  assign n49665 = ~n6345 & n16853 ;
  assign n49666 = n4675 & ~n21597 ;
  assign n49667 = n47805 ^ n28306 ^ 1'b0 ;
  assign n49668 = ( ~n30205 & n33601 ) | ( ~n30205 & n49667 ) | ( n33601 & n49667 ) ;
  assign n49669 = n20145 & ~n26120 ;
  assign n49670 = n2133 & ~n22793 ;
  assign n49671 = n33 & n49670 ;
  assign n49672 = n9639 & n34673 ;
  assign n49673 = ~n11118 & n26288 ;
  assign n49674 = n13541 ^ n4924 ^ 1'b0 ;
  assign n49675 = n2202 ^ n637 ^ 1'b0 ;
  assign n49676 = n39608 ^ n14927 ^ 1'b0 ;
  assign n49677 = n49675 & n49676 ;
  assign n49678 = n23183 ^ n920 ^ 1'b0 ;
  assign n49679 = ~n9795 & n49678 ;
  assign n49680 = n1539 | n30476 ;
  assign n49681 = n15686 ^ n10552 ^ 1'b0 ;
  assign n49682 = n17558 & ~n49681 ;
  assign n49683 = n27907 ^ n19766 ^ 1'b0 ;
  assign n49684 = n25402 | n25651 ;
  assign n49685 = n17433 | n49684 ;
  assign n49686 = n49685 ^ n28493 ^ 1'b0 ;
  assign n49687 = n7582 & ~n48217 ;
  assign n49688 = n1157 & n31415 ;
  assign n49689 = n21488 & n30328 ;
  assign n49690 = n49689 ^ n20544 ^ 1'b0 ;
  assign n49691 = n6846 | n13920 ;
  assign n49692 = n49691 ^ n16398 ^ 1'b0 ;
  assign n49693 = n16433 ^ n3235 ^ 1'b0 ;
  assign n49694 = n11747 & ~n12654 ;
  assign n49695 = n49694 ^ n28623 ^ 1'b0 ;
  assign n49696 = n11187 & ~n49695 ;
  assign n49697 = ~n3442 & n27703 ;
  assign n49698 = ( n9047 & n42255 ) | ( n9047 & n49697 ) | ( n42255 & n49697 ) ;
  assign n49699 = n14149 ^ n5048 ^ 1'b0 ;
  assign n49700 = n7823 | n49699 ;
  assign n49701 = n49700 ^ n9770 ^ 1'b0 ;
  assign n49702 = n44266 | n47584 ;
  assign n49703 = ( n9609 & ~n16197 ) | ( n9609 & n26301 ) | ( ~n16197 & n26301 ) ;
  assign n49704 = n49703 ^ n10795 ^ 1'b0 ;
  assign n49705 = n6754 ^ n3760 ^ 1'b0 ;
  assign n49706 = n49704 & n49705 ;
  assign n49707 = n13695 & n35925 ;
  assign n49708 = ~n7531 & n49707 ;
  assign n49709 = n8217 | n30949 ;
  assign n49710 = n10632 | n23020 ;
  assign n49711 = n49710 ^ n18648 ^ 1'b0 ;
  assign n49717 = n11257 | n36385 ;
  assign n49718 = n7075 & ~n49717 ;
  assign n49719 = n33017 & ~n49718 ;
  assign n49714 = n3909 & ~n4870 ;
  assign n49715 = n49714 ^ n21391 ^ 1'b0 ;
  assign n49713 = x6 & n26021 ;
  assign n49716 = n49715 ^ n49713 ^ 1'b0 ;
  assign n49712 = ~n33049 & n40731 ;
  assign n49720 = n49719 ^ n49716 ^ n49712 ;
  assign n49721 = n12022 | n29635 ;
  assign n49722 = ( n3665 & n6375 ) | ( n3665 & ~n25296 ) | ( n6375 & ~n25296 ) ;
  assign n49723 = n8595 & ~n9650 ;
  assign n49724 = ~n49722 & n49723 ;
  assign n49725 = n49724 ^ n21505 ^ 1'b0 ;
  assign n49726 = ~n12731 & n49725 ;
  assign n49727 = n49726 ^ n11768 ^ 1'b0 ;
  assign n49728 = ~n3542 & n21208 ;
  assign n49729 = n49728 ^ n39538 ^ 1'b0 ;
  assign n49730 = n20283 | n38627 ;
  assign n49731 = ( n12224 & ~n30543 ) | ( n12224 & n42793 ) | ( ~n30543 & n42793 ) ;
  assign n49732 = n13771 & n32205 ;
  assign n49733 = n3779 | n49732 ;
  assign n49734 = n49733 ^ n3489 ^ 1'b0 ;
  assign n49735 = ~n49731 & n49734 ;
  assign n49736 = n8660 & ~n30440 ;
  assign n49737 = n8612 | n23822 ;
  assign n49738 = n4344 & ~n49737 ;
  assign n49739 = n49738 ^ n22599 ^ n1568 ;
  assign n49740 = n7423 & n28389 ;
  assign n49741 = n12160 & n49740 ;
  assign n49742 = n7182 & ~n49741 ;
  assign n49743 = n7913 ^ n6421 ^ 1'b0 ;
  assign n49744 = n290 & n19830 ;
  assign n49745 = ~n6930 & n49744 ;
  assign n49746 = n49743 & n49745 ;
  assign n49747 = n8310 ^ n2137 ^ 1'b0 ;
  assign n49748 = n23541 & ~n27976 ;
  assign n49749 = n1701 & n16053 ;
  assign n49750 = n49749 ^ n831 ^ 1'b0 ;
  assign n49753 = n4420 ^ n1741 ^ 1'b0 ;
  assign n49754 = n6262 | n49753 ;
  assign n49755 = n3586 & n49754 ;
  assign n49751 = n11738 & ~n32185 ;
  assign n49752 = n49751 ^ n4997 ^ 1'b0 ;
  assign n49756 = n49755 ^ n49752 ^ 1'b0 ;
  assign n49757 = n31080 & ~n49756 ;
  assign n49758 = n6033 | n13108 ;
  assign n49759 = ~n20189 & n35674 ;
  assign n49760 = ( n1367 & n34163 ) | ( n1367 & n49759 ) | ( n34163 & n49759 ) ;
  assign n49761 = n25407 & n34732 ;
  assign n49762 = ~n17542 & n49761 ;
  assign n49763 = n49762 ^ n29233 ^ 1'b0 ;
  assign n49764 = n1371 & n21023 ;
  assign n49765 = n49764 ^ n2519 ^ 1'b0 ;
  assign n49766 = n37047 | n40238 ;
  assign n49767 = n12763 | n49766 ;
  assign n49768 = ~n9776 & n33013 ;
  assign n49769 = n49768 ^ n24770 ^ 1'b0 ;
  assign n49770 = n28038 ^ n13308 ^ n3218 ;
  assign n49771 = ( ~n1800 & n2140 ) | ( ~n1800 & n36636 ) | ( n2140 & n36636 ) ;
  assign n49772 = ( n26123 & ~n49770 ) | ( n26123 & n49771 ) | ( ~n49770 & n49771 ) ;
  assign n49773 = n10937 ^ n2029 ^ 1'b0 ;
  assign n49774 = n7486 | n49773 ;
  assign n49775 = ~n15926 & n49774 ;
  assign n49776 = n15539 | n33753 ;
  assign n49777 = n49775 | n49776 ;
  assign n49778 = n1081 & ~n3693 ;
  assign n49779 = n49778 ^ n10421 ^ n1993 ;
  assign n49780 = n749 | n21174 ;
  assign n49781 = n3195 & n10257 ;
  assign n49782 = n30393 | n49781 ;
  assign n49783 = n49782 ^ n11039 ^ 1'b0 ;
  assign n49784 = n45553 ^ n44584 ^ n18441 ;
  assign n49785 = n2989 & n41684 ;
  assign n49786 = n11945 ^ n302 ^ 1'b0 ;
  assign n49787 = n8965 & ~n49786 ;
  assign n49788 = n44994 & ~n49787 ;
  assign n49789 = n49788 ^ n10070 ^ 1'b0 ;
  assign n49790 = n36754 | n49789 ;
  assign n49791 = n49790 ^ n9707 ^ 1'b0 ;
  assign n49792 = n39582 & n49791 ;
  assign n49793 = n20992 ^ n17410 ^ 1'b0 ;
  assign n49794 = ~n21145 & n33468 ;
  assign n49795 = n48791 ^ n7405 ^ 1'b0 ;
  assign n49796 = n30809 | n49795 ;
  assign n49797 = n39607 ^ n38104 ^ 1'b0 ;
  assign n49798 = ( ~n695 & n2566 ) | ( ~n695 & n49797 ) | ( n2566 & n49797 ) ;
  assign n49799 = n9763 ^ n8655 ^ n6091 ;
  assign n49800 = n23324 & n31171 ;
  assign n49801 = ~n49799 & n49800 ;
  assign n49802 = n7637 | n49801 ;
  assign n49803 = ( n365 & ~n19876 ) | ( n365 & n49802 ) | ( ~n19876 & n49802 ) ;
  assign n49804 = n1645 | n48925 ;
  assign n49805 = n15716 ^ n4946 ^ 1'b0 ;
  assign n49806 = n21650 & ~n49805 ;
  assign n49807 = n17797 & n37537 ;
  assign n49808 = n49807 ^ n10595 ^ 1'b0 ;
  assign n49809 = n498 & ~n33391 ;
  assign n49810 = n36687 & n49809 ;
  assign n49811 = n3435 ^ n2492 ^ 1'b0 ;
  assign n49812 = n43474 | n49811 ;
  assign n49813 = n49812 ^ n8135 ^ 1'b0 ;
  assign n49814 = n25817 & ~n49813 ;
  assign n49815 = n1525 & n1545 ;
  assign n49816 = n32375 & n49815 ;
  assign n49817 = n4303 & n11515 ;
  assign n49818 = n31925 & n49817 ;
  assign n49819 = n2368 & ~n4279 ;
  assign n49820 = n27724 ^ n17253 ^ 1'b0 ;
  assign n49821 = n28695 ^ n19116 ^ 1'b0 ;
  assign n49822 = ( n49819 & n49820 ) | ( n49819 & ~n49821 ) | ( n49820 & ~n49821 ) ;
  assign n49823 = n9781 & ~n20012 ;
  assign n49825 = n18416 ^ n2533 ^ 1'b0 ;
  assign n49826 = n21092 & n49825 ;
  assign n49824 = n6198 & n9588 ;
  assign n49827 = n49826 ^ n49824 ^ 1'b0 ;
  assign n49829 = n860 | n13383 ;
  assign n49830 = n21587 & ~n49829 ;
  assign n49828 = n16247 ^ n10500 ^ 1'b0 ;
  assign n49831 = n49830 ^ n49828 ^ 1'b0 ;
  assign n49832 = n23780 | n49831 ;
  assign n49833 = ~n27955 & n49832 ;
  assign n49834 = n9364 | n42665 ;
  assign n49835 = n49833 & ~n49834 ;
  assign n49836 = n9792 | n19186 ;
  assign n49837 = n49836 ^ n4311 ^ 1'b0 ;
  assign n49838 = ~n16736 & n49837 ;
  assign n49839 = n48824 ^ n4008 ^ 1'b0 ;
  assign n49840 = ~n16190 & n49839 ;
  assign n49842 = n2408 & ~n17226 ;
  assign n49841 = ~n11868 & n24255 ;
  assign n49843 = n49842 ^ n49841 ^ 1'b0 ;
  assign n49844 = n9682 & ~n27888 ;
  assign n49845 = ~n7071 & n28121 ;
  assign n49846 = n767 & n49845 ;
  assign n49847 = n1031 & n23351 ;
  assign n49848 = n49847 ^ n4357 ^ 1'b0 ;
  assign n49849 = n8560 & ~n21315 ;
  assign n49850 = n18597 | n19302 ;
  assign n49851 = n18511 | n49850 ;
  assign n49852 = n39020 ^ n24559 ^ 1'b0 ;
  assign n49853 = n49851 & n49852 ;
  assign n49855 = n29912 ^ n19195 ^ 1'b0 ;
  assign n49856 = n45042 & ~n49855 ;
  assign n49857 = n3003 & n38766 ;
  assign n49858 = ~n49856 & n49857 ;
  assign n49854 = ~n10092 & n11177 ;
  assign n49859 = n49858 ^ n49854 ^ 1'b0 ;
  assign n49860 = n4113 | n38419 ;
  assign n49861 = n44996 | n49860 ;
  assign n49862 = ~n31 & n4677 ;
  assign n49863 = n49862 ^ n29544 ^ 1'b0 ;
  assign n49864 = n10717 | n26208 ;
  assign n49865 = n1093 & ~n49864 ;
  assign n49866 = ~n17659 & n49865 ;
  assign n49867 = ~n10711 & n40076 ;
  assign n49868 = ~n28557 & n49867 ;
  assign n49869 = n49868 ^ n37169 ^ 1'b0 ;
  assign n49870 = ( n11852 & ~n27251 ) | ( n11852 & n38965 ) | ( ~n27251 & n38965 ) ;
  assign n49871 = n8870 ^ n1251 ^ 1'b0 ;
  assign n49872 = n9643 & ~n11786 ;
  assign n49873 = n16002 ^ n15103 ^ 1'b0 ;
  assign n49874 = ~n2856 & n49873 ;
  assign n49875 = n14580 | n39873 ;
  assign n49876 = n49875 ^ n9753 ^ 1'b0 ;
  assign n49877 = n33670 ^ n11460 ^ 1'b0 ;
  assign n49878 = n26708 & ~n41334 ;
  assign n49879 = n22654 & n34786 ;
  assign n49880 = n49879 ^ n8595 ^ 1'b0 ;
  assign n49881 = n22607 & ~n24262 ;
  assign n49882 = n16252 & ~n20580 ;
  assign n49883 = ~n4059 & n49882 ;
  assign n49884 = n42883 ^ n8338 ^ 1'b0 ;
  assign n49885 = n30841 ^ n27624 ^ n25553 ;
  assign n49886 = n2155 | n18159 ;
  assign n49887 = n49886 ^ n21402 ^ 1'b0 ;
  assign n49888 = n3818 & ~n49887 ;
  assign n49889 = n38144 & n39176 ;
  assign n49890 = ~n24991 & n49889 ;
  assign n49891 = n7316 ^ n2664 ^ 1'b0 ;
  assign n49892 = n49891 ^ n18041 ^ n5877 ;
  assign n49893 = n3473 & ~n24324 ;
  assign n49894 = n509 | n42569 ;
  assign n49903 = n38772 ^ n19892 ^ 1'b0 ;
  assign n49900 = n31758 ^ n1664 ^ 1'b0 ;
  assign n49901 = n17326 & ~n49900 ;
  assign n49895 = n758 & ~n15623 ;
  assign n49896 = n49895 ^ n11238 ^ 1'b0 ;
  assign n49897 = n26882 & ~n49896 ;
  assign n49898 = n21784 & n49897 ;
  assign n49899 = n37144 & ~n49898 ;
  assign n49902 = n49901 ^ n49899 ^ 1'b0 ;
  assign n49904 = n49903 ^ n49902 ^ n18342 ;
  assign n49905 = n9470 | n33370 ;
  assign n49906 = n49905 ^ n23580 ^ 1'b0 ;
  assign n49907 = ~n1732 & n7924 ;
  assign n49908 = ~n17642 & n49907 ;
  assign n49909 = n11731 & n25454 ;
  assign n49910 = n24059 & n49909 ;
  assign n49911 = n28941 | n33906 ;
  assign n49912 = n15934 | n21052 ;
  assign n49913 = n15851 ^ n2537 ^ 1'b0 ;
  assign n49914 = ( ~n11947 & n49912 ) | ( ~n11947 & n49913 ) | ( n49912 & n49913 ) ;
  assign n49915 = n7755 & n49914 ;
  assign n49916 = n13109 & n34360 ;
  assign n49917 = ~n5305 & n29757 ;
  assign n49918 = n49917 ^ n1395 ^ 1'b0 ;
  assign n49919 = n49918 ^ n18890 ^ 1'b0 ;
  assign n49920 = ~n49916 & n49919 ;
  assign n49921 = ( ~n8494 & n14739 ) | ( ~n8494 & n17350 ) | ( n14739 & n17350 ) ;
  assign n49922 = n49921 ^ n3777 ^ 1'b0 ;
  assign n49923 = n15528 ^ n880 ^ 1'b0 ;
  assign n49924 = n2046 | n49923 ;
  assign n49925 = n49924 ^ n44202 ^ n20506 ;
  assign n49926 = ( n5032 & n43943 ) | ( n5032 & n49925 ) | ( n43943 & n49925 ) ;
  assign n49927 = n16712 & ~n44882 ;
  assign n49928 = n49927 ^ n29655 ^ 1'b0 ;
  assign n49929 = n34710 ^ n26405 ^ n2136 ;
  assign n49930 = n1981 & ~n7521 ;
  assign n49931 = n19946 ^ n3665 ^ 1'b0 ;
  assign n49932 = n49930 & n49931 ;
  assign n49933 = ~n16280 & n49932 ;
  assign n49934 = n31240 & n49933 ;
  assign n49935 = n32715 ^ n26276 ^ 1'b0 ;
  assign n49936 = n15792 | n32364 ;
  assign n49937 = n11524 | n49936 ;
  assign n49938 = n41278 ^ n19438 ^ n5866 ;
  assign n49939 = n170 & n15877 ;
  assign n49940 = n16828 & ~n36528 ;
  assign n49941 = n49940 ^ n35 ^ 1'b0 ;
  assign n49942 = n1838 & ~n49941 ;
  assign n49943 = n34688 ^ n20445 ^ 1'b0 ;
  assign n49944 = n9193 & n49943 ;
  assign n49945 = ( n1047 & n22610 ) | ( n1047 & n38870 ) | ( n22610 & n38870 ) ;
  assign n49946 = ~n1960 & n49945 ;
  assign n49947 = n6474 | n14629 ;
  assign n49948 = ~n1238 & n7319 ;
  assign n49949 = n1238 & n49948 ;
  assign n49950 = n351 & n49949 ;
  assign n49951 = n49950 ^ n42668 ^ 1'b0 ;
  assign n49952 = ( n12163 & n49947 ) | ( n12163 & ~n49951 ) | ( n49947 & ~n49951 ) ;
  assign n49953 = n49952 ^ n45313 ^ 1'b0 ;
  assign n49954 = n23067 & n49953 ;
  assign n49955 = n34349 ^ n13437 ^ 1'b0 ;
  assign n49956 = n21926 & ~n49955 ;
  assign n49957 = n46398 & ~n49956 ;
  assign n49958 = n21779 | n29619 ;
  assign n49959 = n34760 | n49958 ;
  assign n49960 = n40726 ^ n24889 ^ 1'b0 ;
  assign n49961 = n11755 | n46944 ;
  assign n49962 = n18888 ^ n8414 ^ 1'b0 ;
  assign n49963 = ( n4079 & n49961 ) | ( n4079 & n49962 ) | ( n49961 & n49962 ) ;
  assign n49964 = n38572 ^ n36388 ^ n31854 ;
  assign n49965 = ~n16336 & n31675 ;
  assign n49966 = ~n28913 & n49965 ;
  assign n49967 = n36948 ^ n14649 ^ 1'b0 ;
  assign n49968 = n41772 & n49967 ;
  assign n49969 = n9700 | n26004 ;
  assign n49970 = n1647 | n13789 ;
  assign n49971 = n49970 ^ n4321 ^ 1'b0 ;
  assign n49972 = n35057 ^ n24744 ^ 1'b0 ;
  assign n49973 = n6528 & n37039 ;
  assign n49974 = ( n3664 & n6095 ) | ( n3664 & ~n7513 ) | ( n6095 & ~n7513 ) ;
  assign n49975 = n49974 ^ n38162 ^ 1'b0 ;
  assign n49976 = n19047 & ~n27902 ;
  assign n49977 = n28170 ^ n19984 ^ 1'b0 ;
  assign n49978 = n32880 | n49977 ;
  assign n49979 = n30069 ^ n9670 ^ n9421 ;
  assign n49980 = n1949 & ~n16891 ;
  assign n49981 = ~n29475 & n49980 ;
  assign n49982 = n8507 | n49981 ;
  assign n49983 = n4072 & n9773 ;
  assign n49984 = n11868 & n49983 ;
  assign n49985 = n49984 ^ n8670 ^ 1'b0 ;
  assign n49986 = ~n29741 & n46956 ;
  assign n49987 = n43603 ^ n3544 ^ 1'b0 ;
  assign n49988 = n18029 | n49987 ;
  assign n49989 = n6964 & ~n49988 ;
  assign n49990 = n32992 & n49989 ;
  assign n49991 = n49990 ^ n12344 ^ 1'b0 ;
  assign n49992 = n39488 ^ n12346 ^ 1'b0 ;
  assign n49993 = n32168 & n49992 ;
  assign n49994 = n48024 ^ n12458 ^ 1'b0 ;
  assign n49995 = n18305 | n49994 ;
  assign n49996 = n24928 & ~n49122 ;
  assign n49997 = n16523 & n34734 ;
  assign n49998 = n20938 & ~n35226 ;
  assign n49999 = n35510 ^ n688 ^ 1'b0 ;
  assign n50000 = n318 & n20391 ;
  assign n50001 = n19747 & n50000 ;
  assign n50002 = n3147 & ~n23785 ;
  assign n50003 = n7008 & n50002 ;
  assign n50004 = n15515 ^ n5747 ^ 1'b0 ;
  assign n50005 = ~n2930 & n50004 ;
  assign n50006 = n44625 ^ n4380 ^ 1'b0 ;
  assign n50007 = n50005 & n50006 ;
  assign n50008 = ( ~n50001 & n50003 ) | ( ~n50001 & n50007 ) | ( n50003 & n50007 ) ;
  assign n50009 = n12323 ^ n8749 ^ 1'b0 ;
  assign n50010 = n4139 & ~n50009 ;
  assign n50011 = n3136 & ~n4122 ;
  assign n50012 = n5863 & n41763 ;
  assign n50013 = ~n22951 & n50012 ;
  assign n50014 = ~n9022 & n12456 ;
  assign n50015 = ~n48024 & n50014 ;
  assign n50016 = n20546 ^ n2923 ^ 1'b0 ;
  assign n50017 = n22756 ^ n571 ^ 1'b0 ;
  assign n50018 = n29294 ^ n6248 ^ 1'b0 ;
  assign n50019 = ~n1024 & n4151 ;
  assign n50020 = n19401 | n50019 ;
  assign n50021 = n19590 & ~n50020 ;
  assign n50022 = n50021 ^ n40773 ^ 1'b0 ;
  assign n50023 = n17845 & ~n25637 ;
  assign n50024 = n50023 ^ n39448 ^ 1'b0 ;
  assign n50025 = n41866 & ~n50024 ;
  assign n50026 = n6236 ^ n492 ^ 1'b0 ;
  assign n50027 = n4971 & ~n50026 ;
  assign n50028 = n8266 | n40279 ;
  assign n50029 = n24747 | n38423 ;
  assign n50030 = ~n19896 & n33065 ;
  assign n50031 = ~n1178 & n34405 ;
  assign n50032 = ~n50030 & n50031 ;
  assign n50033 = n20233 ^ n7921 ^ 1'b0 ;
  assign n50034 = n24491 ^ n13878 ^ 1'b0 ;
  assign n50035 = n14034 | n27164 ;
  assign n50036 = n43190 ^ n16458 ^ 1'b0 ;
  assign n50037 = n50036 ^ n17887 ^ n2161 ;
  assign n50038 = ~n2489 & n5592 ;
  assign n50039 = n50038 ^ n25316 ^ 1'b0 ;
  assign n50040 = n8195 & ~n50039 ;
  assign n50041 = ~n8387 & n50040 ;
  assign n50042 = n9122 ^ n445 ^ 1'b0 ;
  assign n50043 = n50042 ^ n28363 ^ 1'b0 ;
  assign n50044 = ~n8405 & n14425 ;
  assign n50045 = ~n10660 & n10971 ;
  assign n50046 = n50045 ^ n6149 ^ 1'b0 ;
  assign n50047 = n7430 | n50046 ;
  assign n50050 = ( ~n5627 & n8232 ) | ( ~n5627 & n16283 ) | ( n8232 & n16283 ) ;
  assign n50048 = n552 & n15592 ;
  assign n50049 = n30727 | n50048 ;
  assign n50051 = n50050 ^ n50049 ^ 1'b0 ;
  assign n50052 = n12533 | n43190 ;
  assign n50053 = n20801 & ~n50052 ;
  assign n50054 = n37723 & ~n50053 ;
  assign n50055 = ~n49961 & n50054 ;
  assign n50056 = ~n2781 & n21480 ;
  assign n50057 = n50056 ^ n43662 ^ 1'b0 ;
  assign n50058 = n30593 | n50057 ;
  assign n50059 = n41181 ^ n3071 ^ 1'b0 ;
  assign n50060 = n12655 ^ n5354 ^ 1'b0 ;
  assign n50061 = n1032 & ~n50060 ;
  assign n50062 = n50061 ^ n45534 ^ 1'b0 ;
  assign n50063 = ( n2895 & ~n4696 ) | ( n2895 & n50062 ) | ( ~n4696 & n50062 ) ;
  assign n50064 = n22385 & n47261 ;
  assign n50065 = ~n33521 & n50064 ;
  assign n50066 = n194 & ~n6345 ;
  assign n50067 = n50066 ^ n34588 ^ n22022 ;
  assign n50068 = n2570 & n22913 ;
  assign n50069 = n11402 & n34901 ;
  assign n50070 = n31530 & n50069 ;
  assign n50071 = n21451 | n29319 ;
  assign n50072 = n22470 ^ n9219 ^ 1'b0 ;
  assign n50073 = n907 & ~n17563 ;
  assign n50074 = ~n50072 & n50073 ;
  assign n50075 = n14657 ^ n130 ^ 1'b0 ;
  assign n50076 = ~n9047 & n50075 ;
  assign n50077 = n37423 & n50076 ;
  assign n50078 = n46362 & n50077 ;
  assign n50079 = n3066 & n10352 ;
  assign n50080 = n20071 & n50079 ;
  assign n50081 = ~n3393 & n50080 ;
  assign n50082 = n1201 | n50081 ;
  assign n50083 = n8610 ^ n6272 ^ 1'b0 ;
  assign n50084 = ~n29458 & n50083 ;
  assign n50086 = n14670 ^ n5284 ^ n4668 ;
  assign n50085 = n2261 & ~n37177 ;
  assign n50087 = n50086 ^ n50085 ^ 1'b0 ;
  assign n50088 = n395 & ~n29279 ;
  assign n50089 = ~n50087 & n50088 ;
  assign n50090 = n50089 ^ n29312 ^ 1'b0 ;
  assign n50091 = ~n19400 & n50090 ;
  assign n50092 = n13193 | n27996 ;
  assign n50093 = ~n8529 & n24365 ;
  assign n50094 = n50093 ^ n6759 ^ 1'b0 ;
  assign n50095 = n25956 ^ n17932 ^ 1'b0 ;
  assign n50096 = n27723 | n38040 ;
  assign n50097 = n30989 | n43956 ;
  assign n50098 = n50097 ^ n6326 ^ 1'b0 ;
  assign n50099 = n7839 ^ n4681 ^ 1'b0 ;
  assign n50100 = n12788 | n34101 ;
  assign n50101 = n17789 & ~n26613 ;
  assign n50102 = ~n28200 & n33049 ;
  assign n50103 = ~n50101 & n50102 ;
  assign n50104 = n28133 & ~n50103 ;
  assign n50105 = n50100 & ~n50104 ;
  assign n50106 = n29900 ^ n11060 ^ 1'b0 ;
  assign n50107 = n376 & ~n18336 ;
  assign n50108 = n50107 ^ n3031 ^ 1'b0 ;
  assign n50109 = n12165 & ~n35516 ;
  assign n50110 = n50109 ^ n39627 ^ 1'b0 ;
  assign n50111 = n15622 ^ n12271 ^ 1'b0 ;
  assign n50112 = n10823 & ~n50111 ;
  assign n50113 = n50112 ^ n40785 ^ 1'b0 ;
  assign n50114 = n12643 & ~n50113 ;
  assign n50115 = n50114 ^ n33638 ^ 1'b0 ;
  assign n50118 = ~n6953 & n9098 ;
  assign n50116 = n27635 | n43487 ;
  assign n50117 = n29389 & ~n50116 ;
  assign n50119 = n50118 ^ n50117 ^ 1'b0 ;
  assign n50120 = n16485 | n41921 ;
  assign n50121 = n29297 & n50120 ;
  assign n50122 = n18244 & n30550 ;
  assign n50125 = n372 & ~n5911 ;
  assign n50126 = n105 & n50125 ;
  assign n50124 = n13524 | n43681 ;
  assign n50127 = n50126 ^ n50124 ^ 1'b0 ;
  assign n50123 = ~n34116 & n41861 ;
  assign n50128 = n50127 ^ n50123 ^ n39484 ;
  assign n50129 = n3566 | n4856 ;
  assign n50131 = n38659 ^ n35751 ^ n14806 ;
  assign n50130 = ~n19737 & n24827 ;
  assign n50132 = n50131 ^ n50130 ^ 1'b0 ;
  assign n50133 = n25025 ^ n4485 ^ 1'b0 ;
  assign n50134 = n12516 ^ n2527 ^ 1'b0 ;
  assign n50135 = n17548 & n50134 ;
  assign n50138 = n15698 | n39856 ;
  assign n50139 = ( ~n9696 & n35380 ) | ( ~n9696 & n50138 ) | ( n35380 & n50138 ) ;
  assign n50136 = n15809 | n23001 ;
  assign n50137 = n11309 & ~n50136 ;
  assign n50140 = n50139 ^ n50137 ^ n1217 ;
  assign n50141 = n40575 ^ n11193 ^ n4321 ;
  assign n50142 = n10556 & ~n50141 ;
  assign n50144 = ~n2265 & n24726 ;
  assign n50143 = n10809 & ~n17022 ;
  assign n50145 = n50144 ^ n50143 ^ 1'b0 ;
  assign n50146 = n20113 ^ n10770 ^ 1'b0 ;
  assign n50147 = ~n50145 & n50146 ;
  assign n50148 = n50147 ^ n3372 ^ 1'b0 ;
  assign n50149 = n41310 ^ n10717 ^ 1'b0 ;
  assign n50150 = n29392 | n50149 ;
  assign n50152 = n24380 ^ n6656 ^ 1'b0 ;
  assign n50151 = n21981 | n25851 ;
  assign n50153 = n50152 ^ n50151 ^ 1'b0 ;
  assign n50154 = ( n737 & ~n12426 ) | ( n737 & n26991 ) | ( ~n12426 & n26991 ) ;
  assign n50155 = n15049 | n23817 ;
  assign n50156 = n3761 | n14066 ;
  assign n50157 = n50156 ^ n1422 ^ 1'b0 ;
  assign n50158 = n15431 ^ n3610 ^ 1'b0 ;
  assign n50159 = ~n46293 & n50158 ;
  assign n50160 = ~n2461 & n50159 ;
  assign n50161 = n20970 ^ n10572 ^ 1'b0 ;
  assign n50162 = ~n5637 & n50161 ;
  assign n50163 = ( ~n15668 & n39615 ) | ( ~n15668 & n50162 ) | ( n39615 & n50162 ) ;
  assign n50164 = n1915 | n31328 ;
  assign n50165 = n50164 ^ n1534 ^ 1'b0 ;
  assign n50166 = n4242 & n50165 ;
  assign n50167 = ~n27819 & n29020 ;
  assign n50168 = ~n45791 & n50104 ;
  assign n50169 = n49322 & n50168 ;
  assign n50170 = ( n4033 & n19799 ) | ( n4033 & ~n35589 ) | ( n19799 & ~n35589 ) ;
  assign n50171 = ~n17869 & n50170 ;
  assign n50172 = n50171 ^ n2346 ^ 1'b0 ;
  assign n50173 = n38630 | n50172 ;
  assign n50174 = ~n21241 & n36187 ;
  assign n50175 = ( ~n6833 & n13097 ) | ( ~n6833 & n33778 ) | ( n13097 & n33778 ) ;
  assign n50176 = n7405 & ~n50175 ;
  assign n50177 = n33708 ^ n31681 ^ 1'b0 ;
  assign n50178 = n28641 ^ n5406 ^ 1'b0 ;
  assign n50179 = ( n2980 & n23491 ) | ( n2980 & ~n50178 ) | ( n23491 & ~n50178 ) ;
  assign n50180 = n4926 ^ n3146 ^ 1'b0 ;
  assign n50181 = n7421 & ~n50180 ;
  assign n50182 = ( ~n7338 & n10403 ) | ( ~n7338 & n50181 ) | ( n10403 & n50181 ) ;
  assign n50183 = ~n34002 & n50182 ;
  assign n50184 = n50183 ^ n45779 ^ 1'b0 ;
  assign n50185 = n46618 ^ n22502 ^ 1'b0 ;
  assign n50186 = n1655 | n13555 ;
  assign n50187 = n582 & n32678 ;
  assign n50188 = n50187 ^ n3721 ^ 1'b0 ;
  assign n50189 = n16532 & n42299 ;
  assign n50190 = n493 | n50189 ;
  assign n50191 = n8879 & ~n12949 ;
  assign n50192 = n9915 & n50191 ;
  assign n50193 = n50192 ^ n10513 ^ 1'b0 ;
  assign n50194 = n9751 & ~n26201 ;
  assign n50195 = n1958 & ~n42200 ;
  assign n50196 = ~n6210 & n50195 ;
  assign n50197 = n231 & n30404 ;
  assign n50198 = n33388 & n50197 ;
  assign n50199 = n25971 ^ n7167 ^ 1'b0 ;
  assign n50200 = ~n1792 & n50199 ;
  assign n50203 = n19365 & n34468 ;
  assign n50201 = n4674 | n12717 ;
  assign n50202 = ~n21993 & n50201 ;
  assign n50204 = n50203 ^ n50202 ^ 1'b0 ;
  assign n50205 = n36542 ^ n33817 ^ n5344 ;
  assign n50206 = n26380 ^ n16554 ^ n1069 ;
  assign n50207 = n8625 & n12495 ;
  assign n50208 = n26476 & n50207 ;
  assign n50209 = n20817 & ~n45689 ;
  assign n50210 = n8188 & n50209 ;
  assign n50211 = n15976 ^ n6485 ^ 1'b0 ;
  assign n50212 = n35911 & n50211 ;
  assign n50213 = n263 | n5155 ;
  assign n50214 = n10055 | n50213 ;
  assign n50215 = n50212 | n50214 ;
  assign n50216 = n4988 | n46833 ;
  assign n50217 = n21954 & n41685 ;
  assign n50218 = ~n29628 & n39837 ;
  assign n50219 = n10187 | n29990 ;
  assign n50220 = n50219 ^ n13698 ^ 1'b0 ;
  assign n50221 = n50220 ^ n19934 ^ 1'b0 ;
  assign n50222 = ~n16651 & n29700 ;
  assign n50223 = n50222 ^ n1802 ^ 1'b0 ;
  assign n50224 = n50030 ^ n38036 ^ 1'b0 ;
  assign n50225 = n4059 | n25245 ;
  assign n50226 = n27277 | n44295 ;
  assign n50227 = ~n36553 & n38792 ;
  assign n50228 = n38697 ^ n24016 ^ 1'b0 ;
  assign n50230 = ~n7475 & n7873 ;
  assign n50229 = n11582 ^ n6662 ^ n494 ;
  assign n50231 = n50230 ^ n50229 ^ 1'b0 ;
  assign n50232 = n4709 & ~n50231 ;
  assign n50233 = ~n8704 & n16591 ;
  assign n50234 = n12596 ^ n8443 ^ 1'b0 ;
  assign n50235 = n508 | n50234 ;
  assign n50236 = ( ~n12109 & n15523 ) | ( ~n12109 & n50235 ) | ( n15523 & n50235 ) ;
  assign n50237 = n38547 ^ n20702 ^ n3447 ;
  assign n50238 = ~n494 & n27654 ;
  assign n50239 = n16319 | n50238 ;
  assign n50240 = n10278 | n14075 ;
  assign n50241 = n15008 ^ n11005 ^ 1'b0 ;
  assign n50242 = n21843 | n50241 ;
  assign n50243 = n7952 & ~n50242 ;
  assign n50244 = ~n50240 & n50243 ;
  assign n50245 = ~n3556 & n26912 ;
  assign n50246 = ~n5158 & n5365 ;
  assign n50247 = n50246 ^ n38048 ^ n2438 ;
  assign n50248 = n15317 & n20333 ;
  assign n50249 = n13883 & ~n33311 ;
  assign n50250 = ~n25217 & n50249 ;
  assign n50251 = n21736 & ~n22689 ;
  assign n50252 = ~n6527 & n12839 ;
  assign n50253 = n50252 ^ n50126 ^ 1'b0 ;
  assign n50254 = n50253 ^ n2940 ^ 1'b0 ;
  assign n50255 = n7067 & n50254 ;
  assign n50256 = n10560 & ~n50255 ;
  assign n50257 = n2584 | n20050 ;
  assign n50258 = n36776 & ~n50257 ;
  assign n50259 = n14243 | n24221 ;
  assign n50260 = n7358 | n50259 ;
  assign n50261 = n30582 ^ n6534 ^ 1'b0 ;
  assign n50262 = n50260 & n50261 ;
  assign n50263 = n24621 ^ n14053 ^ 1'b0 ;
  assign n50264 = ~n7568 & n21636 ;
  assign n50265 = n50264 ^ n31998 ^ 1'b0 ;
  assign n50266 = n43466 ^ n29784 ^ n6813 ;
  assign n50267 = ( n12053 & n16809 ) | ( n12053 & n50266 ) | ( n16809 & n50266 ) ;
  assign n50268 = n18246 | n50267 ;
  assign n50269 = ~n5459 & n11077 ;
  assign n50270 = n50269 ^ n13578 ^ 1'b0 ;
  assign n50271 = n50270 ^ n35257 ^ n465 ;
  assign n50272 = ( n37828 & ~n44065 ) | ( n37828 & n50271 ) | ( ~n44065 & n50271 ) ;
  assign n50273 = ( n7569 & ~n11757 ) | ( n7569 & n11810 ) | ( ~n11757 & n11810 ) ;
  assign n50274 = ~n4032 & n25379 ;
  assign n50275 = ~n22035 & n24480 ;
  assign n50276 = n4248 | n5580 ;
  assign n50277 = n6300 & ~n50276 ;
  assign n50278 = n12799 | n31524 ;
  assign n50279 = ( n4246 & n50277 ) | ( n4246 & n50278 ) | ( n50277 & n50278 ) ;
  assign n50280 = n13665 & n41280 ;
  assign n50281 = n3790 & n18516 ;
  assign n50282 = n50281 ^ n45276 ^ 1'b0 ;
  assign n50284 = n27404 ^ n24992 ^ 1'b0 ;
  assign n50285 = ~n33538 & n50284 ;
  assign n50283 = ~n8244 & n14808 ;
  assign n50286 = n50285 ^ n50283 ^ 1'b0 ;
  assign n50287 = n10343 | n16811 ;
  assign n50288 = n50287 ^ n14989 ^ 1'b0 ;
  assign n50289 = ~n33257 & n50288 ;
  assign n50290 = n50289 ^ n15096 ^ 1'b0 ;
  assign n50291 = n3761 | n50290 ;
  assign n50292 = n50291 ^ n695 ^ 1'b0 ;
  assign n50293 = n7958 | n12055 ;
  assign n50294 = n2650 | n50293 ;
  assign n50295 = n1300 & ~n24207 ;
  assign n50296 = ~n50294 & n50295 ;
  assign n50297 = ~n50292 & n50296 ;
  assign n50301 = n24930 & ~n25385 ;
  assign n50298 = n10107 ^ n6704 ^ 1'b0 ;
  assign n50299 = n28161 | n50298 ;
  assign n50300 = n50299 ^ n36821 ^ n8313 ;
  assign n50302 = n50301 ^ n50300 ^ 1'b0 ;
  assign n50303 = n12456 | n44176 ;
  assign n50304 = ( n619 & n2602 ) | ( n619 & n50303 ) | ( n2602 & n50303 ) ;
  assign n50305 = n9267 ^ n2367 ^ 1'b0 ;
  assign n50306 = ~n29142 & n50305 ;
  assign n50307 = ~n173 & n5776 ;
  assign n50308 = ~n9219 & n50307 ;
  assign n50309 = ~n6283 & n50308 ;
  assign n50310 = n50309 ^ n42211 ^ n6267 ;
  assign n50311 = n1542 & n50310 ;
  assign n50312 = n2801 & ~n32898 ;
  assign n50313 = ~n14577 & n50312 ;
  assign n50314 = n667 & ~n10839 ;
  assign n50315 = n4870 & n4968 ;
  assign n50316 = ( n18516 & n20163 ) | ( n18516 & ~n36302 ) | ( n20163 & ~n36302 ) ;
  assign n50317 = n840 & ~n12098 ;
  assign n50318 = n50317 ^ n11175 ^ 1'b0 ;
  assign n50319 = n45633 ^ n9148 ^ 1'b0 ;
  assign n50320 = n6856 ^ n5374 ^ 1'b0 ;
  assign n50321 = n205 & n33515 ;
  assign n50322 = ~n13937 & n38085 ;
  assign n50323 = ~n30557 & n50322 ;
  assign n50324 = n18986 & n30391 ;
  assign n50326 = n17321 & n20370 ;
  assign n50325 = n18617 & n46099 ;
  assign n50327 = n50326 ^ n50325 ^ 1'b0 ;
  assign n50328 = ~n4015 & n38880 ;
  assign n50329 = n1868 | n1988 ;
  assign n50330 = n4718 | n18966 ;
  assign n50331 = n71 | n1378 ;
  assign n50332 = n50330 & ~n50331 ;
  assign n50333 = n2048 ^ n436 ^ 1'b0 ;
  assign n50334 = n18867 | n50333 ;
  assign n50335 = n39945 ^ n7052 ^ 1'b0 ;
  assign n50336 = ~n20520 & n43250 ;
  assign n50337 = n50336 ^ n344 ^ 1'b0 ;
  assign n50338 = n11342 & n18647 ;
  assign n50339 = n15393 & n50338 ;
  assign n50340 = n11105 | n43835 ;
  assign n50341 = n50339 & ~n50340 ;
  assign n50342 = ~n15562 & n24776 ;
  assign n50343 = ~n1853 & n2231 ;
  assign n50344 = n50343 ^ n39020 ^ 1'b0 ;
  assign n50346 = n13559 & ~n14757 ;
  assign n50345 = n5453 & ~n22948 ;
  assign n50347 = n50346 ^ n50345 ^ 1'b0 ;
  assign n50348 = n45363 ^ n30897 ^ 1'b0 ;
  assign n50349 = n26064 ^ n22872 ^ 1'b0 ;
  assign n50350 = n50120 ^ n6551 ^ 1'b0 ;
  assign n50351 = ~n8554 & n21192 ;
  assign n50352 = n9926 & ~n33017 ;
  assign n50353 = n810 & n11384 ;
  assign n50354 = ~n50352 & n50353 ;
  assign n50355 = ~n6899 & n17387 ;
  assign n50356 = n12038 | n35226 ;
  assign n50357 = n50355 & n50356 ;
  assign n50358 = n42442 | n50357 ;
  assign n50359 = n50358 ^ n29407 ^ 1'b0 ;
  assign n50360 = n3131 & n19619 ;
  assign n50361 = n13061 & ~n50360 ;
  assign n50362 = n20281 & n50361 ;
  assign n50363 = ~n20433 & n27963 ;
  assign n50364 = n50363 ^ n15392 ^ 1'b0 ;
  assign n50365 = ~n50362 & n50364 ;
  assign n50366 = ( n1066 & n8283 ) | ( n1066 & ~n27871 ) | ( n8283 & ~n27871 ) ;
  assign n50367 = n50366 ^ n7278 ^ 1'b0 ;
  assign n50368 = n45228 & n48576 ;
  assign n50369 = n1897 & n10106 ;
  assign n50370 = n50369 ^ n30676 ^ n1880 ;
  assign n50371 = n31872 ^ n27106 ^ n9139 ;
  assign n50372 = ~n4010 & n43270 ;
  assign n50373 = n50372 ^ n34719 ^ 1'b0 ;
  assign n50374 = n27568 | n38122 ;
  assign n50375 = n50374 ^ n37746 ^ 1'b0 ;
  assign n50376 = n7899 ^ n5109 ^ 1'b0 ;
  assign n50377 = n40869 & ~n50376 ;
  assign n50378 = n50377 ^ n17730 ^ 1'b0 ;
  assign n50379 = n9356 & ~n50378 ;
  assign n50380 = n12305 | n48886 ;
  assign n50382 = n8589 ^ n801 ^ 1'b0 ;
  assign n50383 = n14386 & n50382 ;
  assign n50381 = n10951 & n41855 ;
  assign n50384 = n50383 ^ n50381 ^ n20046 ;
  assign n50385 = n24200 ^ n23490 ^ 1'b0 ;
  assign n50386 = n1523 | n32274 ;
  assign n50390 = n24837 ^ n4170 ^ 1'b0 ;
  assign n50391 = n9983 & ~n50390 ;
  assign n50387 = n18578 ^ n12466 ^ 1'b0 ;
  assign n50388 = n31298 & ~n50387 ;
  assign n50389 = ~n32598 & n50388 ;
  assign n50392 = n50391 ^ n50389 ^ 1'b0 ;
  assign n50393 = n5540 ^ n3544 ^ 1'b0 ;
  assign n50394 = n41840 & ~n50393 ;
  assign n50395 = n29983 & ~n50394 ;
  assign n50396 = ( n3364 & ~n6917 ) | ( n3364 & n11859 ) | ( ~n6917 & n11859 ) ;
  assign n50397 = n50396 ^ n44488 ^ n42169 ;
  assign n50398 = n9468 | n20271 ;
  assign n50399 = n50397 | n50398 ;
  assign n50400 = n5507 ^ n4477 ^ 1'b0 ;
  assign n50401 = n1591 & n50400 ;
  assign n50402 = n3669 & n50401 ;
  assign n50403 = ~n50399 & n50402 ;
  assign n50404 = n9088 ^ n3731 ^ 1'b0 ;
  assign n50405 = n22654 & ~n24335 ;
  assign n50407 = n2317 & n43735 ;
  assign n50406 = ~n17620 & n23399 ;
  assign n50408 = n50407 ^ n50406 ^ n3970 ;
  assign n50409 = n16637 ^ n9964 ^ 1'b0 ;
  assign n50410 = n20239 & n50409 ;
  assign n50411 = n15650 | n46224 ;
  assign n50412 = n7734 ^ n5664 ^ 1'b0 ;
  assign n50413 = ~n4036 & n17899 ;
  assign n50414 = n50413 ^ n8117 ^ 1'b0 ;
  assign n50415 = ~n50412 & n50414 ;
  assign n50416 = n12299 & n26562 ;
  assign n50417 = n18442 & n50416 ;
  assign n50418 = n27886 ^ n6344 ^ 1'b0 ;
  assign n50419 = n28785 & n50418 ;
  assign n50420 = n50419 ^ n26168 ^ 1'b0 ;
  assign n50421 = n48840 & n50420 ;
  assign n50423 = ~n25124 & n46675 ;
  assign n50424 = n50423 ^ n690 ^ 1'b0 ;
  assign n50422 = n33670 ^ n17903 ^ 1'b0 ;
  assign n50425 = n50424 ^ n50422 ^ 1'b0 ;
  assign n50426 = n34846 ^ n7087 ^ 1'b0 ;
  assign n50427 = n29918 ^ n677 ^ 1'b0 ;
  assign n50428 = ~n27094 & n50427 ;
  assign n50429 = ( n25160 & n30397 ) | ( n25160 & ~n50428 ) | ( n30397 & ~n50428 ) ;
  assign n50430 = n50429 ^ n34729 ^ n15635 ;
  assign n50431 = n1306 | n16718 ;
  assign n50432 = n50430 | n50431 ;
  assign n50433 = n9421 | n26532 ;
  assign n50434 = n44966 & ~n50433 ;
  assign n50435 = n3970 ^ n125 ^ 1'b0 ;
  assign n50436 = n11056 | n38712 ;
  assign n50437 = n14985 ^ n11951 ^ 1'b0 ;
  assign n50438 = ~n4406 & n50437 ;
  assign n50439 = n50438 ^ n47181 ^ 1'b0 ;
  assign n50440 = n21253 ^ n4583 ^ 1'b0 ;
  assign n50441 = ~n5783 & n46726 ;
  assign n50442 = n26550 ^ n11383 ^ 1'b0 ;
  assign n50443 = ~n50441 & n50442 ;
  assign n50444 = n50443 ^ n37469 ^ 1'b0 ;
  assign n50445 = n6292 & ~n8341 ;
  assign n50446 = n20041 & n50445 ;
  assign n50447 = n28070 | n50446 ;
  assign n50448 = n1997 | n20602 ;
  assign n50449 = n11246 & ~n50448 ;
  assign n50450 = n11613 | n43155 ;
  assign n50451 = n50450 ^ n47000 ^ 1'b0 ;
  assign n50452 = ~n32252 & n50451 ;
  assign n50454 = n35682 & n39089 ;
  assign n50455 = n50454 ^ n14555 ^ 1'b0 ;
  assign n50453 = n1627 & ~n22619 ;
  assign n50456 = n50455 ^ n50453 ^ 1'b0 ;
  assign n50457 = ~n27914 & n38167 ;
  assign n50458 = n24696 & n50457 ;
  assign n50459 = n3762 & n13926 ;
  assign n50460 = ~n7542 & n16283 ;
  assign n50461 = n4264 & ~n14487 ;
  assign n50462 = n50461 ^ n3060 ^ 1'b0 ;
  assign n50463 = n12588 & ~n50462 ;
  assign n50464 = n50463 ^ n20880 ^ 1'b0 ;
  assign n50465 = n30612 ^ n2461 ^ 1'b0 ;
  assign n50466 = n19846 | n38828 ;
  assign n50467 = n50466 ^ n18619 ^ 1'b0 ;
  assign n50468 = n3617 | n50467 ;
  assign n50469 = n11095 & ~n50468 ;
  assign n50470 = n45363 & n50469 ;
  assign n50471 = n49732 ^ n18502 ^ 1'b0 ;
  assign n50472 = n18019 ^ n14053 ^ 1'b0 ;
  assign n50473 = n6994 ^ n6472 ^ 1'b0 ;
  assign n50474 = n47001 | n50473 ;
  assign n50475 = ~n29164 & n49787 ;
  assign n50476 = ~n24953 & n50475 ;
  assign n50477 = n24755 & n31549 ;
  assign n50478 = n48780 & n50477 ;
  assign n50479 = n50478 ^ n50100 ^ n28941 ;
  assign n50481 = ( n6858 & n21593 ) | ( n6858 & n36507 ) | ( n21593 & n36507 ) ;
  assign n50480 = n15509 & n39686 ;
  assign n50482 = n50481 ^ n50480 ^ 1'b0 ;
  assign n50483 = n28938 ^ n27087 ^ 1'b0 ;
  assign n50484 = n1528 & n31329 ;
  assign n50485 = n26164 ^ n6405 ^ 1'b0 ;
  assign n50486 = ~n5815 & n20706 ;
  assign n50487 = n50485 & n50486 ;
  assign n50488 = n13737 & ~n21531 ;
  assign n50489 = n1083 & ~n17707 ;
  assign n50490 = n13406 | n21881 ;
  assign n50491 = n14866 & ~n50490 ;
  assign n50492 = n50491 ^ n24084 ^ 1'b0 ;
  assign n50493 = n29810 ^ n29032 ^ 1'b0 ;
  assign n50494 = n20460 ^ n8640 ^ 1'b0 ;
  assign n50495 = n8230 ^ n1323 ^ 1'b0 ;
  assign n50501 = n49787 ^ n15332 ^ 1'b0 ;
  assign n50496 = n6203 ^ n1753 ^ 1'b0 ;
  assign n50497 = ~n15051 & n50496 ;
  assign n50498 = n14614 & ~n50497 ;
  assign n50499 = n9084 | n50498 ;
  assign n50500 = n50499 ^ n13755 ^ 1'b0 ;
  assign n50502 = n50501 ^ n50500 ^ 1'b0 ;
  assign n50503 = n4636 & ~n20143 ;
  assign y0 = x3 ;
  assign y1 = x9 ;
  assign y2 = x10 ;
  assign y3 = ~n13 ;
  assign y4 = ~n15 ;
  assign y5 = ~n17 ;
  assign y6 = ~n19 ;
  assign y7 = ~n20 ;
  assign y8 = ~n21 ;
  assign y9 = ~1'b0 ;
  assign y10 = ~n31 ;
  assign y11 = ~n35 ;
  assign y12 = n36 ;
  assign y13 = n38 ;
  assign y14 = n49 ;
  assign y15 = n51 ;
  assign y16 = n58 ;
  assign y17 = n63 ;
  assign y18 = ~n69 ;
  assign y19 = ~1'b0 ;
  assign y20 = ~n71 ;
  assign y21 = n73 ;
  assign y22 = n74 ;
  assign y23 = ~1'b0 ;
  assign y24 = n76 ;
  assign y25 = x6 ;
  assign y26 = n83 ;
  assign y27 = ~n85 ;
  assign y28 = n91 ;
  assign y29 = ~n93 ;
  assign y30 = ~1'b0 ;
  assign y31 = ~1'b0 ;
  assign y32 = ~n100 ;
  assign y33 = ~n104 ;
  assign y34 = ~1'b0 ;
  assign y35 = n56 ;
  assign y36 = ~1'b0 ;
  assign y37 = ~n106 ;
  assign y38 = ~n112 ;
  assign y39 = ~1'b0 ;
  assign y40 = n113 ;
  assign y41 = ~n119 ;
  assign y42 = ~1'b0 ;
  assign y43 = ~1'b0 ;
  assign y44 = ~n122 ;
  assign y45 = n124 ;
  assign y46 = ~1'b0 ;
  assign y47 = n126 ;
  assign y48 = ~1'b0 ;
  assign y49 = ~n127 ;
  assign y50 = ~1'b0 ;
  assign y51 = n129 ;
  assign y52 = ~n131 ;
  assign y53 = n132 ;
  assign y54 = ~1'b0 ;
  assign y55 = ~n136 ;
  assign y56 = ~n140 ;
  assign y57 = ~n142 ;
  assign y58 = n144 ;
  assign y59 = ~1'b0 ;
  assign y60 = ~n148 ;
  assign y61 = ~n150 ;
  assign y62 = ~n154 ;
  assign y63 = n160 ;
  assign y64 = ~n162 ;
  assign y65 = ~1'b0 ;
  assign y66 = n164 ;
  assign y67 = n171 ;
  assign y68 = ~n177 ;
  assign y69 = n182 ;
  assign y70 = 1'b0 ;
  assign y71 = ~1'b0 ;
  assign y72 = ~n183 ;
  assign y73 = ~n184 ;
  assign y74 = ~1'b0 ;
  assign y75 = ~1'b0 ;
  assign y76 = ~n189 ;
  assign y77 = ~n191 ;
  assign y78 = ~n195 ;
  assign y79 = ~1'b0 ;
  assign y80 = ~n152 ;
  assign y81 = ~n202 ;
  assign y82 = ~n207 ;
  assign y83 = n212 ;
  assign y84 = n216 ;
  assign y85 = ~n219 ;
  assign y86 = n220 ;
  assign y87 = ~1'b0 ;
  assign y88 = n225 ;
  assign y89 = n231 ;
  assign y90 = n233 ;
  assign y91 = ~n234 ;
  assign y92 = n237 ;
  assign y93 = n239 ;
  assign y94 = ~n244 ;
  assign y95 = n246 ;
  assign y96 = n249 ;
  assign y97 = ~n250 ;
  assign y98 = n254 ;
  assign y99 = ~1'b0 ;
  assign y100 = n259 ;
  assign y101 = ~1'b0 ;
  assign y102 = n260 ;
  assign y103 = n264 ;
  assign y104 = ~n265 ;
  assign y105 = n267 ;
  assign y106 = n269 ;
  assign y107 = n271 ;
  assign y108 = ~n275 ;
  assign y109 = ~1'b0 ;
  assign y110 = ~n277 ;
  assign y111 = n279 ;
  assign y112 = n282 ;
  assign y113 = ~1'b0 ;
  assign y114 = n286 ;
  assign y115 = ~n291 ;
  assign y116 = n292 ;
  assign y117 = ~n296 ;
  assign y118 = ~1'b0 ;
  assign y119 = ~1'b0 ;
  assign y120 = ~n297 ;
  assign y121 = n299 ;
  assign y122 = n301 ;
  assign y123 = n306 ;
  assign y124 = ~n309 ;
  assign y125 = ~n312 ;
  assign y126 = ~n316 ;
  assign y127 = ~n325 ;
  assign y128 = ~1'b0 ;
  assign y129 = 1'b0 ;
  assign y130 = n331 ;
  assign y131 = n334 ;
  assign y132 = ~n335 ;
  assign y133 = n336 ;
  assign y134 = n338 ;
  assign y135 = ~n347 ;
  assign y136 = n349 ;
  assign y137 = ~n352 ;
  assign y138 = n358 ;
  assign y139 = ~n362 ;
  assign y140 = ~n366 ;
  assign y141 = n367 ;
  assign y142 = ~n368 ;
  assign y143 = n376 ;
  assign y144 = ~1'b0 ;
  assign y145 = ~1'b0 ;
  assign y146 = ~n379 ;
  assign y147 = n382 ;
  assign y148 = n388 ;
  assign y149 = ~1'b0 ;
  assign y150 = ~n393 ;
  assign y151 = ~1'b0 ;
  assign y152 = ~1'b0 ;
  assign y153 = ~n362 ;
  assign y154 = ~1'b0 ;
  assign y155 = ~1'b0 ;
  assign y156 = ~1'b0 ;
  assign y157 = ~n397 ;
  assign y158 = n401 ;
  assign y159 = ~n403 ;
  assign y160 = ~1'b0 ;
  assign y161 = ~n404 ;
  assign y162 = ~n411 ;
  assign y163 = ~1'b0 ;
  assign y164 = n412 ;
  assign y165 = n419 ;
  assign y166 = ~n423 ;
  assign y167 = n425 ;
  assign y168 = n434 ;
  assign y169 = ~1'b0 ;
  assign y170 = n438 ;
  assign y171 = ~n445 ;
  assign y172 = ~n448 ;
  assign y173 = ~1'b0 ;
  assign y174 = ~1'b0 ;
  assign y175 = ~n450 ;
  assign y176 = ~n451 ;
  assign y177 = ~n452 ;
  assign y178 = n453 ;
  assign y179 = ~n454 ;
  assign y180 = ~1'b0 ;
  assign y181 = ~n456 ;
  assign y182 = ~n461 ;
  assign y183 = ~n466 ;
  assign y184 = ~1'b0 ;
  assign y185 = ~1'b0 ;
  assign y186 = ~n468 ;
  assign y187 = ~1'b0 ;
  assign y188 = n470 ;
  assign y189 = n472 ;
  assign y190 = n477 ;
  assign y191 = n479 ;
  assign y192 = n482 ;
  assign y193 = n484 ;
  assign y194 = n488 ;
  assign y195 = ~1'b0 ;
  assign y196 = n451 ;
  assign y197 = n489 ;
  assign y198 = n493 ;
  assign y199 = ~n495 ;
  assign y200 = n502 ;
  assign y201 = n505 ;
  assign y202 = ~1'b0 ;
  assign y203 = ~n506 ;
  assign y204 = ~n508 ;
  assign y205 = ~n188 ;
  assign y206 = ~n510 ;
  assign y207 = n517 ;
  assign y208 = n521 ;
  assign y209 = ~1'b0 ;
  assign y210 = ~n523 ;
  assign y211 = n525 ;
  assign y212 = n527 ;
  assign y213 = n528 ;
  assign y214 = n533 ;
  assign y215 = ~n31 ;
  assign y216 = n535 ;
  assign y217 = ~1'b0 ;
  assign y218 = 1'b0 ;
  assign y219 = n542 ;
  assign y220 = n543 ;
  assign y221 = n545 ;
  assign y222 = n547 ;
  assign y223 = n549 ;
  assign y224 = ~n553 ;
  assign y225 = ~1'b0 ;
  assign y226 = ~1'b0 ;
  assign y227 = ~n316 ;
  assign y228 = ~1'b0 ;
  assign y229 = n560 ;
  assign y230 = ~n563 ;
  assign y231 = ~n571 ;
  assign y232 = n574 ;
  assign y233 = ~n582 ;
  assign y234 = ~1'b0 ;
  assign y235 = ~n584 ;
  assign y236 = ~n588 ;
  assign y237 = ~1'b0 ;
  assign y238 = ~n591 ;
  assign y239 = ~1'b0 ;
  assign y240 = ~n593 ;
  assign y241 = n595 ;
  assign y242 = ~n296 ;
  assign y243 = ~1'b0 ;
  assign y244 = ~1'b0 ;
  assign y245 = ~n597 ;
  assign y246 = n598 ;
  assign y247 = n604 ;
  assign y248 = ~1'b0 ;
  assign y249 = ~n607 ;
  assign y250 = ~n582 ;
  assign y251 = n608 ;
  assign y252 = ~1'b0 ;
  assign y253 = n220 ;
  assign y254 = ~n609 ;
  assign y255 = n612 ;
  assign y256 = ~1'b0 ;
  assign y257 = ~n592 ;
  assign y258 = ~n614 ;
  assign y259 = n615 ;
  assign y260 = ~n617 ;
  assign y261 = ~n622 ;
  assign y262 = n625 ;
  assign y263 = n466 ;
  assign y264 = ~n627 ;
  assign y265 = ~n634 ;
  assign y266 = n635 ;
  assign y267 = ~1'b0 ;
  assign y268 = n637 ;
  assign y269 = ~n641 ;
  assign y270 = ~x11 ;
  assign y271 = n340 ;
  assign y272 = n647 ;
  assign y273 = n652 ;
  assign y274 = ~1'b0 ;
  assign y275 = ~1'b0 ;
  assign y276 = ~n659 ;
  assign y277 = ~n667 ;
  assign y278 = ~1'b0 ;
  assign y279 = ~n671 ;
  assign y280 = ~1'b0 ;
  assign y281 = n675 ;
  assign y282 = ~1'b0 ;
  assign y283 = n677 ;
  assign y284 = ~1'b0 ;
  assign y285 = ~n682 ;
  assign y286 = ~n683 ;
  assign y287 = n687 ;
  assign y288 = n694 ;
  assign y289 = n696 ;
  assign y290 = ~n698 ;
  assign y291 = n701 ;
  assign y292 = n703 ;
  assign y293 = n704 ;
  assign y294 = ~1'b0 ;
  assign y295 = n706 ;
  assign y296 = n708 ;
  assign y297 = n710 ;
  assign y298 = n716 ;
  assign y299 = ~1'b0 ;
  assign y300 = ~n717 ;
  assign y301 = n721 ;
  assign y302 = ~n584 ;
  assign y303 = ~n510 ;
  assign y304 = 1'b0 ;
  assign y305 = ~n727 ;
  assign y306 = n729 ;
  assign y307 = 1'b0 ;
  assign y308 = ~n732 ;
  assign y309 = n734 ;
  assign y310 = ~n135 ;
  assign y311 = 1'b0 ;
  assign y312 = n736 ;
  assign y313 = ~n740 ;
  assign y314 = ~n741 ;
  assign y315 = n742 ;
  assign y316 = n745 ;
  assign y317 = n625 ;
  assign y318 = ~1'b0 ;
  assign y319 = ~1'b0 ;
  assign y320 = ~n747 ;
  assign y321 = ~n751 ;
  assign y322 = ~n752 ;
  assign y323 = ~1'b0 ;
  assign y324 = ~n753 ;
  assign y325 = n758 ;
  assign y326 = n764 ;
  assign y327 = ~1'b0 ;
  assign y328 = n766 ;
  assign y329 = ~n768 ;
  assign y330 = ~n770 ;
  assign y331 = ~1'b0 ;
  assign y332 = ~n773 ;
  assign y333 = ~n777 ;
  assign y334 = ~n778 ;
  assign y335 = ~n749 ;
  assign y336 = ~n780 ;
  assign y337 = n781 ;
  assign y338 = n786 ;
  assign y339 = ~n787 ;
  assign y340 = n790 ;
  assign y341 = ~n792 ;
  assign y342 = ~n225 ;
  assign y343 = ~n798 ;
  assign y344 = ~1'b0 ;
  assign y345 = ~n805 ;
  assign y346 = n806 ;
  assign y347 = ~1'b0 ;
  assign y348 = ~n808 ;
  assign y349 = n819 ;
  assign y350 = n820 ;
  assign y351 = ~1'b0 ;
  assign y352 = ~1'b0 ;
  assign y353 = ~1'b0 ;
  assign y354 = ~1'b0 ;
  assign y355 = ~1'b0 ;
  assign y356 = n821 ;
  assign y357 = ~1'b0 ;
  assign y358 = ~n825 ;
  assign y359 = ~1'b0 ;
  assign y360 = ~1'b0 ;
  assign y361 = ~1'b0 ;
  assign y362 = n827 ;
  assign y363 = n828 ;
  assign y364 = 1'b0 ;
  assign y365 = n829 ;
  assign y366 = ~n831 ;
  assign y367 = ~n832 ;
  assign y368 = n833 ;
  assign y369 = ~n840 ;
  assign y370 = n841 ;
  assign y371 = ~1'b0 ;
  assign y372 = ~n844 ;
  assign y373 = ~1'b0 ;
  assign y374 = ~n846 ;
  assign y375 = ~1'b0 ;
  assign y376 = ~1'b0 ;
  assign y377 = ~n850 ;
  assign y378 = ~1'b0 ;
  assign y379 = ~1'b0 ;
  assign y380 = 1'b0 ;
  assign y381 = ~n851 ;
  assign y382 = ~1'b0 ;
  assign y383 = ~1'b0 ;
  assign y384 = ~n854 ;
  assign y385 = ~n860 ;
  assign y386 = ~1'b0 ;
  assign y387 = n861 ;
  assign y388 = ~1'b0 ;
  assign y389 = n862 ;
  assign y390 = ~n864 ;
  assign y391 = ~n304 ;
  assign y392 = ~1'b0 ;
  assign y393 = ~1'b0 ;
  assign y394 = ~1'b0 ;
  assign y395 = ~n867 ;
  assign y396 = n875 ;
  assign y397 = n877 ;
  assign y398 = ~n878 ;
  assign y399 = ~1'b0 ;
  assign y400 = ~n880 ;
  assign y401 = 1'b0 ;
  assign y402 = n884 ;
  assign y403 = n886 ;
  assign y404 = ~n890 ;
  assign y405 = ~n891 ;
  assign y406 = ~n896 ;
  assign y407 = n209 ;
  assign y408 = ~n796 ;
  assign y409 = ~n901 ;
  assign y410 = ~1'b0 ;
  assign y411 = n904 ;
  assign y412 = ~n907 ;
  assign y413 = ~1'b0 ;
  assign y414 = ~n911 ;
  assign y415 = ~1'b0 ;
  assign y416 = ~n915 ;
  assign y417 = n379 ;
  assign y418 = ~1'b0 ;
  assign y419 = ~n917 ;
  assign y420 = n920 ;
  assign y421 = ~n922 ;
  assign y422 = ~1'b0 ;
  assign y423 = ~n927 ;
  assign y424 = n929 ;
  assign y425 = n932 ;
  assign y426 = ~n938 ;
  assign y427 = ~1'b0 ;
  assign y428 = ~1'b0 ;
  assign y429 = ~1'b0 ;
  assign y430 = n404 ;
  assign y431 = n949 ;
  assign y432 = 1'b0 ;
  assign y433 = n950 ;
  assign y434 = 1'b0 ;
  assign y435 = ~1'b0 ;
  assign y436 = n954 ;
  assign y437 = ~n959 ;
  assign y438 = ~n965 ;
  assign y439 = ~n717 ;
  assign y440 = n967 ;
  assign y441 = ~n968 ;
  assign y442 = n277 ;
  assign y443 = ~1'b0 ;
  assign y444 = n972 ;
  assign y445 = ~1'b0 ;
  assign y446 = ~n560 ;
  assign y447 = n974 ;
  assign y448 = ~1'b0 ;
  assign y449 = n975 ;
  assign y450 = ~n976 ;
  assign y451 = ~1'b0 ;
  assign y452 = n984 ;
  assign y453 = n985 ;
  assign y454 = ~1'b0 ;
  assign y455 = ~n988 ;
  assign y456 = ~1'b0 ;
  assign y457 = ~n989 ;
  assign y458 = ~n993 ;
  assign y459 = n998 ;
  assign y460 = ~n1000 ;
  assign y461 = ~n1003 ;
  assign y462 = n1004 ;
  assign y463 = n1007 ;
  assign y464 = ~1'b0 ;
  assign y465 = n1010 ;
  assign y466 = n1021 ;
  assign y467 = ~n1024 ;
  assign y468 = n1025 ;
  assign y469 = ~n1029 ;
  assign y470 = ~1'b0 ;
  assign y471 = n1032 ;
  assign y472 = n1038 ;
  assign y473 = ~n1040 ;
  assign y474 = ~n1042 ;
  assign y475 = n1056 ;
  assign y476 = ~n1057 ;
  assign y477 = 1'b0 ;
  assign y478 = ~1'b0 ;
  assign y479 = ~1'b0 ;
  assign y480 = n1063 ;
  assign y481 = n1065 ;
  assign y482 = ~n841 ;
  assign y483 = ~n737 ;
  assign y484 = ~1'b0 ;
  assign y485 = ~1'b0 ;
  assign y486 = ~n1066 ;
  assign y487 = n1071 ;
  assign y488 = ~n1073 ;
  assign y489 = ~n1077 ;
  assign y490 = n1078 ;
  assign y491 = n305 ;
  assign y492 = ~n1083 ;
  assign y493 = ~n1085 ;
  assign y494 = ~n1087 ;
  assign y495 = ~1'b0 ;
  assign y496 = ~n1089 ;
  assign y497 = ~1'b0 ;
  assign y498 = ~1'b0 ;
  assign y499 = n1090 ;
  assign y500 = n1094 ;
  assign y501 = ~n1095 ;
  assign y502 = ~1'b0 ;
  assign y503 = n1104 ;
  assign y504 = n1105 ;
  assign y505 = ~n1111 ;
  assign y506 = n619 ;
  assign y507 = n1114 ;
  assign y508 = ~1'b0 ;
  assign y509 = n1116 ;
  assign y510 = n1118 ;
  assign y511 = ~1'b0 ;
  assign y512 = ~1'b0 ;
  assign y513 = ~1'b0 ;
  assign y514 = ~n263 ;
  assign y515 = n1121 ;
  assign y516 = ~n1123 ;
  assign y517 = ~n286 ;
  assign y518 = n220 ;
  assign y519 = n1124 ;
  assign y520 = n1128 ;
  assign y521 = n1130 ;
  assign y522 = ~n1131 ;
  assign y523 = n1134 ;
  assign y524 = ~n1136 ;
  assign y525 = n1141 ;
  assign y526 = n1144 ;
  assign y527 = 1'b0 ;
  assign y528 = ~n1145 ;
  assign y529 = n1154 ;
  assign y530 = ~1'b0 ;
  assign y531 = n253 ;
  assign y532 = n1157 ;
  assign y533 = n1161 ;
  assign y534 = ~1'b0 ;
  assign y535 = n1165 ;
  assign y536 = ~n1167 ;
  assign y537 = ~1'b0 ;
  assign y538 = ~n1173 ;
  assign y539 = ~1'b0 ;
  assign y540 = ~n1177 ;
  assign y541 = ~1'b0 ;
  assign y542 = n1179 ;
  assign y543 = ~n1186 ;
  assign y544 = ~1'b0 ;
  assign y545 = n1190 ;
  assign y546 = n1192 ;
  assign y547 = ~n1196 ;
  assign y548 = ~1'b0 ;
  assign y549 = ~n1199 ;
  assign y550 = n182 ;
  assign y551 = ~1'b0 ;
  assign y552 = ~n1210 ;
  assign y553 = n1211 ;
  assign y554 = n1213 ;
  assign y555 = ~n1215 ;
  assign y556 = ~1'b0 ;
  assign y557 = ~1'b0 ;
  assign y558 = n1216 ;
  assign y559 = n488 ;
  assign y560 = ~1'b0 ;
  assign y561 = ~1'b0 ;
  assign y562 = ~1'b0 ;
  assign y563 = n1226 ;
  assign y564 = n1227 ;
  assign y565 = n1230 ;
  assign y566 = ~n1231 ;
  assign y567 = n1234 ;
  assign y568 = ~1'b0 ;
  assign y569 = ~n1237 ;
  assign y570 = ~n1238 ;
  assign y571 = ~n1241 ;
  assign y572 = n1243 ;
  assign y573 = ~n1245 ;
  assign y574 = ~n1247 ;
  assign y575 = ~1'b0 ;
  assign y576 = ~n1251 ;
  assign y577 = n1254 ;
  assign y578 = ~1'b0 ;
  assign y579 = ~n1261 ;
  assign y580 = n1264 ;
  assign y581 = n1266 ;
  assign y582 = ~n1267 ;
  assign y583 = ~n1269 ;
  assign y584 = 1'b0 ;
  assign y585 = ~1'b0 ;
  assign y586 = ~1'b0 ;
  assign y587 = ~n1271 ;
  assign y588 = n1276 ;
  assign y589 = ~1'b0 ;
  assign y590 = n1283 ;
  assign y591 = ~n1284 ;
  assign y592 = ~n481 ;
  assign y593 = ~n1291 ;
  assign y594 = n1297 ;
  assign y595 = ~n1299 ;
  assign y596 = ~1'b0 ;
  assign y597 = n1300 ;
  assign y598 = ~1'b0 ;
  assign y599 = ~1'b0 ;
  assign y600 = n1301 ;
  assign y601 = 1'b0 ;
  assign y602 = ~n1305 ;
  assign y603 = n1307 ;
  assign y604 = n1308 ;
  assign y605 = n1310 ;
  assign y606 = n1313 ;
  assign y607 = ~n1315 ;
  assign y608 = n1316 ;
  assign y609 = n1320 ;
  assign y610 = n1321 ;
  assign y611 = 1'b0 ;
  assign y612 = n905 ;
  assign y613 = n1322 ;
  assign y614 = ~n1323 ;
  assign y615 = n270 ;
  assign y616 = n1326 ;
  assign y617 = ~n1329 ;
  assign y618 = ~1'b0 ;
  assign y619 = ~1'b0 ;
  assign y620 = ~1'b0 ;
  assign y621 = ~1'b0 ;
  assign y622 = ~1'b0 ;
  assign y623 = ~n1331 ;
  assign y624 = ~1'b0 ;
  assign y625 = n1335 ;
  assign y626 = n1337 ;
  assign y627 = n1340 ;
  assign y628 = ~n1342 ;
  assign y629 = ~n1344 ;
  assign y630 = n1345 ;
  assign y631 = ~n1346 ;
  assign y632 = ~1'b0 ;
  assign y633 = ~1'b0 ;
  assign y634 = ~n1349 ;
  assign y635 = ~1'b0 ;
  assign y636 = n1352 ;
  assign y637 = ~n1353 ;
  assign y638 = n1355 ;
  assign y639 = n1360 ;
  assign y640 = ~n1361 ;
  assign y641 = ~1'b0 ;
  assign y642 = ~1'b0 ;
  assign y643 = n1365 ;
  assign y644 = ~1'b0 ;
  assign y645 = ~1'b0 ;
  assign y646 = n1370 ;
  assign y647 = ~n1372 ;
  assign y648 = ~n1377 ;
  assign y649 = n1379 ;
  assign y650 = ~n1381 ;
  assign y651 = ~1'b0 ;
  assign y652 = ~1'b0 ;
  assign y653 = ~1'b0 ;
  assign y654 = ~n1385 ;
  assign y655 = ~1'b0 ;
  assign y656 = ~n1386 ;
  assign y657 = ~n1390 ;
  assign y658 = ~1'b0 ;
  assign y659 = ~n1395 ;
  assign y660 = ~1'b0 ;
  assign y661 = ~n1312 ;
  assign y662 = 1'b0 ;
  assign y663 = ~n1398 ;
  assign y664 = n1400 ;
  assign y665 = ~n1403 ;
  assign y666 = n1409 ;
  assign y667 = n1410 ;
  assign y668 = ~n1411 ;
  assign y669 = ~1'b0 ;
  assign y670 = ~n1418 ;
  assign y671 = n924 ;
  assign y672 = ~n1419 ;
  assign y673 = ~1'b0 ;
  assign y674 = ~n1424 ;
  assign y675 = ~1'b0 ;
  assign y676 = ~n1426 ;
  assign y677 = ~1'b0 ;
  assign y678 = ~1'b0 ;
  assign y679 = n1428 ;
  assign y680 = ~n1430 ;
  assign y681 = ~1'b0 ;
  assign y682 = n1435 ;
  assign y683 = ~n140 ;
  assign y684 = ~1'b0 ;
  assign y685 = ~1'b0 ;
  assign y686 = ~n1437 ;
  assign y687 = n1398 ;
  assign y688 = ~1'b0 ;
  assign y689 = n1439 ;
  assign y690 = ~n1442 ;
  assign y691 = ~1'b0 ;
  assign y692 = n798 ;
  assign y693 = ~n1445 ;
  assign y694 = n1451 ;
  assign y695 = 1'b0 ;
  assign y696 = ~1'b0 ;
  assign y697 = n1453 ;
  assign y698 = ~1'b0 ;
  assign y699 = ~n1454 ;
  assign y700 = ~1'b0 ;
  assign y701 = ~n1461 ;
  assign y702 = n1462 ;
  assign y703 = ~n1469 ;
  assign y704 = n372 ;
  assign y705 = ~1'b0 ;
  assign y706 = ~1'b0 ;
  assign y707 = n1481 ;
  assign y708 = ~1'b0 ;
  assign y709 = n1484 ;
  assign y710 = n1485 ;
  assign y711 = n105 ;
  assign y712 = ~1'b0 ;
  assign y713 = ~n1208 ;
  assign y714 = n733 ;
  assign y715 = ~1'b0 ;
  assign y716 = ~n1491 ;
  assign y717 = ~1'b0 ;
  assign y718 = ~n982 ;
  assign y719 = n1215 ;
  assign y720 = n1497 ;
  assign y721 = ~n1499 ;
  assign y722 = ~n1501 ;
  assign y723 = n1502 ;
  assign y724 = ~1'b0 ;
  assign y725 = ~1'b0 ;
  assign y726 = 1'b0 ;
  assign y727 = n1504 ;
  assign y728 = n1505 ;
  assign y729 = ~1'b0 ;
  assign y730 = ~n1506 ;
  assign y731 = n225 ;
  assign y732 = n1507 ;
  assign y733 = ~n1511 ;
  assign y734 = n1513 ;
  assign y735 = ~n1514 ;
  assign y736 = n1516 ;
  assign y737 = ~n1517 ;
  assign y738 = ~n1520 ;
  assign y739 = ~n1522 ;
  assign y740 = n1525 ;
  assign y741 = ~1'b0 ;
  assign y742 = n1528 ;
  assign y743 = ~n1531 ;
  assign y744 = ~1'b0 ;
  assign y745 = ~1'b0 ;
  assign y746 = ~n1535 ;
  assign y747 = ~n1538 ;
  assign y748 = ~1'b0 ;
  assign y749 = ~n1539 ;
  assign y750 = n1548 ;
  assign y751 = ~n1398 ;
  assign y752 = ~1'b0 ;
  assign y753 = n1552 ;
  assign y754 = ~1'b0 ;
  assign y755 = ~1'b0 ;
  assign y756 = n846 ;
  assign y757 = 1'b0 ;
  assign y758 = ~n1560 ;
  assign y759 = n1561 ;
  assign y760 = ~n1563 ;
  assign y761 = ~n1567 ;
  assign y762 = ~1'b0 ;
  assign y763 = ~1'b0 ;
  assign y764 = ~n1542 ;
  assign y765 = ~n1573 ;
  assign y766 = ~1'b0 ;
  assign y767 = n1576 ;
  assign y768 = n1578 ;
  assign y769 = n1591 ;
  assign y770 = ~1'b0 ;
  assign y771 = ~n1594 ;
  assign y772 = ~1'b0 ;
  assign y773 = ~1'b0 ;
  assign y774 = ~1'b0 ;
  assign y775 = ~1'b0 ;
  assign y776 = ~n1598 ;
  assign y777 = ~n1599 ;
  assign y778 = n1603 ;
  assign y779 = n1605 ;
  assign y780 = ~1'b0 ;
  assign y781 = n1608 ;
  assign y782 = ~n1609 ;
  assign y783 = ~1'b0 ;
  assign y784 = ~n1611 ;
  assign y785 = ~1'b0 ;
  assign y786 = n1618 ;
  assign y787 = n1620 ;
  assign y788 = ~1'b0 ;
  assign y789 = ~n997 ;
  assign y790 = ~n1624 ;
  assign y791 = n1625 ;
  assign y792 = ~n1627 ;
  assign y793 = ~1'b0 ;
  assign y794 = ~n1629 ;
  assign y795 = n1631 ;
  assign y796 = n1635 ;
  assign y797 = ~1'b0 ;
  assign y798 = n1636 ;
  assign y799 = ~1'b0 ;
  assign y800 = n1637 ;
  assign y801 = n1649 ;
  assign y802 = ~n1650 ;
  assign y803 = n1653 ;
  assign y804 = 1'b0 ;
  assign y805 = n1654 ;
  assign y806 = ~n1655 ;
  assign y807 = ~1'b0 ;
  assign y808 = ~n1656 ;
  assign y809 = ~n1657 ;
  assign y810 = ~1'b0 ;
  assign y811 = n1658 ;
  assign y812 = n1663 ;
  assign y813 = ~n1664 ;
  assign y814 = ~1'b0 ;
  assign y815 = ~n1672 ;
  assign y816 = ~1'b0 ;
  assign y817 = n1439 ;
  assign y818 = ~1'b0 ;
  assign y819 = ~n1674 ;
  assign y820 = ~1'b0 ;
  assign y821 = ~n1684 ;
  assign y822 = n344 ;
  assign y823 = n1689 ;
  assign y824 = n1690 ;
  assign y825 = ~n1691 ;
  assign y826 = n1699 ;
  assign y827 = ~n1700 ;
  assign y828 = n1701 ;
  assign y829 = ~n1703 ;
  assign y830 = n1715 ;
  assign y831 = ~n1716 ;
  assign y832 = ~1'b0 ;
  assign y833 = ~n1720 ;
  assign y834 = ~1'b0 ;
  assign y835 = n1721 ;
  assign y836 = ~n1728 ;
  assign y837 = ~n1385 ;
  assign y838 = n1729 ;
  assign y839 = n1739 ;
  assign y840 = ~1'b0 ;
  assign y841 = ~1'b0 ;
  assign y842 = ~1'b0 ;
  assign y843 = ~n1741 ;
  assign y844 = ~1'b0 ;
  assign y845 = n1743 ;
  assign y846 = ~n1749 ;
  assign y847 = n395 ;
  assign y848 = n1752 ;
  assign y849 = ~n1758 ;
  assign y850 = n1760 ;
  assign y851 = ~n1764 ;
  assign y852 = ~n1765 ;
  assign y853 = ~1'b0 ;
  assign y854 = n1769 ;
  assign y855 = ~n1771 ;
  assign y856 = ~n1775 ;
  assign y857 = ~n1779 ;
  assign y858 = ~1'b0 ;
  assign y859 = ~n1781 ;
  assign y860 = ~n1783 ;
  assign y861 = ~1'b0 ;
  assign y862 = ~n1788 ;
  assign y863 = n1353 ;
  assign y864 = n1791 ;
  assign y865 = ~1'b0 ;
  assign y866 = ~n1792 ;
  assign y867 = ~1'b0 ;
  assign y868 = n1800 ;
  assign y869 = n1802 ;
  assign y870 = n1804 ;
  assign y871 = ~n1808 ;
  assign y872 = n1809 ;
  assign y873 = ~1'b0 ;
  assign y874 = ~1'b0 ;
  assign y875 = ~1'b0 ;
  assign y876 = ~n1811 ;
  assign y877 = n1814 ;
  assign y878 = ~n1469 ;
  assign y879 = n1816 ;
  assign y880 = ~n1819 ;
  assign y881 = n1823 ;
  assign y882 = n1829 ;
  assign y883 = ~n1830 ;
  assign y884 = ~n1832 ;
  assign y885 = n1834 ;
  assign y886 = ~1'b0 ;
  assign y887 = ~n1835 ;
  assign y888 = ~1'b0 ;
  assign y889 = ~n1837 ;
  assign y890 = ~n1838 ;
  assign y891 = n1841 ;
  assign y892 = ~n1842 ;
  assign y893 = ~n1845 ;
  assign y894 = 1'b0 ;
  assign y895 = ~n1848 ;
  assign y896 = n1849 ;
  assign y897 = ~1'b0 ;
  assign y898 = ~1'b0 ;
  assign y899 = ~1'b0 ;
  assign y900 = ~n1851 ;
  assign y901 = ~n1858 ;
  assign y902 = n1863 ;
  assign y903 = ~1'b0 ;
  assign y904 = ~n1872 ;
  assign y905 = ~1'b0 ;
  assign y906 = 1'b0 ;
  assign y907 = ~n1875 ;
  assign y908 = n1876 ;
  assign y909 = n1882 ;
  assign y910 = ~n1883 ;
  assign y911 = ~1'b0 ;
  assign y912 = n1884 ;
  assign y913 = ~n1892 ;
  assign y914 = ~n1893 ;
  assign y915 = ~1'b0 ;
  assign y916 = ~1'b0 ;
  assign y917 = ~n1896 ;
  assign y918 = 1'b0 ;
  assign y919 = n1902 ;
  assign y920 = ~n1510 ;
  assign y921 = ~1'b0 ;
  assign y922 = ~1'b0 ;
  assign y923 = ~1'b0 ;
  assign y924 = ~n1907 ;
  assign y925 = n1910 ;
  assign y926 = ~n1911 ;
  assign y927 = ~n208 ;
  assign y928 = n1915 ;
  assign y929 = ~1'b0 ;
  assign y930 = ~n1918 ;
  assign y931 = ~1'b0 ;
  assign y932 = ~n831 ;
  assign y933 = ~1'b0 ;
  assign y934 = n1921 ;
  assign y935 = ~1'b0 ;
  assign y936 = n1329 ;
  assign y937 = ~n1924 ;
  assign y938 = ~n1925 ;
  assign y939 = ~1'b0 ;
  assign y940 = n1929 ;
  assign y941 = ~n1932 ;
  assign y942 = ~n1935 ;
  assign y943 = n996 ;
  assign y944 = ~1'b0 ;
  assign y945 = ~1'b0 ;
  assign y946 = n209 ;
  assign y947 = n1941 ;
  assign y948 = ~n1945 ;
  assign y949 = n1947 ;
  assign y950 = ~n1949 ;
  assign y951 = ~1'b0 ;
  assign y952 = ~n1958 ;
  assign y953 = ~1'b0 ;
  assign y954 = ~n1966 ;
  assign y955 = ~1'b0 ;
  assign y956 = 1'b0 ;
  assign y957 = n1968 ;
  assign y958 = ~1'b0 ;
  assign y959 = ~n1973 ;
  assign y960 = ~n1976 ;
  assign y961 = n1980 ;
  assign y962 = n1981 ;
  assign y963 = ~n1985 ;
  assign y964 = ~1'b0 ;
  assign y965 = ~n1986 ;
  assign y966 = ~n1987 ;
  assign y967 = n1988 ;
  assign y968 = n1989 ;
  assign y969 = ~n1993 ;
  assign y970 = ~1'b0 ;
  assign y971 = ~n1999 ;
  assign y972 = ~1'b0 ;
  assign y973 = ~1'b0 ;
  assign y974 = n1010 ;
  assign y975 = ~n2002 ;
  assign y976 = n2007 ;
  assign y977 = ~1'b0 ;
  assign y978 = ~1'b0 ;
  assign y979 = ~n2008 ;
  assign y980 = ~n2010 ;
  assign y981 = ~n2017 ;
  assign y982 = ~n2019 ;
  assign y983 = ~1'b0 ;
  assign y984 = ~n2022 ;
  assign y985 = ~1'b0 ;
  assign y986 = n2023 ;
  assign y987 = ~1'b0 ;
  assign y988 = n2024 ;
  assign y989 = ~n2030 ;
  assign y990 = ~n2032 ;
  assign y991 = n2033 ;
  assign y992 = ~n2034 ;
  assign y993 = ~n2039 ;
  assign y994 = ~n2041 ;
  assign y995 = n2044 ;
  assign y996 = ~1'b0 ;
  assign y997 = n2045 ;
  assign y998 = ~n2046 ;
  assign y999 = ~n2048 ;
  assign y1000 = ~1'b0 ;
  assign y1001 = ~n1584 ;
  assign y1002 = 1'b0 ;
  assign y1003 = ~n2050 ;
  assign y1004 = n2055 ;
  assign y1005 = ~1'b0 ;
  assign y1006 = ~1'b0 ;
  assign y1007 = 1'b0 ;
  assign y1008 = ~n2060 ;
  assign y1009 = n2061 ;
  assign y1010 = ~1'b0 ;
  assign y1011 = n2063 ;
  assign y1012 = n2066 ;
  assign y1013 = n2077 ;
  assign y1014 = n2080 ;
  assign y1015 = n2085 ;
  assign y1016 = n2087 ;
  assign y1017 = n2091 ;
  assign y1018 = ~1'b0 ;
  assign y1019 = n2093 ;
  assign y1020 = ~1'b0 ;
  assign y1021 = ~n2094 ;
  assign y1022 = n2098 ;
  assign y1023 = n2102 ;
  assign y1024 = ~1'b0 ;
  assign y1025 = ~n2103 ;
  assign y1026 = n2106 ;
  assign y1027 = n2108 ;
  assign y1028 = ~n1080 ;
  assign y1029 = ~1'b0 ;
  assign y1030 = ~n2109 ;
  assign y1031 = ~n2110 ;
  assign y1032 = ~1'b0 ;
  assign y1033 = ~1'b0 ;
  assign y1034 = ~n2112 ;
  assign y1035 = n2116 ;
  assign y1036 = n261 ;
  assign y1037 = ~1'b0 ;
  assign y1038 = n2120 ;
  assign y1039 = n2127 ;
  assign y1040 = n2128 ;
  assign y1041 = n2129 ;
  assign y1042 = ~1'b0 ;
  assign y1043 = ~n2097 ;
  assign y1044 = n390 ;
  assign y1045 = ~n2134 ;
  assign y1046 = ~1'b0 ;
  assign y1047 = ~n2136 ;
  assign y1048 = ~1'b0 ;
  assign y1049 = n2138 ;
  assign y1050 = ~1'b0 ;
  assign y1051 = ~n826 ;
  assign y1052 = n2141 ;
  assign y1053 = ~1'b0 ;
  assign y1054 = n2145 ;
  assign y1055 = ~1'b0 ;
  assign y1056 = ~1'b0 ;
  assign y1057 = n2146 ;
  assign y1058 = ~1'b0 ;
  assign y1059 = n2148 ;
  assign y1060 = n2154 ;
  assign y1061 = ~1'b0 ;
  assign y1062 = n2155 ;
  assign y1063 = ~n2157 ;
  assign y1064 = ~1'b0 ;
  assign y1065 = ~1'b0 ;
  assign y1066 = n2158 ;
  assign y1067 = ~n291 ;
  assign y1068 = n2159 ;
  assign y1069 = ~1'b0 ;
  assign y1070 = ~n468 ;
  assign y1071 = ~x5 ;
  assign y1072 = ~1'b0 ;
  assign y1073 = ~n2168 ;
  assign y1074 = ~n2170 ;
  assign y1075 = ~n2175 ;
  assign y1076 = ~1'b0 ;
  assign y1077 = n2176 ;
  assign y1078 = ~n2184 ;
  assign y1079 = ~1'b0 ;
  assign y1080 = ~1'b0 ;
  assign y1081 = ~1'b0 ;
  assign y1082 = n2186 ;
  assign y1083 = ~1'b0 ;
  assign y1084 = ~n2195 ;
  assign y1085 = n2203 ;
  assign y1086 = ~n1460 ;
  assign y1087 = n1264 ;
  assign y1088 = ~n423 ;
  assign y1089 = ~1'b0 ;
  assign y1090 = ~1'b0 ;
  assign y1091 = ~n2204 ;
  assign y1092 = ~1'b0 ;
  assign y1093 = n2207 ;
  assign y1094 = ~1'b0 ;
  assign y1095 = ~n2210 ;
  assign y1096 = n2211 ;
  assign y1097 = n2212 ;
  assign y1098 = ~n2214 ;
  assign y1099 = ~1'b0 ;
  assign y1100 = ~n2217 ;
  assign y1101 = ~1'b0 ;
  assign y1102 = ~n2223 ;
  assign y1103 = ~n2227 ;
  assign y1104 = n2229 ;
  assign y1105 = n2230 ;
  assign y1106 = n2231 ;
  assign y1107 = n2233 ;
  assign y1108 = ~n2235 ;
  assign y1109 = ~n2240 ;
  assign y1110 = ~1'b0 ;
  assign y1111 = ~n2244 ;
  assign y1112 = ~1'b0 ;
  assign y1113 = n2246 ;
  assign y1114 = n2247 ;
  assign y1115 = ~1'b0 ;
  assign y1116 = ~n2250 ;
  assign y1117 = ~1'b0 ;
  assign y1118 = 1'b0 ;
  assign y1119 = n2252 ;
  assign y1120 = ~1'b0 ;
  assign y1121 = ~n2253 ;
  assign y1122 = n2256 ;
  assign y1123 = n2261 ;
  assign y1124 = ~1'b0 ;
  assign y1125 = ~n2265 ;
  assign y1126 = n2270 ;
  assign y1127 = ~1'b0 ;
  assign y1128 = ~n2279 ;
  assign y1129 = ~n1066 ;
  assign y1130 = ~1'b0 ;
  assign y1131 = n2286 ;
  assign y1132 = ~n2288 ;
  assign y1133 = ~1'b0 ;
  assign y1134 = ~n2291 ;
  assign y1135 = n2308 ;
  assign y1136 = ~1'b0 ;
  assign y1137 = n2309 ;
  assign y1138 = ~n2311 ;
  assign y1139 = ~1'b0 ;
  assign y1140 = n2313 ;
  assign y1141 = ~n2316 ;
  assign y1142 = ~1'b0 ;
  assign y1143 = n2319 ;
  assign y1144 = ~1'b0 ;
  assign y1145 = ~n2320 ;
  assign y1146 = ~1'b0 ;
  assign y1147 = n2321 ;
  assign y1148 = n2328 ;
  assign y1149 = n2331 ;
  assign y1150 = ~1'b0 ;
  assign y1151 = ~n2334 ;
  assign y1152 = ~1'b0 ;
  assign y1153 = n2335 ;
  assign y1154 = n2336 ;
  assign y1155 = ~1'b0 ;
  assign y1156 = ~n2340 ;
  assign y1157 = ~1'b0 ;
  assign y1158 = n2341 ;
  assign y1159 = ~n1941 ;
  assign y1160 = ~1'b0 ;
  assign y1161 = ~1'b0 ;
  assign y1162 = ~1'b0 ;
  assign y1163 = n2349 ;
  assign y1164 = ~1'b0 ;
  assign y1165 = n2351 ;
  assign y1166 = n2353 ;
  assign y1167 = ~1'b0 ;
  assign y1168 = ~n2362 ;
  assign y1169 = ~1'b0 ;
  assign y1170 = n2366 ;
  assign y1171 = ~1'b0 ;
  assign y1172 = ~1'b0 ;
  assign y1173 = ~1'b0 ;
  assign y1174 = n1150 ;
  assign y1175 = ~n2367 ;
  assign y1176 = ~1'b0 ;
  assign y1177 = ~n2349 ;
  assign y1178 = n2371 ;
  assign y1179 = n2374 ;
  assign y1180 = ~n2376 ;
  assign y1181 = ~1'b0 ;
  assign y1182 = ~n2381 ;
  assign y1183 = ~n2382 ;
  assign y1184 = n2292 ;
  assign y1185 = ~1'b0 ;
  assign y1186 = ~1'b0 ;
  assign y1187 = ~1'b0 ;
  assign y1188 = 1'b0 ;
  assign y1189 = ~1'b0 ;
  assign y1190 = ~n2386 ;
  assign y1191 = n2387 ;
  assign y1192 = ~n2393 ;
  assign y1193 = ~n2399 ;
  assign y1194 = ~n2401 ;
  assign y1195 = ~1'b0 ;
  assign y1196 = ~n2406 ;
  assign y1197 = n666 ;
  assign y1198 = n2411 ;
  assign y1199 = ~n2423 ;
  assign y1200 = n2426 ;
  assign y1201 = n2428 ;
  assign y1202 = ~n2431 ;
  assign y1203 = n565 ;
  assign y1204 = 1'b0 ;
  assign y1205 = ~n1865 ;
  assign y1206 = ~1'b0 ;
  assign y1207 = ~n2433 ;
  assign y1208 = ~1'b0 ;
  assign y1209 = n2437 ;
  assign y1210 = ~1'b0 ;
  assign y1211 = n2442 ;
  assign y1212 = ~1'b0 ;
  assign y1213 = n2443 ;
  assign y1214 = ~n2446 ;
  assign y1215 = ~1'b0 ;
  assign y1216 = ~1'b0 ;
  assign y1217 = n2448 ;
  assign y1218 = ~n2451 ;
  assign y1219 = n2452 ;
  assign y1220 = n2456 ;
  assign y1221 = 1'b0 ;
  assign y1222 = ~1'b0 ;
  assign y1223 = ~1'b0 ;
  assign y1224 = ~n2458 ;
  assign y1225 = ~n854 ;
  assign y1226 = n1075 ;
  assign y1227 = n2462 ;
  assign y1228 = n2465 ;
  assign y1229 = ~n2467 ;
  assign y1230 = ~1'b0 ;
  assign y1231 = ~n2469 ;
  assign y1232 = ~1'b0 ;
  assign y1233 = ~1'b0 ;
  assign y1234 = ~1'b0 ;
  assign y1235 = ~1'b0 ;
  assign y1236 = n93 ;
  assign y1237 = n2472 ;
  assign y1238 = ~n2474 ;
  assign y1239 = ~1'b0 ;
  assign y1240 = n968 ;
  assign y1241 = ~n2476 ;
  assign y1242 = ~n2478 ;
  assign y1243 = n2480 ;
  assign y1244 = ~1'b0 ;
  assign y1245 = 1'b0 ;
  assign y1246 = 1'b0 ;
  assign y1247 = ~1'b0 ;
  assign y1248 = ~1'b0 ;
  assign y1249 = ~n2483 ;
  assign y1250 = n2488 ;
  assign y1251 = n2489 ;
  assign y1252 = n1419 ;
  assign y1253 = ~1'b0 ;
  assign y1254 = ~n1582 ;
  assign y1255 = ~1'b0 ;
  assign y1256 = n477 ;
  assign y1257 = ~n2492 ;
  assign y1258 = n2494 ;
  assign y1259 = ~n2498 ;
  assign y1260 = ~1'b0 ;
  assign y1261 = ~n2500 ;
  assign y1262 = n2502 ;
  assign y1263 = ~1'b0 ;
  assign y1264 = ~n2504 ;
  assign y1265 = ~n2507 ;
  assign y1266 = ~n2510 ;
  assign y1267 = ~1'b0 ;
  assign y1268 = n2512 ;
  assign y1269 = ~n2513 ;
  assign y1270 = ~1'b0 ;
  assign y1271 = n2518 ;
  assign y1272 = ~n2521 ;
  assign y1273 = n2523 ;
  assign y1274 = ~1'b0 ;
  assign y1275 = ~1'b0 ;
  assign y1276 = n2531 ;
  assign y1277 = n2532 ;
  assign y1278 = ~n2535 ;
  assign y1279 = ~1'b0 ;
  assign y1280 = ~n2539 ;
  assign y1281 = ~1'b0 ;
  assign y1282 = n2543 ;
  assign y1283 = n1276 ;
  assign y1284 = ~n2547 ;
  assign y1285 = ~n2549 ;
  assign y1286 = ~n2551 ;
  assign y1287 = ~1'b0 ;
  assign y1288 = ~1'b0 ;
  assign y1289 = ~n2554 ;
  assign y1290 = n2555 ;
  assign y1291 = ~n2560 ;
  assign y1292 = ~1'b0 ;
  assign y1293 = n768 ;
  assign y1294 = n2563 ;
  assign y1295 = n2564 ;
  assign y1296 = ~1'b0 ;
  assign y1297 = ~n2566 ;
  assign y1298 = n2568 ;
  assign y1299 = ~1'b0 ;
  assign y1300 = n2569 ;
  assign y1301 = n2571 ;
  assign y1302 = n2225 ;
  assign y1303 = 1'b0 ;
  assign y1304 = n2578 ;
  assign y1305 = 1'b0 ;
  assign y1306 = ~n2581 ;
  assign y1307 = n2587 ;
  assign y1308 = ~n2588 ;
  assign y1309 = ~1'b0 ;
  assign y1310 = n2403 ;
  assign y1311 = n2593 ;
  assign y1312 = ~1'b0 ;
  assign y1313 = n1528 ;
  assign y1314 = ~n2594 ;
  assign y1315 = ~n2397 ;
  assign y1316 = ~1'b0 ;
  assign y1317 = n2595 ;
  assign y1318 = ~n2601 ;
  assign y1319 = n1254 ;
  assign y1320 = ~n2612 ;
  assign y1321 = ~n2618 ;
  assign y1322 = n2619 ;
  assign y1323 = ~1'b0 ;
  assign y1324 = ~1'b0 ;
  assign y1325 = ~1'b0 ;
  assign y1326 = ~n2623 ;
  assign y1327 = n2626 ;
  assign y1328 = ~n2627 ;
  assign y1329 = ~1'b0 ;
  assign y1330 = n2630 ;
  assign y1331 = ~1'b0 ;
  assign y1332 = ~n2634 ;
  assign y1333 = ~n2635 ;
  assign y1334 = n2637 ;
  assign y1335 = ~n2638 ;
  assign y1336 = n23 ;
  assign y1337 = n2639 ;
  assign y1338 = 1'b0 ;
  assign y1339 = n2641 ;
  assign y1340 = ~1'b0 ;
  assign y1341 = ~1'b0 ;
  assign y1342 = n2644 ;
  assign y1343 = n48 ;
  assign y1344 = ~n2647 ;
  assign y1345 = ~n2648 ;
  assign y1346 = n2649 ;
  assign y1347 = n582 ;
  assign y1348 = n2650 ;
  assign y1349 = ~1'b0 ;
  assign y1350 = ~1'b0 ;
  assign y1351 = n2653 ;
  assign y1352 = ~n2657 ;
  assign y1353 = ~1'b0 ;
  assign y1354 = n2660 ;
  assign y1355 = n2662 ;
  assign y1356 = ~1'b0 ;
  assign y1357 = n2663 ;
  assign y1358 = ~1'b0 ;
  assign y1359 = n1907 ;
  assign y1360 = ~1'b0 ;
  assign y1361 = ~1'b0 ;
  assign y1362 = ~1'b0 ;
  assign y1363 = n2665 ;
  assign y1364 = n2669 ;
  assign y1365 = ~1'b0 ;
  assign y1366 = n2670 ;
  assign y1367 = ~1'b0 ;
  assign y1368 = n2671 ;
  assign y1369 = ~n2674 ;
  assign y1370 = ~n2678 ;
  assign y1371 = ~1'b0 ;
  assign y1372 = ~n2680 ;
  assign y1373 = n2682 ;
  assign y1374 = n2684 ;
  assign y1375 = ~1'b0 ;
  assign y1376 = 1'b0 ;
  assign y1377 = n2686 ;
  assign y1378 = ~n2689 ;
  assign y1379 = ~1'b0 ;
  assign y1380 = n2693 ;
  assign y1381 = ~1'b0 ;
  assign y1382 = ~1'b0 ;
  assign y1383 = n2698 ;
  assign y1384 = n2706 ;
  assign y1385 = n2709 ;
  assign y1386 = ~1'b0 ;
  assign y1387 = ~1'b0 ;
  assign y1388 = n2711 ;
  assign y1389 = ~n2713 ;
  assign y1390 = ~1'b0 ;
  assign y1391 = ~n2716 ;
  assign y1392 = ~1'b0 ;
  assign y1393 = ~n2719 ;
  assign y1394 = n2727 ;
  assign y1395 = ~n2728 ;
  assign y1396 = ~n2733 ;
  assign y1397 = n2735 ;
  assign y1398 = ~n2736 ;
  assign y1399 = ~1'b0 ;
  assign y1400 = n2746 ;
  assign y1401 = n1392 ;
  assign y1402 = ~1'b0 ;
  assign y1403 = ~n2753 ;
  assign y1404 = n2755 ;
  assign y1405 = ~1'b0 ;
  assign y1406 = ~1'b0 ;
  assign y1407 = n2760 ;
  assign y1408 = ~n2762 ;
  assign y1409 = n2763 ;
  assign y1410 = ~n2767 ;
  assign y1411 = ~1'b0 ;
  assign y1412 = ~1'b0 ;
  assign y1413 = ~n2769 ;
  assign y1414 = ~n2770 ;
  assign y1415 = ~n2771 ;
  assign y1416 = n2772 ;
  assign y1417 = n2775 ;
  assign y1418 = ~1'b0 ;
  assign y1419 = ~n2776 ;
  assign y1420 = ~n2779 ;
  assign y1421 = 1'b0 ;
  assign y1422 = ~n2787 ;
  assign y1423 = ~n2791 ;
  assign y1424 = ~n2794 ;
  assign y1425 = ~n2802 ;
  assign y1426 = ~n2805 ;
  assign y1427 = n2807 ;
  assign y1428 = n2813 ;
  assign y1429 = ~n2815 ;
  assign y1430 = ~1'b0 ;
  assign y1431 = ~n2818 ;
  assign y1432 = ~1'b0 ;
  assign y1433 = n2821 ;
  assign y1434 = ~1'b0 ;
  assign y1435 = n2822 ;
  assign y1436 = ~n2831 ;
  assign y1437 = ~n2838 ;
  assign y1438 = ~n2843 ;
  assign y1439 = ~n2066 ;
  assign y1440 = n2845 ;
  assign y1441 = ~n2846 ;
  assign y1442 = n2847 ;
  assign y1443 = ~n2848 ;
  assign y1444 = ~1'b0 ;
  assign y1445 = ~n2849 ;
  assign y1446 = ~n2852 ;
  assign y1447 = n2854 ;
  assign y1448 = ~n2855 ;
  assign y1449 = ~n2857 ;
  assign y1450 = ~n2860 ;
  assign y1451 = ~n2862 ;
  assign y1452 = ~n2865 ;
  assign y1453 = ~n2869 ;
  assign y1454 = n2874 ;
  assign y1455 = n2875 ;
  assign y1456 = ~n2576 ;
  assign y1457 = ~1'b0 ;
  assign y1458 = ~1'b0 ;
  assign y1459 = ~1'b0 ;
  assign y1460 = n2876 ;
  assign y1461 = ~n1943 ;
  assign y1462 = ~1'b0 ;
  assign y1463 = ~1'b0 ;
  assign y1464 = ~n2891 ;
  assign y1465 = ~1'b0 ;
  assign y1466 = n2893 ;
  assign y1467 = n2899 ;
  assign y1468 = n2900 ;
  assign y1469 = ~n2901 ;
  assign y1470 = ~n2904 ;
  assign y1471 = n2905 ;
  assign y1472 = ~n2906 ;
  assign y1473 = ~1'b0 ;
  assign y1474 = n2907 ;
  assign y1475 = n2914 ;
  assign y1476 = ~n2916 ;
  assign y1477 = n2917 ;
  assign y1478 = ~1'b0 ;
  assign y1479 = ~n2919 ;
  assign y1480 = n2922 ;
  assign y1481 = ~n2923 ;
  assign y1482 = ~n2924 ;
  assign y1483 = n2925 ;
  assign y1484 = ~n2929 ;
  assign y1485 = ~n2930 ;
  assign y1486 = n2932 ;
  assign y1487 = ~n2938 ;
  assign y1488 = ~n2943 ;
  assign y1489 = ~n2948 ;
  assign y1490 = ~1'b0 ;
  assign y1491 = ~n2951 ;
  assign y1492 = n2952 ;
  assign y1493 = ~n2954 ;
  assign y1494 = ~n2955 ;
  assign y1495 = n2960 ;
  assign y1496 = ~n2966 ;
  assign y1497 = ~1'b0 ;
  assign y1498 = ~1'b0 ;
  assign y1499 = ~n2967 ;
  assign y1500 = n2976 ;
  assign y1501 = ~n959 ;
  assign y1502 = ~n2978 ;
  assign y1503 = ~1'b0 ;
  assign y1504 = ~n2981 ;
  assign y1505 = ~1'b0 ;
  assign y1506 = ~1'b0 ;
  assign y1507 = ~n2983 ;
  assign y1508 = ~1'b0 ;
  assign y1509 = n2986 ;
  assign y1510 = ~1'b0 ;
  assign y1511 = ~1'b0 ;
  assign y1512 = n2998 ;
  assign y1513 = ~1'b0 ;
  assign y1514 = ~1'b0 ;
  assign y1515 = n3003 ;
  assign y1516 = ~n3008 ;
  assign y1517 = n3012 ;
  assign y1518 = n3013 ;
  assign y1519 = ~n3017 ;
  assign y1520 = ~n788 ;
  assign y1521 = ~n3020 ;
  assign y1522 = ~1'b0 ;
  assign y1523 = ~n3025 ;
  assign y1524 = ~n3026 ;
  assign y1525 = ~1'b0 ;
  assign y1526 = ~n1582 ;
  assign y1527 = ~1'b0 ;
  assign y1528 = n3027 ;
  assign y1529 = ~n3030 ;
  assign y1530 = ~n3033 ;
  assign y1531 = ~n3034 ;
  assign y1532 = ~n3039 ;
  assign y1533 = n27 ;
  assign y1534 = n3041 ;
  assign y1535 = ~n3044 ;
  assign y1536 = ~n3047 ;
  assign y1537 = ~1'b0 ;
  assign y1538 = ~n3050 ;
  assign y1539 = ~n3054 ;
  assign y1540 = ~n3063 ;
  assign y1541 = ~1'b0 ;
  assign y1542 = ~1'b0 ;
  assign y1543 = n3066 ;
  assign y1544 = ~1'b0 ;
  assign y1545 = n241 ;
  assign y1546 = ~1'b0 ;
  assign y1547 = n3068 ;
  assign y1548 = ~n682 ;
  assign y1549 = n3070 ;
  assign y1550 = ~1'b0 ;
  assign y1551 = n2922 ;
  assign y1552 = n2216 ;
  assign y1553 = n3080 ;
  assign y1554 = ~1'b0 ;
  assign y1555 = n3083 ;
  assign y1556 = n3090 ;
  assign y1557 = ~n3091 ;
  assign y1558 = n3094 ;
  assign y1559 = 1'b0 ;
  assign y1560 = ~n533 ;
  assign y1561 = ~n3096 ;
  assign y1562 = ~n3101 ;
  assign y1563 = ~1'b0 ;
  assign y1564 = ~1'b0 ;
  assign y1565 = n532 ;
  assign y1566 = ~1'b0 ;
  assign y1567 = ~n3110 ;
  assign y1568 = n1816 ;
  assign y1569 = ~n3111 ;
  assign y1570 = n3112 ;
  assign y1571 = ~n3113 ;
  assign y1572 = ~n3114 ;
  assign y1573 = ~n3115 ;
  assign y1574 = n3119 ;
  assign y1575 = ~n3122 ;
  assign y1576 = n3123 ;
  assign y1577 = ~n3124 ;
  assign y1578 = ~n3127 ;
  assign y1579 = n3131 ;
  assign y1580 = ~n3133 ;
  assign y1581 = n3140 ;
  assign y1582 = ~1'b0 ;
  assign y1583 = n3141 ;
  assign y1584 = ~n3142 ;
  assign y1585 = n3143 ;
  assign y1586 = n3147 ;
  assign y1587 = ~n3153 ;
  assign y1588 = ~n3157 ;
  assign y1589 = n3158 ;
  assign y1590 = n3163 ;
  assign y1591 = n2859 ;
  assign y1592 = n3178 ;
  assign y1593 = ~1'b0 ;
  assign y1594 = n3179 ;
  assign y1595 = ~1'b0 ;
  assign y1596 = n1202 ;
  assign y1597 = n3186 ;
  assign y1598 = ~n3187 ;
  assign y1599 = ~n3197 ;
  assign y1600 = n3199 ;
  assign y1601 = ~n3202 ;
  assign y1602 = n3206 ;
  assign y1603 = ~1'b0 ;
  assign y1604 = n3105 ;
  assign y1605 = ~1'b0 ;
  assign y1606 = ~1'b0 ;
  assign y1607 = n3207 ;
  assign y1608 = ~n3211 ;
  assign y1609 = n3213 ;
  assign y1610 = n3216 ;
  assign y1611 = ~1'b0 ;
  assign y1612 = ~n3219 ;
  assign y1613 = ~1'b0 ;
  assign y1614 = ~n3225 ;
  assign y1615 = n3226 ;
  assign y1616 = n3227 ;
  assign y1617 = n3228 ;
  assign y1618 = n3229 ;
  assign y1619 = n3235 ;
  assign y1620 = ~n3236 ;
  assign y1621 = n3239 ;
  assign y1622 = n3240 ;
  assign y1623 = ~n3243 ;
  assign y1624 = ~n3250 ;
  assign y1625 = n3251 ;
  assign y1626 = n2653 ;
  assign y1627 = ~1'b0 ;
  assign y1628 = ~n2094 ;
  assign y1629 = ~1'b0 ;
  assign y1630 = n3259 ;
  assign y1631 = ~1'b0 ;
  assign y1632 = ~1'b0 ;
  assign y1633 = 1'b0 ;
  assign y1634 = ~n3268 ;
  assign y1635 = ~n3270 ;
  assign y1636 = ~n3271 ;
  assign y1637 = ~n2787 ;
  assign y1638 = ~n3274 ;
  assign y1639 = n3276 ;
  assign y1640 = ~1'b0 ;
  assign y1641 = n3285 ;
  assign y1642 = ~n3287 ;
  assign y1643 = n3290 ;
  assign y1644 = 1'b0 ;
  assign y1645 = n3293 ;
  assign y1646 = 1'b0 ;
  assign y1647 = ~n3297 ;
  assign y1648 = ~n3299 ;
  assign y1649 = n3302 ;
  assign y1650 = n3307 ;
  assign y1651 = ~n1908 ;
  assign y1652 = ~n3308 ;
  assign y1653 = ~n3313 ;
  assign y1654 = ~1'b0 ;
  assign y1655 = ~n3318 ;
  assign y1656 = ~n3320 ;
  assign y1657 = ~1'b0 ;
  assign y1658 = ~n3328 ;
  assign y1659 = n3330 ;
  assign y1660 = n3334 ;
  assign y1661 = n3339 ;
  assign y1662 = n3341 ;
  assign y1663 = ~n3345 ;
  assign y1664 = ~n3347 ;
  assign y1665 = ~1'b0 ;
  assign y1666 = ~1'b0 ;
  assign y1667 = ~n3349 ;
  assign y1668 = ~1'b0 ;
  assign y1669 = n3351 ;
  assign y1670 = n3352 ;
  assign y1671 = n3353 ;
  assign y1672 = ~1'b0 ;
  assign y1673 = n492 ;
  assign y1674 = ~n3358 ;
  assign y1675 = ~1'b0 ;
  assign y1676 = ~n1455 ;
  assign y1677 = ~1'b0 ;
  assign y1678 = ~n3364 ;
  assign y1679 = ~n3371 ;
  assign y1680 = ~n3372 ;
  assign y1681 = n3374 ;
  assign y1682 = ~1'b0 ;
  assign y1683 = ~1'b0 ;
  assign y1684 = ~n3375 ;
  assign y1685 = n3377 ;
  assign y1686 = n3378 ;
  assign y1687 = n3379 ;
  assign y1688 = ~1'b0 ;
  assign y1689 = ~n342 ;
  assign y1690 = ~1'b0 ;
  assign y1691 = ~n3386 ;
  assign y1692 = ~n3389 ;
  assign y1693 = ~n3397 ;
  assign y1694 = n3402 ;
  assign y1695 = n3403 ;
  assign y1696 = ~1'b0 ;
  assign y1697 = n3408 ;
  assign y1698 = n3410 ;
  assign y1699 = ~1'b0 ;
  assign y1700 = ~1'b0 ;
  assign y1701 = ~n3413 ;
  assign y1702 = ~n3414 ;
  assign y1703 = n535 ;
  assign y1704 = ~1'b0 ;
  assign y1705 = ~1'b0 ;
  assign y1706 = ~1'b0 ;
  assign y1707 = ~n3417 ;
  assign y1708 = n3418 ;
  assign y1709 = ~1'b0 ;
  assign y1710 = n3422 ;
  assign y1711 = n1513 ;
  assign y1712 = n3428 ;
  assign y1713 = n1073 ;
  assign y1714 = n3429 ;
  assign y1715 = ~1'b0 ;
  assign y1716 = ~n3432 ;
  assign y1717 = ~1'b0 ;
  assign y1718 = 1'b0 ;
  assign y1719 = n3435 ;
  assign y1720 = ~n3439 ;
  assign y1721 = ~1'b0 ;
  assign y1722 = ~1'b0 ;
  assign y1723 = ~1'b0 ;
  assign y1724 = n3440 ;
  assign y1725 = n3441 ;
  assign y1726 = ~1'b0 ;
  assign y1727 = ~n3443 ;
  assign y1728 = ~n3235 ;
  assign y1729 = ~n3445 ;
  assign y1730 = ~n3448 ;
  assign y1731 = n3451 ;
  assign y1732 = ~1'b0 ;
  assign y1733 = ~1'b0 ;
  assign y1734 = ~1'b0 ;
  assign y1735 = ~n3453 ;
  assign y1736 = n3459 ;
  assign y1737 = ~n3465 ;
  assign y1738 = ~n1517 ;
  assign y1739 = ~1'b0 ;
  assign y1740 = ~n3466 ;
  assign y1741 = n3467 ;
  assign y1742 = n3469 ;
  assign y1743 = n3470 ;
  assign y1744 = n3471 ;
  assign y1745 = ~n3474 ;
  assign y1746 = n3475 ;
  assign y1747 = ~1'b0 ;
  assign y1748 = ~1'b0 ;
  assign y1749 = ~n3477 ;
  assign y1750 = n3483 ;
  assign y1751 = n3486 ;
  assign y1752 = ~n3488 ;
  assign y1753 = ~1'b0 ;
  assign y1754 = ~n3489 ;
  assign y1755 = ~1'b0 ;
  assign y1756 = 1'b0 ;
  assign y1757 = n3490 ;
  assign y1758 = ~1'b0 ;
  assign y1759 = n3494 ;
  assign y1760 = n3496 ;
  assign y1761 = ~1'b0 ;
  assign y1762 = ~n3501 ;
  assign y1763 = n3502 ;
  assign y1764 = ~n3505 ;
  assign y1765 = ~n1369 ;
  assign y1766 = ~1'b0 ;
  assign y1767 = n3510 ;
  assign y1768 = ~n3512 ;
  assign y1769 = ~n3519 ;
  assign y1770 = ~n3520 ;
  assign y1771 = ~1'b0 ;
  assign y1772 = ~n3522 ;
  assign y1773 = ~n3524 ;
  assign y1774 = ~n3529 ;
  assign y1775 = n3533 ;
  assign y1776 = ~1'b0 ;
  assign y1777 = ~n3535 ;
  assign y1778 = n3536 ;
  assign y1779 = ~n3539 ;
  assign y1780 = n2317 ;
  assign y1781 = n3349 ;
  assign y1782 = n3543 ;
  assign y1783 = ~1'b0 ;
  assign y1784 = ~n3545 ;
  assign y1785 = ~n3549 ;
  assign y1786 = ~n3550 ;
  assign y1787 = n3556 ;
  assign y1788 = ~n3558 ;
  assign y1789 = ~n3560 ;
  assign y1790 = ~n3567 ;
  assign y1791 = n3568 ;
  assign y1792 = n3572 ;
  assign y1793 = ~1'b0 ;
  assign y1794 = ~1'b0 ;
  assign y1795 = ~n3573 ;
  assign y1796 = n749 ;
  assign y1797 = ~1'b0 ;
  assign y1798 = ~n3574 ;
  assign y1799 = n3576 ;
  assign y1800 = 1'b0 ;
  assign y1801 = n3577 ;
  assign y1802 = ~n3579 ;
  assign y1803 = n3580 ;
  assign y1804 = n3583 ;
  assign y1805 = ~1'b0 ;
  assign y1806 = n3588 ;
  assign y1807 = n3591 ;
  assign y1808 = ~n61 ;
  assign y1809 = ~n3598 ;
  assign y1810 = n3599 ;
  assign y1811 = n3600 ;
  assign y1812 = ~n3603 ;
  assign y1813 = n3611 ;
  assign y1814 = ~1'b0 ;
  assign y1815 = ~n3612 ;
  assign y1816 = ~1'b0 ;
  assign y1817 = n3614 ;
  assign y1818 = n2637 ;
  assign y1819 = n3617 ;
  assign y1820 = ~n3618 ;
  assign y1821 = ~1'b0 ;
  assign y1822 = ~n3622 ;
  assign y1823 = n3623 ;
  assign y1824 = n3628 ;
  assign y1825 = n1284 ;
  assign y1826 = n3631 ;
  assign y1827 = n1083 ;
  assign y1828 = n3635 ;
  assign y1829 = ~1'b0 ;
  assign y1830 = ~n3636 ;
  assign y1831 = ~1'b0 ;
  assign y1832 = n3637 ;
  assign y1833 = 1'b0 ;
  assign y1834 = n3643 ;
  assign y1835 = ~n3652 ;
  assign y1836 = ~n3658 ;
  assign y1837 = ~n2645 ;
  assign y1838 = n3662 ;
  assign y1839 = ~1'b0 ;
  assign y1840 = ~n3663 ;
  assign y1841 = ~n3665 ;
  assign y1842 = ~1'b0 ;
  assign y1843 = n3668 ;
  assign y1844 = n3669 ;
  assign y1845 = ~1'b0 ;
  assign y1846 = ~1'b0 ;
  assign y1847 = ~n3672 ;
  assign y1848 = ~1'b0 ;
  assign y1849 = 1'b0 ;
  assign y1850 = ~n3674 ;
  assign y1851 = n3676 ;
  assign y1852 = n466 ;
  assign y1853 = ~n3682 ;
  assign y1854 = ~n3687 ;
  assign y1855 = ~n3690 ;
  assign y1856 = n3691 ;
  assign y1857 = 1'b0 ;
  assign y1858 = ~1'b0 ;
  assign y1859 = ~1'b0 ;
  assign y1860 = ~1'b0 ;
  assign y1861 = ~n3696 ;
  assign y1862 = ~n3700 ;
  assign y1863 = ~1'b0 ;
  assign y1864 = n86 ;
  assign y1865 = ~1'b0 ;
  assign y1866 = n3703 ;
  assign y1867 = ~n3708 ;
  assign y1868 = ~n3716 ;
  assign y1869 = 1'b0 ;
  assign y1870 = n3718 ;
  assign y1871 = ~n3723 ;
  assign y1872 = ~n3724 ;
  assign y1873 = ~1'b0 ;
  assign y1874 = ~n3725 ;
  assign y1875 = 1'b0 ;
  assign y1876 = ~1'b0 ;
  assign y1877 = ~n3726 ;
  assign y1878 = ~1'b0 ;
  assign y1879 = n3730 ;
  assign y1880 = n3731 ;
  assign y1881 = n3735 ;
  assign y1882 = ~1'b0 ;
  assign y1883 = ~n3736 ;
  assign y1884 = ~1'b0 ;
  assign y1885 = ~1'b0 ;
  assign y1886 = ~1'b0 ;
  assign y1887 = ~n3740 ;
  assign y1888 = ~n3741 ;
  assign y1889 = ~n3753 ;
  assign y1890 = ~n3755 ;
  assign y1891 = n3757 ;
  assign y1892 = ~n3758 ;
  assign y1893 = ~n3761 ;
  assign y1894 = ~1'b0 ;
  assign y1895 = n3763 ;
  assign y1896 = n3766 ;
  assign y1897 = ~n3779 ;
  assign y1898 = n3780 ;
  assign y1899 = 1'b0 ;
  assign y1900 = ~1'b0 ;
  assign y1901 = ~n3783 ;
  assign y1902 = ~n3792 ;
  assign y1903 = n3794 ;
  assign y1904 = n3798 ;
  assign y1905 = ~n3805 ;
  assign y1906 = n3807 ;
  assign y1907 = 1'b0 ;
  assign y1908 = ~n3809 ;
  assign y1909 = ~n3813 ;
  assign y1910 = ~1'b0 ;
  assign y1911 = n3827 ;
  assign y1912 = n2873 ;
  assign y1913 = ~1'b0 ;
  assign y1914 = ~1'b0 ;
  assign y1915 = n3833 ;
  assign y1916 = ~1'b0 ;
  assign y1917 = ~n3842 ;
  assign y1918 = n3848 ;
  assign y1919 = ~n3852 ;
  assign y1920 = ~1'b0 ;
  assign y1921 = n3853 ;
  assign y1922 = 1'b0 ;
  assign y1923 = ~n3856 ;
  assign y1924 = ~n3861 ;
  assign y1925 = n3864 ;
  assign y1926 = 1'b0 ;
  assign y1927 = ~n3873 ;
  assign y1928 = ~n3875 ;
  assign y1929 = ~1'b0 ;
  assign y1930 = ~1'b0 ;
  assign y1931 = n3876 ;
  assign y1932 = ~n3882 ;
  assign y1933 = n3884 ;
  assign y1934 = n3885 ;
  assign y1935 = ~n3886 ;
  assign y1936 = ~n3890 ;
  assign y1937 = n3891 ;
  assign y1938 = n3893 ;
  assign y1939 = ~n3894 ;
  assign y1940 = n3896 ;
  assign y1941 = ~1'b0 ;
  assign y1942 = n2539 ;
  assign y1943 = ~1'b0 ;
  assign y1944 = n3897 ;
  assign y1945 = ~1'b0 ;
  assign y1946 = ~1'b0 ;
  assign y1947 = n3011 ;
  assign y1948 = n3899 ;
  assign y1949 = 1'b0 ;
  assign y1950 = ~1'b0 ;
  assign y1951 = ~1'b0 ;
  assign y1952 = ~1'b0 ;
  assign y1953 = ~n3901 ;
  assign y1954 = n3903 ;
  assign y1955 = ~1'b0 ;
  assign y1956 = ~n3904 ;
  assign y1957 = ~n3911 ;
  assign y1958 = ~1'b0 ;
  assign y1959 = n3218 ;
  assign y1960 = ~n3912 ;
  assign y1961 = 1'b0 ;
  assign y1962 = ~n3913 ;
  assign y1963 = ~n3917 ;
  assign y1964 = ~1'b0 ;
  assign y1965 = ~1'b0 ;
  assign y1966 = ~1'b0 ;
  assign y1967 = n3920 ;
  assign y1968 = ~1'b0 ;
  assign y1969 = ~1'b0 ;
  assign y1970 = n2202 ;
  assign y1971 = n3891 ;
  assign y1972 = ~1'b0 ;
  assign y1973 = n2605 ;
  assign y1974 = ~n3921 ;
  assign y1975 = ~1'b0 ;
  assign y1976 = ~n3923 ;
  assign y1977 = ~1'b0 ;
  assign y1978 = ~1'b0 ;
  assign y1979 = n3924 ;
  assign y1980 = ~1'b0 ;
  assign y1981 = ~n3927 ;
  assign y1982 = ~n3932 ;
  assign y1983 = ~n1584 ;
  assign y1984 = ~1'b0 ;
  assign y1985 = ~n3934 ;
  assign y1986 = n3428 ;
  assign y1987 = n1081 ;
  assign y1988 = ~1'b0 ;
  assign y1989 = ~n3937 ;
  assign y1990 = n3944 ;
  assign y1991 = 1'b0 ;
  assign y1992 = ~n3950 ;
  assign y1993 = ~n3951 ;
  assign y1994 = n3952 ;
  assign y1995 = ~1'b0 ;
  assign y1996 = ~1'b0 ;
  assign y1997 = ~n3953 ;
  assign y1998 = n3955 ;
  assign y1999 = ~n3959 ;
  assign y2000 = ~n1161 ;
  assign y2001 = ~1'b0 ;
  assign y2002 = ~1'b0 ;
  assign y2003 = ~n3962 ;
  assign y2004 = n423 ;
  assign y2005 = ~n3966 ;
  assign y2006 = ~n3971 ;
  assign y2007 = ~1'b0 ;
  assign y2008 = n839 ;
  assign y2009 = ~1'b0 ;
  assign y2010 = ~n3972 ;
  assign y2011 = ~n3974 ;
  assign y2012 = ~1'b0 ;
  assign y2013 = ~n3979 ;
  assign y2014 = ~1'b0 ;
  assign y2015 = n3980 ;
  assign y2016 = n3982 ;
  assign y2017 = n3983 ;
  assign y2018 = ~n3985 ;
  assign y2019 = n3987 ;
  assign y2020 = 1'b0 ;
  assign y2021 = ~n3990 ;
  assign y2022 = ~n808 ;
  assign y2023 = ~n3992 ;
  assign y2024 = ~1'b0 ;
  assign y2025 = ~1'b0 ;
  assign y2026 = ~1'b0 ;
  assign y2027 = ~n3993 ;
  assign y2028 = ~n4000 ;
  assign y2029 = 1'b0 ;
  assign y2030 = n4001 ;
  assign y2031 = ~n4004 ;
  assign y2032 = ~1'b0 ;
  assign y2033 = ~n4005 ;
  assign y2034 = n4006 ;
  assign y2035 = ~n4009 ;
  assign y2036 = ~1'b0 ;
  assign y2037 = ~n4010 ;
  assign y2038 = ~n4015 ;
  assign y2039 = ~1'b0 ;
  assign y2040 = ~1'b0 ;
  assign y2041 = ~n4017 ;
  assign y2042 = ~1'b0 ;
  assign y2043 = ~n4019 ;
  assign y2044 = n4022 ;
  assign y2045 = ~1'b0 ;
  assign y2046 = ~n4025 ;
  assign y2047 = ~1'b0 ;
  assign y2048 = ~1'b0 ;
  assign y2049 = n4026 ;
  assign y2050 = ~1'b0 ;
  assign y2051 = n4030 ;
  assign y2052 = n4036 ;
  assign y2053 = ~n4039 ;
  assign y2054 = n4050 ;
  assign y2055 = ~n4051 ;
  assign y2056 = n4054 ;
  assign y2057 = n4058 ;
  assign y2058 = ~1'b0 ;
  assign y2059 = ~n4061 ;
  assign y2060 = ~1'b0 ;
  assign y2061 = ~1'b0 ;
  assign y2062 = ~n4063 ;
  assign y2063 = n4065 ;
  assign y2064 = ~1'b0 ;
  assign y2065 = n4066 ;
  assign y2066 = ~n4072 ;
  assign y2067 = ~1'b0 ;
  assign y2068 = ~n4075 ;
  assign y2069 = n1511 ;
  assign y2070 = ~1'b0 ;
  assign y2071 = n4079 ;
  assign y2072 = ~n4080 ;
  assign y2073 = 1'b0 ;
  assign y2074 = n4083 ;
  assign y2075 = n4084 ;
  assign y2076 = ~n4087 ;
  assign y2077 = ~1'b0 ;
  assign y2078 = n4089 ;
  assign y2079 = ~1'b0 ;
  assign y2080 = n4090 ;
  assign y2081 = ~1'b0 ;
  assign y2082 = n4092 ;
  assign y2083 = ~n4097 ;
  assign y2084 = n2206 ;
  assign y2085 = n4098 ;
  assign y2086 = n4100 ;
  assign y2087 = ~1'b0 ;
  assign y2088 = ~1'b0 ;
  assign y2089 = ~1'b0 ;
  assign y2090 = n4101 ;
  assign y2091 = ~n4105 ;
  assign y2092 = ~1'b0 ;
  assign y2093 = ~n4108 ;
  assign y2094 = ~n4111 ;
  assign y2095 = n4113 ;
  assign y2096 = n4114 ;
  assign y2097 = ~n4119 ;
  assign y2098 = ~1'b0 ;
  assign y2099 = ~1'b0 ;
  assign y2100 = ~1'b0 ;
  assign y2101 = ~1'b0 ;
  assign y2102 = ~n4122 ;
  assign y2103 = ~n4123 ;
  assign y2104 = ~1'b0 ;
  assign y2105 = n4125 ;
  assign y2106 = ~n4126 ;
  assign y2107 = ~n4132 ;
  assign y2108 = ~1'b0 ;
  assign y2109 = ~n2229 ;
  assign y2110 = ~n4135 ;
  assign y2111 = ~1'b0 ;
  assign y2112 = ~n4138 ;
  assign y2113 = ~n2041 ;
  assign y2114 = ~n4139 ;
  assign y2115 = ~1'b0 ;
  assign y2116 = ~1'b0 ;
  assign y2117 = ~n4147 ;
  assign y2118 = ~n4154 ;
  assign y2119 = ~1'b0 ;
  assign y2120 = ~n4155 ;
  assign y2121 = n4163 ;
  assign y2122 = ~1'b0 ;
  assign y2123 = n4166 ;
  assign y2124 = 1'b0 ;
  assign y2125 = ~n4167 ;
  assign y2126 = ~1'b0 ;
  assign y2127 = n4170 ;
  assign y2128 = ~n4171 ;
  assign y2129 = n4174 ;
  assign y2130 = ~n4178 ;
  assign y2131 = n4179 ;
  assign y2132 = ~n4183 ;
  assign y2133 = ~n4185 ;
  assign y2134 = n4187 ;
  assign y2135 = ~n4191 ;
  assign y2136 = n4193 ;
  assign y2137 = n4194 ;
  assign y2138 = ~1'b0 ;
  assign y2139 = n4199 ;
  assign y2140 = n4201 ;
  assign y2141 = ~1'b0 ;
  assign y2142 = ~n4205 ;
  assign y2143 = ~1'b0 ;
  assign y2144 = ~n4206 ;
  assign y2145 = ~n4211 ;
  assign y2146 = n4213 ;
  assign y2147 = ~1'b0 ;
  assign y2148 = ~1'b0 ;
  assign y2149 = n4214 ;
  assign y2150 = ~n4215 ;
  assign y2151 = ~1'b0 ;
  assign y2152 = ~1'b0 ;
  assign y2153 = ~n4220 ;
  assign y2154 = ~n4221 ;
  assign y2155 = ~1'b0 ;
  assign y2156 = n4226 ;
  assign y2157 = ~1'b0 ;
  assign y2158 = n1853 ;
  assign y2159 = ~1'b0 ;
  assign y2160 = n4231 ;
  assign y2161 = n1660 ;
  assign y2162 = ~n4234 ;
  assign y2163 = ~n4235 ;
  assign y2164 = ~1'b0 ;
  assign y2165 = ~1'b0 ;
  assign y2166 = ~1'b0 ;
  assign y2167 = n4236 ;
  assign y2168 = ~n4238 ;
  assign y2169 = ~n4240 ;
  assign y2170 = n4241 ;
  assign y2171 = ~n4248 ;
  assign y2172 = n4250 ;
  assign y2173 = n4251 ;
  assign y2174 = n4252 ;
  assign y2175 = n4256 ;
  assign y2176 = n4257 ;
  assign y2177 = ~1'b0 ;
  assign y2178 = n4260 ;
  assign y2179 = ~1'b0 ;
  assign y2180 = n4261 ;
  assign y2181 = n4264 ;
  assign y2182 = ~1'b0 ;
  assign y2183 = n4268 ;
  assign y2184 = ~n4269 ;
  assign y2185 = ~1'b0 ;
  assign y2186 = ~n4270 ;
  assign y2187 = ~n4271 ;
  assign y2188 = ~n4274 ;
  assign y2189 = ~n4276 ;
  assign y2190 = ~1'b0 ;
  assign y2191 = ~n4278 ;
  assign y2192 = ~1'b0 ;
  assign y2193 = ~1'b0 ;
  assign y2194 = n4279 ;
  assign y2195 = ~1'b0 ;
  assign y2196 = n4284 ;
  assign y2197 = ~n4285 ;
  assign y2198 = ~n4289 ;
  assign y2199 = ~n4294 ;
  assign y2200 = ~1'b0 ;
  assign y2201 = 1'b0 ;
  assign y2202 = ~1'b0 ;
  assign y2203 = ~1'b0 ;
  assign y2204 = ~n4295 ;
  assign y2205 = ~n4296 ;
  assign y2206 = n4299 ;
  assign y2207 = n4309 ;
  assign y2208 = ~1'b0 ;
  assign y2209 = ~n4312 ;
  assign y2210 = n4313 ;
  assign y2211 = n4315 ;
  assign y2212 = ~n4317 ;
  assign y2213 = ~n4322 ;
  assign y2214 = n4324 ;
  assign y2215 = n4325 ;
  assign y2216 = ~1'b0 ;
  assign y2217 = ~1'b0 ;
  assign y2218 = n4326 ;
  assign y2219 = ~n4327 ;
  assign y2220 = n4329 ;
  assign y2221 = n3052 ;
  assign y2222 = ~n4332 ;
  assign y2223 = ~1'b0 ;
  assign y2224 = ~1'b0 ;
  assign y2225 = n3193 ;
  assign y2226 = ~n4335 ;
  assign y2227 = ~n4338 ;
  assign y2228 = ~n4343 ;
  assign y2229 = ~n4346 ;
  assign y2230 = n4347 ;
  assign y2231 = ~n4348 ;
  assign y2232 = n4349 ;
  assign y2233 = ~1'b0 ;
  assign y2234 = n4350 ;
  assign y2235 = ~n4353 ;
  assign y2236 = n4355 ;
  assign y2237 = ~n4357 ;
  assign y2238 = ~n4361 ;
  assign y2239 = ~1'b0 ;
  assign y2240 = n3731 ;
  assign y2241 = ~n4364 ;
  assign y2242 = n4366 ;
  assign y2243 = ~n4367 ;
  assign y2244 = n4370 ;
  assign y2245 = n4372 ;
  assign y2246 = ~1'b0 ;
  assign y2247 = n4377 ;
  assign y2248 = n4378 ;
  assign y2249 = ~1'b0 ;
  assign y2250 = ~n4380 ;
  assign y2251 = ~1'b0 ;
  assign y2252 = ~n4381 ;
  assign y2253 = ~n4384 ;
  assign y2254 = n163 ;
  assign y2255 = ~1'b0 ;
  assign y2256 = ~1'b0 ;
  assign y2257 = n4386 ;
  assign y2258 = ~n4388 ;
  assign y2259 = ~n4389 ;
  assign y2260 = ~1'b0 ;
  assign y2261 = ~1'b0 ;
  assign y2262 = ~n4391 ;
  assign y2263 = ~n4392 ;
  assign y2264 = ~1'b0 ;
  assign y2265 = ~1'b0 ;
  assign y2266 = ~n4395 ;
  assign y2267 = ~1'b0 ;
  assign y2268 = ~n4402 ;
  assign y2269 = ~n4403 ;
  assign y2270 = ~n4406 ;
  assign y2271 = n4407 ;
  assign y2272 = n3258 ;
  assign y2273 = 1'b0 ;
  assign y2274 = ~1'b0 ;
  assign y2275 = n1918 ;
  assign y2276 = ~n4409 ;
  assign y2277 = ~n4410 ;
  assign y2278 = ~1'b0 ;
  assign y2279 = ~1'b0 ;
  assign y2280 = ~n4415 ;
  assign y2281 = n4416 ;
  assign y2282 = ~1'b0 ;
  assign y2283 = ~1'b0 ;
  assign y2284 = ~n4418 ;
  assign y2285 = ~n4420 ;
  assign y2286 = ~n4422 ;
  assign y2287 = ~1'b0 ;
  assign y2288 = ~1'b0 ;
  assign y2289 = ~n4425 ;
  assign y2290 = n4428 ;
  assign y2291 = n4432 ;
  assign y2292 = n4435 ;
  assign y2293 = ~n4436 ;
  assign y2294 = ~n1834 ;
  assign y2295 = ~n4438 ;
  assign y2296 = ~n4442 ;
  assign y2297 = ~n4446 ;
  assign y2298 = ~n4447 ;
  assign y2299 = n4448 ;
  assign y2300 = ~1'b0 ;
  assign y2301 = ~n4449 ;
  assign y2302 = ~n4451 ;
  assign y2303 = ~1'b0 ;
  assign y2304 = n4455 ;
  assign y2305 = n4457 ;
  assign y2306 = ~n4459 ;
  assign y2307 = ~n2387 ;
  assign y2308 = n4470 ;
  assign y2309 = 1'b0 ;
  assign y2310 = n4479 ;
  assign y2311 = ~n4480 ;
  assign y2312 = n4481 ;
  assign y2313 = ~n4485 ;
  assign y2314 = ~n4486 ;
  assign y2315 = ~n4491 ;
  assign y2316 = ~1'b0 ;
  assign y2317 = n4492 ;
  assign y2318 = n3003 ;
  assign y2319 = ~n4495 ;
  assign y2320 = ~n4496 ;
  assign y2321 = ~n4497 ;
  assign y2322 = ~n4499 ;
  assign y2323 = n4501 ;
  assign y2324 = ~1'b0 ;
  assign y2325 = n3774 ;
  assign y2326 = n4505 ;
  assign y2327 = n4506 ;
  assign y2328 = 1'b0 ;
  assign y2329 = ~n4512 ;
  assign y2330 = n4518 ;
  assign y2331 = n4525 ;
  assign y2332 = ~n4526 ;
  assign y2333 = n3867 ;
  assign y2334 = n4532 ;
  assign y2335 = ~n4535 ;
  assign y2336 = n4537 ;
  assign y2337 = ~1'b0 ;
  assign y2338 = n412 ;
  assign y2339 = n4544 ;
  assign y2340 = n4553 ;
  assign y2341 = ~1'b0 ;
  assign y2342 = ~n200 ;
  assign y2343 = ~1'b0 ;
  assign y2344 = ~n4554 ;
  assign y2345 = ~1'b0 ;
  assign y2346 = n4556 ;
  assign y2347 = ~1'b0 ;
  assign y2348 = ~n4559 ;
  assign y2349 = ~n4555 ;
  assign y2350 = 1'b0 ;
  assign y2351 = ~n4560 ;
  assign y2352 = ~n592 ;
  assign y2353 = ~n4561 ;
  assign y2354 = n4562 ;
  assign y2355 = ~1'b0 ;
  assign y2356 = ~1'b0 ;
  assign y2357 = n4563 ;
  assign y2358 = n4564 ;
  assign y2359 = n4569 ;
  assign y2360 = ~1'b0 ;
  assign y2361 = ~n2562 ;
  assign y2362 = ~n4578 ;
  assign y2363 = ~1'b0 ;
  assign y2364 = ~n4585 ;
  assign y2365 = ~n4586 ;
  assign y2366 = 1'b0 ;
  assign y2367 = n4587 ;
  assign y2368 = ~n4593 ;
  assign y2369 = n4597 ;
  assign y2370 = n4605 ;
  assign y2371 = n4608 ;
  assign y2372 = n4619 ;
  assign y2373 = ~n4629 ;
  assign y2374 = ~n2140 ;
  assign y2375 = n4631 ;
  assign y2376 = ~1'b0 ;
  assign y2377 = ~n4634 ;
  assign y2378 = n4635 ;
  assign y2379 = ~1'b0 ;
  assign y2380 = ~1'b0 ;
  assign y2381 = n4636 ;
  assign y2382 = n4639 ;
  assign y2383 = ~1'b0 ;
  assign y2384 = ~n4643 ;
  assign y2385 = n4644 ;
  assign y2386 = n4646 ;
  assign y2387 = ~n4648 ;
  assign y2388 = ~n4650 ;
  assign y2389 = ~n4653 ;
  assign y2390 = ~1'b0 ;
  assign y2391 = ~1'b0 ;
  assign y2392 = ~n4664 ;
  assign y2393 = ~1'b0 ;
  assign y2394 = ~n4666 ;
  assign y2395 = n4667 ;
  assign y2396 = ~n4672 ;
  assign y2397 = ~1'b0 ;
  assign y2398 = ~1'b0 ;
  assign y2399 = ~n4676 ;
  assign y2400 = n2721 ;
  assign y2401 = ~n4679 ;
  assign y2402 = ~1'b0 ;
  assign y2403 = ~n4681 ;
  assign y2404 = ~n4691 ;
  assign y2405 = ~1'b0 ;
  assign y2406 = ~n1226 ;
  assign y2407 = ~n4698 ;
  assign y2408 = n4700 ;
  assign y2409 = n4704 ;
  assign y2410 = ~1'b0 ;
  assign y2411 = ~1'b0 ;
  assign y2412 = n4711 ;
  assign y2413 = n4720 ;
  assign y2414 = ~1'b0 ;
  assign y2415 = ~1'b0 ;
  assign y2416 = n4722 ;
  assign y2417 = ~n4724 ;
  assign y2418 = n4733 ;
  assign y2419 = n4734 ;
  assign y2420 = n4738 ;
  assign y2421 = ~n4741 ;
  assign y2422 = n4744 ;
  assign y2423 = ~n4745 ;
  assign y2424 = ~n4750 ;
  assign y2425 = n4753 ;
  assign y2426 = ~1'b0 ;
  assign y2427 = n4761 ;
  assign y2428 = n4774 ;
  assign y2429 = n4775 ;
  assign y2430 = n4778 ;
  assign y2431 = ~n4784 ;
  assign y2432 = ~1'b0 ;
  assign y2433 = n3115 ;
  assign y2434 = n4787 ;
  assign y2435 = n4790 ;
  assign y2436 = ~n4796 ;
  assign y2437 = ~1'b0 ;
  assign y2438 = n2193 ;
  assign y2439 = ~n4797 ;
  assign y2440 = ~1'b0 ;
  assign y2441 = ~n4800 ;
  assign y2442 = ~n4802 ;
  assign y2443 = ~1'b0 ;
  assign y2444 = ~n4804 ;
  assign y2445 = ~1'b0 ;
  assign y2446 = ~n4808 ;
  assign y2447 = ~n4813 ;
  assign y2448 = n4814 ;
  assign y2449 = n4817 ;
  assign y2450 = ~n4824 ;
  assign y2451 = ~1'b0 ;
  assign y2452 = ~1'b0 ;
  assign y2453 = ~n4827 ;
  assign y2454 = ~n4832 ;
  assign y2455 = ~1'b0 ;
  assign y2456 = ~1'b0 ;
  assign y2457 = ~n470 ;
  assign y2458 = ~1'b0 ;
  assign y2459 = ~n4841 ;
  assign y2460 = ~1'b0 ;
  assign y2461 = n4843 ;
  assign y2462 = ~1'b0 ;
  assign y2463 = n3379 ;
  assign y2464 = ~n4848 ;
  assign y2465 = n4857 ;
  assign y2466 = ~n4858 ;
  assign y2467 = ~n4860 ;
  assign y2468 = ~n2359 ;
  assign y2469 = ~1'b0 ;
  assign y2470 = n2494 ;
  assign y2471 = ~n4862 ;
  assign y2472 = ~1'b0 ;
  assign y2473 = ~1'b0 ;
  assign y2474 = n4863 ;
  assign y2475 = ~n4865 ;
  assign y2476 = ~n4866 ;
  assign y2477 = 1'b0 ;
  assign y2478 = ~n4870 ;
  assign y2479 = n4873 ;
  assign y2480 = n3227 ;
  assign y2481 = n4877 ;
  assign y2482 = ~n4883 ;
  assign y2483 = ~n4884 ;
  assign y2484 = ~1'b0 ;
  assign y2485 = ~1'b0 ;
  assign y2486 = ~n4886 ;
  assign y2487 = n4888 ;
  assign y2488 = ~n4893 ;
  assign y2489 = ~n4899 ;
  assign y2490 = ~n4902 ;
  assign y2491 = ~1'b0 ;
  assign y2492 = ~1'b0 ;
  assign y2493 = n4903 ;
  assign y2494 = ~n4905 ;
  assign y2495 = ~1'b0 ;
  assign y2496 = n4909 ;
  assign y2497 = 1'b0 ;
  assign y2498 = n4917 ;
  assign y2499 = n4919 ;
  assign y2500 = n4921 ;
  assign y2501 = n3962 ;
  assign y2502 = n4928 ;
  assign y2503 = ~n4935 ;
  assign y2504 = n4938 ;
  assign y2505 = n4940 ;
  assign y2506 = ~1'b0 ;
  assign y2507 = n4941 ;
  assign y2508 = ~1'b0 ;
  assign y2509 = ~n4942 ;
  assign y2510 = n4947 ;
  assign y2511 = ~n4948 ;
  assign y2512 = ~n4955 ;
  assign y2513 = ~n4969 ;
  assign y2514 = ~1'b0 ;
  assign y2515 = ~n4970 ;
  assign y2516 = ~n4971 ;
  assign y2517 = ~1'b0 ;
  assign y2518 = ~n4973 ;
  assign y2519 = ~1'b0 ;
  assign y2520 = ~1'b0 ;
  assign y2521 = ~n4975 ;
  assign y2522 = ~n4976 ;
  assign y2523 = ~1'b0 ;
  assign y2524 = ~1'b0 ;
  assign y2525 = n4977 ;
  assign y2526 = n4979 ;
  assign y2527 = n4980 ;
  assign y2528 = ~n4981 ;
  assign y2529 = n4982 ;
  assign y2530 = ~1'b0 ;
  assign y2531 = ~n4989 ;
  assign y2532 = ~1'b0 ;
  assign y2533 = ~1'b0 ;
  assign y2534 = ~1'b0 ;
  assign y2535 = ~1'b0 ;
  assign y2536 = n582 ;
  assign y2537 = n4991 ;
  assign y2538 = ~1'b0 ;
  assign y2539 = ~n4995 ;
  assign y2540 = n5003 ;
  assign y2541 = ~n5005 ;
  assign y2542 = ~1'b0 ;
  assign y2543 = n5012 ;
  assign y2544 = ~n5015 ;
  assign y2545 = n5018 ;
  assign y2546 = n5022 ;
  assign y2547 = n5023 ;
  assign y2548 = ~1'b0 ;
  assign y2549 = n5025 ;
  assign y2550 = n5027 ;
  assign y2551 = ~1'b0 ;
  assign y2552 = ~n5028 ;
  assign y2553 = ~n5036 ;
  assign y2554 = ~n5040 ;
  assign y2555 = ~n5042 ;
  assign y2556 = n5045 ;
  assign y2557 = ~n5048 ;
  assign y2558 = n1111 ;
  assign y2559 = n5052 ;
  assign y2560 = ~n5055 ;
  assign y2561 = ~n5057 ;
  assign y2562 = ~1'b0 ;
  assign y2563 = n2087 ;
  assign y2564 = n5058 ;
  assign y2565 = ~1'b0 ;
  assign y2566 = n5059 ;
  assign y2567 = ~n934 ;
  assign y2568 = ~1'b0 ;
  assign y2569 = n3940 ;
  assign y2570 = ~n5064 ;
  assign y2571 = ~1'b0 ;
  assign y2572 = ~n5065 ;
  assign y2573 = ~1'b0 ;
  assign y2574 = ~n5070 ;
  assign y2575 = ~n3917 ;
  assign y2576 = ~n5072 ;
  assign y2577 = ~1'b0 ;
  assign y2578 = ~1'b0 ;
  assign y2579 = n5077 ;
  assign y2580 = ~n5078 ;
  assign y2581 = ~1'b0 ;
  assign y2582 = n5079 ;
  assign y2583 = n5081 ;
  assign y2584 = n5091 ;
  assign y2585 = ~n5093 ;
  assign y2586 = ~1'b0 ;
  assign y2587 = ~n5095 ;
  assign y2588 = ~n5101 ;
  assign y2589 = ~1'b0 ;
  assign y2590 = ~n5103 ;
  assign y2591 = ~1'b0 ;
  assign y2592 = n5106 ;
  assign y2593 = ~1'b0 ;
  assign y2594 = ~n5108 ;
  assign y2595 = ~1'b0 ;
  assign y2596 = n5118 ;
  assign y2597 = n5131 ;
  assign y2598 = n5138 ;
  assign y2599 = n5139 ;
  assign y2600 = n5141 ;
  assign y2601 = ~n5143 ;
  assign y2602 = ~1'b0 ;
  assign y2603 = ~1'b0 ;
  assign y2604 = ~1'b0 ;
  assign y2605 = ~1'b0 ;
  assign y2606 = n5144 ;
  assign y2607 = n5147 ;
  assign y2608 = ~n5157 ;
  assign y2609 = ~1'b0 ;
  assign y2610 = ~n5160 ;
  assign y2611 = n5161 ;
  assign y2612 = n5163 ;
  assign y2613 = n5165 ;
  assign y2614 = ~n5166 ;
  assign y2615 = n5167 ;
  assign y2616 = 1'b0 ;
  assign y2617 = ~n5172 ;
  assign y2618 = ~n2802 ;
  assign y2619 = ~1'b0 ;
  assign y2620 = 1'b0 ;
  assign y2621 = n5175 ;
  assign y2622 = ~1'b0 ;
  assign y2623 = ~n5178 ;
  assign y2624 = n5181 ;
  assign y2625 = ~n5182 ;
  assign y2626 = n5184 ;
  assign y2627 = ~1'b0 ;
  assign y2628 = n5195 ;
  assign y2629 = ~1'b0 ;
  assign y2630 = ~n5199 ;
  assign y2631 = n5200 ;
  assign y2632 = ~1'b0 ;
  assign y2633 = ~1'b0 ;
  assign y2634 = ~1'b0 ;
  assign y2635 = n5201 ;
  assign y2636 = ~1'b0 ;
  assign y2637 = n5206 ;
  assign y2638 = n5209 ;
  assign y2639 = ~1'b0 ;
  assign y2640 = 1'b0 ;
  assign y2641 = ~1'b0 ;
  assign y2642 = n5212 ;
  assign y2643 = ~1'b0 ;
  assign y2644 = n5214 ;
  assign y2645 = ~1'b0 ;
  assign y2646 = n5216 ;
  assign y2647 = ~n5218 ;
  assign y2648 = n5221 ;
  assign y2649 = ~n5224 ;
  assign y2650 = n5227 ;
  assign y2651 = ~n5232 ;
  assign y2652 = n3114 ;
  assign y2653 = ~1'b0 ;
  assign y2654 = n5235 ;
  assign y2655 = n5244 ;
  assign y2656 = ~n5245 ;
  assign y2657 = ~1'b0 ;
  assign y2658 = ~n5250 ;
  assign y2659 = ~1'b0 ;
  assign y2660 = n2763 ;
  assign y2661 = n5254 ;
  assign y2662 = n5256 ;
  assign y2663 = ~n5257 ;
  assign y2664 = ~n5258 ;
  assign y2665 = n5259 ;
  assign y2666 = ~n5260 ;
  assign y2667 = ~n5264 ;
  assign y2668 = n5268 ;
  assign y2669 = ~1'b0 ;
  assign y2670 = ~1'b0 ;
  assign y2671 = n5270 ;
  assign y2672 = ~n5277 ;
  assign y2673 = ~n5279 ;
  assign y2674 = ~1'b0 ;
  assign y2675 = ~n5284 ;
  assign y2676 = ~n5285 ;
  assign y2677 = ~n5286 ;
  assign y2678 = n5290 ;
  assign y2679 = 1'b0 ;
  assign y2680 = ~n5292 ;
  assign y2681 = n5296 ;
  assign y2682 = ~1'b0 ;
  assign y2683 = ~n5297 ;
  assign y2684 = n5298 ;
  assign y2685 = ~n5300 ;
  assign y2686 = ~1'b0 ;
  assign y2687 = ~1'b0 ;
  assign y2688 = ~1'b0 ;
  assign y2689 = n910 ;
  assign y2690 = ~n5305 ;
  assign y2691 = ~1'b0 ;
  assign y2692 = ~n5308 ;
  assign y2693 = ~1'b0 ;
  assign y2694 = ~n5310 ;
  assign y2695 = ~n5311 ;
  assign y2696 = ~1'b0 ;
  assign y2697 = n5313 ;
  assign y2698 = ~1'b0 ;
  assign y2699 = ~1'b0 ;
  assign y2700 = ~n5314 ;
  assign y2701 = ~1'b0 ;
  assign y2702 = n1182 ;
  assign y2703 = ~n1732 ;
  assign y2704 = ~1'b0 ;
  assign y2705 = ~n5316 ;
  assign y2706 = n5319 ;
  assign y2707 = n5324 ;
  assign y2708 = ~1'b0 ;
  assign y2709 = n5332 ;
  assign y2710 = n3646 ;
  assign y2711 = ~n5340 ;
  assign y2712 = n5346 ;
  assign y2713 = ~1'b0 ;
  assign y2714 = n5349 ;
  assign y2715 = n5360 ;
  assign y2716 = ~n5362 ;
  assign y2717 = n5366 ;
  assign y2718 = n5367 ;
  assign y2719 = ~n5368 ;
  assign y2720 = ~n5374 ;
  assign y2721 = ~n5377 ;
  assign y2722 = ~1'b0 ;
  assign y2723 = ~n1079 ;
  assign y2724 = ~n5381 ;
  assign y2725 = ~n5382 ;
  assign y2726 = n5385 ;
  assign y2727 = ~1'b0 ;
  assign y2728 = n3564 ;
  assign y2729 = ~1'b0 ;
  assign y2730 = ~1'b0 ;
  assign y2731 = ~n5387 ;
  assign y2732 = ~1'b0 ;
  assign y2733 = ~n5390 ;
  assign y2734 = ~1'b0 ;
  assign y2735 = ~n5391 ;
  assign y2736 = n5394 ;
  assign y2737 = ~n5401 ;
  assign y2738 = n5402 ;
  assign y2739 = n5404 ;
  assign y2740 = ~n5411 ;
  assign y2741 = ~1'b0 ;
  assign y2742 = ~1'b0 ;
  assign y2743 = n5413 ;
  assign y2744 = ~n5414 ;
  assign y2745 = ~n5419 ;
  assign y2746 = ~n5425 ;
  assign y2747 = ~1'b0 ;
  assign y2748 = n5426 ;
  assign y2749 = ~n5438 ;
  assign y2750 = ~n5052 ;
  assign y2751 = ~n5441 ;
  assign y2752 = n5442 ;
  assign y2753 = n5445 ;
  assign y2754 = ~1'b0 ;
  assign y2755 = ~1'b0 ;
  assign y2756 = ~1'b0 ;
  assign y2757 = n5446 ;
  assign y2758 = ~n5447 ;
  assign y2759 = ~1'b0 ;
  assign y2760 = n5449 ;
  assign y2761 = ~n5451 ;
  assign y2762 = n5452 ;
  assign y2763 = n5453 ;
  assign y2764 = 1'b0 ;
  assign y2765 = n5455 ;
  assign y2766 = ~n5456 ;
  assign y2767 = n5461 ;
  assign y2768 = n5464 ;
  assign y2769 = ~1'b0 ;
  assign y2770 = ~1'b0 ;
  assign y2771 = ~1'b0 ;
  assign y2772 = ~n5465 ;
  assign y2773 = ~n2540 ;
  assign y2774 = n5466 ;
  assign y2775 = n5467 ;
  assign y2776 = ~n5471 ;
  assign y2777 = n5472 ;
  assign y2778 = 1'b0 ;
  assign y2779 = ~n5474 ;
  assign y2780 = n5479 ;
  assign y2781 = n5482 ;
  assign y2782 = ~n1539 ;
  assign y2783 = n5485 ;
  assign y2784 = ~1'b0 ;
  assign y2785 = ~n5487 ;
  assign y2786 = ~1'b0 ;
  assign y2787 = ~n5336 ;
  assign y2788 = n5489 ;
  assign y2789 = n5490 ;
  assign y2790 = ~1'b0 ;
  assign y2791 = n5493 ;
  assign y2792 = ~n5501 ;
  assign y2793 = n5505 ;
  assign y2794 = ~n304 ;
  assign y2795 = ~n5507 ;
  assign y2796 = ~n5508 ;
  assign y2797 = n5510 ;
  assign y2798 = ~n5514 ;
  assign y2799 = ~n3537 ;
  assign y2800 = n5523 ;
  assign y2801 = n5525 ;
  assign y2802 = ~1'b0 ;
  assign y2803 = ~1'b0 ;
  assign y2804 = n5528 ;
  assign y2805 = n5395 ;
  assign y2806 = ~1'b0 ;
  assign y2807 = ~n5531 ;
  assign y2808 = ~n5535 ;
  assign y2809 = ~n5539 ;
  assign y2810 = n5540 ;
  assign y2811 = ~1'b0 ;
  assign y2812 = ~1'b0 ;
  assign y2813 = ~n5543 ;
  assign y2814 = n5544 ;
  assign y2815 = ~1'b0 ;
  assign y2816 = ~n5546 ;
  assign y2817 = ~n5547 ;
  assign y2818 = n5549 ;
  assign y2819 = ~1'b0 ;
  assign y2820 = ~n5551 ;
  assign y2821 = ~n5552 ;
  assign y2822 = ~1'b0 ;
  assign y2823 = ~1'b0 ;
  assign y2824 = ~1'b0 ;
  assign y2825 = n2173 ;
  assign y2826 = ~n5555 ;
  assign y2827 = n5557 ;
  assign y2828 = n5562 ;
  assign y2829 = n5563 ;
  assign y2830 = ~n5566 ;
  assign y2831 = ~1'b0 ;
  assign y2832 = n5570 ;
  assign y2833 = ~n5571 ;
  assign y2834 = ~1'b0 ;
  assign y2835 = ~n5573 ;
  assign y2836 = n5574 ;
  assign y2837 = ~1'b0 ;
  assign y2838 = n5575 ;
  assign y2839 = ~1'b0 ;
  assign y2840 = ~1'b0 ;
  assign y2841 = ~1'b0 ;
  assign y2842 = ~n4976 ;
  assign y2843 = n5576 ;
  assign y2844 = ~n5579 ;
  assign y2845 = ~1'b0 ;
  assign y2846 = ~1'b0 ;
  assign y2847 = ~1'b0 ;
  assign y2848 = ~1'b0 ;
  assign y2849 = ~n5581 ;
  assign y2850 = ~n5584 ;
  assign y2851 = ~1'b0 ;
  assign y2852 = ~1'b0 ;
  assign y2853 = n1471 ;
  assign y2854 = ~1'b0 ;
  assign y2855 = n5587 ;
  assign y2856 = ~1'b0 ;
  assign y2857 = ~1'b0 ;
  assign y2858 = n5591 ;
  assign y2859 = n2899 ;
  assign y2860 = ~1'b0 ;
  assign y2861 = ~n5592 ;
  assign y2862 = n5593 ;
  assign y2863 = n5594 ;
  assign y2864 = ~n5600 ;
  assign y2865 = ~1'b0 ;
  assign y2866 = ~n5607 ;
  assign y2867 = ~1'b0 ;
  assign y2868 = n5609 ;
  assign y2869 = n5615 ;
  assign y2870 = ~1'b0 ;
  assign y2871 = ~1'b0 ;
  assign y2872 = ~1'b0 ;
  assign y2873 = n5619 ;
  assign y2874 = n5621 ;
  assign y2875 = ~1'b0 ;
  assign y2876 = ~n5623 ;
  assign y2877 = n5624 ;
  assign y2878 = ~n5630 ;
  assign y2879 = ~1'b0 ;
  assign y2880 = n5632 ;
  assign y2881 = n4267 ;
  assign y2882 = ~1'b0 ;
  assign y2883 = ~n5636 ;
  assign y2884 = n5639 ;
  assign y2885 = n1772 ;
  assign y2886 = ~1'b0 ;
  assign y2887 = n5642 ;
  assign y2888 = ~n5645 ;
  assign y2889 = n5647 ;
  assign y2890 = n5649 ;
  assign y2891 = ~n5651 ;
  assign y2892 = n5655 ;
  assign y2893 = n5664 ;
  assign y2894 = ~n5668 ;
  assign y2895 = ~1'b0 ;
  assign y2896 = ~1'b0 ;
  assign y2897 = n5672 ;
  assign y2898 = ~1'b0 ;
  assign y2899 = n5673 ;
  assign y2900 = ~n320 ;
  assign y2901 = ~1'b0 ;
  assign y2902 = n5675 ;
  assign y2903 = n5676 ;
  assign y2904 = ~n5677 ;
  assign y2905 = ~1'b0 ;
  assign y2906 = ~n5680 ;
  assign y2907 = ~n5684 ;
  assign y2908 = ~1'b0 ;
  assign y2909 = ~1'b0 ;
  assign y2910 = ~n3058 ;
  assign y2911 = ~1'b0 ;
  assign y2912 = ~n5685 ;
  assign y2913 = ~n5686 ;
  assign y2914 = ~n5687 ;
  assign y2915 = n5691 ;
  assign y2916 = ~n5695 ;
  assign y2917 = ~n5699 ;
  assign y2918 = n302 ;
  assign y2919 = 1'b0 ;
  assign y2920 = n5700 ;
  assign y2921 = ~n5704 ;
  assign y2922 = ~n5706 ;
  assign y2923 = ~1'b0 ;
  assign y2924 = ~n5710 ;
  assign y2925 = ~n5717 ;
  assign y2926 = ~1'b0 ;
  assign y2927 = n4832 ;
  assign y2928 = ~1'b0 ;
  assign y2929 = ~1'b0 ;
  assign y2930 = ~n5724 ;
  assign y2931 = n5726 ;
  assign y2932 = ~n5730 ;
  assign y2933 = ~1'b0 ;
  assign y2934 = ~n5731 ;
  assign y2935 = ~n302 ;
  assign y2936 = n5734 ;
  assign y2937 = ~n5739 ;
  assign y2938 = ~n5743 ;
  assign y2939 = ~n5745 ;
  assign y2940 = ~n5749 ;
  assign y2941 = ~n5750 ;
  assign y2942 = n5751 ;
  assign y2943 = ~1'b0 ;
  assign y2944 = n5753 ;
  assign y2945 = ~n5760 ;
  assign y2946 = n5762 ;
  assign y2947 = ~n5763 ;
  assign y2948 = ~1'b0 ;
  assign y2949 = ~1'b0 ;
  assign y2950 = n5767 ;
  assign y2951 = n5768 ;
  assign y2952 = 1'b0 ;
  assign y2953 = ~1'b0 ;
  assign y2954 = n5771 ;
  assign y2955 = n5773 ;
  assign y2956 = n5783 ;
  assign y2957 = ~1'b0 ;
  assign y2958 = ~n5785 ;
  assign y2959 = n5789 ;
  assign y2960 = n5793 ;
  assign y2961 = ~n5795 ;
  assign y2962 = n5797 ;
  assign y2963 = n5799 ;
  assign y2964 = ~n5801 ;
  assign y2965 = ~n5803 ;
  assign y2966 = n3445 ;
  assign y2967 = ~1'b0 ;
  assign y2968 = ~1'b0 ;
  assign y2969 = n5807 ;
  assign y2970 = ~n5810 ;
  assign y2971 = n5812 ;
  assign y2972 = ~n5814 ;
  assign y2973 = n5816 ;
  assign y2974 = ~1'b0 ;
  assign y2975 = n5818 ;
  assign y2976 = ~n5819 ;
  assign y2977 = 1'b0 ;
  assign y2978 = ~1'b0 ;
  assign y2979 = ~n5829 ;
  assign y2980 = ~n5832 ;
  assign y2981 = n5835 ;
  assign y2982 = ~1'b0 ;
  assign y2983 = ~1'b0 ;
  assign y2984 = ~n4461 ;
  assign y2985 = ~n4139 ;
  assign y2986 = ~n5836 ;
  assign y2987 = ~1'b0 ;
  assign y2988 = n5845 ;
  assign y2989 = ~1'b0 ;
  assign y2990 = n5847 ;
  assign y2991 = ~1'b0 ;
  assign y2992 = n5849 ;
  assign y2993 = n5850 ;
  assign y2994 = ~1'b0 ;
  assign y2995 = n5851 ;
  assign y2996 = ~1'b0 ;
  assign y2997 = ~1'b0 ;
  assign y2998 = ~1'b0 ;
  assign y2999 = ~1'b0 ;
  assign y3000 = ~n4533 ;
  assign y3001 = n5857 ;
  assign y3002 = ~n5861 ;
  assign y3003 = ~1'b0 ;
  assign y3004 = n5863 ;
  assign y3005 = n5864 ;
  assign y3006 = n40 ;
  assign y3007 = ~1'b0 ;
  assign y3008 = n2275 ;
  assign y3009 = ~1'b0 ;
  assign y3010 = n5867 ;
  assign y3011 = ~n5868 ;
  assign y3012 = n5871 ;
  assign y3013 = ~n5873 ;
  assign y3014 = ~n5877 ;
  assign y3015 = n2815 ;
  assign y3016 = n5879 ;
  assign y3017 = ~n5880 ;
  assign y3018 = ~n5890 ;
  assign y3019 = 1'b0 ;
  assign y3020 = ~n5896 ;
  assign y3021 = ~1'b0 ;
  assign y3022 = ~1'b0 ;
  assign y3023 = ~n5897 ;
  assign y3024 = ~1'b0 ;
  assign y3025 = ~1'b0 ;
  assign y3026 = ~1'b0 ;
  assign y3027 = n5908 ;
  assign y3028 = n5912 ;
  assign y3029 = n5915 ;
  assign y3030 = n5917 ;
  assign y3031 = ~1'b0 ;
  assign y3032 = n5921 ;
  assign y3033 = ~n5932 ;
  assign y3034 = n5933 ;
  assign y3035 = n5936 ;
  assign y3036 = n5945 ;
  assign y3037 = n5946 ;
  assign y3038 = 1'b0 ;
  assign y3039 = ~1'b0 ;
  assign y3040 = ~n5948 ;
  assign y3041 = n5950 ;
  assign y3042 = ~n5953 ;
  assign y3043 = ~n5956 ;
  assign y3044 = ~n5958 ;
  assign y3045 = ~1'b0 ;
  assign y3046 = n5967 ;
  assign y3047 = ~1'b0 ;
  assign y3048 = ~n5969 ;
  assign y3049 = ~1'b0 ;
  assign y3050 = n5970 ;
  assign y3051 = ~1'b0 ;
  assign y3052 = n5971 ;
  assign y3053 = n5974 ;
  assign y3054 = n5978 ;
  assign y3055 = n5980 ;
  assign y3056 = 1'b0 ;
  assign y3057 = ~1'b0 ;
  assign y3058 = ~n3088 ;
  assign y3059 = n5982 ;
  assign y3060 = n5984 ;
  assign y3061 = ~1'b0 ;
  assign y3062 = ~n5986 ;
  assign y3063 = ~1'b0 ;
  assign y3064 = n5989 ;
  assign y3065 = ~n5994 ;
  assign y3066 = n5995 ;
  assign y3067 = n6000 ;
  assign y3068 = n6001 ;
  assign y3069 = ~n6002 ;
  assign y3070 = ~1'b0 ;
  assign y3071 = n6007 ;
  assign y3072 = n6009 ;
  assign y3073 = ~n6015 ;
  assign y3074 = n6016 ;
  assign y3075 = n6018 ;
  assign y3076 = n6019 ;
  assign y3077 = n6024 ;
  assign y3078 = n6026 ;
  assign y3079 = ~1'b0 ;
  assign y3080 = n6032 ;
  assign y3081 = ~1'b0 ;
  assign y3082 = n6033 ;
  assign y3083 = ~n6035 ;
  assign y3084 = ~n6036 ;
  assign y3085 = ~n6038 ;
  assign y3086 = ~n6039 ;
  assign y3087 = ~1'b0 ;
  assign y3088 = ~n6043 ;
  assign y3089 = ~n83 ;
  assign y3090 = ~n6051 ;
  assign y3091 = ~n6052 ;
  assign y3092 = n6054 ;
  assign y3093 = n322 ;
  assign y3094 = n6058 ;
  assign y3095 = n6060 ;
  assign y3096 = n6063 ;
  assign y3097 = n1411 ;
  assign y3098 = ~1'b0 ;
  assign y3099 = ~n6069 ;
  assign y3100 = n6070 ;
  assign y3101 = ~n6074 ;
  assign y3102 = ~n3710 ;
  assign y3103 = ~1'b0 ;
  assign y3104 = n6079 ;
  assign y3105 = ~n6080 ;
  assign y3106 = n6081 ;
  assign y3107 = ~n6082 ;
  assign y3108 = n6083 ;
  assign y3109 = n6094 ;
  assign y3110 = n6098 ;
  assign y3111 = ~n6100 ;
  assign y3112 = ~1'b0 ;
  assign y3113 = ~n6102 ;
  assign y3114 = ~1'b0 ;
  assign y3115 = ~n6106 ;
  assign y3116 = ~1'b0 ;
  assign y3117 = ~n4485 ;
  assign y3118 = ~n2363 ;
  assign y3119 = ~n6111 ;
  assign y3120 = n6112 ;
  assign y3121 = ~1'b0 ;
  assign y3122 = ~n2791 ;
  assign y3123 = n6121 ;
  assign y3124 = ~n6124 ;
  assign y3125 = ~n6126 ;
  assign y3126 = n6127 ;
  assign y3127 = ~n6128 ;
  assign y3128 = ~n6131 ;
  assign y3129 = ~n6135 ;
  assign y3130 = ~n1635 ;
  assign y3131 = n3314 ;
  assign y3132 = ~n6136 ;
  assign y3133 = n6140 ;
  assign y3134 = ~n6142 ;
  assign y3135 = n1057 ;
  assign y3136 = ~n6147 ;
  assign y3137 = ~1'b0 ;
  assign y3138 = ~n6154 ;
  assign y3139 = n6156 ;
  assign y3140 = ~1'b0 ;
  assign y3141 = ~1'b0 ;
  assign y3142 = ~1'b0 ;
  assign y3143 = n2663 ;
  assign y3144 = ~n6159 ;
  assign y3145 = ~n6162 ;
  assign y3146 = n6164 ;
  assign y3147 = n6165 ;
  assign y3148 = ~n6166 ;
  assign y3149 = ~n6168 ;
  assign y3150 = n6175 ;
  assign y3151 = ~n6177 ;
  assign y3152 = ~n6180 ;
  assign y3153 = ~1'b0 ;
  assign y3154 = n6181 ;
  assign y3155 = n6183 ;
  assign y3156 = ~n6184 ;
  assign y3157 = ~n6189 ;
  assign y3158 = ~n6190 ;
  assign y3159 = ~n6195 ;
  assign y3160 = ~n6205 ;
  assign y3161 = ~1'b0 ;
  assign y3162 = ~1'b0 ;
  assign y3163 = n6215 ;
  assign y3164 = ~1'b0 ;
  assign y3165 = n6216 ;
  assign y3166 = ~n6217 ;
  assign y3167 = n774 ;
  assign y3168 = ~n6218 ;
  assign y3169 = ~n6221 ;
  assign y3170 = ~n4666 ;
  assign y3171 = ~n6225 ;
  assign y3172 = n6227 ;
  assign y3173 = n6229 ;
  assign y3174 = n6230 ;
  assign y3175 = ~1'b0 ;
  assign y3176 = ~1'b0 ;
  assign y3177 = ~1'b0 ;
  assign y3178 = ~1'b0 ;
  assign y3179 = ~n6234 ;
  assign y3180 = ~n6235 ;
  assign y3181 = n6236 ;
  assign y3182 = ~n6238 ;
  assign y3183 = ~n6241 ;
  assign y3184 = n6250 ;
  assign y3185 = ~n727 ;
  assign y3186 = ~1'b0 ;
  assign y3187 = ~1'b0 ;
  assign y3188 = ~1'b0 ;
  assign y3189 = ~n6252 ;
  assign y3190 = ~1'b0 ;
  assign y3191 = ~n6255 ;
  assign y3192 = ~n6216 ;
  assign y3193 = ~n6256 ;
  assign y3194 = n6257 ;
  assign y3195 = ~1'b0 ;
  assign y3196 = n6258 ;
  assign y3197 = ~n6261 ;
  assign y3198 = ~n6262 ;
  assign y3199 = ~n6265 ;
  assign y3200 = ~n6267 ;
  assign y3201 = ~n6271 ;
  assign y3202 = n6272 ;
  assign y3203 = ~n6273 ;
  assign y3204 = ~1'b0 ;
  assign y3205 = ~n5458 ;
  assign y3206 = n6100 ;
  assign y3207 = n6275 ;
  assign y3208 = ~n6277 ;
  assign y3209 = ~1'b0 ;
  assign y3210 = 1'b0 ;
  assign y3211 = n6279 ;
  assign y3212 = ~1'b0 ;
  assign y3213 = n6280 ;
  assign y3214 = ~n6283 ;
  assign y3215 = n6287 ;
  assign y3216 = n6290 ;
  assign y3217 = ~1'b0 ;
  assign y3218 = n5464 ;
  assign y3219 = ~n6293 ;
  assign y3220 = n6296 ;
  assign y3221 = ~n6299 ;
  assign y3222 = ~n6300 ;
  assign y3223 = ~1'b0 ;
  assign y3224 = ~n6307 ;
  assign y3225 = ~1'b0 ;
  assign y3226 = ~1'b0 ;
  assign y3227 = ~1'b0 ;
  assign y3228 = ~1'b0 ;
  assign y3229 = ~n6308 ;
  assign y3230 = ~n6310 ;
  assign y3231 = n6314 ;
  assign y3232 = ~1'b0 ;
  assign y3233 = ~1'b0 ;
  assign y3234 = ~n6316 ;
  assign y3235 = n6320 ;
  assign y3236 = ~1'b0 ;
  assign y3237 = ~n6332 ;
  assign y3238 = ~n6335 ;
  assign y3239 = ~n6338 ;
  assign y3240 = ~n6340 ;
  assign y3241 = ~n6343 ;
  assign y3242 = n6344 ;
  assign y3243 = ~n6348 ;
  assign y3244 = ~1'b0 ;
  assign y3245 = n5104 ;
  assign y3246 = ~n6350 ;
  assign y3247 = ~1'b0 ;
  assign y3248 = n6354 ;
  assign y3249 = n6254 ;
  assign y3250 = ~n6356 ;
  assign y3251 = ~n6365 ;
  assign y3252 = n6368 ;
  assign y3253 = ~n6370 ;
  assign y3254 = ~1'b0 ;
  assign y3255 = n6372 ;
  assign y3256 = ~1'b0 ;
  assign y3257 = n6376 ;
  assign y3258 = ~n6377 ;
  assign y3259 = ~1'b0 ;
  assign y3260 = 1'b0 ;
  assign y3261 = ~1'b0 ;
  assign y3262 = ~1'b0 ;
  assign y3263 = ~n3243 ;
  assign y3264 = ~1'b0 ;
  assign y3265 = n1845 ;
  assign y3266 = ~n6381 ;
  assign y3267 = 1'b0 ;
  assign y3268 = n6383 ;
  assign y3269 = n6389 ;
  assign y3270 = ~n6393 ;
  assign y3271 = ~1'b0 ;
  assign y3272 = ~n6397 ;
  assign y3273 = ~n6398 ;
  assign y3274 = ~n6404 ;
  assign y3275 = n6405 ;
  assign y3276 = n6406 ;
  assign y3277 = ~n6409 ;
  assign y3278 = ~n6410 ;
  assign y3279 = ~n6413 ;
  assign y3280 = ~n6415 ;
  assign y3281 = n6417 ;
  assign y3282 = ~n6423 ;
  assign y3283 = ~n466 ;
  assign y3284 = ~n6424 ;
  assign y3285 = n6426 ;
  assign y3286 = ~n1269 ;
  assign y3287 = ~n6429 ;
  assign y3288 = ~n6430 ;
  assign y3289 = ~1'b0 ;
  assign y3290 = ~n6431 ;
  assign y3291 = n1453 ;
  assign y3292 = n6433 ;
  assign y3293 = n6434 ;
  assign y3294 = ~1'b0 ;
  assign y3295 = ~n6435 ;
  assign y3296 = ~1'b0 ;
  assign y3297 = ~n6439 ;
  assign y3298 = ~1'b0 ;
  assign y3299 = ~n1083 ;
  assign y3300 = ~1'b0 ;
  assign y3301 = ~n6441 ;
  assign y3302 = ~n6442 ;
  assign y3303 = ~n6447 ;
  assign y3304 = ~n6454 ;
  assign y3305 = n6455 ;
  assign y3306 = ~1'b0 ;
  assign y3307 = n6456 ;
  assign y3308 = ~n6457 ;
  assign y3309 = n6458 ;
  assign y3310 = ~n2185 ;
  assign y3311 = ~1'b0 ;
  assign y3312 = ~1'b0 ;
  assign y3313 = ~1'b0 ;
  assign y3314 = ~n6463 ;
  assign y3315 = ~1'b0 ;
  assign y3316 = ~n6468 ;
  assign y3317 = n6473 ;
  assign y3318 = ~1'b0 ;
  assign y3319 = 1'b0 ;
  assign y3320 = ~n6482 ;
  assign y3321 = n6483 ;
  assign y3322 = ~1'b0 ;
  assign y3323 = ~n6486 ;
  assign y3324 = n6492 ;
  assign y3325 = ~1'b0 ;
  assign y3326 = ~1'b0 ;
  assign y3327 = ~1'b0 ;
  assign y3328 = n6504 ;
  assign y3329 = ~n6507 ;
  assign y3330 = n4104 ;
  assign y3331 = n6509 ;
  assign y3332 = 1'b0 ;
  assign y3333 = ~1'b0 ;
  assign y3334 = ~n6511 ;
  assign y3335 = ~n6523 ;
  assign y3336 = ~1'b0 ;
  assign y3337 = n6524 ;
  assign y3338 = ~1'b0 ;
  assign y3339 = n6530 ;
  assign y3340 = ~n6537 ;
  assign y3341 = n6540 ;
  assign y3342 = ~n6553 ;
  assign y3343 = ~1'b0 ;
  assign y3344 = 1'b0 ;
  assign y3345 = ~n6557 ;
  assign y3346 = ~n6102 ;
  assign y3347 = ~n6566 ;
  assign y3348 = ~1'b0 ;
  assign y3349 = n6570 ;
  assign y3350 = ~n5803 ;
  assign y3351 = n6572 ;
  assign y3352 = ~1'b0 ;
  assign y3353 = n6573 ;
  assign y3354 = ~1'b0 ;
  assign y3355 = ~n6574 ;
  assign y3356 = ~1'b0 ;
  assign y3357 = ~n2755 ;
  assign y3358 = ~n6576 ;
  assign y3359 = ~n6580 ;
  assign y3360 = ~1'b0 ;
  assign y3361 = ~n6581 ;
  assign y3362 = n6585 ;
  assign y3363 = ~1'b0 ;
  assign y3364 = ~n6588 ;
  assign y3365 = n6595 ;
  assign y3366 = ~1'b0 ;
  assign y3367 = ~n6599 ;
  assign y3368 = ~n6601 ;
  assign y3369 = n6604 ;
  assign y3370 = ~n6605 ;
  assign y3371 = ~n6608 ;
  assign y3372 = ~n6610 ;
  assign y3373 = ~n6613 ;
  assign y3374 = n6616 ;
  assign y3375 = n2473 ;
  assign y3376 = ~1'b0 ;
  assign y3377 = ~1'b0 ;
  assign y3378 = n6617 ;
  assign y3379 = n6619 ;
  assign y3380 = n6621 ;
  assign y3381 = ~1'b0 ;
  assign y3382 = 1'b0 ;
  assign y3383 = n6628 ;
  assign y3384 = ~1'b0 ;
  assign y3385 = ~n6630 ;
  assign y3386 = ~n6631 ;
  assign y3387 = ~n564 ;
  assign y3388 = n6632 ;
  assign y3389 = ~n6633 ;
  assign y3390 = ~n6638 ;
  assign y3391 = ~n6641 ;
  assign y3392 = n6643 ;
  assign y3393 = n6645 ;
  assign y3394 = n6646 ;
  assign y3395 = n6650 ;
  assign y3396 = n6653 ;
  assign y3397 = n6656 ;
  assign y3398 = ~n6657 ;
  assign y3399 = ~1'b0 ;
  assign y3400 = n138 ;
  assign y3401 = ~n6662 ;
  assign y3402 = ~n6665 ;
  assign y3403 = n6667 ;
  assign y3404 = n6669 ;
  assign y3405 = n6670 ;
  assign y3406 = ~1'b0 ;
  assign y3407 = ~n6675 ;
  assign y3408 = ~n6678 ;
  assign y3409 = ~1'b0 ;
  assign y3410 = ~n6680 ;
  assign y3411 = ~1'b0 ;
  assign y3412 = ~1'b0 ;
  assign y3413 = ~1'b0 ;
  assign y3414 = ~n6681 ;
  assign y3415 = ~1'b0 ;
  assign y3416 = ~n6683 ;
  assign y3417 = ~n6685 ;
  assign y3418 = n6687 ;
  assign y3419 = ~n6692 ;
  assign y3420 = ~1'b0 ;
  assign y3421 = n6695 ;
  assign y3422 = ~n6697 ;
  assign y3423 = ~1'b0 ;
  assign y3424 = n6699 ;
  assign y3425 = ~1'b0 ;
  assign y3426 = ~n6700 ;
  assign y3427 = ~n6702 ;
  assign y3428 = ~n6704 ;
  assign y3429 = ~1'b0 ;
  assign y3430 = n6707 ;
  assign y3431 = ~n6712 ;
  assign y3432 = ~1'b0 ;
  assign y3433 = ~1'b0 ;
  assign y3434 = ~n6713 ;
  assign y3435 = ~1'b0 ;
  assign y3436 = n6716 ;
  assign y3437 = n6717 ;
  assign y3438 = n6720 ;
  assign y3439 = ~1'b0 ;
  assign y3440 = ~n6726 ;
  assign y3441 = ~n6731 ;
  assign y3442 = n6732 ;
  assign y3443 = ~n6736 ;
  assign y3444 = n6738 ;
  assign y3445 = ~1'b0 ;
  assign y3446 = ~n6742 ;
  assign y3447 = ~n6747 ;
  assign y3448 = ~n6749 ;
  assign y3449 = ~1'b0 ;
  assign y3450 = ~n6750 ;
  assign y3451 = ~n6751 ;
  assign y3452 = ~n6754 ;
  assign y3453 = ~n6759 ;
  assign y3454 = n4224 ;
  assign y3455 = ~n6760 ;
  assign y3456 = n6761 ;
  assign y3457 = ~n6763 ;
  assign y3458 = ~1'b0 ;
  assign y3459 = n6764 ;
  assign y3460 = ~n6765 ;
  assign y3461 = ~n6766 ;
  assign y3462 = n6769 ;
  assign y3463 = ~1'b0 ;
  assign y3464 = n6770 ;
  assign y3465 = ~n6774 ;
  assign y3466 = n6775 ;
  assign y3467 = ~1'b0 ;
  assign y3468 = ~n6777 ;
  assign y3469 = ~n6779 ;
  assign y3470 = ~1'b0 ;
  assign y3471 = n2980 ;
  assign y3472 = n6780 ;
  assign y3473 = n6785 ;
  assign y3474 = ~1'b0 ;
  assign y3475 = ~1'b0 ;
  assign y3476 = ~n6787 ;
  assign y3477 = ~n6797 ;
  assign y3478 = ~n6804 ;
  assign y3479 = n6809 ;
  assign y3480 = ~n6814 ;
  assign y3481 = ~n6815 ;
  assign y3482 = ~n56 ;
  assign y3483 = ~n6818 ;
  assign y3484 = ~1'b0 ;
  assign y3485 = n6824 ;
  assign y3486 = ~n6825 ;
  assign y3487 = ~1'b0 ;
  assign y3488 = ~1'b0 ;
  assign y3489 = ~n6829 ;
  assign y3490 = ~1'b0 ;
  assign y3491 = ~n3083 ;
  assign y3492 = ~1'b0 ;
  assign y3493 = ~n6832 ;
  assign y3494 = ~n6833 ;
  assign y3495 = ~1'b0 ;
  assign y3496 = ~n6836 ;
  assign y3497 = ~n6841 ;
  assign y3498 = ~1'b0 ;
  assign y3499 = ~1'b0 ;
  assign y3500 = ~n6844 ;
  assign y3501 = ~n4856 ;
  assign y3502 = n6847 ;
  assign y3503 = n6850 ;
  assign y3504 = ~n6851 ;
  assign y3505 = n6852 ;
  assign y3506 = ~n6855 ;
  assign y3507 = ~n6863 ;
  assign y3508 = ~n98 ;
  assign y3509 = ~1'b0 ;
  assign y3510 = ~1'b0 ;
  assign y3511 = ~1'b0 ;
  assign y3512 = ~1'b0 ;
  assign y3513 = n6869 ;
  assign y3514 = ~n6874 ;
  assign y3515 = n6876 ;
  assign y3516 = ~n6878 ;
  assign y3517 = ~n6886 ;
  assign y3518 = ~1'b0 ;
  assign y3519 = n6890 ;
  assign y3520 = ~1'b0 ;
  assign y3521 = ~n6891 ;
  assign y3522 = n6896 ;
  assign y3523 = n6898 ;
  assign y3524 = ~1'b0 ;
  assign y3525 = ~n6901 ;
  assign y3526 = ~1'b0 ;
  assign y3527 = ~1'b0 ;
  assign y3528 = n6902 ;
  assign y3529 = n6906 ;
  assign y3530 = ~1'b0 ;
  assign y3531 = n2048 ;
  assign y3532 = n6907 ;
  assign y3533 = ~1'b0 ;
  assign y3534 = ~1'b0 ;
  assign y3535 = n6910 ;
  assign y3536 = ~n6911 ;
  assign y3537 = ~n6919 ;
  assign y3538 = ~1'b0 ;
  assign y3539 = n6924 ;
  assign y3540 = n6925 ;
  assign y3541 = ~n6926 ;
  assign y3542 = ~n6928 ;
  assign y3543 = ~n6930 ;
  assign y3544 = n6935 ;
  assign y3545 = ~n6939 ;
  assign y3546 = n6940 ;
  assign y3547 = ~n6941 ;
  assign y3548 = ~1'b0 ;
  assign y3549 = ~n6942 ;
  assign y3550 = ~n6943 ;
  assign y3551 = n6944 ;
  assign y3552 = n6945 ;
  assign y3553 = ~n6946 ;
  assign y3554 = ~n6948 ;
  assign y3555 = ~n6949 ;
  assign y3556 = n6950 ;
  assign y3557 = ~n6951 ;
  assign y3558 = n6955 ;
  assign y3559 = ~n6959 ;
  assign y3560 = n6963 ;
  assign y3561 = n5547 ;
  assign y3562 = ~1'b0 ;
  assign y3563 = ~1'b0 ;
  assign y3564 = n6964 ;
  assign y3565 = ~n6966 ;
  assign y3566 = n1377 ;
  assign y3567 = ~1'b0 ;
  assign y3568 = n6972 ;
  assign y3569 = n6978 ;
  assign y3570 = ~n6981 ;
  assign y3571 = ~1'b0 ;
  assign y3572 = ~n6982 ;
  assign y3573 = ~n6985 ;
  assign y3574 = ~n6986 ;
  assign y3575 = ~1'b0 ;
  assign y3576 = ~n6989 ;
  assign y3577 = ~1'b0 ;
  assign y3578 = n6990 ;
  assign y3579 = ~1'b0 ;
  assign y3580 = n6996 ;
  assign y3581 = n6999 ;
  assign y3582 = ~n7003 ;
  assign y3583 = ~1'b0 ;
  assign y3584 = ~n6598 ;
  assign y3585 = n7010 ;
  assign y3586 = ~n7012 ;
  assign y3587 = n7020 ;
  assign y3588 = n7022 ;
  assign y3589 = ~1'b0 ;
  assign y3590 = ~n7023 ;
  assign y3591 = ~n7029 ;
  assign y3592 = ~n6048 ;
  assign y3593 = ~1'b0 ;
  assign y3594 = ~1'b0 ;
  assign y3595 = ~n7030 ;
  assign y3596 = ~n7034 ;
  assign y3597 = ~1'b0 ;
  assign y3598 = n7036 ;
  assign y3599 = 1'b0 ;
  assign y3600 = n7038 ;
  assign y3601 = ~1'b0 ;
  assign y3602 = ~1'b0 ;
  assign y3603 = 1'b0 ;
  assign y3604 = n7041 ;
  assign y3605 = ~n7047 ;
  assign y3606 = n7053 ;
  assign y3607 = ~1'b0 ;
  assign y3608 = n7061 ;
  assign y3609 = ~n7063 ;
  assign y3610 = n7073 ;
  assign y3611 = n7076 ;
  assign y3612 = ~1'b0 ;
  assign y3613 = ~n7078 ;
  assign y3614 = n1918 ;
  assign y3615 = ~1'b0 ;
  assign y3616 = ~n7079 ;
  assign y3617 = ~n7080 ;
  assign y3618 = ~n5443 ;
  assign y3619 = ~1'b0 ;
  assign y3620 = n7081 ;
  assign y3621 = n7084 ;
  assign y3622 = n7086 ;
  assign y3623 = ~n2146 ;
  assign y3624 = ~n7088 ;
  assign y3625 = ~1'b0 ;
  assign y3626 = ~n7089 ;
  assign y3627 = n6934 ;
  assign y3628 = ~1'b0 ;
  assign y3629 = 1'b0 ;
  assign y3630 = ~1'b0 ;
  assign y3631 = ~n7093 ;
  assign y3632 = ~1'b0 ;
  assign y3633 = n7095 ;
  assign y3634 = n7104 ;
  assign y3635 = ~n7106 ;
  assign y3636 = n7107 ;
  assign y3637 = ~n7108 ;
  assign y3638 = n7118 ;
  assign y3639 = ~1'b0 ;
  assign y3640 = 1'b0 ;
  assign y3641 = ~1'b0 ;
  assign y3642 = n4468 ;
  assign y3643 = ~1'b0 ;
  assign y3644 = ~1'b0 ;
  assign y3645 = ~1'b0 ;
  assign y3646 = 1'b0 ;
  assign y3647 = ~1'b0 ;
  assign y3648 = n7121 ;
  assign y3649 = ~n7124 ;
  assign y3650 = n7125 ;
  assign y3651 = ~1'b0 ;
  assign y3652 = n7127 ;
  assign y3653 = ~1'b0 ;
  assign y3654 = ~n7128 ;
  assign y3655 = ~1'b0 ;
  assign y3656 = ~1'b0 ;
  assign y3657 = ~1'b0 ;
  assign y3658 = ~n4094 ;
  assign y3659 = ~n7131 ;
  assign y3660 = ~1'b0 ;
  assign y3661 = n7132 ;
  assign y3662 = n7133 ;
  assign y3663 = ~n2381 ;
  assign y3664 = ~n7135 ;
  assign y3665 = n7136 ;
  assign y3666 = ~n7139 ;
  assign y3667 = ~n7140 ;
  assign y3668 = ~n7142 ;
  assign y3669 = ~1'b0 ;
  assign y3670 = ~n7143 ;
  assign y3671 = n7146 ;
  assign y3672 = ~n7150 ;
  assign y3673 = ~1'b0 ;
  assign y3674 = ~n7151 ;
  assign y3675 = ~n7153 ;
  assign y3676 = n7154 ;
  assign y3677 = n7160 ;
  assign y3678 = n269 ;
  assign y3679 = 1'b0 ;
  assign y3680 = n7164 ;
  assign y3681 = ~n7165 ;
  assign y3682 = ~n7169 ;
  assign y3683 = ~n7172 ;
  assign y3684 = ~n7175 ;
  assign y3685 = n7182 ;
  assign y3686 = n7189 ;
  assign y3687 = ~n7195 ;
  assign y3688 = n7197 ;
  assign y3689 = n7199 ;
  assign y3690 = ~n7200 ;
  assign y3691 = n7207 ;
  assign y3692 = ~1'b0 ;
  assign y3693 = n7209 ;
  assign y3694 = ~n7232 ;
  assign y3695 = n7234 ;
  assign y3696 = n7236 ;
  assign y3697 = n7238 ;
  assign y3698 = n7239 ;
  assign y3699 = ~1'b0 ;
  assign y3700 = n7240 ;
  assign y3701 = ~n7242 ;
  assign y3702 = ~1'b0 ;
  assign y3703 = n7243 ;
  assign y3704 = ~1'b0 ;
  assign y3705 = n7248 ;
  assign y3706 = n7254 ;
  assign y3707 = n7257 ;
  assign y3708 = ~n7262 ;
  assign y3709 = ~1'b0 ;
  assign y3710 = ~1'b0 ;
  assign y3711 = n5328 ;
  assign y3712 = ~n7265 ;
  assign y3713 = n7268 ;
  assign y3714 = ~1'b0 ;
  assign y3715 = n7269 ;
  assign y3716 = ~n7272 ;
  assign y3717 = n7275 ;
  assign y3718 = ~n7276 ;
  assign y3719 = n5399 ;
  assign y3720 = n7278 ;
  assign y3721 = ~n7287 ;
  assign y3722 = 1'b0 ;
  assign y3723 = ~n7288 ;
  assign y3724 = 1'b0 ;
  assign y3725 = ~n7289 ;
  assign y3726 = ~n7292 ;
  assign y3727 = 1'b0 ;
  assign y3728 = ~n7293 ;
  assign y3729 = n7294 ;
  assign y3730 = ~1'b0 ;
  assign y3731 = ~1'b0 ;
  assign y3732 = n7297 ;
  assign y3733 = n7300 ;
  assign y3734 = ~n7302 ;
  assign y3735 = ~n7305 ;
  assign y3736 = ~n7307 ;
  assign y3737 = n7308 ;
  assign y3738 = ~1'b0 ;
  assign y3739 = ~1'b0 ;
  assign y3740 = ~n7309 ;
  assign y3741 = ~n1897 ;
  assign y3742 = n3962 ;
  assign y3743 = ~n7313 ;
  assign y3744 = n7314 ;
  assign y3745 = ~n7317 ;
  assign y3746 = n7321 ;
  assign y3747 = ~1'b0 ;
  assign y3748 = ~n1066 ;
  assign y3749 = ~1'b0 ;
  assign y3750 = n7324 ;
  assign y3751 = n4720 ;
  assign y3752 = n7333 ;
  assign y3753 = n7347 ;
  assign y3754 = ~1'b0 ;
  assign y3755 = ~1'b0 ;
  assign y3756 = n7348 ;
  assign y3757 = ~1'b0 ;
  assign y3758 = ~n7349 ;
  assign y3759 = n7350 ;
  assign y3760 = n7351 ;
  assign y3761 = ~1'b0 ;
  assign y3762 = 1'b0 ;
  assign y3763 = ~n7360 ;
  assign y3764 = ~n7366 ;
  assign y3765 = n7367 ;
  assign y3766 = ~n7368 ;
  assign y3767 = ~n2989 ;
  assign y3768 = ~n7369 ;
  assign y3769 = ~n7370 ;
  assign y3770 = ~1'b0 ;
  assign y3771 = ~n1853 ;
  assign y3772 = ~n7374 ;
  assign y3773 = n7375 ;
  assign y3774 = n7376 ;
  assign y3775 = n7379 ;
  assign y3776 = ~1'b0 ;
  assign y3777 = ~1'b0 ;
  assign y3778 = ~n7382 ;
  assign y3779 = ~n2532 ;
  assign y3780 = n7383 ;
  assign y3781 = ~n7388 ;
  assign y3782 = n7389 ;
  assign y3783 = ~1'b0 ;
  assign y3784 = n7391 ;
  assign y3785 = ~1'b0 ;
  assign y3786 = n7394 ;
  assign y3787 = n7397 ;
  assign y3788 = n7400 ;
  assign y3789 = ~1'b0 ;
  assign y3790 = n7403 ;
  assign y3791 = ~n7404 ;
  assign y3792 = n7405 ;
  assign y3793 = n7410 ;
  assign y3794 = ~1'b0 ;
  assign y3795 = n7414 ;
  assign y3796 = n7418 ;
  assign y3797 = n5685 ;
  assign y3798 = ~1'b0 ;
  assign y3799 = n7422 ;
  assign y3800 = ~1'b0 ;
  assign y3801 = n7423 ;
  assign y3802 = ~1'b0 ;
  assign y3803 = n7427 ;
  assign y3804 = ~n7430 ;
  assign y3805 = ~1'b0 ;
  assign y3806 = ~n7441 ;
  assign y3807 = n7442 ;
  assign y3808 = ~1'b0 ;
  assign y3809 = ~1'b0 ;
  assign y3810 = ~n7446 ;
  assign y3811 = n7447 ;
  assign y3812 = n7451 ;
  assign y3813 = ~n7454 ;
  assign y3814 = ~n7455 ;
  assign y3815 = n7457 ;
  assign y3816 = ~1'b0 ;
  assign y3817 = n7458 ;
  assign y3818 = ~n7459 ;
  assign y3819 = n7464 ;
  assign y3820 = ~n7466 ;
  assign y3821 = ~n7467 ;
  assign y3822 = ~1'b0 ;
  assign y3823 = ~n7475 ;
  assign y3824 = ~n7477 ;
  assign y3825 = ~1'b0 ;
  assign y3826 = ~1'b0 ;
  assign y3827 = ~1'b0 ;
  assign y3828 = 1'b0 ;
  assign y3829 = ~n7479 ;
  assign y3830 = ~1'b0 ;
  assign y3831 = ~n7480 ;
  assign y3832 = ~n188 ;
  assign y3833 = ~1'b0 ;
  assign y3834 = ~n7482 ;
  assign y3835 = ~1'b0 ;
  assign y3836 = ~n7484 ;
  assign y3837 = n7485 ;
  assign y3838 = n7488 ;
  assign y3839 = ~n7491 ;
  assign y3840 = n7492 ;
  assign y3841 = n7494 ;
  assign y3842 = ~n7497 ;
  assign y3843 = ~n7498 ;
  assign y3844 = n7499 ;
  assign y3845 = ~1'b0 ;
  assign y3846 = ~n7500 ;
  assign y3847 = ~n7501 ;
  assign y3848 = ~n7507 ;
  assign y3849 = ~1'b0 ;
  assign y3850 = ~n7518 ;
  assign y3851 = ~n7521 ;
  assign y3852 = ~1'b0 ;
  assign y3853 = ~1'b0 ;
  assign y3854 = ~1'b0 ;
  assign y3855 = n7522 ;
  assign y3856 = n7523 ;
  assign y3857 = n7528 ;
  assign y3858 = ~1'b0 ;
  assign y3859 = n5755 ;
  assign y3860 = ~1'b0 ;
  assign y3861 = ~1'b0 ;
  assign y3862 = ~n7529 ;
  assign y3863 = ~n7531 ;
  assign y3864 = n7532 ;
  assign y3865 = n7537 ;
  assign y3866 = ~1'b0 ;
  assign y3867 = n7538 ;
  assign y3868 = ~n7542 ;
  assign y3869 = ~n7545 ;
  assign y3870 = ~n7546 ;
  assign y3871 = n7549 ;
  assign y3872 = ~1'b0 ;
  assign y3873 = n7554 ;
  assign y3874 = ~n7558 ;
  assign y3875 = ~1'b0 ;
  assign y3876 = n7564 ;
  assign y3877 = ~n7565 ;
  assign y3878 = ~n7567 ;
  assign y3879 = ~n7568 ;
  assign y3880 = ~n1771 ;
  assign y3881 = ~n7570 ;
  assign y3882 = ~1'b0 ;
  assign y3883 = ~1'b0 ;
  assign y3884 = n7578 ;
  assign y3885 = n7581 ;
  assign y3886 = n7582 ;
  assign y3887 = n7583 ;
  assign y3888 = ~1'b0 ;
  assign y3889 = ~n7586 ;
  assign y3890 = n7589 ;
  assign y3891 = n7590 ;
  assign y3892 = ~n7593 ;
  assign y3893 = n459 ;
  assign y3894 = ~1'b0 ;
  assign y3895 = ~n7598 ;
  assign y3896 = ~1'b0 ;
  assign y3897 = ~1'b0 ;
  assign y3898 = ~1'b0 ;
  assign y3899 = ~1'b0 ;
  assign y3900 = ~n7606 ;
  assign y3901 = ~n7607 ;
  assign y3902 = ~n7611 ;
  assign y3903 = n7613 ;
  assign y3904 = n7616 ;
  assign y3905 = ~n7618 ;
  assign y3906 = n5381 ;
  assign y3907 = ~n7624 ;
  assign y3908 = n7631 ;
  assign y3909 = n7632 ;
  assign y3910 = ~n7633 ;
  assign y3911 = ~n7635 ;
  assign y3912 = ~n7639 ;
  assign y3913 = ~n7643 ;
  assign y3914 = n7645 ;
  assign y3915 = ~1'b0 ;
  assign y3916 = ~1'b0 ;
  assign y3917 = ~1'b0 ;
  assign y3918 = n7647 ;
  assign y3919 = n7652 ;
  assign y3920 = n7656 ;
  assign y3921 = n7658 ;
  assign y3922 = n7665 ;
  assign y3923 = ~1'b0 ;
  assign y3924 = ~n7666 ;
  assign y3925 = ~1'b0 ;
  assign y3926 = ~n7669 ;
  assign y3927 = n7670 ;
  assign y3928 = ~1'b0 ;
  assign y3929 = ~n7673 ;
  assign y3930 = n7676 ;
  assign y3931 = ~1'b0 ;
  assign y3932 = ~n7682 ;
  assign y3933 = n7686 ;
  assign y3934 = n7690 ;
  assign y3935 = ~n7691 ;
  assign y3936 = n7693 ;
  assign y3937 = ~1'b0 ;
  assign y3938 = ~n7695 ;
  assign y3939 = n7699 ;
  assign y3940 = ~n7702 ;
  assign y3941 = n7704 ;
  assign y3942 = n7705 ;
  assign y3943 = ~1'b0 ;
  assign y3944 = ~n7707 ;
  assign y3945 = ~n7710 ;
  assign y3946 = ~1'b0 ;
  assign y3947 = ~n7713 ;
  assign y3948 = n7720 ;
  assign y3949 = ~n7721 ;
  assign y3950 = 1'b0 ;
  assign y3951 = ~n7724 ;
  assign y3952 = n7726 ;
  assign y3953 = ~1'b0 ;
  assign y3954 = n3547 ;
  assign y3955 = ~1'b0 ;
  assign y3956 = ~n7730 ;
  assign y3957 = n7731 ;
  assign y3958 = n7734 ;
  assign y3959 = ~1'b0 ;
  assign y3960 = ~n7735 ;
  assign y3961 = n7737 ;
  assign y3962 = n7746 ;
  assign y3963 = ~n7752 ;
  assign y3964 = ~n7753 ;
  assign y3965 = n7755 ;
  assign y3966 = n7756 ;
  assign y3967 = n7758 ;
  assign y3968 = ~1'b0 ;
  assign y3969 = n6878 ;
  assign y3970 = ~1'b0 ;
  assign y3971 = n7761 ;
  assign y3972 = n7768 ;
  assign y3973 = ~n7773 ;
  assign y3974 = ~n7776 ;
  assign y3975 = ~n7779 ;
  assign y3976 = ~n7786 ;
  assign y3977 = ~n3050 ;
  assign y3978 = 1'b0 ;
  assign y3979 = ~1'b0 ;
  assign y3980 = ~1'b0 ;
  assign y3981 = n7788 ;
  assign y3982 = n7791 ;
  assign y3983 = n3349 ;
  assign y3984 = n7793 ;
  assign y3985 = n7795 ;
  assign y3986 = ~n7802 ;
  assign y3987 = n7806 ;
  assign y3988 = 1'b0 ;
  assign y3989 = ~1'b0 ;
  assign y3990 = ~n7809 ;
  assign y3991 = ~n7814 ;
  assign y3992 = n7816 ;
  assign y3993 = n7822 ;
  assign y3994 = ~1'b0 ;
  assign y3995 = ~n7824 ;
  assign y3996 = ~n7825 ;
  assign y3997 = ~n7827 ;
  assign y3998 = n5150 ;
  assign y3999 = ~n7829 ;
  assign y4000 = ~n7831 ;
  assign y4001 = ~n7833 ;
  assign y4002 = ~n7841 ;
  assign y4003 = n4846 ;
  assign y4004 = ~1'b0 ;
  assign y4005 = ~1'b0 ;
  assign y4006 = n7843 ;
  assign y4007 = n7844 ;
  assign y4008 = ~n7846 ;
  assign y4009 = ~n7847 ;
  assign y4010 = n7848 ;
  assign y4011 = ~1'b0 ;
  assign y4012 = ~n7850 ;
  assign y4013 = n7851 ;
  assign y4014 = ~n7855 ;
  assign y4015 = ~1'b0 ;
  assign y4016 = n3343 ;
  assign y4017 = n7857 ;
  assign y4018 = ~1'b0 ;
  assign y4019 = n6714 ;
  assign y4020 = ~n7861 ;
  assign y4021 = n7864 ;
  assign y4022 = ~1'b0 ;
  assign y4023 = ~1'b0 ;
  assign y4024 = n7871 ;
  assign y4025 = n7878 ;
  assign y4026 = n7886 ;
  assign y4027 = ~n7889 ;
  assign y4028 = ~1'b0 ;
  assign y4029 = ~n7897 ;
  assign y4030 = ~n7898 ;
  assign y4031 = n7899 ;
  assign y4032 = 1'b0 ;
  assign y4033 = n7902 ;
  assign y4034 = ~n6764 ;
  assign y4035 = ~1'b0 ;
  assign y4036 = n7906 ;
  assign y4037 = ~1'b0 ;
  assign y4038 = ~1'b0 ;
  assign y4039 = n7913 ;
  assign y4040 = n7914 ;
  assign y4041 = ~1'b0 ;
  assign y4042 = ~1'b0 ;
  assign y4043 = ~n7917 ;
  assign y4044 = n7919 ;
  assign y4045 = ~n5027 ;
  assign y4046 = ~n572 ;
  assign y4047 = ~1'b0 ;
  assign y4048 = ~1'b0 ;
  assign y4049 = n7924 ;
  assign y4050 = ~1'b0 ;
  assign y4051 = ~1'b0 ;
  assign y4052 = n7932 ;
  assign y4053 = ~n7933 ;
  assign y4054 = ~n7934 ;
  assign y4055 = n7935 ;
  assign y4056 = n7937 ;
  assign y4057 = ~1'b0 ;
  assign y4058 = ~n7939 ;
  assign y4059 = ~n7940 ;
  assign y4060 = n7941 ;
  assign y4061 = ~n7947 ;
  assign y4062 = n7951 ;
  assign y4063 = n7952 ;
  assign y4064 = ~n7953 ;
  assign y4065 = ~n7955 ;
  assign y4066 = ~n7957 ;
  assign y4067 = ~1'b0 ;
  assign y4068 = ~n3476 ;
  assign y4069 = ~1'b0 ;
  assign y4070 = ~1'b0 ;
  assign y4071 = ~n7960 ;
  assign y4072 = ~n7964 ;
  assign y4073 = ~n4632 ;
  assign y4074 = ~1'b0 ;
  assign y4075 = ~n7965 ;
  assign y4076 = ~1'b0 ;
  assign y4077 = ~n7967 ;
  assign y4078 = ~1'b0 ;
  assign y4079 = ~1'b0 ;
  assign y4080 = ~1'b0 ;
  assign y4081 = ~1'b0 ;
  assign y4082 = ~1'b0 ;
  assign y4083 = n7971 ;
  assign y4084 = ~n7977 ;
  assign y4085 = ~n7978 ;
  assign y4086 = n7981 ;
  assign y4087 = n7982 ;
  assign y4088 = ~n7984 ;
  assign y4089 = ~1'b0 ;
  assign y4090 = ~n7987 ;
  assign y4091 = n7989 ;
  assign y4092 = n7990 ;
  assign y4093 = ~n7994 ;
  assign y4094 = ~n7996 ;
  assign y4095 = ~1'b0 ;
  assign y4096 = ~n7998 ;
  assign y4097 = ~n7999 ;
  assign y4098 = ~n8003 ;
  assign y4099 = n8007 ;
  assign y4100 = n8008 ;
  assign y4101 = n8010 ;
  assign y4102 = ~1'b0 ;
  assign y4103 = ~n4679 ;
  assign y4104 = ~n8011 ;
  assign y4105 = n7604 ;
  assign y4106 = n8014 ;
  assign y4107 = ~n8018 ;
  assign y4108 = n8019 ;
  assign y4109 = ~1'b0 ;
  assign y4110 = ~n8020 ;
  assign y4111 = n8022 ;
  assign y4112 = ~n8032 ;
  assign y4113 = ~n559 ;
  assign y4114 = n8033 ;
  assign y4115 = ~n8036 ;
  assign y4116 = ~n8039 ;
  assign y4117 = ~1'b0 ;
  assign y4118 = ~n8042 ;
  assign y4119 = ~n8043 ;
  assign y4120 = ~1'b0 ;
  assign y4121 = ~1'b0 ;
  assign y4122 = n3408 ;
  assign y4123 = n8047 ;
  assign y4124 = n8049 ;
  assign y4125 = ~1'b0 ;
  assign y4126 = n8053 ;
  assign y4127 = ~n2498 ;
  assign y4128 = n8061 ;
  assign y4129 = ~n8066 ;
  assign y4130 = ~n8071 ;
  assign y4131 = ~n7627 ;
  assign y4132 = ~n8072 ;
  assign y4133 = ~1'b0 ;
  assign y4134 = ~n8076 ;
  assign y4135 = n8077 ;
  assign y4136 = ~1'b0 ;
  assign y4137 = ~n8078 ;
  assign y4138 = n8079 ;
  assign y4139 = n8089 ;
  assign y4140 = ~1'b0 ;
  assign y4141 = n8093 ;
  assign y4142 = ~n8099 ;
  assign y4143 = n2671 ;
  assign y4144 = n8100 ;
  assign y4145 = ~n8101 ;
  assign y4146 = ~1'b0 ;
  assign y4147 = n8104 ;
  assign y4148 = n8107 ;
  assign y4149 = ~n8115 ;
  assign y4150 = ~1'b0 ;
  assign y4151 = n8117 ;
  assign y4152 = n8118 ;
  assign y4153 = ~1'b0 ;
  assign y4154 = n8126 ;
  assign y4155 = ~1'b0 ;
  assign y4156 = n8127 ;
  assign y4157 = ~1'b0 ;
  assign y4158 = ~1'b0 ;
  assign y4159 = ~n8128 ;
  assign y4160 = n8129 ;
  assign y4161 = ~1'b0 ;
  assign y4162 = ~1'b0 ;
  assign y4163 = n631 ;
  assign y4164 = n8130 ;
  assign y4165 = n8134 ;
  assign y4166 = n8135 ;
  assign y4167 = 1'b0 ;
  assign y4168 = ~n8136 ;
  assign y4169 = ~n8138 ;
  assign y4170 = ~n8139 ;
  assign y4171 = ~n8141 ;
  assign y4172 = ~n8142 ;
  assign y4173 = n8147 ;
  assign y4174 = n5856 ;
  assign y4175 = ~1'b0 ;
  assign y4176 = ~n8148 ;
  assign y4177 = n8152 ;
  assign y4178 = ~n8153 ;
  assign y4179 = ~1'b0 ;
  assign y4180 = 1'b0 ;
  assign y4181 = ~n8154 ;
  assign y4182 = ~n8156 ;
  assign y4183 = 1'b0 ;
  assign y4184 = ~n3934 ;
  assign y4185 = ~n8166 ;
  assign y4186 = ~n8171 ;
  assign y4187 = ~n8173 ;
  assign y4188 = n8174 ;
  assign y4189 = ~1'b0 ;
  assign y4190 = ~1'b0 ;
  assign y4191 = ~n8183 ;
  assign y4192 = ~n8187 ;
  assign y4193 = ~n8192 ;
  assign y4194 = ~1'b0 ;
  assign y4195 = ~1'b0 ;
  assign y4196 = n8195 ;
  assign y4197 = n8198 ;
  assign y4198 = 1'b0 ;
  assign y4199 = ~1'b0 ;
  assign y4200 = n8199 ;
  assign y4201 = ~n8200 ;
  assign y4202 = ~1'b0 ;
  assign y4203 = ~n4040 ;
  assign y4204 = ~1'b0 ;
  assign y4205 = ~n8201 ;
  assign y4206 = ~n8209 ;
  assign y4207 = n8211 ;
  assign y4208 = ~n2812 ;
  assign y4209 = ~1'b0 ;
  assign y4210 = n8212 ;
  assign y4211 = n8215 ;
  assign y4212 = n8216 ;
  assign y4213 = ~1'b0 ;
  assign y4214 = ~1'b0 ;
  assign y4215 = n8219 ;
  assign y4216 = n8220 ;
  assign y4217 = n8224 ;
  assign y4218 = n5513 ;
  assign y4219 = ~n8225 ;
  assign y4220 = ~1'b0 ;
  assign y4221 = n7368 ;
  assign y4222 = ~1'b0 ;
  assign y4223 = ~n8228 ;
  assign y4224 = n8229 ;
  assign y4225 = n8236 ;
  assign y4226 = n8208 ;
  assign y4227 = n8242 ;
  assign y4228 = ~n8243 ;
  assign y4229 = ~n8244 ;
  assign y4230 = ~n8246 ;
  assign y4231 = ~n8251 ;
  assign y4232 = ~n8252 ;
  assign y4233 = ~1'b0 ;
  assign y4234 = ~1'b0 ;
  assign y4235 = ~1'b0 ;
  assign y4236 = ~1'b0 ;
  assign y4237 = ~n8253 ;
  assign y4238 = ~n8258 ;
  assign y4239 = ~1'b0 ;
  assign y4240 = ~n8259 ;
  assign y4241 = ~n3182 ;
  assign y4242 = ~1'b0 ;
  assign y4243 = ~1'b0 ;
  assign y4244 = ~1'b0 ;
  assign y4245 = ~n8262 ;
  assign y4246 = n8265 ;
  assign y4247 = ~1'b0 ;
  assign y4248 = n8267 ;
  assign y4249 = ~n8269 ;
  assign y4250 = ~n8270 ;
  assign y4251 = ~1'b0 ;
  assign y4252 = ~n400 ;
  assign y4253 = ~1'b0 ;
  assign y4254 = ~n8276 ;
  assign y4255 = ~n8277 ;
  assign y4256 = ~1'b0 ;
  assign y4257 = ~1'b0 ;
  assign y4258 = ~n8278 ;
  assign y4259 = ~1'b0 ;
  assign y4260 = ~1'b0 ;
  assign y4261 = ~1'b0 ;
  assign y4262 = ~1'b0 ;
  assign y4263 = n8281 ;
  assign y4264 = ~n8282 ;
  assign y4265 = ~1'b0 ;
  assign y4266 = n8283 ;
  assign y4267 = n8286 ;
  assign y4268 = n8288 ;
  assign y4269 = ~n8292 ;
  assign y4270 = ~1'b0 ;
  assign y4271 = 1'b0 ;
  assign y4272 = ~n8293 ;
  assign y4273 = n8296 ;
  assign y4274 = ~1'b0 ;
  assign y4275 = ~1'b0 ;
  assign y4276 = n1703 ;
  assign y4277 = n8301 ;
  assign y4278 = n8302 ;
  assign y4279 = ~n8309 ;
  assign y4280 = ~1'b0 ;
  assign y4281 = ~1'b0 ;
  assign y4282 = ~1'b0 ;
  assign y4283 = ~n8310 ;
  assign y4284 = ~n8314 ;
  assign y4285 = ~1'b0 ;
  assign y4286 = ~1'b0 ;
  assign y4287 = ~n8317 ;
  assign y4288 = ~n8321 ;
  assign y4289 = ~n8324 ;
  assign y4290 = n8326 ;
  assign y4291 = ~n8327 ;
  assign y4292 = ~n8330 ;
  assign y4293 = ~n8334 ;
  assign y4294 = ~n8341 ;
  assign y4295 = n7653 ;
  assign y4296 = ~1'b0 ;
  assign y4297 = ~1'b0 ;
  assign y4298 = n8342 ;
  assign y4299 = n8344 ;
  assign y4300 = ~n8349 ;
  assign y4301 = n8350 ;
  assign y4302 = n8351 ;
  assign y4303 = ~1'b0 ;
  assign y4304 = n8354 ;
  assign y4305 = ~1'b0 ;
  assign y4306 = n8357 ;
  assign y4307 = n5492 ;
  assign y4308 = n8359 ;
  assign y4309 = ~1'b0 ;
  assign y4310 = ~n8362 ;
  assign y4311 = n8366 ;
  assign y4312 = n6358 ;
  assign y4313 = n8367 ;
  assign y4314 = ~n8372 ;
  assign y4315 = ~n8373 ;
  assign y4316 = ~n8378 ;
  assign y4317 = ~1'b0 ;
  assign y4318 = ~n8380 ;
  assign y4319 = n8381 ;
  assign y4320 = ~n8383 ;
  assign y4321 = ~n8392 ;
  assign y4322 = ~1'b0 ;
  assign y4323 = ~1'b0 ;
  assign y4324 = ~n8393 ;
  assign y4325 = ~1'b0 ;
  assign y4326 = n8396 ;
  assign y4327 = ~n8404 ;
  assign y4328 = ~1'b0 ;
  assign y4329 = ~1'b0 ;
  assign y4330 = n8407 ;
  assign y4331 = ~1'b0 ;
  assign y4332 = ~1'b0 ;
  assign y4333 = 1'b0 ;
  assign y4334 = n8408 ;
  assign y4335 = ~1'b0 ;
  assign y4336 = ~n8411 ;
  assign y4337 = ~1'b0 ;
  assign y4338 = ~1'b0 ;
  assign y4339 = n8412 ;
  assign y4340 = n8413 ;
  assign y4341 = n8416 ;
  assign y4342 = ~n8419 ;
  assign y4343 = ~1'b0 ;
  assign y4344 = n8423 ;
  assign y4345 = n8426 ;
  assign y4346 = n8427 ;
  assign y4347 = ~n8433 ;
  assign y4348 = ~n8435 ;
  assign y4349 = n8438 ;
  assign y4350 = 1'b0 ;
  assign y4351 = n8441 ;
  assign y4352 = ~n8445 ;
  assign y4353 = ~1'b0 ;
  assign y4354 = ~1'b0 ;
  assign y4355 = ~n8446 ;
  assign y4356 = n874 ;
  assign y4357 = n8449 ;
  assign y4358 = n8450 ;
  assign y4359 = n8452 ;
  assign y4360 = ~n8454 ;
  assign y4361 = n8457 ;
  assign y4362 = ~1'b0 ;
  assign y4363 = 1'b0 ;
  assign y4364 = ~n150 ;
  assign y4365 = ~n8461 ;
  assign y4366 = ~n7825 ;
  assign y4367 = n8463 ;
  assign y4368 = n8468 ;
  assign y4369 = ~n8476 ;
  assign y4370 = ~1'b0 ;
  assign y4371 = ~n8481 ;
  assign y4372 = ~1'b0 ;
  assign y4373 = n1387 ;
  assign y4374 = ~n8485 ;
  assign y4375 = ~1'b0 ;
  assign y4376 = ~1'b0 ;
  assign y4377 = ~1'b0 ;
  assign y4378 = ~n8489 ;
  assign y4379 = ~n8490 ;
  assign y4380 = ~n8491 ;
  assign y4381 = ~n506 ;
  assign y4382 = ~1'b0 ;
  assign y4383 = ~n4267 ;
  assign y4384 = ~1'b0 ;
  assign y4385 = n3851 ;
  assign y4386 = n8494 ;
  assign y4387 = ~n8502 ;
  assign y4388 = n8503 ;
  assign y4389 = ~n8506 ;
  assign y4390 = n8510 ;
  assign y4391 = 1'b0 ;
  assign y4392 = n8514 ;
  assign y4393 = ~1'b0 ;
  assign y4394 = n8515 ;
  assign y4395 = ~1'b0 ;
  assign y4396 = ~1'b0 ;
  assign y4397 = 1'b0 ;
  assign y4398 = n8518 ;
  assign y4399 = n8521 ;
  assign y4400 = ~1'b0 ;
  assign y4401 = n8525 ;
  assign y4402 = ~1'b0 ;
  assign y4403 = n7718 ;
  assign y4404 = ~n8526 ;
  assign y4405 = n8527 ;
  assign y4406 = ~1'b0 ;
  assign y4407 = n8529 ;
  assign y4408 = n8532 ;
  assign y4409 = ~1'b0 ;
  assign y4410 = ~1'b0 ;
  assign y4411 = ~n8536 ;
  assign y4412 = ~n8542 ;
  assign y4413 = n8543 ;
  assign y4414 = ~1'b0 ;
  assign y4415 = n8547 ;
  assign y4416 = ~1'b0 ;
  assign y4417 = ~1'b0 ;
  assign y4418 = ~1'b0 ;
  assign y4419 = n8548 ;
  assign y4420 = 1'b0 ;
  assign y4421 = ~1'b0 ;
  assign y4422 = ~n8551 ;
  assign y4423 = ~1'b0 ;
  assign y4424 = n8552 ;
  assign y4425 = ~1'b0 ;
  assign y4426 = ~n8553 ;
  assign y4427 = ~n8554 ;
  assign y4428 = ~n8555 ;
  assign y4429 = ~1'b0 ;
  assign y4430 = ~n8563 ;
  assign y4431 = ~1'b0 ;
  assign y4432 = ~n8565 ;
  assign y4433 = ~1'b0 ;
  assign y4434 = ~1'b0 ;
  assign y4435 = ~n8566 ;
  assign y4436 = n8568 ;
  assign y4437 = ~n8573 ;
  assign y4438 = n8584 ;
  assign y4439 = n1802 ;
  assign y4440 = ~n8589 ;
  assign y4441 = n8592 ;
  assign y4442 = ~1'b0 ;
  assign y4443 = ~1'b0 ;
  assign y4444 = ~1'b0 ;
  assign y4445 = ~n8594 ;
  assign y4446 = ~1'b0 ;
  assign y4447 = ~1'b0 ;
  assign y4448 = n8595 ;
  assign y4449 = ~n8599 ;
  assign y4450 = ~n8600 ;
  assign y4451 = n8603 ;
  assign y4452 = ~n8607 ;
  assign y4453 = n8611 ;
  assign y4454 = ~1'b0 ;
  assign y4455 = ~1'b0 ;
  assign y4456 = n8613 ;
  assign y4457 = ~1'b0 ;
  assign y4458 = ~n8614 ;
  assign y4459 = ~1'b0 ;
  assign y4460 = n8618 ;
  assign y4461 = ~1'b0 ;
  assign y4462 = ~n8620 ;
  assign y4463 = n8621 ;
  assign y4464 = ~n8624 ;
  assign y4465 = n8629 ;
  assign y4466 = ~1'b0 ;
  assign y4467 = n8631 ;
  assign y4468 = n8637 ;
  assign y4469 = ~1'b0 ;
  assign y4470 = n8144 ;
  assign y4471 = ~n8640 ;
  assign y4472 = n8646 ;
  assign y4473 = ~1'b0 ;
  assign y4474 = ~1'b0 ;
  assign y4475 = 1'b0 ;
  assign y4476 = n8650 ;
  assign y4477 = n8656 ;
  assign y4478 = n8663 ;
  assign y4479 = 1'b0 ;
  assign y4480 = ~n8665 ;
  assign y4481 = n8667 ;
  assign y4482 = ~1'b0 ;
  assign y4483 = n8672 ;
  assign y4484 = n2346 ;
  assign y4485 = n8675 ;
  assign y4486 = ~n8677 ;
  assign y4487 = n8681 ;
  assign y4488 = ~1'b0 ;
  assign y4489 = ~n8684 ;
  assign y4490 = n8686 ;
  assign y4491 = ~n8688 ;
  assign y4492 = n8697 ;
  assign y4493 = n8704 ;
  assign y4494 = ~n8705 ;
  assign y4495 = ~n6586 ;
  assign y4496 = 1'b0 ;
  assign y4497 = ~1'b0 ;
  assign y4498 = ~1'b0 ;
  assign y4499 = ~n8708 ;
  assign y4500 = ~n8710 ;
  assign y4501 = n8712 ;
  assign y4502 = ~n8715 ;
  assign y4503 = n8716 ;
  assign y4504 = n8717 ;
  assign y4505 = ~1'b0 ;
  assign y4506 = ~n8720 ;
  assign y4507 = ~n8721 ;
  assign y4508 = n8727 ;
  assign y4509 = ~n8734 ;
  assign y4510 = ~1'b0 ;
  assign y4511 = ~n8735 ;
  assign y4512 = ~1'b0 ;
  assign y4513 = n421 ;
  assign y4514 = n8737 ;
  assign y4515 = n8741 ;
  assign y4516 = n8747 ;
  assign y4517 = n4046 ;
  assign y4518 = n8749 ;
  assign y4519 = ~1'b0 ;
  assign y4520 = ~1'b0 ;
  assign y4521 = ~n8750 ;
  assign y4522 = n8754 ;
  assign y4523 = ~n8758 ;
  assign y4524 = ~n8759 ;
  assign y4525 = n8763 ;
  assign y4526 = ~1'b0 ;
  assign y4527 = n8766 ;
  assign y4528 = ~1'b0 ;
  assign y4529 = n8774 ;
  assign y4530 = n8781 ;
  assign y4531 = n8782 ;
  assign y4532 = ~n2649 ;
  assign y4533 = ~n8784 ;
  assign y4534 = n8788 ;
  assign y4535 = ~1'b0 ;
  assign y4536 = ~1'b0 ;
  assign y4537 = ~n8789 ;
  assign y4538 = ~1'b0 ;
  assign y4539 = n8797 ;
  assign y4540 = ~n8798 ;
  assign y4541 = ~n8802 ;
  assign y4542 = n8806 ;
  assign y4543 = ~1'b0 ;
  assign y4544 = ~1'b0 ;
  assign y4545 = n8807 ;
  assign y4546 = ~n7804 ;
  assign y4547 = n8812 ;
  assign y4548 = ~1'b0 ;
  assign y4549 = n8817 ;
  assign y4550 = ~1'b0 ;
  assign y4551 = n8823 ;
  assign y4552 = ~1'b0 ;
  assign y4553 = n8824 ;
  assign y4554 = n8826 ;
  assign y4555 = ~1'b0 ;
  assign y4556 = ~1'b0 ;
  assign y4557 = ~1'b0 ;
  assign y4558 = ~n8830 ;
  assign y4559 = n8834 ;
  assign y4560 = n8836 ;
  assign y4561 = ~n8838 ;
  assign y4562 = 1'b0 ;
  assign y4563 = 1'b0 ;
  assign y4564 = ~n8842 ;
  assign y4565 = ~1'b0 ;
  assign y4566 = n8844 ;
  assign y4567 = ~1'b0 ;
  assign y4568 = ~1'b0 ;
  assign y4569 = ~1'b0 ;
  assign y4570 = ~n5562 ;
  assign y4571 = n8845 ;
  assign y4572 = ~n8850 ;
  assign y4573 = ~1'b0 ;
  assign y4574 = 1'b0 ;
  assign y4575 = n8860 ;
  assign y4576 = ~n8862 ;
  assign y4577 = n8871 ;
  assign y4578 = ~1'b0 ;
  assign y4579 = ~1'b0 ;
  assign y4580 = ~n8876 ;
  assign y4581 = ~n8878 ;
  assign y4582 = n5982 ;
  assign y4583 = n8883 ;
  assign y4584 = ~1'b0 ;
  assign y4585 = ~1'b0 ;
  assign y4586 = n8884 ;
  assign y4587 = ~1'b0 ;
  assign y4588 = n8886 ;
  assign y4589 = ~n8891 ;
  assign y4590 = ~n8893 ;
  assign y4591 = ~n8898 ;
  assign y4592 = ~n8903 ;
  assign y4593 = ~n8905 ;
  assign y4594 = ~1'b0 ;
  assign y4595 = ~n8906 ;
  assign y4596 = n8907 ;
  assign y4597 = n8913 ;
  assign y4598 = ~n8918 ;
  assign y4599 = ~n8919 ;
  assign y4600 = n8920 ;
  assign y4601 = n8924 ;
  assign y4602 = ~1'b0 ;
  assign y4603 = n1983 ;
  assign y4604 = ~1'b0 ;
  assign y4605 = ~1'b0 ;
  assign y4606 = n8934 ;
  assign y4607 = ~1'b0 ;
  assign y4608 = ~1'b0 ;
  assign y4609 = ~1'b0 ;
  assign y4610 = ~n8937 ;
  assign y4611 = n8943 ;
  assign y4612 = n3472 ;
  assign y4613 = ~1'b0 ;
  assign y4614 = n8945 ;
  assign y4615 = ~1'b0 ;
  assign y4616 = n8946 ;
  assign y4617 = ~n8950 ;
  assign y4618 = ~1'b0 ;
  assign y4619 = ~n8951 ;
  assign y4620 = n8952 ;
  assign y4621 = n8954 ;
  assign y4622 = n8957 ;
  assign y4623 = ~1'b0 ;
  assign y4624 = ~n8958 ;
  assign y4625 = ~1'b0 ;
  assign y4626 = n8959 ;
  assign y4627 = ~n8962 ;
  assign y4628 = ~n8963 ;
  assign y4629 = ~1'b0 ;
  assign y4630 = n8965 ;
  assign y4631 = ~n8971 ;
  assign y4632 = ~1'b0 ;
  assign y4633 = ~n8972 ;
  assign y4634 = ~1'b0 ;
  assign y4635 = ~n8974 ;
  assign y4636 = ~n8977 ;
  assign y4637 = n8978 ;
  assign y4638 = ~1'b0 ;
  assign y4639 = ~n8980 ;
  assign y4640 = n4636 ;
  assign y4641 = ~1'b0 ;
  assign y4642 = ~1'b0 ;
  assign y4643 = ~1'b0 ;
  assign y4644 = n8981 ;
  assign y4645 = n564 ;
  assign y4646 = n8991 ;
  assign y4647 = n5684 ;
  assign y4648 = ~n8993 ;
  assign y4649 = ~n8997 ;
  assign y4650 = n8998 ;
  assign y4651 = n9000 ;
  assign y4652 = ~n9006 ;
  assign y4653 = ~n9008 ;
  assign y4654 = ~n9009 ;
  assign y4655 = ~1'b0 ;
  assign y4656 = n4408 ;
  assign y4657 = ~n9014 ;
  assign y4658 = ~n9018 ;
  assign y4659 = n9022 ;
  assign y4660 = 1'b0 ;
  assign y4661 = ~1'b0 ;
  assign y4662 = n9024 ;
  assign y4663 = ~1'b0 ;
  assign y4664 = ~1'b0 ;
  assign y4665 = ~n9029 ;
  assign y4666 = n9030 ;
  assign y4667 = ~n9031 ;
  assign y4668 = ~1'b0 ;
  assign y4669 = n9033 ;
  assign y4670 = ~1'b0 ;
  assign y4671 = n5501 ;
  assign y4672 = n9036 ;
  assign y4673 = n9038 ;
  assign y4674 = ~n9041 ;
  assign y4675 = ~1'b0 ;
  assign y4676 = n9043 ;
  assign y4677 = n9044 ;
  assign y4678 = ~n9046 ;
  assign y4679 = ~n9047 ;
  assign y4680 = 1'b0 ;
  assign y4681 = ~n7177 ;
  assign y4682 = n9048 ;
  assign y4683 = n9051 ;
  assign y4684 = ~1'b0 ;
  assign y4685 = 1'b0 ;
  assign y4686 = n9053 ;
  assign y4687 = n9058 ;
  assign y4688 = n9059 ;
  assign y4689 = ~n9060 ;
  assign y4690 = n9062 ;
  assign y4691 = ~1'b0 ;
  assign y4692 = n9065 ;
  assign y4693 = n9069 ;
  assign y4694 = n9070 ;
  assign y4695 = ~n9074 ;
  assign y4696 = ~n1914 ;
  assign y4697 = ~1'b0 ;
  assign y4698 = n9076 ;
  assign y4699 = ~1'b0 ;
  assign y4700 = n9077 ;
  assign y4701 = n9083 ;
  assign y4702 = ~n9084 ;
  assign y4703 = ~1'b0 ;
  assign y4704 = ~n7285 ;
  assign y4705 = ~1'b0 ;
  assign y4706 = ~n9085 ;
  assign y4707 = ~1'b0 ;
  assign y4708 = ~n5973 ;
  assign y4709 = n9086 ;
  assign y4710 = ~1'b0 ;
  assign y4711 = ~n9089 ;
  assign y4712 = ~1'b0 ;
  assign y4713 = n9091 ;
  assign y4714 = n9094 ;
  assign y4715 = ~n8376 ;
  assign y4716 = n9095 ;
  assign y4717 = ~1'b0 ;
  assign y4718 = ~n9098 ;
  assign y4719 = ~n9106 ;
  assign y4720 = ~n9107 ;
  assign y4721 = n9111 ;
  assign y4722 = ~n9126 ;
  assign y4723 = ~n9135 ;
  assign y4724 = n9137 ;
  assign y4725 = ~n9140 ;
  assign y4726 = n9143 ;
  assign y4727 = n9146 ;
  assign y4728 = ~n9148 ;
  assign y4729 = ~1'b0 ;
  assign y4730 = ~1'b0 ;
  assign y4731 = ~1'b0 ;
  assign y4732 = n9165 ;
  assign y4733 = ~n56 ;
  assign y4734 = ~n9169 ;
  assign y4735 = ~n9170 ;
  assign y4736 = 1'b0 ;
  assign y4737 = ~1'b0 ;
  assign y4738 = ~n9173 ;
  assign y4739 = ~n8091 ;
  assign y4740 = n3225 ;
  assign y4741 = ~n9177 ;
  assign y4742 = ~n3060 ;
  assign y4743 = ~n3974 ;
  assign y4744 = ~1'b0 ;
  assign y4745 = ~1'b0 ;
  assign y4746 = ~1'b0 ;
  assign y4747 = ~1'b0 ;
  assign y4748 = n9178 ;
  assign y4749 = ~n9180 ;
  assign y4750 = n9182 ;
  assign y4751 = ~1'b0 ;
  assign y4752 = n5662 ;
  assign y4753 = ~1'b0 ;
  assign y4754 = 1'b0 ;
  assign y4755 = ~1'b0 ;
  assign y4756 = n9184 ;
  assign y4757 = n9191 ;
  assign y4758 = n9192 ;
  assign y4759 = n9195 ;
  assign y4760 = n9196 ;
  assign y4761 = n9201 ;
  assign y4762 = n9203 ;
  assign y4763 = n9205 ;
  assign y4764 = 1'b0 ;
  assign y4765 = n9207 ;
  assign y4766 = n9208 ;
  assign y4767 = ~1'b0 ;
  assign y4768 = ~n9212 ;
  assign y4769 = ~n9215 ;
  assign y4770 = n9216 ;
  assign y4771 = 1'b0 ;
  assign y4772 = n9220 ;
  assign y4773 = n9225 ;
  assign y4774 = n9227 ;
  assign y4775 = ~n9232 ;
  assign y4776 = ~1'b0 ;
  assign y4777 = n9238 ;
  assign y4778 = ~n9239 ;
  assign y4779 = ~n9241 ;
  assign y4780 = ~1'b0 ;
  assign y4781 = ~n9244 ;
  assign y4782 = ~1'b0 ;
  assign y4783 = n4075 ;
  assign y4784 = ~1'b0 ;
  assign y4785 = n9245 ;
  assign y4786 = ~n9250 ;
  assign y4787 = n9251 ;
  assign y4788 = n9253 ;
  assign y4789 = ~n9254 ;
  assign y4790 = n9256 ;
  assign y4791 = ~n9258 ;
  assign y4792 = ~n9260 ;
  assign y4793 = ~1'b0 ;
  assign y4794 = ~1'b0 ;
  assign y4795 = n9263 ;
  assign y4796 = ~n9266 ;
  assign y4797 = n9267 ;
  assign y4798 = n9268 ;
  assign y4799 = ~1'b0 ;
  assign y4800 = n9269 ;
  assign y4801 = 1'b0 ;
  assign y4802 = n9273 ;
  assign y4803 = n9276 ;
  assign y4804 = ~n9282 ;
  assign y4805 = n2309 ;
  assign y4806 = 1'b0 ;
  assign y4807 = ~n9284 ;
  assign y4808 = ~n9287 ;
  assign y4809 = ~1'b0 ;
  assign y4810 = ~1'b0 ;
  assign y4811 = n9288 ;
  assign y4812 = ~n9290 ;
  assign y4813 = ~n9292 ;
  assign y4814 = ~n9307 ;
  assign y4815 = ~1'b0 ;
  assign y4816 = n9314 ;
  assign y4817 = n9316 ;
  assign y4818 = n3660 ;
  assign y4819 = ~1'b0 ;
  assign y4820 = ~n9317 ;
  assign y4821 = ~1'b0 ;
  assign y4822 = ~n9323 ;
  assign y4823 = ~n9325 ;
  assign y4824 = n9326 ;
  assign y4825 = ~n9330 ;
  assign y4826 = n9334 ;
  assign y4827 = ~1'b0 ;
  assign y4828 = ~1'b0 ;
  assign y4829 = n9335 ;
  assign y4830 = n9336 ;
  assign y4831 = n9337 ;
  assign y4832 = n9338 ;
  assign y4833 = 1'b0 ;
  assign y4834 = n9339 ;
  assign y4835 = ~n9341 ;
  assign y4836 = ~1'b0 ;
  assign y4837 = ~1'b0 ;
  assign y4838 = ~n9344 ;
  assign y4839 = n9353 ;
  assign y4840 = ~n9356 ;
  assign y4841 = ~n9363 ;
  assign y4842 = ~n9364 ;
  assign y4843 = ~n9366 ;
  assign y4844 = n9368 ;
  assign y4845 = ~n9369 ;
  assign y4846 = n9376 ;
  assign y4847 = n9378 ;
  assign y4848 = ~n9380 ;
  assign y4849 = ~n9381 ;
  assign y4850 = n3035 ;
  assign y4851 = n9386 ;
  assign y4852 = ~n9390 ;
  assign y4853 = ~n9393 ;
  assign y4854 = ~n9399 ;
  assign y4855 = ~1'b0 ;
  assign y4856 = ~1'b0 ;
  assign y4857 = n4082 ;
  assign y4858 = n9404 ;
  assign y4859 = ~n6808 ;
  assign y4860 = ~n9411 ;
  assign y4861 = ~n9414 ;
  assign y4862 = n9417 ;
  assign y4863 = n9419 ;
  assign y4864 = ~n9421 ;
  assign y4865 = ~n9426 ;
  assign y4866 = ~1'b0 ;
  assign y4867 = n9427 ;
  assign y4868 = n9428 ;
  assign y4869 = ~n9430 ;
  assign y4870 = ~n9434 ;
  assign y4871 = n9437 ;
  assign y4872 = n9439 ;
  assign y4873 = n9440 ;
  assign y4874 = ~1'b0 ;
  assign y4875 = ~n9441 ;
  assign y4876 = ~1'b0 ;
  assign y4877 = ~1'b0 ;
  assign y4878 = n9442 ;
  assign y4879 = n9445 ;
  assign y4880 = ~1'b0 ;
  assign y4881 = ~1'b0 ;
  assign y4882 = ~n9465 ;
  assign y4883 = ~1'b0 ;
  assign y4884 = ~n9467 ;
  assign y4885 = ~n9468 ;
  assign y4886 = ~1'b0 ;
  assign y4887 = ~n9473 ;
  assign y4888 = ~n3968 ;
  assign y4889 = ~1'b0 ;
  assign y4890 = ~n9476 ;
  assign y4891 = n4780 ;
  assign y4892 = n9478 ;
  assign y4893 = ~1'b0 ;
  assign y4894 = ~1'b0 ;
  assign y4895 = ~1'b0 ;
  assign y4896 = ~n9481 ;
  assign y4897 = ~n9483 ;
  assign y4898 = ~n9484 ;
  assign y4899 = ~n9485 ;
  assign y4900 = ~n9486 ;
  assign y4901 = ~n9489 ;
  assign y4902 = ~n9493 ;
  assign y4903 = ~n9495 ;
  assign y4904 = ~1'b0 ;
  assign y4905 = ~n9500 ;
  assign y4906 = ~1'b0 ;
  assign y4907 = n5438 ;
  assign y4908 = n9502 ;
  assign y4909 = ~n9503 ;
  assign y4910 = ~n9507 ;
  assign y4911 = ~n9513 ;
  assign y4912 = ~1'b0 ;
  assign y4913 = ~n9515 ;
  assign y4914 = ~n9521 ;
  assign y4915 = ~n9523 ;
  assign y4916 = ~1'b0 ;
  assign y4917 = ~1'b0 ;
  assign y4918 = n9530 ;
  assign y4919 = ~1'b0 ;
  assign y4920 = ~n9534 ;
  assign y4921 = ~n9538 ;
  assign y4922 = ~n9539 ;
  assign y4923 = n9543 ;
  assign y4924 = ~1'b0 ;
  assign y4925 = ~n9544 ;
  assign y4926 = n9550 ;
  assign y4927 = ~1'b0 ;
  assign y4928 = ~n9552 ;
  assign y4929 = n9553 ;
  assign y4930 = ~1'b0 ;
  assign y4931 = ~1'b0 ;
  assign y4932 = ~1'b0 ;
  assign y4933 = n9559 ;
  assign y4934 = n9560 ;
  assign y4935 = ~1'b0 ;
  assign y4936 = ~1'b0 ;
  assign y4937 = ~n9570 ;
  assign y4938 = ~1'b0 ;
  assign y4939 = ~n9572 ;
  assign y4940 = ~n9574 ;
  assign y4941 = ~n9584 ;
  assign y4942 = ~n9585 ;
  assign y4943 = n9589 ;
  assign y4944 = n9590 ;
  assign y4945 = ~n9593 ;
  assign y4946 = n9597 ;
  assign y4947 = n9598 ;
  assign y4948 = ~n9599 ;
  assign y4949 = n9601 ;
  assign y4950 = ~n9602 ;
  assign y4951 = n9604 ;
  assign y4952 = n9608 ;
  assign y4953 = ~1'b0 ;
  assign y4954 = ~n9609 ;
  assign y4955 = n9611 ;
  assign y4956 = ~n9615 ;
  assign y4957 = ~1'b0 ;
  assign y4958 = ~n9616 ;
  assign y4959 = ~n9625 ;
  assign y4960 = ~1'b0 ;
  assign y4961 = 1'b0 ;
  assign y4962 = 1'b0 ;
  assign y4963 = ~1'b0 ;
  assign y4964 = ~n9629 ;
  assign y4965 = 1'b0 ;
  assign y4966 = ~n9632 ;
  assign y4967 = ~n9636 ;
  assign y4968 = n9639 ;
  assign y4969 = ~1'b0 ;
  assign y4970 = n9641 ;
  assign y4971 = ~1'b0 ;
  assign y4972 = ~1'b0 ;
  assign y4973 = ~1'b0 ;
  assign y4974 = ~1'b0 ;
  assign y4975 = n9645 ;
  assign y4976 = n9648 ;
  assign y4977 = 1'b0 ;
  assign y4978 = n7126 ;
  assign y4979 = n9655 ;
  assign y4980 = ~1'b0 ;
  assign y4981 = n9660 ;
  assign y4982 = ~1'b0 ;
  assign y4983 = n9662 ;
  assign y4984 = n9663 ;
  assign y4985 = n9664 ;
  assign y4986 = ~1'b0 ;
  assign y4987 = n9665 ;
  assign y4988 = ~1'b0 ;
  assign y4989 = ~n9667 ;
  assign y4990 = ~n9668 ;
  assign y4991 = n9672 ;
  assign y4992 = n9674 ;
  assign y4993 = n9676 ;
  assign y4994 = ~n9678 ;
  assign y4995 = ~n967 ;
  assign y4996 = ~n9684 ;
  assign y4997 = ~n9687 ;
  assign y4998 = ~n9693 ;
  assign y4999 = ~n9696 ;
  assign y5000 = ~n9697 ;
  assign y5001 = ~n7335 ;
  assign y5002 = ~1'b0 ;
  assign y5003 = 1'b0 ;
  assign y5004 = ~n9698 ;
  assign y5005 = 1'b0 ;
  assign y5006 = n9699 ;
  assign y5007 = ~n9704 ;
  assign y5008 = 1'b0 ;
  assign y5009 = n9706 ;
  assign y5010 = ~1'b0 ;
  assign y5011 = ~1'b0 ;
  assign y5012 = ~n9709 ;
  assign y5013 = n9710 ;
  assign y5014 = n9714 ;
  assign y5015 = ~n9719 ;
  assign y5016 = ~1'b0 ;
  assign y5017 = ~1'b0 ;
  assign y5018 = n9726 ;
  assign y5019 = ~1'b0 ;
  assign y5020 = ~1'b0 ;
  assign y5021 = n9729 ;
  assign y5022 = n9731 ;
  assign y5023 = ~n9732 ;
  assign y5024 = n9733 ;
  assign y5025 = ~n9743 ;
  assign y5026 = ~1'b0 ;
  assign y5027 = ~1'b0 ;
  assign y5028 = ~1'b0 ;
  assign y5029 = ~n7405 ;
  assign y5030 = ~n9749 ;
  assign y5031 = ~n9758 ;
  assign y5032 = n9761 ;
  assign y5033 = ~n9765 ;
  assign y5034 = ~n9769 ;
  assign y5035 = ~n9776 ;
  assign y5036 = ~1'b0 ;
  assign y5037 = ~1'b0 ;
  assign y5038 = n3867 ;
  assign y5039 = ~1'b0 ;
  assign y5040 = n9777 ;
  assign y5041 = ~n9783 ;
  assign y5042 = 1'b0 ;
  assign y5043 = n9784 ;
  assign y5044 = ~1'b0 ;
  assign y5045 = n9787 ;
  assign y5046 = n9788 ;
  assign y5047 = ~n9789 ;
  assign y5048 = n2658 ;
  assign y5049 = ~1'b0 ;
  assign y5050 = n9790 ;
  assign y5051 = n2619 ;
  assign y5052 = ~1'b0 ;
  assign y5053 = ~n9794 ;
  assign y5054 = ~1'b0 ;
  assign y5055 = ~1'b0 ;
  assign y5056 = n9799 ;
  assign y5057 = ~n9816 ;
  assign y5058 = ~1'b0 ;
  assign y5059 = ~n9819 ;
  assign y5060 = ~1'b0 ;
  assign y5061 = n9827 ;
  assign y5062 = n9832 ;
  assign y5063 = ~n9833 ;
  assign y5064 = ~n9836 ;
  assign y5065 = ~n9837 ;
  assign y5066 = ~n9850 ;
  assign y5067 = n9855 ;
  assign y5068 = ~n9863 ;
  assign y5069 = ~n9867 ;
  assign y5070 = ~n9874 ;
  assign y5071 = ~1'b0 ;
  assign y5072 = ~n9878 ;
  assign y5073 = n9880 ;
  assign y5074 = ~n3992 ;
  assign y5075 = ~1'b0 ;
  assign y5076 = ~1'b0 ;
  assign y5077 = ~n9883 ;
  assign y5078 = ~n9884 ;
  assign y5079 = ~1'b0 ;
  assign y5080 = ~1'b0 ;
  assign y5081 = ~n9886 ;
  assign y5082 = ~n9891 ;
  assign y5083 = n9893 ;
  assign y5084 = n9898 ;
  assign y5085 = ~1'b0 ;
  assign y5086 = ~1'b0 ;
  assign y5087 = ~1'b0 ;
  assign y5088 = ~n9899 ;
  assign y5089 = ~1'b0 ;
  assign y5090 = n9901 ;
  assign y5091 = ~1'b0 ;
  assign y5092 = n9907 ;
  assign y5093 = ~n9908 ;
  assign y5094 = ~n9910 ;
  assign y5095 = ~1'b0 ;
  assign y5096 = ~n9922 ;
  assign y5097 = n9923 ;
  assign y5098 = ~n9925 ;
  assign y5099 = n9927 ;
  assign y5100 = ~n9929 ;
  assign y5101 = n9933 ;
  assign y5102 = ~1'b0 ;
  assign y5103 = ~n9934 ;
  assign y5104 = ~n9940 ;
  assign y5105 = ~n9943 ;
  assign y5106 = n9945 ;
  assign y5107 = ~n9948 ;
  assign y5108 = n9953 ;
  assign y5109 = ~1'b0 ;
  assign y5110 = ~1'b0 ;
  assign y5111 = n9962 ;
  assign y5112 = ~n9965 ;
  assign y5113 = ~n9967 ;
  assign y5114 = n9969 ;
  assign y5115 = n9973 ;
  assign y5116 = ~1'b0 ;
  assign y5117 = 1'b0 ;
  assign y5118 = 1'b0 ;
  assign y5119 = ~n7257 ;
  assign y5120 = ~n9974 ;
  assign y5121 = ~n1778 ;
  assign y5122 = n9975 ;
  assign y5123 = n9977 ;
  assign y5124 = n9979 ;
  assign y5125 = ~1'b0 ;
  assign y5126 = n9983 ;
  assign y5127 = ~n9987 ;
  assign y5128 = ~1'b0 ;
  assign y5129 = ~n9990 ;
  assign y5130 = n9994 ;
  assign y5131 = ~n9996 ;
  assign y5132 = ~n10001 ;
  assign y5133 = n10002 ;
  assign y5134 = ~1'b0 ;
  assign y5135 = ~n10004 ;
  assign y5136 = n10005 ;
  assign y5137 = ~n10007 ;
  assign y5138 = ~n10015 ;
  assign y5139 = n10016 ;
  assign y5140 = ~n10018 ;
  assign y5141 = ~n10019 ;
  assign y5142 = n10022 ;
  assign y5143 = ~1'b0 ;
  assign y5144 = n10029 ;
  assign y5145 = n10031 ;
  assign y5146 = n10034 ;
  assign y5147 = ~n10037 ;
  assign y5148 = n7413 ;
  assign y5149 = n10040 ;
  assign y5150 = n10041 ;
  assign y5151 = ~n10042 ;
  assign y5152 = n10044 ;
  assign y5153 = ~1'b0 ;
  assign y5154 = n10045 ;
  assign y5155 = ~1'b0 ;
  assign y5156 = ~1'b0 ;
  assign y5157 = ~n10051 ;
  assign y5158 = n10054 ;
  assign y5159 = ~n10055 ;
  assign y5160 = ~1'b0 ;
  assign y5161 = ~1'b0 ;
  assign y5162 = ~1'b0 ;
  assign y5163 = ~n10056 ;
  assign y5164 = ~n10057 ;
  assign y5165 = ~n10061 ;
  assign y5166 = n10066 ;
  assign y5167 = n10070 ;
  assign y5168 = ~n10071 ;
  assign y5169 = ~n10073 ;
  assign y5170 = ~1'b0 ;
  assign y5171 = ~1'b0 ;
  assign y5172 = ~1'b0 ;
  assign y5173 = 1'b0 ;
  assign y5174 = ~1'b0 ;
  assign y5175 = ~1'b0 ;
  assign y5176 = ~n10075 ;
  assign y5177 = ~n10076 ;
  assign y5178 = n10078 ;
  assign y5179 = ~1'b0 ;
  assign y5180 = n10081 ;
  assign y5181 = n10084 ;
  assign y5182 = ~1'b0 ;
  assign y5183 = ~n10086 ;
  assign y5184 = ~1'b0 ;
  assign y5185 = ~n10087 ;
  assign y5186 = ~1'b0 ;
  assign y5187 = ~1'b0 ;
  assign y5188 = n4395 ;
  assign y5189 = n10089 ;
  assign y5190 = ~n10092 ;
  assign y5191 = ~n10093 ;
  assign y5192 = ~n10105 ;
  assign y5193 = n10106 ;
  assign y5194 = ~n10108 ;
  assign y5195 = n10111 ;
  assign y5196 = n10114 ;
  assign y5197 = ~1'b0 ;
  assign y5198 = n4589 ;
  assign y5199 = n10118 ;
  assign y5200 = ~n10119 ;
  assign y5201 = ~1'b0 ;
  assign y5202 = n10120 ;
  assign y5203 = n10123 ;
  assign y5204 = ~1'b0 ;
  assign y5205 = ~n1055 ;
  assign y5206 = ~1'b0 ;
  assign y5207 = ~1'b0 ;
  assign y5208 = n4461 ;
  assign y5209 = ~1'b0 ;
  assign y5210 = n10126 ;
  assign y5211 = ~1'b0 ;
  assign y5212 = ~n10129 ;
  assign y5213 = n10133 ;
  assign y5214 = ~1'b0 ;
  assign y5215 = n10134 ;
  assign y5216 = ~n10135 ;
  assign y5217 = ~1'b0 ;
  assign y5218 = n10136 ;
  assign y5219 = ~n10137 ;
  assign y5220 = n10140 ;
  assign y5221 = ~n10142 ;
  assign y5222 = ~1'b0 ;
  assign y5223 = ~n10143 ;
  assign y5224 = ~n10145 ;
  assign y5225 = n10146 ;
  assign y5226 = ~n10147 ;
  assign y5227 = n10150 ;
  assign y5228 = ~1'b0 ;
  assign y5229 = n10152 ;
  assign y5230 = ~n10153 ;
  assign y5231 = ~1'b0 ;
  assign y5232 = ~1'b0 ;
  assign y5233 = ~1'b0 ;
  assign y5234 = n10157 ;
  assign y5235 = n10160 ;
  assign y5236 = ~1'b0 ;
  assign y5237 = n10162 ;
  assign y5238 = n10166 ;
  assign y5239 = ~1'b0 ;
  assign y5240 = ~n10167 ;
  assign y5241 = ~1'b0 ;
  assign y5242 = ~1'b0 ;
  assign y5243 = ~1'b0 ;
  assign y5244 = ~n10170 ;
  assign y5245 = ~n10171 ;
  assign y5246 = ~1'b0 ;
  assign y5247 = n10178 ;
  assign y5248 = n10180 ;
  assign y5249 = ~n10182 ;
  assign y5250 = ~n10187 ;
  assign y5251 = ~n10188 ;
  assign y5252 = ~n10189 ;
  assign y5253 = ~1'b0 ;
  assign y5254 = n10191 ;
  assign y5255 = ~n10193 ;
  assign y5256 = ~n10195 ;
  assign y5257 = n10196 ;
  assign y5258 = ~1'b0 ;
  assign y5259 = n10197 ;
  assign y5260 = n10198 ;
  assign y5261 = ~n10203 ;
  assign y5262 = n10205 ;
  assign y5263 = n10207 ;
  assign y5264 = ~1'b0 ;
  assign y5265 = ~1'b0 ;
  assign y5266 = ~n10208 ;
  assign y5267 = n10210 ;
  assign y5268 = n10212 ;
  assign y5269 = n7265 ;
  assign y5270 = ~1'b0 ;
  assign y5271 = ~n10213 ;
  assign y5272 = ~n10221 ;
  assign y5273 = ~n8725 ;
  assign y5274 = ~1'b0 ;
  assign y5275 = n10223 ;
  assign y5276 = n10225 ;
  assign y5277 = ~n10228 ;
  assign y5278 = ~1'b0 ;
  assign y5279 = ~n4039 ;
  assign y5280 = n10230 ;
  assign y5281 = ~1'b0 ;
  assign y5282 = ~n10232 ;
  assign y5283 = ~n10234 ;
  assign y5284 = ~n10235 ;
  assign y5285 = n10238 ;
  assign y5286 = ~n10239 ;
  assign y5287 = n10241 ;
  assign y5288 = ~1'b0 ;
  assign y5289 = ~n10242 ;
  assign y5290 = ~1'b0 ;
  assign y5291 = ~1'b0 ;
  assign y5292 = ~n10244 ;
  assign y5293 = n7520 ;
  assign y5294 = n10245 ;
  assign y5295 = ~n4993 ;
  assign y5296 = ~1'b0 ;
  assign y5297 = ~1'b0 ;
  assign y5298 = ~1'b0 ;
  assign y5299 = ~n10248 ;
  assign y5300 = ~n10249 ;
  assign y5301 = n10257 ;
  assign y5302 = ~n10259 ;
  assign y5303 = 1'b0 ;
  assign y5304 = ~n10263 ;
  assign y5305 = n10265 ;
  assign y5306 = ~n10267 ;
  assign y5307 = ~n10268 ;
  assign y5308 = ~n10271 ;
  assign y5309 = ~n10274 ;
  assign y5310 = ~1'b0 ;
  assign y5311 = ~1'b0 ;
  assign y5312 = ~n10275 ;
  assign y5313 = n10277 ;
  assign y5314 = ~1'b0 ;
  assign y5315 = ~n10280 ;
  assign y5316 = n10281 ;
  assign y5317 = ~n10283 ;
  assign y5318 = ~1'b0 ;
  assign y5319 = ~1'b0 ;
  assign y5320 = ~n10284 ;
  assign y5321 = ~n10286 ;
  assign y5322 = ~1'b0 ;
  assign y5323 = n10288 ;
  assign y5324 = ~n10289 ;
  assign y5325 = ~n10294 ;
  assign y5326 = ~n10295 ;
  assign y5327 = n10297 ;
  assign y5328 = ~1'b0 ;
  assign y5329 = n10302 ;
  assign y5330 = ~1'b0 ;
  assign y5331 = n10303 ;
  assign y5332 = ~1'b0 ;
  assign y5333 = ~n10306 ;
  assign y5334 = ~1'b0 ;
  assign y5335 = ~n10307 ;
  assign y5336 = ~n10314 ;
  assign y5337 = ~n10315 ;
  assign y5338 = ~n657 ;
  assign y5339 = ~1'b0 ;
  assign y5340 = n10317 ;
  assign y5341 = ~n10321 ;
  assign y5342 = n10323 ;
  assign y5343 = n10327 ;
  assign y5344 = ~1'b0 ;
  assign y5345 = ~n10329 ;
  assign y5346 = n10335 ;
  assign y5347 = ~1'b0 ;
  assign y5348 = ~n10340 ;
  assign y5349 = n10343 ;
  assign y5350 = ~1'b0 ;
  assign y5351 = n10345 ;
  assign y5352 = ~n10347 ;
  assign y5353 = n3259 ;
  assign y5354 = ~n10354 ;
  assign y5355 = ~1'b0 ;
  assign y5356 = n10361 ;
  assign y5357 = ~n10363 ;
  assign y5358 = n10365 ;
  assign y5359 = ~1'b0 ;
  assign y5360 = 1'b0 ;
  assign y5361 = ~1'b0 ;
  assign y5362 = ~n10366 ;
  assign y5363 = n10367 ;
  assign y5364 = ~n4707 ;
  assign y5365 = ~n10368 ;
  assign y5366 = ~1'b0 ;
  assign y5367 = ~n10369 ;
  assign y5368 = ~n10376 ;
  assign y5369 = n10381 ;
  assign y5370 = ~n10387 ;
  assign y5371 = ~n7316 ;
  assign y5372 = ~1'b0 ;
  assign y5373 = ~n10389 ;
  assign y5374 = n10391 ;
  assign y5375 = ~1'b0 ;
  assign y5376 = n10393 ;
  assign y5377 = ~1'b0 ;
  assign y5378 = ~n10399 ;
  assign y5379 = n10405 ;
  assign y5380 = ~n10406 ;
  assign y5381 = ~n10407 ;
  assign y5382 = ~n10411 ;
  assign y5383 = ~n10412 ;
  assign y5384 = ~1'b0 ;
  assign y5385 = ~n10415 ;
  assign y5386 = ~1'b0 ;
  assign y5387 = n10420 ;
  assign y5388 = ~n4317 ;
  assign y5389 = n10423 ;
  assign y5390 = n10425 ;
  assign y5391 = n10426 ;
  assign y5392 = n10431 ;
  assign y5393 = ~1'b0 ;
  assign y5394 = ~1'b0 ;
  assign y5395 = n10432 ;
  assign y5396 = n10433 ;
  assign y5397 = ~1'b0 ;
  assign y5398 = ~n6749 ;
  assign y5399 = ~n10436 ;
  assign y5400 = n10437 ;
  assign y5401 = ~n10439 ;
  assign y5402 = ~n6215 ;
  assign y5403 = ~1'b0 ;
  assign y5404 = ~n10443 ;
  assign y5405 = ~n10445 ;
  assign y5406 = ~1'b0 ;
  assign y5407 = ~n4531 ;
  assign y5408 = ~n10447 ;
  assign y5409 = n10451 ;
  assign y5410 = n10457 ;
  assign y5411 = n10462 ;
  assign y5412 = ~1'b0 ;
  assign y5413 = ~n10468 ;
  assign y5414 = ~1'b0 ;
  assign y5415 = n10470 ;
  assign y5416 = ~1'b0 ;
  assign y5417 = ~1'b0 ;
  assign y5418 = ~1'b0 ;
  assign y5419 = n10480 ;
  assign y5420 = n10483 ;
  assign y5421 = n10484 ;
  assign y5422 = 1'b0 ;
  assign y5423 = n10488 ;
  assign y5424 = n10489 ;
  assign y5425 = ~n10491 ;
  assign y5426 = n10493 ;
  assign y5427 = n10495 ;
  assign y5428 = ~n10499 ;
  assign y5429 = ~1'b0 ;
  assign y5430 = ~1'b0 ;
  assign y5431 = n10501 ;
  assign y5432 = ~n10505 ;
  assign y5433 = ~1'b0 ;
  assign y5434 = ~1'b0 ;
  assign y5435 = ~1'b0 ;
  assign y5436 = ~n10514 ;
  assign y5437 = ~n10516 ;
  assign y5438 = ~1'b0 ;
  assign y5439 = n10521 ;
  assign y5440 = n10522 ;
  assign y5441 = n10524 ;
  assign y5442 = n8482 ;
  assign y5443 = ~1'b0 ;
  assign y5444 = ~1'b0 ;
  assign y5445 = ~1'b0 ;
  assign y5446 = n9724 ;
  assign y5447 = ~n10527 ;
  assign y5448 = ~1'b0 ;
  assign y5449 = ~n10528 ;
  assign y5450 = ~n10529 ;
  assign y5451 = n10530 ;
  assign y5452 = ~n10533 ;
  assign y5453 = ~1'b0 ;
  assign y5454 = n10534 ;
  assign y5455 = ~n10536 ;
  assign y5456 = n10538 ;
  assign y5457 = ~1'b0 ;
  assign y5458 = 1'b0 ;
  assign y5459 = ~n10539 ;
  assign y5460 = ~n10543 ;
  assign y5461 = ~1'b0 ;
  assign y5462 = ~1'b0 ;
  assign y5463 = ~n10545 ;
  assign y5464 = n10548 ;
  assign y5465 = ~1'b0 ;
  assign y5466 = ~1'b0 ;
  assign y5467 = ~n10559 ;
  assign y5468 = n10560 ;
  assign y5469 = n8365 ;
  assign y5470 = ~n4142 ;
  assign y5471 = ~1'b0 ;
  assign y5472 = ~n10564 ;
  assign y5473 = ~1'b0 ;
  assign y5474 = n10565 ;
  assign y5475 = ~n10570 ;
  assign y5476 = n10582 ;
  assign y5477 = n10586 ;
  assign y5478 = n10587 ;
  assign y5479 = ~1'b0 ;
  assign y5480 = n10593 ;
  assign y5481 = n5755 ;
  assign y5482 = ~1'b0 ;
  assign y5483 = ~n10596 ;
  assign y5484 = n10598 ;
  assign y5485 = ~1'b0 ;
  assign y5486 = ~n10600 ;
  assign y5487 = ~1'b0 ;
  assign y5488 = n1479 ;
  assign y5489 = n10601 ;
  assign y5490 = ~n10606 ;
  assign y5491 = n10609 ;
  assign y5492 = ~1'b0 ;
  assign y5493 = ~n10612 ;
  assign y5494 = ~1'b0 ;
  assign y5495 = n10618 ;
  assign y5496 = n10620 ;
  assign y5497 = n10622 ;
  assign y5498 = ~n10632 ;
  assign y5499 = ~1'b0 ;
  assign y5500 = ~n10638 ;
  assign y5501 = ~1'b0 ;
  assign y5502 = ~n10649 ;
  assign y5503 = ~n10652 ;
  assign y5504 = ~n10653 ;
  assign y5505 = ~n10656 ;
  assign y5506 = ~n10657 ;
  assign y5507 = ~1'b0 ;
  assign y5508 = n10658 ;
  assign y5509 = 1'b0 ;
  assign y5510 = ~n10662 ;
  assign y5511 = ~n10667 ;
  assign y5512 = ~n10672 ;
  assign y5513 = ~1'b0 ;
  assign y5514 = ~n10673 ;
  assign y5515 = ~1'b0 ;
  assign y5516 = ~1'b0 ;
  assign y5517 = ~n10674 ;
  assign y5518 = ~n10678 ;
  assign y5519 = n10682 ;
  assign y5520 = ~1'b0 ;
  assign y5521 = ~1'b0 ;
  assign y5522 = ~n10684 ;
  assign y5523 = ~1'b0 ;
  assign y5524 = n10688 ;
  assign y5525 = n10692 ;
  assign y5526 = ~n10701 ;
  assign y5527 = n10703 ;
  assign y5528 = ~n10705 ;
  assign y5529 = ~n10711 ;
  assign y5530 = n10713 ;
  assign y5531 = ~1'b0 ;
  assign y5532 = ~1'b0 ;
  assign y5533 = ~n10716 ;
  assign y5534 = n10719 ;
  assign y5535 = n10720 ;
  assign y5536 = n10728 ;
  assign y5537 = ~1'b0 ;
  assign y5538 = ~n10731 ;
  assign y5539 = ~n10733 ;
  assign y5540 = 1'b0 ;
  assign y5541 = n2946 ;
  assign y5542 = n10735 ;
  assign y5543 = n10737 ;
  assign y5544 = n10739 ;
  assign y5545 = ~1'b0 ;
  assign y5546 = ~1'b0 ;
  assign y5547 = ~1'b0 ;
  assign y5548 = ~n10743 ;
  assign y5549 = ~n10745 ;
  assign y5550 = ~1'b0 ;
  assign y5551 = ~1'b0 ;
  assign y5552 = ~n10748 ;
  assign y5553 = ~1'b0 ;
  assign y5554 = n10753 ;
  assign y5555 = n10756 ;
  assign y5556 = n7116 ;
  assign y5557 = ~n10759 ;
  assign y5558 = n10761 ;
  assign y5559 = ~1'b0 ;
  assign y5560 = ~n10762 ;
  assign y5561 = n10764 ;
  assign y5562 = n10767 ;
  assign y5563 = 1'b0 ;
  assign y5564 = n10770 ;
  assign y5565 = n10774 ;
  assign y5566 = ~n10776 ;
  assign y5567 = ~1'b0 ;
  assign y5568 = n1325 ;
  assign y5569 = ~1'b0 ;
  assign y5570 = ~n4732 ;
  assign y5571 = ~n10780 ;
  assign y5572 = n10782 ;
  assign y5573 = ~1'b0 ;
  assign y5574 = ~n10784 ;
  assign y5575 = n10785 ;
  assign y5576 = ~n10788 ;
  assign y5577 = ~1'b0 ;
  assign y5578 = n10792 ;
  assign y5579 = ~n10795 ;
  assign y5580 = 1'b0 ;
  assign y5581 = ~n10796 ;
  assign y5582 = ~n10801 ;
  assign y5583 = ~1'b0 ;
  assign y5584 = n8163 ;
  assign y5585 = ~1'b0 ;
  assign y5586 = n10803 ;
  assign y5587 = ~n10807 ;
  assign y5588 = n10809 ;
  assign y5589 = n10812 ;
  assign y5590 = ~1'b0 ;
  assign y5591 = ~n10814 ;
  assign y5592 = ~1'b0 ;
  assign y5593 = n10815 ;
  assign y5594 = n10816 ;
  assign y5595 = n10819 ;
  assign y5596 = ~n10825 ;
  assign y5597 = ~1'b0 ;
  assign y5598 = ~n10829 ;
  assign y5599 = ~n10832 ;
  assign y5600 = ~n10834 ;
  assign y5601 = ~n10839 ;
  assign y5602 = ~n10847 ;
  assign y5603 = ~n10848 ;
  assign y5604 = ~n10850 ;
  assign y5605 = n10851 ;
  assign y5606 = ~n10856 ;
  assign y5607 = ~1'b0 ;
  assign y5608 = ~n6124 ;
  assign y5609 = ~1'b0 ;
  assign y5610 = ~n10861 ;
  assign y5611 = ~1'b0 ;
  assign y5612 = ~1'b0 ;
  assign y5613 = ~1'b0 ;
  assign y5614 = n10862 ;
  assign y5615 = ~1'b0 ;
  assign y5616 = ~1'b0 ;
  assign y5617 = ~1'b0 ;
  assign y5618 = n10863 ;
  assign y5619 = ~1'b0 ;
  assign y5620 = ~n10868 ;
  assign y5621 = ~1'b0 ;
  assign y5622 = ~1'b0 ;
  assign y5623 = ~1'b0 ;
  assign y5624 = n10870 ;
  assign y5625 = ~n10881 ;
  assign y5626 = n10882 ;
  assign y5627 = ~1'b0 ;
  assign y5628 = n10883 ;
  assign y5629 = ~n10885 ;
  assign y5630 = n10886 ;
  assign y5631 = ~n10891 ;
  assign y5632 = n2079 ;
  assign y5633 = ~1'b0 ;
  assign y5634 = n10892 ;
  assign y5635 = ~1'b0 ;
  assign y5636 = ~1'b0 ;
  assign y5637 = ~1'b0 ;
  assign y5638 = n10894 ;
  assign y5639 = ~n10900 ;
  assign y5640 = ~1'b0 ;
  assign y5641 = ~n10901 ;
  assign y5642 = ~n10902 ;
  assign y5643 = n10903 ;
  assign y5644 = n10905 ;
  assign y5645 = n10907 ;
  assign y5646 = n10909 ;
  assign y5647 = ~n10910 ;
  assign y5648 = ~n10914 ;
  assign y5649 = n10931 ;
  assign y5650 = ~n10937 ;
  assign y5651 = ~n10946 ;
  assign y5652 = ~1'b0 ;
  assign y5653 = ~n10950 ;
  assign y5654 = ~1'b0 ;
  assign y5655 = n10951 ;
  assign y5656 = ~1'b0 ;
  assign y5657 = ~1'b0 ;
  assign y5658 = n10957 ;
  assign y5659 = n10958 ;
  assign y5660 = ~1'b0 ;
  assign y5661 = n10959 ;
  assign y5662 = ~n10961 ;
  assign y5663 = ~n10962 ;
  assign y5664 = ~n10964 ;
  assign y5665 = n10967 ;
  assign y5666 = ~1'b0 ;
  assign y5667 = ~n10968 ;
  assign y5668 = ~1'b0 ;
  assign y5669 = ~n10975 ;
  assign y5670 = ~1'b0 ;
  assign y5671 = ~n10976 ;
  assign y5672 = ~1'b0 ;
  assign y5673 = ~1'b0 ;
  assign y5674 = ~1'b0 ;
  assign y5675 = ~n10980 ;
  assign y5676 = n10994 ;
  assign y5677 = n10997 ;
  assign y5678 = ~1'b0 ;
  assign y5679 = ~1'b0 ;
  assign y5680 = ~1'b0 ;
  assign y5681 = ~1'b0 ;
  assign y5682 = n10998 ;
  assign y5683 = n11000 ;
  assign y5684 = ~1'b0 ;
  assign y5685 = n11001 ;
  assign y5686 = n11006 ;
  assign y5687 = ~1'b0 ;
  assign y5688 = ~n11008 ;
  assign y5689 = ~1'b0 ;
  assign y5690 = ~n11011 ;
  assign y5691 = n11014 ;
  assign y5692 = 1'b0 ;
  assign y5693 = 1'b0 ;
  assign y5694 = ~1'b0 ;
  assign y5695 = ~n11020 ;
  assign y5696 = ~1'b0 ;
  assign y5697 = ~n11021 ;
  assign y5698 = ~1'b0 ;
  assign y5699 = n11023 ;
  assign y5700 = ~n11027 ;
  assign y5701 = n11033 ;
  assign y5702 = ~n11034 ;
  assign y5703 = n1047 ;
  assign y5704 = ~n11035 ;
  assign y5705 = ~n11037 ;
  assign y5706 = n11038 ;
  assign y5707 = n11046 ;
  assign y5708 = n11048 ;
  assign y5709 = ~n11050 ;
  assign y5710 = ~1'b0 ;
  assign y5711 = ~n11054 ;
  assign y5712 = ~1'b0 ;
  assign y5713 = ~n11056 ;
  assign y5714 = n11062 ;
  assign y5715 = n11063 ;
  assign y5716 = ~1'b0 ;
  assign y5717 = n11064 ;
  assign y5718 = ~1'b0 ;
  assign y5719 = ~1'b0 ;
  assign y5720 = n11065 ;
  assign y5721 = n11066 ;
  assign y5722 = ~n11070 ;
  assign y5723 = ~n11072 ;
  assign y5724 = n11081 ;
  assign y5725 = ~n11083 ;
  assign y5726 = ~n11085 ;
  assign y5727 = n11087 ;
  assign y5728 = 1'b0 ;
  assign y5729 = ~n2093 ;
  assign y5730 = n11095 ;
  assign y5731 = ~n11098 ;
  assign y5732 = ~1'b0 ;
  assign y5733 = ~1'b0 ;
  assign y5734 = n11100 ;
  assign y5735 = ~n11102 ;
  assign y5736 = 1'b0 ;
  assign y5737 = ~1'b0 ;
  assign y5738 = ~n11105 ;
  assign y5739 = ~n11113 ;
  assign y5740 = n11115 ;
  assign y5741 = n11117 ;
  assign y5742 = ~n11118 ;
  assign y5743 = ~n11119 ;
  assign y5744 = ~n11122 ;
  assign y5745 = n11127 ;
  assign y5746 = ~n11129 ;
  assign y5747 = ~1'b0 ;
  assign y5748 = ~1'b0 ;
  assign y5749 = ~n11131 ;
  assign y5750 = ~n11137 ;
  assign y5751 = n11138 ;
  assign y5752 = ~1'b0 ;
  assign y5753 = 1'b0 ;
  assign y5754 = ~n11140 ;
  assign y5755 = ~n10093 ;
  assign y5756 = ~n11142 ;
  assign y5757 = n11144 ;
  assign y5758 = ~n11147 ;
  assign y5759 = ~1'b0 ;
  assign y5760 = n11148 ;
  assign y5761 = n11152 ;
  assign y5762 = ~1'b0 ;
  assign y5763 = ~1'b0 ;
  assign y5764 = ~n11154 ;
  assign y5765 = ~1'b0 ;
  assign y5766 = 1'b0 ;
  assign y5767 = ~1'b0 ;
  assign y5768 = ~1'b0 ;
  assign y5769 = ~n11155 ;
  assign y5770 = n11162 ;
  assign y5771 = ~n11165 ;
  assign y5772 = n11166 ;
  assign y5773 = n11174 ;
  assign y5774 = n5549 ;
  assign y5775 = n11176 ;
  assign y5776 = ~1'b0 ;
  assign y5777 = n11177 ;
  assign y5778 = n11180 ;
  assign y5779 = n11183 ;
  assign y5780 = ~1'b0 ;
  assign y5781 = n11184 ;
  assign y5782 = n11187 ;
  assign y5783 = ~1'b0 ;
  assign y5784 = ~1'b0 ;
  assign y5785 = ~1'b0 ;
  assign y5786 = n11192 ;
  assign y5787 = n11194 ;
  assign y5788 = ~n11201 ;
  assign y5789 = ~n11202 ;
  assign y5790 = ~n11204 ;
  assign y5791 = ~n11211 ;
  assign y5792 = ~n11217 ;
  assign y5793 = n11222 ;
  assign y5794 = ~1'b0 ;
  assign y5795 = ~1'b0 ;
  assign y5796 = ~1'b0 ;
  assign y5797 = ~n11223 ;
  assign y5798 = ~1'b0 ;
  assign y5799 = ~n4357 ;
  assign y5800 = ~n11228 ;
  assign y5801 = ~n11230 ;
  assign y5802 = ~n11232 ;
  assign y5803 = ~n11238 ;
  assign y5804 = ~1'b0 ;
  assign y5805 = n11243 ;
  assign y5806 = 1'b0 ;
  assign y5807 = ~n7529 ;
  assign y5808 = ~n11244 ;
  assign y5809 = n11246 ;
  assign y5810 = ~1'b0 ;
  assign y5811 = n11249 ;
  assign y5812 = 1'b0 ;
  assign y5813 = ~1'b0 ;
  assign y5814 = ~1'b0 ;
  assign y5815 = ~n11253 ;
  assign y5816 = ~n11255 ;
  assign y5817 = 1'b0 ;
  assign y5818 = ~1'b0 ;
  assign y5819 = n11256 ;
  assign y5820 = ~n11257 ;
  assign y5821 = n11258 ;
  assign y5822 = ~1'b0 ;
  assign y5823 = ~1'b0 ;
  assign y5824 = ~1'b0 ;
  assign y5825 = ~n11260 ;
  assign y5826 = ~n4569 ;
  assign y5827 = ~n11266 ;
  assign y5828 = ~n11270 ;
  assign y5829 = ~n11273 ;
  assign y5830 = ~n11274 ;
  assign y5831 = ~1'b0 ;
  assign y5832 = ~n11281 ;
  assign y5833 = ~n11285 ;
  assign y5834 = n765 ;
  assign y5835 = n11287 ;
  assign y5836 = n11290 ;
  assign y5837 = n11294 ;
  assign y5838 = ~n11295 ;
  assign y5839 = ~1'b0 ;
  assign y5840 = n11297 ;
  assign y5841 = n11299 ;
  assign y5842 = n11306 ;
  assign y5843 = ~n11308 ;
  assign y5844 = ~1'b0 ;
  assign y5845 = ~1'b0 ;
  assign y5846 = ~1'b0 ;
  assign y5847 = n11313 ;
  assign y5848 = 1'b0 ;
  assign y5849 = ~n11314 ;
  assign y5850 = n11318 ;
  assign y5851 = ~1'b0 ;
  assign y5852 = n1938 ;
  assign y5853 = n11321 ;
  assign y5854 = n11322 ;
  assign y5855 = ~n11323 ;
  assign y5856 = n11325 ;
  assign y5857 = ~n11329 ;
  assign y5858 = ~1'b0 ;
  assign y5859 = n11331 ;
  assign y5860 = n11334 ;
  assign y5861 = ~n11339 ;
  assign y5862 = n11341 ;
  assign y5863 = ~1'b0 ;
  assign y5864 = n11346 ;
  assign y5865 = n11349 ;
  assign y5866 = ~1'b0 ;
  assign y5867 = ~n11353 ;
  assign y5868 = ~1'b0 ;
  assign y5869 = ~1'b0 ;
  assign y5870 = n11358 ;
  assign y5871 = n11362 ;
  assign y5872 = n11363 ;
  assign y5873 = ~n11364 ;
  assign y5874 = ~n11366 ;
  assign y5875 = n11369 ;
  assign y5876 = n11372 ;
  assign y5877 = ~1'b0 ;
  assign y5878 = ~1'b0 ;
  assign y5879 = ~1'b0 ;
  assign y5880 = ~n11375 ;
  assign y5881 = ~n11377 ;
  assign y5882 = n11384 ;
  assign y5883 = ~1'b0 ;
  assign y5884 = ~n11387 ;
  assign y5885 = ~1'b0 ;
  assign y5886 = n11388 ;
  assign y5887 = n11389 ;
  assign y5888 = ~n11390 ;
  assign y5889 = ~n11394 ;
  assign y5890 = ~1'b0 ;
  assign y5891 = ~n11396 ;
  assign y5892 = ~n11397 ;
  assign y5893 = ~n11399 ;
  assign y5894 = ~1'b0 ;
  assign y5895 = ~1'b0 ;
  assign y5896 = 1'b0 ;
  assign y5897 = n11402 ;
  assign y5898 = ~n11405 ;
  assign y5899 = ~1'b0 ;
  assign y5900 = ~1'b0 ;
  assign y5901 = n5866 ;
  assign y5902 = ~n5391 ;
  assign y5903 = ~1'b0 ;
  assign y5904 = ~n6271 ;
  assign y5905 = n11407 ;
  assign y5906 = ~n11412 ;
  assign y5907 = n11416 ;
  assign y5908 = n11417 ;
  assign y5909 = n11418 ;
  assign y5910 = ~n11421 ;
  assign y5911 = n4641 ;
  assign y5912 = n11426 ;
  assign y5913 = n11428 ;
  assign y5914 = ~n11429 ;
  assign y5915 = ~n11431 ;
  assign y5916 = ~1'b0 ;
  assign y5917 = ~1'b0 ;
  assign y5918 = ~n11434 ;
  assign y5919 = n8720 ;
  assign y5920 = n11435 ;
  assign y5921 = ~1'b0 ;
  assign y5922 = n11436 ;
  assign y5923 = ~n11438 ;
  assign y5924 = n11400 ;
  assign y5925 = ~n11439 ;
  assign y5926 = ~1'b0 ;
  assign y5927 = ~1'b0 ;
  assign y5928 = n11440 ;
  assign y5929 = ~1'b0 ;
  assign y5930 = n11445 ;
  assign y5931 = ~n11446 ;
  assign y5932 = n11447 ;
  assign y5933 = ~1'b0 ;
  assign y5934 = ~1'b0 ;
  assign y5935 = ~1'b0 ;
  assign y5936 = n11451 ;
  assign y5937 = n11452 ;
  assign y5938 = ~n11453 ;
  assign y5939 = n11454 ;
  assign y5940 = ~n11460 ;
  assign y5941 = n11461 ;
  assign y5942 = n11462 ;
  assign y5943 = n11466 ;
  assign y5944 = ~n11467 ;
  assign y5945 = ~1'b0 ;
  assign y5946 = ~1'b0 ;
  assign y5947 = ~n11468 ;
  assign y5948 = ~n11474 ;
  assign y5949 = ~n11476 ;
  assign y5950 = ~1'b0 ;
  assign y5951 = n11477 ;
  assign y5952 = n11480 ;
  assign y5953 = ~1'b0 ;
  assign y5954 = ~1'b0 ;
  assign y5955 = 1'b0 ;
  assign y5956 = n11482 ;
  assign y5957 = 1'b0 ;
  assign y5958 = ~n11483 ;
  assign y5959 = n11484 ;
  assign y5960 = ~1'b0 ;
  assign y5961 = n11485 ;
  assign y5962 = ~1'b0 ;
  assign y5963 = ~1'b0 ;
  assign y5964 = 1'b0 ;
  assign y5965 = n11486 ;
  assign y5966 = ~1'b0 ;
  assign y5967 = ~n11487 ;
  assign y5968 = ~n11489 ;
  assign y5969 = ~n11496 ;
  assign y5970 = ~1'b0 ;
  assign y5971 = n11499 ;
  assign y5972 = n1269 ;
  assign y5973 = n11502 ;
  assign y5974 = n11503 ;
  assign y5975 = ~n11504 ;
  assign y5976 = 1'b0 ;
  assign y5977 = ~1'b0 ;
  assign y5978 = n11506 ;
  assign y5979 = n11508 ;
  assign y5980 = ~n11511 ;
  assign y5981 = ~n11514 ;
  assign y5982 = n11518 ;
  assign y5983 = n11530 ;
  assign y5984 = n11532 ;
  assign y5985 = ~n10449 ;
  assign y5986 = ~1'b0 ;
  assign y5987 = ~1'b0 ;
  assign y5988 = ~n11533 ;
  assign y5989 = n11534 ;
  assign y5990 = ~n11536 ;
  assign y5991 = n11540 ;
  assign y5992 = n11541 ;
  assign y5993 = ~1'b0 ;
  assign y5994 = 1'b0 ;
  assign y5995 = ~1'b0 ;
  assign y5996 = n10616 ;
  assign y5997 = ~n11543 ;
  assign y5998 = ~1'b0 ;
  assign y5999 = ~n11549 ;
  assign y6000 = ~1'b0 ;
  assign y6001 = ~1'b0 ;
  assign y6002 = n11550 ;
  assign y6003 = ~n5215 ;
  assign y6004 = ~1'b0 ;
  assign y6005 = 1'b0 ;
  assign y6006 = ~n11551 ;
  assign y6007 = n11555 ;
  assign y6008 = ~n11557 ;
  assign y6009 = ~1'b0 ;
  assign y6010 = ~n11559 ;
  assign y6011 = ~n11560 ;
  assign y6012 = ~1'b0 ;
  assign y6013 = ~n11563 ;
  assign y6014 = ~n11564 ;
  assign y6015 = ~n11567 ;
  assign y6016 = n11570 ;
  assign y6017 = ~1'b0 ;
  assign y6018 = n5420 ;
  assign y6019 = ~1'b0 ;
  assign y6020 = n11580 ;
  assign y6021 = ~n11582 ;
  assign y6022 = n11583 ;
  assign y6023 = n11584 ;
  assign y6024 = ~1'b0 ;
  assign y6025 = ~n11589 ;
  assign y6026 = ~n11591 ;
  assign y6027 = n11593 ;
  assign y6028 = ~1'b0 ;
  assign y6029 = n11595 ;
  assign y6030 = ~1'b0 ;
  assign y6031 = ~n11600 ;
  assign y6032 = ~n11602 ;
  assign y6033 = ~n11607 ;
  assign y6034 = ~1'b0 ;
  assign y6035 = ~n11608 ;
  assign y6036 = ~n11610 ;
  assign y6037 = ~1'b0 ;
  assign y6038 = ~1'b0 ;
  assign y6039 = ~1'b0 ;
  assign y6040 = ~n11612 ;
  assign y6041 = ~1'b0 ;
  assign y6042 = ~1'b0 ;
  assign y6043 = ~n11613 ;
  assign y6044 = ~n11620 ;
  assign y6045 = ~n11621 ;
  assign y6046 = n11624 ;
  assign y6047 = n11625 ;
  assign y6048 = n11633 ;
  assign y6049 = ~n4357 ;
  assign y6050 = ~n11636 ;
  assign y6051 = n11640 ;
  assign y6052 = ~1'b0 ;
  assign y6053 = n6880 ;
  assign y6054 = ~n11642 ;
  assign y6055 = n11644 ;
  assign y6056 = ~n11651 ;
  assign y6057 = ~1'b0 ;
  assign y6058 = n11653 ;
  assign y6059 = ~n11656 ;
  assign y6060 = ~n11657 ;
  assign y6061 = ~1'b0 ;
  assign y6062 = ~n11659 ;
  assign y6063 = n11662 ;
  assign y6064 = ~n11667 ;
  assign y6065 = n11671 ;
  assign y6066 = ~1'b0 ;
  assign y6067 = ~n11676 ;
  assign y6068 = n10616 ;
  assign y6069 = ~n11688 ;
  assign y6070 = ~1'b0 ;
  assign y6071 = n11690 ;
  assign y6072 = n11692 ;
  assign y6073 = n11696 ;
  assign y6074 = n11697 ;
  assign y6075 = 1'b0 ;
  assign y6076 = ~1'b0 ;
  assign y6077 = n11698 ;
  assign y6078 = ~n11701 ;
  assign y6079 = ~n11702 ;
  assign y6080 = ~n11705 ;
  assign y6081 = n11715 ;
  assign y6082 = n11717 ;
  assign y6083 = ~n11721 ;
  assign y6084 = ~n11724 ;
  assign y6085 = ~1'b0 ;
  assign y6086 = ~n11727 ;
  assign y6087 = ~n11729 ;
  assign y6088 = ~n11732 ;
  assign y6089 = n1256 ;
  assign y6090 = ~n754 ;
  assign y6091 = ~n11735 ;
  assign y6092 = ~1'b0 ;
  assign y6093 = n11740 ;
  assign y6094 = ~n11741 ;
  assign y6095 = ~n10881 ;
  assign y6096 = ~n11743 ;
  assign y6097 = n8233 ;
  assign y6098 = ~n11744 ;
  assign y6099 = ~n11745 ;
  assign y6100 = ~n11749 ;
  assign y6101 = ~n11750 ;
  assign y6102 = ~n11751 ;
  assign y6103 = n10001 ;
  assign y6104 = ~1'b0 ;
  assign y6105 = ~n11752 ;
  assign y6106 = ~n11754 ;
  assign y6107 = ~1'b0 ;
  assign y6108 = ~1'b0 ;
  assign y6109 = ~n11759 ;
  assign y6110 = ~n11760 ;
  assign y6111 = n11761 ;
  assign y6112 = ~n11763 ;
  assign y6113 = ~1'b0 ;
  assign y6114 = ~1'b0 ;
  assign y6115 = ~1'b0 ;
  assign y6116 = ~1'b0 ;
  assign y6117 = n11764 ;
  assign y6118 = ~1'b0 ;
  assign y6119 = n11766 ;
  assign y6120 = ~n11771 ;
  assign y6121 = ~1'b0 ;
  assign y6122 = ~n11774 ;
  assign y6123 = n11776 ;
  assign y6124 = ~n11782 ;
  assign y6125 = n11783 ;
  assign y6126 = n11786 ;
  assign y6127 = n11789 ;
  assign y6128 = 1'b0 ;
  assign y6129 = n11791 ;
  assign y6130 = n11794 ;
  assign y6131 = n11795 ;
  assign y6132 = n11796 ;
  assign y6133 = n11798 ;
  assign y6134 = ~1'b0 ;
  assign y6135 = ~1'b0 ;
  assign y6136 = n11800 ;
  assign y6137 = ~n11801 ;
  assign y6138 = ~n11805 ;
  assign y6139 = ~n11809 ;
  assign y6140 = n11811 ;
  assign y6141 = n11812 ;
  assign y6142 = n11813 ;
  assign y6143 = ~n11815 ;
  assign y6144 = n11818 ;
  assign y6145 = ~n11822 ;
  assign y6146 = ~1'b0 ;
  assign y6147 = ~n11829 ;
  assign y6148 = ~n11831 ;
  assign y6149 = ~n3207 ;
  assign y6150 = ~n339 ;
  assign y6151 = ~n11832 ;
  assign y6152 = ~1'b0 ;
  assign y6153 = ~1'b0 ;
  assign y6154 = ~1'b0 ;
  assign y6155 = n11836 ;
  assign y6156 = n11841 ;
  assign y6157 = ~n11847 ;
  assign y6158 = n8970 ;
  assign y6159 = n11848 ;
  assign y6160 = ~1'b0 ;
  assign y6161 = ~1'b0 ;
  assign y6162 = ~1'b0 ;
  assign y6163 = n11849 ;
  assign y6164 = n11853 ;
  assign y6165 = ~1'b0 ;
  assign y6166 = ~1'b0 ;
  assign y6167 = ~n11854 ;
  assign y6168 = ~1'b0 ;
  assign y6169 = ~n11857 ;
  assign y6170 = ~n11858 ;
  assign y6171 = n11860 ;
  assign y6172 = ~n11861 ;
  assign y6173 = ~n11862 ;
  assign y6174 = ~1'b0 ;
  assign y6175 = ~1'b0 ;
  assign y6176 = ~1'b0 ;
  assign y6177 = n11868 ;
  assign y6178 = n11869 ;
  assign y6179 = n11872 ;
  assign y6180 = n11873 ;
  assign y6181 = ~1'b0 ;
  assign y6182 = ~1'b0 ;
  assign y6183 = ~n11874 ;
  assign y6184 = ~n3082 ;
  assign y6185 = n11879 ;
  assign y6186 = ~n11883 ;
  assign y6187 = n11884 ;
  assign y6188 = ~n11891 ;
  assign y6189 = ~1'b0 ;
  assign y6190 = ~n11898 ;
  assign y6191 = ~n11899 ;
  assign y6192 = ~1'b0 ;
  assign y6193 = ~n11906 ;
  assign y6194 = ~n11914 ;
  assign y6195 = n11917 ;
  assign y6196 = ~1'b0 ;
  assign y6197 = ~1'b0 ;
  assign y6198 = n11918 ;
  assign y6199 = ~1'b0 ;
  assign y6200 = n11923 ;
  assign y6201 = n11931 ;
  assign y6202 = n11935 ;
  assign y6203 = ~n11937 ;
  assign y6204 = ~n11938 ;
  assign y6205 = ~n11939 ;
  assign y6206 = ~n11943 ;
  assign y6207 = n11947 ;
  assign y6208 = n11948 ;
  assign y6209 = ~1'b0 ;
  assign y6210 = ~n11951 ;
  assign y6211 = ~n8853 ;
  assign y6212 = ~n11956 ;
  assign y6213 = ~1'b0 ;
  assign y6214 = n57 ;
  assign y6215 = ~n11958 ;
  assign y6216 = ~n2989 ;
  assign y6217 = ~n11959 ;
  assign y6218 = ~1'b0 ;
  assign y6219 = ~1'b0 ;
  assign y6220 = ~1'b0 ;
  assign y6221 = n11960 ;
  assign y6222 = ~1'b0 ;
  assign y6223 = ~n11967 ;
  assign y6224 = ~n11968 ;
  assign y6225 = n11969 ;
  assign y6226 = n11971 ;
  assign y6227 = n11972 ;
  assign y6228 = ~1'b0 ;
  assign y6229 = ~n11975 ;
  assign y6230 = ~1'b0 ;
  assign y6231 = ~n11978 ;
  assign y6232 = n11980 ;
  assign y6233 = n11998 ;
  assign y6234 = ~1'b0 ;
  assign y6235 = n11999 ;
  assign y6236 = n12000 ;
  assign y6237 = n12003 ;
  assign y6238 = ~n12004 ;
  assign y6239 = n9369 ;
  assign y6240 = ~n448 ;
  assign y6241 = ~n12006 ;
  assign y6242 = ~1'b0 ;
  assign y6243 = ~n12007 ;
  assign y6244 = ~n12009 ;
  assign y6245 = ~n12011 ;
  assign y6246 = n12026 ;
  assign y6247 = n12030 ;
  assign y6248 = ~n12032 ;
  assign y6249 = ~n12034 ;
  assign y6250 = ~1'b0 ;
  assign y6251 = ~1'b0 ;
  assign y6252 = ~n12036 ;
  assign y6253 = n12037 ;
  assign y6254 = ~n7626 ;
  assign y6255 = ~1'b0 ;
  assign y6256 = ~n12038 ;
  assign y6257 = ~n9098 ;
  assign y6258 = n12040 ;
  assign y6259 = ~n12043 ;
  assign y6260 = ~n12046 ;
  assign y6261 = ~n12053 ;
  assign y6262 = n12056 ;
  assign y6263 = n12058 ;
  assign y6264 = n9208 ;
  assign y6265 = n12060 ;
  assign y6266 = ~n12065 ;
  assign y6267 = n12078 ;
  assign y6268 = ~n4567 ;
  assign y6269 = ~n12079 ;
  assign y6270 = ~n12081 ;
  assign y6271 = n12082 ;
  assign y6272 = ~n12086 ;
  assign y6273 = ~n7375 ;
  assign y6274 = ~n12091 ;
  assign y6275 = ~1'b0 ;
  assign y6276 = ~1'b0 ;
  assign y6277 = ~1'b0 ;
  assign y6278 = n12092 ;
  assign y6279 = ~1'b0 ;
  assign y6280 = ~n12095 ;
  assign y6281 = ~n676 ;
  assign y6282 = ~n12099 ;
  assign y6283 = n12101 ;
  assign y6284 = n12104 ;
  assign y6285 = ~n12106 ;
  assign y6286 = n12107 ;
  assign y6287 = 1'b0 ;
  assign y6288 = ~n12113 ;
  assign y6289 = n12114 ;
  assign y6290 = ~n12117 ;
  assign y6291 = ~1'b0 ;
  assign y6292 = ~n12119 ;
  assign y6293 = n12122 ;
  assign y6294 = n12123 ;
  assign y6295 = ~n12132 ;
  assign y6296 = ~1'b0 ;
  assign y6297 = n11908 ;
  assign y6298 = ~1'b0 ;
  assign y6299 = n12133 ;
  assign y6300 = n8659 ;
  assign y6301 = n12134 ;
  assign y6302 = n2835 ;
  assign y6303 = ~n12138 ;
  assign y6304 = ~n12141 ;
  assign y6305 = n12144 ;
  assign y6306 = ~1'b0 ;
  assign y6307 = ~n12145 ;
  assign y6308 = ~n12154 ;
  assign y6309 = ~n12155 ;
  assign y6310 = ~n12156 ;
  assign y6311 = ~n12160 ;
  assign y6312 = ~n6502 ;
  assign y6313 = n12162 ;
  assign y6314 = n12165 ;
  assign y6315 = ~n12166 ;
  assign y6316 = n12168 ;
  assign y6317 = ~n8452 ;
  assign y6318 = ~n12171 ;
  assign y6319 = ~n12175 ;
  assign y6320 = n12176 ;
  assign y6321 = n12177 ;
  assign y6322 = ~n12179 ;
  assign y6323 = ~n12180 ;
  assign y6324 = n12181 ;
  assign y6325 = ~1'b0 ;
  assign y6326 = n12187 ;
  assign y6327 = ~n12189 ;
  assign y6328 = ~n12196 ;
  assign y6329 = n10277 ;
  assign y6330 = ~n12197 ;
  assign y6331 = ~n4510 ;
  assign y6332 = ~1'b0 ;
  assign y6333 = ~1'b0 ;
  assign y6334 = ~1'b0 ;
  assign y6335 = n12198 ;
  assign y6336 = ~1'b0 ;
  assign y6337 = ~n12201 ;
  assign y6338 = ~1'b0 ;
  assign y6339 = n12208 ;
  assign y6340 = ~1'b0 ;
  assign y6341 = ~1'b0 ;
  assign y6342 = n12215 ;
  assign y6343 = ~n12217 ;
  assign y6344 = n12222 ;
  assign y6345 = n12225 ;
  assign y6346 = n1360 ;
  assign y6347 = n12230 ;
  assign y6348 = n12234 ;
  assign y6349 = ~1'b0 ;
  assign y6350 = 1'b0 ;
  assign y6351 = ~n12236 ;
  assign y6352 = n12237 ;
  assign y6353 = n12238 ;
  assign y6354 = n12244 ;
  assign y6355 = ~n12253 ;
  assign y6356 = n12264 ;
  assign y6357 = ~1'b0 ;
  assign y6358 = ~1'b0 ;
  assign y6359 = 1'b0 ;
  assign y6360 = n12270 ;
  assign y6361 = n12271 ;
  assign y6362 = n12274 ;
  assign y6363 = ~n12279 ;
  assign y6364 = ~1'b0 ;
  assign y6365 = ~1'b0 ;
  assign y6366 = ~n12282 ;
  assign y6367 = ~1'b0 ;
  assign y6368 = n8433 ;
  assign y6369 = ~n12283 ;
  assign y6370 = ~1'b0 ;
  assign y6371 = ~n12285 ;
  assign y6372 = ~1'b0 ;
  assign y6373 = n12288 ;
  assign y6374 = ~n12289 ;
  assign y6375 = n2801 ;
  assign y6376 = ~1'b0 ;
  assign y6377 = n12291 ;
  assign y6378 = ~1'b0 ;
  assign y6379 = ~1'b0 ;
  assign y6380 = n12294 ;
  assign y6381 = ~n12297 ;
  assign y6382 = ~1'b0 ;
  assign y6383 = n12298 ;
  assign y6384 = ~n12300 ;
  assign y6385 = ~1'b0 ;
  assign y6386 = ~n12301 ;
  assign y6387 = ~1'b0 ;
  assign y6388 = ~n12305 ;
  assign y6389 = ~n12307 ;
  assign y6390 = ~n12317 ;
  assign y6391 = n12319 ;
  assign y6392 = n12321 ;
  assign y6393 = n12322 ;
  assign y6394 = ~1'b0 ;
  assign y6395 = n12324 ;
  assign y6396 = ~1'b0 ;
  assign y6397 = ~n12326 ;
  assign y6398 = n12330 ;
  assign y6399 = n12333 ;
  assign y6400 = n12338 ;
  assign y6401 = ~n261 ;
  assign y6402 = ~n12340 ;
  assign y6403 = n12343 ;
  assign y6404 = ~n12344 ;
  assign y6405 = n12347 ;
  assign y6406 = n12350 ;
  assign y6407 = ~n12354 ;
  assign y6408 = ~n12356 ;
  assign y6409 = n12358 ;
  assign y6410 = ~n12360 ;
  assign y6411 = n12361 ;
  assign y6412 = n12364 ;
  assign y6413 = ~1'b0 ;
  assign y6414 = ~1'b0 ;
  assign y6415 = ~n12365 ;
  assign y6416 = n12369 ;
  assign y6417 = n12371 ;
  assign y6418 = ~1'b0 ;
  assign y6419 = n12374 ;
  assign y6420 = ~1'b0 ;
  assign y6421 = n12375 ;
  assign y6422 = ~n12376 ;
  assign y6423 = ~1'b0 ;
  assign y6424 = ~n12382 ;
  assign y6425 = ~n12383 ;
  assign y6426 = n12387 ;
  assign y6427 = n12391 ;
  assign y6428 = n12395 ;
  assign y6429 = ~n12405 ;
  assign y6430 = ~n9546 ;
  assign y6431 = ~n12406 ;
  assign y6432 = 1'b0 ;
  assign y6433 = ~n12407 ;
  assign y6434 = ~1'b0 ;
  assign y6435 = 1'b0 ;
  assign y6436 = ~1'b0 ;
  assign y6437 = n12408 ;
  assign y6438 = ~1'b0 ;
  assign y6439 = n12411 ;
  assign y6440 = ~n12413 ;
  assign y6441 = ~n12415 ;
  assign y6442 = ~1'b0 ;
  assign y6443 = ~1'b0 ;
  assign y6444 = ~n12418 ;
  assign y6445 = n12419 ;
  assign y6446 = ~n12421 ;
  assign y6447 = ~n12425 ;
  assign y6448 = ~1'b0 ;
  assign y6449 = ~n12428 ;
  assign y6450 = n12433 ;
  assign y6451 = ~1'b0 ;
  assign y6452 = n12438 ;
  assign y6453 = ~1'b0 ;
  assign y6454 = ~n12444 ;
  assign y6455 = ~n12446 ;
  assign y6456 = ~1'b0 ;
  assign y6457 = n12448 ;
  assign y6458 = n12451 ;
  assign y6459 = ~1'b0 ;
  assign y6460 = n12456 ;
  assign y6461 = ~n12458 ;
  assign y6462 = ~n12460 ;
  assign y6463 = n12461 ;
  assign y6464 = ~1'b0 ;
  assign y6465 = ~1'b0 ;
  assign y6466 = ~n12463 ;
  assign y6467 = ~n12466 ;
  assign y6468 = n12470 ;
  assign y6469 = n12477 ;
  assign y6470 = ~n12482 ;
  assign y6471 = ~1'b0 ;
  assign y6472 = n12483 ;
  assign y6473 = n12485 ;
  assign y6474 = 1'b0 ;
  assign y6475 = n12488 ;
  assign y6476 = n12490 ;
  assign y6477 = n12495 ;
  assign y6478 = ~n12496 ;
  assign y6479 = ~1'b0 ;
  assign y6480 = ~1'b0 ;
  assign y6481 = ~n12497 ;
  assign y6482 = ~1'b0 ;
  assign y6483 = ~1'b0 ;
  assign y6484 = ~n12499 ;
  assign y6485 = n12510 ;
  assign y6486 = 1'b0 ;
  assign y6487 = ~1'b0 ;
  assign y6488 = ~1'b0 ;
  assign y6489 = ~n12517 ;
  assign y6490 = n12519 ;
  assign y6491 = ~1'b0 ;
  assign y6492 = n12520 ;
  assign y6493 = ~n12521 ;
  assign y6494 = ~n12523 ;
  assign y6495 = ~n12531 ;
  assign y6496 = ~n12533 ;
  assign y6497 = ~1'b0 ;
  assign y6498 = n12534 ;
  assign y6499 = ~n12535 ;
  assign y6500 = ~n12543 ;
  assign y6501 = ~1'b0 ;
  assign y6502 = n12546 ;
  assign y6503 = n6551 ;
  assign y6504 = n12547 ;
  assign y6505 = ~n12548 ;
  assign y6506 = n12553 ;
  assign y6507 = ~1'b0 ;
  assign y6508 = 1'b0 ;
  assign y6509 = ~n12555 ;
  assign y6510 = ~n12559 ;
  assign y6511 = n12562 ;
  assign y6512 = ~n12565 ;
  assign y6513 = n12566 ;
  assign y6514 = ~1'b0 ;
  assign y6515 = ~1'b0 ;
  assign y6516 = n12568 ;
  assign y6517 = n12572 ;
  assign y6518 = n12580 ;
  assign y6519 = ~1'b0 ;
  assign y6520 = n2195 ;
  assign y6521 = ~1'b0 ;
  assign y6522 = n1615 ;
  assign y6523 = ~n12583 ;
  assign y6524 = n12585 ;
  assign y6525 = n12586 ;
  assign y6526 = ~1'b0 ;
  assign y6527 = n12588 ;
  assign y6528 = ~1'b0 ;
  assign y6529 = ~1'b0 ;
  assign y6530 = ~n12592 ;
  assign y6531 = n12593 ;
  assign y6532 = ~n12595 ;
  assign y6533 = n12598 ;
  assign y6534 = ~1'b0 ;
  assign y6535 = n9584 ;
  assign y6536 = ~1'b0 ;
  assign y6537 = n9606 ;
  assign y6538 = n12602 ;
  assign y6539 = ~1'b0 ;
  assign y6540 = ~1'b0 ;
  assign y6541 = ~n12611 ;
  assign y6542 = ~n12612 ;
  assign y6543 = ~n12614 ;
  assign y6544 = n12622 ;
  assign y6545 = n12623 ;
  assign y6546 = ~1'b0 ;
  assign y6547 = n12626 ;
  assign y6548 = n12630 ;
  assign y6549 = n12632 ;
  assign y6550 = n12633 ;
  assign y6551 = ~n12635 ;
  assign y6552 = ~1'b0 ;
  assign y6553 = ~n12636 ;
  assign y6554 = n12638 ;
  assign y6555 = n12643 ;
  assign y6556 = ~1'b0 ;
  assign y6557 = ~1'b0 ;
  assign y6558 = n12644 ;
  assign y6559 = ~n9247 ;
  assign y6560 = n12646 ;
  assign y6561 = ~n12649 ;
  assign y6562 = ~n12651 ;
  assign y6563 = ~n12652 ;
  assign y6564 = n12653 ;
  assign y6565 = n12658 ;
  assign y6566 = n12660 ;
  assign y6567 = ~n12662 ;
  assign y6568 = n12669 ;
  assign y6569 = ~1'b0 ;
  assign y6570 = 1'b0 ;
  assign y6571 = ~n12671 ;
  assign y6572 = ~n12675 ;
  assign y6573 = ~n12678 ;
  assign y6574 = ~1'b0 ;
  assign y6575 = ~n12679 ;
  assign y6576 = ~n12680 ;
  assign y6577 = ~1'b0 ;
  assign y6578 = n12681 ;
  assign y6579 = n12682 ;
  assign y6580 = n12683 ;
  assign y6581 = ~n812 ;
  assign y6582 = ~n12689 ;
  assign y6583 = ~n12694 ;
  assign y6584 = ~1'b0 ;
  assign y6585 = ~1'b0 ;
  assign y6586 = n5566 ;
  assign y6587 = ~n12698 ;
  assign y6588 = n11243 ;
  assign y6589 = ~n4593 ;
  assign y6590 = n12700 ;
  assign y6591 = ~1'b0 ;
  assign y6592 = n10298 ;
  assign y6593 = ~n12702 ;
  assign y6594 = n2934 ;
  assign y6595 = n12704 ;
  assign y6596 = n12705 ;
  assign y6597 = ~n12712 ;
  assign y6598 = ~1'b0 ;
  assign y6599 = n12713 ;
  assign y6600 = ~n12716 ;
  assign y6601 = ~n12723 ;
  assign y6602 = ~n12727 ;
  assign y6603 = ~n12731 ;
  assign y6604 = n12733 ;
  assign y6605 = n12735 ;
  assign y6606 = n12738 ;
  assign y6607 = ~n12742 ;
  assign y6608 = ~n12746 ;
  assign y6609 = n12747 ;
  assign y6610 = ~n12755 ;
  assign y6611 = n12758 ;
  assign y6612 = ~n12762 ;
  assign y6613 = ~1'b0 ;
  assign y6614 = ~1'b0 ;
  assign y6615 = n12767 ;
  assign y6616 = ~1'b0 ;
  assign y6617 = ~1'b0 ;
  assign y6618 = ~n12770 ;
  assign y6619 = ~1'b0 ;
  assign y6620 = n8436 ;
  assign y6621 = ~1'b0 ;
  assign y6622 = n12777 ;
  assign y6623 = ~1'b0 ;
  assign y6624 = ~1'b0 ;
  assign y6625 = ~n12779 ;
  assign y6626 = ~n6981 ;
  assign y6627 = n12781 ;
  assign y6628 = ~1'b0 ;
  assign y6629 = ~1'b0 ;
  assign y6630 = n11458 ;
  assign y6631 = ~n12782 ;
  assign y6632 = ~n12784 ;
  assign y6633 = n12788 ;
  assign y6634 = n12790 ;
  assign y6635 = ~n10211 ;
  assign y6636 = ~1'b0 ;
  assign y6637 = ~1'b0 ;
  assign y6638 = ~1'b0 ;
  assign y6639 = ~n12791 ;
  assign y6640 = n12794 ;
  assign y6641 = ~n1167 ;
  assign y6642 = n12796 ;
  assign y6643 = ~n12800 ;
  assign y6644 = ~1'b0 ;
  assign y6645 = ~n12802 ;
  assign y6646 = ~n12804 ;
  assign y6647 = ~n12805 ;
  assign y6648 = ~n12809 ;
  assign y6649 = ~n12814 ;
  assign y6650 = n12815 ;
  assign y6651 = n12816 ;
  assign y6652 = ~1'b0 ;
  assign y6653 = n453 ;
  assign y6654 = n12823 ;
  assign y6655 = ~n12825 ;
  assign y6656 = n12826 ;
  assign y6657 = n12830 ;
  assign y6658 = ~1'b0 ;
  assign y6659 = ~n2610 ;
  assign y6660 = ~n12833 ;
  assign y6661 = n1908 ;
  assign y6662 = ~1'b0 ;
  assign y6663 = ~1'b0 ;
  assign y6664 = n12835 ;
  assign y6665 = ~1'b0 ;
  assign y6666 = n12836 ;
  assign y6667 = ~n12837 ;
  assign y6668 = ~1'b0 ;
  assign y6669 = ~n12847 ;
  assign y6670 = ~n12853 ;
  assign y6671 = ~1'b0 ;
  assign y6672 = ~n12858 ;
  assign y6673 = ~n12867 ;
  assign y6674 = n12871 ;
  assign y6675 = ~n12873 ;
  assign y6676 = ~1'b0 ;
  assign y6677 = ~n12875 ;
  assign y6678 = ~n12878 ;
  assign y6679 = n12879 ;
  assign y6680 = 1'b0 ;
  assign y6681 = ~n12883 ;
  assign y6682 = ~n12885 ;
  assign y6683 = ~1'b0 ;
  assign y6684 = ~1'b0 ;
  assign y6685 = ~n12889 ;
  assign y6686 = n1251 ;
  assign y6687 = n12893 ;
  assign y6688 = ~1'b0 ;
  assign y6689 = 1'b0 ;
  assign y6690 = ~n12896 ;
  assign y6691 = ~n12897 ;
  assign y6692 = ~n12903 ;
  assign y6693 = ~n12911 ;
  assign y6694 = n12913 ;
  assign y6695 = ~1'b0 ;
  assign y6696 = ~1'b0 ;
  assign y6697 = ~n1517 ;
  assign y6698 = ~n5809 ;
  assign y6699 = ~1'b0 ;
  assign y6700 = ~1'b0 ;
  assign y6701 = n12914 ;
  assign y6702 = ~n12916 ;
  assign y6703 = 1'b0 ;
  assign y6704 = ~1'b0 ;
  assign y6705 = ~1'b0 ;
  assign y6706 = n4242 ;
  assign y6707 = ~n12917 ;
  assign y6708 = ~n10059 ;
  assign y6709 = ~n12920 ;
  assign y6710 = ~1'b0 ;
  assign y6711 = ~1'b0 ;
  assign y6712 = 1'b0 ;
  assign y6713 = n12925 ;
  assign y6714 = ~1'b0 ;
  assign y6715 = 1'b0 ;
  assign y6716 = n12929 ;
  assign y6717 = ~n12930 ;
  assign y6718 = ~1'b0 ;
  assign y6719 = n3600 ;
  assign y6720 = n12931 ;
  assign y6721 = ~n12937 ;
  assign y6722 = n12938 ;
  assign y6723 = ~n7804 ;
  assign y6724 = ~n12939 ;
  assign y6725 = n12942 ;
  assign y6726 = ~n12944 ;
  assign y6727 = 1'b0 ;
  assign y6728 = ~n12945 ;
  assign y6729 = ~1'b0 ;
  assign y6730 = ~n12947 ;
  assign y6731 = ~n12949 ;
  assign y6732 = ~n12952 ;
  assign y6733 = n12964 ;
  assign y6734 = ~1'b0 ;
  assign y6735 = ~n9363 ;
  assign y6736 = n12966 ;
  assign y6737 = n11458 ;
  assign y6738 = ~1'b0 ;
  assign y6739 = ~n12967 ;
  assign y6740 = ~n12968 ;
  assign y6741 = ~1'b0 ;
  assign y6742 = ~n12969 ;
  assign y6743 = n12970 ;
  assign y6744 = n12972 ;
  assign y6745 = n12974 ;
  assign y6746 = n12977 ;
  assign y6747 = n12984 ;
  assign y6748 = n4041 ;
  assign y6749 = ~1'b0 ;
  assign y6750 = n12986 ;
  assign y6751 = n12987 ;
  assign y6752 = ~1'b0 ;
  assign y6753 = n12991 ;
  assign y6754 = n13000 ;
  assign y6755 = ~1'b0 ;
  assign y6756 = ~1'b0 ;
  assign y6757 = n13008 ;
  assign y6758 = ~n13010 ;
  assign y6759 = n13013 ;
  assign y6760 = ~1'b0 ;
  assign y6761 = n13015 ;
  assign y6762 = n13017 ;
  assign y6763 = ~1'b0 ;
  assign y6764 = n13018 ;
  assign y6765 = ~1'b0 ;
  assign y6766 = n13019 ;
  assign y6767 = n13023 ;
  assign y6768 = ~1'b0 ;
  assign y6769 = ~n2415 ;
  assign y6770 = ~n13030 ;
  assign y6771 = n13035 ;
  assign y6772 = n13036 ;
  assign y6773 = ~n13041 ;
  assign y6774 = n13046 ;
  assign y6775 = n13053 ;
  assign y6776 = ~1'b0 ;
  assign y6777 = ~1'b0 ;
  assign y6778 = ~n13060 ;
  assign y6779 = n13061 ;
  assign y6780 = ~n2154 ;
  assign y6781 = ~1'b0 ;
  assign y6782 = ~n13062 ;
  assign y6783 = n13063 ;
  assign y6784 = ~1'b0 ;
  assign y6785 = ~1'b0 ;
  assign y6786 = ~1'b0 ;
  assign y6787 = n13066 ;
  assign y6788 = n13073 ;
  assign y6789 = n13075 ;
  assign y6790 = ~n3226 ;
  assign y6791 = ~n13077 ;
  assign y6792 = ~1'b0 ;
  assign y6793 = n13079 ;
  assign y6794 = n13080 ;
  assign y6795 = ~n13081 ;
  assign y6796 = ~n13082 ;
  assign y6797 = ~n13086 ;
  assign y6798 = ~1'b0 ;
  assign y6799 = ~1'b0 ;
  assign y6800 = ~n13089 ;
  assign y6801 = ~1'b0 ;
  assign y6802 = ~n13092 ;
  assign y6803 = n13094 ;
  assign y6804 = n13095 ;
  assign y6805 = ~1'b0 ;
  assign y6806 = ~n13096 ;
  assign y6807 = n5756 ;
  assign y6808 = ~1'b0 ;
  assign y6809 = ~n13102 ;
  assign y6810 = n13103 ;
  assign y6811 = ~1'b0 ;
  assign y6812 = 1'b0 ;
  assign y6813 = ~n13110 ;
  assign y6814 = n13112 ;
  assign y6815 = ~1'b0 ;
  assign y6816 = n13114 ;
  assign y6817 = ~n13115 ;
  assign y6818 = ~n13117 ;
  assign y6819 = ~1'b0 ;
  assign y6820 = ~n13120 ;
  assign y6821 = n13123 ;
  assign y6822 = ~n13125 ;
  assign y6823 = n13126 ;
  assign y6824 = ~1'b0 ;
  assign y6825 = ~1'b0 ;
  assign y6826 = ~n13129 ;
  assign y6827 = ~1'b0 ;
  assign y6828 = n13131 ;
  assign y6829 = ~n13133 ;
  assign y6830 = 1'b0 ;
  assign y6831 = ~1'b0 ;
  assign y6832 = n13137 ;
  assign y6833 = ~1'b0 ;
  assign y6834 = ~n13138 ;
  assign y6835 = n13140 ;
  assign y6836 = ~1'b0 ;
  assign y6837 = ~1'b0 ;
  assign y6838 = ~1'b0 ;
  assign y6839 = ~n13143 ;
  assign y6840 = ~n13144 ;
  assign y6841 = ~n13146 ;
  assign y6842 = ~n13165 ;
  assign y6843 = ~1'b0 ;
  assign y6844 = ~1'b0 ;
  assign y6845 = ~1'b0 ;
  assign y6846 = ~n13167 ;
  assign y6847 = n13168 ;
  assign y6848 = n13171 ;
  assign y6849 = ~n13172 ;
  assign y6850 = ~1'b0 ;
  assign y6851 = ~1'b0 ;
  assign y6852 = ~1'b0 ;
  assign y6853 = ~n13173 ;
  assign y6854 = ~1'b0 ;
  assign y6855 = ~1'b0 ;
  assign y6856 = ~n13176 ;
  assign y6857 = ~n13177 ;
  assign y6858 = ~n13179 ;
  assign y6859 = n13181 ;
  assign y6860 = ~1'b0 ;
  assign y6861 = ~1'b0 ;
  assign y6862 = ~1'b0 ;
  assign y6863 = ~n13182 ;
  assign y6864 = ~1'b0 ;
  assign y6865 = n13184 ;
  assign y6866 = ~1'b0 ;
  assign y6867 = ~1'b0 ;
  assign y6868 = n12593 ;
  assign y6869 = n13185 ;
  assign y6870 = n6917 ;
  assign y6871 = n13188 ;
  assign y6872 = 1'b0 ;
  assign y6873 = ~n13192 ;
  assign y6874 = n13194 ;
  assign y6875 = ~1'b0 ;
  assign y6876 = ~n13202 ;
  assign y6877 = ~n13203 ;
  assign y6878 = ~1'b0 ;
  assign y6879 = ~n13204 ;
  assign y6880 = ~1'b0 ;
  assign y6881 = ~n13207 ;
  assign y6882 = ~n13208 ;
  assign y6883 = ~n13210 ;
  assign y6884 = ~1'b0 ;
  assign y6885 = n13216 ;
  assign y6886 = n13218 ;
  assign y6887 = ~n13224 ;
  assign y6888 = ~1'b0 ;
  assign y6889 = ~n13230 ;
  assign y6890 = ~n13231 ;
  assign y6891 = ~n13234 ;
  assign y6892 = n7556 ;
  assign y6893 = ~n13236 ;
  assign y6894 = n13237 ;
  assign y6895 = n13242 ;
  assign y6896 = ~1'b0 ;
  assign y6897 = n8926 ;
  assign y6898 = ~n13246 ;
  assign y6899 = n13247 ;
  assign y6900 = n13248 ;
  assign y6901 = n13249 ;
  assign y6902 = n13254 ;
  assign y6903 = ~n13255 ;
  assign y6904 = n13256 ;
  assign y6905 = ~1'b0 ;
  assign y6906 = ~n13257 ;
  assign y6907 = ~1'b0 ;
  assign y6908 = ~n13259 ;
  assign y6909 = ~1'b0 ;
  assign y6910 = ~n6762 ;
  assign y6911 = ~n1035 ;
  assign y6912 = ~1'b0 ;
  assign y6913 = n13261 ;
  assign y6914 = ~1'b0 ;
  assign y6915 = n13262 ;
  assign y6916 = ~n13263 ;
  assign y6917 = n13269 ;
  assign y6918 = n13270 ;
  assign y6919 = n13274 ;
  assign y6920 = ~1'b0 ;
  assign y6921 = ~n13277 ;
  assign y6922 = n13285 ;
  assign y6923 = ~n13292 ;
  assign y6924 = x7 ;
  assign y6925 = n13295 ;
  assign y6926 = n13296 ;
  assign y6927 = ~n13302 ;
  assign y6928 = ~1'b0 ;
  assign y6929 = n13303 ;
  assign y6930 = ~n13306 ;
  assign y6931 = n13308 ;
  assign y6932 = ~1'b0 ;
  assign y6933 = n13314 ;
  assign y6934 = n5613 ;
  assign y6935 = ~n13317 ;
  assign y6936 = n790 ;
  assign y6937 = ~n13274 ;
  assign y6938 = ~n13320 ;
  assign y6939 = n13322 ;
  assign y6940 = n12825 ;
  assign y6941 = n13323 ;
  assign y6942 = ~1'b0 ;
  assign y6943 = ~n13325 ;
  assign y6944 = ~n13327 ;
  assign y6945 = ~1'b0 ;
  assign y6946 = n13328 ;
  assign y6947 = n13330 ;
  assign y6948 = ~1'b0 ;
  assign y6949 = n13332 ;
  assign y6950 = ~1'b0 ;
  assign y6951 = ~1'b0 ;
  assign y6952 = n13335 ;
  assign y6953 = ~1'b0 ;
  assign y6954 = ~n13338 ;
  assign y6955 = 1'b0 ;
  assign y6956 = n13340 ;
  assign y6957 = n13345 ;
  assign y6958 = ~n12637 ;
  assign y6959 = n13346 ;
  assign y6960 = ~n13349 ;
  assign y6961 = n13350 ;
  assign y6962 = n13354 ;
  assign y6963 = ~n13356 ;
  assign y6964 = n13357 ;
  assign y6965 = n10357 ;
  assign y6966 = ~n13358 ;
  assign y6967 = ~n13361 ;
  assign y6968 = ~1'b0 ;
  assign y6969 = ~1'b0 ;
  assign y6970 = ~n13364 ;
  assign y6971 = n13366 ;
  assign y6972 = n13373 ;
  assign y6973 = n13377 ;
  assign y6974 = ~n13379 ;
  assign y6975 = ~n13381 ;
  assign y6976 = ~n13385 ;
  assign y6977 = n13386 ;
  assign y6978 = n10792 ;
  assign y6979 = ~n13388 ;
  assign y6980 = ~n13390 ;
  assign y6981 = ~1'b0 ;
  assign y6982 = n10146 ;
  assign y6983 = ~n13391 ;
  assign y6984 = ~n13392 ;
  assign y6985 = ~n13394 ;
  assign y6986 = ~1'b0 ;
  assign y6987 = n13395 ;
  assign y6988 = ~1'b0 ;
  assign y6989 = n13399 ;
  assign y6990 = ~1'b0 ;
  assign y6991 = n13400 ;
  assign y6992 = n13408 ;
  assign y6993 = ~n4044 ;
  assign y6994 = ~1'b0 ;
  assign y6995 = ~1'b0 ;
  assign y6996 = ~n13413 ;
  assign y6997 = ~1'b0 ;
  assign y6998 = n13415 ;
  assign y6999 = n13417 ;
  assign y7000 = ~1'b0 ;
  assign y7001 = 1'b0 ;
  assign y7002 = ~n13419 ;
  assign y7003 = ~1'b0 ;
  assign y7004 = ~1'b0 ;
  assign y7005 = n13422 ;
  assign y7006 = ~1'b0 ;
  assign y7007 = ~n13424 ;
  assign y7008 = n13425 ;
  assign y7009 = n13427 ;
  assign y7010 = ~n13430 ;
  assign y7011 = ~1'b0 ;
  assign y7012 = ~1'b0 ;
  assign y7013 = n13434 ;
  assign y7014 = n13436 ;
  assign y7015 = n13437 ;
  assign y7016 = ~1'b0 ;
  assign y7017 = n13440 ;
  assign y7018 = ~n13441 ;
  assign y7019 = ~1'b0 ;
  assign y7020 = n13442 ;
  assign y7021 = ~1'b0 ;
  assign y7022 = n13443 ;
  assign y7023 = ~1'b0 ;
  assign y7024 = ~n13447 ;
  assign y7025 = ~n13454 ;
  assign y7026 = ~1'b0 ;
  assign y7027 = ~n13458 ;
  assign y7028 = n13460 ;
  assign y7029 = ~n12735 ;
  assign y7030 = n3049 ;
  assign y7031 = n13463 ;
  assign y7032 = ~n13464 ;
  assign y7033 = ~1'b0 ;
  assign y7034 = ~1'b0 ;
  assign y7035 = ~1'b0 ;
  assign y7036 = ~n13470 ;
  assign y7037 = ~n13471 ;
  assign y7038 = n13473 ;
  assign y7039 = n13474 ;
  assign y7040 = ~n13478 ;
  assign y7041 = ~n13479 ;
  assign y7042 = ~n13481 ;
  assign y7043 = ~n13482 ;
  assign y7044 = ~1'b0 ;
  assign y7045 = ~1'b0 ;
  assign y7046 = ~1'b0 ;
  assign y7047 = ~1'b0 ;
  assign y7048 = ~n13485 ;
  assign y7049 = n13487 ;
  assign y7050 = n13489 ;
  assign y7051 = ~n13500 ;
  assign y7052 = n13501 ;
  assign y7053 = n13503 ;
  assign y7054 = n13508 ;
  assign y7055 = ~1'b0 ;
  assign y7056 = ~n13511 ;
  assign y7057 = n13520 ;
  assign y7058 = ~n13523 ;
  assign y7059 = ~n13524 ;
  assign y7060 = ~n13527 ;
  assign y7061 = n13528 ;
  assign y7062 = n13535 ;
  assign y7063 = ~n13539 ;
  assign y7064 = ~1'b0 ;
  assign y7065 = n13545 ;
  assign y7066 = ~1'b0 ;
  assign y7067 = ~n3071 ;
  assign y7068 = ~1'b0 ;
  assign y7069 = ~n13549 ;
  assign y7070 = ~1'b0 ;
  assign y7071 = ~n13550 ;
  assign y7072 = ~1'b0 ;
  assign y7073 = ~n13561 ;
  assign y7074 = 1'b0 ;
  assign y7075 = ~n13562 ;
  assign y7076 = ~n6465 ;
  assign y7077 = ~1'b0 ;
  assign y7078 = n13569 ;
  assign y7079 = ~1'b0 ;
  assign y7080 = ~1'b0 ;
  assign y7081 = ~n13573 ;
  assign y7082 = ~1'b0 ;
  assign y7083 = ~1'b0 ;
  assign y7084 = ~n13575 ;
  assign y7085 = ~n13579 ;
  assign y7086 = n13581 ;
  assign y7087 = n13583 ;
  assign y7088 = ~n13586 ;
  assign y7089 = ~n13589 ;
  assign y7090 = n13590 ;
  assign y7091 = n13592 ;
  assign y7092 = ~n13596 ;
  assign y7093 = ~n13598 ;
  assign y7094 = ~n13601 ;
  assign y7095 = ~n13606 ;
  assign y7096 = n13607 ;
  assign y7097 = ~n13611 ;
  assign y7098 = ~n12985 ;
  assign y7099 = n10166 ;
  assign y7100 = ~1'b0 ;
  assign y7101 = n13612 ;
  assign y7102 = n13613 ;
  assign y7103 = n13614 ;
  assign y7104 = ~1'b0 ;
  assign y7105 = ~1'b0 ;
  assign y7106 = ~1'b0 ;
  assign y7107 = n4931 ;
  assign y7108 = ~1'b0 ;
  assign y7109 = ~1'b0 ;
  assign y7110 = n13615 ;
  assign y7111 = ~1'b0 ;
  assign y7112 = ~n13617 ;
  assign y7113 = ~1'b0 ;
  assign y7114 = n13620 ;
  assign y7115 = ~1'b0 ;
  assign y7116 = ~1'b0 ;
  assign y7117 = ~n13623 ;
  assign y7118 = n2955 ;
  assign y7119 = ~1'b0 ;
  assign y7120 = ~1'b0 ;
  assign y7121 = n13625 ;
  assign y7122 = n13628 ;
  assign y7123 = ~n2185 ;
  assign y7124 = n13630 ;
  assign y7125 = n13634 ;
  assign y7126 = n13636 ;
  assign y7127 = ~n13637 ;
  assign y7128 = n13638 ;
  assign y7129 = ~n13639 ;
  assign y7130 = ~n13660 ;
  assign y7131 = ~1'b0 ;
  assign y7132 = n13661 ;
  assign y7133 = n13663 ;
  assign y7134 = ~n13665 ;
  assign y7135 = ~1'b0 ;
  assign y7136 = ~n13670 ;
  assign y7137 = ~n13673 ;
  assign y7138 = ~1'b0 ;
  assign y7139 = n13676 ;
  assign y7140 = ~1'b0 ;
  assign y7141 = n13677 ;
  assign y7142 = n13678 ;
  assign y7143 = ~n13684 ;
  assign y7144 = ~n13688 ;
  assign y7145 = 1'b0 ;
  assign y7146 = n13690 ;
  assign y7147 = ~1'b0 ;
  assign y7148 = ~n10403 ;
  assign y7149 = n13691 ;
  assign y7150 = ~1'b0 ;
  assign y7151 = ~n13692 ;
  assign y7152 = ~1'b0 ;
  assign y7153 = ~1'b0 ;
  assign y7154 = ~n13693 ;
  assign y7155 = ~n13694 ;
  assign y7156 = ~1'b0 ;
  assign y7157 = ~1'b0 ;
  assign y7158 = ~n4384 ;
  assign y7159 = 1'b0 ;
  assign y7160 = n13696 ;
  assign y7161 = ~1'b0 ;
  assign y7162 = ~n13701 ;
  assign y7163 = ~1'b0 ;
  assign y7164 = ~n13707 ;
  assign y7165 = ~n13710 ;
  assign y7166 = n13714 ;
  assign y7167 = ~1'b0 ;
  assign y7168 = ~n13719 ;
  assign y7169 = ~n13723 ;
  assign y7170 = n13724 ;
  assign y7171 = ~n13730 ;
  assign y7172 = ~1'b0 ;
  assign y7173 = ~1'b0 ;
  assign y7174 = n13732 ;
  assign y7175 = ~n13734 ;
  assign y7176 = n13735 ;
  assign y7177 = ~n13736 ;
  assign y7178 = ~1'b0 ;
  assign y7179 = ~n6256 ;
  assign y7180 = ~n13737 ;
  assign y7181 = ~n13740 ;
  assign y7182 = ~1'b0 ;
  assign y7183 = ~1'b0 ;
  assign y7184 = ~n13742 ;
  assign y7185 = ~n13743 ;
  assign y7186 = ~1'b0 ;
  assign y7187 = n13744 ;
  assign y7188 = n12576 ;
  assign y7189 = ~n13747 ;
  assign y7190 = 1'b0 ;
  assign y7191 = n13748 ;
  assign y7192 = ~n13750 ;
  assign y7193 = 1'b0 ;
  assign y7194 = ~n13751 ;
  assign y7195 = ~n13754 ;
  assign y7196 = n13755 ;
  assign y7197 = ~1'b0 ;
  assign y7198 = ~n13756 ;
  assign y7199 = ~1'b0 ;
  assign y7200 = n13760 ;
  assign y7201 = ~1'b0 ;
  assign y7202 = ~n13761 ;
  assign y7203 = ~n13762 ;
  assign y7204 = n13763 ;
  assign y7205 = ~n13769 ;
  assign y7206 = ~n13771 ;
  assign y7207 = 1'b0 ;
  assign y7208 = ~1'b0 ;
  assign y7209 = ~n13774 ;
  assign y7210 = ~n13778 ;
  assign y7211 = n13786 ;
  assign y7212 = ~1'b0 ;
  assign y7213 = ~n13789 ;
  assign y7214 = ~n13795 ;
  assign y7215 = ~n13800 ;
  assign y7216 = ~1'b0 ;
  assign y7217 = 1'b0 ;
  assign y7218 = n13803 ;
  assign y7219 = n13805 ;
  assign y7220 = ~n13806 ;
  assign y7221 = n13808 ;
  assign y7222 = n3197 ;
  assign y7223 = ~1'b0 ;
  assign y7224 = n13818 ;
  assign y7225 = ~1'b0 ;
  assign y7226 = ~1'b0 ;
  assign y7227 = ~n13820 ;
  assign y7228 = n10603 ;
  assign y7229 = ~1'b0 ;
  assign y7230 = ~1'b0 ;
  assign y7231 = n13823 ;
  assign y7232 = n13825 ;
  assign y7233 = ~n13827 ;
  assign y7234 = 1'b0 ;
  assign y7235 = n13828 ;
  assign y7236 = ~1'b0 ;
  assign y7237 = ~n2732 ;
  assign y7238 = ~n13829 ;
  assign y7239 = ~n13831 ;
  assign y7240 = n12747 ;
  assign y7241 = ~n13832 ;
  assign y7242 = n13835 ;
  assign y7243 = ~1'b0 ;
  assign y7244 = ~n13838 ;
  assign y7245 = ~1'b0 ;
  assign y7246 = ~n13840 ;
  assign y7247 = n13848 ;
  assign y7248 = ~1'b0 ;
  assign y7249 = ~n13849 ;
  assign y7250 = n13851 ;
  assign y7251 = ~1'b0 ;
  assign y7252 = n13854 ;
  assign y7253 = ~n13857 ;
  assign y7254 = n13860 ;
  assign y7255 = ~n13861 ;
  assign y7256 = ~1'b0 ;
  assign y7257 = ~n1469 ;
  assign y7258 = n13862 ;
  assign y7259 = n13863 ;
  assign y7260 = n13866 ;
  assign y7261 = ~1'b0 ;
  assign y7262 = ~n13869 ;
  assign y7263 = n13871 ;
  assign y7264 = ~n13875 ;
  assign y7265 = n13883 ;
  assign y7266 = ~n10364 ;
  assign y7267 = n13885 ;
  assign y7268 = ~n13889 ;
  assign y7269 = ~1'b0 ;
  assign y7270 = ~n13891 ;
  assign y7271 = ~n13893 ;
  assign y7272 = ~n13895 ;
  assign y7273 = ~n13896 ;
  assign y7274 = ~n13899 ;
  assign y7275 = n13900 ;
  assign y7276 = n13904 ;
  assign y7277 = n13907 ;
  assign y7278 = ~1'b0 ;
  assign y7279 = ~n13911 ;
  assign y7280 = ~1'b0 ;
  assign y7281 = ~1'b0 ;
  assign y7282 = ~1'b0 ;
  assign y7283 = ~n13912 ;
  assign y7284 = n13913 ;
  assign y7285 = ~n13915 ;
  assign y7286 = 1'b0 ;
  assign y7287 = ~1'b0 ;
  assign y7288 = n13916 ;
  assign y7289 = ~n13918 ;
  assign y7290 = n13919 ;
  assign y7291 = n13924 ;
  assign y7292 = ~n13925 ;
  assign y7293 = n13926 ;
  assign y7294 = ~1'b0 ;
  assign y7295 = ~n13927 ;
  assign y7296 = n13933 ;
  assign y7297 = ~1'b0 ;
  assign y7298 = n13934 ;
  assign y7299 = ~1'b0 ;
  assign y7300 = ~n13937 ;
  assign y7301 = n13939 ;
  assign y7302 = ~1'b0 ;
  assign y7303 = ~1'b0 ;
  assign y7304 = n13943 ;
  assign y7305 = n13944 ;
  assign y7306 = ~n13946 ;
  assign y7307 = n13949 ;
  assign y7308 = ~n13951 ;
  assign y7309 = ~1'b0 ;
  assign y7310 = n7624 ;
  assign y7311 = ~n13956 ;
  assign y7312 = n10031 ;
  assign y7313 = 1'b0 ;
  assign y7314 = ~1'b0 ;
  assign y7315 = n13960 ;
  assign y7316 = 1'b0 ;
  assign y7317 = ~n13490 ;
  assign y7318 = ~1'b0 ;
  assign y7319 = ~n13965 ;
  assign y7320 = ~n13968 ;
  assign y7321 = ~n8145 ;
  assign y7322 = ~1'b0 ;
  assign y7323 = ~n13971 ;
  assign y7324 = ~n13981 ;
  assign y7325 = ~n13984 ;
  assign y7326 = ~1'b0 ;
  assign y7327 = n13985 ;
  assign y7328 = ~n13986 ;
  assign y7329 = ~n13988 ;
  assign y7330 = ~n13990 ;
  assign y7331 = n11727 ;
  assign y7332 = ~n13991 ;
  assign y7333 = n14003 ;
  assign y7334 = 1'b0 ;
  assign y7335 = n14006 ;
  assign y7336 = n14010 ;
  assign y7337 = ~n14011 ;
  assign y7338 = n3837 ;
  assign y7339 = ~n14012 ;
  assign y7340 = ~1'b0 ;
  assign y7341 = ~n14013 ;
  assign y7342 = ~1'b0 ;
  assign y7343 = n14024 ;
  assign y7344 = n14028 ;
  assign y7345 = ~n14029 ;
  assign y7346 = ~n14030 ;
  assign y7347 = n14032 ;
  assign y7348 = ~n14038 ;
  assign y7349 = ~n14039 ;
  assign y7350 = ~1'b0 ;
  assign y7351 = 1'b0 ;
  assign y7352 = ~1'b0 ;
  assign y7353 = ~1'b0 ;
  assign y7354 = 1'b0 ;
  assign y7355 = ~1'b0 ;
  assign y7356 = ~1'b0 ;
  assign y7357 = n14041 ;
  assign y7358 = n214 ;
  assign y7359 = 1'b0 ;
  assign y7360 = ~n14042 ;
  assign y7361 = ~1'b0 ;
  assign y7362 = ~1'b0 ;
  assign y7363 = ~n14044 ;
  assign y7364 = n4952 ;
  assign y7365 = ~1'b0 ;
  assign y7366 = ~1'b0 ;
  assign y7367 = n14045 ;
  assign y7368 = ~n14046 ;
  assign y7369 = ~1'b0 ;
  assign y7370 = n14050 ;
  assign y7371 = n14054 ;
  assign y7372 = ~1'b0 ;
  assign y7373 = ~1'b0 ;
  assign y7374 = n14057 ;
  assign y7375 = ~1'b0 ;
  assign y7376 = ~n14064 ;
  assign y7377 = ~1'b0 ;
  assign y7378 = n14066 ;
  assign y7379 = ~n14067 ;
  assign y7380 = n14068 ;
  assign y7381 = n13594 ;
  assign y7382 = ~1'b0 ;
  assign y7383 = ~1'b0 ;
  assign y7384 = ~n14069 ;
  assign y7385 = n8034 ;
  assign y7386 = ~n14070 ;
  assign y7387 = ~1'b0 ;
  assign y7388 = ~n14073 ;
  assign y7389 = ~n14075 ;
  assign y7390 = ~1'b0 ;
  assign y7391 = ~1'b0 ;
  assign y7392 = ~n14078 ;
  assign y7393 = ~n11353 ;
  assign y7394 = ~n14081 ;
  assign y7395 = n14083 ;
  assign y7396 = n14086 ;
  assign y7397 = n14088 ;
  assign y7398 = 1'b0 ;
  assign y7399 = ~n14089 ;
  assign y7400 = ~n14093 ;
  assign y7401 = ~n14095 ;
  assign y7402 = ~n14104 ;
  assign y7403 = ~n14108 ;
  assign y7404 = ~1'b0 ;
  assign y7405 = n14111 ;
  assign y7406 = n14114 ;
  assign y7407 = ~n14115 ;
  assign y7408 = n14116 ;
  assign y7409 = ~1'b0 ;
  assign y7410 = ~n14117 ;
  assign y7411 = n14121 ;
  assign y7412 = ~1'b0 ;
  assign y7413 = ~1'b0 ;
  assign y7414 = ~n14122 ;
  assign y7415 = n5396 ;
  assign y7416 = ~n14124 ;
  assign y7417 = ~n14125 ;
  assign y7418 = ~n14126 ;
  assign y7419 = ~1'b0 ;
  assign y7420 = ~1'b0 ;
  assign y7421 = ~1'b0 ;
  assign y7422 = ~1'b0 ;
  assign y7423 = ~n14127 ;
  assign y7424 = ~n14129 ;
  assign y7425 = ~n14132 ;
  assign y7426 = ~n14134 ;
  assign y7427 = ~n9377 ;
  assign y7428 = ~n14135 ;
  assign y7429 = ~n14136 ;
  assign y7430 = ~1'b0 ;
  assign y7431 = ~1'b0 ;
  assign y7432 = ~n14137 ;
  assign y7433 = n14142 ;
  assign y7434 = n14145 ;
  assign y7435 = ~n14146 ;
  assign y7436 = ~1'b0 ;
  assign y7437 = n14148 ;
  assign y7438 = ~1'b0 ;
  assign y7439 = ~n14158 ;
  assign y7440 = n14160 ;
  assign y7441 = n14161 ;
  assign y7442 = n13254 ;
  assign y7443 = ~n14165 ;
  assign y7444 = ~n14166 ;
  assign y7445 = n14167 ;
  assign y7446 = ~n14169 ;
  assign y7447 = ~1'b0 ;
  assign y7448 = ~1'b0 ;
  assign y7449 = ~n14170 ;
  assign y7450 = ~1'b0 ;
  assign y7451 = n14173 ;
  assign y7452 = ~n14175 ;
  assign y7453 = n14188 ;
  assign y7454 = ~n2403 ;
  assign y7455 = ~n14196 ;
  assign y7456 = ~n14197 ;
  assign y7457 = n14210 ;
  assign y7458 = ~1'b0 ;
  assign y7459 = ~1'b0 ;
  assign y7460 = n14213 ;
  assign y7461 = ~1'b0 ;
  assign y7462 = ~1'b0 ;
  assign y7463 = ~n14219 ;
  assign y7464 = n14220 ;
  assign y7465 = n14227 ;
  assign y7466 = n4506 ;
  assign y7467 = ~1'b0 ;
  assign y7468 = ~1'b0 ;
  assign y7469 = ~1'b0 ;
  assign y7470 = n2382 ;
  assign y7471 = n1288 ;
  assign y7472 = ~1'b0 ;
  assign y7473 = n14228 ;
  assign y7474 = ~n14229 ;
  assign y7475 = ~n14230 ;
  assign y7476 = 1'b0 ;
  assign y7477 = n14231 ;
  assign y7478 = n14233 ;
  assign y7479 = ~n14236 ;
  assign y7480 = n14237 ;
  assign y7481 = n14242 ;
  assign y7482 = ~n6494 ;
  assign y7483 = ~n14244 ;
  assign y7484 = n14247 ;
  assign y7485 = ~n4808 ;
  assign y7486 = n14249 ;
  assign y7487 = ~n14251 ;
  assign y7488 = ~n14252 ;
  assign y7489 = n14253 ;
  assign y7490 = n14254 ;
  assign y7491 = ~n14255 ;
  assign y7492 = ~1'b0 ;
  assign y7493 = ~n14258 ;
  assign y7494 = ~n14260 ;
  assign y7495 = ~n12860 ;
  assign y7496 = ~n10716 ;
  assign y7497 = ~n14261 ;
  assign y7498 = ~n14262 ;
  assign y7499 = ~n14266 ;
  assign y7500 = ~n11221 ;
  assign y7501 = ~n2635 ;
  assign y7502 = n14274 ;
  assign y7503 = n8124 ;
  assign y7504 = n14276 ;
  assign y7505 = 1'b0 ;
  assign y7506 = ~1'b0 ;
  assign y7507 = ~1'b0 ;
  assign y7508 = ~n14279 ;
  assign y7509 = n291 ;
  assign y7510 = ~1'b0 ;
  assign y7511 = ~1'b0 ;
  assign y7512 = ~n14280 ;
  assign y7513 = ~n14281 ;
  assign y7514 = n14282 ;
  assign y7515 = n14285 ;
  assign y7516 = ~n14286 ;
  assign y7517 = ~n14287 ;
  assign y7518 = ~1'b0 ;
  assign y7519 = ~n14293 ;
  assign y7520 = n14295 ;
  assign y7521 = n14299 ;
  assign y7522 = n14302 ;
  assign y7523 = ~1'b0 ;
  assign y7524 = ~1'b0 ;
  assign y7525 = ~1'b0 ;
  assign y7526 = n14307 ;
  assign y7527 = ~n14311 ;
  assign y7528 = n14312 ;
  assign y7529 = n14317 ;
  assign y7530 = ~n14320 ;
  assign y7531 = n14322 ;
  assign y7532 = ~1'b0 ;
  assign y7533 = ~n3132 ;
  assign y7534 = ~n14327 ;
  assign y7535 = n14329 ;
  assign y7536 = n9852 ;
  assign y7537 = ~n14330 ;
  assign y7538 = n14333 ;
  assign y7539 = ~1'b0 ;
  assign y7540 = ~n14334 ;
  assign y7541 = ~n14335 ;
  assign y7542 = n14338 ;
  assign y7543 = ~1'b0 ;
  assign y7544 = n14340 ;
  assign y7545 = 1'b0 ;
  assign y7546 = ~n14342 ;
  assign y7547 = n14344 ;
  assign y7548 = ~1'b0 ;
  assign y7549 = n14347 ;
  assign y7550 = ~1'b0 ;
  assign y7551 = ~n14350 ;
  assign y7552 = ~n14352 ;
  assign y7553 = n14354 ;
  assign y7554 = n14360 ;
  assign y7555 = ~n14362 ;
  assign y7556 = n14366 ;
  assign y7557 = n14368 ;
  assign y7558 = n14372 ;
  assign y7559 = ~n3985 ;
  assign y7560 = ~1'b0 ;
  assign y7561 = ~1'b0 ;
  assign y7562 = ~n14373 ;
  assign y7563 = n14374 ;
  assign y7564 = n14379 ;
  assign y7565 = ~1'b0 ;
  assign y7566 = ~1'b0 ;
  assign y7567 = n14382 ;
  assign y7568 = n14384 ;
  assign y7569 = ~1'b0 ;
  assign y7570 = ~1'b0 ;
  assign y7571 = ~1'b0 ;
  assign y7572 = n14386 ;
  assign y7573 = ~n14387 ;
  assign y7574 = n14389 ;
  assign y7575 = ~1'b0 ;
  assign y7576 = ~n14390 ;
  assign y7577 = n12008 ;
  assign y7578 = ~1'b0 ;
  assign y7579 = ~1'b0 ;
  assign y7580 = ~1'b0 ;
  assign y7581 = ~n14392 ;
  assign y7582 = ~n14394 ;
  assign y7583 = ~1'b0 ;
  assign y7584 = n14396 ;
  assign y7585 = ~n14398 ;
  assign y7586 = n14402 ;
  assign y7587 = ~1'b0 ;
  assign y7588 = 1'b0 ;
  assign y7589 = n14403 ;
  assign y7590 = ~n2129 ;
  assign y7591 = n14404 ;
  assign y7592 = n14405 ;
  assign y7593 = ~1'b0 ;
  assign y7594 = ~1'b0 ;
  assign y7595 = ~n14410 ;
  assign y7596 = n14412 ;
  assign y7597 = n11676 ;
  assign y7598 = n14416 ;
  assign y7599 = ~1'b0 ;
  assign y7600 = ~1'b0 ;
  assign y7601 = ~n14417 ;
  assign y7602 = ~1'b0 ;
  assign y7603 = n14420 ;
  assign y7604 = ~n14422 ;
  assign y7605 = n14433 ;
  assign y7606 = ~1'b0 ;
  assign y7607 = ~n14435 ;
  assign y7608 = ~1'b0 ;
  assign y7609 = ~n14438 ;
  assign y7610 = ~1'b0 ;
  assign y7611 = n14441 ;
  assign y7612 = ~n14442 ;
  assign y7613 = ~n14444 ;
  assign y7614 = n14448 ;
  assign y7615 = n14450 ;
  assign y7616 = ~n14451 ;
  assign y7617 = ~n14458 ;
  assign y7618 = ~n14459 ;
  assign y7619 = n14460 ;
  assign y7620 = ~n14464 ;
  assign y7621 = ~1'b0 ;
  assign y7622 = n14465 ;
  assign y7623 = ~1'b0 ;
  assign y7624 = ~1'b0 ;
  assign y7625 = n14469 ;
  assign y7626 = n2101 ;
  assign y7627 = n14473 ;
  assign y7628 = ~1'b0 ;
  assign y7629 = ~1'b0 ;
  assign y7630 = n14475 ;
  assign y7631 = n14480 ;
  assign y7632 = n14484 ;
  assign y7633 = ~n14485 ;
  assign y7634 = ~n14486 ;
  assign y7635 = ~1'b0 ;
  assign y7636 = ~1'b0 ;
  assign y7637 = ~n14491 ;
  assign y7638 = 1'b0 ;
  assign y7639 = n14493 ;
  assign y7640 = ~1'b0 ;
  assign y7641 = n3166 ;
  assign y7642 = n14495 ;
  assign y7643 = ~1'b0 ;
  assign y7644 = n14498 ;
  assign y7645 = ~n14500 ;
  assign y7646 = n14502 ;
  assign y7647 = ~n14507 ;
  assign y7648 = ~n14511 ;
  assign y7649 = ~n14514 ;
  assign y7650 = ~1'b0 ;
  assign y7651 = 1'b0 ;
  assign y7652 = n14519 ;
  assign y7653 = ~n14525 ;
  assign y7654 = n14527 ;
  assign y7655 = ~n14529 ;
  assign y7656 = ~n14532 ;
  assign y7657 = ~1'b0 ;
  assign y7658 = ~1'b0 ;
  assign y7659 = ~1'b0 ;
  assign y7660 = ~n14536 ;
  assign y7661 = ~n14537 ;
  assign y7662 = ~n14538 ;
  assign y7663 = n14540 ;
  assign y7664 = ~1'b0 ;
  assign y7665 = ~n14542 ;
  assign y7666 = n7494 ;
  assign y7667 = n14543 ;
  assign y7668 = n14546 ;
  assign y7669 = ~1'b0 ;
  assign y7670 = ~n14550 ;
  assign y7671 = n14552 ;
  assign y7672 = ~n14556 ;
  assign y7673 = ~1'b0 ;
  assign y7674 = n14559 ;
  assign y7675 = ~n14560 ;
  assign y7676 = n14561 ;
  assign y7677 = ~n14568 ;
  assign y7678 = n3633 ;
  assign y7679 = ~1'b0 ;
  assign y7680 = ~1'b0 ;
  assign y7681 = n14578 ;
  assign y7682 = ~n14579 ;
  assign y7683 = ~1'b0 ;
  assign y7684 = ~1'b0 ;
  assign y7685 = ~n14580 ;
  assign y7686 = ~1'b0 ;
  assign y7687 = ~n14582 ;
  assign y7688 = ~n14593 ;
  assign y7689 = n14595 ;
  assign y7690 = n2923 ;
  assign y7691 = ~n14596 ;
  assign y7692 = ~n14597 ;
  assign y7693 = n14600 ;
  assign y7694 = ~n14601 ;
  assign y7695 = n14603 ;
  assign y7696 = ~n14607 ;
  assign y7697 = n14608 ;
  assign y7698 = ~1'b0 ;
  assign y7699 = n14611 ;
  assign y7700 = n14612 ;
  assign y7701 = n14613 ;
  assign y7702 = n14614 ;
  assign y7703 = n14616 ;
  assign y7704 = ~1'b0 ;
  assign y7705 = ~n14620 ;
  assign y7706 = n14624 ;
  assign y7707 = ~n14634 ;
  assign y7708 = ~n14636 ;
  assign y7709 = n14644 ;
  assign y7710 = n14648 ;
  assign y7711 = ~n14649 ;
  assign y7712 = n14652 ;
  assign y7713 = n14653 ;
  assign y7714 = ~n14250 ;
  assign y7715 = n14657 ;
  assign y7716 = n14662 ;
  assign y7717 = n14665 ;
  assign y7718 = n14670 ;
  assign y7719 = n14674 ;
  assign y7720 = n14675 ;
  assign y7721 = ~1'b0 ;
  assign y7722 = ~n14676 ;
  assign y7723 = n14679 ;
  assign y7724 = n14684 ;
  assign y7725 = ~1'b0 ;
  assign y7726 = ~n14685 ;
  assign y7727 = ~1'b0 ;
  assign y7728 = ~1'b0 ;
  assign y7729 = ~n14686 ;
  assign y7730 = ~n14689 ;
  assign y7731 = n14693 ;
  assign y7732 = n14696 ;
  assign y7733 = ~1'b0 ;
  assign y7734 = ~n14697 ;
  assign y7735 = ~n8342 ;
  assign y7736 = ~n14706 ;
  assign y7737 = ~n14708 ;
  assign y7738 = ~n3637 ;
  assign y7739 = ~n14720 ;
  assign y7740 = ~1'b0 ;
  assign y7741 = ~n14722 ;
  assign y7742 = ~n14724 ;
  assign y7743 = ~1'b0 ;
  assign y7744 = n14730 ;
  assign y7745 = ~n14731 ;
  assign y7746 = ~1'b0 ;
  assign y7747 = ~1'b0 ;
  assign y7748 = ~n14735 ;
  assign y7749 = ~n14739 ;
  assign y7750 = ~n14740 ;
  assign y7751 = ~n14741 ;
  assign y7752 = ~1'b0 ;
  assign y7753 = ~n14746 ;
  assign y7754 = n14748 ;
  assign y7755 = ~n14753 ;
  assign y7756 = n14754 ;
  assign y7757 = ~1'b0 ;
  assign y7758 = n14760 ;
  assign y7759 = n14761 ;
  assign y7760 = 1'b0 ;
  assign y7761 = ~n14763 ;
  assign y7762 = n14765 ;
  assign y7763 = n11666 ;
  assign y7764 = ~1'b0 ;
  assign y7765 = n14770 ;
  assign y7766 = 1'b0 ;
  assign y7767 = ~n14772 ;
  assign y7768 = ~1'b0 ;
  assign y7769 = ~n14774 ;
  assign y7770 = ~n14776 ;
  assign y7771 = n14782 ;
  assign y7772 = n14790 ;
  assign y7773 = ~n14791 ;
  assign y7774 = ~1'b0 ;
  assign y7775 = ~1'b0 ;
  assign y7776 = n14792 ;
  assign y7777 = ~n14795 ;
  assign y7778 = n14796 ;
  assign y7779 = ~1'b0 ;
  assign y7780 = n14804 ;
  assign y7781 = n14805 ;
  assign y7782 = ~n14808 ;
  assign y7783 = ~n14810 ;
  assign y7784 = n14812 ;
  assign y7785 = ~1'b0 ;
  assign y7786 = ~n14815 ;
  assign y7787 = ~n14817 ;
  assign y7788 = ~n14818 ;
  assign y7789 = ~n14819 ;
  assign y7790 = n14824 ;
  assign y7791 = n14825 ;
  assign y7792 = n11360 ;
  assign y7793 = ~1'b0 ;
  assign y7794 = n14827 ;
  assign y7795 = n14829 ;
  assign y7796 = ~n14832 ;
  assign y7797 = n623 ;
  assign y7798 = ~1'b0 ;
  assign y7799 = ~n13205 ;
  assign y7800 = ~n3761 ;
  assign y7801 = ~n14837 ;
  assign y7802 = ~n14839 ;
  assign y7803 = n14842 ;
  assign y7804 = n14845 ;
  assign y7805 = n14846 ;
  assign y7806 = ~1'b0 ;
  assign y7807 = n14853 ;
  assign y7808 = ~1'b0 ;
  assign y7809 = n14856 ;
  assign y7810 = ~n14857 ;
  assign y7811 = ~1'b0 ;
  assign y7812 = n14867 ;
  assign y7813 = 1'b0 ;
  assign y7814 = n4213 ;
  assign y7815 = n4433 ;
  assign y7816 = n14870 ;
  assign y7817 = n14872 ;
  assign y7818 = ~1'b0 ;
  assign y7819 = ~n5221 ;
  assign y7820 = ~n14873 ;
  assign y7821 = ~n14877 ;
  assign y7822 = ~1'b0 ;
  assign y7823 = ~1'b0 ;
  assign y7824 = ~1'b0 ;
  assign y7825 = ~n14880 ;
  assign y7826 = n14885 ;
  assign y7827 = n14889 ;
  assign y7828 = n14890 ;
  assign y7829 = ~1'b0 ;
  assign y7830 = n7609 ;
  assign y7831 = n14891 ;
  assign y7832 = ~n14899 ;
  assign y7833 = ~n14902 ;
  assign y7834 = ~n14904 ;
  assign y7835 = ~1'b0 ;
  assign y7836 = ~n10391 ;
  assign y7837 = n14907 ;
  assign y7838 = ~1'b0 ;
  assign y7839 = ~1'b0 ;
  assign y7840 = n3676 ;
  assign y7841 = ~1'b0 ;
  assign y7842 = ~1'b0 ;
  assign y7843 = ~1'b0 ;
  assign y7844 = ~n14910 ;
  assign y7845 = ~n801 ;
  assign y7846 = ~1'b0 ;
  assign y7847 = ~1'b0 ;
  assign y7848 = ~n9419 ;
  assign y7849 = 1'b0 ;
  assign y7850 = n14915 ;
  assign y7851 = 1'b0 ;
  assign y7852 = ~n14916 ;
  assign y7853 = n428 ;
  assign y7854 = ~n14918 ;
  assign y7855 = n14920 ;
  assign y7856 = ~n14922 ;
  assign y7857 = ~n14923 ;
  assign y7858 = n6749 ;
  assign y7859 = n2478 ;
  assign y7860 = n14925 ;
  assign y7861 = ~n14926 ;
  assign y7862 = n14927 ;
  assign y7863 = ~n14928 ;
  assign y7864 = 1'b0 ;
  assign y7865 = ~n14930 ;
  assign y7866 = n14931 ;
  assign y7867 = n14932 ;
  assign y7868 = n9151 ;
  assign y7869 = n7182 ;
  assign y7870 = ~1'b0 ;
  assign y7871 = ~n14933 ;
  assign y7872 = ~n14934 ;
  assign y7873 = n14941 ;
  assign y7874 = n14944 ;
  assign y7875 = ~1'b0 ;
  assign y7876 = n14947 ;
  assign y7877 = n14950 ;
  assign y7878 = ~n14952 ;
  assign y7879 = ~1'b0 ;
  assign y7880 = 1'b0 ;
  assign y7881 = 1'b0 ;
  assign y7882 = ~n14953 ;
  assign y7883 = n7405 ;
  assign y7884 = n14954 ;
  assign y7885 = ~1'b0 ;
  assign y7886 = ~n14955 ;
  assign y7887 = ~1'b0 ;
  assign y7888 = ~n14957 ;
  assign y7889 = n14958 ;
  assign y7890 = n14959 ;
  assign y7891 = ~n14961 ;
  assign y7892 = ~n14969 ;
  assign y7893 = ~n14973 ;
  assign y7894 = n14976 ;
  assign y7895 = 1'b0 ;
  assign y7896 = n14979 ;
  assign y7897 = ~n14985 ;
  assign y7898 = 1'b0 ;
  assign y7899 = ~1'b0 ;
  assign y7900 = ~n14989 ;
  assign y7901 = ~1'b0 ;
  assign y7902 = n14991 ;
  assign y7903 = n7390 ;
  assign y7904 = 1'b0 ;
  assign y7905 = ~1'b0 ;
  assign y7906 = ~n14994 ;
  assign y7907 = n14997 ;
  assign y7908 = n14999 ;
  assign y7909 = ~n12860 ;
  assign y7910 = ~n15001 ;
  assign y7911 = n15002 ;
  assign y7912 = ~n4883 ;
  assign y7913 = ~1'b0 ;
  assign y7914 = ~n15003 ;
  assign y7915 = ~1'b0 ;
  assign y7916 = n15005 ;
  assign y7917 = ~n15008 ;
  assign y7918 = n15009 ;
  assign y7919 = n15013 ;
  assign y7920 = ~1'b0 ;
  assign y7921 = ~n15015 ;
  assign y7922 = ~n15016 ;
  assign y7923 = n15019 ;
  assign y7924 = ~1'b0 ;
  assign y7925 = ~1'b0 ;
  assign y7926 = n15020 ;
  assign y7927 = ~n15022 ;
  assign y7928 = ~1'b0 ;
  assign y7929 = ~n15025 ;
  assign y7930 = n15027 ;
  assign y7931 = ~n15029 ;
  assign y7932 = n15030 ;
  assign y7933 = n15031 ;
  assign y7934 = ~1'b0 ;
  assign y7935 = ~1'b0 ;
  assign y7936 = ~n15032 ;
  assign y7937 = n15038 ;
  assign y7938 = ~1'b0 ;
  assign y7939 = ~1'b0 ;
  assign y7940 = ~n15043 ;
  assign y7941 = ~1'b0 ;
  assign y7942 = ~n15048 ;
  assign y7943 = n15050 ;
  assign y7944 = n15052 ;
  assign y7945 = ~1'b0 ;
  assign y7946 = n15053 ;
  assign y7947 = n15054 ;
  assign y7948 = n15055 ;
  assign y7949 = ~1'b0 ;
  assign y7950 = n15056 ;
  assign y7951 = ~n15064 ;
  assign y7952 = ~n15070 ;
  assign y7953 = ~n15071 ;
  assign y7954 = ~n15075 ;
  assign y7955 = n15078 ;
  assign y7956 = ~n15081 ;
  assign y7957 = n11312 ;
  assign y7958 = ~1'b0 ;
  assign y7959 = n6271 ;
  assign y7960 = ~1'b0 ;
  assign y7961 = ~1'b0 ;
  assign y7962 = n15084 ;
  assign y7963 = n15086 ;
  assign y7964 = ~1'b0 ;
  assign y7965 = n15087 ;
  assign y7966 = n15090 ;
  assign y7967 = ~n15092 ;
  assign y7968 = n15098 ;
  assign y7969 = n5796 ;
  assign y7970 = ~n15099 ;
  assign y7971 = ~1'b0 ;
  assign y7972 = ~n15105 ;
  assign y7973 = n7027 ;
  assign y7974 = n15106 ;
  assign y7975 = n15108 ;
  assign y7976 = ~1'b0 ;
  assign y7977 = n15112 ;
  assign y7978 = n15115 ;
  assign y7979 = ~n15117 ;
  assign y7980 = n15123 ;
  assign y7981 = ~n15126 ;
  assign y7982 = ~n15127 ;
  assign y7983 = 1'b0 ;
  assign y7984 = ~1'b0 ;
  assign y7985 = n15129 ;
  assign y7986 = ~1'b0 ;
  assign y7987 = ~n15132 ;
  assign y7988 = ~1'b0 ;
  assign y7989 = ~n15133 ;
  assign y7990 = ~n15136 ;
  assign y7991 = n15145 ;
  assign y7992 = ~n15150 ;
  assign y7993 = ~n15157 ;
  assign y7994 = ~n15159 ;
  assign y7995 = n6170 ;
  assign y7996 = ~n15164 ;
  assign y7997 = ~n15168 ;
  assign y7998 = n15170 ;
  assign y7999 = n15174 ;
  assign y8000 = ~1'b0 ;
  assign y8001 = n15178 ;
  assign y8002 = ~1'b0 ;
  assign y8003 = ~n15180 ;
  assign y8004 = ~n15183 ;
  assign y8005 = n15187 ;
  assign y8006 = ~n15188 ;
  assign y8007 = n15189 ;
  assign y8008 = ~1'b0 ;
  assign y8009 = ~1'b0 ;
  assign y8010 = ~n15190 ;
  assign y8011 = n15191 ;
  assign y8012 = ~1'b0 ;
  assign y8013 = ~1'b0 ;
  assign y8014 = n15192 ;
  assign y8015 = ~n15193 ;
  assign y8016 = n15195 ;
  assign y8017 = n15200 ;
  assign y8018 = ~n15206 ;
  assign y8019 = ~n15209 ;
  assign y8020 = ~n15210 ;
  assign y8021 = n15214 ;
  assign y8022 = ~1'b0 ;
  assign y8023 = ~n15218 ;
  assign y8024 = ~1'b0 ;
  assign y8025 = n15220 ;
  assign y8026 = ~1'b0 ;
  assign y8027 = n15221 ;
  assign y8028 = n15222 ;
  assign y8029 = ~1'b0 ;
  assign y8030 = ~1'b0 ;
  assign y8031 = n15226 ;
  assign y8032 = n15228 ;
  assign y8033 = ~n15230 ;
  assign y8034 = ~n15235 ;
  assign y8035 = ~n15238 ;
  assign y8036 = n15240 ;
  assign y8037 = n15244 ;
  assign y8038 = n15246 ;
  assign y8039 = ~1'b0 ;
  assign y8040 = 1'b0 ;
  assign y8041 = n15250 ;
  assign y8042 = ~n15253 ;
  assign y8043 = n15256 ;
  assign y8044 = n15257 ;
  assign y8045 = 1'b0 ;
  assign y8046 = ~1'b0 ;
  assign y8047 = n15259 ;
  assign y8048 = ~n6937 ;
  assign y8049 = ~n15260 ;
  assign y8050 = n2486 ;
  assign y8051 = n8299 ;
  assign y8052 = ~1'b0 ;
  assign y8053 = ~n15261 ;
  assign y8054 = 1'b0 ;
  assign y8055 = n15262 ;
  assign y8056 = ~n15263 ;
  assign y8057 = ~n15265 ;
  assign y8058 = n15267 ;
  assign y8059 = ~1'b0 ;
  assign y8060 = n15268 ;
  assign y8061 = n15270 ;
  assign y8062 = n15271 ;
  assign y8063 = ~n3724 ;
  assign y8064 = ~1'b0 ;
  assign y8065 = ~1'b0 ;
  assign y8066 = ~1'b0 ;
  assign y8067 = ~n15274 ;
  assign y8068 = ~1'b0 ;
  assign y8069 = ~n15275 ;
  assign y8070 = n15278 ;
  assign y8071 = n11242 ;
  assign y8072 = ~n15281 ;
  assign y8073 = ~n15287 ;
  assign y8074 = ~1'b0 ;
  assign y8075 = n12395 ;
  assign y8076 = ~n15290 ;
  assign y8077 = ~n7836 ;
  assign y8078 = ~n15291 ;
  assign y8079 = ~n15298 ;
  assign y8080 = ~n15299 ;
  assign y8081 = ~n15300 ;
  assign y8082 = n15307 ;
  assign y8083 = ~n15310 ;
  assign y8084 = n15313 ;
  assign y8085 = ~n15316 ;
  assign y8086 = ~1'b0 ;
  assign y8087 = n15318 ;
  assign y8088 = ~n15321 ;
  assign y8089 = ~1'b0 ;
  assign y8090 = n15322 ;
  assign y8091 = n15326 ;
  assign y8092 = ~1'b0 ;
  assign y8093 = ~n11102 ;
  assign y8094 = n15328 ;
  assign y8095 = n15331 ;
  assign y8096 = ~n15336 ;
  assign y8097 = ~1'b0 ;
  assign y8098 = ~n15337 ;
  assign y8099 = ~1'b0 ;
  assign y8100 = ~n15338 ;
  assign y8101 = ~n15339 ;
  assign y8102 = n15341 ;
  assign y8103 = ~1'b0 ;
  assign y8104 = ~1'b0 ;
  assign y8105 = n3842 ;
  assign y8106 = n15342 ;
  assign y8107 = ~n15344 ;
  assign y8108 = ~n15347 ;
  assign y8109 = ~1'b0 ;
  assign y8110 = ~1'b0 ;
  assign y8111 = ~1'b0 ;
  assign y8112 = ~1'b0 ;
  assign y8113 = ~1'b0 ;
  assign y8114 = ~1'b0 ;
  assign y8115 = ~1'b0 ;
  assign y8116 = n15352 ;
  assign y8117 = ~n15354 ;
  assign y8118 = 1'b0 ;
  assign y8119 = n15356 ;
  assign y8120 = ~1'b0 ;
  assign y8121 = ~n15364 ;
  assign y8122 = ~n15365 ;
  assign y8123 = ~n13200 ;
  assign y8124 = ~n15371 ;
  assign y8125 = ~n15374 ;
  assign y8126 = 1'b0 ;
  assign y8127 = ~n15377 ;
  assign y8128 = ~1'b0 ;
  assign y8129 = ~1'b0 ;
  assign y8130 = ~n15387 ;
  assign y8131 = ~n15392 ;
  assign y8132 = ~n13566 ;
  assign y8133 = ~1'b0 ;
  assign y8134 = ~1'b0 ;
  assign y8135 = ~1'b0 ;
  assign y8136 = ~1'b0 ;
  assign y8137 = ~1'b0 ;
  assign y8138 = ~1'b0 ;
  assign y8139 = ~1'b0 ;
  assign y8140 = n15393 ;
  assign y8141 = ~n15396 ;
  assign y8142 = ~1'b0 ;
  assign y8143 = ~1'b0 ;
  assign y8144 = ~1'b0 ;
  assign y8145 = n15399 ;
  assign y8146 = ~n15401 ;
  assign y8147 = ~n15403 ;
  assign y8148 = ~1'b0 ;
  assign y8149 = n15404 ;
  assign y8150 = ~n15407 ;
  assign y8151 = ~n15409 ;
  assign y8152 = ~n7808 ;
  assign y8153 = 1'b0 ;
  assign y8154 = ~n13142 ;
  assign y8155 = ~n15411 ;
  assign y8156 = n15412 ;
  assign y8157 = ~1'b0 ;
  assign y8158 = ~n15417 ;
  assign y8159 = ~n15420 ;
  assign y8160 = n15424 ;
  assign y8161 = n15427 ;
  assign y8162 = ~n15429 ;
  assign y8163 = n15433 ;
  assign y8164 = n15435 ;
  assign y8165 = n11550 ;
  assign y8166 = n15436 ;
  assign y8167 = n15437 ;
  assign y8168 = ~n15438 ;
  assign y8169 = ~n15443 ;
  assign y8170 = ~n15444 ;
  assign y8171 = ~1'b0 ;
  assign y8172 = ~n15447 ;
  assign y8173 = ~1'b0 ;
  assign y8174 = n15448 ;
  assign y8175 = ~n15451 ;
  assign y8176 = n15455 ;
  assign y8177 = n15462 ;
  assign y8178 = ~n15465 ;
  assign y8179 = ~1'b0 ;
  assign y8180 = n15468 ;
  assign y8181 = n15471 ;
  assign y8182 = n15473 ;
  assign y8183 = ~1'b0 ;
  assign y8184 = n15479 ;
  assign y8185 = n15481 ;
  assign y8186 = ~1'b0 ;
  assign y8187 = n15483 ;
  assign y8188 = ~1'b0 ;
  assign y8189 = ~1'b0 ;
  assign y8190 = ~n15484 ;
  assign y8191 = n6274 ;
  assign y8192 = ~1'b0 ;
  assign y8193 = n15485 ;
  assign y8194 = n15488 ;
  assign y8195 = n15489 ;
  assign y8196 = ~n15493 ;
  assign y8197 = ~1'b0 ;
  assign y8198 = ~n15495 ;
  assign y8199 = ~1'b0 ;
  assign y8200 = ~n15497 ;
  assign y8201 = n15499 ;
  assign y8202 = ~n15501 ;
  assign y8203 = n15502 ;
  assign y8204 = n11535 ;
  assign y8205 = ~n15506 ;
  assign y8206 = ~1'b0 ;
  assign y8207 = ~n15507 ;
  assign y8208 = n15508 ;
  assign y8209 = ~n15509 ;
  assign y8210 = ~1'b0 ;
  assign y8211 = ~n15512 ;
  assign y8212 = n15513 ;
  assign y8213 = n4044 ;
  assign y8214 = 1'b0 ;
  assign y8215 = ~n11037 ;
  assign y8216 = ~1'b0 ;
  assign y8217 = ~n15515 ;
  assign y8218 = ~1'b0 ;
  assign y8219 = n15520 ;
  assign y8220 = ~1'b0 ;
  assign y8221 = ~n15404 ;
  assign y8222 = n15521 ;
  assign y8223 = n15522 ;
  assign y8224 = ~1'b0 ;
  assign y8225 = n13896 ;
  assign y8226 = n15524 ;
  assign y8227 = n15525 ;
  assign y8228 = ~n15526 ;
  assign y8229 = ~n15533 ;
  assign y8230 = ~n15539 ;
  assign y8231 = n15544 ;
  assign y8232 = n15545 ;
  assign y8233 = n14642 ;
  assign y8234 = ~n15547 ;
  assign y8235 = ~n15548 ;
  assign y8236 = ~1'b0 ;
  assign y8237 = n15550 ;
  assign y8238 = ~1'b0 ;
  assign y8239 = ~n15557 ;
  assign y8240 = ~1'b0 ;
  assign y8241 = ~1'b0 ;
  assign y8242 = n15558 ;
  assign y8243 = ~1'b0 ;
  assign y8244 = ~1'b0 ;
  assign y8245 = 1'b0 ;
  assign y8246 = ~1'b0 ;
  assign y8247 = n15562 ;
  assign y8248 = n15567 ;
  assign y8249 = ~n15571 ;
  assign y8250 = ~1'b0 ;
  assign y8251 = ~n15575 ;
  assign y8252 = 1'b0 ;
  assign y8253 = ~1'b0 ;
  assign y8254 = ~n15584 ;
  assign y8255 = n12533 ;
  assign y8256 = ~n15585 ;
  assign y8257 = n15586 ;
  assign y8258 = ~1'b0 ;
  assign y8259 = ~1'b0 ;
  assign y8260 = n15588 ;
  assign y8261 = ~n15594 ;
  assign y8262 = n15598 ;
  assign y8263 = ~n15599 ;
  assign y8264 = ~n15603 ;
  assign y8265 = ~n15606 ;
  assign y8266 = ~n15609 ;
  assign y8267 = ~n911 ;
  assign y8268 = ~1'b0 ;
  assign y8269 = ~n15611 ;
  assign y8270 = ~n15614 ;
  assign y8271 = ~1'b0 ;
  assign y8272 = ~n15616 ;
  assign y8273 = ~n2905 ;
  assign y8274 = n15617 ;
  assign y8275 = ~1'b0 ;
  assign y8276 = ~n15618 ;
  assign y8277 = ~1'b0 ;
  assign y8278 = ~1'b0 ;
  assign y8279 = ~n15619 ;
  assign y8280 = n15620 ;
  assign y8281 = ~1'b0 ;
  assign y8282 = ~n15622 ;
  assign y8283 = n15623 ;
  assign y8284 = n15636 ;
  assign y8285 = ~1'b0 ;
  assign y8286 = n15230 ;
  assign y8287 = ~n11701 ;
  assign y8288 = ~1'b0 ;
  assign y8289 = n15638 ;
  assign y8290 = ~n15639 ;
  assign y8291 = ~n15644 ;
  assign y8292 = ~n15646 ;
  assign y8293 = n6871 ;
  assign y8294 = ~n15648 ;
  assign y8295 = ~1'b0 ;
  assign y8296 = n15649 ;
  assign y8297 = n15659 ;
  assign y8298 = n15661 ;
  assign y8299 = ~n15662 ;
  assign y8300 = n15664 ;
  assign y8301 = ~1'b0 ;
  assign y8302 = 1'b0 ;
  assign y8303 = ~n15665 ;
  assign y8304 = n15674 ;
  assign y8305 = n15681 ;
  assign y8306 = n15687 ;
  assign y8307 = ~1'b0 ;
  assign y8308 = ~1'b0 ;
  assign y8309 = ~n15689 ;
  assign y8310 = n15690 ;
  assign y8311 = ~1'b0 ;
  assign y8312 = ~n13424 ;
  assign y8313 = ~1'b0 ;
  assign y8314 = ~1'b0 ;
  assign y8315 = 1'b0 ;
  assign y8316 = ~n15698 ;
  assign y8317 = ~1'b0 ;
  assign y8318 = ~1'b0 ;
  assign y8319 = 1'b0 ;
  assign y8320 = n15700 ;
  assign y8321 = ~n15702 ;
  assign y8322 = ~1'b0 ;
  assign y8323 = ~n15703 ;
  assign y8324 = ~1'b0 ;
  assign y8325 = ~1'b0 ;
  assign y8326 = ~n15705 ;
  assign y8327 = ~n15708 ;
  assign y8328 = ~n15710 ;
  assign y8329 = n15712 ;
  assign y8330 = n15715 ;
  assign y8331 = n15716 ;
  assign y8332 = ~1'b0 ;
  assign y8333 = ~1'b0 ;
  assign y8334 = ~1'b0 ;
  assign y8335 = ~1'b0 ;
  assign y8336 = ~1'b0 ;
  assign y8337 = ~n15718 ;
  assign y8338 = n15719 ;
  assign y8339 = ~1'b0 ;
  assign y8340 = ~1'b0 ;
  assign y8341 = n15723 ;
  assign y8342 = ~1'b0 ;
  assign y8343 = n15725 ;
  assign y8344 = n15728 ;
  assign y8345 = ~n15734 ;
  assign y8346 = ~n15424 ;
  assign y8347 = ~n1392 ;
  assign y8348 = ~n15736 ;
  assign y8349 = n15737 ;
  assign y8350 = n15742 ;
  assign y8351 = ~n15745 ;
  assign y8352 = ~1'b0 ;
  assign y8353 = ~n4937 ;
  assign y8354 = ~n15750 ;
  assign y8355 = ~n15756 ;
  assign y8356 = ~1'b0 ;
  assign y8357 = ~n15759 ;
  assign y8358 = n15760 ;
  assign y8359 = ~n15761 ;
  assign y8360 = ~1'b0 ;
  assign y8361 = ~1'b0 ;
  assign y8362 = ~1'b0 ;
  assign y8363 = ~1'b0 ;
  assign y8364 = n15765 ;
  assign y8365 = ~1'b0 ;
  assign y8366 = n15771 ;
  assign y8367 = ~1'b0 ;
  assign y8368 = ~1'b0 ;
  assign y8369 = ~1'b0 ;
  assign y8370 = n15775 ;
  assign y8371 = ~n15784 ;
  assign y8372 = ~n15788 ;
  assign y8373 = n15789 ;
  assign y8374 = n15790 ;
  assign y8375 = 1'b0 ;
  assign y8376 = n15795 ;
  assign y8377 = ~1'b0 ;
  assign y8378 = ~1'b0 ;
  assign y8379 = ~n15799 ;
  assign y8380 = ~n15801 ;
  assign y8381 = ~1'b0 ;
  assign y8382 = ~1'b0 ;
  assign y8383 = ~n15809 ;
  assign y8384 = ~1'b0 ;
  assign y8385 = n10855 ;
  assign y8386 = ~n15813 ;
  assign y8387 = ~1'b0 ;
  assign y8388 = ~n15815 ;
  assign y8389 = ~n15822 ;
  assign y8390 = n15831 ;
  assign y8391 = ~1'b0 ;
  assign y8392 = ~1'b0 ;
  assign y8393 = n15833 ;
  assign y8394 = n15834 ;
  assign y8395 = ~n15836 ;
  assign y8396 = n10595 ;
  assign y8397 = n15844 ;
  assign y8398 = ~n15845 ;
  assign y8399 = n15847 ;
  assign y8400 = n15863 ;
  assign y8401 = n15865 ;
  assign y8402 = ~n15867 ;
  assign y8403 = ~1'b0 ;
  assign y8404 = n15869 ;
  assign y8405 = ~n15870 ;
  assign y8406 = ~n15873 ;
  assign y8407 = n15874 ;
  assign y8408 = ~1'b0 ;
  assign y8409 = ~n15879 ;
  assign y8410 = ~1'b0 ;
  assign y8411 = ~n7062 ;
  assign y8412 = n15881 ;
  assign y8413 = n15882 ;
  assign y8414 = ~n15883 ;
  assign y8415 = ~1'b0 ;
  assign y8416 = n15887 ;
  assign y8417 = ~n666 ;
  assign y8418 = ~n15888 ;
  assign y8419 = ~n15889 ;
  assign y8420 = ~n15890 ;
  assign y8421 = ~1'b0 ;
  assign y8422 = ~1'b0 ;
  assign y8423 = ~1'b0 ;
  assign y8424 = n15892 ;
  assign y8425 = n15893 ;
  assign y8426 = ~n15900 ;
  assign y8427 = ~n15902 ;
  assign y8428 = ~n15905 ;
  assign y8429 = 1'b0 ;
  assign y8430 = ~1'b0 ;
  assign y8431 = n15909 ;
  assign y8432 = ~n15916 ;
  assign y8433 = ~n15926 ;
  assign y8434 = n15928 ;
  assign y8435 = ~n15929 ;
  assign y8436 = ~1'b0 ;
  assign y8437 = ~1'b0 ;
  assign y8438 = ~1'b0 ;
  assign y8439 = ~1'b0 ;
  assign y8440 = ~1'b0 ;
  assign y8441 = n15931 ;
  assign y8442 = ~1'b0 ;
  assign y8443 = ~1'b0 ;
  assign y8444 = n15938 ;
  assign y8445 = 1'b0 ;
  assign y8446 = ~1'b0 ;
  assign y8447 = ~n15939 ;
  assign y8448 = ~1'b0 ;
  assign y8449 = ~n15945 ;
  assign y8450 = ~n15948 ;
  assign y8451 = ~n15950 ;
  assign y8452 = n15953 ;
  assign y8453 = ~1'b0 ;
  assign y8454 = n15956 ;
  assign y8455 = n15957 ;
  assign y8456 = ~1'b0 ;
  assign y8457 = ~n15958 ;
  assign y8458 = n15963 ;
  assign y8459 = n15964 ;
  assign y8460 = ~n15974 ;
  assign y8461 = ~1'b0 ;
  assign y8462 = ~n15976 ;
  assign y8463 = ~n15978 ;
  assign y8464 = ~1'b0 ;
  assign y8465 = ~n15990 ;
  assign y8466 = n15992 ;
  assign y8467 = n15997 ;
  assign y8468 = n16000 ;
  assign y8469 = ~n16002 ;
  assign y8470 = n16003 ;
  assign y8471 = ~1'b0 ;
  assign y8472 = n16006 ;
  assign y8473 = ~1'b0 ;
  assign y8474 = ~n16008 ;
  assign y8475 = ~1'b0 ;
  assign y8476 = ~1'b0 ;
  assign y8477 = ~n9943 ;
  assign y8478 = n16010 ;
  assign y8479 = ~1'b0 ;
  assign y8480 = n16012 ;
  assign y8481 = n16017 ;
  assign y8482 = 1'b0 ;
  assign y8483 = n16018 ;
  assign y8484 = ~1'b0 ;
  assign y8485 = ~1'b0 ;
  assign y8486 = n16019 ;
  assign y8487 = ~n16023 ;
  assign y8488 = n16025 ;
  assign y8489 = n7623 ;
  assign y8490 = n16026 ;
  assign y8491 = n16028 ;
  assign y8492 = ~n16030 ;
  assign y8493 = ~n16031 ;
  assign y8494 = n16033 ;
  assign y8495 = n4039 ;
  assign y8496 = ~n16035 ;
  assign y8497 = ~n16039 ;
  assign y8498 = n16040 ;
  assign y8499 = ~n16041 ;
  assign y8500 = ~1'b0 ;
  assign y8501 = ~n16042 ;
  assign y8502 = ~1'b0 ;
  assign y8503 = ~1'b0 ;
  assign y8504 = ~n16044 ;
  assign y8505 = n2565 ;
  assign y8506 = ~n16047 ;
  assign y8507 = ~1'b0 ;
  assign y8508 = ~1'b0 ;
  assign y8509 = n16052 ;
  assign y8510 = ~1'b0 ;
  assign y8511 = n12458 ;
  assign y8512 = n16064 ;
  assign y8513 = n16067 ;
  assign y8514 = n16068 ;
  assign y8515 = n16070 ;
  assign y8516 = 1'b0 ;
  assign y8517 = n16071 ;
  assign y8518 = ~n16073 ;
  assign y8519 = ~1'b0 ;
  assign y8520 = ~1'b0 ;
  assign y8521 = ~1'b0 ;
  assign y8522 = n16077 ;
  assign y8523 = ~n16083 ;
  assign y8524 = n16085 ;
  assign y8525 = n16092 ;
  assign y8526 = ~n16099 ;
  assign y8527 = n16104 ;
  assign y8528 = n10976 ;
  assign y8529 = ~n16106 ;
  assign y8530 = ~1'b0 ;
  assign y8531 = ~n16107 ;
  assign y8532 = ~1'b0 ;
  assign y8533 = ~n16108 ;
  assign y8534 = n16118 ;
  assign y8535 = n16124 ;
  assign y8536 = ~n16126 ;
  assign y8537 = ~n16128 ;
  assign y8538 = ~1'b0 ;
  assign y8539 = n16129 ;
  assign y8540 = n16131 ;
  assign y8541 = n16133 ;
  assign y8542 = n16135 ;
  assign y8543 = n16137 ;
  assign y8544 = ~n16141 ;
  assign y8545 = ~n16142 ;
  assign y8546 = ~n16143 ;
  assign y8547 = n16145 ;
  assign y8548 = ~n16146 ;
  assign y8549 = ~1'b0 ;
  assign y8550 = ~1'b0 ;
  assign y8551 = ~1'b0 ;
  assign y8552 = 1'b0 ;
  assign y8553 = ~n16147 ;
  assign y8554 = n16152 ;
  assign y8555 = n16153 ;
  assign y8556 = ~n16159 ;
  assign y8557 = ~n16160 ;
  assign y8558 = n16163 ;
  assign y8559 = ~1'b0 ;
  assign y8560 = ~n6623 ;
  assign y8561 = n16168 ;
  assign y8562 = ~n16169 ;
  assign y8563 = ~1'b0 ;
  assign y8564 = ~1'b0 ;
  assign y8565 = ~1'b0 ;
  assign y8566 = n16170 ;
  assign y8567 = ~1'b0 ;
  assign y8568 = n16171 ;
  assign y8569 = ~n16172 ;
  assign y8570 = n16173 ;
  assign y8571 = ~1'b0 ;
  assign y8572 = n16175 ;
  assign y8573 = n16176 ;
  assign y8574 = ~1'b0 ;
  assign y8575 = n10137 ;
  assign y8576 = n16177 ;
  assign y8577 = n16179 ;
  assign y8578 = n16180 ;
  assign y8579 = ~n16181 ;
  assign y8580 = ~n16195 ;
  assign y8581 = ~1'b0 ;
  assign y8582 = ~1'b0 ;
  assign y8583 = ~n16199 ;
  assign y8584 = ~1'b0 ;
  assign y8585 = n16202 ;
  assign y8586 = ~n16203 ;
  assign y8587 = ~n16206 ;
  assign y8588 = n4914 ;
  assign y8589 = ~1'b0 ;
  assign y8590 = ~n16207 ;
  assign y8591 = n16209 ;
  assign y8592 = n12408 ;
  assign y8593 = n16213 ;
  assign y8594 = n16215 ;
  assign y8595 = ~n16216 ;
  assign y8596 = n16219 ;
  assign y8597 = ~n16220 ;
  assign y8598 = ~n16224 ;
  assign y8599 = ~n16227 ;
  assign y8600 = ~1'b0 ;
  assign y8601 = ~1'b0 ;
  assign y8602 = ~1'b0 ;
  assign y8603 = ~n16229 ;
  assign y8604 = ~n16230 ;
  assign y8605 = n16231 ;
  assign y8606 = ~n16233 ;
  assign y8607 = ~n16240 ;
  assign y8608 = n16244 ;
  assign y8609 = ~n16245 ;
  assign y8610 = ~n16247 ;
  assign y8611 = n16253 ;
  assign y8612 = ~1'b0 ;
  assign y8613 = n16255 ;
  assign y8614 = ~1'b0 ;
  assign y8615 = ~n16256 ;
  assign y8616 = n16257 ;
  assign y8617 = ~n16260 ;
  assign y8618 = ~n16262 ;
  assign y8619 = ~1'b0 ;
  assign y8620 = n16265 ;
  assign y8621 = ~1'b0 ;
  assign y8622 = 1'b0 ;
  assign y8623 = ~1'b0 ;
  assign y8624 = ~n16267 ;
  assign y8625 = ~1'b0 ;
  assign y8626 = n16268 ;
  assign y8627 = n16272 ;
  assign y8628 = ~n16275 ;
  assign y8629 = ~n16279 ;
  assign y8630 = ~1'b0 ;
  assign y8631 = ~1'b0 ;
  assign y8632 = ~n16280 ;
  assign y8633 = n16281 ;
  assign y8634 = n16282 ;
  assign y8635 = ~n16284 ;
  assign y8636 = n3489 ;
  assign y8637 = n16290 ;
  assign y8638 = n16291 ;
  assign y8639 = ~n16294 ;
  assign y8640 = n16299 ;
  assign y8641 = n16301 ;
  assign y8642 = ~1'b0 ;
  assign y8643 = ~1'b0 ;
  assign y8644 = n16302 ;
  assign y8645 = ~1'b0 ;
  assign y8646 = ~1'b0 ;
  assign y8647 = ~1'b0 ;
  assign y8648 = ~1'b0 ;
  assign y8649 = n16305 ;
  assign y8650 = ~n16306 ;
  assign y8651 = ~n16310 ;
  assign y8652 = 1'b0 ;
  assign y8653 = 1'b0 ;
  assign y8654 = ~1'b0 ;
  assign y8655 = 1'b0 ;
  assign y8656 = ~n1852 ;
  assign y8657 = ~1'b0 ;
  assign y8658 = ~n16313 ;
  assign y8659 = n16314 ;
  assign y8660 = n16315 ;
  assign y8661 = n16318 ;
  assign y8662 = ~n16319 ;
  assign y8663 = ~1'b0 ;
  assign y8664 = ~n2872 ;
  assign y8665 = ~1'b0 ;
  assign y8666 = ~n16320 ;
  assign y8667 = ~n16322 ;
  assign y8668 = ~1'b0 ;
  assign y8669 = n16328 ;
  assign y8670 = 1'b0 ;
  assign y8671 = ~1'b0 ;
  assign y8672 = ~1'b0 ;
  assign y8673 = 1'b0 ;
  assign y8674 = ~n16330 ;
  assign y8675 = ~1'b0 ;
  assign y8676 = ~n16332 ;
  assign y8677 = ~n16334 ;
  assign y8678 = ~n16337 ;
  assign y8679 = ~n16338 ;
  assign y8680 = n4960 ;
  assign y8681 = ~1'b0 ;
  assign y8682 = ~n16342 ;
  assign y8683 = n16346 ;
  assign y8684 = n16351 ;
  assign y8685 = n14560 ;
  assign y8686 = ~n16356 ;
  assign y8687 = ~1'b0 ;
  assign y8688 = ~n16358 ;
  assign y8689 = ~n16362 ;
  assign y8690 = n16364 ;
  assign y8691 = ~n16365 ;
  assign y8692 = n16371 ;
  assign y8693 = ~n16376 ;
  assign y8694 = ~n16377 ;
  assign y8695 = ~1'b0 ;
  assign y8696 = n16385 ;
  assign y8697 = ~1'b0 ;
  assign y8698 = n16390 ;
  assign y8699 = ~1'b0 ;
  assign y8700 = ~n16392 ;
  assign y8701 = ~n7665 ;
  assign y8702 = ~n16393 ;
  assign y8703 = n16395 ;
  assign y8704 = n16397 ;
  assign y8705 = ~1'b0 ;
  assign y8706 = n16398 ;
  assign y8707 = n16401 ;
  assign y8708 = ~1'b0 ;
  assign y8709 = ~n16404 ;
  assign y8710 = ~1'b0 ;
  assign y8711 = ~n16405 ;
  assign y8712 = n16410 ;
  assign y8713 = n16411 ;
  assign y8714 = n16412 ;
  assign y8715 = ~1'b0 ;
  assign y8716 = ~n16413 ;
  assign y8717 = ~n5380 ;
  assign y8718 = n8208 ;
  assign y8719 = ~1'b0 ;
  assign y8720 = ~n16415 ;
  assign y8721 = n16419 ;
  assign y8722 = n16422 ;
  assign y8723 = ~n16424 ;
  assign y8724 = n16426 ;
  assign y8725 = n16427 ;
  assign y8726 = n16428 ;
  assign y8727 = n16433 ;
  assign y8728 = ~n16435 ;
  assign y8729 = n16436 ;
  assign y8730 = ~1'b0 ;
  assign y8731 = ~1'b0 ;
  assign y8732 = ~1'b0 ;
  assign y8733 = ~1'b0 ;
  assign y8734 = n16439 ;
  assign y8735 = ~1'b0 ;
  assign y8736 = ~1'b0 ;
  assign y8737 = ~1'b0 ;
  assign y8738 = ~n16440 ;
  assign y8739 = ~n16447 ;
  assign y8740 = ~n16450 ;
  assign y8741 = ~1'b0 ;
  assign y8742 = ~1'b0 ;
  assign y8743 = ~n16453 ;
  assign y8744 = n16463 ;
  assign y8745 = n16465 ;
  assign y8746 = n16466 ;
  assign y8747 = ~n16467 ;
  assign y8748 = ~n16468 ;
  assign y8749 = ~1'b0 ;
  assign y8750 = ~n16470 ;
  assign y8751 = n16471 ;
  assign y8752 = ~1'b0 ;
  assign y8753 = n16472 ;
  assign y8754 = ~n16473 ;
  assign y8755 = n1119 ;
  assign y8756 = n16483 ;
  assign y8757 = ~n16487 ;
  assign y8758 = ~n16491 ;
  assign y8759 = ~1'b0 ;
  assign y8760 = n16496 ;
  assign y8761 = ~n16501 ;
  assign y8762 = ~n16504 ;
  assign y8763 = n16505 ;
  assign y8764 = ~1'b0 ;
  assign y8765 = ~1'b0 ;
  assign y8766 = ~n16507 ;
  assign y8767 = ~1'b0 ;
  assign y8768 = ~n16508 ;
  assign y8769 = ~n16509 ;
  assign y8770 = n16514 ;
  assign y8771 = ~n16515 ;
  assign y8772 = ~n16516 ;
  assign y8773 = ~n16517 ;
  assign y8774 = ~n16520 ;
  assign y8775 = ~1'b0 ;
  assign y8776 = ~1'b0 ;
  assign y8777 = n16521 ;
  assign y8778 = ~1'b0 ;
  assign y8779 = ~n16526 ;
  assign y8780 = n16530 ;
  assign y8781 = ~n16532 ;
  assign y8782 = ~n11942 ;
  assign y8783 = ~1'b0 ;
  assign y8784 = n16534 ;
  assign y8785 = ~n16535 ;
  assign y8786 = ~n16542 ;
  assign y8787 = ~n16543 ;
  assign y8788 = ~1'b0 ;
  assign y8789 = ~n16544 ;
  assign y8790 = ~1'b0 ;
  assign y8791 = ~1'b0 ;
  assign y8792 = ~n16552 ;
  assign y8793 = ~1'b0 ;
  assign y8794 = n16555 ;
  assign y8795 = n16556 ;
  assign y8796 = ~1'b0 ;
  assign y8797 = ~n2583 ;
  assign y8798 = ~n2391 ;
  assign y8799 = n16559 ;
  assign y8800 = n16560 ;
  assign y8801 = ~1'b0 ;
  assign y8802 = n16561 ;
  assign y8803 = n16566 ;
  assign y8804 = ~1'b0 ;
  assign y8805 = ~n16570 ;
  assign y8806 = n16575 ;
  assign y8807 = ~n13998 ;
  assign y8808 = ~n6155 ;
  assign y8809 = 1'b0 ;
  assign y8810 = ~1'b0 ;
  assign y8811 = n16576 ;
  assign y8812 = ~n16579 ;
  assign y8813 = ~1'b0 ;
  assign y8814 = ~n16590 ;
  assign y8815 = ~1'b0 ;
  assign y8816 = ~1'b0 ;
  assign y8817 = ~n16596 ;
  assign y8818 = ~1'b0 ;
  assign y8819 = ~n16597 ;
  assign y8820 = ~n16598 ;
  assign y8821 = ~1'b0 ;
  assign y8822 = n16602 ;
  assign y8823 = ~1'b0 ;
  assign y8824 = n16608 ;
  assign y8825 = 1'b0 ;
  assign y8826 = ~1'b0 ;
  assign y8827 = ~n16609 ;
  assign y8828 = ~n16610 ;
  assign y8829 = ~1'b0 ;
  assign y8830 = n16612 ;
  assign y8831 = n2004 ;
  assign y8832 = ~n16617 ;
  assign y8833 = ~n1300 ;
  assign y8834 = n16621 ;
  assign y8835 = ~1'b0 ;
  assign y8836 = n16627 ;
  assign y8837 = n5559 ;
  assign y8838 = ~n14950 ;
  assign y8839 = ~n16632 ;
  assign y8840 = ~n16637 ;
  assign y8841 = n16640 ;
  assign y8842 = ~1'b0 ;
  assign y8843 = n16644 ;
  assign y8844 = ~n3347 ;
  assign y8845 = ~n5119 ;
  assign y8846 = n16645 ;
  assign y8847 = ~1'b0 ;
  assign y8848 = ~1'b0 ;
  assign y8849 = 1'b0 ;
  assign y8850 = ~n16647 ;
  assign y8851 = ~1'b0 ;
  assign y8852 = ~1'b0 ;
  assign y8853 = n16653 ;
  assign y8854 = ~n16660 ;
  assign y8855 = ~n16661 ;
  assign y8856 = n16665 ;
  assign y8857 = n16666 ;
  assign y8858 = ~n16669 ;
  assign y8859 = ~1'b0 ;
  assign y8860 = ~1'b0 ;
  assign y8861 = ~n16670 ;
  assign y8862 = n16671 ;
  assign y8863 = n16672 ;
  assign y8864 = n16674 ;
  assign y8865 = ~1'b0 ;
  assign y8866 = n16676 ;
  assign y8867 = ~1'b0 ;
  assign y8868 = ~n16677 ;
  assign y8869 = ~n16678 ;
  assign y8870 = n16682 ;
  assign y8871 = ~1'b0 ;
  assign y8872 = ~1'b0 ;
  assign y8873 = ~n16686 ;
  assign y8874 = ~n16688 ;
  assign y8875 = n16689 ;
  assign y8876 = n16693 ;
  assign y8877 = ~n16695 ;
  assign y8878 = ~n16701 ;
  assign y8879 = n16702 ;
  assign y8880 = ~n16706 ;
  assign y8881 = ~n16707 ;
  assign y8882 = n16711 ;
  assign y8883 = n16713 ;
  assign y8884 = ~n16716 ;
  assign y8885 = ~1'b0 ;
  assign y8886 = ~n16718 ;
  assign y8887 = ~n16721 ;
  assign y8888 = ~1'b0 ;
  assign y8889 = n16726 ;
  assign y8890 = ~1'b0 ;
  assign y8891 = ~n16727 ;
  assign y8892 = ~n16729 ;
  assign y8893 = ~n16731 ;
  assign y8894 = n7877 ;
  assign y8895 = n16732 ;
  assign y8896 = ~n16733 ;
  assign y8897 = ~n16736 ;
  assign y8898 = ~n16738 ;
  assign y8899 = ~n16740 ;
  assign y8900 = ~1'b0 ;
  assign y8901 = n16749 ;
  assign y8902 = n16754 ;
  assign y8903 = ~n15484 ;
  assign y8904 = ~1'b0 ;
  assign y8905 = ~1'b0 ;
  assign y8906 = ~n12516 ;
  assign y8907 = ~n16757 ;
  assign y8908 = n16758 ;
  assign y8909 = n16762 ;
  assign y8910 = n16764 ;
  assign y8911 = n9440 ;
  assign y8912 = ~1'b0 ;
  assign y8913 = n16765 ;
  assign y8914 = ~1'b0 ;
  assign y8915 = ~n16767 ;
  assign y8916 = n16768 ;
  assign y8917 = n16787 ;
  assign y8918 = n16791 ;
  assign y8919 = ~n9319 ;
  assign y8920 = ~n16792 ;
  assign y8921 = n15596 ;
  assign y8922 = ~1'b0 ;
  assign y8923 = ~1'b0 ;
  assign y8924 = n16793 ;
  assign y8925 = ~n16800 ;
  assign y8926 = n16802 ;
  assign y8927 = n16804 ;
  assign y8928 = ~n16808 ;
  assign y8929 = n16810 ;
  assign y8930 = n14252 ;
  assign y8931 = ~n16811 ;
  assign y8932 = n13015 ;
  assign y8933 = n16817 ;
  assign y8934 = ~n16820 ;
  assign y8935 = ~n16821 ;
  assign y8936 = n12592 ;
  assign y8937 = n16823 ;
  assign y8938 = ~n16825 ;
  assign y8939 = n16827 ;
  assign y8940 = ~n16829 ;
  assign y8941 = ~1'b0 ;
  assign y8942 = ~1'b0 ;
  assign y8943 = n16835 ;
  assign y8944 = ~1'b0 ;
  assign y8945 = ~1'b0 ;
  assign y8946 = ~n16838 ;
  assign y8947 = ~1'b0 ;
  assign y8948 = ~1'b0 ;
  assign y8949 = ~n16840 ;
  assign y8950 = ~1'b0 ;
  assign y8951 = n16842 ;
  assign y8952 = n16843 ;
  assign y8953 = ~1'b0 ;
  assign y8954 = ~n16844 ;
  assign y8955 = n16847 ;
  assign y8956 = n16849 ;
  assign y8957 = ~1'b0 ;
  assign y8958 = n16850 ;
  assign y8959 = 1'b0 ;
  assign y8960 = n16853 ;
  assign y8961 = ~n16854 ;
  assign y8962 = ~1'b0 ;
  assign y8963 = ~n16856 ;
  assign y8964 = ~1'b0 ;
  assign y8965 = n16859 ;
  assign y8966 = ~1'b0 ;
  assign y8967 = n16863 ;
  assign y8968 = n16865 ;
  assign y8969 = n10711 ;
  assign y8970 = ~1'b0 ;
  assign y8971 = ~1'b0 ;
  assign y8972 = ~n16869 ;
  assign y8973 = ~1'b0 ;
  assign y8974 = ~1'b0 ;
  assign y8975 = ~n2805 ;
  assign y8976 = ~n16878 ;
  assign y8977 = ~n16880 ;
  assign y8978 = ~1'b0 ;
  assign y8979 = 1'b0 ;
  assign y8980 = n16881 ;
  assign y8981 = ~n1431 ;
  assign y8982 = ~n11793 ;
  assign y8983 = ~n16882 ;
  assign y8984 = n16883 ;
  assign y8985 = ~n16887 ;
  assign y8986 = n16888 ;
  assign y8987 = 1'b0 ;
  assign y8988 = ~1'b0 ;
  assign y8989 = ~n16889 ;
  assign y8990 = n16890 ;
  assign y8991 = ~1'b0 ;
  assign y8992 = ~n16894 ;
  assign y8993 = ~n16908 ;
  assign y8994 = n16915 ;
  assign y8995 = ~1'b0 ;
  assign y8996 = n16916 ;
  assign y8997 = ~n16918 ;
  assign y8998 = n16922 ;
  assign y8999 = ~1'b0 ;
  assign y9000 = ~1'b0 ;
  assign y9001 = n16924 ;
  assign y9002 = ~1'b0 ;
  assign y9003 = ~1'b0 ;
  assign y9004 = ~1'b0 ;
  assign y9005 = ~1'b0 ;
  assign y9006 = n16928 ;
  assign y9007 = ~1'b0 ;
  assign y9008 = ~1'b0 ;
  assign y9009 = n16933 ;
  assign y9010 = ~1'b0 ;
  assign y9011 = n16936 ;
  assign y9012 = ~1'b0 ;
  assign y9013 = n16939 ;
  assign y9014 = ~1'b0 ;
  assign y9015 = n16945 ;
  assign y9016 = ~1'b0 ;
  assign y9017 = ~1'b0 ;
  assign y9018 = ~n16946 ;
  assign y9019 = ~n16947 ;
  assign y9020 = ~n16950 ;
  assign y9021 = n16951 ;
  assign y9022 = ~n16954 ;
  assign y9023 = n16956 ;
  assign y9024 = n16959 ;
  assign y9025 = ~1'b0 ;
  assign y9026 = ~n16960 ;
  assign y9027 = ~n16962 ;
  assign y9028 = ~n16963 ;
  assign y9029 = ~1'b0 ;
  assign y9030 = ~n16966 ;
  assign y9031 = n16969 ;
  assign y9032 = n16975 ;
  assign y9033 = ~1'b0 ;
  assign y9034 = ~1'b0 ;
  assign y9035 = ~1'b0 ;
  assign y9036 = ~1'b0 ;
  assign y9037 = ~n16976 ;
  assign y9038 = n16980 ;
  assign y9039 = n16983 ;
  assign y9040 = n16984 ;
  assign y9041 = n16987 ;
  assign y9042 = ~n16992 ;
  assign y9043 = ~n16996 ;
  assign y9044 = ~n15619 ;
  assign y9045 = n16999 ;
  assign y9046 = ~1'b0 ;
  assign y9047 = ~1'b0 ;
  assign y9048 = ~1'b0 ;
  assign y9049 = n1943 ;
  assign y9050 = n17000 ;
  assign y9051 = ~n17001 ;
  assign y9052 = n17002 ;
  assign y9053 = n17005 ;
  assign y9054 = n17007 ;
  assign y9055 = ~n17010 ;
  assign y9056 = ~n5071 ;
  assign y9057 = ~n17011 ;
  assign y9058 = ~1'b0 ;
  assign y9059 = ~n17012 ;
  assign y9060 = ~n10403 ;
  assign y9061 = n9471 ;
  assign y9062 = ~n17013 ;
  assign y9063 = ~n17014 ;
  assign y9064 = n17015 ;
  assign y9065 = ~n17021 ;
  assign y9066 = ~n547 ;
  assign y9067 = ~n17023 ;
  assign y9068 = ~n17024 ;
  assign y9069 = ~n17034 ;
  assign y9070 = n17038 ;
  assign y9071 = ~1'b0 ;
  assign y9072 = ~n17040 ;
  assign y9073 = ~n17042 ;
  assign y9074 = n17043 ;
  assign y9075 = n17044 ;
  assign y9076 = n17045 ;
  assign y9077 = n17054 ;
  assign y9078 = ~n17057 ;
  assign y9079 = ~n17061 ;
  assign y9080 = n17063 ;
  assign y9081 = ~1'b0 ;
  assign y9082 = ~n17064 ;
  assign y9083 = ~n17066 ;
  assign y9084 = ~1'b0 ;
  assign y9085 = ~1'b0 ;
  assign y9086 = ~n17068 ;
  assign y9087 = n17070 ;
  assign y9088 = n17074 ;
  assign y9089 = ~n367 ;
  assign y9090 = ~1'b0 ;
  assign y9091 = n17079 ;
  assign y9092 = ~n17080 ;
  assign y9093 = ~n17081 ;
  assign y9094 = ~n17085 ;
  assign y9095 = n17086 ;
  assign y9096 = n17090 ;
  assign y9097 = n17092 ;
  assign y9098 = ~n17095 ;
  assign y9099 = ~n17098 ;
  assign y9100 = ~1'b0 ;
  assign y9101 = n17100 ;
  assign y9102 = ~n17102 ;
  assign y9103 = n17103 ;
  assign y9104 = n9276 ;
  assign y9105 = ~n17106 ;
  assign y9106 = ~1'b0 ;
  assign y9107 = ~n17121 ;
  assign y9108 = ~n17122 ;
  assign y9109 = ~1'b0 ;
  assign y9110 = n17124 ;
  assign y9111 = ~n17126 ;
  assign y9112 = n17128 ;
  assign y9113 = n17129 ;
  assign y9114 = n17131 ;
  assign y9115 = ~1'b0 ;
  assign y9116 = ~1'b0 ;
  assign y9117 = ~1'b0 ;
  assign y9118 = ~1'b0 ;
  assign y9119 = n17132 ;
  assign y9120 = ~1'b0 ;
  assign y9121 = n17134 ;
  assign y9122 = 1'b0 ;
  assign y9123 = ~n17139 ;
  assign y9124 = ~1'b0 ;
  assign y9125 = ~n3558 ;
  assign y9126 = ~n17140 ;
  assign y9127 = n17145 ;
  assign y9128 = ~1'b0 ;
  assign y9129 = ~1'b0 ;
  assign y9130 = n17146 ;
  assign y9131 = ~n17148 ;
  assign y9132 = ~n17150 ;
  assign y9133 = n17153 ;
  assign y9134 = ~n785 ;
  assign y9135 = ~n17155 ;
  assign y9136 = ~1'b0 ;
  assign y9137 = n17156 ;
  assign y9138 = ~1'b0 ;
  assign y9139 = ~1'b0 ;
  assign y9140 = ~n17157 ;
  assign y9141 = n17160 ;
  assign y9142 = n17164 ;
  assign y9143 = n17165 ;
  assign y9144 = n17169 ;
  assign y9145 = ~1'b0 ;
  assign y9146 = ~1'b0 ;
  assign y9147 = ~n17171 ;
  assign y9148 = ~n17174 ;
  assign y9149 = ~n17175 ;
  assign y9150 = ~n17180 ;
  assign y9151 = ~n17183 ;
  assign y9152 = n17184 ;
  assign y9153 = ~1'b0 ;
  assign y9154 = n17185 ;
  assign y9155 = ~n17187 ;
  assign y9156 = ~1'b0 ;
  assign y9157 = ~n8704 ;
  assign y9158 = ~n13554 ;
  assign y9159 = n17193 ;
  assign y9160 = ~n17198 ;
  assign y9161 = n17199 ;
  assign y9162 = ~n17201 ;
  assign y9163 = ~n17203 ;
  assign y9164 = ~n17204 ;
  assign y9165 = ~1'b0 ;
  assign y9166 = ~n17207 ;
  assign y9167 = ~n17208 ;
  assign y9168 = ~n17220 ;
  assign y9169 = ~1'b0 ;
  assign y9170 = ~n17226 ;
  assign y9171 = ~1'b0 ;
  assign y9172 = ~n17228 ;
  assign y9173 = ~1'b0 ;
  assign y9174 = ~1'b0 ;
  assign y9175 = ~n17230 ;
  assign y9176 = ~n17232 ;
  assign y9177 = ~n17233 ;
  assign y9178 = ~n17235 ;
  assign y9179 = ~1'b0 ;
  assign y9180 = ~n17237 ;
  assign y9181 = ~1'b0 ;
  assign y9182 = n17242 ;
  assign y9183 = n17246 ;
  assign y9184 = n17249 ;
  assign y9185 = n17253 ;
  assign y9186 = ~1'b0 ;
  assign y9187 = n17254 ;
  assign y9188 = ~1'b0 ;
  assign y9189 = ~n17258 ;
  assign y9190 = n17259 ;
  assign y9191 = n17264 ;
  assign y9192 = n17266 ;
  assign y9193 = ~n17268 ;
  assign y9194 = ~1'b0 ;
  assign y9195 = n17272 ;
  assign y9196 = 1'b0 ;
  assign y9197 = ~1'b0 ;
  assign y9198 = ~1'b0 ;
  assign y9199 = ~n9194 ;
  assign y9200 = ~1'b0 ;
  assign y9201 = ~1'b0 ;
  assign y9202 = ~1'b0 ;
  assign y9203 = n17274 ;
  assign y9204 = ~1'b0 ;
  assign y9205 = ~1'b0 ;
  assign y9206 = ~n17278 ;
  assign y9207 = n17285 ;
  assign y9208 = n17287 ;
  assign y9209 = ~1'b0 ;
  assign y9210 = ~n17293 ;
  assign y9211 = ~1'b0 ;
  assign y9212 = 1'b0 ;
  assign y9213 = n17295 ;
  assign y9214 = n17303 ;
  assign y9215 = ~n5158 ;
  assign y9216 = ~n17306 ;
  assign y9217 = n17312 ;
  assign y9218 = ~n17313 ;
  assign y9219 = n17314 ;
  assign y9220 = ~1'b0 ;
  assign y9221 = ~n13973 ;
  assign y9222 = ~1'b0 ;
  assign y9223 = 1'b0 ;
  assign y9224 = ~n17323 ;
  assign y9225 = n3881 ;
  assign y9226 = ~1'b0 ;
  assign y9227 = ~1'b0 ;
  assign y9228 = ~1'b0 ;
  assign y9229 = ~1'b0 ;
  assign y9230 = ~n17327 ;
  assign y9231 = ~1'b0 ;
  assign y9232 = ~n17330 ;
  assign y9233 = n8289 ;
  assign y9234 = ~1'b0 ;
  assign y9235 = ~1'b0 ;
  assign y9236 = n17331 ;
  assign y9237 = ~n8787 ;
  assign y9238 = n17333 ;
  assign y9239 = n3510 ;
  assign y9240 = ~n7655 ;
  assign y9241 = ~1'b0 ;
  assign y9242 = ~n17336 ;
  assign y9243 = n17338 ;
  assign y9244 = ~1'b0 ;
  assign y9245 = n4328 ;
  assign y9246 = n17339 ;
  assign y9247 = ~n17343 ;
  assign y9248 = n17345 ;
  assign y9249 = n5768 ;
  assign y9250 = ~1'b0 ;
  assign y9251 = n17348 ;
  assign y9252 = ~n17352 ;
  assign y9253 = n17355 ;
  assign y9254 = ~n17357 ;
  assign y9255 = n17360 ;
  assign y9256 = ~n17363 ;
  assign y9257 = 1'b0 ;
  assign y9258 = ~n17367 ;
  assign y9259 = ~n17368 ;
  assign y9260 = ~n136 ;
  assign y9261 = ~1'b0 ;
  assign y9262 = ~n17375 ;
  assign y9263 = n17377 ;
  assign y9264 = n17378 ;
  assign y9265 = n17379 ;
  assign y9266 = n6856 ;
  assign y9267 = 1'b0 ;
  assign y9268 = ~1'b0 ;
  assign y9269 = n17383 ;
  assign y9270 = ~n17384 ;
  assign y9271 = n17385 ;
  assign y9272 = n17387 ;
  assign y9273 = ~n17388 ;
  assign y9274 = n17390 ;
  assign y9275 = ~n17394 ;
  assign y9276 = ~n17395 ;
  assign y9277 = ~1'b0 ;
  assign y9278 = n17399 ;
  assign y9279 = ~1'b0 ;
  assign y9280 = n17400 ;
  assign y9281 = ~n17402 ;
  assign y9282 = n16707 ;
  assign y9283 = ~n17409 ;
  assign y9284 = ~n17410 ;
  assign y9285 = n17411 ;
  assign y9286 = ~1'b0 ;
  assign y9287 = ~n17412 ;
  assign y9288 = ~n17415 ;
  assign y9289 = n17416 ;
  assign y9290 = ~n17418 ;
  assign y9291 = ~1'b0 ;
  assign y9292 = ~1'b0 ;
  assign y9293 = ~1'b0 ;
  assign y9294 = n17420 ;
  assign y9295 = n17421 ;
  assign y9296 = ~1'b0 ;
  assign y9297 = n12280 ;
  assign y9298 = ~1'b0 ;
  assign y9299 = ~n17429 ;
  assign y9300 = n17431 ;
  assign y9301 = n17432 ;
  assign y9302 = ~n17433 ;
  assign y9303 = ~n17437 ;
  assign y9304 = ~1'b0 ;
  assign y9305 = n17441 ;
  assign y9306 = ~1'b0 ;
  assign y9307 = ~1'b0 ;
  assign y9308 = ~n17448 ;
  assign y9309 = ~1'b0 ;
  assign y9310 = ~n17453 ;
  assign y9311 = ~n17455 ;
  assign y9312 = ~1'b0 ;
  assign y9313 = ~1'b0 ;
  assign y9314 = ~n17457 ;
  assign y9315 = ~n17461 ;
  assign y9316 = n17463 ;
  assign y9317 = ~1'b0 ;
  assign y9318 = ~n17468 ;
  assign y9319 = ~n17474 ;
  assign y9320 = ~1'b0 ;
  assign y9321 = ~1'b0 ;
  assign y9322 = ~1'b0 ;
  assign y9323 = ~n17476 ;
  assign y9324 = ~n17486 ;
  assign y9325 = ~1'b0 ;
  assign y9326 = n17487 ;
  assign y9327 = n17490 ;
  assign y9328 = ~n17497 ;
  assign y9329 = ~n8904 ;
  assign y9330 = 1'b0 ;
  assign y9331 = ~n17500 ;
  assign y9332 = ~n17503 ;
  assign y9333 = n17506 ;
  assign y9334 = ~n17509 ;
  assign y9335 = ~1'b0 ;
  assign y9336 = ~n17510 ;
  assign y9337 = ~1'b0 ;
  assign y9338 = n17511 ;
  assign y9339 = ~1'b0 ;
  assign y9340 = ~1'b0 ;
  assign y9341 = ~1'b0 ;
  assign y9342 = ~1'b0 ;
  assign y9343 = n17513 ;
  assign y9344 = ~1'b0 ;
  assign y9345 = n17514 ;
  assign y9346 = n16335 ;
  assign y9347 = n17516 ;
  assign y9348 = ~1'b0 ;
  assign y9349 = ~1'b0 ;
  assign y9350 = ~n17518 ;
  assign y9351 = ~1'b0 ;
  assign y9352 = 1'b0 ;
  assign y9353 = 1'b0 ;
  assign y9354 = n17526 ;
  assign y9355 = ~n17531 ;
  assign y9356 = ~n17535 ;
  assign y9357 = ~n17543 ;
  assign y9358 = 1'b0 ;
  assign y9359 = n17544 ;
  assign y9360 = ~1'b0 ;
  assign y9361 = ~n17546 ;
  assign y9362 = n17549 ;
  assign y9363 = ~n17551 ;
  assign y9364 = ~1'b0 ;
  assign y9365 = n17554 ;
  assign y9366 = ~n17557 ;
  assign y9367 = 1'b0 ;
  assign y9368 = ~n14598 ;
  assign y9369 = ~1'b0 ;
  assign y9370 = ~1'b0 ;
  assign y9371 = 1'b0 ;
  assign y9372 = ~n17558 ;
  assign y9373 = ~n17560 ;
  assign y9374 = ~n17563 ;
  assign y9375 = ~1'b0 ;
  assign y9376 = ~n17564 ;
  assign y9377 = ~n17567 ;
  assign y9378 = ~n17571 ;
  assign y9379 = ~1'b0 ;
  assign y9380 = ~1'b0 ;
  assign y9381 = ~n17573 ;
  assign y9382 = ~1'b0 ;
  assign y9383 = ~1'b0 ;
  assign y9384 = ~n17577 ;
  assign y9385 = n17579 ;
  assign y9386 = ~1'b0 ;
  assign y9387 = ~n17580 ;
  assign y9388 = ~1'b0 ;
  assign y9389 = n17583 ;
  assign y9390 = n17586 ;
  assign y9391 = 1'b0 ;
  assign y9392 = ~n17587 ;
  assign y9393 = ~n17596 ;
  assign y9394 = n17601 ;
  assign y9395 = n17604 ;
  assign y9396 = n17612 ;
  assign y9397 = ~n17615 ;
  assign y9398 = ~1'b0 ;
  assign y9399 = ~1'b0 ;
  assign y9400 = ~n17616 ;
  assign y9401 = ~1'b0 ;
  assign y9402 = ~1'b0 ;
  assign y9403 = n17618 ;
  assign y9404 = ~n17622 ;
  assign y9405 = ~n17624 ;
  assign y9406 = ~1'b0 ;
  assign y9407 = ~n17626 ;
  assign y9408 = ~n17634 ;
  assign y9409 = ~n17635 ;
  assign y9410 = ~1'b0 ;
  assign y9411 = n17637 ;
  assign y9412 = n17638 ;
  assign y9413 = ~1'b0 ;
  assign y9414 = ~n10670 ;
  assign y9415 = ~1'b0 ;
  assign y9416 = ~1'b0 ;
  assign y9417 = ~n17639 ;
  assign y9418 = n17640 ;
  assign y9419 = ~1'b0 ;
  assign y9420 = ~n17642 ;
  assign y9421 = ~1'b0 ;
  assign y9422 = n17643 ;
  assign y9423 = ~n17647 ;
  assign y9424 = n17648 ;
  assign y9425 = n4888 ;
  assign y9426 = ~n17652 ;
  assign y9427 = ~1'b0 ;
  assign y9428 = ~n17655 ;
  assign y9429 = ~1'b0 ;
  assign y9430 = n17656 ;
  assign y9431 = n17657 ;
  assign y9432 = ~1'b0 ;
  assign y9433 = ~1'b0 ;
  assign y9434 = n17658 ;
  assign y9435 = n4348 ;
  assign y9436 = n17661 ;
  assign y9437 = n17664 ;
  assign y9438 = n17665 ;
  assign y9439 = n13377 ;
  assign y9440 = n17666 ;
  assign y9441 = n17669 ;
  assign y9442 = ~1'b0 ;
  assign y9443 = ~n17670 ;
  assign y9444 = n17673 ;
  assign y9445 = ~1'b0 ;
  assign y9446 = n17678 ;
  assign y9447 = ~1'b0 ;
  assign y9448 = ~n17679 ;
  assign y9449 = ~n17680 ;
  assign y9450 = n7089 ;
  assign y9451 = n17681 ;
  assign y9452 = ~1'b0 ;
  assign y9453 = ~n16010 ;
  assign y9454 = ~n17683 ;
  assign y9455 = n17684 ;
  assign y9456 = n17688 ;
  assign y9457 = ~n17691 ;
  assign y9458 = n17693 ;
  assign y9459 = ~n17694 ;
  assign y9460 = ~n13355 ;
  assign y9461 = ~1'b0 ;
  assign y9462 = ~1'b0 ;
  assign y9463 = ~1'b0 ;
  assign y9464 = ~n17695 ;
  assign y9465 = ~n17696 ;
  assign y9466 = ~1'b0 ;
  assign y9467 = ~1'b0 ;
  assign y9468 = ~n8529 ;
  assign y9469 = ~n17698 ;
  assign y9470 = ~n17702 ;
  assign y9471 = n17706 ;
  assign y9472 = n15206 ;
  assign y9473 = n17709 ;
  assign y9474 = ~1'b0 ;
  assign y9475 = n17715 ;
  assign y9476 = n17721 ;
  assign y9477 = n17727 ;
  assign y9478 = ~1'b0 ;
  assign y9479 = ~1'b0 ;
  assign y9480 = ~1'b0 ;
  assign y9481 = ~n17729 ;
  assign y9482 = n17731 ;
  assign y9483 = n17739 ;
  assign y9484 = ~1'b0 ;
  assign y9485 = ~n17743 ;
  assign y9486 = ~n17746 ;
  assign y9487 = ~1'b0 ;
  assign y9488 = ~n17747 ;
  assign y9489 = ~1'b0 ;
  assign y9490 = ~n17751 ;
  assign y9491 = ~1'b0 ;
  assign y9492 = ~n17760 ;
  assign y9493 = ~n17763 ;
  assign y9494 = ~n17767 ;
  assign y9495 = ~n17769 ;
  assign y9496 = ~n17770 ;
  assign y9497 = ~n17773 ;
  assign y9498 = ~n17774 ;
  assign y9499 = ~n17775 ;
  assign y9500 = ~n16002 ;
  assign y9501 = ~n17779 ;
  assign y9502 = n17783 ;
  assign y9503 = ~1'b0 ;
  assign y9504 = n17785 ;
  assign y9505 = n17787 ;
  assign y9506 = ~n124 ;
  assign y9507 = ~1'b0 ;
  assign y9508 = n17789 ;
  assign y9509 = ~n17797 ;
  assign y9510 = ~n17798 ;
  assign y9511 = ~n17800 ;
  assign y9512 = ~1'b0 ;
  assign y9513 = ~1'b0 ;
  assign y9514 = n14853 ;
  assign y9515 = n17804 ;
  assign y9516 = ~n7008 ;
  assign y9517 = ~1'b0 ;
  assign y9518 = n17802 ;
  assign y9519 = ~n17805 ;
  assign y9520 = n17806 ;
  assign y9521 = n17807 ;
  assign y9522 = n17809 ;
  assign y9523 = n17816 ;
  assign y9524 = n17820 ;
  assign y9525 = ~n2097 ;
  assign y9526 = 1'b0 ;
  assign y9527 = ~n17821 ;
  assign y9528 = ~1'b0 ;
  assign y9529 = ~1'b0 ;
  assign y9530 = n17825 ;
  assign y9531 = ~1'b0 ;
  assign y9532 = ~n17827 ;
  assign y9533 = ~1'b0 ;
  assign y9534 = n4545 ;
  assign y9535 = ~n17828 ;
  assign y9536 = ~1'b0 ;
  assign y9537 = 1'b0 ;
  assign y9538 = n17834 ;
  assign y9539 = ~n17839 ;
  assign y9540 = n17841 ;
  assign y9541 = ~1'b0 ;
  assign y9542 = ~1'b0 ;
  assign y9543 = n17850 ;
  assign y9544 = ~n17853 ;
  assign y9545 = n17858 ;
  assign y9546 = n14082 ;
  assign y9547 = ~1'b0 ;
  assign y9548 = ~1'b0 ;
  assign y9549 = n17859 ;
  assign y9550 = ~1'b0 ;
  assign y9551 = n11193 ;
  assign y9552 = ~1'b0 ;
  assign y9553 = ~1'b0 ;
  assign y9554 = ~n6099 ;
  assign y9555 = ~n17860 ;
  assign y9556 = ~1'b0 ;
  assign y9557 = n17862 ;
  assign y9558 = ~n17864 ;
  assign y9559 = ~n17868 ;
  assign y9560 = ~n17869 ;
  assign y9561 = ~n17879 ;
  assign y9562 = ~1'b0 ;
  assign y9563 = ~1'b0 ;
  assign y9564 = n17881 ;
  assign y9565 = n17886 ;
  assign y9566 = n17888 ;
  assign y9567 = ~1'b0 ;
  assign y9568 = ~n17891 ;
  assign y9569 = n17310 ;
  assign y9570 = ~n17892 ;
  assign y9571 = ~n17893 ;
  assign y9572 = ~1'b0 ;
  assign y9573 = n16714 ;
  assign y9574 = ~1'b0 ;
  assign y9575 = n17897 ;
  assign y9576 = n17901 ;
  assign y9577 = n17902 ;
  assign y9578 = n17904 ;
  assign y9579 = ~n17913 ;
  assign y9580 = ~1'b0 ;
  assign y9581 = ~n17917 ;
  assign y9582 = ~1'b0 ;
  assign y9583 = ~1'b0 ;
  assign y9584 = ~n17922 ;
  assign y9585 = n17926 ;
  assign y9586 = ~n17929 ;
  assign y9587 = ~1'b0 ;
  assign y9588 = n17931 ;
  assign y9589 = ~n17932 ;
  assign y9590 = n17934 ;
  assign y9591 = n17936 ;
  assign y9592 = ~n17937 ;
  assign y9593 = n17939 ;
  assign y9594 = ~n17940 ;
  assign y9595 = n17943 ;
  assign y9596 = ~1'b0 ;
  assign y9597 = ~1'b0 ;
  assign y9598 = ~1'b0 ;
  assign y9599 = n17945 ;
  assign y9600 = ~1'b0 ;
  assign y9601 = n17946 ;
  assign y9602 = ~n17961 ;
  assign y9603 = n17962 ;
  assign y9604 = n17963 ;
  assign y9605 = n17965 ;
  assign y9606 = n17966 ;
  assign y9607 = ~1'b0 ;
  assign y9608 = ~n17968 ;
  assign y9609 = n17969 ;
  assign y9610 = 1'b0 ;
  assign y9611 = ~1'b0 ;
  assign y9612 = ~n17972 ;
  assign y9613 = n17974 ;
  assign y9614 = ~n17978 ;
  assign y9615 = ~1'b0 ;
  assign y9616 = n17980 ;
  assign y9617 = n17981 ;
  assign y9618 = ~1'b0 ;
  assign y9619 = n4702 ;
  assign y9620 = n17982 ;
  assign y9621 = ~1'b0 ;
  assign y9622 = ~1'b0 ;
  assign y9623 = ~1'b0 ;
  assign y9624 = ~1'b0 ;
  assign y9625 = ~n17983 ;
  assign y9626 = ~n17984 ;
  assign y9627 = ~1'b0 ;
  assign y9628 = n17986 ;
  assign y9629 = ~n17987 ;
  assign y9630 = n17990 ;
  assign y9631 = n17992 ;
  assign y9632 = ~n17996 ;
  assign y9633 = ~n17998 ;
  assign y9634 = ~1'b0 ;
  assign y9635 = ~n18002 ;
  assign y9636 = 1'b0 ;
  assign y9637 = ~n18004 ;
  assign y9638 = n18006 ;
  assign y9639 = n18007 ;
  assign y9640 = ~n18010 ;
  assign y9641 = ~n18013 ;
  assign y9642 = ~1'b0 ;
  assign y9643 = ~n18014 ;
  assign y9644 = ~n18016 ;
  assign y9645 = n18017 ;
  assign y9646 = ~n18018 ;
  assign y9647 = ~n18019 ;
  assign y9648 = ~1'b0 ;
  assign y9649 = ~1'b0 ;
  assign y9650 = ~1'b0 ;
  assign y9651 = ~n18021 ;
  assign y9652 = ~1'b0 ;
  assign y9653 = n18024 ;
  assign y9654 = n18025 ;
  assign y9655 = ~n18027 ;
  assign y9656 = n18033 ;
  assign y9657 = ~n18034 ;
  assign y9658 = n18035 ;
  assign y9659 = ~n18037 ;
  assign y9660 = ~1'b0 ;
  assign y9661 = ~n18039 ;
  assign y9662 = n5001 ;
  assign y9663 = ~1'b0 ;
  assign y9664 = ~1'b0 ;
  assign y9665 = ~1'b0 ;
  assign y9666 = ~n18042 ;
  assign y9667 = n18049 ;
  assign y9668 = n18050 ;
  assign y9669 = ~n18051 ;
  assign y9670 = n18052 ;
  assign y9671 = ~1'b0 ;
  assign y9672 = ~n18055 ;
  assign y9673 = ~n7342 ;
  assign y9674 = n18059 ;
  assign y9675 = ~n18070 ;
  assign y9676 = ~n18076 ;
  assign y9677 = n18084 ;
  assign y9678 = ~1'b0 ;
  assign y9679 = ~1'b0 ;
  assign y9680 = ~n18087 ;
  assign y9681 = ~1'b0 ;
  assign y9682 = ~n18089 ;
  assign y9683 = n18091 ;
  assign y9684 = ~n18092 ;
  assign y9685 = ~n18099 ;
  assign y9686 = ~n18100 ;
  assign y9687 = n18104 ;
  assign y9688 = n18108 ;
  assign y9689 = ~1'b0 ;
  assign y9690 = ~n18110 ;
  assign y9691 = ~1'b0 ;
  assign y9692 = ~n18115 ;
  assign y9693 = ~1'b0 ;
  assign y9694 = ~1'b0 ;
  assign y9695 = n18117 ;
  assign y9696 = n18125 ;
  assign y9697 = n18126 ;
  assign y9698 = ~n18132 ;
  assign y9699 = n18134 ;
  assign y9700 = ~n18136 ;
  assign y9701 = ~n18138 ;
  assign y9702 = n18140 ;
  assign y9703 = ~n18144 ;
  assign y9704 = n18146 ;
  assign y9705 = ~1'b0 ;
  assign y9706 = ~1'b0 ;
  assign y9707 = ~n8421 ;
  assign y9708 = n18147 ;
  assign y9709 = ~1'b0 ;
  assign y9710 = ~n18149 ;
  assign y9711 = ~n18152 ;
  assign y9712 = n18158 ;
  assign y9713 = n18162 ;
  assign y9714 = n18164 ;
  assign y9715 = ~n18166 ;
  assign y9716 = n18169 ;
  assign y9717 = ~n15060 ;
  assign y9718 = ~1'b0 ;
  assign y9719 = ~n18171 ;
  assign y9720 = ~n18173 ;
  assign y9721 = ~1'b0 ;
  assign y9722 = ~1'b0 ;
  assign y9723 = ~n18178 ;
  assign y9724 = ~n18181 ;
  assign y9725 = ~n18183 ;
  assign y9726 = ~n2460 ;
  assign y9727 = n18185 ;
  assign y9728 = ~n18186 ;
  assign y9729 = ~n18192 ;
  assign y9730 = ~n18194 ;
  assign y9731 = n333 ;
  assign y9732 = n8705 ;
  assign y9733 = ~n18197 ;
  assign y9734 = n18200 ;
  assign y9735 = 1'b0 ;
  assign y9736 = ~n18205 ;
  assign y9737 = ~n18207 ;
  assign y9738 = ~n18208 ;
  assign y9739 = ~1'b0 ;
  assign y9740 = n18210 ;
  assign y9741 = ~n15804 ;
  assign y9742 = ~1'b0 ;
  assign y9743 = n18213 ;
  assign y9744 = ~n18220 ;
  assign y9745 = ~n18226 ;
  assign y9746 = n18227 ;
  assign y9747 = ~1'b0 ;
  assign y9748 = ~n18229 ;
  assign y9749 = ~n18236 ;
  assign y9750 = n18240 ;
  assign y9751 = ~n18242 ;
  assign y9752 = n812 ;
  assign y9753 = n18245 ;
  assign y9754 = ~n12510 ;
  assign y9755 = ~1'b0 ;
  assign y9756 = ~1'b0 ;
  assign y9757 = ~1'b0 ;
  assign y9758 = ~1'b0 ;
  assign y9759 = ~n18246 ;
  assign y9760 = ~1'b0 ;
  assign y9761 = ~1'b0 ;
  assign y9762 = ~1'b0 ;
  assign y9763 = ~n12228 ;
  assign y9764 = ~1'b0 ;
  assign y9765 = ~n18248 ;
  assign y9766 = ~1'b0 ;
  assign y9767 = n18249 ;
  assign y9768 = ~n18250 ;
  assign y9769 = ~n18252 ;
  assign y9770 = ~1'b0 ;
  assign y9771 = n18256 ;
  assign y9772 = ~n18258 ;
  assign y9773 = n18261 ;
  assign y9774 = ~n18264 ;
  assign y9775 = ~n18268 ;
  assign y9776 = ~n18270 ;
  assign y9777 = ~1'b0 ;
  assign y9778 = ~1'b0 ;
  assign y9779 = ~n18271 ;
  assign y9780 = ~n18272 ;
  assign y9781 = ~1'b0 ;
  assign y9782 = ~n18274 ;
  assign y9783 = ~1'b0 ;
  assign y9784 = 1'b0 ;
  assign y9785 = ~n18276 ;
  assign y9786 = ~1'b0 ;
  assign y9787 = ~n18281 ;
  assign y9788 = ~1'b0 ;
  assign y9789 = n18283 ;
  assign y9790 = ~1'b0 ;
  assign y9791 = ~n18288 ;
  assign y9792 = ~1'b0 ;
  assign y9793 = n18289 ;
  assign y9794 = ~n18291 ;
  assign y9795 = n13626 ;
  assign y9796 = 1'b0 ;
  assign y9797 = n18299 ;
  assign y9798 = ~1'b0 ;
  assign y9799 = n18304 ;
  assign y9800 = ~1'b0 ;
  assign y9801 = ~1'b0 ;
  assign y9802 = ~1'b0 ;
  assign y9803 = ~n18308 ;
  assign y9804 = n18309 ;
  assign y9805 = ~1'b0 ;
  assign y9806 = ~n18317 ;
  assign y9807 = n18322 ;
  assign y9808 = n7653 ;
  assign y9809 = ~1'b0 ;
  assign y9810 = ~n18327 ;
  assign y9811 = n18329 ;
  assign y9812 = n18332 ;
  assign y9813 = ~n362 ;
  assign y9814 = ~n18335 ;
  assign y9815 = n18338 ;
  assign y9816 = ~n18343 ;
  assign y9817 = ~1'b0 ;
  assign y9818 = ~n18345 ;
  assign y9819 = n18352 ;
  assign y9820 = n18353 ;
  assign y9821 = ~n18357 ;
  assign y9822 = ~1'b0 ;
  assign y9823 = ~1'b0 ;
  assign y9824 = ~1'b0 ;
  assign y9825 = n18360 ;
  assign y9826 = ~1'b0 ;
  assign y9827 = 1'b0 ;
  assign y9828 = ~1'b0 ;
  assign y9829 = n2581 ;
  assign y9830 = ~1'b0 ;
  assign y9831 = n18364 ;
  assign y9832 = ~1'b0 ;
  assign y9833 = ~n18368 ;
  assign y9834 = ~1'b0 ;
  assign y9835 = n18369 ;
  assign y9836 = ~1'b0 ;
  assign y9837 = n18372 ;
  assign y9838 = n18374 ;
  assign y9839 = ~1'b0 ;
  assign y9840 = n18378 ;
  assign y9841 = n18379 ;
  assign y9842 = ~1'b0 ;
  assign y9843 = n18381 ;
  assign y9844 = ~1'b0 ;
  assign y9845 = ~1'b0 ;
  assign y9846 = ~1'b0 ;
  assign y9847 = ~n18385 ;
  assign y9848 = ~n18386 ;
  assign y9849 = n18388 ;
  assign y9850 = ~n10968 ;
  assign y9851 = ~1'b0 ;
  assign y9852 = ~1'b0 ;
  assign y9853 = ~1'b0 ;
  assign y9854 = n18390 ;
  assign y9855 = ~1'b0 ;
  assign y9856 = 1'b0 ;
  assign y9857 = ~1'b0 ;
  assign y9858 = ~n18398 ;
  assign y9859 = ~n18399 ;
  assign y9860 = ~1'b0 ;
  assign y9861 = ~n18404 ;
  assign y9862 = ~1'b0 ;
  assign y9863 = 1'b0 ;
  assign y9864 = n18407 ;
  assign y9865 = ~1'b0 ;
  assign y9866 = ~n1178 ;
  assign y9867 = n18410 ;
  assign y9868 = ~1'b0 ;
  assign y9869 = n18411 ;
  assign y9870 = n18413 ;
  assign y9871 = ~1'b0 ;
  assign y9872 = ~n18414 ;
  assign y9873 = n18420 ;
  assign y9874 = n18423 ;
  assign y9875 = n18429 ;
  assign y9876 = n13520 ;
  assign y9877 = n18430 ;
  assign y9878 = ~n18433 ;
  assign y9879 = n18439 ;
  assign y9880 = n18442 ;
  assign y9881 = n18443 ;
  assign y9882 = ~n17684 ;
  assign y9883 = n18449 ;
  assign y9884 = ~1'b0 ;
  assign y9885 = n18450 ;
  assign y9886 = n18452 ;
  assign y9887 = n18453 ;
  assign y9888 = ~n18454 ;
  assign y9889 = n18455 ;
  assign y9890 = ~n18460 ;
  assign y9891 = n282 ;
  assign y9892 = ~n18465 ;
  assign y9893 = n18468 ;
  assign y9894 = n18470 ;
  assign y9895 = n18472 ;
  assign y9896 = ~1'b0 ;
  assign y9897 = ~1'b0 ;
  assign y9898 = ~1'b0 ;
  assign y9899 = n18473 ;
  assign y9900 = ~n18475 ;
  assign y9901 = ~n18477 ;
  assign y9902 = ~n18480 ;
  assign y9903 = ~n18485 ;
  assign y9904 = ~n18488 ;
  assign y9905 = ~1'b0 ;
  assign y9906 = n18489 ;
  assign y9907 = n18500 ;
  assign y9908 = n18502 ;
  assign y9909 = ~n7110 ;
  assign y9910 = ~n18505 ;
  assign y9911 = n18506 ;
  assign y9912 = ~n18507 ;
  assign y9913 = n18508 ;
  assign y9914 = ~n18510 ;
  assign y9915 = n18514 ;
  assign y9916 = n18520 ;
  assign y9917 = ~n18523 ;
  assign y9918 = n18529 ;
  assign y9919 = n11934 ;
  assign y9920 = ~1'b0 ;
  assign y9921 = ~n18530 ;
  assign y9922 = ~1'b0 ;
  assign y9923 = ~1'b0 ;
  assign y9924 = ~1'b0 ;
  assign y9925 = ~1'b0 ;
  assign y9926 = n18533 ;
  assign y9927 = ~1'b0 ;
  assign y9928 = ~n18538 ;
  assign y9929 = ~1'b0 ;
  assign y9930 = n18542 ;
  assign y9931 = 1'b0 ;
  assign y9932 = n18549 ;
  assign y9933 = ~n18550 ;
  assign y9934 = ~n18551 ;
  assign y9935 = ~n18554 ;
  assign y9936 = ~1'b0 ;
  assign y9937 = n18556 ;
  assign y9938 = n18558 ;
  assign y9939 = n18559 ;
  assign y9940 = n18560 ;
  assign y9941 = ~n18561 ;
  assign y9942 = ~n18562 ;
  assign y9943 = ~1'b0 ;
  assign y9944 = ~1'b0 ;
  assign y9945 = ~1'b0 ;
  assign y9946 = ~1'b0 ;
  assign y9947 = ~1'b0 ;
  assign y9948 = ~n18564 ;
  assign y9949 = n18565 ;
  assign y9950 = n18583 ;
  assign y9951 = ~1'b0 ;
  assign y9952 = ~1'b0 ;
  assign y9953 = n18585 ;
  assign y9954 = ~n18588 ;
  assign y9955 = ~n18589 ;
  assign y9956 = 1'b0 ;
  assign y9957 = ~n18591 ;
  assign y9958 = ~n18593 ;
  assign y9959 = ~1'b0 ;
  assign y9960 = ~1'b0 ;
  assign y9961 = 1'b0 ;
  assign y9962 = ~1'b0 ;
  assign y9963 = ~n18594 ;
  assign y9964 = ~n18597 ;
  assign y9965 = n18599 ;
  assign y9966 = ~n18600 ;
  assign y9967 = ~1'b0 ;
  assign y9968 = n11572 ;
  assign y9969 = ~n18602 ;
  assign y9970 = ~n18603 ;
  assign y9971 = ~n18607 ;
  assign y9972 = ~n18608 ;
  assign y9973 = n18610 ;
  assign y9974 = ~n18612 ;
  assign y9975 = ~n18620 ;
  assign y9976 = ~n18622 ;
  assign y9977 = ~n18625 ;
  assign y9978 = n18634 ;
  assign y9979 = n18636 ;
  assign y9980 = ~1'b0 ;
  assign y9981 = ~1'b0 ;
  assign y9982 = 1'b0 ;
  assign y9983 = n18637 ;
  assign y9984 = ~1'b0 ;
  assign y9985 = ~n18643 ;
  assign y9986 = ~n18645 ;
  assign y9987 = n18652 ;
  assign y9988 = 1'b0 ;
  assign y9989 = ~n18654 ;
  assign y9990 = ~n18659 ;
  assign y9991 = ~1'b0 ;
  assign y9992 = n18664 ;
  assign y9993 = ~n18665 ;
  assign y9994 = ~n18667 ;
  assign y9995 = ~n18670 ;
  assign y9996 = ~n18671 ;
  assign y9997 = 1'b0 ;
  assign y9998 = ~n18672 ;
  assign y9999 = n18673 ;
  assign y10000 = ~1'b0 ;
  assign y10001 = ~1'b0 ;
  assign y10002 = ~1'b0 ;
  assign y10003 = n18676 ;
  assign y10004 = n18677 ;
  assign y10005 = ~1'b0 ;
  assign y10006 = ~1'b0 ;
  assign y10007 = n18678 ;
  assign y10008 = ~1'b0 ;
  assign y10009 = ~1'b0 ;
  assign y10010 = n18681 ;
  assign y10011 = ~1'b0 ;
  assign y10012 = n18685 ;
  assign y10013 = ~1'b0 ;
  assign y10014 = ~1'b0 ;
  assign y10015 = ~n18695 ;
  assign y10016 = n18699 ;
  assign y10017 = n18704 ;
  assign y10018 = n18709 ;
  assign y10019 = n1157 ;
  assign y10020 = ~n3181 ;
  assign y10021 = ~n18712 ;
  assign y10022 = ~n18714 ;
  assign y10023 = n18719 ;
  assign y10024 = n3061 ;
  assign y10025 = n18721 ;
  assign y10026 = ~1'b0 ;
  assign y10027 = ~n10728 ;
  assign y10028 = ~1'b0 ;
  assign y10029 = n18729 ;
  assign y10030 = n18732 ;
  assign y10031 = ~n18736 ;
  assign y10032 = n18738 ;
  assign y10033 = ~n18739 ;
  assign y10034 = ~n18740 ;
  assign y10035 = ~1'b0 ;
  assign y10036 = ~n18741 ;
  assign y10037 = n18743 ;
  assign y10038 = ~1'b0 ;
  assign y10039 = n18748 ;
  assign y10040 = ~n18753 ;
  assign y10041 = ~1'b0 ;
  assign y10042 = ~1'b0 ;
  assign y10043 = n18754 ;
  assign y10044 = ~1'b0 ;
  assign y10045 = n18757 ;
  assign y10046 = ~n18759 ;
  assign y10047 = n18760 ;
  assign y10048 = n18761 ;
  assign y10049 = n18764 ;
  assign y10050 = n18767 ;
  assign y10051 = n18768 ;
  assign y10052 = ~n18770 ;
  assign y10053 = n18774 ;
  assign y10054 = n18778 ;
  assign y10055 = ~1'b0 ;
  assign y10056 = ~n18782 ;
  assign y10057 = 1'b0 ;
  assign y10058 = ~n14385 ;
  assign y10059 = ~n18784 ;
  assign y10060 = ~n18786 ;
  assign y10061 = ~1'b0 ;
  assign y10062 = n18793 ;
  assign y10063 = ~n18794 ;
  assign y10064 = ~1'b0 ;
  assign y10065 = n18796 ;
  assign y10066 = n18801 ;
  assign y10067 = n18803 ;
  assign y10068 = n18804 ;
  assign y10069 = ~n18807 ;
  assign y10070 = ~n18810 ;
  assign y10071 = n18811 ;
  assign y10072 = ~n18812 ;
  assign y10073 = ~n18815 ;
  assign y10074 = 1'b0 ;
  assign y10075 = n18823 ;
  assign y10076 = ~n18824 ;
  assign y10077 = n4962 ;
  assign y10078 = ~n18827 ;
  assign y10079 = n18833 ;
  assign y10080 = ~1'b0 ;
  assign y10081 = n18836 ;
  assign y10082 = ~1'b0 ;
  assign y10083 = ~n18837 ;
  assign y10084 = ~n18841 ;
  assign y10085 = ~1'b0 ;
  assign y10086 = ~n3442 ;
  assign y10087 = ~n18844 ;
  assign y10088 = ~1'b0 ;
  assign y10089 = n18846 ;
  assign y10090 = n18847 ;
  assign y10091 = n18848 ;
  assign y10092 = ~1'b0 ;
  assign y10093 = ~1'b0 ;
  assign y10094 = ~n18854 ;
  assign y10095 = n18856 ;
  assign y10096 = n18858 ;
  assign y10097 = ~n18860 ;
  assign y10098 = ~n18864 ;
  assign y10099 = ~n18867 ;
  assign y10100 = 1'b0 ;
  assign y10101 = ~n18870 ;
  assign y10102 = ~1'b0 ;
  assign y10103 = ~n9536 ;
  assign y10104 = ~1'b0 ;
  assign y10105 = ~n18878 ;
  assign y10106 = n18882 ;
  assign y10107 = n18884 ;
  assign y10108 = n18889 ;
  assign y10109 = n18890 ;
  assign y10110 = n12215 ;
  assign y10111 = ~1'b0 ;
  assign y10112 = ~1'b0 ;
  assign y10113 = ~n18892 ;
  assign y10114 = ~n18894 ;
  assign y10115 = ~n18895 ;
  assign y10116 = ~n18897 ;
  assign y10117 = ~n3012 ;
  assign y10118 = ~n18900 ;
  assign y10119 = ~n18902 ;
  assign y10120 = ~n18905 ;
  assign y10121 = ~n18907 ;
  assign y10122 = 1'b0 ;
  assign y10123 = ~1'b0 ;
  assign y10124 = n18910 ;
  assign y10125 = n18912 ;
  assign y10126 = ~n18913 ;
  assign y10127 = ~1'b0 ;
  assign y10128 = n18917 ;
  assign y10129 = ~n18918 ;
  assign y10130 = ~n11954 ;
  assign y10131 = ~n18923 ;
  assign y10132 = ~n18925 ;
  assign y10133 = ~n18927 ;
  assign y10134 = ~n18929 ;
  assign y10135 = n18930 ;
  assign y10136 = ~n18934 ;
  assign y10137 = ~n18938 ;
  assign y10138 = ~1'b0 ;
  assign y10139 = ~n18940 ;
  assign y10140 = n18943 ;
  assign y10141 = ~1'b0 ;
  assign y10142 = n18948 ;
  assign y10143 = ~n18954 ;
  assign y10144 = n18955 ;
  assign y10145 = ~n18956 ;
  assign y10146 = ~n18957 ;
  assign y10147 = ~1'b0 ;
  assign y10148 = n18960 ;
  assign y10149 = ~1'b0 ;
  assign y10150 = n18965 ;
  assign y10151 = n18966 ;
  assign y10152 = ~n18971 ;
  assign y10153 = n18980 ;
  assign y10154 = ~n18982 ;
  assign y10155 = ~n18988 ;
  assign y10156 = ~n18989 ;
  assign y10157 = ~1'b0 ;
  assign y10158 = n18990 ;
  assign y10159 = ~1'b0 ;
  assign y10160 = ~n14846 ;
  assign y10161 = n18991 ;
  assign y10162 = n18992 ;
  assign y10163 = ~1'b0 ;
  assign y10164 = ~n18994 ;
  assign y10165 = ~n3392 ;
  assign y10166 = n18995 ;
  assign y10167 = ~n18996 ;
  assign y10168 = 1'b0 ;
  assign y10169 = ~n18999 ;
  assign y10170 = ~n19001 ;
  assign y10171 = ~n19004 ;
  assign y10172 = ~1'b0 ;
  assign y10173 = ~n19006 ;
  assign y10174 = n19013 ;
  assign y10175 = ~1'b0 ;
  assign y10176 = ~1'b0 ;
  assign y10177 = ~1'b0 ;
  assign y10178 = ~n19016 ;
  assign y10179 = ~n19024 ;
  assign y10180 = n19027 ;
  assign y10181 = ~1'b0 ;
  assign y10182 = ~n19028 ;
  assign y10183 = ~1'b0 ;
  assign y10184 = ~n19034 ;
  assign y10185 = ~1'b0 ;
  assign y10186 = ~n19036 ;
  assign y10187 = ~1'b0 ;
  assign y10188 = ~n19037 ;
  assign y10189 = ~1'b0 ;
  assign y10190 = ~n19038 ;
  assign y10191 = n12322 ;
  assign y10192 = n19040 ;
  assign y10193 = ~n19046 ;
  assign y10194 = n19054 ;
  assign y10195 = ~n19056 ;
  assign y10196 = n19060 ;
  assign y10197 = ~n19063 ;
  assign y10198 = n19067 ;
  assign y10199 = n19072 ;
  assign y10200 = n19073 ;
  assign y10201 = ~n19074 ;
  assign y10202 = n1469 ;
  assign y10203 = ~n19076 ;
  assign y10204 = ~1'b0 ;
  assign y10205 = ~n19078 ;
  assign y10206 = n12275 ;
  assign y10207 = ~n19079 ;
  assign y10208 = ~n19081 ;
  assign y10209 = n19084 ;
  assign y10210 = n19085 ;
  assign y10211 = ~1'b0 ;
  assign y10212 = ~n19086 ;
  assign y10213 = ~1'b0 ;
  assign y10214 = ~1'b0 ;
  assign y10215 = 1'b0 ;
  assign y10216 = ~n19094 ;
  assign y10217 = ~1'b0 ;
  assign y10218 = n19095 ;
  assign y10219 = ~n19097 ;
  assign y10220 = n19098 ;
  assign y10221 = ~n19100 ;
  assign y10222 = n19105 ;
  assign y10223 = n19107 ;
  assign y10224 = n19109 ;
  assign y10225 = n19116 ;
  assign y10226 = ~1'b0 ;
  assign y10227 = n1323 ;
  assign y10228 = ~n19120 ;
  assign y10229 = ~1'b0 ;
  assign y10230 = ~n19126 ;
  assign y10231 = n19128 ;
  assign y10232 = ~n19129 ;
  assign y10233 = ~n19131 ;
  assign y10234 = n19136 ;
  assign y10235 = ~1'b0 ;
  assign y10236 = n19143 ;
  assign y10237 = ~1'b0 ;
  assign y10238 = ~n19149 ;
  assign y10239 = ~n19153 ;
  assign y10240 = n3909 ;
  assign y10241 = ~1'b0 ;
  assign y10242 = n19158 ;
  assign y10243 = ~1'b0 ;
  assign y10244 = ~1'b0 ;
  assign y10245 = ~n19159 ;
  assign y10246 = ~1'b0 ;
  assign y10247 = n19160 ;
  assign y10248 = n19161 ;
  assign y10249 = n19172 ;
  assign y10250 = ~n19173 ;
  assign y10251 = ~n13205 ;
  assign y10252 = ~n19178 ;
  assign y10253 = ~n19184 ;
  assign y10254 = ~1'b0 ;
  assign y10255 = 1'b0 ;
  assign y10256 = n19188 ;
  assign y10257 = ~1'b0 ;
  assign y10258 = ~1'b0 ;
  assign y10259 = n19189 ;
  assign y10260 = ~1'b0 ;
  assign y10261 = n19190 ;
  assign y10262 = ~n19191 ;
  assign y10263 = n19200 ;
  assign y10264 = ~1'b0 ;
  assign y10265 = ~n19206 ;
  assign y10266 = n19208 ;
  assign y10267 = ~n19212 ;
  assign y10268 = ~1'b0 ;
  assign y10269 = n19214 ;
  assign y10270 = n19216 ;
  assign y10271 = ~1'b0 ;
  assign y10272 = ~n19218 ;
  assign y10273 = n19219 ;
  assign y10274 = ~n15034 ;
  assign y10275 = 1'b0 ;
  assign y10276 = ~n19220 ;
  assign y10277 = n19221 ;
  assign y10278 = ~n19228 ;
  assign y10279 = ~n19229 ;
  assign y10280 = n19231 ;
  assign y10281 = ~n19233 ;
  assign y10282 = ~1'b0 ;
  assign y10283 = ~n19234 ;
  assign y10284 = n19235 ;
  assign y10285 = ~1'b0 ;
  assign y10286 = ~1'b0 ;
  assign y10287 = ~1'b0 ;
  assign y10288 = ~n19237 ;
  assign y10289 = n3572 ;
  assign y10290 = ~n19238 ;
  assign y10291 = ~1'b0 ;
  assign y10292 = ~1'b0 ;
  assign y10293 = ~n19240 ;
  assign y10294 = ~1'b0 ;
  assign y10295 = n19243 ;
  assign y10296 = ~n19246 ;
  assign y10297 = ~1'b0 ;
  assign y10298 = ~1'b0 ;
  assign y10299 = ~1'b0 ;
  assign y10300 = 1'b0 ;
  assign y10301 = ~n19247 ;
  assign y10302 = ~1'b0 ;
  assign y10303 = ~n19248 ;
  assign y10304 = ~1'b0 ;
  assign y10305 = ~1'b0 ;
  assign y10306 = n5519 ;
  assign y10307 = ~n19251 ;
  assign y10308 = ~1'b0 ;
  assign y10309 = n19252 ;
  assign y10310 = ~1'b0 ;
  assign y10311 = ~n19254 ;
  assign y10312 = ~n19255 ;
  assign y10313 = n19257 ;
  assign y10314 = n19261 ;
  assign y10315 = ~1'b0 ;
  assign y10316 = ~n19263 ;
  assign y10317 = n19265 ;
  assign y10318 = ~1'b0 ;
  assign y10319 = ~1'b0 ;
  assign y10320 = ~n19268 ;
  assign y10321 = ~n19269 ;
  assign y10322 = n19270 ;
  assign y10323 = ~n19275 ;
  assign y10324 = ~1'b0 ;
  assign y10325 = ~1'b0 ;
  assign y10326 = ~1'b0 ;
  assign y10327 = ~1'b0 ;
  assign y10328 = ~1'b0 ;
  assign y10329 = ~1'b0 ;
  assign y10330 = ~n13529 ;
  assign y10331 = n5497 ;
  assign y10332 = n19281 ;
  assign y10333 = ~n19287 ;
  assign y10334 = n19288 ;
  assign y10335 = ~1'b0 ;
  assign y10336 = ~1'b0 ;
  assign y10337 = ~n19289 ;
  assign y10338 = ~n19293 ;
  assign y10339 = n19300 ;
  assign y10340 = n19304 ;
  assign y10341 = n19308 ;
  assign y10342 = ~1'b0 ;
  assign y10343 = ~1'b0 ;
  assign y10344 = 1'b0 ;
  assign y10345 = ~1'b0 ;
  assign y10346 = n19310 ;
  assign y10347 = n19311 ;
  assign y10348 = ~1'b0 ;
  assign y10349 = n19317 ;
  assign y10350 = n19318 ;
  assign y10351 = n19321 ;
  assign y10352 = n19322 ;
  assign y10353 = ~1'b0 ;
  assign y10354 = n19325 ;
  assign y10355 = n19327 ;
  assign y10356 = ~n19336 ;
  assign y10357 = n19341 ;
  assign y10358 = n19345 ;
  assign y10359 = n19349 ;
  assign y10360 = ~n19353 ;
  assign y10361 = ~n19354 ;
  assign y10362 = ~n19356 ;
  assign y10363 = ~1'b0 ;
  assign y10364 = n19358 ;
  assign y10365 = n12673 ;
  assign y10366 = ~1'b0 ;
  assign y10367 = ~n19359 ;
  assign y10368 = ~n2650 ;
  assign y10369 = ~n19362 ;
  assign y10370 = n19367 ;
  assign y10371 = ~n10755 ;
  assign y10372 = n19370 ;
  assign y10373 = ~1'b0 ;
  assign y10374 = ~n12860 ;
  assign y10375 = n19372 ;
  assign y10376 = n19374 ;
  assign y10377 = n19376 ;
  assign y10378 = ~1'b0 ;
  assign y10379 = ~1'b0 ;
  assign y10380 = ~n19377 ;
  assign y10381 = ~1'b0 ;
  assign y10382 = ~1'b0 ;
  assign y10383 = ~n19378 ;
  assign y10384 = n1430 ;
  assign y10385 = 1'b0 ;
  assign y10386 = ~1'b0 ;
  assign y10387 = ~1'b0 ;
  assign y10388 = n19383 ;
  assign y10389 = n15614 ;
  assign y10390 = ~1'b0 ;
  assign y10391 = 1'b0 ;
  assign y10392 = n19385 ;
  assign y10393 = ~n19386 ;
  assign y10394 = n19390 ;
  assign y10395 = n19392 ;
  assign y10396 = n19394 ;
  assign y10397 = ~n19395 ;
  assign y10398 = n19396 ;
  assign y10399 = ~n19401 ;
  assign y10400 = ~1'b0 ;
  assign y10401 = ~n19406 ;
  assign y10402 = n19407 ;
  assign y10403 = ~1'b0 ;
  assign y10404 = ~n19412 ;
  assign y10405 = ~1'b0 ;
  assign y10406 = ~1'b0 ;
  assign y10407 = ~1'b0 ;
  assign y10408 = ~1'b0 ;
  assign y10409 = ~1'b0 ;
  assign y10410 = n19414 ;
  assign y10411 = 1'b0 ;
  assign y10412 = n19419 ;
  assign y10413 = n19422 ;
  assign y10414 = ~n19425 ;
  assign y10415 = ~1'b0 ;
  assign y10416 = ~1'b0 ;
  assign y10417 = ~n19430 ;
  assign y10418 = n19439 ;
  assign y10419 = ~n19440 ;
  assign y10420 = ~n19442 ;
  assign y10421 = ~n17262 ;
  assign y10422 = n19445 ;
  assign y10423 = ~1'b0 ;
  assign y10424 = ~1'b0 ;
  assign y10425 = ~n19448 ;
  assign y10426 = ~n19452 ;
  assign y10427 = n19453 ;
  assign y10428 = ~n19458 ;
  assign y10429 = ~1'b0 ;
  assign y10430 = n6060 ;
  assign y10431 = ~1'b0 ;
  assign y10432 = ~n19461 ;
  assign y10433 = ~1'b0 ;
  assign y10434 = 1'b0 ;
  assign y10435 = ~n19466 ;
  assign y10436 = n19469 ;
  assign y10437 = ~n19471 ;
  assign y10438 = ~n19473 ;
  assign y10439 = ~1'b0 ;
  assign y10440 = ~1'b0 ;
  assign y10441 = n19477 ;
  assign y10442 = n19478 ;
  assign y10443 = ~1'b0 ;
  assign y10444 = n19485 ;
  assign y10445 = ~1'b0 ;
  assign y10446 = ~1'b0 ;
  assign y10447 = ~n13520 ;
  assign y10448 = n19486 ;
  assign y10449 = ~1'b0 ;
  assign y10450 = n19491 ;
  assign y10451 = n19492 ;
  assign y10452 = ~n19493 ;
  assign y10453 = ~1'b0 ;
  assign y10454 = n19495 ;
  assign y10455 = ~1'b0 ;
  assign y10456 = ~n19498 ;
  assign y10457 = ~1'b0 ;
  assign y10458 = ~1'b0 ;
  assign y10459 = n19499 ;
  assign y10460 = ~n19500 ;
  assign y10461 = ~n19502 ;
  assign y10462 = ~n8012 ;
  assign y10463 = n19507 ;
  assign y10464 = ~n19514 ;
  assign y10465 = n19515 ;
  assign y10466 = ~n19518 ;
  assign y10467 = n19519 ;
  assign y10468 = ~1'b0 ;
  assign y10469 = n19523 ;
  assign y10470 = n19525 ;
  assign y10471 = n19529 ;
  assign y10472 = n19536 ;
  assign y10473 = n19538 ;
  assign y10474 = n19542 ;
  assign y10475 = ~n19543 ;
  assign y10476 = 1'b0 ;
  assign y10477 = ~1'b0 ;
  assign y10478 = ~n19544 ;
  assign y10479 = ~n19550 ;
  assign y10480 = ~1'b0 ;
  assign y10481 = ~1'b0 ;
  assign y10482 = n16931 ;
  assign y10483 = n19551 ;
  assign y10484 = ~n19554 ;
  assign y10485 = ~1'b0 ;
  assign y10486 = ~n19560 ;
  assign y10487 = ~n19564 ;
  assign y10488 = ~n19568 ;
  assign y10489 = ~1'b0 ;
  assign y10490 = ~n19569 ;
  assign y10491 = ~n19571 ;
  assign y10492 = n19573 ;
  assign y10493 = ~1'b0 ;
  assign y10494 = 1'b0 ;
  assign y10495 = ~n2415 ;
  assign y10496 = ~n19576 ;
  assign y10497 = ~1'b0 ;
  assign y10498 = ~n19579 ;
  assign y10499 = ~1'b0 ;
  assign y10500 = n6198 ;
  assign y10501 = n19581 ;
  assign y10502 = 1'b0 ;
  assign y10503 = ~n19586 ;
  assign y10504 = ~n19587 ;
  assign y10505 = ~n19588 ;
  assign y10506 = ~1'b0 ;
  assign y10507 = n19591 ;
  assign y10508 = ~n19598 ;
  assign y10509 = ~n19600 ;
  assign y10510 = ~1'b0 ;
  assign y10511 = n19601 ;
  assign y10512 = n19602 ;
  assign y10513 = n19603 ;
  assign y10514 = ~n19607 ;
  assign y10515 = ~1'b0 ;
  assign y10516 = ~1'b0 ;
  assign y10517 = ~1'b0 ;
  assign y10518 = ~n12415 ;
  assign y10519 = ~1'b0 ;
  assign y10520 = ~n19608 ;
  assign y10521 = ~n19609 ;
  assign y10522 = n19611 ;
  assign y10523 = n19613 ;
  assign y10524 = n19615 ;
  assign y10525 = ~n19624 ;
  assign y10526 = ~1'b0 ;
  assign y10527 = ~1'b0 ;
  assign y10528 = n19626 ;
  assign y10529 = ~1'b0 ;
  assign y10530 = ~1'b0 ;
  assign y10531 = ~1'b0 ;
  assign y10532 = n18466 ;
  assign y10533 = n19631 ;
  assign y10534 = ~n9931 ;
  assign y10535 = ~n19634 ;
  assign y10536 = ~n19635 ;
  assign y10537 = ~n19640 ;
  assign y10538 = n19643 ;
  assign y10539 = ~n19644 ;
  assign y10540 = ~1'b0 ;
  assign y10541 = ~n19650 ;
  assign y10542 = ~n19653 ;
  assign y10543 = ~1'b0 ;
  assign y10544 = n19655 ;
  assign y10545 = ~1'b0 ;
  assign y10546 = ~1'b0 ;
  assign y10547 = ~1'b0 ;
  assign y10548 = ~n19661 ;
  assign y10549 = ~n19662 ;
  assign y10550 = ~n19664 ;
  assign y10551 = n19667 ;
  assign y10552 = 1'b0 ;
  assign y10553 = ~n19672 ;
  assign y10554 = ~n19674 ;
  assign y10555 = ~1'b0 ;
  assign y10556 = ~n19675 ;
  assign y10557 = n19677 ;
  assign y10558 = ~n19681 ;
  assign y10559 = ~1'b0 ;
  assign y10560 = ~n19683 ;
  assign y10561 = n19685 ;
  assign y10562 = 1'b0 ;
  assign y10563 = n19687 ;
  assign y10564 = ~n19693 ;
  assign y10565 = ~n19699 ;
  assign y10566 = 1'b0 ;
  assign y10567 = n19701 ;
  assign y10568 = ~1'b0 ;
  assign y10569 = ~1'b0 ;
  assign y10570 = ~1'b0 ;
  assign y10571 = ~n19702 ;
  assign y10572 = ~1'b0 ;
  assign y10573 = ~1'b0 ;
  assign y10574 = ~1'b0 ;
  assign y10575 = ~1'b0 ;
  assign y10576 = n19703 ;
  assign y10577 = n19710 ;
  assign y10578 = 1'b0 ;
  assign y10579 = ~1'b0 ;
  assign y10580 = ~n19712 ;
  assign y10581 = n19713 ;
  assign y10582 = ~1'b0 ;
  assign y10583 = ~n16479 ;
  assign y10584 = ~n19718 ;
  assign y10585 = ~n19721 ;
  assign y10586 = ~n3637 ;
  assign y10587 = n19723 ;
  assign y10588 = ~1'b0 ;
  assign y10589 = ~n19725 ;
  assign y10590 = ~1'b0 ;
  assign y10591 = 1'b0 ;
  assign y10592 = n19726 ;
  assign y10593 = n19727 ;
  assign y10594 = n9232 ;
  assign y10595 = ~1'b0 ;
  assign y10596 = n19729 ;
  assign y10597 = n14598 ;
  assign y10598 = ~n19732 ;
  assign y10599 = 1'b0 ;
  assign y10600 = ~n19734 ;
  assign y10601 = ~n19737 ;
  assign y10602 = ~n19738 ;
  assign y10603 = ~1'b0 ;
  assign y10604 = ~n19740 ;
  assign y10605 = n19744 ;
  assign y10606 = ~1'b0 ;
  assign y10607 = 1'b0 ;
  assign y10608 = ~1'b0 ;
  assign y10609 = ~1'b0 ;
  assign y10610 = n19745 ;
  assign y10611 = n19749 ;
  assign y10612 = ~n19750 ;
  assign y10613 = n19752 ;
  assign y10614 = n2789 ;
  assign y10615 = ~1'b0 ;
  assign y10616 = ~1'b0 ;
  assign y10617 = ~1'b0 ;
  assign y10618 = ~n19753 ;
  assign y10619 = ~n19754 ;
  assign y10620 = ~1'b0 ;
  assign y10621 = ~1'b0 ;
  assign y10622 = n19756 ;
  assign y10623 = ~n19757 ;
  assign y10624 = ~1'b0 ;
  assign y10625 = n19759 ;
  assign y10626 = n19760 ;
  assign y10627 = ~n19764 ;
  assign y10628 = ~n19767 ;
  assign y10629 = ~1'b0 ;
  assign y10630 = n19769 ;
  assign y10631 = ~n19775 ;
  assign y10632 = n19776 ;
  assign y10633 = n19778 ;
  assign y10634 = ~1'b0 ;
  assign y10635 = 1'b0 ;
  assign y10636 = ~1'b0 ;
  assign y10637 = n19780 ;
  assign y10638 = n19787 ;
  assign y10639 = ~n19788 ;
  assign y10640 = ~n19789 ;
  assign y10641 = ~1'b0 ;
  assign y10642 = ~n19791 ;
  assign y10643 = ~n19795 ;
  assign y10644 = 1'b0 ;
  assign y10645 = ~n19796 ;
  assign y10646 = n19799 ;
  assign y10647 = n19801 ;
  assign y10648 = ~n12261 ;
  assign y10649 = ~n19802 ;
  assign y10650 = ~n19804 ;
  assign y10651 = ~n19807 ;
  assign y10652 = ~n19809 ;
  assign y10653 = n19810 ;
  assign y10654 = n19811 ;
  assign y10655 = ~1'b0 ;
  assign y10656 = n4677 ;
  assign y10657 = ~1'b0 ;
  assign y10658 = n19813 ;
  assign y10659 = ~n19816 ;
  assign y10660 = n19820 ;
  assign y10661 = ~1'b0 ;
  assign y10662 = n19824 ;
  assign y10663 = n19826 ;
  assign y10664 = ~n19828 ;
  assign y10665 = n18502 ;
  assign y10666 = ~n19829 ;
  assign y10667 = ~1'b0 ;
  assign y10668 = n10804 ;
  assign y10669 = n19830 ;
  assign y10670 = ~n19836 ;
  assign y10671 = n19839 ;
  assign y10672 = ~1'b0 ;
  assign y10673 = ~1'b0 ;
  assign y10674 = ~1'b0 ;
  assign y10675 = ~1'b0 ;
  assign y10676 = ~n19843 ;
  assign y10677 = ~n12520 ;
  assign y10678 = ~n19846 ;
  assign y10679 = ~1'b0 ;
  assign y10680 = ~n19847 ;
  assign y10681 = ~n19849 ;
  assign y10682 = n19854 ;
  assign y10683 = ~n19875 ;
  assign y10684 = ~1'b0 ;
  assign y10685 = ~1'b0 ;
  assign y10686 = n19880 ;
  assign y10687 = n5130 ;
  assign y10688 = ~n11553 ;
  assign y10689 = ~1'b0 ;
  assign y10690 = ~n19881 ;
  assign y10691 = n19882 ;
  assign y10692 = n3896 ;
  assign y10693 = n19884 ;
  assign y10694 = n12588 ;
  assign y10695 = ~1'b0 ;
  assign y10696 = ~n19886 ;
  assign y10697 = ~1'b0 ;
  assign y10698 = n19890 ;
  assign y10699 = n19891 ;
  assign y10700 = n19892 ;
  assign y10701 = ~n19895 ;
  assign y10702 = n19896 ;
  assign y10703 = ~n19902 ;
  assign y10704 = ~n19905 ;
  assign y10705 = ~n19906 ;
  assign y10706 = ~1'b0 ;
  assign y10707 = n5901 ;
  assign y10708 = ~1'b0 ;
  assign y10709 = n19907 ;
  assign y10710 = ~n19908 ;
  assign y10711 = n19909 ;
  assign y10712 = ~n19910 ;
  assign y10713 = ~1'b0 ;
  assign y10714 = n19915 ;
  assign y10715 = ~n19916 ;
  assign y10716 = ~n19918 ;
  assign y10717 = ~n19919 ;
  assign y10718 = ~n19925 ;
  assign y10719 = ~1'b0 ;
  assign y10720 = ~n19926 ;
  assign y10721 = ~1'b0 ;
  assign y10722 = ~1'b0 ;
  assign y10723 = ~1'b0 ;
  assign y10724 = n19927 ;
  assign y10725 = ~n19929 ;
  assign y10726 = ~n74 ;
  assign y10727 = ~1'b0 ;
  assign y10728 = ~1'b0 ;
  assign y10729 = ~n19930 ;
  assign y10730 = 1'b0 ;
  assign y10731 = ~n19932 ;
  assign y10732 = 1'b0 ;
  assign y10733 = n19935 ;
  assign y10734 = ~n19937 ;
  assign y10735 = n19941 ;
  assign y10736 = n19942 ;
  assign y10737 = n19943 ;
  assign y10738 = n19947 ;
  assign y10739 = ~1'b0 ;
  assign y10740 = n19949 ;
  assign y10741 = ~1'b0 ;
  assign y10742 = n19958 ;
  assign y10743 = n19961 ;
  assign y10744 = ~1'b0 ;
  assign y10745 = n19964 ;
  assign y10746 = ~n19969 ;
  assign y10747 = ~n19976 ;
  assign y10748 = ~n19980 ;
  assign y10749 = n19981 ;
  assign y10750 = n19983 ;
  assign y10751 = ~1'b0 ;
  assign y10752 = n19984 ;
  assign y10753 = ~n19987 ;
  assign y10754 = n19989 ;
  assign y10755 = ~1'b0 ;
  assign y10756 = ~1'b0 ;
  assign y10757 = n16015 ;
  assign y10758 = n19991 ;
  assign y10759 = n19992 ;
  assign y10760 = n20001 ;
  assign y10761 = ~n938 ;
  assign y10762 = n20004 ;
  assign y10763 = ~1'b0 ;
  assign y10764 = ~1'b0 ;
  assign y10765 = ~1'b0 ;
  assign y10766 = ~n20007 ;
  assign y10767 = n20008 ;
  assign y10768 = n20011 ;
  assign y10769 = ~1'b0 ;
  assign y10770 = ~n20019 ;
  assign y10771 = ~1'b0 ;
  assign y10772 = n20020 ;
  assign y10773 = n20022 ;
  assign y10774 = ~1'b0 ;
  assign y10775 = ~1'b0 ;
  assign y10776 = n20024 ;
  assign y10777 = n1469 ;
  assign y10778 = ~n2324 ;
  assign y10779 = ~n20025 ;
  assign y10780 = ~1'b0 ;
  assign y10781 = ~n20026 ;
  assign y10782 = ~n20027 ;
  assign y10783 = ~1'b0 ;
  assign y10784 = n20030 ;
  assign y10785 = ~1'b0 ;
  assign y10786 = ~1'b0 ;
  assign y10787 = n20046 ;
  assign y10788 = ~1'b0 ;
  assign y10789 = ~n20047 ;
  assign y10790 = n20051 ;
  assign y10791 = n20059 ;
  assign y10792 = ~1'b0 ;
  assign y10793 = n20060 ;
  assign y10794 = ~1'b0 ;
  assign y10795 = ~n20065 ;
  assign y10796 = ~1'b0 ;
  assign y10797 = ~n20069 ;
  assign y10798 = ~n20070 ;
  assign y10799 = ~1'b0 ;
  assign y10800 = n20073 ;
  assign y10801 = ~1'b0 ;
  assign y10802 = n20075 ;
  assign y10803 = ~n20077 ;
  assign y10804 = n20078 ;
  assign y10805 = n20082 ;
  assign y10806 = n20083 ;
  assign y10807 = ~n20084 ;
  assign y10808 = ~n20088 ;
  assign y10809 = ~1'b0 ;
  assign y10810 = n20090 ;
  assign y10811 = n20092 ;
  assign y10812 = 1'b0 ;
  assign y10813 = ~n20097 ;
  assign y10814 = ~n20099 ;
  assign y10815 = n20108 ;
  assign y10816 = n17554 ;
  assign y10817 = ~1'b0 ;
  assign y10818 = 1'b0 ;
  assign y10819 = ~1'b0 ;
  assign y10820 = 1'b0 ;
  assign y10821 = n20112 ;
  assign y10822 = n20114 ;
  assign y10823 = n20116 ;
  assign y10824 = n20117 ;
  assign y10825 = n8117 ;
  assign y10826 = n20120 ;
  assign y10827 = ~n20122 ;
  assign y10828 = n20123 ;
  assign y10829 = ~n20131 ;
  assign y10830 = n20137 ;
  assign y10831 = n2478 ;
  assign y10832 = n20138 ;
  assign y10833 = ~1'b0 ;
  assign y10834 = ~n20139 ;
  assign y10835 = ~1'b0 ;
  assign y10836 = ~1'b0 ;
  assign y10837 = n20140 ;
  assign y10838 = ~n20141 ;
  assign y10839 = n20142 ;
  assign y10840 = ~n20148 ;
  assign y10841 = ~n20150 ;
  assign y10842 = n20151 ;
  assign y10843 = ~1'b0 ;
  assign y10844 = n20154 ;
  assign y10845 = ~1'b0 ;
  assign y10846 = n20155 ;
  assign y10847 = ~1'b0 ;
  assign y10848 = ~n20162 ;
  assign y10849 = ~1'b0 ;
  assign y10850 = ~1'b0 ;
  assign y10851 = n13692 ;
  assign y10852 = n20171 ;
  assign y10853 = 1'b0 ;
  assign y10854 = ~1'b0 ;
  assign y10855 = n19512 ;
  assign y10856 = ~n20172 ;
  assign y10857 = 1'b0 ;
  assign y10858 = n20175 ;
  assign y10859 = ~1'b0 ;
  assign y10860 = ~1'b0 ;
  assign y10861 = ~n20176 ;
  assign y10862 = ~1'b0 ;
  assign y10863 = ~n20177 ;
  assign y10864 = n20185 ;
  assign y10865 = n20189 ;
  assign y10866 = n20193 ;
  assign y10867 = ~1'b0 ;
  assign y10868 = ~1'b0 ;
  assign y10869 = n20198 ;
  assign y10870 = ~1'b0 ;
  assign y10871 = ~1'b0 ;
  assign y10872 = n20204 ;
  assign y10873 = ~1'b0 ;
  assign y10874 = ~n20205 ;
  assign y10875 = ~n20209 ;
  assign y10876 = ~n20220 ;
  assign y10877 = ~n20221 ;
  assign y10878 = n20222 ;
  assign y10879 = ~n20225 ;
  assign y10880 = n20228 ;
  assign y10881 = ~1'b0 ;
  assign y10882 = ~1'b0 ;
  assign y10883 = n20229 ;
  assign y10884 = ~n20234 ;
  assign y10885 = n20237 ;
  assign y10886 = n20239 ;
  assign y10887 = ~1'b0 ;
  assign y10888 = ~n20247 ;
  assign y10889 = ~n2361 ;
  assign y10890 = n20249 ;
  assign y10891 = ~n20252 ;
  assign y10892 = ~1'b0 ;
  assign y10893 = ~n20255 ;
  assign y10894 = n20258 ;
  assign y10895 = n20259 ;
  assign y10896 = n20263 ;
  assign y10897 = 1'b0 ;
  assign y10898 = n20270 ;
  assign y10899 = ~n20271 ;
  assign y10900 = ~n20276 ;
  assign y10901 = ~n20277 ;
  assign y10902 = 1'b0 ;
  assign y10903 = ~1'b0 ;
  assign y10904 = n20278 ;
  assign y10905 = n2233 ;
  assign y10906 = ~n20280 ;
  assign y10907 = ~n20282 ;
  assign y10908 = ~n8217 ;
  assign y10909 = ~n20283 ;
  assign y10910 = ~n20287 ;
  assign y10911 = n20288 ;
  assign y10912 = n20289 ;
  assign y10913 = n20291 ;
  assign y10914 = 1'b0 ;
  assign y10915 = n20292 ;
  assign y10916 = n20294 ;
  assign y10917 = ~1'b0 ;
  assign y10918 = n20295 ;
  assign y10919 = ~n20296 ;
  assign y10920 = ~1'b0 ;
  assign y10921 = ~n20297 ;
  assign y10922 = ~1'b0 ;
  assign y10923 = ~n20299 ;
  assign y10924 = 1'b0 ;
  assign y10925 = ~n20301 ;
  assign y10926 = n20307 ;
  assign y10927 = n20308 ;
  assign y10928 = ~1'b0 ;
  assign y10929 = ~n20309 ;
  assign y10930 = ~n20311 ;
  assign y10931 = 1'b0 ;
  assign y10932 = ~n20317 ;
  assign y10933 = ~1'b0 ;
  assign y10934 = ~1'b0 ;
  assign y10935 = ~1'b0 ;
  assign y10936 = ~1'b0 ;
  assign y10937 = n20318 ;
  assign y10938 = ~1'b0 ;
  assign y10939 = 1'b0 ;
  assign y10940 = n20320 ;
  assign y10941 = ~n20289 ;
  assign y10942 = ~1'b0 ;
  assign y10943 = ~n20323 ;
  assign y10944 = ~1'b0 ;
  assign y10945 = ~1'b0 ;
  assign y10946 = ~n20327 ;
  assign y10947 = ~1'b0 ;
  assign y10948 = n20328 ;
  assign y10949 = n20329 ;
  assign y10950 = ~1'b0 ;
  assign y10951 = n6665 ;
  assign y10952 = ~1'b0 ;
  assign y10953 = ~1'b0 ;
  assign y10954 = ~n20335 ;
  assign y10955 = ~n20336 ;
  assign y10956 = ~n20341 ;
  assign y10957 = n20342 ;
  assign y10958 = ~n20345 ;
  assign y10959 = ~1'b0 ;
  assign y10960 = n20346 ;
  assign y10961 = ~n8879 ;
  assign y10962 = n20347 ;
  assign y10963 = ~n20351 ;
  assign y10964 = ~1'b0 ;
  assign y10965 = n20357 ;
  assign y10966 = ~n20363 ;
  assign y10967 = ~n20366 ;
  assign y10968 = ~1'b0 ;
  assign y10969 = ~n20368 ;
  assign y10970 = ~1'b0 ;
  assign y10971 = n4517 ;
  assign y10972 = ~1'b0 ;
  assign y10973 = ~n20373 ;
  assign y10974 = ~n20376 ;
  assign y10975 = n3443 ;
  assign y10976 = ~1'b0 ;
  assign y10977 = ~1'b0 ;
  assign y10978 = n20378 ;
  assign y10979 = ~n20379 ;
  assign y10980 = 1'b0 ;
  assign y10981 = ~n20380 ;
  assign y10982 = ~1'b0 ;
  assign y10983 = ~1'b0 ;
  assign y10984 = n20382 ;
  assign y10985 = ~1'b0 ;
  assign y10986 = n20386 ;
  assign y10987 = n798 ;
  assign y10988 = n774 ;
  assign y10989 = n20388 ;
  assign y10990 = ~1'b0 ;
  assign y10991 = ~1'b0 ;
  assign y10992 = ~1'b0 ;
  assign y10993 = n20390 ;
  assign y10994 = ~n800 ;
  assign y10995 = n20391 ;
  assign y10996 = n20394 ;
  assign y10997 = ~n20395 ;
  assign y10998 = n20401 ;
  assign y10999 = n20406 ;
  assign y11000 = ~1'b0 ;
  assign y11001 = n20407 ;
  assign y11002 = ~1'b0 ;
  assign y11003 = n20411 ;
  assign y11004 = ~1'b0 ;
  assign y11005 = ~1'b0 ;
  assign y11006 = n20412 ;
  assign y11007 = n20414 ;
  assign y11008 = ~1'b0 ;
  assign y11009 = n10103 ;
  assign y11010 = ~n20415 ;
  assign y11011 = ~1'b0 ;
  assign y11012 = n7427 ;
  assign y11013 = n20417 ;
  assign y11014 = ~n20418 ;
  assign y11015 = n20422 ;
  assign y11016 = n20426 ;
  assign y11017 = ~1'b0 ;
  assign y11018 = ~1'b0 ;
  assign y11019 = n20428 ;
  assign y11020 = ~1'b0 ;
  assign y11021 = n20435 ;
  assign y11022 = ~n20437 ;
  assign y11023 = n20438 ;
  assign y11024 = ~1'b0 ;
  assign y11025 = ~1'b0 ;
  assign y11026 = 1'b0 ;
  assign y11027 = n20441 ;
  assign y11028 = ~n20444 ;
  assign y11029 = n20445 ;
  assign y11030 = n20448 ;
  assign y11031 = ~1'b0 ;
  assign y11032 = ~n20451 ;
  assign y11033 = ~n20452 ;
  assign y11034 = ~n17968 ;
  assign y11035 = n20453 ;
  assign y11036 = ~n20454 ;
  assign y11037 = ~n7040 ;
  assign y11038 = n20462 ;
  assign y11039 = ~1'b0 ;
  assign y11040 = ~1'b0 ;
  assign y11041 = ~1'b0 ;
  assign y11042 = ~n20463 ;
  assign y11043 = n20465 ;
  assign y11044 = ~n20474 ;
  assign y11045 = n20475 ;
  assign y11046 = n20476 ;
  assign y11047 = n20479 ;
  assign y11048 = n20481 ;
  assign y11049 = ~1'b0 ;
  assign y11050 = ~1'b0 ;
  assign y11051 = n20483 ;
  assign y11052 = ~n20484 ;
  assign y11053 = ~n9268 ;
  assign y11054 = n20485 ;
  assign y11055 = n20491 ;
  assign y11056 = ~n20494 ;
  assign y11057 = ~n20500 ;
  assign y11058 = ~1'b0 ;
  assign y11059 = ~1'b0 ;
  assign y11060 = ~1'b0 ;
  assign y11061 = ~1'b0 ;
  assign y11062 = 1'b0 ;
  assign y11063 = n20501 ;
  assign y11064 = n4245 ;
  assign y11065 = ~1'b0 ;
  assign y11066 = ~1'b0 ;
  assign y11067 = ~1'b0 ;
  assign y11068 = ~n20503 ;
  assign y11069 = ~n20504 ;
  assign y11070 = n20507 ;
  assign y11071 = ~1'b0 ;
  assign y11072 = ~1'b0 ;
  assign y11073 = ~n20510 ;
  assign y11074 = ~n4939 ;
  assign y11075 = n20516 ;
  assign y11076 = ~1'b0 ;
  assign y11077 = 1'b0 ;
  assign y11078 = ~n20524 ;
  assign y11079 = ~n968 ;
  assign y11080 = ~1'b0 ;
  assign y11081 = n20526 ;
  assign y11082 = ~n20527 ;
  assign y11083 = n20528 ;
  assign y11084 = n20531 ;
  assign y11085 = n20537 ;
  assign y11086 = ~n20542 ;
  assign y11087 = n20543 ;
  assign y11088 = ~n20548 ;
  assign y11089 = ~n20552 ;
  assign y11090 = n20553 ;
  assign y11091 = n20557 ;
  assign y11092 = n20558 ;
  assign y11093 = n20562 ;
  assign y11094 = 1'b0 ;
  assign y11095 = ~1'b0 ;
  assign y11096 = ~n20563 ;
  assign y11097 = ~1'b0 ;
  assign y11098 = n20564 ;
  assign y11099 = ~n20566 ;
  assign y11100 = ~n20569 ;
  assign y11101 = n15316 ;
  assign y11102 = ~n20570 ;
  assign y11103 = ~n20572 ;
  assign y11104 = ~n20576 ;
  assign y11105 = ~1'b0 ;
  assign y11106 = ~n20580 ;
  assign y11107 = n5057 ;
  assign y11108 = ~1'b0 ;
  assign y11109 = ~1'b0 ;
  assign y11110 = ~n20582 ;
  assign y11111 = n20587 ;
  assign y11112 = ~n20588 ;
  assign y11113 = n20590 ;
  assign y11114 = ~n20591 ;
  assign y11115 = ~n20592 ;
  assign y11116 = ~1'b0 ;
  assign y11117 = n20594 ;
  assign y11118 = n13407 ;
  assign y11119 = ~1'b0 ;
  assign y11120 = ~1'b0 ;
  assign y11121 = ~1'b0 ;
  assign y11122 = n8101 ;
  assign y11123 = ~n20595 ;
  assign y11124 = n20596 ;
  assign y11125 = ~1'b0 ;
  assign y11126 = ~1'b0 ;
  assign y11127 = ~n20597 ;
  assign y11128 = n20602 ;
  assign y11129 = n20603 ;
  assign y11130 = n20605 ;
  assign y11131 = ~n20612 ;
  assign y11132 = ~n20613 ;
  assign y11133 = ~1'b0 ;
  assign y11134 = n20614 ;
  assign y11135 = ~n20615 ;
  assign y11136 = ~n20621 ;
  assign y11137 = ~1'b0 ;
  assign y11138 = n20623 ;
  assign y11139 = n20627 ;
  assign y11140 = ~n20630 ;
  assign y11141 = ~1'b0 ;
  assign y11142 = ~n20632 ;
  assign y11143 = 1'b0 ;
  assign y11144 = ~n20635 ;
  assign y11145 = n20637 ;
  assign y11146 = ~1'b0 ;
  assign y11147 = n20638 ;
  assign y11148 = ~n20639 ;
  assign y11149 = n20640 ;
  assign y11150 = ~n20641 ;
  assign y11151 = ~1'b0 ;
  assign y11152 = ~1'b0 ;
  assign y11153 = ~n20643 ;
  assign y11154 = ~n7933 ;
  assign y11155 = ~n20647 ;
  assign y11156 = ~1'b0 ;
  assign y11157 = ~n15938 ;
  assign y11158 = n20653 ;
  assign y11159 = n20655 ;
  assign y11160 = ~1'b0 ;
  assign y11161 = ~n20658 ;
  assign y11162 = ~1'b0 ;
  assign y11163 = n20671 ;
  assign y11164 = n20672 ;
  assign y11165 = ~1'b0 ;
  assign y11166 = ~1'b0 ;
  assign y11167 = ~n20673 ;
  assign y11168 = ~n20674 ;
  assign y11169 = ~n15934 ;
  assign y11170 = ~1'b0 ;
  assign y11171 = ~1'b0 ;
  assign y11172 = n6428 ;
  assign y11173 = ~n20675 ;
  assign y11174 = ~1'b0 ;
  assign y11175 = ~n20676 ;
  assign y11176 = ~1'b0 ;
  assign y11177 = ~n20679 ;
  assign y11178 = ~1'b0 ;
  assign y11179 = n20682 ;
  assign y11180 = n20686 ;
  assign y11181 = n20687 ;
  assign y11182 = n9945 ;
  assign y11183 = n20695 ;
  assign y11184 = ~1'b0 ;
  assign y11185 = ~n20699 ;
  assign y11186 = n20706 ;
  assign y11187 = ~n20713 ;
  assign y11188 = n20714 ;
  assign y11189 = ~1'b0 ;
  assign y11190 = n20718 ;
  assign y11191 = n20721 ;
  assign y11192 = ~1'b0 ;
  assign y11193 = ~1'b0 ;
  assign y11194 = ~1'b0 ;
  assign y11195 = n20728 ;
  assign y11196 = n20731 ;
  assign y11197 = n20735 ;
  assign y11198 = 1'b0 ;
  assign y11199 = ~1'b0 ;
  assign y11200 = ~n20738 ;
  assign y11201 = ~1'b0 ;
  assign y11202 = ~1'b0 ;
  assign y11203 = ~n20742 ;
  assign y11204 = ~n20745 ;
  assign y11205 = 1'b0 ;
  assign y11206 = ~1'b0 ;
  assign y11207 = 1'b0 ;
  assign y11208 = n20747 ;
  assign y11209 = n20751 ;
  assign y11210 = n20753 ;
  assign y11211 = n20756 ;
  assign y11212 = ~n20757 ;
  assign y11213 = ~1'b0 ;
  assign y11214 = 1'b0 ;
  assign y11215 = ~1'b0 ;
  assign y11216 = ~1'b0 ;
  assign y11217 = ~1'b0 ;
  assign y11218 = ~n20760 ;
  assign y11219 = ~1'b0 ;
  assign y11220 = ~n20761 ;
  assign y11221 = n20766 ;
  assign y11222 = ~n20768 ;
  assign y11223 = ~n20770 ;
  assign y11224 = n20773 ;
  assign y11225 = 1'b0 ;
  assign y11226 = n20774 ;
  assign y11227 = n20776 ;
  assign y11228 = n20780 ;
  assign y11229 = n20781 ;
  assign y11230 = n20783 ;
  assign y11231 = ~n20786 ;
  assign y11232 = ~1'b0 ;
  assign y11233 = 1'b0 ;
  assign y11234 = ~n20787 ;
  assign y11235 = ~n20788 ;
  assign y11236 = n20789 ;
  assign y11237 = ~n20463 ;
  assign y11238 = ~1'b0 ;
  assign y11239 = n15928 ;
  assign y11240 = ~n20791 ;
  assign y11241 = ~n20801 ;
  assign y11242 = ~n2186 ;
  assign y11243 = n20805 ;
  assign y11244 = ~n20806 ;
  assign y11245 = ~n8150 ;
  assign y11246 = ~n20816 ;
  assign y11247 = n20817 ;
  assign y11248 = ~n20819 ;
  assign y11249 = ~1'b0 ;
  assign y11250 = ~1'b0 ;
  assign y11251 = ~n20821 ;
  assign y11252 = ~n20823 ;
  assign y11253 = n7100 ;
  assign y11254 = ~n20826 ;
  assign y11255 = n20829 ;
  assign y11256 = ~1'b0 ;
  assign y11257 = ~n1434 ;
  assign y11258 = n20832 ;
  assign y11259 = ~n20833 ;
  assign y11260 = n20843 ;
  assign y11261 = ~n20844 ;
  assign y11262 = n20846 ;
  assign y11263 = ~1'b0 ;
  assign y11264 = ~n20848 ;
  assign y11265 = ~1'b0 ;
  assign y11266 = ~n20849 ;
  assign y11267 = ~1'b0 ;
  assign y11268 = ~n20851 ;
  assign y11269 = n20856 ;
  assign y11270 = ~1'b0 ;
  assign y11271 = ~n20862 ;
  assign y11272 = ~n20867 ;
  assign y11273 = ~1'b0 ;
  assign y11274 = n20874 ;
  assign y11275 = ~n20877 ;
  assign y11276 = n20879 ;
  assign y11277 = n20881 ;
  assign y11278 = 1'b0 ;
  assign y11279 = ~1'b0 ;
  assign y11280 = n20882 ;
  assign y11281 = ~1'b0 ;
  assign y11282 = ~1'b0 ;
  assign y11283 = n20901 ;
  assign y11284 = n20902 ;
  assign y11285 = ~1'b0 ;
  assign y11286 = ~1'b0 ;
  assign y11287 = ~n20906 ;
  assign y11288 = ~n20907 ;
  assign y11289 = n3820 ;
  assign y11290 = ~n20911 ;
  assign y11291 = ~n20912 ;
  assign y11292 = ~1'b0 ;
  assign y11293 = ~1'b0 ;
  assign y11294 = n20913 ;
  assign y11295 = ~n20915 ;
  assign y11296 = ~1'b0 ;
  assign y11297 = ~n20916 ;
  assign y11298 = n20922 ;
  assign y11299 = n2012 ;
  assign y11300 = ~n20923 ;
  assign y11301 = n20924 ;
  assign y11302 = ~1'b0 ;
  assign y11303 = ~1'b0 ;
  assign y11304 = ~n20927 ;
  assign y11305 = ~n20928 ;
  assign y11306 = ~n20931 ;
  assign y11307 = ~n20935 ;
  assign y11308 = ~1'b0 ;
  assign y11309 = n20940 ;
  assign y11310 = ~1'b0 ;
  assign y11311 = n20946 ;
  assign y11312 = n20947 ;
  assign y11313 = ~n20949 ;
  assign y11314 = ~n20951 ;
  assign y11315 = n20954 ;
  assign y11316 = ~1'b0 ;
  assign y11317 = ~n20957 ;
  assign y11318 = ~1'b0 ;
  assign y11319 = ~n20960 ;
  assign y11320 = n20961 ;
  assign y11321 = ~n20964 ;
  assign y11322 = n20967 ;
  assign y11323 = n5662 ;
  assign y11324 = ~n20970 ;
  assign y11325 = ~n20972 ;
  assign y11326 = ~1'b0 ;
  assign y11327 = n20982 ;
  assign y11328 = ~1'b0 ;
  assign y11329 = ~1'b0 ;
  assign y11330 = ~1'b0 ;
  assign y11331 = n20983 ;
  assign y11332 = ~n20984 ;
  assign y11333 = ~n20985 ;
  assign y11334 = n12790 ;
  assign y11335 = ~n15944 ;
  assign y11336 = n20988 ;
  assign y11337 = ~n20989 ;
  assign y11338 = ~1'b0 ;
  assign y11339 = ~n20994 ;
  assign y11340 = n20995 ;
  assign y11341 = n20998 ;
  assign y11342 = n21001 ;
  assign y11343 = ~1'b0 ;
  assign y11344 = ~1'b0 ;
  assign y11345 = ~1'b0 ;
  assign y11346 = ~n1539 ;
  assign y11347 = ~1'b0 ;
  assign y11348 = ~n21004 ;
  assign y11349 = n17095 ;
  assign y11350 = ~n21005 ;
  assign y11351 = ~n16314 ;
  assign y11352 = ~1'b0 ;
  assign y11353 = n21010 ;
  assign y11354 = ~n21011 ;
  assign y11355 = ~n21013 ;
  assign y11356 = ~1'b0 ;
  assign y11357 = n21019 ;
  assign y11358 = n21023 ;
  assign y11359 = ~n21024 ;
  assign y11360 = ~1'b0 ;
  assign y11361 = ~1'b0 ;
  assign y11362 = n21026 ;
  assign y11363 = ~1'b0 ;
  assign y11364 = ~n21027 ;
  assign y11365 = n21028 ;
  assign y11366 = ~n21034 ;
  assign y11367 = ~n21038 ;
  assign y11368 = ~n21047 ;
  assign y11369 = n21050 ;
  assign y11370 = ~n21058 ;
  assign y11371 = ~n21059 ;
  assign y11372 = ~n21062 ;
  assign y11373 = ~n21071 ;
  assign y11374 = ~1'b0 ;
  assign y11375 = ~n21076 ;
  assign y11376 = ~n21084 ;
  assign y11377 = n12513 ;
  assign y11378 = n21086 ;
  assign y11379 = ~1'b0 ;
  assign y11380 = ~1'b0 ;
  assign y11381 = n21089 ;
  assign y11382 = n19360 ;
  assign y11383 = n21092 ;
  assign y11384 = n21095 ;
  assign y11385 = n21102 ;
  assign y11386 = ~n20617 ;
  assign y11387 = n21104 ;
  assign y11388 = ~n21108 ;
  assign y11389 = ~1'b0 ;
  assign y11390 = n21109 ;
  assign y11391 = ~1'b0 ;
  assign y11392 = ~n21114 ;
  assign y11393 = n21115 ;
  assign y11394 = n21116 ;
  assign y11395 = n21117 ;
  assign y11396 = ~1'b0 ;
  assign y11397 = n12897 ;
  assign y11398 = ~1'b0 ;
  assign y11399 = ~1'b0 ;
  assign y11400 = n21119 ;
  assign y11401 = n21121 ;
  assign y11402 = n21126 ;
  assign y11403 = ~n8503 ;
  assign y11404 = ~1'b0 ;
  assign y11405 = ~n21129 ;
  assign y11406 = ~n21131 ;
  assign y11407 = 1'b0 ;
  assign y11408 = n21133 ;
  assign y11409 = n21134 ;
  assign y11410 = ~1'b0 ;
  assign y11411 = ~n21137 ;
  assign y11412 = ~1'b0 ;
  assign y11413 = ~1'b0 ;
  assign y11414 = ~n21139 ;
  assign y11415 = ~1'b0 ;
  assign y11416 = 1'b0 ;
  assign y11417 = ~1'b0 ;
  assign y11418 = ~1'b0 ;
  assign y11419 = n21142 ;
  assign y11420 = ~1'b0 ;
  assign y11421 = ~n21144 ;
  assign y11422 = ~n21145 ;
  assign y11423 = ~1'b0 ;
  assign y11424 = ~1'b0 ;
  assign y11425 = ~n21148 ;
  assign y11426 = ~1'b0 ;
  assign y11427 = ~n21149 ;
  assign y11428 = ~1'b0 ;
  assign y11429 = n21151 ;
  assign y11430 = n21153 ;
  assign y11431 = ~n16394 ;
  assign y11432 = n20974 ;
  assign y11433 = 1'b0 ;
  assign y11434 = ~1'b0 ;
  assign y11435 = ~1'b0 ;
  assign y11436 = ~1'b0 ;
  assign y11437 = ~n21154 ;
  assign y11438 = ~n21158 ;
  assign y11439 = n21160 ;
  assign y11440 = ~1'b0 ;
  assign y11441 = ~1'b0 ;
  assign y11442 = n21162 ;
  assign y11443 = ~1'b0 ;
  assign y11444 = ~1'b0 ;
  assign y11445 = ~1'b0 ;
  assign y11446 = ~n21166 ;
  assign y11447 = ~1'b0 ;
  assign y11448 = n21174 ;
  assign y11449 = ~1'b0 ;
  assign y11450 = ~1'b0 ;
  assign y11451 = n21175 ;
  assign y11452 = ~1'b0 ;
  assign y11453 = ~n3833 ;
  assign y11454 = ~1'b0 ;
  assign y11455 = ~n21179 ;
  assign y11456 = ~1'b0 ;
  assign y11457 = ~1'b0 ;
  assign y11458 = ~n21181 ;
  assign y11459 = ~n21182 ;
  assign y11460 = n21191 ;
  assign y11461 = n1346 ;
  assign y11462 = ~n21194 ;
  assign y11463 = n8773 ;
  assign y11464 = ~n10513 ;
  assign y11465 = n2231 ;
  assign y11466 = n21195 ;
  assign y11467 = n21201 ;
  assign y11468 = 1'b0 ;
  assign y11469 = n21203 ;
  assign y11470 = n21204 ;
  assign y11471 = ~1'b0 ;
  assign y11472 = ~1'b0 ;
  assign y11473 = ~1'b0 ;
  assign y11474 = ~n21207 ;
  assign y11475 = n21208 ;
  assign y11476 = n21209 ;
  assign y11477 = n105 ;
  assign y11478 = ~n21210 ;
  assign y11479 = ~1'b0 ;
  assign y11480 = n21214 ;
  assign y11481 = ~1'b0 ;
  assign y11482 = ~n21215 ;
  assign y11483 = n21216 ;
  assign y11484 = ~1'b0 ;
  assign y11485 = ~1'b0 ;
  assign y11486 = ~n21218 ;
  assign y11487 = n21219 ;
  assign y11488 = ~1'b0 ;
  assign y11489 = n21223 ;
  assign y11490 = ~1'b0 ;
  assign y11491 = ~n21225 ;
  assign y11492 = ~n21226 ;
  assign y11493 = n21227 ;
  assign y11494 = n21233 ;
  assign y11495 = ~1'b0 ;
  assign y11496 = n21235 ;
  assign y11497 = ~1'b0 ;
  assign y11498 = 1'b0 ;
  assign y11499 = n21236 ;
  assign y11500 = n21242 ;
  assign y11501 = n21243 ;
  assign y11502 = ~n21244 ;
  assign y11503 = ~1'b0 ;
  assign y11504 = ~n21246 ;
  assign y11505 = ~1'b0 ;
  assign y11506 = ~n21250 ;
  assign y11507 = ~n21254 ;
  assign y11508 = ~1'b0 ;
  assign y11509 = n9290 ;
  assign y11510 = n5106 ;
  assign y11511 = n21257 ;
  assign y11512 = ~1'b0 ;
  assign y11513 = n21263 ;
  assign y11514 = ~1'b0 ;
  assign y11515 = ~1'b0 ;
  assign y11516 = ~n21266 ;
  assign y11517 = ~1'b0 ;
  assign y11518 = ~n21268 ;
  assign y11519 = ~1'b0 ;
  assign y11520 = ~1'b0 ;
  assign y11521 = ~1'b0 ;
  assign y11522 = ~n3235 ;
  assign y11523 = ~n21269 ;
  assign y11524 = ~n21272 ;
  assign y11525 = ~1'b0 ;
  assign y11526 = n21274 ;
  assign y11527 = ~1'b0 ;
  assign y11528 = ~n21276 ;
  assign y11529 = n21281 ;
  assign y11530 = ~n21284 ;
  assign y11531 = ~1'b0 ;
  assign y11532 = ~1'b0 ;
  assign y11533 = n21285 ;
  assign y11534 = ~1'b0 ;
  assign y11535 = n10958 ;
  assign y11536 = n21286 ;
  assign y11537 = ~1'b0 ;
  assign y11538 = n3315 ;
  assign y11539 = ~1'b0 ;
  assign y11540 = ~n21292 ;
  assign y11541 = n21294 ;
  assign y11542 = ~1'b0 ;
  assign y11543 = n21295 ;
  assign y11544 = ~1'b0 ;
  assign y11545 = n21297 ;
  assign y11546 = n21298 ;
  assign y11547 = n21299 ;
  assign y11548 = ~1'b0 ;
  assign y11549 = ~n21300 ;
  assign y11550 = n21301 ;
  assign y11551 = ~n21305 ;
  assign y11552 = ~n9240 ;
  assign y11553 = 1'b0 ;
  assign y11554 = n21306 ;
  assign y11555 = ~1'b0 ;
  assign y11556 = ~n21307 ;
  assign y11557 = ~n21311 ;
  assign y11558 = ~1'b0 ;
  assign y11559 = ~1'b0 ;
  assign y11560 = ~1'b0 ;
  assign y11561 = ~n21321 ;
  assign y11562 = 1'b0 ;
  assign y11563 = ~1'b0 ;
  assign y11564 = ~n21323 ;
  assign y11565 = ~1'b0 ;
  assign y11566 = ~1'b0 ;
  assign y11567 = ~1'b0 ;
  assign y11568 = ~1'b0 ;
  assign y11569 = ~1'b0 ;
  assign y11570 = ~n21328 ;
  assign y11571 = ~n21330 ;
  assign y11572 = ~n21343 ;
  assign y11573 = ~n21346 ;
  assign y11574 = ~1'b0 ;
  assign y11575 = n21347 ;
  assign y11576 = 1'b0 ;
  assign y11577 = ~n21351 ;
  assign y11578 = n8010 ;
  assign y11579 = 1'b0 ;
  assign y11580 = ~n21357 ;
  assign y11581 = n21365 ;
  assign y11582 = ~1'b0 ;
  assign y11583 = ~n21368 ;
  assign y11584 = n21369 ;
  assign y11585 = n5933 ;
  assign y11586 = n21375 ;
  assign y11587 = n21376 ;
  assign y11588 = ~1'b0 ;
  assign y11589 = ~n21379 ;
  assign y11590 = ~n21381 ;
  assign y11591 = n21383 ;
  assign y11592 = n3351 ;
  assign y11593 = n15719 ;
  assign y11594 = n21388 ;
  assign y11595 = ~n21389 ;
  assign y11596 = ~n21397 ;
  assign y11597 = n21400 ;
  assign y11598 = n21404 ;
  assign y11599 = ~1'b0 ;
  assign y11600 = ~1'b0 ;
  assign y11601 = ~n21408 ;
  assign y11602 = ~n21409 ;
  assign y11603 = ~n21412 ;
  assign y11604 = n10162 ;
  assign y11605 = n21413 ;
  assign y11606 = 1'b0 ;
  assign y11607 = n21414 ;
  assign y11608 = n21416 ;
  assign y11609 = n21417 ;
  assign y11610 = ~n21420 ;
  assign y11611 = n21422 ;
  assign y11612 = n21424 ;
  assign y11613 = n21426 ;
  assign y11614 = ~n1553 ;
  assign y11615 = ~1'b0 ;
  assign y11616 = ~n21431 ;
  assign y11617 = ~n21435 ;
  assign y11618 = n21438 ;
  assign y11619 = 1'b0 ;
  assign y11620 = n21439 ;
  assign y11621 = ~n21440 ;
  assign y11622 = ~n21443 ;
  assign y11623 = ~n21453 ;
  assign y11624 = ~n21454 ;
  assign y11625 = n21457 ;
  assign y11626 = ~n21464 ;
  assign y11627 = n21467 ;
  assign y11628 = n21469 ;
  assign y11629 = ~n21470 ;
  assign y11630 = n13953 ;
  assign y11631 = n21472 ;
  assign y11632 = ~n21474 ;
  assign y11633 = n21476 ;
  assign y11634 = ~n21482 ;
  assign y11635 = ~n21484 ;
  assign y11636 = n21485 ;
  assign y11637 = n21486 ;
  assign y11638 = ~1'b0 ;
  assign y11639 = ~1'b0 ;
  assign y11640 = n21487 ;
  assign y11641 = n21488 ;
  assign y11642 = ~1'b0 ;
  assign y11643 = ~n21489 ;
  assign y11644 = n21491 ;
  assign y11645 = n21495 ;
  assign y11646 = ~1'b0 ;
  assign y11647 = n21499 ;
  assign y11648 = ~n21501 ;
  assign y11649 = n21502 ;
  assign y11650 = ~n21505 ;
  assign y11651 = ~1'b0 ;
  assign y11652 = n21506 ;
  assign y11653 = ~1'b0 ;
  assign y11654 = ~n21508 ;
  assign y11655 = ~1'b0 ;
  assign y11656 = ~n21509 ;
  assign y11657 = n21511 ;
  assign y11658 = n21512 ;
  assign y11659 = ~n21514 ;
  assign y11660 = ~1'b0 ;
  assign y11661 = ~1'b0 ;
  assign y11662 = ~n21522 ;
  assign y11663 = ~n21525 ;
  assign y11664 = ~1'b0 ;
  assign y11665 = n21527 ;
  assign y11666 = ~n21529 ;
  assign y11667 = ~n21539 ;
  assign y11668 = n21542 ;
  assign y11669 = ~1'b0 ;
  assign y11670 = ~n21544 ;
  assign y11671 = ~n21546 ;
  assign y11672 = ~n21551 ;
  assign y11673 = ~1'b0 ;
  assign y11674 = ~1'b0 ;
  assign y11675 = n21552 ;
  assign y11676 = ~n21554 ;
  assign y11677 = ~n21556 ;
  assign y11678 = n21560 ;
  assign y11679 = ~1'b0 ;
  assign y11680 = n11001 ;
  assign y11681 = ~n21562 ;
  assign y11682 = ~n21571 ;
  assign y11683 = ~n21576 ;
  assign y11684 = n21581 ;
  assign y11685 = n21582 ;
  assign y11686 = ~n7109 ;
  assign y11687 = ~n21584 ;
  assign y11688 = n20031 ;
  assign y11689 = ~1'b0 ;
  assign y11690 = ~n21587 ;
  assign y11691 = ~n21592 ;
  assign y11692 = ~1'b0 ;
  assign y11693 = ~n21594 ;
  assign y11694 = n21596 ;
  assign y11695 = ~1'b0 ;
  assign y11696 = n21599 ;
  assign y11697 = ~1'b0 ;
  assign y11698 = ~1'b0 ;
  assign y11699 = ~n21600 ;
  assign y11700 = n21602 ;
  assign y11701 = n9542 ;
  assign y11702 = ~n17493 ;
  assign y11703 = ~n18875 ;
  assign y11704 = ~1'b0 ;
  assign y11705 = ~n21604 ;
  assign y11706 = ~n21607 ;
  assign y11707 = ~1'b0 ;
  assign y11708 = 1'b0 ;
  assign y11709 = ~n21608 ;
  assign y11710 = ~1'b0 ;
  assign y11711 = n21612 ;
  assign y11712 = ~n4039 ;
  assign y11713 = n620 ;
  assign y11714 = ~1'b0 ;
  assign y11715 = ~1'b0 ;
  assign y11716 = n21617 ;
  assign y11717 = ~n21624 ;
  assign y11718 = ~1'b0 ;
  assign y11719 = n21626 ;
  assign y11720 = ~n21628 ;
  assign y11721 = ~1'b0 ;
  assign y11722 = ~1'b0 ;
  assign y11723 = ~n21632 ;
  assign y11724 = ~n7209 ;
  assign y11725 = ~n21637 ;
  assign y11726 = n21638 ;
  assign y11727 = n21641 ;
  assign y11728 = ~n21643 ;
  assign y11729 = n21644 ;
  assign y11730 = ~1'b0 ;
  assign y11731 = ~n21652 ;
  assign y11732 = n21655 ;
  assign y11733 = ~n21659 ;
  assign y11734 = ~1'b0 ;
  assign y11735 = ~n21662 ;
  assign y11736 = ~1'b0 ;
  assign y11737 = ~n21665 ;
  assign y11738 = n21668 ;
  assign y11739 = ~n21670 ;
  assign y11740 = ~1'b0 ;
  assign y11741 = ~n21672 ;
  assign y11742 = ~n21675 ;
  assign y11743 = n21678 ;
  assign y11744 = ~1'b0 ;
  assign y11745 = ~n21680 ;
  assign y11746 = ~n21681 ;
  assign y11747 = n21683 ;
  assign y11748 = ~n21685 ;
  assign y11749 = ~1'b0 ;
  assign y11750 = n21690 ;
  assign y11751 = ~n21701 ;
  assign y11752 = n21702 ;
  assign y11753 = n21704 ;
  assign y11754 = n21705 ;
  assign y11755 = ~n15226 ;
  assign y11756 = ~n21707 ;
  assign y11757 = ~n21711 ;
  assign y11758 = ~n21716 ;
  assign y11759 = ~n21719 ;
  assign y11760 = ~1'b0 ;
  assign y11761 = ~1'b0 ;
  assign y11762 = ~1'b0 ;
  assign y11763 = ~1'b0 ;
  assign y11764 = ~n21725 ;
  assign y11765 = ~n21727 ;
  assign y11766 = n21730 ;
  assign y11767 = ~n21731 ;
  assign y11768 = ~1'b0 ;
  assign y11769 = n21735 ;
  assign y11770 = ~n21738 ;
  assign y11771 = ~n21743 ;
  assign y11772 = ~n21744 ;
  assign y11773 = ~1'b0 ;
  assign y11774 = ~n21746 ;
  assign y11775 = n21747 ;
  assign y11776 = ~n21749 ;
  assign y11777 = ~n21757 ;
  assign y11778 = ~1'b0 ;
  assign y11779 = ~n21758 ;
  assign y11780 = ~n21761 ;
  assign y11781 = ~1'b0 ;
  assign y11782 = ~n2080 ;
  assign y11783 = ~1'b0 ;
  assign y11784 = ~n21772 ;
  assign y11785 = n21777 ;
  assign y11786 = ~n21778 ;
  assign y11787 = n7825 ;
  assign y11788 = ~n21779 ;
  assign y11789 = ~n21780 ;
  assign y11790 = ~1'b0 ;
  assign y11791 = ~n21781 ;
  assign y11792 = ~n21782 ;
  assign y11793 = n11055 ;
  assign y11794 = ~1'b0 ;
  assign y11795 = ~1'b0 ;
  assign y11796 = ~1'b0 ;
  assign y11797 = n21789 ;
  assign y11798 = ~1'b0 ;
  assign y11799 = n21791 ;
  assign y11800 = ~n21794 ;
  assign y11801 = n21797 ;
  assign y11802 = n21798 ;
  assign y11803 = ~1'b0 ;
  assign y11804 = ~1'b0 ;
  assign y11805 = ~n21800 ;
  assign y11806 = ~1'b0 ;
  assign y11807 = ~1'b0 ;
  assign y11808 = n21801 ;
  assign y11809 = ~1'b0 ;
  assign y11810 = ~1'b0 ;
  assign y11811 = ~1'b0 ;
  assign y11812 = ~n21802 ;
  assign y11813 = ~n17281 ;
  assign y11814 = ~n21804 ;
  assign y11815 = 1'b0 ;
  assign y11816 = n21805 ;
  assign y11817 = ~1'b0 ;
  assign y11818 = n21806 ;
  assign y11819 = n21809 ;
  assign y11820 = ~1'b0 ;
  assign y11821 = ~n21812 ;
  assign y11822 = n21818 ;
  assign y11823 = ~1'b0 ;
  assign y11824 = n21819 ;
  assign y11825 = ~1'b0 ;
  assign y11826 = ~n21820 ;
  assign y11827 = ~n21821 ;
  assign y11828 = n21822 ;
  assign y11829 = n21825 ;
  assign y11830 = ~1'b0 ;
  assign y11831 = ~n21826 ;
  assign y11832 = ~n21830 ;
  assign y11833 = ~1'b0 ;
  assign y11834 = ~n21834 ;
  assign y11835 = ~1'b0 ;
  assign y11836 = n21844 ;
  assign y11837 = ~n1325 ;
  assign y11838 = ~1'b0 ;
  assign y11839 = n21846 ;
  assign y11840 = n21848 ;
  assign y11841 = ~1'b0 ;
  assign y11842 = n21852 ;
  assign y11843 = ~1'b0 ;
  assign y11844 = n21853 ;
  assign y11845 = n21855 ;
  assign y11846 = ~1'b0 ;
  assign y11847 = ~n8881 ;
  assign y11848 = ~n21861 ;
  assign y11849 = ~1'b0 ;
  assign y11850 = ~1'b0 ;
  assign y11851 = ~n21869 ;
  assign y11852 = ~1'b0 ;
  assign y11853 = ~n21872 ;
  assign y11854 = ~n21874 ;
  assign y11855 = ~1'b0 ;
  assign y11856 = ~n21875 ;
  assign y11857 = ~n21878 ;
  assign y11858 = ~n21881 ;
  assign y11859 = n21882 ;
  assign y11860 = n11662 ;
  assign y11861 = ~1'b0 ;
  assign y11862 = n21883 ;
  assign y11863 = n6527 ;
  assign y11864 = ~n21885 ;
  assign y11865 = ~1'b0 ;
  assign y11866 = ~n19818 ;
  assign y11867 = ~1'b0 ;
  assign y11868 = n21886 ;
  assign y11869 = ~1'b0 ;
  assign y11870 = n21889 ;
  assign y11871 = ~1'b0 ;
  assign y11872 = n21890 ;
  assign y11873 = n21892 ;
  assign y11874 = ~n21893 ;
  assign y11875 = ~1'b0 ;
  assign y11876 = n21894 ;
  assign y11877 = ~1'b0 ;
  assign y11878 = ~n21896 ;
  assign y11879 = ~n21897 ;
  assign y11880 = ~1'b0 ;
  assign y11881 = ~n21899 ;
  assign y11882 = ~1'b0 ;
  assign y11883 = n21900 ;
  assign y11884 = n18740 ;
  assign y11885 = ~n21905 ;
  assign y11886 = n21909 ;
  assign y11887 = n21911 ;
  assign y11888 = ~1'b0 ;
  assign y11889 = n11477 ;
  assign y11890 = ~n21912 ;
  assign y11891 = n21913 ;
  assign y11892 = n21923 ;
  assign y11893 = ~1'b0 ;
  assign y11894 = ~1'b0 ;
  assign y11895 = n21931 ;
  assign y11896 = ~1'b0 ;
  assign y11897 = ~1'b0 ;
  assign y11898 = n21932 ;
  assign y11899 = ~n21938 ;
  assign y11900 = n21940 ;
  assign y11901 = n21944 ;
  assign y11902 = ~1'b0 ;
  assign y11903 = n21950 ;
  assign y11904 = ~1'b0 ;
  assign y11905 = n21952 ;
  assign y11906 = ~n21953 ;
  assign y11907 = ~1'b0 ;
  assign y11908 = ~n21960 ;
  assign y11909 = ~1'b0 ;
  assign y11910 = n21962 ;
  assign y11911 = ~1'b0 ;
  assign y11912 = n21964 ;
  assign y11913 = ~n21965 ;
  assign y11914 = ~n21969 ;
  assign y11915 = n21970 ;
  assign y11916 = ~n21980 ;
  assign y11917 = ~n21984 ;
  assign y11918 = ~n12799 ;
  assign y11919 = n21985 ;
  assign y11920 = n21987 ;
  assign y11921 = ~1'b0 ;
  assign y11922 = ~n21989 ;
  assign y11923 = ~1'b0 ;
  assign y11924 = n21990 ;
  assign y11925 = n2415 ;
  assign y11926 = ~n21992 ;
  assign y11927 = ~n21993 ;
  assign y11928 = ~1'b0 ;
  assign y11929 = n21995 ;
  assign y11930 = ~n22000 ;
  assign y11931 = ~1'b0 ;
  assign y11932 = ~1'b0 ;
  assign y11933 = n22001 ;
  assign y11934 = ~n22002 ;
  assign y11935 = ~1'b0 ;
  assign y11936 = ~n5911 ;
  assign y11937 = ~n22004 ;
  assign y11938 = ~n22009 ;
  assign y11939 = ~1'b0 ;
  assign y11940 = ~1'b0 ;
  assign y11941 = ~n22015 ;
  assign y11942 = ~n3713 ;
  assign y11943 = n22021 ;
  assign y11944 = n22027 ;
  assign y11945 = ~1'b0 ;
  assign y11946 = n22028 ;
  assign y11947 = ~1'b0 ;
  assign y11948 = ~n22031 ;
  assign y11949 = n17065 ;
  assign y11950 = ~n20992 ;
  assign y11951 = ~n22033 ;
  assign y11952 = ~1'b0 ;
  assign y11953 = ~1'b0 ;
  assign y11954 = ~1'b0 ;
  assign y11955 = ~1'b0 ;
  assign y11956 = ~1'b0 ;
  assign y11957 = ~n22034 ;
  assign y11958 = ~n22036 ;
  assign y11959 = ~1'b0 ;
  assign y11960 = ~1'b0 ;
  assign y11961 = ~1'b0 ;
  assign y11962 = ~1'b0 ;
  assign y11963 = n22037 ;
  assign y11964 = ~n22039 ;
  assign y11965 = ~1'b0 ;
  assign y11966 = ~1'b0 ;
  assign y11967 = n22040 ;
  assign y11968 = ~1'b0 ;
  assign y11969 = ~n22041 ;
  assign y11970 = ~n22047 ;
  assign y11971 = n22048 ;
  assign y11972 = n22050 ;
  assign y11973 = ~1'b0 ;
  assign y11974 = n22051 ;
  assign y11975 = n12363 ;
  assign y11976 = ~n22054 ;
  assign y11977 = n22063 ;
  assign y11978 = ~n22068 ;
  assign y11979 = n22070 ;
  assign y11980 = ~1'b0 ;
  assign y11981 = 1'b0 ;
  assign y11982 = n22077 ;
  assign y11983 = n22081 ;
  assign y11984 = ~n22086 ;
  assign y11985 = ~1'b0 ;
  assign y11986 = ~1'b0 ;
  assign y11987 = ~1'b0 ;
  assign y11988 = n22090 ;
  assign y11989 = ~1'b0 ;
  assign y11990 = ~n22091 ;
  assign y11991 = n6472 ;
  assign y11992 = ~1'b0 ;
  assign y11993 = ~n22095 ;
  assign y11994 = n22097 ;
  assign y11995 = ~1'b0 ;
  assign y11996 = n22098 ;
  assign y11997 = 1'b0 ;
  assign y11998 = n22099 ;
  assign y11999 = ~1'b0 ;
  assign y12000 = ~n22102 ;
  assign y12001 = 1'b0 ;
  assign y12002 = n22105 ;
  assign y12003 = n22106 ;
  assign y12004 = n22108 ;
  assign y12005 = ~1'b0 ;
  assign y12006 = n22110 ;
  assign y12007 = n22114 ;
  assign y12008 = ~1'b0 ;
  assign y12009 = 1'b0 ;
  assign y12010 = n22115 ;
  assign y12011 = ~1'b0 ;
  assign y12012 = ~n22119 ;
  assign y12013 = n22121 ;
  assign y12014 = ~n22123 ;
  assign y12015 = ~n22124 ;
  assign y12016 = ~1'b0 ;
  assign y12017 = ~n22127 ;
  assign y12018 = ~n1592 ;
  assign y12019 = ~n22128 ;
  assign y12020 = ~1'b0 ;
  assign y12021 = n22134 ;
  assign y12022 = n22138 ;
  assign y12023 = ~n22140 ;
  assign y12024 = ~n22141 ;
  assign y12025 = ~1'b0 ;
  assign y12026 = ~1'b0 ;
  assign y12027 = n22143 ;
  assign y12028 = n22144 ;
  assign y12029 = ~n22152 ;
  assign y12030 = ~1'b0 ;
  assign y12031 = n22156 ;
  assign y12032 = ~1'b0 ;
  assign y12033 = ~n22163 ;
  assign y12034 = n22175 ;
  assign y12035 = n22179 ;
  assign y12036 = ~n3772 ;
  assign y12037 = ~n22180 ;
  assign y12038 = ~1'b0 ;
  assign y12039 = ~1'b0 ;
  assign y12040 = n22181 ;
  assign y12041 = n22182 ;
  assign y12042 = n22183 ;
  assign y12043 = ~1'b0 ;
  assign y12044 = n22184 ;
  assign y12045 = n22187 ;
  assign y12046 = ~n22189 ;
  assign y12047 = ~1'b0 ;
  assign y12048 = n2661 ;
  assign y12049 = ~n22190 ;
  assign y12050 = ~n2610 ;
  assign y12051 = ~1'b0 ;
  assign y12052 = ~1'b0 ;
  assign y12053 = ~1'b0 ;
  assign y12054 = ~1'b0 ;
  assign y12055 = n22194 ;
  assign y12056 = n695 ;
  assign y12057 = ~1'b0 ;
  assign y12058 = ~n22199 ;
  assign y12059 = ~1'b0 ;
  assign y12060 = ~1'b0 ;
  assign y12061 = n162 ;
  assign y12062 = n22202 ;
  assign y12063 = ~1'b0 ;
  assign y12064 = n22204 ;
  assign y12065 = 1'b0 ;
  assign y12066 = ~n22205 ;
  assign y12067 = ~1'b0 ;
  assign y12068 = n22206 ;
  assign y12069 = ~1'b0 ;
  assign y12070 = ~1'b0 ;
  assign y12071 = ~n22207 ;
  assign y12072 = ~1'b0 ;
  assign y12073 = n22211 ;
  assign y12074 = n22212 ;
  assign y12075 = ~1'b0 ;
  assign y12076 = ~1'b0 ;
  assign y12077 = 1'b0 ;
  assign y12078 = 1'b0 ;
  assign y12079 = ~1'b0 ;
  assign y12080 = ~n22216 ;
  assign y12081 = ~n22230 ;
  assign y12082 = ~n22233 ;
  assign y12083 = n22235 ;
  assign y12084 = n22236 ;
  assign y12085 = ~n13601 ;
  assign y12086 = ~n22237 ;
  assign y12087 = ~1'b0 ;
  assign y12088 = 1'b0 ;
  assign y12089 = n7512 ;
  assign y12090 = ~n22240 ;
  assign y12091 = ~1'b0 ;
  assign y12092 = n22243 ;
  assign y12093 = n22248 ;
  assign y12094 = ~n22249 ;
  assign y12095 = ~n22250 ;
  assign y12096 = n22254 ;
  assign y12097 = ~1'b0 ;
  assign y12098 = n22256 ;
  assign y12099 = ~1'b0 ;
  assign y12100 = ~1'b0 ;
  assign y12101 = ~n22259 ;
  assign y12102 = ~1'b0 ;
  assign y12103 = n22260 ;
  assign y12104 = ~n557 ;
  assign y12105 = ~n22261 ;
  assign y12106 = n22265 ;
  assign y12107 = ~1'b0 ;
  assign y12108 = n7265 ;
  assign y12109 = ~n22266 ;
  assign y12110 = n1749 ;
  assign y12111 = n22267 ;
  assign y12112 = ~1'b0 ;
  assign y12113 = ~n22269 ;
  assign y12114 = ~1'b0 ;
  assign y12115 = ~n22271 ;
  assign y12116 = ~n22277 ;
  assign y12117 = n22278 ;
  assign y12118 = ~n22279 ;
  assign y12119 = ~1'b0 ;
  assign y12120 = ~n22281 ;
  assign y12121 = ~n22284 ;
  assign y12122 = ~n22285 ;
  assign y12123 = ~1'b0 ;
  assign y12124 = ~n16847 ;
  assign y12125 = ~1'b0 ;
  assign y12126 = ~1'b0 ;
  assign y12127 = ~n22291 ;
  assign y12128 = ~1'b0 ;
  assign y12129 = ~n22299 ;
  assign y12130 = n22302 ;
  assign y12131 = ~n22303 ;
  assign y12132 = ~1'b0 ;
  assign y12133 = n22305 ;
  assign y12134 = ~n22310 ;
  assign y12135 = ~n22312 ;
  assign y12136 = ~1'b0 ;
  assign y12137 = ~1'b0 ;
  assign y12138 = ~n22316 ;
  assign y12139 = ~1'b0 ;
  assign y12140 = ~n22318 ;
  assign y12141 = n22319 ;
  assign y12142 = ~n22321 ;
  assign y12143 = ~1'b0 ;
  assign y12144 = ~n22323 ;
  assign y12145 = ~n22328 ;
  assign y12146 = n22335 ;
  assign y12147 = ~n22338 ;
  assign y12148 = n19769 ;
  assign y12149 = ~1'b0 ;
  assign y12150 = ~1'b0 ;
  assign y12151 = ~n22342 ;
  assign y12152 = ~1'b0 ;
  assign y12153 = ~n22343 ;
  assign y12154 = ~1'b0 ;
  assign y12155 = n22350 ;
  assign y12156 = ~n22351 ;
  assign y12157 = n22354 ;
  assign y12158 = n22357 ;
  assign y12159 = ~1'b0 ;
  assign y12160 = n22358 ;
  assign y12161 = ~1'b0 ;
  assign y12162 = ~1'b0 ;
  assign y12163 = n22360 ;
  assign y12164 = ~1'b0 ;
  assign y12165 = ~n22362 ;
  assign y12166 = n22366 ;
  assign y12167 = ~n22372 ;
  assign y12168 = n22374 ;
  assign y12169 = n22377 ;
  assign y12170 = ~n22381 ;
  assign y12171 = n19446 ;
  assign y12172 = ~n22393 ;
  assign y12173 = ~n22394 ;
  assign y12174 = n21892 ;
  assign y12175 = ~n22395 ;
  assign y12176 = n22397 ;
  assign y12177 = n22398 ;
  assign y12178 = ~n22401 ;
  assign y12179 = n22405 ;
  assign y12180 = n22406 ;
  assign y12181 = ~1'b0 ;
  assign y12182 = n22409 ;
  assign y12183 = n5916 ;
  assign y12184 = ~n22411 ;
  assign y12185 = ~1'b0 ;
  assign y12186 = n22412 ;
  assign y12187 = n6535 ;
  assign y12188 = ~1'b0 ;
  assign y12189 = ~1'b0 ;
  assign y12190 = ~n22413 ;
  assign y12191 = n22415 ;
  assign y12192 = ~n22416 ;
  assign y12193 = ~1'b0 ;
  assign y12194 = n22417 ;
  assign y12195 = n22420 ;
  assign y12196 = n22424 ;
  assign y12197 = ~1'b0 ;
  assign y12198 = ~n22430 ;
  assign y12199 = ~1'b0 ;
  assign y12200 = n22431 ;
  assign y12201 = 1'b0 ;
  assign y12202 = ~n22433 ;
  assign y12203 = n22447 ;
  assign y12204 = n22450 ;
  assign y12205 = ~n22451 ;
  assign y12206 = ~n22453 ;
  assign y12207 = ~n22456 ;
  assign y12208 = ~n22465 ;
  assign y12209 = n22466 ;
  assign y12210 = ~n11069 ;
  assign y12211 = ~1'b0 ;
  assign y12212 = ~1'b0 ;
  assign y12213 = n22471 ;
  assign y12214 = ~n22474 ;
  assign y12215 = ~n22476 ;
  assign y12216 = ~n22478 ;
  assign y12217 = ~1'b0 ;
  assign y12218 = n22482 ;
  assign y12219 = ~n22484 ;
  assign y12220 = n22486 ;
  assign y12221 = ~1'b0 ;
  assign y12222 = ~n22488 ;
  assign y12223 = ~n22495 ;
  assign y12224 = ~1'b0 ;
  assign y12225 = n22497 ;
  assign y12226 = n21269 ;
  assign y12227 = ~n22501 ;
  assign y12228 = ~1'b0 ;
  assign y12229 = n22504 ;
  assign y12230 = n22509 ;
  assign y12231 = ~n22511 ;
  assign y12232 = ~n22514 ;
  assign y12233 = ~1'b0 ;
  assign y12234 = ~1'b0 ;
  assign y12235 = ~n22515 ;
  assign y12236 = ~n22516 ;
  assign y12237 = n22517 ;
  assign y12238 = ~1'b0 ;
  assign y12239 = ~1'b0 ;
  assign y12240 = ~n22522 ;
  assign y12241 = ~n22523 ;
  assign y12242 = n22525 ;
  assign y12243 = ~1'b0 ;
  assign y12244 = n22530 ;
  assign y12245 = ~1'b0 ;
  assign y12246 = ~n22533 ;
  assign y12247 = ~n13218 ;
  assign y12248 = ~1'b0 ;
  assign y12249 = ~1'b0 ;
  assign y12250 = n5562 ;
  assign y12251 = ~n22535 ;
  assign y12252 = n22537 ;
  assign y12253 = ~1'b0 ;
  assign y12254 = ~n22540 ;
  assign y12255 = n6023 ;
  assign y12256 = ~1'b0 ;
  assign y12257 = ~n22543 ;
  assign y12258 = ~n22547 ;
  assign y12259 = ~n22549 ;
  assign y12260 = n22553 ;
  assign y12261 = ~n22560 ;
  assign y12262 = ~1'b0 ;
  assign y12263 = ~n22564 ;
  assign y12264 = n22572 ;
  assign y12265 = n22576 ;
  assign y12266 = n22579 ;
  assign y12267 = ~1'b0 ;
  assign y12268 = ~1'b0 ;
  assign y12269 = n22580 ;
  assign y12270 = n22584 ;
  assign y12271 = ~1'b0 ;
  assign y12272 = n22588 ;
  assign y12273 = ~n22590 ;
  assign y12274 = n22593 ;
  assign y12275 = n22594 ;
  assign y12276 = ~1'b0 ;
  assign y12277 = ~n13399 ;
  assign y12278 = ~n22597 ;
  assign y12279 = ~1'b0 ;
  assign y12280 = n22604 ;
  assign y12281 = n22606 ;
  assign y12282 = ~1'b0 ;
  assign y12283 = ~1'b0 ;
  assign y12284 = ~n22611 ;
  assign y12285 = ~1'b0 ;
  assign y12286 = ~1'b0 ;
  assign y12287 = n22612 ;
  assign y12288 = n22614 ;
  assign y12289 = ~n22616 ;
  assign y12290 = n22621 ;
  assign y12291 = ~n22622 ;
  assign y12292 = ~1'b0 ;
  assign y12293 = ~1'b0 ;
  assign y12294 = n22623 ;
  assign y12295 = n22625 ;
  assign y12296 = ~n22627 ;
  assign y12297 = ~1'b0 ;
  assign y12298 = ~1'b0 ;
  assign y12299 = ~1'b0 ;
  assign y12300 = ~1'b0 ;
  assign y12301 = ~1'b0 ;
  assign y12302 = 1'b0 ;
  assign y12303 = ~n21781 ;
  assign y12304 = ~n22628 ;
  assign y12305 = 1'b0 ;
  assign y12306 = ~n22630 ;
  assign y12307 = n22635 ;
  assign y12308 = ~1'b0 ;
  assign y12309 = n22636 ;
  assign y12310 = ~n22638 ;
  assign y12311 = n22640 ;
  assign y12312 = ~n22645 ;
  assign y12313 = n22648 ;
  assign y12314 = n22656 ;
  assign y12315 = ~1'b0 ;
  assign y12316 = ~n22662 ;
  assign y12317 = ~1'b0 ;
  assign y12318 = ~n22665 ;
  assign y12319 = n20469 ;
  assign y12320 = n22667 ;
  assign y12321 = ~1'b0 ;
  assign y12322 = ~1'b0 ;
  assign y12323 = n22669 ;
  assign y12324 = ~1'b0 ;
  assign y12325 = ~1'b0 ;
  assign y12326 = ~n22670 ;
  assign y12327 = ~1'b0 ;
  assign y12328 = ~1'b0 ;
  assign y12329 = ~1'b0 ;
  assign y12330 = n22671 ;
  assign y12331 = ~n22672 ;
  assign y12332 = n11698 ;
  assign y12333 = ~1'b0 ;
  assign y12334 = n22674 ;
  assign y12335 = ~n22675 ;
  assign y12336 = ~n22678 ;
  assign y12337 = ~n22680 ;
  assign y12338 = n22681 ;
  assign y12339 = 1'b0 ;
  assign y12340 = n22687 ;
  assign y12341 = ~1'b0 ;
  assign y12342 = ~1'b0 ;
  assign y12343 = 1'b0 ;
  assign y12344 = ~1'b0 ;
  assign y12345 = ~n22693 ;
  assign y12346 = n22695 ;
  assign y12347 = n22701 ;
  assign y12348 = n22702 ;
  assign y12349 = ~1'b0 ;
  assign y12350 = ~1'b0 ;
  assign y12351 = ~1'b0 ;
  assign y12352 = 1'b0 ;
  assign y12353 = ~n22703 ;
  assign y12354 = n22706 ;
  assign y12355 = ~n22708 ;
  assign y12356 = ~1'b0 ;
  assign y12357 = n11759 ;
  assign y12358 = ~n22711 ;
  assign y12359 = n22717 ;
  assign y12360 = ~1'b0 ;
  assign y12361 = n22724 ;
  assign y12362 = n22727 ;
  assign y12363 = n22730 ;
  assign y12364 = ~n22735 ;
  assign y12365 = ~1'b0 ;
  assign y12366 = ~1'b0 ;
  assign y12367 = ~n22736 ;
  assign y12368 = n22748 ;
  assign y12369 = ~1'b0 ;
  assign y12370 = ~n22749 ;
  assign y12371 = ~1'b0 ;
  assign y12372 = n22753 ;
  assign y12373 = ~n22756 ;
  assign y12374 = ~n22763 ;
  assign y12375 = n22764 ;
  assign y12376 = ~1'b0 ;
  assign y12377 = ~n22768 ;
  assign y12378 = ~n22769 ;
  assign y12379 = ~1'b0 ;
  assign y12380 = ~n4707 ;
  assign y12381 = ~n1306 ;
  assign y12382 = n22772 ;
  assign y12383 = n22775 ;
  assign y12384 = n22777 ;
  assign y12385 = ~n22778 ;
  assign y12386 = n8142 ;
  assign y12387 = ~n22779 ;
  assign y12388 = n22780 ;
  assign y12389 = ~n22782 ;
  assign y12390 = ~n22786 ;
  assign y12391 = ~n22787 ;
  assign y12392 = ~n22789 ;
  assign y12393 = ~1'b0 ;
  assign y12394 = ~1'b0 ;
  assign y12395 = ~1'b0 ;
  assign y12396 = n22792 ;
  assign y12397 = n22793 ;
  assign y12398 = ~n22795 ;
  assign y12399 = ~n22800 ;
  assign y12400 = ~1'b0 ;
  assign y12401 = n22803 ;
  assign y12402 = ~1'b0 ;
  assign y12403 = n22804 ;
  assign y12404 = ~n22808 ;
  assign y12405 = ~n22810 ;
  assign y12406 = ~n22812 ;
  assign y12407 = ~n22816 ;
  assign y12408 = ~n22818 ;
  assign y12409 = ~n22820 ;
  assign y12410 = ~1'b0 ;
  assign y12411 = ~n22823 ;
  assign y12412 = ~1'b0 ;
  assign y12413 = n22826 ;
  assign y12414 = n22827 ;
  assign y12415 = n22828 ;
  assign y12416 = n22830 ;
  assign y12417 = n22831 ;
  assign y12418 = ~1'b0 ;
  assign y12419 = n22833 ;
  assign y12420 = n22836 ;
  assign y12421 = ~n22839 ;
  assign y12422 = ~n22840 ;
  assign y12423 = ~n22841 ;
  assign y12424 = ~1'b0 ;
  assign y12425 = n22846 ;
  assign y12426 = n22847 ;
  assign y12427 = ~n12807 ;
  assign y12428 = n22848 ;
  assign y12429 = ~1'b0 ;
  assign y12430 = n22850 ;
  assign y12431 = ~1'b0 ;
  assign y12432 = n4328 ;
  assign y12433 = ~1'b0 ;
  assign y12434 = ~1'b0 ;
  assign y12435 = ~1'b0 ;
  assign y12436 = ~1'b0 ;
  assign y12437 = ~1'b0 ;
  assign y12438 = ~n22851 ;
  assign y12439 = ~1'b0 ;
  assign y12440 = 1'b0 ;
  assign y12441 = ~n22853 ;
  assign y12442 = ~1'b0 ;
  assign y12443 = n2235 ;
  assign y12444 = ~n10177 ;
  assign y12445 = n22854 ;
  assign y12446 = ~n22855 ;
  assign y12447 = n22856 ;
  assign y12448 = ~1'b0 ;
  assign y12449 = n22859 ;
  assign y12450 = ~n22862 ;
  assign y12451 = n22863 ;
  assign y12452 = ~n22864 ;
  assign y12453 = n22868 ;
  assign y12454 = ~1'b0 ;
  assign y12455 = ~n22869 ;
  assign y12456 = ~1'b0 ;
  assign y12457 = ~1'b0 ;
  assign y12458 = ~1'b0 ;
  assign y12459 = n22870 ;
  assign y12460 = ~1'b0 ;
  assign y12461 = ~1'b0 ;
  assign y12462 = 1'b0 ;
  assign y12463 = n22872 ;
  assign y12464 = n22875 ;
  assign y12465 = ~n22877 ;
  assign y12466 = ~1'b0 ;
  assign y12467 = n22881 ;
  assign y12468 = n22882 ;
  assign y12469 = ~n22887 ;
  assign y12470 = ~1'b0 ;
  assign y12471 = n22890 ;
  assign y12472 = ~n22893 ;
  assign y12473 = ~1'b0 ;
  assign y12474 = 1'b0 ;
  assign y12475 = n22894 ;
  assign y12476 = n22895 ;
  assign y12477 = n22896 ;
  assign y12478 = n22902 ;
  assign y12479 = n22905 ;
  assign y12480 = n22906 ;
  assign y12481 = n14234 ;
  assign y12482 = n22911 ;
  assign y12483 = n22913 ;
  assign y12484 = n17481 ;
  assign y12485 = ~n22917 ;
  assign y12486 = ~n22919 ;
  assign y12487 = n22920 ;
  assign y12488 = n22921 ;
  assign y12489 = 1'b0 ;
  assign y12490 = ~1'b0 ;
  assign y12491 = ~1'b0 ;
  assign y12492 = ~n22924 ;
  assign y12493 = ~1'b0 ;
  assign y12494 = ~1'b0 ;
  assign y12495 = ~n22925 ;
  assign y12496 = n22931 ;
  assign y12497 = ~n22934 ;
  assign y12498 = n3897 ;
  assign y12499 = n22935 ;
  assign y12500 = n22938 ;
  assign y12501 = ~n22941 ;
  assign y12502 = ~1'b0 ;
  assign y12503 = ~1'b0 ;
  assign y12504 = n22950 ;
  assign y12505 = ~n22953 ;
  assign y12506 = ~n5633 ;
  assign y12507 = ~n22956 ;
  assign y12508 = n22964 ;
  assign y12509 = ~n22968 ;
  assign y12510 = ~1'b0 ;
  assign y12511 = ~n22971 ;
  assign y12512 = ~n22972 ;
  assign y12513 = ~n22978 ;
  assign y12514 = ~n18077 ;
  assign y12515 = n22979 ;
  assign y12516 = n7806 ;
  assign y12517 = ~1'b0 ;
  assign y12518 = n22980 ;
  assign y12519 = ~n22982 ;
  assign y12520 = ~n22985 ;
  assign y12521 = ~n22991 ;
  assign y12522 = n22994 ;
  assign y12523 = ~1'b0 ;
  assign y12524 = n22995 ;
  assign y12525 = n22996 ;
  assign y12526 = ~n22998 ;
  assign y12527 = n23003 ;
  assign y12528 = ~n23005 ;
  assign y12529 = ~1'b0 ;
  assign y12530 = ~n23010 ;
  assign y12531 = ~1'b0 ;
  assign y12532 = n23015 ;
  assign y12533 = ~n16110 ;
  assign y12534 = ~n23017 ;
  assign y12535 = ~1'b0 ;
  assign y12536 = n1143 ;
  assign y12537 = ~1'b0 ;
  assign y12538 = n16795 ;
  assign y12539 = n23023 ;
  assign y12540 = ~1'b0 ;
  assign y12541 = ~n23025 ;
  assign y12542 = n23030 ;
  assign y12543 = n23031 ;
  assign y12544 = 1'b0 ;
  assign y12545 = n23033 ;
  assign y12546 = ~n23038 ;
  assign y12547 = ~n5961 ;
  assign y12548 = ~n23040 ;
  assign y12549 = n23042 ;
  assign y12550 = n23052 ;
  assign y12551 = ~1'b0 ;
  assign y12552 = ~n23053 ;
  assign y12553 = ~1'b0 ;
  assign y12554 = ~n23054 ;
  assign y12555 = n23055 ;
  assign y12556 = ~n13638 ;
  assign y12557 = n23060 ;
  assign y12558 = n10352 ;
  assign y12559 = 1'b0 ;
  assign y12560 = 1'b0 ;
  assign y12561 = n23062 ;
  assign y12562 = ~n23067 ;
  assign y12563 = ~n23071 ;
  assign y12564 = n23073 ;
  assign y12565 = n23074 ;
  assign y12566 = ~1'b0 ;
  assign y12567 = ~n23076 ;
  assign y12568 = ~n3093 ;
  assign y12569 = ~1'b0 ;
  assign y12570 = ~n9704 ;
  assign y12571 = n23077 ;
  assign y12572 = ~n23080 ;
  assign y12573 = ~1'b0 ;
  assign y12574 = ~n23082 ;
  assign y12575 = ~n23084 ;
  assign y12576 = ~n16669 ;
  assign y12577 = ~n23088 ;
  assign y12578 = ~n23089 ;
  assign y12579 = ~n23090 ;
  assign y12580 = ~n23094 ;
  assign y12581 = ~n23100 ;
  assign y12582 = ~n23104 ;
  assign y12583 = ~n23106 ;
  assign y12584 = ~n23109 ;
  assign y12585 = n23110 ;
  assign y12586 = n23115 ;
  assign y12587 = ~n23116 ;
  assign y12588 = ~1'b0 ;
  assign y12589 = ~1'b0 ;
  assign y12590 = ~n23117 ;
  assign y12591 = n23122 ;
  assign y12592 = ~1'b0 ;
  assign y12593 = ~n23123 ;
  assign y12594 = n23124 ;
  assign y12595 = n23130 ;
  assign y12596 = ~1'b0 ;
  assign y12597 = ~1'b0 ;
  assign y12598 = ~1'b0 ;
  assign y12599 = n23134 ;
  assign y12600 = 1'b0 ;
  assign y12601 = ~n23140 ;
  assign y12602 = n23143 ;
  assign y12603 = n6756 ;
  assign y12604 = ~n23145 ;
  assign y12605 = ~1'b0 ;
  assign y12606 = n23147 ;
  assign y12607 = ~n23148 ;
  assign y12608 = ~1'b0 ;
  assign y12609 = ~1'b0 ;
  assign y12610 = 1'b0 ;
  assign y12611 = ~n12651 ;
  assign y12612 = n23151 ;
  assign y12613 = ~n23154 ;
  assign y12614 = n23155 ;
  assign y12615 = ~1'b0 ;
  assign y12616 = n23158 ;
  assign y12617 = ~n23160 ;
  assign y12618 = ~n13356 ;
  assign y12619 = ~n23162 ;
  assign y12620 = ~1'b0 ;
  assign y12621 = n23163 ;
  assign y12622 = ~n23164 ;
  assign y12623 = ~n23165 ;
  assign y12624 = ~n10238 ;
  assign y12625 = ~n23166 ;
  assign y12626 = ~1'b0 ;
  assign y12627 = ~n23169 ;
  assign y12628 = ~n23170 ;
  assign y12629 = ~n6869 ;
  assign y12630 = n23172 ;
  assign y12631 = n23173 ;
  assign y12632 = n23175 ;
  assign y12633 = ~n23176 ;
  assign y12634 = n23179 ;
  assign y12635 = n23182 ;
  assign y12636 = ~1'b0 ;
  assign y12637 = ~n23192 ;
  assign y12638 = n23193 ;
  assign y12639 = n23194 ;
  assign y12640 = n23195 ;
  assign y12641 = n23196 ;
  assign y12642 = ~1'b0 ;
  assign y12643 = ~n23198 ;
  assign y12644 = ~1'b0 ;
  assign y12645 = ~1'b0 ;
  assign y12646 = ~1'b0 ;
  assign y12647 = ~1'b0 ;
  assign y12648 = ~1'b0 ;
  assign y12649 = ~n23200 ;
  assign y12650 = ~n23205 ;
  assign y12651 = ~1'b0 ;
  assign y12652 = ~1'b0 ;
  assign y12653 = ~1'b0 ;
  assign y12654 = n23211 ;
  assign y12655 = ~1'b0 ;
  assign y12656 = 1'b0 ;
  assign y12657 = ~n9630 ;
  assign y12658 = ~n23213 ;
  assign y12659 = ~n23217 ;
  assign y12660 = ~n23220 ;
  assign y12661 = ~n23222 ;
  assign y12662 = n23225 ;
  assign y12663 = ~1'b0 ;
  assign y12664 = n23231 ;
  assign y12665 = n15746 ;
  assign y12666 = n23232 ;
  assign y12667 = ~n23237 ;
  assign y12668 = ~1'b0 ;
  assign y12669 = ~n13859 ;
  assign y12670 = n23238 ;
  assign y12671 = ~n19924 ;
  assign y12672 = n23240 ;
  assign y12673 = ~1'b0 ;
  assign y12674 = ~1'b0 ;
  assign y12675 = n7335 ;
  assign y12676 = n23242 ;
  assign y12677 = n23243 ;
  assign y12678 = ~n23244 ;
  assign y12679 = n23247 ;
  assign y12680 = ~1'b0 ;
  assign y12681 = ~n23249 ;
  assign y12682 = n23256 ;
  assign y12683 = n23260 ;
  assign y12684 = n23263 ;
  assign y12685 = n23266 ;
  assign y12686 = n23273 ;
  assign y12687 = n12030 ;
  assign y12688 = n23278 ;
  assign y12689 = ~1'b0 ;
  assign y12690 = ~n23285 ;
  assign y12691 = ~n23288 ;
  assign y12692 = n23289 ;
  assign y12693 = ~1'b0 ;
  assign y12694 = n23291 ;
  assign y12695 = ~1'b0 ;
  assign y12696 = n23294 ;
  assign y12697 = ~n23297 ;
  assign y12698 = n23299 ;
  assign y12699 = n23301 ;
  assign y12700 = ~1'b0 ;
  assign y12701 = ~n23303 ;
  assign y12702 = ~1'b0 ;
  assign y12703 = ~n23306 ;
  assign y12704 = ~n23311 ;
  assign y12705 = ~1'b0 ;
  assign y12706 = ~1'b0 ;
  assign y12707 = n23313 ;
  assign y12708 = n23314 ;
  assign y12709 = ~n23316 ;
  assign y12710 = n23325 ;
  assign y12711 = ~1'b0 ;
  assign y12712 = ~n23327 ;
  assign y12713 = n9945 ;
  assign y12714 = ~n6841 ;
  assign y12715 = n23328 ;
  assign y12716 = ~n23329 ;
  assign y12717 = ~1'b0 ;
  assign y12718 = ~n23335 ;
  assign y12719 = ~n23336 ;
  assign y12720 = ~n23340 ;
  assign y12721 = ~1'b0 ;
  assign y12722 = ~n23348 ;
  assign y12723 = ~1'b0 ;
  assign y12724 = n23350 ;
  assign y12725 = ~n23352 ;
  assign y12726 = ~1'b0 ;
  assign y12727 = ~1'b0 ;
  assign y12728 = n2812 ;
  assign y12729 = ~n5668 ;
  assign y12730 = n23353 ;
  assign y12731 = ~n23356 ;
  assign y12732 = n23358 ;
  assign y12733 = ~1'b0 ;
  assign y12734 = ~n23359 ;
  assign y12735 = ~1'b0 ;
  assign y12736 = ~n23369 ;
  assign y12737 = n23370 ;
  assign y12738 = n23375 ;
  assign y12739 = ~n19647 ;
  assign y12740 = ~1'b0 ;
  assign y12741 = n23379 ;
  assign y12742 = n23380 ;
  assign y12743 = ~n23381 ;
  assign y12744 = ~1'b0 ;
  assign y12745 = ~n23383 ;
  assign y12746 = n23385 ;
  assign y12747 = ~n23387 ;
  assign y12748 = ~1'b0 ;
  assign y12749 = n23391 ;
  assign y12750 = ~n23392 ;
  assign y12751 = ~1'b0 ;
  assign y12752 = ~n16673 ;
  assign y12753 = ~1'b0 ;
  assign y12754 = ~n23393 ;
  assign y12755 = ~n23397 ;
  assign y12756 = ~1'b0 ;
  assign y12757 = ~n21382 ;
  assign y12758 = ~1'b0 ;
  assign y12759 = ~1'b0 ;
  assign y12760 = ~1'b0 ;
  assign y12761 = n23399 ;
  assign y12762 = n23400 ;
  assign y12763 = ~n23405 ;
  assign y12764 = ~n23421 ;
  assign y12765 = ~n23424 ;
  assign y12766 = n2232 ;
  assign y12767 = ~n23425 ;
  assign y12768 = ~1'b0 ;
  assign y12769 = 1'b0 ;
  assign y12770 = ~n23428 ;
  assign y12771 = ~n23430 ;
  assign y12772 = ~1'b0 ;
  assign y12773 = ~1'b0 ;
  assign y12774 = ~1'b0 ;
  assign y12775 = n23432 ;
  assign y12776 = ~1'b0 ;
  assign y12777 = ~1'b0 ;
  assign y12778 = ~n23437 ;
  assign y12779 = ~n23441 ;
  assign y12780 = n23444 ;
  assign y12781 = ~n23446 ;
  assign y12782 = ~n21878 ;
  assign y12783 = n23451 ;
  assign y12784 = n23455 ;
  assign y12785 = ~n23457 ;
  assign y12786 = ~n23461 ;
  assign y12787 = n23468 ;
  assign y12788 = ~n23472 ;
  assign y12789 = ~1'b0 ;
  assign y12790 = 1'b0 ;
  assign y12791 = n23473 ;
  assign y12792 = n23474 ;
  assign y12793 = ~n23476 ;
  assign y12794 = n23478 ;
  assign y12795 = ~1'b0 ;
  assign y12796 = n6716 ;
  assign y12797 = ~n23480 ;
  assign y12798 = 1'b0 ;
  assign y12799 = n23481 ;
  assign y12800 = ~n23484 ;
  assign y12801 = ~n15495 ;
  assign y12802 = ~1'b0 ;
  assign y12803 = ~n23500 ;
  assign y12804 = n23505 ;
  assign y12805 = ~n23508 ;
  assign y12806 = n23514 ;
  assign y12807 = n23518 ;
  assign y12808 = ~n23524 ;
  assign y12809 = ~1'b0 ;
  assign y12810 = n23525 ;
  assign y12811 = n23529 ;
  assign y12812 = n23531 ;
  assign y12813 = n23537 ;
  assign y12814 = ~n23539 ;
  assign y12815 = ~1'b0 ;
  assign y12816 = ~1'b0 ;
  assign y12817 = ~n23540 ;
  assign y12818 = ~n23544 ;
  assign y12819 = 1'b0 ;
  assign y12820 = n23547 ;
  assign y12821 = ~n956 ;
  assign y12822 = n23549 ;
  assign y12823 = ~1'b0 ;
  assign y12824 = ~n23557 ;
  assign y12825 = ~1'b0 ;
  assign y12826 = n23563 ;
  assign y12827 = ~1'b0 ;
  assign y12828 = ~1'b0 ;
  assign y12829 = ~1'b0 ;
  assign y12830 = ~n23564 ;
  assign y12831 = ~1'b0 ;
  assign y12832 = ~n23566 ;
  assign y12833 = n23567 ;
  assign y12834 = n23568 ;
  assign y12835 = n23571 ;
  assign y12836 = ~n23575 ;
  assign y12837 = n23580 ;
  assign y12838 = n23582 ;
  assign y12839 = 1'b0 ;
  assign y12840 = ~1'b0 ;
  assign y12841 = ~n23585 ;
  assign y12842 = ~1'b0 ;
  assign y12843 = ~1'b0 ;
  assign y12844 = ~n23586 ;
  assign y12845 = ~n23587 ;
  assign y12846 = ~1'b0 ;
  assign y12847 = ~n12050 ;
  assign y12848 = ~n23588 ;
  assign y12849 = ~n23593 ;
  assign y12850 = ~n23597 ;
  assign y12851 = n23598 ;
  assign y12852 = n23599 ;
  assign y12853 = ~n23604 ;
  assign y12854 = 1'b0 ;
  assign y12855 = ~1'b0 ;
  assign y12856 = ~n11847 ;
  assign y12857 = ~n23607 ;
  assign y12858 = n23610 ;
  assign y12859 = ~n23611 ;
  assign y12860 = ~1'b0 ;
  assign y12861 = ~1'b0 ;
  assign y12862 = ~1'b0 ;
  assign y12863 = ~1'b0 ;
  assign y12864 = ~1'b0 ;
  assign y12865 = ~n23612 ;
  assign y12866 = ~1'b0 ;
  assign y12867 = n23616 ;
  assign y12868 = ~n23617 ;
  assign y12869 = ~n23619 ;
  assign y12870 = n23623 ;
  assign y12871 = n23624 ;
  assign y12872 = ~1'b0 ;
  assign y12873 = ~n2044 ;
  assign y12874 = ~1'b0 ;
  assign y12875 = n23625 ;
  assign y12876 = ~1'b0 ;
  assign y12877 = ~1'b0 ;
  assign y12878 = n23631 ;
  assign y12879 = n23638 ;
  assign y12880 = ~n23639 ;
  assign y12881 = ~1'b0 ;
  assign y12882 = n23646 ;
  assign y12883 = n23649 ;
  assign y12884 = n23656 ;
  assign y12885 = n277 ;
  assign y12886 = n23659 ;
  assign y12887 = ~1'b0 ;
  assign y12888 = ~n23661 ;
  assign y12889 = ~n8970 ;
  assign y12890 = ~n23663 ;
  assign y12891 = n23664 ;
  assign y12892 = ~n23665 ;
  assign y12893 = n23666 ;
  assign y12894 = ~n23668 ;
  assign y12895 = n23674 ;
  assign y12896 = ~1'b0 ;
  assign y12897 = ~n23680 ;
  assign y12898 = ~n23682 ;
  assign y12899 = ~1'b0 ;
  assign y12900 = ~1'b0 ;
  assign y12901 = ~n23686 ;
  assign y12902 = ~n23690 ;
  assign y12903 = ~n23691 ;
  assign y12904 = n23692 ;
  assign y12905 = ~1'b0 ;
  assign y12906 = n23695 ;
  assign y12907 = ~n23696 ;
  assign y12908 = n23700 ;
  assign y12909 = ~1'b0 ;
  assign y12910 = n23712 ;
  assign y12911 = 1'b0 ;
  assign y12912 = ~1'b0 ;
  assign y12913 = n23715 ;
  assign y12914 = ~n22756 ;
  assign y12915 = ~1'b0 ;
  assign y12916 = n23716 ;
  assign y12917 = n23717 ;
  assign y12918 = n23718 ;
  assign y12919 = ~1'b0 ;
  assign y12920 = n23719 ;
  assign y12921 = ~n23720 ;
  assign y12922 = n23726 ;
  assign y12923 = 1'b0 ;
  assign y12924 = ~n23729 ;
  assign y12925 = ~n23731 ;
  assign y12926 = ~1'b0 ;
  assign y12927 = ~1'b0 ;
  assign y12928 = ~1'b0 ;
  assign y12929 = n23734 ;
  assign y12930 = ~n23739 ;
  assign y12931 = ~n3991 ;
  assign y12932 = ~n23741 ;
  assign y12933 = ~n14305 ;
  assign y12934 = n23742 ;
  assign y12935 = ~n23744 ;
  assign y12936 = ~1'b0 ;
  assign y12937 = n23747 ;
  assign y12938 = ~1'b0 ;
  assign y12939 = ~n23764 ;
  assign y12940 = n23768 ;
  assign y12941 = ~n23777 ;
  assign y12942 = n23778 ;
  assign y12943 = ~n23779 ;
  assign y12944 = n23781 ;
  assign y12945 = ~1'b0 ;
  assign y12946 = 1'b0 ;
  assign y12947 = ~n23783 ;
  assign y12948 = ~1'b0 ;
  assign y12949 = ~1'b0 ;
  assign y12950 = 1'b0 ;
  assign y12951 = n23788 ;
  assign y12952 = ~n23792 ;
  assign y12953 = ~1'b0 ;
  assign y12954 = ~n23794 ;
  assign y12955 = ~n23795 ;
  assign y12956 = 1'b0 ;
  assign y12957 = ~n23799 ;
  assign y12958 = n23801 ;
  assign y12959 = ~1'b0 ;
  assign y12960 = n23805 ;
  assign y12961 = ~n23814 ;
  assign y12962 = ~n23819 ;
  assign y12963 = n12285 ;
  assign y12964 = ~1'b0 ;
  assign y12965 = ~n23822 ;
  assign y12966 = 1'b0 ;
  assign y12967 = n23825 ;
  assign y12968 = ~1'b0 ;
  assign y12969 = 1'b0 ;
  assign y12970 = ~1'b0 ;
  assign y12971 = ~1'b0 ;
  assign y12972 = ~n23826 ;
  assign y12973 = ~1'b0 ;
  assign y12974 = ~n23828 ;
  assign y12975 = ~1'b0 ;
  assign y12976 = n23829 ;
  assign y12977 = n23830 ;
  assign y12978 = n23832 ;
  assign y12979 = n8102 ;
  assign y12980 = n23833 ;
  assign y12981 = n23841 ;
  assign y12982 = ~n23845 ;
  assign y12983 = n23847 ;
  assign y12984 = ~n23849 ;
  assign y12985 = n23851 ;
  assign y12986 = ~n23861 ;
  assign y12987 = n23862 ;
  assign y12988 = n23864 ;
  assign y12989 = n23867 ;
  assign y12990 = 1'b0 ;
  assign y12991 = ~n23869 ;
  assign y12992 = n21954 ;
  assign y12993 = ~n23873 ;
  assign y12994 = ~1'b0 ;
  assign y12995 = n23874 ;
  assign y12996 = n23878 ;
  assign y12997 = ~n23879 ;
  assign y12998 = ~n23882 ;
  assign y12999 = ~n23888 ;
  assign y13000 = ~1'b0 ;
  assign y13001 = ~n23889 ;
  assign y13002 = ~1'b0 ;
  assign y13003 = n23894 ;
  assign y13004 = 1'b0 ;
  assign y13005 = ~1'b0 ;
  assign y13006 = ~n23896 ;
  assign y13007 = ~n23899 ;
  assign y13008 = ~n23902 ;
  assign y13009 = ~1'b0 ;
  assign y13010 = ~n23904 ;
  assign y13011 = ~n23905 ;
  assign y13012 = n23907 ;
  assign y13013 = n23909 ;
  assign y13014 = ~1'b0 ;
  assign y13015 = ~1'b0 ;
  assign y13016 = ~1'b0 ;
  assign y13017 = ~n23910 ;
  assign y13018 = ~1'b0 ;
  assign y13019 = n23911 ;
  assign y13020 = n23912 ;
  assign y13021 = ~1'b0 ;
  assign y13022 = ~1'b0 ;
  assign y13023 = n23913 ;
  assign y13024 = n23916 ;
  assign y13025 = ~n23917 ;
  assign y13026 = n7464 ;
  assign y13027 = ~n23925 ;
  assign y13028 = ~n23926 ;
  assign y13029 = n20068 ;
  assign y13030 = n23929 ;
  assign y13031 = ~1'b0 ;
  assign y13032 = ~1'b0 ;
  assign y13033 = n23934 ;
  assign y13034 = ~1'b0 ;
  assign y13035 = n23943 ;
  assign y13036 = ~n23945 ;
  assign y13037 = n23951 ;
  assign y13038 = ~1'b0 ;
  assign y13039 = ~n23952 ;
  assign y13040 = ~n23954 ;
  assign y13041 = ~1'b0 ;
  assign y13042 = ~n23957 ;
  assign y13043 = ~n23960 ;
  assign y13044 = ~1'b0 ;
  assign y13045 = ~n23961 ;
  assign y13046 = ~n23965 ;
  assign y13047 = ~n23968 ;
  assign y13048 = n23971 ;
  assign y13049 = ~n19362 ;
  assign y13050 = ~1'b0 ;
  assign y13051 = ~n23973 ;
  assign y13052 = ~1'b0 ;
  assign y13053 = ~n23975 ;
  assign y13054 = n23978 ;
  assign y13055 = ~n24004 ;
  assign y13056 = ~1'b0 ;
  assign y13057 = ~n24007 ;
  assign y13058 = ~n24009 ;
  assign y13059 = ~n24011 ;
  assign y13060 = ~n24013 ;
  assign y13061 = ~1'b0 ;
  assign y13062 = ~1'b0 ;
  assign y13063 = n24016 ;
  assign y13064 = n24017 ;
  assign y13065 = ~1'b0 ;
  assign y13066 = n798 ;
  assign y13067 = n24019 ;
  assign y13068 = ~n24020 ;
  assign y13069 = ~1'b0 ;
  assign y13070 = ~1'b0 ;
  assign y13071 = ~n24025 ;
  assign y13072 = ~n24029 ;
  assign y13073 = n24030 ;
  assign y13074 = ~1'b0 ;
  assign y13075 = ~1'b0 ;
  assign y13076 = 1'b0 ;
  assign y13077 = ~n24032 ;
  assign y13078 = ~n5282 ;
  assign y13079 = ~n22408 ;
  assign y13080 = ~1'b0 ;
  assign y13081 = ~1'b0 ;
  assign y13082 = ~n24038 ;
  assign y13083 = ~n24039 ;
  assign y13084 = n24045 ;
  assign y13085 = n24046 ;
  assign y13086 = ~n24047 ;
  assign y13087 = ~1'b0 ;
  assign y13088 = n24048 ;
  assign y13089 = n24049 ;
  assign y13090 = n24050 ;
  assign y13091 = n24053 ;
  assign y13092 = ~n24055 ;
  assign y13093 = ~n24057 ;
  assign y13094 = n24061 ;
  assign y13095 = ~1'b0 ;
  assign y13096 = n24063 ;
  assign y13097 = ~n24066 ;
  assign y13098 = ~1'b0 ;
  assign y13099 = n24067 ;
  assign y13100 = ~n24069 ;
  assign y13101 = ~1'b0 ;
  assign y13102 = n24072 ;
  assign y13103 = ~1'b0 ;
  assign y13104 = n24074 ;
  assign y13105 = ~n24076 ;
  assign y13106 = ~1'b0 ;
  assign y13107 = ~n24078 ;
  assign y13108 = n24081 ;
  assign y13109 = n24082 ;
  assign y13110 = ~1'b0 ;
  assign y13111 = ~1'b0 ;
  assign y13112 = ~n24086 ;
  assign y13113 = n24091 ;
  assign y13114 = n24096 ;
  assign y13115 = n24097 ;
  assign y13116 = ~1'b0 ;
  assign y13117 = n24099 ;
  assign y13118 = n24105 ;
  assign y13119 = ~1'b0 ;
  assign y13120 = n24109 ;
  assign y13121 = ~n24114 ;
  assign y13122 = ~1'b0 ;
  assign y13123 = ~1'b0 ;
  assign y13124 = n390 ;
  assign y13125 = ~n24115 ;
  assign y13126 = ~1'b0 ;
  assign y13127 = ~n24116 ;
  assign y13128 = ~1'b0 ;
  assign y13129 = n24120 ;
  assign y13130 = ~n24122 ;
  assign y13131 = n24123 ;
  assign y13132 = n24124 ;
  assign y13133 = n24125 ;
  assign y13134 = n24126 ;
  assign y13135 = ~n24128 ;
  assign y13136 = ~1'b0 ;
  assign y13137 = ~1'b0 ;
  assign y13138 = ~n24130 ;
  assign y13139 = n24139 ;
  assign y13140 = n24140 ;
  assign y13141 = ~n24141 ;
  assign y13142 = n19062 ;
  assign y13143 = n24143 ;
  assign y13144 = n24144 ;
  assign y13145 = n24145 ;
  assign y13146 = n24146 ;
  assign y13147 = ~n24150 ;
  assign y13148 = ~n24151 ;
  assign y13149 = ~1'b0 ;
  assign y13150 = n24152 ;
  assign y13151 = ~n24153 ;
  assign y13152 = n24154 ;
  assign y13153 = ~n21062 ;
  assign y13154 = ~n24166 ;
  assign y13155 = ~n24167 ;
  assign y13156 = n24168 ;
  assign y13157 = ~n24170 ;
  assign y13158 = n24173 ;
  assign y13159 = ~n24174 ;
  assign y13160 = ~n24175 ;
  assign y13161 = ~n24177 ;
  assign y13162 = ~1'b0 ;
  assign y13163 = ~n24183 ;
  assign y13164 = ~1'b0 ;
  assign y13165 = ~n15556 ;
  assign y13166 = ~1'b0 ;
  assign y13167 = ~1'b0 ;
  assign y13168 = n6988 ;
  assign y13169 = n24186 ;
  assign y13170 = n24189 ;
  assign y13171 = ~n24191 ;
  assign y13172 = ~1'b0 ;
  assign y13173 = ~n24192 ;
  assign y13174 = ~n24196 ;
  assign y13175 = n24202 ;
  assign y13176 = ~n24203 ;
  assign y13177 = ~1'b0 ;
  assign y13178 = ~1'b0 ;
  assign y13179 = ~n24209 ;
  assign y13180 = ~n24216 ;
  assign y13181 = ~1'b0 ;
  assign y13182 = ~n24221 ;
  assign y13183 = ~1'b0 ;
  assign y13184 = ~n24222 ;
  assign y13185 = n24226 ;
  assign y13186 = ~n5526 ;
  assign y13187 = n24230 ;
  assign y13188 = ~1'b0 ;
  assign y13189 = n24231 ;
  assign y13190 = ~n24233 ;
  assign y13191 = ~1'b0 ;
  assign y13192 = ~n24234 ;
  assign y13193 = ~1'b0 ;
  assign y13194 = ~n24236 ;
  assign y13195 = n24238 ;
  assign y13196 = n24240 ;
  assign y13197 = n24246 ;
  assign y13198 = ~n24247 ;
  assign y13199 = ~n24252 ;
  assign y13200 = ~1'b0 ;
  assign y13201 = ~n24260 ;
  assign y13202 = n10245 ;
  assign y13203 = n24261 ;
  assign y13204 = ~1'b0 ;
  assign y13205 = ~n24262 ;
  assign y13206 = ~n24265 ;
  assign y13207 = n1205 ;
  assign y13208 = ~n24268 ;
  assign y13209 = ~n24275 ;
  assign y13210 = n24277 ;
  assign y13211 = n24279 ;
  assign y13212 = ~1'b0 ;
  assign y13213 = n24280 ;
  assign y13214 = ~1'b0 ;
  assign y13215 = n14749 ;
  assign y13216 = n24282 ;
  assign y13217 = ~1'b0 ;
  assign y13218 = n24284 ;
  assign y13219 = n24286 ;
  assign y13220 = ~1'b0 ;
  assign y13221 = n24289 ;
  assign y13222 = ~n24291 ;
  assign y13223 = ~n24295 ;
  assign y13224 = ~n24297 ;
  assign y13225 = ~n24299 ;
  assign y13226 = ~1'b0 ;
  assign y13227 = ~1'b0 ;
  assign y13228 = n24301 ;
  assign y13229 = n24302 ;
  assign y13230 = ~1'b0 ;
  assign y13231 = ~1'b0 ;
  assign y13232 = ~1'b0 ;
  assign y13233 = n24307 ;
  assign y13234 = ~n24308 ;
  assign y13235 = 1'b0 ;
  assign y13236 = n24312 ;
  assign y13237 = n24313 ;
  assign y13238 = ~n24315 ;
  assign y13239 = ~n24317 ;
  assign y13240 = ~1'b0 ;
  assign y13241 = ~1'b0 ;
  assign y13242 = ~n24322 ;
  assign y13243 = n24324 ;
  assign y13244 = ~1'b0 ;
  assign y13245 = ~1'b0 ;
  assign y13246 = n24329 ;
  assign y13247 = ~n24330 ;
  assign y13248 = ~1'b0 ;
  assign y13249 = ~n23120 ;
  assign y13250 = n15680 ;
  assign y13251 = n24332 ;
  assign y13252 = n24336 ;
  assign y13253 = ~1'b0 ;
  assign y13254 = ~n24341 ;
  assign y13255 = ~n24342 ;
  assign y13256 = n968 ;
  assign y13257 = ~1'b0 ;
  assign y13258 = ~n24345 ;
  assign y13259 = n24348 ;
  assign y13260 = n24350 ;
  assign y13261 = ~n24362 ;
  assign y13262 = ~n24363 ;
  assign y13263 = ~n24367 ;
  assign y13264 = n2883 ;
  assign y13265 = ~n24372 ;
  assign y13266 = ~n24378 ;
  assign y13267 = ~n24381 ;
  assign y13268 = ~n24382 ;
  assign y13269 = ~n24383 ;
  assign y13270 = n24384 ;
  assign y13271 = ~n24385 ;
  assign y13272 = n24386 ;
  assign y13273 = ~n24389 ;
  assign y13274 = n24393 ;
  assign y13275 = ~n24395 ;
  assign y13276 = n24396 ;
  assign y13277 = ~1'b0 ;
  assign y13278 = n24397 ;
  assign y13279 = n24400 ;
  assign y13280 = n24403 ;
  assign y13281 = ~1'b0 ;
  assign y13282 = n24408 ;
  assign y13283 = ~n24410 ;
  assign y13284 = ~1'b0 ;
  assign y13285 = n24417 ;
  assign y13286 = ~n24420 ;
  assign y13287 = ~1'b0 ;
  assign y13288 = ~n24422 ;
  assign y13289 = n24425 ;
  assign y13290 = n19884 ;
  assign y13291 = ~n24426 ;
  assign y13292 = ~n24430 ;
  assign y13293 = ~n24432 ;
  assign y13294 = ~n24433 ;
  assign y13295 = ~n24436 ;
  assign y13296 = ~n24440 ;
  assign y13297 = ~1'b0 ;
  assign y13298 = ~1'b0 ;
  assign y13299 = ~n24441 ;
  assign y13300 = ~n24443 ;
  assign y13301 = ~n24446 ;
  assign y13302 = ~n24448 ;
  assign y13303 = ~1'b0 ;
  assign y13304 = n8468 ;
  assign y13305 = ~n24450 ;
  assign y13306 = ~1'b0 ;
  assign y13307 = n24451 ;
  assign y13308 = ~n24452 ;
  assign y13309 = 1'b0 ;
  assign y13310 = n11170 ;
  assign y13311 = n24456 ;
  assign y13312 = n24458 ;
  assign y13313 = n24459 ;
  assign y13314 = ~n24464 ;
  assign y13315 = ~1'b0 ;
  assign y13316 = ~n1973 ;
  assign y13317 = n24466 ;
  assign y13318 = n24469 ;
  assign y13319 = ~n24470 ;
  assign y13320 = ~1'b0 ;
  assign y13321 = n24471 ;
  assign y13322 = ~1'b0 ;
  assign y13323 = n24474 ;
  assign y13324 = n24475 ;
  assign y13325 = n24477 ;
  assign y13326 = ~n24483 ;
  assign y13327 = n24485 ;
  assign y13328 = ~1'b0 ;
  assign y13329 = n24486 ;
  assign y13330 = n24487 ;
  assign y13331 = ~1'b0 ;
  assign y13332 = n24493 ;
  assign y13333 = ~1'b0 ;
  assign y13334 = ~n10477 ;
  assign y13335 = ~n24494 ;
  assign y13336 = ~1'b0 ;
  assign y13337 = n24495 ;
  assign y13338 = ~n24497 ;
  assign y13339 = n24498 ;
  assign y13340 = n24499 ;
  assign y13341 = ~n24502 ;
  assign y13342 = ~n24504 ;
  assign y13343 = n24505 ;
  assign y13344 = n24513 ;
  assign y13345 = n24520 ;
  assign y13346 = n21803 ;
  assign y13347 = n20425 ;
  assign y13348 = n24521 ;
  assign y13349 = n24524 ;
  assign y13350 = ~n4831 ;
  assign y13351 = n24526 ;
  assign y13352 = ~1'b0 ;
  assign y13353 = n24532 ;
  assign y13354 = n24533 ;
  assign y13355 = ~1'b0 ;
  assign y13356 = ~1'b0 ;
  assign y13357 = ~n24534 ;
  assign y13358 = n24538 ;
  assign y13359 = n24539 ;
  assign y13360 = 1'b0 ;
  assign y13361 = n24541 ;
  assign y13362 = ~n24542 ;
  assign y13363 = ~1'b0 ;
  assign y13364 = ~n24544 ;
  assign y13365 = ~n24545 ;
  assign y13366 = n24549 ;
  assign y13367 = 1'b0 ;
  assign y13368 = ~n16770 ;
  assign y13369 = n24550 ;
  assign y13370 = n24551 ;
  assign y13371 = n24553 ;
  assign y13372 = n24559 ;
  assign y13373 = ~n12053 ;
  assign y13374 = n24561 ;
  assign y13375 = ~1'b0 ;
  assign y13376 = ~1'b0 ;
  assign y13377 = 1'b0 ;
  assign y13378 = n24570 ;
  assign y13379 = n24571 ;
  assign y13380 = n24588 ;
  assign y13381 = ~n2572 ;
  assign y13382 = ~n24590 ;
  assign y13383 = n24592 ;
  assign y13384 = ~1'b0 ;
  assign y13385 = n24593 ;
  assign y13386 = 1'b0 ;
  assign y13387 = ~1'b0 ;
  assign y13388 = n24597 ;
  assign y13389 = ~n24599 ;
  assign y13390 = ~n24600 ;
  assign y13391 = ~n24601 ;
  assign y13392 = ~1'b0 ;
  assign y13393 = n5108 ;
  assign y13394 = ~n12485 ;
  assign y13395 = ~n24610 ;
  assign y13396 = ~1'b0 ;
  assign y13397 = ~1'b0 ;
  assign y13398 = ~1'b0 ;
  assign y13399 = n24612 ;
  assign y13400 = n16234 ;
  assign y13401 = n24614 ;
  assign y13402 = ~n24617 ;
  assign y13403 = ~1'b0 ;
  assign y13404 = ~n24619 ;
  assign y13405 = ~1'b0 ;
  assign y13406 = n24622 ;
  assign y13407 = ~n24628 ;
  assign y13408 = ~n4422 ;
  assign y13409 = n6912 ;
  assign y13410 = ~1'b0 ;
  assign y13411 = ~1'b0 ;
  assign y13412 = ~1'b0 ;
  assign y13413 = n13285 ;
  assign y13414 = ~n24630 ;
  assign y13415 = ~n24633 ;
  assign y13416 = ~n24635 ;
  assign y13417 = ~1'b0 ;
  assign y13418 = n24638 ;
  assign y13419 = ~n24640 ;
  assign y13420 = ~n24643 ;
  assign y13421 = ~n24646 ;
  assign y13422 = n24647 ;
  assign y13423 = ~n24648 ;
  assign y13424 = n24651 ;
  assign y13425 = n2179 ;
  assign y13426 = ~n24653 ;
  assign y13427 = ~1'b0 ;
  assign y13428 = n24655 ;
  assign y13429 = n24656 ;
  assign y13430 = ~1'b0 ;
  assign y13431 = ~1'b0 ;
  assign y13432 = ~1'b0 ;
  assign y13433 = n24657 ;
  assign y13434 = ~1'b0 ;
  assign y13435 = ~n24658 ;
  assign y13436 = n24660 ;
  assign y13437 = ~n24671 ;
  assign y13438 = n24672 ;
  assign y13439 = ~n15839 ;
  assign y13440 = ~n24675 ;
  assign y13441 = n24677 ;
  assign y13442 = 1'b0 ;
  assign y13443 = ~n24681 ;
  assign y13444 = ~1'b0 ;
  assign y13445 = n24682 ;
  assign y13446 = n24685 ;
  assign y13447 = ~n24690 ;
  assign y13448 = ~n24698 ;
  assign y13449 = n24699 ;
  assign y13450 = n24706 ;
  assign y13451 = ~n15071 ;
  assign y13452 = n24711 ;
  assign y13453 = n24712 ;
  assign y13454 = ~1'b0 ;
  assign y13455 = ~1'b0 ;
  assign y13456 = ~1'b0 ;
  assign y13457 = n24713 ;
  assign y13458 = n24714 ;
  assign y13459 = n24716 ;
  assign y13460 = ~n24722 ;
  assign y13461 = n24723 ;
  assign y13462 = ~1'b0 ;
  assign y13463 = n24731 ;
  assign y13464 = n19595 ;
  assign y13465 = ~1'b0 ;
  assign y13466 = n24736 ;
  assign y13467 = n24739 ;
  assign y13468 = n24741 ;
  assign y13469 = ~n24742 ;
  assign y13470 = 1'b0 ;
  assign y13471 = n24743 ;
  assign y13472 = ~n24745 ;
  assign y13473 = ~1'b0 ;
  assign y13474 = ~1'b0 ;
  assign y13475 = n24747 ;
  assign y13476 = ~n9703 ;
  assign y13477 = ~n14542 ;
  assign y13478 = ~n24751 ;
  assign y13479 = ~1'b0 ;
  assign y13480 = n24755 ;
  assign y13481 = ~n24756 ;
  assign y13482 = n24759 ;
  assign y13483 = ~n24760 ;
  assign y13484 = n150 ;
  assign y13485 = ~n24762 ;
  assign y13486 = n24764 ;
  assign y13487 = ~n24766 ;
  assign y13488 = ~1'b0 ;
  assign y13489 = ~1'b0 ;
  assign y13490 = n24773 ;
  assign y13491 = n24778 ;
  assign y13492 = ~1'b0 ;
  assign y13493 = ~1'b0 ;
  assign y13494 = ~n24779 ;
  assign y13495 = ~1'b0 ;
  assign y13496 = n24782 ;
  assign y13497 = n24784 ;
  assign y13498 = ~n24787 ;
  assign y13499 = ~1'b0 ;
  assign y13500 = ~n24794 ;
  assign y13501 = ~1'b0 ;
  assign y13502 = n24795 ;
  assign y13503 = ~n24798 ;
  assign y13504 = ~1'b0 ;
  assign y13505 = ~n24802 ;
  assign y13506 = ~n24805 ;
  assign y13507 = n16295 ;
  assign y13508 = ~n24807 ;
  assign y13509 = ~1'b0 ;
  assign y13510 = 1'b0 ;
  assign y13511 = ~1'b0 ;
  assign y13512 = ~1'b0 ;
  assign y13513 = ~1'b0 ;
  assign y13514 = ~1'b0 ;
  assign y13515 = ~n24808 ;
  assign y13516 = n24811 ;
  assign y13517 = n24812 ;
  assign y13518 = n24813 ;
  assign y13519 = ~1'b0 ;
  assign y13520 = n24815 ;
  assign y13521 = ~1'b0 ;
  assign y13522 = ~1'b0 ;
  assign y13523 = ~1'b0 ;
  assign y13524 = ~1'b0 ;
  assign y13525 = ~1'b0 ;
  assign y13526 = n24816 ;
  assign y13527 = n24820 ;
  assign y13528 = ~1'b0 ;
  assign y13529 = n24821 ;
  assign y13530 = ~n24823 ;
  assign y13531 = ~n24825 ;
  assign y13532 = ~n24826 ;
  assign y13533 = ~n15674 ;
  assign y13534 = ~n24829 ;
  assign y13535 = ~1'b0 ;
  assign y13536 = ~1'b0 ;
  assign y13537 = n24834 ;
  assign y13538 = ~n24835 ;
  assign y13539 = ~1'b0 ;
  assign y13540 = ~1'b0 ;
  assign y13541 = ~1'b0 ;
  assign y13542 = ~n24836 ;
  assign y13543 = n24844 ;
  assign y13544 = ~1'b0 ;
  assign y13545 = n24846 ;
  assign y13546 = n24850 ;
  assign y13547 = ~1'b0 ;
  assign y13548 = ~n9163 ;
  assign y13549 = n18307 ;
  assign y13550 = ~n24851 ;
  assign y13551 = n24853 ;
  assign y13552 = ~1'b0 ;
  assign y13553 = n3319 ;
  assign y13554 = ~1'b0 ;
  assign y13555 = n24856 ;
  assign y13556 = ~1'b0 ;
  assign y13557 = ~n24857 ;
  assign y13558 = n24858 ;
  assign y13559 = ~1'b0 ;
  assign y13560 = n24863 ;
  assign y13561 = ~n24867 ;
  assign y13562 = ~1'b0 ;
  assign y13563 = ~n24872 ;
  assign y13564 = ~n24874 ;
  assign y13565 = n24876 ;
  assign y13566 = ~n24878 ;
  assign y13567 = ~1'b0 ;
  assign y13568 = n24881 ;
  assign y13569 = n24882 ;
  assign y13570 = n24883 ;
  assign y13571 = ~1'b0 ;
  assign y13572 = ~1'b0 ;
  assign y13573 = n24885 ;
  assign y13574 = ~n24887 ;
  assign y13575 = ~n24888 ;
  assign y13576 = n24891 ;
  assign y13577 = ~1'b0 ;
  assign y13578 = ~n11295 ;
  assign y13579 = n24892 ;
  assign y13580 = ~1'b0 ;
  assign y13581 = ~n24893 ;
  assign y13582 = ~n24903 ;
  assign y13583 = n24905 ;
  assign y13584 = n24908 ;
  assign y13585 = ~1'b0 ;
  assign y13586 = ~n24909 ;
  assign y13587 = n24910 ;
  assign y13588 = ~n24915 ;
  assign y13589 = n24917 ;
  assign y13590 = n24927 ;
  assign y13591 = ~n24928 ;
  assign y13592 = ~1'b0 ;
  assign y13593 = ~n24929 ;
  assign y13594 = ~n24930 ;
  assign y13595 = ~n24931 ;
  assign y13596 = ~n24933 ;
  assign y13597 = ~n24935 ;
  assign y13598 = ~n24944 ;
  assign y13599 = ~1'b0 ;
  assign y13600 = ~1'b0 ;
  assign y13601 = ~1'b0 ;
  assign y13602 = n24945 ;
  assign y13603 = ~n24950 ;
  assign y13604 = ~n24952 ;
  assign y13605 = ~1'b0 ;
  assign y13606 = n24953 ;
  assign y13607 = ~1'b0 ;
  assign y13608 = n24954 ;
  assign y13609 = ~n24957 ;
  assign y13610 = ~1'b0 ;
  assign y13611 = ~n24958 ;
  assign y13612 = ~1'b0 ;
  assign y13613 = n24959 ;
  assign y13614 = ~n24963 ;
  assign y13615 = 1'b0 ;
  assign y13616 = ~1'b0 ;
  assign y13617 = ~n8904 ;
  assign y13618 = ~n24964 ;
  assign y13619 = ~n24965 ;
  assign y13620 = n24967 ;
  assign y13621 = ~1'b0 ;
  assign y13622 = n24971 ;
  assign y13623 = ~1'b0 ;
  assign y13624 = n24972 ;
  assign y13625 = ~n4919 ;
  assign y13626 = n24973 ;
  assign y13627 = ~n24976 ;
  assign y13628 = ~n2321 ;
  assign y13629 = n24977 ;
  assign y13630 = n24978 ;
  assign y13631 = ~1'b0 ;
  assign y13632 = ~1'b0 ;
  assign y13633 = n24982 ;
  assign y13634 = ~n24983 ;
  assign y13635 = ~1'b0 ;
  assign y13636 = n24986 ;
  assign y13637 = n3114 ;
  assign y13638 = n24988 ;
  assign y13639 = ~n24992 ;
  assign y13640 = ~1'b0 ;
  assign y13641 = ~n1582 ;
  assign y13642 = n24994 ;
  assign y13643 = ~n15246 ;
  assign y13644 = ~n24996 ;
  assign y13645 = n16507 ;
  assign y13646 = ~1'b0 ;
  assign y13647 = 1'b0 ;
  assign y13648 = ~1'b0 ;
  assign y13649 = ~1'b0 ;
  assign y13650 = ~n24997 ;
  assign y13651 = ~1'b0 ;
  assign y13652 = ~1'b0 ;
  assign y13653 = n24999 ;
  assign y13654 = ~n25001 ;
  assign y13655 = ~1'b0 ;
  assign y13656 = ~1'b0 ;
  assign y13657 = ~1'b0 ;
  assign y13658 = ~n25004 ;
  assign y13659 = n25007 ;
  assign y13660 = ~1'b0 ;
  assign y13661 = n25012 ;
  assign y13662 = ~1'b0 ;
  assign y13663 = ~n25016 ;
  assign y13664 = ~1'b0 ;
  assign y13665 = n25017 ;
  assign y13666 = ~n25018 ;
  assign y13667 = ~n263 ;
  assign y13668 = n25019 ;
  assign y13669 = ~n25023 ;
  assign y13670 = ~1'b0 ;
  assign y13671 = ~n25027 ;
  assign y13672 = ~n25028 ;
  assign y13673 = ~1'b0 ;
  assign y13674 = ~1'b0 ;
  assign y13675 = ~n25029 ;
  assign y13676 = ~n25031 ;
  assign y13677 = n25032 ;
  assign y13678 = ~n25033 ;
  assign y13679 = n25036 ;
  assign y13680 = ~n25039 ;
  assign y13681 = ~n25041 ;
  assign y13682 = n25042 ;
  assign y13683 = ~n25046 ;
  assign y13684 = n25047 ;
  assign y13685 = ~n25048 ;
  assign y13686 = ~1'b0 ;
  assign y13687 = ~n25050 ;
  assign y13688 = ~n25052 ;
  assign y13689 = n25055 ;
  assign y13690 = ~n25058 ;
  assign y13691 = ~n25060 ;
  assign y13692 = n25061 ;
  assign y13693 = ~n25062 ;
  assign y13694 = ~1'b0 ;
  assign y13695 = ~1'b0 ;
  assign y13696 = n25064 ;
  assign y13697 = n25065 ;
  assign y13698 = ~n25068 ;
  assign y13699 = n25069 ;
  assign y13700 = n25072 ;
  assign y13701 = ~n25073 ;
  assign y13702 = ~n25077 ;
  assign y13703 = ~1'b0 ;
  assign y13704 = ~n25078 ;
  assign y13705 = ~1'b0 ;
  assign y13706 = ~1'b0 ;
  assign y13707 = ~1'b0 ;
  assign y13708 = ~n25082 ;
  assign y13709 = n20714 ;
  assign y13710 = ~1'b0 ;
  assign y13711 = ~n25083 ;
  assign y13712 = ~1'b0 ;
  assign y13713 = ~1'b0 ;
  assign y13714 = n25086 ;
  assign y13715 = ~n25087 ;
  assign y13716 = n25089 ;
  assign y13717 = ~1'b0 ;
  assign y13718 = ~1'b0 ;
  assign y13719 = 1'b0 ;
  assign y13720 = ~1'b0 ;
  assign y13721 = n14456 ;
  assign y13722 = ~1'b0 ;
  assign y13723 = ~n25091 ;
  assign y13724 = ~1'b0 ;
  assign y13725 = n25092 ;
  assign y13726 = ~1'b0 ;
  assign y13727 = ~n25098 ;
  assign y13728 = n8495 ;
  assign y13729 = ~n25102 ;
  assign y13730 = n25107 ;
  assign y13731 = ~1'b0 ;
  assign y13732 = ~n25109 ;
  assign y13733 = n25115 ;
  assign y13734 = ~n25117 ;
  assign y13735 = ~1'b0 ;
  assign y13736 = ~1'b0 ;
  assign y13737 = ~n25120 ;
  assign y13738 = ~n25122 ;
  assign y13739 = ~1'b0 ;
  assign y13740 = ~n25124 ;
  assign y13741 = ~1'b0 ;
  assign y13742 = ~n25126 ;
  assign y13743 = n25127 ;
  assign y13744 = ~n25128 ;
  assign y13745 = n25129 ;
  assign y13746 = ~n25137 ;
  assign y13747 = n25140 ;
  assign y13748 = ~1'b0 ;
  assign y13749 = n25141 ;
  assign y13750 = n25144 ;
  assign y13751 = ~n25148 ;
  assign y13752 = n25151 ;
  assign y13753 = ~n25152 ;
  assign y13754 = ~1'b0 ;
  assign y13755 = ~n25155 ;
  assign y13756 = n25157 ;
  assign y13757 = ~1'b0 ;
  assign y13758 = n25158 ;
  assign y13759 = ~1'b0 ;
  assign y13760 = ~n25161 ;
  assign y13761 = n3823 ;
  assign y13762 = ~1'b0 ;
  assign y13763 = ~1'b0 ;
  assign y13764 = ~n25164 ;
  assign y13765 = ~1'b0 ;
  assign y13766 = ~n25166 ;
  assign y13767 = ~1'b0 ;
  assign y13768 = n25168 ;
  assign y13769 = n2940 ;
  assign y13770 = n25171 ;
  assign y13771 = n25174 ;
  assign y13772 = ~n25175 ;
  assign y13773 = n25182 ;
  assign y13774 = ~n25184 ;
  assign y13775 = ~n25186 ;
  assign y13776 = n12516 ;
  assign y13777 = ~n25188 ;
  assign y13778 = n7530 ;
  assign y13779 = n25189 ;
  assign y13780 = 1'b0 ;
  assign y13781 = n25193 ;
  assign y13782 = ~n13473 ;
  assign y13783 = ~n25194 ;
  assign y13784 = ~n25199 ;
  assign y13785 = ~1'b0 ;
  assign y13786 = ~n25205 ;
  assign y13787 = ~n25207 ;
  assign y13788 = ~1'b0 ;
  assign y13789 = ~n15997 ;
  assign y13790 = ~1'b0 ;
  assign y13791 = ~n1205 ;
  assign y13792 = n25210 ;
  assign y13793 = ~n25212 ;
  assign y13794 = n25214 ;
  assign y13795 = n25218 ;
  assign y13796 = ~1'b0 ;
  assign y13797 = ~n25223 ;
  assign y13798 = ~n25224 ;
  assign y13799 = ~1'b0 ;
  assign y13800 = ~n25230 ;
  assign y13801 = ~n25231 ;
  assign y13802 = ~n25232 ;
  assign y13803 = ~n25234 ;
  assign y13804 = ~n25236 ;
  assign y13805 = ~1'b0 ;
  assign y13806 = ~1'b0 ;
  assign y13807 = ~1'b0 ;
  assign y13808 = 1'b0 ;
  assign y13809 = 1'b0 ;
  assign y13810 = n25237 ;
  assign y13811 = n25241 ;
  assign y13812 = ~1'b0 ;
  assign y13813 = ~n25257 ;
  assign y13814 = ~n25258 ;
  assign y13815 = ~1'b0 ;
  assign y13816 = ~n25259 ;
  assign y13817 = ~n3414 ;
  assign y13818 = ~1'b0 ;
  assign y13819 = ~n1605 ;
  assign y13820 = n25263 ;
  assign y13821 = ~n25269 ;
  assign y13822 = n25270 ;
  assign y13823 = n25271 ;
  assign y13824 = ~1'b0 ;
  assign y13825 = ~n25273 ;
  assign y13826 = n25279 ;
  assign y13827 = n25282 ;
  assign y13828 = ~n25284 ;
  assign y13829 = ~n25291 ;
  assign y13830 = ~n25292 ;
  assign y13831 = ~1'b0 ;
  assign y13832 = n9122 ;
  assign y13833 = ~n6020 ;
  assign y13834 = ~n25293 ;
  assign y13835 = ~n25294 ;
  assign y13836 = n25299 ;
  assign y13837 = ~1'b0 ;
  assign y13838 = 1'b0 ;
  assign y13839 = ~1'b0 ;
  assign y13840 = n25301 ;
  assign y13841 = n25305 ;
  assign y13842 = ~n25309 ;
  assign y13843 = ~n25312 ;
  assign y13844 = n25315 ;
  assign y13845 = n25316 ;
  assign y13846 = ~1'b0 ;
  assign y13847 = ~1'b0 ;
  assign y13848 = ~1'b0 ;
  assign y13849 = ~1'b0 ;
  assign y13850 = ~1'b0 ;
  assign y13851 = n25318 ;
  assign y13852 = ~1'b0 ;
  assign y13853 = n25320 ;
  assign y13854 = n25322 ;
  assign y13855 = ~1'b0 ;
  assign y13856 = ~n25323 ;
  assign y13857 = ~n25325 ;
  assign y13858 = ~n25328 ;
  assign y13859 = ~n25333 ;
  assign y13860 = ~n25336 ;
  assign y13861 = ~1'b0 ;
  assign y13862 = ~1'b0 ;
  assign y13863 = n25337 ;
  assign y13864 = ~n25342 ;
  assign y13865 = ~1'b0 ;
  assign y13866 = ~n25345 ;
  assign y13867 = n25349 ;
  assign y13868 = ~1'b0 ;
  assign y13869 = ~1'b0 ;
  assign y13870 = ~n25351 ;
  assign y13871 = n25355 ;
  assign y13872 = ~1'b0 ;
  assign y13873 = n25356 ;
  assign y13874 = n25360 ;
  assign y13875 = n25364 ;
  assign y13876 = n25365 ;
  assign y13877 = ~n25367 ;
  assign y13878 = ~1'b0 ;
  assign y13879 = ~n25374 ;
  assign y13880 = ~n25375 ;
  assign y13881 = n25378 ;
  assign y13882 = n25381 ;
  assign y13883 = ~1'b0 ;
  assign y13884 = n25393 ;
  assign y13885 = ~n25394 ;
  assign y13886 = ~1'b0 ;
  assign y13887 = ~n25395 ;
  assign y13888 = ~1'b0 ;
  assign y13889 = n25397 ;
  assign y13890 = ~1'b0 ;
  assign y13891 = ~1'b0 ;
  assign y13892 = ~n25401 ;
  assign y13893 = n25404 ;
  assign y13894 = ~n25405 ;
  assign y13895 = ~n25408 ;
  assign y13896 = n25410 ;
  assign y13897 = n25412 ;
  assign y13898 = ~1'b0 ;
  assign y13899 = n25413 ;
  assign y13900 = ~1'b0 ;
  assign y13901 = n25414 ;
  assign y13902 = ~n25415 ;
  assign y13903 = n25417 ;
  assign y13904 = n25418 ;
  assign y13905 = n25420 ;
  assign y13906 = 1'b0 ;
  assign y13907 = n25421 ;
  assign y13908 = n25424 ;
  assign y13909 = 1'b0 ;
  assign y13910 = ~1'b0 ;
  assign y13911 = n25427 ;
  assign y13912 = ~n25433 ;
  assign y13913 = ~1'b0 ;
  assign y13914 = ~n25444 ;
  assign y13915 = n25446 ;
  assign y13916 = ~1'b0 ;
  assign y13917 = n25451 ;
  assign y13918 = n25454 ;
  assign y13919 = ~n25456 ;
  assign y13920 = ~n25459 ;
  assign y13921 = ~n3802 ;
  assign y13922 = n8331 ;
  assign y13923 = n25461 ;
  assign y13924 = ~1'b0 ;
  assign y13925 = ~1'b0 ;
  assign y13926 = ~1'b0 ;
  assign y13927 = n25464 ;
  assign y13928 = ~n25466 ;
  assign y13929 = ~n25468 ;
  assign y13930 = ~n25471 ;
  assign y13931 = ~1'b0 ;
  assign y13932 = ~1'b0 ;
  assign y13933 = ~1'b0 ;
  assign y13934 = ~1'b0 ;
  assign y13935 = n25473 ;
  assign y13936 = ~1'b0 ;
  assign y13937 = ~n25474 ;
  assign y13938 = ~n8819 ;
  assign y13939 = ~n25478 ;
  assign y13940 = n25480 ;
  assign y13941 = ~1'b0 ;
  assign y13942 = n25486 ;
  assign y13943 = ~n10935 ;
  assign y13944 = n25489 ;
  assign y13945 = ~1'b0 ;
  assign y13946 = ~1'b0 ;
  assign y13947 = n16926 ;
  assign y13948 = ~n25490 ;
  assign y13949 = ~1'b0 ;
  assign y13950 = n25491 ;
  assign y13951 = ~1'b0 ;
  assign y13952 = n311 ;
  assign y13953 = ~n25492 ;
  assign y13954 = ~1'b0 ;
  assign y13955 = n25498 ;
  assign y13956 = n11530 ;
  assign y13957 = ~1'b0 ;
  assign y13958 = ~1'b0 ;
  assign y13959 = ~1'b0 ;
  assign y13960 = ~1'b0 ;
  assign y13961 = ~n25503 ;
  assign y13962 = n25507 ;
  assign y13963 = ~n901 ;
  assign y13964 = ~n25508 ;
  assign y13965 = ~1'b0 ;
  assign y13966 = ~1'b0 ;
  assign y13967 = ~1'b0 ;
  assign y13968 = n25509 ;
  assign y13969 = ~1'b0 ;
  assign y13970 = ~1'b0 ;
  assign y13971 = ~1'b0 ;
  assign y13972 = ~n25512 ;
  assign y13973 = ~1'b0 ;
  assign y13974 = n25514 ;
  assign y13975 = n25518 ;
  assign y13976 = ~1'b0 ;
  assign y13977 = n25522 ;
  assign y13978 = ~n25523 ;
  assign y13979 = ~1'b0 ;
  assign y13980 = ~n24423 ;
  assign y13981 = ~n25524 ;
  assign y13982 = n25528 ;
  assign y13983 = n25530 ;
  assign y13984 = 1'b0 ;
  assign y13985 = ~1'b0 ;
  assign y13986 = ~n25531 ;
  assign y13987 = n25532 ;
  assign y13988 = n14577 ;
  assign y13989 = ~n25534 ;
  assign y13990 = ~1'b0 ;
  assign y13991 = n25536 ;
  assign y13992 = ~n25540 ;
  assign y13993 = ~1'b0 ;
  assign y13994 = ~n25548 ;
  assign y13995 = ~1'b0 ;
  assign y13996 = ~n4103 ;
  assign y13997 = n15109 ;
  assign y13998 = n25550 ;
  assign y13999 = n25551 ;
  assign y14000 = ~n25552 ;
  assign y14001 = ~1'b0 ;
  assign y14002 = n25557 ;
  assign y14003 = ~n25558 ;
  assign y14004 = ~n1590 ;
  assign y14005 = ~n25560 ;
  assign y14006 = n6366 ;
  assign y14007 = n25561 ;
  assign y14008 = n25564 ;
  assign y14009 = n25569 ;
  assign y14010 = ~1'b0 ;
  assign y14011 = ~1'b0 ;
  assign y14012 = ~n4370 ;
  assign y14013 = n25570 ;
  assign y14014 = n25574 ;
  assign y14015 = ~n25576 ;
  assign y14016 = n25577 ;
  assign y14017 = ~1'b0 ;
  assign y14018 = ~1'b0 ;
  assign y14019 = ~1'b0 ;
  assign y14020 = ~n25596 ;
  assign y14021 = ~1'b0 ;
  assign y14022 = n25598 ;
  assign y14023 = ~n25599 ;
  assign y14024 = n25601 ;
  assign y14025 = ~n25609 ;
  assign y14026 = n22843 ;
  assign y14027 = ~1'b0 ;
  assign y14028 = ~1'b0 ;
  assign y14029 = ~1'b0 ;
  assign y14030 = n25611 ;
  assign y14031 = n25612 ;
  assign y14032 = n25618 ;
  assign y14033 = ~n9851 ;
  assign y14034 = n25619 ;
  assign y14035 = n25621 ;
  assign y14036 = n25623 ;
  assign y14037 = ~1'b0 ;
  assign y14038 = n25625 ;
  assign y14039 = 1'b0 ;
  assign y14040 = ~n25628 ;
  assign y14041 = n25633 ;
  assign y14042 = ~n25634 ;
  assign y14043 = ~1'b0 ;
  assign y14044 = ~n25640 ;
  assign y14045 = n25645 ;
  assign y14046 = ~1'b0 ;
  assign y14047 = ~1'b0 ;
  assign y14048 = ~n25647 ;
  assign y14049 = 1'b0 ;
  assign y14050 = ~n25648 ;
  assign y14051 = n25649 ;
  assign y14052 = n25651 ;
  assign y14053 = n25653 ;
  assign y14054 = ~1'b0 ;
  assign y14055 = ~n25662 ;
  assign y14056 = 1'b0 ;
  assign y14057 = ~n25666 ;
  assign y14058 = ~1'b0 ;
  assign y14059 = ~1'b0 ;
  assign y14060 = ~1'b0 ;
  assign y14061 = ~n25670 ;
  assign y14062 = ~n25675 ;
  assign y14063 = n25676 ;
  assign y14064 = ~1'b0 ;
  assign y14065 = n25677 ;
  assign y14066 = ~n25682 ;
  assign y14067 = ~1'b0 ;
  assign y14068 = n25687 ;
  assign y14069 = n25690 ;
  assign y14070 = ~1'b0 ;
  assign y14071 = ~1'b0 ;
  assign y14072 = n25691 ;
  assign y14073 = ~1'b0 ;
  assign y14074 = ~n25696 ;
  assign y14075 = ~1'b0 ;
  assign y14076 = ~n25699 ;
  assign y14077 = ~1'b0 ;
  assign y14078 = n1814 ;
  assign y14079 = n25700 ;
  assign y14080 = n25702 ;
  assign y14081 = n25707 ;
  assign y14082 = ~n25708 ;
  assign y14083 = ~n25709 ;
  assign y14084 = ~1'b0 ;
  assign y14085 = ~n25712 ;
  assign y14086 = n25715 ;
  assign y14087 = ~n25720 ;
  assign y14088 = ~n25722 ;
  assign y14089 = ~1'b0 ;
  assign y14090 = ~n25727 ;
  assign y14091 = ~1'b0 ;
  assign y14092 = n25735 ;
  assign y14093 = ~n8365 ;
  assign y14094 = ~1'b0 ;
  assign y14095 = ~n25737 ;
  assign y14096 = ~1'b0 ;
  assign y14097 = ~n511 ;
  assign y14098 = n25740 ;
  assign y14099 = ~1'b0 ;
  assign y14100 = n11563 ;
  assign y14101 = ~n25741 ;
  assign y14102 = n25747 ;
  assign y14103 = ~1'b0 ;
  assign y14104 = ~1'b0 ;
  assign y14105 = ~1'b0 ;
  assign y14106 = ~n25750 ;
  assign y14107 = n25752 ;
  assign y14108 = ~n25754 ;
  assign y14109 = ~1'b0 ;
  assign y14110 = ~n25756 ;
  assign y14111 = n25760 ;
  assign y14112 = n25761 ;
  assign y14113 = ~n25762 ;
  assign y14114 = ~1'b0 ;
  assign y14115 = ~1'b0 ;
  assign y14116 = ~n25763 ;
  assign y14117 = n25766 ;
  assign y14118 = ~n25769 ;
  assign y14119 = ~1'b0 ;
  assign y14120 = n25771 ;
  assign y14121 = n17201 ;
  assign y14122 = ~1'b0 ;
  assign y14123 = n7763 ;
  assign y14124 = ~n25772 ;
  assign y14125 = n16048 ;
  assign y14126 = ~1'b0 ;
  assign y14127 = n25773 ;
  assign y14128 = n23908 ;
  assign y14129 = ~n25780 ;
  assign y14130 = n1786 ;
  assign y14131 = ~n25784 ;
  assign y14132 = ~n13787 ;
  assign y14133 = ~1'b0 ;
  assign y14134 = n25786 ;
  assign y14135 = n25789 ;
  assign y14136 = n25796 ;
  assign y14137 = n25799 ;
  assign y14138 = n25801 ;
  assign y14139 = ~n25805 ;
  assign y14140 = ~n25808 ;
  assign y14141 = n25809 ;
  assign y14142 = n25810 ;
  assign y14143 = ~1'b0 ;
  assign y14144 = ~n25812 ;
  assign y14145 = ~1'b0 ;
  assign y14146 = n25819 ;
  assign y14147 = ~1'b0 ;
  assign y14148 = ~1'b0 ;
  assign y14149 = ~n25820 ;
  assign y14150 = n25829 ;
  assign y14151 = ~1'b0 ;
  assign y14152 = ~1'b0 ;
  assign y14153 = ~n25831 ;
  assign y14154 = ~1'b0 ;
  assign y14155 = ~1'b0 ;
  assign y14156 = n25848 ;
  assign y14157 = ~1'b0 ;
  assign y14158 = ~1'b0 ;
  assign y14159 = ~1'b0 ;
  assign y14160 = ~n24326 ;
  assign y14161 = ~1'b0 ;
  assign y14162 = ~n8555 ;
  assign y14163 = ~n25849 ;
  assign y14164 = ~1'b0 ;
  assign y14165 = ~1'b0 ;
  assign y14166 = ~1'b0 ;
  assign y14167 = ~1'b0 ;
  assign y14168 = n25850 ;
  assign y14169 = ~n25853 ;
  assign y14170 = ~n25857 ;
  assign y14171 = ~n25858 ;
  assign y14172 = ~1'b0 ;
  assign y14173 = ~1'b0 ;
  assign y14174 = ~1'b0 ;
  assign y14175 = ~1'b0 ;
  assign y14176 = ~1'b0 ;
  assign y14177 = ~n25859 ;
  assign y14178 = 1'b0 ;
  assign y14179 = ~1'b0 ;
  assign y14180 = ~1'b0 ;
  assign y14181 = n25860 ;
  assign y14182 = ~n25865 ;
  assign y14183 = ~n25455 ;
  assign y14184 = ~1'b0 ;
  assign y14185 = ~n25867 ;
  assign y14186 = ~1'b0 ;
  assign y14187 = n25868 ;
  assign y14188 = ~1'b0 ;
  assign y14189 = n25876 ;
  assign y14190 = ~n25877 ;
  assign y14191 = ~n25879 ;
  assign y14192 = n25884 ;
  assign y14193 = n25887 ;
  assign y14194 = ~1'b0 ;
  assign y14195 = n25888 ;
  assign y14196 = ~1'b0 ;
  assign y14197 = ~n25893 ;
  assign y14198 = ~n25896 ;
  assign y14199 = ~1'b0 ;
  assign y14200 = n25899 ;
  assign y14201 = ~1'b0 ;
  assign y14202 = n25901 ;
  assign y14203 = ~1'b0 ;
  assign y14204 = ~n25902 ;
  assign y14205 = ~1'b0 ;
  assign y14206 = ~1'b0 ;
  assign y14207 = ~n25903 ;
  assign y14208 = n25904 ;
  assign y14209 = n25905 ;
  assign y14210 = n25906 ;
  assign y14211 = n25908 ;
  assign y14212 = ~1'b0 ;
  assign y14213 = ~1'b0 ;
  assign y14214 = ~n25909 ;
  assign y14215 = n25910 ;
  assign y14216 = n25911 ;
  assign y14217 = ~n25914 ;
  assign y14218 = ~1'b0 ;
  assign y14219 = ~n25921 ;
  assign y14220 = ~n25922 ;
  assign y14221 = n25924 ;
  assign y14222 = ~1'b0 ;
  assign y14223 = ~n25925 ;
  assign y14224 = ~n25926 ;
  assign y14225 = ~n25931 ;
  assign y14226 = ~n25935 ;
  assign y14227 = ~n25937 ;
  assign y14228 = ~n25938 ;
  assign y14229 = n17123 ;
  assign y14230 = ~1'b0 ;
  assign y14231 = n25941 ;
  assign y14232 = ~1'b0 ;
  assign y14233 = n15712 ;
  assign y14234 = ~n25943 ;
  assign y14235 = ~1'b0 ;
  assign y14236 = ~n2387 ;
  assign y14237 = ~n25944 ;
  assign y14238 = ~n25945 ;
  assign y14239 = n25946 ;
  assign y14240 = ~n25951 ;
  assign y14241 = ~1'b0 ;
  assign y14242 = ~1'b0 ;
  assign y14243 = ~n20335 ;
  assign y14244 = n25955 ;
  assign y14245 = ~n25957 ;
  assign y14246 = ~1'b0 ;
  assign y14247 = n25960 ;
  assign y14248 = ~n25962 ;
  assign y14249 = ~n25963 ;
  assign y14250 = ~1'b0 ;
  assign y14251 = n25964 ;
  assign y14252 = ~1'b0 ;
  assign y14253 = ~1'b0 ;
  assign y14254 = ~n25969 ;
  assign y14255 = ~1'b0 ;
  assign y14256 = ~1'b0 ;
  assign y14257 = n25972 ;
  assign y14258 = n540 ;
  assign y14259 = ~n25975 ;
  assign y14260 = ~1'b0 ;
  assign y14261 = n25976 ;
  assign y14262 = ~n4666 ;
  assign y14263 = ~1'b0 ;
  assign y14264 = ~n25977 ;
  assign y14265 = ~1'b0 ;
  assign y14266 = ~1'b0 ;
  assign y14267 = n25980 ;
  assign y14268 = n25983 ;
  assign y14269 = ~1'b0 ;
  assign y14270 = ~n25995 ;
  assign y14271 = n15925 ;
  assign y14272 = n25997 ;
  assign y14273 = n26000 ;
  assign y14274 = ~n26004 ;
  assign y14275 = ~1'b0 ;
  assign y14276 = n26007 ;
  assign y14277 = ~n26008 ;
  assign y14278 = n26009 ;
  assign y14279 = n26011 ;
  assign y14280 = ~n26012 ;
  assign y14281 = ~1'b0 ;
  assign y14282 = ~1'b0 ;
  assign y14283 = ~1'b0 ;
  assign y14284 = n11813 ;
  assign y14285 = n26015 ;
  assign y14286 = ~1'b0 ;
  assign y14287 = ~n26019 ;
  assign y14288 = n26022 ;
  assign y14289 = ~1'b0 ;
  assign y14290 = ~1'b0 ;
  assign y14291 = n26026 ;
  assign y14292 = n26027 ;
  assign y14293 = n26028 ;
  assign y14294 = n26030 ;
  assign y14295 = 1'b0 ;
  assign y14296 = n26032 ;
  assign y14297 = ~n26035 ;
  assign y14298 = n26041 ;
  assign y14299 = 1'b0 ;
  assign y14300 = ~1'b0 ;
  assign y14301 = ~1'b0 ;
  assign y14302 = ~n26042 ;
  assign y14303 = ~1'b0 ;
  assign y14304 = n25351 ;
  assign y14305 = ~1'b0 ;
  assign y14306 = n26044 ;
  assign y14307 = ~1'b0 ;
  assign y14308 = ~n13734 ;
  assign y14309 = ~n26050 ;
  assign y14310 = ~n26051 ;
  assign y14311 = n26059 ;
  assign y14312 = ~n26062 ;
  assign y14313 = ~1'b0 ;
  assign y14314 = ~1'b0 ;
  assign y14315 = ~1'b0 ;
  assign y14316 = ~1'b0 ;
  assign y14317 = ~1'b0 ;
  assign y14318 = ~1'b0 ;
  assign y14319 = n13096 ;
  assign y14320 = n26063 ;
  assign y14321 = ~n26070 ;
  assign y14322 = n26074 ;
  assign y14323 = ~n26075 ;
  assign y14324 = ~n26076 ;
  assign y14325 = ~n26085 ;
  assign y14326 = ~n26093 ;
  assign y14327 = ~1'b0 ;
  assign y14328 = n26095 ;
  assign y14329 = n26097 ;
  assign y14330 = ~n26103 ;
  assign y14331 = ~1'b0 ;
  assign y14332 = ~n26104 ;
  assign y14333 = n26105 ;
  assign y14334 = ~n26106 ;
  assign y14335 = n18910 ;
  assign y14336 = n26108 ;
  assign y14337 = n26109 ;
  assign y14338 = ~n26111 ;
  assign y14339 = n26112 ;
  assign y14340 = ~n1644 ;
  assign y14341 = n26113 ;
  assign y14342 = n26115 ;
  assign y14343 = ~n26116 ;
  assign y14344 = ~1'b0 ;
  assign y14345 = ~n5008 ;
  assign y14346 = ~1'b0 ;
  assign y14347 = 1'b0 ;
  assign y14348 = n26121 ;
  assign y14349 = ~n26122 ;
  assign y14350 = ~1'b0 ;
  assign y14351 = n26124 ;
  assign y14352 = ~n26127 ;
  assign y14353 = ~n26128 ;
  assign y14354 = ~1'b0 ;
  assign y14355 = ~n20233 ;
  assign y14356 = n26129 ;
  assign y14357 = n26131 ;
  assign y14358 = ~1'b0 ;
  assign y14359 = ~1'b0 ;
  assign y14360 = ~n26133 ;
  assign y14361 = ~n26134 ;
  assign y14362 = n26136 ;
  assign y14363 = ~n26137 ;
  assign y14364 = ~n7755 ;
  assign y14365 = ~1'b0 ;
  assign y14366 = ~n26140 ;
  assign y14367 = n26141 ;
  assign y14368 = n26142 ;
  assign y14369 = ~n26143 ;
  assign y14370 = n26151 ;
  assign y14371 = n21534 ;
  assign y14372 = ~n26152 ;
  assign y14373 = n26154 ;
  assign y14374 = n26156 ;
  assign y14375 = ~n26162 ;
  assign y14376 = n26163 ;
  assign y14377 = n26166 ;
  assign y14378 = n26168 ;
  assign y14379 = n26171 ;
  assign y14380 = ~1'b0 ;
  assign y14381 = n26172 ;
  assign y14382 = n26176 ;
  assign y14383 = ~n26181 ;
  assign y14384 = n26184 ;
  assign y14385 = ~1'b0 ;
  assign y14386 = ~1'b0 ;
  assign y14387 = n26185 ;
  assign y14388 = n26187 ;
  assign y14389 = n26190 ;
  assign y14390 = ~1'b0 ;
  assign y14391 = ~1'b0 ;
  assign y14392 = ~n17433 ;
  assign y14393 = 1'b0 ;
  assign y14394 = ~1'b0 ;
  assign y14395 = ~1'b0 ;
  assign y14396 = ~1'b0 ;
  assign y14397 = ~n26195 ;
  assign y14398 = ~n26198 ;
  assign y14399 = ~n26199 ;
  assign y14400 = ~n26201 ;
  assign y14401 = ~1'b0 ;
  assign y14402 = ~n26204 ;
  assign y14403 = ~n26206 ;
  assign y14404 = ~n26209 ;
  assign y14405 = n26214 ;
  assign y14406 = ~1'b0 ;
  assign y14407 = ~n26216 ;
  assign y14408 = ~n4226 ;
  assign y14409 = ~1'b0 ;
  assign y14410 = ~1'b0 ;
  assign y14411 = ~1'b0 ;
  assign y14412 = ~n10950 ;
  assign y14413 = 1'b0 ;
  assign y14414 = n26219 ;
  assign y14415 = ~n26221 ;
  assign y14416 = n26227 ;
  assign y14417 = ~n26237 ;
  assign y14418 = ~1'b0 ;
  assign y14419 = ~n26241 ;
  assign y14420 = ~n26242 ;
  assign y14421 = ~n8239 ;
  assign y14422 = ~1'b0 ;
  assign y14423 = ~1'b0 ;
  assign y14424 = n26244 ;
  assign y14425 = ~1'b0 ;
  assign y14426 = ~n26245 ;
  assign y14427 = ~1'b0 ;
  assign y14428 = 1'b0 ;
  assign y14429 = ~1'b0 ;
  assign y14430 = ~n9377 ;
  assign y14431 = n26251 ;
  assign y14432 = n26253 ;
  assign y14433 = ~n21004 ;
  assign y14434 = ~1'b0 ;
  assign y14435 = 1'b0 ;
  assign y14436 = n26259 ;
  assign y14437 = ~n26272 ;
  assign y14438 = n26276 ;
  assign y14439 = ~n26279 ;
  assign y14440 = ~n26281 ;
  assign y14441 = ~n26283 ;
  assign y14442 = n26285 ;
  assign y14443 = n25408 ;
  assign y14444 = n26290 ;
  assign y14445 = n26291 ;
  assign y14446 = ~n26295 ;
  assign y14447 = ~n26296 ;
  assign y14448 = ~1'b0 ;
  assign y14449 = n6702 ;
  assign y14450 = n26303 ;
  assign y14451 = n3472 ;
  assign y14452 = ~n26304 ;
  assign y14453 = ~1'b0 ;
  assign y14454 = ~n26306 ;
  assign y14455 = ~1'b0 ;
  assign y14456 = ~1'b0 ;
  assign y14457 = n26307 ;
  assign y14458 = ~1'b0 ;
  assign y14459 = ~n26311 ;
  assign y14460 = ~1'b0 ;
  assign y14461 = ~n26317 ;
  assign y14462 = n26321 ;
  assign y14463 = ~1'b0 ;
  assign y14464 = ~n26325 ;
  assign y14465 = n26327 ;
  assign y14466 = n26328 ;
  assign y14467 = n26332 ;
  assign y14468 = ~1'b0 ;
  assign y14469 = n26333 ;
  assign y14470 = ~1'b0 ;
  assign y14471 = n26335 ;
  assign y14472 = ~n26337 ;
  assign y14473 = n26338 ;
  assign y14474 = ~1'b0 ;
  assign y14475 = ~1'b0 ;
  assign y14476 = ~n26341 ;
  assign y14477 = ~n26342 ;
  assign y14478 = ~1'b0 ;
  assign y14479 = ~1'b0 ;
  assign y14480 = n26344 ;
  assign y14481 = ~n26348 ;
  assign y14482 = n26349 ;
  assign y14483 = ~n26351 ;
  assign y14484 = ~n26352 ;
  assign y14485 = 1'b0 ;
  assign y14486 = ~1'b0 ;
  assign y14487 = ~1'b0 ;
  assign y14488 = n820 ;
  assign y14489 = ~n26354 ;
  assign y14490 = ~n26355 ;
  assign y14491 = n26363 ;
  assign y14492 = ~n26366 ;
  assign y14493 = ~1'b0 ;
  assign y14494 = ~n26371 ;
  assign y14495 = ~1'b0 ;
  assign y14496 = n26373 ;
  assign y14497 = n26374 ;
  assign y14498 = n10389 ;
  assign y14499 = ~1'b0 ;
  assign y14500 = n26375 ;
  assign y14501 = n26379 ;
  assign y14502 = ~n26385 ;
  assign y14503 = n26387 ;
  assign y14504 = n26388 ;
  assign y14505 = n26389 ;
  assign y14506 = ~n26391 ;
  assign y14507 = ~1'b0 ;
  assign y14508 = n26397 ;
  assign y14509 = n26408 ;
  assign y14510 = ~n26409 ;
  assign y14511 = n6794 ;
  assign y14512 = ~n26410 ;
  assign y14513 = 1'b0 ;
  assign y14514 = ~1'b0 ;
  assign y14515 = ~1'b0 ;
  assign y14516 = ~n26415 ;
  assign y14517 = n26418 ;
  assign y14518 = n11285 ;
  assign y14519 = ~1'b0 ;
  assign y14520 = n26420 ;
  assign y14521 = ~1'b0 ;
  assign y14522 = ~1'b0 ;
  assign y14523 = ~1'b0 ;
  assign y14524 = n26421 ;
  assign y14525 = ~1'b0 ;
  assign y14526 = ~n26426 ;
  assign y14527 = ~n26433 ;
  assign y14528 = ~n26434 ;
  assign y14529 = n26448 ;
  assign y14530 = n26449 ;
  assign y14531 = ~n26455 ;
  assign y14532 = ~n11759 ;
  assign y14533 = ~1'b0 ;
  assign y14534 = n26456 ;
  assign y14535 = n22161 ;
  assign y14536 = ~n8761 ;
  assign y14537 = n26457 ;
  assign y14538 = ~n26459 ;
  assign y14539 = ~1'b0 ;
  assign y14540 = ~1'b0 ;
  assign y14541 = ~1'b0 ;
  assign y14542 = ~n26466 ;
  assign y14543 = ~1'b0 ;
  assign y14544 = n26468 ;
  assign y14545 = ~n26469 ;
  assign y14546 = ~n26471 ;
  assign y14547 = ~1'b0 ;
  assign y14548 = ~n26473 ;
  assign y14549 = n17294 ;
  assign y14550 = ~n26475 ;
  assign y14551 = ~1'b0 ;
  assign y14552 = ~n26478 ;
  assign y14553 = ~n26484 ;
  assign y14554 = ~1'b0 ;
  assign y14555 = ~n26485 ;
  assign y14556 = n26486 ;
  assign y14557 = n26487 ;
  assign y14558 = n26489 ;
  assign y14559 = ~n26490 ;
  assign y14560 = n26492 ;
  assign y14561 = ~1'b0 ;
  assign y14562 = ~n26493 ;
  assign y14563 = n26494 ;
  assign y14564 = ~1'b0 ;
  assign y14565 = n26496 ;
  assign y14566 = n26498 ;
  assign y14567 = n26502 ;
  assign y14568 = ~n26504 ;
  assign y14569 = ~n9267 ;
  assign y14570 = ~n17640 ;
  assign y14571 = ~n26505 ;
  assign y14572 = ~1'b0 ;
  assign y14573 = n4991 ;
  assign y14574 = ~1'b0 ;
  assign y14575 = ~1'b0 ;
  assign y14576 = ~1'b0 ;
  assign y14577 = ~n26506 ;
  assign y14578 = n26514 ;
  assign y14579 = n8738 ;
  assign y14580 = n15135 ;
  assign y14581 = n26516 ;
  assign y14582 = ~n12217 ;
  assign y14583 = n12197 ;
  assign y14584 = ~1'b0 ;
  assign y14585 = ~n26519 ;
  assign y14586 = n19991 ;
  assign y14587 = ~1'b0 ;
  assign y14588 = n26522 ;
  assign y14589 = ~1'b0 ;
  assign y14590 = n26524 ;
  assign y14591 = ~1'b0 ;
  assign y14592 = ~n26525 ;
  assign y14593 = ~1'b0 ;
  assign y14594 = ~1'b0 ;
  assign y14595 = ~1'b0 ;
  assign y14596 = n26527 ;
  assign y14597 = ~1'b0 ;
  assign y14598 = n26529 ;
  assign y14599 = ~1'b0 ;
  assign y14600 = n26531 ;
  assign y14601 = ~n14458 ;
  assign y14602 = ~1'b0 ;
  assign y14603 = ~1'b0 ;
  assign y14604 = n26537 ;
  assign y14605 = ~1'b0 ;
  assign y14606 = ~n26541 ;
  assign y14607 = ~1'b0 ;
  assign y14608 = n26545 ;
  assign y14609 = n26546 ;
  assign y14610 = n26550 ;
  assign y14611 = ~1'b0 ;
  assign y14612 = n26556 ;
  assign y14613 = n26559 ;
  assign y14614 = n26562 ;
  assign y14615 = ~n26564 ;
  assign y14616 = ~n26566 ;
  assign y14617 = ~1'b0 ;
  assign y14618 = 1'b0 ;
  assign y14619 = n26572 ;
  assign y14620 = ~1'b0 ;
  assign y14621 = n26574 ;
  assign y14622 = n26575 ;
  assign y14623 = n26584 ;
  assign y14624 = ~n1201 ;
  assign y14625 = ~1'b0 ;
  assign y14626 = ~1'b0 ;
  assign y14627 = ~n1176 ;
  assign y14628 = ~n26585 ;
  assign y14629 = n26586 ;
  assign y14630 = ~n26587 ;
  assign y14631 = ~n26588 ;
  assign y14632 = ~n26589 ;
  assign y14633 = n26593 ;
  assign y14634 = n26597 ;
  assign y14635 = ~1'b0 ;
  assign y14636 = n26598 ;
  assign y14637 = ~1'b0 ;
  assign y14638 = ~1'b0 ;
  assign y14639 = ~1'b0 ;
  assign y14640 = ~n26599 ;
  assign y14641 = ~n10425 ;
  assign y14642 = n26600 ;
  assign y14643 = ~n26602 ;
  assign y14644 = ~1'b0 ;
  assign y14645 = ~n26606 ;
  assign y14646 = ~n26607 ;
  assign y14647 = n26610 ;
  assign y14648 = ~n26612 ;
  assign y14649 = ~1'b0 ;
  assign y14650 = ~n26616 ;
  assign y14651 = ~n26618 ;
  assign y14652 = ~1'b0 ;
  assign y14653 = ~n26619 ;
  assign y14654 = ~1'b0 ;
  assign y14655 = n19281 ;
  assign y14656 = ~1'b0 ;
  assign y14657 = n18383 ;
  assign y14658 = n26620 ;
  assign y14659 = ~n26621 ;
  assign y14660 = n26624 ;
  assign y14661 = ~1'b0 ;
  assign y14662 = n26625 ;
  assign y14663 = n26627 ;
  assign y14664 = ~n26630 ;
  assign y14665 = ~1'b0 ;
  assign y14666 = ~1'b0 ;
  assign y14667 = ~n26632 ;
  assign y14668 = n26639 ;
  assign y14669 = ~n26641 ;
  assign y14670 = n26644 ;
  assign y14671 = n26651 ;
  assign y14672 = n26653 ;
  assign y14673 = n9731 ;
  assign y14674 = n26657 ;
  assign y14675 = n26660 ;
  assign y14676 = n26662 ;
  assign y14677 = n26664 ;
  assign y14678 = ~1'b0 ;
  assign y14679 = n26668 ;
  assign y14680 = ~1'b0 ;
  assign y14681 = ~1'b0 ;
  assign y14682 = ~n26670 ;
  assign y14683 = n26673 ;
  assign y14684 = ~n26676 ;
  assign y14685 = ~1'b0 ;
  assign y14686 = ~n26677 ;
  assign y14687 = ~n26678 ;
  assign y14688 = ~1'b0 ;
  assign y14689 = n26679 ;
  assign y14690 = ~n26684 ;
  assign y14691 = n26686 ;
  assign y14692 = ~1'b0 ;
  assign y14693 = ~n26688 ;
  assign y14694 = ~n26693 ;
  assign y14695 = n26695 ;
  assign y14696 = n26698 ;
  assign y14697 = ~1'b0 ;
  assign y14698 = ~n26704 ;
  assign y14699 = ~1'b0 ;
  assign y14700 = ~n26712 ;
  assign y14701 = ~1'b0 ;
  assign y14702 = n26716 ;
  assign y14703 = ~n26720 ;
  assign y14704 = n26722 ;
  assign y14705 = ~n26723 ;
  assign y14706 = n26724 ;
  assign y14707 = ~1'b0 ;
  assign y14708 = ~n26725 ;
  assign y14709 = ~1'b0 ;
  assign y14710 = n26731 ;
  assign y14711 = ~1'b0 ;
  assign y14712 = n26732 ;
  assign y14713 = ~n26737 ;
  assign y14714 = ~1'b0 ;
  assign y14715 = ~1'b0 ;
  assign y14716 = n26738 ;
  assign y14717 = n26739 ;
  assign y14718 = ~n26740 ;
  assign y14719 = ~1'b0 ;
  assign y14720 = n26745 ;
  assign y14721 = ~1'b0 ;
  assign y14722 = ~1'b0 ;
  assign y14723 = n26746 ;
  assign y14724 = n26750 ;
  assign y14725 = ~n26751 ;
  assign y14726 = ~n26752 ;
  assign y14727 = n26754 ;
  assign y14728 = ~n26760 ;
  assign y14729 = n26761 ;
  assign y14730 = ~1'b0 ;
  assign y14731 = n26763 ;
  assign y14732 = ~n26768 ;
  assign y14733 = n22600 ;
  assign y14734 = ~1'b0 ;
  assign y14735 = n26773 ;
  assign y14736 = ~n26774 ;
  assign y14737 = 1'b0 ;
  assign y14738 = n26775 ;
  assign y14739 = n26778 ;
  assign y14740 = ~n26779 ;
  assign y14741 = ~n26782 ;
  assign y14742 = n26789 ;
  assign y14743 = ~1'b0 ;
  assign y14744 = n26790 ;
  assign y14745 = ~n26792 ;
  assign y14746 = ~1'b0 ;
  assign y14747 = ~n468 ;
  assign y14748 = n26798 ;
  assign y14749 = n26072 ;
  assign y14750 = ~n26801 ;
  assign y14751 = ~n26803 ;
  assign y14752 = ~n26807 ;
  assign y14753 = ~1'b0 ;
  assign y14754 = n26814 ;
  assign y14755 = n26820 ;
  assign y14756 = ~1'b0 ;
  assign y14757 = n26821 ;
  assign y14758 = n4001 ;
  assign y14759 = ~1'b0 ;
  assign y14760 = n26822 ;
  assign y14761 = n11442 ;
  assign y14762 = n26824 ;
  assign y14763 = ~1'b0 ;
  assign y14764 = n26825 ;
  assign y14765 = n26826 ;
  assign y14766 = ~1'b0 ;
  assign y14767 = n26829 ;
  assign y14768 = ~1'b0 ;
  assign y14769 = n15660 ;
  assign y14770 = n26830 ;
  assign y14771 = ~1'b0 ;
  assign y14772 = ~n26834 ;
  assign y14773 = n26835 ;
  assign y14774 = ~n26836 ;
  assign y14775 = n26839 ;
  assign y14776 = ~n26844 ;
  assign y14777 = ~1'b0 ;
  assign y14778 = n22599 ;
  assign y14779 = ~n26846 ;
  assign y14780 = ~1'b0 ;
  assign y14781 = ~1'b0 ;
  assign y14782 = ~n26848 ;
  assign y14783 = n26851 ;
  assign y14784 = ~n8141 ;
  assign y14785 = 1'b0 ;
  assign y14786 = ~n22671 ;
  assign y14787 = ~n26854 ;
  assign y14788 = ~n26858 ;
  assign y14789 = ~n26863 ;
  assign y14790 = ~1'b0 ;
  assign y14791 = ~n26865 ;
  assign y14792 = n26874 ;
  assign y14793 = n26875 ;
  assign y14794 = ~n26876 ;
  assign y14795 = ~n26878 ;
  assign y14796 = n26879 ;
  assign y14797 = n26881 ;
  assign y14798 = ~n21191 ;
  assign y14799 = ~n3547 ;
  assign y14800 = n26882 ;
  assign y14801 = n26885 ;
  assign y14802 = n10828 ;
  assign y14803 = n26889 ;
  assign y14804 = ~n11269 ;
  assign y14805 = ~n26890 ;
  assign y14806 = ~n26892 ;
  assign y14807 = ~1'b0 ;
  assign y14808 = ~1'b0 ;
  assign y14809 = ~n26895 ;
  assign y14810 = n26898 ;
  assign y14811 = ~1'b0 ;
  assign y14812 = ~1'b0 ;
  assign y14813 = ~n26899 ;
  assign y14814 = n26901 ;
  assign y14815 = ~n26902 ;
  assign y14816 = ~1'b0 ;
  assign y14817 = ~1'b0 ;
  assign y14818 = ~n26905 ;
  assign y14819 = ~n26907 ;
  assign y14820 = n24384 ;
  assign y14821 = ~n26910 ;
  assign y14822 = n26912 ;
  assign y14823 = n26915 ;
  assign y14824 = n1227 ;
  assign y14825 = ~1'b0 ;
  assign y14826 = ~n26917 ;
  assign y14827 = ~n26919 ;
  assign y14828 = ~1'b0 ;
  assign y14829 = n26922 ;
  assign y14830 = ~n26923 ;
  assign y14831 = n26924 ;
  assign y14832 = ~1'b0 ;
  assign y14833 = ~1'b0 ;
  assign y14834 = n26927 ;
  assign y14835 = n26930 ;
  assign y14836 = n26931 ;
  assign y14837 = ~n26935 ;
  assign y14838 = ~n26938 ;
  assign y14839 = ~n220 ;
  assign y14840 = n26007 ;
  assign y14841 = n26946 ;
  assign y14842 = n26948 ;
  assign y14843 = 1'b0 ;
  assign y14844 = 1'b0 ;
  assign y14845 = n26949 ;
  assign y14846 = ~1'b0 ;
  assign y14847 = ~1'b0 ;
  assign y14848 = n26951 ;
  assign y14849 = n26952 ;
  assign y14850 = n26959 ;
  assign y14851 = ~n26960 ;
  assign y14852 = n26962 ;
  assign y14853 = n8503 ;
  assign y14854 = n26965 ;
  assign y14855 = ~n26969 ;
  assign y14856 = ~1'b0 ;
  assign y14857 = ~1'b0 ;
  assign y14858 = n26972 ;
  assign y14859 = ~n16563 ;
  assign y14860 = ~1'b0 ;
  assign y14861 = ~1'b0 ;
  assign y14862 = n26974 ;
  assign y14863 = n26975 ;
  assign y14864 = ~n26980 ;
  assign y14865 = ~n26986 ;
  assign y14866 = ~1'b0 ;
  assign y14867 = ~1'b0 ;
  assign y14868 = ~n26987 ;
  assign y14869 = ~1'b0 ;
  assign y14870 = 1'b0 ;
  assign y14871 = ~n26988 ;
  assign y14872 = ~1'b0 ;
  assign y14873 = ~1'b0 ;
  assign y14874 = n26989 ;
  assign y14875 = ~1'b0 ;
  assign y14876 = ~1'b0 ;
  assign y14877 = ~1'b0 ;
  assign y14878 = n26992 ;
  assign y14879 = ~n3031 ;
  assign y14880 = ~n14378 ;
  assign y14881 = ~n26995 ;
  assign y14882 = ~n27000 ;
  assign y14883 = ~1'b0 ;
  assign y14884 = ~1'b0 ;
  assign y14885 = n7902 ;
  assign y14886 = ~1'b0 ;
  assign y14887 = ~1'b0 ;
  assign y14888 = n27002 ;
  assign y14889 = ~1'b0 ;
  assign y14890 = n27004 ;
  assign y14891 = n27005 ;
  assign y14892 = n27011 ;
  assign y14893 = n376 ;
  assign y14894 = n10552 ;
  assign y14895 = n27013 ;
  assign y14896 = ~n2453 ;
  assign y14897 = ~n27015 ;
  assign y14898 = ~n27017 ;
  assign y14899 = n27018 ;
  assign y14900 = ~n27021 ;
  assign y14901 = n27025 ;
  assign y14902 = ~n27026 ;
  assign y14903 = ~n27027 ;
  assign y14904 = ~1'b0 ;
  assign y14905 = ~1'b0 ;
  assign y14906 = n27032 ;
  assign y14907 = ~n25759 ;
  assign y14908 = n27034 ;
  assign y14909 = n27035 ;
  assign y14910 = ~n27040 ;
  assign y14911 = n27045 ;
  assign y14912 = ~n6399 ;
  assign y14913 = n27048 ;
  assign y14914 = n27051 ;
  assign y14915 = 1'b0 ;
  assign y14916 = n27055 ;
  assign y14917 = n17940 ;
  assign y14918 = 1'b0 ;
  assign y14919 = n27056 ;
  assign y14920 = ~1'b0 ;
  assign y14921 = n27058 ;
  assign y14922 = n27062 ;
  assign y14923 = n27063 ;
  assign y14924 = n27065 ;
  assign y14925 = ~n27068 ;
  assign y14926 = n27072 ;
  assign y14927 = ~n27074 ;
  assign y14928 = 1'b0 ;
  assign y14929 = n27077 ;
  assign y14930 = n27078 ;
  assign y14931 = 1'b0 ;
  assign y14932 = ~n27083 ;
  assign y14933 = n27085 ;
  assign y14934 = n27087 ;
  assign y14935 = ~n27090 ;
  assign y14936 = ~n27096 ;
  assign y14937 = n27097 ;
  assign y14938 = n27098 ;
  assign y14939 = n25981 ;
  assign y14940 = ~1'b0 ;
  assign y14941 = ~1'b0 ;
  assign y14942 = n27101 ;
  assign y14943 = ~n27107 ;
  assign y14944 = ~n27111 ;
  assign y14945 = ~n27113 ;
  assign y14946 = ~n27116 ;
  assign y14947 = n27121 ;
  assign y14948 = ~1'b0 ;
  assign y14949 = ~n27123 ;
  assign y14950 = n14658 ;
  assign y14951 = n27125 ;
  assign y14952 = n27127 ;
  assign y14953 = ~n27128 ;
  assign y14954 = n27131 ;
  assign y14955 = n27133 ;
  assign y14956 = ~n27134 ;
  assign y14957 = ~1'b0 ;
  assign y14958 = n27135 ;
  assign y14959 = n27136 ;
  assign y14960 = ~1'b0 ;
  assign y14961 = n27138 ;
  assign y14962 = ~n27140 ;
  assign y14963 = n21460 ;
  assign y14964 = n27141 ;
  assign y14965 = ~n27143 ;
  assign y14966 = ~n27157 ;
  assign y14967 = ~n27158 ;
  assign y14968 = ~1'b0 ;
  assign y14969 = n27169 ;
  assign y14970 = ~n27171 ;
  assign y14971 = n27174 ;
  assign y14972 = ~n27176 ;
  assign y14973 = n27179 ;
  assign y14974 = 1'b0 ;
  assign y14975 = ~1'b0 ;
  assign y14976 = n16257 ;
  assign y14977 = ~n27182 ;
  assign y14978 = ~1'b0 ;
  assign y14979 = ~1'b0 ;
  assign y14980 = ~1'b0 ;
  assign y14981 = ~1'b0 ;
  assign y14982 = n27184 ;
  assign y14983 = ~n27190 ;
  assign y14984 = n27197 ;
  assign y14985 = ~1'b0 ;
  assign y14986 = ~n27200 ;
  assign y14987 = ~1'b0 ;
  assign y14988 = ~n27202 ;
  assign y14989 = ~n27203 ;
  assign y14990 = ~1'b0 ;
  assign y14991 = ~1'b0 ;
  assign y14992 = ~n27204 ;
  assign y14993 = n27211 ;
  assign y14994 = ~1'b0 ;
  assign y14995 = ~n27216 ;
  assign y14996 = ~n27224 ;
  assign y14997 = ~n27225 ;
  assign y14998 = ~1'b0 ;
  assign y14999 = n27226 ;
  assign y15000 = ~1'b0 ;
  assign y15001 = ~n27232 ;
  assign y15002 = ~1'b0 ;
  assign y15003 = ~1'b0 ;
  assign y15004 = ~1'b0 ;
  assign y15005 = n26 ;
  assign y15006 = 1'b0 ;
  assign y15007 = ~n27233 ;
  assign y15008 = ~n27234 ;
  assign y15009 = ~1'b0 ;
  assign y15010 = ~1'b0 ;
  assign y15011 = n27240 ;
  assign y15012 = ~n27246 ;
  assign y15013 = ~1'b0 ;
  assign y15014 = n27249 ;
  assign y15015 = ~1'b0 ;
  assign y15016 = ~1'b0 ;
  assign y15017 = ~n27250 ;
  assign y15018 = ~1'b0 ;
  assign y15019 = ~n799 ;
  assign y15020 = 1'b0 ;
  assign y15021 = ~1'b0 ;
  assign y15022 = ~n27254 ;
  assign y15023 = ~n27257 ;
  assign y15024 = ~n27258 ;
  assign y15025 = ~1'b0 ;
  assign y15026 = n27259 ;
  assign y15027 = ~n27261 ;
  assign y15028 = n27269 ;
  assign y15029 = ~n27270 ;
  assign y15030 = ~1'b0 ;
  assign y15031 = ~1'b0 ;
  assign y15032 = ~n27273 ;
  assign y15033 = n27275 ;
  assign y15034 = n27279 ;
  assign y15035 = ~n27281 ;
  assign y15036 = n27285 ;
  assign y15037 = n27290 ;
  assign y15038 = n27292 ;
  assign y15039 = ~n24927 ;
  assign y15040 = n27293 ;
  assign y15041 = ~n27299 ;
  assign y15042 = n27300 ;
  assign y15043 = ~1'b0 ;
  assign y15044 = n5507 ;
  assign y15045 = ~1'b0 ;
  assign y15046 = n27306 ;
  assign y15047 = ~1'b0 ;
  assign y15048 = ~1'b0 ;
  assign y15049 = ~n27309 ;
  assign y15050 = n27311 ;
  assign y15051 = ~1'b0 ;
  assign y15052 = n27312 ;
  assign y15053 = ~n27314 ;
  assign y15054 = ~1'b0 ;
  assign y15055 = ~n27315 ;
  assign y15056 = ~n27319 ;
  assign y15057 = ~n27320 ;
  assign y15058 = ~1'b0 ;
  assign y15059 = n27323 ;
  assign y15060 = n27324 ;
  assign y15061 = ~n27329 ;
  assign y15062 = n27331 ;
  assign y15063 = 1'b0 ;
  assign y15064 = ~n27332 ;
  assign y15065 = n11979 ;
  assign y15066 = 1'b0 ;
  assign y15067 = n27333 ;
  assign y15068 = ~1'b0 ;
  assign y15069 = ~n14424 ;
  assign y15070 = ~n27337 ;
  assign y15071 = n27338 ;
  assign y15072 = ~n27340 ;
  assign y15073 = n27341 ;
  assign y15074 = ~n27343 ;
  assign y15075 = ~n27346 ;
  assign y15076 = n27349 ;
  assign y15077 = ~n27350 ;
  assign y15078 = ~n27352 ;
  assign y15079 = n9731 ;
  assign y15080 = ~1'b0 ;
  assign y15081 = ~n27360 ;
  assign y15082 = n27362 ;
  assign y15083 = ~n27369 ;
  assign y15084 = ~n27380 ;
  assign y15085 = ~1'b0 ;
  assign y15086 = n27382 ;
  assign y15087 = ~1'b0 ;
  assign y15088 = ~1'b0 ;
  assign y15089 = 1'b0 ;
  assign y15090 = ~n27383 ;
  assign y15091 = n21061 ;
  assign y15092 = n27385 ;
  assign y15093 = n27386 ;
  assign y15094 = n27387 ;
  assign y15095 = ~n27389 ;
  assign y15096 = ~1'b0 ;
  assign y15097 = ~1'b0 ;
  assign y15098 = ~1'b0 ;
  assign y15099 = ~1'b0 ;
  assign y15100 = ~1'b0 ;
  assign y15101 = ~n27392 ;
  assign y15102 = n27394 ;
  assign y15103 = ~n27396 ;
  assign y15104 = ~n27397 ;
  assign y15105 = n27402 ;
  assign y15106 = ~1'b0 ;
  assign y15107 = ~n27403 ;
  assign y15108 = n27406 ;
  assign y15109 = ~n27410 ;
  assign y15110 = n27414 ;
  assign y15111 = n27416 ;
  assign y15112 = ~1'b0 ;
  assign y15113 = ~n27421 ;
  assign y15114 = ~1'b0 ;
  assign y15115 = ~1'b0 ;
  assign y15116 = n27423 ;
  assign y15117 = ~1'b0 ;
  assign y15118 = ~1'b0 ;
  assign y15119 = ~n27425 ;
  assign y15120 = ~1'b0 ;
  assign y15121 = ~n27428 ;
  assign y15122 = n27431 ;
  assign y15123 = n27437 ;
  assign y15124 = ~1'b0 ;
  assign y15125 = ~1'b0 ;
  assign y15126 = ~n27443 ;
  assign y15127 = ~1'b0 ;
  assign y15128 = ~n27447 ;
  assign y15129 = n27448 ;
  assign y15130 = ~1'b0 ;
  assign y15131 = n27449 ;
  assign y15132 = n27451 ;
  assign y15133 = n23792 ;
  assign y15134 = ~1'b0 ;
  assign y15135 = ~1'b0 ;
  assign y15136 = ~n27453 ;
  assign y15137 = ~1'b0 ;
  assign y15138 = ~n27454 ;
  assign y15139 = ~n27455 ;
  assign y15140 = n27460 ;
  assign y15141 = n27461 ;
  assign y15142 = ~1'b0 ;
  assign y15143 = ~1'b0 ;
  assign y15144 = ~1'b0 ;
  assign y15145 = ~n27464 ;
  assign y15146 = n27471 ;
  assign y15147 = ~1'b0 ;
  assign y15148 = n20756 ;
  assign y15149 = ~n27472 ;
  assign y15150 = n27476 ;
  assign y15151 = ~1'b0 ;
  assign y15152 = 1'b0 ;
  assign y15153 = n2159 ;
  assign y15154 = ~n27477 ;
  assign y15155 = ~1'b0 ;
  assign y15156 = n27480 ;
  assign y15157 = ~n27482 ;
  assign y15158 = ~n27485 ;
  assign y15159 = n27486 ;
  assign y15160 = ~n27489 ;
  assign y15161 = n27492 ;
  assign y15162 = n27495 ;
  assign y15163 = ~1'b0 ;
  assign y15164 = 1'b0 ;
  assign y15165 = ~1'b0 ;
  assign y15166 = n27497 ;
  assign y15167 = ~1'b0 ;
  assign y15168 = ~1'b0 ;
  assign y15169 = ~n27504 ;
  assign y15170 = ~n27506 ;
  assign y15171 = ~n27507 ;
  assign y15172 = n27508 ;
  assign y15173 = ~n27511 ;
  assign y15174 = ~1'b0 ;
  assign y15175 = n27514 ;
  assign y15176 = n27521 ;
  assign y15177 = ~1'b0 ;
  assign y15178 = n4757 ;
  assign y15179 = n27522 ;
  assign y15180 = ~1'b0 ;
  assign y15181 = ~n10532 ;
  assign y15182 = n27523 ;
  assign y15183 = ~1'b0 ;
  assign y15184 = ~n27525 ;
  assign y15185 = n27527 ;
  assign y15186 = ~1'b0 ;
  assign y15187 = 1'b0 ;
  assign y15188 = ~1'b0 ;
  assign y15189 = ~1'b0 ;
  assign y15190 = n27529 ;
  assign y15191 = ~1'b0 ;
  assign y15192 = ~n27531 ;
  assign y15193 = n27534 ;
  assign y15194 = n27535 ;
  assign y15195 = ~1'b0 ;
  assign y15196 = ~n27536 ;
  assign y15197 = ~n27538 ;
  assign y15198 = ~1'b0 ;
  assign y15199 = n27541 ;
  assign y15200 = ~n27543 ;
  assign y15201 = n27545 ;
  assign y15202 = n27548 ;
  assign y15203 = n27549 ;
  assign y15204 = ~n27550 ;
  assign y15205 = ~n27552 ;
  assign y15206 = ~n27553 ;
  assign y15207 = n27559 ;
  assign y15208 = n27561 ;
  assign y15209 = ~1'b0 ;
  assign y15210 = ~n27563 ;
  assign y15211 = ~n27565 ;
  assign y15212 = ~1'b0 ;
  assign y15213 = ~n27568 ;
  assign y15214 = ~1'b0 ;
  assign y15215 = n13311 ;
  assign y15216 = n27569 ;
  assign y15217 = ~n27573 ;
  assign y15218 = ~1'b0 ;
  assign y15219 = ~n27575 ;
  assign y15220 = n27576 ;
  assign y15221 = ~1'b0 ;
  assign y15222 = ~1'b0 ;
  assign y15223 = n5547 ;
  assign y15224 = ~n27580 ;
  assign y15225 = ~1'b0 ;
  assign y15226 = n1157 ;
  assign y15227 = ~n27584 ;
  assign y15228 = ~1'b0 ;
  assign y15229 = n27589 ;
  assign y15230 = n27592 ;
  assign y15231 = ~1'b0 ;
  assign y15232 = ~1'b0 ;
  assign y15233 = n27593 ;
  assign y15234 = n27595 ;
  assign y15235 = ~1'b0 ;
  assign y15236 = ~1'b0 ;
  assign y15237 = ~n27597 ;
  assign y15238 = n27601 ;
  assign y15239 = n27602 ;
  assign y15240 = 1'b0 ;
  assign y15241 = ~n27604 ;
  assign y15242 = ~n27605 ;
  assign y15243 = ~1'b0 ;
  assign y15244 = n27611 ;
  assign y15245 = n27613 ;
  assign y15246 = n27614 ;
  assign y15247 = n27619 ;
  assign y15248 = ~1'b0 ;
  assign y15249 = n27623 ;
  assign y15250 = ~n27631 ;
  assign y15251 = n27633 ;
  assign y15252 = ~1'b0 ;
  assign y15253 = n27640 ;
  assign y15254 = 1'b0 ;
  assign y15255 = n27643 ;
  assign y15256 = n27644 ;
  assign y15257 = ~n27653 ;
  assign y15258 = ~1'b0 ;
  assign y15259 = n27657 ;
  assign y15260 = n27659 ;
  assign y15261 = ~n27664 ;
  assign y15262 = ~1'b0 ;
  assign y15263 = ~1'b0 ;
  assign y15264 = ~n27666 ;
  assign y15265 = ~n27670 ;
  assign y15266 = ~n25774 ;
  assign y15267 = ~n27672 ;
  assign y15268 = ~1'b0 ;
  assign y15269 = ~1'b0 ;
  assign y15270 = n27678 ;
  assign y15271 = ~1'b0 ;
  assign y15272 = ~n27680 ;
  assign y15273 = ~n27681 ;
  assign y15274 = n27684 ;
  assign y15275 = ~n27685 ;
  assign y15276 = n27688 ;
  assign y15277 = ~n27696 ;
  assign y15278 = 1'b0 ;
  assign y15279 = ~n27702 ;
  assign y15280 = ~1'b0 ;
  assign y15281 = ~n27707 ;
  assign y15282 = ~1'b0 ;
  assign y15283 = ~1'b0 ;
  assign y15284 = ~1'b0 ;
  assign y15285 = ~1'b0 ;
  assign y15286 = n27713 ;
  assign y15287 = ~1'b0 ;
  assign y15288 = ~n27715 ;
  assign y15289 = n27716 ;
  assign y15290 = ~1'b0 ;
  assign y15291 = ~n27717 ;
  assign y15292 = ~1'b0 ;
  assign y15293 = ~1'b0 ;
  assign y15294 = n27718 ;
  assign y15295 = n27720 ;
  assign y15296 = ~1'b0 ;
  assign y15297 = n27721 ;
  assign y15298 = ~n27726 ;
  assign y15299 = n27729 ;
  assign y15300 = n15424 ;
  assign y15301 = ~1'b0 ;
  assign y15302 = n27730 ;
  assign y15303 = ~n27731 ;
  assign y15304 = ~1'b0 ;
  assign y15305 = ~1'b0 ;
  assign y15306 = ~1'b0 ;
  assign y15307 = n27733 ;
  assign y15308 = ~1'b0 ;
  assign y15309 = ~n27735 ;
  assign y15310 = ~1'b0 ;
  assign y15311 = ~1'b0 ;
  assign y15312 = ~n27737 ;
  assign y15313 = n27744 ;
  assign y15314 = ~1'b0 ;
  assign y15315 = ~n27746 ;
  assign y15316 = ~n27750 ;
  assign y15317 = ~1'b0 ;
  assign y15318 = ~1'b0 ;
  assign y15319 = ~n27751 ;
  assign y15320 = ~1'b0 ;
  assign y15321 = n10544 ;
  assign y15322 = n27752 ;
  assign y15323 = ~n27753 ;
  assign y15324 = ~n27762 ;
  assign y15325 = ~1'b0 ;
  assign y15326 = n27765 ;
  assign y15327 = ~1'b0 ;
  assign y15328 = ~1'b0 ;
  assign y15329 = ~n27766 ;
  assign y15330 = 1'b0 ;
  assign y15331 = ~n27767 ;
  assign y15332 = ~1'b0 ;
  assign y15333 = n27769 ;
  assign y15334 = ~1'b0 ;
  assign y15335 = ~n27771 ;
  assign y15336 = n27773 ;
  assign y15337 = 1'b0 ;
  assign y15338 = 1'b0 ;
  assign y15339 = ~1'b0 ;
  assign y15340 = ~1'b0 ;
  assign y15341 = ~n27776 ;
  assign y15342 = n27777 ;
  assign y15343 = ~n27778 ;
  assign y15344 = ~1'b0 ;
  assign y15345 = n27783 ;
  assign y15346 = ~n27785 ;
  assign y15347 = n27792 ;
  assign y15348 = ~n27793 ;
  assign y15349 = n27796 ;
  assign y15350 = ~1'b0 ;
  assign y15351 = n27798 ;
  assign y15352 = ~1'b0 ;
  assign y15353 = ~n4119 ;
  assign y15354 = ~1'b0 ;
  assign y15355 = ~1'b0 ;
  assign y15356 = ~1'b0 ;
  assign y15357 = n27799 ;
  assign y15358 = 1'b0 ;
  assign y15359 = ~n27800 ;
  assign y15360 = ~n3097 ;
  assign y15361 = n27802 ;
  assign y15362 = ~1'b0 ;
  assign y15363 = ~1'b0 ;
  assign y15364 = ~1'b0 ;
  assign y15365 = ~n27806 ;
  assign y15366 = ~n24580 ;
  assign y15367 = ~n27807 ;
  assign y15368 = ~n27811 ;
  assign y15369 = ~n27812 ;
  assign y15370 = n27813 ;
  assign y15371 = ~n27814 ;
  assign y15372 = ~n27815 ;
  assign y15373 = ~1'b0 ;
  assign y15374 = ~n15897 ;
  assign y15375 = ~n27817 ;
  assign y15376 = n27821 ;
  assign y15377 = ~n27824 ;
  assign y15378 = ~n27825 ;
  assign y15379 = ~n27827 ;
  assign y15380 = ~n12237 ;
  assign y15381 = ~n27829 ;
  assign y15382 = n27830 ;
  assign y15383 = ~n27833 ;
  assign y15384 = 1'b0 ;
  assign y15385 = n27836 ;
  assign y15386 = ~n27841 ;
  assign y15387 = n27843 ;
  assign y15388 = ~1'b0 ;
  assign y15389 = ~1'b0 ;
  assign y15390 = ~1'b0 ;
  assign y15391 = n27846 ;
  assign y15392 = n27847 ;
  assign y15393 = ~n27853 ;
  assign y15394 = 1'b0 ;
  assign y15395 = ~n4653 ;
  assign y15396 = ~n27856 ;
  assign y15397 = ~n16751 ;
  assign y15398 = ~n19524 ;
  assign y15399 = ~n27857 ;
  assign y15400 = n27860 ;
  assign y15401 = ~n27866 ;
  assign y15402 = ~n27868 ;
  assign y15403 = n27874 ;
  assign y15404 = n27876 ;
  assign y15405 = n27878 ;
  assign y15406 = ~1'b0 ;
  assign y15407 = n27881 ;
  assign y15408 = ~1'b0 ;
  assign y15409 = ~n27883 ;
  assign y15410 = n27886 ;
  assign y15411 = n27889 ;
  assign y15412 = ~1'b0 ;
  assign y15413 = ~1'b0 ;
  assign y15414 = n27895 ;
  assign y15415 = ~1'b0 ;
  assign y15416 = ~n27899 ;
  assign y15417 = ~n27900 ;
  assign y15418 = ~1'b0 ;
  assign y15419 = ~n27904 ;
  assign y15420 = n24500 ;
  assign y15421 = ~1'b0 ;
  assign y15422 = n27913 ;
  assign y15423 = ~1'b0 ;
  assign y15424 = ~n27914 ;
  assign y15425 = n1300 ;
  assign y15426 = ~n27916 ;
  assign y15427 = ~1'b0 ;
  assign y15428 = ~1'b0 ;
  assign y15429 = n27917 ;
  assign y15430 = ~n27918 ;
  assign y15431 = n27922 ;
  assign y15432 = ~n27923 ;
  assign y15433 = ~1'b0 ;
  assign y15434 = ~1'b0 ;
  assign y15435 = ~n27925 ;
  assign y15436 = ~n25269 ;
  assign y15437 = ~n27929 ;
  assign y15438 = ~n27934 ;
  assign y15439 = ~n27935 ;
  assign y15440 = ~n27939 ;
  assign y15441 = n27940 ;
  assign y15442 = n27945 ;
  assign y15443 = ~n12807 ;
  assign y15444 = n27948 ;
  assign y15445 = ~1'b0 ;
  assign y15446 = n27949 ;
  assign y15447 = ~1'b0 ;
  assign y15448 = n27951 ;
  assign y15449 = ~n27954 ;
  assign y15450 = ~1'b0 ;
  assign y15451 = 1'b0 ;
  assign y15452 = ~1'b0 ;
  assign y15453 = n27956 ;
  assign y15454 = ~1'b0 ;
  assign y15455 = n27959 ;
  assign y15456 = ~1'b0 ;
  assign y15457 = ~n27960 ;
  assign y15458 = ~n27962 ;
  assign y15459 = ~1'b0 ;
  assign y15460 = n27964 ;
  assign y15461 = n27970 ;
  assign y15462 = ~1'b0 ;
  assign y15463 = ~n27972 ;
  assign y15464 = ~n8399 ;
  assign y15465 = ~n27976 ;
  assign y15466 = ~n27977 ;
  assign y15467 = ~n27982 ;
  assign y15468 = 1'b0 ;
  assign y15469 = n27984 ;
  assign y15470 = n27987 ;
  assign y15471 = n27989 ;
  assign y15472 = n6273 ;
  assign y15473 = ~n27991 ;
  assign y15474 = ~n27992 ;
  assign y15475 = ~1'b0 ;
  assign y15476 = n2316 ;
  assign y15477 = ~n27993 ;
  assign y15478 = ~1'b0 ;
  assign y15479 = n27995 ;
  assign y15480 = n20101 ;
  assign y15481 = ~n26692 ;
  assign y15482 = ~1'b0 ;
  assign y15483 = ~n28001 ;
  assign y15484 = ~n28005 ;
  assign y15485 = n28019 ;
  assign y15486 = ~1'b0 ;
  assign y15487 = ~n28020 ;
  assign y15488 = ~1'b0 ;
  assign y15489 = ~1'b0 ;
  assign y15490 = ~1'b0 ;
  assign y15491 = ~1'b0 ;
  assign y15492 = ~1'b0 ;
  assign y15493 = ~n24537 ;
  assign y15494 = ~n28023 ;
  assign y15495 = ~1'b0 ;
  assign y15496 = ~1'b0 ;
  assign y15497 = ~1'b0 ;
  assign y15498 = 1'b0 ;
  assign y15499 = ~n28025 ;
  assign y15500 = ~1'b0 ;
  assign y15501 = ~1'b0 ;
  assign y15502 = ~1'b0 ;
  assign y15503 = n28026 ;
  assign y15504 = ~1'b0 ;
  assign y15505 = ~1'b0 ;
  assign y15506 = ~1'b0 ;
  assign y15507 = ~1'b0 ;
  assign y15508 = ~1'b0 ;
  assign y15509 = n28027 ;
  assign y15510 = ~1'b0 ;
  assign y15511 = ~1'b0 ;
  assign y15512 = ~n28032 ;
  assign y15513 = ~1'b0 ;
  assign y15514 = ~n28035 ;
  assign y15515 = ~1'b0 ;
  assign y15516 = ~n28037 ;
  assign y15517 = ~1'b0 ;
  assign y15518 = ~n28039 ;
  assign y15519 = n28040 ;
  assign y15520 = n28041 ;
  assign y15521 = ~1'b0 ;
  assign y15522 = ~n28043 ;
  assign y15523 = n28045 ;
  assign y15524 = ~n28048 ;
  assign y15525 = 1'b0 ;
  assign y15526 = ~1'b0 ;
  assign y15527 = ~1'b0 ;
  assign y15528 = ~n5417 ;
  assign y15529 = n28050 ;
  assign y15530 = ~n17198 ;
  assign y15531 = ~1'b0 ;
  assign y15532 = ~1'b0 ;
  assign y15533 = n28055 ;
  assign y15534 = n344 ;
  assign y15535 = n28057 ;
  assign y15536 = ~n28059 ;
  assign y15537 = ~n18895 ;
  assign y15538 = n13801 ;
  assign y15539 = n28061 ;
  assign y15540 = ~1'b0 ;
  assign y15541 = ~n28062 ;
  assign y15542 = n28063 ;
  assign y15543 = n28064 ;
  assign y15544 = n28066 ;
  assign y15545 = ~1'b0 ;
  assign y15546 = ~1'b0 ;
  assign y15547 = ~n28072 ;
  assign y15548 = n28075 ;
  assign y15549 = ~n28077 ;
  assign y15550 = ~n28081 ;
  assign y15551 = n7265 ;
  assign y15552 = ~1'b0 ;
  assign y15553 = n28088 ;
  assign y15554 = n28094 ;
  assign y15555 = ~n28096 ;
  assign y15556 = n28100 ;
  assign y15557 = n28102 ;
  assign y15558 = n13048 ;
  assign y15559 = n28106 ;
  assign y15560 = ~1'b0 ;
  assign y15561 = n2653 ;
  assign y15562 = n28109 ;
  assign y15563 = ~1'b0 ;
  assign y15564 = ~1'b0 ;
  assign y15565 = ~1'b0 ;
  assign y15566 = n28110 ;
  assign y15567 = ~n28112 ;
  assign y15568 = ~1'b0 ;
  assign y15569 = n28113 ;
  assign y15570 = ~n28115 ;
  assign y15571 = ~n28119 ;
  assign y15572 = n28121 ;
  assign y15573 = ~1'b0 ;
  assign y15574 = ~n28124 ;
  assign y15575 = ~1'b0 ;
  assign y15576 = ~1'b0 ;
  assign y15577 = ~1'b0 ;
  assign y15578 = ~n28127 ;
  assign y15579 = n28128 ;
  assign y15580 = ~n21868 ;
  assign y15581 = n28131 ;
  assign y15582 = ~1'b0 ;
  assign y15583 = n1804 ;
  assign y15584 = ~n28132 ;
  assign y15585 = ~n7972 ;
  assign y15586 = ~n28134 ;
  assign y15587 = n28135 ;
  assign y15588 = n28141 ;
  assign y15589 = ~n28144 ;
  assign y15590 = n28145 ;
  assign y15591 = ~1'b0 ;
  assign y15592 = n28150 ;
  assign y15593 = ~n28151 ;
  assign y15594 = ~1'b0 ;
  assign y15595 = ~1'b0 ;
  assign y15596 = 1'b0 ;
  assign y15597 = ~n1080 ;
  assign y15598 = ~n28153 ;
  assign y15599 = n28159 ;
  assign y15600 = n28160 ;
  assign y15601 = n28164 ;
  assign y15602 = ~n28166 ;
  assign y15603 = ~1'b0 ;
  assign y15604 = ~1'b0 ;
  assign y15605 = ~1'b0 ;
  assign y15606 = ~1'b0 ;
  assign y15607 = ~1'b0 ;
  assign y15608 = ~n28173 ;
  assign y15609 = ~n28175 ;
  assign y15610 = n28177 ;
  assign y15611 = n6827 ;
  assign y15612 = ~n28179 ;
  assign y15613 = n28182 ;
  assign y15614 = 1'b0 ;
  assign y15615 = ~n28185 ;
  assign y15616 = n28187 ;
  assign y15617 = n28188 ;
  assign y15618 = ~1'b0 ;
  assign y15619 = ~n28190 ;
  assign y15620 = ~1'b0 ;
  assign y15621 = n1545 ;
  assign y15622 = 1'b0 ;
  assign y15623 = ~n28192 ;
  assign y15624 = ~n28193 ;
  assign y15625 = ~n6984 ;
  assign y15626 = n28198 ;
  assign y15627 = ~n28200 ;
  assign y15628 = n28201 ;
  assign y15629 = ~1'b0 ;
  assign y15630 = ~n28203 ;
  assign y15631 = n5178 ;
  assign y15632 = ~1'b0 ;
  assign y15633 = n28204 ;
  assign y15634 = ~n28205 ;
  assign y15635 = ~1'b0 ;
  assign y15636 = ~1'b0 ;
  assign y15637 = ~1'b0 ;
  assign y15638 = n28211 ;
  assign y15639 = ~n28217 ;
  assign y15640 = n28219 ;
  assign y15641 = n28220 ;
  assign y15642 = ~1'b0 ;
  assign y15643 = ~1'b0 ;
  assign y15644 = n511 ;
  assign y15645 = 1'b0 ;
  assign y15646 = ~1'b0 ;
  assign y15647 = ~n28222 ;
  assign y15648 = ~n28224 ;
  assign y15649 = ~1'b0 ;
  assign y15650 = n28227 ;
  assign y15651 = ~n28233 ;
  assign y15652 = ~n28236 ;
  assign y15653 = ~1'b0 ;
  assign y15654 = ~n28239 ;
  assign y15655 = n28246 ;
  assign y15656 = n20831 ;
  assign y15657 = n28253 ;
  assign y15658 = ~1'b0 ;
  assign y15659 = n28258 ;
  assign y15660 = n28262 ;
  assign y15661 = ~n28265 ;
  assign y15662 = ~n28267 ;
  assign y15663 = n28268 ;
  assign y15664 = n28270 ;
  assign y15665 = ~n6946 ;
  assign y15666 = n28276 ;
  assign y15667 = n8814 ;
  assign y15668 = ~n28277 ;
  assign y15669 = n28280 ;
  assign y15670 = n28281 ;
  assign y15671 = n28283 ;
  assign y15672 = ~n28285 ;
  assign y15673 = ~n28287 ;
  assign y15674 = ~n28288 ;
  assign y15675 = ~n28292 ;
  assign y15676 = n28298 ;
  assign y15677 = n28299 ;
  assign y15678 = ~n28305 ;
  assign y15679 = ~n28308 ;
  assign y15680 = ~1'b0 ;
  assign y15681 = ~n28314 ;
  assign y15682 = n28317 ;
  assign y15683 = ~1'b0 ;
  assign y15684 = ~n28320 ;
  assign y15685 = ~1'b0 ;
  assign y15686 = ~n28321 ;
  assign y15687 = ~1'b0 ;
  assign y15688 = ~1'b0 ;
  assign y15689 = ~n28324 ;
  assign y15690 = ~1'b0 ;
  assign y15691 = ~1'b0 ;
  assign y15692 = n8662 ;
  assign y15693 = ~n28325 ;
  assign y15694 = ~n11758 ;
  assign y15695 = n28327 ;
  assign y15696 = n28329 ;
  assign y15697 = ~n28331 ;
  assign y15698 = ~1'b0 ;
  assign y15699 = ~1'b0 ;
  assign y15700 = n28332 ;
  assign y15701 = 1'b0 ;
  assign y15702 = ~n28335 ;
  assign y15703 = ~1'b0 ;
  assign y15704 = ~n28341 ;
  assign y15705 = ~1'b0 ;
  assign y15706 = n28347 ;
  assign y15707 = n12878 ;
  assign y15708 = ~n28351 ;
  assign y15709 = n28355 ;
  assign y15710 = n26729 ;
  assign y15711 = n28363 ;
  assign y15712 = ~n28366 ;
  assign y15713 = ~1'b0 ;
  assign y15714 = ~n28367 ;
  assign y15715 = ~1'b0 ;
  assign y15716 = ~1'b0 ;
  assign y15717 = ~1'b0 ;
  assign y15718 = ~n28369 ;
  assign y15719 = n28370 ;
  assign y15720 = 1'b0 ;
  assign y15721 = ~1'b0 ;
  assign y15722 = ~n28373 ;
  assign y15723 = ~n24886 ;
  assign y15724 = ~1'b0 ;
  assign y15725 = n28377 ;
  assign y15726 = ~n3535 ;
  assign y15727 = n4040 ;
  assign y15728 = n28379 ;
  assign y15729 = ~n28386 ;
  assign y15730 = ~n28387 ;
  assign y15731 = ~1'b0 ;
  assign y15732 = n28390 ;
  assign y15733 = n28392 ;
  assign y15734 = n28393 ;
  assign y15735 = ~n28397 ;
  assign y15736 = n28405 ;
  assign y15737 = ~n28408 ;
  assign y15738 = ~1'b0 ;
  assign y15739 = n28410 ;
  assign y15740 = n28412 ;
  assign y15741 = ~1'b0 ;
  assign y15742 = 1'b0 ;
  assign y15743 = n28414 ;
  assign y15744 = ~n28418 ;
  assign y15745 = ~1'b0 ;
  assign y15746 = ~1'b0 ;
  assign y15747 = ~1'b0 ;
  assign y15748 = n28419 ;
  assign y15749 = n28423 ;
  assign y15750 = n28424 ;
  assign y15751 = ~n28425 ;
  assign y15752 = ~1'b0 ;
  assign y15753 = n28427 ;
  assign y15754 = n28429 ;
  assign y15755 = n28431 ;
  assign y15756 = ~n28433 ;
  assign y15757 = n28434 ;
  assign y15758 = ~n28440 ;
  assign y15759 = n28442 ;
  assign y15760 = n28443 ;
  assign y15761 = ~1'b0 ;
  assign y15762 = n28444 ;
  assign y15763 = n28445 ;
  assign y15764 = n28447 ;
  assign y15765 = ~n28451 ;
  assign y15766 = ~n28454 ;
  assign y15767 = n28455 ;
  assign y15768 = ~n28460 ;
  assign y15769 = n28461 ;
  assign y15770 = ~1'b0 ;
  assign y15771 = n28470 ;
  assign y15772 = ~1'b0 ;
  assign y15773 = n28474 ;
  assign y15774 = n28475 ;
  assign y15775 = n28478 ;
  assign y15776 = ~1'b0 ;
  assign y15777 = ~n28480 ;
  assign y15778 = ~1'b0 ;
  assign y15779 = n28482 ;
  assign y15780 = ~1'b0 ;
  assign y15781 = n28484 ;
  assign y15782 = ~n28485 ;
  assign y15783 = n28487 ;
  assign y15784 = ~n28488 ;
  assign y15785 = ~1'b0 ;
  assign y15786 = ~n28491 ;
  assign y15787 = ~n28492 ;
  assign y15788 = n28496 ;
  assign y15789 = ~1'b0 ;
  assign y15790 = ~n16468 ;
  assign y15791 = ~n28498 ;
  assign y15792 = ~n28502 ;
  assign y15793 = n28503 ;
  assign y15794 = ~n28505 ;
  assign y15795 = ~n28506 ;
  assign y15796 = ~n28508 ;
  assign y15797 = ~n28515 ;
  assign y15798 = ~n8406 ;
  assign y15799 = n28516 ;
  assign y15800 = ~n28521 ;
  assign y15801 = ~n28524 ;
  assign y15802 = n28525 ;
  assign y15803 = ~n28526 ;
  assign y15804 = ~1'b0 ;
  assign y15805 = n28527 ;
  assign y15806 = ~1'b0 ;
  assign y15807 = ~n28528 ;
  assign y15808 = n28529 ;
  assign y15809 = n28534 ;
  assign y15810 = ~n28537 ;
  assign y15811 = n28542 ;
  assign y15812 = ~1'b0 ;
  assign y15813 = n28546 ;
  assign y15814 = n28550 ;
  assign y15815 = n28552 ;
  assign y15816 = ~1'b0 ;
  assign y15817 = ~1'b0 ;
  assign y15818 = ~1'b0 ;
  assign y15819 = ~n1477 ;
  assign y15820 = ~n28553 ;
  assign y15821 = ~n28557 ;
  assign y15822 = n28558 ;
  assign y15823 = 1'b0 ;
  assign y15824 = ~1'b0 ;
  assign y15825 = ~n28559 ;
  assign y15826 = ~1'b0 ;
  assign y15827 = n28560 ;
  assign y15828 = ~1'b0 ;
  assign y15829 = ~n28562 ;
  assign y15830 = n28563 ;
  assign y15831 = ~1'b0 ;
  assign y15832 = ~1'b0 ;
  assign y15833 = n28564 ;
  assign y15834 = ~1'b0 ;
  assign y15835 = 1'b0 ;
  assign y15836 = ~1'b0 ;
  assign y15837 = ~n28565 ;
  assign y15838 = n28567 ;
  assign y15839 = ~1'b0 ;
  assign y15840 = n28575 ;
  assign y15841 = ~n28577 ;
  assign y15842 = n28581 ;
  assign y15843 = ~n28582 ;
  assign y15844 = ~n28584 ;
  assign y15845 = ~1'b0 ;
  assign y15846 = 1'b0 ;
  assign y15847 = n25231 ;
  assign y15848 = n28585 ;
  assign y15849 = ~1'b0 ;
  assign y15850 = ~1'b0 ;
  assign y15851 = ~n28587 ;
  assign y15852 = n28591 ;
  assign y15853 = n28593 ;
  assign y15854 = ~n28596 ;
  assign y15855 = n28599 ;
  assign y15856 = n28602 ;
  assign y15857 = ~n28604 ;
  assign y15858 = ~n8273 ;
  assign y15859 = n28609 ;
  assign y15860 = n28611 ;
  assign y15861 = ~n5142 ;
  assign y15862 = ~1'b0 ;
  assign y15863 = n28612 ;
  assign y15864 = ~n21982 ;
  assign y15865 = ~1'b0 ;
  assign y15866 = ~1'b0 ;
  assign y15867 = ~n28613 ;
  assign y15868 = ~1'b0 ;
  assign y15869 = ~n28614 ;
  assign y15870 = n28619 ;
  assign y15871 = ~1'b0 ;
  assign y15872 = n28620 ;
  assign y15873 = n28622 ;
  assign y15874 = ~1'b0 ;
  assign y15875 = ~1'b0 ;
  assign y15876 = ~n28624 ;
  assign y15877 = 1'b0 ;
  assign y15878 = ~n3592 ;
  assign y15879 = ~1'b0 ;
  assign y15880 = ~n28626 ;
  assign y15881 = ~n28628 ;
  assign y15882 = ~n28632 ;
  assign y15883 = ~n28633 ;
  assign y15884 = n28634 ;
  assign y15885 = ~n28636 ;
  assign y15886 = ~n28639 ;
  assign y15887 = ~n28640 ;
  assign y15888 = ~n28644 ;
  assign y15889 = 1'b0 ;
  assign y15890 = ~n28645 ;
  assign y15891 = n28666 ;
  assign y15892 = n28667 ;
  assign y15893 = ~1'b0 ;
  assign y15894 = n28674 ;
  assign y15895 = ~1'b0 ;
  assign y15896 = ~n28676 ;
  assign y15897 = ~n28680 ;
  assign y15898 = n28685 ;
  assign y15899 = ~n28690 ;
  assign y15900 = 1'b0 ;
  assign y15901 = ~1'b0 ;
  assign y15902 = n4570 ;
  assign y15903 = ~1'b0 ;
  assign y15904 = ~n28697 ;
  assign y15905 = ~n28699 ;
  assign y15906 = ~n28700 ;
  assign y15907 = n28703 ;
  assign y15908 = ~n28704 ;
  assign y15909 = ~1'b0 ;
  assign y15910 = ~1'b0 ;
  assign y15911 = n28706 ;
  assign y15912 = ~n28708 ;
  assign y15913 = ~1'b0 ;
  assign y15914 = ~n28713 ;
  assign y15915 = ~1'b0 ;
  assign y15916 = n28716 ;
  assign y15917 = ~1'b0 ;
  assign y15918 = ~1'b0 ;
  assign y15919 = ~n28718 ;
  assign y15920 = ~n28719 ;
  assign y15921 = ~n28723 ;
  assign y15922 = ~n28725 ;
  assign y15923 = ~n28728 ;
  assign y15924 = ~n28729 ;
  assign y15925 = n28732 ;
  assign y15926 = n28734 ;
  assign y15927 = n28736 ;
  assign y15928 = ~n28737 ;
  assign y15929 = ~n28741 ;
  assign y15930 = ~1'b0 ;
  assign y15931 = n28742 ;
  assign y15932 = ~n28743 ;
  assign y15933 = n28745 ;
  assign y15934 = ~1'b0 ;
  assign y15935 = ~1'b0 ;
  assign y15936 = ~n28747 ;
  assign y15937 = ~n28751 ;
  assign y15938 = n28755 ;
  assign y15939 = ~n28758 ;
  assign y15940 = ~n28761 ;
  assign y15941 = n28763 ;
  assign y15942 = ~n28776 ;
  assign y15943 = n28777 ;
  assign y15944 = ~1'b0 ;
  assign y15945 = ~n28782 ;
  assign y15946 = ~n16325 ;
  assign y15947 = n5070 ;
  assign y15948 = ~1'b0 ;
  assign y15949 = n28787 ;
  assign y15950 = ~n28789 ;
  assign y15951 = ~n28793 ;
  assign y15952 = ~n28794 ;
  assign y15953 = n28798 ;
  assign y15954 = n28804 ;
  assign y15955 = ~1'b0 ;
  assign y15956 = n28805 ;
  assign y15957 = ~1'b0 ;
  assign y15958 = ~n28806 ;
  assign y15959 = ~n22798 ;
  assign y15960 = n28808 ;
  assign y15961 = n28810 ;
  assign y15962 = n28818 ;
  assign y15963 = n28820 ;
  assign y15964 = ~1'b0 ;
  assign y15965 = n28826 ;
  assign y15966 = n28827 ;
  assign y15967 = ~n28828 ;
  assign y15968 = n28831 ;
  assign y15969 = ~1'b0 ;
  assign y15970 = ~n28833 ;
  assign y15971 = ~1'b0 ;
  assign y15972 = n28834 ;
  assign y15973 = n28836 ;
  assign y15974 = n28840 ;
  assign y15975 = n28845 ;
  assign y15976 = ~1'b0 ;
  assign y15977 = ~n28847 ;
  assign y15978 = ~1'b0 ;
  assign y15979 = ~n28849 ;
  assign y15980 = ~n28853 ;
  assign y15981 = ~n10626 ;
  assign y15982 = n28856 ;
  assign y15983 = n28858 ;
  assign y15984 = 1'b0 ;
  assign y15985 = n28862 ;
  assign y15986 = n28875 ;
  assign y15987 = ~1'b0 ;
  assign y15988 = n28879 ;
  assign y15989 = ~n28880 ;
  assign y15990 = ~n28887 ;
  assign y15991 = n28888 ;
  assign y15992 = ~n28890 ;
  assign y15993 = ~n28892 ;
  assign y15994 = n28894 ;
  assign y15995 = n28896 ;
  assign y15996 = ~1'b0 ;
  assign y15997 = n28897 ;
  assign y15998 = n28899 ;
  assign y15999 = n28901 ;
  assign y16000 = n28903 ;
  assign y16001 = ~n28904 ;
  assign y16002 = ~1'b0 ;
  assign y16003 = n28906 ;
  assign y16004 = ~1'b0 ;
  assign y16005 = ~1'b0 ;
  assign y16006 = ~1'b0 ;
  assign y16007 = ~n28910 ;
  assign y16008 = n28911 ;
  assign y16009 = ~n28918 ;
  assign y16010 = n28921 ;
  assign y16011 = ~n28924 ;
  assign y16012 = n28925 ;
  assign y16013 = ~1'b0 ;
  assign y16014 = ~n26496 ;
  assign y16015 = ~n28926 ;
  assign y16016 = n28927 ;
  assign y16017 = ~n28928 ;
  assign y16018 = n28931 ;
  assign y16019 = n28933 ;
  assign y16020 = n28934 ;
  assign y16021 = ~1'b0 ;
  assign y16022 = n28935 ;
  assign y16023 = ~1'b0 ;
  assign y16024 = ~1'b0 ;
  assign y16025 = ~1'b0 ;
  assign y16026 = ~n28936 ;
  assign y16027 = n28939 ;
  assign y16028 = ~n28940 ;
  assign y16029 = n11542 ;
  assign y16030 = n28943 ;
  assign y16031 = ~1'b0 ;
  assign y16032 = ~1'b0 ;
  assign y16033 = ~1'b0 ;
  assign y16034 = ~n28945 ;
  assign y16035 = n28946 ;
  assign y16036 = n28947 ;
  assign y16037 = ~1'b0 ;
  assign y16038 = ~n28948 ;
  assign y16039 = ~1'b0 ;
  assign y16040 = ~n28952 ;
  assign y16041 = ~n28957 ;
  assign y16042 = n28959 ;
  assign y16043 = ~n28964 ;
  assign y16044 = ~n28965 ;
  assign y16045 = ~n1830 ;
  assign y16046 = ~1'b0 ;
  assign y16047 = n28966 ;
  assign y16048 = ~n28967 ;
  assign y16049 = n28975 ;
  assign y16050 = 1'b0 ;
  assign y16051 = n28978 ;
  assign y16052 = ~n28980 ;
  assign y16053 = ~n28983 ;
  assign y16054 = n28984 ;
  assign y16055 = ~1'b0 ;
  assign y16056 = ~n28985 ;
  assign y16057 = ~1'b0 ;
  assign y16058 = ~n28987 ;
  assign y16059 = ~n14158 ;
  assign y16060 = n812 ;
  assign y16061 = ~n28990 ;
  assign y16062 = ~1'b0 ;
  assign y16063 = ~n6296 ;
  assign y16064 = n28991 ;
  assign y16065 = ~n28992 ;
  assign y16066 = ~n11305 ;
  assign y16067 = ~n28998 ;
  assign y16068 = n29002 ;
  assign y16069 = n29006 ;
  assign y16070 = n29008 ;
  assign y16071 = n29012 ;
  assign y16072 = ~1'b0 ;
  assign y16073 = ~1'b0 ;
  assign y16074 = ~n29015 ;
  assign y16075 = n29017 ;
  assign y16076 = n29019 ;
  assign y16077 = ~n29020 ;
  assign y16078 = n29023 ;
  assign y16079 = ~1'b0 ;
  assign y16080 = ~n29027 ;
  assign y16081 = ~n29029 ;
  assign y16082 = ~1'b0 ;
  assign y16083 = ~n13167 ;
  assign y16084 = ~1'b0 ;
  assign y16085 = ~1'b0 ;
  assign y16086 = ~n29030 ;
  assign y16087 = ~n29031 ;
  assign y16088 = n29036 ;
  assign y16089 = ~n29040 ;
  assign y16090 = ~n29051 ;
  assign y16091 = ~n11694 ;
  assign y16092 = ~n15963 ;
  assign y16093 = ~1'b0 ;
  assign y16094 = ~1'b0 ;
  assign y16095 = n29054 ;
  assign y16096 = 1'b0 ;
  assign y16097 = ~1'b0 ;
  assign y16098 = n29056 ;
  assign y16099 = ~n29058 ;
  assign y16100 = ~n29062 ;
  assign y16101 = n29063 ;
  assign y16102 = ~n29064 ;
  assign y16103 = n2871 ;
  assign y16104 = 1'b0 ;
  assign y16105 = ~n29065 ;
  assign y16106 = ~n29067 ;
  assign y16107 = ~1'b0 ;
  assign y16108 = n29069 ;
  assign y16109 = n29070 ;
  assign y16110 = n14750 ;
  assign y16111 = ~n29072 ;
  assign y16112 = ~1'b0 ;
  assign y16113 = ~1'b0 ;
  assign y16114 = ~n29075 ;
  assign y16115 = ~n29079 ;
  assign y16116 = ~1'b0 ;
  assign y16117 = ~n29087 ;
  assign y16118 = 1'b0 ;
  assign y16119 = ~1'b0 ;
  assign y16120 = ~1'b0 ;
  assign y16121 = ~1'b0 ;
  assign y16122 = ~n29088 ;
  assign y16123 = ~1'b0 ;
  assign y16124 = n29089 ;
  assign y16125 = ~1'b0 ;
  assign y16126 = ~n29093 ;
  assign y16127 = n29096 ;
  assign y16128 = n29097 ;
  assign y16129 = ~1'b0 ;
  assign y16130 = n29098 ;
  assign y16131 = n29100 ;
  assign y16132 = ~n29101 ;
  assign y16133 = ~n29109 ;
  assign y16134 = n29125 ;
  assign y16135 = n29127 ;
  assign y16136 = ~n7528 ;
  assign y16137 = ~1'b0 ;
  assign y16138 = ~n29128 ;
  assign y16139 = ~1'b0 ;
  assign y16140 = ~n29129 ;
  assign y16141 = ~1'b0 ;
  assign y16142 = n29130 ;
  assign y16143 = ~n29131 ;
  assign y16144 = n29135 ;
  assign y16145 = ~1'b0 ;
  assign y16146 = ~n29146 ;
  assign y16147 = ~n29147 ;
  assign y16148 = ~n29148 ;
  assign y16149 = ~n29149 ;
  assign y16150 = n29150 ;
  assign y16151 = ~n29151 ;
  assign y16152 = ~n29152 ;
  assign y16153 = ~n29153 ;
  assign y16154 = ~1'b0 ;
  assign y16155 = ~n29154 ;
  assign y16156 = ~1'b0 ;
  assign y16157 = n29161 ;
  assign y16158 = ~n29164 ;
  assign y16159 = n29165 ;
  assign y16160 = n29170 ;
  assign y16161 = n29173 ;
  assign y16162 = ~n29177 ;
  assign y16163 = ~1'b0 ;
  assign y16164 = ~1'b0 ;
  assign y16165 = ~n29197 ;
  assign y16166 = ~1'b0 ;
  assign y16167 = ~n29201 ;
  assign y16168 = n29203 ;
  assign y16169 = n29205 ;
  assign y16170 = ~n29207 ;
  assign y16171 = n856 ;
  assign y16172 = ~n124 ;
  assign y16173 = n29209 ;
  assign y16174 = ~1'b0 ;
  assign y16175 = n29210 ;
  assign y16176 = n11870 ;
  assign y16177 = ~n29216 ;
  assign y16178 = n29220 ;
  assign y16179 = ~n29222 ;
  assign y16180 = ~1'b0 ;
  assign y16181 = ~n29225 ;
  assign y16182 = ~n29227 ;
  assign y16183 = ~1'b0 ;
  assign y16184 = n29228 ;
  assign y16185 = ~1'b0 ;
  assign y16186 = n29230 ;
  assign y16187 = ~1'b0 ;
  assign y16188 = n29231 ;
  assign y16189 = ~n24620 ;
  assign y16190 = ~1'b0 ;
  assign y16191 = ~1'b0 ;
  assign y16192 = ~n1517 ;
  assign y16193 = ~n29233 ;
  assign y16194 = 1'b0 ;
  assign y16195 = n29237 ;
  assign y16196 = ~n29238 ;
  assign y16197 = ~n29239 ;
  assign y16198 = ~n29242 ;
  assign y16199 = n29250 ;
  assign y16200 = ~1'b0 ;
  assign y16201 = ~1'b0 ;
  assign y16202 = ~n29251 ;
  assign y16203 = n29258 ;
  assign y16204 = n29273 ;
  assign y16205 = ~1'b0 ;
  assign y16206 = n29208 ;
  assign y16207 = n29277 ;
  assign y16208 = n29284 ;
  assign y16209 = n29288 ;
  assign y16210 = 1'b0 ;
  assign y16211 = n29292 ;
  assign y16212 = ~n9769 ;
  assign y16213 = n29295 ;
  assign y16214 = ~1'b0 ;
  assign y16215 = n29297 ;
  assign y16216 = n29298 ;
  assign y16217 = ~n29299 ;
  assign y16218 = ~1'b0 ;
  assign y16219 = ~n29300 ;
  assign y16220 = ~n13114 ;
  assign y16221 = 1'b0 ;
  assign y16222 = ~n29302 ;
  assign y16223 = ~1'b0 ;
  assign y16224 = n29308 ;
  assign y16225 = ~n29311 ;
  assign y16226 = ~n29312 ;
  assign y16227 = ~1'b0 ;
  assign y16228 = ~n29316 ;
  assign y16229 = ~1'b0 ;
  assign y16230 = n29321 ;
  assign y16231 = ~1'b0 ;
  assign y16232 = ~1'b0 ;
  assign y16233 = n29322 ;
  assign y16234 = ~n29328 ;
  assign y16235 = ~1'b0 ;
  assign y16236 = ~n29330 ;
  assign y16237 = n29333 ;
  assign y16238 = ~n29335 ;
  assign y16239 = ~1'b0 ;
  assign y16240 = ~n29339 ;
  assign y16241 = n29341 ;
  assign y16242 = ~1'b0 ;
  assign y16243 = n29343 ;
  assign y16244 = ~1'b0 ;
  assign y16245 = ~n29344 ;
  assign y16246 = ~n29345 ;
  assign y16247 = n29348 ;
  assign y16248 = ~1'b0 ;
  assign y16249 = n29350 ;
  assign y16250 = ~1'b0 ;
  assign y16251 = ~n2468 ;
  assign y16252 = ~n29353 ;
  assign y16253 = ~n29357 ;
  assign y16254 = ~n29362 ;
  assign y16255 = ~n29366 ;
  assign y16256 = ~1'b0 ;
  assign y16257 = ~n29367 ;
  assign y16258 = n29368 ;
  assign y16259 = ~1'b0 ;
  assign y16260 = ~n29370 ;
  assign y16261 = n29373 ;
  assign y16262 = ~n29374 ;
  assign y16263 = 1'b0 ;
  assign y16264 = n29376 ;
  assign y16265 = n29377 ;
  assign y16266 = ~1'b0 ;
  assign y16267 = ~1'b0 ;
  assign y16268 = ~n19159 ;
  assign y16269 = 1'b0 ;
  assign y16270 = ~1'b0 ;
  assign y16271 = n292 ;
  assign y16272 = ~n16716 ;
  assign y16273 = n29378 ;
  assign y16274 = ~n29383 ;
  assign y16275 = ~1'b0 ;
  assign y16276 = ~1'b0 ;
  assign y16277 = ~n29387 ;
  assign y16278 = n29388 ;
  assign y16279 = ~1'b0 ;
  assign y16280 = n29389 ;
  assign y16281 = ~1'b0 ;
  assign y16282 = ~n19941 ;
  assign y16283 = n29390 ;
  assign y16284 = ~n29398 ;
  assign y16285 = ~n29399 ;
  assign y16286 = n29400 ;
  assign y16287 = ~n29404 ;
  assign y16288 = ~n29405 ;
  assign y16289 = ~n29410 ;
  assign y16290 = n29412 ;
  assign y16291 = ~n17201 ;
  assign y16292 = ~n29413 ;
  assign y16293 = ~n29415 ;
  assign y16294 = ~1'b0 ;
  assign y16295 = n29420 ;
  assign y16296 = n29422 ;
  assign y16297 = ~n29424 ;
  assign y16298 = ~n29425 ;
  assign y16299 = n25152 ;
  assign y16300 = ~n25138 ;
  assign y16301 = n29426 ;
  assign y16302 = ~n29428 ;
  assign y16303 = ~n6283 ;
  assign y16304 = n29429 ;
  assign y16305 = ~n29430 ;
  assign y16306 = ~n29432 ;
  assign y16307 = ~n29434 ;
  assign y16308 = n29436 ;
  assign y16309 = ~n29437 ;
  assign y16310 = ~1'b0 ;
  assign y16311 = ~n29439 ;
  assign y16312 = ~1'b0 ;
  assign y16313 = ~n29440 ;
  assign y16314 = ~1'b0 ;
  assign y16315 = ~1'b0 ;
  assign y16316 = ~n29444 ;
  assign y16317 = ~n22740 ;
  assign y16318 = ~n29446 ;
  assign y16319 = 1'b0 ;
  assign y16320 = ~n29449 ;
  assign y16321 = n712 ;
  assign y16322 = n29452 ;
  assign y16323 = n7077 ;
  assign y16324 = ~1'b0 ;
  assign y16325 = ~1'b0 ;
  assign y16326 = ~n29453 ;
  assign y16327 = n29455 ;
  assign y16328 = ~n29459 ;
  assign y16329 = ~n29463 ;
  assign y16330 = ~n29465 ;
  assign y16331 = ~n29473 ;
  assign y16332 = ~1'b0 ;
  assign y16333 = ~n29475 ;
  assign y16334 = ~1'b0 ;
  assign y16335 = ~n29478 ;
  assign y16336 = ~n29480 ;
  assign y16337 = n29485 ;
  assign y16338 = ~1'b0 ;
  assign y16339 = ~1'b0 ;
  assign y16340 = ~1'b0 ;
  assign y16341 = n29489 ;
  assign y16342 = n29496 ;
  assign y16343 = ~1'b0 ;
  assign y16344 = ~1'b0 ;
  assign y16345 = ~1'b0 ;
  assign y16346 = ~n29501 ;
  assign y16347 = ~1'b0 ;
  assign y16348 = ~1'b0 ;
  assign y16349 = ~n29503 ;
  assign y16350 = ~1'b0 ;
  assign y16351 = ~1'b0 ;
  assign y16352 = 1'b0 ;
  assign y16353 = ~n29504 ;
  assign y16354 = n9740 ;
  assign y16355 = ~1'b0 ;
  assign y16356 = ~n29505 ;
  assign y16357 = 1'b0 ;
  assign y16358 = ~1'b0 ;
  assign y16359 = n29506 ;
  assign y16360 = n29509 ;
  assign y16361 = ~n29510 ;
  assign y16362 = ~1'b0 ;
  assign y16363 = n29512 ;
  assign y16364 = ~1'b0 ;
  assign y16365 = n29521 ;
  assign y16366 = ~1'b0 ;
  assign y16367 = ~1'b0 ;
  assign y16368 = n29522 ;
  assign y16369 = ~1'b0 ;
  assign y16370 = ~n29524 ;
  assign y16371 = n29525 ;
  assign y16372 = ~1'b0 ;
  assign y16373 = ~n29526 ;
  assign y16374 = n29527 ;
  assign y16375 = ~1'b0 ;
  assign y16376 = ~n29528 ;
  assign y16377 = n29532 ;
  assign y16378 = ~n29534 ;
  assign y16379 = 1'b0 ;
  assign y16380 = n29536 ;
  assign y16381 = n29540 ;
  assign y16382 = ~n29543 ;
  assign y16383 = n29544 ;
  assign y16384 = ~n29545 ;
  assign y16385 = n29546 ;
  assign y16386 = ~n29551 ;
  assign y16387 = n29552 ;
  assign y16388 = n29554 ;
  assign y16389 = n29555 ;
  assign y16390 = ~1'b0 ;
  assign y16391 = ~1'b0 ;
  assign y16392 = ~n29556 ;
  assign y16393 = n29558 ;
  assign y16394 = ~n23541 ;
  assign y16395 = 1'b0 ;
  assign y16396 = n29559 ;
  assign y16397 = n29560 ;
  assign y16398 = n15509 ;
  assign y16399 = ~n29565 ;
  assign y16400 = n29573 ;
  assign y16401 = n29575 ;
  assign y16402 = n29576 ;
  assign y16403 = ~1'b0 ;
  assign y16404 = ~n29580 ;
  assign y16405 = n29581 ;
  assign y16406 = ~n29583 ;
  assign y16407 = ~n29584 ;
  assign y16408 = ~n1251 ;
  assign y16409 = ~n29585 ;
  assign y16410 = n29589 ;
  assign y16411 = ~n29593 ;
  assign y16412 = ~n29597 ;
  assign y16413 = 1'b0 ;
  assign y16414 = ~n29599 ;
  assign y16415 = ~1'b0 ;
  assign y16416 = ~n29601 ;
  assign y16417 = ~n29606 ;
  assign y16418 = ~n29610 ;
  assign y16419 = ~1'b0 ;
  assign y16420 = n29612 ;
  assign y16421 = n29613 ;
  assign y16422 = ~n29618 ;
  assign y16423 = ~1'b0 ;
  assign y16424 = ~n23926 ;
  assign y16425 = n29621 ;
  assign y16426 = n29622 ;
  assign y16427 = ~1'b0 ;
  assign y16428 = n29623 ;
  assign y16429 = ~n29625 ;
  assign y16430 = n29626 ;
  assign y16431 = n29633 ;
  assign y16432 = n29638 ;
  assign y16433 = ~n29642 ;
  assign y16434 = n29643 ;
  assign y16435 = ~n12541 ;
  assign y16436 = n29645 ;
  assign y16437 = ~1'b0 ;
  assign y16438 = ~n29646 ;
  assign y16439 = ~n29658 ;
  assign y16440 = ~n29659 ;
  assign y16441 = n19032 ;
  assign y16442 = ~n29661 ;
  assign y16443 = ~1'b0 ;
  assign y16444 = n29666 ;
  assign y16445 = n29667 ;
  assign y16446 = ~n29670 ;
  assign y16447 = ~n29671 ;
  assign y16448 = ~n29673 ;
  assign y16449 = ~n29684 ;
  assign y16450 = n29685 ;
  assign y16451 = ~1'b0 ;
  assign y16452 = n29686 ;
  assign y16453 = n29687 ;
  assign y16454 = ~n29691 ;
  assign y16455 = n29692 ;
  assign y16456 = ~n29697 ;
  assign y16457 = n29700 ;
  assign y16458 = ~1'b0 ;
  assign y16459 = ~n29701 ;
  assign y16460 = n29706 ;
  assign y16461 = ~n29708 ;
  assign y16462 = ~n29711 ;
  assign y16463 = ~n29715 ;
  assign y16464 = n29717 ;
  assign y16465 = n23451 ;
  assign y16466 = ~1'b0 ;
  assign y16467 = ~1'b0 ;
  assign y16468 = ~1'b0 ;
  assign y16469 = ~n29723 ;
  assign y16470 = ~1'b0 ;
  assign y16471 = ~n29731 ;
  assign y16472 = ~n29732 ;
  assign y16473 = ~n29734 ;
  assign y16474 = n1528 ;
  assign y16475 = ~n29739 ;
  assign y16476 = ~1'b0 ;
  assign y16477 = ~n3592 ;
  assign y16478 = ~1'b0 ;
  assign y16479 = n29740 ;
  assign y16480 = ~1'b0 ;
  assign y16481 = n29745 ;
  assign y16482 = ~n29746 ;
  assign y16483 = n29748 ;
  assign y16484 = n29750 ;
  assign y16485 = ~n5316 ;
  assign y16486 = ~n29752 ;
  assign y16487 = n29754 ;
  assign y16488 = ~1'b0 ;
  assign y16489 = ~n29755 ;
  assign y16490 = n29757 ;
  assign y16491 = ~n29759 ;
  assign y16492 = n29761 ;
  assign y16493 = ~n29762 ;
  assign y16494 = n18547 ;
  assign y16495 = ~n29765 ;
  assign y16496 = n29766 ;
  assign y16497 = 1'b0 ;
  assign y16498 = ~n29768 ;
  assign y16499 = n29770 ;
  assign y16500 = ~n29771 ;
  assign y16501 = ~1'b0 ;
  assign y16502 = ~1'b0 ;
  assign y16503 = n29772 ;
  assign y16504 = n29775 ;
  assign y16505 = ~n29776 ;
  assign y16506 = ~1'b0 ;
  assign y16507 = ~1'b0 ;
  assign y16508 = n29782 ;
  assign y16509 = n29784 ;
  assign y16510 = ~n29789 ;
  assign y16511 = ~1'b0 ;
  assign y16512 = ~n23387 ;
  assign y16513 = ~n29792 ;
  assign y16514 = ~n29813 ;
  assign y16515 = ~n29814 ;
  assign y16516 = ~1'b0 ;
  assign y16517 = ~n29815 ;
  assign y16518 = ~n29817 ;
  assign y16519 = ~1'b0 ;
  assign y16520 = ~n29821 ;
  assign y16521 = ~n29822 ;
  assign y16522 = ~1'b0 ;
  assign y16523 = n29828 ;
  assign y16524 = ~1'b0 ;
  assign y16525 = ~1'b0 ;
  assign y16526 = n29830 ;
  assign y16527 = ~1'b0 ;
  assign y16528 = n29831 ;
  assign y16529 = n29833 ;
  assign y16530 = ~n29836 ;
  assign y16531 = ~n29837 ;
  assign y16532 = ~n29838 ;
  assign y16533 = ~1'b0 ;
  assign y16534 = ~1'b0 ;
  assign y16535 = ~n29841 ;
  assign y16536 = n29843 ;
  assign y16537 = n29844 ;
  assign y16538 = n29339 ;
  assign y16539 = ~n29845 ;
  assign y16540 = ~n29850 ;
  assign y16541 = ~1'b0 ;
  assign y16542 = ~1'b0 ;
  assign y16543 = ~1'b0 ;
  assign y16544 = ~1'b0 ;
  assign y16545 = n29851 ;
  assign y16546 = ~1'b0 ;
  assign y16547 = ~1'b0 ;
  assign y16548 = ~1'b0 ;
  assign y16549 = ~n29855 ;
  assign y16550 = n29859 ;
  assign y16551 = ~n29861 ;
  assign y16552 = 1'b0 ;
  assign y16553 = ~n29862 ;
  assign y16554 = ~1'b0 ;
  assign y16555 = n10596 ;
  assign y16556 = n29863 ;
  assign y16557 = ~1'b0 ;
  assign y16558 = ~1'b0 ;
  assign y16559 = ~1'b0 ;
  assign y16560 = ~n29865 ;
  assign y16561 = ~n29866 ;
  assign y16562 = n29868 ;
  assign y16563 = ~1'b0 ;
  assign y16564 = n29869 ;
  assign y16565 = 1'b0 ;
  assign y16566 = n29314 ;
  assign y16567 = ~1'b0 ;
  assign y16568 = n26076 ;
  assign y16569 = ~n29871 ;
  assign y16570 = ~1'b0 ;
  assign y16571 = n29872 ;
  assign y16572 = n12582 ;
  assign y16573 = ~1'b0 ;
  assign y16574 = ~n29874 ;
  assign y16575 = ~n29876 ;
  assign y16576 = ~1'b0 ;
  assign y16577 = ~n29877 ;
  assign y16578 = n29880 ;
  assign y16579 = n29881 ;
  assign y16580 = ~1'b0 ;
  assign y16581 = ~n29883 ;
  assign y16582 = ~n29886 ;
  assign y16583 = ~1'b0 ;
  assign y16584 = ~n29887 ;
  assign y16585 = ~n29888 ;
  assign y16586 = ~1'b0 ;
  assign y16587 = n29889 ;
  assign y16588 = ~1'b0 ;
  assign y16589 = ~1'b0 ;
  assign y16590 = ~n29890 ;
  assign y16591 = ~1'b0 ;
  assign y16592 = ~1'b0 ;
  assign y16593 = ~1'b0 ;
  assign y16594 = ~1'b0 ;
  assign y16595 = n29894 ;
  assign y16596 = n29898 ;
  assign y16597 = ~n29899 ;
  assign y16598 = 1'b0 ;
  assign y16599 = n29901 ;
  assign y16600 = ~n29902 ;
  assign y16601 = n29911 ;
  assign y16602 = ~n29912 ;
  assign y16603 = n29914 ;
  assign y16604 = ~n29915 ;
  assign y16605 = ~n29918 ;
  assign y16606 = n29919 ;
  assign y16607 = n29921 ;
  assign y16608 = ~1'b0 ;
  assign y16609 = n29922 ;
  assign y16610 = n29925 ;
  assign y16611 = ~n29926 ;
  assign y16612 = ~n29929 ;
  assign y16613 = ~1'b0 ;
  assign y16614 = n29931 ;
  assign y16615 = ~n29935 ;
  assign y16616 = ~n29938 ;
  assign y16617 = ~n13393 ;
  assign y16618 = n11316 ;
  assign y16619 = n10320 ;
  assign y16620 = ~n29940 ;
  assign y16621 = n29941 ;
  assign y16622 = ~n29943 ;
  assign y16623 = ~1'b0 ;
  assign y16624 = ~n29947 ;
  assign y16625 = ~1'b0 ;
  assign y16626 = ~n29951 ;
  assign y16627 = ~n29956 ;
  assign y16628 = n29958 ;
  assign y16629 = n29960 ;
  assign y16630 = ~1'b0 ;
  assign y16631 = n29961 ;
  assign y16632 = n29965 ;
  assign y16633 = ~n29970 ;
  assign y16634 = ~n29971 ;
  assign y16635 = ~1'b0 ;
  assign y16636 = n29972 ;
  assign y16637 = 1'b0 ;
  assign y16638 = n29973 ;
  assign y16639 = ~n29979 ;
  assign y16640 = n29980 ;
  assign y16641 = ~n29982 ;
  assign y16642 = ~1'b0 ;
  assign y16643 = ~1'b0 ;
  assign y16644 = ~1'b0 ;
  assign y16645 = ~n29984 ;
  assign y16646 = 1'b0 ;
  assign y16647 = ~1'b0 ;
  assign y16648 = ~n29985 ;
  assign y16649 = ~n26743 ;
  assign y16650 = n29627 ;
  assign y16651 = ~n29986 ;
  assign y16652 = ~n4644 ;
  assign y16653 = ~1'b0 ;
  assign y16654 = ~1'b0 ;
  assign y16655 = 1'b0 ;
  assign y16656 = ~n29989 ;
  assign y16657 = ~n29990 ;
  assign y16658 = ~n29992 ;
  assign y16659 = n29937 ;
  assign y16660 = ~1'b0 ;
  assign y16661 = n29999 ;
  assign y16662 = ~n30006 ;
  assign y16663 = ~n30010 ;
  assign y16664 = ~1'b0 ;
  assign y16665 = ~n6025 ;
  assign y16666 = ~n30011 ;
  assign y16667 = ~n30012 ;
  assign y16668 = ~1'b0 ;
  assign y16669 = ~n30015 ;
  assign y16670 = ~n19196 ;
  assign y16671 = ~1'b0 ;
  assign y16672 = n30019 ;
  assign y16673 = n30020 ;
  assign y16674 = ~n30021 ;
  assign y16675 = n30022 ;
  assign y16676 = ~n30023 ;
  assign y16677 = ~1'b0 ;
  assign y16678 = n30025 ;
  assign y16679 = ~1'b0 ;
  assign y16680 = ~n30027 ;
  assign y16681 = n30029 ;
  assign y16682 = ~1'b0 ;
  assign y16683 = n30032 ;
  assign y16684 = n30033 ;
  assign y16685 = ~1'b0 ;
  assign y16686 = n30039 ;
  assign y16687 = n30047 ;
  assign y16688 = n30050 ;
  assign y16689 = ~1'b0 ;
  assign y16690 = ~n30053 ;
  assign y16691 = ~1'b0 ;
  assign y16692 = n30041 ;
  assign y16693 = n30055 ;
  assign y16694 = n30057 ;
  assign y16695 = ~1'b0 ;
  assign y16696 = ~1'b0 ;
  assign y16697 = ~n30065 ;
  assign y16698 = ~1'b0 ;
  assign y16699 = n30073 ;
  assign y16700 = n17600 ;
  assign y16701 = ~1'b0 ;
  assign y16702 = n30074 ;
  assign y16703 = 1'b0 ;
  assign y16704 = ~1'b0 ;
  assign y16705 = ~n30076 ;
  assign y16706 = ~1'b0 ;
  assign y16707 = ~n30079 ;
  assign y16708 = ~1'b0 ;
  assign y16709 = ~1'b0 ;
  assign y16710 = ~1'b0 ;
  assign y16711 = ~n30081 ;
  assign y16712 = n30083 ;
  assign y16713 = ~n30084 ;
  assign y16714 = ~n30086 ;
  assign y16715 = ~1'b0 ;
  assign y16716 = ~1'b0 ;
  assign y16717 = ~n30088 ;
  assign y16718 = 1'b0 ;
  assign y16719 = ~n30090 ;
  assign y16720 = ~n30092 ;
  assign y16721 = ~n30095 ;
  assign y16722 = ~1'b0 ;
  assign y16723 = n30097 ;
  assign y16724 = ~n30099 ;
  assign y16725 = ~n30106 ;
  assign y16726 = n30108 ;
  assign y16727 = n30110 ;
  assign y16728 = ~1'b0 ;
  assign y16729 = ~1'b0 ;
  assign y16730 = ~1'b0 ;
  assign y16731 = n9203 ;
  assign y16732 = ~n30112 ;
  assign y16733 = ~n15792 ;
  assign y16734 = ~n30117 ;
  assign y16735 = n30118 ;
  assign y16736 = ~n30123 ;
  assign y16737 = n30124 ;
  assign y16738 = ~1'b0 ;
  assign y16739 = n30126 ;
  assign y16740 = n30128 ;
  assign y16741 = ~1'b0 ;
  assign y16742 = ~1'b0 ;
  assign y16743 = ~1'b0 ;
  assign y16744 = ~n30130 ;
  assign y16745 = n30131 ;
  assign y16746 = ~1'b0 ;
  assign y16747 = ~1'b0 ;
  assign y16748 = n30132 ;
  assign y16749 = ~n30136 ;
  assign y16750 = n30137 ;
  assign y16751 = ~n30138 ;
  assign y16752 = ~1'b0 ;
  assign y16753 = ~n17363 ;
  assign y16754 = ~1'b0 ;
  assign y16755 = ~1'b0 ;
  assign y16756 = ~n30144 ;
  assign y16757 = ~n30146 ;
  assign y16758 = n30150 ;
  assign y16759 = ~1'b0 ;
  assign y16760 = n30152 ;
  assign y16761 = ~1'b0 ;
  assign y16762 = ~1'b0 ;
  assign y16763 = n30155 ;
  assign y16764 = ~n22558 ;
  assign y16765 = ~n30157 ;
  assign y16766 = n2348 ;
  assign y16767 = ~1'b0 ;
  assign y16768 = ~1'b0 ;
  assign y16769 = ~n30165 ;
  assign y16770 = ~n30167 ;
  assign y16771 = n7558 ;
  assign y16772 = ~1'b0 ;
  assign y16773 = n30168 ;
  assign y16774 = n30169 ;
  assign y16775 = ~1'b0 ;
  assign y16776 = n30170 ;
  assign y16777 = ~n30175 ;
  assign y16778 = n30176 ;
  assign y16779 = n30177 ;
  assign y16780 = ~1'b0 ;
  assign y16781 = ~n30179 ;
  assign y16782 = ~n30180 ;
  assign y16783 = ~1'b0 ;
  assign y16784 = n30182 ;
  assign y16785 = ~n30184 ;
  assign y16786 = ~n30186 ;
  assign y16787 = ~n30190 ;
  assign y16788 = ~1'b0 ;
  assign y16789 = ~n30195 ;
  assign y16790 = ~n30197 ;
  assign y16791 = ~n30198 ;
  assign y16792 = ~n30202 ;
  assign y16793 = ~n30203 ;
  assign y16794 = n30204 ;
  assign y16795 = ~n30209 ;
  assign y16796 = ~1'b0 ;
  assign y16797 = ~n30213 ;
  assign y16798 = n30217 ;
  assign y16799 = ~n30220 ;
  assign y16800 = ~n25181 ;
  assign y16801 = ~n30221 ;
  assign y16802 = ~n30222 ;
  assign y16803 = ~n30223 ;
  assign y16804 = n30226 ;
  assign y16805 = ~n30228 ;
  assign y16806 = ~n30230 ;
  assign y16807 = n30238 ;
  assign y16808 = ~1'b0 ;
  assign y16809 = n30242 ;
  assign y16810 = ~n30243 ;
  assign y16811 = ~1'b0 ;
  assign y16812 = n23481 ;
  assign y16813 = n30244 ;
  assign y16814 = n30247 ;
  assign y16815 = ~1'b0 ;
  assign y16816 = ~1'b0 ;
  assign y16817 = ~1'b0 ;
  assign y16818 = ~1'b0 ;
  assign y16819 = ~n30251 ;
  assign y16820 = ~1'b0 ;
  assign y16821 = n9576 ;
  assign y16822 = n30255 ;
  assign y16823 = ~1'b0 ;
  assign y16824 = n30260 ;
  assign y16825 = ~n22183 ;
  assign y16826 = n30264 ;
  assign y16827 = n30265 ;
  assign y16828 = n30267 ;
  assign y16829 = ~n30270 ;
  assign y16830 = n30273 ;
  assign y16831 = n30274 ;
  assign y16832 = n30278 ;
  assign y16833 = ~1'b0 ;
  assign y16834 = ~1'b0 ;
  assign y16835 = ~n30279 ;
  assign y16836 = ~n30281 ;
  assign y16837 = ~1'b0 ;
  assign y16838 = n3233 ;
  assign y16839 = ~1'b0 ;
  assign y16840 = ~n30284 ;
  assign y16841 = n30285 ;
  assign y16842 = ~n30287 ;
  assign y16843 = ~n30290 ;
  assign y16844 = n30292 ;
  assign y16845 = ~n30293 ;
  assign y16846 = ~1'b0 ;
  assign y16847 = n30294 ;
  assign y16848 = ~1'b0 ;
  assign y16849 = ~n18324 ;
  assign y16850 = ~n30299 ;
  assign y16851 = n30301 ;
  assign y16852 = ~n30304 ;
  assign y16853 = ~n30308 ;
  assign y16854 = n18635 ;
  assign y16855 = ~n30314 ;
  assign y16856 = ~n30315 ;
  assign y16857 = ~n30317 ;
  assign y16858 = ~n30319 ;
  assign y16859 = ~n30324 ;
  assign y16860 = ~n30326 ;
  assign y16861 = n30329 ;
  assign y16862 = ~n30330 ;
  assign y16863 = ~n30332 ;
  assign y16864 = ~n30333 ;
  assign y16865 = ~1'b0 ;
  assign y16866 = ~n30335 ;
  assign y16867 = ~n30342 ;
  assign y16868 = n30343 ;
  assign y16869 = ~n30346 ;
  assign y16870 = n30351 ;
  assign y16871 = ~1'b0 ;
  assign y16872 = ~1'b0 ;
  assign y16873 = n30353 ;
  assign y16874 = ~1'b0 ;
  assign y16875 = n30356 ;
  assign y16876 = n30360 ;
  assign y16877 = ~1'b0 ;
  assign y16878 = ~n30362 ;
  assign y16879 = ~n30364 ;
  assign y16880 = ~1'b0 ;
  assign y16881 = n30366 ;
  assign y16882 = ~1'b0 ;
  assign y16883 = ~n30369 ;
  assign y16884 = n30372 ;
  assign y16885 = n30375 ;
  assign y16886 = ~n30377 ;
  assign y16887 = n30382 ;
  assign y16888 = n30383 ;
  assign y16889 = ~n30384 ;
  assign y16890 = 1'b0 ;
  assign y16891 = n30385 ;
  assign y16892 = ~n30390 ;
  assign y16893 = ~n30393 ;
  assign y16894 = ~1'b0 ;
  assign y16895 = n30395 ;
  assign y16896 = ~n30396 ;
  assign y16897 = n30397 ;
  assign y16898 = ~n30398 ;
  assign y16899 = ~n30404 ;
  assign y16900 = n30408 ;
  assign y16901 = ~n30409 ;
  assign y16902 = n30410 ;
  assign y16903 = ~n30412 ;
  assign y16904 = ~1'b0 ;
  assign y16905 = ~n30413 ;
  assign y16906 = ~n30415 ;
  assign y16907 = n30418 ;
  assign y16908 = n30419 ;
  assign y16909 = ~n15086 ;
  assign y16910 = n30426 ;
  assign y16911 = n30427 ;
  assign y16912 = n2562 ;
  assign y16913 = ~1'b0 ;
  assign y16914 = ~1'b0 ;
  assign y16915 = ~n1112 ;
  assign y16916 = ~1'b0 ;
  assign y16917 = ~1'b0 ;
  assign y16918 = ~n22935 ;
  assign y16919 = ~n30435 ;
  assign y16920 = ~1'b0 ;
  assign y16921 = n30438 ;
  assign y16922 = ~n30441 ;
  assign y16923 = ~n30443 ;
  assign y16924 = n30444 ;
  assign y16925 = ~n30445 ;
  assign y16926 = n30448 ;
  assign y16927 = ~1'b0 ;
  assign y16928 = n30449 ;
  assign y16929 = n30450 ;
  assign y16930 = ~n30451 ;
  assign y16931 = n30453 ;
  assign y16932 = ~n30462 ;
  assign y16933 = ~1'b0 ;
  assign y16934 = ~n30466 ;
  assign y16935 = ~1'b0 ;
  assign y16936 = ~1'b0 ;
  assign y16937 = n30468 ;
  assign y16938 = n30469 ;
  assign y16939 = ~n30472 ;
  assign y16940 = ~n30473 ;
  assign y16941 = ~n30474 ;
  assign y16942 = n30478 ;
  assign y16943 = ~n30480 ;
  assign y16944 = ~1'b0 ;
  assign y16945 = ~n30486 ;
  assign y16946 = ~n30487 ;
  assign y16947 = ~n30488 ;
  assign y16948 = n30490 ;
  assign y16949 = ~1'b0 ;
  assign y16950 = ~1'b0 ;
  assign y16951 = ~1'b0 ;
  assign y16952 = n30495 ;
  assign y16953 = n30501 ;
  assign y16954 = ~n30502 ;
  assign y16955 = ~1'b0 ;
  assign y16956 = n525 ;
  assign y16957 = ~1'b0 ;
  assign y16958 = 1'b0 ;
  assign y16959 = n30506 ;
  assign y16960 = ~n30512 ;
  assign y16961 = ~1'b0 ;
  assign y16962 = ~n9037 ;
  assign y16963 = ~n30514 ;
  assign y16964 = n30515 ;
  assign y16965 = ~1'b0 ;
  assign y16966 = n30517 ;
  assign y16967 = n30520 ;
  assign y16968 = n30523 ;
  assign y16969 = ~n10736 ;
  assign y16970 = ~1'b0 ;
  assign y16971 = ~1'b0 ;
  assign y16972 = ~1'b0 ;
  assign y16973 = n30524 ;
  assign y16974 = n30533 ;
  assign y16975 = ~n30538 ;
  assign y16976 = ~1'b0 ;
  assign y16977 = ~n30540 ;
  assign y16978 = ~n30541 ;
  assign y16979 = n30542 ;
  assign y16980 = ~n30545 ;
  assign y16981 = ~n25867 ;
  assign y16982 = n30548 ;
  assign y16983 = ~1'b0 ;
  assign y16984 = ~n30549 ;
  assign y16985 = n30552 ;
  assign y16986 = n30553 ;
  assign y16987 = ~n30554 ;
  assign y16988 = ~n30555 ;
  assign y16989 = ~n13251 ;
  assign y16990 = n30558 ;
  assign y16991 = ~n30561 ;
  assign y16992 = ~n30564 ;
  assign y16993 = ~1'b0 ;
  assign y16994 = n30565 ;
  assign y16995 = n17482 ;
  assign y16996 = ~1'b0 ;
  assign y16997 = n30566 ;
  assign y16998 = ~1'b0 ;
  assign y16999 = n30568 ;
  assign y17000 = ~1'b0 ;
  assign y17001 = ~1'b0 ;
  assign y17002 = ~n6437 ;
  assign y17003 = ~n30569 ;
  assign y17004 = ~n30571 ;
  assign y17005 = n30573 ;
  assign y17006 = ~1'b0 ;
  assign y17007 = 1'b0 ;
  assign y17008 = n30575 ;
  assign y17009 = n23063 ;
  assign y17010 = ~1'b0 ;
  assign y17011 = ~n30579 ;
  assign y17012 = n30580 ;
  assign y17013 = n30582 ;
  assign y17014 = ~1'b0 ;
  assign y17015 = ~n30584 ;
  assign y17016 = n30585 ;
  assign y17017 = n30588 ;
  assign y17018 = ~n30591 ;
  assign y17019 = n30593 ;
  assign y17020 = ~1'b0 ;
  assign y17021 = ~n21331 ;
  assign y17022 = n30594 ;
  assign y17023 = n30596 ;
  assign y17024 = ~n30609 ;
  assign y17025 = n30610 ;
  assign y17026 = n30618 ;
  assign y17027 = n30620 ;
  assign y17028 = n15319 ;
  assign y17029 = ~n30622 ;
  assign y17030 = ~1'b0 ;
  assign y17031 = ~1'b0 ;
  assign y17032 = n30625 ;
  assign y17033 = n30626 ;
  assign y17034 = ~n30628 ;
  assign y17035 = ~1'b0 ;
  assign y17036 = ~1'b0 ;
  assign y17037 = ~n30629 ;
  assign y17038 = ~n30634 ;
  assign y17039 = ~1'b0 ;
  assign y17040 = 1'b0 ;
  assign y17041 = ~n30635 ;
  assign y17042 = ~1'b0 ;
  assign y17043 = n30637 ;
  assign y17044 = ~1'b0 ;
  assign y17045 = n30639 ;
  assign y17046 = n30642 ;
  assign y17047 = ~n30644 ;
  assign y17048 = n30656 ;
  assign y17049 = ~n30664 ;
  assign y17050 = ~n30665 ;
  assign y17051 = ~n30666 ;
  assign y17052 = ~n27261 ;
  assign y17053 = n30668 ;
  assign y17054 = ~n30674 ;
  assign y17055 = n30678 ;
  assign y17056 = ~n30681 ;
  assign y17057 = ~1'b0 ;
  assign y17058 = n30682 ;
  assign y17059 = n30683 ;
  assign y17060 = ~n30686 ;
  assign y17061 = n30690 ;
  assign y17062 = n30692 ;
  assign y17063 = ~n30696 ;
  assign y17064 = ~n30698 ;
  assign y17065 = 1'b0 ;
  assign y17066 = ~n16314 ;
  assign y17067 = 1'b0 ;
  assign y17068 = n30699 ;
  assign y17069 = ~n30701 ;
  assign y17070 = ~1'b0 ;
  assign y17071 = ~1'b0 ;
  assign y17072 = n30704 ;
  assign y17073 = ~n30705 ;
  assign y17074 = n30710 ;
  assign y17075 = n30711 ;
  assign y17076 = ~n30712 ;
  assign y17077 = n30714 ;
  assign y17078 = ~1'b0 ;
  assign y17079 = ~n30726 ;
  assign y17080 = ~n30727 ;
  assign y17081 = ~n30729 ;
  assign y17082 = ~n30731 ;
  assign y17083 = ~1'b0 ;
  assign y17084 = ~n30735 ;
  assign y17085 = n30738 ;
  assign y17086 = n30743 ;
  assign y17087 = n30750 ;
  assign y17088 = n30751 ;
  assign y17089 = n17253 ;
  assign y17090 = 1'b0 ;
  assign y17091 = ~1'b0 ;
  assign y17092 = ~1'b0 ;
  assign y17093 = ~1'b0 ;
  assign y17094 = n30754 ;
  assign y17095 = n30755 ;
  assign y17096 = ~1'b0 ;
  assign y17097 = n30761 ;
  assign y17098 = ~n30765 ;
  assign y17099 = 1'b0 ;
  assign y17100 = ~n30767 ;
  assign y17101 = n30771 ;
  assign y17102 = n30773 ;
  assign y17103 = n30779 ;
  assign y17104 = n30783 ;
  assign y17105 = n30784 ;
  assign y17106 = n30785 ;
  assign y17107 = ~n30788 ;
  assign y17108 = ~n30790 ;
  assign y17109 = ~1'b0 ;
  assign y17110 = n30791 ;
  assign y17111 = ~1'b0 ;
  assign y17112 = n30792 ;
  assign y17113 = n30794 ;
  assign y17114 = ~1'b0 ;
  assign y17115 = n30795 ;
  assign y17116 = ~1'b0 ;
  assign y17117 = n30802 ;
  assign y17118 = ~1'b0 ;
  assign y17119 = ~1'b0 ;
  assign y17120 = ~n30803 ;
  assign y17121 = ~n30807 ;
  assign y17122 = ~n30813 ;
  assign y17123 = ~n30819 ;
  assign y17124 = n30821 ;
  assign y17125 = n30822 ;
  assign y17126 = n30825 ;
  assign y17127 = n30826 ;
  assign y17128 = n30828 ;
  assign y17129 = n30829 ;
  assign y17130 = ~n30832 ;
  assign y17131 = n30834 ;
  assign y17132 = n30835 ;
  assign y17133 = ~1'b0 ;
  assign y17134 = ~1'b0 ;
  assign y17135 = n30836 ;
  assign y17136 = ~1'b0 ;
  assign y17137 = n30837 ;
  assign y17138 = ~n30838 ;
  assign y17139 = ~1'b0 ;
  assign y17140 = ~n30839 ;
  assign y17141 = ~n30845 ;
  assign y17142 = ~1'b0 ;
  assign y17143 = ~n30846 ;
  assign y17144 = 1'b0 ;
  assign y17145 = ~1'b0 ;
  assign y17146 = ~n30851 ;
  assign y17147 = ~n30852 ;
  assign y17148 = ~n30853 ;
  assign y17149 = ~1'b0 ;
  assign y17150 = ~1'b0 ;
  assign y17151 = n30858 ;
  assign y17152 = ~1'b0 ;
  assign y17153 = n30861 ;
  assign y17154 = n30864 ;
  assign y17155 = ~n30870 ;
  assign y17156 = ~1'b0 ;
  assign y17157 = n30875 ;
  assign y17158 = ~1'b0 ;
  assign y17159 = n30877 ;
  assign y17160 = ~n30881 ;
  assign y17161 = n27327 ;
  assign y17162 = ~1'b0 ;
  assign y17163 = ~n30882 ;
  assign y17164 = ~1'b0 ;
  assign y17165 = n30888 ;
  assign y17166 = n30890 ;
  assign y17167 = ~n30891 ;
  assign y17168 = ~n30893 ;
  assign y17169 = n30895 ;
  assign y17170 = ~1'b0 ;
  assign y17171 = ~1'b0 ;
  assign y17172 = ~n30897 ;
  assign y17173 = ~n30900 ;
  assign y17174 = ~n30901 ;
  assign y17175 = n30902 ;
  assign y17176 = n30903 ;
  assign y17177 = ~1'b0 ;
  assign y17178 = ~1'b0 ;
  assign y17179 = ~n30908 ;
  assign y17180 = ~1'b0 ;
  assign y17181 = ~n30910 ;
  assign y17182 = n30915 ;
  assign y17183 = ~1'b0 ;
  assign y17184 = ~1'b0 ;
  assign y17185 = n12326 ;
  assign y17186 = n7504 ;
  assign y17187 = n30917 ;
  assign y17188 = ~1'b0 ;
  assign y17189 = ~n30920 ;
  assign y17190 = n30926 ;
  assign y17191 = ~1'b0 ;
  assign y17192 = ~1'b0 ;
  assign y17193 = ~1'b0 ;
  assign y17194 = n30928 ;
  assign y17195 = ~1'b0 ;
  assign y17196 = n30931 ;
  assign y17197 = ~1'b0 ;
  assign y17198 = n30934 ;
  assign y17199 = ~n30940 ;
  assign y17200 = ~n30943 ;
  assign y17201 = n11789 ;
  assign y17202 = n30944 ;
  assign y17203 = n30945 ;
  assign y17204 = ~1'b0 ;
  assign y17205 = ~1'b0 ;
  assign y17206 = ~1'b0 ;
  assign y17207 = n29857 ;
  assign y17208 = ~1'b0 ;
  assign y17209 = n30947 ;
  assign y17210 = ~n30948 ;
  assign y17211 = ~n30957 ;
  assign y17212 = ~n30958 ;
  assign y17213 = ~1'b0 ;
  assign y17214 = ~n30961 ;
  assign y17215 = n30962 ;
  assign y17216 = ~n30964 ;
  assign y17217 = n30965 ;
  assign y17218 = n30966 ;
  assign y17219 = ~n30967 ;
  assign y17220 = n30969 ;
  assign y17221 = ~n30970 ;
  assign y17222 = ~1'b0 ;
  assign y17223 = n30971 ;
  assign y17224 = n30972 ;
  assign y17225 = ~1'b0 ;
  assign y17226 = ~1'b0 ;
  assign y17227 = ~1'b0 ;
  assign y17228 = n30974 ;
  assign y17229 = n30976 ;
  assign y17230 = n30979 ;
  assign y17231 = ~n30980 ;
  assign y17232 = ~1'b0 ;
  assign y17233 = ~1'b0 ;
  assign y17234 = ~1'b0 ;
  assign y17235 = n28280 ;
  assign y17236 = n30986 ;
  assign y17237 = ~n30987 ;
  assign y17238 = ~1'b0 ;
  assign y17239 = ~n30988 ;
  assign y17240 = ~n5930 ;
  assign y17241 = ~n30989 ;
  assign y17242 = ~1'b0 ;
  assign y17243 = n31001 ;
  assign y17244 = ~1'b0 ;
  assign y17245 = ~1'b0 ;
  assign y17246 = ~n31005 ;
  assign y17247 = ~n31009 ;
  assign y17248 = n31011 ;
  assign y17249 = ~n31014 ;
  assign y17250 = ~1'b0 ;
  assign y17251 = ~n31016 ;
  assign y17252 = ~1'b0 ;
  assign y17253 = ~1'b0 ;
  assign y17254 = ~n31018 ;
  assign y17255 = ~1'b0 ;
  assign y17256 = n31019 ;
  assign y17257 = ~n31020 ;
  assign y17258 = n31025 ;
  assign y17259 = ~n31029 ;
  assign y17260 = ~n31033 ;
  assign y17261 = ~1'b0 ;
  assign y17262 = n31034 ;
  assign y17263 = ~n31035 ;
  assign y17264 = ~1'b0 ;
  assign y17265 = n31038 ;
  assign y17266 = ~n31041 ;
  assign y17267 = n31043 ;
  assign y17268 = ~1'b0 ;
  assign y17269 = ~1'b0 ;
  assign y17270 = ~1'b0 ;
  assign y17271 = n31046 ;
  assign y17272 = ~1'b0 ;
  assign y17273 = ~n31048 ;
  assign y17274 = n21806 ;
  assign y17275 = ~n31050 ;
  assign y17276 = n31053 ;
  assign y17277 = n31055 ;
  assign y17278 = ~n31062 ;
  assign y17279 = ~1'b0 ;
  assign y17280 = ~n31063 ;
  assign y17281 = 1'b0 ;
  assign y17282 = n31064 ;
  assign y17283 = n10171 ;
  assign y17284 = 1'b0 ;
  assign y17285 = ~1'b0 ;
  assign y17286 = ~1'b0 ;
  assign y17287 = n31066 ;
  assign y17288 = ~n31068 ;
  assign y17289 = ~n31074 ;
  assign y17290 = ~n31076 ;
  assign y17291 = ~1'b0 ;
  assign y17292 = n31078 ;
  assign y17293 = ~n31082 ;
  assign y17294 = ~n31084 ;
  assign y17295 = ~1'b0 ;
  assign y17296 = ~1'b0 ;
  assign y17297 = n31087 ;
  assign y17298 = ~n31088 ;
  assign y17299 = ~n31090 ;
  assign y17300 = ~n31094 ;
  assign y17301 = ~1'b0 ;
  assign y17302 = ~n31100 ;
  assign y17303 = ~n31101 ;
  assign y17304 = ~n31104 ;
  assign y17305 = ~1'b0 ;
  assign y17306 = 1'b0 ;
  assign y17307 = ~1'b0 ;
  assign y17308 = ~1'b0 ;
  assign y17309 = ~1'b0 ;
  assign y17310 = ~1'b0 ;
  assign y17311 = n31106 ;
  assign y17312 = ~1'b0 ;
  assign y17313 = n31107 ;
  assign y17314 = n31109 ;
  assign y17315 = n31110 ;
  assign y17316 = ~1'b0 ;
  assign y17317 = ~n31113 ;
  assign y17318 = n31115 ;
  assign y17319 = ~n31117 ;
  assign y17320 = ~1'b0 ;
  assign y17321 = ~n31118 ;
  assign y17322 = ~n31119 ;
  assign y17323 = n21145 ;
  assign y17324 = ~1'b0 ;
  assign y17325 = ~n31122 ;
  assign y17326 = n31127 ;
  assign y17327 = ~1'b0 ;
  assign y17328 = n31130 ;
  assign y17329 = ~n31132 ;
  assign y17330 = ~1'b0 ;
  assign y17331 = ~1'b0 ;
  assign y17332 = n31133 ;
  assign y17333 = ~n31136 ;
  assign y17334 = n31141 ;
  assign y17335 = n31143 ;
  assign y17336 = n31145 ;
  assign y17337 = ~n4377 ;
  assign y17338 = ~1'b0 ;
  assign y17339 = ~n31147 ;
  assign y17340 = ~1'b0 ;
  assign y17341 = n31162 ;
  assign y17342 = ~n31168 ;
  assign y17343 = n31173 ;
  assign y17344 = ~n31175 ;
  assign y17345 = ~1'b0 ;
  assign y17346 = n31178 ;
  assign y17347 = ~n13687 ;
  assign y17348 = ~n31185 ;
  assign y17349 = n31189 ;
  assign y17350 = ~1'b0 ;
  assign y17351 = ~1'b0 ;
  assign y17352 = ~1'b0 ;
  assign y17353 = ~n31194 ;
  assign y17354 = ~n31195 ;
  assign y17355 = ~1'b0 ;
  assign y17356 = n31200 ;
  assign y17357 = n10684 ;
  assign y17358 = n31202 ;
  assign y17359 = ~n31204 ;
  assign y17360 = ~1'b0 ;
  assign y17361 = n31211 ;
  assign y17362 = ~1'b0 ;
  assign y17363 = n31212 ;
  assign y17364 = ~n31215 ;
  assign y17365 = ~1'b0 ;
  assign y17366 = ~n31219 ;
  assign y17367 = n31221 ;
  assign y17368 = ~1'b0 ;
  assign y17369 = ~1'b0 ;
  assign y17370 = n31222 ;
  assign y17371 = n11514 ;
  assign y17372 = ~n31223 ;
  assign y17373 = n31224 ;
  assign y17374 = ~1'b0 ;
  assign y17375 = ~n31229 ;
  assign y17376 = ~n31232 ;
  assign y17377 = ~n31236 ;
  assign y17378 = ~n31246 ;
  assign y17379 = ~n31249 ;
  assign y17380 = n31252 ;
  assign y17381 = n31253 ;
  assign y17382 = ~n31256 ;
  assign y17383 = ~n31259 ;
  assign y17384 = n31260 ;
  assign y17385 = n31266 ;
  assign y17386 = ~n31268 ;
  assign y17387 = n31270 ;
  assign y17388 = n31271 ;
  assign y17389 = n31272 ;
  assign y17390 = n31274 ;
  assign y17391 = ~1'b0 ;
  assign y17392 = ~1'b0 ;
  assign y17393 = ~n31278 ;
  assign y17394 = n31279 ;
  assign y17395 = ~n31281 ;
  assign y17396 = ~n31290 ;
  assign y17397 = ~1'b0 ;
  assign y17398 = n31292 ;
  assign y17399 = n31293 ;
  assign y17400 = n31294 ;
  assign y17401 = 1'b0 ;
  assign y17402 = ~n31300 ;
  assign y17403 = n31302 ;
  assign y17404 = n31304 ;
  assign y17405 = ~n31306 ;
  assign y17406 = n31308 ;
  assign y17407 = n31310 ;
  assign y17408 = n3166 ;
  assign y17409 = ~1'b0 ;
  assign y17410 = n31314 ;
  assign y17411 = ~n6488 ;
  assign y17412 = n31315 ;
  assign y17413 = n16298 ;
  assign y17414 = n31319 ;
  assign y17415 = ~n31326 ;
  assign y17416 = ~n31328 ;
  assign y17417 = ~n31332 ;
  assign y17418 = n31336 ;
  assign y17419 = n31337 ;
  assign y17420 = 1'b0 ;
  assign y17421 = ~n31344 ;
  assign y17422 = n31347 ;
  assign y17423 = ~n31349 ;
  assign y17424 = 1'b0 ;
  assign y17425 = n31350 ;
  assign y17426 = n31353 ;
  assign y17427 = n31359 ;
  assign y17428 = n31361 ;
  assign y17429 = ~n31364 ;
  assign y17430 = ~1'b0 ;
  assign y17431 = n31366 ;
  assign y17432 = ~n31368 ;
  assign y17433 = ~n31371 ;
  assign y17434 = ~n31372 ;
  assign y17435 = ~n31374 ;
  assign y17436 = n31375 ;
  assign y17437 = ~n7207 ;
  assign y17438 = ~n31379 ;
  assign y17439 = ~1'b0 ;
  assign y17440 = ~n31382 ;
  assign y17441 = n31384 ;
  assign y17442 = n31385 ;
  assign y17443 = n31386 ;
  assign y17444 = ~n31388 ;
  assign y17445 = n31390 ;
  assign y17446 = ~1'b0 ;
  assign y17447 = ~n31393 ;
  assign y17448 = n18392 ;
  assign y17449 = ~1'b0 ;
  assign y17450 = ~1'b0 ;
  assign y17451 = ~1'b0 ;
  assign y17452 = ~n31395 ;
  assign y17453 = n31398 ;
  assign y17454 = n31400 ;
  assign y17455 = n31402 ;
  assign y17456 = ~1'b0 ;
  assign y17457 = ~n31405 ;
  assign y17458 = ~n31416 ;
  assign y17459 = n31417 ;
  assign y17460 = ~1'b0 ;
  assign y17461 = n26555 ;
  assign y17462 = n31418 ;
  assign y17463 = n31420 ;
  assign y17464 = n31422 ;
  assign y17465 = ~1'b0 ;
  assign y17466 = ~n31427 ;
  assign y17467 = ~1'b0 ;
  assign y17468 = ~n31428 ;
  assign y17469 = n17027 ;
  assign y17470 = ~1'b0 ;
  assign y17471 = ~n25034 ;
  assign y17472 = ~n31430 ;
  assign y17473 = ~1'b0 ;
  assign y17474 = n31432 ;
  assign y17475 = n31434 ;
  assign y17476 = n31435 ;
  assign y17477 = n31437 ;
  assign y17478 = ~1'b0 ;
  assign y17479 = ~n31441 ;
  assign y17480 = ~1'b0 ;
  assign y17481 = n31446 ;
  assign y17482 = n31447 ;
  assign y17483 = ~1'b0 ;
  assign y17484 = ~n31452 ;
  assign y17485 = ~1'b0 ;
  assign y17486 = ~1'b0 ;
  assign y17487 = ~n31454 ;
  assign y17488 = n31459 ;
  assign y17489 = ~n31461 ;
  assign y17490 = ~1'b0 ;
  assign y17491 = ~n7429 ;
  assign y17492 = n31463 ;
  assign y17493 = ~1'b0 ;
  assign y17494 = ~1'b0 ;
  assign y17495 = n31472 ;
  assign y17496 = n31475 ;
  assign y17497 = ~1'b0 ;
  assign y17498 = n1363 ;
  assign y17499 = ~1'b0 ;
  assign y17500 = ~1'b0 ;
  assign y17501 = n31478 ;
  assign y17502 = ~1'b0 ;
  assign y17503 = ~1'b0 ;
  assign y17504 = ~1'b0 ;
  assign y17505 = n31485 ;
  assign y17506 = ~n31490 ;
  assign y17507 = ~n31492 ;
  assign y17508 = ~n31495 ;
  assign y17509 = n31496 ;
  assign y17510 = ~n31501 ;
  assign y17511 = ~1'b0 ;
  assign y17512 = n31504 ;
  assign y17513 = ~n31505 ;
  assign y17514 = n23966 ;
  assign y17515 = ~n31508 ;
  assign y17516 = ~n13342 ;
  assign y17517 = n31509 ;
  assign y17518 = n31511 ;
  assign y17519 = 1'b0 ;
  assign y17520 = ~1'b0 ;
  assign y17521 = n31517 ;
  assign y17522 = n12391 ;
  assign y17523 = n31523 ;
  assign y17524 = ~1'b0 ;
  assign y17525 = n31524 ;
  assign y17526 = ~n31528 ;
  assign y17527 = n31533 ;
  assign y17528 = n31535 ;
  assign y17529 = ~1'b0 ;
  assign y17530 = ~n31541 ;
  assign y17531 = n31542 ;
  assign y17532 = n31543 ;
  assign y17533 = n31544 ;
  assign y17534 = ~n31546 ;
  assign y17535 = ~1'b0 ;
  assign y17536 = ~1'b0 ;
  assign y17537 = n31547 ;
  assign y17538 = n31551 ;
  assign y17539 = ~n31556 ;
  assign y17540 = n31558 ;
  assign y17541 = ~1'b0 ;
  assign y17542 = n31559 ;
  assign y17543 = 1'b0 ;
  assign y17544 = ~1'b0 ;
  assign y17545 = n31560 ;
  assign y17546 = ~1'b0 ;
  assign y17547 = ~1'b0 ;
  assign y17548 = n31561 ;
  assign y17549 = ~1'b0 ;
  assign y17550 = ~n31562 ;
  assign y17551 = n31567 ;
  assign y17552 = n31569 ;
  assign y17553 = 1'b0 ;
  assign y17554 = ~n31579 ;
  assign y17555 = ~n5497 ;
  assign y17556 = n31582 ;
  assign y17557 = 1'b0 ;
  assign y17558 = ~1'b0 ;
  assign y17559 = n31584 ;
  assign y17560 = n31585 ;
  assign y17561 = n31586 ;
  assign y17562 = ~1'b0 ;
  assign y17563 = n31587 ;
  assign y17564 = ~n31589 ;
  assign y17565 = ~n31593 ;
  assign y17566 = ~1'b0 ;
  assign y17567 = ~1'b0 ;
  assign y17568 = ~n31595 ;
  assign y17569 = ~n31596 ;
  assign y17570 = ~1'b0 ;
  assign y17571 = n31600 ;
  assign y17572 = n31604 ;
  assign y17573 = ~n31607 ;
  assign y17574 = ~n31611 ;
  assign y17575 = ~n31612 ;
  assign y17576 = ~n31615 ;
  assign y17577 = ~n31616 ;
  assign y17578 = ~n31618 ;
  assign y17579 = ~n31619 ;
  assign y17580 = ~n31621 ;
  assign y17581 = n31624 ;
  assign y17582 = ~1'b0 ;
  assign y17583 = ~1'b0 ;
  assign y17584 = ~1'b0 ;
  assign y17585 = ~n31628 ;
  assign y17586 = 1'b0 ;
  assign y17587 = n31631 ;
  assign y17588 = ~n710 ;
  assign y17589 = n31632 ;
  assign y17590 = n31634 ;
  assign y17591 = ~n31636 ;
  assign y17592 = n31637 ;
  assign y17593 = 1'b0 ;
  assign y17594 = n4461 ;
  assign y17595 = ~1'b0 ;
  assign y17596 = n31641 ;
  assign y17597 = ~n31644 ;
  assign y17598 = n31648 ;
  assign y17599 = ~1'b0 ;
  assign y17600 = n31649 ;
  assign y17601 = ~1'b0 ;
  assign y17602 = n31650 ;
  assign y17603 = ~1'b0 ;
  assign y17604 = ~1'b0 ;
  assign y17605 = ~n5811 ;
  assign y17606 = n31651 ;
  assign y17607 = n31653 ;
  assign y17608 = n31655 ;
  assign y17609 = n31656 ;
  assign y17610 = n31659 ;
  assign y17611 = ~n31670 ;
  assign y17612 = n31675 ;
  assign y17613 = ~1'b0 ;
  assign y17614 = n31676 ;
  assign y17615 = ~1'b0 ;
  assign y17616 = 1'b0 ;
  assign y17617 = ~n31678 ;
  assign y17618 = ~1'b0 ;
  assign y17619 = ~n31680 ;
  assign y17620 = ~1'b0 ;
  assign y17621 = ~n31684 ;
  assign y17622 = ~n31685 ;
  assign y17623 = ~n12687 ;
  assign y17624 = n31686 ;
  assign y17625 = ~1'b0 ;
  assign y17626 = n31704 ;
  assign y17627 = ~n31707 ;
  assign y17628 = ~1'b0 ;
  assign y17629 = ~1'b0 ;
  assign y17630 = n31708 ;
  assign y17631 = ~n31709 ;
  assign y17632 = ~1'b0 ;
  assign y17633 = ~1'b0 ;
  assign y17634 = ~1'b0 ;
  assign y17635 = ~n31710 ;
  assign y17636 = ~1'b0 ;
  assign y17637 = ~n31712 ;
  assign y17638 = n25361 ;
  assign y17639 = n31714 ;
  assign y17640 = ~1'b0 ;
  assign y17641 = ~n31717 ;
  assign y17642 = n31719 ;
  assign y17643 = ~n31722 ;
  assign y17644 = ~1'b0 ;
  assign y17645 = ~n31726 ;
  assign y17646 = n31731 ;
  assign y17647 = n31732 ;
  assign y17648 = n31734 ;
  assign y17649 = ~1'b0 ;
  assign y17650 = ~1'b0 ;
  assign y17651 = ~1'b0 ;
  assign y17652 = n31737 ;
  assign y17653 = ~n31738 ;
  assign y17654 = ~n31739 ;
  assign y17655 = n31740 ;
  assign y17656 = ~n31742 ;
  assign y17657 = n31745 ;
  assign y17658 = ~n31751 ;
  assign y17659 = ~n31752 ;
  assign y17660 = n31753 ;
  assign y17661 = ~n31759 ;
  assign y17662 = ~1'b0 ;
  assign y17663 = ~n31763 ;
  assign y17664 = ~n31764 ;
  assign y17665 = n31765 ;
  assign y17666 = n31769 ;
  assign y17667 = n31770 ;
  assign y17668 = ~1'b0 ;
  assign y17669 = ~n31773 ;
  assign y17670 = ~n31774 ;
  assign y17671 = ~1'b0 ;
  assign y17672 = n31780 ;
  assign y17673 = n31783 ;
  assign y17674 = n31784 ;
  assign y17675 = 1'b0 ;
  assign y17676 = n31787 ;
  assign y17677 = n31791 ;
  assign y17678 = n31792 ;
  assign y17679 = n31799 ;
  assign y17680 = ~n31801 ;
  assign y17681 = ~n31802 ;
  assign y17682 = n31804 ;
  assign y17683 = 1'b0 ;
  assign y17684 = ~1'b0 ;
  assign y17685 = ~1'b0 ;
  assign y17686 = ~n31806 ;
  assign y17687 = ~n31807 ;
  assign y17688 = ~n31809 ;
  assign y17689 = n31811 ;
  assign y17690 = ~1'b0 ;
  assign y17691 = n31814 ;
  assign y17692 = n31820 ;
  assign y17693 = ~1'b0 ;
  assign y17694 = ~n31822 ;
  assign y17695 = ~1'b0 ;
  assign y17696 = ~n31826 ;
  assign y17697 = ~n31828 ;
  assign y17698 = ~n31830 ;
  assign y17699 = n31832 ;
  assign y17700 = ~1'b0 ;
  assign y17701 = n31835 ;
  assign y17702 = ~n30008 ;
  assign y17703 = ~1'b0 ;
  assign y17704 = ~1'b0 ;
  assign y17705 = ~n31837 ;
  assign y17706 = ~n31838 ;
  assign y17707 = ~n31840 ;
  assign y17708 = ~n31843 ;
  assign y17709 = n31844 ;
  assign y17710 = ~1'b0 ;
  assign y17711 = ~n31845 ;
  assign y17712 = ~n31846 ;
  assign y17713 = n31847 ;
  assign y17714 = n31855 ;
  assign y17715 = ~n31856 ;
  assign y17716 = n31857 ;
  assign y17717 = ~n31861 ;
  assign y17718 = ~1'b0 ;
  assign y17719 = ~n31864 ;
  assign y17720 = ~1'b0 ;
  assign y17721 = ~n31866 ;
  assign y17722 = n7999 ;
  assign y17723 = n31868 ;
  assign y17724 = ~n31869 ;
  assign y17725 = ~n31871 ;
  assign y17726 = ~1'b0 ;
  assign y17727 = ~1'b0 ;
  assign y17728 = n31873 ;
  assign y17729 = n31874 ;
  assign y17730 = n31876 ;
  assign y17731 = n31877 ;
  assign y17732 = ~n31886 ;
  assign y17733 = n31889 ;
  assign y17734 = n31892 ;
  assign y17735 = ~1'b0 ;
  assign y17736 = ~1'b0 ;
  assign y17737 = n31894 ;
  assign y17738 = n31896 ;
  assign y17739 = 1'b0 ;
  assign y17740 = ~1'b0 ;
  assign y17741 = n31900 ;
  assign y17742 = ~n31904 ;
  assign y17743 = ~n31905 ;
  assign y17744 = ~1'b0 ;
  assign y17745 = n31908 ;
  assign y17746 = ~n31909 ;
  assign y17747 = ~1'b0 ;
  assign y17748 = ~n31911 ;
  assign y17749 = n1119 ;
  assign y17750 = ~n31913 ;
  assign y17751 = n25289 ;
  assign y17752 = ~1'b0 ;
  assign y17753 = ~1'b0 ;
  assign y17754 = ~n31915 ;
  assign y17755 = ~1'b0 ;
  assign y17756 = 1'b0 ;
  assign y17757 = ~n31916 ;
  assign y17758 = ~1'b0 ;
  assign y17759 = ~1'b0 ;
  assign y17760 = ~n31922 ;
  assign y17761 = ~1'b0 ;
  assign y17762 = n31924 ;
  assign y17763 = ~n31926 ;
  assign y17764 = ~1'b0 ;
  assign y17765 = ~n31928 ;
  assign y17766 = ~n31930 ;
  assign y17767 = ~n31934 ;
  assign y17768 = ~n31935 ;
  assign y17769 = n31937 ;
  assign y17770 = n31941 ;
  assign y17771 = n31945 ;
  assign y17772 = ~n31946 ;
  assign y17773 = ~1'b0 ;
  assign y17774 = ~n31949 ;
  assign y17775 = ~1'b0 ;
  assign y17776 = ~1'b0 ;
  assign y17777 = ~n31950 ;
  assign y17778 = ~n31953 ;
  assign y17779 = ~1'b0 ;
  assign y17780 = ~n31955 ;
  assign y17781 = ~1'b0 ;
  assign y17782 = ~1'b0 ;
  assign y17783 = ~1'b0 ;
  assign y17784 = ~1'b0 ;
  assign y17785 = ~1'b0 ;
  assign y17786 = ~n31958 ;
  assign y17787 = ~1'b0 ;
  assign y17788 = n31964 ;
  assign y17789 = ~1'b0 ;
  assign y17790 = ~1'b0 ;
  assign y17791 = ~1'b0 ;
  assign y17792 = n31966 ;
  assign y17793 = n31967 ;
  assign y17794 = ~n31968 ;
  assign y17795 = ~1'b0 ;
  assign y17796 = n31971 ;
  assign y17797 = n31974 ;
  assign y17798 = ~n31976 ;
  assign y17799 = ~1'b0 ;
  assign y17800 = n31979 ;
  assign y17801 = n31981 ;
  assign y17802 = ~1'b0 ;
  assign y17803 = n31982 ;
  assign y17804 = ~1'b0 ;
  assign y17805 = ~n24583 ;
  assign y17806 = n31983 ;
  assign y17807 = ~n31984 ;
  assign y17808 = ~1'b0 ;
  assign y17809 = n14122 ;
  assign y17810 = n31985 ;
  assign y17811 = ~n22974 ;
  assign y17812 = ~n31987 ;
  assign y17813 = ~1'b0 ;
  assign y17814 = ~1'b0 ;
  assign y17815 = ~n31989 ;
  assign y17816 = ~1'b0 ;
  assign y17817 = ~1'b0 ;
  assign y17818 = n31990 ;
  assign y17819 = ~n31992 ;
  assign y17820 = n31994 ;
  assign y17821 = n31995 ;
  assign y17822 = ~n31996 ;
  assign y17823 = ~n13860 ;
  assign y17824 = n31997 ;
  assign y17825 = n32001 ;
  assign y17826 = ~n32003 ;
  assign y17827 = ~n32005 ;
  assign y17828 = 1'b0 ;
  assign y17829 = ~n32006 ;
  assign y17830 = ~1'b0 ;
  assign y17831 = ~1'b0 ;
  assign y17832 = ~1'b0 ;
  assign y17833 = ~n32007 ;
  assign y17834 = ~n32008 ;
  assign y17835 = n13551 ;
  assign y17836 = n32012 ;
  assign y17837 = n32022 ;
  assign y17838 = n32024 ;
  assign y17839 = n32026 ;
  assign y17840 = ~n32028 ;
  assign y17841 = n32035 ;
  assign y17842 = ~1'b0 ;
  assign y17843 = ~n32036 ;
  assign y17844 = ~n32040 ;
  assign y17845 = n32041 ;
  assign y17846 = n32042 ;
  assign y17847 = ~1'b0 ;
  assign y17848 = 1'b0 ;
  assign y17849 = n32043 ;
  assign y17850 = ~n32045 ;
  assign y17851 = n32050 ;
  assign y17852 = ~1'b0 ;
  assign y17853 = n1434 ;
  assign y17854 = ~n32054 ;
  assign y17855 = ~1'b0 ;
  assign y17856 = ~n32057 ;
  assign y17857 = ~1'b0 ;
  assign y17858 = n32061 ;
  assign y17859 = ~n32063 ;
  assign y17860 = n32064 ;
  assign y17861 = ~n32065 ;
  assign y17862 = ~n32067 ;
  assign y17863 = ~n32068 ;
  assign y17864 = 1'b0 ;
  assign y17865 = ~n32073 ;
  assign y17866 = 1'b0 ;
  assign y17867 = ~n30121 ;
  assign y17868 = ~1'b0 ;
  assign y17869 = ~n32076 ;
  assign y17870 = ~n32077 ;
  assign y17871 = n32083 ;
  assign y17872 = n32089 ;
  assign y17873 = ~n9755 ;
  assign y17874 = n31953 ;
  assign y17875 = n32091 ;
  assign y17876 = ~n32093 ;
  assign y17877 = 1'b0 ;
  assign y17878 = n14226 ;
  assign y17879 = ~n7297 ;
  assign y17880 = n32095 ;
  assign y17881 = ~1'b0 ;
  assign y17882 = ~1'b0 ;
  assign y17883 = ~1'b0 ;
  assign y17884 = ~n32099 ;
  assign y17885 = n21993 ;
  assign y17886 = ~1'b0 ;
  assign y17887 = n32102 ;
  assign y17888 = n17251 ;
  assign y17889 = ~1'b0 ;
  assign y17890 = 1'b0 ;
  assign y17891 = ~1'b0 ;
  assign y17892 = ~1'b0 ;
  assign y17893 = ~1'b0 ;
  assign y17894 = n32103 ;
  assign y17895 = ~1'b0 ;
  assign y17896 = n32108 ;
  assign y17897 = ~n32109 ;
  assign y17898 = ~1'b0 ;
  assign y17899 = ~n32110 ;
  assign y17900 = n23264 ;
  assign y17901 = ~1'b0 ;
  assign y17902 = ~1'b0 ;
  assign y17903 = 1'b0 ;
  assign y17904 = n32111 ;
  assign y17905 = n32113 ;
  assign y17906 = n32114 ;
  assign y17907 = 1'b0 ;
  assign y17908 = ~n32115 ;
  assign y17909 = ~n32121 ;
  assign y17910 = ~1'b0 ;
  assign y17911 = n32124 ;
  assign y17912 = ~n32128 ;
  assign y17913 = n32131 ;
  assign y17914 = n32134 ;
  assign y17915 = n32136 ;
  assign y17916 = 1'b0 ;
  assign y17917 = n32139 ;
  assign y17918 = n32141 ;
  assign y17919 = ~n32142 ;
  assign y17920 = ~1'b0 ;
  assign y17921 = ~n32143 ;
  assign y17922 = n32144 ;
  assign y17923 = n26743 ;
  assign y17924 = ~n32146 ;
  assign y17925 = n32148 ;
  assign y17926 = n32149 ;
  assign y17927 = n32150 ;
  assign y17928 = ~n32152 ;
  assign y17929 = n32153 ;
  assign y17930 = n32154 ;
  assign y17931 = ~1'b0 ;
  assign y17932 = ~1'b0 ;
  assign y17933 = ~n13013 ;
  assign y17934 = ~1'b0 ;
  assign y17935 = n32155 ;
  assign y17936 = ~1'b0 ;
  assign y17937 = ~n32156 ;
  assign y17938 = ~1'b0 ;
  assign y17939 = ~1'b0 ;
  assign y17940 = n5336 ;
  assign y17941 = ~n32158 ;
  assign y17942 = ~n32160 ;
  assign y17943 = ~n32161 ;
  assign y17944 = ~n32162 ;
  assign y17945 = ~n32170 ;
  assign y17946 = n32175 ;
  assign y17947 = 1'b0 ;
  assign y17948 = ~n32177 ;
  assign y17949 = n32178 ;
  assign y17950 = n32181 ;
  assign y17951 = ~1'b0 ;
  assign y17952 = ~1'b0 ;
  assign y17953 = ~1'b0 ;
  assign y17954 = ~1'b0 ;
  assign y17955 = ~n32183 ;
  assign y17956 = ~n32184 ;
  assign y17957 = ~1'b0 ;
  assign y17958 = ~n32186 ;
  assign y17959 = ~n32187 ;
  assign y17960 = n32188 ;
  assign y17961 = n32190 ;
  assign y17962 = ~1'b0 ;
  assign y17963 = ~1'b0 ;
  assign y17964 = ~1'b0 ;
  assign y17965 = ~n231 ;
  assign y17966 = ~1'b0 ;
  assign y17967 = ~n32193 ;
  assign y17968 = n32194 ;
  assign y17969 = n32195 ;
  assign y17970 = ~1'b0 ;
  assign y17971 = ~n15195 ;
  assign y17972 = ~1'b0 ;
  assign y17973 = ~n32200 ;
  assign y17974 = n32204 ;
  assign y17975 = n32207 ;
  assign y17976 = n32214 ;
  assign y17977 = ~1'b0 ;
  assign y17978 = ~n32224 ;
  assign y17979 = ~1'b0 ;
  assign y17980 = ~n32231 ;
  assign y17981 = ~1'b0 ;
  assign y17982 = ~1'b0 ;
  assign y17983 = n32233 ;
  assign y17984 = ~n32242 ;
  assign y17985 = ~n32243 ;
  assign y17986 = ~n32244 ;
  assign y17987 = n32245 ;
  assign y17988 = ~n32248 ;
  assign y17989 = ~1'b0 ;
  assign y17990 = ~1'b0 ;
  assign y17991 = n32249 ;
  assign y17992 = ~n32254 ;
  assign y17993 = ~1'b0 ;
  assign y17994 = ~n32257 ;
  assign y17995 = ~1'b0 ;
  assign y17996 = ~1'b0 ;
  assign y17997 = n32261 ;
  assign y17998 = n32266 ;
  assign y17999 = ~n32269 ;
  assign y18000 = ~1'b0 ;
  assign y18001 = n32270 ;
  assign y18002 = ~1'b0 ;
  assign y18003 = n32274 ;
  assign y18004 = ~1'b0 ;
  assign y18005 = ~n32279 ;
  assign y18006 = ~n32281 ;
  assign y18007 = ~n32283 ;
  assign y18008 = ~n32287 ;
  assign y18009 = ~n32288 ;
  assign y18010 = n32290 ;
  assign y18011 = ~1'b0 ;
  assign y18012 = ~1'b0 ;
  assign y18013 = ~n32292 ;
  assign y18014 = ~1'b0 ;
  assign y18015 = ~n32296 ;
  assign y18016 = ~n32297 ;
  assign y18017 = ~n32299 ;
  assign y18018 = ~1'b0 ;
  assign y18019 = ~n32301 ;
  assign y18020 = ~n32302 ;
  assign y18021 = n32305 ;
  assign y18022 = ~n32306 ;
  assign y18023 = ~1'b0 ;
  assign y18024 = n32307 ;
  assign y18025 = 1'b0 ;
  assign y18026 = ~n32312 ;
  assign y18027 = n32315 ;
  assign y18028 = ~1'b0 ;
  assign y18029 = n3325 ;
  assign y18030 = ~1'b0 ;
  assign y18031 = ~n49 ;
  assign y18032 = ~1'b0 ;
  assign y18033 = ~1'b0 ;
  assign y18034 = ~n32316 ;
  assign y18035 = ~1'b0 ;
  assign y18036 = n32318 ;
  assign y18037 = n6865 ;
  assign y18038 = 1'b0 ;
  assign y18039 = n24621 ;
  assign y18040 = ~n32320 ;
  assign y18041 = n32325 ;
  assign y18042 = n32327 ;
  assign y18043 = ~1'b0 ;
  assign y18044 = ~1'b0 ;
  assign y18045 = n32328 ;
  assign y18046 = ~1'b0 ;
  assign y18047 = n32336 ;
  assign y18048 = ~1'b0 ;
  assign y18049 = n32339 ;
  assign y18050 = ~n32340 ;
  assign y18051 = ~n32342 ;
  assign y18052 = n32343 ;
  assign y18053 = ~n32347 ;
  assign y18054 = ~1'b0 ;
  assign y18055 = ~n32348 ;
  assign y18056 = ~n32350 ;
  assign y18057 = n24023 ;
  assign y18058 = n24007 ;
  assign y18059 = n32354 ;
  assign y18060 = n32355 ;
  assign y18061 = n32361 ;
  assign y18062 = ~n6941 ;
  assign y18063 = ~n32365 ;
  assign y18064 = ~1'b0 ;
  assign y18065 = ~1'b0 ;
  assign y18066 = 1'b0 ;
  assign y18067 = ~1'b0 ;
  assign y18068 = n32370 ;
  assign y18069 = ~1'b0 ;
  assign y18070 = n32371 ;
  assign y18071 = n32373 ;
  assign y18072 = n32377 ;
  assign y18073 = n32378 ;
  assign y18074 = n32385 ;
  assign y18075 = n32386 ;
  assign y18076 = n32387 ;
  assign y18077 = n32388 ;
  assign y18078 = n22454 ;
  assign y18079 = n32390 ;
  assign y18080 = ~1'b0 ;
  assign y18081 = n16909 ;
  assign y18082 = ~1'b0 ;
  assign y18083 = ~n32391 ;
  assign y18084 = n32392 ;
  assign y18085 = n32394 ;
  assign y18086 = n32396 ;
  assign y18087 = ~1'b0 ;
  assign y18088 = ~1'b0 ;
  assign y18089 = n32397 ;
  assign y18090 = ~1'b0 ;
  assign y18091 = ~n32398 ;
  assign y18092 = ~1'b0 ;
  assign y18093 = n32399 ;
  assign y18094 = ~n32400 ;
  assign y18095 = ~1'b0 ;
  assign y18096 = ~1'b0 ;
  assign y18097 = ~n16947 ;
  assign y18098 = ~1'b0 ;
  assign y18099 = ~n32401 ;
  assign y18100 = n32404 ;
  assign y18101 = ~n32406 ;
  assign y18102 = ~1'b0 ;
  assign y18103 = n32407 ;
  assign y18104 = ~n32408 ;
  assign y18105 = ~n1325 ;
  assign y18106 = ~1'b0 ;
  assign y18107 = ~1'b0 ;
  assign y18108 = ~n32409 ;
  assign y18109 = ~n32413 ;
  assign y18110 = n32415 ;
  assign y18111 = n32417 ;
  assign y18112 = n32420 ;
  assign y18113 = n32421 ;
  assign y18114 = ~1'b0 ;
  assign y18115 = n32423 ;
  assign y18116 = ~n27432 ;
  assign y18117 = ~n32426 ;
  assign y18118 = ~n32427 ;
  assign y18119 = ~1'b0 ;
  assign y18120 = n25449 ;
  assign y18121 = ~n32430 ;
  assign y18122 = ~1'b0 ;
  assign y18123 = n32431 ;
  assign y18124 = ~n32432 ;
  assign y18125 = ~1'b0 ;
  assign y18126 = ~1'b0 ;
  assign y18127 = ~n32447 ;
  assign y18128 = n32448 ;
  assign y18129 = n32452 ;
  assign y18130 = ~1'b0 ;
  assign y18131 = n32453 ;
  assign y18132 = n32456 ;
  assign y18133 = n32460 ;
  assign y18134 = n32461 ;
  assign y18135 = ~n12669 ;
  assign y18136 = ~1'b0 ;
  assign y18137 = ~n32463 ;
  assign y18138 = ~1'b0 ;
  assign y18139 = n32464 ;
  assign y18140 = n32468 ;
  assign y18141 = n5082 ;
  assign y18142 = n32471 ;
  assign y18143 = n32472 ;
  assign y18144 = n32475 ;
  assign y18145 = ~1'b0 ;
  assign y18146 = ~n29587 ;
  assign y18147 = ~1'b0 ;
  assign y18148 = ~n32477 ;
  assign y18149 = n32481 ;
  assign y18150 = ~n32482 ;
  assign y18151 = ~n5136 ;
  assign y18152 = n32483 ;
  assign y18153 = 1'b0 ;
  assign y18154 = n32485 ;
  assign y18155 = ~n32486 ;
  assign y18156 = ~n32489 ;
  assign y18157 = ~1'b0 ;
  assign y18158 = ~1'b0 ;
  assign y18159 = ~n32490 ;
  assign y18160 = ~n32492 ;
  assign y18161 = n32494 ;
  assign y18162 = n32499 ;
  assign y18163 = ~n32506 ;
  assign y18164 = ~n32507 ;
  assign y18165 = n32508 ;
  assign y18166 = n8620 ;
  assign y18167 = 1'b0 ;
  assign y18168 = n32518 ;
  assign y18169 = ~n32519 ;
  assign y18170 = n32522 ;
  assign y18171 = ~n32524 ;
  assign y18172 = n32526 ;
  assign y18173 = ~1'b0 ;
  assign y18174 = ~n32527 ;
  assign y18175 = ~n32528 ;
  assign y18176 = ~n32531 ;
  assign y18177 = n32532 ;
  assign y18178 = ~n32533 ;
  assign y18179 = ~n32534 ;
  assign y18180 = n32535 ;
  assign y18181 = n32544 ;
  assign y18182 = n32546 ;
  assign y18183 = ~n32553 ;
  assign y18184 = ~1'b0 ;
  assign y18185 = ~n32554 ;
  assign y18186 = ~1'b0 ;
  assign y18187 = n13708 ;
  assign y18188 = n32557 ;
  assign y18189 = ~n32559 ;
  assign y18190 = n32561 ;
  assign y18191 = ~n32562 ;
  assign y18192 = n32564 ;
  assign y18193 = ~n32565 ;
  assign y18194 = n32570 ;
  assign y18195 = n32572 ;
  assign y18196 = ~1'b0 ;
  assign y18197 = n32575 ;
  assign y18198 = n32576 ;
  assign y18199 = ~1'b0 ;
  assign y18200 = n32579 ;
  assign y18201 = ~n32580 ;
  assign y18202 = n32581 ;
  assign y18203 = ~1'b0 ;
  assign y18204 = ~1'b0 ;
  assign y18205 = ~1'b0 ;
  assign y18206 = n5137 ;
  assign y18207 = ~1'b0 ;
  assign y18208 = ~n32584 ;
  assign y18209 = ~1'b0 ;
  assign y18210 = ~n32591 ;
  assign y18211 = ~n32595 ;
  assign y18212 = ~1'b0 ;
  assign y18213 = ~n32598 ;
  assign y18214 = ~n32601 ;
  assign y18215 = ~n32602 ;
  assign y18216 = ~1'b0 ;
  assign y18217 = ~n32606 ;
  assign y18218 = ~1'b0 ;
  assign y18219 = n32607 ;
  assign y18220 = n32608 ;
  assign y18221 = n32612 ;
  assign y18222 = ~1'b0 ;
  assign y18223 = n32613 ;
  assign y18224 = n32615 ;
  assign y18225 = ~n32616 ;
  assign y18226 = ~1'b0 ;
  assign y18227 = n32620 ;
  assign y18228 = ~1'b0 ;
  assign y18229 = ~1'b0 ;
  assign y18230 = ~n32621 ;
  assign y18231 = n32622 ;
  assign y18232 = n32625 ;
  assign y18233 = ~1'b0 ;
  assign y18234 = ~1'b0 ;
  assign y18235 = n32630 ;
  assign y18236 = n32632 ;
  assign y18237 = ~1'b0 ;
  assign y18238 = n32634 ;
  assign y18239 = ~n32636 ;
  assign y18240 = ~n32638 ;
  assign y18241 = ~n32640 ;
  assign y18242 = ~1'b0 ;
  assign y18243 = n3061 ;
  assign y18244 = n32643 ;
  assign y18245 = ~1'b0 ;
  assign y18246 = ~1'b0 ;
  assign y18247 = ~1'b0 ;
  assign y18248 = n32644 ;
  assign y18249 = n32645 ;
  assign y18250 = ~n32646 ;
  assign y18251 = ~1'b0 ;
  assign y18252 = n32650 ;
  assign y18253 = ~1'b0 ;
  assign y18254 = n32653 ;
  assign y18255 = n22636 ;
  assign y18256 = n32654 ;
  assign y18257 = ~n32657 ;
  assign y18258 = ~n32661 ;
  assign y18259 = ~1'b0 ;
  assign y18260 = ~1'b0 ;
  assign y18261 = 1'b0 ;
  assign y18262 = ~1'b0 ;
  assign y18263 = n32662 ;
  assign y18264 = n32666 ;
  assign y18265 = n32670 ;
  assign y18266 = n32674 ;
  assign y18267 = ~n32676 ;
  assign y18268 = n32679 ;
  assign y18269 = ~1'b0 ;
  assign y18270 = 1'b0 ;
  assign y18271 = ~1'b0 ;
  assign y18272 = n32689 ;
  assign y18273 = ~1'b0 ;
  assign y18274 = ~n32690 ;
  assign y18275 = n15535 ;
  assign y18276 = ~1'b0 ;
  assign y18277 = ~n32692 ;
  assign y18278 = 1'b0 ;
  assign y18279 = n32695 ;
  assign y18280 = n32696 ;
  assign y18281 = n17962 ;
  assign y18282 = ~n6036 ;
  assign y18283 = ~1'b0 ;
  assign y18284 = ~1'b0 ;
  assign y18285 = ~n32698 ;
  assign y18286 = n32700 ;
  assign y18287 = n32701 ;
  assign y18288 = ~n32702 ;
  assign y18289 = n32705 ;
  assign y18290 = ~n32710 ;
  assign y18291 = n32711 ;
  assign y18292 = ~1'b0 ;
  assign y18293 = ~n32713 ;
  assign y18294 = ~1'b0 ;
  assign y18295 = ~1'b0 ;
  assign y18296 = ~1'b0 ;
  assign y18297 = ~n32714 ;
  assign y18298 = ~1'b0 ;
  assign y18299 = ~1'b0 ;
  assign y18300 = ~1'b0 ;
  assign y18301 = ~n32715 ;
  assign y18302 = n32719 ;
  assign y18303 = ~n32721 ;
  assign y18304 = ~1'b0 ;
  assign y18305 = ~1'b0 ;
  assign y18306 = ~1'b0 ;
  assign y18307 = ~n32725 ;
  assign y18308 = ~n32728 ;
  assign y18309 = n32734 ;
  assign y18310 = ~n32736 ;
  assign y18311 = ~n32737 ;
  assign y18312 = n32738 ;
  assign y18313 = n32740 ;
  assign y18314 = ~1'b0 ;
  assign y18315 = ~1'b0 ;
  assign y18316 = n32742 ;
  assign y18317 = ~1'b0 ;
  assign y18318 = ~n32745 ;
  assign y18319 = n12813 ;
  assign y18320 = ~n32746 ;
  assign y18321 = ~1'b0 ;
  assign y18322 = ~1'b0 ;
  assign y18323 = ~n32749 ;
  assign y18324 = ~n32751 ;
  assign y18325 = n32754 ;
  assign y18326 = ~1'b0 ;
  assign y18327 = ~n32757 ;
  assign y18328 = ~n32758 ;
  assign y18329 = n32760 ;
  assign y18330 = n23355 ;
  assign y18331 = 1'b0 ;
  assign y18332 = n17861 ;
  assign y18333 = ~n32763 ;
  assign y18334 = n19931 ;
  assign y18335 = ~n32764 ;
  assign y18336 = ~1'b0 ;
  assign y18337 = ~n32766 ;
  assign y18338 = ~1'b0 ;
  assign y18339 = n32767 ;
  assign y18340 = ~1'b0 ;
  assign y18341 = ~n32772 ;
  assign y18342 = n32773 ;
  assign y18343 = n32778 ;
  assign y18344 = ~n32779 ;
  assign y18345 = ~1'b0 ;
  assign y18346 = n32785 ;
  assign y18347 = ~n32786 ;
  assign y18348 = ~1'b0 ;
  assign y18349 = n32788 ;
  assign y18350 = n32790 ;
  assign y18351 = ~1'b0 ;
  assign y18352 = n32791 ;
  assign y18353 = n32792 ;
  assign y18354 = n32795 ;
  assign y18355 = n32796 ;
  assign y18356 = n32803 ;
  assign y18357 = ~n32809 ;
  assign y18358 = ~1'b0 ;
  assign y18359 = ~1'b0 ;
  assign y18360 = ~n32817 ;
  assign y18361 = ~n32819 ;
  assign y18362 = ~n32822 ;
  assign y18363 = ~1'b0 ;
  assign y18364 = ~1'b0 ;
  assign y18365 = ~1'b0 ;
  assign y18366 = n32823 ;
  assign y18367 = 1'b0 ;
  assign y18368 = ~n32825 ;
  assign y18369 = ~1'b0 ;
  assign y18370 = n32826 ;
  assign y18371 = ~1'b0 ;
  assign y18372 = ~1'b0 ;
  assign y18373 = ~n32827 ;
  assign y18374 = ~n32828 ;
  assign y18375 = n32832 ;
  assign y18376 = ~n32833 ;
  assign y18377 = ~1'b0 ;
  assign y18378 = ~1'b0 ;
  assign y18379 = ~1'b0 ;
  assign y18380 = n32835 ;
  assign y18381 = 1'b0 ;
  assign y18382 = ~n32838 ;
  assign y18383 = n32842 ;
  assign y18384 = n32844 ;
  assign y18385 = ~n32845 ;
  assign y18386 = n32846 ;
  assign y18387 = ~1'b0 ;
  assign y18388 = ~n32854 ;
  assign y18389 = ~1'b0 ;
  assign y18390 = ~n32858 ;
  assign y18391 = ~n32861 ;
  assign y18392 = ~n32863 ;
  assign y18393 = ~n32866 ;
  assign y18394 = ~n32869 ;
  assign y18395 = ~n32871 ;
  assign y18396 = n32875 ;
  assign y18397 = n32882 ;
  assign y18398 = ~1'b0 ;
  assign y18399 = n32884 ;
  assign y18400 = n32885 ;
  assign y18401 = n32888 ;
  assign y18402 = ~n32895 ;
  assign y18403 = ~n9865 ;
  assign y18404 = n32896 ;
  assign y18405 = ~1'b0 ;
  assign y18406 = ~1'b0 ;
  assign y18407 = ~n32905 ;
  assign y18408 = ~1'b0 ;
  assign y18409 = ~n8624 ;
  assign y18410 = ~1'b0 ;
  assign y18411 = n32909 ;
  assign y18412 = ~n32910 ;
  assign y18413 = ~1'b0 ;
  assign y18414 = n32911 ;
  assign y18415 = ~1'b0 ;
  assign y18416 = ~n32914 ;
  assign y18417 = n32916 ;
  assign y18418 = ~n6930 ;
  assign y18419 = ~1'b0 ;
  assign y18420 = n32918 ;
  assign y18421 = n32923 ;
  assign y18422 = ~n32927 ;
  assign y18423 = ~n24568 ;
  assign y18424 = ~1'b0 ;
  assign y18425 = n32928 ;
  assign y18426 = ~n32929 ;
  assign y18427 = ~n32930 ;
  assign y18428 = ~1'b0 ;
  assign y18429 = ~1'b0 ;
  assign y18430 = ~n32932 ;
  assign y18431 = ~1'b0 ;
  assign y18432 = ~n32937 ;
  assign y18433 = n32938 ;
  assign y18434 = ~n32943 ;
  assign y18435 = n32947 ;
  assign y18436 = n32949 ;
  assign y18437 = ~1'b0 ;
  assign y18438 = ~1'b0 ;
  assign y18439 = ~n32950 ;
  assign y18440 = n32952 ;
  assign y18441 = ~1'b0 ;
  assign y18442 = ~n32956 ;
  assign y18443 = n32962 ;
  assign y18444 = 1'b0 ;
  assign y18445 = ~1'b0 ;
  assign y18446 = ~1'b0 ;
  assign y18447 = ~n32963 ;
  assign y18448 = ~1'b0 ;
  assign y18449 = n32965 ;
  assign y18450 = n32967 ;
  assign y18451 = 1'b0 ;
  assign y18452 = n32973 ;
  assign y18453 = ~1'b0 ;
  assign y18454 = n32976 ;
  assign y18455 = ~n32977 ;
  assign y18456 = n32978 ;
  assign y18457 = ~n32980 ;
  assign y18458 = n32981 ;
  assign y18459 = ~n32982 ;
  assign y18460 = ~1'b0 ;
  assign y18461 = n3039 ;
  assign y18462 = ~1'b0 ;
  assign y18463 = 1'b0 ;
  assign y18464 = ~n32986 ;
  assign y18465 = ~1'b0 ;
  assign y18466 = ~n32987 ;
  assign y18467 = n32993 ;
  assign y18468 = n32997 ;
  assign y18469 = ~1'b0 ;
  assign y18470 = n33005 ;
  assign y18471 = ~1'b0 ;
  assign y18472 = ~n33007 ;
  assign y18473 = 1'b0 ;
  assign y18474 = ~1'b0 ;
  assign y18475 = ~1'b0 ;
  assign y18476 = ~n33011 ;
  assign y18477 = n33012 ;
  assign y18478 = n33013 ;
  assign y18479 = ~1'b0 ;
  assign y18480 = ~n33015 ;
  assign y18481 = n33018 ;
  assign y18482 = ~1'b0 ;
  assign y18483 = n33021 ;
  assign y18484 = ~n33023 ;
  assign y18485 = ~n33026 ;
  assign y18486 = n33027 ;
  assign y18487 = ~n33028 ;
  assign y18488 = n33032 ;
  assign y18489 = n33036 ;
  assign y18490 = ~n33038 ;
  assign y18491 = n33039 ;
  assign y18492 = n33040 ;
  assign y18493 = ~1'b0 ;
  assign y18494 = ~1'b0 ;
  assign y18495 = n33043 ;
  assign y18496 = ~n33046 ;
  assign y18497 = n33047 ;
  assign y18498 = ~n16841 ;
  assign y18499 = ~n33048 ;
  assign y18500 = n33049 ;
  assign y18501 = ~n33054 ;
  assign y18502 = ~1'b0 ;
  assign y18503 = ~1'b0 ;
  assign y18504 = n845 ;
  assign y18505 = n33058 ;
  assign y18506 = n33059 ;
  assign y18507 = ~n13981 ;
  assign y18508 = ~n33060 ;
  assign y18509 = ~n33061 ;
  assign y18510 = n33064 ;
  assign y18511 = n33067 ;
  assign y18512 = ~1'b0 ;
  assign y18513 = n33069 ;
  assign y18514 = ~n33072 ;
  assign y18515 = n33079 ;
  assign y18516 = ~n33083 ;
  assign y18517 = 1'b0 ;
  assign y18518 = ~1'b0 ;
  assign y18519 = ~n33089 ;
  assign y18520 = ~n30708 ;
  assign y18521 = ~1'b0 ;
  assign y18522 = n33090 ;
  assign y18523 = ~1'b0 ;
  assign y18524 = ~n33096 ;
  assign y18525 = ~1'b0 ;
  assign y18526 = ~1'b0 ;
  assign y18527 = n33097 ;
  assign y18528 = ~n33104 ;
  assign y18529 = ~1'b0 ;
  assign y18530 = n33107 ;
  assign y18531 = ~1'b0 ;
  assign y18532 = n33111 ;
  assign y18533 = n33117 ;
  assign y18534 = ~1'b0 ;
  assign y18535 = ~1'b0 ;
  assign y18536 = ~1'b0 ;
  assign y18537 = n33118 ;
  assign y18538 = 1'b0 ;
  assign y18539 = ~1'b0 ;
  assign y18540 = ~n33123 ;
  assign y18541 = ~1'b0 ;
  assign y18542 = ~1'b0 ;
  assign y18543 = ~n8751 ;
  assign y18544 = ~n33126 ;
  assign y18545 = ~1'b0 ;
  assign y18546 = ~n33133 ;
  assign y18547 = ~1'b0 ;
  assign y18548 = ~n5566 ;
  assign y18549 = ~n33136 ;
  assign y18550 = n33137 ;
  assign y18551 = ~n33138 ;
  assign y18552 = 1'b0 ;
  assign y18553 = n33141 ;
  assign y18554 = ~n33144 ;
  assign y18555 = n33146 ;
  assign y18556 = ~n33147 ;
  assign y18557 = n33148 ;
  assign y18558 = n33150 ;
  assign y18559 = ~n33155 ;
  assign y18560 = ~n33156 ;
  assign y18561 = n33158 ;
  assign y18562 = ~1'b0 ;
  assign y18563 = ~1'b0 ;
  assign y18564 = n33159 ;
  assign y18565 = n33161 ;
  assign y18566 = ~1'b0 ;
  assign y18567 = ~n33163 ;
  assign y18568 = ~n22756 ;
  assign y18569 = ~n33165 ;
  assign y18570 = n33172 ;
  assign y18571 = ~1'b0 ;
  assign y18572 = n33174 ;
  assign y18573 = n1020 ;
  assign y18574 = ~1'b0 ;
  assign y18575 = ~1'b0 ;
  assign y18576 = ~1'b0 ;
  assign y18577 = ~n33175 ;
  assign y18578 = n33176 ;
  assign y18579 = ~n33177 ;
  assign y18580 = ~1'b0 ;
  assign y18581 = ~n33179 ;
  assign y18582 = ~1'b0 ;
  assign y18583 = ~1'b0 ;
  assign y18584 = n33181 ;
  assign y18585 = ~n33185 ;
  assign y18586 = n33186 ;
  assign y18587 = ~n33193 ;
  assign y18588 = ~n33195 ;
  assign y18589 = ~n33198 ;
  assign y18590 = ~n33200 ;
  assign y18591 = ~1'b0 ;
  assign y18592 = n33201 ;
  assign y18593 = 1'b0 ;
  assign y18594 = ~n33207 ;
  assign y18595 = ~n33209 ;
  assign y18596 = ~n33210 ;
  assign y18597 = n33215 ;
  assign y18598 = ~n33216 ;
  assign y18599 = n33218 ;
  assign y18600 = ~1'b0 ;
  assign y18601 = ~1'b0 ;
  assign y18602 = ~n26104 ;
  assign y18603 = n33223 ;
  assign y18604 = ~n33225 ;
  assign y18605 = ~1'b0 ;
  assign y18606 = n33227 ;
  assign y18607 = ~n33228 ;
  assign y18608 = ~n18522 ;
  assign y18609 = ~n33229 ;
  assign y18610 = n33231 ;
  assign y18611 = ~1'b0 ;
  assign y18612 = ~n33233 ;
  assign y18613 = n33236 ;
  assign y18614 = ~1'b0 ;
  assign y18615 = n33237 ;
  assign y18616 = ~1'b0 ;
  assign y18617 = n33238 ;
  assign y18618 = 1'b0 ;
  assign y18619 = ~n33241 ;
  assign y18620 = ~n33242 ;
  assign y18621 = n33244 ;
  assign y18622 = ~1'b0 ;
  assign y18623 = ~n33246 ;
  assign y18624 = ~1'b0 ;
  assign y18625 = ~n33248 ;
  assign y18626 = ~n33250 ;
  assign y18627 = ~n33251 ;
  assign y18628 = n33253 ;
  assign y18629 = ~1'b0 ;
  assign y18630 = ~n33255 ;
  assign y18631 = ~n33259 ;
  assign y18632 = ~n33260 ;
  assign y18633 = ~n33261 ;
  assign y18634 = ~n33263 ;
  assign y18635 = ~n33264 ;
  assign y18636 = n33268 ;
  assign y18637 = n33272 ;
  assign y18638 = ~1'b0 ;
  assign y18639 = ~1'b0 ;
  assign y18640 = ~n33273 ;
  assign y18641 = ~1'b0 ;
  assign y18642 = n33279 ;
  assign y18643 = ~1'b0 ;
  assign y18644 = n33286 ;
  assign y18645 = ~n33291 ;
  assign y18646 = ~1'b0 ;
  assign y18647 = n33294 ;
  assign y18648 = ~1'b0 ;
  assign y18649 = n33295 ;
  assign y18650 = ~n33297 ;
  assign y18651 = ~1'b0 ;
  assign y18652 = n33300 ;
  assign y18653 = ~n33307 ;
  assign y18654 = ~1'b0 ;
  assign y18655 = ~1'b0 ;
  assign y18656 = ~n33308 ;
  assign y18657 = n33309 ;
  assign y18658 = n14841 ;
  assign y18659 = n33312 ;
  assign y18660 = ~n33313 ;
  assign y18661 = ~n33315 ;
  assign y18662 = n33318 ;
  assign y18663 = ~1'b0 ;
  assign y18664 = n33320 ;
  assign y18665 = n33321 ;
  assign y18666 = ~n33324 ;
  assign y18667 = n33326 ;
  assign y18668 = ~n33327 ;
  assign y18669 = ~n33328 ;
  assign y18670 = ~1'b0 ;
  assign y18671 = ~1'b0 ;
  assign y18672 = ~n19771 ;
  assign y18673 = ~1'b0 ;
  assign y18674 = ~1'b0 ;
  assign y18675 = n33331 ;
  assign y18676 = n33333 ;
  assign y18677 = n33335 ;
  assign y18678 = n33337 ;
  assign y18679 = ~n33339 ;
  assign y18680 = ~1'b0 ;
  assign y18681 = ~n33340 ;
  assign y18682 = ~n33343 ;
  assign y18683 = ~n2192 ;
  assign y18684 = n33345 ;
  assign y18685 = ~1'b0 ;
  assign y18686 = n33347 ;
  assign y18687 = ~n33348 ;
  assign y18688 = ~n33349 ;
  assign y18689 = n33355 ;
  assign y18690 = n23944 ;
  assign y18691 = ~n33356 ;
  assign y18692 = ~1'b0 ;
  assign y18693 = ~1'b0 ;
  assign y18694 = ~1'b0 ;
  assign y18695 = ~n33359 ;
  assign y18696 = n33361 ;
  assign y18697 = ~n33368 ;
  assign y18698 = ~n33370 ;
  assign y18699 = ~1'b0 ;
  assign y18700 = n33371 ;
  assign y18701 = n33372 ;
  assign y18702 = ~1'b0 ;
  assign y18703 = n33375 ;
  assign y18704 = ~1'b0 ;
  assign y18705 = n33377 ;
  assign y18706 = ~1'b0 ;
  assign y18707 = ~1'b0 ;
  assign y18708 = n33378 ;
  assign y18709 = n2631 ;
  assign y18710 = ~n33380 ;
  assign y18711 = ~1'b0 ;
  assign y18712 = ~1'b0 ;
  assign y18713 = ~n33381 ;
  assign y18714 = ~n33383 ;
  assign y18715 = n33384 ;
  assign y18716 = n33386 ;
  assign y18717 = n33387 ;
  assign y18718 = ~n33391 ;
  assign y18719 = ~n33392 ;
  assign y18720 = ~1'b0 ;
  assign y18721 = 1'b0 ;
  assign y18722 = ~n33395 ;
  assign y18723 = ~1'b0 ;
  assign y18724 = ~1'b0 ;
  assign y18725 = n33402 ;
  assign y18726 = n33405 ;
  assign y18727 = n33407 ;
  assign y18728 = ~n33410 ;
  assign y18729 = n33411 ;
  assign y18730 = n33412 ;
  assign y18731 = ~n33416 ;
  assign y18732 = ~1'b0 ;
  assign y18733 = n33417 ;
  assign y18734 = ~1'b0 ;
  assign y18735 = n5321 ;
  assign y18736 = n33419 ;
  assign y18737 = ~n33421 ;
  assign y18738 = ~1'b0 ;
  assign y18739 = ~1'b0 ;
  assign y18740 = ~n33422 ;
  assign y18741 = ~n33424 ;
  assign y18742 = n33431 ;
  assign y18743 = ~n33432 ;
  assign y18744 = ~1'b0 ;
  assign y18745 = n33435 ;
  assign y18746 = ~1'b0 ;
  assign y18747 = ~n33436 ;
  assign y18748 = ~n33438 ;
  assign y18749 = n33439 ;
  assign y18750 = n33441 ;
  assign y18751 = ~n33444 ;
  assign y18752 = ~n32104 ;
  assign y18753 = ~n33447 ;
  assign y18754 = 1'b0 ;
  assign y18755 = ~1'b0 ;
  assign y18756 = ~n33449 ;
  assign y18757 = n33450 ;
  assign y18758 = ~n33452 ;
  assign y18759 = ~n33454 ;
  assign y18760 = ~n33455 ;
  assign y18761 = ~1'b0 ;
  assign y18762 = ~1'b0 ;
  assign y18763 = 1'b0 ;
  assign y18764 = ~1'b0 ;
  assign y18765 = ~n33462 ;
  assign y18766 = ~1'b0 ;
  assign y18767 = ~n33463 ;
  assign y18768 = n33464 ;
  assign y18769 = n33465 ;
  assign y18770 = ~n8591 ;
  assign y18771 = ~n33467 ;
  assign y18772 = n33469 ;
  assign y18773 = n33471 ;
  assign y18774 = n33475 ;
  assign y18775 = ~n33476 ;
  assign y18776 = n33478 ;
  assign y18777 = n33479 ;
  assign y18778 = ~1'b0 ;
  assign y18779 = ~n33482 ;
  assign y18780 = ~1'b0 ;
  assign y18781 = n28706 ;
  assign y18782 = n33483 ;
  assign y18783 = ~n33488 ;
  assign y18784 = ~1'b0 ;
  assign y18785 = 1'b0 ;
  assign y18786 = 1'b0 ;
  assign y18787 = n33493 ;
  assign y18788 = n33494 ;
  assign y18789 = n33496 ;
  assign y18790 = ~n975 ;
  assign y18791 = ~1'b0 ;
  assign y18792 = ~n33497 ;
  assign y18793 = ~n33504 ;
  assign y18794 = ~1'b0 ;
  assign y18795 = ~1'b0 ;
  assign y18796 = ~n33509 ;
  assign y18797 = n33511 ;
  assign y18798 = ~1'b0 ;
  assign y18799 = n33512 ;
  assign y18800 = n33514 ;
  assign y18801 = n33516 ;
  assign y18802 = ~n33517 ;
  assign y18803 = ~n33518 ;
  assign y18804 = ~n33520 ;
  assign y18805 = ~1'b0 ;
  assign y18806 = ~n33492 ;
  assign y18807 = ~1'b0 ;
  assign y18808 = n33341 ;
  assign y18809 = n33522 ;
  assign y18810 = n33523 ;
  assign y18811 = 1'b0 ;
  assign y18812 = ~1'b0 ;
  assign y18813 = ~n33528 ;
  assign y18814 = ~1'b0 ;
  assign y18815 = ~n33530 ;
  assign y18816 = ~1'b0 ;
  assign y18817 = ~n33531 ;
  assign y18818 = n33533 ;
  assign y18819 = n33534 ;
  assign y18820 = n33535 ;
  assign y18821 = ~n33537 ;
  assign y18822 = n33539 ;
  assign y18823 = ~n8273 ;
  assign y18824 = ~n33540 ;
  assign y18825 = ~n33546 ;
  assign y18826 = ~n33547 ;
  assign y18827 = n33551 ;
  assign y18828 = ~n33553 ;
  assign y18829 = n33556 ;
  assign y18830 = ~1'b0 ;
  assign y18831 = n33558 ;
  assign y18832 = ~n5963 ;
  assign y18833 = ~n33559 ;
  assign y18834 = ~n33563 ;
  assign y18835 = 1'b0 ;
  assign y18836 = ~1'b0 ;
  assign y18837 = ~1'b0 ;
  assign y18838 = ~n33570 ;
  assign y18839 = n33574 ;
  assign y18840 = ~n33575 ;
  assign y18841 = ~1'b0 ;
  assign y18842 = ~n33579 ;
  assign y18843 = ~n33580 ;
  assign y18844 = ~1'b0 ;
  assign y18845 = n33581 ;
  assign y18846 = n33583 ;
  assign y18847 = ~1'b0 ;
  assign y18848 = ~1'b0 ;
  assign y18849 = n33584 ;
  assign y18850 = ~1'b0 ;
  assign y18851 = ~1'b0 ;
  assign y18852 = n33586 ;
  assign y18853 = ~n33591 ;
  assign y18854 = ~n33595 ;
  assign y18855 = n33599 ;
  assign y18856 = n33600 ;
  assign y18857 = ~1'b0 ;
  assign y18858 = ~1'b0 ;
  assign y18859 = ~n33603 ;
  assign y18860 = ~1'b0 ;
  assign y18861 = ~n33604 ;
  assign y18862 = n33605 ;
  assign y18863 = n33606 ;
  assign y18864 = ~n14885 ;
  assign y18865 = ~1'b0 ;
  assign y18866 = n33611 ;
  assign y18867 = ~n33612 ;
  assign y18868 = n33616 ;
  assign y18869 = ~1'b0 ;
  assign y18870 = n33618 ;
  assign y18871 = ~n33619 ;
  assign y18872 = ~n33623 ;
  assign y18873 = n33624 ;
  assign y18874 = ~n33626 ;
  assign y18875 = n33633 ;
  assign y18876 = n33634 ;
  assign y18877 = n33636 ;
  assign y18878 = ~n33637 ;
  assign y18879 = n33639 ;
  assign y18880 = n33643 ;
  assign y18881 = ~n33646 ;
  assign y18882 = ~1'b0 ;
  assign y18883 = ~1'b0 ;
  assign y18884 = 1'b0 ;
  assign y18885 = ~1'b0 ;
  assign y18886 = n33647 ;
  assign y18887 = ~n33648 ;
  assign y18888 = n4939 ;
  assign y18889 = n33649 ;
  assign y18890 = n33651 ;
  assign y18891 = ~1'b0 ;
  assign y18892 = ~n33653 ;
  assign y18893 = ~1'b0 ;
  assign y18894 = n33654 ;
  assign y18895 = ~n33655 ;
  assign y18896 = ~1'b0 ;
  assign y18897 = ~n20547 ;
  assign y18898 = n4341 ;
  assign y18899 = n33657 ;
  assign y18900 = ~1'b0 ;
  assign y18901 = ~n33658 ;
  assign y18902 = ~n33662 ;
  assign y18903 = ~1'b0 ;
  assign y18904 = ~n33666 ;
  assign y18905 = ~1'b0 ;
  assign y18906 = ~1'b0 ;
  assign y18907 = ~1'b0 ;
  assign y18908 = ~1'b0 ;
  assign y18909 = n33673 ;
  assign y18910 = ~n16853 ;
  assign y18911 = ~1'b0 ;
  assign y18912 = ~n33675 ;
  assign y18913 = n33678 ;
  assign y18914 = ~1'b0 ;
  assign y18915 = ~n33681 ;
  assign y18916 = ~n33685 ;
  assign y18917 = ~n33691 ;
  assign y18918 = n33693 ;
  assign y18919 = ~1'b0 ;
  assign y18920 = ~n33696 ;
  assign y18921 = ~n33698 ;
  assign y18922 = n33701 ;
  assign y18923 = n33702 ;
  assign y18924 = ~n33705 ;
  assign y18925 = n33707 ;
  assign y18926 = n33708 ;
  assign y18927 = ~n33711 ;
  assign y18928 = ~n33712 ;
  assign y18929 = ~1'b0 ;
  assign y18930 = ~n33717 ;
  assign y18931 = ~1'b0 ;
  assign y18932 = ~1'b0 ;
  assign y18933 = ~1'b0 ;
  assign y18934 = ~n10089 ;
  assign y18935 = n33719 ;
  assign y18936 = n33720 ;
  assign y18937 = ~n33726 ;
  assign y18938 = ~n33728 ;
  assign y18939 = ~n33730 ;
  assign y18940 = ~n33731 ;
  assign y18941 = ~1'b0 ;
  assign y18942 = ~1'b0 ;
  assign y18943 = ~1'b0 ;
  assign y18944 = ~1'b0 ;
  assign y18945 = ~n33740 ;
  assign y18946 = ~1'b0 ;
  assign y18947 = n33742 ;
  assign y18948 = ~1'b0 ;
  assign y18949 = ~n33744 ;
  assign y18950 = n33745 ;
  assign y18951 = n4004 ;
  assign y18952 = ~1'b0 ;
  assign y18953 = 1'b0 ;
  assign y18954 = ~n33747 ;
  assign y18955 = ~n33751 ;
  assign y18956 = 1'b0 ;
  assign y18957 = n33752 ;
  assign y18958 = n33754 ;
  assign y18959 = n33757 ;
  assign y18960 = n33760 ;
  assign y18961 = n33761 ;
  assign y18962 = n33764 ;
  assign y18963 = ~1'b0 ;
  assign y18964 = ~1'b0 ;
  assign y18965 = ~1'b0 ;
  assign y18966 = ~n33768 ;
  assign y18967 = n33769 ;
  assign y18968 = ~1'b0 ;
  assign y18969 = n33770 ;
  assign y18970 = n33771 ;
  assign y18971 = n17412 ;
  assign y18972 = ~n33774 ;
  assign y18973 = ~1'b0 ;
  assign y18974 = ~n33776 ;
  assign y18975 = ~1'b0 ;
  assign y18976 = ~1'b0 ;
  assign y18977 = ~n33784 ;
  assign y18978 = ~n33786 ;
  assign y18979 = ~n27301 ;
  assign y18980 = n33788 ;
  assign y18981 = ~1'b0 ;
  assign y18982 = n22231 ;
  assign y18983 = ~n33789 ;
  assign y18984 = ~1'b0 ;
  assign y18985 = 1'b0 ;
  assign y18986 = ~n33790 ;
  assign y18987 = n33791 ;
  assign y18988 = ~n33793 ;
  assign y18989 = ~1'b0 ;
  assign y18990 = n33798 ;
  assign y18991 = ~n33799 ;
  assign y18992 = n33801 ;
  assign y18993 = ~n33802 ;
  assign y18994 = ~1'b0 ;
  assign y18995 = n33803 ;
  assign y18996 = ~1'b0 ;
  assign y18997 = n7036 ;
  assign y18998 = ~1'b0 ;
  assign y18999 = ~1'b0 ;
  assign y19000 = ~1'b0 ;
  assign y19001 = ~n33804 ;
  assign y19002 = n33809 ;
  assign y19003 = n33814 ;
  assign y19004 = ~n33816 ;
  assign y19005 = ~1'b0 ;
  assign y19006 = ~1'b0 ;
  assign y19007 = n33822 ;
  assign y19008 = n33823 ;
  assign y19009 = 1'b0 ;
  assign y19010 = n33824 ;
  assign y19011 = ~n33825 ;
  assign y19012 = ~n33826 ;
  assign y19013 = n33827 ;
  assign y19014 = n33831 ;
  assign y19015 = ~n33832 ;
  assign y19016 = ~1'b0 ;
  assign y19017 = n33835 ;
  assign y19018 = ~n10965 ;
  assign y19019 = ~n14916 ;
  assign y19020 = n33838 ;
  assign y19021 = n33839 ;
  assign y19022 = n33840 ;
  assign y19023 = ~n33842 ;
  assign y19024 = n33844 ;
  assign y19025 = ~n33845 ;
  assign y19026 = ~n16291 ;
  assign y19027 = n33847 ;
  assign y19028 = n33848 ;
  assign y19029 = ~1'b0 ;
  assign y19030 = ~n33851 ;
  assign y19031 = n33855 ;
  assign y19032 = ~1'b0 ;
  assign y19033 = n33856 ;
  assign y19034 = n33858 ;
  assign y19035 = n33860 ;
  assign y19036 = ~n33862 ;
  assign y19037 = n33864 ;
  assign y19038 = ~n18126 ;
  assign y19039 = ~n33866 ;
  assign y19040 = ~n33868 ;
  assign y19041 = ~n33869 ;
  assign y19042 = ~1'b0 ;
  assign y19043 = ~n33873 ;
  assign y19044 = n33875 ;
  assign y19045 = n33877 ;
  assign y19046 = ~1'b0 ;
  assign y19047 = n16562 ;
  assign y19048 = ~1'b0 ;
  assign y19049 = ~n33878 ;
  assign y19050 = n33880 ;
  assign y19051 = ~n33882 ;
  assign y19052 = ~1'b0 ;
  assign y19053 = n33883 ;
  assign y19054 = n16221 ;
  assign y19055 = ~1'b0 ;
  assign y19056 = n27899 ;
  assign y19057 = n33887 ;
  assign y19058 = ~1'b0 ;
  assign y19059 = ~n33892 ;
  assign y19060 = n33893 ;
  assign y19061 = ~1'b0 ;
  assign y19062 = ~n33895 ;
  assign y19063 = 1'b0 ;
  assign y19064 = ~1'b0 ;
  assign y19065 = ~1'b0 ;
  assign y19066 = ~n33896 ;
  assign y19067 = ~1'b0 ;
  assign y19068 = n33901 ;
  assign y19069 = ~n33903 ;
  assign y19070 = ~n23078 ;
  assign y19071 = ~n33908 ;
  assign y19072 = n9631 ;
  assign y19073 = ~n33910 ;
  assign y19074 = n452 ;
  assign y19075 = ~1'b0 ;
  assign y19076 = ~1'b0 ;
  assign y19077 = n33912 ;
  assign y19078 = ~1'b0 ;
  assign y19079 = n33914 ;
  assign y19080 = ~n11561 ;
  assign y19081 = ~n24467 ;
  assign y19082 = n33915 ;
  assign y19083 = n33916 ;
  assign y19084 = n13503 ;
  assign y19085 = ~1'b0 ;
  assign y19086 = ~n33919 ;
  assign y19087 = ~1'b0 ;
  assign y19088 = 1'b0 ;
  assign y19089 = ~1'b0 ;
  assign y19090 = n33923 ;
  assign y19091 = n33926 ;
  assign y19092 = ~n33932 ;
  assign y19093 = ~n33934 ;
  assign y19094 = ~n33939 ;
  assign y19095 = n33941 ;
  assign y19096 = ~n33943 ;
  assign y19097 = ~n33946 ;
  assign y19098 = ~1'b0 ;
  assign y19099 = ~1'b0 ;
  assign y19100 = ~n33949 ;
  assign y19101 = ~1'b0 ;
  assign y19102 = n33950 ;
  assign y19103 = ~n33953 ;
  assign y19104 = ~n33956 ;
  assign y19105 = ~n33960 ;
  assign y19106 = n33964 ;
  assign y19107 = ~n33965 ;
  assign y19108 = ~n33966 ;
  assign y19109 = n12843 ;
  assign y19110 = n33969 ;
  assign y19111 = ~1'b0 ;
  assign y19112 = n33973 ;
  assign y19113 = ~1'b0 ;
  assign y19114 = ~1'b0 ;
  assign y19115 = ~n33974 ;
  assign y19116 = ~1'b0 ;
  assign y19117 = ~n33976 ;
  assign y19118 = n33977 ;
  assign y19119 = ~n33979 ;
  assign y19120 = ~1'b0 ;
  assign y19121 = ~n33984 ;
  assign y19122 = ~n33985 ;
  assign y19123 = ~n12239 ;
  assign y19124 = ~n33987 ;
  assign y19125 = ~n33990 ;
  assign y19126 = n33995 ;
  assign y19127 = ~1'b0 ;
  assign y19128 = ~1'b0 ;
  assign y19129 = ~1'b0 ;
  assign y19130 = ~1'b0 ;
  assign y19131 = n33998 ;
  assign y19132 = ~1'b0 ;
  assign y19133 = n33999 ;
  assign y19134 = ~1'b0 ;
  assign y19135 = n34000 ;
  assign y19136 = ~n34003 ;
  assign y19137 = ~n34005 ;
  assign y19138 = n8879 ;
  assign y19139 = ~1'b0 ;
  assign y19140 = ~n34007 ;
  assign y19141 = 1'b0 ;
  assign y19142 = ~n2203 ;
  assign y19143 = ~n34008 ;
  assign y19144 = ~1'b0 ;
  assign y19145 = ~n34012 ;
  assign y19146 = ~n34016 ;
  assign y19147 = n34018 ;
  assign y19148 = ~n34020 ;
  assign y19149 = ~n34021 ;
  assign y19150 = n28130 ;
  assign y19151 = ~n34023 ;
  assign y19152 = n34025 ;
  assign y19153 = n34026 ;
  assign y19154 = n19668 ;
  assign y19155 = n34027 ;
  assign y19156 = ~n34028 ;
  assign y19157 = ~1'b0 ;
  assign y19158 = n34038 ;
  assign y19159 = n34042 ;
  assign y19160 = ~n34043 ;
  assign y19161 = n34045 ;
  assign y19162 = n34046 ;
  assign y19163 = n34047 ;
  assign y19164 = ~n34050 ;
  assign y19165 = n34053 ;
  assign y19166 = n34055 ;
  assign y19167 = n34058 ;
  assign y19168 = ~1'b0 ;
  assign y19169 = ~1'b0 ;
  assign y19170 = n21981 ;
  assign y19171 = ~n34062 ;
  assign y19172 = ~1'b0 ;
  assign y19173 = ~n34063 ;
  assign y19174 = ~n34064 ;
  assign y19175 = ~1'b0 ;
  assign y19176 = ~1'b0 ;
  assign y19177 = ~1'b0 ;
  assign y19178 = n34065 ;
  assign y19179 = n34066 ;
  assign y19180 = ~1'b0 ;
  assign y19181 = ~1'b0 ;
  assign y19182 = ~1'b0 ;
  assign y19183 = ~1'b0 ;
  assign y19184 = ~n34069 ;
  assign y19185 = ~n34074 ;
  assign y19186 = ~n29443 ;
  assign y19187 = n34083 ;
  assign y19188 = ~n34085 ;
  assign y19189 = ~1'b0 ;
  assign y19190 = n34086 ;
  assign y19191 = ~1'b0 ;
  assign y19192 = ~n20631 ;
  assign y19193 = ~1'b0 ;
  assign y19194 = n34087 ;
  assign y19195 = ~n34091 ;
  assign y19196 = ~1'b0 ;
  assign y19197 = ~n34093 ;
  assign y19198 = ~n34096 ;
  assign y19199 = ~1'b0 ;
  assign y19200 = ~n34100 ;
  assign y19201 = ~n34101 ;
  assign y19202 = n34104 ;
  assign y19203 = ~n34109 ;
  assign y19204 = n34111 ;
  assign y19205 = n34113 ;
  assign y19206 = ~1'b0 ;
  assign y19207 = ~n34116 ;
  assign y19208 = ~1'b0 ;
  assign y19209 = ~n34118 ;
  assign y19210 = n34127 ;
  assign y19211 = ~n34128 ;
  assign y19212 = ~1'b0 ;
  assign y19213 = n34129 ;
  assign y19214 = n34131 ;
  assign y19215 = n34132 ;
  assign y19216 = n34133 ;
  assign y19217 = n34134 ;
  assign y19218 = ~n34137 ;
  assign y19219 = ~1'b0 ;
  assign y19220 = ~n34138 ;
  assign y19221 = ~1'b0 ;
  assign y19222 = n9194 ;
  assign y19223 = 1'b0 ;
  assign y19224 = n34139 ;
  assign y19225 = n34142 ;
  assign y19226 = ~1'b0 ;
  assign y19227 = ~n7768 ;
  assign y19228 = ~n34145 ;
  assign y19229 = n5863 ;
  assign y19230 = ~1'b0 ;
  assign y19231 = ~1'b0 ;
  assign y19232 = ~1'b0 ;
  assign y19233 = ~n8106 ;
  assign y19234 = ~1'b0 ;
  assign y19235 = n34158 ;
  assign y19236 = ~n34160 ;
  assign y19237 = ~1'b0 ;
  assign y19238 = n34161 ;
  assign y19239 = ~1'b0 ;
  assign y19240 = ~1'b0 ;
  assign y19241 = ~1'b0 ;
  assign y19242 = n7495 ;
  assign y19243 = ~1'b0 ;
  assign y19244 = ~1'b0 ;
  assign y19245 = n34165 ;
  assign y19246 = n34167 ;
  assign y19247 = n34168 ;
  assign y19248 = n34169 ;
  assign y19249 = ~n34172 ;
  assign y19250 = n34173 ;
  assign y19251 = n34175 ;
  assign y19252 = ~1'b0 ;
  assign y19253 = ~n34181 ;
  assign y19254 = ~1'b0 ;
  assign y19255 = ~1'b0 ;
  assign y19256 = ~1'b0 ;
  assign y19257 = ~n34182 ;
  assign y19258 = ~1'b0 ;
  assign y19259 = ~1'b0 ;
  assign y19260 = n34183 ;
  assign y19261 = ~n34185 ;
  assign y19262 = 1'b0 ;
  assign y19263 = ~n34187 ;
  assign y19264 = n10217 ;
  assign y19265 = ~n34188 ;
  assign y19266 = n31384 ;
  assign y19267 = ~n34189 ;
  assign y19268 = n34191 ;
  assign y19269 = n34194 ;
  assign y19270 = n34195 ;
  assign y19271 = n22969 ;
  assign y19272 = n34199 ;
  assign y19273 = ~1'b0 ;
  assign y19274 = n34200 ;
  assign y19275 = n34201 ;
  assign y19276 = ~1'b0 ;
  assign y19277 = ~n34202 ;
  assign y19278 = ~n5874 ;
  assign y19279 = ~1'b0 ;
  assign y19280 = n27782 ;
  assign y19281 = ~n34203 ;
  assign y19282 = ~n34204 ;
  assign y19283 = ~n34206 ;
  assign y19284 = 1'b0 ;
  assign y19285 = ~n34207 ;
  assign y19286 = ~1'b0 ;
  assign y19287 = ~n34208 ;
  assign y19288 = ~1'b0 ;
  assign y19289 = ~n34212 ;
  assign y19290 = n34217 ;
  assign y19291 = ~1'b0 ;
  assign y19292 = n34219 ;
  assign y19293 = ~1'b0 ;
  assign y19294 = n34220 ;
  assign y19295 = ~n34223 ;
  assign y19296 = n9477 ;
  assign y19297 = ~n34224 ;
  assign y19298 = n34226 ;
  assign y19299 = n34228 ;
  assign y19300 = ~n34230 ;
  assign y19301 = ~n4207 ;
  assign y19302 = ~1'b0 ;
  assign y19303 = n31496 ;
  assign y19304 = ~n34232 ;
  assign y19305 = n34233 ;
  assign y19306 = n34236 ;
  assign y19307 = n34241 ;
  assign y19308 = ~n34242 ;
  assign y19309 = ~1'b0 ;
  assign y19310 = n34243 ;
  assign y19311 = ~n34244 ;
  assign y19312 = ~1'b0 ;
  assign y19313 = n34245 ;
  assign y19314 = ~1'b0 ;
  assign y19315 = ~1'b0 ;
  assign y19316 = n34247 ;
  assign y19317 = ~1'b0 ;
  assign y19318 = 1'b0 ;
  assign y19319 = ~1'b0 ;
  assign y19320 = ~1'b0 ;
  assign y19321 = ~1'b0 ;
  assign y19322 = ~1'b0 ;
  assign y19323 = ~1'b0 ;
  assign y19324 = ~n34251 ;
  assign y19325 = ~1'b0 ;
  assign y19326 = ~1'b0 ;
  assign y19327 = ~1'b0 ;
  assign y19328 = ~1'b0 ;
  assign y19329 = ~n34252 ;
  assign y19330 = ~n34255 ;
  assign y19331 = n34257 ;
  assign y19332 = ~n34258 ;
  assign y19333 = n34261 ;
  assign y19334 = ~n34262 ;
  assign y19335 = ~n34266 ;
  assign y19336 = ~1'b0 ;
  assign y19337 = ~n34268 ;
  assign y19338 = n34269 ;
  assign y19339 = ~1'b0 ;
  assign y19340 = n34275 ;
  assign y19341 = ~n34279 ;
  assign y19342 = n34282 ;
  assign y19343 = ~n34283 ;
  assign y19344 = ~n8138 ;
  assign y19345 = ~1'b0 ;
  assign y19346 = n34284 ;
  assign y19347 = ~1'b0 ;
  assign y19348 = ~n34285 ;
  assign y19349 = ~1'b0 ;
  assign y19350 = ~1'b0 ;
  assign y19351 = ~n34286 ;
  assign y19352 = 1'b0 ;
  assign y19353 = n34287 ;
  assign y19354 = n34288 ;
  assign y19355 = ~n34293 ;
  assign y19356 = 1'b0 ;
  assign y19357 = ~n25245 ;
  assign y19358 = ~n34297 ;
  assign y19359 = ~n34301 ;
  assign y19360 = n34307 ;
  assign y19361 = ~1'b0 ;
  assign y19362 = ~n34308 ;
  assign y19363 = ~n34314 ;
  assign y19364 = ~n34315 ;
  assign y19365 = n34317 ;
  assign y19366 = ~1'b0 ;
  assign y19367 = ~1'b0 ;
  assign y19368 = n34318 ;
  assign y19369 = ~n12553 ;
  assign y19370 = n34319 ;
  assign y19371 = n34320 ;
  assign y19372 = n8570 ;
  assign y19373 = n34322 ;
  assign y19374 = n34330 ;
  assign y19375 = ~n34332 ;
  assign y19376 = n34335 ;
  assign y19377 = n34336 ;
  assign y19378 = ~n34338 ;
  assign y19379 = n34339 ;
  assign y19380 = ~1'b0 ;
  assign y19381 = ~n34343 ;
  assign y19382 = ~1'b0 ;
  assign y19383 = n34344 ;
  assign y19384 = n34345 ;
  assign y19385 = ~1'b0 ;
  assign y19386 = ~n34346 ;
  assign y19387 = ~n34347 ;
  assign y19388 = ~1'b0 ;
  assign y19389 = n34351 ;
  assign y19390 = ~n34352 ;
  assign y19391 = ~1'b0 ;
  assign y19392 = n9424 ;
  assign y19393 = ~1'b0 ;
  assign y19394 = ~n34353 ;
  assign y19395 = n34354 ;
  assign y19396 = n34355 ;
  assign y19397 = ~n34357 ;
  assign y19398 = ~1'b0 ;
  assign y19399 = n34359 ;
  assign y19400 = ~n34361 ;
  assign y19401 = ~1'b0 ;
  assign y19402 = n34366 ;
  assign y19403 = n34368 ;
  assign y19404 = n34388 ;
  assign y19405 = ~n34391 ;
  assign y19406 = ~n34393 ;
  assign y19407 = ~n34394 ;
  assign y19408 = 1'b0 ;
  assign y19409 = n34395 ;
  assign y19410 = 1'b0 ;
  assign y19411 = ~n34397 ;
  assign y19412 = ~n2663 ;
  assign y19413 = ~n34398 ;
  assign y19414 = ~1'b0 ;
  assign y19415 = ~n34400 ;
  assign y19416 = n34402 ;
  assign y19417 = ~n34403 ;
  assign y19418 = ~n34410 ;
  assign y19419 = ~n34414 ;
  assign y19420 = n34415 ;
  assign y19421 = ~1'b0 ;
  assign y19422 = n34423 ;
  assign y19423 = n34424 ;
  assign y19424 = n34426 ;
  assign y19425 = ~1'b0 ;
  assign y19426 = n34437 ;
  assign y19427 = ~n34438 ;
  assign y19428 = n34440 ;
  assign y19429 = ~1'b0 ;
  assign y19430 = ~1'b0 ;
  assign y19431 = ~1'b0 ;
  assign y19432 = ~n34441 ;
  assign y19433 = ~1'b0 ;
  assign y19434 = ~n34443 ;
  assign y19435 = ~n34444 ;
  assign y19436 = ~n34447 ;
  assign y19437 = ~n34451 ;
  assign y19438 = 1'b0 ;
  assign y19439 = ~n34453 ;
  assign y19440 = ~1'b0 ;
  assign y19441 = ~1'b0 ;
  assign y19442 = ~n34456 ;
  assign y19443 = ~n34457 ;
  assign y19444 = n34463 ;
  assign y19445 = ~n34464 ;
  assign y19446 = n34466 ;
  assign y19447 = ~1'b0 ;
  assign y19448 = ~n34473 ;
  assign y19449 = ~n34475 ;
  assign y19450 = ~n34478 ;
  assign y19451 = n34483 ;
  assign y19452 = ~n34490 ;
  assign y19453 = ~n34491 ;
  assign y19454 = n34499 ;
  assign y19455 = ~n34502 ;
  assign y19456 = n34504 ;
  assign y19457 = n2283 ;
  assign y19458 = ~n34510 ;
  assign y19459 = ~n34514 ;
  assign y19460 = n34515 ;
  assign y19461 = ~1'b0 ;
  assign y19462 = ~n34517 ;
  assign y19463 = n34519 ;
  assign y19464 = n34521 ;
  assign y19465 = n34523 ;
  assign y19466 = ~n477 ;
  assign y19467 = n34524 ;
  assign y19468 = n34525 ;
  assign y19469 = ~1'b0 ;
  assign y19470 = ~1'b0 ;
  assign y19471 = ~n34531 ;
  assign y19472 = n34532 ;
  assign y19473 = ~1'b0 ;
  assign y19474 = n34533 ;
  assign y19475 = ~1'b0 ;
  assign y19476 = ~n34535 ;
  assign y19477 = ~n34537 ;
  assign y19478 = n34538 ;
  assign y19479 = n34539 ;
  assign y19480 = ~1'b0 ;
  assign y19481 = ~1'b0 ;
  assign y19482 = ~1'b0 ;
  assign y19483 = ~n15478 ;
  assign y19484 = n34540 ;
  assign y19485 = n34541 ;
  assign y19486 = n34542 ;
  assign y19487 = ~n34543 ;
  assign y19488 = n34546 ;
  assign y19489 = n34548 ;
  assign y19490 = ~1'b0 ;
  assign y19491 = ~n34550 ;
  assign y19492 = n34551 ;
  assign y19493 = n34555 ;
  assign y19494 = n34556 ;
  assign y19495 = n34561 ;
  assign y19496 = ~n34562 ;
  assign y19497 = ~1'b0 ;
  assign y19498 = n34564 ;
  assign y19499 = n34565 ;
  assign y19500 = ~1'b0 ;
  assign y19501 = ~1'b0 ;
  assign y19502 = n34566 ;
  assign y19503 = ~n34568 ;
  assign y19504 = ~n34569 ;
  assign y19505 = n34570 ;
  assign y19506 = n34575 ;
  assign y19507 = n34577 ;
  assign y19508 = ~n34581 ;
  assign y19509 = ~n34590 ;
  assign y19510 = ~n34593 ;
  assign y19511 = n25114 ;
  assign y19512 = n34596 ;
  assign y19513 = ~1'b0 ;
  assign y19514 = n34597 ;
  assign y19515 = ~1'b0 ;
  assign y19516 = ~n34600 ;
  assign y19517 = ~1'b0 ;
  assign y19518 = n34603 ;
  assign y19519 = n34604 ;
  assign y19520 = ~n34608 ;
  assign y19521 = ~1'b0 ;
  assign y19522 = n34610 ;
  assign y19523 = 1'b0 ;
  assign y19524 = ~n34611 ;
  assign y19525 = n21192 ;
  assign y19526 = ~n34612 ;
  assign y19527 = n34614 ;
  assign y19528 = ~1'b0 ;
  assign y19529 = ~1'b0 ;
  assign y19530 = ~1'b0 ;
  assign y19531 = ~1'b0 ;
  assign y19532 = ~1'b0 ;
  assign y19533 = ~n34615 ;
  assign y19534 = ~n17030 ;
  assign y19535 = ~1'b0 ;
  assign y19536 = ~1'b0 ;
  assign y19537 = n34616 ;
  assign y19538 = ~1'b0 ;
  assign y19539 = n34617 ;
  assign y19540 = ~1'b0 ;
  assign y19541 = ~1'b0 ;
  assign y19542 = ~1'b0 ;
  assign y19543 = ~n34618 ;
  assign y19544 = n34619 ;
  assign y19545 = n34622 ;
  assign y19546 = n34628 ;
  assign y19547 = 1'b0 ;
  assign y19548 = ~n34630 ;
  assign y19549 = ~1'b0 ;
  assign y19550 = ~1'b0 ;
  assign y19551 = ~1'b0 ;
  assign y19552 = n34633 ;
  assign y19553 = ~n34634 ;
  assign y19554 = n34638 ;
  assign y19555 = ~n34643 ;
  assign y19556 = ~n27514 ;
  assign y19557 = ~1'b0 ;
  assign y19558 = ~1'b0 ;
  assign y19559 = ~n28070 ;
  assign y19560 = ~n34645 ;
  assign y19561 = n34646 ;
  assign y19562 = n34647 ;
  assign y19563 = n34650 ;
  assign y19564 = ~1'b0 ;
  assign y19565 = ~1'b0 ;
  assign y19566 = ~n34654 ;
  assign y19567 = n34655 ;
  assign y19568 = ~n34656 ;
  assign y19569 = ~n34658 ;
  assign y19570 = ~1'b0 ;
  assign y19571 = n34660 ;
  assign y19572 = ~n34664 ;
  assign y19573 = ~n34667 ;
  assign y19574 = ~1'b0 ;
  assign y19575 = ~n34669 ;
  assign y19576 = ~1'b0 ;
  assign y19577 = ~n34670 ;
  assign y19578 = ~n34671 ;
  assign y19579 = ~1'b0 ;
  assign y19580 = n34680 ;
  assign y19581 = ~n34684 ;
  assign y19582 = ~1'b0 ;
  assign y19583 = ~n34687 ;
  assign y19584 = n34689 ;
  assign y19585 = ~1'b0 ;
  assign y19586 = ~1'b0 ;
  assign y19587 = ~n34691 ;
  assign y19588 = ~1'b0 ;
  assign y19589 = ~n34693 ;
  assign y19590 = 1'b0 ;
  assign y19591 = n34700 ;
  assign y19592 = ~n34707 ;
  assign y19593 = ~1'b0 ;
  assign y19594 = ~n443 ;
  assign y19595 = ~n34712 ;
  assign y19596 = n34715 ;
  assign y19597 = ~1'b0 ;
  assign y19598 = ~n34716 ;
  assign y19599 = n34717 ;
  assign y19600 = n34718 ;
  assign y19601 = ~n34721 ;
  assign y19602 = ~n34722 ;
  assign y19603 = ~n34725 ;
  assign y19604 = n34728 ;
  assign y19605 = ~n33906 ;
  assign y19606 = n34730 ;
  assign y19607 = n34732 ;
  assign y19608 = ~n34733 ;
  assign y19609 = n34734 ;
  assign y19610 = ~1'b0 ;
  assign y19611 = ~n34735 ;
  assign y19612 = ~n34736 ;
  assign y19613 = ~n34738 ;
  assign y19614 = ~1'b0 ;
  assign y19615 = ~n28172 ;
  assign y19616 = n34741 ;
  assign y19617 = n23948 ;
  assign y19618 = n34745 ;
  assign y19619 = ~1'b0 ;
  assign y19620 = n34746 ;
  assign y19621 = ~1'b0 ;
  assign y19622 = n34747 ;
  assign y19623 = ~1'b0 ;
  assign y19624 = ~1'b0 ;
  assign y19625 = ~n34748 ;
  assign y19626 = n34752 ;
  assign y19627 = n34755 ;
  assign y19628 = ~n31051 ;
  assign y19629 = ~1'b0 ;
  assign y19630 = ~n34756 ;
  assign y19631 = n34757 ;
  assign y19632 = ~1'b0 ;
  assign y19633 = ~1'b0 ;
  assign y19634 = ~1'b0 ;
  assign y19635 = ~n16978 ;
  assign y19636 = ~n34758 ;
  assign y19637 = ~1'b0 ;
  assign y19638 = ~n4229 ;
  assign y19639 = ~n34762 ;
  assign y19640 = ~1'b0 ;
  assign y19641 = ~n34763 ;
  assign y19642 = ~n34765 ;
  assign y19643 = ~n34768 ;
  assign y19644 = ~n34771 ;
  assign y19645 = ~n34773 ;
  assign y19646 = ~1'b0 ;
  assign y19647 = ~1'b0 ;
  assign y19648 = ~n34774 ;
  assign y19649 = ~n34775 ;
  assign y19650 = 1'b0 ;
  assign y19651 = n34778 ;
  assign y19652 = ~n34784 ;
  assign y19653 = ~n34785 ;
  assign y19654 = ~n34786 ;
  assign y19655 = 1'b0 ;
  assign y19656 = ~n34793 ;
  assign y19657 = n34796 ;
  assign y19658 = ~n34797 ;
  assign y19659 = ~n34799 ;
  assign y19660 = n34800 ;
  assign y19661 = 1'b0 ;
  assign y19662 = ~n14384 ;
  assign y19663 = ~n34801 ;
  assign y19664 = ~n34805 ;
  assign y19665 = ~1'b0 ;
  assign y19666 = ~n34806 ;
  assign y19667 = ~n34808 ;
  assign y19668 = n34809 ;
  assign y19669 = ~n34811 ;
  assign y19670 = 1'b0 ;
  assign y19671 = 1'b0 ;
  assign y19672 = n34812 ;
  assign y19673 = ~n34817 ;
  assign y19674 = ~n34823 ;
  assign y19675 = ~1'b0 ;
  assign y19676 = n34824 ;
  assign y19677 = ~n34826 ;
  assign y19678 = n34829 ;
  assign y19679 = n22158 ;
  assign y19680 = ~n34839 ;
  assign y19681 = ~n34840 ;
  assign y19682 = ~n15229 ;
  assign y19683 = ~n34842 ;
  assign y19684 = n34843 ;
  assign y19685 = n34845 ;
  assign y19686 = ~n34848 ;
  assign y19687 = ~1'b0 ;
  assign y19688 = ~1'b0 ;
  assign y19689 = ~1'b0 ;
  assign y19690 = ~n34851 ;
  assign y19691 = ~1'b0 ;
  assign y19692 = n34853 ;
  assign y19693 = n34854 ;
  assign y19694 = n34856 ;
  assign y19695 = ~n34857 ;
  assign y19696 = n34859 ;
  assign y19697 = ~n34861 ;
  assign y19698 = ~n34863 ;
  assign y19699 = ~1'b0 ;
  assign y19700 = ~1'b0 ;
  assign y19701 = ~1'b0 ;
  assign y19702 = ~n34864 ;
  assign y19703 = ~1'b0 ;
  assign y19704 = ~n34866 ;
  assign y19705 = ~1'b0 ;
  assign y19706 = ~n34870 ;
  assign y19707 = ~1'b0 ;
  assign y19708 = ~n34873 ;
  assign y19709 = ~1'b0 ;
  assign y19710 = n34877 ;
  assign y19711 = ~1'b0 ;
  assign y19712 = n34879 ;
  assign y19713 = ~1'b0 ;
  assign y19714 = ~n34881 ;
  assign y19715 = n7866 ;
  assign y19716 = n34882 ;
  assign y19717 = ~1'b0 ;
  assign y19718 = ~1'b0 ;
  assign y19719 = ~n34885 ;
  assign y19720 = ~n34887 ;
  assign y19721 = n34890 ;
  assign y19722 = ~n34891 ;
  assign y19723 = ~n34893 ;
  assign y19724 = ~n34896 ;
  assign y19725 = 1'b0 ;
  assign y19726 = ~1'b0 ;
  assign y19727 = ~1'b0 ;
  assign y19728 = ~n34904 ;
  assign y19729 = ~n34906 ;
  assign y19730 = ~1'b0 ;
  assign y19731 = ~n34908 ;
  assign y19732 = ~n34910 ;
  assign y19733 = n34914 ;
  assign y19734 = ~n34918 ;
  assign y19735 = n19192 ;
  assign y19736 = 1'b0 ;
  assign y19737 = ~1'b0 ;
  assign y19738 = ~n34922 ;
  assign y19739 = n34929 ;
  assign y19740 = n34932 ;
  assign y19741 = ~1'b0 ;
  assign y19742 = ~1'b0 ;
  assign y19743 = n34934 ;
  assign y19744 = ~n34935 ;
  assign y19745 = ~n15550 ;
  assign y19746 = n5497 ;
  assign y19747 = ~1'b0 ;
  assign y19748 = ~n34939 ;
  assign y19749 = n34942 ;
  assign y19750 = n34951 ;
  assign y19751 = 1'b0 ;
  assign y19752 = 1'b0 ;
  assign y19753 = n34956 ;
  assign y19754 = ~n34958 ;
  assign y19755 = ~n34959 ;
  assign y19756 = ~1'b0 ;
  assign y19757 = ~1'b0 ;
  assign y19758 = ~n34960 ;
  assign y19759 = ~1'b0 ;
  assign y19760 = n34965 ;
  assign y19761 = ~n34967 ;
  assign y19762 = ~1'b0 ;
  assign y19763 = n34968 ;
  assign y19764 = ~1'b0 ;
  assign y19765 = ~1'b0 ;
  assign y19766 = ~1'b0 ;
  assign y19767 = n34969 ;
  assign y19768 = ~n34971 ;
  assign y19769 = n34972 ;
  assign y19770 = ~n2829 ;
  assign y19771 = n29402 ;
  assign y19772 = ~n34975 ;
  assign y19773 = n34978 ;
  assign y19774 = ~n34980 ;
  assign y19775 = n436 ;
  assign y19776 = n34982 ;
  assign y19777 = n34986 ;
  assign y19778 = n34987 ;
  assign y19779 = ~n34988 ;
  assign y19780 = ~n34989 ;
  assign y19781 = ~n34990 ;
  assign y19782 = ~n34991 ;
  assign y19783 = ~n34994 ;
  assign y19784 = ~n34999 ;
  assign y19785 = ~n35003 ;
  assign y19786 = n35004 ;
  assign y19787 = n35007 ;
  assign y19788 = ~1'b0 ;
  assign y19789 = ~1'b0 ;
  assign y19790 = ~n17094 ;
  assign y19791 = n35008 ;
  assign y19792 = ~1'b0 ;
  assign y19793 = ~1'b0 ;
  assign y19794 = ~1'b0 ;
  assign y19795 = ~n35010 ;
  assign y19796 = ~n61 ;
  assign y19797 = ~1'b0 ;
  assign y19798 = ~1'b0 ;
  assign y19799 = ~n35014 ;
  assign y19800 = ~1'b0 ;
  assign y19801 = ~n35015 ;
  assign y19802 = n35017 ;
  assign y19803 = ~n5953 ;
  assign y19804 = ~n35018 ;
  assign y19805 = ~1'b0 ;
  assign y19806 = n35020 ;
  assign y19807 = ~n35027 ;
  assign y19808 = n35029 ;
  assign y19809 = ~n35030 ;
  assign y19810 = ~1'b0 ;
  assign y19811 = ~1'b0 ;
  assign y19812 = ~n35031 ;
  assign y19813 = ~n35032 ;
  assign y19814 = ~1'b0 ;
  assign y19815 = n8284 ;
  assign y19816 = ~n26571 ;
  assign y19817 = ~n35033 ;
  assign y19818 = ~1'b0 ;
  assign y19819 = ~1'b0 ;
  assign y19820 = n35034 ;
  assign y19821 = ~n18006 ;
  assign y19822 = n35035 ;
  assign y19823 = n35036 ;
  assign y19824 = ~n35038 ;
  assign y19825 = ~n35041 ;
  assign y19826 = ~n35042 ;
  assign y19827 = ~n35044 ;
  assign y19828 = ~1'b0 ;
  assign y19829 = ~n17035 ;
  assign y19830 = ~n35045 ;
  assign y19831 = n35046 ;
  assign y19832 = ~n35048 ;
  assign y19833 = 1'b0 ;
  assign y19834 = ~n35053 ;
  assign y19835 = ~n35054 ;
  assign y19836 = n3280 ;
  assign y19837 = ~n35056 ;
  assign y19838 = n35061 ;
  assign y19839 = n35065 ;
  assign y19840 = ~n35067 ;
  assign y19841 = ~1'b0 ;
  assign y19842 = ~n35070 ;
  assign y19843 = ~1'b0 ;
  assign y19844 = ~n35071 ;
  assign y19845 = ~n35075 ;
  assign y19846 = n35078 ;
  assign y19847 = ~n35080 ;
  assign y19848 = n35081 ;
  assign y19849 = ~n35088 ;
  assign y19850 = n35089 ;
  assign y19851 = 1'b0 ;
  assign y19852 = ~n35090 ;
  assign y19853 = n35092 ;
  assign y19854 = n35093 ;
  assign y19855 = n35094 ;
  assign y19856 = ~n35095 ;
  assign y19857 = ~n35099 ;
  assign y19858 = ~n35100 ;
  assign y19859 = ~n35104 ;
  assign y19860 = ~n35106 ;
  assign y19861 = ~n35107 ;
  assign y19862 = n35110 ;
  assign y19863 = ~1'b0 ;
  assign y19864 = ~1'b0 ;
  assign y19865 = ~1'b0 ;
  assign y19866 = 1'b0 ;
  assign y19867 = ~1'b0 ;
  assign y19868 = n35115 ;
  assign y19869 = n35116 ;
  assign y19870 = ~n35122 ;
  assign y19871 = 1'b0 ;
  assign y19872 = n35126 ;
  assign y19873 = ~1'b0 ;
  assign y19874 = n35130 ;
  assign y19875 = ~n35131 ;
  assign y19876 = ~1'b0 ;
  assign y19877 = n35133 ;
  assign y19878 = 1'b0 ;
  assign y19879 = ~n35137 ;
  assign y19880 = ~1'b0 ;
  assign y19881 = ~1'b0 ;
  assign y19882 = n35138 ;
  assign y19883 = ~n35143 ;
  assign y19884 = ~n16435 ;
  assign y19885 = ~1'b0 ;
  assign y19886 = ~1'b0 ;
  assign y19887 = ~n18727 ;
  assign y19888 = ~n6080 ;
  assign y19889 = ~1'b0 ;
  assign y19890 = ~n35145 ;
  assign y19891 = ~1'b0 ;
  assign y19892 = n35146 ;
  assign y19893 = ~1'b0 ;
  assign y19894 = ~n35151 ;
  assign y19895 = n6043 ;
  assign y19896 = ~n19418 ;
  assign y19897 = n1422 ;
  assign y19898 = n35154 ;
  assign y19899 = n35157 ;
  assign y19900 = ~n35158 ;
  assign y19901 = n35160 ;
  assign y19902 = ~n35161 ;
  assign y19903 = ~1'b0 ;
  assign y19904 = ~n19705 ;
  assign y19905 = n35165 ;
  assign y19906 = ~1'b0 ;
  assign y19907 = ~1'b0 ;
  assign y19908 = n35166 ;
  assign y19909 = ~1'b0 ;
  assign y19910 = ~1'b0 ;
  assign y19911 = n35169 ;
  assign y19912 = ~1'b0 ;
  assign y19913 = n35170 ;
  assign y19914 = ~n35172 ;
  assign y19915 = n35173 ;
  assign y19916 = ~1'b0 ;
  assign y19917 = ~n35174 ;
  assign y19918 = n19158 ;
  assign y19919 = n35176 ;
  assign y19920 = ~n35177 ;
  assign y19921 = ~n35179 ;
  assign y19922 = n35180 ;
  assign y19923 = n35181 ;
  assign y19924 = 1'b0 ;
  assign y19925 = n35183 ;
  assign y19926 = n3489 ;
  assign y19927 = n35185 ;
  assign y19928 = ~1'b0 ;
  assign y19929 = ~1'b0 ;
  assign y19930 = n35197 ;
  assign y19931 = n35200 ;
  assign y19932 = ~n35201 ;
  assign y19933 = ~1'b0 ;
  assign y19934 = ~n35202 ;
  assign y19935 = n35204 ;
  assign y19936 = n35207 ;
  assign y19937 = ~1'b0 ;
  assign y19938 = ~1'b0 ;
  assign y19939 = ~n35211 ;
  assign y19940 = ~n35212 ;
  assign y19941 = ~1'b0 ;
  assign y19942 = n14649 ;
  assign y19943 = n35214 ;
  assign y19944 = 1'b0 ;
  assign y19945 = ~1'b0 ;
  assign y19946 = n35215 ;
  assign y19947 = ~1'b0 ;
  assign y19948 = n35217 ;
  assign y19949 = ~n35219 ;
  assign y19950 = ~n35221 ;
  assign y19951 = ~1'b0 ;
  assign y19952 = n35223 ;
  assign y19953 = ~n34218 ;
  assign y19954 = ~n35224 ;
  assign y19955 = ~n35228 ;
  assign y19956 = ~n35231 ;
  assign y19957 = ~n3595 ;
  assign y19958 = n35233 ;
  assign y19959 = ~1'b0 ;
  assign y19960 = n35234 ;
  assign y19961 = n35237 ;
  assign y19962 = n35238 ;
  assign y19963 = n35239 ;
  assign y19964 = n35241 ;
  assign y19965 = ~1'b0 ;
  assign y19966 = ~n35243 ;
  assign y19967 = ~n35244 ;
  assign y19968 = ~n35248 ;
  assign y19969 = n35251 ;
  assign y19970 = n35259 ;
  assign y19971 = ~1'b0 ;
  assign y19972 = n35262 ;
  assign y19973 = n35264 ;
  assign y19974 = ~n31048 ;
  assign y19975 = n35267 ;
  assign y19976 = ~n35270 ;
  assign y19977 = ~n35271 ;
  assign y19978 = n35272 ;
  assign y19979 = n35274 ;
  assign y19980 = n35277 ;
  assign y19981 = n35283 ;
  assign y19982 = 1'b0 ;
  assign y19983 = ~n35287 ;
  assign y19984 = ~1'b0 ;
  assign y19985 = ~n35288 ;
  assign y19986 = ~n35292 ;
  assign y19987 = n35294 ;
  assign y19988 = ~1'b0 ;
  assign y19989 = ~n35298 ;
  assign y19990 = n35303 ;
  assign y19991 = n35304 ;
  assign y19992 = n16636 ;
  assign y19993 = ~1'b0 ;
  assign y19994 = ~n708 ;
  assign y19995 = n35313 ;
  assign y19996 = ~n35318 ;
  assign y19997 = n35319 ;
  assign y19998 = ~n35321 ;
  assign y19999 = ~n35322 ;
  assign y20000 = ~1'b0 ;
  assign y20001 = ~1'b0 ;
  assign y20002 = ~1'b0 ;
  assign y20003 = n35323 ;
  assign y20004 = n35325 ;
  assign y20005 = ~n35326 ;
  assign y20006 = ~1'b0 ;
  assign y20007 = n35330 ;
  assign y20008 = ~n35331 ;
  assign y20009 = ~n19543 ;
  assign y20010 = ~n21865 ;
  assign y20011 = ~n35337 ;
  assign y20012 = ~n35344 ;
  assign y20013 = ~1'b0 ;
  assign y20014 = n35345 ;
  assign y20015 = n35347 ;
  assign y20016 = ~1'b0 ;
  assign y20017 = ~1'b0 ;
  assign y20018 = ~1'b0 ;
  assign y20019 = ~n35349 ;
  assign y20020 = 1'b0 ;
  assign y20021 = n35354 ;
  assign y20022 = n23571 ;
  assign y20023 = 1'b0 ;
  assign y20024 = ~n22131 ;
  assign y20025 = ~1'b0 ;
  assign y20026 = ~1'b0 ;
  assign y20027 = n35360 ;
  assign y20028 = n35362 ;
  assign y20029 = ~1'b0 ;
  assign y20030 = ~1'b0 ;
  assign y20031 = n35364 ;
  assign y20032 = ~1'b0 ;
  assign y20033 = ~1'b0 ;
  assign y20034 = ~n35365 ;
  assign y20035 = ~n35368 ;
  assign y20036 = ~1'b0 ;
  assign y20037 = n35373 ;
  assign y20038 = n35374 ;
  assign y20039 = ~n35379 ;
  assign y20040 = ~n35382 ;
  assign y20041 = ~n35385 ;
  assign y20042 = n35390 ;
  assign y20043 = n35392 ;
  assign y20044 = n35394 ;
  assign y20045 = ~n7089 ;
  assign y20046 = ~1'b0 ;
  assign y20047 = ~1'b0 ;
  assign y20048 = ~n30751 ;
  assign y20049 = n35396 ;
  assign y20050 = ~n35398 ;
  assign y20051 = ~1'b0 ;
  assign y20052 = ~1'b0 ;
  assign y20053 = ~1'b0 ;
  assign y20054 = n35401 ;
  assign y20055 = ~1'b0 ;
  assign y20056 = ~n35403 ;
  assign y20057 = ~n35408 ;
  assign y20058 = n20641 ;
  assign y20059 = ~1'b0 ;
  assign y20060 = ~n35411 ;
  assign y20061 = ~n35416 ;
  assign y20062 = ~n35418 ;
  assign y20063 = n35422 ;
  assign y20064 = n35423 ;
  assign y20065 = n16709 ;
  assign y20066 = 1'b0 ;
  assign y20067 = n35424 ;
  assign y20068 = ~n35428 ;
  assign y20069 = n35433 ;
  assign y20070 = n35435 ;
  assign y20071 = ~n19949 ;
  assign y20072 = n35436 ;
  assign y20073 = ~n35437 ;
  assign y20074 = n35439 ;
  assign y20075 = ~n35440 ;
  assign y20076 = ~1'b0 ;
  assign y20077 = ~1'b0 ;
  assign y20078 = n35443 ;
  assign y20079 = n35445 ;
  assign y20080 = n35446 ;
  assign y20081 = ~n35447 ;
  assign y20082 = n35450 ;
  assign y20083 = n33214 ;
  assign y20084 = ~n35451 ;
  assign y20085 = ~n35457 ;
  assign y20086 = ~1'b0 ;
  assign y20087 = n35462 ;
  assign y20088 = ~n35464 ;
  assign y20089 = ~n35466 ;
  assign y20090 = ~1'b0 ;
  assign y20091 = ~1'b0 ;
  assign y20092 = n35472 ;
  assign y20093 = ~1'b0 ;
  assign y20094 = ~n35477 ;
  assign y20095 = 1'b0 ;
  assign y20096 = n35479 ;
  assign y20097 = ~1'b0 ;
  assign y20098 = ~n35480 ;
  assign y20099 = ~n35482 ;
  assign y20100 = n35485 ;
  assign y20101 = n35486 ;
  assign y20102 = n35487 ;
  assign y20103 = ~1'b0 ;
  assign y20104 = ~n35490 ;
  assign y20105 = n35491 ;
  assign y20106 = ~1'b0 ;
  assign y20107 = n24926 ;
  assign y20108 = ~1'b0 ;
  assign y20109 = n35492 ;
  assign y20110 = n3416 ;
  assign y20111 = ~1'b0 ;
  assign y20112 = ~1'b0 ;
  assign y20113 = ~1'b0 ;
  assign y20114 = ~1'b0 ;
  assign y20115 = n35495 ;
  assign y20116 = ~n35498 ;
  assign y20117 = ~1'b0 ;
  assign y20118 = ~1'b0 ;
  assign y20119 = n35500 ;
  assign y20120 = n35508 ;
  assign y20121 = n7234 ;
  assign y20122 = n35509 ;
  assign y20123 = ~n18087 ;
  assign y20124 = ~n21468 ;
  assign y20125 = ~n35512 ;
  assign y20126 = ~1'b0 ;
  assign y20127 = ~1'b0 ;
  assign y20128 = 1'b0 ;
  assign y20129 = ~1'b0 ;
  assign y20130 = ~1'b0 ;
  assign y20131 = n35514 ;
  assign y20132 = n35517 ;
  assign y20133 = n35519 ;
  assign y20134 = ~1'b0 ;
  assign y20135 = ~1'b0 ;
  assign y20136 = n35521 ;
  assign y20137 = ~1'b0 ;
  assign y20138 = n35523 ;
  assign y20139 = n35526 ;
  assign y20140 = n35531 ;
  assign y20141 = n35532 ;
  assign y20142 = ~n35539 ;
  assign y20143 = n35382 ;
  assign y20144 = ~1'b0 ;
  assign y20145 = 1'b0 ;
  assign y20146 = ~n6200 ;
  assign y20147 = n35544 ;
  assign y20148 = n35546 ;
  assign y20149 = ~1'b0 ;
  assign y20150 = ~1'b0 ;
  assign y20151 = n35548 ;
  assign y20152 = ~n35549 ;
  assign y20153 = ~n35552 ;
  assign y20154 = ~1'b0 ;
  assign y20155 = n35555 ;
  assign y20156 = ~1'b0 ;
  assign y20157 = ~n35557 ;
  assign y20158 = ~1'b0 ;
  assign y20159 = n35561 ;
  assign y20160 = ~n35569 ;
  assign y20161 = n35574 ;
  assign y20162 = ~n35575 ;
  assign y20163 = n35577 ;
  assign y20164 = ~n35583 ;
  assign y20165 = ~1'b0 ;
  assign y20166 = n35587 ;
  assign y20167 = n35591 ;
  assign y20168 = ~n35600 ;
  assign y20169 = n35601 ;
  assign y20170 = ~1'b0 ;
  assign y20171 = ~1'b0 ;
  assign y20172 = ~1'b0 ;
  assign y20173 = ~1'b0 ;
  assign y20174 = n35604 ;
  assign y20175 = ~1'b0 ;
  assign y20176 = n35611 ;
  assign y20177 = ~n35612 ;
  assign y20178 = n35615 ;
  assign y20179 = ~n35620 ;
  assign y20180 = n35622 ;
  assign y20181 = ~n35627 ;
  assign y20182 = n35628 ;
  assign y20183 = ~1'b0 ;
  assign y20184 = ~n10302 ;
  assign y20185 = n35636 ;
  assign y20186 = ~n8404 ;
  assign y20187 = ~n35639 ;
  assign y20188 = ~1'b0 ;
  assign y20189 = ~1'b0 ;
  assign y20190 = ~n35641 ;
  assign y20191 = ~1'b0 ;
  assign y20192 = ~1'b0 ;
  assign y20193 = ~1'b0 ;
  assign y20194 = ~n28172 ;
  assign y20195 = n35643 ;
  assign y20196 = n35644 ;
  assign y20197 = ~n35646 ;
  assign y20198 = ~n35647 ;
  assign y20199 = ~n35651 ;
  assign y20200 = ~n35655 ;
  assign y20201 = ~n15331 ;
  assign y20202 = ~1'b0 ;
  assign y20203 = 1'b0 ;
  assign y20204 = ~n35658 ;
  assign y20205 = n35660 ;
  assign y20206 = n35662 ;
  assign y20207 = ~1'b0 ;
  assign y20208 = ~1'b0 ;
  assign y20209 = ~1'b0 ;
  assign y20210 = ~1'b0 ;
  assign y20211 = n35667 ;
  assign y20212 = n35668 ;
  assign y20213 = n35670 ;
  assign y20214 = ~n17325 ;
  assign y20215 = 1'b0 ;
  assign y20216 = ~1'b0 ;
  assign y20217 = ~1'b0 ;
  assign y20218 = ~n35671 ;
  assign y20219 = ~n35672 ;
  assign y20220 = ~1'b0 ;
  assign y20221 = ~n35673 ;
  assign y20222 = n35675 ;
  assign y20223 = ~1'b0 ;
  assign y20224 = n35678 ;
  assign y20225 = ~n35679 ;
  assign y20226 = n35681 ;
  assign y20227 = n35682 ;
  assign y20228 = n3061 ;
  assign y20229 = ~n35685 ;
  assign y20230 = n35686 ;
  assign y20231 = n8961 ;
  assign y20232 = ~n35689 ;
  assign y20233 = n35693 ;
  assign y20234 = ~1'b0 ;
  assign y20235 = n35696 ;
  assign y20236 = ~n35698 ;
  assign y20237 = n35701 ;
  assign y20238 = ~1'b0 ;
  assign y20239 = n35703 ;
  assign y20240 = ~1'b0 ;
  assign y20241 = ~1'b0 ;
  assign y20242 = ~n35705 ;
  assign y20243 = ~1'b0 ;
  assign y20244 = ~n35708 ;
  assign y20245 = ~1'b0 ;
  assign y20246 = ~n35714 ;
  assign y20247 = ~n35716 ;
  assign y20248 = ~n35718 ;
  assign y20249 = n35719 ;
  assign y20250 = ~1'b0 ;
  assign y20251 = n35723 ;
  assign y20252 = n35724 ;
  assign y20253 = n35726 ;
  assign y20254 = n35727 ;
  assign y20255 = ~1'b0 ;
  assign y20256 = ~n35729 ;
  assign y20257 = n35737 ;
  assign y20258 = ~n35738 ;
  assign y20259 = ~n20158 ;
  assign y20260 = ~n35743 ;
  assign y20261 = n20346 ;
  assign y20262 = ~n35747 ;
  assign y20263 = ~1'b0 ;
  assign y20264 = n35749 ;
  assign y20265 = n35752 ;
  assign y20266 = ~1'b0 ;
  assign y20267 = ~n5350 ;
  assign y20268 = n35755 ;
  assign y20269 = ~n35758 ;
  assign y20270 = n35759 ;
  assign y20271 = ~n35763 ;
  assign y20272 = ~n35765 ;
  assign y20273 = n35766 ;
  assign y20274 = ~n35785 ;
  assign y20275 = ~n35790 ;
  assign y20276 = n35792 ;
  assign y20277 = ~n35794 ;
  assign y20278 = n35799 ;
  assign y20279 = ~n35804 ;
  assign y20280 = ~1'b0 ;
  assign y20281 = ~n35806 ;
  assign y20282 = n35808 ;
  assign y20283 = n35809 ;
  assign y20284 = ~n35811 ;
  assign y20285 = ~1'b0 ;
  assign y20286 = ~n14453 ;
  assign y20287 = ~1'b0 ;
  assign y20288 = ~n35812 ;
  assign y20289 = n35818 ;
  assign y20290 = ~n35825 ;
  assign y20291 = ~n35826 ;
  assign y20292 = ~n35827 ;
  assign y20293 = n35829 ;
  assign y20294 = ~n35831 ;
  assign y20295 = n35833 ;
  assign y20296 = ~1'b0 ;
  assign y20297 = ~n35837 ;
  assign y20298 = ~1'b0 ;
  assign y20299 = ~1'b0 ;
  assign y20300 = ~1'b0 ;
  assign y20301 = ~n35843 ;
  assign y20302 = ~n35847 ;
  assign y20303 = ~1'b0 ;
  assign y20304 = ~n35849 ;
  assign y20305 = ~1'b0 ;
  assign y20306 = n35850 ;
  assign y20307 = ~n28724 ;
  assign y20308 = ~1'b0 ;
  assign y20309 = ~n35852 ;
  assign y20310 = n21663 ;
  assign y20311 = n35855 ;
  assign y20312 = n35863 ;
  assign y20313 = ~n35866 ;
  assign y20314 = ~n35868 ;
  assign y20315 = ~1'b0 ;
  assign y20316 = ~1'b0 ;
  assign y20317 = n35869 ;
  assign y20318 = ~n35872 ;
  assign y20319 = ~1'b0 ;
  assign y20320 = ~1'b0 ;
  assign y20321 = n18246 ;
  assign y20322 = ~1'b0 ;
  assign y20323 = ~n31951 ;
  assign y20324 = ~1'b0 ;
  assign y20325 = ~n20458 ;
  assign y20326 = ~n35877 ;
  assign y20327 = n35879 ;
  assign y20328 = n35881 ;
  assign y20329 = ~1'b0 ;
  assign y20330 = ~1'b0 ;
  assign y20331 = ~1'b0 ;
  assign y20332 = n35882 ;
  assign y20333 = n35883 ;
  assign y20334 = ~n35893 ;
  assign y20335 = n35901 ;
  assign y20336 = ~1'b0 ;
  assign y20337 = ~1'b0 ;
  assign y20338 = 1'b0 ;
  assign y20339 = ~n35902 ;
  assign y20340 = ~n35903 ;
  assign y20341 = ~1'b0 ;
  assign y20342 = ~n35906 ;
  assign y20343 = ~1'b0 ;
  assign y20344 = ~n35914 ;
  assign y20345 = ~n35916 ;
  assign y20346 = n35919 ;
  assign y20347 = ~1'b0 ;
  assign y20348 = n35924 ;
  assign y20349 = ~n35927 ;
  assign y20350 = ~n35929 ;
  assign y20351 = 1'b0 ;
  assign y20352 = ~1'b0 ;
  assign y20353 = ~1'b0 ;
  assign y20354 = ~n226 ;
  assign y20355 = n35933 ;
  assign y20356 = ~n35934 ;
  assign y20357 = ~1'b0 ;
  assign y20358 = ~n35941 ;
  assign y20359 = n35942 ;
  assign y20360 = ~n35947 ;
  assign y20361 = ~n35948 ;
  assign y20362 = ~n35950 ;
  assign y20363 = ~1'b0 ;
  assign y20364 = ~n35951 ;
  assign y20365 = ~1'b0 ;
  assign y20366 = n35954 ;
  assign y20367 = 1'b0 ;
  assign y20368 = ~n35957 ;
  assign y20369 = n35961 ;
  assign y20370 = n35964 ;
  assign y20371 = ~n35965 ;
  assign y20372 = ~1'b0 ;
  assign y20373 = ~1'b0 ;
  assign y20374 = n35973 ;
  assign y20375 = n29338 ;
  assign y20376 = ~1'b0 ;
  assign y20377 = n35975 ;
  assign y20378 = ~1'b0 ;
  assign y20379 = n35976 ;
  assign y20380 = n35980 ;
  assign y20381 = ~1'b0 ;
  assign y20382 = ~1'b0 ;
  assign y20383 = ~1'b0 ;
  assign y20384 = ~n30374 ;
  assign y20385 = n35981 ;
  assign y20386 = ~1'b0 ;
  assign y20387 = ~n35987 ;
  assign y20388 = ~1'b0 ;
  assign y20389 = ~1'b0 ;
  assign y20390 = ~n35992 ;
  assign y20391 = ~1'b0 ;
  assign y20392 = n35994 ;
  assign y20393 = n35995 ;
  assign y20394 = ~1'b0 ;
  assign y20395 = n35998 ;
  assign y20396 = ~n36004 ;
  assign y20397 = ~n36005 ;
  assign y20398 = ~n36006 ;
  assign y20399 = n36007 ;
  assign y20400 = 1'b0 ;
  assign y20401 = ~1'b0 ;
  assign y20402 = n36009 ;
  assign y20403 = 1'b0 ;
  assign y20404 = n36011 ;
  assign y20405 = ~1'b0 ;
  assign y20406 = ~n36016 ;
  assign y20407 = n36019 ;
  assign y20408 = n36021 ;
  assign y20409 = ~n36032 ;
  assign y20410 = ~1'b0 ;
  assign y20411 = ~1'b0 ;
  assign y20412 = 1'b0 ;
  assign y20413 = ~n36038 ;
  assign y20414 = ~n36039 ;
  assign y20415 = n36043 ;
  assign y20416 = n36044 ;
  assign y20417 = n36045 ;
  assign y20418 = ~n36048 ;
  assign y20419 = ~1'b0 ;
  assign y20420 = ~n36050 ;
  assign y20421 = ~1'b0 ;
  assign y20422 = ~n34450 ;
  assign y20423 = n36053 ;
  assign y20424 = n36056 ;
  assign y20425 = ~1'b0 ;
  assign y20426 = ~n36063 ;
  assign y20427 = ~1'b0 ;
  assign y20428 = ~n36066 ;
  assign y20429 = ~n36068 ;
  assign y20430 = n36071 ;
  assign y20431 = n36073 ;
  assign y20432 = ~n36074 ;
  assign y20433 = 1'b0 ;
  assign y20434 = ~n36075 ;
  assign y20435 = ~1'b0 ;
  assign y20436 = n36077 ;
  assign y20437 = ~n36080 ;
  assign y20438 = n36082 ;
  assign y20439 = ~n36083 ;
  assign y20440 = ~1'b0 ;
  assign y20441 = n4216 ;
  assign y20442 = n36084 ;
  assign y20443 = ~n36087 ;
  assign y20444 = n36093 ;
  assign y20445 = ~n36095 ;
  assign y20446 = n10153 ;
  assign y20447 = ~n36100 ;
  assign y20448 = n36101 ;
  assign y20449 = ~n26888 ;
  assign y20450 = ~1'b0 ;
  assign y20451 = ~1'b0 ;
  assign y20452 = ~1'b0 ;
  assign y20453 = ~n36102 ;
  assign y20454 = ~1'b0 ;
  assign y20455 = ~n36103 ;
  assign y20456 = n36104 ;
  assign y20457 = ~1'b0 ;
  assign y20458 = ~n36106 ;
  assign y20459 = ~1'b0 ;
  assign y20460 = ~n20740 ;
  assign y20461 = ~n36107 ;
  assign y20462 = ~n36110 ;
  assign y20463 = ~n36113 ;
  assign y20464 = ~n36118 ;
  assign y20465 = n36120 ;
  assign y20466 = ~1'b0 ;
  assign y20467 = ~n36124 ;
  assign y20468 = ~1'b0 ;
  assign y20469 = n36128 ;
  assign y20470 = n36131 ;
  assign y20471 = ~n36136 ;
  assign y20472 = n28699 ;
  assign y20473 = n36139 ;
  assign y20474 = ~1'b0 ;
  assign y20475 = ~1'b0 ;
  assign y20476 = n36141 ;
  assign y20477 = n23033 ;
  assign y20478 = ~1'b0 ;
  assign y20479 = ~n36142 ;
  assign y20480 = ~n36143 ;
  assign y20481 = ~n36147 ;
  assign y20482 = n36149 ;
  assign y20483 = n36152 ;
  assign y20484 = ~1'b0 ;
  assign y20485 = ~n36155 ;
  assign y20486 = n36164 ;
  assign y20487 = ~n36166 ;
  assign y20488 = ~n36167 ;
  assign y20489 = n14385 ;
  assign y20490 = 1'b0 ;
  assign y20491 = n36170 ;
  assign y20492 = ~n36180 ;
  assign y20493 = n36181 ;
  assign y20494 = n36185 ;
  assign y20495 = n36187 ;
  assign y20496 = ~n36189 ;
  assign y20497 = ~1'b0 ;
  assign y20498 = ~1'b0 ;
  assign y20499 = ~n36191 ;
  assign y20500 = ~n36194 ;
  assign y20501 = n36196 ;
  assign y20502 = ~1'b0 ;
  assign y20503 = ~n10330 ;
  assign y20504 = ~1'b0 ;
  assign y20505 = n36200 ;
  assign y20506 = ~1'b0 ;
  assign y20507 = n36203 ;
  assign y20508 = n36205 ;
  assign y20509 = ~n36207 ;
  assign y20510 = n36210 ;
  assign y20511 = ~1'b0 ;
  assign y20512 = ~1'b0 ;
  assign y20513 = n36212 ;
  assign y20514 = ~n36213 ;
  assign y20515 = n36214 ;
  assign y20516 = ~1'b0 ;
  assign y20517 = ~1'b0 ;
  assign y20518 = ~n36218 ;
  assign y20519 = ~n36221 ;
  assign y20520 = n36225 ;
  assign y20521 = ~n36227 ;
  assign y20522 = ~1'b0 ;
  assign y20523 = n36228 ;
  assign y20524 = ~n36230 ;
  assign y20525 = ~n36231 ;
  assign y20526 = ~1'b0 ;
  assign y20527 = n36233 ;
  assign y20528 = ~1'b0 ;
  assign y20529 = ~1'b0 ;
  assign y20530 = n22712 ;
  assign y20531 = ~1'b0 ;
  assign y20532 = ~n36234 ;
  assign y20533 = ~n36238 ;
  assign y20534 = ~n36240 ;
  assign y20535 = ~n36242 ;
  assign y20536 = ~n36243 ;
  assign y20537 = n26060 ;
  assign y20538 = ~n36246 ;
  assign y20539 = ~1'b0 ;
  assign y20540 = ~1'b0 ;
  assign y20541 = ~1'b0 ;
  assign y20542 = n36248 ;
  assign y20543 = ~1'b0 ;
  assign y20544 = ~1'b0 ;
  assign y20545 = n36251 ;
  assign y20546 = ~1'b0 ;
  assign y20547 = ~n36275 ;
  assign y20548 = n36277 ;
  assign y20549 = ~n36281 ;
  assign y20550 = n36283 ;
  assign y20551 = ~n25281 ;
  assign y20552 = ~1'b0 ;
  assign y20553 = n36284 ;
  assign y20554 = n36285 ;
  assign y20555 = 1'b0 ;
  assign y20556 = ~1'b0 ;
  assign y20557 = n36287 ;
  assign y20558 = ~1'b0 ;
  assign y20559 = n36289 ;
  assign y20560 = ~1'b0 ;
  assign y20561 = ~n36291 ;
  assign y20562 = ~n36294 ;
  assign y20563 = ~n36299 ;
  assign y20564 = ~1'b0 ;
  assign y20565 = ~1'b0 ;
  assign y20566 = n36304 ;
  assign y20567 = ~1'b0 ;
  assign y20568 = ~n36306 ;
  assign y20569 = n36308 ;
  assign y20570 = n36309 ;
  assign y20571 = ~1'b0 ;
  assign y20572 = ~1'b0 ;
  assign y20573 = ~n36310 ;
  assign y20574 = ~1'b0 ;
  assign y20575 = n36311 ;
  assign y20576 = ~n36313 ;
  assign y20577 = n36316 ;
  assign y20578 = ~n36318 ;
  assign y20579 = ~1'b0 ;
  assign y20580 = ~n36321 ;
  assign y20581 = ~1'b0 ;
  assign y20582 = ~n36322 ;
  assign y20583 = ~n36323 ;
  assign y20584 = ~n36325 ;
  assign y20585 = n36329 ;
  assign y20586 = n36331 ;
  assign y20587 = n36332 ;
  assign y20588 = ~n36336 ;
  assign y20589 = n24986 ;
  assign y20590 = n36338 ;
  assign y20591 = ~1'b0 ;
  assign y20592 = n36340 ;
  assign y20593 = n36343 ;
  assign y20594 = n36344 ;
  assign y20595 = ~n36346 ;
  assign y20596 = ~1'b0 ;
  assign y20597 = ~1'b0 ;
  assign y20598 = n5077 ;
  assign y20599 = ~1'b0 ;
  assign y20600 = ~n33869 ;
  assign y20601 = n36348 ;
  assign y20602 = n36350 ;
  assign y20603 = ~n36354 ;
  assign y20604 = ~n17329 ;
  assign y20605 = n15829 ;
  assign y20606 = n36355 ;
  assign y20607 = ~1'b0 ;
  assign y20608 = ~1'b0 ;
  assign y20609 = ~1'b0 ;
  assign y20610 = ~n36359 ;
  assign y20611 = ~n36360 ;
  assign y20612 = ~n36364 ;
  assign y20613 = ~1'b0 ;
  assign y20614 = n36365 ;
  assign y20615 = n36366 ;
  assign y20616 = n36368 ;
  assign y20617 = ~1'b0 ;
  assign y20618 = n15581 ;
  assign y20619 = ~1'b0 ;
  assign y20620 = ~1'b0 ;
  assign y20621 = ~1'b0 ;
  assign y20622 = ~n36369 ;
  assign y20623 = n36370 ;
  assign y20624 = ~n36371 ;
  assign y20625 = n36373 ;
  assign y20626 = ~1'b0 ;
  assign y20627 = n25340 ;
  assign y20628 = ~n36375 ;
  assign y20629 = n36376 ;
  assign y20630 = ~1'b0 ;
  assign y20631 = ~n36381 ;
  assign y20632 = 1'b0 ;
  assign y20633 = ~n36383 ;
  assign y20634 = ~n36387 ;
  assign y20635 = ~1'b0 ;
  assign y20636 = n36390 ;
  assign y20637 = ~1'b0 ;
  assign y20638 = ~n36392 ;
  assign y20639 = ~1'b0 ;
  assign y20640 = ~n36395 ;
  assign y20641 = ~n36400 ;
  assign y20642 = ~1'b0 ;
  assign y20643 = n36409 ;
  assign y20644 = ~1'b0 ;
  assign y20645 = ~1'b0 ;
  assign y20646 = ~n36411 ;
  assign y20647 = ~1'b0 ;
  assign y20648 = ~n36415 ;
  assign y20649 = n36417 ;
  assign y20650 = ~1'b0 ;
  assign y20651 = ~n36419 ;
  assign y20652 = ~1'b0 ;
  assign y20653 = ~n36422 ;
  assign y20654 = ~n36424 ;
  assign y20655 = ~1'b0 ;
  assign y20656 = n36425 ;
  assign y20657 = n36427 ;
  assign y20658 = ~n36428 ;
  assign y20659 = ~n36429 ;
  assign y20660 = ~1'b0 ;
  assign y20661 = ~1'b0 ;
  assign y20662 = n33196 ;
  assign y20663 = n36432 ;
  assign y20664 = ~1'b0 ;
  assign y20665 = n36445 ;
  assign y20666 = n36446 ;
  assign y20667 = ~1'b0 ;
  assign y20668 = n25598 ;
  assign y20669 = n36447 ;
  assign y20670 = ~1'b0 ;
  assign y20671 = n36449 ;
  assign y20672 = n36451 ;
  assign y20673 = n36452 ;
  assign y20674 = ~1'b0 ;
  assign y20675 = ~n36457 ;
  assign y20676 = ~1'b0 ;
  assign y20677 = ~1'b0 ;
  assign y20678 = ~n36459 ;
  assign y20679 = ~n36462 ;
  assign y20680 = ~n36466 ;
  assign y20681 = n4801 ;
  assign y20682 = n36471 ;
  assign y20683 = n36473 ;
  assign y20684 = n36478 ;
  assign y20685 = ~n11302 ;
  assign y20686 = n36481 ;
  assign y20687 = ~n36482 ;
  assign y20688 = n36484 ;
  assign y20689 = n36490 ;
  assign y20690 = ~n36491 ;
  assign y20691 = ~1'b0 ;
  assign y20692 = n10719 ;
  assign y20693 = ~n30608 ;
  assign y20694 = ~n36494 ;
  assign y20695 = ~n36495 ;
  assign y20696 = ~n36496 ;
  assign y20697 = ~n36497 ;
  assign y20698 = ~1'b0 ;
  assign y20699 = n36498 ;
  assign y20700 = ~n36499 ;
  assign y20701 = ~1'b0 ;
  assign y20702 = ~n36502 ;
  assign y20703 = ~1'b0 ;
  assign y20704 = ~n36506 ;
  assign y20705 = n36509 ;
  assign y20706 = ~1'b0 ;
  assign y20707 = ~1'b0 ;
  assign y20708 = n36511 ;
  assign y20709 = ~1'b0 ;
  assign y20710 = ~1'b0 ;
  assign y20711 = ~n36512 ;
  assign y20712 = ~n36514 ;
  assign y20713 = ~n36516 ;
  assign y20714 = n36519 ;
  assign y20715 = ~1'b0 ;
  assign y20716 = ~1'b0 ;
  assign y20717 = n36520 ;
  assign y20718 = ~n36521 ;
  assign y20719 = ~1'b0 ;
  assign y20720 = ~n36522 ;
  assign y20721 = n36525 ;
  assign y20722 = ~1'b0 ;
  assign y20723 = ~1'b0 ;
  assign y20724 = ~1'b0 ;
  assign y20725 = ~1'b0 ;
  assign y20726 = ~n17702 ;
  assign y20727 = ~n36529 ;
  assign y20728 = ~1'b0 ;
  assign y20729 = ~n36533 ;
  assign y20730 = n36536 ;
  assign y20731 = ~1'b0 ;
  assign y20732 = n29074 ;
  assign y20733 = ~1'b0 ;
  assign y20734 = ~1'b0 ;
  assign y20735 = n36537 ;
  assign y20736 = n36538 ;
  assign y20737 = ~1'b0 ;
  assign y20738 = ~n36539 ;
  assign y20739 = ~1'b0 ;
  assign y20740 = ~1'b0 ;
  assign y20741 = n36541 ;
  assign y20742 = ~n36546 ;
  assign y20743 = ~n36547 ;
  assign y20744 = n36550 ;
  assign y20745 = 1'b0 ;
  assign y20746 = ~1'b0 ;
  assign y20747 = ~1'b0 ;
  assign y20748 = ~1'b0 ;
  assign y20749 = n36552 ;
  assign y20750 = ~n36555 ;
  assign y20751 = ~1'b0 ;
  assign y20752 = 1'b0 ;
  assign y20753 = ~1'b0 ;
  assign y20754 = ~n36556 ;
  assign y20755 = n36557 ;
  assign y20756 = ~n36562 ;
  assign y20757 = ~n16809 ;
  assign y20758 = n36564 ;
  assign y20759 = n36567 ;
  assign y20760 = ~n36571 ;
  assign y20761 = ~n31290 ;
  assign y20762 = ~n36572 ;
  assign y20763 = ~1'b0 ;
  assign y20764 = ~n36576 ;
  assign y20765 = n36577 ;
  assign y20766 = ~n36579 ;
  assign y20767 = ~1'b0 ;
  assign y20768 = ~1'b0 ;
  assign y20769 = ~1'b0 ;
  assign y20770 = ~1'b0 ;
  assign y20771 = ~n36580 ;
  assign y20772 = ~n36581 ;
  assign y20773 = ~n36582 ;
  assign y20774 = n36583 ;
  assign y20775 = ~n36585 ;
  assign y20776 = ~1'b0 ;
  assign y20777 = ~n36588 ;
  assign y20778 = n36591 ;
  assign y20779 = ~n36594 ;
  assign y20780 = 1'b0 ;
  assign y20781 = ~1'b0 ;
  assign y20782 = ~1'b0 ;
  assign y20783 = ~n36596 ;
  assign y20784 = n36597 ;
  assign y20785 = n36598 ;
  assign y20786 = ~n36599 ;
  assign y20787 = n36600 ;
  assign y20788 = ~n36605 ;
  assign y20789 = ~1'b0 ;
  assign y20790 = ~n36607 ;
  assign y20791 = n20349 ;
  assign y20792 = n36610 ;
  assign y20793 = ~1'b0 ;
  assign y20794 = n36613 ;
  assign y20795 = ~n36615 ;
  assign y20796 = ~n36622 ;
  assign y20797 = n36623 ;
  assign y20798 = ~1'b0 ;
  assign y20799 = n36627 ;
  assign y20800 = ~n36628 ;
  assign y20801 = n12528 ;
  assign y20802 = ~1'b0 ;
  assign y20803 = ~1'b0 ;
  assign y20804 = ~n36630 ;
  assign y20805 = ~1'b0 ;
  assign y20806 = ~n36635 ;
  assign y20807 = n36640 ;
  assign y20808 = ~1'b0 ;
  assign y20809 = ~1'b0 ;
  assign y20810 = ~n36645 ;
  assign y20811 = ~1'b0 ;
  assign y20812 = n36646 ;
  assign y20813 = n36648 ;
  assign y20814 = ~1'b0 ;
  assign y20815 = n36653 ;
  assign y20816 = n36654 ;
  assign y20817 = ~1'b0 ;
  assign y20818 = 1'b0 ;
  assign y20819 = ~n36656 ;
  assign y20820 = ~1'b0 ;
  assign y20821 = ~1'b0 ;
  assign y20822 = ~n36661 ;
  assign y20823 = n36664 ;
  assign y20824 = ~1'b0 ;
  assign y20825 = ~1'b0 ;
  assign y20826 = ~n36668 ;
  assign y20827 = ~n36671 ;
  assign y20828 = ~1'b0 ;
  assign y20829 = n36673 ;
  assign y20830 = ~1'b0 ;
  assign y20831 = n36674 ;
  assign y20832 = ~1'b0 ;
  assign y20833 = ~n36678 ;
  assign y20834 = ~1'b0 ;
  assign y20835 = ~n36680 ;
  assign y20836 = ~n36684 ;
  assign y20837 = n36685 ;
  assign y20838 = ~n36689 ;
  assign y20839 = ~n36690 ;
  assign y20840 = n2391 ;
  assign y20841 = ~n36691 ;
  assign y20842 = ~1'b0 ;
  assign y20843 = n36695 ;
  assign y20844 = n36697 ;
  assign y20845 = ~n36699 ;
  assign y20846 = n36704 ;
  assign y20847 = ~n36711 ;
  assign y20848 = ~1'b0 ;
  assign y20849 = ~1'b0 ;
  assign y20850 = 1'b0 ;
  assign y20851 = ~n36714 ;
  assign y20852 = ~n36716 ;
  assign y20853 = n36718 ;
  assign y20854 = n36723 ;
  assign y20855 = n36726 ;
  assign y20856 = ~1'b0 ;
  assign y20857 = n36728 ;
  assign y20858 = n36729 ;
  assign y20859 = ~1'b0 ;
  assign y20860 = ~n36730 ;
  assign y20861 = ~n25476 ;
  assign y20862 = n36734 ;
  assign y20863 = ~1'b0 ;
  assign y20864 = 1'b0 ;
  assign y20865 = n36737 ;
  assign y20866 = ~n36740 ;
  assign y20867 = ~1'b0 ;
  assign y20868 = ~n8242 ;
  assign y20869 = n36741 ;
  assign y20870 = ~1'b0 ;
  assign y20871 = n36742 ;
  assign y20872 = n36744 ;
  assign y20873 = ~n36745 ;
  assign y20874 = ~1'b0 ;
  assign y20875 = ~1'b0 ;
  assign y20876 = ~n36746 ;
  assign y20877 = n36748 ;
  assign y20878 = n3924 ;
  assign y20879 = n36751 ;
  assign y20880 = ~n36753 ;
  assign y20881 = 1'b0 ;
  assign y20882 = n36755 ;
  assign y20883 = n36756 ;
  assign y20884 = n6133 ;
  assign y20885 = ~n36759 ;
  assign y20886 = n10376 ;
  assign y20887 = ~1'b0 ;
  assign y20888 = ~n7824 ;
  assign y20889 = ~n17434 ;
  assign y20890 = ~n36760 ;
  assign y20891 = ~1'b0 ;
  assign y20892 = n36764 ;
  assign y20893 = ~n36765 ;
  assign y20894 = ~n36767 ;
  assign y20895 = ~n36770 ;
  assign y20896 = ~n36773 ;
  assign y20897 = n36776 ;
  assign y20898 = ~1'b0 ;
  assign y20899 = n36778 ;
  assign y20900 = ~n36780 ;
  assign y20901 = n36784 ;
  assign y20902 = ~n36785 ;
  assign y20903 = ~n36786 ;
  assign y20904 = n36787 ;
  assign y20905 = ~n36788 ;
  assign y20906 = n36789 ;
  assign y20907 = ~1'b0 ;
  assign y20908 = ~n36793 ;
  assign y20909 = ~n19626 ;
  assign y20910 = n36795 ;
  assign y20911 = ~n36798 ;
  assign y20912 = ~n36802 ;
  assign y20913 = ~1'b0 ;
  assign y20914 = ~n36803 ;
  assign y20915 = ~n36806 ;
  assign y20916 = n36809 ;
  assign y20917 = ~1'b0 ;
  assign y20918 = ~1'b0 ;
  assign y20919 = ~n36815 ;
  assign y20920 = ~n7111 ;
  assign y20921 = n34357 ;
  assign y20922 = n36817 ;
  assign y20923 = n36818 ;
  assign y20924 = n36821 ;
  assign y20925 = n36823 ;
  assign y20926 = n19045 ;
  assign y20927 = ~n36825 ;
  assign y20928 = ~n36830 ;
  assign y20929 = ~n36834 ;
  assign y20930 = ~1'b0 ;
  assign y20931 = 1'b0 ;
  assign y20932 = n36836 ;
  assign y20933 = ~n36838 ;
  assign y20934 = n36839 ;
  assign y20935 = ~n36840 ;
  assign y20936 = n27586 ;
  assign y20937 = ~n36842 ;
  assign y20938 = n36844 ;
  assign y20939 = ~n36846 ;
  assign y20940 = n36848 ;
  assign y20941 = n36849 ;
  assign y20942 = ~n36851 ;
  assign y20943 = ~n36854 ;
  assign y20944 = n36856 ;
  assign y20945 = ~n36861 ;
  assign y20946 = ~n36864 ;
  assign y20947 = n36866 ;
  assign y20948 = n36868 ;
  assign y20949 = ~1'b0 ;
  assign y20950 = n36870 ;
  assign y20951 = ~1'b0 ;
  assign y20952 = ~n36874 ;
  assign y20953 = ~1'b0 ;
  assign y20954 = ~n36875 ;
  assign y20955 = ~n36877 ;
  assign y20956 = n36880 ;
  assign y20957 = ~1'b0 ;
  assign y20958 = ~n36886 ;
  assign y20959 = ~1'b0 ;
  assign y20960 = ~n36887 ;
  assign y20961 = n36891 ;
  assign y20962 = n36892 ;
  assign y20963 = n36895 ;
  assign y20964 = 1'b0 ;
  assign y20965 = n35444 ;
  assign y20966 = ~1'b0 ;
  assign y20967 = ~1'b0 ;
  assign y20968 = ~n36899 ;
  assign y20969 = ~1'b0 ;
  assign y20970 = ~n36901 ;
  assign y20971 = n36906 ;
  assign y20972 = 1'b0 ;
  assign y20973 = ~1'b0 ;
  assign y20974 = n36913 ;
  assign y20975 = n36918 ;
  assign y20976 = ~1'b0 ;
  assign y20977 = ~n7010 ;
  assign y20978 = ~n36921 ;
  assign y20979 = n3384 ;
  assign y20980 = ~n2363 ;
  assign y20981 = ~n36922 ;
  assign y20982 = ~n36925 ;
  assign y20983 = ~n36929 ;
  assign y20984 = n36931 ;
  assign y20985 = n36932 ;
  assign y20986 = n36935 ;
  assign y20987 = ~n36936 ;
  assign y20988 = n36939 ;
  assign y20989 = n36940 ;
  assign y20990 = ~n36941 ;
  assign y20991 = ~1'b0 ;
  assign y20992 = ~n6396 ;
  assign y20993 = n36942 ;
  assign y20994 = n36945 ;
  assign y20995 = n36965 ;
  assign y20996 = ~n36970 ;
  assign y20997 = 1'b0 ;
  assign y20998 = n36971 ;
  assign y20999 = ~n36974 ;
  assign y21000 = n36979 ;
  assign y21001 = ~n36980 ;
  assign y21002 = ~1'b0 ;
  assign y21003 = ~n36981 ;
  assign y21004 = n36983 ;
  assign y21005 = ~1'b0 ;
  assign y21006 = 1'b0 ;
  assign y21007 = n8827 ;
  assign y21008 = ~1'b0 ;
  assign y21009 = ~1'b0 ;
  assign y21010 = ~1'b0 ;
  assign y21011 = n36994 ;
  assign y21012 = ~1'b0 ;
  assign y21013 = ~1'b0 ;
  assign y21014 = ~1'b0 ;
  assign y21015 = ~n36998 ;
  assign y21016 = n37002 ;
  assign y21017 = ~n37003 ;
  assign y21018 = ~n37010 ;
  assign y21019 = n37012 ;
  assign y21020 = ~n37015 ;
  assign y21021 = ~1'b0 ;
  assign y21022 = ~1'b0 ;
  assign y21023 = ~n37017 ;
  assign y21024 = ~1'b0 ;
  assign y21025 = ~1'b0 ;
  assign y21026 = ~1'b0 ;
  assign y21027 = n37022 ;
  assign y21028 = ~n37024 ;
  assign y21029 = ~n37025 ;
  assign y21030 = ~1'b0 ;
  assign y21031 = ~n37028 ;
  assign y21032 = ~n37029 ;
  assign y21033 = ~n37032 ;
  assign y21034 = n37033 ;
  assign y21035 = n37035 ;
  assign y21036 = ~1'b0 ;
  assign y21037 = ~n37040 ;
  assign y21038 = ~n37042 ;
  assign y21039 = ~n37043 ;
  assign y21040 = n18941 ;
  assign y21041 = n37045 ;
  assign y21042 = n2131 ;
  assign y21043 = ~1'b0 ;
  assign y21044 = ~1'b0 ;
  assign y21045 = ~1'b0 ;
  assign y21046 = ~n37051 ;
  assign y21047 = n37054 ;
  assign y21048 = n37056 ;
  assign y21049 = ~n37057 ;
  assign y21050 = ~n37058 ;
  assign y21051 = n37062 ;
  assign y21052 = n37063 ;
  assign y21053 = n15166 ;
  assign y21054 = ~1'b0 ;
  assign y21055 = ~1'b0 ;
  assign y21056 = ~n37065 ;
  assign y21057 = ~n37067 ;
  assign y21058 = n37070 ;
  assign y21059 = ~1'b0 ;
  assign y21060 = n1700 ;
  assign y21061 = ~n37072 ;
  assign y21062 = 1'b0 ;
  assign y21063 = ~1'b0 ;
  assign y21064 = ~1'b0 ;
  assign y21065 = ~1'b0 ;
  assign y21066 = n12541 ;
  assign y21067 = ~1'b0 ;
  assign y21068 = ~n37076 ;
  assign y21069 = n37077 ;
  assign y21070 = ~n37080 ;
  assign y21071 = ~1'b0 ;
  assign y21072 = ~1'b0 ;
  assign y21073 = ~n37082 ;
  assign y21074 = n37085 ;
  assign y21075 = ~n37087 ;
  assign y21076 = 1'b0 ;
  assign y21077 = n37090 ;
  assign y21078 = ~n37092 ;
  assign y21079 = ~n37093 ;
  assign y21080 = ~1'b0 ;
  assign y21081 = n37094 ;
  assign y21082 = ~n37096 ;
  assign y21083 = n37103 ;
  assign y21084 = ~n927 ;
  assign y21085 = n37104 ;
  assign y21086 = ~n23707 ;
  assign y21087 = n37106 ;
  assign y21088 = n37108 ;
  assign y21089 = ~1'b0 ;
  assign y21090 = n37111 ;
  assign y21091 = n37112 ;
  assign y21092 = n15736 ;
  assign y21093 = ~n37113 ;
  assign y21094 = ~n37117 ;
  assign y21095 = n37126 ;
  assign y21096 = ~n37129 ;
  assign y21097 = n37131 ;
  assign y21098 = n37133 ;
  assign y21099 = ~n37134 ;
  assign y21100 = ~n37136 ;
  assign y21101 = ~1'b0 ;
  assign y21102 = ~n37138 ;
  assign y21103 = n37144 ;
  assign y21104 = 1'b0 ;
  assign y21105 = n20138 ;
  assign y21106 = ~n37146 ;
  assign y21107 = n37147 ;
  assign y21108 = n37148 ;
  assign y21109 = n9453 ;
  assign y21110 = ~1'b0 ;
  assign y21111 = ~1'b0 ;
  assign y21112 = ~n37151 ;
  assign y21113 = ~1'b0 ;
  assign y21114 = n37153 ;
  assign y21115 = n37154 ;
  assign y21116 = n37155 ;
  assign y21117 = n37157 ;
  assign y21118 = ~n37158 ;
  assign y21119 = n37159 ;
  assign y21120 = ~n37162 ;
  assign y21121 = ~n37163 ;
  assign y21122 = ~1'b0 ;
  assign y21123 = ~n37167 ;
  assign y21124 = n37168 ;
  assign y21125 = n37171 ;
  assign y21126 = ~1'b0 ;
  assign y21127 = n37173 ;
  assign y21128 = ~n32449 ;
  assign y21129 = n37175 ;
  assign y21130 = ~1'b0 ;
  assign y21131 = n37176 ;
  assign y21132 = n24923 ;
  assign y21133 = ~1'b0 ;
  assign y21134 = ~n37178 ;
  assign y21135 = n18653 ;
  assign y21136 = n37181 ;
  assign y21137 = 1'b0 ;
  assign y21138 = ~n7063 ;
  assign y21139 = n37182 ;
  assign y21140 = n37184 ;
  assign y21141 = n37185 ;
  assign y21142 = ~n37187 ;
  assign y21143 = n37189 ;
  assign y21144 = ~n37195 ;
  assign y21145 = n37201 ;
  assign y21146 = ~1'b0 ;
  assign y21147 = ~n37202 ;
  assign y21148 = ~n37203 ;
  assign y21149 = ~n37204 ;
  assign y21150 = ~1'b0 ;
  assign y21151 = ~n19480 ;
  assign y21152 = ~n37205 ;
  assign y21153 = ~n37206 ;
  assign y21154 = ~n37207 ;
  assign y21155 = ~1'b0 ;
  assign y21156 = 1'b0 ;
  assign y21157 = ~1'b0 ;
  assign y21158 = ~n37209 ;
  assign y21159 = 1'b0 ;
  assign y21160 = ~1'b0 ;
  assign y21161 = ~n15538 ;
  assign y21162 = ~1'b0 ;
  assign y21163 = n37211 ;
  assign y21164 = ~n37214 ;
  assign y21165 = ~n37220 ;
  assign y21166 = ~1'b0 ;
  assign y21167 = ~n37221 ;
  assign y21168 = ~n37224 ;
  assign y21169 = n37229 ;
  assign y21170 = n37233 ;
  assign y21171 = ~n37235 ;
  assign y21172 = ~1'b0 ;
  assign y21173 = ~1'b0 ;
  assign y21174 = ~1'b0 ;
  assign y21175 = ~1'b0 ;
  assign y21176 = ~1'b0 ;
  assign y21177 = ~n37236 ;
  assign y21178 = ~n37238 ;
  assign y21179 = ~1'b0 ;
  assign y21180 = ~1'b0 ;
  assign y21181 = n37241 ;
  assign y21182 = ~1'b0 ;
  assign y21183 = ~n37243 ;
  assign y21184 = ~1'b0 ;
  assign y21185 = ~n37244 ;
  assign y21186 = n37247 ;
  assign y21187 = ~1'b0 ;
  assign y21188 = ~n37250 ;
  assign y21189 = n37252 ;
  assign y21190 = ~n37257 ;
  assign y21191 = ~n37260 ;
  assign y21192 = ~n37263 ;
  assign y21193 = ~1'b0 ;
  assign y21194 = ~n37266 ;
  assign y21195 = ~1'b0 ;
  assign y21196 = 1'b0 ;
  assign y21197 = n37272 ;
  assign y21198 = n37274 ;
  assign y21199 = ~1'b0 ;
  assign y21200 = ~n37280 ;
  assign y21201 = ~1'b0 ;
  assign y21202 = n37281 ;
  assign y21203 = n37284 ;
  assign y21204 = n37285 ;
  assign y21205 = ~1'b0 ;
  assign y21206 = ~n37289 ;
  assign y21207 = ~n37296 ;
  assign y21208 = n24755 ;
  assign y21209 = n37297 ;
  assign y21210 = ~n37298 ;
  assign y21211 = ~1'b0 ;
  assign y21212 = ~n37300 ;
  assign y21213 = n37302 ;
  assign y21214 = n22893 ;
  assign y21215 = ~n37304 ;
  assign y21216 = ~n2933 ;
  assign y21217 = n37308 ;
  assign y21218 = ~1'b0 ;
  assign y21219 = n37309 ;
  assign y21220 = ~n37311 ;
  assign y21221 = ~n37315 ;
  assign y21222 = ~1'b0 ;
  assign y21223 = ~1'b0 ;
  assign y21224 = 1'b0 ;
  assign y21225 = ~n37317 ;
  assign y21226 = ~n37319 ;
  assign y21227 = ~n37321 ;
  assign y21228 = n37323 ;
  assign y21229 = n37324 ;
  assign y21230 = ~n37325 ;
  assign y21231 = n37326 ;
  assign y21232 = ~n37328 ;
  assign y21233 = n37329 ;
  assign y21234 = n37332 ;
  assign y21235 = n37334 ;
  assign y21236 = n37336 ;
  assign y21237 = ~n37337 ;
  assign y21238 = ~n37338 ;
  assign y21239 = ~1'b0 ;
  assign y21240 = ~n37339 ;
  assign y21241 = n37340 ;
  assign y21242 = ~1'b0 ;
  assign y21243 = n37343 ;
  assign y21244 = ~1'b0 ;
  assign y21245 = ~n37344 ;
  assign y21246 = n37347 ;
  assign y21247 = n37350 ;
  assign y21248 = ~1'b0 ;
  assign y21249 = n37351 ;
  assign y21250 = n37352 ;
  assign y21251 = n37354 ;
  assign y21252 = ~1'b0 ;
  assign y21253 = n37355 ;
  assign y21254 = n24371 ;
  assign y21255 = n37356 ;
  assign y21256 = n37358 ;
  assign y21257 = n37359 ;
  assign y21258 = ~1'b0 ;
  assign y21259 = 1'b0 ;
  assign y21260 = n37361 ;
  assign y21261 = ~n37363 ;
  assign y21262 = ~n37364 ;
  assign y21263 = ~n37370 ;
  assign y21264 = n37372 ;
  assign y21265 = n37373 ;
  assign y21266 = ~1'b0 ;
  assign y21267 = ~1'b0 ;
  assign y21268 = n37378 ;
  assign y21269 = n37379 ;
  assign y21270 = n36797 ;
  assign y21271 = ~n37382 ;
  assign y21272 = n37383 ;
  assign y21273 = n37385 ;
  assign y21274 = ~n129 ;
  assign y21275 = ~n37387 ;
  assign y21276 = n37388 ;
  assign y21277 = ~1'b0 ;
  assign y21278 = ~n37391 ;
  assign y21279 = n24073 ;
  assign y21280 = n37392 ;
  assign y21281 = 1'b0 ;
  assign y21282 = ~1'b0 ;
  assign y21283 = n37395 ;
  assign y21284 = n37398 ;
  assign y21285 = n37399 ;
  assign y21286 = ~1'b0 ;
  assign y21287 = ~1'b0 ;
  assign y21288 = n37401 ;
  assign y21289 = ~1'b0 ;
  assign y21290 = n37403 ;
  assign y21291 = ~1'b0 ;
  assign y21292 = ~1'b0 ;
  assign y21293 = ~n2668 ;
  assign y21294 = ~n37405 ;
  assign y21295 = ~n37410 ;
  assign y21296 = ~n37412 ;
  assign y21297 = n37413 ;
  assign y21298 = ~n37415 ;
  assign y21299 = n37417 ;
  assign y21300 = ~n37420 ;
  assign y21301 = n37423 ;
  assign y21302 = n37425 ;
  assign y21303 = ~1'b0 ;
  assign y21304 = ~n37429 ;
  assign y21305 = ~n37439 ;
  assign y21306 = ~n37445 ;
  assign y21307 = ~1'b0 ;
  assign y21308 = ~1'b0 ;
  assign y21309 = ~n37447 ;
  assign y21310 = ~n37450 ;
  assign y21311 = ~n37451 ;
  assign y21312 = 1'b0 ;
  assign y21313 = n37452 ;
  assign y21314 = n37455 ;
  assign y21315 = ~n37460 ;
  assign y21316 = ~1'b0 ;
  assign y21317 = n2638 ;
  assign y21318 = ~n37461 ;
  assign y21319 = ~1'b0 ;
  assign y21320 = ~n21960 ;
  assign y21321 = n37464 ;
  assign y21322 = ~1'b0 ;
  assign y21323 = n37465 ;
  assign y21324 = ~1'b0 ;
  assign y21325 = ~n37466 ;
  assign y21326 = ~1'b0 ;
  assign y21327 = n37471 ;
  assign y21328 = ~1'b0 ;
  assign y21329 = ~1'b0 ;
  assign y21330 = ~n15319 ;
  assign y21331 = ~n37473 ;
  assign y21332 = n37475 ;
  assign y21333 = n37476 ;
  assign y21334 = ~1'b0 ;
  assign y21335 = ~1'b0 ;
  assign y21336 = n37477 ;
  assign y21337 = ~1'b0 ;
  assign y21338 = ~n37479 ;
  assign y21339 = ~1'b0 ;
  assign y21340 = n37482 ;
  assign y21341 = ~n37487 ;
  assign y21342 = ~n37490 ;
  assign y21343 = n37492 ;
  assign y21344 = ~1'b0 ;
  assign y21345 = n37493 ;
  assign y21346 = ~1'b0 ;
  assign y21347 = n37494 ;
  assign y21348 = ~n37499 ;
  assign y21349 = ~1'b0 ;
  assign y21350 = ~n19271 ;
  assign y21351 = ~n37501 ;
  assign y21352 = ~1'b0 ;
  assign y21353 = n1210 ;
  assign y21354 = n6709 ;
  assign y21355 = n37505 ;
  assign y21356 = n37506 ;
  assign y21357 = ~n37507 ;
  assign y21358 = n37508 ;
  assign y21359 = ~n37512 ;
  assign y21360 = ~n37513 ;
  assign y21361 = n37516 ;
  assign y21362 = ~1'b0 ;
  assign y21363 = n37517 ;
  assign y21364 = ~1'b0 ;
  assign y21365 = ~1'b0 ;
  assign y21366 = n37520 ;
  assign y21367 = ~n37524 ;
  assign y21368 = n37525 ;
  assign y21369 = ~1'b0 ;
  assign y21370 = n37528 ;
  assign y21371 = ~1'b0 ;
  assign y21372 = ~n37530 ;
  assign y21373 = n13013 ;
  assign y21374 = ~1'b0 ;
  assign y21375 = ~n37532 ;
  assign y21376 = ~1'b0 ;
  assign y21377 = ~n37533 ;
  assign y21378 = 1'b0 ;
  assign y21379 = ~n37534 ;
  assign y21380 = ~1'b0 ;
  assign y21381 = ~1'b0 ;
  assign y21382 = ~1'b0 ;
  assign y21383 = ~1'b0 ;
  assign y21384 = ~n37535 ;
  assign y21385 = ~n12550 ;
  assign y21386 = ~n37536 ;
  assign y21387 = ~1'b0 ;
  assign y21388 = n37540 ;
  assign y21389 = n37544 ;
  assign y21390 = ~1'b0 ;
  assign y21391 = ~1'b0 ;
  assign y21392 = n37547 ;
  assign y21393 = ~n37549 ;
  assign y21394 = ~n37551 ;
  assign y21395 = ~1'b0 ;
  assign y21396 = n37555 ;
  assign y21397 = n5114 ;
  assign y21398 = ~n37556 ;
  assign y21399 = ~n37557 ;
  assign y21400 = n37560 ;
  assign y21401 = n3246 ;
  assign y21402 = n2552 ;
  assign y21403 = n37563 ;
  assign y21404 = ~n37569 ;
  assign y21405 = ~n37572 ;
  assign y21406 = n37574 ;
  assign y21407 = n37579 ;
  assign y21408 = ~n37581 ;
  assign y21409 = ~1'b0 ;
  assign y21410 = ~n37583 ;
  assign y21411 = 1'b0 ;
  assign y21412 = ~n37586 ;
  assign y21413 = ~1'b0 ;
  assign y21414 = ~1'b0 ;
  assign y21415 = ~1'b0 ;
  assign y21416 = n37590 ;
  assign y21417 = n26604 ;
  assign y21418 = ~n37591 ;
  assign y21419 = n21241 ;
  assign y21420 = n37593 ;
  assign y21421 = n14276 ;
  assign y21422 = n37595 ;
  assign y21423 = ~1'b0 ;
  assign y21424 = ~1'b0 ;
  assign y21425 = ~1'b0 ;
  assign y21426 = ~n37596 ;
  assign y21427 = ~n37598 ;
  assign y21428 = n37599 ;
  assign y21429 = n30367 ;
  assign y21430 = ~1'b0 ;
  assign y21431 = ~n37600 ;
  assign y21432 = n37603 ;
  assign y21433 = ~n6084 ;
  assign y21434 = ~n37607 ;
  assign y21435 = ~n37610 ;
  assign y21436 = ~1'b0 ;
  assign y21437 = n37612 ;
  assign y21438 = ~1'b0 ;
  assign y21439 = ~n37615 ;
  assign y21440 = n34397 ;
  assign y21441 = ~1'b0 ;
  assign y21442 = ~n37617 ;
  assign y21443 = ~n37619 ;
  assign y21444 = 1'b0 ;
  assign y21445 = n37620 ;
  assign y21446 = ~1'b0 ;
  assign y21447 = 1'b0 ;
  assign y21448 = n37628 ;
  assign y21449 = ~n37630 ;
  assign y21450 = ~n37631 ;
  assign y21451 = ~1'b0 ;
  assign y21452 = ~n37634 ;
  assign y21453 = n37635 ;
  assign y21454 = n30659 ;
  assign y21455 = n37640 ;
  assign y21456 = ~1'b0 ;
  assign y21457 = 1'b0 ;
  assign y21458 = n37643 ;
  assign y21459 = ~1'b0 ;
  assign y21460 = n37645 ;
  assign y21461 = n37647 ;
  assign y21462 = 1'b0 ;
  assign y21463 = n37648 ;
  assign y21464 = ~1'b0 ;
  assign y21465 = n1416 ;
  assign y21466 = ~n37649 ;
  assign y21467 = ~1'b0 ;
  assign y21468 = 1'b0 ;
  assign y21469 = n37654 ;
  assign y21470 = ~1'b0 ;
  assign y21471 = ~n24261 ;
  assign y21472 = ~n37657 ;
  assign y21473 = ~n37659 ;
  assign y21474 = ~n37662 ;
  assign y21475 = ~n37669 ;
  assign y21476 = ~1'b0 ;
  assign y21477 = ~1'b0 ;
  assign y21478 = n37670 ;
  assign y21479 = ~n37674 ;
  assign y21480 = n37677 ;
  assign y21481 = 1'b0 ;
  assign y21482 = ~n37679 ;
  assign y21483 = ~n37687 ;
  assign y21484 = n37689 ;
  assign y21485 = 1'b0 ;
  assign y21486 = n37690 ;
  assign y21487 = n37696 ;
  assign y21488 = n35820 ;
  assign y21489 = ~1'b0 ;
  assign y21490 = ~n37703 ;
  assign y21491 = n37704 ;
  assign y21492 = ~n35389 ;
  assign y21493 = ~n37705 ;
  assign y21494 = ~n37707 ;
  assign y21495 = n37709 ;
  assign y21496 = n37711 ;
  assign y21497 = ~n20068 ;
  assign y21498 = n37712 ;
  assign y21499 = ~n37718 ;
  assign y21500 = n37719 ;
  assign y21501 = n32207 ;
  assign y21502 = ~1'b0 ;
  assign y21503 = ~1'b0 ;
  assign y21504 = n37723 ;
  assign y21505 = n12013 ;
  assign y21506 = n37730 ;
  assign y21507 = n37731 ;
  assign y21508 = ~1'b0 ;
  assign y21509 = n36812 ;
  assign y21510 = ~n37733 ;
  assign y21511 = ~n37736 ;
  assign y21512 = ~1'b0 ;
  assign y21513 = n37737 ;
  assign y21514 = ~n37738 ;
  assign y21515 = ~n37742 ;
  assign y21516 = n37744 ;
  assign y21517 = n37745 ;
  assign y21518 = n37749 ;
  assign y21519 = ~n34769 ;
  assign y21520 = n37751 ;
  assign y21521 = n37752 ;
  assign y21522 = n37755 ;
  assign y21523 = n37762 ;
  assign y21524 = n37765 ;
  assign y21525 = ~1'b0 ;
  assign y21526 = 1'b0 ;
  assign y21527 = ~1'b0 ;
  assign y21528 = ~n37771 ;
  assign y21529 = ~n11159 ;
  assign y21530 = ~1'b0 ;
  assign y21531 = n37775 ;
  assign y21532 = ~1'b0 ;
  assign y21533 = ~n37777 ;
  assign y21534 = n37780 ;
  assign y21535 = ~1'b0 ;
  assign y21536 = ~1'b0 ;
  assign y21537 = ~n37786 ;
  assign y21538 = n37787 ;
  assign y21539 = ~1'b0 ;
  assign y21540 = 1'b0 ;
  assign y21541 = ~n37789 ;
  assign y21542 = ~n37794 ;
  assign y21543 = ~1'b0 ;
  assign y21544 = n37796 ;
  assign y21545 = ~n37797 ;
  assign y21546 = n5410 ;
  assign y21547 = ~n37798 ;
  assign y21548 = ~1'b0 ;
  assign y21549 = n37801 ;
  assign y21550 = ~1'b0 ;
  assign y21551 = ~n37805 ;
  assign y21552 = ~n37807 ;
  assign y21553 = n37810 ;
  assign y21554 = ~n37812 ;
  assign y21555 = ~n37814 ;
  assign y21556 = ~n37816 ;
  assign y21557 = n37821 ;
  assign y21558 = n37822 ;
  assign y21559 = ~n37826 ;
  assign y21560 = ~n820 ;
  assign y21561 = n37827 ;
  assign y21562 = ~1'b0 ;
  assign y21563 = ~n37830 ;
  assign y21564 = 1'b0 ;
  assign y21565 = n37832 ;
  assign y21566 = ~1'b0 ;
  assign y21567 = ~n37834 ;
  assign y21568 = ~1'b0 ;
  assign y21569 = ~n37835 ;
  assign y21570 = ~n37839 ;
  assign y21571 = n14480 ;
  assign y21572 = n37840 ;
  assign y21573 = n37841 ;
  assign y21574 = n37843 ;
  assign y21575 = ~1'b0 ;
  assign y21576 = n37845 ;
  assign y21577 = ~1'b0 ;
  assign y21578 = ~n37846 ;
  assign y21579 = n37852 ;
  assign y21580 = n37855 ;
  assign y21581 = n37856 ;
  assign y21582 = ~n37863 ;
  assign y21583 = n37864 ;
  assign y21584 = ~n37866 ;
  assign y21585 = ~n37867 ;
  assign y21586 = n37868 ;
  assign y21587 = ~n14493 ;
  assign y21588 = ~1'b0 ;
  assign y21589 = ~1'b0 ;
  assign y21590 = n37874 ;
  assign y21591 = ~1'b0 ;
  assign y21592 = n37876 ;
  assign y21593 = ~n37879 ;
  assign y21594 = ~1'b0 ;
  assign y21595 = ~n37881 ;
  assign y21596 = n1054 ;
  assign y21597 = ~n6669 ;
  assign y21598 = ~1'b0 ;
  assign y21599 = n37884 ;
  assign y21600 = ~n37885 ;
  assign y21601 = n37887 ;
  assign y21602 = ~1'b0 ;
  assign y21603 = n37890 ;
  assign y21604 = n37894 ;
  assign y21605 = ~1'b0 ;
  assign y21606 = n37897 ;
  assign y21607 = ~1'b0 ;
  assign y21608 = ~1'b0 ;
  assign y21609 = ~n37898 ;
  assign y21610 = ~1'b0 ;
  assign y21611 = n36670 ;
  assign y21612 = n37899 ;
  assign y21613 = ~n37900 ;
  assign y21614 = n37901 ;
  assign y21615 = ~1'b0 ;
  assign y21616 = n37908 ;
  assign y21617 = n37910 ;
  assign y21618 = ~1'b0 ;
  assign y21619 = ~1'b0 ;
  assign y21620 = n37912 ;
  assign y21621 = ~n37913 ;
  assign y21622 = ~1'b0 ;
  assign y21623 = n37914 ;
  assign y21624 = ~1'b0 ;
  assign y21625 = n37917 ;
  assign y21626 = ~n37919 ;
  assign y21627 = n37920 ;
  assign y21628 = n37922 ;
  assign y21629 = ~n37923 ;
  assign y21630 = ~1'b0 ;
  assign y21631 = ~n37925 ;
  assign y21632 = ~n37928 ;
  assign y21633 = ~1'b0 ;
  assign y21634 = ~1'b0 ;
  assign y21635 = n37929 ;
  assign y21636 = ~1'b0 ;
  assign y21637 = n37931 ;
  assign y21638 = ~1'b0 ;
  assign y21639 = n37936 ;
  assign y21640 = ~n37938 ;
  assign y21641 = n37940 ;
  assign y21642 = ~n37941 ;
  assign y21643 = n37943 ;
  assign y21644 = ~n37944 ;
  assign y21645 = n37946 ;
  assign y21646 = ~1'b0 ;
  assign y21647 = ~1'b0 ;
  assign y21648 = ~n37947 ;
  assign y21649 = ~n34745 ;
  assign y21650 = ~n37950 ;
  assign y21651 = n37954 ;
  assign y21652 = ~n37955 ;
  assign y21653 = n37956 ;
  assign y21654 = n37962 ;
  assign y21655 = n37963 ;
  assign y21656 = n37968 ;
  assign y21657 = n37972 ;
  assign y21658 = n37973 ;
  assign y21659 = ~1'b0 ;
  assign y21660 = ~1'b0 ;
  assign y21661 = ~n37976 ;
  assign y21662 = n37979 ;
  assign y21663 = ~n4148 ;
  assign y21664 = ~n37981 ;
  assign y21665 = ~1'b0 ;
  assign y21666 = n37982 ;
  assign y21667 = ~1'b0 ;
  assign y21668 = ~1'b0 ;
  assign y21669 = n37984 ;
  assign y21670 = ~n37987 ;
  assign y21671 = ~n37990 ;
  assign y21672 = ~1'b0 ;
  assign y21673 = n37993 ;
  assign y21674 = n12889 ;
  assign y21675 = ~n37996 ;
  assign y21676 = ~n38000 ;
  assign y21677 = n38002 ;
  assign y21678 = n38007 ;
  assign y21679 = ~n38009 ;
  assign y21680 = ~1'b0 ;
  assign y21681 = ~1'b0 ;
  assign y21682 = ~1'b0 ;
  assign y21683 = ~1'b0 ;
  assign y21684 = n38014 ;
  assign y21685 = ~n38017 ;
  assign y21686 = ~n38019 ;
  assign y21687 = ~1'b0 ;
  assign y21688 = ~n38022 ;
  assign y21689 = ~1'b0 ;
  assign y21690 = 1'b0 ;
  assign y21691 = ~n38023 ;
  assign y21692 = ~1'b0 ;
  assign y21693 = ~1'b0 ;
  assign y21694 = ~1'b0 ;
  assign y21695 = ~n20073 ;
  assign y21696 = ~n31821 ;
  assign y21697 = ~n3928 ;
  assign y21698 = n4501 ;
  assign y21699 = ~1'b0 ;
  assign y21700 = ~1'b0 ;
  assign y21701 = ~n38026 ;
  assign y21702 = ~n38028 ;
  assign y21703 = ~1'b0 ;
  assign y21704 = n38029 ;
  assign y21705 = n38030 ;
  assign y21706 = ~1'b0 ;
  assign y21707 = ~n38031 ;
  assign y21708 = ~n861 ;
  assign y21709 = ~n38032 ;
  assign y21710 = ~n136 ;
  assign y21711 = ~1'b0 ;
  assign y21712 = ~n38036 ;
  assign y21713 = ~1'b0 ;
  assign y21714 = ~1'b0 ;
  assign y21715 = ~n38045 ;
  assign y21716 = ~n38050 ;
  assign y21717 = ~1'b0 ;
  assign y21718 = ~1'b0 ;
  assign y21719 = ~n38052 ;
  assign y21720 = n38057 ;
  assign y21721 = n17190 ;
  assign y21722 = ~n38058 ;
  assign y21723 = ~n38060 ;
  assign y21724 = ~1'b0 ;
  assign y21725 = n38061 ;
  assign y21726 = ~n38066 ;
  assign y21727 = ~1'b0 ;
  assign y21728 = ~n38067 ;
  assign y21729 = ~n38070 ;
  assign y21730 = 1'b0 ;
  assign y21731 = ~1'b0 ;
  assign y21732 = n28726 ;
  assign y21733 = ~n38071 ;
  assign y21734 = ~n38072 ;
  assign y21735 = ~1'b0 ;
  assign y21736 = n38074 ;
  assign y21737 = n38076 ;
  assign y21738 = ~n38078 ;
  assign y21739 = 1'b0 ;
  assign y21740 = ~1'b0 ;
  assign y21741 = ~1'b0 ;
  assign y21742 = ~1'b0 ;
  assign y21743 = ~1'b0 ;
  assign y21744 = ~1'b0 ;
  assign y21745 = n38079 ;
  assign y21746 = ~1'b0 ;
  assign y21747 = ~n38082 ;
  assign y21748 = ~1'b0 ;
  assign y21749 = n38083 ;
  assign y21750 = n38090 ;
  assign y21751 = ~n38094 ;
  assign y21752 = ~n38095 ;
  assign y21753 = ~n38100 ;
  assign y21754 = ~n38101 ;
  assign y21755 = ~n38103 ;
  assign y21756 = ~1'b0 ;
  assign y21757 = n34818 ;
  assign y21758 = ~n38104 ;
  assign y21759 = ~1'b0 ;
  assign y21760 = n38106 ;
  assign y21761 = ~n38109 ;
  assign y21762 = ~1'b0 ;
  assign y21763 = ~n38110 ;
  assign y21764 = n8264 ;
  assign y21765 = n38112 ;
  assign y21766 = n12916 ;
  assign y21767 = n38114 ;
  assign y21768 = ~n38115 ;
  assign y21769 = n38117 ;
  assign y21770 = ~n10903 ;
  assign y21771 = n38119 ;
  assign y21772 = ~n38121 ;
  assign y21773 = n38123 ;
  assign y21774 = n38125 ;
  assign y21775 = ~1'b0 ;
  assign y21776 = n38126 ;
  assign y21777 = ~n38130 ;
  assign y21778 = ~n38133 ;
  assign y21779 = n38141 ;
  assign y21780 = ~1'b0 ;
  assign y21781 = ~n38142 ;
  assign y21782 = n38146 ;
  assign y21783 = ~1'b0 ;
  assign y21784 = n18209 ;
  assign y21785 = ~1'b0 ;
  assign y21786 = ~1'b0 ;
  assign y21787 = n38147 ;
  assign y21788 = n38148 ;
  assign y21789 = ~n38150 ;
  assign y21790 = ~n38154 ;
  assign y21791 = ~n38156 ;
  assign y21792 = n38158 ;
  assign y21793 = ~n38159 ;
  assign y21794 = ~n38163 ;
  assign y21795 = ~n38164 ;
  assign y21796 = n38166 ;
  assign y21797 = ~n38171 ;
  assign y21798 = ~n38177 ;
  assign y21799 = ~n38183 ;
  assign y21800 = ~n38186 ;
  assign y21801 = 1'b0 ;
  assign y21802 = ~1'b0 ;
  assign y21803 = ~1'b0 ;
  assign y21804 = n38189 ;
  assign y21805 = ~n38192 ;
  assign y21806 = ~n38196 ;
  assign y21807 = n38199 ;
  assign y21808 = n38201 ;
  assign y21809 = ~n38202 ;
  assign y21810 = ~n38204 ;
  assign y21811 = ~n38220 ;
  assign y21812 = ~1'b0 ;
  assign y21813 = ~n38226 ;
  assign y21814 = n38227 ;
  assign y21815 = n38229 ;
  assign y21816 = n38238 ;
  assign y21817 = n14478 ;
  assign y21818 = ~n38239 ;
  assign y21819 = ~n38241 ;
  assign y21820 = n38243 ;
  assign y21821 = ~1'b0 ;
  assign y21822 = ~1'b0 ;
  assign y21823 = n38244 ;
  assign y21824 = ~1'b0 ;
  assign y21825 = n38245 ;
  assign y21826 = n38246 ;
  assign y21827 = ~n38247 ;
  assign y21828 = n38248 ;
  assign y21829 = n35952 ;
  assign y21830 = n38251 ;
  assign y21831 = n38252 ;
  assign y21832 = ~n38254 ;
  assign y21833 = ~n38255 ;
  assign y21834 = n38256 ;
  assign y21835 = ~n38258 ;
  assign y21836 = n38263 ;
  assign y21837 = ~n38270 ;
  assign y21838 = ~1'b0 ;
  assign y21839 = ~n38271 ;
  assign y21840 = ~n38277 ;
  assign y21841 = ~1'b0 ;
  assign y21842 = ~1'b0 ;
  assign y21843 = ~n38281 ;
  assign y21844 = ~1'b0 ;
  assign y21845 = ~1'b0 ;
  assign y21846 = n38282 ;
  assign y21847 = ~1'b0 ;
  assign y21848 = ~1'b0 ;
  assign y21849 = ~n38287 ;
  assign y21850 = ~n38289 ;
  assign y21851 = ~n38290 ;
  assign y21852 = ~n38291 ;
  assign y21853 = ~n4578 ;
  assign y21854 = ~1'b0 ;
  assign y21855 = ~n38295 ;
  assign y21856 = n38298 ;
  assign y21857 = n38299 ;
  assign y21858 = ~n15241 ;
  assign y21859 = ~n38301 ;
  assign y21860 = ~n21729 ;
  assign y21861 = ~1'b0 ;
  assign y21862 = n38302 ;
  assign y21863 = n38304 ;
  assign y21864 = ~n38306 ;
  assign y21865 = ~1'b0 ;
  assign y21866 = n29965 ;
  assign y21867 = ~n31141 ;
  assign y21868 = ~n38308 ;
  assign y21869 = ~n38309 ;
  assign y21870 = n38310 ;
  assign y21871 = ~1'b0 ;
  assign y21872 = ~n38313 ;
  assign y21873 = n38316 ;
  assign y21874 = ~1'b0 ;
  assign y21875 = n38317 ;
  assign y21876 = ~n38319 ;
  assign y21877 = ~1'b0 ;
  assign y21878 = ~n38322 ;
  assign y21879 = ~n38323 ;
  assign y21880 = n38326 ;
  assign y21881 = n38327 ;
  assign y21882 = ~n38332 ;
  assign y21883 = n38333 ;
  assign y21884 = ~1'b0 ;
  assign y21885 = ~n38334 ;
  assign y21886 = n38337 ;
  assign y21887 = ~n38340 ;
  assign y21888 = n38346 ;
  assign y21889 = n18080 ;
  assign y21890 = n38347 ;
  assign y21891 = ~n38348 ;
  assign y21892 = ~1'b0 ;
  assign y21893 = n38354 ;
  assign y21894 = n38357 ;
  assign y21895 = 1'b0 ;
  assign y21896 = ~n38363 ;
  assign y21897 = ~n21718 ;
  assign y21898 = 1'b0 ;
  assign y21899 = ~1'b0 ;
  assign y21900 = n38364 ;
  assign y21901 = ~1'b0 ;
  assign y21902 = ~1'b0 ;
  assign y21903 = ~n38366 ;
  assign y21904 = ~1'b0 ;
  assign y21905 = ~1'b0 ;
  assign y21906 = ~n35646 ;
  assign y21907 = ~1'b0 ;
  assign y21908 = ~1'b0 ;
  assign y21909 = 1'b0 ;
  assign y21910 = ~1'b0 ;
  assign y21911 = ~n38369 ;
  assign y21912 = n38370 ;
  assign y21913 = ~n38373 ;
  assign y21914 = ~1'b0 ;
  assign y21915 = n20150 ;
  assign y21916 = ~1'b0 ;
  assign y21917 = ~n38375 ;
  assign y21918 = ~1'b0 ;
  assign y21919 = n38382 ;
  assign y21920 = n38388 ;
  assign y21921 = n38389 ;
  assign y21922 = n38393 ;
  assign y21923 = ~n38396 ;
  assign y21924 = n38397 ;
  assign y21925 = n38400 ;
  assign y21926 = ~1'b0 ;
  assign y21927 = ~n38401 ;
  assign y21928 = ~n38402 ;
  assign y21929 = n38404 ;
  assign y21930 = ~n38405 ;
  assign y21931 = ~1'b0 ;
  assign y21932 = n38406 ;
  assign y21933 = n38410 ;
  assign y21934 = ~n38412 ;
  assign y21935 = ~n38415 ;
  assign y21936 = ~n38417 ;
  assign y21937 = 1'b0 ;
  assign y21938 = 1'b0 ;
  assign y21939 = 1'b0 ;
  assign y21940 = ~n38419 ;
  assign y21941 = n38420 ;
  assign y21942 = n38422 ;
  assign y21943 = ~n38423 ;
  assign y21944 = ~1'b0 ;
  assign y21945 = ~n38425 ;
  assign y21946 = n38427 ;
  assign y21947 = ~1'b0 ;
  assign y21948 = n25800 ;
  assign y21949 = ~1'b0 ;
  assign y21950 = ~n38428 ;
  assign y21951 = ~n38432 ;
  assign y21952 = n38433 ;
  assign y21953 = ~n38439 ;
  assign y21954 = ~1'b0 ;
  assign y21955 = n38440 ;
  assign y21956 = ~1'b0 ;
  assign y21957 = ~1'b0 ;
  assign y21958 = n38442 ;
  assign y21959 = n38446 ;
  assign y21960 = n38448 ;
  assign y21961 = n38450 ;
  assign y21962 = ~1'b0 ;
  assign y21963 = ~n38454 ;
  assign y21964 = ~1'b0 ;
  assign y21965 = ~n33019 ;
  assign y21966 = ~1'b0 ;
  assign y21967 = ~n38464 ;
  assign y21968 = n38465 ;
  assign y21969 = n38468 ;
  assign y21970 = ~n38470 ;
  assign y21971 = n38471 ;
  assign y21972 = ~1'b0 ;
  assign y21973 = ~1'b0 ;
  assign y21974 = n38472 ;
  assign y21975 = ~n38474 ;
  assign y21976 = ~n27302 ;
  assign y21977 = ~n38475 ;
  assign y21978 = ~n104 ;
  assign y21979 = ~n38476 ;
  assign y21980 = ~1'b0 ;
  assign y21981 = ~n38477 ;
  assign y21982 = 1'b0 ;
  assign y21983 = ~n38479 ;
  assign y21984 = ~n1690 ;
  assign y21985 = ~n38487 ;
  assign y21986 = ~n4360 ;
  assign y21987 = ~n38494 ;
  assign y21988 = n38495 ;
  assign y21989 = ~1'b0 ;
  assign y21990 = ~1'b0 ;
  assign y21991 = ~n38499 ;
  assign y21992 = ~1'b0 ;
  assign y21993 = n38502 ;
  assign y21994 = ~1'b0 ;
  assign y21995 = ~n38504 ;
  assign y21996 = ~n38508 ;
  assign y21997 = ~n38509 ;
  assign y21998 = ~n38514 ;
  assign y21999 = n38517 ;
  assign y22000 = ~n38519 ;
  assign y22001 = ~1'b0 ;
  assign y22002 = ~1'b0 ;
  assign y22003 = n21877 ;
  assign y22004 = ~1'b0 ;
  assign y22005 = ~n38522 ;
  assign y22006 = ~1'b0 ;
  assign y22007 = ~n38523 ;
  assign y22008 = n38524 ;
  assign y22009 = n38525 ;
  assign y22010 = ~1'b0 ;
  assign y22011 = ~1'b0 ;
  assign y22012 = ~1'b0 ;
  assign y22013 = ~1'b0 ;
  assign y22014 = ~n38530 ;
  assign y22015 = ~n38534 ;
  assign y22016 = n34327 ;
  assign y22017 = n38537 ;
  assign y22018 = ~n38538 ;
  assign y22019 = ~1'b0 ;
  assign y22020 = n38539 ;
  assign y22021 = n38540 ;
  assign y22022 = n38548 ;
  assign y22023 = ~n38551 ;
  assign y22024 = ~n38554 ;
  assign y22025 = ~1'b0 ;
  assign y22026 = ~n38559 ;
  assign y22027 = ~n38560 ;
  assign y22028 = ~n38561 ;
  assign y22029 = n38562 ;
  assign y22030 = n38566 ;
  assign y22031 = n38567 ;
  assign y22032 = ~n28139 ;
  assign y22033 = ~1'b0 ;
  assign y22034 = ~n38573 ;
  assign y22035 = ~1'b0 ;
  assign y22036 = n38574 ;
  assign y22037 = n1769 ;
  assign y22038 = n38580 ;
  assign y22039 = ~n38583 ;
  assign y22040 = n34601 ;
  assign y22041 = ~1'b0 ;
  assign y22042 = ~n38584 ;
  assign y22043 = 1'b0 ;
  assign y22044 = ~1'b0 ;
  assign y22045 = n38588 ;
  assign y22046 = n38593 ;
  assign y22047 = ~n38595 ;
  assign y22048 = ~n38596 ;
  assign y22049 = n38597 ;
  assign y22050 = ~1'b0 ;
  assign y22051 = ~1'b0 ;
  assign y22052 = ~1'b0 ;
  assign y22053 = ~1'b0 ;
  assign y22054 = ~n38601 ;
  assign y22055 = n38603 ;
  assign y22056 = ~n38605 ;
  assign y22057 = ~1'b0 ;
  assign y22058 = ~n38608 ;
  assign y22059 = ~n9797 ;
  assign y22060 = n38609 ;
  assign y22061 = ~n38610 ;
  assign y22062 = n38612 ;
  assign y22063 = n38615 ;
  assign y22064 = ~n38620 ;
  assign y22065 = ~n17938 ;
  assign y22066 = ~n38621 ;
  assign y22067 = ~n38623 ;
  assign y22068 = n38629 ;
  assign y22069 = ~n38630 ;
  assign y22070 = ~n16663 ;
  assign y22071 = n38631 ;
  assign y22072 = n38632 ;
  assign y22073 = ~n38634 ;
  assign y22074 = ~1'b0 ;
  assign y22075 = ~1'b0 ;
  assign y22076 = ~1'b0 ;
  assign y22077 = ~n38635 ;
  assign y22078 = n38638 ;
  assign y22079 = ~n38641 ;
  assign y22080 = ~1'b0 ;
  assign y22081 = ~1'b0 ;
  assign y22082 = n38642 ;
  assign y22083 = n38647 ;
  assign y22084 = ~n38651 ;
  assign y22085 = ~1'b0 ;
  assign y22086 = ~n38653 ;
  assign y22087 = ~n38654 ;
  assign y22088 = n38656 ;
  assign y22089 = ~n38657 ;
  assign y22090 = ~n38658 ;
  assign y22091 = ~1'b0 ;
  assign y22092 = ~n38664 ;
  assign y22093 = ~1'b0 ;
  assign y22094 = n38665 ;
  assign y22095 = 1'b0 ;
  assign y22096 = n38671 ;
  assign y22097 = n38672 ;
  assign y22098 = ~n38673 ;
  assign y22099 = ~n38675 ;
  assign y22100 = ~1'b0 ;
  assign y22101 = 1'b0 ;
  assign y22102 = ~n38676 ;
  assign y22103 = ~n26824 ;
  assign y22104 = ~1'b0 ;
  assign y22105 = n38680 ;
  assign y22106 = n38681 ;
  assign y22107 = 1'b0 ;
  assign y22108 = ~1'b0 ;
  assign y22109 = n38683 ;
  assign y22110 = ~1'b0 ;
  assign y22111 = ~1'b0 ;
  assign y22112 = ~n38688 ;
  assign y22113 = n38690 ;
  assign y22114 = ~1'b0 ;
  assign y22115 = ~n11520 ;
  assign y22116 = 1'b0 ;
  assign y22117 = n38691 ;
  assign y22118 = n38694 ;
  assign y22119 = n38698 ;
  assign y22120 = n38706 ;
  assign y22121 = n5695 ;
  assign y22122 = ~n13632 ;
  assign y22123 = ~n38708 ;
  assign y22124 = ~1'b0 ;
  assign y22125 = n38710 ;
  assign y22126 = ~1'b0 ;
  assign y22127 = ~1'b0 ;
  assign y22128 = ~n38714 ;
  assign y22129 = n38715 ;
  assign y22130 = ~n38717 ;
  assign y22131 = n38720 ;
  assign y22132 = ~n38724 ;
  assign y22133 = n38725 ;
  assign y22134 = ~n38734 ;
  assign y22135 = ~1'b0 ;
  assign y22136 = ~n38738 ;
  assign y22137 = n38743 ;
  assign y22138 = n6292 ;
  assign y22139 = ~1'b0 ;
  assign y22140 = ~n38745 ;
  assign y22141 = n38750 ;
  assign y22142 = ~1'b0 ;
  assign y22143 = ~1'b0 ;
  assign y22144 = ~1'b0 ;
  assign y22145 = ~n38752 ;
  assign y22146 = ~1'b0 ;
  assign y22147 = ~1'b0 ;
  assign y22148 = n38753 ;
  assign y22149 = ~1'b0 ;
  assign y22150 = n38756 ;
  assign y22151 = ~1'b0 ;
  assign y22152 = n38758 ;
  assign y22153 = n38761 ;
  assign y22154 = ~n38765 ;
  assign y22155 = n38767 ;
  assign y22156 = ~1'b0 ;
  assign y22157 = ~n38770 ;
  assign y22158 = ~n38774 ;
  assign y22159 = n38778 ;
  assign y22160 = ~n38780 ;
  assign y22161 = ~1'b0 ;
  assign y22162 = n38783 ;
  assign y22163 = ~n38784 ;
  assign y22164 = ~n10854 ;
  assign y22165 = ~n19564 ;
  assign y22166 = ~1'b0 ;
  assign y22167 = ~n38793 ;
  assign y22168 = ~n38795 ;
  assign y22169 = ~1'b0 ;
  assign y22170 = n38796 ;
  assign y22171 = ~n38799 ;
  assign y22172 = n38800 ;
  assign y22173 = ~n1763 ;
  assign y22174 = ~n38801 ;
  assign y22175 = n38807 ;
  assign y22176 = n38811 ;
  assign y22177 = ~1'b0 ;
  assign y22178 = ~1'b0 ;
  assign y22179 = n38816 ;
  assign y22180 = ~n38826 ;
  assign y22181 = ~n38828 ;
  assign y22182 = n38833 ;
  assign y22183 = ~1'b0 ;
  assign y22184 = ~n38835 ;
  assign y22185 = ~n38836 ;
  assign y22186 = ~1'b0 ;
  assign y22187 = ~n8843 ;
  assign y22188 = ~n38837 ;
  assign y22189 = ~n38838 ;
  assign y22190 = ~n38840 ;
  assign y22191 = n38841 ;
  assign y22192 = ~n38849 ;
  assign y22193 = ~1'b0 ;
  assign y22194 = ~n38850 ;
  assign y22195 = n38853 ;
  assign y22196 = n38854 ;
  assign y22197 = n38855 ;
  assign y22198 = ~n38857 ;
  assign y22199 = ~n38859 ;
  assign y22200 = ~1'b0 ;
  assign y22201 = ~1'b0 ;
  assign y22202 = ~n38861 ;
  assign y22203 = ~n38865 ;
  assign y22204 = ~n38868 ;
  assign y22205 = ~n38873 ;
  assign y22206 = ~n6968 ;
  assign y22207 = ~1'b0 ;
  assign y22208 = n38876 ;
  assign y22209 = n38882 ;
  assign y22210 = ~1'b0 ;
  assign y22211 = ~1'b0 ;
  assign y22212 = n38883 ;
  assign y22213 = ~n20272 ;
  assign y22214 = ~n38884 ;
  assign y22215 = ~1'b0 ;
  assign y22216 = ~1'b0 ;
  assign y22217 = ~n38889 ;
  assign y22218 = ~n38890 ;
  assign y22219 = ~n38893 ;
  assign y22220 = ~n38894 ;
  assign y22221 = ~n38895 ;
  assign y22222 = n38896 ;
  assign y22223 = n38897 ;
  assign y22224 = ~1'b0 ;
  assign y22225 = ~1'b0 ;
  assign y22226 = n38903 ;
  assign y22227 = n38904 ;
  assign y22228 = ~n38910 ;
  assign y22229 = n782 ;
  assign y22230 = ~1'b0 ;
  assign y22231 = ~n38911 ;
  assign y22232 = n38912 ;
  assign y22233 = ~n38913 ;
  assign y22234 = ~n36409 ;
  assign y22235 = ~1'b0 ;
  assign y22236 = n38919 ;
  assign y22237 = ~1'b0 ;
  assign y22238 = ~n38921 ;
  assign y22239 = ~n38923 ;
  assign y22240 = n32139 ;
  assign y22241 = ~1'b0 ;
  assign y22242 = n38925 ;
  assign y22243 = ~1'b0 ;
  assign y22244 = ~n38929 ;
  assign y22245 = ~n38931 ;
  assign y22246 = ~n38932 ;
  assign y22247 = n38933 ;
  assign y22248 = ~n38936 ;
  assign y22249 = n38938 ;
  assign y22250 = ~1'b0 ;
  assign y22251 = ~1'b0 ;
  assign y22252 = ~n38940 ;
  assign y22253 = n38941 ;
  assign y22254 = ~n38944 ;
  assign y22255 = n38947 ;
  assign y22256 = ~1'b0 ;
  assign y22257 = ~n38948 ;
  assign y22258 = 1'b0 ;
  assign y22259 = ~1'b0 ;
  assign y22260 = ~n38950 ;
  assign y22261 = ~n38952 ;
  assign y22262 = ~1'b0 ;
  assign y22263 = n38953 ;
  assign y22264 = n38955 ;
  assign y22265 = ~n38958 ;
  assign y22266 = n38959 ;
  assign y22267 = ~n38960 ;
  assign y22268 = ~1'b0 ;
  assign y22269 = ~n38961 ;
  assign y22270 = ~n38962 ;
  assign y22271 = n38963 ;
  assign y22272 = n38966 ;
  assign y22273 = n38971 ;
  assign y22274 = ~1'b0 ;
  assign y22275 = ~n38975 ;
  assign y22276 = ~1'b0 ;
  assign y22277 = n38977 ;
  assign y22278 = ~n38979 ;
  assign y22279 = ~n38983 ;
  assign y22280 = ~n38984 ;
  assign y22281 = n38986 ;
  assign y22282 = n38988 ;
  assign y22283 = ~n38990 ;
  assign y22284 = n38992 ;
  assign y22285 = n38993 ;
  assign y22286 = n38994 ;
  assign y22287 = n38995 ;
  assign y22288 = ~1'b0 ;
  assign y22289 = ~n38996 ;
  assign y22290 = n38997 ;
  assign y22291 = ~n38999 ;
  assign y22292 = ~1'b0 ;
  assign y22293 = n39003 ;
  assign y22294 = ~n39005 ;
  assign y22295 = ~1'b0 ;
  assign y22296 = n39012 ;
  assign y22297 = ~1'b0 ;
  assign y22298 = ~n39013 ;
  assign y22299 = ~n20488 ;
  assign y22300 = ~n39014 ;
  assign y22301 = n39015 ;
  assign y22302 = 1'b0 ;
  assign y22303 = ~n39016 ;
  assign y22304 = n39017 ;
  assign y22305 = n39019 ;
  assign y22306 = ~1'b0 ;
  assign y22307 = ~1'b0 ;
  assign y22308 = ~n39028 ;
  assign y22309 = ~n19993 ;
  assign y22310 = ~1'b0 ;
  assign y22311 = n39030 ;
  assign y22312 = ~1'b0 ;
  assign y22313 = n39031 ;
  assign y22314 = ~n39035 ;
  assign y22315 = ~n39041 ;
  assign y22316 = ~n39043 ;
  assign y22317 = n39045 ;
  assign y22318 = n39047 ;
  assign y22319 = n39048 ;
  assign y22320 = n3225 ;
  assign y22321 = n39050 ;
  assign y22322 = ~1'b0 ;
  assign y22323 = ~n39052 ;
  assign y22324 = ~n39053 ;
  assign y22325 = n14534 ;
  assign y22326 = ~n10428 ;
  assign y22327 = ~n39054 ;
  assign y22328 = ~1'b0 ;
  assign y22329 = ~n39058 ;
  assign y22330 = ~1'b0 ;
  assign y22331 = 1'b0 ;
  assign y22332 = ~1'b0 ;
  assign y22333 = n39062 ;
  assign y22334 = n39065 ;
  assign y22335 = ~n1075 ;
  assign y22336 = n39066 ;
  assign y22337 = ~1'b0 ;
  assign y22338 = ~1'b0 ;
  assign y22339 = ~n39069 ;
  assign y22340 = ~n39073 ;
  assign y22341 = n39074 ;
  assign y22342 = n39075 ;
  assign y22343 = 1'b0 ;
  assign y22344 = ~n39077 ;
  assign y22345 = ~n39081 ;
  assign y22346 = ~1'b0 ;
  assign y22347 = ~1'b0 ;
  assign y22348 = ~n39086 ;
  assign y22349 = ~1'b0 ;
  assign y22350 = n8634 ;
  assign y22351 = ~n39088 ;
  assign y22352 = n11216 ;
  assign y22353 = ~1'b0 ;
  assign y22354 = n39089 ;
  assign y22355 = ~1'b0 ;
  assign y22356 = n39091 ;
  assign y22357 = ~1'b0 ;
  assign y22358 = ~1'b0 ;
  assign y22359 = ~1'b0 ;
  assign y22360 = n30845 ;
  assign y22361 = ~1'b0 ;
  assign y22362 = ~1'b0 ;
  assign y22363 = ~n13063 ;
  assign y22364 = ~n39095 ;
  assign y22365 = 1'b0 ;
  assign y22366 = ~n32046 ;
  assign y22367 = ~n39096 ;
  assign y22368 = ~n39098 ;
  assign y22369 = ~n39100 ;
  assign y22370 = n39103 ;
  assign y22371 = n39104 ;
  assign y22372 = ~n39107 ;
  assign y22373 = ~n39108 ;
  assign y22374 = n39109 ;
  assign y22375 = ~n39111 ;
  assign y22376 = ~1'b0 ;
  assign y22377 = ~n39114 ;
  assign y22378 = ~n39115 ;
  assign y22379 = n7913 ;
  assign y22380 = n26347 ;
  assign y22381 = ~n39119 ;
  assign y22382 = n39120 ;
  assign y22383 = ~n39125 ;
  assign y22384 = n39126 ;
  assign y22385 = ~1'b0 ;
  assign y22386 = ~n39130 ;
  assign y22387 = n39133 ;
  assign y22388 = n39138 ;
  assign y22389 = n3823 ;
  assign y22390 = ~n39140 ;
  assign y22391 = ~1'b0 ;
  assign y22392 = ~1'b0 ;
  assign y22393 = ~n39143 ;
  assign y22394 = ~n39144 ;
  assign y22395 = n39147 ;
  assign y22396 = ~n39149 ;
  assign y22397 = ~1'b0 ;
  assign y22398 = ~n16445 ;
  assign y22399 = ~1'b0 ;
  assign y22400 = ~n39156 ;
  assign y22401 = n39158 ;
  assign y22402 = n1771 ;
  assign y22403 = n39160 ;
  assign y22404 = ~1'b0 ;
  assign y22405 = n39162 ;
  assign y22406 = ~n39163 ;
  assign y22407 = ~n39167 ;
  assign y22408 = n39169 ;
  assign y22409 = n39170 ;
  assign y22410 = n39176 ;
  assign y22411 = ~n39178 ;
  assign y22412 = n39180 ;
  assign y22413 = ~1'b0 ;
  assign y22414 = ~n24149 ;
  assign y22415 = n39181 ;
  assign y22416 = ~1'b0 ;
  assign y22417 = ~n35581 ;
  assign y22418 = 1'b0 ;
  assign y22419 = 1'b0 ;
  assign y22420 = ~n39183 ;
  assign y22421 = n23971 ;
  assign y22422 = ~n39184 ;
  assign y22423 = n35099 ;
  assign y22424 = ~1'b0 ;
  assign y22425 = ~1'b0 ;
  assign y22426 = n39186 ;
  assign y22427 = n39187 ;
  assign y22428 = n39188 ;
  assign y22429 = ~n39189 ;
  assign y22430 = ~n4372 ;
  assign y22431 = ~1'b0 ;
  assign y22432 = n39191 ;
  assign y22433 = n39193 ;
  assign y22434 = ~1'b0 ;
  assign y22435 = ~n16534 ;
  assign y22436 = 1'b0 ;
  assign y22437 = ~n39195 ;
  assign y22438 = ~1'b0 ;
  assign y22439 = n21872 ;
  assign y22440 = n39196 ;
  assign y22441 = n9390 ;
  assign y22442 = ~n39198 ;
  assign y22443 = 1'b0 ;
  assign y22444 = ~n39199 ;
  assign y22445 = n3550 ;
  assign y22446 = ~1'b0 ;
  assign y22447 = ~1'b0 ;
  assign y22448 = ~1'b0 ;
  assign y22449 = ~1'b0 ;
  assign y22450 = n39201 ;
  assign y22451 = 1'b0 ;
  assign y22452 = ~n39202 ;
  assign y22453 = 1'b0 ;
  assign y22454 = ~n39204 ;
  assign y22455 = ~n3034 ;
  assign y22456 = ~1'b0 ;
  assign y22457 = ~1'b0 ;
  assign y22458 = n39205 ;
  assign y22459 = n39207 ;
  assign y22460 = ~1'b0 ;
  assign y22461 = ~1'b0 ;
  assign y22462 = ~n4451 ;
  assign y22463 = ~n39211 ;
  assign y22464 = ~n39213 ;
  assign y22465 = n39217 ;
  assign y22466 = 1'b0 ;
  assign y22467 = ~n39223 ;
  assign y22468 = 1'b0 ;
  assign y22469 = ~n39225 ;
  assign y22470 = ~n39226 ;
  assign y22471 = n39227 ;
  assign y22472 = ~1'b0 ;
  assign y22473 = ~n39228 ;
  assign y22474 = ~1'b0 ;
  assign y22475 = n39232 ;
  assign y22476 = ~n10702 ;
  assign y22477 = ~n39236 ;
  assign y22478 = ~1'b0 ;
  assign y22479 = ~n39237 ;
  assign y22480 = ~1'b0 ;
  assign y22481 = ~n39239 ;
  assign y22482 = ~n39241 ;
  assign y22483 = ~n39243 ;
  assign y22484 = ~n39244 ;
  assign y22485 = n39246 ;
  assign y22486 = ~1'b0 ;
  assign y22487 = n39249 ;
  assign y22488 = n39257 ;
  assign y22489 = n39259 ;
  assign y22490 = ~1'b0 ;
  assign y22491 = n39261 ;
  assign y22492 = ~1'b0 ;
  assign y22493 = ~1'b0 ;
  assign y22494 = ~n39263 ;
  assign y22495 = ~n39265 ;
  assign y22496 = ~1'b0 ;
  assign y22497 = ~1'b0 ;
  assign y22498 = ~n39266 ;
  assign y22499 = ~1'b0 ;
  assign y22500 = ~n39267 ;
  assign y22501 = ~n39269 ;
  assign y22502 = n20917 ;
  assign y22503 = n39273 ;
  assign y22504 = ~n39276 ;
  assign y22505 = n39281 ;
  assign y22506 = 1'b0 ;
  assign y22507 = ~n39283 ;
  assign y22508 = 1'b0 ;
  assign y22509 = ~n39284 ;
  assign y22510 = ~n39290 ;
  assign y22511 = n39294 ;
  assign y22512 = n39297 ;
  assign y22513 = ~n39300 ;
  assign y22514 = ~n39302 ;
  assign y22515 = n39304 ;
  assign y22516 = n39305 ;
  assign y22517 = ~n39307 ;
  assign y22518 = ~1'b0 ;
  assign y22519 = ~n39308 ;
  assign y22520 = n39309 ;
  assign y22521 = 1'b0 ;
  assign y22522 = ~1'b0 ;
  assign y22523 = n22881 ;
  assign y22524 = ~n39312 ;
  assign y22525 = ~n39314 ;
  assign y22526 = ~n39315 ;
  assign y22527 = ~n39317 ;
  assign y22528 = ~1'b0 ;
  assign y22529 = n39318 ;
  assign y22530 = n39319 ;
  assign y22531 = n39321 ;
  assign y22532 = ~1'b0 ;
  assign y22533 = ~n39323 ;
  assign y22534 = ~1'b0 ;
  assign y22535 = n39328 ;
  assign y22536 = n39329 ;
  assign y22537 = n39334 ;
  assign y22538 = ~n39338 ;
  assign y22539 = ~1'b0 ;
  assign y22540 = n39343 ;
  assign y22541 = ~1'b0 ;
  assign y22542 = ~n39344 ;
  assign y22543 = ~n881 ;
  assign y22544 = ~1'b0 ;
  assign y22545 = ~n39347 ;
  assign y22546 = n39348 ;
  assign y22547 = ~1'b0 ;
  assign y22548 = ~1'b0 ;
  assign y22549 = ~1'b0 ;
  assign y22550 = n39350 ;
  assign y22551 = n39352 ;
  assign y22552 = n39353 ;
  assign y22553 = ~n39354 ;
  assign y22554 = ~n39355 ;
  assign y22555 = ~1'b0 ;
  assign y22556 = n39356 ;
  assign y22557 = ~n39358 ;
  assign y22558 = ~1'b0 ;
  assign y22559 = n32934 ;
  assign y22560 = ~n39363 ;
  assign y22561 = ~1'b0 ;
  assign y22562 = ~n39368 ;
  assign y22563 = ~1'b0 ;
  assign y22564 = n39370 ;
  assign y22565 = ~n39374 ;
  assign y22566 = ~1'b0 ;
  assign y22567 = n39375 ;
  assign y22568 = ~1'b0 ;
  assign y22569 = ~1'b0 ;
  assign y22570 = n39376 ;
  assign y22571 = n39381 ;
  assign y22572 = ~n39388 ;
  assign y22573 = ~n13293 ;
  assign y22574 = 1'b0 ;
  assign y22575 = n39389 ;
  assign y22576 = ~n39390 ;
  assign y22577 = ~n39392 ;
  assign y22578 = ~n39393 ;
  assign y22579 = ~1'b0 ;
  assign y22580 = ~1'b0 ;
  assign y22581 = ~1'b0 ;
  assign y22582 = ~n39404 ;
  assign y22583 = n39407 ;
  assign y22584 = ~n39408 ;
  assign y22585 = n2927 ;
  assign y22586 = ~n39409 ;
  assign y22587 = ~n39410 ;
  assign y22588 = n39414 ;
  assign y22589 = ~n28699 ;
  assign y22590 = n39418 ;
  assign y22591 = ~n39420 ;
  assign y22592 = ~1'b0 ;
  assign y22593 = ~n39424 ;
  assign y22594 = n39426 ;
  assign y22595 = ~1'b0 ;
  assign y22596 = n39427 ;
  assign y22597 = n39428 ;
  assign y22598 = ~n9795 ;
  assign y22599 = ~1'b0 ;
  assign y22600 = ~1'b0 ;
  assign y22601 = ~n39429 ;
  assign y22602 = n39431 ;
  assign y22603 = ~n39433 ;
  assign y22604 = ~n39434 ;
  assign y22605 = n39440 ;
  assign y22606 = n39444 ;
  assign y22607 = ~n39446 ;
  assign y22608 = 1'b0 ;
  assign y22609 = ~1'b0 ;
  assign y22610 = ~n39452 ;
  assign y22611 = ~n39454 ;
  assign y22612 = 1'b0 ;
  assign y22613 = ~n39459 ;
  assign y22614 = n39464 ;
  assign y22615 = n39466 ;
  assign y22616 = ~1'b0 ;
  assign y22617 = n39468 ;
  assign y22618 = n39470 ;
  assign y22619 = ~n39472 ;
  assign y22620 = n39475 ;
  assign y22621 = ~n39477 ;
  assign y22622 = ~n39483 ;
  assign y22623 = ~1'b0 ;
  assign y22624 = n39486 ;
  assign y22625 = n39488 ;
  assign y22626 = ~n39495 ;
  assign y22627 = ~1'b0 ;
  assign y22628 = n39497 ;
  assign y22629 = n39501 ;
  assign y22630 = ~n39502 ;
  assign y22631 = ~n39504 ;
  assign y22632 = ~1'b0 ;
  assign y22633 = n39506 ;
  assign y22634 = n39507 ;
  assign y22635 = ~1'b0 ;
  assign y22636 = ~1'b0 ;
  assign y22637 = ~n39510 ;
  assign y22638 = n39511 ;
  assign y22639 = ~n39512 ;
  assign y22640 = ~1'b0 ;
  assign y22641 = ~n39513 ;
  assign y22642 = ~1'b0 ;
  assign y22643 = ~1'b0 ;
  assign y22644 = ~n39517 ;
  assign y22645 = ~n976 ;
  assign y22646 = n39519 ;
  assign y22647 = n39520 ;
  assign y22648 = ~n39523 ;
  assign y22649 = ~1'b0 ;
  assign y22650 = ~1'b0 ;
  assign y22651 = ~1'b0 ;
  assign y22652 = ~n39528 ;
  assign y22653 = n39530 ;
  assign y22654 = n39531 ;
  assign y22655 = ~n39532 ;
  assign y22656 = ~n39534 ;
  assign y22657 = ~1'b0 ;
  assign y22658 = n39535 ;
  assign y22659 = ~n39540 ;
  assign y22660 = n39542 ;
  assign y22661 = n39543 ;
  assign y22662 = ~1'b0 ;
  assign y22663 = n39544 ;
  assign y22664 = ~n39545 ;
  assign y22665 = 1'b0 ;
  assign y22666 = n39547 ;
  assign y22667 = n39549 ;
  assign y22668 = ~n39551 ;
  assign y22669 = ~n21935 ;
  assign y22670 = ~1'b0 ;
  assign y22671 = ~1'b0 ;
  assign y22672 = ~1'b0 ;
  assign y22673 = n39555 ;
  assign y22674 = n4317 ;
  assign y22675 = ~n39044 ;
  assign y22676 = ~1'b0 ;
  assign y22677 = n39556 ;
  assign y22678 = ~1'b0 ;
  assign y22679 = ~1'b0 ;
  assign y22680 = n39558 ;
  assign y22681 = ~n39559 ;
  assign y22682 = ~1'b0 ;
  assign y22683 = ~1'b0 ;
  assign y22684 = ~n39560 ;
  assign y22685 = ~1'b0 ;
  assign y22686 = ~1'b0 ;
  assign y22687 = ~n39564 ;
  assign y22688 = n26991 ;
  assign y22689 = ~n39566 ;
  assign y22690 = ~n39570 ;
  assign y22691 = n39572 ;
  assign y22692 = ~1'b0 ;
  assign y22693 = ~1'b0 ;
  assign y22694 = ~1'b0 ;
  assign y22695 = n39576 ;
  assign y22696 = n39583 ;
  assign y22697 = ~1'b0 ;
  assign y22698 = n39584 ;
  assign y22699 = ~1'b0 ;
  assign y22700 = ~1'b0 ;
  assign y22701 = ~n39586 ;
  assign y22702 = n39588 ;
  assign y22703 = n39595 ;
  assign y22704 = n39596 ;
  assign y22705 = n39598 ;
  assign y22706 = n39599 ;
  assign y22707 = 1'b0 ;
  assign y22708 = ~n38281 ;
  assign y22709 = ~1'b0 ;
  assign y22710 = n39601 ;
  assign y22711 = 1'b0 ;
  assign y22712 = n39602 ;
  assign y22713 = ~n39603 ;
  assign y22714 = ~1'b0 ;
  assign y22715 = n39605 ;
  assign y22716 = n39611 ;
  assign y22717 = ~n39613 ;
  assign y22718 = ~n39617 ;
  assign y22719 = n20868 ;
  assign y22720 = ~1'b0 ;
  assign y22721 = ~n39618 ;
  assign y22722 = ~n39620 ;
  assign y22723 = ~1'b0 ;
  assign y22724 = n39621 ;
  assign y22725 = n39622 ;
  assign y22726 = ~n39624 ;
  assign y22727 = n22399 ;
  assign y22728 = ~n39628 ;
  assign y22729 = n39631 ;
  assign y22730 = n39634 ;
  assign y22731 = n39635 ;
  assign y22732 = n39636 ;
  assign y22733 = ~n39640 ;
  assign y22734 = ~n39641 ;
  assign y22735 = ~1'b0 ;
  assign y22736 = ~1'b0 ;
  assign y22737 = ~1'b0 ;
  assign y22738 = ~1'b0 ;
  assign y22739 = ~n39642 ;
  assign y22740 = ~n39645 ;
  assign y22741 = n39647 ;
  assign y22742 = ~n39648 ;
  assign y22743 = ~1'b0 ;
  assign y22744 = ~n39650 ;
  assign y22745 = ~n39654 ;
  assign y22746 = ~1'b0 ;
  assign y22747 = n33452 ;
  assign y22748 = n39655 ;
  assign y22749 = n2637 ;
  assign y22750 = ~1'b0 ;
  assign y22751 = ~n39657 ;
  assign y22752 = ~n39661 ;
  assign y22753 = ~1'b0 ;
  assign y22754 = ~1'b0 ;
  assign y22755 = ~n39665 ;
  assign y22756 = ~n39670 ;
  assign y22757 = ~n39674 ;
  assign y22758 = n39676 ;
  assign y22759 = n39679 ;
  assign y22760 = ~n10955 ;
  assign y22761 = n39683 ;
  assign y22762 = ~n39684 ;
  assign y22763 = n15544 ;
  assign y22764 = ~n39689 ;
  assign y22765 = 1'b0 ;
  assign y22766 = n39692 ;
  assign y22767 = n39694 ;
  assign y22768 = ~n39696 ;
  assign y22769 = ~n17840 ;
  assign y22770 = ~1'b0 ;
  assign y22771 = n39698 ;
  assign y22772 = n39699 ;
  assign y22773 = ~1'b0 ;
  assign y22774 = n39700 ;
  assign y22775 = ~1'b0 ;
  assign y22776 = ~1'b0 ;
  assign y22777 = n39702 ;
  assign y22778 = n39704 ;
  assign y22779 = n39706 ;
  assign y22780 = ~1'b0 ;
  assign y22781 = ~1'b0 ;
  assign y22782 = ~1'b0 ;
  assign y22783 = n39710 ;
  assign y22784 = ~1'b0 ;
  assign y22785 = ~1'b0 ;
  assign y22786 = n39711 ;
  assign y22787 = n39714 ;
  assign y22788 = ~1'b0 ;
  assign y22789 = ~1'b0 ;
  assign y22790 = n39715 ;
  assign y22791 = n10348 ;
  assign y22792 = ~n39716 ;
  assign y22793 = ~1'b0 ;
  assign y22794 = ~1'b0 ;
  assign y22795 = ~n39717 ;
  assign y22796 = 1'b0 ;
  assign y22797 = ~n39719 ;
  assign y22798 = ~1'b0 ;
  assign y22799 = n39725 ;
  assign y22800 = ~n39726 ;
  assign y22801 = ~1'b0 ;
  assign y22802 = ~1'b0 ;
  assign y22803 = ~1'b0 ;
  assign y22804 = n39732 ;
  assign y22805 = ~1'b0 ;
  assign y22806 = ~n39738 ;
  assign y22807 = ~1'b0 ;
  assign y22808 = ~n39740 ;
  assign y22809 = ~n39741 ;
  assign y22810 = n39743 ;
  assign y22811 = ~1'b0 ;
  assign y22812 = 1'b0 ;
  assign y22813 = 1'b0 ;
  assign y22814 = ~1'b0 ;
  assign y22815 = ~n39745 ;
  assign y22816 = ~1'b0 ;
  assign y22817 = 1'b0 ;
  assign y22818 = n39747 ;
  assign y22819 = 1'b0 ;
  assign y22820 = n39748 ;
  assign y22821 = n39749 ;
  assign y22822 = ~n39750 ;
  assign y22823 = ~1'b0 ;
  assign y22824 = ~1'b0 ;
  assign y22825 = 1'b0 ;
  assign y22826 = ~1'b0 ;
  assign y22827 = n39751 ;
  assign y22828 = ~1'b0 ;
  assign y22829 = ~n39752 ;
  assign y22830 = n39753 ;
  assign y22831 = n13916 ;
  assign y22832 = ~n39755 ;
  assign y22833 = ~n39756 ;
  assign y22834 = n14750 ;
  assign y22835 = ~1'b0 ;
  assign y22836 = ~n39757 ;
  assign y22837 = ~1'b0 ;
  assign y22838 = n39759 ;
  assign y22839 = ~1'b0 ;
  assign y22840 = n39760 ;
  assign y22841 = n39761 ;
  assign y22842 = ~n39766 ;
  assign y22843 = n39768 ;
  assign y22844 = n39770 ;
  assign y22845 = n39773 ;
  assign y22846 = ~1'b0 ;
  assign y22847 = n39774 ;
  assign y22848 = ~1'b0 ;
  assign y22849 = ~1'b0 ;
  assign y22850 = ~n39777 ;
  assign y22851 = ~n39779 ;
  assign y22852 = ~1'b0 ;
  assign y22853 = n39782 ;
  assign y22854 = ~1'b0 ;
  assign y22855 = n39784 ;
  assign y22856 = ~n22935 ;
  assign y22857 = ~1'b0 ;
  assign y22858 = ~1'b0 ;
  assign y22859 = ~n39786 ;
  assign y22860 = n39788 ;
  assign y22861 = ~1'b0 ;
  assign y22862 = n39793 ;
  assign y22863 = ~1'b0 ;
  assign y22864 = ~1'b0 ;
  assign y22865 = n39799 ;
  assign y22866 = n39801 ;
  assign y22867 = ~n39804 ;
  assign y22868 = ~1'b0 ;
  assign y22869 = n39805 ;
  assign y22870 = n39806 ;
  assign y22871 = ~1'b0 ;
  assign y22872 = ~1'b0 ;
  assign y22873 = ~n39809 ;
  assign y22874 = n39811 ;
  assign y22875 = n25555 ;
  assign y22876 = ~1'b0 ;
  assign y22877 = n39812 ;
  assign y22878 = ~n39814 ;
  assign y22879 = ~n39815 ;
  assign y22880 = n39819 ;
  assign y22881 = ~n39822 ;
  assign y22882 = ~1'b0 ;
  assign y22883 = ~1'b0 ;
  assign y22884 = ~1'b0 ;
  assign y22885 = ~1'b0 ;
  assign y22886 = ~n39824 ;
  assign y22887 = ~n39827 ;
  assign y22888 = ~1'b0 ;
  assign y22889 = ~1'b0 ;
  assign y22890 = ~n39829 ;
  assign y22891 = ~1'b0 ;
  assign y22892 = n39833 ;
  assign y22893 = n757 ;
  assign y22894 = n39835 ;
  assign y22895 = ~n39838 ;
  assign y22896 = n26240 ;
  assign y22897 = ~1'b0 ;
  assign y22898 = n39840 ;
  assign y22899 = ~n39845 ;
  assign y22900 = ~n39846 ;
  assign y22901 = n39850 ;
  assign y22902 = ~1'b0 ;
  assign y22903 = ~1'b0 ;
  assign y22904 = n39853 ;
  assign y22905 = ~n39855 ;
  assign y22906 = ~n39858 ;
  assign y22907 = 1'b0 ;
  assign y22908 = n29871 ;
  assign y22909 = n39860 ;
  assign y22910 = 1'b0 ;
  assign y22911 = ~n39866 ;
  assign y22912 = n39876 ;
  assign y22913 = n39878 ;
  assign y22914 = ~n39880 ;
  assign y22915 = ~1'b0 ;
  assign y22916 = ~1'b0 ;
  assign y22917 = ~n39881 ;
  assign y22918 = 1'b0 ;
  assign y22919 = n39882 ;
  assign y22920 = ~n39885 ;
  assign y22921 = ~1'b0 ;
  assign y22922 = ~1'b0 ;
  assign y22923 = n39888 ;
  assign y22924 = ~n39891 ;
  assign y22925 = ~n39892 ;
  assign y22926 = ~n39893 ;
  assign y22927 = ~1'b0 ;
  assign y22928 = ~n39896 ;
  assign y22929 = ~1'b0 ;
  assign y22930 = n39898 ;
  assign y22931 = ~n39901 ;
  assign y22932 = ~1'b0 ;
  assign y22933 = n39903 ;
  assign y22934 = ~1'b0 ;
  assign y22935 = n39904 ;
  assign y22936 = ~n39905 ;
  assign y22937 = n39906 ;
  assign y22938 = ~1'b0 ;
  assign y22939 = n39907 ;
  assign y22940 = ~n14226 ;
  assign y22941 = ~1'b0 ;
  assign y22942 = n39908 ;
  assign y22943 = ~1'b0 ;
  assign y22944 = n27616 ;
  assign y22945 = ~n39911 ;
  assign y22946 = n39914 ;
  assign y22947 = ~n39916 ;
  assign y22948 = n39917 ;
  assign y22949 = n39918 ;
  assign y22950 = ~1'b0 ;
  assign y22951 = n39921 ;
  assign y22952 = ~n39922 ;
  assign y22953 = n11696 ;
  assign y22954 = ~n39927 ;
  assign y22955 = ~n39929 ;
  assign y22956 = ~n18066 ;
  assign y22957 = n39930 ;
  assign y22958 = ~1'b0 ;
  assign y22959 = ~1'b0 ;
  assign y22960 = ~n39932 ;
  assign y22961 = n39942 ;
  assign y22962 = ~n39946 ;
  assign y22963 = n39947 ;
  assign y22964 = ~1'b0 ;
  assign y22965 = ~n39950 ;
  assign y22966 = ~n39952 ;
  assign y22967 = n39956 ;
  assign y22968 = ~n11614 ;
  assign y22969 = n23859 ;
  assign y22970 = ~1'b0 ;
  assign y22971 = ~1'b0 ;
  assign y22972 = ~n39958 ;
  assign y22973 = ~n39959 ;
  assign y22974 = n39960 ;
  assign y22975 = n39961 ;
  assign y22976 = ~1'b0 ;
  assign y22977 = ~n39962 ;
  assign y22978 = ~1'b0 ;
  assign y22979 = 1'b0 ;
  assign y22980 = ~n39964 ;
  assign y22981 = ~1'b0 ;
  assign y22982 = n39966 ;
  assign y22983 = n39969 ;
  assign y22984 = n39973 ;
  assign y22985 = ~1'b0 ;
  assign y22986 = ~1'b0 ;
  assign y22987 = ~n39975 ;
  assign y22988 = ~n39976 ;
  assign y22989 = ~1'b0 ;
  assign y22990 = ~n39978 ;
  assign y22991 = ~n39980 ;
  assign y22992 = ~1'b0 ;
  assign y22993 = n39983 ;
  assign y22994 = ~n39986 ;
  assign y22995 = ~1'b0 ;
  assign y22996 = n39989 ;
  assign y22997 = ~n39990 ;
  assign y22998 = ~n39992 ;
  assign y22999 = ~1'b0 ;
  assign y23000 = ~1'b0 ;
  assign y23001 = n39993 ;
  assign y23002 = ~n39995 ;
  assign y23003 = ~1'b0 ;
  assign y23004 = ~1'b0 ;
  assign y23005 = ~1'b0 ;
  assign y23006 = n39996 ;
  assign y23007 = n39999 ;
  assign y23008 = ~n40001 ;
  assign y23009 = ~n7979 ;
  assign y23010 = n40006 ;
  assign y23011 = n40008 ;
  assign y23012 = n40009 ;
  assign y23013 = ~1'b0 ;
  assign y23014 = n40010 ;
  assign y23015 = ~1'b0 ;
  assign y23016 = ~1'b0 ;
  assign y23017 = ~1'b0 ;
  assign y23018 = n40011 ;
  assign y23019 = n40013 ;
  assign y23020 = ~1'b0 ;
  assign y23021 = ~n40017 ;
  assign y23022 = n40018 ;
  assign y23023 = ~1'b0 ;
  assign y23024 = ~1'b0 ;
  assign y23025 = ~n40021 ;
  assign y23026 = ~1'b0 ;
  assign y23027 = n13961 ;
  assign y23028 = n40022 ;
  assign y23029 = ~1'b0 ;
  assign y23030 = n40023 ;
  assign y23031 = n40024 ;
  assign y23032 = ~n40025 ;
  assign y23033 = ~n40028 ;
  assign y23034 = ~1'b0 ;
  assign y23035 = n40031 ;
  assign y23036 = ~n40032 ;
  assign y23037 = ~1'b0 ;
  assign y23038 = ~1'b0 ;
  assign y23039 = n40034 ;
  assign y23040 = ~1'b0 ;
  assign y23041 = ~n40035 ;
  assign y23042 = ~n40037 ;
  assign y23043 = ~n40038 ;
  assign y23044 = ~n40043 ;
  assign y23045 = n40046 ;
  assign y23046 = ~n40048 ;
  assign y23047 = n40054 ;
  assign y23048 = n40056 ;
  assign y23049 = ~n40057 ;
  assign y23050 = ~1'b0 ;
  assign y23051 = ~1'b0 ;
  assign y23052 = ~1'b0 ;
  assign y23053 = ~1'b0 ;
  assign y23054 = n40058 ;
  assign y23055 = n40061 ;
  assign y23056 = ~n40063 ;
  assign y23057 = ~n40067 ;
  assign y23058 = ~1'b0 ;
  assign y23059 = n40071 ;
  assign y23060 = n40072 ;
  assign y23061 = n40081 ;
  assign y23062 = n40084 ;
  assign y23063 = n40086 ;
  assign y23064 = n40087 ;
  assign y23065 = ~1'b0 ;
  assign y23066 = ~n40091 ;
  assign y23067 = ~n40097 ;
  assign y23068 = ~n40099 ;
  assign y23069 = ~n40102 ;
  assign y23070 = ~1'b0 ;
  assign y23071 = ~1'b0 ;
  assign y23072 = n40103 ;
  assign y23073 = ~n40107 ;
  assign y23074 = n40109 ;
  assign y23075 = n40111 ;
  assign y23076 = ~1'b0 ;
  assign y23077 = ~1'b0 ;
  assign y23078 = n40113 ;
  assign y23079 = ~n40114 ;
  assign y23080 = ~1'b0 ;
  assign y23081 = ~n40116 ;
  assign y23082 = 1'b0 ;
  assign y23083 = ~1'b0 ;
  assign y23084 = n40117 ;
  assign y23085 = n27721 ;
  assign y23086 = ~1'b0 ;
  assign y23087 = ~n40124 ;
  assign y23088 = ~n40126 ;
  assign y23089 = n40128 ;
  assign y23090 = ~n40130 ;
  assign y23091 = ~n40132 ;
  assign y23092 = ~1'b0 ;
  assign y23093 = ~n40135 ;
  assign y23094 = n40136 ;
  assign y23095 = ~1'b0 ;
  assign y23096 = ~n24057 ;
  assign y23097 = ~1'b0 ;
  assign y23098 = ~n40139 ;
  assign y23099 = n40140 ;
  assign y23100 = n40142 ;
  assign y23101 = ~1'b0 ;
  assign y23102 = ~1'b0 ;
  assign y23103 = n40143 ;
  assign y23104 = ~n29964 ;
  assign y23105 = n40145 ;
  assign y23106 = ~n18424 ;
  assign y23107 = n40147 ;
  assign y23108 = n40149 ;
  assign y23109 = ~1'b0 ;
  assign y23110 = ~n12763 ;
  assign y23111 = ~1'b0 ;
  assign y23112 = ~1'b0 ;
  assign y23113 = n40150 ;
  assign y23114 = ~n40151 ;
  assign y23115 = ~n40152 ;
  assign y23116 = n40154 ;
  assign y23117 = n40157 ;
  assign y23118 = n40158 ;
  assign y23119 = n40161 ;
  assign y23120 = ~1'b0 ;
  assign y23121 = 1'b0 ;
  assign y23122 = n40162 ;
  assign y23123 = 1'b0 ;
  assign y23124 = ~n40163 ;
  assign y23125 = ~1'b0 ;
  assign y23126 = ~1'b0 ;
  assign y23127 = ~n40164 ;
  assign y23128 = ~n40169 ;
  assign y23129 = ~n40171 ;
  assign y23130 = ~1'b0 ;
  assign y23131 = ~1'b0 ;
  assign y23132 = ~n40172 ;
  assign y23133 = n40173 ;
  assign y23134 = ~n40178 ;
  assign y23135 = n40181 ;
  assign y23136 = n9765 ;
  assign y23137 = ~1'b0 ;
  assign y23138 = ~1'b0 ;
  assign y23139 = ~1'b0 ;
  assign y23140 = ~n40183 ;
  assign y23141 = n21836 ;
  assign y23142 = ~1'b0 ;
  assign y23143 = ~n40185 ;
  assign y23144 = ~1'b0 ;
  assign y23145 = ~n40189 ;
  assign y23146 = ~n40191 ;
  assign y23147 = ~1'b0 ;
  assign y23148 = ~1'b0 ;
  assign y23149 = ~n40192 ;
  assign y23150 = ~n40193 ;
  assign y23151 = ~1'b0 ;
  assign y23152 = ~n40194 ;
  assign y23153 = n40196 ;
  assign y23154 = ~n40198 ;
  assign y23155 = ~1'b0 ;
  assign y23156 = ~1'b0 ;
  assign y23157 = ~n40200 ;
  assign y23158 = n40203 ;
  assign y23159 = ~n40204 ;
  assign y23160 = ~1'b0 ;
  assign y23161 = ~n40205 ;
  assign y23162 = ~1'b0 ;
  assign y23163 = ~1'b0 ;
  assign y23164 = ~1'b0 ;
  assign y23165 = ~n40207 ;
  assign y23166 = ~n40210 ;
  assign y23167 = n40211 ;
  assign y23168 = ~n14044 ;
  assign y23169 = ~n29374 ;
  assign y23170 = n40214 ;
  assign y23171 = n40217 ;
  assign y23172 = ~n40218 ;
  assign y23173 = n40219 ;
  assign y23174 = ~1'b0 ;
  assign y23175 = n40220 ;
  assign y23176 = n40226 ;
  assign y23177 = ~1'b0 ;
  assign y23178 = n18834 ;
  assign y23179 = ~1'b0 ;
  assign y23180 = ~n40229 ;
  assign y23181 = ~n36848 ;
  assign y23182 = n40231 ;
  assign y23183 = ~n36941 ;
  assign y23184 = n40233 ;
  assign y23185 = 1'b0 ;
  assign y23186 = ~n40237 ;
  assign y23187 = ~n40238 ;
  assign y23188 = ~1'b0 ;
  assign y23189 = ~n40239 ;
  assign y23190 = ~1'b0 ;
  assign y23191 = n40240 ;
  assign y23192 = ~1'b0 ;
  assign y23193 = ~1'b0 ;
  assign y23194 = ~n40241 ;
  assign y23195 = ~1'b0 ;
  assign y23196 = ~n40246 ;
  assign y23197 = ~n40247 ;
  assign y23198 = ~n40249 ;
  assign y23199 = ~n40250 ;
  assign y23200 = ~1'b0 ;
  assign y23201 = n6774 ;
  assign y23202 = ~1'b0 ;
  assign y23203 = n28220 ;
  assign y23204 = ~1'b0 ;
  assign y23205 = n40254 ;
  assign y23206 = n40258 ;
  assign y23207 = n40261 ;
  assign y23208 = n40265 ;
  assign y23209 = ~n40267 ;
  assign y23210 = ~1'b0 ;
  assign y23211 = n40268 ;
  assign y23212 = ~1'b0 ;
  assign y23213 = ~1'b0 ;
  assign y23214 = ~1'b0 ;
  assign y23215 = n40272 ;
  assign y23216 = ~1'b0 ;
  assign y23217 = n40274 ;
  assign y23218 = 1'b0 ;
  assign y23219 = ~n40277 ;
  assign y23220 = ~n40280 ;
  assign y23221 = ~n40281 ;
  assign y23222 = n6933 ;
  assign y23223 = ~1'b0 ;
  assign y23224 = n40283 ;
  assign y23225 = ~1'b0 ;
  assign y23226 = n40288 ;
  assign y23227 = ~1'b0 ;
  assign y23228 = ~n40289 ;
  assign y23229 = n40290 ;
  assign y23230 = ~n40296 ;
  assign y23231 = ~1'b0 ;
  assign y23232 = n40297 ;
  assign y23233 = ~1'b0 ;
  assign y23234 = ~n40299 ;
  assign y23235 = ~1'b0 ;
  assign y23236 = n40300 ;
  assign y23237 = ~n40302 ;
  assign y23238 = n40306 ;
  assign y23239 = ~n40308 ;
  assign y23240 = ~1'b0 ;
  assign y23241 = ~n40310 ;
  assign y23242 = ~n40314 ;
  assign y23243 = ~n40316 ;
  assign y23244 = ~n40317 ;
  assign y23245 = n26098 ;
  assign y23246 = ~n40318 ;
  assign y23247 = ~n40319 ;
  assign y23248 = n40321 ;
  assign y23249 = ~1'b0 ;
  assign y23250 = ~1'b0 ;
  assign y23251 = ~n40322 ;
  assign y23252 = ~n23065 ;
  assign y23253 = ~1'b0 ;
  assign y23254 = ~1'b0 ;
  assign y23255 = n40323 ;
  assign y23256 = ~n40330 ;
  assign y23257 = ~n40331 ;
  assign y23258 = n40332 ;
  assign y23259 = ~n40335 ;
  assign y23260 = ~1'b0 ;
  assign y23261 = n40337 ;
  assign y23262 = ~n40338 ;
  assign y23263 = ~n40342 ;
  assign y23264 = ~n21034 ;
  assign y23265 = ~n40346 ;
  assign y23266 = ~1'b0 ;
  assign y23267 = ~n40352 ;
  assign y23268 = n40356 ;
  assign y23269 = ~n40359 ;
  assign y23270 = n40361 ;
  assign y23271 = ~1'b0 ;
  assign y23272 = n40362 ;
  assign y23273 = ~n6256 ;
  assign y23274 = n40366 ;
  assign y23275 = ~1'b0 ;
  assign y23276 = ~n40369 ;
  assign y23277 = ~n40372 ;
  assign y23278 = ~1'b0 ;
  assign y23279 = ~1'b0 ;
  assign y23280 = ~1'b0 ;
  assign y23281 = n25092 ;
  assign y23282 = ~1'b0 ;
  assign y23283 = ~1'b0 ;
  assign y23284 = n40374 ;
  assign y23285 = ~1'b0 ;
  assign y23286 = n40379 ;
  assign y23287 = ~n40383 ;
  assign y23288 = ~n40388 ;
  assign y23289 = ~1'b0 ;
  assign y23290 = ~n40390 ;
  assign y23291 = ~n40392 ;
  assign y23292 = n40394 ;
  assign y23293 = ~1'b0 ;
  assign y23294 = ~n40395 ;
  assign y23295 = ~n22598 ;
  assign y23296 = n40396 ;
  assign y23297 = ~n40398 ;
  assign y23298 = n40402 ;
  assign y23299 = n40404 ;
  assign y23300 = ~n25389 ;
  assign y23301 = ~1'b0 ;
  assign y23302 = ~n40405 ;
  assign y23303 = n40408 ;
  assign y23304 = ~n40409 ;
  assign y23305 = ~1'b0 ;
  assign y23306 = ~1'b0 ;
  assign y23307 = ~1'b0 ;
  assign y23308 = ~1'b0 ;
  assign y23309 = ~n40410 ;
  assign y23310 = ~1'b0 ;
  assign y23311 = ~n40411 ;
  assign y23312 = ~n6114 ;
  assign y23313 = ~1'b0 ;
  assign y23314 = ~n40413 ;
  assign y23315 = n40414 ;
  assign y23316 = n14817 ;
  assign y23317 = ~1'b0 ;
  assign y23318 = ~1'b0 ;
  assign y23319 = ~1'b0 ;
  assign y23320 = n40419 ;
  assign y23321 = n40421 ;
  assign y23322 = ~n40423 ;
  assign y23323 = 1'b0 ;
  assign y23324 = ~n40424 ;
  assign y23325 = ~n40427 ;
  assign y23326 = ~n40431 ;
  assign y23327 = ~1'b0 ;
  assign y23328 = ~n40436 ;
  assign y23329 = n40437 ;
  assign y23330 = n40440 ;
  assign y23331 = n40448 ;
  assign y23332 = n40451 ;
  assign y23333 = n40453 ;
  assign y23334 = ~n25968 ;
  assign y23335 = ~1'b0 ;
  assign y23336 = n40457 ;
  assign y23337 = ~n40458 ;
  assign y23338 = ~n40459 ;
  assign y23339 = ~n40460 ;
  assign y23340 = ~n31010 ;
  assign y23341 = ~1'b0 ;
  assign y23342 = ~n40464 ;
  assign y23343 = n40465 ;
  assign y23344 = n28032 ;
  assign y23345 = ~1'b0 ;
  assign y23346 = n40468 ;
  assign y23347 = ~n40469 ;
  assign y23348 = ~n40470 ;
  assign y23349 = ~n40472 ;
  assign y23350 = n40473 ;
  assign y23351 = n40478 ;
  assign y23352 = 1'b0 ;
  assign y23353 = n40482 ;
  assign y23354 = n40484 ;
  assign y23355 = ~n40485 ;
  assign y23356 = ~n40488 ;
  assign y23357 = ~1'b0 ;
  assign y23358 = ~n40489 ;
  assign y23359 = ~1'b0 ;
  assign y23360 = n34264 ;
  assign y23361 = ~1'b0 ;
  assign y23362 = ~n40490 ;
  assign y23363 = n15938 ;
  assign y23364 = n40493 ;
  assign y23365 = ~1'b0 ;
  assign y23366 = ~1'b0 ;
  assign y23367 = ~1'b0 ;
  assign y23368 = ~1'b0 ;
  assign y23369 = n40494 ;
  assign y23370 = n40498 ;
  assign y23371 = ~n40505 ;
  assign y23372 = ~1'b0 ;
  assign y23373 = n40507 ;
  assign y23374 = n40508 ;
  assign y23375 = ~n40513 ;
  assign y23376 = ~n40516 ;
  assign y23377 = ~n40521 ;
  assign y23378 = n35101 ;
  assign y23379 = ~1'b0 ;
  assign y23380 = ~1'b0 ;
  assign y23381 = n40524 ;
  assign y23382 = n40525 ;
  assign y23383 = n40526 ;
  assign y23384 = ~n40527 ;
  assign y23385 = ~n40528 ;
  assign y23386 = ~n40530 ;
  assign y23387 = ~1'b0 ;
  assign y23388 = ~1'b0 ;
  assign y23389 = ~1'b0 ;
  assign y23390 = n11338 ;
  assign y23391 = n40534 ;
  assign y23392 = ~n40535 ;
  assign y23393 = n40537 ;
  assign y23394 = n40539 ;
  assign y23395 = n40541 ;
  assign y23396 = n40544 ;
  assign y23397 = ~1'b0 ;
  assign y23398 = ~n40547 ;
  assign y23399 = ~n40551 ;
  assign y23400 = ~n40554 ;
  assign y23401 = ~n155 ;
  assign y23402 = ~n3063 ;
  assign y23403 = ~n40557 ;
  assign y23404 = 1'b0 ;
  assign y23405 = n40558 ;
  assign y23406 = ~1'b0 ;
  assign y23407 = ~1'b0 ;
  assign y23408 = ~1'b0 ;
  assign y23409 = n40560 ;
  assign y23410 = n40562 ;
  assign y23411 = n40564 ;
  assign y23412 = ~1'b0 ;
  assign y23413 = ~n40569 ;
  assign y23414 = n3646 ;
  assign y23415 = ~n33009 ;
  assign y23416 = n40572 ;
  assign y23417 = n40574 ;
  assign y23418 = ~n40581 ;
  assign y23419 = ~n40582 ;
  assign y23420 = ~n40583 ;
  assign y23421 = ~1'b0 ;
  assign y23422 = n40590 ;
  assign y23423 = n40592 ;
  assign y23424 = ~n40594 ;
  assign y23425 = ~1'b0 ;
  assign y23426 = ~n40596 ;
  assign y23427 = n40609 ;
  assign y23428 = ~n40612 ;
  assign y23429 = ~1'b0 ;
  assign y23430 = ~n40613 ;
  assign y23431 = n11008 ;
  assign y23432 = n40615 ;
  assign y23433 = ~n40620 ;
  assign y23434 = ~1'b0 ;
  assign y23435 = n17735 ;
  assign y23436 = ~1'b0 ;
  assign y23437 = ~1'b0 ;
  assign y23438 = ~n40621 ;
  assign y23439 = n40623 ;
  assign y23440 = ~1'b0 ;
  assign y23441 = ~1'b0 ;
  assign y23442 = ~1'b0 ;
  assign y23443 = ~n40624 ;
  assign y23444 = ~1'b0 ;
  assign y23445 = ~1'b0 ;
  assign y23446 = n40627 ;
  assign y23447 = ~n40630 ;
  assign y23448 = ~n40637 ;
  assign y23449 = ~1'b0 ;
  assign y23450 = ~n40639 ;
  assign y23451 = n40641 ;
  assign y23452 = ~n2380 ;
  assign y23453 = n40642 ;
  assign y23454 = ~n40643 ;
  assign y23455 = ~n40647 ;
  assign y23456 = ~n40648 ;
  assign y23457 = n40652 ;
  assign y23458 = ~1'b0 ;
  assign y23459 = n40654 ;
  assign y23460 = ~n40657 ;
  assign y23461 = ~1'b0 ;
  assign y23462 = ~1'b0 ;
  assign y23463 = ~n40658 ;
  assign y23464 = n40659 ;
  assign y23465 = ~1'b0 ;
  assign y23466 = ~1'b0 ;
  assign y23467 = n40663 ;
  assign y23468 = ~1'b0 ;
  assign y23469 = ~n40678 ;
  assign y23470 = ~n40679 ;
  assign y23471 = ~1'b0 ;
  assign y23472 = n11485 ;
  assign y23473 = n38345 ;
  assign y23474 = 1'b0 ;
  assign y23475 = n40680 ;
  assign y23476 = ~n40682 ;
  assign y23477 = n40687 ;
  assign y23478 = ~1'b0 ;
  assign y23479 = ~n8425 ;
  assign y23480 = ~1'b0 ;
  assign y23481 = ~n40688 ;
  assign y23482 = n40690 ;
  assign y23483 = ~n40691 ;
  assign y23484 = ~n19164 ;
  assign y23485 = ~n40692 ;
  assign y23486 = ~1'b0 ;
  assign y23487 = ~1'b0 ;
  assign y23488 = n40693 ;
  assign y23489 = n40694 ;
  assign y23490 = ~1'b0 ;
  assign y23491 = ~n40698 ;
  assign y23492 = ~n40703 ;
  assign y23493 = ~1'b0 ;
  assign y23494 = ~1'b0 ;
  assign y23495 = n40705 ;
  assign y23496 = ~n40708 ;
  assign y23497 = n40710 ;
  assign y23498 = ~n40713 ;
  assign y23499 = 1'b0 ;
  assign y23500 = ~1'b0 ;
  assign y23501 = n40718 ;
  assign y23502 = ~1'b0 ;
  assign y23503 = n40721 ;
  assign y23504 = ~n40722 ;
  assign y23505 = n40723 ;
  assign y23506 = ~n40728 ;
  assign y23507 = n40730 ;
  assign y23508 = ~n40735 ;
  assign y23509 = ~n40738 ;
  assign y23510 = ~n40739 ;
  assign y23511 = ~1'b0 ;
  assign y23512 = n40742 ;
  assign y23513 = ~n40745 ;
  assign y23514 = ~n40746 ;
  assign y23515 = ~n40749 ;
  assign y23516 = ~n40752 ;
  assign y23517 = ~n40756 ;
  assign y23518 = ~1'b0 ;
  assign y23519 = n40758 ;
  assign y23520 = n40761 ;
  assign y23521 = ~n40763 ;
  assign y23522 = n6663 ;
  assign y23523 = n40766 ;
  assign y23524 = ~1'b0 ;
  assign y23525 = ~n40767 ;
  assign y23526 = ~n40769 ;
  assign y23527 = ~1'b0 ;
  assign y23528 = 1'b0 ;
  assign y23529 = n40771 ;
  assign y23530 = n40772 ;
  assign y23531 = ~1'b0 ;
  assign y23532 = ~n40773 ;
  assign y23533 = n40774 ;
  assign y23534 = ~1'b0 ;
  assign y23535 = ~1'b0 ;
  assign y23536 = n40775 ;
  assign y23537 = n40777 ;
  assign y23538 = n40779 ;
  assign y23539 = n40784 ;
  assign y23540 = n40786 ;
  assign y23541 = ~1'b0 ;
  assign y23542 = ~1'b0 ;
  assign y23543 = n340 ;
  assign y23544 = ~n40790 ;
  assign y23545 = ~n40792 ;
  assign y23546 = ~n22900 ;
  assign y23547 = ~1'b0 ;
  assign y23548 = n8227 ;
  assign y23549 = n40795 ;
  assign y23550 = ~n24079 ;
  assign y23551 = ~n40801 ;
  assign y23552 = ~n40805 ;
  assign y23553 = ~n40806 ;
  assign y23554 = ~n40808 ;
  assign y23555 = ~n40817 ;
  assign y23556 = 1'b0 ;
  assign y23557 = n40818 ;
  assign y23558 = n40821 ;
  assign y23559 = ~n40823 ;
  assign y23560 = ~n30343 ;
  assign y23561 = n40825 ;
  assign y23562 = ~n9167 ;
  assign y23563 = n40826 ;
  assign y23564 = ~n40827 ;
  assign y23565 = ~n40829 ;
  assign y23566 = ~n40839 ;
  assign y23567 = ~n40840 ;
  assign y23568 = ~1'b0 ;
  assign y23569 = ~n40843 ;
  assign y23570 = ~n26024 ;
  assign y23571 = ~1'b0 ;
  assign y23572 = ~1'b0 ;
  assign y23573 = n40844 ;
  assign y23574 = n40845 ;
  assign y23575 = ~1'b0 ;
  assign y23576 = ~n15096 ;
  assign y23577 = ~1'b0 ;
  assign y23578 = n40849 ;
  assign y23579 = n40854 ;
  assign y23580 = n40855 ;
  assign y23581 = ~n40856 ;
  assign y23582 = n40857 ;
  assign y23583 = ~1'b0 ;
  assign y23584 = ~n40859 ;
  assign y23585 = ~n40864 ;
  assign y23586 = ~1'b0 ;
  assign y23587 = ~1'b0 ;
  assign y23588 = ~n40866 ;
  assign y23589 = n40871 ;
  assign y23590 = n40873 ;
  assign y23591 = ~1'b0 ;
  assign y23592 = ~1'b0 ;
  assign y23593 = n40874 ;
  assign y23594 = 1'b0 ;
  assign y23595 = ~n40875 ;
  assign y23596 = ~1'b0 ;
  assign y23597 = ~n40881 ;
  assign y23598 = n40882 ;
  assign y23599 = ~n40883 ;
  assign y23600 = ~1'b0 ;
  assign y23601 = ~n40887 ;
  assign y23602 = ~n4379 ;
  assign y23603 = ~1'b0 ;
  assign y23604 = n40888 ;
  assign y23605 = n40891 ;
  assign y23606 = ~1'b0 ;
  assign y23607 = ~1'b0 ;
  assign y23608 = ~n40893 ;
  assign y23609 = ~1'b0 ;
  assign y23610 = ~n40894 ;
  assign y23611 = ~1'b0 ;
  assign y23612 = n40896 ;
  assign y23613 = ~n40898 ;
  assign y23614 = n40900 ;
  assign y23615 = ~n40902 ;
  assign y23616 = ~n40903 ;
  assign y23617 = ~1'b0 ;
  assign y23618 = n40905 ;
  assign y23619 = ~n40907 ;
  assign y23620 = ~n40908 ;
  assign y23621 = ~1'b0 ;
  assign y23622 = ~n40909 ;
  assign y23623 = n40910 ;
  assign y23624 = n2050 ;
  assign y23625 = n40911 ;
  assign y23626 = ~n40913 ;
  assign y23627 = ~n40915 ;
  assign y23628 = n40916 ;
  assign y23629 = n40918 ;
  assign y23630 = ~1'b0 ;
  assign y23631 = ~1'b0 ;
  assign y23632 = ~n40920 ;
  assign y23633 = ~1'b0 ;
  assign y23634 = ~1'b0 ;
  assign y23635 = ~1'b0 ;
  assign y23636 = ~n40923 ;
  assign y23637 = n40924 ;
  assign y23638 = ~1'b0 ;
  assign y23639 = ~n40927 ;
  assign y23640 = n40928 ;
  assign y23641 = n40929 ;
  assign y23642 = ~1'b0 ;
  assign y23643 = ~n40930 ;
  assign y23644 = n40933 ;
  assign y23645 = n40935 ;
  assign y23646 = ~n40937 ;
  assign y23647 = ~1'b0 ;
  assign y23648 = ~n40939 ;
  assign y23649 = ~1'b0 ;
  assign y23650 = ~1'b0 ;
  assign y23651 = n40941 ;
  assign y23652 = ~1'b0 ;
  assign y23653 = ~1'b0 ;
  assign y23654 = ~n40943 ;
  assign y23655 = ~n40944 ;
  assign y23656 = ~1'b0 ;
  assign y23657 = ~n40947 ;
  assign y23658 = ~1'b0 ;
  assign y23659 = n40949 ;
  assign y23660 = ~1'b0 ;
  assign y23661 = ~1'b0 ;
  assign y23662 = ~1'b0 ;
  assign y23663 = ~1'b0 ;
  assign y23664 = n28099 ;
  assign y23665 = ~n40950 ;
  assign y23666 = n40951 ;
  assign y23667 = n40952 ;
  assign y23668 = n40955 ;
  assign y23669 = ~n40960 ;
  assign y23670 = ~1'b0 ;
  assign y23671 = n40964 ;
  assign y23672 = ~n40965 ;
  assign y23673 = n40969 ;
  assign y23674 = ~n40971 ;
  assign y23675 = ~n40973 ;
  assign y23676 = n40974 ;
  assign y23677 = ~1'b0 ;
  assign y23678 = n40977 ;
  assign y23679 = ~n40983 ;
  assign y23680 = n40984 ;
  assign y23681 = ~1'b0 ;
  assign y23682 = n40985 ;
  assign y23683 = n40987 ;
  assign y23684 = ~1'b0 ;
  assign y23685 = n40990 ;
  assign y23686 = ~n40992 ;
  assign y23687 = n40993 ;
  assign y23688 = ~n32268 ;
  assign y23689 = ~1'b0 ;
  assign y23690 = n40671 ;
  assign y23691 = n40994 ;
  assign y23692 = ~1'b0 ;
  assign y23693 = n40996 ;
  assign y23694 = ~n40999 ;
  assign y23695 = ~1'b0 ;
  assign y23696 = n41001 ;
  assign y23697 = ~1'b0 ;
  assign y23698 = ~1'b0 ;
  assign y23699 = n41002 ;
  assign y23700 = ~n41003 ;
  assign y23701 = ~n41005 ;
  assign y23702 = ~n41009 ;
  assign y23703 = n41010 ;
  assign y23704 = ~n41012 ;
  assign y23705 = ~n41016 ;
  assign y23706 = ~1'b0 ;
  assign y23707 = ~1'b0 ;
  assign y23708 = ~1'b0 ;
  assign y23709 = 1'b0 ;
  assign y23710 = ~n41018 ;
  assign y23711 = n41020 ;
  assign y23712 = ~1'b0 ;
  assign y23713 = ~n41023 ;
  assign y23714 = ~n41024 ;
  assign y23715 = n41026 ;
  assign y23716 = ~1'b0 ;
  assign y23717 = ~n41029 ;
  assign y23718 = n41031 ;
  assign y23719 = n41032 ;
  assign y23720 = ~n41034 ;
  assign y23721 = ~n41036 ;
  assign y23722 = ~n41037 ;
  assign y23723 = ~n41038 ;
  assign y23724 = ~1'b0 ;
  assign y23725 = ~1'b0 ;
  assign y23726 = n41040 ;
  assign y23727 = ~n41044 ;
  assign y23728 = ~n41046 ;
  assign y23729 = n41048 ;
  assign y23730 = n41052 ;
  assign y23731 = ~n41053 ;
  assign y23732 = ~n41054 ;
  assign y23733 = ~n41055 ;
  assign y23734 = ~1'b0 ;
  assign y23735 = ~n41058 ;
  assign y23736 = ~1'b0 ;
  assign y23737 = n35622 ;
  assign y23738 = 1'b0 ;
  assign y23739 = ~n41061 ;
  assign y23740 = n41062 ;
  assign y23741 = ~n565 ;
  assign y23742 = n41064 ;
  assign y23743 = ~1'b0 ;
  assign y23744 = n41065 ;
  assign y23745 = 1'b0 ;
  assign y23746 = n41067 ;
  assign y23747 = ~1'b0 ;
  assign y23748 = n41071 ;
  assign y23749 = ~n41072 ;
  assign y23750 = n41076 ;
  assign y23751 = ~1'b0 ;
  assign y23752 = ~n41077 ;
  assign y23753 = ~1'b0 ;
  assign y23754 = ~n41079 ;
  assign y23755 = n41080 ;
  assign y23756 = n41084 ;
  assign y23757 = ~n41085 ;
  assign y23758 = ~1'b0 ;
  assign y23759 = n41086 ;
  assign y23760 = ~1'b0 ;
  assign y23761 = n41088 ;
  assign y23762 = ~1'b0 ;
  assign y23763 = n41091 ;
  assign y23764 = n41093 ;
  assign y23765 = ~n41095 ;
  assign y23766 = ~n41096 ;
  assign y23767 = ~n41098 ;
  assign y23768 = ~1'b0 ;
  assign y23769 = ~n41100 ;
  assign y23770 = ~n41102 ;
  assign y23771 = ~n41103 ;
  assign y23772 = ~1'b0 ;
  assign y23773 = ~1'b0 ;
  assign y23774 = ~1'b0 ;
  assign y23775 = ~n41107 ;
  assign y23776 = ~1'b0 ;
  assign y23777 = ~n41108 ;
  assign y23778 = ~1'b0 ;
  assign y23779 = ~n41110 ;
  assign y23780 = ~1'b0 ;
  assign y23781 = n41113 ;
  assign y23782 = ~n41114 ;
  assign y23783 = n34696 ;
  assign y23784 = n41115 ;
  assign y23785 = ~1'b0 ;
  assign y23786 = ~n41118 ;
  assign y23787 = ~1'b0 ;
  assign y23788 = ~n41121 ;
  assign y23789 = ~1'b0 ;
  assign y23790 = n41123 ;
  assign y23791 = ~1'b0 ;
  assign y23792 = ~n41126 ;
  assign y23793 = ~n41129 ;
  assign y23794 = ~n41132 ;
  assign y23795 = n41138 ;
  assign y23796 = ~1'b0 ;
  assign y23797 = n41144 ;
  assign y23798 = n28901 ;
  assign y23799 = ~1'b0 ;
  assign y23800 = ~1'b0 ;
  assign y23801 = n41145 ;
  assign y23802 = n41146 ;
  assign y23803 = ~n41147 ;
  assign y23804 = ~1'b0 ;
  assign y23805 = ~1'b0 ;
  assign y23806 = ~n41149 ;
  assign y23807 = n32113 ;
  assign y23808 = n6895 ;
  assign y23809 = ~1'b0 ;
  assign y23810 = n41156 ;
  assign y23811 = ~n41157 ;
  assign y23812 = n41158 ;
  assign y23813 = ~n41162 ;
  assign y23814 = ~1'b0 ;
  assign y23815 = ~1'b0 ;
  assign y23816 = n41163 ;
  assign y23817 = n16192 ;
  assign y23818 = ~1'b0 ;
  assign y23819 = ~n41166 ;
  assign y23820 = ~n3763 ;
  assign y23821 = n41168 ;
  assign y23822 = 1'b0 ;
  assign y23823 = n41170 ;
  assign y23824 = ~1'b0 ;
  assign y23825 = ~n41172 ;
  assign y23826 = n41173 ;
  assign y23827 = n41174 ;
  assign y23828 = ~1'b0 ;
  assign y23829 = n41175 ;
  assign y23830 = ~1'b0 ;
  assign y23831 = n41176 ;
  assign y23832 = ~n41179 ;
  assign y23833 = ~n41182 ;
  assign y23834 = ~n9215 ;
  assign y23835 = n41184 ;
  assign y23836 = ~1'b0 ;
  assign y23837 = ~1'b0 ;
  assign y23838 = ~1'b0 ;
  assign y23839 = ~n41185 ;
  assign y23840 = ~1'b0 ;
  assign y23841 = ~n41187 ;
  assign y23842 = n41189 ;
  assign y23843 = n41194 ;
  assign y23844 = n41195 ;
  assign y23845 = n41197 ;
  assign y23846 = ~n41199 ;
  assign y23847 = ~1'b0 ;
  assign y23848 = ~1'b0 ;
  assign y23849 = n41200 ;
  assign y23850 = n41203 ;
  assign y23851 = ~n41204 ;
  assign y23852 = n41208 ;
  assign y23853 = ~n41211 ;
  assign y23854 = ~1'b0 ;
  assign y23855 = n41213 ;
  assign y23856 = n28812 ;
  assign y23857 = ~n41214 ;
  assign y23858 = ~n41217 ;
  assign y23859 = n41221 ;
  assign y23860 = ~1'b0 ;
  assign y23861 = ~n41224 ;
  assign y23862 = ~1'b0 ;
  assign y23863 = n41225 ;
  assign y23864 = n41226 ;
  assign y23865 = ~n41228 ;
  assign y23866 = n25097 ;
  assign y23867 = ~n41231 ;
  assign y23868 = n41236 ;
  assign y23869 = ~n41237 ;
  assign y23870 = n41238 ;
  assign y23871 = n41248 ;
  assign y23872 = ~1'b0 ;
  assign y23873 = ~1'b0 ;
  assign y23874 = ~1'b0 ;
  assign y23875 = n41250 ;
  assign y23876 = ~n23490 ;
  assign y23877 = ~1'b0 ;
  assign y23878 = n41251 ;
  assign y23879 = n41253 ;
  assign y23880 = ~n22524 ;
  assign y23881 = ~n41254 ;
  assign y23882 = n41256 ;
  assign y23883 = n41258 ;
  assign y23884 = n41259 ;
  assign y23885 = ~n41263 ;
  assign y23886 = 1'b0 ;
  assign y23887 = ~1'b0 ;
  assign y23888 = ~n41268 ;
  assign y23889 = ~n41269 ;
  assign y23890 = ~n1907 ;
  assign y23891 = ~1'b0 ;
  assign y23892 = ~n41270 ;
  assign y23893 = ~n41271 ;
  assign y23894 = ~n41275 ;
  assign y23895 = n41281 ;
  assign y23896 = 1'b0 ;
  assign y23897 = ~n41282 ;
  assign y23898 = ~1'b0 ;
  assign y23899 = n41283 ;
  assign y23900 = ~n8974 ;
  assign y23901 = ~1'b0 ;
  assign y23902 = ~1'b0 ;
  assign y23903 = ~n41285 ;
  assign y23904 = n41286 ;
  assign y23905 = n41288 ;
  assign y23906 = ~n41291 ;
  assign y23907 = ~1'b0 ;
  assign y23908 = ~1'b0 ;
  assign y23909 = ~n41292 ;
  assign y23910 = ~1'b0 ;
  assign y23911 = ~n41296 ;
  assign y23912 = n41298 ;
  assign y23913 = ~n41299 ;
  assign y23914 = n41302 ;
  assign y23915 = ~1'b0 ;
  assign y23916 = ~1'b0 ;
  assign y23917 = n41303 ;
  assign y23918 = ~n41305 ;
  assign y23919 = n5328 ;
  assign y23920 = n41307 ;
  assign y23921 = 1'b0 ;
  assign y23922 = ~1'b0 ;
  assign y23923 = ~n41308 ;
  assign y23924 = ~1'b0 ;
  assign y23925 = ~1'b0 ;
  assign y23926 = n41310 ;
  assign y23927 = n41314 ;
  assign y23928 = n41319 ;
  assign y23929 = ~n16360 ;
  assign y23930 = n41321 ;
  assign y23931 = ~1'b0 ;
  assign y23932 = ~1'b0 ;
  assign y23933 = ~n41328 ;
  assign y23934 = ~1'b0 ;
  assign y23935 = n41329 ;
  assign y23936 = n41330 ;
  assign y23937 = n41331 ;
  assign y23938 = ~n41332 ;
  assign y23939 = ~1'b0 ;
  assign y23940 = ~1'b0 ;
  assign y23941 = n38776 ;
  assign y23942 = ~1'b0 ;
  assign y23943 = ~n41334 ;
  assign y23944 = ~n41335 ;
  assign y23945 = ~n41339 ;
  assign y23946 = n41340 ;
  assign y23947 = n41341 ;
  assign y23948 = ~n41342 ;
  assign y23949 = 1'b0 ;
  assign y23950 = ~n41343 ;
  assign y23951 = ~n41348 ;
  assign y23952 = n41350 ;
  assign y23953 = ~1'b0 ;
  assign y23954 = ~n41355 ;
  assign y23955 = ~n41357 ;
  assign y23956 = n41359 ;
  assign y23957 = n41361 ;
  assign y23958 = n41364 ;
  assign y23959 = ~1'b0 ;
  assign y23960 = n41365 ;
  assign y23961 = n41366 ;
  assign y23962 = ~1'b0 ;
  assign y23963 = ~n41367 ;
  assign y23964 = n41368 ;
  assign y23965 = ~1'b0 ;
  assign y23966 = ~1'b0 ;
  assign y23967 = ~1'b0 ;
  assign y23968 = ~n41372 ;
  assign y23969 = ~1'b0 ;
  assign y23970 = n41375 ;
  assign y23971 = ~1'b0 ;
  assign y23972 = ~1'b0 ;
  assign y23973 = ~n41377 ;
  assign y23974 = n41378 ;
  assign y23975 = ~n41380 ;
  assign y23976 = ~1'b0 ;
  assign y23977 = ~n41383 ;
  assign y23978 = ~n41387 ;
  assign y23979 = 1'b0 ;
  assign y23980 = ~1'b0 ;
  assign y23981 = ~1'b0 ;
  assign y23982 = n41391 ;
  assign y23983 = n41397 ;
  assign y23984 = ~n17066 ;
  assign y23985 = ~n41401 ;
  assign y23986 = ~n41404 ;
  assign y23987 = n41407 ;
  assign y23988 = ~1'b0 ;
  assign y23989 = n41409 ;
  assign y23990 = ~n41411 ;
  assign y23991 = n41413 ;
  assign y23992 = ~1'b0 ;
  assign y23993 = n41414 ;
  assign y23994 = n41419 ;
  assign y23995 = n41423 ;
  assign y23996 = ~1'b0 ;
  assign y23997 = ~n41428 ;
  assign y23998 = 1'b0 ;
  assign y23999 = ~n41431 ;
  assign y24000 = n41438 ;
  assign y24001 = ~n41443 ;
  assign y24002 = n41444 ;
  assign y24003 = n41446 ;
  assign y24004 = ~n41447 ;
  assign y24005 = ~n41448 ;
  assign y24006 = ~1'b0 ;
  assign y24007 = ~n36622 ;
  assign y24008 = ~n41454 ;
  assign y24009 = ~n41456 ;
  assign y24010 = n41457 ;
  assign y24011 = ~n41460 ;
  assign y24012 = n41462 ;
  assign y24013 = 1'b0 ;
  assign y24014 = ~n41463 ;
  assign y24015 = ~n41464 ;
  assign y24016 = ~1'b0 ;
  assign y24017 = n41465 ;
  assign y24018 = ~n41468 ;
  assign y24019 = n41475 ;
  assign y24020 = n41478 ;
  assign y24021 = ~n41479 ;
  assign y24022 = ~n41481 ;
  assign y24023 = ~n41489 ;
  assign y24024 = n41491 ;
  assign y24025 = ~n41492 ;
  assign y24026 = ~n41498 ;
  assign y24027 = ~n18565 ;
  assign y24028 = ~n36468 ;
  assign y24029 = ~1'b0 ;
  assign y24030 = n41500 ;
  assign y24031 = n41503 ;
  assign y24032 = ~n5604 ;
  assign y24033 = n11378 ;
  assign y24034 = n41504 ;
  assign y24035 = ~n41505 ;
  assign y24036 = ~1'b0 ;
  assign y24037 = ~1'b0 ;
  assign y24038 = ~n41509 ;
  assign y24039 = ~1'b0 ;
  assign y24040 = ~n41511 ;
  assign y24041 = ~n41514 ;
  assign y24042 = ~1'b0 ;
  assign y24043 = n41515 ;
  assign y24044 = ~n41517 ;
  assign y24045 = ~n18458 ;
  assign y24046 = ~n41519 ;
  assign y24047 = n41521 ;
  assign y24048 = ~n41523 ;
  assign y24049 = n41526 ;
  assign y24050 = 1'b0 ;
  assign y24051 = n41527 ;
  assign y24052 = n41531 ;
  assign y24053 = 1'b0 ;
  assign y24054 = ~1'b0 ;
  assign y24055 = ~1'b0 ;
  assign y24056 = ~1'b0 ;
  assign y24057 = n41534 ;
  assign y24058 = n41535 ;
  assign y24059 = n41536 ;
  assign y24060 = ~n18080 ;
  assign y24061 = n41540 ;
  assign y24062 = n41547 ;
  assign y24063 = n41549 ;
  assign y24064 = ~1'b0 ;
  assign y24065 = ~n41551 ;
  assign y24066 = n41554 ;
  assign y24067 = n41556 ;
  assign y24068 = ~n40495 ;
  assign y24069 = n40442 ;
  assign y24070 = ~n41559 ;
  assign y24071 = ~n41561 ;
  assign y24072 = n41563 ;
  assign y24073 = ~1'b0 ;
  assign y24074 = ~1'b0 ;
  assign y24075 = ~n41565 ;
  assign y24076 = n3930 ;
  assign y24077 = ~1'b0 ;
  assign y24078 = n41566 ;
  assign y24079 = ~1'b0 ;
  assign y24080 = ~n41567 ;
  assign y24081 = ~1'b0 ;
  assign y24082 = ~n41568 ;
  assign y24083 = n41572 ;
  assign y24084 = ~n41575 ;
  assign y24085 = ~1'b0 ;
  assign y24086 = ~1'b0 ;
  assign y24087 = ~n41577 ;
  assign y24088 = ~1'b0 ;
  assign y24089 = ~n41583 ;
  assign y24090 = n41050 ;
  assign y24091 = ~n41585 ;
  assign y24092 = ~1'b0 ;
  assign y24093 = ~n41586 ;
  assign y24094 = ~1'b0 ;
  assign y24095 = ~1'b0 ;
  assign y24096 = ~1'b0 ;
  assign y24097 = n41591 ;
  assign y24098 = n31932 ;
  assign y24099 = ~n41594 ;
  assign y24100 = n4960 ;
  assign y24101 = n41596 ;
  assign y24102 = ~n4718 ;
  assign y24103 = ~n41598 ;
  assign y24104 = ~1'b0 ;
  assign y24105 = ~1'b0 ;
  assign y24106 = ~n41603 ;
  assign y24107 = ~n41604 ;
  assign y24108 = n41607 ;
  assign y24109 = n41610 ;
  assign y24110 = ~n41612 ;
  assign y24111 = ~1'b0 ;
  assign y24112 = ~n41615 ;
  assign y24113 = ~n41623 ;
  assign y24114 = ~1'b0 ;
  assign y24115 = n13042 ;
  assign y24116 = ~n41624 ;
  assign y24117 = ~1'b0 ;
  assign y24118 = ~1'b0 ;
  assign y24119 = ~1'b0 ;
  assign y24120 = ~1'b0 ;
  assign y24121 = n41625 ;
  assign y24122 = ~1'b0 ;
  assign y24123 = ~1'b0 ;
  assign y24124 = n41629 ;
  assign y24125 = n41632 ;
  assign y24126 = ~n41638 ;
  assign y24127 = ~n41640 ;
  assign y24128 = ~1'b0 ;
  assign y24129 = ~n41641 ;
  assign y24130 = ~n41642 ;
  assign y24131 = ~n41643 ;
  assign y24132 = ~n41645 ;
  assign y24133 = ~n41647 ;
  assign y24134 = 1'b0 ;
  assign y24135 = ~1'b0 ;
  assign y24136 = ~n41648 ;
  assign y24137 = ~1'b0 ;
  assign y24138 = ~1'b0 ;
  assign y24139 = n41650 ;
  assign y24140 = ~1'b0 ;
  assign y24141 = ~1'b0 ;
  assign y24142 = ~1'b0 ;
  assign y24143 = ~n1251 ;
  assign y24144 = ~n41654 ;
  assign y24145 = ~n41659 ;
  assign y24146 = ~n41660 ;
  assign y24147 = ~n11891 ;
  assign y24148 = ~n41662 ;
  assign y24149 = ~1'b0 ;
  assign y24150 = n41663 ;
  assign y24151 = ~n41664 ;
  assign y24152 = ~n41666 ;
  assign y24153 = n6185 ;
  assign y24154 = ~n41667 ;
  assign y24155 = ~1'b0 ;
  assign y24156 = ~n41668 ;
  assign y24157 = ~n41669 ;
  assign y24158 = n22256 ;
  assign y24159 = ~n41670 ;
  assign y24160 = ~1'b0 ;
  assign y24161 = n41671 ;
  assign y24162 = ~1'b0 ;
  assign y24163 = ~n34630 ;
  assign y24164 = ~1'b0 ;
  assign y24165 = n41672 ;
  assign y24166 = ~n41674 ;
  assign y24167 = ~1'b0 ;
  assign y24168 = ~1'b0 ;
  assign y24169 = ~n41675 ;
  assign y24170 = ~n41678 ;
  assign y24171 = n41680 ;
  assign y24172 = n41681 ;
  assign y24173 = n41682 ;
  assign y24174 = ~n41688 ;
  assign y24175 = ~n41689 ;
  assign y24176 = n41690 ;
  assign y24177 = ~n41691 ;
  assign y24178 = n41693 ;
  assign y24179 = ~n41695 ;
  assign y24180 = ~1'b0 ;
  assign y24181 = ~n41697 ;
  assign y24182 = ~n41700 ;
  assign y24183 = n41703 ;
  assign y24184 = ~n41705 ;
  assign y24185 = ~n41708 ;
  assign y24186 = n41710 ;
  assign y24187 = n41713 ;
  assign y24188 = n41714 ;
  assign y24189 = n41716 ;
  assign y24190 = ~1'b0 ;
  assign y24191 = ~n41717 ;
  assign y24192 = n25726 ;
  assign y24193 = n41718 ;
  assign y24194 = n41719 ;
  assign y24195 = n19468 ;
  assign y24196 = ~1'b0 ;
  assign y24197 = n41722 ;
  assign y24198 = ~n41724 ;
  assign y24199 = n14593 ;
  assign y24200 = ~1'b0 ;
  assign y24201 = ~n41725 ;
  assign y24202 = ~1'b0 ;
  assign y24203 = ~n41727 ;
  assign y24204 = ~n41728 ;
  assign y24205 = ~1'b0 ;
  assign y24206 = ~1'b0 ;
  assign y24207 = n41729 ;
  assign y24208 = ~1'b0 ;
  assign y24209 = ~1'b0 ;
  assign y24210 = ~1'b0 ;
  assign y24211 = ~1'b0 ;
  assign y24212 = n41731 ;
  assign y24213 = ~n41732 ;
  assign y24214 = n41733 ;
  assign y24215 = ~1'b0 ;
  assign y24216 = ~1'b0 ;
  assign y24217 = ~n41735 ;
  assign y24218 = ~1'b0 ;
  assign y24219 = ~1'b0 ;
  assign y24220 = ~1'b0 ;
  assign y24221 = 1'b0 ;
  assign y24222 = n41738 ;
  assign y24223 = n41740 ;
  assign y24224 = n41741 ;
  assign y24225 = ~n41748 ;
  assign y24226 = ~n41752 ;
  assign y24227 = n41754 ;
  assign y24228 = ~1'b0 ;
  assign y24229 = n41759 ;
  assign y24230 = ~1'b0 ;
  assign y24231 = ~n41760 ;
  assign y24232 = n35704 ;
  assign y24233 = ~1'b0 ;
  assign y24234 = ~n41768 ;
  assign y24235 = ~n41775 ;
  assign y24236 = ~1'b0 ;
  assign y24237 = n41778 ;
  assign y24238 = n41779 ;
  assign y24239 = ~n41781 ;
  assign y24240 = n41786 ;
  assign y24241 = n41787 ;
  assign y24242 = ~1'b0 ;
  assign y24243 = ~1'b0 ;
  assign y24244 = ~n41791 ;
  assign y24245 = ~1'b0 ;
  assign y24246 = ~n41792 ;
  assign y24247 = n41793 ;
  assign y24248 = ~n16032 ;
  assign y24249 = ~1'b0 ;
  assign y24250 = n19759 ;
  assign y24251 = n41794 ;
  assign y24252 = ~1'b0 ;
  assign y24253 = 1'b0 ;
  assign y24254 = n41796 ;
  assign y24255 = ~1'b0 ;
  assign y24256 = ~1'b0 ;
  assign y24257 = n41797 ;
  assign y24258 = ~1'b0 ;
  assign y24259 = ~n41798 ;
  assign y24260 = n28960 ;
  assign y24261 = ~n41800 ;
  assign y24262 = ~n30989 ;
  assign y24263 = n41801 ;
  assign y24264 = n41802 ;
  assign y24265 = ~1'b0 ;
  assign y24266 = n41804 ;
  assign y24267 = ~n41806 ;
  assign y24268 = ~1'b0 ;
  assign y24269 = ~n41809 ;
  assign y24270 = n41810 ;
  assign y24271 = n41812 ;
  assign y24272 = n41814 ;
  assign y24273 = ~n27168 ;
  assign y24274 = n41815 ;
  assign y24275 = n41821 ;
  assign y24276 = n22218 ;
  assign y24277 = ~1'b0 ;
  assign y24278 = ~1'b0 ;
  assign y24279 = ~n41824 ;
  assign y24280 = ~1'b0 ;
  assign y24281 = ~n41828 ;
  assign y24282 = ~1'b0 ;
  assign y24283 = n41831 ;
  assign y24284 = n41833 ;
  assign y24285 = n41836 ;
  assign y24286 = 1'b0 ;
  assign y24287 = ~n41837 ;
  assign y24288 = n41845 ;
  assign y24289 = ~n41852 ;
  assign y24290 = n41853 ;
  assign y24291 = n41858 ;
  assign y24292 = ~n41862 ;
  assign y24293 = ~n41868 ;
  assign y24294 = ~n41869 ;
  assign y24295 = n41870 ;
  assign y24296 = ~n41872 ;
  assign y24297 = ~n41878 ;
  assign y24298 = ~n41880 ;
  assign y24299 = n41881 ;
  assign y24300 = ~1'b0 ;
  assign y24301 = n41883 ;
  assign y24302 = ~1'b0 ;
  assign y24303 = ~n41888 ;
  assign y24304 = ~1'b0 ;
  assign y24305 = ~n41889 ;
  assign y24306 = n41891 ;
  assign y24307 = n41892 ;
  assign y24308 = n41896 ;
  assign y24309 = ~1'b0 ;
  assign y24310 = ~n41900 ;
  assign y24311 = ~n41903 ;
  assign y24312 = 1'b0 ;
  assign y24313 = n41905 ;
  assign y24314 = n41909 ;
  assign y24315 = n41913 ;
  assign y24316 = n41915 ;
  assign y24317 = ~1'b0 ;
  assign y24318 = ~n41920 ;
  assign y24319 = ~n41925 ;
  assign y24320 = n41926 ;
  assign y24321 = n41927 ;
  assign y24322 = ~n41929 ;
  assign y24323 = n41932 ;
  assign y24324 = n41933 ;
  assign y24325 = n41934 ;
  assign y24326 = ~1'b0 ;
  assign y24327 = ~n41935 ;
  assign y24328 = n41939 ;
  assign y24329 = ~n41941 ;
  assign y24330 = ~1'b0 ;
  assign y24331 = ~n41947 ;
  assign y24332 = n41949 ;
  assign y24333 = n41951 ;
  assign y24334 = ~n41952 ;
  assign y24335 = n41954 ;
  assign y24336 = n41955 ;
  assign y24337 = ~1'b0 ;
  assign y24338 = ~1'b0 ;
  assign y24339 = ~1'b0 ;
  assign y24340 = ~1'b0 ;
  assign y24341 = ~1'b0 ;
  assign y24342 = ~1'b0 ;
  assign y24343 = n41958 ;
  assign y24344 = n41959 ;
  assign y24345 = ~n41961 ;
  assign y24346 = ~n41962 ;
  assign y24347 = n41964 ;
  assign y24348 = 1'b0 ;
  assign y24349 = ~n41971 ;
  assign y24350 = ~1'b0 ;
  assign y24351 = ~n41974 ;
  assign y24352 = ~n41976 ;
  assign y24353 = ~n41977 ;
  assign y24354 = n41979 ;
  assign y24355 = n41982 ;
  assign y24356 = ~1'b0 ;
  assign y24357 = ~1'b0 ;
  assign y24358 = ~n41983 ;
  assign y24359 = n41985 ;
  assign y24360 = ~1'b0 ;
  assign y24361 = ~n41986 ;
  assign y24362 = ~1'b0 ;
  assign y24363 = ~1'b0 ;
  assign y24364 = n41989 ;
  assign y24365 = n41995 ;
  assign y24366 = ~n41997 ;
  assign y24367 = n41999 ;
  assign y24368 = ~n42001 ;
  assign y24369 = n42002 ;
  assign y24370 = ~n42006 ;
  assign y24371 = ~1'b0 ;
  assign y24372 = ~n42008 ;
  assign y24373 = ~n42010 ;
  assign y24374 = n42011 ;
  assign y24375 = ~n42015 ;
  assign y24376 = 1'b0 ;
  assign y24377 = ~1'b0 ;
  assign y24378 = n42019 ;
  assign y24379 = n42020 ;
  assign y24380 = ~1'b0 ;
  assign y24381 = ~1'b0 ;
  assign y24382 = ~1'b0 ;
  assign y24383 = n42023 ;
  assign y24384 = ~1'b0 ;
  assign y24385 = ~n42027 ;
  assign y24386 = n42029 ;
  assign y24387 = n42038 ;
  assign y24388 = ~1'b0 ;
  assign y24389 = n34818 ;
  assign y24390 = n42040 ;
  assign y24391 = ~1'b0 ;
  assign y24392 = ~n42041 ;
  assign y24393 = n42046 ;
  assign y24394 = ~1'b0 ;
  assign y24395 = ~n42048 ;
  assign y24396 = ~1'b0 ;
  assign y24397 = ~n2292 ;
  assign y24398 = n42050 ;
  assign y24399 = n42051 ;
  assign y24400 = n42052 ;
  assign y24401 = ~1'b0 ;
  assign y24402 = ~1'b0 ;
  assign y24403 = ~1'b0 ;
  assign y24404 = n38373 ;
  assign y24405 = ~1'b0 ;
  assign y24406 = ~n42059 ;
  assign y24407 = n42062 ;
  assign y24408 = ~1'b0 ;
  assign y24409 = ~1'b0 ;
  assign y24410 = ~1'b0 ;
  assign y24411 = n42065 ;
  assign y24412 = n42067 ;
  assign y24413 = n42071 ;
  assign y24414 = n42074 ;
  assign y24415 = ~n42075 ;
  assign y24416 = n42076 ;
  assign y24417 = ~n42080 ;
  assign y24418 = ~n39356 ;
  assign y24419 = ~n42081 ;
  assign y24420 = n42083 ;
  assign y24421 = ~1'b0 ;
  assign y24422 = ~1'b0 ;
  assign y24423 = ~n42087 ;
  assign y24424 = n42088 ;
  assign y24425 = ~n42091 ;
  assign y24426 = 1'b0 ;
  assign y24427 = ~1'b0 ;
  assign y24428 = n26535 ;
  assign y24429 = ~1'b0 ;
  assign y24430 = ~n42092 ;
  assign y24431 = ~n42093 ;
  assign y24432 = ~n42094 ;
  assign y24433 = ~1'b0 ;
  assign y24434 = ~1'b0 ;
  assign y24435 = ~1'b0 ;
  assign y24436 = 1'b0 ;
  assign y24437 = ~n42098 ;
  assign y24438 = ~n42104 ;
  assign y24439 = ~n42107 ;
  assign y24440 = n42109 ;
  assign y24441 = ~n42113 ;
  assign y24442 = n42114 ;
  assign y24443 = ~1'b0 ;
  assign y24444 = n25069 ;
  assign y24445 = ~1'b0 ;
  assign y24446 = ~1'b0 ;
  assign y24447 = n42115 ;
  assign y24448 = n33582 ;
  assign y24449 = ~n42118 ;
  assign y24450 = ~n42119 ;
  assign y24451 = ~n42120 ;
  assign y24452 = ~n39267 ;
  assign y24453 = ~1'b0 ;
  assign y24454 = n42121 ;
  assign y24455 = ~n42123 ;
  assign y24456 = ~n5041 ;
  assign y24457 = ~1'b0 ;
  assign y24458 = ~1'b0 ;
  assign y24459 = ~n42125 ;
  assign y24460 = n42128 ;
  assign y24461 = ~n42129 ;
  assign y24462 = n42130 ;
  assign y24463 = n42133 ;
  assign y24464 = 1'b0 ;
  assign y24465 = ~n42136 ;
  assign y24466 = ~1'b0 ;
  assign y24467 = ~n42139 ;
  assign y24468 = n42140 ;
  assign y24469 = n42141 ;
  assign y24470 = n18514 ;
  assign y24471 = n42142 ;
  assign y24472 = ~n1736 ;
  assign y24473 = ~n42144 ;
  assign y24474 = ~n42150 ;
  assign y24475 = ~n42152 ;
  assign y24476 = n42155 ;
  assign y24477 = ~n32562 ;
  assign y24478 = ~1'b0 ;
  assign y24479 = ~1'b0 ;
  assign y24480 = ~n42156 ;
  assign y24481 = ~n42157 ;
  assign y24482 = ~n42158 ;
  assign y24483 = ~n42160 ;
  assign y24484 = ~n42164 ;
  assign y24485 = ~1'b0 ;
  assign y24486 = ~n42166 ;
  assign y24487 = ~1'b0 ;
  assign y24488 = ~1'b0 ;
  assign y24489 = ~1'b0 ;
  assign y24490 = ~n42170 ;
  assign y24491 = ~n42174 ;
  assign y24492 = ~n42177 ;
  assign y24493 = n42182 ;
  assign y24494 = 1'b0 ;
  assign y24495 = ~n42186 ;
  assign y24496 = n42187 ;
  assign y24497 = n42189 ;
  assign y24498 = ~1'b0 ;
  assign y24499 = ~1'b0 ;
  assign y24500 = n5692 ;
  assign y24501 = n42190 ;
  assign y24502 = ~n42191 ;
  assign y24503 = n42193 ;
  assign y24504 = ~n42194 ;
  assign y24505 = ~1'b0 ;
  assign y24506 = ~1'b0 ;
  assign y24507 = n42198 ;
  assign y24508 = ~n42199 ;
  assign y24509 = ~n42200 ;
  assign y24510 = ~n36631 ;
  assign y24511 = ~1'b0 ;
  assign y24512 = ~1'b0 ;
  assign y24513 = n42204 ;
  assign y24514 = ~1'b0 ;
  assign y24515 = ~1'b0 ;
  assign y24516 = ~n11402 ;
  assign y24517 = n42208 ;
  assign y24518 = ~n42209 ;
  assign y24519 = ~n42214 ;
  assign y24520 = 1'b0 ;
  assign y24521 = ~n42215 ;
  assign y24522 = ~n42217 ;
  assign y24523 = ~1'b0 ;
  assign y24524 = ~n42218 ;
  assign y24525 = ~1'b0 ;
  assign y24526 = n20945 ;
  assign y24527 = ~n42221 ;
  assign y24528 = ~n42228 ;
  assign y24529 = ~1'b0 ;
  assign y24530 = ~n42230 ;
  assign y24531 = ~n42231 ;
  assign y24532 = ~n9886 ;
  assign y24533 = ~1'b0 ;
  assign y24534 = ~1'b0 ;
  assign y24535 = ~1'b0 ;
  assign y24536 = ~1'b0 ;
  assign y24537 = ~1'b0 ;
  assign y24538 = n8324 ;
  assign y24539 = ~n42234 ;
  assign y24540 = ~n42236 ;
  assign y24541 = n42237 ;
  assign y24542 = n42239 ;
  assign y24543 = ~1'b0 ;
  assign y24544 = ~n42238 ;
  assign y24545 = ~n42240 ;
  assign y24546 = ~1'b0 ;
  assign y24547 = n42245 ;
  assign y24548 = ~n42249 ;
  assign y24549 = ~n42251 ;
  assign y24550 = ~n12356 ;
  assign y24551 = n42259 ;
  assign y24552 = ~n42261 ;
  assign y24553 = ~n42262 ;
  assign y24554 = ~n42263 ;
  assign y24555 = ~n42268 ;
  assign y24556 = n42270 ;
  assign y24557 = ~n42271 ;
  assign y24558 = ~n42273 ;
  assign y24559 = n34131 ;
  assign y24560 = ~n42275 ;
  assign y24561 = ~1'b0 ;
  assign y24562 = n42283 ;
  assign y24563 = ~n42285 ;
  assign y24564 = ~n42288 ;
  assign y24565 = n42289 ;
  assign y24566 = ~1'b0 ;
  assign y24567 = n42290 ;
  assign y24568 = ~1'b0 ;
  assign y24569 = ~n42293 ;
  assign y24570 = ~n42294 ;
  assign y24571 = n42301 ;
  assign y24572 = ~1'b0 ;
  assign y24573 = ~n42303 ;
  assign y24574 = ~1'b0 ;
  assign y24575 = 1'b0 ;
  assign y24576 = n42305 ;
  assign y24577 = ~1'b0 ;
  assign y24578 = n42306 ;
  assign y24579 = ~1'b0 ;
  assign y24580 = ~1'b0 ;
  assign y24581 = n42308 ;
  assign y24582 = ~1'b0 ;
  assign y24583 = n8884 ;
  assign y24584 = n42311 ;
  assign y24585 = ~n42314 ;
  assign y24586 = ~1'b0 ;
  assign y24587 = ~n42317 ;
  assign y24588 = n42320 ;
  assign y24589 = ~n42321 ;
  assign y24590 = ~1'b0 ;
  assign y24591 = ~n29482 ;
  assign y24592 = ~1'b0 ;
  assign y24593 = ~n42323 ;
  assign y24594 = n42325 ;
  assign y24595 = ~1'b0 ;
  assign y24596 = ~n42330 ;
  assign y24597 = ~1'b0 ;
  assign y24598 = ~n42331 ;
  assign y24599 = n42334 ;
  assign y24600 = n42337 ;
  assign y24601 = ~n42341 ;
  assign y24602 = n42342 ;
  assign y24603 = ~1'b0 ;
  assign y24604 = ~n42343 ;
  assign y24605 = n42345 ;
  assign y24606 = ~1'b0 ;
  assign y24607 = ~n42347 ;
  assign y24608 = ~1'b0 ;
  assign y24609 = ~1'b0 ;
  assign y24610 = ~n42348 ;
  assign y24611 = ~n42353 ;
  assign y24612 = ~n2962 ;
  assign y24613 = ~n42354 ;
  assign y24614 = ~1'b0 ;
  assign y24615 = ~n42358 ;
  assign y24616 = ~1'b0 ;
  assign y24617 = ~n42360 ;
  assign y24618 = ~1'b0 ;
  assign y24619 = ~1'b0 ;
  assign y24620 = n42361 ;
  assign y24621 = ~1'b0 ;
  assign y24622 = n42363 ;
  assign y24623 = n42364 ;
  assign y24624 = ~1'b0 ;
  assign y24625 = ~1'b0 ;
  assign y24626 = ~1'b0 ;
  assign y24627 = ~n2424 ;
  assign y24628 = ~1'b0 ;
  assign y24629 = ~n42366 ;
  assign y24630 = n42367 ;
  assign y24631 = ~n42370 ;
  assign y24632 = ~1'b0 ;
  assign y24633 = n42377 ;
  assign y24634 = ~1'b0 ;
  assign y24635 = ~1'b0 ;
  assign y24636 = n42380 ;
  assign y24637 = n42381 ;
  assign y24638 = ~1'b0 ;
  assign y24639 = n42382 ;
  assign y24640 = n18544 ;
  assign y24641 = ~n42387 ;
  assign y24642 = ~n42390 ;
  assign y24643 = ~1'b0 ;
  assign y24644 = ~n42393 ;
  assign y24645 = ~1'b0 ;
  assign y24646 = n42397 ;
  assign y24647 = ~1'b0 ;
  assign y24648 = ~n42402 ;
  assign y24649 = n42403 ;
  assign y24650 = n42404 ;
  assign y24651 = ~1'b0 ;
  assign y24652 = n42405 ;
  assign y24653 = ~n42408 ;
  assign y24654 = n42409 ;
  assign y24655 = ~1'b0 ;
  assign y24656 = 1'b0 ;
  assign y24657 = ~1'b0 ;
  assign y24658 = n42410 ;
  assign y24659 = n42412 ;
  assign y24660 = ~1'b0 ;
  assign y24661 = ~n33429 ;
  assign y24662 = ~n42415 ;
  assign y24663 = n42420 ;
  assign y24664 = ~n42422 ;
  assign y24665 = ~n42426 ;
  assign y24666 = n42427 ;
  assign y24667 = ~n42428 ;
  assign y24668 = n42430 ;
  assign y24669 = ~n42431 ;
  assign y24670 = ~1'b0 ;
  assign y24671 = n42432 ;
  assign y24672 = ~n28020 ;
  assign y24673 = 1'b0 ;
  assign y24674 = n42434 ;
  assign y24675 = ~1'b0 ;
  assign y24676 = ~1'b0 ;
  assign y24677 = ~n42435 ;
  assign y24678 = n42437 ;
  assign y24679 = n42440 ;
  assign y24680 = n42441 ;
  assign y24681 = ~1'b0 ;
  assign y24682 = ~n42442 ;
  assign y24683 = ~n42445 ;
  assign y24684 = ~n42446 ;
  assign y24685 = ~n42450 ;
  assign y24686 = ~n42451 ;
  assign y24687 = n42452 ;
  assign y24688 = n42453 ;
  assign y24689 = ~n42457 ;
  assign y24690 = ~1'b0 ;
  assign y24691 = n42458 ;
  assign y24692 = ~n42461 ;
  assign y24693 = ~n42463 ;
  assign y24694 = ~1'b0 ;
  assign y24695 = n42466 ;
  assign y24696 = ~n42467 ;
  assign y24697 = n2356 ;
  assign y24698 = ~1'b0 ;
  assign y24699 = ~1'b0 ;
  assign y24700 = ~n42469 ;
  assign y24701 = ~n16120 ;
  assign y24702 = ~1'b0 ;
  assign y24703 = n42472 ;
  assign y24704 = n42473 ;
  assign y24705 = n42476 ;
  assign y24706 = ~n42482 ;
  assign y24707 = ~n27498 ;
  assign y24708 = ~n42489 ;
  assign y24709 = ~n42491 ;
  assign y24710 = ~n42492 ;
  assign y24711 = ~n42496 ;
  assign y24712 = n20695 ;
  assign y24713 = n42502 ;
  assign y24714 = n42504 ;
  assign y24715 = ~n42505 ;
  assign y24716 = ~1'b0 ;
  assign y24717 = ~1'b0 ;
  assign y24718 = ~n42506 ;
  assign y24719 = ~1'b0 ;
  assign y24720 = ~1'b0 ;
  assign y24721 = ~n42510 ;
  assign y24722 = ~1'b0 ;
  assign y24723 = ~1'b0 ;
  assign y24724 = ~1'b0 ;
  assign y24725 = ~n2971 ;
  assign y24726 = ~n42514 ;
  assign y24727 = ~n42515 ;
  assign y24728 = 1'b0 ;
  assign y24729 = ~n42516 ;
  assign y24730 = ~1'b0 ;
  assign y24731 = ~1'b0 ;
  assign y24732 = n42518 ;
  assign y24733 = ~n34302 ;
  assign y24734 = ~1'b0 ;
  assign y24735 = n42519 ;
  assign y24736 = n7734 ;
  assign y24737 = n42520 ;
  assign y24738 = 1'b0 ;
  assign y24739 = ~n42524 ;
  assign y24740 = n8963 ;
  assign y24741 = n42530 ;
  assign y24742 = ~n42533 ;
  assign y24743 = ~n42534 ;
  assign y24744 = ~1'b0 ;
  assign y24745 = ~1'b0 ;
  assign y24746 = n42535 ;
  assign y24747 = n42538 ;
  assign y24748 = ~n42543 ;
  assign y24749 = ~n42547 ;
  assign y24750 = ~1'b0 ;
  assign y24751 = ~n8639 ;
  assign y24752 = n42548 ;
  assign y24753 = ~1'b0 ;
  assign y24754 = ~n42552 ;
  assign y24755 = 1'b0 ;
  assign y24756 = ~1'b0 ;
  assign y24757 = n42556 ;
  assign y24758 = ~n42559 ;
  assign y24759 = ~1'b0 ;
  assign y24760 = ~1'b0 ;
  assign y24761 = ~n42561 ;
  assign y24762 = ~n42562 ;
  assign y24763 = ~n42563 ;
  assign y24764 = ~n42564 ;
  assign y24765 = ~n42568 ;
  assign y24766 = ~n42569 ;
  assign y24767 = ~n34249 ;
  assign y24768 = ~n27349 ;
  assign y24769 = ~1'b0 ;
  assign y24770 = ~1'b0 ;
  assign y24771 = ~1'b0 ;
  assign y24772 = ~n42570 ;
  assign y24773 = ~n42571 ;
  assign y24774 = n42579 ;
  assign y24775 = ~1'b0 ;
  assign y24776 = n42580 ;
  assign y24777 = ~1'b0 ;
  assign y24778 = ~1'b0 ;
  assign y24779 = ~n35581 ;
  assign y24780 = n42581 ;
  assign y24781 = n42582 ;
  assign y24782 = ~n42583 ;
  assign y24783 = ~1'b0 ;
  assign y24784 = ~1'b0 ;
  assign y24785 = ~1'b0 ;
  assign y24786 = ~n42587 ;
  assign y24787 = ~n42591 ;
  assign y24788 = n42593 ;
  assign y24789 = ~n42595 ;
  assign y24790 = ~n42600 ;
  assign y24791 = ~1'b0 ;
  assign y24792 = ~1'b0 ;
  assign y24793 = ~n42602 ;
  assign y24794 = ~n42604 ;
  assign y24795 = n42605 ;
  assign y24796 = ~1'b0 ;
  assign y24797 = n42606 ;
  assign y24798 = n42608 ;
  assign y24799 = ~1'b0 ;
  assign y24800 = 1'b0 ;
  assign y24801 = ~1'b0 ;
  assign y24802 = ~n42612 ;
  assign y24803 = ~1'b0 ;
  assign y24804 = ~n3124 ;
  assign y24805 = ~1'b0 ;
  assign y24806 = ~1'b0 ;
  assign y24807 = ~n42619 ;
  assign y24808 = ~n42621 ;
  assign y24809 = n42622 ;
  assign y24810 = ~n42625 ;
  assign y24811 = ~n42627 ;
  assign y24812 = n42632 ;
  assign y24813 = ~n42634 ;
  assign y24814 = 1'b0 ;
  assign y24815 = n42635 ;
  assign y24816 = ~n42636 ;
  assign y24817 = n42637 ;
  assign y24818 = ~n11655 ;
  assign y24819 = ~1'b0 ;
  assign y24820 = ~1'b0 ;
  assign y24821 = n42638 ;
  assign y24822 = ~n42639 ;
  assign y24823 = ~n21297 ;
  assign y24824 = n42642 ;
  assign y24825 = ~n13011 ;
  assign y24826 = ~n42643 ;
  assign y24827 = ~n42646 ;
  assign y24828 = n42650 ;
  assign y24829 = ~n42651 ;
  assign y24830 = n42654 ;
  assign y24831 = ~1'b0 ;
  assign y24832 = ~n42655 ;
  assign y24833 = ~1'b0 ;
  assign y24834 = ~1'b0 ;
  assign y24835 = n42658 ;
  assign y24836 = ~n42660 ;
  assign y24837 = ~n42661 ;
  assign y24838 = ~n16185 ;
  assign y24839 = n42667 ;
  assign y24840 = ~n42669 ;
  assign y24841 = n5145 ;
  assign y24842 = n42670 ;
  assign y24843 = n42673 ;
  assign y24844 = ~1'b0 ;
  assign y24845 = n42674 ;
  assign y24846 = ~n42677 ;
  assign y24847 = 1'b0 ;
  assign y24848 = ~1'b0 ;
  assign y24849 = n42678 ;
  assign y24850 = n42679 ;
  assign y24851 = n42680 ;
  assign y24852 = n42681 ;
  assign y24853 = ~n42683 ;
  assign y24854 = ~n21438 ;
  assign y24855 = ~1'b0 ;
  assign y24856 = ~1'b0 ;
  assign y24857 = n42685 ;
  assign y24858 = n42687 ;
  assign y24859 = ~n42695 ;
  assign y24860 = ~1'b0 ;
  assign y24861 = ~1'b0 ;
  assign y24862 = ~1'b0 ;
  assign y24863 = ~n42697 ;
  assign y24864 = ~1'b0 ;
  assign y24865 = n42701 ;
  assign y24866 = ~1'b0 ;
  assign y24867 = n42702 ;
  assign y24868 = n42707 ;
  assign y24869 = ~n42710 ;
  assign y24870 = n42711 ;
  assign y24871 = ~n42712 ;
  assign y24872 = ~1'b0 ;
  assign y24873 = ~n42713 ;
  assign y24874 = ~n42716 ;
  assign y24875 = ~n2981 ;
  assign y24876 = n42717 ;
  assign y24877 = ~n42719 ;
  assign y24878 = ~n11485 ;
  assign y24879 = ~n42720 ;
  assign y24880 = ~n5222 ;
  assign y24881 = n42721 ;
  assign y24882 = 1'b0 ;
  assign y24883 = n42722 ;
  assign y24884 = n42726 ;
  assign y24885 = ~n42728 ;
  assign y24886 = ~1'b0 ;
  assign y24887 = n42732 ;
  assign y24888 = ~1'b0 ;
  assign y24889 = ~n42733 ;
  assign y24890 = ~n42734 ;
  assign y24891 = ~1'b0 ;
  assign y24892 = ~1'b0 ;
  assign y24893 = n42736 ;
  assign y24894 = ~1'b0 ;
  assign y24895 = ~n42739 ;
  assign y24896 = 1'b0 ;
  assign y24897 = ~n42740 ;
  assign y24898 = n42741 ;
  assign y24899 = ~n42742 ;
  assign y24900 = ~n42747 ;
  assign y24901 = ~n831 ;
  assign y24902 = n42748 ;
  assign y24903 = ~1'b0 ;
  assign y24904 = ~n42750 ;
  assign y24905 = n42751 ;
  assign y24906 = ~1'b0 ;
  assign y24907 = ~n16411 ;
  assign y24908 = n42752 ;
  assign y24909 = ~n42757 ;
  assign y24910 = n42759 ;
  assign y24911 = n34111 ;
  assign y24912 = ~n3314 ;
  assign y24913 = n42761 ;
  assign y24914 = n42765 ;
  assign y24915 = ~1'b0 ;
  assign y24916 = n27773 ;
  assign y24917 = ~n42766 ;
  assign y24918 = n42770 ;
  assign y24919 = n42771 ;
  assign y24920 = ~1'b0 ;
  assign y24921 = ~1'b0 ;
  assign y24922 = ~1'b0 ;
  assign y24923 = ~n33973 ;
  assign y24924 = ~n7994 ;
  assign y24925 = ~n42772 ;
  assign y24926 = n42774 ;
  assign y24927 = n42775 ;
  assign y24928 = ~n42776 ;
  assign y24929 = n42777 ;
  assign y24930 = ~n42779 ;
  assign y24931 = n42781 ;
  assign y24932 = n16021 ;
  assign y24933 = n42782 ;
  assign y24934 = ~n42783 ;
  assign y24935 = n42785 ;
  assign y24936 = n42786 ;
  assign y24937 = ~n42789 ;
  assign y24938 = n42792 ;
  assign y24939 = ~1'b0 ;
  assign y24940 = ~n42796 ;
  assign y24941 = ~1'b0 ;
  assign y24942 = 1'b0 ;
  assign y24943 = ~n42803 ;
  assign y24944 = n10790 ;
  assign y24945 = ~n42809 ;
  assign y24946 = ~1'b0 ;
  assign y24947 = n42810 ;
  assign y24948 = ~1'b0 ;
  assign y24949 = n42811 ;
  assign y24950 = ~1'b0 ;
  assign y24951 = ~n42814 ;
  assign y24952 = n42816 ;
  assign y24953 = ~n15028 ;
  assign y24954 = ~n42817 ;
  assign y24955 = n42823 ;
  assign y24956 = n42825 ;
  assign y24957 = n42826 ;
  assign y24958 = ~n42828 ;
  assign y24959 = ~1'b0 ;
  assign y24960 = ~n42830 ;
  assign y24961 = ~1'b0 ;
  assign y24962 = n42834 ;
  assign y24963 = ~1'b0 ;
  assign y24964 = ~n42836 ;
  assign y24965 = ~n42842 ;
  assign y24966 = ~n42844 ;
  assign y24967 = ~1'b0 ;
  assign y24968 = n42846 ;
  assign y24969 = ~1'b0 ;
  assign y24970 = ~n42878 ;
  assign y24971 = n42879 ;
  assign y24972 = ~1'b0 ;
  assign y24973 = n42881 ;
  assign y24974 = ~1'b0 ;
  assign y24975 = n42884 ;
  assign y24976 = ~1'b0 ;
  assign y24977 = ~n42886 ;
  assign y24978 = ~1'b0 ;
  assign y24979 = n42887 ;
  assign y24980 = n42888 ;
  assign y24981 = n42890 ;
  assign y24982 = ~1'b0 ;
  assign y24983 = ~n42892 ;
  assign y24984 = n16179 ;
  assign y24985 = ~1'b0 ;
  assign y24986 = ~1'b0 ;
  assign y24987 = ~1'b0 ;
  assign y24988 = n42893 ;
  assign y24989 = ~n42896 ;
  assign y24990 = n42900 ;
  assign y24991 = n31903 ;
  assign y24992 = ~n42902 ;
  assign y24993 = 1'b0 ;
  assign y24994 = ~1'b0 ;
  assign y24995 = ~1'b0 ;
  assign y24996 = n42903 ;
  assign y24997 = n42911 ;
  assign y24998 = ~n42912 ;
  assign y24999 = ~n42913 ;
  assign y25000 = ~n17412 ;
  assign y25001 = n42914 ;
  assign y25002 = ~n22073 ;
  assign y25003 = ~1'b0 ;
  assign y25004 = n42915 ;
  assign y25005 = ~n42917 ;
  assign y25006 = ~1'b0 ;
  assign y25007 = ~n42919 ;
  assign y25008 = n42920 ;
  assign y25009 = ~1'b0 ;
  assign y25010 = ~n42924 ;
  assign y25011 = ~n42929 ;
  assign y25012 = 1'b0 ;
  assign y25013 = ~n42931 ;
  assign y25014 = n42933 ;
  assign y25015 = ~1'b0 ;
  assign y25016 = ~1'b0 ;
  assign y25017 = ~1'b0 ;
  assign y25018 = n42935 ;
  assign y25019 = ~1'b0 ;
  assign y25020 = n42937 ;
  assign y25021 = ~1'b0 ;
  assign y25022 = ~n42941 ;
  assign y25023 = ~1'b0 ;
  assign y25024 = n42944 ;
  assign y25025 = ~n42946 ;
  assign y25026 = n42948 ;
  assign y25027 = n42949 ;
  assign y25028 = ~n42957 ;
  assign y25029 = n42962 ;
  assign y25030 = 1'b0 ;
  assign y25031 = n42963 ;
  assign y25032 = ~n42966 ;
  assign y25033 = ~1'b0 ;
  assign y25034 = n42967 ;
  assign y25035 = ~n42972 ;
  assign y25036 = ~1'b0 ;
  assign y25037 = ~n42973 ;
  assign y25038 = ~n42977 ;
  assign y25039 = ~n42978 ;
  assign y25040 = ~n42983 ;
  assign y25041 = ~1'b0 ;
  assign y25042 = ~1'b0 ;
  assign y25043 = n42984 ;
  assign y25044 = ~1'b0 ;
  assign y25045 = ~1'b0 ;
  assign y25046 = ~n15147 ;
  assign y25047 = ~1'b0 ;
  assign y25048 = ~1'b0 ;
  assign y25049 = ~n42985 ;
  assign y25050 = ~n42987 ;
  assign y25051 = ~n42988 ;
  assign y25052 = ~n42990 ;
  assign y25053 = ~1'b0 ;
  assign y25054 = n42991 ;
  assign y25055 = ~n42992 ;
  assign y25056 = n42994 ;
  assign y25057 = n42997 ;
  assign y25058 = ~n43004 ;
  assign y25059 = n43007 ;
  assign y25060 = ~1'b0 ;
  assign y25061 = n43008 ;
  assign y25062 = n24810 ;
  assign y25063 = ~n43010 ;
  assign y25064 = ~1'b0 ;
  assign y25065 = ~n43011 ;
  assign y25066 = ~1'b0 ;
  assign y25067 = ~n43012 ;
  assign y25068 = ~n43014 ;
  assign y25069 = ~n43015 ;
  assign y25070 = n43016 ;
  assign y25071 = ~1'b0 ;
  assign y25072 = n43017 ;
  assign y25073 = ~n43021 ;
  assign y25074 = ~n43022 ;
  assign y25075 = ~1'b0 ;
  assign y25076 = ~n43025 ;
  assign y25077 = ~1'b0 ;
  assign y25078 = ~1'b0 ;
  assign y25079 = ~1'b0 ;
  assign y25080 = ~n43027 ;
  assign y25081 = n43029 ;
  assign y25082 = n43030 ;
  assign y25083 = n43033 ;
  assign y25084 = n43034 ;
  assign y25085 = ~1'b0 ;
  assign y25086 = ~n43035 ;
  assign y25087 = 1'b0 ;
  assign y25088 = ~1'b0 ;
  assign y25089 = n43038 ;
  assign y25090 = ~1'b0 ;
  assign y25091 = ~1'b0 ;
  assign y25092 = ~1'b0 ;
  assign y25093 = ~n43040 ;
  assign y25094 = n43043 ;
  assign y25095 = ~1'b0 ;
  assign y25096 = ~1'b0 ;
  assign y25097 = n43046 ;
  assign y25098 = n43047 ;
  assign y25099 = ~1'b0 ;
  assign y25100 = ~1'b0 ;
  assign y25101 = ~n43048 ;
  assign y25102 = ~n43050 ;
  assign y25103 = n43052 ;
  assign y25104 = ~n27680 ;
  assign y25105 = n43055 ;
  assign y25106 = ~n43057 ;
  assign y25107 = ~1'b0 ;
  assign y25108 = n43067 ;
  assign y25109 = ~1'b0 ;
  assign y25110 = ~n43069 ;
  assign y25111 = ~n11500 ;
  assign y25112 = n43070 ;
  assign y25113 = ~1'b0 ;
  assign y25114 = ~1'b0 ;
  assign y25115 = ~n43071 ;
  assign y25116 = n43073 ;
  assign y25117 = ~n43077 ;
  assign y25118 = ~n37386 ;
  assign y25119 = ~n43079 ;
  assign y25120 = n43081 ;
  assign y25121 = n43082 ;
  assign y25122 = ~n43088 ;
  assign y25123 = n43091 ;
  assign y25124 = n43092 ;
  assign y25125 = n43094 ;
  assign y25126 = ~1'b0 ;
  assign y25127 = ~n43095 ;
  assign y25128 = ~1'b0 ;
  assign y25129 = 1'b0 ;
  assign y25130 = ~n43103 ;
  assign y25131 = ~n43104 ;
  assign y25132 = ~n43107 ;
  assign y25133 = ~1'b0 ;
  assign y25134 = n43108 ;
  assign y25135 = ~1'b0 ;
  assign y25136 = ~1'b0 ;
  assign y25137 = ~n43117 ;
  assign y25138 = ~1'b0 ;
  assign y25139 = ~n43122 ;
  assign y25140 = ~n43125 ;
  assign y25141 = ~1'b0 ;
  assign y25142 = ~n43145 ;
  assign y25143 = ~n43148 ;
  assign y25144 = ~n43150 ;
  assign y25145 = ~1'b0 ;
  assign y25146 = ~n43152 ;
  assign y25147 = n8802 ;
  assign y25148 = ~n43156 ;
  assign y25149 = n43158 ;
  assign y25150 = ~1'b0 ;
  assign y25151 = ~n43161 ;
  assign y25152 = n43164 ;
  assign y25153 = ~n43167 ;
  assign y25154 = n43169 ;
  assign y25155 = n43170 ;
  assign y25156 = ~n43173 ;
  assign y25157 = n43176 ;
  assign y25158 = n4814 ;
  assign y25159 = n43180 ;
  assign y25160 = ~n43181 ;
  assign y25161 = ~n43183 ;
  assign y25162 = ~n6156 ;
  assign y25163 = ~1'b0 ;
  assign y25164 = ~n40630 ;
  assign y25165 = n43184 ;
  assign y25166 = ~1'b0 ;
  assign y25167 = ~n43185 ;
  assign y25168 = n28705 ;
  assign y25169 = ~1'b0 ;
  assign y25170 = ~n43186 ;
  assign y25171 = n43188 ;
  assign y25172 = ~n43189 ;
  assign y25173 = ~n43193 ;
  assign y25174 = ~1'b0 ;
  assign y25175 = ~n43194 ;
  assign y25176 = ~n43195 ;
  assign y25177 = n43203 ;
  assign y25178 = n43206 ;
  assign y25179 = ~1'b0 ;
  assign y25180 = ~n43207 ;
  assign y25181 = ~n43211 ;
  assign y25182 = ~n43214 ;
  assign y25183 = n43216 ;
  assign y25184 = ~1'b0 ;
  assign y25185 = 1'b0 ;
  assign y25186 = ~n41720 ;
  assign y25187 = n43217 ;
  assign y25188 = ~n43218 ;
  assign y25189 = ~n43219 ;
  assign y25190 = ~n43221 ;
  assign y25191 = ~n3790 ;
  assign y25192 = n43222 ;
  assign y25193 = n43223 ;
  assign y25194 = ~1'b0 ;
  assign y25195 = ~n43225 ;
  assign y25196 = ~n43226 ;
  assign y25197 = ~n43227 ;
  assign y25198 = ~n43228 ;
  assign y25199 = ~n43230 ;
  assign y25200 = n43231 ;
  assign y25201 = n43235 ;
  assign y25202 = ~n43236 ;
  assign y25203 = ~n43237 ;
  assign y25204 = 1'b0 ;
  assign y25205 = ~1'b0 ;
  assign y25206 = ~n11336 ;
  assign y25207 = n43239 ;
  assign y25208 = n43241 ;
  assign y25209 = n43242 ;
  assign y25210 = ~1'b0 ;
  assign y25211 = n43243 ;
  assign y25212 = ~1'b0 ;
  assign y25213 = n43244 ;
  assign y25214 = n43247 ;
  assign y25215 = n43248 ;
  assign y25216 = 1'b0 ;
  assign y25217 = ~1'b0 ;
  assign y25218 = n43249 ;
  assign y25219 = n43254 ;
  assign y25220 = ~n43255 ;
  assign y25221 = ~n43257 ;
  assign y25222 = ~n43259 ;
  assign y25223 = n43260 ;
  assign y25224 = ~1'b0 ;
  assign y25225 = 1'b0 ;
  assign y25226 = ~1'b0 ;
  assign y25227 = ~1'b0 ;
  assign y25228 = ~1'b0 ;
  assign y25229 = n43262 ;
  assign y25230 = n43264 ;
  assign y25231 = ~1'b0 ;
  assign y25232 = n43267 ;
  assign y25233 = ~n43271 ;
  assign y25234 = n43275 ;
  assign y25235 = ~1'b0 ;
  assign y25236 = ~1'b0 ;
  assign y25237 = ~1'b0 ;
  assign y25238 = ~1'b0 ;
  assign y25239 = n43276 ;
  assign y25240 = ~1'b0 ;
  assign y25241 = n43277 ;
  assign y25242 = ~1'b0 ;
  assign y25243 = n43279 ;
  assign y25244 = ~n43280 ;
  assign y25245 = n43281 ;
  assign y25246 = n43283 ;
  assign y25247 = ~1'b0 ;
  assign y25248 = n43286 ;
  assign y25249 = ~n43287 ;
  assign y25250 = ~1'b0 ;
  assign y25251 = ~n42523 ;
  assign y25252 = ~n1693 ;
  assign y25253 = n43297 ;
  assign y25254 = n43299 ;
  assign y25255 = n43300 ;
  assign y25256 = ~1'b0 ;
  assign y25257 = ~n43301 ;
  assign y25258 = ~1'b0 ;
  assign y25259 = n43303 ;
  assign y25260 = n43305 ;
  assign y25261 = ~1'b0 ;
  assign y25262 = ~1'b0 ;
  assign y25263 = n43306 ;
  assign y25264 = ~1'b0 ;
  assign y25265 = ~1'b0 ;
  assign y25266 = ~n43310 ;
  assign y25267 = n43315 ;
  assign y25268 = n43317 ;
  assign y25269 = ~1'b0 ;
  assign y25270 = ~n43319 ;
  assign y25271 = ~n28140 ;
  assign y25272 = n43320 ;
  assign y25273 = ~n43323 ;
  assign y25274 = n43324 ;
  assign y25275 = ~n43327 ;
  assign y25276 = ~1'b0 ;
  assign y25277 = ~1'b0 ;
  assign y25278 = n43330 ;
  assign y25279 = ~n33299 ;
  assign y25280 = ~1'b0 ;
  assign y25281 = n43332 ;
  assign y25282 = 1'b0 ;
  assign y25283 = n43333 ;
  assign y25284 = n43334 ;
  assign y25285 = n32542 ;
  assign y25286 = ~n43336 ;
  assign y25287 = ~n43338 ;
  assign y25288 = n43340 ;
  assign y25289 = ~1'b0 ;
  assign y25290 = ~n43342 ;
  assign y25291 = n43344 ;
  assign y25292 = ~1'b0 ;
  assign y25293 = ~1'b0 ;
  assign y25294 = ~n24324 ;
  assign y25295 = ~1'b0 ;
  assign y25296 = ~1'b0 ;
  assign y25297 = ~n43345 ;
  assign y25298 = n43346 ;
  assign y25299 = 1'b0 ;
  assign y25300 = n43348 ;
  assign y25301 = 1'b0 ;
  assign y25302 = ~1'b0 ;
  assign y25303 = ~n2087 ;
  assign y25304 = ~1'b0 ;
  assign y25305 = n43349 ;
  assign y25306 = ~n43351 ;
  assign y25307 = ~n43354 ;
  assign y25308 = ~n43355 ;
  assign y25309 = ~1'b0 ;
  assign y25310 = ~n43356 ;
  assign y25311 = ~1'b0 ;
  assign y25312 = n43357 ;
  assign y25313 = ~n43359 ;
  assign y25314 = n43361 ;
  assign y25315 = ~1'b0 ;
  assign y25316 = ~n43362 ;
  assign y25317 = n43365 ;
  assign y25318 = ~1'b0 ;
  assign y25319 = n43368 ;
  assign y25320 = ~n43370 ;
  assign y25321 = ~1'b0 ;
  assign y25322 = ~n43371 ;
  assign y25323 = ~1'b0 ;
  assign y25324 = n43372 ;
  assign y25325 = ~1'b0 ;
  assign y25326 = n43373 ;
  assign y25327 = ~n43374 ;
  assign y25328 = ~1'b0 ;
  assign y25329 = ~n43375 ;
  assign y25330 = ~n43376 ;
  assign y25331 = ~n43378 ;
  assign y25332 = n43383 ;
  assign y25333 = ~n43385 ;
  assign y25334 = ~n43389 ;
  assign y25335 = n43390 ;
  assign y25336 = ~1'b0 ;
  assign y25337 = n43391 ;
  assign y25338 = ~n43392 ;
  assign y25339 = ~1'b0 ;
  assign y25340 = n43393 ;
  assign y25341 = n43396 ;
  assign y25342 = ~n43399 ;
  assign y25343 = ~n43401 ;
  assign y25344 = n43403 ;
  assign y25345 = n43404 ;
  assign y25346 = ~n43405 ;
  assign y25347 = n43407 ;
  assign y25348 = n43410 ;
  assign y25349 = ~n43412 ;
  assign y25350 = ~n43413 ;
  assign y25351 = ~n43414 ;
  assign y25352 = ~1'b0 ;
  assign y25353 = ~1'b0 ;
  assign y25354 = n43415 ;
  assign y25355 = ~1'b0 ;
  assign y25356 = ~1'b0 ;
  assign y25357 = n43416 ;
  assign y25358 = ~n43417 ;
  assign y25359 = ~n22596 ;
  assign y25360 = ~n35312 ;
  assign y25361 = n43418 ;
  assign y25362 = ~1'b0 ;
  assign y25363 = ~1'b0 ;
  assign y25364 = ~1'b0 ;
  assign y25365 = n43419 ;
  assign y25366 = ~1'b0 ;
  assign y25367 = n43420 ;
  assign y25368 = ~1'b0 ;
  assign y25369 = ~1'b0 ;
  assign y25370 = ~1'b0 ;
  assign y25371 = ~n43421 ;
  assign y25372 = ~n43425 ;
  assign y25373 = n43426 ;
  assign y25374 = ~n43427 ;
  assign y25375 = n43429 ;
  assign y25376 = n43433 ;
  assign y25377 = ~n43434 ;
  assign y25378 = ~1'b0 ;
  assign y25379 = n43436 ;
  assign y25380 = n13557 ;
  assign y25381 = ~n14867 ;
  assign y25382 = n43437 ;
  assign y25383 = n13971 ;
  assign y25384 = n43438 ;
  assign y25385 = n18861 ;
  assign y25386 = ~n43440 ;
  assign y25387 = ~n43456 ;
  assign y25388 = n43461 ;
  assign y25389 = n43464 ;
  assign y25390 = ~1'b0 ;
  assign y25391 = ~n43465 ;
  assign y25392 = n43467 ;
  assign y25393 = n39045 ;
  assign y25394 = n43470 ;
  assign y25395 = ~n43472 ;
  assign y25396 = n43476 ;
  assign y25397 = ~n43477 ;
  assign y25398 = ~n43485 ;
  assign y25399 = n43489 ;
  assign y25400 = ~n43490 ;
  assign y25401 = ~1'b0 ;
  assign y25402 = ~n43491 ;
  assign y25403 = ~n43493 ;
  assign y25404 = ~1'b0 ;
  assign y25405 = n7739 ;
  assign y25406 = ~1'b0 ;
  assign y25407 = ~1'b0 ;
  assign y25408 = ~n4546 ;
  assign y25409 = n43496 ;
  assign y25410 = ~1'b0 ;
  assign y25411 = n43498 ;
  assign y25412 = ~n43500 ;
  assign y25413 = ~1'b0 ;
  assign y25414 = ~n43501 ;
  assign y25415 = ~n43504 ;
  assign y25416 = ~n43506 ;
  assign y25417 = ~n18270 ;
  assign y25418 = 1'b0 ;
  assign y25419 = n43507 ;
  assign y25420 = ~n43510 ;
  assign y25421 = ~n3586 ;
  assign y25422 = ~1'b0 ;
  assign y25423 = ~1'b0 ;
  assign y25424 = ~n43511 ;
  assign y25425 = ~n43513 ;
  assign y25426 = ~n43521 ;
  assign y25427 = ~1'b0 ;
  assign y25428 = ~n43522 ;
  assign y25429 = n43523 ;
  assign y25430 = ~n43524 ;
  assign y25431 = ~1'b0 ;
  assign y25432 = 1'b0 ;
  assign y25433 = ~1'b0 ;
  assign y25434 = ~n43525 ;
  assign y25435 = n43527 ;
  assign y25436 = n43529 ;
  assign y25437 = n20798 ;
  assign y25438 = n22794 ;
  assign y25439 = 1'b0 ;
  assign y25440 = n43531 ;
  assign y25441 = n43533 ;
  assign y25442 = ~1'b0 ;
  assign y25443 = ~1'b0 ;
  assign y25444 = ~1'b0 ;
  assign y25445 = ~n40077 ;
  assign y25446 = n43535 ;
  assign y25447 = ~1'b0 ;
  assign y25448 = ~n43539 ;
  assign y25449 = ~n43542 ;
  assign y25450 = ~n43543 ;
  assign y25451 = n43544 ;
  assign y25452 = ~n43545 ;
  assign y25453 = ~1'b0 ;
  assign y25454 = ~1'b0 ;
  assign y25455 = ~1'b0 ;
  assign y25456 = ~1'b0 ;
  assign y25457 = n43547 ;
  assign y25458 = ~n43548 ;
  assign y25459 = ~n43549 ;
  assign y25460 = n152 ;
  assign y25461 = ~1'b0 ;
  assign y25462 = n43552 ;
  assign y25463 = ~n43554 ;
  assign y25464 = ~n43556 ;
  assign y25465 = n43558 ;
  assign y25466 = ~n43559 ;
  assign y25467 = n43561 ;
  assign y25468 = ~n43562 ;
  assign y25469 = n43567 ;
  assign y25470 = ~n3445 ;
  assign y25471 = n43569 ;
  assign y25472 = ~1'b0 ;
  assign y25473 = 1'b0 ;
  assign y25474 = n43572 ;
  assign y25475 = ~n43573 ;
  assign y25476 = ~n43574 ;
  assign y25477 = n43576 ;
  assign y25478 = ~1'b0 ;
  assign y25479 = ~n43577 ;
  assign y25480 = ~1'b0 ;
  assign y25481 = n43579 ;
  assign y25482 = n43580 ;
  assign y25483 = ~n43582 ;
  assign y25484 = ~n43585 ;
  assign y25485 = n43588 ;
  assign y25486 = ~1'b0 ;
  assign y25487 = ~1'b0 ;
  assign y25488 = ~1'b0 ;
  assign y25489 = n43589 ;
  assign y25490 = n43594 ;
  assign y25491 = ~n43595 ;
  assign y25492 = ~n43596 ;
  assign y25493 = ~1'b0 ;
  assign y25494 = n43598 ;
  assign y25495 = n43599 ;
  assign y25496 = n35956 ;
  assign y25497 = ~n43601 ;
  assign y25498 = ~n43605 ;
  assign y25499 = n43607 ;
  assign y25500 = ~1'b0 ;
  assign y25501 = n2776 ;
  assign y25502 = ~1'b0 ;
  assign y25503 = n43609 ;
  assign y25504 = n43611 ;
  assign y25505 = ~n43614 ;
  assign y25506 = ~1'b0 ;
  assign y25507 = ~1'b0 ;
  assign y25508 = ~n43615 ;
  assign y25509 = 1'b0 ;
  assign y25510 = n43620 ;
  assign y25511 = ~1'b0 ;
  assign y25512 = ~1'b0 ;
  assign y25513 = 1'b0 ;
  assign y25514 = ~n43622 ;
  assign y25515 = ~n19032 ;
  assign y25516 = n43630 ;
  assign y25517 = n22828 ;
  assign y25518 = n43631 ;
  assign y25519 = ~n43637 ;
  assign y25520 = ~1'b0 ;
  assign y25521 = ~n43638 ;
  assign y25522 = ~1'b0 ;
  assign y25523 = ~n43640 ;
  assign y25524 = n43641 ;
  assign y25525 = ~n42731 ;
  assign y25526 = n43642 ;
  assign y25527 = ~n43643 ;
  assign y25528 = ~n43644 ;
  assign y25529 = n43645 ;
  assign y25530 = n43647 ;
  assign y25531 = ~n43650 ;
  assign y25532 = n43651 ;
  assign y25533 = ~n43652 ;
  assign y25534 = ~n43653 ;
  assign y25535 = ~1'b0 ;
  assign y25536 = n43654 ;
  assign y25537 = n2250 ;
  assign y25538 = ~1'b0 ;
  assign y25539 = n43658 ;
  assign y25540 = n43659 ;
  assign y25541 = ~n43660 ;
  assign y25542 = ~1'b0 ;
  assign y25543 = ~n43662 ;
  assign y25544 = n43663 ;
  assign y25545 = ~n43664 ;
  assign y25546 = n43665 ;
  assign y25547 = n43670 ;
  assign y25548 = ~1'b0 ;
  assign y25549 = n43674 ;
  assign y25550 = ~n43680 ;
  assign y25551 = n43682 ;
  assign y25552 = ~n43687 ;
  assign y25553 = ~n19433 ;
  assign y25554 = ~1'b0 ;
  assign y25555 = n43688 ;
  assign y25556 = ~1'b0 ;
  assign y25557 = ~n43689 ;
  assign y25558 = ~1'b0 ;
  assign y25559 = ~n43691 ;
  assign y25560 = ~1'b0 ;
  assign y25561 = ~1'b0 ;
  assign y25562 = ~n43692 ;
  assign y25563 = ~n43693 ;
  assign y25564 = ~1'b0 ;
  assign y25565 = ~n43697 ;
  assign y25566 = ~1'b0 ;
  assign y25567 = ~1'b0 ;
  assign y25568 = n43698 ;
  assign y25569 = ~n43701 ;
  assign y25570 = ~1'b0 ;
  assign y25571 = ~n43702 ;
  assign y25572 = n3073 ;
  assign y25573 = n43704 ;
  assign y25574 = ~1'b0 ;
  assign y25575 = n43706 ;
  assign y25576 = ~1'b0 ;
  assign y25577 = ~n43710 ;
  assign y25578 = ~n43712 ;
  assign y25579 = ~n33447 ;
  assign y25580 = ~n43715 ;
  assign y25581 = ~1'b0 ;
  assign y25582 = n43716 ;
  assign y25583 = ~1'b0 ;
  assign y25584 = ~n43717 ;
  assign y25585 = ~1'b0 ;
  assign y25586 = ~1'b0 ;
  assign y25587 = n43721 ;
  assign y25588 = ~1'b0 ;
  assign y25589 = n43725 ;
  assign y25590 = ~n43731 ;
  assign y25591 = ~1'b0 ;
  assign y25592 = ~n43733 ;
  assign y25593 = n43736 ;
  assign y25594 = ~n33890 ;
  assign y25595 = n43738 ;
  assign y25596 = ~n43740 ;
  assign y25597 = ~n43743 ;
  assign y25598 = ~1'b0 ;
  assign y25599 = ~n43744 ;
  assign y25600 = ~n43745 ;
  assign y25601 = n43747 ;
  assign y25602 = n43749 ;
  assign y25603 = n43751 ;
  assign y25604 = ~1'b0 ;
  assign y25605 = ~1'b0 ;
  assign y25606 = ~1'b0 ;
  assign y25607 = ~n43753 ;
  assign y25608 = n43756 ;
  assign y25609 = ~1'b0 ;
  assign y25610 = ~n43757 ;
  assign y25611 = ~1'b0 ;
  assign y25612 = ~1'b0 ;
  assign y25613 = ~n43761 ;
  assign y25614 = ~n43763 ;
  assign y25615 = ~n1347 ;
  assign y25616 = ~n43764 ;
  assign y25617 = ~1'b0 ;
  assign y25618 = ~1'b0 ;
  assign y25619 = ~1'b0 ;
  assign y25620 = ~n43768 ;
  assign y25621 = ~n43773 ;
  assign y25622 = ~n43775 ;
  assign y25623 = n43776 ;
  assign y25624 = n43778 ;
  assign y25625 = ~1'b0 ;
  assign y25626 = n43781 ;
  assign y25627 = ~n43786 ;
  assign y25628 = n43787 ;
  assign y25629 = ~n43789 ;
  assign y25630 = n43790 ;
  assign y25631 = n43791 ;
  assign y25632 = ~1'b0 ;
  assign y25633 = ~1'b0 ;
  assign y25634 = n20174 ;
  assign y25635 = ~n43792 ;
  assign y25636 = n43794 ;
  assign y25637 = ~n43798 ;
  assign y25638 = ~1'b0 ;
  assign y25639 = n43799 ;
  assign y25640 = n43802 ;
  assign y25641 = ~n43806 ;
  assign y25642 = n43807 ;
  assign y25643 = ~n43809 ;
  assign y25644 = ~1'b0 ;
  assign y25645 = ~n43810 ;
  assign y25646 = ~n43811 ;
  assign y25647 = n41777 ;
  assign y25648 = n43818 ;
  assign y25649 = ~1'b0 ;
  assign y25650 = ~1'b0 ;
  assign y25651 = ~n17207 ;
  assign y25652 = n43820 ;
  assign y25653 = n43823 ;
  assign y25654 = ~n12873 ;
  assign y25655 = ~1'b0 ;
  assign y25656 = ~1'b0 ;
  assign y25657 = n43825 ;
  assign y25658 = ~1'b0 ;
  assign y25659 = ~n43826 ;
  assign y25660 = n43827 ;
  assign y25661 = ~1'b0 ;
  assign y25662 = ~1'b0 ;
  assign y25663 = n32521 ;
  assign y25664 = ~1'b0 ;
  assign y25665 = n43828 ;
  assign y25666 = ~1'b0 ;
  assign y25667 = ~1'b0 ;
  assign y25668 = ~1'b0 ;
  assign y25669 = ~n37378 ;
  assign y25670 = ~n43829 ;
  assign y25671 = ~n43831 ;
  assign y25672 = n25937 ;
  assign y25673 = n43832 ;
  assign y25674 = 1'b0 ;
  assign y25675 = ~n43833 ;
  assign y25676 = n43837 ;
  assign y25677 = ~1'b0 ;
  assign y25678 = ~1'b0 ;
  assign y25679 = ~n43839 ;
  assign y25680 = ~1'b0 ;
  assign y25681 = n43840 ;
  assign y25682 = ~n43841 ;
  assign y25683 = n43860 ;
  assign y25684 = ~n1217 ;
  assign y25685 = 1'b0 ;
  assign y25686 = ~n43861 ;
  assign y25687 = ~1'b0 ;
  assign y25688 = ~n37136 ;
  assign y25689 = ~n43862 ;
  assign y25690 = ~n43864 ;
  assign y25691 = n43866 ;
  assign y25692 = ~n43868 ;
  assign y25693 = ~n43869 ;
  assign y25694 = ~n43870 ;
  assign y25695 = ~1'b0 ;
  assign y25696 = n43871 ;
  assign y25697 = ~1'b0 ;
  assign y25698 = n43872 ;
  assign y25699 = ~n43874 ;
  assign y25700 = n11827 ;
  assign y25701 = n43878 ;
  assign y25702 = ~n43879 ;
  assign y25703 = n43884 ;
  assign y25704 = ~1'b0 ;
  assign y25705 = ~n43888 ;
  assign y25706 = n4386 ;
  assign y25707 = n43890 ;
  assign y25708 = ~1'b0 ;
  assign y25709 = n43891 ;
  assign y25710 = n15373 ;
  assign y25711 = n43898 ;
  assign y25712 = ~1'b0 ;
  assign y25713 = ~n43908 ;
  assign y25714 = ~1'b0 ;
  assign y25715 = ~1'b0 ;
  assign y25716 = ~n43909 ;
  assign y25717 = n43911 ;
  assign y25718 = ~n43914 ;
  assign y25719 = n43917 ;
  assign y25720 = ~n43920 ;
  assign y25721 = ~1'b0 ;
  assign y25722 = ~n43923 ;
  assign y25723 = ~n43926 ;
  assign y25724 = ~n43930 ;
  assign y25725 = ~1'b0 ;
  assign y25726 = ~1'b0 ;
  assign y25727 = ~n43931 ;
  assign y25728 = ~n43933 ;
  assign y25729 = ~1'b0 ;
  assign y25730 = n43934 ;
  assign y25731 = ~n2867 ;
  assign y25732 = ~1'b0 ;
  assign y25733 = ~n43936 ;
  assign y25734 = ~n43938 ;
  assign y25735 = n43940 ;
  assign y25736 = ~n43946 ;
  assign y25737 = n43949 ;
  assign y25738 = ~n43950 ;
  assign y25739 = n43954 ;
  assign y25740 = ~n43959 ;
  assign y25741 = ~1'b0 ;
  assign y25742 = ~n4734 ;
  assign y25743 = ~n43960 ;
  assign y25744 = n43961 ;
  assign y25745 = ~1'b0 ;
  assign y25746 = ~1'b0 ;
  assign y25747 = ~n43964 ;
  assign y25748 = ~n43965 ;
  assign y25749 = ~n43967 ;
  assign y25750 = ~1'b0 ;
  assign y25751 = ~1'b0 ;
  assign y25752 = ~n43969 ;
  assign y25753 = ~n43973 ;
  assign y25754 = ~1'b0 ;
  assign y25755 = ~n63 ;
  assign y25756 = ~1'b0 ;
  assign y25757 = n43976 ;
  assign y25758 = n43978 ;
  assign y25759 = n26648 ;
  assign y25760 = ~n43982 ;
  assign y25761 = ~n43983 ;
  assign y25762 = ~1'b0 ;
  assign y25763 = ~1'b0 ;
  assign y25764 = n43986 ;
  assign y25765 = n43989 ;
  assign y25766 = ~n43993 ;
  assign y25767 = n43995 ;
  assign y25768 = n43996 ;
  assign y25769 = n43998 ;
  assign y25770 = ~n44002 ;
  assign y25771 = ~1'b0 ;
  assign y25772 = ~1'b0 ;
  assign y25773 = ~1'b0 ;
  assign y25774 = ~n44005 ;
  assign y25775 = ~1'b0 ;
  assign y25776 = ~1'b0 ;
  assign y25777 = ~n44006 ;
  assign y25778 = ~1'b0 ;
  assign y25779 = n44008 ;
  assign y25780 = n44016 ;
  assign y25781 = ~n44017 ;
  assign y25782 = ~1'b0 ;
  assign y25783 = ~n44018 ;
  assign y25784 = n44021 ;
  assign y25785 = ~n44022 ;
  assign y25786 = ~n44024 ;
  assign y25787 = ~1'b0 ;
  assign y25788 = n44026 ;
  assign y25789 = 1'b0 ;
  assign y25790 = n44028 ;
  assign y25791 = ~1'b0 ;
  assign y25792 = ~1'b0 ;
  assign y25793 = n44031 ;
  assign y25794 = ~n44032 ;
  assign y25795 = ~n44034 ;
  assign y25796 = 1'b0 ;
  assign y25797 = ~n44037 ;
  assign y25798 = ~1'b0 ;
  assign y25799 = ~1'b0 ;
  assign y25800 = n44040 ;
  assign y25801 = n44041 ;
  assign y25802 = n44046 ;
  assign y25803 = ~n44049 ;
  assign y25804 = ~n44051 ;
  assign y25805 = ~1'b0 ;
  assign y25806 = n44052 ;
  assign y25807 = ~n44053 ;
  assign y25808 = ~1'b0 ;
  assign y25809 = ~1'b0 ;
  assign y25810 = n44054 ;
  assign y25811 = n44057 ;
  assign y25812 = ~1'b0 ;
  assign y25813 = n44058 ;
  assign y25814 = ~1'b0 ;
  assign y25815 = n44063 ;
  assign y25816 = n44064 ;
  assign y25817 = ~1'b0 ;
  assign y25818 = n44067 ;
  assign y25819 = ~n44070 ;
  assign y25820 = n44072 ;
  assign y25821 = n44077 ;
  assign y25822 = ~n44079 ;
  assign y25823 = ~1'b0 ;
  assign y25824 = n44081 ;
  assign y25825 = ~1'b0 ;
  assign y25826 = ~1'b0 ;
  assign y25827 = 1'b0 ;
  assign y25828 = ~n44084 ;
  assign y25829 = ~n6415 ;
  assign y25830 = ~n44085 ;
  assign y25831 = ~1'b0 ;
  assign y25832 = ~1'b0 ;
  assign y25833 = ~1'b0 ;
  assign y25834 = ~1'b0 ;
  assign y25835 = ~1'b0 ;
  assign y25836 = ~n44088 ;
  assign y25837 = ~1'b0 ;
  assign y25838 = ~n44089 ;
  assign y25839 = ~1'b0 ;
  assign y25840 = ~n44090 ;
  assign y25841 = n44091 ;
  assign y25842 = ~n44092 ;
  assign y25843 = n44093 ;
  assign y25844 = ~1'b0 ;
  assign y25845 = ~n44094 ;
  assign y25846 = ~n44095 ;
  assign y25847 = ~n44096 ;
  assign y25848 = n44098 ;
  assign y25849 = ~n44100 ;
  assign y25850 = ~n44103 ;
  assign y25851 = ~n43252 ;
  assign y25852 = ~1'b0 ;
  assign y25853 = n44104 ;
  assign y25854 = ~1'b0 ;
  assign y25855 = n44106 ;
  assign y25856 = ~n44108 ;
  assign y25857 = ~1'b0 ;
  assign y25858 = ~n3107 ;
  assign y25859 = ~n44109 ;
  assign y25860 = ~1'b0 ;
  assign y25861 = ~n44110 ;
  assign y25862 = ~n44112 ;
  assign y25863 = n44113 ;
  assign y25864 = ~n44114 ;
  assign y25865 = ~n44116 ;
  assign y25866 = ~1'b0 ;
  assign y25867 = ~n44117 ;
  assign y25868 = ~1'b0 ;
  assign y25869 = ~n3950 ;
  assign y25870 = n44164 ;
  assign y25871 = n36861 ;
  assign y25872 = ~n44166 ;
  assign y25873 = n44167 ;
  assign y25874 = ~n39826 ;
  assign y25875 = ~1'b0 ;
  assign y25876 = ~n44169 ;
  assign y25877 = n44170 ;
  assign y25878 = n44175 ;
  assign y25879 = ~1'b0 ;
  assign y25880 = ~n44178 ;
  assign y25881 = 1'b0 ;
  assign y25882 = ~n44179 ;
  assign y25883 = ~n44180 ;
  assign y25884 = ~n44184 ;
  assign y25885 = n44188 ;
  assign y25886 = ~1'b0 ;
  assign y25887 = ~1'b0 ;
  assign y25888 = ~n44190 ;
  assign y25889 = n18276 ;
  assign y25890 = n44195 ;
  assign y25891 = ~n44196 ;
  assign y25892 = n44199 ;
  assign y25893 = n44200 ;
  assign y25894 = ~n44205 ;
  assign y25895 = ~1'b0 ;
  assign y25896 = ~1'b0 ;
  assign y25897 = 1'b0 ;
  assign y25898 = ~n44206 ;
  assign y25899 = ~n44208 ;
  assign y25900 = ~n44214 ;
  assign y25901 = ~n44217 ;
  assign y25902 = ~n44220 ;
  assign y25903 = ~1'b0 ;
  assign y25904 = n34141 ;
  assign y25905 = n44222 ;
  assign y25906 = n44223 ;
  assign y25907 = ~1'b0 ;
  assign y25908 = n44228 ;
  assign y25909 = ~1'b0 ;
  assign y25910 = n44230 ;
  assign y25911 = ~n44234 ;
  assign y25912 = n44236 ;
  assign y25913 = ~1'b0 ;
  assign y25914 = ~1'b0 ;
  assign y25915 = ~1'b0 ;
  assign y25916 = ~1'b0 ;
  assign y25917 = ~1'b0 ;
  assign y25918 = 1'b0 ;
  assign y25919 = ~n44242 ;
  assign y25920 = n44243 ;
  assign y25921 = n44244 ;
  assign y25922 = n44245 ;
  assign y25923 = ~n44251 ;
  assign y25924 = ~n44253 ;
  assign y25925 = ~n44254 ;
  assign y25926 = ~1'b0 ;
  assign y25927 = n44256 ;
  assign y25928 = ~1'b0 ;
  assign y25929 = ~n44259 ;
  assign y25930 = n44263 ;
  assign y25931 = n5188 ;
  assign y25932 = 1'b0 ;
  assign y25933 = ~n44264 ;
  assign y25934 = ~n44267 ;
  assign y25935 = ~1'b0 ;
  assign y25936 = n44269 ;
  assign y25937 = ~n44273 ;
  assign y25938 = 1'b0 ;
  assign y25939 = 1'b0 ;
  assign y25940 = ~1'b0 ;
  assign y25941 = ~1'b0 ;
  assign y25942 = n7116 ;
  assign y25943 = ~n44274 ;
  assign y25944 = ~n44277 ;
  assign y25945 = n44280 ;
  assign y25946 = n44282 ;
  assign y25947 = ~1'b0 ;
  assign y25948 = n44284 ;
  assign y25949 = ~n20295 ;
  assign y25950 = n44285 ;
  assign y25951 = ~n44288 ;
  assign y25952 = ~n44291 ;
  assign y25953 = n44296 ;
  assign y25954 = ~n44297 ;
  assign y25955 = ~1'b0 ;
  assign y25956 = ~n44298 ;
  assign y25957 = n44302 ;
  assign y25958 = ~n44303 ;
  assign y25959 = ~n44306 ;
  assign y25960 = ~1'b0 ;
  assign y25961 = n44307 ;
  assign y25962 = ~n44308 ;
  assign y25963 = 1'b0 ;
  assign y25964 = ~1'b0 ;
  assign y25965 = ~n44311 ;
  assign y25966 = ~1'b0 ;
  assign y25967 = ~n44312 ;
  assign y25968 = n44313 ;
  assign y25969 = ~n44315 ;
  assign y25970 = n823 ;
  assign y25971 = ~n44317 ;
  assign y25972 = ~1'b0 ;
  assign y25973 = n44318 ;
  assign y25974 = ~n44319 ;
  assign y25975 = ~n44320 ;
  assign y25976 = 1'b0 ;
  assign y25977 = ~1'b0 ;
  assign y25978 = ~1'b0 ;
  assign y25979 = 1'b0 ;
  assign y25980 = ~n44322 ;
  assign y25981 = ~1'b0 ;
  assign y25982 = n44323 ;
  assign y25983 = ~n1237 ;
  assign y25984 = n44328 ;
  assign y25985 = ~n44330 ;
  assign y25986 = n31217 ;
  assign y25987 = n44331 ;
  assign y25988 = n44334 ;
  assign y25989 = ~n44335 ;
  assign y25990 = ~n44337 ;
  assign y25991 = ~1'b0 ;
  assign y25992 = ~n34011 ;
  assign y25993 = n44338 ;
  assign y25994 = n44339 ;
  assign y25995 = ~n44343 ;
  assign y25996 = ~1'b0 ;
  assign y25997 = ~n44344 ;
  assign y25998 = ~n44347 ;
  assign y25999 = n44351 ;
  assign y26000 = n44352 ;
  assign y26001 = ~1'b0 ;
  assign y26002 = n44354 ;
  assign y26003 = n44357 ;
  assign y26004 = ~n44359 ;
  assign y26005 = 1'b0 ;
  assign y26006 = n44360 ;
  assign y26007 = ~1'b0 ;
  assign y26008 = n44361 ;
  assign y26009 = ~n27418 ;
  assign y26010 = ~1'b0 ;
  assign y26011 = n44366 ;
  assign y26012 = n44367 ;
  assign y26013 = ~n39690 ;
  assign y26014 = ~n44368 ;
  assign y26015 = ~n44369 ;
  assign y26016 = ~n44393 ;
  assign y26017 = ~1'b0 ;
  assign y26018 = ~1'b0 ;
  assign y26019 = ~1'b0 ;
  assign y26020 = ~1'b0 ;
  assign y26021 = n44394 ;
  assign y26022 = n44396 ;
  assign y26023 = ~n44397 ;
  assign y26024 = ~n44399 ;
  assign y26025 = n44400 ;
  assign y26026 = ~n22781 ;
  assign y26027 = ~n44401 ;
  assign y26028 = ~n44403 ;
  assign y26029 = n44404 ;
  assign y26030 = ~1'b0 ;
  assign y26031 = ~1'b0 ;
  assign y26032 = ~1'b0 ;
  assign y26033 = n44405 ;
  assign y26034 = n44409 ;
  assign y26035 = n29960 ;
  assign y26036 = n44411 ;
  assign y26037 = ~1'b0 ;
  assign y26038 = n44414 ;
  assign y26039 = n44419 ;
  assign y26040 = ~n44421 ;
  assign y26041 = n44422 ;
  assign y26042 = 1'b0 ;
  assign y26043 = n44424 ;
  assign y26044 = n44426 ;
  assign y26045 = ~1'b0 ;
  assign y26046 = n44428 ;
  assign y26047 = ~1'b0 ;
  assign y26048 = n44429 ;
  assign y26049 = ~1'b0 ;
  assign y26050 = ~n44438 ;
  assign y26051 = n42004 ;
  assign y26052 = n44439 ;
  assign y26053 = ~1'b0 ;
  assign y26054 = n44441 ;
  assign y26055 = ~n44449 ;
  assign y26056 = n44451 ;
  assign y26057 = ~n44453 ;
  assign y26058 = ~1'b0 ;
  assign y26059 = ~n44455 ;
  assign y26060 = ~1'b0 ;
  assign y26061 = ~n44457 ;
  assign y26062 = ~n5886 ;
  assign y26063 = ~1'b0 ;
  assign y26064 = ~n44458 ;
  assign y26065 = n44460 ;
  assign y26066 = ~1'b0 ;
  assign y26067 = ~n44461 ;
  assign y26068 = ~n44463 ;
  assign y26069 = ~1'b0 ;
  assign y26070 = ~n44465 ;
  assign y26071 = ~1'b0 ;
  assign y26072 = n38962 ;
  assign y26073 = ~n44467 ;
  assign y26074 = ~1'b0 ;
  assign y26075 = ~1'b0 ;
  assign y26076 = ~n44469 ;
  assign y26077 = n44470 ;
  assign y26078 = ~n44471 ;
  assign y26079 = n44478 ;
  assign y26080 = ~n44482 ;
  assign y26081 = ~n7357 ;
  assign y26082 = n44483 ;
  assign y26083 = ~n44484 ;
  assign y26084 = n44487 ;
  assign y26085 = n44490 ;
  assign y26086 = n44493 ;
  assign y26087 = n44497 ;
  assign y26088 = n44498 ;
  assign y26089 = ~1'b0 ;
  assign y26090 = ~1'b0 ;
  assign y26091 = n44500 ;
  assign y26092 = ~n44501 ;
  assign y26093 = ~n44503 ;
  assign y26094 = ~1'b0 ;
  assign y26095 = n44505 ;
  assign y26096 = ~n24768 ;
  assign y26097 = ~n44506 ;
  assign y26098 = ~n44510 ;
  assign y26099 = ~n44512 ;
  assign y26100 = ~n44514 ;
  assign y26101 = ~1'b0 ;
  assign y26102 = n44515 ;
  assign y26103 = ~n44517 ;
  assign y26104 = ~n44518 ;
  assign y26105 = n42487 ;
  assign y26106 = n44520 ;
  assign y26107 = ~1'b0 ;
  assign y26108 = ~1'b0 ;
  assign y26109 = ~1'b0 ;
  assign y26110 = n44521 ;
  assign y26111 = ~1'b0 ;
  assign y26112 = ~n13819 ;
  assign y26113 = ~n44523 ;
  assign y26114 = ~n44524 ;
  assign y26115 = n44528 ;
  assign y26116 = n12640 ;
  assign y26117 = n44532 ;
  assign y26118 = ~1'b0 ;
  assign y26119 = n44536 ;
  assign y26120 = ~n44541 ;
  assign y26121 = ~1'b0 ;
  assign y26122 = ~1'b0 ;
  assign y26123 = ~n38973 ;
  assign y26124 = ~1'b0 ;
  assign y26125 = n44542 ;
  assign y26126 = n44543 ;
  assign y26127 = ~n44548 ;
  assign y26128 = ~n44550 ;
  assign y26129 = n5061 ;
  assign y26130 = ~1'b0 ;
  assign y26131 = n44551 ;
  assign y26132 = ~1'b0 ;
  assign y26133 = n44557 ;
  assign y26134 = ~n44558 ;
  assign y26135 = ~n44559 ;
  assign y26136 = n44565 ;
  assign y26137 = ~n44566 ;
  assign y26138 = ~n30951 ;
  assign y26139 = n44570 ;
  assign y26140 = ~n9076 ;
  assign y26141 = ~n26488 ;
  assign y26142 = n44571 ;
  assign y26143 = ~n44573 ;
  assign y26144 = ~n44576 ;
  assign y26145 = ~1'b0 ;
  assign y26146 = ~1'b0 ;
  assign y26147 = ~n44577 ;
  assign y26148 = ~n44578 ;
  assign y26149 = ~1'b0 ;
  assign y26150 = n44580 ;
  assign y26151 = ~1'b0 ;
  assign y26152 = n44583 ;
  assign y26153 = ~1'b0 ;
  assign y26154 = n44585 ;
  assign y26155 = ~n44586 ;
  assign y26156 = ~1'b0 ;
  assign y26157 = n44587 ;
  assign y26158 = ~n37928 ;
  assign y26159 = ~1'b0 ;
  assign y26160 = ~n44591 ;
  assign y26161 = ~1'b0 ;
  assign y26162 = n44592 ;
  assign y26163 = ~1'b0 ;
  assign y26164 = ~n44597 ;
  assign y26165 = ~1'b0 ;
  assign y26166 = ~1'b0 ;
  assign y26167 = ~1'b0 ;
  assign y26168 = n44598 ;
  assign y26169 = ~n44600 ;
  assign y26170 = 1'b0 ;
  assign y26171 = n44601 ;
  assign y26172 = ~n44603 ;
  assign y26173 = n44610 ;
  assign y26174 = n44615 ;
  assign y26175 = n44619 ;
  assign y26176 = ~1'b0 ;
  assign y26177 = ~1'b0 ;
  assign y26178 = n44620 ;
  assign y26179 = n36202 ;
  assign y26180 = 1'b0 ;
  assign y26181 = ~n44622 ;
  assign y26182 = n44627 ;
  assign y26183 = ~n44628 ;
  assign y26184 = n26384 ;
  assign y26185 = ~1'b0 ;
  assign y26186 = n44629 ;
  assign y26187 = ~1'b0 ;
  assign y26188 = ~n44644 ;
  assign y26189 = n44646 ;
  assign y26190 = ~1'b0 ;
  assign y26191 = ~1'b0 ;
  assign y26192 = ~n44647 ;
  assign y26193 = ~1'b0 ;
  assign y26194 = ~1'b0 ;
  assign y26195 = ~n44649 ;
  assign y26196 = n44651 ;
  assign y26197 = ~1'b0 ;
  assign y26198 = ~n44655 ;
  assign y26199 = n44656 ;
  assign y26200 = ~1'b0 ;
  assign y26201 = n4919 ;
  assign y26202 = n44658 ;
  assign y26203 = n44659 ;
  assign y26204 = ~n44661 ;
  assign y26205 = n44664 ;
  assign y26206 = ~1'b0 ;
  assign y26207 = n44666 ;
  assign y26208 = n44670 ;
  assign y26209 = n44674 ;
  assign y26210 = ~1'b0 ;
  assign y26211 = ~n44678 ;
  assign y26212 = ~n44681 ;
  assign y26213 = ~1'b0 ;
  assign y26214 = ~n25612 ;
  assign y26215 = ~n44683 ;
  assign y26216 = ~1'b0 ;
  assign y26217 = n44685 ;
  assign y26218 = ~1'b0 ;
  assign y26219 = ~1'b0 ;
  assign y26220 = ~n44686 ;
  assign y26221 = n44689 ;
  assign y26222 = n44692 ;
  assign y26223 = ~n44694 ;
  assign y26224 = ~1'b0 ;
  assign y26225 = n44699 ;
  assign y26226 = n44706 ;
  assign y26227 = ~1'b0 ;
  assign y26228 = n44711 ;
  assign y26229 = ~n44716 ;
  assign y26230 = ~1'b0 ;
  assign y26231 = n44719 ;
  assign y26232 = ~1'b0 ;
  assign y26233 = ~n44723 ;
  assign y26234 = ~1'b0 ;
  assign y26235 = ~1'b0 ;
  assign y26236 = n44724 ;
  assign y26237 = ~1'b0 ;
  assign y26238 = n44727 ;
  assign y26239 = n44729 ;
  assign y26240 = ~n44730 ;
  assign y26241 = ~1'b0 ;
  assign y26242 = ~n44732 ;
  assign y26243 = n44733 ;
  assign y26244 = ~n44737 ;
  assign y26245 = n44740 ;
  assign y26246 = ~n44741 ;
  assign y26247 = 1'b0 ;
  assign y26248 = ~n44743 ;
  assign y26249 = ~n10359 ;
  assign y26250 = ~n44747 ;
  assign y26251 = ~1'b0 ;
  assign y26252 = ~1'b0 ;
  assign y26253 = ~1'b0 ;
  assign y26254 = ~1'b0 ;
  assign y26255 = n44749 ;
  assign y26256 = ~1'b0 ;
  assign y26257 = ~1'b0 ;
  assign y26258 = ~1'b0 ;
  assign y26259 = ~n44750 ;
  assign y26260 = ~n44751 ;
  assign y26261 = n44753 ;
  assign y26262 = ~n24329 ;
  assign y26263 = ~n15111 ;
  assign y26264 = ~n44754 ;
  assign y26265 = 1'b0 ;
  assign y26266 = ~1'b0 ;
  assign y26267 = ~n44757 ;
  assign y26268 = n44758 ;
  assign y26269 = n44759 ;
  assign y26270 = ~n44761 ;
  assign y26271 = ~n44763 ;
  assign y26272 = ~n44765 ;
  assign y26273 = n44767 ;
  assign y26274 = n44771 ;
  assign y26275 = ~n44773 ;
  assign y26276 = ~1'b0 ;
  assign y26277 = n44774 ;
  assign y26278 = ~1'b0 ;
  assign y26279 = n44777 ;
  assign y26280 = ~1'b0 ;
  assign y26281 = n44779 ;
  assign y26282 = n44780 ;
  assign y26283 = n44783 ;
  assign y26284 = n44785 ;
  assign y26285 = ~n44787 ;
  assign y26286 = ~n44788 ;
  assign y26287 = n44792 ;
  assign y26288 = n5149 ;
  assign y26289 = n35335 ;
  assign y26290 = ~n26112 ;
  assign y26291 = ~1'b0 ;
  assign y26292 = n44793 ;
  assign y26293 = n44794 ;
  assign y26294 = n44796 ;
  assign y26295 = 1'b0 ;
  assign y26296 = ~1'b0 ;
  assign y26297 = ~1'b0 ;
  assign y26298 = ~1'b0 ;
  assign y26299 = 1'b0 ;
  assign y26300 = ~n44800 ;
  assign y26301 = n44802 ;
  assign y26302 = n44803 ;
  assign y26303 = ~1'b0 ;
  assign y26304 = ~1'b0 ;
  assign y26305 = ~n44808 ;
  assign y26306 = ~1'b0 ;
  assign y26307 = n44812 ;
  assign y26308 = ~n44814 ;
  assign y26309 = ~n44815 ;
  assign y26310 = ~1'b0 ;
  assign y26311 = n44817 ;
  assign y26312 = ~n44819 ;
  assign y26313 = ~1'b0 ;
  assign y26314 = ~n18016 ;
  assign y26315 = n4843 ;
  assign y26316 = ~1'b0 ;
  assign y26317 = 1'b0 ;
  assign y26318 = ~n44822 ;
  assign y26319 = ~1'b0 ;
  assign y26320 = n4179 ;
  assign y26321 = ~n44826 ;
  assign y26322 = ~1'b0 ;
  assign y26323 = ~n44827 ;
  assign y26324 = ~n10953 ;
  assign y26325 = ~n44828 ;
  assign y26326 = ~1'b0 ;
  assign y26327 = ~1'b0 ;
  assign y26328 = ~1'b0 ;
  assign y26329 = 1'b0 ;
  assign y26330 = ~n44829 ;
  assign y26331 = ~n44834 ;
  assign y26332 = n44835 ;
  assign y26333 = ~n44837 ;
  assign y26334 = n44839 ;
  assign y26335 = ~1'b0 ;
  assign y26336 = ~n44842 ;
  assign y26337 = n44843 ;
  assign y26338 = n44846 ;
  assign y26339 = ~n40583 ;
  assign y26340 = n44849 ;
  assign y26341 = n44850 ;
  assign y26342 = n44851 ;
  assign y26343 = ~n44853 ;
  assign y26344 = n44854 ;
  assign y26345 = ~1'b0 ;
  assign y26346 = n44856 ;
  assign y26347 = n44857 ;
  assign y26348 = n44858 ;
  assign y26349 = ~1'b0 ;
  assign y26350 = ~1'b0 ;
  assign y26351 = n44860 ;
  assign y26352 = n44862 ;
  assign y26353 = ~n822 ;
  assign y26354 = ~n44863 ;
  assign y26355 = ~1'b0 ;
  assign y26356 = ~n44865 ;
  assign y26357 = n37398 ;
  assign y26358 = ~1'b0 ;
  assign y26359 = ~n44867 ;
  assign y26360 = n44872 ;
  assign y26361 = ~1'b0 ;
  assign y26362 = ~1'b0 ;
  assign y26363 = n44873 ;
  assign y26364 = ~1'b0 ;
  assign y26365 = ~n30933 ;
  assign y26366 = ~1'b0 ;
  assign y26367 = ~n44875 ;
  assign y26368 = ~1'b0 ;
  assign y26369 = ~1'b0 ;
  assign y26370 = ~1'b0 ;
  assign y26371 = ~n9854 ;
  assign y26372 = ~1'b0 ;
  assign y26373 = ~n44880 ;
  assign y26374 = ~1'b0 ;
  assign y26375 = ~n44882 ;
  assign y26376 = n44889 ;
  assign y26377 = n44894 ;
  assign y26378 = ~n44897 ;
  assign y26379 = n44899 ;
  assign y26380 = ~n28697 ;
  assign y26381 = ~n44903 ;
  assign y26382 = ~1'b0 ;
  assign y26383 = ~1'b0 ;
  assign y26384 = ~n44904 ;
  assign y26385 = n44905 ;
  assign y26386 = ~n44906 ;
  assign y26387 = ~n44907 ;
  assign y26388 = ~1'b0 ;
  assign y26389 = n44908 ;
  assign y26390 = ~1'b0 ;
  assign y26391 = n44911 ;
  assign y26392 = n44913 ;
  assign y26393 = ~n44914 ;
  assign y26394 = ~n44915 ;
  assign y26395 = ~n44921 ;
  assign y26396 = ~n26565 ;
  assign y26397 = ~1'b0 ;
  assign y26398 = ~n44922 ;
  assign y26399 = ~n44925 ;
  assign y26400 = ~1'b0 ;
  assign y26401 = ~n44928 ;
  assign y26402 = ~n44929 ;
  assign y26403 = n44930 ;
  assign y26404 = ~1'b0 ;
  assign y26405 = ~1'b0 ;
  assign y26406 = ~1'b0 ;
  assign y26407 = ~1'b0 ;
  assign y26408 = ~1'b0 ;
  assign y26409 = 1'b0 ;
  assign y26410 = ~n44933 ;
  assign y26411 = n44938 ;
  assign y26412 = n44939 ;
  assign y26413 = n44940 ;
  assign y26414 = ~n44944 ;
  assign y26415 = ~n44946 ;
  assign y26416 = ~1'b0 ;
  assign y26417 = ~n10499 ;
  assign y26418 = ~n44950 ;
  assign y26419 = ~1'b0 ;
  assign y26420 = ~n44951 ;
  assign y26421 = ~n44956 ;
  assign y26422 = ~1'b0 ;
  assign y26423 = ~n28618 ;
  assign y26424 = n44961 ;
  assign y26425 = ~1'b0 ;
  assign y26426 = ~n44971 ;
  assign y26427 = ~n44975 ;
  assign y26428 = n44981 ;
  assign y26429 = ~n44985 ;
  assign y26430 = n44987 ;
  assign y26431 = n44988 ;
  assign y26432 = n44989 ;
  assign y26433 = ~1'b0 ;
  assign y26434 = n44990 ;
  assign y26435 = ~1'b0 ;
  assign y26436 = ~1'b0 ;
  assign y26437 = ~1'b0 ;
  assign y26438 = ~1'b0 ;
  assign y26439 = ~n28556 ;
  assign y26440 = ~n44991 ;
  assign y26441 = ~1'b0 ;
  assign y26442 = n44993 ;
  assign y26443 = ~n44995 ;
  assign y26444 = ~1'b0 ;
  assign y26445 = ~n44997 ;
  assign y26446 = n44999 ;
  assign y26447 = ~n45000 ;
  assign y26448 = ~1'b0 ;
  assign y26449 = ~1'b0 ;
  assign y26450 = n45001 ;
  assign y26451 = n45002 ;
  assign y26452 = ~1'b0 ;
  assign y26453 = ~1'b0 ;
  assign y26454 = ~1'b0 ;
  assign y26455 = ~n26573 ;
  assign y26456 = ~1'b0 ;
  assign y26457 = n45004 ;
  assign y26458 = ~1'b0 ;
  assign y26459 = ~n17686 ;
  assign y26460 = ~n45006 ;
  assign y26461 = ~1'b0 ;
  assign y26462 = ~1'b0 ;
  assign y26463 = ~n45009 ;
  assign y26464 = ~n45013 ;
  assign y26465 = ~n41028 ;
  assign y26466 = ~1'b0 ;
  assign y26467 = ~1'b0 ;
  assign y26468 = ~1'b0 ;
  assign y26469 = n45014 ;
  assign y26470 = ~n45015 ;
  assign y26471 = ~1'b0 ;
  assign y26472 = ~n45018 ;
  assign y26473 = ~1'b0 ;
  assign y26474 = n45019 ;
  assign y26475 = n45021 ;
  assign y26476 = n45022 ;
  assign y26477 = n45024 ;
  assign y26478 = ~1'b0 ;
  assign y26479 = ~1'b0 ;
  assign y26480 = 1'b0 ;
  assign y26481 = n45025 ;
  assign y26482 = ~n45027 ;
  assign y26483 = ~n8253 ;
  assign y26484 = n45028 ;
  assign y26485 = n45030 ;
  assign y26486 = ~n45036 ;
  assign y26487 = ~1'b0 ;
  assign y26488 = n45038 ;
  assign y26489 = n45039 ;
  assign y26490 = ~n45040 ;
  assign y26491 = n45044 ;
  assign y26492 = n45045 ;
  assign y26493 = ~n45050 ;
  assign y26494 = n45054 ;
  assign y26495 = ~n45056 ;
  assign y26496 = ~n45057 ;
  assign y26497 = ~1'b0 ;
  assign y26498 = ~n45060 ;
  assign y26499 = ~1'b0 ;
  assign y26500 = n45063 ;
  assign y26501 = ~n45065 ;
  assign y26502 = ~1'b0 ;
  assign y26503 = ~n45067 ;
  assign y26504 = ~n45068 ;
  assign y26505 = n45069 ;
  assign y26506 = ~n45072 ;
  assign y26507 = ~1'b0 ;
  assign y26508 = ~1'b0 ;
  assign y26509 = ~n45076 ;
  assign y26510 = n45078 ;
  assign y26511 = n45079 ;
  assign y26512 = ~n30819 ;
  assign y26513 = ~n45080 ;
  assign y26514 = n45081 ;
  assign y26515 = n45087 ;
  assign y26516 = n45088 ;
  assign y26517 = ~1'b0 ;
  assign y26518 = ~n45092 ;
  assign y26519 = ~n45094 ;
  assign y26520 = ~n45098 ;
  assign y26521 = ~1'b0 ;
  assign y26522 = ~n45100 ;
  assign y26523 = ~1'b0 ;
  assign y26524 = ~n45104 ;
  assign y26525 = ~n45105 ;
  assign y26526 = n45106 ;
  assign y26527 = ~1'b0 ;
  assign y26528 = ~n45107 ;
  assign y26529 = ~1'b0 ;
  assign y26530 = ~n45111 ;
  assign y26531 = ~n45112 ;
  assign y26532 = n45115 ;
  assign y26533 = n45116 ;
  assign y26534 = n45117 ;
  assign y26535 = ~1'b0 ;
  assign y26536 = ~n45118 ;
  assign y26537 = ~1'b0 ;
  assign y26538 = ~1'b0 ;
  assign y26539 = ~1'b0 ;
  assign y26540 = n45119 ;
  assign y26541 = n45121 ;
  assign y26542 = ~n45125 ;
  assign y26543 = n45128 ;
  assign y26544 = n45129 ;
  assign y26545 = 1'b0 ;
  assign y26546 = 1'b0 ;
  assign y26547 = ~n45132 ;
  assign y26548 = ~1'b0 ;
  assign y26549 = ~n45134 ;
  assign y26550 = ~n45137 ;
  assign y26551 = ~1'b0 ;
  assign y26552 = ~1'b0 ;
  assign y26553 = n45142 ;
  assign y26554 = n45144 ;
  assign y26555 = ~1'b0 ;
  assign y26556 = ~1'b0 ;
  assign y26557 = n45146 ;
  assign y26558 = n45148 ;
  assign y26559 = ~1'b0 ;
  assign y26560 = n45150 ;
  assign y26561 = n45153 ;
  assign y26562 = n45156 ;
  assign y26563 = 1'b0 ;
  assign y26564 = n45158 ;
  assign y26565 = ~n45163 ;
  assign y26566 = ~n45169 ;
  assign y26567 = n45170 ;
  assign y26568 = 1'b0 ;
  assign y26569 = ~1'b0 ;
  assign y26570 = n45171 ;
  assign y26571 = n45172 ;
  assign y26572 = ~n45173 ;
  assign y26573 = ~n45175 ;
  assign y26574 = ~1'b0 ;
  assign y26575 = n45178 ;
  assign y26576 = ~1'b0 ;
  assign y26577 = ~1'b0 ;
  assign y26578 = ~n14830 ;
  assign y26579 = ~n45181 ;
  assign y26580 = n45182 ;
  assign y26581 = n45192 ;
  assign y26582 = ~n302 ;
  assign y26583 = ~n45193 ;
  assign y26584 = ~1'b0 ;
  assign y26585 = n45194 ;
  assign y26586 = ~1'b0 ;
  assign y26587 = ~1'b0 ;
  assign y26588 = ~n45197 ;
  assign y26589 = ~1'b0 ;
  assign y26590 = n45199 ;
  assign y26591 = ~1'b0 ;
  assign y26592 = n45202 ;
  assign y26593 = n45204 ;
  assign y26594 = n45205 ;
  assign y26595 = ~n45208 ;
  assign y26596 = n45210 ;
  assign y26597 = ~n45211 ;
  assign y26598 = ~1'b0 ;
  assign y26599 = ~1'b0 ;
  assign y26600 = n45212 ;
  assign y26601 = n5181 ;
  assign y26602 = ~1'b0 ;
  assign y26603 = 1'b0 ;
  assign y26604 = ~n45215 ;
  assign y26605 = n45217 ;
  assign y26606 = n45220 ;
  assign y26607 = ~n45222 ;
  assign y26608 = ~1'b0 ;
  assign y26609 = ~1'b0 ;
  assign y26610 = ~1'b0 ;
  assign y26611 = ~n45223 ;
  assign y26612 = ~1'b0 ;
  assign y26613 = ~n45225 ;
  assign y26614 = ~n45231 ;
  assign y26615 = n45237 ;
  assign y26616 = ~1'b0 ;
  assign y26617 = ~1'b0 ;
  assign y26618 = ~1'b0 ;
  assign y26619 = ~1'b0 ;
  assign y26620 = n45238 ;
  assign y26621 = n45239 ;
  assign y26622 = n45240 ;
  assign y26623 = 1'b0 ;
  assign y26624 = n45245 ;
  assign y26625 = n45251 ;
  assign y26626 = ~1'b0 ;
  assign y26627 = ~1'b0 ;
  assign y26628 = n45255 ;
  assign y26629 = ~1'b0 ;
  assign y26630 = ~n12480 ;
  assign y26631 = ~n45258 ;
  assign y26632 = ~n45260 ;
  assign y26633 = ~1'b0 ;
  assign y26634 = ~1'b0 ;
  assign y26635 = n45262 ;
  assign y26636 = n45263 ;
  assign y26637 = ~n45264 ;
  assign y26638 = ~1'b0 ;
  assign y26639 = ~n45265 ;
  assign y26640 = n45267 ;
  assign y26641 = 1'b0 ;
  assign y26642 = n45268 ;
  assign y26643 = ~1'b0 ;
  assign y26644 = ~1'b0 ;
  assign y26645 = ~n45269 ;
  assign y26646 = ~1'b0 ;
  assign y26647 = n45271 ;
  assign y26648 = ~1'b0 ;
  assign y26649 = ~1'b0 ;
  assign y26650 = ~n45272 ;
  assign y26651 = n45275 ;
  assign y26652 = ~n45277 ;
  assign y26653 = ~n45279 ;
  assign y26654 = ~n45284 ;
  assign y26655 = n45286 ;
  assign y26656 = ~1'b0 ;
  assign y26657 = n45287 ;
  assign y26658 = ~n23435 ;
  assign y26659 = ~n45291 ;
  assign y26660 = ~1'b0 ;
  assign y26661 = n45293 ;
  assign y26662 = ~1'b0 ;
  assign y26663 = ~1'b0 ;
  assign y26664 = ~n45294 ;
  assign y26665 = ~n45299 ;
  assign y26666 = ~n45301 ;
  assign y26667 = n45304 ;
  assign y26668 = 1'b0 ;
  assign y26669 = ~n45307 ;
  assign y26670 = n45309 ;
  assign y26671 = n1991 ;
  assign y26672 = ~n45313 ;
  assign y26673 = ~1'b0 ;
  assign y26674 = ~1'b0 ;
  assign y26675 = ~1'b0 ;
  assign y26676 = n16854 ;
  assign y26677 = n45316 ;
  assign y26678 = ~n45317 ;
  assign y26679 = ~n10835 ;
  assign y26680 = ~n45318 ;
  assign y26681 = ~n45322 ;
  assign y26682 = n45324 ;
  assign y26683 = ~n45326 ;
  assign y26684 = ~1'b0 ;
  assign y26685 = ~1'b0 ;
  assign y26686 = n45327 ;
  assign y26687 = ~1'b0 ;
  assign y26688 = ~1'b0 ;
  assign y26689 = ~n45328 ;
  assign y26690 = n45330 ;
  assign y26691 = ~n45331 ;
  assign y26692 = ~1'b0 ;
  assign y26693 = ~n45335 ;
  assign y26694 = n6622 ;
  assign y26695 = n10141 ;
  assign y26696 = 1'b0 ;
  assign y26697 = ~1'b0 ;
  assign y26698 = n45336 ;
  assign y26699 = ~1'b0 ;
  assign y26700 = 1'b0 ;
  assign y26701 = ~1'b0 ;
  assign y26702 = ~1'b0 ;
  assign y26703 = n45338 ;
  assign y26704 = n45340 ;
  assign y26705 = n45344 ;
  assign y26706 = ~n45345 ;
  assign y26707 = ~n45346 ;
  assign y26708 = ~n45347 ;
  assign y26709 = n45350 ;
  assign y26710 = ~n45352 ;
  assign y26711 = ~1'b0 ;
  assign y26712 = n6613 ;
  assign y26713 = ~1'b0 ;
  assign y26714 = ~1'b0 ;
  assign y26715 = ~n45353 ;
  assign y26716 = ~1'b0 ;
  assign y26717 = ~1'b0 ;
  assign y26718 = ~n45354 ;
  assign y26719 = n45355 ;
  assign y26720 = ~n45356 ;
  assign y26721 = ~1'b0 ;
  assign y26722 = n45357 ;
  assign y26723 = ~1'b0 ;
  assign y26724 = n4629 ;
  assign y26725 = ~n45360 ;
  assign y26726 = ~1'b0 ;
  assign y26727 = n45361 ;
  assign y26728 = n45365 ;
  assign y26729 = ~n45368 ;
  assign y26730 = n33507 ;
  assign y26731 = ~n45371 ;
  assign y26732 = ~1'b0 ;
  assign y26733 = n45375 ;
  assign y26734 = ~1'b0 ;
  assign y26735 = ~n28606 ;
  assign y26736 = ~n45377 ;
  assign y26737 = ~n45382 ;
  assign y26738 = ~n21066 ;
  assign y26739 = ~n681 ;
  assign y26740 = n45384 ;
  assign y26741 = n45387 ;
  assign y26742 = ~1'b0 ;
  assign y26743 = ~n45389 ;
  assign y26744 = n45393 ;
  assign y26745 = ~1'b0 ;
  assign y26746 = ~n45399 ;
  assign y26747 = n45401 ;
  assign y26748 = ~n45402 ;
  assign y26749 = n45404 ;
  assign y26750 = n45406 ;
  assign y26751 = ~1'b0 ;
  assign y26752 = n45408 ;
  assign y26753 = ~1'b0 ;
  assign y26754 = n45411 ;
  assign y26755 = ~n45413 ;
  assign y26756 = n45414 ;
  assign y26757 = n28878 ;
  assign y26758 = ~1'b0 ;
  assign y26759 = ~n45418 ;
  assign y26760 = n45421 ;
  assign y26761 = n45423 ;
  assign y26762 = ~1'b0 ;
  assign y26763 = n1446 ;
  assign y26764 = ~1'b0 ;
  assign y26765 = n45427 ;
  assign y26766 = ~n45431 ;
  assign y26767 = ~n45432 ;
  assign y26768 = ~n45434 ;
  assign y26769 = ~1'b0 ;
  assign y26770 = ~n45436 ;
  assign y26771 = n45437 ;
  assign y26772 = n45442 ;
  assign y26773 = n45444 ;
  assign y26774 = ~n45446 ;
  assign y26775 = ~n45450 ;
  assign y26776 = n45453 ;
  assign y26777 = ~n45457 ;
  assign y26778 = ~n45460 ;
  assign y26779 = ~1'b0 ;
  assign y26780 = ~n29407 ;
  assign y26781 = ~n45461 ;
  assign y26782 = 1'b0 ;
  assign y26783 = n45463 ;
  assign y26784 = n45464 ;
  assign y26785 = ~n45466 ;
  assign y26786 = ~n45467 ;
  assign y26787 = ~n45469 ;
  assign y26788 = n45471 ;
  assign y26789 = ~n45479 ;
  assign y26790 = n45483 ;
  assign y26791 = ~n45488 ;
  assign y26792 = ~1'b0 ;
  assign y26793 = ~1'b0 ;
  assign y26794 = ~n45489 ;
  assign y26795 = ~n45490 ;
  assign y26796 = ~n45491 ;
  assign y26797 = n38320 ;
  assign y26798 = n45494 ;
  assign y26799 = ~n45496 ;
  assign y26800 = ~1'b0 ;
  assign y26801 = n45500 ;
  assign y26802 = ~1'b0 ;
  assign y26803 = 1'b0 ;
  assign y26804 = n45501 ;
  assign y26805 = n45503 ;
  assign y26806 = ~1'b0 ;
  assign y26807 = ~1'b0 ;
  assign y26808 = ~n45506 ;
  assign y26809 = ~1'b0 ;
  assign y26810 = ~1'b0 ;
  assign y26811 = ~1'b0 ;
  assign y26812 = ~1'b0 ;
  assign y26813 = ~1'b0 ;
  assign y26814 = ~n45512 ;
  assign y26815 = ~1'b0 ;
  assign y26816 = ~1'b0 ;
  assign y26817 = ~n45517 ;
  assign y26818 = n45519 ;
  assign y26819 = ~n45522 ;
  assign y26820 = ~1'b0 ;
  assign y26821 = ~1'b0 ;
  assign y26822 = n45524 ;
  assign y26823 = ~n45526 ;
  assign y26824 = n45528 ;
  assign y26825 = ~1'b0 ;
  assign y26826 = ~1'b0 ;
  assign y26827 = n45530 ;
  assign y26828 = n45532 ;
  assign y26829 = 1'b0 ;
  assign y26830 = n45534 ;
  assign y26831 = ~1'b0 ;
  assign y26832 = n45542 ;
  assign y26833 = ~1'b0 ;
  assign y26834 = ~1'b0 ;
  assign y26835 = n45543 ;
  assign y26836 = ~1'b0 ;
  assign y26837 = ~n31361 ;
  assign y26838 = 1'b0 ;
  assign y26839 = 1'b0 ;
  assign y26840 = ~1'b0 ;
  assign y26841 = n45544 ;
  assign y26842 = n45545 ;
  assign y26843 = n45547 ;
  assign y26844 = n45548 ;
  assign y26845 = n4616 ;
  assign y26846 = ~n45550 ;
  assign y26847 = n45551 ;
  assign y26848 = ~1'b0 ;
  assign y26849 = n45555 ;
  assign y26850 = n45556 ;
  assign y26851 = ~n23208 ;
  assign y26852 = ~1'b0 ;
  assign y26853 = ~n45557 ;
  assign y26854 = ~n45558 ;
  assign y26855 = n45559 ;
  assign y26856 = ~1'b0 ;
  assign y26857 = ~1'b0 ;
  assign y26858 = ~1'b0 ;
  assign y26859 = ~1'b0 ;
  assign y26860 = n45561 ;
  assign y26861 = 1'b0 ;
  assign y26862 = ~n45562 ;
  assign y26863 = n45563 ;
  assign y26864 = ~n7067 ;
  assign y26865 = ~n45565 ;
  assign y26866 = ~1'b0 ;
  assign y26867 = n45566 ;
  assign y26868 = ~1'b0 ;
  assign y26869 = n45570 ;
  assign y26870 = ~1'b0 ;
  assign y26871 = ~1'b0 ;
  assign y26872 = ~n45571 ;
  assign y26873 = ~n45572 ;
  assign y26874 = ~n45575 ;
  assign y26875 = ~n45576 ;
  assign y26876 = ~1'b0 ;
  assign y26877 = ~1'b0 ;
  assign y26878 = ~n45577 ;
  assign y26879 = n45578 ;
  assign y26880 = ~1'b0 ;
  assign y26881 = n45579 ;
  assign y26882 = ~n45581 ;
  assign y26883 = ~n45588 ;
  assign y26884 = ~n45589 ;
  assign y26885 = n45590 ;
  assign y26886 = ~n2833 ;
  assign y26887 = n45593 ;
  assign y26888 = ~n45595 ;
  assign y26889 = x5 ;
  assign y26890 = ~1'b0 ;
  assign y26891 = ~n45597 ;
  assign y26892 = ~n2408 ;
  assign y26893 = ~n45598 ;
  assign y26894 = ~n43750 ;
  assign y26895 = ~n45599 ;
  assign y26896 = n45605 ;
  assign y26897 = ~1'b0 ;
  assign y26898 = n45608 ;
  assign y26899 = ~n45615 ;
  assign y26900 = n45616 ;
  assign y26901 = ~n45620 ;
  assign y26902 = n1419 ;
  assign y26903 = ~n45623 ;
  assign y26904 = ~n45625 ;
  assign y26905 = n45628 ;
  assign y26906 = ~1'b0 ;
  assign y26907 = n45632 ;
  assign y26908 = ~1'b0 ;
  assign y26909 = n45636 ;
  assign y26910 = ~n45638 ;
  assign y26911 = ~n13092 ;
  assign y26912 = ~1'b0 ;
  assign y26913 = ~n44740 ;
  assign y26914 = ~1'b0 ;
  assign y26915 = ~n45642 ;
  assign y26916 = ~1'b0 ;
  assign y26917 = n45643 ;
  assign y26918 = ~n45644 ;
  assign y26919 = ~n16253 ;
  assign y26920 = n10399 ;
  assign y26921 = ~1'b0 ;
  assign y26922 = ~1'b0 ;
  assign y26923 = ~1'b0 ;
  assign y26924 = n45646 ;
  assign y26925 = n45648 ;
  assign y26926 = ~1'b0 ;
  assign y26927 = n45650 ;
  assign y26928 = ~1'b0 ;
  assign y26929 = ~1'b0 ;
  assign y26930 = ~n45653 ;
  assign y26931 = ~1'b0 ;
  assign y26932 = n45655 ;
  assign y26933 = ~n45657 ;
  assign y26934 = n45658 ;
  assign y26935 = ~1'b0 ;
  assign y26936 = n45661 ;
  assign y26937 = n45662 ;
  assign y26938 = ~n45670 ;
  assign y26939 = ~1'b0 ;
  assign y26940 = ~n45673 ;
  assign y26941 = ~1'b0 ;
  assign y26942 = ~1'b0 ;
  assign y26943 = n45675 ;
  assign y26944 = ~n45676 ;
  assign y26945 = n45679 ;
  assign y26946 = n45683 ;
  assign y26947 = n45684 ;
  assign y26948 = ~1'b0 ;
  assign y26949 = ~1'b0 ;
  assign y26950 = ~1'b0 ;
  assign y26951 = n45686 ;
  assign y26952 = ~1'b0 ;
  assign y26953 = n45687 ;
  assign y26954 = ~n45688 ;
  assign y26955 = ~n45690 ;
  assign y26956 = n45693 ;
  assign y26957 = ~n45697 ;
  assign y26958 = ~n45699 ;
  assign y26959 = n45702 ;
  assign y26960 = ~n45705 ;
  assign y26961 = 1'b0 ;
  assign y26962 = n45706 ;
  assign y26963 = n45708 ;
  assign y26964 = ~1'b0 ;
  assign y26965 = ~n45709 ;
  assign y26966 = ~n45710 ;
  assign y26967 = n45711 ;
  assign y26968 = ~n45712 ;
  assign y26969 = ~1'b0 ;
  assign y26970 = 1'b0 ;
  assign y26971 = n45715 ;
  assign y26972 = ~n45719 ;
  assign y26973 = ~n39576 ;
  assign y26974 = ~1'b0 ;
  assign y26975 = ~1'b0 ;
  assign y26976 = ~n45721 ;
  assign y26977 = ~1'b0 ;
  assign y26978 = ~n45724 ;
  assign y26979 = n45727 ;
  assign y26980 = ~1'b0 ;
  assign y26981 = ~1'b0 ;
  assign y26982 = ~n45729 ;
  assign y26983 = ~n45732 ;
  assign y26984 = ~n45733 ;
  assign y26985 = ~n45734 ;
  assign y26986 = 1'b0 ;
  assign y26987 = n45735 ;
  assign y26988 = ~1'b0 ;
  assign y26989 = ~1'b0 ;
  assign y26990 = ~1'b0 ;
  assign y26991 = n45736 ;
  assign y26992 = ~n45741 ;
  assign y26993 = n45742 ;
  assign y26994 = n45745 ;
  assign y26995 = ~n45746 ;
  assign y26996 = ~n45752 ;
  assign y26997 = n45754 ;
  assign y26998 = ~1'b0 ;
  assign y26999 = ~1'b0 ;
  assign y27000 = ~1'b0 ;
  assign y27001 = ~n45755 ;
  assign y27002 = ~1'b0 ;
  assign y27003 = n45756 ;
  assign y27004 = ~n45757 ;
  assign y27005 = ~n45759 ;
  assign y27006 = n45762 ;
  assign y27007 = ~n45763 ;
  assign y27008 = ~1'b0 ;
  assign y27009 = n45764 ;
  assign y27010 = n45767 ;
  assign y27011 = ~1'b0 ;
  assign y27012 = n45770 ;
  assign y27013 = ~n45775 ;
  assign y27014 = n45776 ;
  assign y27015 = n45777 ;
  assign y27016 = ~1'b0 ;
  assign y27017 = ~1'b0 ;
  assign y27018 = ~1'b0 ;
  assign y27019 = ~1'b0 ;
  assign y27020 = ~1'b0 ;
  assign y27021 = ~n45779 ;
  assign y27022 = ~1'b0 ;
  assign y27023 = ~n24860 ;
  assign y27024 = n45780 ;
  assign y27025 = n45781 ;
  assign y27026 = ~1'b0 ;
  assign y27027 = n45787 ;
  assign y27028 = ~1'b0 ;
  assign y27029 = ~n45788 ;
  assign y27030 = n45789 ;
  assign y27031 = ~1'b0 ;
  assign y27032 = ~n45791 ;
  assign y27033 = n45794 ;
  assign y27034 = ~n45802 ;
  assign y27035 = ~n45804 ;
  assign y27036 = n3790 ;
  assign y27037 = ~1'b0 ;
  assign y27038 = ~n23948 ;
  assign y27039 = 1'b0 ;
  assign y27040 = ~1'b0 ;
  assign y27041 = ~1'b0 ;
  assign y27042 = n45806 ;
  assign y27043 = ~n45810 ;
  assign y27044 = n45812 ;
  assign y27045 = ~n45816 ;
  assign y27046 = ~1'b0 ;
  assign y27047 = ~1'b0 ;
  assign y27048 = ~1'b0 ;
  assign y27049 = ~n45818 ;
  assign y27050 = ~n45819 ;
  assign y27051 = ~1'b0 ;
  assign y27052 = ~n45828 ;
  assign y27053 = ~n45832 ;
  assign y27054 = ~1'b0 ;
  assign y27055 = ~n45833 ;
  assign y27056 = n45836 ;
  assign y27057 = ~1'b0 ;
  assign y27058 = ~n45840 ;
  assign y27059 = ~1'b0 ;
  assign y27060 = ~n4787 ;
  assign y27061 = ~n45842 ;
  assign y27062 = n45846 ;
  assign y27063 = n45850 ;
  assign y27064 = ~n45851 ;
  assign y27065 = n45852 ;
  assign y27066 = ~n45853 ;
  assign y27067 = n45858 ;
  assign y27068 = n45862 ;
  assign y27069 = n45864 ;
  assign y27070 = n45865 ;
  assign y27071 = ~1'b0 ;
  assign y27072 = n45866 ;
  assign y27073 = n24398 ;
  assign y27074 = ~n45867 ;
  assign y27075 = ~1'b0 ;
  assign y27076 = n45868 ;
  assign y27077 = n14676 ;
  assign y27078 = ~1'b0 ;
  assign y27079 = ~1'b0 ;
  assign y27080 = ~1'b0 ;
  assign y27081 = ~n45869 ;
  assign y27082 = ~n45870 ;
  assign y27083 = ~n45874 ;
  assign y27084 = ~1'b0 ;
  assign y27085 = ~n45876 ;
  assign y27086 = ~1'b0 ;
  assign y27087 = n45880 ;
  assign y27088 = n45881 ;
  assign y27089 = ~1'b0 ;
  assign y27090 = ~n3082 ;
  assign y27091 = ~n45883 ;
  assign y27092 = ~n45888 ;
  assign y27093 = ~1'b0 ;
  assign y27094 = n45899 ;
  assign y27095 = ~1'b0 ;
  assign y27096 = ~1'b0 ;
  assign y27097 = n45900 ;
  assign y27098 = n45901 ;
  assign y27099 = n45902 ;
  assign y27100 = n2201 ;
  assign y27101 = ~1'b0 ;
  assign y27102 = n45905 ;
  assign y27103 = ~1'b0 ;
  assign y27104 = n27321 ;
  assign y27105 = ~n45910 ;
  assign y27106 = ~1'b0 ;
  assign y27107 = n45914 ;
  assign y27108 = n45915 ;
  assign y27109 = ~n45917 ;
  assign y27110 = ~1'b0 ;
  assign y27111 = ~1'b0 ;
  assign y27112 = ~n45918 ;
  assign y27113 = ~n45919 ;
  assign y27114 = ~1'b0 ;
  assign y27115 = n45921 ;
  assign y27116 = ~1'b0 ;
  assign y27117 = n45925 ;
  assign y27118 = ~n45932 ;
  assign y27119 = ~1'b0 ;
  assign y27120 = ~1'b0 ;
  assign y27121 = ~1'b0 ;
  assign y27122 = n45937 ;
  assign y27123 = n45941 ;
  assign y27124 = ~n45943 ;
  assign y27125 = ~1'b0 ;
  assign y27126 = n45945 ;
  assign y27127 = n45947 ;
  assign y27128 = ~n30357 ;
  assign y27129 = ~n45950 ;
  assign y27130 = n45951 ;
  assign y27131 = n45957 ;
  assign y27132 = n45958 ;
  assign y27133 = ~1'b0 ;
  assign y27134 = ~n9222 ;
  assign y27135 = ~n45963 ;
  assign y27136 = 1'b0 ;
  assign y27137 = ~n45966 ;
  assign y27138 = ~n45968 ;
  assign y27139 = n1217 ;
  assign y27140 = ~1'b0 ;
  assign y27141 = ~1'b0 ;
  assign y27142 = n45972 ;
  assign y27143 = n45977 ;
  assign y27144 = ~1'b0 ;
  assign y27145 = n45981 ;
  assign y27146 = ~n45982 ;
  assign y27147 = n45983 ;
  assign y27148 = ~n45984 ;
  assign y27149 = ~1'b0 ;
  assign y27150 = ~1'b0 ;
  assign y27151 = ~n45986 ;
  assign y27152 = ~n45991 ;
  assign y27153 = ~n45993 ;
  assign y27154 = ~1'b0 ;
  assign y27155 = ~1'b0 ;
  assign y27156 = n45996 ;
  assign y27157 = ~1'b0 ;
  assign y27158 = n46000 ;
  assign y27159 = n46009 ;
  assign y27160 = ~1'b0 ;
  assign y27161 = n46011 ;
  assign y27162 = n46013 ;
  assign y27163 = ~n46016 ;
  assign y27164 = n46019 ;
  assign y27165 = ~1'b0 ;
  assign y27166 = ~1'b0 ;
  assign y27167 = n46022 ;
  assign y27168 = n46023 ;
  assign y27169 = n46024 ;
  assign y27170 = ~1'b0 ;
  assign y27171 = n46026 ;
  assign y27172 = ~1'b0 ;
  assign y27173 = ~n46027 ;
  assign y27174 = n46028 ;
  assign y27175 = n46029 ;
  assign y27176 = ~1'b0 ;
  assign y27177 = n40286 ;
  assign y27178 = n46032 ;
  assign y27179 = n46033 ;
  assign y27180 = n46035 ;
  assign y27181 = ~n46039 ;
  assign y27182 = ~n46042 ;
  assign y27183 = ~n46043 ;
  assign y27184 = ~n46047 ;
  assign y27185 = n46050 ;
  assign y27186 = 1'b0 ;
  assign y27187 = ~1'b0 ;
  assign y27188 = ~1'b0 ;
  assign y27189 = n46052 ;
  assign y27190 = ~n46054 ;
  assign y27191 = ~n46056 ;
  assign y27192 = n34114 ;
  assign y27193 = ~n46057 ;
  assign y27194 = n46059 ;
  assign y27195 = ~1'b0 ;
  assign y27196 = n46061 ;
  assign y27197 = ~n46063 ;
  assign y27198 = ~n46069 ;
  assign y27199 = n46072 ;
  assign y27200 = ~1'b0 ;
  assign y27201 = n46075 ;
  assign y27202 = n46076 ;
  assign y27203 = ~1'b0 ;
  assign y27204 = ~n17313 ;
  assign y27205 = ~n46078 ;
  assign y27206 = n46079 ;
  assign y27207 = n46080 ;
  assign y27208 = n46082 ;
  assign y27209 = ~n46084 ;
  assign y27210 = ~n3428 ;
  assign y27211 = n31015 ;
  assign y27212 = ~1'b0 ;
  assign y27213 = n19044 ;
  assign y27214 = ~n46086 ;
  assign y27215 = ~n46088 ;
  assign y27216 = n46090 ;
  assign y27217 = ~1'b0 ;
  assign y27218 = 1'b0 ;
  assign y27219 = ~n46092 ;
  assign y27220 = ~n40380 ;
  assign y27221 = n27200 ;
  assign y27222 = ~1'b0 ;
  assign y27223 = n46093 ;
  assign y27224 = n46095 ;
  assign y27225 = n46097 ;
  assign y27226 = ~1'b0 ;
  assign y27227 = ~n46098 ;
  assign y27228 = n46099 ;
  assign y27229 = n39632 ;
  assign y27230 = n46101 ;
  assign y27231 = n46102 ;
  assign y27232 = ~n46103 ;
  assign y27233 = ~1'b0 ;
  assign y27234 = n46105 ;
  assign y27235 = n46107 ;
  assign y27236 = n2574 ;
  assign y27237 = ~1'b0 ;
  assign y27238 = ~n46109 ;
  assign y27239 = ~1'b0 ;
  assign y27240 = n46005 ;
  assign y27241 = n46110 ;
  assign y27242 = n46111 ;
  assign y27243 = n46112 ;
  assign y27244 = ~n46117 ;
  assign y27245 = ~1'b0 ;
  assign y27246 = ~1'b0 ;
  assign y27247 = n42975 ;
  assign y27248 = ~1'b0 ;
  assign y27249 = ~n46118 ;
  assign y27250 = n46121 ;
  assign y27251 = ~n46123 ;
  assign y27252 = n46124 ;
  assign y27253 = ~n46125 ;
  assign y27254 = ~1'b0 ;
  assign y27255 = ~n46129 ;
  assign y27256 = ~1'b0 ;
  assign y27257 = n46134 ;
  assign y27258 = ~1'b0 ;
  assign y27259 = ~1'b0 ;
  assign y27260 = ~1'b0 ;
  assign y27261 = ~n46138 ;
  assign y27262 = ~n42516 ;
  assign y27263 = n46140 ;
  assign y27264 = n46142 ;
  assign y27265 = n46144 ;
  assign y27266 = ~1'b0 ;
  assign y27267 = n46147 ;
  assign y27268 = n46148 ;
  assign y27269 = ~n46149 ;
  assign y27270 = ~1'b0 ;
  assign y27271 = ~1'b0 ;
  assign y27272 = ~n46152 ;
  assign y27273 = n11269 ;
  assign y27274 = ~1'b0 ;
  assign y27275 = n46154 ;
  assign y27276 = n46155 ;
  assign y27277 = n46156 ;
  assign y27278 = n46158 ;
  assign y27279 = ~n6997 ;
  assign y27280 = ~n29248 ;
  assign y27281 = n46162 ;
  assign y27282 = ~1'b0 ;
  assign y27283 = ~1'b0 ;
  assign y27284 = ~1'b0 ;
  assign y27285 = n46165 ;
  assign y27286 = n46170 ;
  assign y27287 = ~1'b0 ;
  assign y27288 = ~1'b0 ;
  assign y27289 = ~n46175 ;
  assign y27290 = ~n46179 ;
  assign y27291 = ~n44239 ;
  assign y27292 = ~n46180 ;
  assign y27293 = 1'b0 ;
  assign y27294 = n46186 ;
  assign y27295 = ~1'b0 ;
  assign y27296 = n26873 ;
  assign y27297 = ~1'b0 ;
  assign y27298 = ~1'b0 ;
  assign y27299 = ~n46190 ;
  assign y27300 = ~1'b0 ;
  assign y27301 = n46193 ;
  assign y27302 = n46196 ;
  assign y27303 = n46202 ;
  assign y27304 = ~1'b0 ;
  assign y27305 = n46203 ;
  assign y27306 = n46204 ;
  assign y27307 = ~n46207 ;
  assign y27308 = 1'b0 ;
  assign y27309 = ~n46209 ;
  assign y27310 = ~1'b0 ;
  assign y27311 = ~1'b0 ;
  assign y27312 = ~n46210 ;
  assign y27313 = n46212 ;
  assign y27314 = ~1'b0 ;
  assign y27315 = n46214 ;
  assign y27316 = n46216 ;
  assign y27317 = ~n46217 ;
  assign y27318 = ~n46218 ;
  assign y27319 = n29914 ;
  assign y27320 = 1'b0 ;
  assign y27321 = n46222 ;
  assign y27322 = n46231 ;
  assign y27323 = ~1'b0 ;
  assign y27324 = ~1'b0 ;
  assign y27325 = ~n46235 ;
  assign y27326 = n46237 ;
  assign y27327 = ~1'b0 ;
  assign y27328 = ~n46241 ;
  assign y27329 = n46242 ;
  assign y27330 = n46243 ;
  assign y27331 = n46245 ;
  assign y27332 = ~1'b0 ;
  assign y27333 = ~n37716 ;
  assign y27334 = n30876 ;
  assign y27335 = ~1'b0 ;
  assign y27336 = ~n46246 ;
  assign y27337 = n46250 ;
  assign y27338 = ~n46251 ;
  assign y27339 = n46253 ;
  assign y27340 = ~1'b0 ;
  assign y27341 = ~n46254 ;
  assign y27342 = ~n46256 ;
  assign y27343 = n46257 ;
  assign y27344 = ~n46259 ;
  assign y27345 = ~n46260 ;
  assign y27346 = n46261 ;
  assign y27347 = ~n46262 ;
  assign y27348 = ~n46263 ;
  assign y27349 = n46264 ;
  assign y27350 = n17114 ;
  assign y27351 = n46267 ;
  assign y27352 = ~1'b0 ;
  assign y27353 = ~1'b0 ;
  assign y27354 = ~n16193 ;
  assign y27355 = ~n46269 ;
  assign y27356 = ~n46273 ;
  assign y27357 = n46275 ;
  assign y27358 = ~n46276 ;
  assign y27359 = ~1'b0 ;
  assign y27360 = ~1'b0 ;
  assign y27361 = n12274 ;
  assign y27362 = ~1'b0 ;
  assign y27363 = n46277 ;
  assign y27364 = 1'b0 ;
  assign y27365 = ~n46278 ;
  assign y27366 = ~1'b0 ;
  assign y27367 = ~n40015 ;
  assign y27368 = ~n46279 ;
  assign y27369 = n46286 ;
  assign y27370 = ~n46287 ;
  assign y27371 = ~n46289 ;
  assign y27372 = ~n46291 ;
  assign y27373 = ~n46293 ;
  assign y27374 = ~1'b0 ;
  assign y27375 = ~1'b0 ;
  assign y27376 = ~1'b0 ;
  assign y27377 = n46296 ;
  assign y27378 = ~n46300 ;
  assign y27379 = ~n46301 ;
  assign y27380 = ~1'b0 ;
  assign y27381 = ~1'b0 ;
  assign y27382 = ~n46304 ;
  assign y27383 = ~1'b0 ;
  assign y27384 = ~n46307 ;
  assign y27385 = ~n46308 ;
  assign y27386 = ~n46309 ;
  assign y27387 = ~n46310 ;
  assign y27388 = n46311 ;
  assign y27389 = n46312 ;
  assign y27390 = n46315 ;
  assign y27391 = ~n46317 ;
  assign y27392 = ~n6512 ;
  assign y27393 = ~n46318 ;
  assign y27394 = n46321 ;
  assign y27395 = ~1'b0 ;
  assign y27396 = ~n46322 ;
  assign y27397 = 1'b0 ;
  assign y27398 = n14731 ;
  assign y27399 = n46324 ;
  assign y27400 = n46325 ;
  assign y27401 = ~1'b0 ;
  assign y27402 = n46328 ;
  assign y27403 = ~n46329 ;
  assign y27404 = ~1'b0 ;
  assign y27405 = ~1'b0 ;
  assign y27406 = ~n46335 ;
  assign y27407 = n46339 ;
  assign y27408 = n46340 ;
  assign y27409 = ~1'b0 ;
  assign y27410 = ~n46345 ;
  assign y27411 = ~1'b0 ;
  assign y27412 = ~1'b0 ;
  assign y27413 = ~n6396 ;
  assign y27414 = ~n46346 ;
  assign y27415 = ~n46347 ;
  assign y27416 = ~n46348 ;
  assign y27417 = ~1'b0 ;
  assign y27418 = n46352 ;
  assign y27419 = ~1'b0 ;
  assign y27420 = 1'b0 ;
  assign y27421 = ~n46355 ;
  assign y27422 = n46358 ;
  assign y27423 = ~n46359 ;
  assign y27424 = ~n46360 ;
  assign y27425 = ~n28199 ;
  assign y27426 = ~1'b0 ;
  assign y27427 = ~n13774 ;
  assign y27428 = ~1'b0 ;
  assign y27429 = ~n46361 ;
  assign y27430 = ~n25091 ;
  assign y27431 = ~n46363 ;
  assign y27432 = ~1'b0 ;
  assign y27433 = ~1'b0 ;
  assign y27434 = n13981 ;
  assign y27435 = n46366 ;
  assign y27436 = n46367 ;
  assign y27437 = ~n46369 ;
  assign y27438 = ~n46374 ;
  assign y27439 = 1'b0 ;
  assign y27440 = n46378 ;
  assign y27441 = n46379 ;
  assign y27442 = ~n23065 ;
  assign y27443 = ~1'b0 ;
  assign y27444 = ~1'b0 ;
  assign y27445 = ~1'b0 ;
  assign y27446 = ~1'b0 ;
  assign y27447 = ~n46380 ;
  assign y27448 = n46381 ;
  assign y27449 = ~1'b0 ;
  assign y27450 = ~1'b0 ;
  assign y27451 = ~1'b0 ;
  assign y27452 = n808 ;
  assign y27453 = ~n46383 ;
  assign y27454 = n46384 ;
  assign y27455 = ~1'b0 ;
  assign y27456 = ~1'b0 ;
  assign y27457 = n46387 ;
  assign y27458 = n46393 ;
  assign y27459 = ~1'b0 ;
  assign y27460 = ~n46395 ;
  assign y27461 = ~n46397 ;
  assign y27462 = n46398 ;
  assign y27463 = ~n46401 ;
  assign y27464 = ~n35428 ;
  assign y27465 = ~1'b0 ;
  assign y27466 = ~1'b0 ;
  assign y27467 = ~n46404 ;
  assign y27468 = ~n15999 ;
  assign y27469 = ~n30521 ;
  assign y27470 = ~1'b0 ;
  assign y27471 = n7589 ;
  assign y27472 = n46411 ;
  assign y27473 = ~1'b0 ;
  assign y27474 = ~1'b0 ;
  assign y27475 = ~n46413 ;
  assign y27476 = ~1'b0 ;
  assign y27477 = ~n39606 ;
  assign y27478 = ~1'b0 ;
  assign y27479 = ~n46415 ;
  assign y27480 = ~n46417 ;
  assign y27481 = ~n46419 ;
  assign y27482 = ~1'b0 ;
  assign y27483 = ~n46421 ;
  assign y27484 = n28438 ;
  assign y27485 = n2570 ;
  assign y27486 = ~n18571 ;
  assign y27487 = ~1'b0 ;
  assign y27488 = n46428 ;
  assign y27489 = ~n46429 ;
  assign y27490 = ~n46431 ;
  assign y27491 = ~1'b0 ;
  assign y27492 = ~1'b0 ;
  assign y27493 = ~n46432 ;
  assign y27494 = ~n6058 ;
  assign y27495 = 1'b0 ;
  assign y27496 = ~n46436 ;
  assign y27497 = ~1'b0 ;
  assign y27498 = ~1'b0 ;
  assign y27499 = n46440 ;
  assign y27500 = ~n10166 ;
  assign y27501 = n46443 ;
  assign y27502 = n46445 ;
  assign y27503 = n46446 ;
  assign y27504 = ~1'b0 ;
  assign y27505 = ~n46447 ;
  assign y27506 = ~n46449 ;
  assign y27507 = ~1'b0 ;
  assign y27508 = n46450 ;
  assign y27509 = ~1'b0 ;
  assign y27510 = ~1'b0 ;
  assign y27511 = ~1'b0 ;
  assign y27512 = ~1'b0 ;
  assign y27513 = n46455 ;
  assign y27514 = n46457 ;
  assign y27515 = ~n46460 ;
  assign y27516 = n45077 ;
  assign y27517 = ~n43804 ;
  assign y27518 = ~1'b0 ;
  assign y27519 = n46461 ;
  assign y27520 = ~n46462 ;
  assign y27521 = 1'b0 ;
  assign y27522 = ~1'b0 ;
  assign y27523 = n46464 ;
  assign y27524 = ~1'b0 ;
  assign y27525 = ~n46465 ;
  assign y27526 = ~1'b0 ;
  assign y27527 = n46471 ;
  assign y27528 = n46477 ;
  assign y27529 = 1'b0 ;
  assign y27530 = ~1'b0 ;
  assign y27531 = ~1'b0 ;
  assign y27532 = n46480 ;
  assign y27533 = ~1'b0 ;
  assign y27534 = n11862 ;
  assign y27535 = ~n46482 ;
  assign y27536 = ~1'b0 ;
  assign y27537 = ~n1868 ;
  assign y27538 = ~1'b0 ;
  assign y27539 = ~1'b0 ;
  assign y27540 = n46486 ;
  assign y27541 = ~1'b0 ;
  assign y27542 = ~1'b0 ;
  assign y27543 = ~1'b0 ;
  assign y27544 = n46487 ;
  assign y27545 = n46488 ;
  assign y27546 = n46494 ;
  assign y27547 = n46496 ;
  assign y27548 = ~1'b0 ;
  assign y27549 = 1'b0 ;
  assign y27550 = ~1'b0 ;
  assign y27551 = n46499 ;
  assign y27552 = ~n46502 ;
  assign y27553 = n46503 ;
  assign y27554 = n11904 ;
  assign y27555 = ~n46504 ;
  assign y27556 = ~1'b0 ;
  assign y27557 = ~n46505 ;
  assign y27558 = ~n46510 ;
  assign y27559 = n46512 ;
  assign y27560 = ~n46514 ;
  assign y27561 = n46516 ;
  assign y27562 = ~1'b0 ;
  assign y27563 = n46520 ;
  assign y27564 = ~n46523 ;
  assign y27565 = n44766 ;
  assign y27566 = n46525 ;
  assign y27567 = ~1'b0 ;
  assign y27568 = ~1'b0 ;
  assign y27569 = ~n46528 ;
  assign y27570 = ~n46529 ;
  assign y27571 = ~n46530 ;
  assign y27572 = ~1'b0 ;
  assign y27573 = ~n46533 ;
  assign y27574 = ~1'b0 ;
  assign y27575 = ~1'b0 ;
  assign y27576 = n46534 ;
  assign y27577 = n30749 ;
  assign y27578 = ~1'b0 ;
  assign y27579 = ~1'b0 ;
  assign y27580 = n46542 ;
  assign y27581 = ~1'b0 ;
  assign y27582 = ~1'b0 ;
  assign y27583 = ~n46543 ;
  assign y27584 = ~n46544 ;
  assign y27585 = ~n46547 ;
  assign y27586 = n22847 ;
  assign y27587 = ~1'b0 ;
  assign y27588 = n46548 ;
  assign y27589 = ~n46550 ;
  assign y27590 = ~n46554 ;
  assign y27591 = ~1'b0 ;
  assign y27592 = ~1'b0 ;
  assign y27593 = n46558 ;
  assign y27594 = n46559 ;
  assign y27595 = ~n46561 ;
  assign y27596 = n46562 ;
  assign y27597 = ~1'b0 ;
  assign y27598 = ~1'b0 ;
  assign y27599 = n46563 ;
  assign y27600 = ~1'b0 ;
  assign y27601 = ~n46565 ;
  assign y27602 = n46566 ;
  assign y27603 = ~n46571 ;
  assign y27604 = ~n46575 ;
  assign y27605 = ~n46579 ;
  assign y27606 = 1'b0 ;
  assign y27607 = n26080 ;
  assign y27608 = ~n46581 ;
  assign y27609 = ~1'b0 ;
  assign y27610 = ~1'b0 ;
  assign y27611 = ~n46583 ;
  assign y27612 = ~n46586 ;
  assign y27613 = n46588 ;
  assign y27614 = ~1'b0 ;
  assign y27615 = 1'b0 ;
  assign y27616 = ~n46590 ;
  assign y27617 = ~1'b0 ;
  assign y27618 = ~n46591 ;
  assign y27619 = ~n46592 ;
  assign y27620 = n23705 ;
  assign y27621 = ~n46602 ;
  assign y27622 = n46605 ;
  assign y27623 = ~n46606 ;
  assign y27624 = ~n46608 ;
  assign y27625 = ~1'b0 ;
  assign y27626 = ~n46611 ;
  assign y27627 = ~n25105 ;
  assign y27628 = n46614 ;
  assign y27629 = ~1'b0 ;
  assign y27630 = n46616 ;
  assign y27631 = ~1'b0 ;
  assign y27632 = ~n46621 ;
  assign y27633 = ~1'b0 ;
  assign y27634 = ~1'b0 ;
  assign y27635 = ~n46622 ;
  assign y27636 = n46623 ;
  assign y27637 = ~n46624 ;
  assign y27638 = n46628 ;
  assign y27639 = ~1'b0 ;
  assign y27640 = ~1'b0 ;
  assign y27641 = ~n46629 ;
  assign y27642 = ~1'b0 ;
  assign y27643 = n46630 ;
  assign y27644 = ~1'b0 ;
  assign y27645 = n46632 ;
  assign y27646 = n18217 ;
  assign y27647 = ~n46634 ;
  assign y27648 = n46636 ;
  assign y27649 = ~n46638 ;
  assign y27650 = ~n46639 ;
  assign y27651 = 1'b0 ;
  assign y27652 = n46641 ;
  assign y27653 = 1'b0 ;
  assign y27654 = n46646 ;
  assign y27655 = n31112 ;
  assign y27656 = ~1'b0 ;
  assign y27657 = ~n46647 ;
  assign y27658 = ~n46649 ;
  assign y27659 = n46653 ;
  assign y27660 = ~n46655 ;
  assign y27661 = ~n46656 ;
  assign y27662 = n46657 ;
  assign y27663 = ~1'b0 ;
  assign y27664 = ~n46660 ;
  assign y27665 = n46662 ;
  assign y27666 = ~n46664 ;
  assign y27667 = 1'b0 ;
  assign y27668 = n46665 ;
  assign y27669 = n5779 ;
  assign y27670 = ~1'b0 ;
  assign y27671 = ~1'b0 ;
  assign y27672 = ~1'b0 ;
  assign y27673 = ~n46666 ;
  assign y27674 = n46668 ;
  assign y27675 = n46671 ;
  assign y27676 = ~n46678 ;
  assign y27677 = n46680 ;
  assign y27678 = n46682 ;
  assign y27679 = n46687 ;
  assign y27680 = n46690 ;
  assign y27681 = ~n46693 ;
  assign y27682 = ~n46694 ;
  assign y27683 = ~1'b0 ;
  assign y27684 = ~n46699 ;
  assign y27685 = ~n46701 ;
  assign y27686 = 1'b0 ;
  assign y27687 = ~n46702 ;
  assign y27688 = ~n46703 ;
  assign y27689 = ~1'b0 ;
  assign y27690 = ~n46704 ;
  assign y27691 = n46706 ;
  assign y27692 = n46709 ;
  assign y27693 = ~1'b0 ;
  assign y27694 = n46711 ;
  assign y27695 = ~n37836 ;
  assign y27696 = ~1'b0 ;
  assign y27697 = ~n20903 ;
  assign y27698 = ~n21289 ;
  assign y27699 = ~n46714 ;
  assign y27700 = ~1'b0 ;
  assign y27701 = n46715 ;
  assign y27702 = ~1'b0 ;
  assign y27703 = ~n46717 ;
  assign y27704 = ~1'b0 ;
  assign y27705 = n46719 ;
  assign y27706 = n46721 ;
  assign y27707 = ~1'b0 ;
  assign y27708 = ~n46722 ;
  assign y27709 = ~1'b0 ;
  assign y27710 = n46723 ;
  assign y27711 = n20289 ;
  assign y27712 = ~1'b0 ;
  assign y27713 = ~1'b0 ;
  assign y27714 = ~n46732 ;
  assign y27715 = 1'b0 ;
  assign y27716 = n46733 ;
  assign y27717 = n46734 ;
  assign y27718 = ~n46735 ;
  assign y27719 = ~1'b0 ;
  assign y27720 = n46737 ;
  assign y27721 = ~n46741 ;
  assign y27722 = ~n31574 ;
  assign y27723 = n46745 ;
  assign y27724 = ~n46747 ;
  assign y27725 = ~n46753 ;
  assign y27726 = n23039 ;
  assign y27727 = ~n46754 ;
  assign y27728 = ~n10340 ;
  assign y27729 = ~1'b0 ;
  assign y27730 = ~n46755 ;
  assign y27731 = ~n46760 ;
  assign y27732 = ~1'b0 ;
  assign y27733 = n46764 ;
  assign y27734 = ~n46765 ;
  assign y27735 = ~1'b0 ;
  assign y27736 = n46766 ;
  assign y27737 = ~n46769 ;
  assign y27738 = ~1'b0 ;
  assign y27739 = n27836 ;
  assign y27740 = ~n46771 ;
  assign y27741 = ~n46777 ;
  assign y27742 = ~1'b0 ;
  assign y27743 = n46779 ;
  assign y27744 = ~1'b0 ;
  assign y27745 = n46780 ;
  assign y27746 = ~1'b0 ;
  assign y27747 = n46783 ;
  assign y27748 = ~n46784 ;
  assign y27749 = n46786 ;
  assign y27750 = ~n46787 ;
  assign y27751 = ~1'b0 ;
  assign y27752 = ~1'b0 ;
  assign y27753 = n46788 ;
  assign y27754 = n46790 ;
  assign y27755 = n46791 ;
  assign y27756 = ~1'b0 ;
  assign y27757 = n22221 ;
  assign y27758 = ~n46792 ;
  assign y27759 = ~n46799 ;
  assign y27760 = n46804 ;
  assign y27761 = 1'b0 ;
  assign y27762 = ~1'b0 ;
  assign y27763 = ~1'b0 ;
  assign y27764 = ~1'b0 ;
  assign y27765 = n46808 ;
  assign y27766 = n46811 ;
  assign y27767 = n46813 ;
  assign y27768 = n46814 ;
  assign y27769 = ~n46831 ;
  assign y27770 = ~1'b0 ;
  assign y27771 = ~1'b0 ;
  assign y27772 = 1'b0 ;
  assign y27773 = n46835 ;
  assign y27774 = ~n19356 ;
  assign y27775 = n46838 ;
  assign y27776 = 1'b0 ;
  assign y27777 = 1'b0 ;
  assign y27778 = ~n46839 ;
  assign y27779 = ~1'b0 ;
  assign y27780 = n46843 ;
  assign y27781 = ~n46848 ;
  assign y27782 = ~n46849 ;
  assign y27783 = ~n46851 ;
  assign y27784 = ~1'b0 ;
  assign y27785 = ~n46853 ;
  assign y27786 = ~1'b0 ;
  assign y27787 = ~n46855 ;
  assign y27788 = ~n46859 ;
  assign y27789 = ~1'b0 ;
  assign y27790 = 1'b0 ;
  assign y27791 = n46862 ;
  assign y27792 = n46863 ;
  assign y27793 = 1'b0 ;
  assign y27794 = n46868 ;
  assign y27795 = ~n46869 ;
  assign y27796 = ~1'b0 ;
  assign y27797 = ~n46870 ;
  assign y27798 = ~n46871 ;
  assign y27799 = n46872 ;
  assign y27800 = ~n46874 ;
  assign y27801 = ~1'b0 ;
  assign y27802 = ~1'b0 ;
  assign y27803 = n46876 ;
  assign y27804 = n46879 ;
  assign y27805 = n46882 ;
  assign y27806 = n46886 ;
  assign y27807 = n46887 ;
  assign y27808 = n46890 ;
  assign y27809 = n46891 ;
  assign y27810 = ~1'b0 ;
  assign y27811 = ~1'b0 ;
  assign y27812 = ~n46893 ;
  assign y27813 = ~n46895 ;
  assign y27814 = ~1'b0 ;
  assign y27815 = n10421 ;
  assign y27816 = ~1'b0 ;
  assign y27817 = ~n46896 ;
  assign y27818 = ~1'b0 ;
  assign y27819 = ~1'b0 ;
  assign y27820 = ~n46902 ;
  assign y27821 = ~n46905 ;
  assign y27822 = ~n46906 ;
  assign y27823 = ~1'b0 ;
  assign y27824 = n46907 ;
  assign y27825 = ~1'b0 ;
  assign y27826 = ~1'b0 ;
  assign y27827 = n46912 ;
  assign y27828 = ~n46913 ;
  assign y27829 = ~n46915 ;
  assign y27830 = ~1'b0 ;
  assign y27831 = 1'b0 ;
  assign y27832 = n46920 ;
  assign y27833 = n46922 ;
  assign y27834 = n32807 ;
  assign y27835 = n46927 ;
  assign y27836 = ~1'b0 ;
  assign y27837 = ~1'b0 ;
  assign y27838 = n46931 ;
  assign y27839 = n45557 ;
  assign y27840 = ~1'b0 ;
  assign y27841 = n4378 ;
  assign y27842 = n46932 ;
  assign y27843 = ~1'b0 ;
  assign y27844 = ~1'b0 ;
  assign y27845 = ~n46935 ;
  assign y27846 = n46936 ;
  assign y27847 = 1'b0 ;
  assign y27848 = ~1'b0 ;
  assign y27849 = ~n46937 ;
  assign y27850 = n10381 ;
  assign y27851 = n46938 ;
  assign y27852 = ~1'b0 ;
  assign y27853 = ~1'b0 ;
  assign y27854 = n46939 ;
  assign y27855 = ~n46945 ;
  assign y27856 = n46946 ;
  assign y27857 = ~n46949 ;
  assign y27858 = ~1'b0 ;
  assign y27859 = ~n46955 ;
  assign y27860 = ~n46956 ;
  assign y27861 = ~n46963 ;
  assign y27862 = n46964 ;
  assign y27863 = ~1'b0 ;
  assign y27864 = ~1'b0 ;
  assign y27865 = ~1'b0 ;
  assign y27866 = ~1'b0 ;
  assign y27867 = n46966 ;
  assign y27868 = n46967 ;
  assign y27869 = n46971 ;
  assign y27870 = ~n46974 ;
  assign y27871 = n46978 ;
  assign y27872 = ~n46979 ;
  assign y27873 = ~1'b0 ;
  assign y27874 = ~n46980 ;
  assign y27875 = n46984 ;
  assign y27876 = n46985 ;
  assign y27877 = ~1'b0 ;
  assign y27878 = ~1'b0 ;
  assign y27879 = ~1'b0 ;
  assign y27880 = n35023 ;
  assign y27881 = n46986 ;
  assign y27882 = n46989 ;
  assign y27883 = ~n46990 ;
  assign y27884 = ~n46992 ;
  assign y27885 = ~n46996 ;
  assign y27886 = n46997 ;
  assign y27887 = n46998 ;
  assign y27888 = ~1'b0 ;
  assign y27889 = n47000 ;
  assign y27890 = ~n45930 ;
  assign y27891 = n47005 ;
  assign y27892 = n47006 ;
  assign y27893 = n47012 ;
  assign y27894 = ~1'b0 ;
  assign y27895 = ~n47015 ;
  assign y27896 = n47016 ;
  assign y27897 = ~n47019 ;
  assign y27898 = n47024 ;
  assign y27899 = ~n14325 ;
  assign y27900 = ~n47027 ;
  assign y27901 = ~1'b0 ;
  assign y27902 = n47030 ;
  assign y27903 = ~n47032 ;
  assign y27904 = ~n11257 ;
  assign y27905 = ~n47035 ;
  assign y27906 = n47036 ;
  assign y27907 = ~1'b0 ;
  assign y27908 = n47041 ;
  assign y27909 = n47042 ;
  assign y27910 = n47043 ;
  assign y27911 = ~n47046 ;
  assign y27912 = ~1'b0 ;
  assign y27913 = ~n47047 ;
  assign y27914 = n47049 ;
  assign y27915 = ~1'b0 ;
  assign y27916 = ~1'b0 ;
  assign y27917 = n1285 ;
  assign y27918 = ~1'b0 ;
  assign y27919 = ~n47051 ;
  assign y27920 = n47055 ;
  assign y27921 = n47057 ;
  assign y27922 = ~1'b0 ;
  assign y27923 = ~n47059 ;
  assign y27924 = ~n47061 ;
  assign y27925 = ~n47063 ;
  assign y27926 = ~1'b0 ;
  assign y27927 = ~n3423 ;
  assign y27928 = n47064 ;
  assign y27929 = n47065 ;
  assign y27930 = ~1'b0 ;
  assign y27931 = n47070 ;
  assign y27932 = n451 ;
  assign y27933 = ~n47072 ;
  assign y27934 = n47078 ;
  assign y27935 = n47087 ;
  assign y27936 = ~1'b0 ;
  assign y27937 = ~n47088 ;
  assign y27938 = ~1'b0 ;
  assign y27939 = n47089 ;
  assign y27940 = n4540 ;
  assign y27941 = ~1'b0 ;
  assign y27942 = ~n47110 ;
  assign y27943 = 1'b0 ;
  assign y27944 = ~1'b0 ;
  assign y27945 = n47111 ;
  assign y27946 = ~n47112 ;
  assign y27947 = ~n47115 ;
  assign y27948 = n47116 ;
  assign y27949 = 1'b0 ;
  assign y27950 = ~n47120 ;
  assign y27951 = ~1'b0 ;
  assign y27952 = n47121 ;
  assign y27953 = ~n47125 ;
  assign y27954 = ~n47126 ;
  assign y27955 = n23688 ;
  assign y27956 = n47129 ;
  assign y27957 = ~n47130 ;
  assign y27958 = ~1'b0 ;
  assign y27959 = n47134 ;
  assign y27960 = n47137 ;
  assign y27961 = ~n47139 ;
  assign y27962 = n47142 ;
  assign y27963 = ~1'b0 ;
  assign y27964 = 1'b0 ;
  assign y27965 = ~1'b0 ;
  assign y27966 = n47144 ;
  assign y27967 = n47145 ;
  assign y27968 = n47149 ;
  assign y27969 = ~1'b0 ;
  assign y27970 = ~1'b0 ;
  assign y27971 = n47151 ;
  assign y27972 = n47155 ;
  assign y27973 = ~n47157 ;
  assign y27974 = n47158 ;
  assign y27975 = n47159 ;
  assign y27976 = ~n47161 ;
  assign y27977 = ~n45979 ;
  assign y27978 = n47163 ;
  assign y27979 = n47164 ;
  assign y27980 = ~n47168 ;
  assign y27981 = 1'b0 ;
  assign y27982 = ~1'b0 ;
  assign y27983 = ~1'b0 ;
  assign y27984 = ~n47170 ;
  assign y27985 = ~1'b0 ;
  assign y27986 = ~n47176 ;
  assign y27987 = n47178 ;
  assign y27988 = ~n47179 ;
  assign y27989 = ~n47180 ;
  assign y27990 = n47183 ;
  assign y27991 = ~1'b0 ;
  assign y27992 = ~n47188 ;
  assign y27993 = n23185 ;
  assign y27994 = n47192 ;
  assign y27995 = n47194 ;
  assign y27996 = n47195 ;
  assign y27997 = ~1'b0 ;
  assign y27998 = n47198 ;
  assign y27999 = n47200 ;
  assign y28000 = ~n47201 ;
  assign y28001 = ~n47203 ;
  assign y28002 = 1'b0 ;
  assign y28003 = n47204 ;
  assign y28004 = ~1'b0 ;
  assign y28005 = ~1'b0 ;
  assign y28006 = ~1'b0 ;
  assign y28007 = ~n5381 ;
  assign y28008 = n47205 ;
  assign y28009 = n21429 ;
  assign y28010 = ~n47209 ;
  assign y28011 = n47214 ;
  assign y28012 = n15819 ;
  assign y28013 = ~n47218 ;
  assign y28014 = n47219 ;
  assign y28015 = n47221 ;
  assign y28016 = ~n47223 ;
  assign y28017 = n47225 ;
  assign y28018 = ~1'b0 ;
  assign y28019 = n47230 ;
  assign y28020 = ~n47238 ;
  assign y28021 = ~n47241 ;
  assign y28022 = n47242 ;
  assign y28023 = ~n47245 ;
  assign y28024 = ~1'b0 ;
  assign y28025 = n47249 ;
  assign y28026 = ~n47251 ;
  assign y28027 = ~1'b0 ;
  assign y28028 = ~1'b0 ;
  assign y28029 = n47252 ;
  assign y28030 = ~n33755 ;
  assign y28031 = n27738 ;
  assign y28032 = ~1'b0 ;
  assign y28033 = ~n47253 ;
  assign y28034 = ~n47254 ;
  assign y28035 = n47255 ;
  assign y28036 = ~n47258 ;
  assign y28037 = n47259 ;
  assign y28038 = ~n47260 ;
  assign y28039 = n47261 ;
  assign y28040 = n47263 ;
  assign y28041 = n47264 ;
  assign y28042 = ~1'b0 ;
  assign y28043 = ~n47266 ;
  assign y28044 = n47268 ;
  assign y28045 = ~1'b0 ;
  assign y28046 = ~n47270 ;
  assign y28047 = n47272 ;
  assign y28048 = n47273 ;
  assign y28049 = 1'b0 ;
  assign y28050 = ~1'b0 ;
  assign y28051 = ~1'b0 ;
  assign y28052 = ~1'b0 ;
  assign y28053 = n46767 ;
  assign y28054 = ~n47275 ;
  assign y28055 = ~1'b0 ;
  assign y28056 = ~n47277 ;
  assign y28057 = ~n47279 ;
  assign y28058 = ~n47280 ;
  assign y28059 = n47281 ;
  assign y28060 = ~n47283 ;
  assign y28061 = ~n47284 ;
  assign y28062 = n25044 ;
  assign y28063 = ~1'b0 ;
  assign y28064 = ~n47285 ;
  assign y28065 = n47286 ;
  assign y28066 = ~1'b0 ;
  assign y28067 = ~n47287 ;
  assign y28068 = n47289 ;
  assign y28069 = ~n47290 ;
  assign y28070 = n47291 ;
  assign y28071 = ~n47294 ;
  assign y28072 = n15887 ;
  assign y28073 = ~1'b0 ;
  assign y28074 = n47295 ;
  assign y28075 = 1'b0 ;
  assign y28076 = ~n47299 ;
  assign y28077 = ~1'b0 ;
  assign y28078 = ~n47301 ;
  assign y28079 = ~n6054 ;
  assign y28080 = ~1'b0 ;
  assign y28081 = ~1'b0 ;
  assign y28082 = ~n47302 ;
  assign y28083 = ~n10381 ;
  assign y28084 = ~n47304 ;
  assign y28085 = ~n47305 ;
  assign y28086 = ~n47307 ;
  assign y28087 = 1'b0 ;
  assign y28088 = ~n47309 ;
  assign y28089 = ~n47311 ;
  assign y28090 = n47312 ;
  assign y28091 = ~n47318 ;
  assign y28092 = ~n47321 ;
  assign y28093 = ~1'b0 ;
  assign y28094 = ~n47327 ;
  assign y28095 = ~n47331 ;
  assign y28096 = ~1'b0 ;
  assign y28097 = ~n47332 ;
  assign y28098 = ~n47333 ;
  assign y28099 = n47334 ;
  assign y28100 = n47335 ;
  assign y28101 = n47336 ;
  assign y28102 = n47338 ;
  assign y28103 = n47339 ;
  assign y28104 = n34615 ;
  assign y28105 = ~n47342 ;
  assign y28106 = ~n47344 ;
  assign y28107 = ~n47348 ;
  assign y28108 = ~1'b0 ;
  assign y28109 = ~1'b0 ;
  assign y28110 = ~n47351 ;
  assign y28111 = ~1'b0 ;
  assign y28112 = ~n47354 ;
  assign y28113 = ~n47356 ;
  assign y28114 = n47359 ;
  assign y28115 = n47363 ;
  assign y28116 = ~1'b0 ;
  assign y28117 = n47366 ;
  assign y28118 = ~1'b0 ;
  assign y28119 = ~n13677 ;
  assign y28120 = n5111 ;
  assign y28121 = n47368 ;
  assign y28122 = ~1'b0 ;
  assign y28123 = ~1'b0 ;
  assign y28124 = n47375 ;
  assign y28125 = 1'b0 ;
  assign y28126 = n47377 ;
  assign y28127 = 1'b0 ;
  assign y28128 = ~1'b0 ;
  assign y28129 = ~n37162 ;
  assign y28130 = ~n47381 ;
  assign y28131 = ~n47385 ;
  assign y28132 = 1'b0 ;
  assign y28133 = ~n47387 ;
  assign y28134 = ~n47393 ;
  assign y28135 = ~n47394 ;
  assign y28136 = 1'b0 ;
  assign y28137 = ~1'b0 ;
  assign y28138 = n47396 ;
  assign y28139 = ~1'b0 ;
  assign y28140 = ~n47397 ;
  assign y28141 = n47401 ;
  assign y28142 = n47403 ;
  assign y28143 = ~n47407 ;
  assign y28144 = ~n47409 ;
  assign y28145 = n47411 ;
  assign y28146 = ~n47412 ;
  assign y28147 = ~n47418 ;
  assign y28148 = ~1'b0 ;
  assign y28149 = ~n47420 ;
  assign y28150 = ~n47431 ;
  assign y28151 = ~n47432 ;
  assign y28152 = n47433 ;
  assign y28153 = 1'b0 ;
  assign y28154 = ~1'b0 ;
  assign y28155 = ~1'b0 ;
  assign y28156 = n47436 ;
  assign y28157 = n47437 ;
  assign y28158 = n47438 ;
  assign y28159 = ~n47439 ;
  assign y28160 = n47441 ;
  assign y28161 = n47457 ;
  assign y28162 = n47460 ;
  assign y28163 = ~n47463 ;
  assign y28164 = n47467 ;
  assign y28165 = ~n25719 ;
  assign y28166 = ~1'b0 ;
  assign y28167 = n47468 ;
  assign y28168 = n47475 ;
  assign y28169 = ~1'b0 ;
  assign y28170 = ~n47476 ;
  assign y28171 = ~1'b0 ;
  assign y28172 = ~n47479 ;
  assign y28173 = ~n47481 ;
  assign y28174 = ~1'b0 ;
  assign y28175 = n47484 ;
  assign y28176 = ~n9108 ;
  assign y28177 = n47485 ;
  assign y28178 = n47489 ;
  assign y28179 = 1'b0 ;
  assign y28180 = 1'b0 ;
  assign y28181 = ~n47490 ;
  assign y28182 = ~n47493 ;
  assign y28183 = n47495 ;
  assign y28184 = n47497 ;
  assign y28185 = n47499 ;
  assign y28186 = n26457 ;
  assign y28187 = n47500 ;
  assign y28188 = ~n47502 ;
  assign y28189 = ~1'b0 ;
  assign y28190 = ~n47504 ;
  assign y28191 = n47506 ;
  assign y28192 = n47507 ;
  assign y28193 = ~n47511 ;
  assign y28194 = n47513 ;
  assign y28195 = ~n47515 ;
  assign y28196 = n47517 ;
  assign y28197 = 1'b0 ;
  assign y28198 = ~n47525 ;
  assign y28199 = ~n47526 ;
  assign y28200 = ~n47528 ;
  assign y28201 = n47532 ;
  assign y28202 = n47533 ;
  assign y28203 = ~n47534 ;
  assign y28204 = ~1'b0 ;
  assign y28205 = ~1'b0 ;
  assign y28206 = ~1'b0 ;
  assign y28207 = ~1'b0 ;
  assign y28208 = n47536 ;
  assign y28209 = ~n47537 ;
  assign y28210 = ~n47538 ;
  assign y28211 = n47540 ;
  assign y28212 = ~n47542 ;
  assign y28213 = ~n47543 ;
  assign y28214 = ~1'b0 ;
  assign y28215 = ~1'b0 ;
  assign y28216 = n47544 ;
  assign y28217 = ~1'b0 ;
  assign y28218 = 1'b0 ;
  assign y28219 = ~1'b0 ;
  assign y28220 = n47545 ;
  assign y28221 = n47549 ;
  assign y28222 = ~1'b0 ;
  assign y28223 = ~1'b0 ;
  assign y28224 = n47553 ;
  assign y28225 = ~1'b0 ;
  assign y28226 = n47554 ;
  assign y28227 = n47561 ;
  assign y28228 = n47564 ;
  assign y28229 = n47570 ;
  assign y28230 = n47571 ;
  assign y28231 = ~n47576 ;
  assign y28232 = ~n47578 ;
  assign y28233 = ~n47583 ;
  assign y28234 = ~1'b0 ;
  assign y28235 = ~1'b0 ;
  assign y28236 = ~1'b0 ;
  assign y28237 = n47588 ;
  assign y28238 = ~1'b0 ;
  assign y28239 = ~1'b0 ;
  assign y28240 = n17674 ;
  assign y28241 = n47592 ;
  assign y28242 = n47593 ;
  assign y28243 = ~n47599 ;
  assign y28244 = ~n47601 ;
  assign y28245 = ~n47602 ;
  assign y28246 = ~n47603 ;
  assign y28247 = 1'b0 ;
  assign y28248 = ~1'b0 ;
  assign y28249 = n47604 ;
  assign y28250 = n47607 ;
  assign y28251 = n47608 ;
  assign y28252 = ~n47610 ;
  assign y28253 = ~1'b0 ;
  assign y28254 = ~1'b0 ;
  assign y28255 = 1'b0 ;
  assign y28256 = n47612 ;
  assign y28257 = ~1'b0 ;
  assign y28258 = n47614 ;
  assign y28259 = n22284 ;
  assign y28260 = ~1'b0 ;
  assign y28261 = ~1'b0 ;
  assign y28262 = ~n47618 ;
  assign y28263 = ~n35585 ;
  assign y28264 = ~n47619 ;
  assign y28265 = n47624 ;
  assign y28266 = ~n47625 ;
  assign y28267 = n47627 ;
  assign y28268 = ~1'b0 ;
  assign y28269 = n47630 ;
  assign y28270 = ~1'b0 ;
  assign y28271 = ~1'b0 ;
  assign y28272 = ~n47632 ;
  assign y28273 = ~1'b0 ;
  assign y28274 = n47639 ;
  assign y28275 = 1'b0 ;
  assign y28276 = ~1'b0 ;
  assign y28277 = n47640 ;
  assign y28278 = ~1'b0 ;
  assign y28279 = ~1'b0 ;
  assign y28280 = ~n47642 ;
  assign y28281 = n47643 ;
  assign y28282 = ~1'b0 ;
  assign y28283 = n46702 ;
  assign y28284 = ~1'b0 ;
  assign y28285 = ~1'b0 ;
  assign y28286 = ~n47646 ;
  assign y28287 = ~1'b0 ;
  assign y28288 = n6024 ;
  assign y28289 = ~1'b0 ;
  assign y28290 = ~n47647 ;
  assign y28291 = n47648 ;
  assign y28292 = ~n47651 ;
  assign y28293 = ~n47652 ;
  assign y28294 = ~1'b0 ;
  assign y28295 = n47655 ;
  assign y28296 = ~1'b0 ;
  assign y28297 = n47657 ;
  assign y28298 = ~1'b0 ;
  assign y28299 = ~1'b0 ;
  assign y28300 = n47661 ;
  assign y28301 = ~n47662 ;
  assign y28302 = ~n47667 ;
  assign y28303 = ~1'b0 ;
  assign y28304 = ~1'b0 ;
  assign y28305 = ~1'b0 ;
  assign y28306 = ~1'b0 ;
  assign y28307 = ~n47669 ;
  assign y28308 = ~1'b0 ;
  assign y28309 = n47672 ;
  assign y28310 = ~1'b0 ;
  assign y28311 = n4772 ;
  assign y28312 = ~n47675 ;
  assign y28313 = n47676 ;
  assign y28314 = ~n47679 ;
  assign y28315 = n47682 ;
  assign y28316 = n47683 ;
  assign y28317 = n47685 ;
  assign y28318 = n47686 ;
  assign y28319 = ~n47690 ;
  assign y28320 = n47691 ;
  assign y28321 = n47696 ;
  assign y28322 = n47699 ;
  assign y28323 = ~n47701 ;
  assign y28324 = ~1'b0 ;
  assign y28325 = ~n47705 ;
  assign y28326 = ~n493 ;
  assign y28327 = ~n47707 ;
  assign y28328 = ~n2492 ;
  assign y28329 = 1'b0 ;
  assign y28330 = ~1'b0 ;
  assign y28331 = ~n47708 ;
  assign y28332 = ~n47710 ;
  assign y28333 = n9453 ;
  assign y28334 = ~n47711 ;
  assign y28335 = n47712 ;
  assign y28336 = ~n47714 ;
  assign y28337 = n6833 ;
  assign y28338 = ~n47716 ;
  assign y28339 = ~n23882 ;
  assign y28340 = n47717 ;
  assign y28341 = ~n47719 ;
  assign y28342 = ~1'b0 ;
  assign y28343 = n47724 ;
  assign y28344 = ~n47725 ;
  assign y28345 = ~1'b0 ;
  assign y28346 = ~n47726 ;
  assign y28347 = n7174 ;
  assign y28348 = ~n47727 ;
  assign y28349 = ~n47733 ;
  assign y28350 = n47735 ;
  assign y28351 = ~1'b0 ;
  assign y28352 = n47736 ;
  assign y28353 = ~n47739 ;
  assign y28354 = n47742 ;
  assign y28355 = ~1'b0 ;
  assign y28356 = ~n47743 ;
  assign y28357 = ~n47745 ;
  assign y28358 = ~1'b0 ;
  assign y28359 = n47747 ;
  assign y28360 = ~n47748 ;
  assign y28361 = ~n47750 ;
  assign y28362 = ~n47752 ;
  assign y28363 = n47754 ;
  assign y28364 = ~n47756 ;
  assign y28365 = ~n47757 ;
  assign y28366 = ~1'b0 ;
  assign y28367 = n47759 ;
  assign y28368 = 1'b0 ;
  assign y28369 = ~n47763 ;
  assign y28370 = n47764 ;
  assign y28371 = ~n47765 ;
  assign y28372 = n47767 ;
  assign y28373 = n47769 ;
  assign y28374 = ~1'b0 ;
  assign y28375 = ~n47770 ;
  assign y28376 = n27100 ;
  assign y28377 = 1'b0 ;
  assign y28378 = ~n47776 ;
  assign y28379 = ~1'b0 ;
  assign y28380 = ~1'b0 ;
  assign y28381 = n47777 ;
  assign y28382 = ~1'b0 ;
  assign y28383 = ~1'b0 ;
  assign y28384 = n47779 ;
  assign y28385 = ~n47781 ;
  assign y28386 = ~n47782 ;
  assign y28387 = ~1'b0 ;
  assign y28388 = n8867 ;
  assign y28389 = ~n15157 ;
  assign y28390 = ~n47784 ;
  assign y28391 = ~n47788 ;
  assign y28392 = ~n47791 ;
  assign y28393 = n47800 ;
  assign y28394 = ~1'b0 ;
  assign y28395 = n47801 ;
  assign y28396 = n47803 ;
  assign y28397 = n47808 ;
  assign y28398 = ~n13293 ;
  assign y28399 = ~n47810 ;
  assign y28400 = ~1'b0 ;
  assign y28401 = ~n47814 ;
  assign y28402 = ~1'b0 ;
  assign y28403 = n47816 ;
  assign y28404 = ~n47817 ;
  assign y28405 = ~n47822 ;
  assign y28406 = ~1'b0 ;
  assign y28407 = ~n47827 ;
  assign y28408 = n47829 ;
  assign y28409 = ~1'b0 ;
  assign y28410 = ~n47830 ;
  assign y28411 = ~1'b0 ;
  assign y28412 = ~1'b0 ;
  assign y28413 = ~n47833 ;
  assign y28414 = ~1'b0 ;
  assign y28415 = n47834 ;
  assign y28416 = n47837 ;
  assign y28417 = ~n47838 ;
  assign y28418 = n47840 ;
  assign y28419 = ~n47842 ;
  assign y28420 = ~n47843 ;
  assign y28421 = ~1'b0 ;
  assign y28422 = n47844 ;
  assign y28423 = n47845 ;
  assign y28424 = ~n47847 ;
  assign y28425 = n47848 ;
  assign y28426 = 1'b0 ;
  assign y28427 = n47850 ;
  assign y28428 = ~n47853 ;
  assign y28429 = ~1'b0 ;
  assign y28430 = n47854 ;
  assign y28431 = n10160 ;
  assign y28432 = n47856 ;
  assign y28433 = ~n47858 ;
  assign y28434 = n47862 ;
  assign y28435 = n47863 ;
  assign y28436 = ~n47865 ;
  assign y28437 = ~1'b0 ;
  assign y28438 = n18960 ;
  assign y28439 = ~n47866 ;
  assign y28440 = ~1'b0 ;
  assign y28441 = ~1'b0 ;
  assign y28442 = n47868 ;
  assign y28443 = ~1'b0 ;
  assign y28444 = ~n47870 ;
  assign y28445 = ~1'b0 ;
  assign y28446 = ~n47875 ;
  assign y28447 = n47876 ;
  assign y28448 = ~1'b0 ;
  assign y28449 = ~n47884 ;
  assign y28450 = ~n34828 ;
  assign y28451 = ~n47886 ;
  assign y28452 = n13460 ;
  assign y28453 = n47887 ;
  assign y28454 = ~n47892 ;
  assign y28455 = ~n47894 ;
  assign y28456 = n14484 ;
  assign y28457 = n47895 ;
  assign y28458 = ~n47896 ;
  assign y28459 = ~1'b0 ;
  assign y28460 = 1'b0 ;
  assign y28461 = ~1'b0 ;
  assign y28462 = n47903 ;
  assign y28463 = n5150 ;
  assign y28464 = n7842 ;
  assign y28465 = ~n47904 ;
  assign y28466 = 1'b0 ;
  assign y28467 = ~1'b0 ;
  assign y28468 = n22263 ;
  assign y28469 = ~n47905 ;
  assign y28470 = ~n47907 ;
  assign y28471 = ~n47908 ;
  assign y28472 = n47910 ;
  assign y28473 = ~n47911 ;
  assign y28474 = ~n47913 ;
  assign y28475 = n47916 ;
  assign y28476 = n47917 ;
  assign y28477 = ~1'b0 ;
  assign y28478 = ~1'b0 ;
  assign y28479 = n47921 ;
  assign y28480 = n47922 ;
  assign y28481 = ~n47925 ;
  assign y28482 = ~1'b0 ;
  assign y28483 = ~n47927 ;
  assign y28484 = n47932 ;
  assign y28485 = ~1'b0 ;
  assign y28486 = ~1'b0 ;
  assign y28487 = ~n47933 ;
  assign y28488 = ~1'b0 ;
  assign y28489 = ~n47934 ;
  assign y28490 = ~n47937 ;
  assign y28491 = ~n47939 ;
  assign y28492 = ~n20812 ;
  assign y28493 = ~1'b0 ;
  assign y28494 = n47942 ;
  assign y28495 = ~n47943 ;
  assign y28496 = ~n47946 ;
  assign y28497 = ~n47949 ;
  assign y28498 = ~n47950 ;
  assign y28499 = ~1'b0 ;
  assign y28500 = n47951 ;
  assign y28501 = ~1'b0 ;
  assign y28502 = ~n47952 ;
  assign y28503 = ~n47953 ;
  assign y28504 = n20945 ;
  assign y28505 = ~n47956 ;
  assign y28506 = n47957 ;
  assign y28507 = n47959 ;
  assign y28508 = ~n47961 ;
  assign y28509 = n28301 ;
  assign y28510 = n47963 ;
  assign y28511 = n11367 ;
  assign y28512 = n47965 ;
  assign y28513 = ~1'b0 ;
  assign y28514 = ~n10499 ;
  assign y28515 = ~n47967 ;
  assign y28516 = n5240 ;
  assign y28517 = n47968 ;
  assign y28518 = ~1'b0 ;
  assign y28519 = n47973 ;
  assign y28520 = n47981 ;
  assign y28521 = ~n47984 ;
  assign y28522 = n47989 ;
  assign y28523 = n47993 ;
  assign y28524 = ~n47994 ;
  assign y28525 = ~n47995 ;
  assign y28526 = ~1'b0 ;
  assign y28527 = ~1'b0 ;
  assign y28528 = ~n47997 ;
  assign y28529 = n48000 ;
  assign y28530 = ~1'b0 ;
  assign y28531 = ~n48001 ;
  assign y28532 = ~n48004 ;
  assign y28533 = ~n48005 ;
  assign y28534 = n48008 ;
  assign y28535 = ~1'b0 ;
  assign y28536 = n48011 ;
  assign y28537 = ~n48015 ;
  assign y28538 = ~n8886 ;
  assign y28539 = ~n48020 ;
  assign y28540 = ~1'b0 ;
  assign y28541 = ~1'b0 ;
  assign y28542 = n48022 ;
  assign y28543 = ~1'b0 ;
  assign y28544 = n48025 ;
  assign y28545 = ~1'b0 ;
  assign y28546 = ~n10749 ;
  assign y28547 = ~n48031 ;
  assign y28548 = ~1'b0 ;
  assign y28549 = n48033 ;
  assign y28550 = ~n48036 ;
  assign y28551 = n48039 ;
  assign y28552 = n48040 ;
  assign y28553 = n48047 ;
  assign y28554 = ~1'b0 ;
  assign y28555 = n48049 ;
  assign y28556 = n48052 ;
  assign y28557 = ~1'b0 ;
  assign y28558 = ~1'b0 ;
  assign y28559 = n9224 ;
  assign y28560 = ~n48054 ;
  assign y28561 = ~1'b0 ;
  assign y28562 = n48055 ;
  assign y28563 = n48056 ;
  assign y28564 = n48057 ;
  assign y28565 = ~1'b0 ;
  assign y28566 = n48060 ;
  assign y28567 = ~n48061 ;
  assign y28568 = ~n48062 ;
  assign y28569 = ~n48065 ;
  assign y28570 = ~n48069 ;
  assign y28571 = ~1'b0 ;
  assign y28572 = n22242 ;
  assign y28573 = 1'b0 ;
  assign y28574 = n48070 ;
  assign y28575 = n48073 ;
  assign y28576 = 1'b0 ;
  assign y28577 = ~n48077 ;
  assign y28578 = n48078 ;
  assign y28579 = ~1'b0 ;
  assign y28580 = n6468 ;
  assign y28581 = ~1'b0 ;
  assign y28582 = ~n48080 ;
  assign y28583 = ~n14885 ;
  assign y28584 = ~n48082 ;
  assign y28585 = ~n48102 ;
  assign y28586 = ~1'b0 ;
  assign y28587 = n48103 ;
  assign y28588 = ~1'b0 ;
  assign y28589 = ~1'b0 ;
  assign y28590 = ~1'b0 ;
  assign y28591 = ~1'b0 ;
  assign y28592 = n48105 ;
  assign y28593 = ~1'b0 ;
  assign y28594 = ~n48106 ;
  assign y28595 = n48110 ;
  assign y28596 = ~1'b0 ;
  assign y28597 = n48111 ;
  assign y28598 = ~n48115 ;
  assign y28599 = 1'b0 ;
  assign y28600 = n3252 ;
  assign y28601 = ~1'b0 ;
  assign y28602 = ~1'b0 ;
  assign y28603 = n48117 ;
  assign y28604 = ~n48121 ;
  assign y28605 = n48122 ;
  assign y28606 = ~1'b0 ;
  assign y28607 = ~1'b0 ;
  assign y28608 = 1'b0 ;
  assign y28609 = ~n48124 ;
  assign y28610 = n43637 ;
  assign y28611 = ~1'b0 ;
  assign y28612 = n48127 ;
  assign y28613 = ~1'b0 ;
  assign y28614 = ~n48128 ;
  assign y28615 = n48131 ;
  assign y28616 = ~1'b0 ;
  assign y28617 = ~1'b0 ;
  assign y28618 = ~n48133 ;
  assign y28619 = ~n14849 ;
  assign y28620 = ~1'b0 ;
  assign y28621 = ~1'b0 ;
  assign y28622 = n48142 ;
  assign y28623 = ~1'b0 ;
  assign y28624 = n48145 ;
  assign y28625 = ~1'b0 ;
  assign y28626 = ~n48147 ;
  assign y28627 = n48152 ;
  assign y28628 = n48157 ;
  assign y28629 = ~n48158 ;
  assign y28630 = ~1'b0 ;
  assign y28631 = 1'b0 ;
  assign y28632 = ~n48160 ;
  assign y28633 = ~1'b0 ;
  assign y28634 = n48162 ;
  assign y28635 = 1'b0 ;
  assign y28636 = ~n48163 ;
  assign y28637 = ~n48166 ;
  assign y28638 = ~n48169 ;
  assign y28639 = ~1'b0 ;
  assign y28640 = ~1'b0 ;
  assign y28641 = ~1'b0 ;
  assign y28642 = 1'b0 ;
  assign y28643 = n10897 ;
  assign y28644 = n48170 ;
  assign y28645 = n48173 ;
  assign y28646 = n48174 ;
  assign y28647 = ~n48175 ;
  assign y28648 = ~n48176 ;
  assign y28649 = n48177 ;
  assign y28650 = ~1'b0 ;
  assign y28651 = ~1'b0 ;
  assign y28652 = ~n48178 ;
  assign y28653 = n48179 ;
  assign y28654 = ~1'b0 ;
  assign y28655 = ~n48181 ;
  assign y28656 = n48182 ;
  assign y28657 = ~n48183 ;
  assign y28658 = ~n48185 ;
  assign y28659 = ~1'b0 ;
  assign y28660 = ~1'b0 ;
  assign y28661 = ~n12403 ;
  assign y28662 = n48190 ;
  assign y28663 = ~1'b0 ;
  assign y28664 = ~1'b0 ;
  assign y28665 = 1'b0 ;
  assign y28666 = ~1'b0 ;
  assign y28667 = ~n48191 ;
  assign y28668 = n48192 ;
  assign y28669 = n48195 ;
  assign y28670 = n48196 ;
  assign y28671 = ~1'b0 ;
  assign y28672 = n48199 ;
  assign y28673 = ~n48202 ;
  assign y28674 = ~1'b0 ;
  assign y28675 = n48207 ;
  assign y28676 = n48208 ;
  assign y28677 = n48209 ;
  assign y28678 = n48210 ;
  assign y28679 = ~1'b0 ;
  assign y28680 = ~n48212 ;
  assign y28681 = 1'b0 ;
  assign y28682 = n48214 ;
  assign y28683 = 1'b0 ;
  assign y28684 = n48215 ;
  assign y28685 = ~n48221 ;
  assign y28686 = ~n48225 ;
  assign y28687 = 1'b0 ;
  assign y28688 = ~n48230 ;
  assign y28689 = ~1'b0 ;
  assign y28690 = ~1'b0 ;
  assign y28691 = 1'b0 ;
  assign y28692 = ~n48231 ;
  assign y28693 = n30102 ;
  assign y28694 = n7933 ;
  assign y28695 = ~n48232 ;
  assign y28696 = ~1'b0 ;
  assign y28697 = 1'b0 ;
  assign y28698 = ~n48237 ;
  assign y28699 = n48238 ;
  assign y28700 = ~1'b0 ;
  assign y28701 = ~1'b0 ;
  assign y28702 = ~n48243 ;
  assign y28703 = n14885 ;
  assign y28704 = ~n48244 ;
  assign y28705 = ~1'b0 ;
  assign y28706 = n48247 ;
  assign y28707 = ~n48248 ;
  assign y28708 = ~1'b0 ;
  assign y28709 = ~n48251 ;
  assign y28710 = 1'b0 ;
  assign y28711 = ~1'b0 ;
  assign y28712 = ~n48253 ;
  assign y28713 = 1'b0 ;
  assign y28714 = ~1'b0 ;
  assign y28715 = ~1'b0 ;
  assign y28716 = ~n48256 ;
  assign y28717 = n48260 ;
  assign y28718 = n48261 ;
  assign y28719 = ~n48263 ;
  assign y28720 = ~n4088 ;
  assign y28721 = ~n48266 ;
  assign y28722 = ~1'b0 ;
  assign y28723 = ~n48267 ;
  assign y28724 = ~n48269 ;
  assign y28725 = n48271 ;
  assign y28726 = ~1'b0 ;
  assign y28727 = ~1'b0 ;
  assign y28728 = ~1'b0 ;
  assign y28729 = 1'b0 ;
  assign y28730 = n27758 ;
  assign y28731 = ~n13100 ;
  assign y28732 = n48272 ;
  assign y28733 = ~n48274 ;
  assign y28734 = ~n48276 ;
  assign y28735 = n33966 ;
  assign y28736 = ~1'b0 ;
  assign y28737 = ~1'b0 ;
  assign y28738 = ~n2728 ;
  assign y28739 = ~1'b0 ;
  assign y28740 = ~n48282 ;
  assign y28741 = ~n48283 ;
  assign y28742 = n48284 ;
  assign y28743 = ~n48289 ;
  assign y28744 = n48290 ;
  assign y28745 = ~1'b0 ;
  assign y28746 = ~1'b0 ;
  assign y28747 = ~1'b0 ;
  assign y28748 = n48292 ;
  assign y28749 = ~1'b0 ;
  assign y28750 = ~n48294 ;
  assign y28751 = ~n48297 ;
  assign y28752 = ~n3064 ;
  assign y28753 = ~n48298 ;
  assign y28754 = ~1'b0 ;
  assign y28755 = ~n48299 ;
  assign y28756 = ~n48303 ;
  assign y28757 = n48305 ;
  assign y28758 = ~n48306 ;
  assign y28759 = ~1'b0 ;
  assign y28760 = ~n48308 ;
  assign y28761 = n48311 ;
  assign y28762 = ~n48313 ;
  assign y28763 = ~1'b0 ;
  assign y28764 = ~n48314 ;
  assign y28765 = n48317 ;
  assign y28766 = n48323 ;
  assign y28767 = ~n48326 ;
  assign y28768 = n19175 ;
  assign y28769 = n48327 ;
  assign y28770 = n48328 ;
  assign y28771 = ~n48330 ;
  assign y28772 = ~n48333 ;
  assign y28773 = ~n48334 ;
  assign y28774 = n48337 ;
  assign y28775 = ~1'b0 ;
  assign y28776 = n48340 ;
  assign y28777 = ~1'b0 ;
  assign y28778 = ~1'b0 ;
  assign y28779 = ~1'b0 ;
  assign y28780 = ~n48341 ;
  assign y28781 = ~n48342 ;
  assign y28782 = ~1'b0 ;
  assign y28783 = n48343 ;
  assign y28784 = ~n48347 ;
  assign y28785 = n2486 ;
  assign y28786 = n48349 ;
  assign y28787 = ~n48351 ;
  assign y28788 = ~n48352 ;
  assign y28789 = n48354 ;
  assign y28790 = ~n48360 ;
  assign y28791 = ~n48362 ;
  assign y28792 = n7997 ;
  assign y28793 = ~n48365 ;
  assign y28794 = n28346 ;
  assign y28795 = ~1'b0 ;
  assign y28796 = n48366 ;
  assign y28797 = ~1'b0 ;
  assign y28798 = n48368 ;
  assign y28799 = ~1'b0 ;
  assign y28800 = ~1'b0 ;
  assign y28801 = n48369 ;
  assign y28802 = ~1'b0 ;
  assign y28803 = n48370 ;
  assign y28804 = n48371 ;
  assign y28805 = ~n48373 ;
  assign y28806 = ~n48374 ;
  assign y28807 = n48376 ;
  assign y28808 = ~n48382 ;
  assign y28809 = ~n48387 ;
  assign y28810 = ~1'b0 ;
  assign y28811 = n48389 ;
  assign y28812 = n48393 ;
  assign y28813 = n48395 ;
  assign y28814 = ~1'b0 ;
  assign y28815 = n48397 ;
  assign y28816 = ~n5168 ;
  assign y28817 = ~1'b0 ;
  assign y28818 = ~n1157 ;
  assign y28819 = n48398 ;
  assign y28820 = ~1'b0 ;
  assign y28821 = ~1'b0 ;
  assign y28822 = n48399 ;
  assign y28823 = n48401 ;
  assign y28824 = n48402 ;
  assign y28825 = n48404 ;
  assign y28826 = 1'b0 ;
  assign y28827 = ~1'b0 ;
  assign y28828 = ~1'b0 ;
  assign y28829 = ~n48407 ;
  assign y28830 = 1'b0 ;
  assign y28831 = n48411 ;
  assign y28832 = n22720 ;
  assign y28833 = n48412 ;
  assign y28834 = ~n5727 ;
  assign y28835 = ~n48413 ;
  assign y28836 = 1'b0 ;
  assign y28837 = ~1'b0 ;
  assign y28838 = ~n23352 ;
  assign y28839 = ~1'b0 ;
  assign y28840 = ~1'b0 ;
  assign y28841 = ~n48415 ;
  assign y28842 = ~n48417 ;
  assign y28843 = ~n48418 ;
  assign y28844 = ~n48419 ;
  assign y28845 = ~n48425 ;
  assign y28846 = ~1'b0 ;
  assign y28847 = ~1'b0 ;
  assign y28848 = ~n7080 ;
  assign y28849 = n48429 ;
  assign y28850 = ~n48430 ;
  assign y28851 = ~1'b0 ;
  assign y28852 = ~n48432 ;
  assign y28853 = n48433 ;
  assign y28854 = ~n48436 ;
  assign y28855 = ~n48441 ;
  assign y28856 = ~n48444 ;
  assign y28857 = n48445 ;
  assign y28858 = ~1'b0 ;
  assign y28859 = 1'b0 ;
  assign y28860 = ~n48447 ;
  assign y28861 = n48448 ;
  assign y28862 = n48449 ;
  assign y28863 = ~n48451 ;
  assign y28864 = ~n48453 ;
  assign y28865 = ~n48455 ;
  assign y28866 = n48458 ;
  assign y28867 = ~1'b0 ;
  assign y28868 = ~n48460 ;
  assign y28869 = ~n48461 ;
  assign y28870 = n48464 ;
  assign y28871 = ~1'b0 ;
  assign y28872 = n48468 ;
  assign y28873 = ~n48470 ;
  assign y28874 = ~1'b0 ;
  assign y28875 = ~n48472 ;
  assign y28876 = n48475 ;
  assign y28877 = n38372 ;
  assign y28878 = n48477 ;
  assign y28879 = ~1'b0 ;
  assign y28880 = ~1'b0 ;
  assign y28881 = ~1'b0 ;
  assign y28882 = ~n48479 ;
  assign y28883 = n48480 ;
  assign y28884 = ~n48481 ;
  assign y28885 = ~1'b0 ;
  assign y28886 = n48487 ;
  assign y28887 = ~n48489 ;
  assign y28888 = ~n48490 ;
  assign y28889 = ~1'b0 ;
  assign y28890 = ~n48492 ;
  assign y28891 = ~n48495 ;
  assign y28892 = ~1'b0 ;
  assign y28893 = ~n37846 ;
  assign y28894 = n48497 ;
  assign y28895 = n48500 ;
  assign y28896 = ~1'b0 ;
  assign y28897 = n48502 ;
  assign y28898 = ~n48504 ;
  assign y28899 = ~1'b0 ;
  assign y28900 = ~n48507 ;
  assign y28901 = ~n48511 ;
  assign y28902 = ~n48513 ;
  assign y28903 = n48514 ;
  assign y28904 = n48515 ;
  assign y28905 = n48517 ;
  assign y28906 = ~1'b0 ;
  assign y28907 = n48520 ;
  assign y28908 = n48521 ;
  assign y28909 = ~n48523 ;
  assign y28910 = n19929 ;
  assign y28911 = n48524 ;
  assign y28912 = n48527 ;
  assign y28913 = n48529 ;
  assign y28914 = n48530 ;
  assign y28915 = n48534 ;
  assign y28916 = ~1'b0 ;
  assign y28917 = ~1'b0 ;
  assign y28918 = n48537 ;
  assign y28919 = n417 ;
  assign y28920 = ~n1914 ;
  assign y28921 = ~n48540 ;
  assign y28922 = ~n48542 ;
  assign y28923 = ~n48544 ;
  assign y28924 = ~1'b0 ;
  assign y28925 = ~1'b0 ;
  assign y28926 = n48545 ;
  assign y28927 = ~1'b0 ;
  assign y28928 = n48547 ;
  assign y28929 = ~n48548 ;
  assign y28930 = ~n48549 ;
  assign y28931 = ~n48551 ;
  assign y28932 = ~n48553 ;
  assign y28933 = ~n9322 ;
  assign y28934 = ~1'b0 ;
  assign y28935 = ~n48555 ;
  assign y28936 = ~1'b0 ;
  assign y28937 = ~1'b0 ;
  assign y28938 = n24543 ;
  assign y28939 = n1969 ;
  assign y28940 = ~n48556 ;
  assign y28941 = ~1'b0 ;
  assign y28942 = 1'b0 ;
  assign y28943 = ~n48558 ;
  assign y28944 = ~n48559 ;
  assign y28945 = ~1'b0 ;
  assign y28946 = 1'b0 ;
  assign y28947 = ~n48561 ;
  assign y28948 = n1904 ;
  assign y28949 = n48562 ;
  assign y28950 = ~n48565 ;
  assign y28951 = n48569 ;
  assign y28952 = ~n48571 ;
  assign y28953 = ~1'b0 ;
  assign y28954 = ~1'b0 ;
  assign y28955 = n48572 ;
  assign y28956 = ~1'b0 ;
  assign y28957 = ~n48578 ;
  assign y28958 = ~1'b0 ;
  assign y28959 = ~n48580 ;
  assign y28960 = ~1'b0 ;
  assign y28961 = n48582 ;
  assign y28962 = n48583 ;
  assign y28963 = ~n48589 ;
  assign y28964 = ~1'b0 ;
  assign y28965 = n48591 ;
  assign y28966 = ~1'b0 ;
  assign y28967 = n48592 ;
  assign y28968 = n48593 ;
  assign y28969 = ~1'b0 ;
  assign y28970 = ~1'b0 ;
  assign y28971 = n13375 ;
  assign y28972 = ~1'b0 ;
  assign y28973 = ~n48594 ;
  assign y28974 = n25644 ;
  assign y28975 = ~n16381 ;
  assign y28976 = n48595 ;
  assign y28977 = ~1'b0 ;
  assign y28978 = n48599 ;
  assign y28979 = ~1'b0 ;
  assign y28980 = n15246 ;
  assign y28981 = ~n48602 ;
  assign y28982 = 1'b0 ;
  assign y28983 = ~n48603 ;
  assign y28984 = ~1'b0 ;
  assign y28985 = n48605 ;
  assign y28986 = n48607 ;
  assign y28987 = ~1'b0 ;
  assign y28988 = ~n48609 ;
  assign y28989 = ~1'b0 ;
  assign y28990 = ~1'b0 ;
  assign y28991 = n48612 ;
  assign y28992 = ~n32009 ;
  assign y28993 = ~1'b0 ;
  assign y28994 = n48614 ;
  assign y28995 = n21009 ;
  assign y28996 = 1'b0 ;
  assign y28997 = ~n48618 ;
  assign y28998 = ~n48620 ;
  assign y28999 = ~n48621 ;
  assign y29000 = ~n48622 ;
  assign y29001 = ~n33347 ;
  assign y29002 = ~1'b0 ;
  assign y29003 = n48625 ;
  assign y29004 = ~n48626 ;
  assign y29005 = ~1'b0 ;
  assign y29006 = ~n48629 ;
  assign y29007 = ~1'b0 ;
  assign y29008 = 1'b0 ;
  assign y29009 = ~n48630 ;
  assign y29010 = ~n48632 ;
  assign y29011 = n48633 ;
  assign y29012 = ~1'b0 ;
  assign y29013 = n48635 ;
  assign y29014 = ~n48638 ;
  assign y29015 = ~n48642 ;
  assign y29016 = n48643 ;
  assign y29017 = ~1'b0 ;
  assign y29018 = ~n48645 ;
  assign y29019 = ~n48646 ;
  assign y29020 = ~n15324 ;
  assign y29021 = n48649 ;
  assign y29022 = ~1'b0 ;
  assign y29023 = n48650 ;
  assign y29024 = ~1'b0 ;
  assign y29025 = ~n20567 ;
  assign y29026 = ~1'b0 ;
  assign y29027 = ~1'b0 ;
  assign y29028 = ~1'b0 ;
  assign y29029 = ~1'b0 ;
  assign y29030 = n48654 ;
  assign y29031 = ~n48655 ;
  assign y29032 = ~n48656 ;
  assign y29033 = ~1'b0 ;
  assign y29034 = ~1'b0 ;
  assign y29035 = ~n48657 ;
  assign y29036 = n5076 ;
  assign y29037 = ~1'b0 ;
  assign y29038 = 1'b0 ;
  assign y29039 = n48658 ;
  assign y29040 = n48661 ;
  assign y29041 = ~1'b0 ;
  assign y29042 = ~1'b0 ;
  assign y29043 = n12594 ;
  assign y29044 = ~1'b0 ;
  assign y29045 = ~1'b0 ;
  assign y29046 = ~n48664 ;
  assign y29047 = 1'b0 ;
  assign y29048 = ~n48666 ;
  assign y29049 = ~n48667 ;
  assign y29050 = n48669 ;
  assign y29051 = n48670 ;
  assign y29052 = ~n48672 ;
  assign y29053 = ~n48673 ;
  assign y29054 = n48675 ;
  assign y29055 = ~1'b0 ;
  assign y29056 = n48676 ;
  assign y29057 = n48678 ;
  assign y29058 = ~n48681 ;
  assign y29059 = ~1'b0 ;
  assign y29060 = n48682 ;
  assign y29061 = n48683 ;
  assign y29062 = ~1'b0 ;
  assign y29063 = n48684 ;
  assign y29064 = n48685 ;
  assign y29065 = n48686 ;
  assign y29066 = ~1'b0 ;
  assign y29067 = ~1'b0 ;
  assign y29068 = n48688 ;
  assign y29069 = ~n48693 ;
  assign y29070 = ~n48694 ;
  assign y29071 = ~1'b0 ;
  assign y29072 = ~1'b0 ;
  assign y29073 = ~1'b0 ;
  assign y29074 = ~1'b0 ;
  assign y29075 = ~n48695 ;
  assign y29076 = ~n48696 ;
  assign y29077 = ~1'b0 ;
  assign y29078 = n48697 ;
  assign y29079 = n48699 ;
  assign y29080 = ~n48700 ;
  assign y29081 = n48701 ;
  assign y29082 = ~1'b0 ;
  assign y29083 = ~n9692 ;
  assign y29084 = n48702 ;
  assign y29085 = ~1'b0 ;
  assign y29086 = n48703 ;
  assign y29087 = ~n31166 ;
  assign y29088 = n48704 ;
  assign y29089 = n48705 ;
  assign y29090 = ~n37275 ;
  assign y29091 = n48707 ;
  assign y29092 = n48708 ;
  assign y29093 = ~n48711 ;
  assign y29094 = ~1'b0 ;
  assign y29095 = ~n48714 ;
  assign y29096 = ~1'b0 ;
  assign y29097 = ~n3449 ;
  assign y29098 = 1'b0 ;
  assign y29099 = ~n13520 ;
  assign y29100 = n48715 ;
  assign y29101 = n48716 ;
  assign y29102 = ~1'b0 ;
  assign y29103 = ~1'b0 ;
  assign y29104 = ~1'b0 ;
  assign y29105 = ~1'b0 ;
  assign y29106 = 1'b0 ;
  assign y29107 = n48717 ;
  assign y29108 = n48719 ;
  assign y29109 = ~1'b0 ;
  assign y29110 = ~1'b0 ;
  assign y29111 = ~n48722 ;
  assign y29112 = n11515 ;
  assign y29113 = ~n48723 ;
  assign y29114 = ~1'b0 ;
  assign y29115 = ~n48729 ;
  assign y29116 = n48731 ;
  assign y29117 = ~n48734 ;
  assign y29118 = ~1'b0 ;
  assign y29119 = ~n48735 ;
  assign y29120 = ~n48736 ;
  assign y29121 = ~n48742 ;
  assign y29122 = n48743 ;
  assign y29123 = ~n48749 ;
  assign y29124 = ~1'b0 ;
  assign y29125 = ~1'b0 ;
  assign y29126 = n48753 ;
  assign y29127 = ~1'b0 ;
  assign y29128 = ~n48756 ;
  assign y29129 = ~1'b0 ;
  assign y29130 = n12450 ;
  assign y29131 = ~n1083 ;
  assign y29132 = n48758 ;
  assign y29133 = ~n48760 ;
  assign y29134 = ~1'b0 ;
  assign y29135 = ~1'b0 ;
  assign y29136 = n48766 ;
  assign y29137 = ~n48771 ;
  assign y29138 = ~n48776 ;
  assign y29139 = ~1'b0 ;
  assign y29140 = ~1'b0 ;
  assign y29141 = ~n48778 ;
  assign y29142 = ~n48780 ;
  assign y29143 = ~1'b0 ;
  assign y29144 = ~1'b0 ;
  assign y29145 = ~n48783 ;
  assign y29146 = ~n48786 ;
  assign y29147 = n48787 ;
  assign y29148 = ~1'b0 ;
  assign y29149 = n48788 ;
  assign y29150 = n48790 ;
  assign y29151 = n48793 ;
  assign y29152 = n48797 ;
  assign y29153 = n48798 ;
  assign y29154 = ~1'b0 ;
  assign y29155 = n48800 ;
  assign y29156 = ~1'b0 ;
  assign y29157 = ~1'b0 ;
  assign y29158 = ~1'b0 ;
  assign y29159 = ~n48802 ;
  assign y29160 = n48807 ;
  assign y29161 = ~n48814 ;
  assign y29162 = ~n48816 ;
  assign y29163 = n48817 ;
  assign y29164 = ~n10568 ;
  assign y29165 = n48818 ;
  assign y29166 = ~n48821 ;
  assign y29167 = n48822 ;
  assign y29168 = ~n48824 ;
  assign y29169 = n48825 ;
  assign y29170 = ~1'b0 ;
  assign y29171 = n48826 ;
  assign y29172 = ~n48828 ;
  assign y29173 = ~n48829 ;
  assign y29174 = ~n48830 ;
  assign y29175 = n48832 ;
  assign y29176 = ~1'b0 ;
  assign y29177 = n48834 ;
  assign y29178 = ~1'b0 ;
  assign y29179 = ~1'b0 ;
  assign y29180 = ~1'b0 ;
  assign y29181 = n48836 ;
  assign y29182 = ~1'b0 ;
  assign y29183 = ~n48837 ;
  assign y29184 = ~1'b0 ;
  assign y29185 = n48839 ;
  assign y29186 = n48842 ;
  assign y29187 = ~n42427 ;
  assign y29188 = ~1'b0 ;
  assign y29189 = ~n48843 ;
  assign y29190 = ~n48845 ;
  assign y29191 = n48846 ;
  assign y29192 = ~n48847 ;
  assign y29193 = ~n48849 ;
  assign y29194 = ~n48853 ;
  assign y29195 = ~n48854 ;
  assign y29196 = n48856 ;
  assign y29197 = ~1'b0 ;
  assign y29198 = ~n48858 ;
  assign y29199 = ~n48863 ;
  assign y29200 = ~n48864 ;
  assign y29201 = n48866 ;
  assign y29202 = ~n48867 ;
  assign y29203 = ~n5535 ;
  assign y29204 = ~1'b0 ;
  assign y29205 = n48869 ;
  assign y29206 = ~n48872 ;
  assign y29207 = n48874 ;
  assign y29208 = ~1'b0 ;
  assign y29209 = ~n48875 ;
  assign y29210 = ~n48881 ;
  assign y29211 = ~n48882 ;
  assign y29212 = ~1'b0 ;
  assign y29213 = ~1'b0 ;
  assign y29214 = n48883 ;
  assign y29215 = ~n48885 ;
  assign y29216 = ~1'b0 ;
  assign y29217 = ~n48887 ;
  assign y29218 = n48888 ;
  assign y29219 = n46016 ;
  assign y29220 = ~n48890 ;
  assign y29221 = ~1'b0 ;
  assign y29222 = ~n48892 ;
  assign y29223 = ~1'b0 ;
  assign y29224 = n48899 ;
  assign y29225 = ~1'b0 ;
  assign y29226 = ~1'b0 ;
  assign y29227 = ~n48900 ;
  assign y29228 = ~n48902 ;
  assign y29229 = n48903 ;
  assign y29230 = ~n48905 ;
  assign y29231 = n48911 ;
  assign y29232 = ~1'b0 ;
  assign y29233 = n48912 ;
  assign y29234 = ~1'b0 ;
  assign y29235 = ~1'b0 ;
  assign y29236 = ~1'b0 ;
  assign y29237 = ~n48914 ;
  assign y29238 = ~n48917 ;
  assign y29239 = ~n48920 ;
  assign y29240 = ~n48921 ;
  assign y29241 = ~n48924 ;
  assign y29242 = n48925 ;
  assign y29243 = ~n6099 ;
  assign y29244 = ~1'b0 ;
  assign y29245 = n48935 ;
  assign y29246 = ~1'b0 ;
  assign y29247 = n48938 ;
  assign y29248 = ~n48939 ;
  assign y29249 = n48942 ;
  assign y29250 = ~1'b0 ;
  assign y29251 = ~1'b0 ;
  assign y29252 = ~n48943 ;
  assign y29253 = ~n48944 ;
  assign y29254 = ~n48946 ;
  assign y29255 = ~n48952 ;
  assign y29256 = ~1'b0 ;
  assign y29257 = ~1'b0 ;
  assign y29258 = ~1'b0 ;
  assign y29259 = ~n48953 ;
  assign y29260 = ~1'b0 ;
  assign y29261 = ~1'b0 ;
  assign y29262 = ~n48958 ;
  assign y29263 = ~1'b0 ;
  assign y29264 = ~n48959 ;
  assign y29265 = n48962 ;
  assign y29266 = ~1'b0 ;
  assign y29267 = ~1'b0 ;
  assign y29268 = ~n48963 ;
  assign y29269 = n48968 ;
  assign y29270 = n48971 ;
  assign y29271 = ~1'b0 ;
  assign y29272 = 1'b0 ;
  assign y29273 = n48975 ;
  assign y29274 = ~1'b0 ;
  assign y29275 = n48978 ;
  assign y29276 = n48984 ;
  assign y29277 = ~1'b0 ;
  assign y29278 = ~n48986 ;
  assign y29279 = ~n48987 ;
  assign y29280 = ~n48988 ;
  assign y29281 = ~n48989 ;
  assign y29282 = ~n48993 ;
  assign y29283 = n49001 ;
  assign y29284 = ~1'b0 ;
  assign y29285 = ~1'b0 ;
  assign y29286 = ~1'b0 ;
  assign y29287 = ~1'b0 ;
  assign y29288 = ~1'b0 ;
  assign y29289 = ~n49003 ;
  assign y29290 = n49004 ;
  assign y29291 = ~n49007 ;
  assign y29292 = 1'b0 ;
  assign y29293 = ~n49013 ;
  assign y29294 = n49019 ;
  assign y29295 = ~n49022 ;
  assign y29296 = ~n49026 ;
  assign y29297 = ~1'b0 ;
  assign y29298 = ~n49028 ;
  assign y29299 = ~n49029 ;
  assign y29300 = ~n49031 ;
  assign y29301 = n49032 ;
  assign y29302 = ~1'b0 ;
  assign y29303 = n49039 ;
  assign y29304 = ~1'b0 ;
  assign y29305 = ~1'b0 ;
  assign y29306 = ~1'b0 ;
  assign y29307 = ~1'b0 ;
  assign y29308 = ~n49041 ;
  assign y29309 = ~n7922 ;
  assign y29310 = ~n49043 ;
  assign y29311 = 1'b0 ;
  assign y29312 = ~1'b0 ;
  assign y29313 = ~n49044 ;
  assign y29314 = ~n49045 ;
  assign y29315 = ~1'b0 ;
  assign y29316 = n49046 ;
  assign y29317 = ~n15036 ;
  assign y29318 = n35617 ;
  assign y29319 = 1'b0 ;
  assign y29320 = ~n49047 ;
  assign y29321 = n49049 ;
  assign y29322 = ~n49050 ;
  assign y29323 = ~n49051 ;
  assign y29324 = n49052 ;
  assign y29325 = ~1'b0 ;
  assign y29326 = ~n49054 ;
  assign y29327 = ~1'b0 ;
  assign y29328 = ~1'b0 ;
  assign y29329 = n49057 ;
  assign y29330 = ~n17744 ;
  assign y29331 = ~1'b0 ;
  assign y29332 = ~1'b0 ;
  assign y29333 = ~n49059 ;
  assign y29334 = n49060 ;
  assign y29335 = ~1'b0 ;
  assign y29336 = ~n49065 ;
  assign y29337 = n49066 ;
  assign y29338 = ~n1438 ;
  assign y29339 = n49069 ;
  assign y29340 = ~1'b0 ;
  assign y29341 = n19840 ;
  assign y29342 = ~n49070 ;
  assign y29343 = ~n49074 ;
  assign y29344 = ~n49075 ;
  assign y29345 = ~1'b0 ;
  assign y29346 = ~n49077 ;
  assign y29347 = ~1'b0 ;
  assign y29348 = n49079 ;
  assign y29349 = ~n49080 ;
  assign y29350 = ~1'b0 ;
  assign y29351 = n49081 ;
  assign y29352 = n49083 ;
  assign y29353 = ~1'b0 ;
  assign y29354 = n49084 ;
  assign y29355 = ~n49086 ;
  assign y29356 = n17189 ;
  assign y29357 = ~n49089 ;
  assign y29358 = ~1'b0 ;
  assign y29359 = n49091 ;
  assign y29360 = ~1'b0 ;
  assign y29361 = n49092 ;
  assign y29362 = n25822 ;
  assign y29363 = n49094 ;
  assign y29364 = ~1'b0 ;
  assign y29365 = ~n49095 ;
  assign y29366 = ~1'b0 ;
  assign y29367 = ~1'b0 ;
  assign y29368 = n49097 ;
  assign y29369 = n49103 ;
  assign y29370 = ~n49106 ;
  assign y29371 = n49107 ;
  assign y29372 = ~n49109 ;
  assign y29373 = n37548 ;
  assign y29374 = n49110 ;
  assign y29375 = n49113 ;
  assign y29376 = n49116 ;
  assign y29377 = n49118 ;
  assign y29378 = ~1'b0 ;
  assign y29379 = ~n49120 ;
  assign y29380 = n49126 ;
  assign y29381 = ~1'b0 ;
  assign y29382 = ~1'b0 ;
  assign y29383 = ~1'b0 ;
  assign y29384 = n49127 ;
  assign y29385 = n49131 ;
  assign y29386 = ~1'b0 ;
  assign y29387 = ~1'b0 ;
  assign y29388 = ~1'b0 ;
  assign y29389 = ~1'b0 ;
  assign y29390 = n49132 ;
  assign y29391 = ~1'b0 ;
  assign y29392 = n49134 ;
  assign y29393 = ~1'b0 ;
  assign y29394 = n49137 ;
  assign y29395 = 1'b0 ;
  assign y29396 = ~1'b0 ;
  assign y29397 = ~1'b0 ;
  assign y29398 = ~n49140 ;
  assign y29399 = ~n49141 ;
  assign y29400 = ~1'b0 ;
  assign y29401 = ~n49146 ;
  assign y29402 = ~n49148 ;
  assign y29403 = ~n49152 ;
  assign y29404 = ~1'b0 ;
  assign y29405 = ~n49154 ;
  assign y29406 = ~n23780 ;
  assign y29407 = ~1'b0 ;
  assign y29408 = ~n49161 ;
  assign y29409 = ~1'b0 ;
  assign y29410 = ~1'b0 ;
  assign y29411 = ~1'b0 ;
  assign y29412 = ~n49162 ;
  assign y29413 = ~1'b0 ;
  assign y29414 = ~1'b0 ;
  assign y29415 = ~1'b0 ;
  assign y29416 = n49163 ;
  assign y29417 = ~n49166 ;
  assign y29418 = ~1'b0 ;
  assign y29419 = ~1'b0 ;
  assign y29420 = ~n49167 ;
  assign y29421 = ~n49168 ;
  assign y29422 = ~1'b0 ;
  assign y29423 = ~1'b0 ;
  assign y29424 = ~1'b0 ;
  assign y29425 = ~1'b0 ;
  assign y29426 = ~n49169 ;
  assign y29427 = ~n49171 ;
  assign y29428 = ~1'b0 ;
  assign y29429 = n49173 ;
  assign y29430 = n49174 ;
  assign y29431 = ~n49175 ;
  assign y29432 = n49176 ;
  assign y29433 = ~n49180 ;
  assign y29434 = ~n49182 ;
  assign y29435 = ~1'b0 ;
  assign y29436 = n49184 ;
  assign y29437 = n49186 ;
  assign y29438 = ~n11524 ;
  assign y29439 = ~1'b0 ;
  assign y29440 = ~1'b0 ;
  assign y29441 = ~n49188 ;
  assign y29442 = ~1'b0 ;
  assign y29443 = ~n49190 ;
  assign y29444 = n49191 ;
  assign y29445 = n49194 ;
  assign y29446 = ~n49195 ;
  assign y29447 = n758 ;
  assign y29448 = ~n49197 ;
  assign y29449 = n29402 ;
  assign y29450 = ~n49200 ;
  assign y29451 = n49201 ;
  assign y29452 = ~n49202 ;
  assign y29453 = n49203 ;
  assign y29454 = ~n49204 ;
  assign y29455 = ~n49207 ;
  assign y29456 = ~1'b0 ;
  assign y29457 = ~n49208 ;
  assign y29458 = n49210 ;
  assign y29459 = ~1'b0 ;
  assign y29460 = n49214 ;
  assign y29461 = ~1'b0 ;
  assign y29462 = ~1'b0 ;
  assign y29463 = ~1'b0 ;
  assign y29464 = n49215 ;
  assign y29465 = ~n49218 ;
  assign y29466 = ~1'b0 ;
  assign y29467 = ~1'b0 ;
  assign y29468 = n14194 ;
  assign y29469 = n49219 ;
  assign y29470 = ~n47998 ;
  assign y29471 = ~n49220 ;
  assign y29472 = 1'b0 ;
  assign y29473 = n49221 ;
  assign y29474 = ~n49224 ;
  assign y29475 = ~1'b0 ;
  assign y29476 = n49225 ;
  assign y29477 = n46911 ;
  assign y29478 = ~1'b0 ;
  assign y29479 = ~1'b0 ;
  assign y29480 = ~n49227 ;
  assign y29481 = ~1'b0 ;
  assign y29482 = ~n49229 ;
  assign y29483 = ~1'b0 ;
  assign y29484 = ~n49230 ;
  assign y29485 = ~n49233 ;
  assign y29486 = n49236 ;
  assign y29487 = ~1'b0 ;
  assign y29488 = n49238 ;
  assign y29489 = ~1'b0 ;
  assign y29490 = n49240 ;
  assign y29491 = n49241 ;
  assign y29492 = n49243 ;
  assign y29493 = n7619 ;
  assign y29494 = ~n49244 ;
  assign y29495 = n49246 ;
  assign y29496 = n49250 ;
  assign y29497 = ~1'b0 ;
  assign y29498 = ~n49251 ;
  assign y29499 = n49252 ;
  assign y29500 = n49255 ;
  assign y29501 = n49256 ;
  assign y29502 = n49257 ;
  assign y29503 = ~1'b0 ;
  assign y29504 = ~1'b0 ;
  assign y29505 = ~1'b0 ;
  assign y29506 = ~1'b0 ;
  assign y29507 = n49258 ;
  assign y29508 = ~1'b0 ;
  assign y29509 = ~n49260 ;
  assign y29510 = ~n49267 ;
  assign y29511 = n49273 ;
  assign y29512 = ~n49276 ;
  assign y29513 = ~n49278 ;
  assign y29514 = n49280 ;
  assign y29515 = ~1'b0 ;
  assign y29516 = n49288 ;
  assign y29517 = ~1'b0 ;
  assign y29518 = n49289 ;
  assign y29519 = n49291 ;
  assign y29520 = ~n49292 ;
  assign y29521 = n49293 ;
  assign y29522 = n49296 ;
  assign y29523 = 1'b0 ;
  assign y29524 = ~1'b0 ;
  assign y29525 = ~n49298 ;
  assign y29526 = n8993 ;
  assign y29527 = ~1'b0 ;
  assign y29528 = ~1'b0 ;
  assign y29529 = ~n49300 ;
  assign y29530 = 1'b0 ;
  assign y29531 = ~1'b0 ;
  assign y29532 = ~n49301 ;
  assign y29533 = n49302 ;
  assign y29534 = ~1'b0 ;
  assign y29535 = ~1'b0 ;
  assign y29536 = ~n49305 ;
  assign y29537 = ~1'b0 ;
  assign y29538 = n49307 ;
  assign y29539 = n41330 ;
  assign y29540 = ~1'b0 ;
  assign y29541 = ~1'b0 ;
  assign y29542 = ~n49309 ;
  assign y29543 = ~n49310 ;
  assign y29544 = n49312 ;
  assign y29545 = ~1'b0 ;
  assign y29546 = ~n49314 ;
  assign y29547 = ~n49316 ;
  assign y29548 = ~1'b0 ;
  assign y29549 = n49318 ;
  assign y29550 = ~n49319 ;
  assign y29551 = n49321 ;
  assign y29552 = ~n49323 ;
  assign y29553 = n1045 ;
  assign y29554 = n49325 ;
  assign y29555 = ~n49328 ;
  assign y29556 = n49332 ;
  assign y29557 = ~1'b0 ;
  assign y29558 = ~n15777 ;
  assign y29559 = ~n49334 ;
  assign y29560 = ~1'b0 ;
  assign y29561 = ~1'b0 ;
  assign y29562 = ~n49336 ;
  assign y29563 = ~n49338 ;
  assign y29564 = n49341 ;
  assign y29565 = n49345 ;
  assign y29566 = n49347 ;
  assign y29567 = ~1'b0 ;
  assign y29568 = n49350 ;
  assign y29569 = ~1'b0 ;
  assign y29570 = ~n49351 ;
  assign y29571 = n29957 ;
  assign y29572 = ~1'b0 ;
  assign y29573 = ~1'b0 ;
  assign y29574 = n49355 ;
  assign y29575 = ~n49356 ;
  assign y29576 = ~n49360 ;
  assign y29577 = ~n49361 ;
  assign y29578 = n49362 ;
  assign y29579 = n49364 ;
  assign y29580 = n49367 ;
  assign y29581 = n49369 ;
  assign y29582 = n49370 ;
  assign y29583 = n49379 ;
  assign y29584 = ~n49381 ;
  assign y29585 = n12582 ;
  assign y29586 = ~n49383 ;
  assign y29587 = n49387 ;
  assign y29588 = ~n49394 ;
  assign y29589 = ~1'b0 ;
  assign y29590 = ~n49396 ;
  assign y29591 = ~1'b0 ;
  assign y29592 = ~n49401 ;
  assign y29593 = n49407 ;
  assign y29594 = ~n49408 ;
  assign y29595 = ~n49409 ;
  assign y29596 = ~n49412 ;
  assign y29597 = ~1'b0 ;
  assign y29598 = n49414 ;
  assign y29599 = ~n49415 ;
  assign y29600 = n49416 ;
  assign y29601 = ~1'b0 ;
  assign y29602 = ~n49417 ;
  assign y29603 = n49418 ;
  assign y29604 = n49419 ;
  assign y29605 = n49421 ;
  assign y29606 = ~n49423 ;
  assign y29607 = n49426 ;
  assign y29608 = ~1'b0 ;
  assign y29609 = ~1'b0 ;
  assign y29610 = ~n49427 ;
  assign y29611 = ~1'b0 ;
  assign y29612 = n49431 ;
  assign y29613 = n49433 ;
  assign y29614 = ~1'b0 ;
  assign y29615 = n49438 ;
  assign y29616 = ~1'b0 ;
  assign y29617 = n49443 ;
  assign y29618 = ~n49444 ;
  assign y29619 = ~n49447 ;
  assign y29620 = 1'b0 ;
  assign y29621 = ~1'b0 ;
  assign y29622 = n49450 ;
  assign y29623 = n49451 ;
  assign y29624 = n49453 ;
  assign y29625 = ~1'b0 ;
  assign y29626 = ~1'b0 ;
  assign y29627 = n49454 ;
  assign y29628 = ~n49463 ;
  assign y29629 = ~n49464 ;
  assign y29630 = ~n49465 ;
  assign y29631 = ~1'b0 ;
  assign y29632 = n17352 ;
  assign y29633 = ~1'b0 ;
  assign y29634 = n45388 ;
  assign y29635 = n49467 ;
  assign y29636 = ~1'b0 ;
  assign y29637 = ~1'b0 ;
  assign y29638 = ~n49468 ;
  assign y29639 = ~n49472 ;
  assign y29640 = n49478 ;
  assign y29641 = ~1'b0 ;
  assign y29642 = ~n49480 ;
  assign y29643 = ~1'b0 ;
  assign y29644 = ~n49482 ;
  assign y29645 = n2540 ;
  assign y29646 = ~1'b0 ;
  assign y29647 = ~n49484 ;
  assign y29648 = n49485 ;
  assign y29649 = n49489 ;
  assign y29650 = n49492 ;
  assign y29651 = ~1'b0 ;
  assign y29652 = n49494 ;
  assign y29653 = ~n49496 ;
  assign y29654 = n3378 ;
  assign y29655 = n49503 ;
  assign y29656 = ~1'b0 ;
  assign y29657 = n49505 ;
  assign y29658 = ~1'b0 ;
  assign y29659 = ~n49506 ;
  assign y29660 = ~n49507 ;
  assign y29661 = ~1'b0 ;
  assign y29662 = n49510 ;
  assign y29663 = n49513 ;
  assign y29664 = ~1'b0 ;
  assign y29665 = n43454 ;
  assign y29666 = n49515 ;
  assign y29667 = n49518 ;
  assign y29668 = ~n49521 ;
  assign y29669 = ~n49525 ;
  assign y29670 = 1'b0 ;
  assign y29671 = n49526 ;
  assign y29672 = n49532 ;
  assign y29673 = ~n49534 ;
  assign y29674 = n49535 ;
  assign y29675 = n49536 ;
  assign y29676 = ~1'b0 ;
  assign y29677 = ~1'b0 ;
  assign y29678 = ~n49538 ;
  assign y29679 = ~1'b0 ;
  assign y29680 = ~1'b0 ;
  assign y29681 = ~n49546 ;
  assign y29682 = ~n522 ;
  assign y29683 = ~1'b0 ;
  assign y29684 = ~n46162 ;
  assign y29685 = n49547 ;
  assign y29686 = ~n49551 ;
  assign y29687 = n49553 ;
  assign y29688 = ~1'b0 ;
  assign y29689 = ~n49554 ;
  assign y29690 = n49557 ;
  assign y29691 = ~n49558 ;
  assign y29692 = n49559 ;
  assign y29693 = ~n49560 ;
  assign y29694 = ~n49561 ;
  assign y29695 = ~n25429 ;
  assign y29696 = 1'b0 ;
  assign y29697 = ~n1065 ;
  assign y29698 = n49563 ;
  assign y29699 = ~n15068 ;
  assign y29700 = ~1'b0 ;
  assign y29701 = ~n49564 ;
  assign y29702 = ~1'b0 ;
  assign y29703 = ~1'b0 ;
  assign y29704 = n49565 ;
  assign y29705 = ~n49569 ;
  assign y29706 = n18731 ;
  assign y29707 = n41841 ;
  assign y29708 = ~1'b0 ;
  assign y29709 = 1'b0 ;
  assign y29710 = ~n49577 ;
  assign y29711 = ~n4357 ;
  assign y29712 = ~n49579 ;
  assign y29713 = ~n49580 ;
  assign y29714 = ~n49582 ;
  assign y29715 = ~n49584 ;
  assign y29716 = ~n49585 ;
  assign y29717 = ~1'b0 ;
  assign y29718 = ~1'b0 ;
  assign y29719 = ~n49589 ;
  assign y29720 = ~1'b0 ;
  assign y29721 = ~n49591 ;
  assign y29722 = ~1'b0 ;
  assign y29723 = ~n49594 ;
  assign y29724 = ~1'b0 ;
  assign y29725 = n49595 ;
  assign y29726 = n49599 ;
  assign y29727 = 1'b0 ;
  assign y29728 = ~n49601 ;
  assign y29729 = n49602 ;
  assign y29730 = ~1'b0 ;
  assign y29731 = ~1'b0 ;
  assign y29732 = ~n49603 ;
  assign y29733 = n49604 ;
  assign y29734 = ~1'b0 ;
  assign y29735 = n49605 ;
  assign y29736 = ~n6563 ;
  assign y29737 = n49607 ;
  assign y29738 = n23768 ;
  assign y29739 = ~1'b0 ;
  assign y29740 = ~1'b0 ;
  assign y29741 = n49613 ;
  assign y29742 = ~n49614 ;
  assign y29743 = n49615 ;
  assign y29744 = ~1'b0 ;
  assign y29745 = ~1'b0 ;
  assign y29746 = ~n49617 ;
  assign y29747 = n49626 ;
  assign y29748 = ~1'b0 ;
  assign y29749 = ~n49627 ;
  assign y29750 = ~n49632 ;
  assign y29751 = ~n49633 ;
  assign y29752 = ~n49635 ;
  assign y29753 = n49636 ;
  assign y29754 = n49638 ;
  assign y29755 = ~1'b0 ;
  assign y29756 = ~1'b0 ;
  assign y29757 = n49639 ;
  assign y29758 = 1'b0 ;
  assign y29759 = ~n49641 ;
  assign y29760 = n49642 ;
  assign y29761 = ~n49645 ;
  assign y29762 = n49647 ;
  assign y29763 = ~n49648 ;
  assign y29764 = ~n49649 ;
  assign y29765 = ~n49652 ;
  assign y29766 = n49653 ;
  assign y29767 = ~1'b0 ;
  assign y29768 = n39630 ;
  assign y29769 = n49656 ;
  assign y29770 = n49660 ;
  assign y29771 = n49662 ;
  assign y29772 = n49664 ;
  assign y29773 = ~1'b0 ;
  assign y29774 = n49665 ;
  assign y29775 = ~1'b0 ;
  assign y29776 = ~1'b0 ;
  assign y29777 = n49666 ;
  assign y29778 = ~n911 ;
  assign y29779 = ~n49668 ;
  assign y29780 = n49669 ;
  assign y29781 = ~n49671 ;
  assign y29782 = ~1'b0 ;
  assign y29783 = ~n6428 ;
  assign y29784 = ~n49672 ;
  assign y29785 = ~1'b0 ;
  assign y29786 = ~1'b0 ;
  assign y29787 = ~1'b0 ;
  assign y29788 = ~1'b0 ;
  assign y29789 = ~n49673 ;
  assign y29790 = ~n49674 ;
  assign y29791 = ~1'b0 ;
  assign y29792 = n27902 ;
  assign y29793 = n49677 ;
  assign y29794 = n49679 ;
  assign y29795 = ~n49680 ;
  assign y29796 = n49682 ;
  assign y29797 = ~n35451 ;
  assign y29798 = n38576 ;
  assign y29799 = n49683 ;
  assign y29800 = n44272 ;
  assign y29801 = n35559 ;
  assign y29802 = n49686 ;
  assign y29803 = n49687 ;
  assign y29804 = ~1'b0 ;
  assign y29805 = 1'b0 ;
  assign y29806 = n49688 ;
  assign y29807 = n49690 ;
  assign y29808 = n49692 ;
  assign y29809 = ~1'b0 ;
  assign y29810 = ~n49693 ;
  assign y29811 = n49696 ;
  assign y29812 = ~n49698 ;
  assign y29813 = n49701 ;
  assign y29814 = n49702 ;
  assign y29815 = n49706 ;
  assign y29816 = ~n49708 ;
  assign y29817 = n49709 ;
  assign y29818 = ~n49711 ;
  assign y29819 = ~1'b0 ;
  assign y29820 = ~1'b0 ;
  assign y29821 = n10826 ;
  assign y29822 = ~n36952 ;
  assign y29823 = ~n49720 ;
  assign y29824 = ~1'b0 ;
  assign y29825 = ~n3651 ;
  assign y29826 = ~n49721 ;
  assign y29827 = ~1'b0 ;
  assign y29828 = ~n49727 ;
  assign y29829 = ~n49729 ;
  assign y29830 = ~n49730 ;
  assign y29831 = n49735 ;
  assign y29832 = ~n49736 ;
  assign y29833 = n49739 ;
  assign y29834 = ~n49742 ;
  assign y29835 = 1'b0 ;
  assign y29836 = ~n49746 ;
  assign y29837 = ~1'b0 ;
  assign y29838 = ~1'b0 ;
  assign y29839 = n49747 ;
  assign y29840 = ~n49748 ;
  assign y29841 = n49750 ;
  assign y29842 = n49757 ;
  assign y29843 = ~n49758 ;
  assign y29844 = n49760 ;
  assign y29845 = ~n49763 ;
  assign y29846 = ~n49765 ;
  assign y29847 = ~1'b0 ;
  assign y29848 = ~1'b0 ;
  assign y29849 = n49767 ;
  assign y29850 = n49769 ;
  assign y29851 = ~1'b0 ;
  assign y29852 = ~1'b0 ;
  assign y29853 = ~1'b0 ;
  assign y29854 = n49772 ;
  assign y29855 = ~n17970 ;
  assign y29856 = n15856 ;
  assign y29857 = n49777 ;
  assign y29858 = ~n49779 ;
  assign y29859 = ~n49780 ;
  assign y29860 = n49783 ;
  assign y29861 = 1'b0 ;
  assign y29862 = n30313 ;
  assign y29863 = ~1'b0 ;
  assign y29864 = 1'b0 ;
  assign y29865 = ~n49784 ;
  assign y29866 = ~n49785 ;
  assign y29867 = 1'b0 ;
  assign y29868 = n49792 ;
  assign y29869 = ~1'b0 ;
  assign y29870 = ~n49793 ;
  assign y29871 = ~1'b0 ;
  assign y29872 = ~n49794 ;
  assign y29873 = ~n49796 ;
  assign y29874 = ~1'b0 ;
  assign y29875 = n49798 ;
  assign y29876 = ~n49803 ;
  assign y29877 = ~n49804 ;
  assign y29878 = ~n49806 ;
  assign y29879 = ~n49808 ;
  assign y29880 = ~1'b0 ;
  assign y29881 = ~n49810 ;
  assign y29882 = n49814 ;
  assign y29883 = ~n49816 ;
  assign y29884 = ~n49571 ;
  assign y29885 = ~1'b0 ;
  assign y29886 = ~n49818 ;
  assign y29887 = ~n49822 ;
  assign y29888 = n49823 ;
  assign y29889 = ~n49827 ;
  assign y29890 = ~n49835 ;
  assign y29891 = n49838 ;
  assign y29892 = ~1'b0 ;
  assign y29893 = n49840 ;
  assign y29894 = ~n45804 ;
  assign y29895 = ~1'b0 ;
  assign y29896 = ~1'b0 ;
  assign y29897 = ~n49843 ;
  assign y29898 = n49844 ;
  assign y29899 = ~n49846 ;
  assign y29900 = ~1'b0 ;
  assign y29901 = ~1'b0 ;
  assign y29902 = n49848 ;
  assign y29903 = ~1'b0 ;
  assign y29904 = ~1'b0 ;
  assign y29905 = ~n49849 ;
  assign y29906 = n49853 ;
  assign y29907 = n49859 ;
  assign y29908 = ~n27524 ;
  assign y29909 = ~1'b0 ;
  assign y29910 = ~1'b0 ;
  assign y29911 = n49861 ;
  assign y29912 = n49863 ;
  assign y29913 = ~n49866 ;
  assign y29914 = n7757 ;
  assign y29915 = ~1'b0 ;
  assign y29916 = ~1'b0 ;
  assign y29917 = ~1'b0 ;
  assign y29918 = n49869 ;
  assign y29919 = n49870 ;
  assign y29920 = n49871 ;
  assign y29921 = 1'b0 ;
  assign y29922 = ~1'b0 ;
  assign y29923 = ~1'b0 ;
  assign y29924 = ~1'b0 ;
  assign y29925 = ~1'b0 ;
  assign y29926 = n49872 ;
  assign y29927 = ~1'b0 ;
  assign y29928 = n49874 ;
  assign y29929 = ~n6256 ;
  assign y29930 = ~1'b0 ;
  assign y29931 = n49876 ;
  assign y29932 = ~1'b0 ;
  assign y29933 = ~1'b0 ;
  assign y29934 = ~n49877 ;
  assign y29935 = n11438 ;
  assign y29936 = ~n49878 ;
  assign y29937 = ~1'b0 ;
  assign y29938 = ~n49880 ;
  assign y29939 = n49881 ;
  assign y29940 = ~n49883 ;
  assign y29941 = ~n49884 ;
  assign y29942 = ~n49885 ;
  assign y29943 = ~n49888 ;
  assign y29944 = ~1'b0 ;
  assign y29945 = ~1'b0 ;
  assign y29946 = ~1'b0 ;
  assign y29947 = ~n49890 ;
  assign y29948 = ~n49892 ;
  assign y29949 = ~1'b0 ;
  assign y29950 = n49893 ;
  assign y29951 = n49894 ;
  assign y29952 = ~n6917 ;
  assign y29953 = ~n49904 ;
  assign y29954 = n49906 ;
  assign y29955 = ~1'b0 ;
  assign y29956 = ~1'b0 ;
  assign y29957 = ~n49908 ;
  assign y29958 = ~n49910 ;
  assign y29959 = n49911 ;
  assign y29960 = ~n49915 ;
  assign y29961 = ~1'b0 ;
  assign y29962 = n49920 ;
  assign y29963 = ~n49922 ;
  assign y29964 = ~n49926 ;
  assign y29965 = 1'b0 ;
  assign y29966 = n49928 ;
  assign y29967 = ~1'b0 ;
  assign y29968 = ~n49929 ;
  assign y29969 = ~n49934 ;
  assign y29970 = n49935 ;
  assign y29971 = n49937 ;
  assign y29972 = ~n2080 ;
  assign y29973 = ~1'b0 ;
  assign y29974 = n14388 ;
  assign y29975 = n49938 ;
  assign y29976 = n49939 ;
  assign y29977 = n49942 ;
  assign y29978 = n49944 ;
  assign y29979 = ~n49946 ;
  assign y29980 = n49954 ;
  assign y29981 = ~n49957 ;
  assign y29982 = n49959 ;
  assign y29983 = ~1'b0 ;
  assign y29984 = ~n49960 ;
  assign y29985 = n49963 ;
  assign y29986 = ~n49964 ;
  assign y29987 = ~1'b0 ;
  assign y29988 = ~1'b0 ;
  assign y29989 = ~1'b0 ;
  assign y29990 = ~n49966 ;
  assign y29991 = ~1'b0 ;
  assign y29992 = n49968 ;
  assign y29993 = n49969 ;
  assign y29994 = ~1'b0 ;
  assign y29995 = ~n49971 ;
  assign y29996 = n49972 ;
  assign y29997 = n49973 ;
  assign y29998 = ~1'b0 ;
  assign y29999 = ~1'b0 ;
  assign y30000 = n49975 ;
  assign y30001 = ~1'b0 ;
  assign y30002 = ~1'b0 ;
  assign y30003 = n49976 ;
  assign y30004 = ~1'b0 ;
  assign y30005 = ~1'b0 ;
  assign y30006 = ~n49978 ;
  assign y30007 = n49979 ;
  assign y30008 = n49982 ;
  assign y30009 = ~1'b0 ;
  assign y30010 = ~n49985 ;
  assign y30011 = 1'b0 ;
  assign y30012 = ~1'b0 ;
  assign y30013 = 1'b0 ;
  assign y30014 = n49986 ;
  assign y30015 = n27087 ;
  assign y30016 = ~n49991 ;
  assign y30017 = n49993 ;
  assign y30018 = ~1'b0 ;
  assign y30019 = n6709 ;
  assign y30020 = n49995 ;
  assign y30021 = ~n49996 ;
  assign y30022 = ~n49997 ;
  assign y30023 = ~1'b0 ;
  assign y30024 = ~1'b0 ;
  assign y30025 = ~1'b0 ;
  assign y30026 = ~n49998 ;
  assign y30027 = ~n49999 ;
  assign y30028 = n50008 ;
  assign y30029 = n31370 ;
  assign y30030 = ~1'b0 ;
  assign y30031 = ~1'b0 ;
  assign y30032 = ~1'b0 ;
  assign y30033 = ~1'b0 ;
  assign y30034 = n50010 ;
  assign y30035 = ~1'b0 ;
  assign y30036 = n50011 ;
  assign y30037 = ~1'b0 ;
  assign y30038 = ~1'b0 ;
  assign y30039 = ~n50013 ;
  assign y30040 = n50015 ;
  assign y30041 = ~1'b0 ;
  assign y30042 = n50016 ;
  assign y30043 = ~n11211 ;
  assign y30044 = ~n50017 ;
  assign y30045 = n50018 ;
  assign y30046 = ~1'b0 ;
  assign y30047 = 1'b0 ;
  assign y30048 = ~n50022 ;
  assign y30049 = ~1'b0 ;
  assign y30050 = n26095 ;
  assign y30051 = n33099 ;
  assign y30052 = n50025 ;
  assign y30053 = 1'b0 ;
  assign y30054 = n50027 ;
  assign y30055 = n20656 ;
  assign y30056 = ~n50028 ;
  assign y30057 = ~n50029 ;
  assign y30058 = ~n50032 ;
  assign y30059 = n50033 ;
  assign y30060 = n50034 ;
  assign y30061 = n50035 ;
  assign y30062 = ~n50037 ;
  assign y30063 = ~n50041 ;
  assign y30064 = ~n50043 ;
  assign y30065 = n50044 ;
  assign y30066 = n50047 ;
  assign y30067 = n50051 ;
  assign y30068 = ~n50055 ;
  assign y30069 = ~1'b0 ;
  assign y30070 = ~n50058 ;
  assign y30071 = n50059 ;
  assign y30072 = ~n8239 ;
  assign y30073 = n50063 ;
  assign y30074 = ~n50065 ;
  assign y30075 = n50067 ;
  assign y30076 = ~1'b0 ;
  assign y30077 = ~1'b0 ;
  assign y30078 = ~n50068 ;
  assign y30079 = ~1'b0 ;
  assign y30080 = ~1'b0 ;
  assign y30081 = ~1'b0 ;
  assign y30082 = n50070 ;
  assign y30083 = n50071 ;
  assign y30084 = ~n36140 ;
  assign y30085 = ~1'b0 ;
  assign y30086 = ~1'b0 ;
  assign y30087 = ~n50074 ;
  assign y30088 = ~n50078 ;
  assign y30089 = ~1'b0 ;
  assign y30090 = n14718 ;
  assign y30091 = ~n50082 ;
  assign y30092 = n50084 ;
  assign y30093 = n50091 ;
  assign y30094 = n50092 ;
  assign y30095 = ~n39288 ;
  assign y30096 = n50094 ;
  assign y30097 = ~1'b0 ;
  assign y30098 = ~1'b0 ;
  assign y30099 = ~n50095 ;
  assign y30100 = ~n50096 ;
  assign y30101 = n50098 ;
  assign y30102 = ~1'b0 ;
  assign y30103 = ~n50099 ;
  assign y30104 = ~1'b0 ;
  assign y30105 = ~n50105 ;
  assign y30106 = ~n50106 ;
  assign y30107 = n50108 ;
  assign y30108 = ~n50110 ;
  assign y30109 = ~n50115 ;
  assign y30110 = ~n50119 ;
  assign y30111 = ~n16359 ;
  assign y30112 = n50121 ;
  assign y30113 = ~1'b0 ;
  assign y30114 = ~1'b0 ;
  assign y30115 = ~1'b0 ;
  assign y30116 = ~n50122 ;
  assign y30117 = n50128 ;
  assign y30118 = ~n50129 ;
  assign y30119 = 1'b0 ;
  assign y30120 = ~n50132 ;
  assign y30121 = n50133 ;
  assign y30122 = ~n4570 ;
  assign y30123 = n51 ;
  assign y30124 = n50135 ;
  assign y30125 = n48540 ;
  assign y30126 = ~n50140 ;
  assign y30127 = ~n50142 ;
  assign y30128 = n38061 ;
  assign y30129 = ~1'b0 ;
  assign y30130 = n50148 ;
  assign y30131 = ~1'b0 ;
  assign y30132 = ~1'b0 ;
  assign y30133 = ~n50150 ;
  assign y30134 = ~1'b0 ;
  assign y30135 = ~1'b0 ;
  assign y30136 = ~1'b0 ;
  assign y30137 = n50153 ;
  assign y30138 = n50154 ;
  assign y30139 = ~1'b0 ;
  assign y30140 = ~1'b0 ;
  assign y30141 = ~n50155 ;
  assign y30142 = n50157 ;
  assign y30143 = ~n8757 ;
  assign y30144 = ~n50160 ;
  assign y30145 = ~1'b0 ;
  assign y30146 = ~1'b0 ;
  assign y30147 = n4942 ;
  assign y30148 = n50163 ;
  assign y30149 = n50166 ;
  assign y30150 = ~1'b0 ;
  assign y30151 = n50167 ;
  assign y30152 = ~n50169 ;
  assign y30153 = 1'b0 ;
  assign y30154 = ~n50173 ;
  assign y30155 = n50174 ;
  assign y30156 = ~n50176 ;
  assign y30157 = ~n50177 ;
  assign y30158 = ~1'b0 ;
  assign y30159 = ~n10003 ;
  assign y30160 = n50179 ;
  assign y30161 = n50184 ;
  assign y30162 = ~n50185 ;
  assign y30163 = ~1'b0 ;
  assign y30164 = ~1'b0 ;
  assign y30165 = ~1'b0 ;
  assign y30166 = ~1'b0 ;
  assign y30167 = ~n50186 ;
  assign y30168 = n50188 ;
  assign y30169 = ~1'b0 ;
  assign y30170 = n50190 ;
  assign y30171 = ~n50193 ;
  assign y30172 = ~n50194 ;
  assign y30173 = ~1'b0 ;
  assign y30174 = ~1'b0 ;
  assign y30175 = ~n50196 ;
  assign y30176 = ~1'b0 ;
  assign y30177 = ~1'b0 ;
  assign y30178 = ~n50198 ;
  assign y30179 = ~n50200 ;
  assign y30180 = ~n50204 ;
  assign y30181 = ~n50205 ;
  assign y30182 = n50206 ;
  assign y30183 = ~1'b0 ;
  assign y30184 = ~n50208 ;
  assign y30185 = ~n50210 ;
  assign y30186 = n50215 ;
  assign y30187 = ~n21535 ;
  assign y30188 = ~n50216 ;
  assign y30189 = ~1'b0 ;
  assign y30190 = ~n50217 ;
  assign y30191 = ~1'b0 ;
  assign y30192 = n50218 ;
  assign y30193 = n50221 ;
  assign y30194 = ~1'b0 ;
  assign y30195 = ~1'b0 ;
  assign y30196 = ~1'b0 ;
  assign y30197 = ~n50223 ;
  assign y30198 = ~1'b0 ;
  assign y30199 = n50224 ;
  assign y30200 = ~1'b0 ;
  assign y30201 = ~1'b0 ;
  assign y30202 = ~n50225 ;
  assign y30203 = ~n50226 ;
  assign y30204 = ~n50227 ;
  assign y30205 = ~1'b0 ;
  assign y30206 = ~n50228 ;
  assign y30207 = ~1'b0 ;
  assign y30208 = ~n50232 ;
  assign y30209 = ~1'b0 ;
  assign y30210 = ~1'b0 ;
  assign y30211 = ~n50233 ;
  assign y30212 = ~n50236 ;
  assign y30213 = ~n50237 ;
  assign y30214 = ~n42353 ;
  assign y30215 = ~n50239 ;
  assign y30216 = ~1'b0 ;
  assign y30217 = ~1'b0 ;
  assign y30218 = ~1'b0 ;
  assign y30219 = ~n50244 ;
  assign y30220 = ~n17940 ;
  assign y30221 = n50245 ;
  assign y30222 = ~1'b0 ;
  assign y30223 = ~n50247 ;
  assign y30224 = ~n50248 ;
  assign y30225 = ~n50250 ;
  assign y30226 = n50251 ;
  assign y30227 = ~n50256 ;
  assign y30228 = ~n50258 ;
  assign y30229 = ~1'b0 ;
  assign y30230 = n50262 ;
  assign y30231 = ~n50263 ;
  assign y30232 = ~n50265 ;
  assign y30233 = ~n50268 ;
  assign y30234 = n50272 ;
  assign y30235 = n50273 ;
  assign y30236 = ~1'b0 ;
  assign y30237 = ~1'b0 ;
  assign y30238 = ~1'b0 ;
  assign y30239 = ~1'b0 ;
  assign y30240 = ~n50274 ;
  assign y30241 = ~1'b0 ;
  assign y30242 = n50021 ;
  assign y30243 = ~1'b0 ;
  assign y30244 = ~n50275 ;
  assign y30245 = ~n50279 ;
  assign y30246 = ~1'b0 ;
  assign y30247 = n1847 ;
  assign y30248 = ~n50280 ;
  assign y30249 = n8513 ;
  assign y30250 = n50282 ;
  assign y30251 = n19436 ;
  assign y30252 = ~n50286 ;
  assign y30253 = n50297 ;
  assign y30254 = ~1'b0 ;
  assign y30255 = n50302 ;
  assign y30256 = n50304 ;
  assign y30257 = ~1'b0 ;
  assign y30258 = ~1'b0 ;
  assign y30259 = n50306 ;
  assign y30260 = n22628 ;
  assign y30261 = n50311 ;
  assign y30262 = ~n50313 ;
  assign y30263 = ~1'b0 ;
  assign y30264 = n50314 ;
  assign y30265 = n50315 ;
  assign y30266 = n50316 ;
  assign y30267 = ~n50318 ;
  assign y30268 = n50319 ;
  assign y30269 = ~n50320 ;
  assign y30270 = ~n50321 ;
  assign y30271 = ~n50323 ;
  assign y30272 = ~n17331 ;
  assign y30273 = ~1'b0 ;
  assign y30274 = ~1'b0 ;
  assign y30275 = ~1'b0 ;
  assign y30276 = ~n21146 ;
  assign y30277 = ~n50324 ;
  assign y30278 = ~n18238 ;
  assign y30279 = ~n50327 ;
  assign y30280 = ~n22571 ;
  assign y30281 = ~n50328 ;
  assign y30282 = ~1'b0 ;
  assign y30283 = n6265 ;
  assign y30284 = ~n50329 ;
  assign y30285 = n11302 ;
  assign y30286 = ~n50332 ;
  assign y30287 = n50334 ;
  assign y30288 = ~n50335 ;
  assign y30289 = ~n50337 ;
  assign y30290 = ~n50341 ;
  assign y30291 = n50342 ;
  assign y30292 = ~1'b0 ;
  assign y30293 = ~n50344 ;
  assign y30294 = ~n50347 ;
  assign y30295 = ~1'b0 ;
  assign y30296 = ~n50348 ;
  assign y30297 = ~1'b0 ;
  assign y30298 = n50349 ;
  assign y30299 = n50350 ;
  assign y30300 = n29975 ;
  assign y30301 = ~n50351 ;
  assign y30302 = ~1'b0 ;
  assign y30303 = ~n50354 ;
  assign y30304 = ~1'b0 ;
  assign y30305 = ~n50359 ;
  assign y30306 = n50365 ;
  assign y30307 = ~n50367 ;
  assign y30308 = n50368 ;
  assign y30309 = ~1'b0 ;
  assign y30310 = n50370 ;
  assign y30311 = n50371 ;
  assign y30312 = ~n50373 ;
  assign y30313 = ~1'b0 ;
  assign y30314 = ~1'b0 ;
  assign y30315 = ~n50375 ;
  assign y30316 = n50379 ;
  assign y30317 = n46326 ;
  assign y30318 = n50380 ;
  assign y30319 = ~1'b0 ;
  assign y30320 = n50384 ;
  assign y30321 = n50385 ;
  assign y30322 = n23377 ;
  assign y30323 = ~1'b0 ;
  assign y30324 = ~n50386 ;
  assign y30325 = ~n50392 ;
  assign y30326 = ~n50395 ;
  assign y30327 = ~1'b0 ;
  assign y30328 = ~n50403 ;
  assign y30329 = ~n50404 ;
  assign y30330 = ~1'b0 ;
  assign y30331 = ~1'b0 ;
  assign y30332 = n50405 ;
  assign y30333 = ~n50408 ;
  assign y30334 = n50410 ;
  assign y30335 = ~n50411 ;
  assign y30336 = ~n9808 ;
  assign y30337 = n50415 ;
  assign y30338 = 1'b0 ;
  assign y30339 = ~n50417 ;
  assign y30340 = ~1'b0 ;
  assign y30341 = n50421 ;
  assign y30342 = ~n50425 ;
  assign y30343 = ~n19164 ;
  assign y30344 = n50426 ;
  assign y30345 = n50432 ;
  assign y30346 = ~n50434 ;
  assign y30347 = ~1'b0 ;
  assign y30348 = ~1'b0 ;
  assign y30349 = n50435 ;
  assign y30350 = ~1'b0 ;
  assign y30351 = ~n50436 ;
  assign y30352 = ~n50439 ;
  assign y30353 = ~n50440 ;
  assign y30354 = ~n50444 ;
  assign y30355 = ~n50447 ;
  assign y30356 = ~1'b0 ;
  assign y30357 = ~n4635 ;
  assign y30358 = n34355 ;
  assign y30359 = 1'b0 ;
  assign y30360 = n50449 ;
  assign y30361 = ~1'b0 ;
  assign y30362 = ~1'b0 ;
  assign y30363 = n50452 ;
  assign y30364 = ~n49165 ;
  assign y30365 = n50456 ;
  assign y30366 = n26719 ;
  assign y30367 = ~1'b0 ;
  assign y30368 = ~1'b0 ;
  assign y30369 = ~n50458 ;
  assign y30370 = ~n42988 ;
  assign y30371 = ~n50459 ;
  assign y30372 = ~1'b0 ;
  assign y30373 = n50460 ;
  assign y30374 = n50464 ;
  assign y30375 = ~n50465 ;
  assign y30376 = ~1'b0 ;
  assign y30377 = ~n50470 ;
  assign y30378 = n50471 ;
  assign y30379 = n3731 ;
  assign y30380 = ~n50472 ;
  assign y30381 = ~1'b0 ;
  assign y30382 = ~1'b0 ;
  assign y30383 = ~n50474 ;
  assign y30384 = ~n50476 ;
  assign y30385 = ~1'b0 ;
  assign y30386 = n50479 ;
  assign y30387 = ~n49791 ;
  assign y30388 = ~n50482 ;
  assign y30389 = n50483 ;
  assign y30390 = ~n50484 ;
  assign y30391 = ~n50487 ;
  assign y30392 = ~1'b0 ;
  assign y30393 = n36876 ;
  assign y30394 = n50488 ;
  assign y30395 = ~n19982 ;
  assign y30396 = ~n50489 ;
  assign y30397 = n20709 ;
  assign y30398 = ~n50492 ;
  assign y30399 = ~n50493 ;
  assign y30400 = ~1'b0 ;
  assign y30401 = ~1'b0 ;
  assign y30402 = ~1'b0 ;
  assign y30403 = ~1'b0 ;
  assign y30404 = ~1'b0 ;
  assign y30405 = ~1'b0 ;
  assign y30406 = ~1'b0 ;
  assign y30407 = ~n50494 ;
  assign y30408 = n50495 ;
  assign y30409 = n50502 ;
  assign y30410 = n50503 ;
  assign y30411 = n7532 ;
  assign y30412 = ~1'b0 ;
endmodule
