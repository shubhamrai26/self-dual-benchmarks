module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 , y256 , y257 , y258 , y259 , y260 , y261 , y262 , y263 , y264 , y265 , y266 , y267 , y268 , y269 , y270 , y271 , y272 , y273 , y274 , y275 , y276 , y277 , y278 , y279 , y280 , y281 , y282 , y283 , y284 , y285 , y286 , y287 , y288 , y289 , y290 , y291 , y292 , y293 , y294 , y295 , y296 , y297 , y298 , y299 , y300 , y301 , y302 , y303 , y304 , y305 , y306 , y307 , y308 , y309 , y310 , y311 , y312 , y313 , y314 , y315 , y316 , y317 , y318 , y319 , y320 , y321 , y322 , y323 , y324 , y325 , y326 , y327 , y328 , y329 , y330 , y331 , y332 , y333 , y334 , y335 , y336 , y337 , y338 , y339 , y340 , y341 , y342 , y343 , y344 , y345 , y346 , y347 , y348 , y349 , y350 , y351 , y352 , y353 , y354 , y355 , y356 , y357 , y358 , y359 , y360 , y361 , y362 , y363 , y364 , y365 , y366 , y367 , y368 , y369 , y370 , y371 , y372 , y373 , y374 , y375 , y376 , y377 , y378 , y379 , y380 , y381 , y382 , y383 , y384 , y385 , y386 , y387 , y388 , y389 , y390 , y391 , y392 , y393 , y394 , y395 , y396 , y397 , y398 , y399 , y400 , y401 , y402 , y403 , y404 , y405 , y406 , y407 , y408 , y409 , y410 , y411 , y412 , y413 , y414 , y415 , y416 , y417 , y418 , y419 , y420 , y421 , y422 , y423 , y424 , y425 , y426 , y427 , y428 , y429 , y430 , y431 , y432 , y433 , y434 , y435 , y436 , y437 , y438 , y439 , y440 , y441 , y442 , y443 , y444 , y445 , y446 , y447 , y448 , y449 , y450 , y451 , y452 , y453 , y454 , y455 , y456 , y457 , y458 , y459 , y460 , y461 , y462 , y463 , y464 , y465 , y466 , y467 , y468 , y469 , y470 , y471 , y472 , y473 , y474 , y475 , y476 , y477 , y478 , y479 , y480 , y481 , y482 , y483 , y484 , y485 , y486 , y487 , y488 , y489 , y490 , y491 , y492 , y493 , y494 , y495 , y496 , y497 , y498 , y499 , y500 , y501 , y502 , y503 , y504 , y505 , y506 , y507 , y508 , y509 , y510 , y511 , y512 , y513 , y514 , y515 , y516 , y517 , y518 , y519 , y520 , y521 , y522 , y523 , y524 , y525 , y526 , y527 , y528 , y529 , y530 , y531 , y532 , y533 , y534 , y535 , y536 , y537 , y538 , y539 , y540 , y541 , y542 , y543 , y544 , y545 , y546 , y547 , y548 , y549 , y550 , y551 , y552 , y553 , y554 , y555 , y556 , y557 , y558 , y559 , y560 , y561 , y562 , y563 , y564 , y565 , y566 , y567 , y568 , y569 , y570 , y571 , y572 , y573 , y574 , y575 , y576 , y577 , y578 , y579 , y580 , y581 , y582 , y583 , y584 , y585 , y586 , y587 , y588 , y589 , y590 , y591 , y592 , y593 , y594 , y595 , y596 , y597 , y598 , y599 , y600 , y601 , y602 , y603 , y604 , y605 , y606 , y607 , y608 , y609 , y610 , y611 , y612 , y613 , y614 , y615 , y616 , y617 , y618 , y619 , y620 , y621 , y622 , y623 , y624 , y625 , y626 , y627 , y628 , y629 , y630 , y631 , y632 , y633 , y634 , y635 , y636 , y637 , y638 , y639 , y640 , y641 , y642 , y643 , y644 , y645 , y646 , y647 , y648 , y649 , y650 , y651 , y652 , y653 , y654 , y655 , y656 , y657 , y658 , y659 , y660 , y661 , y662 , y663 , y664 , y665 , y666 , y667 , y668 , y669 , y670 , y671 , y672 , y673 , y674 , y675 , y676 , y677 , y678 , y679 , y680 , y681 , y682 , y683 , y684 , y685 , y686 , y687 , y688 , y689 , y690 , y691 , y692 , y693 , y694 , y695 , y696 , y697 , y698 , y699 , y700 , y701 , y702 , y703 , y704 , y705 , y706 , y707 , y708 , y709 , y710 , y711 , y712 , y713 , y714 , y715 , y716 , y717 , y718 , y719 , y720 , y721 , y722 , y723 , y724 , y725 , y726 , y727 , y728 , y729 , y730 , y731 , y732 , y733 , y734 , y735 , y736 , y737 , y738 , y739 , y740 , y741 , y742 , y743 , y744 , y745 , y746 , y747 , y748 , y749 , y750 , y751 , y752 , y753 , y754 , y755 , y756 , y757 , y758 , y759 , y760 , y761 , y762 , y763 , y764 , y765 , y766 , y767 , y768 , y769 , y770 , y771 , y772 , y773 , y774 , y775 , y776 , y777 , y778 , y779 , y780 , y781 , y782 , y783 , y784 , y785 , y786 , y787 , y788 , y789 , y790 , y791 , y792 , y793 , y794 , y795 , y796 , y797 , y798 , y799 , y800 , y801 , y802 , y803 , y804 , y805 , y806 , y807 , y808 , y809 , y810 , y811 , y812 , y813 , y814 , y815 , y816 , y817 , y818 , y819 , y820 , y821 , y822 , y823 , y824 , y825 , y826 , y827 , y828 , y829 , y830 , y831 , y832 , y833 , y834 , y835 , y836 , y837 , y838 , y839 , y840 , y841 , y842 , y843 , y844 , y845 , y846 , y847 , y848 , y849 , y850 , y851 , y852 , y853 , y854 , y855 , y856 , y857 , y858 , y859 , y860 , y861 , y862 , y863 , y864 , y865 , y866 , y867 , y868 , y869 , y870 , y871 , y872 , y873 , y874 , y875 , y876 , y877 , y878 , y879 , y880 , y881 , y882 , y883 , y884 , y885 , y886 , y887 , y888 , y889 , y890 , y891 , y892 , y893 , y894 , y895 , y896 , y897 , y898 , y899 , y900 , y901 , y902 , y903 , y904 , y905 , y906 , y907 , y908 , y909 , y910 , y911 , y912 , y913 , y914 , y915 , y916 , y917 , y918 , y919 , y920 , y921 , y922 , y923 , y924 , y925 , y926 , y927 , y928 , y929 , y930 , y931 , y932 , y933 , y934 , y935 , y936 , y937 , y938 , y939 , y940 , y941 , y942 , y943 , y944 , y945 , y946 , y947 , y948 , y949 , y950 , y951 , y952 , y953 , y954 , y955 , y956 , y957 , y958 , y959 , y960 , y961 , y962 , y963 , y964 , y965 , y966 , y967 , y968 , y969 , y970 , y971 , y972 , y973 , y974 , y975 , y976 , y977 , y978 , y979 , y980 , y981 , y982 , y983 , y984 , y985 , y986 , y987 , y988 , y989 , y990 , y991 , y992 , y993 , y994 , y995 , y996 , y997 , y998 , y999 , y1000 , y1001 , y1002 , y1003 , y1004 , y1005 , y1006 , y1007 , y1008 , y1009 , y1010 , y1011 , y1012 , y1013 , y1014 , y1015 , y1016 , y1017 , y1018 , y1019 , y1020 , y1021 , y1022 , y1023 , y1024 , y1025 , y1026 , y1027 , y1028 , y1029 , y1030 , y1031 , y1032 , y1033 , y1034 , y1035 , y1036 , y1037 , y1038 , y1039 , y1040 , y1041 , y1042 , y1043 , y1044 , y1045 , y1046 , y1047 , y1048 , y1049 , y1050 , y1051 , y1052 , y1053 , y1054 , y1055 , y1056 , y1057 , y1058 , y1059 , y1060 , y1061 , y1062 , y1063 , y1064 , y1065 , y1066 , y1067 , y1068 , y1069 , y1070 , y1071 , y1072 , y1073 , y1074 , y1075 , y1076 , y1077 , y1078 , y1079 , y1080 , y1081 , y1082 , y1083 , y1084 , y1085 , y1086 , y1087 , y1088 , y1089 , y1090 , y1091 , y1092 , y1093 , y1094 , y1095 , y1096 , y1097 , y1098 , y1099 , y1100 , y1101 , y1102 , y1103 , y1104 , y1105 , y1106 , y1107 , y1108 , y1109 , y1110 , y1111 , y1112 , y1113 , y1114 , y1115 , y1116 , y1117 , y1118 , y1119 , y1120 , y1121 , y1122 , y1123 , y1124 , y1125 , y1126 , y1127 , y1128 , y1129 , y1130 , y1131 , y1132 , y1133 , y1134 , y1135 , y1136 , y1137 , y1138 , y1139 , y1140 , y1141 , y1142 , y1143 , y1144 , y1145 , y1146 , y1147 , y1148 , y1149 , y1150 , y1151 , y1152 , y1153 , y1154 , y1155 , y1156 , y1157 , y1158 , y1159 , y1160 , y1161 , y1162 , y1163 , y1164 , y1165 , y1166 , y1167 , y1168 , y1169 , y1170 , y1171 , y1172 , y1173 , y1174 , y1175 , y1176 , y1177 , y1178 , y1179 , y1180 , y1181 , y1182 , y1183 , y1184 , y1185 , y1186 , y1187 , y1188 , y1189 , y1190 , y1191 , y1192 , y1193 , y1194 , y1195 , y1196 , y1197 , y1198 , y1199 , y1200 , y1201 , y1202 , y1203 , y1204 , y1205 , y1206 , y1207 , y1208 , y1209 , y1210 , y1211 , y1212 , y1213 , y1214 , y1215 , y1216 , y1217 , y1218 , y1219 , y1220 , y1221 , y1222 , y1223 , y1224 , y1225 , y1226 , y1227 , y1228 , y1229 , y1230 , y1231 , y1232 , y1233 , y1234 , y1235 , y1236 , y1237 , y1238 , y1239 , y1240 , y1241 , y1242 , y1243 , y1244 , y1245 , y1246 , y1247 , y1248 , y1249 , y1250 , y1251 , y1252 , y1253 , y1254 , y1255 , y1256 , y1257 , y1258 , y1259 , y1260 , y1261 , y1262 , y1263 , y1264 , y1265 , y1266 , y1267 , y1268 , y1269 , y1270 , y1271 , y1272 , y1273 , y1274 , y1275 , y1276 , y1277 , y1278 , y1279 , y1280 , y1281 , y1282 , y1283 , y1284 , y1285 , y1286 , y1287 , y1288 , y1289 , y1290 , y1291 , y1292 , y1293 , y1294 , y1295 , y1296 , y1297 , y1298 , y1299 , y1300 , y1301 , y1302 , y1303 , y1304 , y1305 , y1306 , y1307 , y1308 , y1309 , y1310 , y1311 , y1312 , y1313 , y1314 , y1315 , y1316 , y1317 , y1318 , y1319 , y1320 , y1321 , y1322 , y1323 , y1324 , y1325 , y1326 , y1327 , y1328 , y1329 , y1330 , y1331 , y1332 , y1333 , y1334 , y1335 , y1336 , y1337 , y1338 , y1339 , y1340 , y1341 , y1342 , y1343 , y1344 , y1345 , y1346 , y1347 , y1348 , y1349 , y1350 , y1351 , y1352 , y1353 , y1354 , y1355 , y1356 , y1357 , y1358 , y1359 , y1360 , y1361 , y1362 , y1363 , y1364 , y1365 , y1366 , y1367 , y1368 , y1369 , y1370 , y1371 , y1372 , y1373 , y1374 , y1375 , y1376 , y1377 , y1378 , y1379 , y1380 , y1381 , y1382 , y1383 , y1384 , y1385 , y1386 , y1387 , y1388 , y1389 , y1390 , y1391 , y1392 , y1393 , y1394 , y1395 , y1396 , y1397 , y1398 , y1399 , y1400 , y1401 , y1402 , y1403 , y1404 , y1405 , y1406 , y1407 , y1408 , y1409 , y1410 , y1411 , y1412 , y1413 , y1414 , y1415 , y1416 , y1417 , y1418 , y1419 , y1420 , y1421 , y1422 , y1423 , y1424 , y1425 , y1426 , y1427 , y1428 , y1429 , y1430 , y1431 , y1432 , y1433 , y1434 , y1435 , y1436 , y1437 , y1438 , y1439 , y1440 , y1441 , y1442 , y1443 , y1444 , y1445 , y1446 , y1447 , y1448 , y1449 , y1450 , y1451 , y1452 , y1453 , y1454 , y1455 , y1456 , y1457 , y1458 , y1459 , y1460 , y1461 , y1462 , y1463 , y1464 , y1465 , y1466 , y1467 , y1468 , y1469 , y1470 , y1471 , y1472 , y1473 , y1474 , y1475 , y1476 , y1477 , y1478 , y1479 , y1480 , y1481 , y1482 , y1483 , y1484 , y1485 , y1486 , y1487 , y1488 , y1489 , y1490 , y1491 , y1492 , y1493 , y1494 , y1495 , y1496 , y1497 , y1498 , y1499 , y1500 , y1501 , y1502 , y1503 , y1504 , y1505 , y1506 , y1507 , y1508 , y1509 , y1510 , y1511 , y1512 , y1513 , y1514 , y1515 , y1516 , y1517 , y1518 , y1519 , y1520 , y1521 , y1522 , y1523 , y1524 , y1525 , y1526 , y1527 , y1528 , y1529 , y1530 , y1531 , y1532 , y1533 , y1534 , y1535 , y1536 , y1537 , y1538 , y1539 , y1540 , y1541 , y1542 , y1543 , y1544 , y1545 , y1546 , y1547 , y1548 , y1549 , y1550 , y1551 , y1552 , y1553 , y1554 , y1555 , y1556 , y1557 , y1558 , y1559 , y1560 , y1561 , y1562 , y1563 , y1564 , y1565 , y1566 , y1567 , y1568 , y1569 , y1570 , y1571 , y1572 , y1573 , y1574 , y1575 , y1576 , y1577 , y1578 , y1579 , y1580 , y1581 , y1582 , y1583 , y1584 , y1585 , y1586 , y1587 , y1588 , y1589 , y1590 , y1591 , y1592 , y1593 , y1594 , y1595 , y1596 , y1597 , y1598 , y1599 , y1600 , y1601 , y1602 , y1603 , y1604 , y1605 , y1606 , y1607 , y1608 , y1609 , y1610 , y1611 , y1612 , y1613 , y1614 , y1615 , y1616 , y1617 , y1618 , y1619 , y1620 , y1621 , y1622 , y1623 , y1624 , y1625 , y1626 , y1627 , y1628 , y1629 , y1630 , y1631 , y1632 , y1633 , y1634 , y1635 , y1636 , y1637 , y1638 , y1639 , y1640 , y1641 , y1642 , y1643 , y1644 , y1645 , y1646 , y1647 , y1648 , y1649 , y1650 , y1651 , y1652 , y1653 , y1654 , y1655 , y1656 , y1657 , y1658 , y1659 , y1660 , y1661 , y1662 , y1663 , y1664 , y1665 , y1666 , y1667 , y1668 , y1669 , y1670 , y1671 , y1672 , y1673 , y1674 , y1675 , y1676 , y1677 , y1678 , y1679 , y1680 , y1681 , y1682 , y1683 , y1684 , y1685 , y1686 , y1687 , y1688 , y1689 , y1690 , y1691 , y1692 , y1693 , y1694 , y1695 , y1696 , y1697 , y1698 , y1699 , y1700 , y1701 , y1702 , y1703 , y1704 , y1705 , y1706 , y1707 , y1708 , y1709 , y1710 , y1711 , y1712 , y1713 , y1714 , y1715 , y1716 , y1717 , y1718 , y1719 , y1720 , y1721 , y1722 , y1723 , y1724 , y1725 , y1726 , y1727 , y1728 , y1729 , y1730 , y1731 , y1732 , y1733 , y1734 , y1735 , y1736 , y1737 , y1738 , y1739 , y1740 , y1741 , y1742 , y1743 , y1744 , y1745 , y1746 , y1747 , y1748 , y1749 , y1750 , y1751 , y1752 , y1753 , y1754 , y1755 , y1756 , y1757 , y1758 , y1759 , y1760 , y1761 , y1762 , y1763 , y1764 , y1765 , y1766 , y1767 , y1768 , y1769 , y1770 , y1771 , y1772 , y1773 , y1774 , y1775 , y1776 , y1777 , y1778 , y1779 , y1780 , y1781 , y1782 , y1783 , y1784 , y1785 , y1786 , y1787 , y1788 , y1789 , y1790 , y1791 , y1792 , y1793 , y1794 , y1795 , y1796 , y1797 , y1798 , y1799 , y1800 , y1801 , y1802 , y1803 , y1804 , y1805 , y1806 , y1807 , y1808 , y1809 , y1810 , y1811 , y1812 , y1813 , y1814 , y1815 , y1816 , y1817 , y1818 , y1819 , y1820 , y1821 , y1822 , y1823 , y1824 , y1825 , y1826 , y1827 , y1828 , y1829 , y1830 , y1831 , y1832 , y1833 , y1834 , y1835 , y1836 , y1837 , y1838 , y1839 , y1840 , y1841 , y1842 , y1843 , y1844 , y1845 , y1846 , y1847 , y1848 , y1849 , y1850 , y1851 , y1852 , y1853 , y1854 , y1855 , y1856 , y1857 , y1858 , y1859 , y1860 , y1861 , y1862 , y1863 , y1864 , y1865 , y1866 , y1867 , y1868 , y1869 , y1870 , y1871 , y1872 , y1873 , y1874 , y1875 , y1876 , y1877 , y1878 , y1879 , y1880 , y1881 , y1882 , y1883 , y1884 , y1885 , y1886 , y1887 , y1888 , y1889 , y1890 , y1891 , y1892 , y1893 , y1894 , y1895 , y1896 , y1897 , y1898 , y1899 , y1900 , y1901 , y1902 , y1903 , y1904 , y1905 , y1906 , y1907 , y1908 , y1909 , y1910 , y1911 , y1912 , y1913 , y1914 , y1915 , y1916 , y1917 , y1918 , y1919 , y1920 , y1921 , y1922 , y1923 , y1924 , y1925 , y1926 , y1927 , y1928 , y1929 , y1930 , y1931 , y1932 , y1933 , y1934 , y1935 , y1936 , y1937 , y1938 , y1939 , y1940 , y1941 , y1942 , y1943 , y1944 , y1945 , y1946 , y1947 , y1948 , y1949 , y1950 , y1951 , y1952 , y1953 , y1954 , y1955 , y1956 , y1957 , y1958 , y1959 , y1960 , y1961 , y1962 , y1963 , y1964 , y1965 , y1966 , y1967 , y1968 , y1969 , y1970 , y1971 , y1972 , y1973 , y1974 , y1975 , y1976 , y1977 , y1978 , y1979 , y1980 , y1981 , y1982 , y1983 , y1984 , y1985 , y1986 , y1987 , y1988 , y1989 , y1990 , y1991 , y1992 , y1993 , y1994 , y1995 , y1996 , y1997 , y1998 , y1999 , y2000 , y2001 , y2002 , y2003 , y2004 , y2005 , y2006 , y2007 , y2008 , y2009 , y2010 , y2011 , y2012 , y2013 , y2014 , y2015 , y2016 , y2017 , y2018 , y2019 , y2020 , y2021 , y2022 , y2023 , y2024 , y2025 , y2026 , y2027 , y2028 , y2029 , y2030 , y2031 , y2032 , y2033 , y2034 , y2035 , y2036 , y2037 , y2038 , y2039 , y2040 , y2041 , y2042 , y2043 , y2044 , y2045 , y2046 , y2047 , y2048 , y2049 , y2050 , y2051 , y2052 , y2053 , y2054 , y2055 , y2056 , y2057 , y2058 , y2059 , y2060 , y2061 , y2062 , y2063 , y2064 , y2065 , y2066 , y2067 , y2068 , y2069 , y2070 , y2071 , y2072 , y2073 , y2074 , y2075 , y2076 , y2077 , y2078 , y2079 , y2080 , y2081 , y2082 , y2083 , y2084 , y2085 , y2086 , y2087 , y2088 , y2089 , y2090 , y2091 , y2092 , y2093 , y2094 , y2095 , y2096 , y2097 , y2098 , y2099 , y2100 , y2101 , y2102 , y2103 , y2104 , y2105 , y2106 , y2107 , y2108 , y2109 , y2110 , y2111 , y2112 , y2113 , y2114 , y2115 , y2116 , y2117 , y2118 , y2119 , y2120 , y2121 , y2122 , y2123 , y2124 , y2125 , y2126 , y2127 , y2128 , y2129 , y2130 , y2131 , y2132 , y2133 , y2134 , y2135 , y2136 , y2137 , y2138 , y2139 , y2140 , y2141 , y2142 , y2143 , y2144 , y2145 , y2146 , y2147 , y2148 , y2149 , y2150 , y2151 , y2152 , y2153 , y2154 , y2155 , y2156 , y2157 , y2158 , y2159 , y2160 , y2161 , y2162 , y2163 , y2164 , y2165 , y2166 , y2167 , y2168 , y2169 , y2170 , y2171 , y2172 , y2173 , y2174 , y2175 , y2176 , y2177 , y2178 , y2179 , y2180 , y2181 , y2182 , y2183 , y2184 , y2185 , y2186 , y2187 , y2188 , y2189 , y2190 , y2191 , y2192 , y2193 , y2194 , y2195 , y2196 , y2197 , y2198 , y2199 , y2200 , y2201 , y2202 , y2203 , y2204 , y2205 , y2206 , y2207 , y2208 , y2209 , y2210 , y2211 , y2212 , y2213 , y2214 , y2215 , y2216 , y2217 , y2218 , y2219 , y2220 , y2221 , y2222 , y2223 , y2224 , y2225 , y2226 , y2227 , y2228 , y2229 , y2230 , y2231 , y2232 , y2233 , y2234 , y2235 , y2236 , y2237 , y2238 , y2239 , y2240 , y2241 , y2242 , y2243 , y2244 , y2245 , y2246 , y2247 , y2248 , y2249 , y2250 , y2251 , y2252 , y2253 , y2254 , y2255 , y2256 , y2257 , y2258 , y2259 , y2260 , y2261 , y2262 , y2263 , y2264 , y2265 , y2266 , y2267 , y2268 , y2269 , y2270 , y2271 , y2272 , y2273 , y2274 , y2275 , y2276 , y2277 , y2278 , y2279 , y2280 , y2281 , y2282 , y2283 , y2284 , y2285 , y2286 , y2287 , y2288 , y2289 , y2290 , y2291 , y2292 , y2293 , y2294 , y2295 , y2296 , y2297 , y2298 , y2299 , y2300 , y2301 , y2302 , y2303 , y2304 , y2305 , y2306 , y2307 , y2308 , y2309 , y2310 , y2311 , y2312 , y2313 , y2314 , y2315 , y2316 , y2317 , y2318 , y2319 , y2320 , y2321 , y2322 , y2323 , y2324 , y2325 , y2326 , y2327 , y2328 , y2329 , y2330 , y2331 , y2332 , y2333 , y2334 , y2335 , y2336 , y2337 , y2338 , y2339 , y2340 , y2341 , y2342 , y2343 , y2344 , y2345 , y2346 , y2347 , y2348 , y2349 , y2350 , y2351 , y2352 , y2353 , y2354 , y2355 , y2356 , y2357 , y2358 , y2359 , y2360 , y2361 , y2362 , y2363 , y2364 , y2365 , y2366 , y2367 , y2368 , y2369 , y2370 , y2371 , y2372 , y2373 , y2374 , y2375 , y2376 , y2377 , y2378 , y2379 , y2380 , y2381 , y2382 , y2383 , y2384 , y2385 , y2386 , y2387 , y2388 , y2389 , y2390 , y2391 , y2392 , y2393 , y2394 , y2395 , y2396 , y2397 , y2398 , y2399 , y2400 , y2401 , y2402 , y2403 , y2404 , y2405 , y2406 , y2407 , y2408 , y2409 , y2410 , y2411 , y2412 , y2413 , y2414 , y2415 , y2416 , y2417 , y2418 , y2419 , y2420 , y2421 , y2422 , y2423 , y2424 , y2425 , y2426 , y2427 , y2428 , y2429 , y2430 , y2431 , y2432 , y2433 , y2434 , y2435 , y2436 , y2437 , y2438 , y2439 , y2440 , y2441 , y2442 , y2443 , y2444 , y2445 , y2446 , y2447 , y2448 , y2449 , y2450 , y2451 , y2452 , y2453 , y2454 , y2455 , y2456 , y2457 , y2458 , y2459 , y2460 , y2461 , y2462 , y2463 , y2464 , y2465 , y2466 , y2467 , y2468 , y2469 , y2470 , y2471 , y2472 , y2473 , y2474 , y2475 , y2476 , y2477 , y2478 , y2479 , y2480 , y2481 , y2482 , y2483 , y2484 , y2485 , y2486 , y2487 , y2488 , y2489 , y2490 , y2491 , y2492 , y2493 , y2494 , y2495 , y2496 , y2497 , y2498 , y2499 , y2500 , y2501 , y2502 , y2503 , y2504 , y2505 , y2506 , y2507 , y2508 , y2509 , y2510 , y2511 , y2512 , y2513 , y2514 , y2515 , y2516 , y2517 , y2518 , y2519 , y2520 , y2521 , y2522 , y2523 , y2524 , y2525 , y2526 , y2527 , y2528 , y2529 , y2530 , y2531 , y2532 , y2533 , y2534 , y2535 , y2536 , y2537 , y2538 , y2539 , y2540 , y2541 , y2542 , y2543 , y2544 , y2545 , y2546 , y2547 , y2548 , y2549 , y2550 , y2551 , y2552 , y2553 , y2554 , y2555 , y2556 , y2557 , y2558 , y2559 , y2560 , y2561 , y2562 , y2563 , y2564 , y2565 , y2566 , y2567 , y2568 , y2569 , y2570 , y2571 , y2572 , y2573 , y2574 , y2575 , y2576 , y2577 , y2578 , y2579 , y2580 , y2581 , y2582 , y2583 , y2584 , y2585 , y2586 , y2587 , y2588 , y2589 , y2590 , y2591 , y2592 , y2593 , y2594 , y2595 , y2596 , y2597 , y2598 , y2599 , y2600 , y2601 , y2602 , y2603 , y2604 , y2605 , y2606 , y2607 , y2608 , y2609 , y2610 , y2611 , y2612 , y2613 , y2614 , y2615 , y2616 , y2617 , y2618 , y2619 , y2620 , y2621 , y2622 , y2623 , y2624 , y2625 , y2626 , y2627 , y2628 , y2629 , y2630 , y2631 , y2632 , y2633 , y2634 , y2635 , y2636 , y2637 , y2638 , y2639 , y2640 , y2641 , y2642 , y2643 , y2644 , y2645 , y2646 , y2647 , y2648 , y2649 , y2650 , y2651 , y2652 , y2653 , y2654 , y2655 , y2656 , y2657 , y2658 , y2659 , y2660 , y2661 , y2662 , y2663 , y2664 , y2665 , y2666 , y2667 , y2668 , y2669 , y2670 , y2671 , y2672 , y2673 , y2674 , y2675 , y2676 , y2677 , y2678 , y2679 , y2680 , y2681 , y2682 , y2683 , y2684 , y2685 , y2686 , y2687 , y2688 , y2689 , y2690 , y2691 , y2692 , y2693 , y2694 , y2695 , y2696 , y2697 , y2698 , y2699 , y2700 , y2701 , y2702 , y2703 , y2704 , y2705 , y2706 , y2707 , y2708 , y2709 , y2710 , y2711 , y2712 , y2713 , y2714 , y2715 , y2716 , y2717 , y2718 , y2719 , y2720 , y2721 , y2722 , y2723 , y2724 , y2725 , y2726 , y2727 , y2728 , y2729 , y2730 , y2731 , y2732 , y2733 , y2734 , y2735 , y2736 , y2737 , y2738 , y2739 , y2740 , y2741 , y2742 , y2743 , y2744 , y2745 , y2746 , y2747 , y2748 , y2749 , y2750 , y2751 , y2752 , y2753 , y2754 , y2755 , y2756 , y2757 , y2758 , y2759 , y2760 , y2761 , y2762 , y2763 , y2764 , y2765 , y2766 , y2767 , y2768 , y2769 , y2770 , y2771 , y2772 , y2773 , y2774 , y2775 , y2776 , y2777 , y2778 , y2779 , y2780 , y2781 , y2782 , y2783 , y2784 , y2785 , y2786 , y2787 , y2788 , y2789 , y2790 , y2791 , y2792 , y2793 , y2794 , y2795 , y2796 , y2797 , y2798 , y2799 , y2800 , y2801 , y2802 , y2803 , y2804 , y2805 , y2806 , y2807 , y2808 , y2809 , y2810 , y2811 , y2812 , y2813 , y2814 , y2815 , y2816 , y2817 , y2818 , y2819 , y2820 , y2821 , y2822 , y2823 , y2824 , y2825 , y2826 , y2827 , y2828 , y2829 , y2830 , y2831 , y2832 , y2833 , y2834 , y2835 , y2836 , y2837 , y2838 , y2839 , y2840 , y2841 , y2842 , y2843 , y2844 , y2845 , y2846 , y2847 , y2848 , y2849 , y2850 , y2851 , y2852 , y2853 , y2854 , y2855 , y2856 , y2857 , y2858 , y2859 , y2860 , y2861 , y2862 , y2863 , y2864 , y2865 , y2866 , y2867 , y2868 , y2869 , y2870 , y2871 , y2872 , y2873 , y2874 , y2875 , y2876 , y2877 , y2878 , y2879 , y2880 , y2881 , y2882 , y2883 , y2884 , y2885 , y2886 , y2887 , y2888 , y2889 , y2890 , y2891 , y2892 , y2893 , y2894 , y2895 , y2896 , y2897 , y2898 , y2899 , y2900 , y2901 , y2902 , y2903 , y2904 , y2905 , y2906 , y2907 , y2908 , y2909 , y2910 , y2911 , y2912 , y2913 , y2914 , y2915 , y2916 , y2917 , y2918 , y2919 , y2920 , y2921 , y2922 , y2923 , y2924 , y2925 , y2926 , y2927 , y2928 , y2929 , y2930 , y2931 , y2932 , y2933 , y2934 , y2935 , y2936 , y2937 , y2938 , y2939 , y2940 , y2941 , y2942 , y2943 , y2944 , y2945 , y2946 , y2947 , y2948 , y2949 , y2950 , y2951 , y2952 , y2953 , y2954 , y2955 , y2956 , y2957 , y2958 , y2959 , y2960 , y2961 , y2962 , y2963 , y2964 , y2965 , y2966 , y2967 , y2968 , y2969 , y2970 , y2971 , y2972 , y2973 , y2974 , y2975 , y2976 , y2977 , y2978 , y2979 , y2980 , y2981 , y2982 , y2983 , y2984 , y2985 , y2986 , y2987 , y2988 , y2989 , y2990 , y2991 , y2992 , y2993 , y2994 , y2995 , y2996 , y2997 , y2998 , y2999 , y3000 , y3001 , y3002 , y3003 , y3004 , y3005 , y3006 , y3007 , y3008 , y3009 , y3010 , y3011 , y3012 , y3013 , y3014 , y3015 , y3016 , y3017 , y3018 , y3019 , y3020 , y3021 , y3022 , y3023 , y3024 , y3025 , y3026 , y3027 , y3028 , y3029 , y3030 , y3031 , y3032 , y3033 , y3034 , y3035 , y3036 , y3037 , y3038 , y3039 , y3040 , y3041 , y3042 , y3043 , y3044 , y3045 , y3046 , y3047 , y3048 , y3049 , y3050 , y3051 , y3052 , y3053 , y3054 , y3055 , y3056 , y3057 , y3058 , y3059 , y3060 , y3061 , y3062 , y3063 , y3064 , y3065 , y3066 , y3067 , y3068 , y3069 , y3070 , y3071 , y3072 , y3073 , y3074 , y3075 , y3076 , y3077 , y3078 , y3079 , y3080 , y3081 , y3082 , y3083 , y3084 , y3085 , y3086 , y3087 , y3088 , y3089 , y3090 , y3091 , y3092 , y3093 , y3094 , y3095 , y3096 , y3097 , y3098 , y3099 , y3100 , y3101 , y3102 , y3103 , y3104 , y3105 , y3106 , y3107 , y3108 , y3109 , y3110 , y3111 , y3112 , y3113 , y3114 , y3115 , y3116 , y3117 , y3118 , y3119 , y3120 , y3121 , y3122 , y3123 , y3124 , y3125 , y3126 , y3127 , y3128 , y3129 , y3130 , y3131 , y3132 , y3133 , y3134 , y3135 , y3136 , y3137 , y3138 , y3139 , y3140 , y3141 , y3142 , y3143 , y3144 , y3145 , y3146 , y3147 , y3148 , y3149 , y3150 , y3151 , y3152 , y3153 , y3154 , y3155 , y3156 , y3157 , y3158 , y3159 , y3160 , y3161 , y3162 , y3163 , y3164 , y3165 , y3166 , y3167 , y3168 , y3169 , y3170 , y3171 , y3172 , y3173 , y3174 , y3175 , y3176 , y3177 , y3178 , y3179 , y3180 , y3181 , y3182 , y3183 , y3184 , y3185 , y3186 , y3187 , y3188 , y3189 , y3190 , y3191 , y3192 , y3193 , y3194 , y3195 , y3196 , y3197 , y3198 , y3199 , y3200 , y3201 , y3202 , y3203 , y3204 , y3205 , y3206 , y3207 , y3208 , y3209 , y3210 , y3211 , y3212 , y3213 , y3214 , y3215 , y3216 , y3217 , y3218 , y3219 , y3220 , y3221 , y3222 , y3223 , y3224 , y3225 , y3226 , y3227 , y3228 , y3229 , y3230 , y3231 , y3232 , y3233 , y3234 , y3235 , y3236 , y3237 , y3238 , y3239 , y3240 , y3241 , y3242 , y3243 , y3244 , y3245 , y3246 , y3247 , y3248 , y3249 , y3250 , y3251 , y3252 , y3253 , y3254 , y3255 , y3256 , y3257 , y3258 , y3259 , y3260 , y3261 , y3262 , y3263 , y3264 , y3265 , y3266 , y3267 , y3268 , y3269 , y3270 , y3271 , y3272 , y3273 , y3274 , y3275 , y3276 , y3277 , y3278 , y3279 , y3280 , y3281 , y3282 , y3283 , y3284 , y3285 , y3286 , y3287 , y3288 , y3289 , y3290 , y3291 , y3292 , y3293 , y3294 , y3295 , y3296 , y3297 , y3298 , y3299 , y3300 , y3301 , y3302 , y3303 , y3304 , y3305 , y3306 , y3307 , y3308 , y3309 , y3310 , y3311 , y3312 , y3313 , y3314 , y3315 , y3316 , y3317 , y3318 , y3319 , y3320 , y3321 , y3322 , y3323 , y3324 , y3325 , y3326 , y3327 , y3328 , y3329 , y3330 , y3331 , y3332 , y3333 , y3334 , y3335 , y3336 , y3337 , y3338 , y3339 , y3340 , y3341 , y3342 , y3343 , y3344 , y3345 , y3346 , y3347 , y3348 , y3349 , y3350 , y3351 , y3352 , y3353 , y3354 , y3355 , y3356 , y3357 , y3358 , y3359 , y3360 , y3361 , y3362 , y3363 , y3364 , y3365 , y3366 , y3367 , y3368 , y3369 , y3370 , y3371 , y3372 , y3373 , y3374 , y3375 , y3376 , y3377 , y3378 , y3379 , y3380 , y3381 , y3382 , y3383 , y3384 , y3385 , y3386 , y3387 , y3388 , y3389 , y3390 , y3391 , y3392 , y3393 , y3394 , y3395 , y3396 , y3397 , y3398 , y3399 , y3400 , y3401 , y3402 , y3403 , y3404 , y3405 , y3406 , y3407 , y3408 , y3409 , y3410 , y3411 , y3412 , y3413 , y3414 , y3415 , y3416 , y3417 , y3418 , y3419 , y3420 , y3421 , y3422 , y3423 , y3424 , y3425 , y3426 , y3427 , y3428 , y3429 , y3430 , y3431 , y3432 , y3433 , y3434 , y3435 , y3436 , y3437 , y3438 , y3439 , y3440 , y3441 , y3442 , y3443 , y3444 , y3445 , y3446 , y3447 , y3448 , y3449 , y3450 , y3451 , y3452 , y3453 , y3454 , y3455 , y3456 , y3457 , y3458 , y3459 , y3460 , y3461 , y3462 , y3463 , y3464 , y3465 , y3466 , y3467 , y3468 , y3469 , y3470 , y3471 , y3472 , y3473 , y3474 , y3475 , y3476 , y3477 , y3478 , y3479 , y3480 , y3481 , y3482 , y3483 , y3484 , y3485 , y3486 , y3487 , y3488 , y3489 , y3490 , y3491 , y3492 , y3493 , y3494 , y3495 , y3496 , y3497 , y3498 , y3499 , y3500 , y3501 , y3502 , y3503 , y3504 , y3505 , y3506 , y3507 , y3508 , y3509 , y3510 , y3511 , y3512 , y3513 , y3514 , y3515 , y3516 , y3517 , y3518 , y3519 , y3520 , y3521 , y3522 , y3523 , y3524 , y3525 , y3526 , y3527 , y3528 , y3529 , y3530 , y3531 , y3532 , y3533 , y3534 , y3535 , y3536 , y3537 , y3538 , y3539 , y3540 , y3541 , y3542 , y3543 , y3544 , y3545 , y3546 , y3547 , y3548 , y3549 , y3550 , y3551 , y3552 , y3553 , y3554 , y3555 , y3556 , y3557 , y3558 , y3559 , y3560 , y3561 , y3562 , y3563 , y3564 , y3565 , y3566 , y3567 , y3568 , y3569 , y3570 , y3571 , y3572 , y3573 , y3574 , y3575 , y3576 , y3577 , y3578 , y3579 , y3580 , y3581 , y3582 , y3583 , y3584 , y3585 , y3586 , y3587 , y3588 , y3589 , y3590 , y3591 , y3592 , y3593 , y3594 , y3595 , y3596 , y3597 , y3598 , y3599 , y3600 , y3601 , y3602 , y3603 , y3604 , y3605 , y3606 , y3607 , y3608 , y3609 , y3610 , y3611 , y3612 , y3613 , y3614 , y3615 , y3616 , y3617 , y3618 , y3619 , y3620 , y3621 , y3622 , y3623 , y3624 , y3625 , y3626 , y3627 , y3628 , y3629 , y3630 , y3631 , y3632 , y3633 , y3634 , y3635 , y3636 , y3637 , y3638 , y3639 , y3640 , y3641 , y3642 , y3643 , y3644 , y3645 , y3646 , y3647 , y3648 , y3649 , y3650 , y3651 , y3652 , y3653 , y3654 , y3655 , y3656 , y3657 , y3658 , y3659 , y3660 , y3661 , y3662 , y3663 , y3664 , y3665 , y3666 , y3667 , y3668 , y3669 , y3670 , y3671 , y3672 , y3673 , y3674 , y3675 , y3676 , y3677 , y3678 , y3679 , y3680 , y3681 , y3682 , y3683 , y3684 , y3685 , y3686 , y3687 , y3688 , y3689 , y3690 , y3691 , y3692 , y3693 , y3694 , y3695 , y3696 , y3697 , y3698 , y3699 , y3700 , y3701 , y3702 , y3703 , y3704 , y3705 , y3706 , y3707 , y3708 , y3709 , y3710 , y3711 , y3712 , y3713 , y3714 , y3715 , y3716 , y3717 , y3718 , y3719 , y3720 , y3721 , y3722 , y3723 , y3724 , y3725 , y3726 , y3727 , y3728 , y3729 , y3730 , y3731 , y3732 , y3733 , y3734 , y3735 , y3736 , y3737 , y3738 , y3739 , y3740 , y3741 , y3742 , y3743 , y3744 , y3745 , y3746 , y3747 , y3748 , y3749 , y3750 , y3751 , y3752 , y3753 , y3754 , y3755 , y3756 , y3757 , y3758 , y3759 , y3760 , y3761 , y3762 , y3763 , y3764 , y3765 , y3766 , y3767 , y3768 , y3769 , y3770 , y3771 , y3772 , y3773 , y3774 , y3775 , y3776 , y3777 , y3778 , y3779 , y3780 , y3781 , y3782 , y3783 , y3784 , y3785 , y3786 , y3787 , y3788 , y3789 , y3790 , y3791 , y3792 , y3793 , y3794 , y3795 , y3796 , y3797 , y3798 , y3799 , y3800 , y3801 , y3802 , y3803 , y3804 , y3805 , y3806 , y3807 , y3808 , y3809 , y3810 , y3811 , y3812 , y3813 , y3814 , y3815 , y3816 , y3817 , y3818 , y3819 , y3820 , y3821 , y3822 , y3823 , y3824 , y3825 , y3826 , y3827 , y3828 , y3829 , y3830 , y3831 , y3832 , y3833 , y3834 , y3835 , y3836 , y3837 , y3838 , y3839 , y3840 , y3841 , y3842 , y3843 , y3844 , y3845 , y3846 , y3847 , y3848 , y3849 , y3850 , y3851 , y3852 , y3853 , y3854 , y3855 , y3856 , y3857 , y3858 , y3859 , y3860 , y3861 , y3862 , y3863 , y3864 , y3865 , y3866 , y3867 , y3868 , y3869 , y3870 , y3871 , y3872 , y3873 , y3874 , y3875 , y3876 , y3877 , y3878 , y3879 , y3880 , y3881 , y3882 , y3883 , y3884 , y3885 , y3886 , y3887 , y3888 , y3889 , y3890 , y3891 , y3892 , y3893 , y3894 , y3895 , y3896 , y3897 , y3898 , y3899 , y3900 , y3901 , y3902 , y3903 , y3904 , y3905 , y3906 , y3907 , y3908 , y3909 , y3910 , y3911 , y3912 , y3913 , y3914 , y3915 , y3916 , y3917 , y3918 , y3919 , y3920 , y3921 , y3922 , y3923 , y3924 , y3925 , y3926 , y3927 , y3928 , y3929 , y3930 , y3931 , y3932 , y3933 , y3934 , y3935 , y3936 , y3937 , y3938 , y3939 , y3940 , y3941 , y3942 , y3943 , y3944 , y3945 , y3946 , y3947 , y3948 , y3949 , y3950 , y3951 , y3952 , y3953 , y3954 , y3955 , y3956 , y3957 , y3958 , y3959 , y3960 , y3961 , y3962 , y3963 , y3964 , y3965 , y3966 , y3967 , y3968 , y3969 , y3970 , y3971 , y3972 , y3973 , y3974 , y3975 , y3976 , y3977 , y3978 , y3979 , y3980 , y3981 , y3982 , y3983 , y3984 , y3985 , y3986 , y3987 , y3988 , y3989 , y3990 , y3991 , y3992 , y3993 , y3994 , y3995 , y3996 , y3997 , y3998 , y3999 , y4000 , y4001 , y4002 , y4003 , y4004 , y4005 , y4006 , y4007 , y4008 , y4009 , y4010 , y4011 , y4012 , y4013 , y4014 , y4015 , y4016 , y4017 , y4018 , y4019 , y4020 , y4021 , y4022 , y4023 , y4024 , y4025 , y4026 , y4027 , y4028 , y4029 , y4030 , y4031 , y4032 , y4033 , y4034 , y4035 , y4036 , y4037 , y4038 , y4039 , y4040 , y4041 , y4042 , y4043 , y4044 , y4045 , y4046 , y4047 , y4048 , y4049 , y4050 , y4051 , y4052 , y4053 , y4054 , y4055 , y4056 , y4057 , y4058 , y4059 , y4060 , y4061 , y4062 , y4063 , y4064 , y4065 , y4066 , y4067 , y4068 , y4069 , y4070 , y4071 , y4072 , y4073 , y4074 , y4075 , y4076 , y4077 , y4078 , y4079 , y4080 , y4081 , y4082 , y4083 , y4084 , y4085 , y4086 , y4087 , y4088 , y4089 , y4090 , y4091 , y4092 , y4093 , y4094 , y4095 , y4096 , y4097 , y4098 , y4099 , y4100 , y4101 , y4102 , y4103 , y4104 , y4105 , y4106 , y4107 , y4108 , y4109 , y4110 , y4111 , y4112 , y4113 , y4114 , y4115 , y4116 , y4117 , y4118 , y4119 , y4120 , y4121 , y4122 , y4123 , y4124 , y4125 , y4126 , y4127 , y4128 , y4129 , y4130 , y4131 , y4132 , y4133 , y4134 , y4135 , y4136 , y4137 , y4138 , y4139 , y4140 , y4141 , y4142 , y4143 , y4144 , y4145 , y4146 , y4147 , y4148 , y4149 , y4150 , y4151 , y4152 , y4153 , y4154 , y4155 , y4156 , y4157 , y4158 , y4159 , y4160 , y4161 , y4162 , y4163 , y4164 , y4165 , y4166 , y4167 , y4168 , y4169 , y4170 , y4171 , y4172 , y4173 , y4174 , y4175 , y4176 , y4177 , y4178 , y4179 , y4180 , y4181 , y4182 , y4183 , y4184 , y4185 , y4186 , y4187 , y4188 , y4189 , y4190 , y4191 , y4192 , y4193 , y4194 , y4195 , y4196 , y4197 , y4198 , y4199 , y4200 , y4201 , y4202 , y4203 , y4204 , y4205 , y4206 , y4207 , y4208 , y4209 , y4210 , y4211 , y4212 , y4213 , y4214 , y4215 , y4216 , y4217 , y4218 , y4219 , y4220 , y4221 , y4222 , y4223 , y4224 , y4225 , y4226 , y4227 , y4228 , y4229 , y4230 , y4231 , y4232 , y4233 , y4234 , y4235 , y4236 , y4237 , y4238 , y4239 , y4240 , y4241 , y4242 , y4243 , y4244 , y4245 , y4246 , y4247 , y4248 , y4249 , y4250 , y4251 , y4252 , y4253 , y4254 , y4255 , y4256 , y4257 , y4258 , y4259 , y4260 , y4261 , y4262 , y4263 , y4264 , y4265 , y4266 , y4267 , y4268 , y4269 , y4270 , y4271 , y4272 , y4273 , y4274 , y4275 , y4276 , y4277 , y4278 , y4279 , y4280 , y4281 , y4282 , y4283 , y4284 , y4285 , y4286 , y4287 , y4288 , y4289 , y4290 , y4291 , y4292 , y4293 , y4294 , y4295 , y4296 , y4297 , y4298 , y4299 , y4300 , y4301 , y4302 , y4303 , y4304 , y4305 , y4306 , y4307 , y4308 , y4309 , y4310 , y4311 , y4312 , y4313 , y4314 , y4315 , y4316 , y4317 , y4318 , y4319 , y4320 , y4321 , y4322 , y4323 , y4324 , y4325 , y4326 , y4327 , y4328 , y4329 , y4330 , y4331 , y4332 , y4333 , y4334 , y4335 , y4336 , y4337 , y4338 , y4339 , y4340 , y4341 , y4342 , y4343 , y4344 , y4345 , y4346 , y4347 , y4348 , y4349 , y4350 , y4351 , y4352 , y4353 , y4354 , y4355 , y4356 , y4357 , y4358 , y4359 , y4360 , y4361 , y4362 , y4363 , y4364 , y4365 , y4366 , y4367 , y4368 , y4369 , y4370 , y4371 , y4372 , y4373 , y4374 , y4375 , y4376 , y4377 , y4378 , y4379 , y4380 , y4381 , y4382 , y4383 , y4384 , y4385 , y4386 , y4387 , y4388 , y4389 , y4390 , y4391 , y4392 , y4393 , y4394 , y4395 , y4396 , y4397 , y4398 , y4399 , y4400 , y4401 , y4402 , y4403 , y4404 , y4405 , y4406 , y4407 , y4408 , y4409 , y4410 , y4411 , y4412 , y4413 , y4414 , y4415 , y4416 , y4417 , y4418 , y4419 , y4420 , y4421 , y4422 , y4423 , y4424 , y4425 , y4426 , y4427 , y4428 , y4429 , y4430 , y4431 , y4432 , y4433 , y4434 , y4435 , y4436 , y4437 , y4438 , y4439 , y4440 , y4441 , y4442 , y4443 , y4444 , y4445 , y4446 , y4447 , y4448 , y4449 , y4450 , y4451 , y4452 , y4453 , y4454 , y4455 , y4456 , y4457 , y4458 , y4459 , y4460 , y4461 , y4462 , y4463 , y4464 , y4465 , y4466 , y4467 , y4468 , y4469 , y4470 , y4471 , y4472 , y4473 , y4474 , y4475 , y4476 , y4477 , y4478 , y4479 , y4480 , y4481 , y4482 , y4483 , y4484 , y4485 , y4486 , y4487 , y4488 , y4489 , y4490 , y4491 , y4492 , y4493 , y4494 , y4495 , y4496 , y4497 , y4498 , y4499 , y4500 , y4501 , y4502 , y4503 , y4504 , y4505 , y4506 , y4507 , y4508 , y4509 , y4510 , y4511 , y4512 , y4513 , y4514 , y4515 , y4516 , y4517 , y4518 , y4519 , y4520 , y4521 , y4522 , y4523 , y4524 , y4525 , y4526 , y4527 , y4528 , y4529 , y4530 , y4531 , y4532 , y4533 , y4534 , y4535 , y4536 , y4537 , y4538 , y4539 , y4540 , y4541 , y4542 , y4543 , y4544 , y4545 , y4546 , y4547 , y4548 , y4549 , y4550 , y4551 , y4552 , y4553 , y4554 , y4555 , y4556 , y4557 , y4558 , y4559 , y4560 , y4561 , y4562 , y4563 , y4564 , y4565 , y4566 , y4567 , y4568 , y4569 , y4570 , y4571 , y4572 , y4573 , y4574 , y4575 , y4576 , y4577 , y4578 , y4579 , y4580 , y4581 , y4582 , y4583 , y4584 , y4585 , y4586 , y4587 , y4588 , y4589 , y4590 , y4591 , y4592 , y4593 , y4594 , y4595 , y4596 , y4597 , y4598 , y4599 , y4600 , y4601 , y4602 , y4603 , y4604 , y4605 , y4606 , y4607 , y4608 , y4609 , y4610 , y4611 , y4612 , y4613 , y4614 , y4615 , y4616 , y4617 , y4618 , y4619 , y4620 , y4621 , y4622 , y4623 , y4624 , y4625 , y4626 , y4627 , y4628 , y4629 , y4630 , y4631 , y4632 , y4633 , y4634 , y4635 , y4636 , y4637 , y4638 , y4639 , y4640 , y4641 , y4642 , y4643 , y4644 , y4645 , y4646 , y4647 , y4648 , y4649 , y4650 , y4651 , y4652 , y4653 , y4654 , y4655 , y4656 , y4657 , y4658 , y4659 , y4660 , y4661 , y4662 , y4663 , y4664 , y4665 , y4666 , y4667 , y4668 , y4669 , y4670 , y4671 , y4672 , y4673 , y4674 , y4675 , y4676 , y4677 , y4678 , y4679 , y4680 , y4681 , y4682 , y4683 , y4684 , y4685 , y4686 , y4687 , y4688 , y4689 , y4690 , y4691 , y4692 , y4693 , y4694 , y4695 , y4696 , y4697 , y4698 , y4699 , y4700 , y4701 , y4702 , y4703 , y4704 , y4705 , y4706 , y4707 , y4708 , y4709 , y4710 , y4711 , y4712 , y4713 , y4714 , y4715 , y4716 , y4717 , y4718 , y4719 , y4720 , y4721 , y4722 , y4723 , y4724 , y4725 , y4726 , y4727 , y4728 , y4729 , y4730 , y4731 , y4732 , y4733 , y4734 , y4735 , y4736 , y4737 , y4738 , y4739 , y4740 , y4741 , y4742 , y4743 , y4744 , y4745 , y4746 , y4747 , y4748 , y4749 , y4750 , y4751 , y4752 , y4753 , y4754 , y4755 , y4756 , y4757 , y4758 , y4759 , y4760 , y4761 , y4762 , y4763 , y4764 , y4765 , y4766 , y4767 , y4768 , y4769 , y4770 , y4771 , y4772 , y4773 , y4774 , y4775 , y4776 , y4777 , y4778 , y4779 , y4780 , y4781 , y4782 , y4783 , y4784 , y4785 , y4786 , y4787 , y4788 , y4789 , y4790 , y4791 , y4792 , y4793 , y4794 , y4795 , y4796 , y4797 , y4798 , y4799 , y4800 , y4801 , y4802 , y4803 , y4804 , y4805 , y4806 , y4807 , y4808 , y4809 , y4810 , y4811 , y4812 , y4813 , y4814 , y4815 , y4816 , y4817 , y4818 , y4819 , y4820 , y4821 , y4822 , y4823 , y4824 , y4825 , y4826 , y4827 , y4828 , y4829 , y4830 , y4831 , y4832 , y4833 , y4834 , y4835 , y4836 , y4837 , y4838 , y4839 , y4840 , y4841 , y4842 , y4843 , y4844 , y4845 , y4846 , y4847 , y4848 , y4849 , y4850 , y4851 , y4852 , y4853 , y4854 , y4855 , y4856 , y4857 , y4858 , y4859 , y4860 , y4861 , y4862 , y4863 , y4864 , y4865 , y4866 , y4867 , y4868 , y4869 , y4870 , y4871 , y4872 , y4873 , y4874 , y4875 , y4876 , y4877 , y4878 , y4879 , y4880 , y4881 , y4882 , y4883 , y4884 , y4885 , y4886 , y4887 , y4888 , y4889 , y4890 , y4891 , y4892 , y4893 , y4894 , y4895 , y4896 , y4897 , y4898 , y4899 , y4900 , y4901 , y4902 , y4903 , y4904 , y4905 , y4906 , y4907 , y4908 , y4909 , y4910 , y4911 , y4912 , y4913 , y4914 , y4915 , y4916 , y4917 , y4918 , y4919 , y4920 , y4921 , y4922 , y4923 , y4924 , y4925 , y4926 , y4927 , y4928 , y4929 , y4930 , y4931 , y4932 , y4933 , y4934 , y4935 , y4936 , y4937 , y4938 , y4939 , y4940 , y4941 , y4942 , y4943 , y4944 , y4945 , y4946 , y4947 , y4948 , y4949 , y4950 , y4951 , y4952 , y4953 , y4954 , y4955 , y4956 , y4957 , y4958 , y4959 , y4960 , y4961 , y4962 , y4963 , y4964 , y4965 , y4966 , y4967 , y4968 , y4969 , y4970 , y4971 , y4972 , y4973 , y4974 , y4975 , y4976 , y4977 , y4978 , y4979 , y4980 , y4981 , y4982 , y4983 , y4984 , y4985 , y4986 , y4987 , y4988 , y4989 , y4990 , y4991 , y4992 , y4993 , y4994 , y4995 , y4996 , y4997 , y4998 , y4999 , y5000 , y5001 , y5002 , y5003 , y5004 , y5005 , y5006 , y5007 , y5008 , y5009 , y5010 , y5011 , y5012 , y5013 , y5014 , y5015 , y5016 , y5017 , y5018 , y5019 , y5020 , y5021 , y5022 , y5023 , y5024 , y5025 , y5026 , y5027 , y5028 , y5029 , y5030 , y5031 , y5032 , y5033 , y5034 , y5035 , y5036 , y5037 , y5038 , y5039 , y5040 , y5041 , y5042 , y5043 , y5044 , y5045 , y5046 , y5047 , y5048 , y5049 , y5050 , y5051 , y5052 , y5053 , y5054 , y5055 , y5056 , y5057 , y5058 , y5059 , y5060 , y5061 , y5062 , y5063 , y5064 , y5065 , y5066 , y5067 , y5068 , y5069 , y5070 , y5071 , y5072 , y5073 , y5074 , y5075 , y5076 , y5077 , y5078 , y5079 , y5080 , y5081 , y5082 , y5083 , y5084 , y5085 , y5086 , y5087 , y5088 , y5089 , y5090 , y5091 , y5092 , y5093 , y5094 , y5095 , y5096 , y5097 , y5098 , y5099 , y5100 , y5101 , y5102 , y5103 , y5104 , y5105 , y5106 , y5107 , y5108 , y5109 , y5110 , y5111 , y5112 , y5113 , y5114 , y5115 , y5116 , y5117 , y5118 , y5119 , y5120 , y5121 , y5122 , y5123 , y5124 , y5125 , y5126 , y5127 , y5128 , y5129 , y5130 , y5131 , y5132 , y5133 , y5134 , y5135 , y5136 , y5137 , y5138 , y5139 , y5140 , y5141 , y5142 , y5143 , y5144 , y5145 , y5146 , y5147 , y5148 , y5149 , y5150 , y5151 , y5152 , y5153 , y5154 , y5155 , y5156 , y5157 , y5158 , y5159 , y5160 , y5161 , y5162 , y5163 , y5164 , y5165 , y5166 , y5167 , y5168 , y5169 , y5170 , y5171 , y5172 , y5173 , y5174 , y5175 , y5176 , y5177 , y5178 , y5179 , y5180 , y5181 , y5182 , y5183 , y5184 , y5185 , y5186 , y5187 , y5188 , y5189 , y5190 , y5191 , y5192 , y5193 , y5194 , y5195 , y5196 , y5197 , y5198 , y5199 , y5200 , y5201 , y5202 , y5203 , y5204 , y5205 , y5206 , y5207 , y5208 , y5209 , y5210 , y5211 , y5212 , y5213 , y5214 , y5215 , y5216 , y5217 , y5218 , y5219 , y5220 , y5221 , y5222 , y5223 , y5224 , y5225 , y5226 , y5227 , y5228 , y5229 , y5230 , y5231 , y5232 , y5233 , y5234 , y5235 , y5236 , y5237 , y5238 , y5239 , y5240 , y5241 , y5242 , y5243 , y5244 , y5245 , y5246 , y5247 , y5248 , y5249 , y5250 , y5251 , y5252 , y5253 , y5254 , y5255 , y5256 , y5257 , y5258 , y5259 , y5260 , y5261 , y5262 , y5263 , y5264 , y5265 , y5266 , y5267 , y5268 , y5269 , y5270 , y5271 , y5272 , y5273 , y5274 , y5275 , y5276 , y5277 , y5278 , y5279 , y5280 , y5281 , y5282 , y5283 , y5284 , y5285 , y5286 , y5287 , y5288 , y5289 , y5290 , y5291 , y5292 , y5293 , y5294 , y5295 , y5296 , y5297 , y5298 , y5299 , y5300 , y5301 , y5302 , y5303 , y5304 , y5305 , y5306 , y5307 , y5308 , y5309 , y5310 , y5311 , y5312 , y5313 , y5314 , y5315 , y5316 , y5317 , y5318 , y5319 , y5320 , y5321 , y5322 , y5323 , y5324 , y5325 , y5326 , y5327 , y5328 , y5329 , y5330 , y5331 , y5332 , y5333 , y5334 , y5335 , y5336 , y5337 , y5338 , y5339 , y5340 , y5341 , y5342 , y5343 , y5344 , y5345 , y5346 , y5347 , y5348 , y5349 , y5350 , y5351 , y5352 , y5353 , y5354 , y5355 , y5356 , y5357 , y5358 , y5359 , y5360 , y5361 , y5362 , y5363 , y5364 , y5365 , y5366 , y5367 , y5368 , y5369 , y5370 , y5371 , y5372 , y5373 , y5374 , y5375 , y5376 , y5377 , y5378 , y5379 , y5380 , y5381 , y5382 , y5383 , y5384 , y5385 , y5386 , y5387 , y5388 , y5389 , y5390 , y5391 , y5392 , y5393 , y5394 , y5395 , y5396 , y5397 , y5398 , y5399 , y5400 , y5401 , y5402 , y5403 , y5404 , y5405 , y5406 , y5407 , y5408 , y5409 , y5410 , y5411 , y5412 , y5413 , y5414 , y5415 , y5416 , y5417 , y5418 , y5419 , y5420 , y5421 , y5422 , y5423 , y5424 , y5425 , y5426 , y5427 , y5428 , y5429 , y5430 , y5431 , y5432 , y5433 , y5434 , y5435 , y5436 , y5437 , y5438 , y5439 , y5440 , y5441 , y5442 , y5443 , y5444 , y5445 , y5446 , y5447 , y5448 , y5449 , y5450 , y5451 , y5452 , y5453 , y5454 , y5455 , y5456 , y5457 , y5458 , y5459 , y5460 , y5461 , y5462 , y5463 , y5464 , y5465 , y5466 , y5467 , y5468 , y5469 , y5470 , y5471 , y5472 , y5473 , y5474 , y5475 , y5476 , y5477 , y5478 , y5479 , y5480 , y5481 , y5482 , y5483 , y5484 , y5485 , y5486 , y5487 , y5488 , y5489 , y5490 , y5491 , y5492 , y5493 , y5494 , y5495 , y5496 , y5497 , y5498 , y5499 , y5500 , y5501 , y5502 , y5503 , y5504 , y5505 , y5506 , y5507 , y5508 , y5509 , y5510 , y5511 , y5512 , y5513 , y5514 , y5515 , y5516 , y5517 , y5518 , y5519 , y5520 , y5521 , y5522 , y5523 , y5524 , y5525 , y5526 , y5527 , y5528 , y5529 , y5530 , y5531 , y5532 , y5533 , y5534 , y5535 , y5536 , y5537 , y5538 , y5539 , y5540 , y5541 , y5542 , y5543 , y5544 , y5545 , y5546 , y5547 , y5548 , y5549 , y5550 , y5551 , y5552 , y5553 , y5554 , y5555 , y5556 , y5557 , y5558 , y5559 , y5560 , y5561 , y5562 , y5563 , y5564 , y5565 , y5566 , y5567 , y5568 , y5569 , y5570 , y5571 , y5572 , y5573 , y5574 , y5575 , y5576 , y5577 , y5578 , y5579 , y5580 , y5581 , y5582 , y5583 , y5584 , y5585 , y5586 , y5587 , y5588 , y5589 , y5590 , y5591 , y5592 , y5593 , y5594 , y5595 , y5596 , y5597 , y5598 , y5599 , y5600 , y5601 , y5602 , y5603 , y5604 , y5605 , y5606 , y5607 , y5608 , y5609 , y5610 , y5611 , y5612 , y5613 , y5614 , y5615 , y5616 , y5617 , y5618 , y5619 , y5620 , y5621 , y5622 , y5623 , y5624 , y5625 , y5626 , y5627 , y5628 , y5629 , y5630 , y5631 , y5632 , y5633 , y5634 , y5635 , y5636 , y5637 , y5638 , y5639 , y5640 , y5641 , y5642 , y5643 , y5644 , y5645 , y5646 , y5647 , y5648 , y5649 , y5650 , y5651 , y5652 , y5653 , y5654 , y5655 , y5656 , y5657 , y5658 , y5659 , y5660 , y5661 , y5662 , y5663 , y5664 , y5665 , y5666 , y5667 , y5668 , y5669 , y5670 , y5671 , y5672 , y5673 , y5674 , y5675 , y5676 , y5677 , y5678 , y5679 , y5680 , y5681 , y5682 , y5683 , y5684 , y5685 , y5686 , y5687 , y5688 , y5689 , y5690 , y5691 , y5692 , y5693 , y5694 , y5695 , y5696 , y5697 , y5698 , y5699 , y5700 , y5701 , y5702 , y5703 , y5704 , y5705 , y5706 , y5707 , y5708 , y5709 , y5710 , y5711 , y5712 , y5713 , y5714 , y5715 , y5716 , y5717 , y5718 , y5719 , y5720 , y5721 , y5722 , y5723 , y5724 , y5725 , y5726 , y5727 , y5728 , y5729 , y5730 , y5731 , y5732 , y5733 , y5734 , y5735 , y5736 , y5737 , y5738 , y5739 , y5740 , y5741 , y5742 , y5743 , y5744 , y5745 , y5746 , y5747 , y5748 , y5749 , y5750 , y5751 , y5752 , y5753 , y5754 , y5755 , y5756 , y5757 , y5758 , y5759 , y5760 , y5761 , y5762 , y5763 , y5764 , y5765 , y5766 , y5767 , y5768 , y5769 , y5770 , y5771 , y5772 , y5773 , y5774 , y5775 , y5776 , y5777 , y5778 , y5779 , y5780 , y5781 , y5782 , y5783 , y5784 , y5785 , y5786 , y5787 , y5788 , y5789 , y5790 , y5791 , y5792 , y5793 , y5794 , y5795 , y5796 , y5797 , y5798 , y5799 , y5800 , y5801 , y5802 , y5803 , y5804 , y5805 , y5806 , y5807 , y5808 , y5809 , y5810 , y5811 , y5812 , y5813 , y5814 , y5815 , y5816 , y5817 , y5818 , y5819 , y5820 , y5821 , y5822 , y5823 , y5824 , y5825 , y5826 , y5827 , y5828 , y5829 , y5830 , y5831 , y5832 , y5833 , y5834 , y5835 , y5836 , y5837 , y5838 , y5839 , y5840 , y5841 , y5842 , y5843 , y5844 , y5845 , y5846 , y5847 , y5848 , y5849 , y5850 , y5851 , y5852 , y5853 , y5854 , y5855 , y5856 , y5857 , y5858 , y5859 , y5860 , y5861 , y5862 , y5863 , y5864 , y5865 , y5866 , y5867 , y5868 , y5869 , y5870 , y5871 , y5872 , y5873 , y5874 , y5875 , y5876 , y5877 , y5878 , y5879 , y5880 , y5881 , y5882 , y5883 , y5884 , y5885 , y5886 , y5887 , y5888 , y5889 , y5890 , y5891 , y5892 , y5893 , y5894 , y5895 , y5896 , y5897 , y5898 , y5899 , y5900 , y5901 , y5902 , y5903 , y5904 , y5905 , y5906 , y5907 , y5908 , y5909 , y5910 , y5911 , y5912 , y5913 , y5914 , y5915 , y5916 , y5917 , y5918 , y5919 , y5920 , y5921 , y5922 , y5923 , y5924 , y5925 , y5926 , y5927 , y5928 , y5929 , y5930 , y5931 , y5932 , y5933 , y5934 , y5935 , y5936 , y5937 , y5938 , y5939 , y5940 , y5941 , y5942 , y5943 , y5944 , y5945 , y5946 , y5947 , y5948 , y5949 , y5950 , y5951 , y5952 , y5953 , y5954 , y5955 , y5956 , y5957 , y5958 , y5959 , y5960 , y5961 , y5962 , y5963 , y5964 , y5965 , y5966 , y5967 , y5968 , y5969 , y5970 , y5971 , y5972 , y5973 , y5974 , y5975 , y5976 , y5977 , y5978 , y5979 , y5980 , y5981 , y5982 , y5983 , y5984 , y5985 , y5986 , y5987 , y5988 , y5989 , y5990 , y5991 , y5992 , y5993 , y5994 , y5995 , y5996 , y5997 , y5998 , y5999 , y6000 , y6001 , y6002 , y6003 , y6004 , y6005 , y6006 , y6007 , y6008 , y6009 , y6010 , y6011 , y6012 , y6013 , y6014 , y6015 , y6016 , y6017 , y6018 , y6019 , y6020 , y6021 , y6022 , y6023 , y6024 , y6025 , y6026 , y6027 , y6028 , y6029 , y6030 , y6031 , y6032 , y6033 , y6034 , y6035 , y6036 , y6037 , y6038 , y6039 , y6040 , y6041 , y6042 , y6043 , y6044 , y6045 , y6046 , y6047 , y6048 , y6049 , y6050 , y6051 , y6052 , y6053 , y6054 , y6055 , y6056 , y6057 , y6058 , y6059 , y6060 , y6061 , y6062 , y6063 , y6064 , y6065 , y6066 , y6067 , y6068 , y6069 , y6070 , y6071 , y6072 , y6073 , y6074 , y6075 , y6076 , y6077 , y6078 , y6079 , y6080 , y6081 , y6082 , y6083 , y6084 , y6085 , y6086 , y6087 , y6088 , y6089 , y6090 , y6091 , y6092 , y6093 , y6094 , y6095 , y6096 , y6097 , y6098 , y6099 , y6100 , y6101 , y6102 , y6103 , y6104 , y6105 , y6106 , y6107 , y6108 , y6109 , y6110 , y6111 , y6112 , y6113 , y6114 , y6115 , y6116 , y6117 , y6118 , y6119 , y6120 , y6121 , y6122 , y6123 , y6124 , y6125 , y6126 , y6127 , y6128 , y6129 , y6130 , y6131 , y6132 , y6133 , y6134 , y6135 , y6136 , y6137 , y6138 , y6139 , y6140 , y6141 , y6142 , y6143 , y6144 , y6145 , y6146 , y6147 , y6148 , y6149 , y6150 , y6151 , y6152 , y6153 , y6154 , y6155 , y6156 , y6157 , y6158 , y6159 , y6160 , y6161 , y6162 , y6163 , y6164 , y6165 , y6166 , y6167 , y6168 , y6169 , y6170 , y6171 , y6172 , y6173 , y6174 , y6175 , y6176 , y6177 , y6178 , y6179 , y6180 , y6181 , y6182 , y6183 , y6184 , y6185 , y6186 , y6187 , y6188 , y6189 , y6190 , y6191 , y6192 , y6193 , y6194 , y6195 , y6196 , y6197 , y6198 , y6199 , y6200 , y6201 , y6202 , y6203 , y6204 , y6205 , y6206 , y6207 , y6208 , y6209 , y6210 , y6211 , y6212 , y6213 , y6214 , y6215 , y6216 , y6217 , y6218 , y6219 , y6220 , y6221 , y6222 , y6223 , y6224 , y6225 , y6226 , y6227 , y6228 , y6229 , y6230 , y6231 , y6232 , y6233 , y6234 , y6235 , y6236 , y6237 , y6238 , y6239 , y6240 , y6241 , y6242 , y6243 , y6244 , y6245 , y6246 , y6247 , y6248 , y6249 , y6250 , y6251 , y6252 , y6253 , y6254 , y6255 , y6256 , y6257 , y6258 , y6259 , y6260 , y6261 , y6262 , y6263 , y6264 , y6265 , y6266 , y6267 , y6268 , y6269 , y6270 , y6271 , y6272 , y6273 , y6274 , y6275 , y6276 , y6277 , y6278 , y6279 , y6280 , y6281 , y6282 , y6283 , y6284 , y6285 , y6286 , y6287 , y6288 , y6289 , y6290 , y6291 , y6292 , y6293 , y6294 , y6295 , y6296 , y6297 , y6298 , y6299 , y6300 , y6301 , y6302 , y6303 , y6304 , y6305 , y6306 , y6307 , y6308 , y6309 , y6310 , y6311 , y6312 , y6313 , y6314 , y6315 , y6316 , y6317 , y6318 , y6319 , y6320 , y6321 , y6322 , y6323 , y6324 , y6325 , y6326 , y6327 , y6328 , y6329 , y6330 , y6331 , y6332 , y6333 , y6334 , y6335 , y6336 , y6337 , y6338 , y6339 , y6340 , y6341 , y6342 , y6343 , y6344 , y6345 , y6346 , y6347 , y6348 , y6349 , y6350 , y6351 , y6352 , y6353 , y6354 , y6355 , y6356 , y6357 , y6358 , y6359 , y6360 , y6361 , y6362 , y6363 , y6364 , y6365 , y6366 , y6367 , y6368 , y6369 , y6370 , y6371 , y6372 , y6373 , y6374 , y6375 , y6376 , y6377 , y6378 , y6379 , y6380 , y6381 , y6382 , y6383 , y6384 , y6385 , y6386 , y6387 , y6388 , y6389 , y6390 , y6391 , y6392 , y6393 , y6394 , y6395 , y6396 , y6397 , y6398 , y6399 , y6400 , y6401 , y6402 , y6403 , y6404 , y6405 , y6406 , y6407 , y6408 , y6409 , y6410 , y6411 , y6412 , y6413 , y6414 , y6415 , y6416 , y6417 , y6418 , y6419 , y6420 , y6421 , y6422 , y6423 , y6424 , y6425 , y6426 , y6427 , y6428 , y6429 , y6430 , y6431 , y6432 , y6433 , y6434 , y6435 , y6436 , y6437 , y6438 , y6439 , y6440 , y6441 , y6442 , y6443 , y6444 , y6445 , y6446 , y6447 , y6448 , y6449 , y6450 , y6451 , y6452 , y6453 , y6454 , y6455 , y6456 , y6457 , y6458 , y6459 , y6460 , y6461 , y6462 , y6463 , y6464 , y6465 , y6466 , y6467 , y6468 , y6469 , y6470 , y6471 , y6472 , y6473 , y6474 , y6475 , y6476 , y6477 , y6478 , y6479 , y6480 , y6481 , y6482 , y6483 , y6484 , y6485 , y6486 , y6487 , y6488 , y6489 , y6490 , y6491 , y6492 , y6493 , y6494 , y6495 , y6496 , y6497 , y6498 , y6499 , y6500 , y6501 , y6502 , y6503 , y6504 , y6505 , y6506 , y6507 , y6508 , y6509 , y6510 , y6511 , y6512 , y6513 , y6514 , y6515 , y6516 , y6517 , y6518 , y6519 , y6520 , y6521 , y6522 , y6523 , y6524 , y6525 , y6526 , y6527 , y6528 , y6529 , y6530 , y6531 , y6532 , y6533 , y6534 , y6535 , y6536 , y6537 , y6538 , y6539 , y6540 , y6541 , y6542 , y6543 , y6544 , y6545 , y6546 , y6547 , y6548 , y6549 , y6550 , y6551 , y6552 , y6553 , y6554 , y6555 , y6556 , y6557 , y6558 , y6559 , y6560 , y6561 , y6562 , y6563 , y6564 , y6565 , y6566 , y6567 , y6568 , y6569 , y6570 , y6571 , y6572 , y6573 , y6574 , y6575 , y6576 , y6577 , y6578 , y6579 , y6580 , y6581 , y6582 , y6583 , y6584 , y6585 , y6586 , y6587 , y6588 , y6589 , y6590 , y6591 , y6592 , y6593 , y6594 , y6595 , y6596 , y6597 , y6598 , y6599 , y6600 , y6601 , y6602 , y6603 , y6604 , y6605 , y6606 , y6607 , y6608 , y6609 , y6610 , y6611 , y6612 , y6613 , y6614 , y6615 , y6616 , y6617 , y6618 , y6619 , y6620 , y6621 , y6622 , y6623 , y6624 , y6625 , y6626 , y6627 , y6628 , y6629 , y6630 , y6631 , y6632 , y6633 , y6634 , y6635 , y6636 , y6637 , y6638 , y6639 , y6640 , y6641 , y6642 , y6643 , y6644 , y6645 , y6646 , y6647 , y6648 , y6649 , y6650 , y6651 , y6652 , y6653 , y6654 , y6655 , y6656 , y6657 , y6658 , y6659 , y6660 , y6661 , y6662 , y6663 , y6664 , y6665 , y6666 , y6667 , y6668 , y6669 , y6670 , y6671 , y6672 , y6673 , y6674 , y6675 , y6676 , y6677 , y6678 , y6679 , y6680 , y6681 , y6682 , y6683 , y6684 , y6685 , y6686 , y6687 , y6688 , y6689 , y6690 , y6691 , y6692 , y6693 , y6694 , y6695 , y6696 , y6697 , y6698 , y6699 , y6700 , y6701 , y6702 , y6703 , y6704 , y6705 , y6706 , y6707 , y6708 , y6709 , y6710 , y6711 , y6712 , y6713 , y6714 , y6715 , y6716 , y6717 , y6718 , y6719 , y6720 , y6721 , y6722 , y6723 , y6724 , y6725 , y6726 , y6727 , y6728 , y6729 , y6730 , y6731 , y6732 , y6733 , y6734 , y6735 , y6736 , y6737 , y6738 , y6739 , y6740 , y6741 , y6742 , y6743 , y6744 , y6745 , y6746 , y6747 , y6748 , y6749 , y6750 , y6751 , y6752 , y6753 , y6754 , y6755 , y6756 , y6757 , y6758 , y6759 , y6760 , y6761 , y6762 , y6763 , y6764 , y6765 , y6766 , y6767 , y6768 , y6769 , y6770 , y6771 , y6772 , y6773 , y6774 , y6775 , y6776 , y6777 , y6778 , y6779 , y6780 , y6781 , y6782 , y6783 , y6784 , y6785 , y6786 , y6787 , y6788 , y6789 , y6790 , y6791 , y6792 , y6793 , y6794 , y6795 , y6796 , y6797 , y6798 , y6799 , y6800 , y6801 , y6802 , y6803 , y6804 , y6805 , y6806 , y6807 , y6808 , y6809 , y6810 , y6811 , y6812 , y6813 , y6814 , y6815 , y6816 , y6817 , y6818 , y6819 , y6820 , y6821 , y6822 , y6823 , y6824 , y6825 , y6826 , y6827 , y6828 , y6829 , y6830 , y6831 , y6832 , y6833 , y6834 , y6835 , y6836 , y6837 , y6838 , y6839 , y6840 , y6841 , y6842 , y6843 , y6844 , y6845 , y6846 , y6847 , y6848 , y6849 , y6850 , y6851 , y6852 , y6853 , y6854 , y6855 , y6856 , y6857 , y6858 , y6859 , y6860 , y6861 , y6862 , y6863 , y6864 , y6865 , y6866 , y6867 , y6868 , y6869 , y6870 , y6871 , y6872 , y6873 , y6874 , y6875 , y6876 , y6877 , y6878 , y6879 , y6880 , y6881 , y6882 , y6883 , y6884 , y6885 , y6886 , y6887 , y6888 , y6889 , y6890 , y6891 , y6892 , y6893 , y6894 , y6895 , y6896 , y6897 , y6898 , y6899 , y6900 , y6901 , y6902 , y6903 , y6904 , y6905 , y6906 , y6907 , y6908 , y6909 , y6910 , y6911 , y6912 , y6913 , y6914 , y6915 , y6916 , y6917 , y6918 , y6919 , y6920 , y6921 , y6922 , y6923 , y6924 , y6925 , y6926 , y6927 , y6928 , y6929 , y6930 , y6931 , y6932 , y6933 , y6934 , y6935 , y6936 , y6937 , y6938 , y6939 , y6940 , y6941 , y6942 , y6943 , y6944 , y6945 , y6946 , y6947 , y6948 , y6949 , y6950 , y6951 , y6952 , y6953 , y6954 , y6955 , y6956 , y6957 , y6958 , y6959 , y6960 , y6961 , y6962 , y6963 , y6964 , y6965 , y6966 , y6967 , y6968 , y6969 , y6970 , y6971 , y6972 , y6973 , y6974 , y6975 , y6976 , y6977 , y6978 , y6979 , y6980 , y6981 , y6982 , y6983 , y6984 , y6985 , y6986 , y6987 , y6988 , y6989 , y6990 , y6991 , y6992 , y6993 , y6994 , y6995 , y6996 , y6997 , y6998 , y6999 , y7000 , y7001 , y7002 , y7003 , y7004 , y7005 , y7006 , y7007 , y7008 , y7009 , y7010 , y7011 , y7012 , y7013 , y7014 , y7015 , y7016 , y7017 , y7018 , y7019 , y7020 , y7021 , y7022 , y7023 , y7024 , y7025 , y7026 , y7027 , y7028 , y7029 , y7030 , y7031 , y7032 , y7033 , y7034 , y7035 , y7036 , y7037 , y7038 , y7039 , y7040 , y7041 , y7042 , y7043 , y7044 , y7045 , y7046 , y7047 , y7048 , y7049 , y7050 , y7051 , y7052 , y7053 , y7054 , y7055 , y7056 , y7057 , y7058 , y7059 , y7060 , y7061 , y7062 , y7063 , y7064 , y7065 , y7066 , y7067 , y7068 , y7069 , y7070 , y7071 , y7072 , y7073 , y7074 , y7075 , y7076 , y7077 , y7078 , y7079 , y7080 , y7081 , y7082 , y7083 , y7084 , y7085 , y7086 , y7087 , y7088 , y7089 , y7090 , y7091 , y7092 , y7093 , y7094 , y7095 , y7096 , y7097 , y7098 , y7099 , y7100 , y7101 , y7102 , y7103 , y7104 , y7105 , y7106 , y7107 , y7108 , y7109 , y7110 , y7111 , y7112 , y7113 , y7114 , y7115 , y7116 , y7117 , y7118 , y7119 , y7120 , y7121 , y7122 , y7123 , y7124 , y7125 , y7126 , y7127 , y7128 , y7129 , y7130 , y7131 , y7132 , y7133 , y7134 , y7135 , y7136 , y7137 , y7138 , y7139 , y7140 , y7141 , y7142 , y7143 , y7144 , y7145 , y7146 , y7147 , y7148 , y7149 , y7150 , y7151 , y7152 , y7153 , y7154 , y7155 , y7156 , y7157 , y7158 , y7159 , y7160 , y7161 , y7162 , y7163 , y7164 , y7165 , y7166 , y7167 , y7168 , y7169 , y7170 , y7171 , y7172 , y7173 , y7174 , y7175 , y7176 , y7177 , y7178 , y7179 , y7180 , y7181 , y7182 , y7183 , y7184 , y7185 , y7186 , y7187 , y7188 , y7189 , y7190 , y7191 , y7192 , y7193 , y7194 , y7195 , y7196 , y7197 , y7198 , y7199 , y7200 , y7201 , y7202 , y7203 , y7204 , y7205 , y7206 , y7207 , y7208 , y7209 , y7210 , y7211 , y7212 , y7213 , y7214 , y7215 , y7216 , y7217 , y7218 , y7219 , y7220 , y7221 , y7222 , y7223 , y7224 , y7225 , y7226 , y7227 , y7228 , y7229 , y7230 , y7231 , y7232 , y7233 , y7234 , y7235 , y7236 , y7237 , y7238 , y7239 , y7240 , y7241 , y7242 , y7243 , y7244 , y7245 , y7246 , y7247 , y7248 , y7249 , y7250 , y7251 , y7252 , y7253 , y7254 , y7255 , y7256 , y7257 , y7258 , y7259 , y7260 , y7261 , y7262 , y7263 , y7264 , y7265 , y7266 , y7267 , y7268 , y7269 , y7270 , y7271 , y7272 , y7273 , y7274 , y7275 , y7276 , y7277 , y7278 , y7279 , y7280 , y7281 , y7282 , y7283 , y7284 , y7285 , y7286 , y7287 , y7288 , y7289 , y7290 , y7291 , y7292 , y7293 , y7294 , y7295 , y7296 , y7297 , y7298 , y7299 , y7300 , y7301 , y7302 , y7303 , y7304 , y7305 , y7306 , y7307 , y7308 , y7309 , y7310 , y7311 , y7312 , y7313 , y7314 , y7315 , y7316 , y7317 , y7318 , y7319 , y7320 , y7321 , y7322 , y7323 , y7324 , y7325 , y7326 , y7327 , y7328 , y7329 , y7330 , y7331 , y7332 , y7333 , y7334 , y7335 , y7336 , y7337 , y7338 , y7339 , y7340 , y7341 , y7342 , y7343 , y7344 , y7345 , y7346 , y7347 , y7348 , y7349 , y7350 , y7351 , y7352 , y7353 , y7354 , y7355 , y7356 , y7357 , y7358 , y7359 , y7360 , y7361 , y7362 , y7363 , y7364 , y7365 , y7366 , y7367 , y7368 , y7369 , y7370 , y7371 , y7372 , y7373 , y7374 , y7375 , y7376 , y7377 , y7378 , y7379 , y7380 , y7381 , y7382 , y7383 , y7384 , y7385 , y7386 , y7387 , y7388 , y7389 , y7390 , y7391 , y7392 , y7393 , y7394 , y7395 , y7396 , y7397 , y7398 , y7399 , y7400 , y7401 , y7402 , y7403 , y7404 , y7405 , y7406 , y7407 , y7408 , y7409 , y7410 , y7411 , y7412 , y7413 , y7414 , y7415 , y7416 , y7417 , y7418 , y7419 , y7420 , y7421 , y7422 , y7423 , y7424 , y7425 , y7426 , y7427 , y7428 , y7429 , y7430 , y7431 , y7432 , y7433 , y7434 , y7435 , y7436 , y7437 , y7438 , y7439 , y7440 , y7441 , y7442 , y7443 , y7444 , y7445 , y7446 , y7447 , y7448 , y7449 , y7450 , y7451 , y7452 , y7453 , y7454 , y7455 , y7456 , y7457 , y7458 , y7459 , y7460 , y7461 , y7462 , y7463 , y7464 , y7465 , y7466 , y7467 , y7468 , y7469 , y7470 , y7471 , y7472 , y7473 , y7474 , y7475 , y7476 , y7477 , y7478 , y7479 , y7480 , y7481 , y7482 , y7483 , y7484 , y7485 , y7486 , y7487 , y7488 , y7489 , y7490 , y7491 , y7492 , y7493 , y7494 , y7495 , y7496 , y7497 , y7498 , y7499 , y7500 , y7501 , y7502 , y7503 , y7504 , y7505 , y7506 , y7507 , y7508 , y7509 , y7510 , y7511 , y7512 , y7513 , y7514 , y7515 , y7516 , y7517 , y7518 , y7519 , y7520 , y7521 , y7522 , y7523 , y7524 , y7525 , y7526 , y7527 , y7528 , y7529 , y7530 , y7531 , y7532 , y7533 , y7534 , y7535 , y7536 , y7537 , y7538 , y7539 , y7540 , y7541 , y7542 , y7543 , y7544 , y7545 , y7546 , y7547 , y7548 , y7549 , y7550 , y7551 , y7552 , y7553 , y7554 , y7555 , y7556 , y7557 , y7558 , y7559 , y7560 , y7561 , y7562 , y7563 , y7564 , y7565 , y7566 , y7567 , y7568 , y7569 , y7570 , y7571 , y7572 , y7573 , y7574 , y7575 , y7576 , y7577 , y7578 , y7579 , y7580 , y7581 , y7582 , y7583 , y7584 , y7585 , y7586 , y7587 , y7588 , y7589 , y7590 , y7591 , y7592 , y7593 , y7594 , y7595 , y7596 , y7597 , y7598 , y7599 , y7600 , y7601 , y7602 , y7603 , y7604 , y7605 , y7606 , y7607 , y7608 , y7609 , y7610 , y7611 , y7612 , y7613 , y7614 , y7615 , y7616 , y7617 , y7618 , y7619 , y7620 , y7621 , y7622 , y7623 , y7624 , y7625 , y7626 , y7627 , y7628 , y7629 , y7630 , y7631 , y7632 , y7633 , y7634 , y7635 , y7636 , y7637 , y7638 , y7639 , y7640 , y7641 , y7642 , y7643 , y7644 , y7645 , y7646 , y7647 , y7648 , y7649 , y7650 , y7651 , y7652 , y7653 , y7654 , y7655 , y7656 , y7657 , y7658 , y7659 , y7660 , y7661 , y7662 , y7663 , y7664 , y7665 , y7666 , y7667 , y7668 , y7669 , y7670 , y7671 , y7672 , y7673 , y7674 , y7675 , y7676 , y7677 , y7678 , y7679 , y7680 , y7681 , y7682 , y7683 , y7684 , y7685 , y7686 , y7687 , y7688 , y7689 , y7690 , y7691 , y7692 , y7693 , y7694 , y7695 , y7696 , y7697 , y7698 , y7699 , y7700 , y7701 , y7702 , y7703 , y7704 , y7705 , y7706 , y7707 , y7708 , y7709 , y7710 , y7711 , y7712 , y7713 , y7714 , y7715 , y7716 , y7717 , y7718 , y7719 , y7720 , y7721 , y7722 , y7723 , y7724 , y7725 , y7726 , y7727 , y7728 , y7729 , y7730 , y7731 , y7732 , y7733 , y7734 , y7735 , y7736 , y7737 , y7738 , y7739 , y7740 , y7741 , y7742 , y7743 , y7744 , y7745 , y7746 , y7747 , y7748 , y7749 , y7750 , y7751 , y7752 , y7753 , y7754 , y7755 , y7756 , y7757 , y7758 , y7759 , y7760 , y7761 , y7762 , y7763 , y7764 , y7765 , y7766 , y7767 , y7768 , y7769 , y7770 , y7771 , y7772 , y7773 , y7774 , y7775 , y7776 , y7777 , y7778 , y7779 , y7780 , y7781 , y7782 , y7783 , y7784 , y7785 , y7786 , y7787 , y7788 , y7789 , y7790 , y7791 , y7792 , y7793 , y7794 , y7795 , y7796 , y7797 , y7798 , y7799 , y7800 , y7801 , y7802 , y7803 , y7804 , y7805 , y7806 , y7807 , y7808 , y7809 , y7810 , y7811 , y7812 , y7813 , y7814 , y7815 , y7816 , y7817 , y7818 , y7819 , y7820 , y7821 , y7822 , y7823 , y7824 , y7825 , y7826 , y7827 , y7828 , y7829 , y7830 , y7831 , y7832 , y7833 , y7834 , y7835 , y7836 , y7837 , y7838 , y7839 , y7840 , y7841 , y7842 , y7843 , y7844 , y7845 , y7846 , y7847 , y7848 , y7849 , y7850 , y7851 , y7852 , y7853 , y7854 , y7855 , y7856 , y7857 , y7858 , y7859 , y7860 , y7861 , y7862 , y7863 , y7864 , y7865 , y7866 , y7867 , y7868 , y7869 , y7870 , y7871 , y7872 , y7873 , y7874 , y7875 , y7876 , y7877 , y7878 , y7879 , y7880 , y7881 , y7882 , y7883 , y7884 , y7885 , y7886 , y7887 , y7888 , y7889 , y7890 , y7891 , y7892 , y7893 , y7894 , y7895 , y7896 , y7897 , y7898 , y7899 , y7900 , y7901 , y7902 , y7903 , y7904 , y7905 , y7906 , y7907 , y7908 , y7909 , y7910 , y7911 , y7912 , y7913 , y7914 , y7915 , y7916 , y7917 , y7918 , y7919 , y7920 , y7921 , y7922 , y7923 , y7924 , y7925 , y7926 , y7927 , y7928 , y7929 , y7930 , y7931 , y7932 , y7933 , y7934 , y7935 , y7936 , y7937 , y7938 , y7939 , y7940 , y7941 , y7942 , y7943 , y7944 , y7945 , y7946 , y7947 , y7948 , y7949 , y7950 , y7951 , y7952 , y7953 , y7954 , y7955 , y7956 , y7957 , y7958 , y7959 , y7960 , y7961 , y7962 , y7963 , y7964 , y7965 , y7966 , y7967 , y7968 , y7969 , y7970 , y7971 , y7972 , y7973 , y7974 , y7975 , y7976 , y7977 , y7978 , y7979 , y7980 , y7981 , y7982 , y7983 , y7984 , y7985 , y7986 , y7987 , y7988 , y7989 , y7990 , y7991 , y7992 , y7993 , y7994 , y7995 , y7996 , y7997 , y7998 , y7999 , y8000 , y8001 , y8002 , y8003 , y8004 , y8005 , y8006 , y8007 , y8008 , y8009 , y8010 , y8011 , y8012 , y8013 , y8014 , y8015 , y8016 , y8017 , y8018 , y8019 , y8020 , y8021 , y8022 , y8023 , y8024 , y8025 , y8026 , y8027 , y8028 , y8029 , y8030 , y8031 , y8032 , y8033 , y8034 , y8035 , y8036 , y8037 , y8038 , y8039 , y8040 , y8041 , y8042 , y8043 , y8044 , y8045 , y8046 , y8047 , y8048 , y8049 , y8050 , y8051 , y8052 , y8053 , y8054 , y8055 , y8056 , y8057 , y8058 , y8059 , y8060 , y8061 , y8062 , y8063 , y8064 , y8065 , y8066 , y8067 , y8068 , y8069 , y8070 , y8071 , y8072 , y8073 , y8074 , y8075 , y8076 , y8077 , y8078 , y8079 , y8080 , y8081 , y8082 , y8083 , y8084 , y8085 , y8086 , y8087 , y8088 , y8089 , y8090 , y8091 , y8092 , y8093 , y8094 , y8095 , y8096 , y8097 , y8098 , y8099 , y8100 , y8101 , y8102 , y8103 , y8104 , y8105 , y8106 , y8107 , y8108 , y8109 , y8110 , y8111 , y8112 , y8113 , y8114 , y8115 , y8116 , y8117 , y8118 , y8119 , y8120 , y8121 , y8122 , y8123 , y8124 , y8125 , y8126 , y8127 , y8128 , y8129 , y8130 , y8131 , y8132 , y8133 , y8134 , y8135 , y8136 , y8137 , y8138 , y8139 , y8140 , y8141 , y8142 , y8143 , y8144 , y8145 , y8146 , y8147 , y8148 , y8149 , y8150 , y8151 , y8152 , y8153 , y8154 , y8155 , y8156 , y8157 , y8158 , y8159 , y8160 , y8161 , y8162 , y8163 , y8164 , y8165 , y8166 , y8167 , y8168 , y8169 , y8170 , y8171 , y8172 , y8173 , y8174 , y8175 , y8176 , y8177 , y8178 , y8179 , y8180 , y8181 , y8182 , y8183 , y8184 , y8185 , y8186 , y8187 , y8188 , y8189 , y8190 , y8191 , y8192 , y8193 , y8194 , y8195 , y8196 , y8197 , y8198 , y8199 , y8200 , y8201 , y8202 , y8203 , y8204 , y8205 , y8206 , y8207 , y8208 , y8209 , y8210 , y8211 , y8212 , y8213 , y8214 , y8215 , y8216 , y8217 , y8218 , y8219 , y8220 , y8221 , y8222 , y8223 , y8224 , y8225 , y8226 , y8227 , y8228 , y8229 , y8230 , y8231 , y8232 , y8233 , y8234 , y8235 , y8236 , y8237 , y8238 , y8239 , y8240 , y8241 , y8242 , y8243 , y8244 , y8245 , y8246 , y8247 , y8248 , y8249 , y8250 , y8251 , y8252 , y8253 , y8254 , y8255 , y8256 , y8257 , y8258 , y8259 , y8260 , y8261 , y8262 , y8263 , y8264 , y8265 , y8266 , y8267 , y8268 , y8269 , y8270 , y8271 , y8272 , y8273 , y8274 , y8275 , y8276 , y8277 , y8278 , y8279 , y8280 , y8281 , y8282 , y8283 , y8284 , y8285 , y8286 , y8287 , y8288 , y8289 , y8290 , y8291 , y8292 , y8293 , y8294 , y8295 , y8296 , y8297 , y8298 , y8299 , y8300 , y8301 , y8302 , y8303 , y8304 , y8305 , y8306 , y8307 , y8308 , y8309 , y8310 , y8311 , y8312 , y8313 , y8314 , y8315 , y8316 , y8317 , y8318 , y8319 , y8320 , y8321 , y8322 , y8323 , y8324 , y8325 , y8326 , y8327 , y8328 , y8329 , y8330 , y8331 , y8332 , y8333 , y8334 , y8335 , y8336 , y8337 , y8338 , y8339 , y8340 , y8341 , y8342 , y8343 , y8344 , y8345 , y8346 , y8347 , y8348 , y8349 , y8350 , y8351 , y8352 , y8353 , y8354 , y8355 , y8356 , y8357 , y8358 , y8359 , y8360 , y8361 , y8362 , y8363 , y8364 , y8365 , y8366 , y8367 , y8368 , y8369 , y8370 , y8371 , y8372 , y8373 , y8374 , y8375 , y8376 , y8377 , y8378 , y8379 , y8380 , y8381 , y8382 , y8383 , y8384 , y8385 , y8386 , y8387 , y8388 , y8389 , y8390 , y8391 , y8392 , y8393 , y8394 , y8395 , y8396 , y8397 , y8398 , y8399 , y8400 , y8401 , y8402 , y8403 , y8404 , y8405 , y8406 , y8407 , y8408 , y8409 , y8410 , y8411 , y8412 , y8413 , y8414 , y8415 , y8416 , y8417 , y8418 , y8419 , y8420 , y8421 , y8422 , y8423 , y8424 , y8425 , y8426 , y8427 , y8428 , y8429 , y8430 , y8431 , y8432 , y8433 , y8434 , y8435 , y8436 , y8437 , y8438 , y8439 , y8440 , y8441 , y8442 , y8443 , y8444 , y8445 , y8446 , y8447 , y8448 , y8449 , y8450 , y8451 , y8452 , y8453 , y8454 , y8455 , y8456 , y8457 , y8458 , y8459 , y8460 , y8461 , y8462 , y8463 , y8464 , y8465 , y8466 , y8467 , y8468 , y8469 , y8470 , y8471 , y8472 , y8473 , y8474 , y8475 , y8476 , y8477 , y8478 , y8479 , y8480 , y8481 , y8482 , y8483 , y8484 , y8485 , y8486 , y8487 , y8488 , y8489 , y8490 , y8491 , y8492 , y8493 , y8494 , y8495 , y8496 , y8497 , y8498 , y8499 , y8500 , y8501 , y8502 , y8503 , y8504 , y8505 , y8506 , y8507 , y8508 , y8509 , y8510 , y8511 , y8512 , y8513 , y8514 , y8515 , y8516 , y8517 , y8518 , y8519 , y8520 , y8521 , y8522 , y8523 , y8524 , y8525 , y8526 , y8527 , y8528 , y8529 , y8530 , y8531 , y8532 , y8533 , y8534 , y8535 , y8536 , y8537 , y8538 , y8539 , y8540 , y8541 , y8542 , y8543 , y8544 , y8545 , y8546 , y8547 , y8548 , y8549 , y8550 , y8551 , y8552 , y8553 , y8554 , y8555 , y8556 , y8557 , y8558 , y8559 , y8560 , y8561 , y8562 , y8563 , y8564 , y8565 , y8566 , y8567 , y8568 , y8569 , y8570 , y8571 , y8572 , y8573 , y8574 , y8575 , y8576 , y8577 , y8578 , y8579 , y8580 , y8581 , y8582 , y8583 , y8584 , y8585 , y8586 , y8587 , y8588 , y8589 , y8590 , y8591 , y8592 , y8593 , y8594 , y8595 , y8596 , y8597 , y8598 , y8599 , y8600 , y8601 , y8602 , y8603 , y8604 , y8605 , y8606 , y8607 , y8608 , y8609 , y8610 , y8611 , y8612 , y8613 , y8614 , y8615 , y8616 , y8617 , y8618 , y8619 , y8620 , y8621 , y8622 , y8623 , y8624 , y8625 , y8626 , y8627 , y8628 , y8629 , y8630 , y8631 , y8632 , y8633 , y8634 , y8635 , y8636 , y8637 , y8638 , y8639 , y8640 , y8641 , y8642 , y8643 , y8644 , y8645 , y8646 , y8647 , y8648 , y8649 , y8650 , y8651 , y8652 , y8653 , y8654 , y8655 , y8656 , y8657 , y8658 , y8659 , y8660 , y8661 , y8662 , y8663 , y8664 , y8665 , y8666 , y8667 , y8668 , y8669 , y8670 , y8671 , y8672 , y8673 , y8674 , y8675 , y8676 , y8677 , y8678 , y8679 , y8680 , y8681 , y8682 , y8683 , y8684 , y8685 , y8686 , y8687 , y8688 , y8689 , y8690 , y8691 , y8692 , y8693 , y8694 , y8695 , y8696 , y8697 , y8698 , y8699 , y8700 , y8701 , y8702 , y8703 , y8704 , y8705 , y8706 , y8707 , y8708 , y8709 , y8710 , y8711 , y8712 , y8713 , y8714 , y8715 , y8716 , y8717 , y8718 , y8719 , y8720 , y8721 , y8722 , y8723 , y8724 , y8725 , y8726 , y8727 , y8728 , y8729 , y8730 , y8731 , y8732 , y8733 , y8734 , y8735 , y8736 , y8737 , y8738 , y8739 , y8740 , y8741 , y8742 , y8743 , y8744 , y8745 , y8746 , y8747 , y8748 , y8749 , y8750 , y8751 , y8752 , y8753 , y8754 , y8755 , y8756 , y8757 , y8758 , y8759 , y8760 , y8761 , y8762 , y8763 , y8764 , y8765 , y8766 , y8767 , y8768 , y8769 , y8770 , y8771 , y8772 , y8773 , y8774 , y8775 , y8776 , y8777 , y8778 , y8779 , y8780 , y8781 , y8782 , y8783 , y8784 , y8785 , y8786 , y8787 , y8788 , y8789 , y8790 , y8791 , y8792 , y8793 , y8794 , y8795 , y8796 , y8797 , y8798 , y8799 , y8800 , y8801 , y8802 , y8803 , y8804 , y8805 , y8806 , y8807 , y8808 , y8809 , y8810 , y8811 , y8812 , y8813 , y8814 , y8815 , y8816 , y8817 , y8818 , y8819 , y8820 , y8821 , y8822 , y8823 , y8824 , y8825 , y8826 , y8827 , y8828 , y8829 , y8830 , y8831 , y8832 , y8833 , y8834 , y8835 , y8836 , y8837 , y8838 , y8839 , y8840 , y8841 , y8842 , y8843 , y8844 , y8845 , y8846 , y8847 , y8848 , y8849 , y8850 , y8851 , y8852 , y8853 , y8854 , y8855 , y8856 , y8857 , y8858 , y8859 , y8860 , y8861 , y8862 , y8863 , y8864 , y8865 , y8866 , y8867 , y8868 , y8869 , y8870 , y8871 , y8872 , y8873 , y8874 , y8875 , y8876 , y8877 , y8878 , y8879 , y8880 , y8881 , y8882 , y8883 , y8884 , y8885 , y8886 , y8887 , y8888 , y8889 , y8890 , y8891 , y8892 , y8893 , y8894 , y8895 , y8896 , y8897 , y8898 , y8899 , y8900 , y8901 , y8902 , y8903 , y8904 , y8905 , y8906 , y8907 , y8908 , y8909 , y8910 , y8911 , y8912 , y8913 , y8914 , y8915 , y8916 , y8917 , y8918 , y8919 , y8920 , y8921 , y8922 , y8923 , y8924 , y8925 , y8926 , y8927 , y8928 , y8929 , y8930 , y8931 , y8932 , y8933 , y8934 , y8935 , y8936 , y8937 , y8938 , y8939 , y8940 , y8941 , y8942 , y8943 , y8944 , y8945 , y8946 , y8947 , y8948 , y8949 , y8950 , y8951 , y8952 , y8953 , y8954 , y8955 , y8956 , y8957 , y8958 , y8959 , y8960 , y8961 , y8962 , y8963 , y8964 , y8965 , y8966 , y8967 , y8968 , y8969 , y8970 , y8971 , y8972 , y8973 , y8974 , y8975 , y8976 , y8977 , y8978 , y8979 , y8980 , y8981 , y8982 , y8983 , y8984 , y8985 , y8986 , y8987 , y8988 , y8989 , y8990 , y8991 , y8992 , y8993 , y8994 , y8995 , y8996 , y8997 , y8998 , y8999 , y9000 , y9001 , y9002 , y9003 , y9004 , y9005 , y9006 , y9007 , y9008 , y9009 , y9010 , y9011 , y9012 , y9013 , y9014 , y9015 , y9016 , y9017 , y9018 , y9019 , y9020 , y9021 , y9022 , y9023 , y9024 , y9025 , y9026 , y9027 , y9028 , y9029 , y9030 , y9031 , y9032 , y9033 , y9034 , y9035 , y9036 , y9037 , y9038 , y9039 , y9040 , y9041 , y9042 , y9043 , y9044 , y9045 , y9046 , y9047 , y9048 , y9049 , y9050 , y9051 , y9052 , y9053 , y9054 , y9055 , y9056 , y9057 , y9058 , y9059 , y9060 , y9061 , y9062 , y9063 , y9064 , y9065 , y9066 , y9067 , y9068 , y9069 , y9070 , y9071 , y9072 , y9073 , y9074 , y9075 , y9076 , y9077 , y9078 , y9079 , y9080 , y9081 , y9082 , y9083 , y9084 , y9085 , y9086 , y9087 , y9088 , y9089 , y9090 , y9091 , y9092 , y9093 , y9094 , y9095 , y9096 , y9097 , y9098 , y9099 , y9100 , y9101 , y9102 , y9103 , y9104 , y9105 , y9106 , y9107 , y9108 , y9109 , y9110 , y9111 , y9112 , y9113 , y9114 , y9115 , y9116 , y9117 , y9118 , y9119 , y9120 , y9121 , y9122 , y9123 , y9124 , y9125 , y9126 , y9127 , y9128 , y9129 , y9130 , y9131 , y9132 , y9133 , y9134 , y9135 , y9136 , y9137 , y9138 , y9139 , y9140 , y9141 , y9142 , y9143 , y9144 , y9145 , y9146 , y9147 , y9148 , y9149 , y9150 , y9151 , y9152 , y9153 , y9154 , y9155 , y9156 , y9157 , y9158 , y9159 , y9160 , y9161 , y9162 , y9163 , y9164 , y9165 , y9166 , y9167 , y9168 , y9169 , y9170 , y9171 , y9172 , y9173 , y9174 , y9175 , y9176 , y9177 , y9178 , y9179 , y9180 , y9181 , y9182 , y9183 , y9184 , y9185 , y9186 , y9187 , y9188 , y9189 , y9190 , y9191 , y9192 , y9193 , y9194 , y9195 , y9196 , y9197 , y9198 , y9199 , y9200 , y9201 , y9202 , y9203 , y9204 , y9205 , y9206 , y9207 , y9208 , y9209 , y9210 , y9211 , y9212 , y9213 , y9214 , y9215 , y9216 , y9217 , y9218 , y9219 , y9220 , y9221 , y9222 , y9223 , y9224 , y9225 , y9226 , y9227 , y9228 , y9229 , y9230 , y9231 , y9232 , y9233 , y9234 , y9235 , y9236 , y9237 , y9238 , y9239 , y9240 , y9241 , y9242 , y9243 , y9244 , y9245 , y9246 , y9247 , y9248 , y9249 , y9250 , y9251 , y9252 , y9253 , y9254 , y9255 , y9256 , y9257 , y9258 , y9259 , y9260 , y9261 , y9262 , y9263 , y9264 , y9265 , y9266 , y9267 , y9268 , y9269 , y9270 , y9271 , y9272 , y9273 , y9274 , y9275 , y9276 , y9277 , y9278 , y9279 , y9280 , y9281 , y9282 , y9283 , y9284 , y9285 , y9286 , y9287 , y9288 , y9289 , y9290 , y9291 , y9292 , y9293 , y9294 , y9295 , y9296 , y9297 , y9298 , y9299 , y9300 , y9301 , y9302 , y9303 , y9304 , y9305 , y9306 , y9307 , y9308 , y9309 , y9310 , y9311 , y9312 , y9313 , y9314 , y9315 , y9316 , y9317 , y9318 , y9319 , y9320 , y9321 , y9322 , y9323 , y9324 , y9325 , y9326 , y9327 , y9328 , y9329 , y9330 , y9331 , y9332 , y9333 , y9334 , y9335 , y9336 , y9337 , y9338 , y9339 , y9340 , y9341 , y9342 , y9343 , y9344 , y9345 , y9346 , y9347 , y9348 , y9349 , y9350 , y9351 , y9352 , y9353 , y9354 , y9355 , y9356 , y9357 , y9358 , y9359 , y9360 , y9361 , y9362 , y9363 , y9364 , y9365 , y9366 , y9367 , y9368 , y9369 , y9370 , y9371 , y9372 , y9373 , y9374 , y9375 , y9376 , y9377 , y9378 , y9379 , y9380 , y9381 , y9382 , y9383 , y9384 , y9385 , y9386 , y9387 , y9388 , y9389 , y9390 , y9391 , y9392 , y9393 , y9394 , y9395 , y9396 , y9397 , y9398 , y9399 , y9400 , y9401 , y9402 , y9403 , y9404 , y9405 , y9406 , y9407 , y9408 , y9409 , y9410 , y9411 , y9412 , y9413 , y9414 , y9415 , y9416 , y9417 , y9418 , y9419 , y9420 , y9421 , y9422 , y9423 , y9424 , y9425 , y9426 , y9427 , y9428 , y9429 , y9430 , y9431 , y9432 , y9433 , y9434 , y9435 , y9436 , y9437 , y9438 , y9439 , y9440 , y9441 , y9442 , y9443 , y9444 , y9445 , y9446 , y9447 , y9448 , y9449 , y9450 , y9451 , y9452 , y9453 , y9454 , y9455 , y9456 , y9457 , y9458 , y9459 , y9460 , y9461 , y9462 , y9463 , y9464 , y9465 , y9466 , y9467 , y9468 , y9469 , y9470 , y9471 , y9472 , y9473 , y9474 , y9475 , y9476 , y9477 , y9478 , y9479 , y9480 , y9481 , y9482 , y9483 , y9484 , y9485 , y9486 , y9487 , y9488 , y9489 , y9490 , y9491 , y9492 , y9493 , y9494 , y9495 , y9496 , y9497 , y9498 , y9499 , y9500 , y9501 , y9502 , y9503 , y9504 , y9505 , y9506 , y9507 , y9508 , y9509 , y9510 , y9511 , y9512 , y9513 , y9514 , y9515 , y9516 , y9517 , y9518 , y9519 , y9520 , y9521 , y9522 , y9523 , y9524 , y9525 , y9526 , y9527 , y9528 , y9529 , y9530 , y9531 , y9532 , y9533 , y9534 , y9535 , y9536 , y9537 , y9538 , y9539 , y9540 , y9541 , y9542 , y9543 , y9544 , y9545 , y9546 , y9547 , y9548 , y9549 , y9550 , y9551 , y9552 , y9553 , y9554 , y9555 , y9556 , y9557 , y9558 , y9559 , y9560 , y9561 , y9562 , y9563 , y9564 , y9565 , y9566 , y9567 , y9568 , y9569 , y9570 , y9571 , y9572 , y9573 , y9574 , y9575 , y9576 , y9577 , y9578 , y9579 , y9580 , y9581 , y9582 , y9583 , y9584 , y9585 , y9586 , y9587 , y9588 , y9589 , y9590 , y9591 , y9592 , y9593 , y9594 , y9595 , y9596 , y9597 , y9598 , y9599 , y9600 , y9601 , y9602 , y9603 , y9604 , y9605 , y9606 , y9607 , y9608 , y9609 , y9610 , y9611 , y9612 , y9613 , y9614 , y9615 , y9616 , y9617 , y9618 , y9619 , y9620 , y9621 , y9622 , y9623 , y9624 , y9625 , y9626 , y9627 , y9628 , y9629 , y9630 , y9631 , y9632 , y9633 , y9634 , y9635 , y9636 , y9637 , y9638 , y9639 , y9640 , y9641 , y9642 , y9643 , y9644 , y9645 , y9646 , y9647 , y9648 , y9649 , y9650 , y9651 , y9652 , y9653 , y9654 , y9655 , y9656 , y9657 , y9658 , y9659 , y9660 , y9661 , y9662 , y9663 , y9664 , y9665 , y9666 , y9667 , y9668 , y9669 , y9670 , y9671 , y9672 , y9673 , y9674 , y9675 , y9676 , y9677 , y9678 , y9679 , y9680 , y9681 , y9682 , y9683 , y9684 , y9685 , y9686 , y9687 , y9688 , y9689 , y9690 , y9691 , y9692 , y9693 , y9694 , y9695 , y9696 , y9697 , y9698 , y9699 , y9700 , y9701 , y9702 , y9703 , y9704 , y9705 , y9706 , y9707 , y9708 , y9709 , y9710 , y9711 , y9712 , y9713 , y9714 , y9715 , y9716 , y9717 , y9718 , y9719 , y9720 , y9721 , y9722 , y9723 , y9724 , y9725 , y9726 , y9727 , y9728 , y9729 , y9730 , y9731 , y9732 , y9733 , y9734 , y9735 , y9736 , y9737 , y9738 , y9739 , y9740 , y9741 , y9742 , y9743 , y9744 , y9745 , y9746 , y9747 , y9748 , y9749 , y9750 , y9751 , y9752 , y9753 , y9754 , y9755 , y9756 , y9757 , y9758 , y9759 , y9760 , y9761 , y9762 , y9763 , y9764 , y9765 , y9766 , y9767 , y9768 , y9769 , y9770 , y9771 , y9772 , y9773 , y9774 , y9775 , y9776 , y9777 , y9778 , y9779 , y9780 , y9781 , y9782 , y9783 , y9784 , y9785 , y9786 , y9787 , y9788 , y9789 , y9790 , y9791 , y9792 , y9793 , y9794 , y9795 , y9796 , y9797 , y9798 , y9799 , y9800 , y9801 , y9802 , y9803 , y9804 , y9805 , y9806 , y9807 , y9808 , y9809 , y9810 , y9811 , y9812 , y9813 , y9814 , y9815 , y9816 , y9817 , y9818 , y9819 , y9820 , y9821 , y9822 , y9823 , y9824 , y9825 , y9826 , y9827 , y9828 , y9829 , y9830 , y9831 , y9832 , y9833 , y9834 , y9835 , y9836 , y9837 , y9838 , y9839 , y9840 , y9841 , y9842 , y9843 , y9844 , y9845 , y9846 , y9847 , y9848 , y9849 , y9850 , y9851 , y9852 , y9853 , y9854 , y9855 , y9856 , y9857 , y9858 , y9859 , y9860 , y9861 , y9862 , y9863 , y9864 , y9865 , y9866 , y9867 , y9868 , y9869 , y9870 , y9871 , y9872 , y9873 , y9874 , y9875 , y9876 , y9877 , y9878 , y9879 , y9880 , y9881 , y9882 , y9883 , y9884 , y9885 , y9886 , y9887 , y9888 , y9889 , y9890 , y9891 , y9892 , y9893 , y9894 , y9895 , y9896 , y9897 , y9898 , y9899 , y9900 , y9901 , y9902 , y9903 , y9904 , y9905 , y9906 , y9907 , y9908 , y9909 , y9910 , y9911 , y9912 , y9913 , y9914 , y9915 , y9916 , y9917 , y9918 , y9919 , y9920 , y9921 , y9922 , y9923 , y9924 , y9925 , y9926 , y9927 , y9928 , y9929 , y9930 , y9931 , y9932 , y9933 , y9934 , y9935 , y9936 , y9937 , y9938 , y9939 , y9940 , y9941 , y9942 , y9943 , y9944 , y9945 , y9946 , y9947 , y9948 , y9949 , y9950 , y9951 , y9952 , y9953 , y9954 , y9955 , y9956 , y9957 , y9958 , y9959 , y9960 , y9961 , y9962 , y9963 , y9964 , y9965 , y9966 , y9967 , y9968 , y9969 , y9970 , y9971 , y9972 , y9973 , y9974 , y9975 , y9976 , y9977 , y9978 , y9979 , y9980 , y9981 , y9982 , y9983 , y9984 , y9985 , y9986 , y9987 , y9988 , y9989 , y9990 , y9991 , y9992 , y9993 , y9994 , y9995 , y9996 , y9997 , y9998 , y9999 , y10000 , y10001 , y10002 , y10003 , y10004 , y10005 , y10006 , y10007 , y10008 , y10009 , y10010 , y10011 , y10012 , y10013 , y10014 , y10015 , y10016 , y10017 , y10018 , y10019 , y10020 , y10021 , y10022 , y10023 , y10024 , y10025 , y10026 , y10027 , y10028 , y10029 , y10030 , y10031 , y10032 , y10033 , y10034 , y10035 , y10036 , y10037 , y10038 , y10039 , y10040 , y10041 , y10042 , y10043 , y10044 , y10045 , y10046 , y10047 , y10048 , y10049 , y10050 , y10051 , y10052 , y10053 , y10054 , y10055 , y10056 , y10057 , y10058 , y10059 , y10060 , y10061 , y10062 , y10063 , y10064 , y10065 , y10066 , y10067 , y10068 , y10069 , y10070 , y10071 , y10072 , y10073 , y10074 , y10075 , y10076 , y10077 , y10078 , y10079 , y10080 , y10081 , y10082 , y10083 , y10084 , y10085 , y10086 , y10087 , y10088 , y10089 , y10090 , y10091 , y10092 , y10093 , y10094 , y10095 , y10096 , y10097 , y10098 , y10099 , y10100 , y10101 , y10102 , y10103 , y10104 , y10105 , y10106 , y10107 , y10108 , y10109 , y10110 , y10111 , y10112 , y10113 , y10114 , y10115 , y10116 , y10117 , y10118 , y10119 , y10120 , y10121 , y10122 , y10123 , y10124 , y10125 , y10126 , y10127 , y10128 , y10129 , y10130 , y10131 , y10132 , y10133 , y10134 , y10135 , y10136 , y10137 , y10138 , y10139 , y10140 , y10141 , y10142 , y10143 , y10144 , y10145 , y10146 , y10147 , y10148 , y10149 , y10150 , y10151 , y10152 , y10153 , y10154 , y10155 , y10156 , y10157 , y10158 , y10159 , y10160 , y10161 , y10162 , y10163 , y10164 , y10165 , y10166 , y10167 , y10168 , y10169 , y10170 , y10171 , y10172 , y10173 , y10174 , y10175 , y10176 , y10177 , y10178 , y10179 , y10180 , y10181 , y10182 , y10183 , y10184 , y10185 , y10186 , y10187 , y10188 , y10189 , y10190 , y10191 , y10192 , y10193 , y10194 , y10195 , y10196 , y10197 , y10198 , y10199 , y10200 , y10201 , y10202 , y10203 , y10204 , y10205 , y10206 , y10207 , y10208 , y10209 , y10210 , y10211 , y10212 , y10213 , y10214 , y10215 , y10216 , y10217 , y10218 , y10219 , y10220 , y10221 , y10222 , y10223 , y10224 , y10225 , y10226 , y10227 , y10228 , y10229 , y10230 , y10231 , y10232 , y10233 , y10234 , y10235 , y10236 , y10237 , y10238 , y10239 , y10240 , y10241 , y10242 , y10243 , y10244 , y10245 , y10246 , y10247 , y10248 , y10249 , y10250 , y10251 , y10252 , y10253 , y10254 , y10255 , y10256 , y10257 , y10258 , y10259 , y10260 , y10261 , y10262 , y10263 , y10264 , y10265 , y10266 , y10267 , y10268 , y10269 , y10270 , y10271 , y10272 , y10273 , y10274 , y10275 , y10276 , y10277 , y10278 , y10279 , y10280 , y10281 , y10282 , y10283 , y10284 , y10285 , y10286 , y10287 , y10288 , y10289 , y10290 , y10291 , y10292 , y10293 , y10294 , y10295 , y10296 , y10297 , y10298 , y10299 , y10300 , y10301 , y10302 , y10303 , y10304 , y10305 , y10306 , y10307 , y10308 , y10309 , y10310 , y10311 , y10312 , y10313 , y10314 , y10315 , y10316 , y10317 , y10318 , y10319 , y10320 , y10321 , y10322 , y10323 , y10324 , y10325 , y10326 , y10327 , y10328 , y10329 , y10330 , y10331 , y10332 , y10333 , y10334 , y10335 , y10336 , y10337 , y10338 , y10339 , y10340 , y10341 , y10342 , y10343 , y10344 , y10345 , y10346 , y10347 , y10348 , y10349 , y10350 , y10351 , y10352 , y10353 , y10354 , y10355 , y10356 , y10357 , y10358 , y10359 , y10360 , y10361 , y10362 , y10363 , y10364 , y10365 , y10366 , y10367 , y10368 , y10369 , y10370 , y10371 , y10372 , y10373 , y10374 , y10375 , y10376 , y10377 , y10378 , y10379 , y10380 , y10381 , y10382 , y10383 , y10384 , y10385 , y10386 , y10387 , y10388 , y10389 , y10390 , y10391 , y10392 , y10393 , y10394 , y10395 , y10396 , y10397 , y10398 , y10399 , y10400 , y10401 , y10402 , y10403 , y10404 , y10405 , y10406 , y10407 , y10408 , y10409 , y10410 , y10411 , y10412 , y10413 , y10414 , y10415 , y10416 , y10417 , y10418 , y10419 , y10420 , y10421 , y10422 , y10423 , y10424 , y10425 , y10426 , y10427 , y10428 , y10429 , y10430 , y10431 , y10432 , y10433 , y10434 , y10435 , y10436 , y10437 , y10438 , y10439 , y10440 , y10441 , y10442 , y10443 , y10444 , y10445 , y10446 , y10447 , y10448 , y10449 , y10450 , y10451 , y10452 , y10453 , y10454 , y10455 , y10456 , y10457 , y10458 , y10459 , y10460 , y10461 , y10462 , y10463 , y10464 , y10465 , y10466 , y10467 , y10468 , y10469 , y10470 , y10471 , y10472 , y10473 , y10474 , y10475 , y10476 , y10477 , y10478 , y10479 , y10480 , y10481 , y10482 , y10483 , y10484 , y10485 , y10486 , y10487 , y10488 , y10489 , y10490 , y10491 , y10492 , y10493 , y10494 , y10495 , y10496 , y10497 , y10498 , y10499 , y10500 , y10501 , y10502 , y10503 , y10504 , y10505 , y10506 , y10507 , y10508 , y10509 , y10510 , y10511 , y10512 , y10513 , y10514 , y10515 , y10516 , y10517 , y10518 , y10519 , y10520 , y10521 , y10522 , y10523 , y10524 , y10525 , y10526 , y10527 , y10528 , y10529 , y10530 , y10531 , y10532 , y10533 , y10534 , y10535 , y10536 , y10537 , y10538 , y10539 , y10540 , y10541 , y10542 , y10543 , y10544 , y10545 , y10546 , y10547 , y10548 , y10549 , y10550 , y10551 , y10552 , y10553 , y10554 , y10555 , y10556 , y10557 , y10558 , y10559 , y10560 , y10561 , y10562 , y10563 , y10564 , y10565 , y10566 , y10567 , y10568 , y10569 , y10570 , y10571 , y10572 , y10573 , y10574 , y10575 , y10576 , y10577 , y10578 , y10579 , y10580 , y10581 , y10582 , y10583 , y10584 , y10585 , y10586 , y10587 , y10588 , y10589 , y10590 , y10591 , y10592 , y10593 , y10594 , y10595 , y10596 , y10597 , y10598 , y10599 , y10600 , y10601 , y10602 , y10603 , y10604 , y10605 , y10606 , y10607 , y10608 , y10609 , y10610 , y10611 , y10612 , y10613 , y10614 , y10615 , y10616 , y10617 , y10618 , y10619 , y10620 , y10621 , y10622 , y10623 , y10624 , y10625 , y10626 , y10627 , y10628 , y10629 , y10630 , y10631 , y10632 , y10633 , y10634 , y10635 , y10636 , y10637 , y10638 , y10639 , y10640 , y10641 , y10642 , y10643 , y10644 , y10645 , y10646 , y10647 , y10648 , y10649 , y10650 , y10651 , y10652 , y10653 , y10654 , y10655 , y10656 , y10657 , y10658 , y10659 , y10660 , y10661 , y10662 , y10663 , y10664 , y10665 , y10666 , y10667 , y10668 , y10669 , y10670 , y10671 , y10672 , y10673 , y10674 , y10675 , y10676 , y10677 , y10678 , y10679 , y10680 , y10681 , y10682 , y10683 , y10684 , y10685 , y10686 , y10687 , y10688 , y10689 , y10690 , y10691 , y10692 , y10693 , y10694 , y10695 , y10696 , y10697 , y10698 , y10699 , y10700 , y10701 , y10702 , y10703 , y10704 , y10705 , y10706 , y10707 , y10708 , y10709 , y10710 , y10711 , y10712 , y10713 , y10714 , y10715 , y10716 , y10717 , y10718 , y10719 , y10720 , y10721 , y10722 , y10723 , y10724 , y10725 , y10726 , y10727 , y10728 , y10729 , y10730 , y10731 , y10732 , y10733 , y10734 , y10735 , y10736 , y10737 , y10738 , y10739 , y10740 , y10741 , y10742 , y10743 , y10744 , y10745 , y10746 , y10747 , y10748 , y10749 , y10750 , y10751 , y10752 , y10753 , y10754 , y10755 , y10756 , y10757 , y10758 , y10759 , y10760 , y10761 , y10762 , y10763 , y10764 , y10765 , y10766 , y10767 , y10768 , y10769 , y10770 , y10771 , y10772 , y10773 , y10774 , y10775 , y10776 , y10777 , y10778 , y10779 , y10780 , y10781 , y10782 , y10783 , y10784 , y10785 , y10786 , y10787 , y10788 , y10789 , y10790 , y10791 , y10792 , y10793 , y10794 , y10795 , y10796 , y10797 , y10798 , y10799 , y10800 , y10801 , y10802 , y10803 , y10804 , y10805 , y10806 , y10807 , y10808 , y10809 , y10810 , y10811 , y10812 , y10813 , y10814 , y10815 , y10816 , y10817 , y10818 , y10819 , y10820 , y10821 , y10822 , y10823 , y10824 , y10825 , y10826 , y10827 , y10828 , y10829 , y10830 , y10831 , y10832 , y10833 , y10834 , y10835 , y10836 , y10837 , y10838 , y10839 , y10840 , y10841 , y10842 , y10843 , y10844 , y10845 , y10846 , y10847 , y10848 , y10849 , y10850 , y10851 , y10852 , y10853 , y10854 , y10855 , y10856 , y10857 , y10858 , y10859 , y10860 , y10861 , y10862 , y10863 , y10864 , y10865 , y10866 , y10867 , y10868 , y10869 , y10870 , y10871 , y10872 , y10873 , y10874 , y10875 , y10876 , y10877 , y10878 , y10879 , y10880 , y10881 , y10882 , y10883 , y10884 , y10885 , y10886 , y10887 , y10888 , y10889 , y10890 , y10891 , y10892 , y10893 , y10894 , y10895 , y10896 , y10897 , y10898 , y10899 , y10900 , y10901 , y10902 , y10903 , y10904 , y10905 , y10906 , y10907 , y10908 , y10909 , y10910 , y10911 , y10912 , y10913 , y10914 , y10915 , y10916 , y10917 , y10918 , y10919 , y10920 , y10921 , y10922 , y10923 , y10924 , y10925 , y10926 , y10927 , y10928 , y10929 , y10930 , y10931 , y10932 , y10933 , y10934 , y10935 , y10936 , y10937 , y10938 , y10939 , y10940 , y10941 , y10942 , y10943 , y10944 , y10945 , y10946 , y10947 , y10948 , y10949 , y10950 , y10951 , y10952 , y10953 , y10954 , y10955 , y10956 , y10957 , y10958 , y10959 , y10960 , y10961 , y10962 , y10963 , y10964 , y10965 , y10966 , y10967 , y10968 , y10969 , y10970 , y10971 , y10972 , y10973 , y10974 , y10975 , y10976 , y10977 , y10978 , y10979 , y10980 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 , y256 , y257 , y258 , y259 , y260 , y261 , y262 , y263 , y264 , y265 , y266 , y267 , y268 , y269 , y270 , y271 , y272 , y273 , y274 , y275 , y276 , y277 , y278 , y279 , y280 , y281 , y282 , y283 , y284 , y285 , y286 , y287 , y288 , y289 , y290 , y291 , y292 , y293 , y294 , y295 , y296 , y297 , y298 , y299 , y300 , y301 , y302 , y303 , y304 , y305 , y306 , y307 , y308 , y309 , y310 , y311 , y312 , y313 , y314 , y315 , y316 , y317 , y318 , y319 , y320 , y321 , y322 , y323 , y324 , y325 , y326 , y327 , y328 , y329 , y330 , y331 , y332 , y333 , y334 , y335 , y336 , y337 , y338 , y339 , y340 , y341 , y342 , y343 , y344 , y345 , y346 , y347 , y348 , y349 , y350 , y351 , y352 , y353 , y354 , y355 , y356 , y357 , y358 , y359 , y360 , y361 , y362 , y363 , y364 , y365 , y366 , y367 , y368 , y369 , y370 , y371 , y372 , y373 , y374 , y375 , y376 , y377 , y378 , y379 , y380 , y381 , y382 , y383 , y384 , y385 , y386 , y387 , y388 , y389 , y390 , y391 , y392 , y393 , y394 , y395 , y396 , y397 , y398 , y399 , y400 , y401 , y402 , y403 , y404 , y405 , y406 , y407 , y408 , y409 , y410 , y411 , y412 , y413 , y414 , y415 , y416 , y417 , y418 , y419 , y420 , y421 , y422 , y423 , y424 , y425 , y426 , y427 , y428 , y429 , y430 , y431 , y432 , y433 , y434 , y435 , y436 , y437 , y438 , y439 , y440 , y441 , y442 , y443 , y444 , y445 , y446 , y447 , y448 , y449 , y450 , y451 , y452 , y453 , y454 , y455 , y456 , y457 , y458 , y459 , y460 , y461 , y462 , y463 , y464 , y465 , y466 , y467 , y468 , y469 , y470 , y471 , y472 , y473 , y474 , y475 , y476 , y477 , y478 , y479 , y480 , y481 , y482 , y483 , y484 , y485 , y486 , y487 , y488 , y489 , y490 , y491 , y492 , y493 , y494 , y495 , y496 , y497 , y498 , y499 , y500 , y501 , y502 , y503 , y504 , y505 , y506 , y507 , y508 , y509 , y510 , y511 , y512 , y513 , y514 , y515 , y516 , y517 , y518 , y519 , y520 , y521 , y522 , y523 , y524 , y525 , y526 , y527 , y528 , y529 , y530 , y531 , y532 , y533 , y534 , y535 , y536 , y537 , y538 , y539 , y540 , y541 , y542 , y543 , y544 , y545 , y546 , y547 , y548 , y549 , y550 , y551 , y552 , y553 , y554 , y555 , y556 , y557 , y558 , y559 , y560 , y561 , y562 , y563 , y564 , y565 , y566 , y567 , y568 , y569 , y570 , y571 , y572 , y573 , y574 , y575 , y576 , y577 , y578 , y579 , y580 , y581 , y582 , y583 , y584 , y585 , y586 , y587 , y588 , y589 , y590 , y591 , y592 , y593 , y594 , y595 , y596 , y597 , y598 , y599 , y600 , y601 , y602 , y603 , y604 , y605 , y606 , y607 , y608 , y609 , y610 , y611 , y612 , y613 , y614 , y615 , y616 , y617 , y618 , y619 , y620 , y621 , y622 , y623 , y624 , y625 , y626 , y627 , y628 , y629 , y630 , y631 , y632 , y633 , y634 , y635 , y636 , y637 , y638 , y639 , y640 , y641 , y642 , y643 , y644 , y645 , y646 , y647 , y648 , y649 , y650 , y651 , y652 , y653 , y654 , y655 , y656 , y657 , y658 , y659 , y660 , y661 , y662 , y663 , y664 , y665 , y666 , y667 , y668 , y669 , y670 , y671 , y672 , y673 , y674 , y675 , y676 , y677 , y678 , y679 , y680 , y681 , y682 , y683 , y684 , y685 , y686 , y687 , y688 , y689 , y690 , y691 , y692 , y693 , y694 , y695 , y696 , y697 , y698 , y699 , y700 , y701 , y702 , y703 , y704 , y705 , y706 , y707 , y708 , y709 , y710 , y711 , y712 , y713 , y714 , y715 , y716 , y717 , y718 , y719 , y720 , y721 , y722 , y723 , y724 , y725 , y726 , y727 , y728 , y729 , y730 , y731 , y732 , y733 , y734 , y735 , y736 , y737 , y738 , y739 , y740 , y741 , y742 , y743 , y744 , y745 , y746 , y747 , y748 , y749 , y750 , y751 , y752 , y753 , y754 , y755 , y756 , y757 , y758 , y759 , y760 , y761 , y762 , y763 , y764 , y765 , y766 , y767 , y768 , y769 , y770 , y771 , y772 , y773 , y774 , y775 , y776 , y777 , y778 , y779 , y780 , y781 , y782 , y783 , y784 , y785 , y786 , y787 , y788 , y789 , y790 , y791 , y792 , y793 , y794 , y795 , y796 , y797 , y798 , y799 , y800 , y801 , y802 , y803 , y804 , y805 , y806 , y807 , y808 , y809 , y810 , y811 , y812 , y813 , y814 , y815 , y816 , y817 , y818 , y819 , y820 , y821 , y822 , y823 , y824 , y825 , y826 , y827 , y828 , y829 , y830 , y831 , y832 , y833 , y834 , y835 , y836 , y837 , y838 , y839 , y840 , y841 , y842 , y843 , y844 , y845 , y846 , y847 , y848 , y849 , y850 , y851 , y852 , y853 , y854 , y855 , y856 , y857 , y858 , y859 , y860 , y861 , y862 , y863 , y864 , y865 , y866 , y867 , y868 , y869 , y870 , y871 , y872 , y873 , y874 , y875 , y876 , y877 , y878 , y879 , y880 , y881 , y882 , y883 , y884 , y885 , y886 , y887 , y888 , y889 , y890 , y891 , y892 , y893 , y894 , y895 , y896 , y897 , y898 , y899 , y900 , y901 , y902 , y903 , y904 , y905 , y906 , y907 , y908 , y909 , y910 , y911 , y912 , y913 , y914 , y915 , y916 , y917 , y918 , y919 , y920 , y921 , y922 , y923 , y924 , y925 , y926 , y927 , y928 , y929 , y930 , y931 , y932 , y933 , y934 , y935 , y936 , y937 , y938 , y939 , y940 , y941 , y942 , y943 , y944 , y945 , y946 , y947 , y948 , y949 , y950 , y951 , y952 , y953 , y954 , y955 , y956 , y957 , y958 , y959 , y960 , y961 , y962 , y963 , y964 , y965 , y966 , y967 , y968 , y969 , y970 , y971 , y972 , y973 , y974 , y975 , y976 , y977 , y978 , y979 , y980 , y981 , y982 , y983 , y984 , y985 , y986 , y987 , y988 , y989 , y990 , y991 , y992 , y993 , y994 , y995 , y996 , y997 , y998 , y999 , y1000 , y1001 , y1002 , y1003 , y1004 , y1005 , y1006 , y1007 , y1008 , y1009 , y1010 , y1011 , y1012 , y1013 , y1014 , y1015 , y1016 , y1017 , y1018 , y1019 , y1020 , y1021 , y1022 , y1023 , y1024 , y1025 , y1026 , y1027 , y1028 , y1029 , y1030 , y1031 , y1032 , y1033 , y1034 , y1035 , y1036 , y1037 , y1038 , y1039 , y1040 , y1041 , y1042 , y1043 , y1044 , y1045 , y1046 , y1047 , y1048 , y1049 , y1050 , y1051 , y1052 , y1053 , y1054 , y1055 , y1056 , y1057 , y1058 , y1059 , y1060 , y1061 , y1062 , y1063 , y1064 , y1065 , y1066 , y1067 , y1068 , y1069 , y1070 , y1071 , y1072 , y1073 , y1074 , y1075 , y1076 , y1077 , y1078 , y1079 , y1080 , y1081 , y1082 , y1083 , y1084 , y1085 , y1086 , y1087 , y1088 , y1089 , y1090 , y1091 , y1092 , y1093 , y1094 , y1095 , y1096 , y1097 , y1098 , y1099 , y1100 , y1101 , y1102 , y1103 , y1104 , y1105 , y1106 , y1107 , y1108 , y1109 , y1110 , y1111 , y1112 , y1113 , y1114 , y1115 , y1116 , y1117 , y1118 , y1119 , y1120 , y1121 , y1122 , y1123 , y1124 , y1125 , y1126 , y1127 , y1128 , y1129 , y1130 , y1131 , y1132 , y1133 , y1134 , y1135 , y1136 , y1137 , y1138 , y1139 , y1140 , y1141 , y1142 , y1143 , y1144 , y1145 , y1146 , y1147 , y1148 , y1149 , y1150 , y1151 , y1152 , y1153 , y1154 , y1155 , y1156 , y1157 , y1158 , y1159 , y1160 , y1161 , y1162 , y1163 , y1164 , y1165 , y1166 , y1167 , y1168 , y1169 , y1170 , y1171 , y1172 , y1173 , y1174 , y1175 , y1176 , y1177 , y1178 , y1179 , y1180 , y1181 , y1182 , y1183 , y1184 , y1185 , y1186 , y1187 , y1188 , y1189 , y1190 , y1191 , y1192 , y1193 , y1194 , y1195 , y1196 , y1197 , y1198 , y1199 , y1200 , y1201 , y1202 , y1203 , y1204 , y1205 , y1206 , y1207 , y1208 , y1209 , y1210 , y1211 , y1212 , y1213 , y1214 , y1215 , y1216 , y1217 , y1218 , y1219 , y1220 , y1221 , y1222 , y1223 , y1224 , y1225 , y1226 , y1227 , y1228 , y1229 , y1230 , y1231 , y1232 , y1233 , y1234 , y1235 , y1236 , y1237 , y1238 , y1239 , y1240 , y1241 , y1242 , y1243 , y1244 , y1245 , y1246 , y1247 , y1248 , y1249 , y1250 , y1251 , y1252 , y1253 , y1254 , y1255 , y1256 , y1257 , y1258 , y1259 , y1260 , y1261 , y1262 , y1263 , y1264 , y1265 , y1266 , y1267 , y1268 , y1269 , y1270 , y1271 , y1272 , y1273 , y1274 , y1275 , y1276 , y1277 , y1278 , y1279 , y1280 , y1281 , y1282 , y1283 , y1284 , y1285 , y1286 , y1287 , y1288 , y1289 , y1290 , y1291 , y1292 , y1293 , y1294 , y1295 , y1296 , y1297 , y1298 , y1299 , y1300 , y1301 , y1302 , y1303 , y1304 , y1305 , y1306 , y1307 , y1308 , y1309 , y1310 , y1311 , y1312 , y1313 , y1314 , y1315 , y1316 , y1317 , y1318 , y1319 , y1320 , y1321 , y1322 , y1323 , y1324 , y1325 , y1326 , y1327 , y1328 , y1329 , y1330 , y1331 , y1332 , y1333 , y1334 , y1335 , y1336 , y1337 , y1338 , y1339 , y1340 , y1341 , y1342 , y1343 , y1344 , y1345 , y1346 , y1347 , y1348 , y1349 , y1350 , y1351 , y1352 , y1353 , y1354 , y1355 , y1356 , y1357 , y1358 , y1359 , y1360 , y1361 , y1362 , y1363 , y1364 , y1365 , y1366 , y1367 , y1368 , y1369 , y1370 , y1371 , y1372 , y1373 , y1374 , y1375 , y1376 , y1377 , y1378 , y1379 , y1380 , y1381 , y1382 , y1383 , y1384 , y1385 , y1386 , y1387 , y1388 , y1389 , y1390 , y1391 , y1392 , y1393 , y1394 , y1395 , y1396 , y1397 , y1398 , y1399 , y1400 , y1401 , y1402 , y1403 , y1404 , y1405 , y1406 , y1407 , y1408 , y1409 , y1410 , y1411 , y1412 , y1413 , y1414 , y1415 , y1416 , y1417 , y1418 , y1419 , y1420 , y1421 , y1422 , y1423 , y1424 , y1425 , y1426 , y1427 , y1428 , y1429 , y1430 , y1431 , y1432 , y1433 , y1434 , y1435 , y1436 , y1437 , y1438 , y1439 , y1440 , y1441 , y1442 , y1443 , y1444 , y1445 , y1446 , y1447 , y1448 , y1449 , y1450 , y1451 , y1452 , y1453 , y1454 , y1455 , y1456 , y1457 , y1458 , y1459 , y1460 , y1461 , y1462 , y1463 , y1464 , y1465 , y1466 , y1467 , y1468 , y1469 , y1470 , y1471 , y1472 , y1473 , y1474 , y1475 , y1476 , y1477 , y1478 , y1479 , y1480 , y1481 , y1482 , y1483 , y1484 , y1485 , y1486 , y1487 , y1488 , y1489 , y1490 , y1491 , y1492 , y1493 , y1494 , y1495 , y1496 , y1497 , y1498 , y1499 , y1500 , y1501 , y1502 , y1503 , y1504 , y1505 , y1506 , y1507 , y1508 , y1509 , y1510 , y1511 , y1512 , y1513 , y1514 , y1515 , y1516 , y1517 , y1518 , y1519 , y1520 , y1521 , y1522 , y1523 , y1524 , y1525 , y1526 , y1527 , y1528 , y1529 , y1530 , y1531 , y1532 , y1533 , y1534 , y1535 , y1536 , y1537 , y1538 , y1539 , y1540 , y1541 , y1542 , y1543 , y1544 , y1545 , y1546 , y1547 , y1548 , y1549 , y1550 , y1551 , y1552 , y1553 , y1554 , y1555 , y1556 , y1557 , y1558 , y1559 , y1560 , y1561 , y1562 , y1563 , y1564 , y1565 , y1566 , y1567 , y1568 , y1569 , y1570 , y1571 , y1572 , y1573 , y1574 , y1575 , y1576 , y1577 , y1578 , y1579 , y1580 , y1581 , y1582 , y1583 , y1584 , y1585 , y1586 , y1587 , y1588 , y1589 , y1590 , y1591 , y1592 , y1593 , y1594 , y1595 , y1596 , y1597 , y1598 , y1599 , y1600 , y1601 , y1602 , y1603 , y1604 , y1605 , y1606 , y1607 , y1608 , y1609 , y1610 , y1611 , y1612 , y1613 , y1614 , y1615 , y1616 , y1617 , y1618 , y1619 , y1620 , y1621 , y1622 , y1623 , y1624 , y1625 , y1626 , y1627 , y1628 , y1629 , y1630 , y1631 , y1632 , y1633 , y1634 , y1635 , y1636 , y1637 , y1638 , y1639 , y1640 , y1641 , y1642 , y1643 , y1644 , y1645 , y1646 , y1647 , y1648 , y1649 , y1650 , y1651 , y1652 , y1653 , y1654 , y1655 , y1656 , y1657 , y1658 , y1659 , y1660 , y1661 , y1662 , y1663 , y1664 , y1665 , y1666 , y1667 , y1668 , y1669 , y1670 , y1671 , y1672 , y1673 , y1674 , y1675 , y1676 , y1677 , y1678 , y1679 , y1680 , y1681 , y1682 , y1683 , y1684 , y1685 , y1686 , y1687 , y1688 , y1689 , y1690 , y1691 , y1692 , y1693 , y1694 , y1695 , y1696 , y1697 , y1698 , y1699 , y1700 , y1701 , y1702 , y1703 , y1704 , y1705 , y1706 , y1707 , y1708 , y1709 , y1710 , y1711 , y1712 , y1713 , y1714 , y1715 , y1716 , y1717 , y1718 , y1719 , y1720 , y1721 , y1722 , y1723 , y1724 , y1725 , y1726 , y1727 , y1728 , y1729 , y1730 , y1731 , y1732 , y1733 , y1734 , y1735 , y1736 , y1737 , y1738 , y1739 , y1740 , y1741 , y1742 , y1743 , y1744 , y1745 , y1746 , y1747 , y1748 , y1749 , y1750 , y1751 , y1752 , y1753 , y1754 , y1755 , y1756 , y1757 , y1758 , y1759 , y1760 , y1761 , y1762 , y1763 , y1764 , y1765 , y1766 , y1767 , y1768 , y1769 , y1770 , y1771 , y1772 , y1773 , y1774 , y1775 , y1776 , y1777 , y1778 , y1779 , y1780 , y1781 , y1782 , y1783 , y1784 , y1785 , y1786 , y1787 , y1788 , y1789 , y1790 , y1791 , y1792 , y1793 , y1794 , y1795 , y1796 , y1797 , y1798 , y1799 , y1800 , y1801 , y1802 , y1803 , y1804 , y1805 , y1806 , y1807 , y1808 , y1809 , y1810 , y1811 , y1812 , y1813 , y1814 , y1815 , y1816 , y1817 , y1818 , y1819 , y1820 , y1821 , y1822 , y1823 , y1824 , y1825 , y1826 , y1827 , y1828 , y1829 , y1830 , y1831 , y1832 , y1833 , y1834 , y1835 , y1836 , y1837 , y1838 , y1839 , y1840 , y1841 , y1842 , y1843 , y1844 , y1845 , y1846 , y1847 , y1848 , y1849 , y1850 , y1851 , y1852 , y1853 , y1854 , y1855 , y1856 , y1857 , y1858 , y1859 , y1860 , y1861 , y1862 , y1863 , y1864 , y1865 , y1866 , y1867 , y1868 , y1869 , y1870 , y1871 , y1872 , y1873 , y1874 , y1875 , y1876 , y1877 , y1878 , y1879 , y1880 , y1881 , y1882 , y1883 , y1884 , y1885 , y1886 , y1887 , y1888 , y1889 , y1890 , y1891 , y1892 , y1893 , y1894 , y1895 , y1896 , y1897 , y1898 , y1899 , y1900 , y1901 , y1902 , y1903 , y1904 , y1905 , y1906 , y1907 , y1908 , y1909 , y1910 , y1911 , y1912 , y1913 , y1914 , y1915 , y1916 , y1917 , y1918 , y1919 , y1920 , y1921 , y1922 , y1923 , y1924 , y1925 , y1926 , y1927 , y1928 , y1929 , y1930 , y1931 , y1932 , y1933 , y1934 , y1935 , y1936 , y1937 , y1938 , y1939 , y1940 , y1941 , y1942 , y1943 , y1944 , y1945 , y1946 , y1947 , y1948 , y1949 , y1950 , y1951 , y1952 , y1953 , y1954 , y1955 , y1956 , y1957 , y1958 , y1959 , y1960 , y1961 , y1962 , y1963 , y1964 , y1965 , y1966 , y1967 , y1968 , y1969 , y1970 , y1971 , y1972 , y1973 , y1974 , y1975 , y1976 , y1977 , y1978 , y1979 , y1980 , y1981 , y1982 , y1983 , y1984 , y1985 , y1986 , y1987 , y1988 , y1989 , y1990 , y1991 , y1992 , y1993 , y1994 , y1995 , y1996 , y1997 , y1998 , y1999 , y2000 , y2001 , y2002 , y2003 , y2004 , y2005 , y2006 , y2007 , y2008 , y2009 , y2010 , y2011 , y2012 , y2013 , y2014 , y2015 , y2016 , y2017 , y2018 , y2019 , y2020 , y2021 , y2022 , y2023 , y2024 , y2025 , y2026 , y2027 , y2028 , y2029 , y2030 , y2031 , y2032 , y2033 , y2034 , y2035 , y2036 , y2037 , y2038 , y2039 , y2040 , y2041 , y2042 , y2043 , y2044 , y2045 , y2046 , y2047 , y2048 , y2049 , y2050 , y2051 , y2052 , y2053 , y2054 , y2055 , y2056 , y2057 , y2058 , y2059 , y2060 , y2061 , y2062 , y2063 , y2064 , y2065 , y2066 , y2067 , y2068 , y2069 , y2070 , y2071 , y2072 , y2073 , y2074 , y2075 , y2076 , y2077 , y2078 , y2079 , y2080 , y2081 , y2082 , y2083 , y2084 , y2085 , y2086 , y2087 , y2088 , y2089 , y2090 , y2091 , y2092 , y2093 , y2094 , y2095 , y2096 , y2097 , y2098 , y2099 , y2100 , y2101 , y2102 , y2103 , y2104 , y2105 , y2106 , y2107 , y2108 , y2109 , y2110 , y2111 , y2112 , y2113 , y2114 , y2115 , y2116 , y2117 , y2118 , y2119 , y2120 , y2121 , y2122 , y2123 , y2124 , y2125 , y2126 , y2127 , y2128 , y2129 , y2130 , y2131 , y2132 , y2133 , y2134 , y2135 , y2136 , y2137 , y2138 , y2139 , y2140 , y2141 , y2142 , y2143 , y2144 , y2145 , y2146 , y2147 , y2148 , y2149 , y2150 , y2151 , y2152 , y2153 , y2154 , y2155 , y2156 , y2157 , y2158 , y2159 , y2160 , y2161 , y2162 , y2163 , y2164 , y2165 , y2166 , y2167 , y2168 , y2169 , y2170 , y2171 , y2172 , y2173 , y2174 , y2175 , y2176 , y2177 , y2178 , y2179 , y2180 , y2181 , y2182 , y2183 , y2184 , y2185 , y2186 , y2187 , y2188 , y2189 , y2190 , y2191 , y2192 , y2193 , y2194 , y2195 , y2196 , y2197 , y2198 , y2199 , y2200 , y2201 , y2202 , y2203 , y2204 , y2205 , y2206 , y2207 , y2208 , y2209 , y2210 , y2211 , y2212 , y2213 , y2214 , y2215 , y2216 , y2217 , y2218 , y2219 , y2220 , y2221 , y2222 , y2223 , y2224 , y2225 , y2226 , y2227 , y2228 , y2229 , y2230 , y2231 , y2232 , y2233 , y2234 , y2235 , y2236 , y2237 , y2238 , y2239 , y2240 , y2241 , y2242 , y2243 , y2244 , y2245 , y2246 , y2247 , y2248 , y2249 , y2250 , y2251 , y2252 , y2253 , y2254 , y2255 , y2256 , y2257 , y2258 , y2259 , y2260 , y2261 , y2262 , y2263 , y2264 , y2265 , y2266 , y2267 , y2268 , y2269 , y2270 , y2271 , y2272 , y2273 , y2274 , y2275 , y2276 , y2277 , y2278 , y2279 , y2280 , y2281 , y2282 , y2283 , y2284 , y2285 , y2286 , y2287 , y2288 , y2289 , y2290 , y2291 , y2292 , y2293 , y2294 , y2295 , y2296 , y2297 , y2298 , y2299 , y2300 , y2301 , y2302 , y2303 , y2304 , y2305 , y2306 , y2307 , y2308 , y2309 , y2310 , y2311 , y2312 , y2313 , y2314 , y2315 , y2316 , y2317 , y2318 , y2319 , y2320 , y2321 , y2322 , y2323 , y2324 , y2325 , y2326 , y2327 , y2328 , y2329 , y2330 , y2331 , y2332 , y2333 , y2334 , y2335 , y2336 , y2337 , y2338 , y2339 , y2340 , y2341 , y2342 , y2343 , y2344 , y2345 , y2346 , y2347 , y2348 , y2349 , y2350 , y2351 , y2352 , y2353 , y2354 , y2355 , y2356 , y2357 , y2358 , y2359 , y2360 , y2361 , y2362 , y2363 , y2364 , y2365 , y2366 , y2367 , y2368 , y2369 , y2370 , y2371 , y2372 , y2373 , y2374 , y2375 , y2376 , y2377 , y2378 , y2379 , y2380 , y2381 , y2382 , y2383 , y2384 , y2385 , y2386 , y2387 , y2388 , y2389 , y2390 , y2391 , y2392 , y2393 , y2394 , y2395 , y2396 , y2397 , y2398 , y2399 , y2400 , y2401 , y2402 , y2403 , y2404 , y2405 , y2406 , y2407 , y2408 , y2409 , y2410 , y2411 , y2412 , y2413 , y2414 , y2415 , y2416 , y2417 , y2418 , y2419 , y2420 , y2421 , y2422 , y2423 , y2424 , y2425 , y2426 , y2427 , y2428 , y2429 , y2430 , y2431 , y2432 , y2433 , y2434 , y2435 , y2436 , y2437 , y2438 , y2439 , y2440 , y2441 , y2442 , y2443 , y2444 , y2445 , y2446 , y2447 , y2448 , y2449 , y2450 , y2451 , y2452 , y2453 , y2454 , y2455 , y2456 , y2457 , y2458 , y2459 , y2460 , y2461 , y2462 , y2463 , y2464 , y2465 , y2466 , y2467 , y2468 , y2469 , y2470 , y2471 , y2472 , y2473 , y2474 , y2475 , y2476 , y2477 , y2478 , y2479 , y2480 , y2481 , y2482 , y2483 , y2484 , y2485 , y2486 , y2487 , y2488 , y2489 , y2490 , y2491 , y2492 , y2493 , y2494 , y2495 , y2496 , y2497 , y2498 , y2499 , y2500 , y2501 , y2502 , y2503 , y2504 , y2505 , y2506 , y2507 , y2508 , y2509 , y2510 , y2511 , y2512 , y2513 , y2514 , y2515 , y2516 , y2517 , y2518 , y2519 , y2520 , y2521 , y2522 , y2523 , y2524 , y2525 , y2526 , y2527 , y2528 , y2529 , y2530 , y2531 , y2532 , y2533 , y2534 , y2535 , y2536 , y2537 , y2538 , y2539 , y2540 , y2541 , y2542 , y2543 , y2544 , y2545 , y2546 , y2547 , y2548 , y2549 , y2550 , y2551 , y2552 , y2553 , y2554 , y2555 , y2556 , y2557 , y2558 , y2559 , y2560 , y2561 , y2562 , y2563 , y2564 , y2565 , y2566 , y2567 , y2568 , y2569 , y2570 , y2571 , y2572 , y2573 , y2574 , y2575 , y2576 , y2577 , y2578 , y2579 , y2580 , y2581 , y2582 , y2583 , y2584 , y2585 , y2586 , y2587 , y2588 , y2589 , y2590 , y2591 , y2592 , y2593 , y2594 , y2595 , y2596 , y2597 , y2598 , y2599 , y2600 , y2601 , y2602 , y2603 , y2604 , y2605 , y2606 , y2607 , y2608 , y2609 , y2610 , y2611 , y2612 , y2613 , y2614 , y2615 , y2616 , y2617 , y2618 , y2619 , y2620 , y2621 , y2622 , y2623 , y2624 , y2625 , y2626 , y2627 , y2628 , y2629 , y2630 , y2631 , y2632 , y2633 , y2634 , y2635 , y2636 , y2637 , y2638 , y2639 , y2640 , y2641 , y2642 , y2643 , y2644 , y2645 , y2646 , y2647 , y2648 , y2649 , y2650 , y2651 , y2652 , y2653 , y2654 , y2655 , y2656 , y2657 , y2658 , y2659 , y2660 , y2661 , y2662 , y2663 , y2664 , y2665 , y2666 , y2667 , y2668 , y2669 , y2670 , y2671 , y2672 , y2673 , y2674 , y2675 , y2676 , y2677 , y2678 , y2679 , y2680 , y2681 , y2682 , y2683 , y2684 , y2685 , y2686 , y2687 , y2688 , y2689 , y2690 , y2691 , y2692 , y2693 , y2694 , y2695 , y2696 , y2697 , y2698 , y2699 , y2700 , y2701 , y2702 , y2703 , y2704 , y2705 , y2706 , y2707 , y2708 , y2709 , y2710 , y2711 , y2712 , y2713 , y2714 , y2715 , y2716 , y2717 , y2718 , y2719 , y2720 , y2721 , y2722 , y2723 , y2724 , y2725 , y2726 , y2727 , y2728 , y2729 , y2730 , y2731 , y2732 , y2733 , y2734 , y2735 , y2736 , y2737 , y2738 , y2739 , y2740 , y2741 , y2742 , y2743 , y2744 , y2745 , y2746 , y2747 , y2748 , y2749 , y2750 , y2751 , y2752 , y2753 , y2754 , y2755 , y2756 , y2757 , y2758 , y2759 , y2760 , y2761 , y2762 , y2763 , y2764 , y2765 , y2766 , y2767 , y2768 , y2769 , y2770 , y2771 , y2772 , y2773 , y2774 , y2775 , y2776 , y2777 , y2778 , y2779 , y2780 , y2781 , y2782 , y2783 , y2784 , y2785 , y2786 , y2787 , y2788 , y2789 , y2790 , y2791 , y2792 , y2793 , y2794 , y2795 , y2796 , y2797 , y2798 , y2799 , y2800 , y2801 , y2802 , y2803 , y2804 , y2805 , y2806 , y2807 , y2808 , y2809 , y2810 , y2811 , y2812 , y2813 , y2814 , y2815 , y2816 , y2817 , y2818 , y2819 , y2820 , y2821 , y2822 , y2823 , y2824 , y2825 , y2826 , y2827 , y2828 , y2829 , y2830 , y2831 , y2832 , y2833 , y2834 , y2835 , y2836 , y2837 , y2838 , y2839 , y2840 , y2841 , y2842 , y2843 , y2844 , y2845 , y2846 , y2847 , y2848 , y2849 , y2850 , y2851 , y2852 , y2853 , y2854 , y2855 , y2856 , y2857 , y2858 , y2859 , y2860 , y2861 , y2862 , y2863 , y2864 , y2865 , y2866 , y2867 , y2868 , y2869 , y2870 , y2871 , y2872 , y2873 , y2874 , y2875 , y2876 , y2877 , y2878 , y2879 , y2880 , y2881 , y2882 , y2883 , y2884 , y2885 , y2886 , y2887 , y2888 , y2889 , y2890 , y2891 , y2892 , y2893 , y2894 , y2895 , y2896 , y2897 , y2898 , y2899 , y2900 , y2901 , y2902 , y2903 , y2904 , y2905 , y2906 , y2907 , y2908 , y2909 , y2910 , y2911 , y2912 , y2913 , y2914 , y2915 , y2916 , y2917 , y2918 , y2919 , y2920 , y2921 , y2922 , y2923 , y2924 , y2925 , y2926 , y2927 , y2928 , y2929 , y2930 , y2931 , y2932 , y2933 , y2934 , y2935 , y2936 , y2937 , y2938 , y2939 , y2940 , y2941 , y2942 , y2943 , y2944 , y2945 , y2946 , y2947 , y2948 , y2949 , y2950 , y2951 , y2952 , y2953 , y2954 , y2955 , y2956 , y2957 , y2958 , y2959 , y2960 , y2961 , y2962 , y2963 , y2964 , y2965 , y2966 , y2967 , y2968 , y2969 , y2970 , y2971 , y2972 , y2973 , y2974 , y2975 , y2976 , y2977 , y2978 , y2979 , y2980 , y2981 , y2982 , y2983 , y2984 , y2985 , y2986 , y2987 , y2988 , y2989 , y2990 , y2991 , y2992 , y2993 , y2994 , y2995 , y2996 , y2997 , y2998 , y2999 , y3000 , y3001 , y3002 , y3003 , y3004 , y3005 , y3006 , y3007 , y3008 , y3009 , y3010 , y3011 , y3012 , y3013 , y3014 , y3015 , y3016 , y3017 , y3018 , y3019 , y3020 , y3021 , y3022 , y3023 , y3024 , y3025 , y3026 , y3027 , y3028 , y3029 , y3030 , y3031 , y3032 , y3033 , y3034 , y3035 , y3036 , y3037 , y3038 , y3039 , y3040 , y3041 , y3042 , y3043 , y3044 , y3045 , y3046 , y3047 , y3048 , y3049 , y3050 , y3051 , y3052 , y3053 , y3054 , y3055 , y3056 , y3057 , y3058 , y3059 , y3060 , y3061 , y3062 , y3063 , y3064 , y3065 , y3066 , y3067 , y3068 , y3069 , y3070 , y3071 , y3072 , y3073 , y3074 , y3075 , y3076 , y3077 , y3078 , y3079 , y3080 , y3081 , y3082 , y3083 , y3084 , y3085 , y3086 , y3087 , y3088 , y3089 , y3090 , y3091 , y3092 , y3093 , y3094 , y3095 , y3096 , y3097 , y3098 , y3099 , y3100 , y3101 , y3102 , y3103 , y3104 , y3105 , y3106 , y3107 , y3108 , y3109 , y3110 , y3111 , y3112 , y3113 , y3114 , y3115 , y3116 , y3117 , y3118 , y3119 , y3120 , y3121 , y3122 , y3123 , y3124 , y3125 , y3126 , y3127 , y3128 , y3129 , y3130 , y3131 , y3132 , y3133 , y3134 , y3135 , y3136 , y3137 , y3138 , y3139 , y3140 , y3141 , y3142 , y3143 , y3144 , y3145 , y3146 , y3147 , y3148 , y3149 , y3150 , y3151 , y3152 , y3153 , y3154 , y3155 , y3156 , y3157 , y3158 , y3159 , y3160 , y3161 , y3162 , y3163 , y3164 , y3165 , y3166 , y3167 , y3168 , y3169 , y3170 , y3171 , y3172 , y3173 , y3174 , y3175 , y3176 , y3177 , y3178 , y3179 , y3180 , y3181 , y3182 , y3183 , y3184 , y3185 , y3186 , y3187 , y3188 , y3189 , y3190 , y3191 , y3192 , y3193 , y3194 , y3195 , y3196 , y3197 , y3198 , y3199 , y3200 , y3201 , y3202 , y3203 , y3204 , y3205 , y3206 , y3207 , y3208 , y3209 , y3210 , y3211 , y3212 , y3213 , y3214 , y3215 , y3216 , y3217 , y3218 , y3219 , y3220 , y3221 , y3222 , y3223 , y3224 , y3225 , y3226 , y3227 , y3228 , y3229 , y3230 , y3231 , y3232 , y3233 , y3234 , y3235 , y3236 , y3237 , y3238 , y3239 , y3240 , y3241 , y3242 , y3243 , y3244 , y3245 , y3246 , y3247 , y3248 , y3249 , y3250 , y3251 , y3252 , y3253 , y3254 , y3255 , y3256 , y3257 , y3258 , y3259 , y3260 , y3261 , y3262 , y3263 , y3264 , y3265 , y3266 , y3267 , y3268 , y3269 , y3270 , y3271 , y3272 , y3273 , y3274 , y3275 , y3276 , y3277 , y3278 , y3279 , y3280 , y3281 , y3282 , y3283 , y3284 , y3285 , y3286 , y3287 , y3288 , y3289 , y3290 , y3291 , y3292 , y3293 , y3294 , y3295 , y3296 , y3297 , y3298 , y3299 , y3300 , y3301 , y3302 , y3303 , y3304 , y3305 , y3306 , y3307 , y3308 , y3309 , y3310 , y3311 , y3312 , y3313 , y3314 , y3315 , y3316 , y3317 , y3318 , y3319 , y3320 , y3321 , y3322 , y3323 , y3324 , y3325 , y3326 , y3327 , y3328 , y3329 , y3330 , y3331 , y3332 , y3333 , y3334 , y3335 , y3336 , y3337 , y3338 , y3339 , y3340 , y3341 , y3342 , y3343 , y3344 , y3345 , y3346 , y3347 , y3348 , y3349 , y3350 , y3351 , y3352 , y3353 , y3354 , y3355 , y3356 , y3357 , y3358 , y3359 , y3360 , y3361 , y3362 , y3363 , y3364 , y3365 , y3366 , y3367 , y3368 , y3369 , y3370 , y3371 , y3372 , y3373 , y3374 , y3375 , y3376 , y3377 , y3378 , y3379 , y3380 , y3381 , y3382 , y3383 , y3384 , y3385 , y3386 , y3387 , y3388 , y3389 , y3390 , y3391 , y3392 , y3393 , y3394 , y3395 , y3396 , y3397 , y3398 , y3399 , y3400 , y3401 , y3402 , y3403 , y3404 , y3405 , y3406 , y3407 , y3408 , y3409 , y3410 , y3411 , y3412 , y3413 , y3414 , y3415 , y3416 , y3417 , y3418 , y3419 , y3420 , y3421 , y3422 , y3423 , y3424 , y3425 , y3426 , y3427 , y3428 , y3429 , y3430 , y3431 , y3432 , y3433 , y3434 , y3435 , y3436 , y3437 , y3438 , y3439 , y3440 , y3441 , y3442 , y3443 , y3444 , y3445 , y3446 , y3447 , y3448 , y3449 , y3450 , y3451 , y3452 , y3453 , y3454 , y3455 , y3456 , y3457 , y3458 , y3459 , y3460 , y3461 , y3462 , y3463 , y3464 , y3465 , y3466 , y3467 , y3468 , y3469 , y3470 , y3471 , y3472 , y3473 , y3474 , y3475 , y3476 , y3477 , y3478 , y3479 , y3480 , y3481 , y3482 , y3483 , y3484 , y3485 , y3486 , y3487 , y3488 , y3489 , y3490 , y3491 , y3492 , y3493 , y3494 , y3495 , y3496 , y3497 , y3498 , y3499 , y3500 , y3501 , y3502 , y3503 , y3504 , y3505 , y3506 , y3507 , y3508 , y3509 , y3510 , y3511 , y3512 , y3513 , y3514 , y3515 , y3516 , y3517 , y3518 , y3519 , y3520 , y3521 , y3522 , y3523 , y3524 , y3525 , y3526 , y3527 , y3528 , y3529 , y3530 , y3531 , y3532 , y3533 , y3534 , y3535 , y3536 , y3537 , y3538 , y3539 , y3540 , y3541 , y3542 , y3543 , y3544 , y3545 , y3546 , y3547 , y3548 , y3549 , y3550 , y3551 , y3552 , y3553 , y3554 , y3555 , y3556 , y3557 , y3558 , y3559 , y3560 , y3561 , y3562 , y3563 , y3564 , y3565 , y3566 , y3567 , y3568 , y3569 , y3570 , y3571 , y3572 , y3573 , y3574 , y3575 , y3576 , y3577 , y3578 , y3579 , y3580 , y3581 , y3582 , y3583 , y3584 , y3585 , y3586 , y3587 , y3588 , y3589 , y3590 , y3591 , y3592 , y3593 , y3594 , y3595 , y3596 , y3597 , y3598 , y3599 , y3600 , y3601 , y3602 , y3603 , y3604 , y3605 , y3606 , y3607 , y3608 , y3609 , y3610 , y3611 , y3612 , y3613 , y3614 , y3615 , y3616 , y3617 , y3618 , y3619 , y3620 , y3621 , y3622 , y3623 , y3624 , y3625 , y3626 , y3627 , y3628 , y3629 , y3630 , y3631 , y3632 , y3633 , y3634 , y3635 , y3636 , y3637 , y3638 , y3639 , y3640 , y3641 , y3642 , y3643 , y3644 , y3645 , y3646 , y3647 , y3648 , y3649 , y3650 , y3651 , y3652 , y3653 , y3654 , y3655 , y3656 , y3657 , y3658 , y3659 , y3660 , y3661 , y3662 , y3663 , y3664 , y3665 , y3666 , y3667 , y3668 , y3669 , y3670 , y3671 , y3672 , y3673 , y3674 , y3675 , y3676 , y3677 , y3678 , y3679 , y3680 , y3681 , y3682 , y3683 , y3684 , y3685 , y3686 , y3687 , y3688 , y3689 , y3690 , y3691 , y3692 , y3693 , y3694 , y3695 , y3696 , y3697 , y3698 , y3699 , y3700 , y3701 , y3702 , y3703 , y3704 , y3705 , y3706 , y3707 , y3708 , y3709 , y3710 , y3711 , y3712 , y3713 , y3714 , y3715 , y3716 , y3717 , y3718 , y3719 , y3720 , y3721 , y3722 , y3723 , y3724 , y3725 , y3726 , y3727 , y3728 , y3729 , y3730 , y3731 , y3732 , y3733 , y3734 , y3735 , y3736 , y3737 , y3738 , y3739 , y3740 , y3741 , y3742 , y3743 , y3744 , y3745 , y3746 , y3747 , y3748 , y3749 , y3750 , y3751 , y3752 , y3753 , y3754 , y3755 , y3756 , y3757 , y3758 , y3759 , y3760 , y3761 , y3762 , y3763 , y3764 , y3765 , y3766 , y3767 , y3768 , y3769 , y3770 , y3771 , y3772 , y3773 , y3774 , y3775 , y3776 , y3777 , y3778 , y3779 , y3780 , y3781 , y3782 , y3783 , y3784 , y3785 , y3786 , y3787 , y3788 , y3789 , y3790 , y3791 , y3792 , y3793 , y3794 , y3795 , y3796 , y3797 , y3798 , y3799 , y3800 , y3801 , y3802 , y3803 , y3804 , y3805 , y3806 , y3807 , y3808 , y3809 , y3810 , y3811 , y3812 , y3813 , y3814 , y3815 , y3816 , y3817 , y3818 , y3819 , y3820 , y3821 , y3822 , y3823 , y3824 , y3825 , y3826 , y3827 , y3828 , y3829 , y3830 , y3831 , y3832 , y3833 , y3834 , y3835 , y3836 , y3837 , y3838 , y3839 , y3840 , y3841 , y3842 , y3843 , y3844 , y3845 , y3846 , y3847 , y3848 , y3849 , y3850 , y3851 , y3852 , y3853 , y3854 , y3855 , y3856 , y3857 , y3858 , y3859 , y3860 , y3861 , y3862 , y3863 , y3864 , y3865 , y3866 , y3867 , y3868 , y3869 , y3870 , y3871 , y3872 , y3873 , y3874 , y3875 , y3876 , y3877 , y3878 , y3879 , y3880 , y3881 , y3882 , y3883 , y3884 , y3885 , y3886 , y3887 , y3888 , y3889 , y3890 , y3891 , y3892 , y3893 , y3894 , y3895 , y3896 , y3897 , y3898 , y3899 , y3900 , y3901 , y3902 , y3903 , y3904 , y3905 , y3906 , y3907 , y3908 , y3909 , y3910 , y3911 , y3912 , y3913 , y3914 , y3915 , y3916 , y3917 , y3918 , y3919 , y3920 , y3921 , y3922 , y3923 , y3924 , y3925 , y3926 , y3927 , y3928 , y3929 , y3930 , y3931 , y3932 , y3933 , y3934 , y3935 , y3936 , y3937 , y3938 , y3939 , y3940 , y3941 , y3942 , y3943 , y3944 , y3945 , y3946 , y3947 , y3948 , y3949 , y3950 , y3951 , y3952 , y3953 , y3954 , y3955 , y3956 , y3957 , y3958 , y3959 , y3960 , y3961 , y3962 , y3963 , y3964 , y3965 , y3966 , y3967 , y3968 , y3969 , y3970 , y3971 , y3972 , y3973 , y3974 , y3975 , y3976 , y3977 , y3978 , y3979 , y3980 , y3981 , y3982 , y3983 , y3984 , y3985 , y3986 , y3987 , y3988 , y3989 , y3990 , y3991 , y3992 , y3993 , y3994 , y3995 , y3996 , y3997 , y3998 , y3999 , y4000 , y4001 , y4002 , y4003 , y4004 , y4005 , y4006 , y4007 , y4008 , y4009 , y4010 , y4011 , y4012 , y4013 , y4014 , y4015 , y4016 , y4017 , y4018 , y4019 , y4020 , y4021 , y4022 , y4023 , y4024 , y4025 , y4026 , y4027 , y4028 , y4029 , y4030 , y4031 , y4032 , y4033 , y4034 , y4035 , y4036 , y4037 , y4038 , y4039 , y4040 , y4041 , y4042 , y4043 , y4044 , y4045 , y4046 , y4047 , y4048 , y4049 , y4050 , y4051 , y4052 , y4053 , y4054 , y4055 , y4056 , y4057 , y4058 , y4059 , y4060 , y4061 , y4062 , y4063 , y4064 , y4065 , y4066 , y4067 , y4068 , y4069 , y4070 , y4071 , y4072 , y4073 , y4074 , y4075 , y4076 , y4077 , y4078 , y4079 , y4080 , y4081 , y4082 , y4083 , y4084 , y4085 , y4086 , y4087 , y4088 , y4089 , y4090 , y4091 , y4092 , y4093 , y4094 , y4095 , y4096 , y4097 , y4098 , y4099 , y4100 , y4101 , y4102 , y4103 , y4104 , y4105 , y4106 , y4107 , y4108 , y4109 , y4110 , y4111 , y4112 , y4113 , y4114 , y4115 , y4116 , y4117 , y4118 , y4119 , y4120 , y4121 , y4122 , y4123 , y4124 , y4125 , y4126 , y4127 , y4128 , y4129 , y4130 , y4131 , y4132 , y4133 , y4134 , y4135 , y4136 , y4137 , y4138 , y4139 , y4140 , y4141 , y4142 , y4143 , y4144 , y4145 , y4146 , y4147 , y4148 , y4149 , y4150 , y4151 , y4152 , y4153 , y4154 , y4155 , y4156 , y4157 , y4158 , y4159 , y4160 , y4161 , y4162 , y4163 , y4164 , y4165 , y4166 , y4167 , y4168 , y4169 , y4170 , y4171 , y4172 , y4173 , y4174 , y4175 , y4176 , y4177 , y4178 , y4179 , y4180 , y4181 , y4182 , y4183 , y4184 , y4185 , y4186 , y4187 , y4188 , y4189 , y4190 , y4191 , y4192 , y4193 , y4194 , y4195 , y4196 , y4197 , y4198 , y4199 , y4200 , y4201 , y4202 , y4203 , y4204 , y4205 , y4206 , y4207 , y4208 , y4209 , y4210 , y4211 , y4212 , y4213 , y4214 , y4215 , y4216 , y4217 , y4218 , y4219 , y4220 , y4221 , y4222 , y4223 , y4224 , y4225 , y4226 , y4227 , y4228 , y4229 , y4230 , y4231 , y4232 , y4233 , y4234 , y4235 , y4236 , y4237 , y4238 , y4239 , y4240 , y4241 , y4242 , y4243 , y4244 , y4245 , y4246 , y4247 , y4248 , y4249 , y4250 , y4251 , y4252 , y4253 , y4254 , y4255 , y4256 , y4257 , y4258 , y4259 , y4260 , y4261 , y4262 , y4263 , y4264 , y4265 , y4266 , y4267 , y4268 , y4269 , y4270 , y4271 , y4272 , y4273 , y4274 , y4275 , y4276 , y4277 , y4278 , y4279 , y4280 , y4281 , y4282 , y4283 , y4284 , y4285 , y4286 , y4287 , y4288 , y4289 , y4290 , y4291 , y4292 , y4293 , y4294 , y4295 , y4296 , y4297 , y4298 , y4299 , y4300 , y4301 , y4302 , y4303 , y4304 , y4305 , y4306 , y4307 , y4308 , y4309 , y4310 , y4311 , y4312 , y4313 , y4314 , y4315 , y4316 , y4317 , y4318 , y4319 , y4320 , y4321 , y4322 , y4323 , y4324 , y4325 , y4326 , y4327 , y4328 , y4329 , y4330 , y4331 , y4332 , y4333 , y4334 , y4335 , y4336 , y4337 , y4338 , y4339 , y4340 , y4341 , y4342 , y4343 , y4344 , y4345 , y4346 , y4347 , y4348 , y4349 , y4350 , y4351 , y4352 , y4353 , y4354 , y4355 , y4356 , y4357 , y4358 , y4359 , y4360 , y4361 , y4362 , y4363 , y4364 , y4365 , y4366 , y4367 , y4368 , y4369 , y4370 , y4371 , y4372 , y4373 , y4374 , y4375 , y4376 , y4377 , y4378 , y4379 , y4380 , y4381 , y4382 , y4383 , y4384 , y4385 , y4386 , y4387 , y4388 , y4389 , y4390 , y4391 , y4392 , y4393 , y4394 , y4395 , y4396 , y4397 , y4398 , y4399 , y4400 , y4401 , y4402 , y4403 , y4404 , y4405 , y4406 , y4407 , y4408 , y4409 , y4410 , y4411 , y4412 , y4413 , y4414 , y4415 , y4416 , y4417 , y4418 , y4419 , y4420 , y4421 , y4422 , y4423 , y4424 , y4425 , y4426 , y4427 , y4428 , y4429 , y4430 , y4431 , y4432 , y4433 , y4434 , y4435 , y4436 , y4437 , y4438 , y4439 , y4440 , y4441 , y4442 , y4443 , y4444 , y4445 , y4446 , y4447 , y4448 , y4449 , y4450 , y4451 , y4452 , y4453 , y4454 , y4455 , y4456 , y4457 , y4458 , y4459 , y4460 , y4461 , y4462 , y4463 , y4464 , y4465 , y4466 , y4467 , y4468 , y4469 , y4470 , y4471 , y4472 , y4473 , y4474 , y4475 , y4476 , y4477 , y4478 , y4479 , y4480 , y4481 , y4482 , y4483 , y4484 , y4485 , y4486 , y4487 , y4488 , y4489 , y4490 , y4491 , y4492 , y4493 , y4494 , y4495 , y4496 , y4497 , y4498 , y4499 , y4500 , y4501 , y4502 , y4503 , y4504 , y4505 , y4506 , y4507 , y4508 , y4509 , y4510 , y4511 , y4512 , y4513 , y4514 , y4515 , y4516 , y4517 , y4518 , y4519 , y4520 , y4521 , y4522 , y4523 , y4524 , y4525 , y4526 , y4527 , y4528 , y4529 , y4530 , y4531 , y4532 , y4533 , y4534 , y4535 , y4536 , y4537 , y4538 , y4539 , y4540 , y4541 , y4542 , y4543 , y4544 , y4545 , y4546 , y4547 , y4548 , y4549 , y4550 , y4551 , y4552 , y4553 , y4554 , y4555 , y4556 , y4557 , y4558 , y4559 , y4560 , y4561 , y4562 , y4563 , y4564 , y4565 , y4566 , y4567 , y4568 , y4569 , y4570 , y4571 , y4572 , y4573 , y4574 , y4575 , y4576 , y4577 , y4578 , y4579 , y4580 , y4581 , y4582 , y4583 , y4584 , y4585 , y4586 , y4587 , y4588 , y4589 , y4590 , y4591 , y4592 , y4593 , y4594 , y4595 , y4596 , y4597 , y4598 , y4599 , y4600 , y4601 , y4602 , y4603 , y4604 , y4605 , y4606 , y4607 , y4608 , y4609 , y4610 , y4611 , y4612 , y4613 , y4614 , y4615 , y4616 , y4617 , y4618 , y4619 , y4620 , y4621 , y4622 , y4623 , y4624 , y4625 , y4626 , y4627 , y4628 , y4629 , y4630 , y4631 , y4632 , y4633 , y4634 , y4635 , y4636 , y4637 , y4638 , y4639 , y4640 , y4641 , y4642 , y4643 , y4644 , y4645 , y4646 , y4647 , y4648 , y4649 , y4650 , y4651 , y4652 , y4653 , y4654 , y4655 , y4656 , y4657 , y4658 , y4659 , y4660 , y4661 , y4662 , y4663 , y4664 , y4665 , y4666 , y4667 , y4668 , y4669 , y4670 , y4671 , y4672 , y4673 , y4674 , y4675 , y4676 , y4677 , y4678 , y4679 , y4680 , y4681 , y4682 , y4683 , y4684 , y4685 , y4686 , y4687 , y4688 , y4689 , y4690 , y4691 , y4692 , y4693 , y4694 , y4695 , y4696 , y4697 , y4698 , y4699 , y4700 , y4701 , y4702 , y4703 , y4704 , y4705 , y4706 , y4707 , y4708 , y4709 , y4710 , y4711 , y4712 , y4713 , y4714 , y4715 , y4716 , y4717 , y4718 , y4719 , y4720 , y4721 , y4722 , y4723 , y4724 , y4725 , y4726 , y4727 , y4728 , y4729 , y4730 , y4731 , y4732 , y4733 , y4734 , y4735 , y4736 , y4737 , y4738 , y4739 , y4740 , y4741 , y4742 , y4743 , y4744 , y4745 , y4746 , y4747 , y4748 , y4749 , y4750 , y4751 , y4752 , y4753 , y4754 , y4755 , y4756 , y4757 , y4758 , y4759 , y4760 , y4761 , y4762 , y4763 , y4764 , y4765 , y4766 , y4767 , y4768 , y4769 , y4770 , y4771 , y4772 , y4773 , y4774 , y4775 , y4776 , y4777 , y4778 , y4779 , y4780 , y4781 , y4782 , y4783 , y4784 , y4785 , y4786 , y4787 , y4788 , y4789 , y4790 , y4791 , y4792 , y4793 , y4794 , y4795 , y4796 , y4797 , y4798 , y4799 , y4800 , y4801 , y4802 , y4803 , y4804 , y4805 , y4806 , y4807 , y4808 , y4809 , y4810 , y4811 , y4812 , y4813 , y4814 , y4815 , y4816 , y4817 , y4818 , y4819 , y4820 , y4821 , y4822 , y4823 , y4824 , y4825 , y4826 , y4827 , y4828 , y4829 , y4830 , y4831 , y4832 , y4833 , y4834 , y4835 , y4836 , y4837 , y4838 , y4839 , y4840 , y4841 , y4842 , y4843 , y4844 , y4845 , y4846 , y4847 , y4848 , y4849 , y4850 , y4851 , y4852 , y4853 , y4854 , y4855 , y4856 , y4857 , y4858 , y4859 , y4860 , y4861 , y4862 , y4863 , y4864 , y4865 , y4866 , y4867 , y4868 , y4869 , y4870 , y4871 , y4872 , y4873 , y4874 , y4875 , y4876 , y4877 , y4878 , y4879 , y4880 , y4881 , y4882 , y4883 , y4884 , y4885 , y4886 , y4887 , y4888 , y4889 , y4890 , y4891 , y4892 , y4893 , y4894 , y4895 , y4896 , y4897 , y4898 , y4899 , y4900 , y4901 , y4902 , y4903 , y4904 , y4905 , y4906 , y4907 , y4908 , y4909 , y4910 , y4911 , y4912 , y4913 , y4914 , y4915 , y4916 , y4917 , y4918 , y4919 , y4920 , y4921 , y4922 , y4923 , y4924 , y4925 , y4926 , y4927 , y4928 , y4929 , y4930 , y4931 , y4932 , y4933 , y4934 , y4935 , y4936 , y4937 , y4938 , y4939 , y4940 , y4941 , y4942 , y4943 , y4944 , y4945 , y4946 , y4947 , y4948 , y4949 , y4950 , y4951 , y4952 , y4953 , y4954 , y4955 , y4956 , y4957 , y4958 , y4959 , y4960 , y4961 , y4962 , y4963 , y4964 , y4965 , y4966 , y4967 , y4968 , y4969 , y4970 , y4971 , y4972 , y4973 , y4974 , y4975 , y4976 , y4977 , y4978 , y4979 , y4980 , y4981 , y4982 , y4983 , y4984 , y4985 , y4986 , y4987 , y4988 , y4989 , y4990 , y4991 , y4992 , y4993 , y4994 , y4995 , y4996 , y4997 , y4998 , y4999 , y5000 , y5001 , y5002 , y5003 , y5004 , y5005 , y5006 , y5007 , y5008 , y5009 , y5010 , y5011 , y5012 , y5013 , y5014 , y5015 , y5016 , y5017 , y5018 , y5019 , y5020 , y5021 , y5022 , y5023 , y5024 , y5025 , y5026 , y5027 , y5028 , y5029 , y5030 , y5031 , y5032 , y5033 , y5034 , y5035 , y5036 , y5037 , y5038 , y5039 , y5040 , y5041 , y5042 , y5043 , y5044 , y5045 , y5046 , y5047 , y5048 , y5049 , y5050 , y5051 , y5052 , y5053 , y5054 , y5055 , y5056 , y5057 , y5058 , y5059 , y5060 , y5061 , y5062 , y5063 , y5064 , y5065 , y5066 , y5067 , y5068 , y5069 , y5070 , y5071 , y5072 , y5073 , y5074 , y5075 , y5076 , y5077 , y5078 , y5079 , y5080 , y5081 , y5082 , y5083 , y5084 , y5085 , y5086 , y5087 , y5088 , y5089 , y5090 , y5091 , y5092 , y5093 , y5094 , y5095 , y5096 , y5097 , y5098 , y5099 , y5100 , y5101 , y5102 , y5103 , y5104 , y5105 , y5106 , y5107 , y5108 , y5109 , y5110 , y5111 , y5112 , y5113 , y5114 , y5115 , y5116 , y5117 , y5118 , y5119 , y5120 , y5121 , y5122 , y5123 , y5124 , y5125 , y5126 , y5127 , y5128 , y5129 , y5130 , y5131 , y5132 , y5133 , y5134 , y5135 , y5136 , y5137 , y5138 , y5139 , y5140 , y5141 , y5142 , y5143 , y5144 , y5145 , y5146 , y5147 , y5148 , y5149 , y5150 , y5151 , y5152 , y5153 , y5154 , y5155 , y5156 , y5157 , y5158 , y5159 , y5160 , y5161 , y5162 , y5163 , y5164 , y5165 , y5166 , y5167 , y5168 , y5169 , y5170 , y5171 , y5172 , y5173 , y5174 , y5175 , y5176 , y5177 , y5178 , y5179 , y5180 , y5181 , y5182 , y5183 , y5184 , y5185 , y5186 , y5187 , y5188 , y5189 , y5190 , y5191 , y5192 , y5193 , y5194 , y5195 , y5196 , y5197 , y5198 , y5199 , y5200 , y5201 , y5202 , y5203 , y5204 , y5205 , y5206 , y5207 , y5208 , y5209 , y5210 , y5211 , y5212 , y5213 , y5214 , y5215 , y5216 , y5217 , y5218 , y5219 , y5220 , y5221 , y5222 , y5223 , y5224 , y5225 , y5226 , y5227 , y5228 , y5229 , y5230 , y5231 , y5232 , y5233 , y5234 , y5235 , y5236 , y5237 , y5238 , y5239 , y5240 , y5241 , y5242 , y5243 , y5244 , y5245 , y5246 , y5247 , y5248 , y5249 , y5250 , y5251 , y5252 , y5253 , y5254 , y5255 , y5256 , y5257 , y5258 , y5259 , y5260 , y5261 , y5262 , y5263 , y5264 , y5265 , y5266 , y5267 , y5268 , y5269 , y5270 , y5271 , y5272 , y5273 , y5274 , y5275 , y5276 , y5277 , y5278 , y5279 , y5280 , y5281 , y5282 , y5283 , y5284 , y5285 , y5286 , y5287 , y5288 , y5289 , y5290 , y5291 , y5292 , y5293 , y5294 , y5295 , y5296 , y5297 , y5298 , y5299 , y5300 , y5301 , y5302 , y5303 , y5304 , y5305 , y5306 , y5307 , y5308 , y5309 , y5310 , y5311 , y5312 , y5313 , y5314 , y5315 , y5316 , y5317 , y5318 , y5319 , y5320 , y5321 , y5322 , y5323 , y5324 , y5325 , y5326 , y5327 , y5328 , y5329 , y5330 , y5331 , y5332 , y5333 , y5334 , y5335 , y5336 , y5337 , y5338 , y5339 , y5340 , y5341 , y5342 , y5343 , y5344 , y5345 , y5346 , y5347 , y5348 , y5349 , y5350 , y5351 , y5352 , y5353 , y5354 , y5355 , y5356 , y5357 , y5358 , y5359 , y5360 , y5361 , y5362 , y5363 , y5364 , y5365 , y5366 , y5367 , y5368 , y5369 , y5370 , y5371 , y5372 , y5373 , y5374 , y5375 , y5376 , y5377 , y5378 , y5379 , y5380 , y5381 , y5382 , y5383 , y5384 , y5385 , y5386 , y5387 , y5388 , y5389 , y5390 , y5391 , y5392 , y5393 , y5394 , y5395 , y5396 , y5397 , y5398 , y5399 , y5400 , y5401 , y5402 , y5403 , y5404 , y5405 , y5406 , y5407 , y5408 , y5409 , y5410 , y5411 , y5412 , y5413 , y5414 , y5415 , y5416 , y5417 , y5418 , y5419 , y5420 , y5421 , y5422 , y5423 , y5424 , y5425 , y5426 , y5427 , y5428 , y5429 , y5430 , y5431 , y5432 , y5433 , y5434 , y5435 , y5436 , y5437 , y5438 , y5439 , y5440 , y5441 , y5442 , y5443 , y5444 , y5445 , y5446 , y5447 , y5448 , y5449 , y5450 , y5451 , y5452 , y5453 , y5454 , y5455 , y5456 , y5457 , y5458 , y5459 , y5460 , y5461 , y5462 , y5463 , y5464 , y5465 , y5466 , y5467 , y5468 , y5469 , y5470 , y5471 , y5472 , y5473 , y5474 , y5475 , y5476 , y5477 , y5478 , y5479 , y5480 , y5481 , y5482 , y5483 , y5484 , y5485 , y5486 , y5487 , y5488 , y5489 , y5490 , y5491 , y5492 , y5493 , y5494 , y5495 , y5496 , y5497 , y5498 , y5499 , y5500 , y5501 , y5502 , y5503 , y5504 , y5505 , y5506 , y5507 , y5508 , y5509 , y5510 , y5511 , y5512 , y5513 , y5514 , y5515 , y5516 , y5517 , y5518 , y5519 , y5520 , y5521 , y5522 , y5523 , y5524 , y5525 , y5526 , y5527 , y5528 , y5529 , y5530 , y5531 , y5532 , y5533 , y5534 , y5535 , y5536 , y5537 , y5538 , y5539 , y5540 , y5541 , y5542 , y5543 , y5544 , y5545 , y5546 , y5547 , y5548 , y5549 , y5550 , y5551 , y5552 , y5553 , y5554 , y5555 , y5556 , y5557 , y5558 , y5559 , y5560 , y5561 , y5562 , y5563 , y5564 , y5565 , y5566 , y5567 , y5568 , y5569 , y5570 , y5571 , y5572 , y5573 , y5574 , y5575 , y5576 , y5577 , y5578 , y5579 , y5580 , y5581 , y5582 , y5583 , y5584 , y5585 , y5586 , y5587 , y5588 , y5589 , y5590 , y5591 , y5592 , y5593 , y5594 , y5595 , y5596 , y5597 , y5598 , y5599 , y5600 , y5601 , y5602 , y5603 , y5604 , y5605 , y5606 , y5607 , y5608 , y5609 , y5610 , y5611 , y5612 , y5613 , y5614 , y5615 , y5616 , y5617 , y5618 , y5619 , y5620 , y5621 , y5622 , y5623 , y5624 , y5625 , y5626 , y5627 , y5628 , y5629 , y5630 , y5631 , y5632 , y5633 , y5634 , y5635 , y5636 , y5637 , y5638 , y5639 , y5640 , y5641 , y5642 , y5643 , y5644 , y5645 , y5646 , y5647 , y5648 , y5649 , y5650 , y5651 , y5652 , y5653 , y5654 , y5655 , y5656 , y5657 , y5658 , y5659 , y5660 , y5661 , y5662 , y5663 , y5664 , y5665 , y5666 , y5667 , y5668 , y5669 , y5670 , y5671 , y5672 , y5673 , y5674 , y5675 , y5676 , y5677 , y5678 , y5679 , y5680 , y5681 , y5682 , y5683 , y5684 , y5685 , y5686 , y5687 , y5688 , y5689 , y5690 , y5691 , y5692 , y5693 , y5694 , y5695 , y5696 , y5697 , y5698 , y5699 , y5700 , y5701 , y5702 , y5703 , y5704 , y5705 , y5706 , y5707 , y5708 , y5709 , y5710 , y5711 , y5712 , y5713 , y5714 , y5715 , y5716 , y5717 , y5718 , y5719 , y5720 , y5721 , y5722 , y5723 , y5724 , y5725 , y5726 , y5727 , y5728 , y5729 , y5730 , y5731 , y5732 , y5733 , y5734 , y5735 , y5736 , y5737 , y5738 , y5739 , y5740 , y5741 , y5742 , y5743 , y5744 , y5745 , y5746 , y5747 , y5748 , y5749 , y5750 , y5751 , y5752 , y5753 , y5754 , y5755 , y5756 , y5757 , y5758 , y5759 , y5760 , y5761 , y5762 , y5763 , y5764 , y5765 , y5766 , y5767 , y5768 , y5769 , y5770 , y5771 , y5772 , y5773 , y5774 , y5775 , y5776 , y5777 , y5778 , y5779 , y5780 , y5781 , y5782 , y5783 , y5784 , y5785 , y5786 , y5787 , y5788 , y5789 , y5790 , y5791 , y5792 , y5793 , y5794 , y5795 , y5796 , y5797 , y5798 , y5799 , y5800 , y5801 , y5802 , y5803 , y5804 , y5805 , y5806 , y5807 , y5808 , y5809 , y5810 , y5811 , y5812 , y5813 , y5814 , y5815 , y5816 , y5817 , y5818 , y5819 , y5820 , y5821 , y5822 , y5823 , y5824 , y5825 , y5826 , y5827 , y5828 , y5829 , y5830 , y5831 , y5832 , y5833 , y5834 , y5835 , y5836 , y5837 , y5838 , y5839 , y5840 , y5841 , y5842 , y5843 , y5844 , y5845 , y5846 , y5847 , y5848 , y5849 , y5850 , y5851 , y5852 , y5853 , y5854 , y5855 , y5856 , y5857 , y5858 , y5859 , y5860 , y5861 , y5862 , y5863 , y5864 , y5865 , y5866 , y5867 , y5868 , y5869 , y5870 , y5871 , y5872 , y5873 , y5874 , y5875 , y5876 , y5877 , y5878 , y5879 , y5880 , y5881 , y5882 , y5883 , y5884 , y5885 , y5886 , y5887 , y5888 , y5889 , y5890 , y5891 , y5892 , y5893 , y5894 , y5895 , y5896 , y5897 , y5898 , y5899 , y5900 , y5901 , y5902 , y5903 , y5904 , y5905 , y5906 , y5907 , y5908 , y5909 , y5910 , y5911 , y5912 , y5913 , y5914 , y5915 , y5916 , y5917 , y5918 , y5919 , y5920 , y5921 , y5922 , y5923 , y5924 , y5925 , y5926 , y5927 , y5928 , y5929 , y5930 , y5931 , y5932 , y5933 , y5934 , y5935 , y5936 , y5937 , y5938 , y5939 , y5940 , y5941 , y5942 , y5943 , y5944 , y5945 , y5946 , y5947 , y5948 , y5949 , y5950 , y5951 , y5952 , y5953 , y5954 , y5955 , y5956 , y5957 , y5958 , y5959 , y5960 , y5961 , y5962 , y5963 , y5964 , y5965 , y5966 , y5967 , y5968 , y5969 , y5970 , y5971 , y5972 , y5973 , y5974 , y5975 , y5976 , y5977 , y5978 , y5979 , y5980 , y5981 , y5982 , y5983 , y5984 , y5985 , y5986 , y5987 , y5988 , y5989 , y5990 , y5991 , y5992 , y5993 , y5994 , y5995 , y5996 , y5997 , y5998 , y5999 , y6000 , y6001 , y6002 , y6003 , y6004 , y6005 , y6006 , y6007 , y6008 , y6009 , y6010 , y6011 , y6012 , y6013 , y6014 , y6015 , y6016 , y6017 , y6018 , y6019 , y6020 , y6021 , y6022 , y6023 , y6024 , y6025 , y6026 , y6027 , y6028 , y6029 , y6030 , y6031 , y6032 , y6033 , y6034 , y6035 , y6036 , y6037 , y6038 , y6039 , y6040 , y6041 , y6042 , y6043 , y6044 , y6045 , y6046 , y6047 , y6048 , y6049 , y6050 , y6051 , y6052 , y6053 , y6054 , y6055 , y6056 , y6057 , y6058 , y6059 , y6060 , y6061 , y6062 , y6063 , y6064 , y6065 , y6066 , y6067 , y6068 , y6069 , y6070 , y6071 , y6072 , y6073 , y6074 , y6075 , y6076 , y6077 , y6078 , y6079 , y6080 , y6081 , y6082 , y6083 , y6084 , y6085 , y6086 , y6087 , y6088 , y6089 , y6090 , y6091 , y6092 , y6093 , y6094 , y6095 , y6096 , y6097 , y6098 , y6099 , y6100 , y6101 , y6102 , y6103 , y6104 , y6105 , y6106 , y6107 , y6108 , y6109 , y6110 , y6111 , y6112 , y6113 , y6114 , y6115 , y6116 , y6117 , y6118 , y6119 , y6120 , y6121 , y6122 , y6123 , y6124 , y6125 , y6126 , y6127 , y6128 , y6129 , y6130 , y6131 , y6132 , y6133 , y6134 , y6135 , y6136 , y6137 , y6138 , y6139 , y6140 , y6141 , y6142 , y6143 , y6144 , y6145 , y6146 , y6147 , y6148 , y6149 , y6150 , y6151 , y6152 , y6153 , y6154 , y6155 , y6156 , y6157 , y6158 , y6159 , y6160 , y6161 , y6162 , y6163 , y6164 , y6165 , y6166 , y6167 , y6168 , y6169 , y6170 , y6171 , y6172 , y6173 , y6174 , y6175 , y6176 , y6177 , y6178 , y6179 , y6180 , y6181 , y6182 , y6183 , y6184 , y6185 , y6186 , y6187 , y6188 , y6189 , y6190 , y6191 , y6192 , y6193 , y6194 , y6195 , y6196 , y6197 , y6198 , y6199 , y6200 , y6201 , y6202 , y6203 , y6204 , y6205 , y6206 , y6207 , y6208 , y6209 , y6210 , y6211 , y6212 , y6213 , y6214 , y6215 , y6216 , y6217 , y6218 , y6219 , y6220 , y6221 , y6222 , y6223 , y6224 , y6225 , y6226 , y6227 , y6228 , y6229 , y6230 , y6231 , y6232 , y6233 , y6234 , y6235 , y6236 , y6237 , y6238 , y6239 , y6240 , y6241 , y6242 , y6243 , y6244 , y6245 , y6246 , y6247 , y6248 , y6249 , y6250 , y6251 , y6252 , y6253 , y6254 , y6255 , y6256 , y6257 , y6258 , y6259 , y6260 , y6261 , y6262 , y6263 , y6264 , y6265 , y6266 , y6267 , y6268 , y6269 , y6270 , y6271 , y6272 , y6273 , y6274 , y6275 , y6276 , y6277 , y6278 , y6279 , y6280 , y6281 , y6282 , y6283 , y6284 , y6285 , y6286 , y6287 , y6288 , y6289 , y6290 , y6291 , y6292 , y6293 , y6294 , y6295 , y6296 , y6297 , y6298 , y6299 , y6300 , y6301 , y6302 , y6303 , y6304 , y6305 , y6306 , y6307 , y6308 , y6309 , y6310 , y6311 , y6312 , y6313 , y6314 , y6315 , y6316 , y6317 , y6318 , y6319 , y6320 , y6321 , y6322 , y6323 , y6324 , y6325 , y6326 , y6327 , y6328 , y6329 , y6330 , y6331 , y6332 , y6333 , y6334 , y6335 , y6336 , y6337 , y6338 , y6339 , y6340 , y6341 , y6342 , y6343 , y6344 , y6345 , y6346 , y6347 , y6348 , y6349 , y6350 , y6351 , y6352 , y6353 , y6354 , y6355 , y6356 , y6357 , y6358 , y6359 , y6360 , y6361 , y6362 , y6363 , y6364 , y6365 , y6366 , y6367 , y6368 , y6369 , y6370 , y6371 , y6372 , y6373 , y6374 , y6375 , y6376 , y6377 , y6378 , y6379 , y6380 , y6381 , y6382 , y6383 , y6384 , y6385 , y6386 , y6387 , y6388 , y6389 , y6390 , y6391 , y6392 , y6393 , y6394 , y6395 , y6396 , y6397 , y6398 , y6399 , y6400 , y6401 , y6402 , y6403 , y6404 , y6405 , y6406 , y6407 , y6408 , y6409 , y6410 , y6411 , y6412 , y6413 , y6414 , y6415 , y6416 , y6417 , y6418 , y6419 , y6420 , y6421 , y6422 , y6423 , y6424 , y6425 , y6426 , y6427 , y6428 , y6429 , y6430 , y6431 , y6432 , y6433 , y6434 , y6435 , y6436 , y6437 , y6438 , y6439 , y6440 , y6441 , y6442 , y6443 , y6444 , y6445 , y6446 , y6447 , y6448 , y6449 , y6450 , y6451 , y6452 , y6453 , y6454 , y6455 , y6456 , y6457 , y6458 , y6459 , y6460 , y6461 , y6462 , y6463 , y6464 , y6465 , y6466 , y6467 , y6468 , y6469 , y6470 , y6471 , y6472 , y6473 , y6474 , y6475 , y6476 , y6477 , y6478 , y6479 , y6480 , y6481 , y6482 , y6483 , y6484 , y6485 , y6486 , y6487 , y6488 , y6489 , y6490 , y6491 , y6492 , y6493 , y6494 , y6495 , y6496 , y6497 , y6498 , y6499 , y6500 , y6501 , y6502 , y6503 , y6504 , y6505 , y6506 , y6507 , y6508 , y6509 , y6510 , y6511 , y6512 , y6513 , y6514 , y6515 , y6516 , y6517 , y6518 , y6519 , y6520 , y6521 , y6522 , y6523 , y6524 , y6525 , y6526 , y6527 , y6528 , y6529 , y6530 , y6531 , y6532 , y6533 , y6534 , y6535 , y6536 , y6537 , y6538 , y6539 , y6540 , y6541 , y6542 , y6543 , y6544 , y6545 , y6546 , y6547 , y6548 , y6549 , y6550 , y6551 , y6552 , y6553 , y6554 , y6555 , y6556 , y6557 , y6558 , y6559 , y6560 , y6561 , y6562 , y6563 , y6564 , y6565 , y6566 , y6567 , y6568 , y6569 , y6570 , y6571 , y6572 , y6573 , y6574 , y6575 , y6576 , y6577 , y6578 , y6579 , y6580 , y6581 , y6582 , y6583 , y6584 , y6585 , y6586 , y6587 , y6588 , y6589 , y6590 , y6591 , y6592 , y6593 , y6594 , y6595 , y6596 , y6597 , y6598 , y6599 , y6600 , y6601 , y6602 , y6603 , y6604 , y6605 , y6606 , y6607 , y6608 , y6609 , y6610 , y6611 , y6612 , y6613 , y6614 , y6615 , y6616 , y6617 , y6618 , y6619 , y6620 , y6621 , y6622 , y6623 , y6624 , y6625 , y6626 , y6627 , y6628 , y6629 , y6630 , y6631 , y6632 , y6633 , y6634 , y6635 , y6636 , y6637 , y6638 , y6639 , y6640 , y6641 , y6642 , y6643 , y6644 , y6645 , y6646 , y6647 , y6648 , y6649 , y6650 , y6651 , y6652 , y6653 , y6654 , y6655 , y6656 , y6657 , y6658 , y6659 , y6660 , y6661 , y6662 , y6663 , y6664 , y6665 , y6666 , y6667 , y6668 , y6669 , y6670 , y6671 , y6672 , y6673 , y6674 , y6675 , y6676 , y6677 , y6678 , y6679 , y6680 , y6681 , y6682 , y6683 , y6684 , y6685 , y6686 , y6687 , y6688 , y6689 , y6690 , y6691 , y6692 , y6693 , y6694 , y6695 , y6696 , y6697 , y6698 , y6699 , y6700 , y6701 , y6702 , y6703 , y6704 , y6705 , y6706 , y6707 , y6708 , y6709 , y6710 , y6711 , y6712 , y6713 , y6714 , y6715 , y6716 , y6717 , y6718 , y6719 , y6720 , y6721 , y6722 , y6723 , y6724 , y6725 , y6726 , y6727 , y6728 , y6729 , y6730 , y6731 , y6732 , y6733 , y6734 , y6735 , y6736 , y6737 , y6738 , y6739 , y6740 , y6741 , y6742 , y6743 , y6744 , y6745 , y6746 , y6747 , y6748 , y6749 , y6750 , y6751 , y6752 , y6753 , y6754 , y6755 , y6756 , y6757 , y6758 , y6759 , y6760 , y6761 , y6762 , y6763 , y6764 , y6765 , y6766 , y6767 , y6768 , y6769 , y6770 , y6771 , y6772 , y6773 , y6774 , y6775 , y6776 , y6777 , y6778 , y6779 , y6780 , y6781 , y6782 , y6783 , y6784 , y6785 , y6786 , y6787 , y6788 , y6789 , y6790 , y6791 , y6792 , y6793 , y6794 , y6795 , y6796 , y6797 , y6798 , y6799 , y6800 , y6801 , y6802 , y6803 , y6804 , y6805 , y6806 , y6807 , y6808 , y6809 , y6810 , y6811 , y6812 , y6813 , y6814 , y6815 , y6816 , y6817 , y6818 , y6819 , y6820 , y6821 , y6822 , y6823 , y6824 , y6825 , y6826 , y6827 , y6828 , y6829 , y6830 , y6831 , y6832 , y6833 , y6834 , y6835 , y6836 , y6837 , y6838 , y6839 , y6840 , y6841 , y6842 , y6843 , y6844 , y6845 , y6846 , y6847 , y6848 , y6849 , y6850 , y6851 , y6852 , y6853 , y6854 , y6855 , y6856 , y6857 , y6858 , y6859 , y6860 , y6861 , y6862 , y6863 , y6864 , y6865 , y6866 , y6867 , y6868 , y6869 , y6870 , y6871 , y6872 , y6873 , y6874 , y6875 , y6876 , y6877 , y6878 , y6879 , y6880 , y6881 , y6882 , y6883 , y6884 , y6885 , y6886 , y6887 , y6888 , y6889 , y6890 , y6891 , y6892 , y6893 , y6894 , y6895 , y6896 , y6897 , y6898 , y6899 , y6900 , y6901 , y6902 , y6903 , y6904 , y6905 , y6906 , y6907 , y6908 , y6909 , y6910 , y6911 , y6912 , y6913 , y6914 , y6915 , y6916 , y6917 , y6918 , y6919 , y6920 , y6921 , y6922 , y6923 , y6924 , y6925 , y6926 , y6927 , y6928 , y6929 , y6930 , y6931 , y6932 , y6933 , y6934 , y6935 , y6936 , y6937 , y6938 , y6939 , y6940 , y6941 , y6942 , y6943 , y6944 , y6945 , y6946 , y6947 , y6948 , y6949 , y6950 , y6951 , y6952 , y6953 , y6954 , y6955 , y6956 , y6957 , y6958 , y6959 , y6960 , y6961 , y6962 , y6963 , y6964 , y6965 , y6966 , y6967 , y6968 , y6969 , y6970 , y6971 , y6972 , y6973 , y6974 , y6975 , y6976 , y6977 , y6978 , y6979 , y6980 , y6981 , y6982 , y6983 , y6984 , y6985 , y6986 , y6987 , y6988 , y6989 , y6990 , y6991 , y6992 , y6993 , y6994 , y6995 , y6996 , y6997 , y6998 , y6999 , y7000 , y7001 , y7002 , y7003 , y7004 , y7005 , y7006 , y7007 , y7008 , y7009 , y7010 , y7011 , y7012 , y7013 , y7014 , y7015 , y7016 , y7017 , y7018 , y7019 , y7020 , y7021 , y7022 , y7023 , y7024 , y7025 , y7026 , y7027 , y7028 , y7029 , y7030 , y7031 , y7032 , y7033 , y7034 , y7035 , y7036 , y7037 , y7038 , y7039 , y7040 , y7041 , y7042 , y7043 , y7044 , y7045 , y7046 , y7047 , y7048 , y7049 , y7050 , y7051 , y7052 , y7053 , y7054 , y7055 , y7056 , y7057 , y7058 , y7059 , y7060 , y7061 , y7062 , y7063 , y7064 , y7065 , y7066 , y7067 , y7068 , y7069 , y7070 , y7071 , y7072 , y7073 , y7074 , y7075 , y7076 , y7077 , y7078 , y7079 , y7080 , y7081 , y7082 , y7083 , y7084 , y7085 , y7086 , y7087 , y7088 , y7089 , y7090 , y7091 , y7092 , y7093 , y7094 , y7095 , y7096 , y7097 , y7098 , y7099 , y7100 , y7101 , y7102 , y7103 , y7104 , y7105 , y7106 , y7107 , y7108 , y7109 , y7110 , y7111 , y7112 , y7113 , y7114 , y7115 , y7116 , y7117 , y7118 , y7119 , y7120 , y7121 , y7122 , y7123 , y7124 , y7125 , y7126 , y7127 , y7128 , y7129 , y7130 , y7131 , y7132 , y7133 , y7134 , y7135 , y7136 , y7137 , y7138 , y7139 , y7140 , y7141 , y7142 , y7143 , y7144 , y7145 , y7146 , y7147 , y7148 , y7149 , y7150 , y7151 , y7152 , y7153 , y7154 , y7155 , y7156 , y7157 , y7158 , y7159 , y7160 , y7161 , y7162 , y7163 , y7164 , y7165 , y7166 , y7167 , y7168 , y7169 , y7170 , y7171 , y7172 , y7173 , y7174 , y7175 , y7176 , y7177 , y7178 , y7179 , y7180 , y7181 , y7182 , y7183 , y7184 , y7185 , y7186 , y7187 , y7188 , y7189 , y7190 , y7191 , y7192 , y7193 , y7194 , y7195 , y7196 , y7197 , y7198 , y7199 , y7200 , y7201 , y7202 , y7203 , y7204 , y7205 , y7206 , y7207 , y7208 , y7209 , y7210 , y7211 , y7212 , y7213 , y7214 , y7215 , y7216 , y7217 , y7218 , y7219 , y7220 , y7221 , y7222 , y7223 , y7224 , y7225 , y7226 , y7227 , y7228 , y7229 , y7230 , y7231 , y7232 , y7233 , y7234 , y7235 , y7236 , y7237 , y7238 , y7239 , y7240 , y7241 , y7242 , y7243 , y7244 , y7245 , y7246 , y7247 , y7248 , y7249 , y7250 , y7251 , y7252 , y7253 , y7254 , y7255 , y7256 , y7257 , y7258 , y7259 , y7260 , y7261 , y7262 , y7263 , y7264 , y7265 , y7266 , y7267 , y7268 , y7269 , y7270 , y7271 , y7272 , y7273 , y7274 , y7275 , y7276 , y7277 , y7278 , y7279 , y7280 , y7281 , y7282 , y7283 , y7284 , y7285 , y7286 , y7287 , y7288 , y7289 , y7290 , y7291 , y7292 , y7293 , y7294 , y7295 , y7296 , y7297 , y7298 , y7299 , y7300 , y7301 , y7302 , y7303 , y7304 , y7305 , y7306 , y7307 , y7308 , y7309 , y7310 , y7311 , y7312 , y7313 , y7314 , y7315 , y7316 , y7317 , y7318 , y7319 , y7320 , y7321 , y7322 , y7323 , y7324 , y7325 , y7326 , y7327 , y7328 , y7329 , y7330 , y7331 , y7332 , y7333 , y7334 , y7335 , y7336 , y7337 , y7338 , y7339 , y7340 , y7341 , y7342 , y7343 , y7344 , y7345 , y7346 , y7347 , y7348 , y7349 , y7350 , y7351 , y7352 , y7353 , y7354 , y7355 , y7356 , y7357 , y7358 , y7359 , y7360 , y7361 , y7362 , y7363 , y7364 , y7365 , y7366 , y7367 , y7368 , y7369 , y7370 , y7371 , y7372 , y7373 , y7374 , y7375 , y7376 , y7377 , y7378 , y7379 , y7380 , y7381 , y7382 , y7383 , y7384 , y7385 , y7386 , y7387 , y7388 , y7389 , y7390 , y7391 , y7392 , y7393 , y7394 , y7395 , y7396 , y7397 , y7398 , y7399 , y7400 , y7401 , y7402 , y7403 , y7404 , y7405 , y7406 , y7407 , y7408 , y7409 , y7410 , y7411 , y7412 , y7413 , y7414 , y7415 , y7416 , y7417 , y7418 , y7419 , y7420 , y7421 , y7422 , y7423 , y7424 , y7425 , y7426 , y7427 , y7428 , y7429 , y7430 , y7431 , y7432 , y7433 , y7434 , y7435 , y7436 , y7437 , y7438 , y7439 , y7440 , y7441 , y7442 , y7443 , y7444 , y7445 , y7446 , y7447 , y7448 , y7449 , y7450 , y7451 , y7452 , y7453 , y7454 , y7455 , y7456 , y7457 , y7458 , y7459 , y7460 , y7461 , y7462 , y7463 , y7464 , y7465 , y7466 , y7467 , y7468 , y7469 , y7470 , y7471 , y7472 , y7473 , y7474 , y7475 , y7476 , y7477 , y7478 , y7479 , y7480 , y7481 , y7482 , y7483 , y7484 , y7485 , y7486 , y7487 , y7488 , y7489 , y7490 , y7491 , y7492 , y7493 , y7494 , y7495 , y7496 , y7497 , y7498 , y7499 , y7500 , y7501 , y7502 , y7503 , y7504 , y7505 , y7506 , y7507 , y7508 , y7509 , y7510 , y7511 , y7512 , y7513 , y7514 , y7515 , y7516 , y7517 , y7518 , y7519 , y7520 , y7521 , y7522 , y7523 , y7524 , y7525 , y7526 , y7527 , y7528 , y7529 , y7530 , y7531 , y7532 , y7533 , y7534 , y7535 , y7536 , y7537 , y7538 , y7539 , y7540 , y7541 , y7542 , y7543 , y7544 , y7545 , y7546 , y7547 , y7548 , y7549 , y7550 , y7551 , y7552 , y7553 , y7554 , y7555 , y7556 , y7557 , y7558 , y7559 , y7560 , y7561 , y7562 , y7563 , y7564 , y7565 , y7566 , y7567 , y7568 , y7569 , y7570 , y7571 , y7572 , y7573 , y7574 , y7575 , y7576 , y7577 , y7578 , y7579 , y7580 , y7581 , y7582 , y7583 , y7584 , y7585 , y7586 , y7587 , y7588 , y7589 , y7590 , y7591 , y7592 , y7593 , y7594 , y7595 , y7596 , y7597 , y7598 , y7599 , y7600 , y7601 , y7602 , y7603 , y7604 , y7605 , y7606 , y7607 , y7608 , y7609 , y7610 , y7611 , y7612 , y7613 , y7614 , y7615 , y7616 , y7617 , y7618 , y7619 , y7620 , y7621 , y7622 , y7623 , y7624 , y7625 , y7626 , y7627 , y7628 , y7629 , y7630 , y7631 , y7632 , y7633 , y7634 , y7635 , y7636 , y7637 , y7638 , y7639 , y7640 , y7641 , y7642 , y7643 , y7644 , y7645 , y7646 , y7647 , y7648 , y7649 , y7650 , y7651 , y7652 , y7653 , y7654 , y7655 , y7656 , y7657 , y7658 , y7659 , y7660 , y7661 , y7662 , y7663 , y7664 , y7665 , y7666 , y7667 , y7668 , y7669 , y7670 , y7671 , y7672 , y7673 , y7674 , y7675 , y7676 , y7677 , y7678 , y7679 , y7680 , y7681 , y7682 , y7683 , y7684 , y7685 , y7686 , y7687 , y7688 , y7689 , y7690 , y7691 , y7692 , y7693 , y7694 , y7695 , y7696 , y7697 , y7698 , y7699 , y7700 , y7701 , y7702 , y7703 , y7704 , y7705 , y7706 , y7707 , y7708 , y7709 , y7710 , y7711 , y7712 , y7713 , y7714 , y7715 , y7716 , y7717 , y7718 , y7719 , y7720 , y7721 , y7722 , y7723 , y7724 , y7725 , y7726 , y7727 , y7728 , y7729 , y7730 , y7731 , y7732 , y7733 , y7734 , y7735 , y7736 , y7737 , y7738 , y7739 , y7740 , y7741 , y7742 , y7743 , y7744 , y7745 , y7746 , y7747 , y7748 , y7749 , y7750 , y7751 , y7752 , y7753 , y7754 , y7755 , y7756 , y7757 , y7758 , y7759 , y7760 , y7761 , y7762 , y7763 , y7764 , y7765 , y7766 , y7767 , y7768 , y7769 , y7770 , y7771 , y7772 , y7773 , y7774 , y7775 , y7776 , y7777 , y7778 , y7779 , y7780 , y7781 , y7782 , y7783 , y7784 , y7785 , y7786 , y7787 , y7788 , y7789 , y7790 , y7791 , y7792 , y7793 , y7794 , y7795 , y7796 , y7797 , y7798 , y7799 , y7800 , y7801 , y7802 , y7803 , y7804 , y7805 , y7806 , y7807 , y7808 , y7809 , y7810 , y7811 , y7812 , y7813 , y7814 , y7815 , y7816 , y7817 , y7818 , y7819 , y7820 , y7821 , y7822 , y7823 , y7824 , y7825 , y7826 , y7827 , y7828 , y7829 , y7830 , y7831 , y7832 , y7833 , y7834 , y7835 , y7836 , y7837 , y7838 , y7839 , y7840 , y7841 , y7842 , y7843 , y7844 , y7845 , y7846 , y7847 , y7848 , y7849 , y7850 , y7851 , y7852 , y7853 , y7854 , y7855 , y7856 , y7857 , y7858 , y7859 , y7860 , y7861 , y7862 , y7863 , y7864 , y7865 , y7866 , y7867 , y7868 , y7869 , y7870 , y7871 , y7872 , y7873 , y7874 , y7875 , y7876 , y7877 , y7878 , y7879 , y7880 , y7881 , y7882 , y7883 , y7884 , y7885 , y7886 , y7887 , y7888 , y7889 , y7890 , y7891 , y7892 , y7893 , y7894 , y7895 , y7896 , y7897 , y7898 , y7899 , y7900 , y7901 , y7902 , y7903 , y7904 , y7905 , y7906 , y7907 , y7908 , y7909 , y7910 , y7911 , y7912 , y7913 , y7914 , y7915 , y7916 , y7917 , y7918 , y7919 , y7920 , y7921 , y7922 , y7923 , y7924 , y7925 , y7926 , y7927 , y7928 , y7929 , y7930 , y7931 , y7932 , y7933 , y7934 , y7935 , y7936 , y7937 , y7938 , y7939 , y7940 , y7941 , y7942 , y7943 , y7944 , y7945 , y7946 , y7947 , y7948 , y7949 , y7950 , y7951 , y7952 , y7953 , y7954 , y7955 , y7956 , y7957 , y7958 , y7959 , y7960 , y7961 , y7962 , y7963 , y7964 , y7965 , y7966 , y7967 , y7968 , y7969 , y7970 , y7971 , y7972 , y7973 , y7974 , y7975 , y7976 , y7977 , y7978 , y7979 , y7980 , y7981 , y7982 , y7983 , y7984 , y7985 , y7986 , y7987 , y7988 , y7989 , y7990 , y7991 , y7992 , y7993 , y7994 , y7995 , y7996 , y7997 , y7998 , y7999 , y8000 , y8001 , y8002 , y8003 , y8004 , y8005 , y8006 , y8007 , y8008 , y8009 , y8010 , y8011 , y8012 , y8013 , y8014 , y8015 , y8016 , y8017 , y8018 , y8019 , y8020 , y8021 , y8022 , y8023 , y8024 , y8025 , y8026 , y8027 , y8028 , y8029 , y8030 , y8031 , y8032 , y8033 , y8034 , y8035 , y8036 , y8037 , y8038 , y8039 , y8040 , y8041 , y8042 , y8043 , y8044 , y8045 , y8046 , y8047 , y8048 , y8049 , y8050 , y8051 , y8052 , y8053 , y8054 , y8055 , y8056 , y8057 , y8058 , y8059 , y8060 , y8061 , y8062 , y8063 , y8064 , y8065 , y8066 , y8067 , y8068 , y8069 , y8070 , y8071 , y8072 , y8073 , y8074 , y8075 , y8076 , y8077 , y8078 , y8079 , y8080 , y8081 , y8082 , y8083 , y8084 , y8085 , y8086 , y8087 , y8088 , y8089 , y8090 , y8091 , y8092 , y8093 , y8094 , y8095 , y8096 , y8097 , y8098 , y8099 , y8100 , y8101 , y8102 , y8103 , y8104 , y8105 , y8106 , y8107 , y8108 , y8109 , y8110 , y8111 , y8112 , y8113 , y8114 , y8115 , y8116 , y8117 , y8118 , y8119 , y8120 , y8121 , y8122 , y8123 , y8124 , y8125 , y8126 , y8127 , y8128 , y8129 , y8130 , y8131 , y8132 , y8133 , y8134 , y8135 , y8136 , y8137 , y8138 , y8139 , y8140 , y8141 , y8142 , y8143 , y8144 , y8145 , y8146 , y8147 , y8148 , y8149 , y8150 , y8151 , y8152 , y8153 , y8154 , y8155 , y8156 , y8157 , y8158 , y8159 , y8160 , y8161 , y8162 , y8163 , y8164 , y8165 , y8166 , y8167 , y8168 , y8169 , y8170 , y8171 , y8172 , y8173 , y8174 , y8175 , y8176 , y8177 , y8178 , y8179 , y8180 , y8181 , y8182 , y8183 , y8184 , y8185 , y8186 , y8187 , y8188 , y8189 , y8190 , y8191 , y8192 , y8193 , y8194 , y8195 , y8196 , y8197 , y8198 , y8199 , y8200 , y8201 , y8202 , y8203 , y8204 , y8205 , y8206 , y8207 , y8208 , y8209 , y8210 , y8211 , y8212 , y8213 , y8214 , y8215 , y8216 , y8217 , y8218 , y8219 , y8220 , y8221 , y8222 , y8223 , y8224 , y8225 , y8226 , y8227 , y8228 , y8229 , y8230 , y8231 , y8232 , y8233 , y8234 , y8235 , y8236 , y8237 , y8238 , y8239 , y8240 , y8241 , y8242 , y8243 , y8244 , y8245 , y8246 , y8247 , y8248 , y8249 , y8250 , y8251 , y8252 , y8253 , y8254 , y8255 , y8256 , y8257 , y8258 , y8259 , y8260 , y8261 , y8262 , y8263 , y8264 , y8265 , y8266 , y8267 , y8268 , y8269 , y8270 , y8271 , y8272 , y8273 , y8274 , y8275 , y8276 , y8277 , y8278 , y8279 , y8280 , y8281 , y8282 , y8283 , y8284 , y8285 , y8286 , y8287 , y8288 , y8289 , y8290 , y8291 , y8292 , y8293 , y8294 , y8295 , y8296 , y8297 , y8298 , y8299 , y8300 , y8301 , y8302 , y8303 , y8304 , y8305 , y8306 , y8307 , y8308 , y8309 , y8310 , y8311 , y8312 , y8313 , y8314 , y8315 , y8316 , y8317 , y8318 , y8319 , y8320 , y8321 , y8322 , y8323 , y8324 , y8325 , y8326 , y8327 , y8328 , y8329 , y8330 , y8331 , y8332 , y8333 , y8334 , y8335 , y8336 , y8337 , y8338 , y8339 , y8340 , y8341 , y8342 , y8343 , y8344 , y8345 , y8346 , y8347 , y8348 , y8349 , y8350 , y8351 , y8352 , y8353 , y8354 , y8355 , y8356 , y8357 , y8358 , y8359 , y8360 , y8361 , y8362 , y8363 , y8364 , y8365 , y8366 , y8367 , y8368 , y8369 , y8370 , y8371 , y8372 , y8373 , y8374 , y8375 , y8376 , y8377 , y8378 , y8379 , y8380 , y8381 , y8382 , y8383 , y8384 , y8385 , y8386 , y8387 , y8388 , y8389 , y8390 , y8391 , y8392 , y8393 , y8394 , y8395 , y8396 , y8397 , y8398 , y8399 , y8400 , y8401 , y8402 , y8403 , y8404 , y8405 , y8406 , y8407 , y8408 , y8409 , y8410 , y8411 , y8412 , y8413 , y8414 , y8415 , y8416 , y8417 , y8418 , y8419 , y8420 , y8421 , y8422 , y8423 , y8424 , y8425 , y8426 , y8427 , y8428 , y8429 , y8430 , y8431 , y8432 , y8433 , y8434 , y8435 , y8436 , y8437 , y8438 , y8439 , y8440 , y8441 , y8442 , y8443 , y8444 , y8445 , y8446 , y8447 , y8448 , y8449 , y8450 , y8451 , y8452 , y8453 , y8454 , y8455 , y8456 , y8457 , y8458 , y8459 , y8460 , y8461 , y8462 , y8463 , y8464 , y8465 , y8466 , y8467 , y8468 , y8469 , y8470 , y8471 , y8472 , y8473 , y8474 , y8475 , y8476 , y8477 , y8478 , y8479 , y8480 , y8481 , y8482 , y8483 , y8484 , y8485 , y8486 , y8487 , y8488 , y8489 , y8490 , y8491 , y8492 , y8493 , y8494 , y8495 , y8496 , y8497 , y8498 , y8499 , y8500 , y8501 , y8502 , y8503 , y8504 , y8505 , y8506 , y8507 , y8508 , y8509 , y8510 , y8511 , y8512 , y8513 , y8514 , y8515 , y8516 , y8517 , y8518 , y8519 , y8520 , y8521 , y8522 , y8523 , y8524 , y8525 , y8526 , y8527 , y8528 , y8529 , y8530 , y8531 , y8532 , y8533 , y8534 , y8535 , y8536 , y8537 , y8538 , y8539 , y8540 , y8541 , y8542 , y8543 , y8544 , y8545 , y8546 , y8547 , y8548 , y8549 , y8550 , y8551 , y8552 , y8553 , y8554 , y8555 , y8556 , y8557 , y8558 , y8559 , y8560 , y8561 , y8562 , y8563 , y8564 , y8565 , y8566 , y8567 , y8568 , y8569 , y8570 , y8571 , y8572 , y8573 , y8574 , y8575 , y8576 , y8577 , y8578 , y8579 , y8580 , y8581 , y8582 , y8583 , y8584 , y8585 , y8586 , y8587 , y8588 , y8589 , y8590 , y8591 , y8592 , y8593 , y8594 , y8595 , y8596 , y8597 , y8598 , y8599 , y8600 , y8601 , y8602 , y8603 , y8604 , y8605 , y8606 , y8607 , y8608 , y8609 , y8610 , y8611 , y8612 , y8613 , y8614 , y8615 , y8616 , y8617 , y8618 , y8619 , y8620 , y8621 , y8622 , y8623 , y8624 , y8625 , y8626 , y8627 , y8628 , y8629 , y8630 , y8631 , y8632 , y8633 , y8634 , y8635 , y8636 , y8637 , y8638 , y8639 , y8640 , y8641 , y8642 , y8643 , y8644 , y8645 , y8646 , y8647 , y8648 , y8649 , y8650 , y8651 , y8652 , y8653 , y8654 , y8655 , y8656 , y8657 , y8658 , y8659 , y8660 , y8661 , y8662 , y8663 , y8664 , y8665 , y8666 , y8667 , y8668 , y8669 , y8670 , y8671 , y8672 , y8673 , y8674 , y8675 , y8676 , y8677 , y8678 , y8679 , y8680 , y8681 , y8682 , y8683 , y8684 , y8685 , y8686 , y8687 , y8688 , y8689 , y8690 , y8691 , y8692 , y8693 , y8694 , y8695 , y8696 , y8697 , y8698 , y8699 , y8700 , y8701 , y8702 , y8703 , y8704 , y8705 , y8706 , y8707 , y8708 , y8709 , y8710 , y8711 , y8712 , y8713 , y8714 , y8715 , y8716 , y8717 , y8718 , y8719 , y8720 , y8721 , y8722 , y8723 , y8724 , y8725 , y8726 , y8727 , y8728 , y8729 , y8730 , y8731 , y8732 , y8733 , y8734 , y8735 , y8736 , y8737 , y8738 , y8739 , y8740 , y8741 , y8742 , y8743 , y8744 , y8745 , y8746 , y8747 , y8748 , y8749 , y8750 , y8751 , y8752 , y8753 , y8754 , y8755 , y8756 , y8757 , y8758 , y8759 , y8760 , y8761 , y8762 , y8763 , y8764 , y8765 , y8766 , y8767 , y8768 , y8769 , y8770 , y8771 , y8772 , y8773 , y8774 , y8775 , y8776 , y8777 , y8778 , y8779 , y8780 , y8781 , y8782 , y8783 , y8784 , y8785 , y8786 , y8787 , y8788 , y8789 , y8790 , y8791 , y8792 , y8793 , y8794 , y8795 , y8796 , y8797 , y8798 , y8799 , y8800 , y8801 , y8802 , y8803 , y8804 , y8805 , y8806 , y8807 , y8808 , y8809 , y8810 , y8811 , y8812 , y8813 , y8814 , y8815 , y8816 , y8817 , y8818 , y8819 , y8820 , y8821 , y8822 , y8823 , y8824 , y8825 , y8826 , y8827 , y8828 , y8829 , y8830 , y8831 , y8832 , y8833 , y8834 , y8835 , y8836 , y8837 , y8838 , y8839 , y8840 , y8841 , y8842 , y8843 , y8844 , y8845 , y8846 , y8847 , y8848 , y8849 , y8850 , y8851 , y8852 , y8853 , y8854 , y8855 , y8856 , y8857 , y8858 , y8859 , y8860 , y8861 , y8862 , y8863 , y8864 , y8865 , y8866 , y8867 , y8868 , y8869 , y8870 , y8871 , y8872 , y8873 , y8874 , y8875 , y8876 , y8877 , y8878 , y8879 , y8880 , y8881 , y8882 , y8883 , y8884 , y8885 , y8886 , y8887 , y8888 , y8889 , y8890 , y8891 , y8892 , y8893 , y8894 , y8895 , y8896 , y8897 , y8898 , y8899 , y8900 , y8901 , y8902 , y8903 , y8904 , y8905 , y8906 , y8907 , y8908 , y8909 , y8910 , y8911 , y8912 , y8913 , y8914 , y8915 , y8916 , y8917 , y8918 , y8919 , y8920 , y8921 , y8922 , y8923 , y8924 , y8925 , y8926 , y8927 , y8928 , y8929 , y8930 , y8931 , y8932 , y8933 , y8934 , y8935 , y8936 , y8937 , y8938 , y8939 , y8940 , y8941 , y8942 , y8943 , y8944 , y8945 , y8946 , y8947 , y8948 , y8949 , y8950 , y8951 , y8952 , y8953 , y8954 , y8955 , y8956 , y8957 , y8958 , y8959 , y8960 , y8961 , y8962 , y8963 , y8964 , y8965 , y8966 , y8967 , y8968 , y8969 , y8970 , y8971 , y8972 , y8973 , y8974 , y8975 , y8976 , y8977 , y8978 , y8979 , y8980 , y8981 , y8982 , y8983 , y8984 , y8985 , y8986 , y8987 , y8988 , y8989 , y8990 , y8991 , y8992 , y8993 , y8994 , y8995 , y8996 , y8997 , y8998 , y8999 , y9000 , y9001 , y9002 , y9003 , y9004 , y9005 , y9006 , y9007 , y9008 , y9009 , y9010 , y9011 , y9012 , y9013 , y9014 , y9015 , y9016 , y9017 , y9018 , y9019 , y9020 , y9021 , y9022 , y9023 , y9024 , y9025 , y9026 , y9027 , y9028 , y9029 , y9030 , y9031 , y9032 , y9033 , y9034 , y9035 , y9036 , y9037 , y9038 , y9039 , y9040 , y9041 , y9042 , y9043 , y9044 , y9045 , y9046 , y9047 , y9048 , y9049 , y9050 , y9051 , y9052 , y9053 , y9054 , y9055 , y9056 , y9057 , y9058 , y9059 , y9060 , y9061 , y9062 , y9063 , y9064 , y9065 , y9066 , y9067 , y9068 , y9069 , y9070 , y9071 , y9072 , y9073 , y9074 , y9075 , y9076 , y9077 , y9078 , y9079 , y9080 , y9081 , y9082 , y9083 , y9084 , y9085 , y9086 , y9087 , y9088 , y9089 , y9090 , y9091 , y9092 , y9093 , y9094 , y9095 , y9096 , y9097 , y9098 , y9099 , y9100 , y9101 , y9102 , y9103 , y9104 , y9105 , y9106 , y9107 , y9108 , y9109 , y9110 , y9111 , y9112 , y9113 , y9114 , y9115 , y9116 , y9117 , y9118 , y9119 , y9120 , y9121 , y9122 , y9123 , y9124 , y9125 , y9126 , y9127 , y9128 , y9129 , y9130 , y9131 , y9132 , y9133 , y9134 , y9135 , y9136 , y9137 , y9138 , y9139 , y9140 , y9141 , y9142 , y9143 , y9144 , y9145 , y9146 , y9147 , y9148 , y9149 , y9150 , y9151 , y9152 , y9153 , y9154 , y9155 , y9156 , y9157 , y9158 , y9159 , y9160 , y9161 , y9162 , y9163 , y9164 , y9165 , y9166 , y9167 , y9168 , y9169 , y9170 , y9171 , y9172 , y9173 , y9174 , y9175 , y9176 , y9177 , y9178 , y9179 , y9180 , y9181 , y9182 , y9183 , y9184 , y9185 , y9186 , y9187 , y9188 , y9189 , y9190 , y9191 , y9192 , y9193 , y9194 , y9195 , y9196 , y9197 , y9198 , y9199 , y9200 , y9201 , y9202 , y9203 , y9204 , y9205 , y9206 , y9207 , y9208 , y9209 , y9210 , y9211 , y9212 , y9213 , y9214 , y9215 , y9216 , y9217 , y9218 , y9219 , y9220 , y9221 , y9222 , y9223 , y9224 , y9225 , y9226 , y9227 , y9228 , y9229 , y9230 , y9231 , y9232 , y9233 , y9234 , y9235 , y9236 , y9237 , y9238 , y9239 , y9240 , y9241 , y9242 , y9243 , y9244 , y9245 , y9246 , y9247 , y9248 , y9249 , y9250 , y9251 , y9252 , y9253 , y9254 , y9255 , y9256 , y9257 , y9258 , y9259 , y9260 , y9261 , y9262 , y9263 , y9264 , y9265 , y9266 , y9267 , y9268 , y9269 , y9270 , y9271 , y9272 , y9273 , y9274 , y9275 , y9276 , y9277 , y9278 , y9279 , y9280 , y9281 , y9282 , y9283 , y9284 , y9285 , y9286 , y9287 , y9288 , y9289 , y9290 , y9291 , y9292 , y9293 , y9294 , y9295 , y9296 , y9297 , y9298 , y9299 , y9300 , y9301 , y9302 , y9303 , y9304 , y9305 , y9306 , y9307 , y9308 , y9309 , y9310 , y9311 , y9312 , y9313 , y9314 , y9315 , y9316 , y9317 , y9318 , y9319 , y9320 , y9321 , y9322 , y9323 , y9324 , y9325 , y9326 , y9327 , y9328 , y9329 , y9330 , y9331 , y9332 , y9333 , y9334 , y9335 , y9336 , y9337 , y9338 , y9339 , y9340 , y9341 , y9342 , y9343 , y9344 , y9345 , y9346 , y9347 , y9348 , y9349 , y9350 , y9351 , y9352 , y9353 , y9354 , y9355 , y9356 , y9357 , y9358 , y9359 , y9360 , y9361 , y9362 , y9363 , y9364 , y9365 , y9366 , y9367 , y9368 , y9369 , y9370 , y9371 , y9372 , y9373 , y9374 , y9375 , y9376 , y9377 , y9378 , y9379 , y9380 , y9381 , y9382 , y9383 , y9384 , y9385 , y9386 , y9387 , y9388 , y9389 , y9390 , y9391 , y9392 , y9393 , y9394 , y9395 , y9396 , y9397 , y9398 , y9399 , y9400 , y9401 , y9402 , y9403 , y9404 , y9405 , y9406 , y9407 , y9408 , y9409 , y9410 , y9411 , y9412 , y9413 , y9414 , y9415 , y9416 , y9417 , y9418 , y9419 , y9420 , y9421 , y9422 , y9423 , y9424 , y9425 , y9426 , y9427 , y9428 , y9429 , y9430 , y9431 , y9432 , y9433 , y9434 , y9435 , y9436 , y9437 , y9438 , y9439 , y9440 , y9441 , y9442 , y9443 , y9444 , y9445 , y9446 , y9447 , y9448 , y9449 , y9450 , y9451 , y9452 , y9453 , y9454 , y9455 , y9456 , y9457 , y9458 , y9459 , y9460 , y9461 , y9462 , y9463 , y9464 , y9465 , y9466 , y9467 , y9468 , y9469 , y9470 , y9471 , y9472 , y9473 , y9474 , y9475 , y9476 , y9477 , y9478 , y9479 , y9480 , y9481 , y9482 , y9483 , y9484 , y9485 , y9486 , y9487 , y9488 , y9489 , y9490 , y9491 , y9492 , y9493 , y9494 , y9495 , y9496 , y9497 , y9498 , y9499 , y9500 , y9501 , y9502 , y9503 , y9504 , y9505 , y9506 , y9507 , y9508 , y9509 , y9510 , y9511 , y9512 , y9513 , y9514 , y9515 , y9516 , y9517 , y9518 , y9519 , y9520 , y9521 , y9522 , y9523 , y9524 , y9525 , y9526 , y9527 , y9528 , y9529 , y9530 , y9531 , y9532 , y9533 , y9534 , y9535 , y9536 , y9537 , y9538 , y9539 , y9540 , y9541 , y9542 , y9543 , y9544 , y9545 , y9546 , y9547 , y9548 , y9549 , y9550 , y9551 , y9552 , y9553 , y9554 , y9555 , y9556 , y9557 , y9558 , y9559 , y9560 , y9561 , y9562 , y9563 , y9564 , y9565 , y9566 , y9567 , y9568 , y9569 , y9570 , y9571 , y9572 , y9573 , y9574 , y9575 , y9576 , y9577 , y9578 , y9579 , y9580 , y9581 , y9582 , y9583 , y9584 , y9585 , y9586 , y9587 , y9588 , y9589 , y9590 , y9591 , y9592 , y9593 , y9594 , y9595 , y9596 , y9597 , y9598 , y9599 , y9600 , y9601 , y9602 , y9603 , y9604 , y9605 , y9606 , y9607 , y9608 , y9609 , y9610 , y9611 , y9612 , y9613 , y9614 , y9615 , y9616 , y9617 , y9618 , y9619 , y9620 , y9621 , y9622 , y9623 , y9624 , y9625 , y9626 , y9627 , y9628 , y9629 , y9630 , y9631 , y9632 , y9633 , y9634 , y9635 , y9636 , y9637 , y9638 , y9639 , y9640 , y9641 , y9642 , y9643 , y9644 , y9645 , y9646 , y9647 , y9648 , y9649 , y9650 , y9651 , y9652 , y9653 , y9654 , y9655 , y9656 , y9657 , y9658 , y9659 , y9660 , y9661 , y9662 , y9663 , y9664 , y9665 , y9666 , y9667 , y9668 , y9669 , y9670 , y9671 , y9672 , y9673 , y9674 , y9675 , y9676 , y9677 , y9678 , y9679 , y9680 , y9681 , y9682 , y9683 , y9684 , y9685 , y9686 , y9687 , y9688 , y9689 , y9690 , y9691 , y9692 , y9693 , y9694 , y9695 , y9696 , y9697 , y9698 , y9699 , y9700 , y9701 , y9702 , y9703 , y9704 , y9705 , y9706 , y9707 , y9708 , y9709 , y9710 , y9711 , y9712 , y9713 , y9714 , y9715 , y9716 , y9717 , y9718 , y9719 , y9720 , y9721 , y9722 , y9723 , y9724 , y9725 , y9726 , y9727 , y9728 , y9729 , y9730 , y9731 , y9732 , y9733 , y9734 , y9735 , y9736 , y9737 , y9738 , y9739 , y9740 , y9741 , y9742 , y9743 , y9744 , y9745 , y9746 , y9747 , y9748 , y9749 , y9750 , y9751 , y9752 , y9753 , y9754 , y9755 , y9756 , y9757 , y9758 , y9759 , y9760 , y9761 , y9762 , y9763 , y9764 , y9765 , y9766 , y9767 , y9768 , y9769 , y9770 , y9771 , y9772 , y9773 , y9774 , y9775 , y9776 , y9777 , y9778 , y9779 , y9780 , y9781 , y9782 , y9783 , y9784 , y9785 , y9786 , y9787 , y9788 , y9789 , y9790 , y9791 , y9792 , y9793 , y9794 , y9795 , y9796 , y9797 , y9798 , y9799 , y9800 , y9801 , y9802 , y9803 , y9804 , y9805 , y9806 , y9807 , y9808 , y9809 , y9810 , y9811 , y9812 , y9813 , y9814 , y9815 , y9816 , y9817 , y9818 , y9819 , y9820 , y9821 , y9822 , y9823 , y9824 , y9825 , y9826 , y9827 , y9828 , y9829 , y9830 , y9831 , y9832 , y9833 , y9834 , y9835 , y9836 , y9837 , y9838 , y9839 , y9840 , y9841 , y9842 , y9843 , y9844 , y9845 , y9846 , y9847 , y9848 , y9849 , y9850 , y9851 , y9852 , y9853 , y9854 , y9855 , y9856 , y9857 , y9858 , y9859 , y9860 , y9861 , y9862 , y9863 , y9864 , y9865 , y9866 , y9867 , y9868 , y9869 , y9870 , y9871 , y9872 , y9873 , y9874 , y9875 , y9876 , y9877 , y9878 , y9879 , y9880 , y9881 , y9882 , y9883 , y9884 , y9885 , y9886 , y9887 , y9888 , y9889 , y9890 , y9891 , y9892 , y9893 , y9894 , y9895 , y9896 , y9897 , y9898 , y9899 , y9900 , y9901 , y9902 , y9903 , y9904 , y9905 , y9906 , y9907 , y9908 , y9909 , y9910 , y9911 , y9912 , y9913 , y9914 , y9915 , y9916 , y9917 , y9918 , y9919 , y9920 , y9921 , y9922 , y9923 , y9924 , y9925 , y9926 , y9927 , y9928 , y9929 , y9930 , y9931 , y9932 , y9933 , y9934 , y9935 , y9936 , y9937 , y9938 , y9939 , y9940 , y9941 , y9942 , y9943 , y9944 , y9945 , y9946 , y9947 , y9948 , y9949 , y9950 , y9951 , y9952 , y9953 , y9954 , y9955 , y9956 , y9957 , y9958 , y9959 , y9960 , y9961 , y9962 , y9963 , y9964 , y9965 , y9966 , y9967 , y9968 , y9969 , y9970 , y9971 , y9972 , y9973 , y9974 , y9975 , y9976 , y9977 , y9978 , y9979 , y9980 , y9981 , y9982 , y9983 , y9984 , y9985 , y9986 , y9987 , y9988 , y9989 , y9990 , y9991 , y9992 , y9993 , y9994 , y9995 , y9996 , y9997 , y9998 , y9999 , y10000 , y10001 , y10002 , y10003 , y10004 , y10005 , y10006 , y10007 , y10008 , y10009 , y10010 , y10011 , y10012 , y10013 , y10014 , y10015 , y10016 , y10017 , y10018 , y10019 , y10020 , y10021 , y10022 , y10023 , y10024 , y10025 , y10026 , y10027 , y10028 , y10029 , y10030 , y10031 , y10032 , y10033 , y10034 , y10035 , y10036 , y10037 , y10038 , y10039 , y10040 , y10041 , y10042 , y10043 , y10044 , y10045 , y10046 , y10047 , y10048 , y10049 , y10050 , y10051 , y10052 , y10053 , y10054 , y10055 , y10056 , y10057 , y10058 , y10059 , y10060 , y10061 , y10062 , y10063 , y10064 , y10065 , y10066 , y10067 , y10068 , y10069 , y10070 , y10071 , y10072 , y10073 , y10074 , y10075 , y10076 , y10077 , y10078 , y10079 , y10080 , y10081 , y10082 , y10083 , y10084 , y10085 , y10086 , y10087 , y10088 , y10089 , y10090 , y10091 , y10092 , y10093 , y10094 , y10095 , y10096 , y10097 , y10098 , y10099 , y10100 , y10101 , y10102 , y10103 , y10104 , y10105 , y10106 , y10107 , y10108 , y10109 , y10110 , y10111 , y10112 , y10113 , y10114 , y10115 , y10116 , y10117 , y10118 , y10119 , y10120 , y10121 , y10122 , y10123 , y10124 , y10125 , y10126 , y10127 , y10128 , y10129 , y10130 , y10131 , y10132 , y10133 , y10134 , y10135 , y10136 , y10137 , y10138 , y10139 , y10140 , y10141 , y10142 , y10143 , y10144 , y10145 , y10146 , y10147 , y10148 , y10149 , y10150 , y10151 , y10152 , y10153 , y10154 , y10155 , y10156 , y10157 , y10158 , y10159 , y10160 , y10161 , y10162 , y10163 , y10164 , y10165 , y10166 , y10167 , y10168 , y10169 , y10170 , y10171 , y10172 , y10173 , y10174 , y10175 , y10176 , y10177 , y10178 , y10179 , y10180 , y10181 , y10182 , y10183 , y10184 , y10185 , y10186 , y10187 , y10188 , y10189 , y10190 , y10191 , y10192 , y10193 , y10194 , y10195 , y10196 , y10197 , y10198 , y10199 , y10200 , y10201 , y10202 , y10203 , y10204 , y10205 , y10206 , y10207 , y10208 , y10209 , y10210 , y10211 , y10212 , y10213 , y10214 , y10215 , y10216 , y10217 , y10218 , y10219 , y10220 , y10221 , y10222 , y10223 , y10224 , y10225 , y10226 , y10227 , y10228 , y10229 , y10230 , y10231 , y10232 , y10233 , y10234 , y10235 , y10236 , y10237 , y10238 , y10239 , y10240 , y10241 , y10242 , y10243 , y10244 , y10245 , y10246 , y10247 , y10248 , y10249 , y10250 , y10251 , y10252 , y10253 , y10254 , y10255 , y10256 , y10257 , y10258 , y10259 , y10260 , y10261 , y10262 , y10263 , y10264 , y10265 , y10266 , y10267 , y10268 , y10269 , y10270 , y10271 , y10272 , y10273 , y10274 , y10275 , y10276 , y10277 , y10278 , y10279 , y10280 , y10281 , y10282 , y10283 , y10284 , y10285 , y10286 , y10287 , y10288 , y10289 , y10290 , y10291 , y10292 , y10293 , y10294 , y10295 , y10296 , y10297 , y10298 , y10299 , y10300 , y10301 , y10302 , y10303 , y10304 , y10305 , y10306 , y10307 , y10308 , y10309 , y10310 , y10311 , y10312 , y10313 , y10314 , y10315 , y10316 , y10317 , y10318 , y10319 , y10320 , y10321 , y10322 , y10323 , y10324 , y10325 , y10326 , y10327 , y10328 , y10329 , y10330 , y10331 , y10332 , y10333 , y10334 , y10335 , y10336 , y10337 , y10338 , y10339 , y10340 , y10341 , y10342 , y10343 , y10344 , y10345 , y10346 , y10347 , y10348 , y10349 , y10350 , y10351 , y10352 , y10353 , y10354 , y10355 , y10356 , y10357 , y10358 , y10359 , y10360 , y10361 , y10362 , y10363 , y10364 , y10365 , y10366 , y10367 , y10368 , y10369 , y10370 , y10371 , y10372 , y10373 , y10374 , y10375 , y10376 , y10377 , y10378 , y10379 , y10380 , y10381 , y10382 , y10383 , y10384 , y10385 , y10386 , y10387 , y10388 , y10389 , y10390 , y10391 , y10392 , y10393 , y10394 , y10395 , y10396 , y10397 , y10398 , y10399 , y10400 , y10401 , y10402 , y10403 , y10404 , y10405 , y10406 , y10407 , y10408 , y10409 , y10410 , y10411 , y10412 , y10413 , y10414 , y10415 , y10416 , y10417 , y10418 , y10419 , y10420 , y10421 , y10422 , y10423 , y10424 , y10425 , y10426 , y10427 , y10428 , y10429 , y10430 , y10431 , y10432 , y10433 , y10434 , y10435 , y10436 , y10437 , y10438 , y10439 , y10440 , y10441 , y10442 , y10443 , y10444 , y10445 , y10446 , y10447 , y10448 , y10449 , y10450 , y10451 , y10452 , y10453 , y10454 , y10455 , y10456 , y10457 , y10458 , y10459 , y10460 , y10461 , y10462 , y10463 , y10464 , y10465 , y10466 , y10467 , y10468 , y10469 , y10470 , y10471 , y10472 , y10473 , y10474 , y10475 , y10476 , y10477 , y10478 , y10479 , y10480 , y10481 , y10482 , y10483 , y10484 , y10485 , y10486 , y10487 , y10488 , y10489 , y10490 , y10491 , y10492 , y10493 , y10494 , y10495 , y10496 , y10497 , y10498 , y10499 , y10500 , y10501 , y10502 , y10503 , y10504 , y10505 , y10506 , y10507 , y10508 , y10509 , y10510 , y10511 , y10512 , y10513 , y10514 , y10515 , y10516 , y10517 , y10518 , y10519 , y10520 , y10521 , y10522 , y10523 , y10524 , y10525 , y10526 , y10527 , y10528 , y10529 , y10530 , y10531 , y10532 , y10533 , y10534 , y10535 , y10536 , y10537 , y10538 , y10539 , y10540 , y10541 , y10542 , y10543 , y10544 , y10545 , y10546 , y10547 , y10548 , y10549 , y10550 , y10551 , y10552 , y10553 , y10554 , y10555 , y10556 , y10557 , y10558 , y10559 , y10560 , y10561 , y10562 , y10563 , y10564 , y10565 , y10566 , y10567 , y10568 , y10569 , y10570 , y10571 , y10572 , y10573 , y10574 , y10575 , y10576 , y10577 , y10578 , y10579 , y10580 , y10581 , y10582 , y10583 , y10584 , y10585 , y10586 , y10587 , y10588 , y10589 , y10590 , y10591 , y10592 , y10593 , y10594 , y10595 , y10596 , y10597 , y10598 , y10599 , y10600 , y10601 , y10602 , y10603 , y10604 , y10605 , y10606 , y10607 , y10608 , y10609 , y10610 , y10611 , y10612 , y10613 , y10614 , y10615 , y10616 , y10617 , y10618 , y10619 , y10620 , y10621 , y10622 , y10623 , y10624 , y10625 , y10626 , y10627 , y10628 , y10629 , y10630 , y10631 , y10632 , y10633 , y10634 , y10635 , y10636 , y10637 , y10638 , y10639 , y10640 , y10641 , y10642 , y10643 , y10644 , y10645 , y10646 , y10647 , y10648 , y10649 , y10650 , y10651 , y10652 , y10653 , y10654 , y10655 , y10656 , y10657 , y10658 , y10659 , y10660 , y10661 , y10662 , y10663 , y10664 , y10665 , y10666 , y10667 , y10668 , y10669 , y10670 , y10671 , y10672 , y10673 , y10674 , y10675 , y10676 , y10677 , y10678 , y10679 , y10680 , y10681 , y10682 , y10683 , y10684 , y10685 , y10686 , y10687 , y10688 , y10689 , y10690 , y10691 , y10692 , y10693 , y10694 , y10695 , y10696 , y10697 , y10698 , y10699 , y10700 , y10701 , y10702 , y10703 , y10704 , y10705 , y10706 , y10707 , y10708 , y10709 , y10710 , y10711 , y10712 , y10713 , y10714 , y10715 , y10716 , y10717 , y10718 , y10719 , y10720 , y10721 , y10722 , y10723 , y10724 , y10725 , y10726 , y10727 , y10728 , y10729 , y10730 , y10731 , y10732 , y10733 , y10734 , y10735 , y10736 , y10737 , y10738 , y10739 , y10740 , y10741 , y10742 , y10743 , y10744 , y10745 , y10746 , y10747 , y10748 , y10749 , y10750 , y10751 , y10752 , y10753 , y10754 , y10755 , y10756 , y10757 , y10758 , y10759 , y10760 , y10761 , y10762 , y10763 , y10764 , y10765 , y10766 , y10767 , y10768 , y10769 , y10770 , y10771 , y10772 , y10773 , y10774 , y10775 , y10776 , y10777 , y10778 , y10779 , y10780 , y10781 , y10782 , y10783 , y10784 , y10785 , y10786 , y10787 , y10788 , y10789 , y10790 , y10791 , y10792 , y10793 , y10794 , y10795 , y10796 , y10797 , y10798 , y10799 , y10800 , y10801 , y10802 , y10803 , y10804 , y10805 , y10806 , y10807 , y10808 , y10809 , y10810 , y10811 , y10812 , y10813 , y10814 , y10815 , y10816 , y10817 , y10818 , y10819 , y10820 , y10821 , y10822 , y10823 , y10824 , y10825 , y10826 , y10827 , y10828 , y10829 , y10830 , y10831 , y10832 , y10833 , y10834 , y10835 , y10836 , y10837 , y10838 , y10839 , y10840 , y10841 , y10842 , y10843 , y10844 , y10845 , y10846 , y10847 , y10848 , y10849 , y10850 , y10851 , y10852 , y10853 , y10854 , y10855 , y10856 , y10857 , y10858 , y10859 , y10860 , y10861 , y10862 , y10863 , y10864 , y10865 , y10866 , y10867 , y10868 , y10869 , y10870 , y10871 , y10872 , y10873 , y10874 , y10875 , y10876 , y10877 , y10878 , y10879 , y10880 , y10881 , y10882 , y10883 , y10884 , y10885 , y10886 , y10887 , y10888 , y10889 , y10890 , y10891 , y10892 , y10893 , y10894 , y10895 , y10896 , y10897 , y10898 , y10899 , y10900 , y10901 , y10902 , y10903 , y10904 , y10905 , y10906 , y10907 , y10908 , y10909 , y10910 , y10911 , y10912 , y10913 , y10914 , y10915 , y10916 , y10917 , y10918 , y10919 , y10920 , y10921 , y10922 , y10923 , y10924 , y10925 , y10926 , y10927 , y10928 , y10929 , y10930 , y10931 , y10932 , y10933 , y10934 , y10935 , y10936 , y10937 , y10938 , y10939 , y10940 , y10941 , y10942 , y10943 , y10944 , y10945 , y10946 , y10947 , y10948 , y10949 , y10950 , y10951 , y10952 , y10953 , y10954 , y10955 , y10956 , y10957 , y10958 , y10959 , y10960 , y10961 , y10962 , y10963 , y10964 , y10965 , y10966 , y10967 , y10968 , y10969 , y10970 , y10971 , y10972 , y10973 , y10974 , y10975 , y10976 , y10977 , y10978 , y10979 , y10980 ;
  wire n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , n18511 , n18512 , n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , n18679 , n18680 , n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , n18709 , n18710 , n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , n18841 , n18842 , n18843 , n18844 , n18845 , n18846 , n18847 , n18848 , n18849 , n18850 , n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , n18870 , n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , n18891 , n18892 , n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , n18910 , n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , n18921 , n18922 , n18923 , n18924 , n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , n18969 , n18970 , n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , n18977 , n18978 , n18979 , n18980 , n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , n18989 , n18990 , n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , n18999 , n19000 , n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , n19017 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , n19029 , n19030 , n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , n19037 , n19038 , n19039 , n19040 , n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , n19049 , n19050 , n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , n19060 , n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , n19067 , n19068 , n19069 , n19070 , n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , n19079 , n19080 , n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , n19089 , n19090 , n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , n19099 , n19100 , n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , n19137 , n19138 , n19139 , n19140 , n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , n19157 , n19158 , n19159 , n19160 , n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , n19167 , n19168 , n19169 , n19170 , n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , n19179 , n19180 , n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , n19189 , n19190 , n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , n19198 , n19199 , n19200 , n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , n19210 , n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , n19217 , n19218 , n19219 , n19220 , n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , n19229 , n19230 , n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , n19239 , n19240 , n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , n19249 , n19250 , n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , n19259 , n19260 , n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , n19279 , n19280 , n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , n19287 , n19288 , n19289 , n19290 , n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , n19297 , n19298 , n19299 , n19300 , n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , n19309 , n19310 , n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , n19319 , n19320 , n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , n19329 , n19330 , n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , n19339 , n19340 , n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , n19359 , n19360 , n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , n19369 , n19370 , n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , n19379 , n19380 , n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19387 , n19388 , n19389 , n19390 , n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , n19400 , n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , n19410 , n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , n19417 , n19418 , n19419 , n19420 , n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , n19440 , n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , n19450 , n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , n19459 , n19460 , n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , n19470 , n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , n19529 , n19530 , n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , n19550 , n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , n19567 , n19568 , n19569 , n19570 , n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , n19587 , n19588 , n19589 , n19590 , n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , n19619 , n19620 , n19621 , n19622 , n19623 , n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , n19670 , n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , n19711 , n19712 , n19713 , n19714 , n19715 , n19716 , n19717 , n19718 , n19719 , n19720 , n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , n19737 , n19738 , n19739 , n19740 , n19741 , n19742 , n19743 , n19744 , n19745 , n19746 , n19747 , n19748 , n19749 , n19750 , n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , n19757 , n19758 , n19759 , n19760 , n19761 , n19762 , n19763 , n19764 , n19765 , n19766 , n19767 , n19768 , n19769 , n19770 , n19771 , n19772 , n19773 , n19774 , n19775 , n19776 , n19777 , n19778 , n19779 , n19780 , n19781 , n19782 , n19783 , n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , n19791 , n19792 , n19793 , n19794 , n19795 , n19796 , n19797 , n19798 , n19799 , n19800 , n19801 , n19802 , n19803 , n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , n19811 , n19812 , n19813 , n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , n19821 , n19822 , n19823 , n19824 , n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , n19831 , n19832 , n19833 , n19834 , n19835 , n19836 , n19837 , n19838 , n19839 , n19840 , n19841 , n19842 , n19843 , n19844 , n19845 , n19846 , n19847 , n19848 , n19849 , n19850 , n19851 , n19852 , n19853 , n19854 , n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , n19861 , n19862 , n19863 , n19864 , n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , n19871 , n19872 , n19873 , n19874 , n19875 , n19876 , n19877 , n19878 , n19879 , n19880 , n19881 , n19882 , n19883 , n19884 , n19885 , n19886 , n19887 , n19888 , n19889 , n19890 , n19891 , n19892 , n19893 , n19894 , n19895 , n19896 , n19897 , n19898 , n19899 , n19900 , n19901 , n19902 , n19903 , n19904 , n19905 , n19906 , n19907 , n19908 , n19909 , n19910 , n19911 , n19912 , n19913 , n19914 , n19915 , n19916 , n19917 , n19918 , n19919 , n19920 , n19921 , n19922 , n19923 , n19924 , n19925 , n19926 , n19927 , n19928 , n19929 , n19930 , n19931 , n19932 , n19933 , n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , n19940 , n19941 , n19942 , n19943 , n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , n19951 , n19952 , n19953 , n19954 , n19955 , n19956 , n19957 , n19958 , n19959 , n19960 , n19961 , n19962 , n19963 , n19964 , n19965 , n19966 , n19967 , n19968 , n19969 , n19970 , n19971 , n19972 , n19973 , n19974 , n19975 , n19976 , n19977 , n19978 , n19979 , n19980 , n19981 , n19982 , n19983 , n19984 , n19985 , n19986 , n19987 , n19988 , n19989 , n19990 , n19991 , n19992 , n19993 , n19994 , n19995 , n19996 , n19997 , n19998 , n19999 , n20000 , n20001 , n20002 , n20003 , n20004 , n20005 , n20006 , n20007 , n20008 , n20009 , n20010 , n20011 , n20012 , n20013 , n20014 , n20015 , n20016 , n20017 , n20018 , n20019 , n20020 , n20021 , n20022 , n20023 , n20024 , n20025 , n20026 , n20027 , n20028 , n20029 , n20030 , n20031 , n20032 , n20033 , n20034 , n20035 , n20036 , n20037 , n20038 , n20039 , n20040 , n20041 , n20042 , n20043 , n20044 , n20045 , n20046 , n20047 , n20048 , n20049 , n20050 , n20051 , n20052 , n20053 , n20054 , n20055 , n20056 , n20057 , n20058 , n20059 , n20060 , n20061 , n20062 , n20063 , n20064 , n20065 , n20066 , n20067 , n20068 , n20069 , n20070 , n20071 , n20072 , n20073 , n20074 , n20075 , n20076 , n20077 , n20078 , n20079 , n20080 , n20081 , n20082 , n20083 , n20084 , n20085 , n20086 , n20087 , n20088 , n20089 , n20090 , n20091 , n20092 , n20093 , n20094 , n20095 , n20096 , n20097 , n20098 , n20099 , n20100 , n20101 , n20102 , n20103 , n20104 , n20105 , n20106 , n20107 , n20108 , n20109 , n20110 , n20111 , n20112 , n20113 , n20114 , n20115 , n20116 , n20117 , n20118 , n20119 , n20120 , n20121 , n20122 , n20123 , n20124 , n20125 , n20126 , n20127 , n20128 , n20129 , n20130 , n20131 , n20132 , n20133 , n20134 , n20135 , n20136 , n20137 , n20138 , n20139 , n20140 , n20141 , n20142 , n20143 , n20144 , n20145 , n20146 , n20147 , n20148 , n20149 , n20150 , n20151 , n20152 , n20153 , n20154 , n20155 , n20156 , n20157 , n20158 , n20159 , n20160 , n20161 , n20162 , n20163 , n20164 , n20165 , n20166 , n20167 , n20168 , n20169 , n20170 , n20171 , n20172 , n20173 , n20174 , n20175 , n20176 , n20177 , n20178 , n20179 , n20180 , n20181 , n20182 , n20183 , n20184 , n20185 , n20186 , n20187 , n20188 , n20189 , n20190 , n20191 , n20192 , n20193 , n20194 , n20195 , n20196 , n20197 , n20198 , n20199 , n20200 , n20201 , n20202 , n20203 , n20204 , n20205 , n20206 , n20207 , n20208 , n20209 , n20210 , n20211 , n20212 , n20213 , n20214 , n20215 , n20216 , n20217 , n20218 , n20219 , n20220 , n20221 , n20222 , n20223 , n20224 , n20225 , n20226 , n20227 , n20228 , n20229 , n20230 , n20231 , n20232 , n20233 , n20234 , n20235 , n20236 , n20237 , n20238 , n20239 , n20240 , n20241 , n20242 , n20243 , n20244 , n20245 , n20246 , n20247 , n20248 , n20249 , n20250 , n20251 , n20252 , n20253 , n20254 , n20255 , n20256 , n20257 , n20258 , n20259 , n20260 , n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , n20267 , n20268 , n20269 , n20270 , n20271 , n20272 , n20273 , n20274 , n20275 , n20276 , n20277 , n20278 , n20279 , n20280 , n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , n20287 , n20288 , n20289 , n20290 , n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , n20297 , n20298 , n20299 , n20300 , n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , n20307 , n20308 , n20309 , n20310 , n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , n20317 , n20318 , n20319 , n20320 , n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , n20327 , n20328 , n20329 , n20330 , n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , n20337 , n20338 , n20339 , n20340 , n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , n20347 , n20348 , n20349 , n20350 , n20351 , n20352 , n20353 , n20354 , n20355 , n20356 , n20357 , n20358 , n20359 , n20360 , n20361 , n20362 , n20363 , n20364 , n20365 , n20366 , n20367 , n20368 , n20369 , n20370 , n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , n20377 , n20378 , n20379 , n20380 , n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , n20389 , n20390 , n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , n20397 , n20398 , n20399 , n20400 , n20401 , n20402 , n20403 , n20404 , n20405 , n20406 , n20407 , n20408 , n20409 , n20410 , n20411 , n20412 , n20413 , n20414 , n20415 , n20416 , n20417 , n20418 , n20419 , n20420 , n20421 , n20422 , n20423 , n20424 , n20425 , n20426 , n20427 , n20428 , n20429 , n20430 , n20431 , n20432 , n20433 , n20434 , n20435 , n20436 , n20437 , n20438 , n20439 , n20440 , n20441 , n20442 , n20443 , n20444 , n20445 , n20446 , n20447 , n20448 , n20449 , n20450 , n20451 , n20452 , n20453 , n20454 , n20455 , n20456 , n20457 , n20458 , n20459 , n20460 , n20461 , n20462 , n20463 , n20464 , n20465 , n20466 , n20467 , n20468 , n20469 , n20470 , n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , n20477 , n20478 , n20479 , n20480 , n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , n20487 , n20488 , n20489 , n20490 , n20491 , n20492 , n20493 , n20494 , n20495 , n20496 , n20497 , n20498 , n20499 , n20500 , n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , n20507 , n20508 , n20509 , n20510 , n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , n20519 , n20520 , n20521 , n20522 , n20523 , n20524 , n20525 , n20526 , n20527 , n20528 , n20529 , n20530 , n20531 , n20532 , n20533 , n20534 , n20535 , n20536 , n20537 , n20538 , n20539 , n20540 , n20541 , n20542 , n20543 , n20544 , n20545 , n20546 , n20547 , n20548 , n20549 , n20550 , n20551 , n20552 , n20553 , n20554 , n20555 , n20556 , n20557 , n20558 , n20559 , n20560 , n20561 , n20562 , n20563 , n20564 , n20565 , n20566 , n20567 , n20568 , n20569 , n20570 , n20571 , n20572 , n20573 , n20574 , n20575 , n20576 , n20577 , n20578 , n20579 , n20580 , n20581 , n20582 , n20583 , n20584 , n20585 , n20586 , n20587 , n20588 , n20589 , n20590 , n20591 , n20592 , n20593 , n20594 , n20595 , n20596 , n20597 , n20598 , n20599 , n20600 , n20601 , n20602 , n20603 , n20604 , n20605 , n20606 , n20607 , n20608 , n20609 , n20610 , n20611 , n20612 , n20613 , n20614 , n20615 , n20616 , n20617 , n20618 , n20619 , n20620 , n20621 , n20622 , n20623 , n20624 , n20625 , n20626 , n20627 , n20628 , n20629 , n20630 , n20631 , n20632 , n20633 , n20634 , n20635 , n20636 , n20637 , n20638 , n20639 , n20640 , n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , n20647 , n20648 , n20649 , n20650 , n20651 , n20652 , n20653 , n20654 , n20655 , n20656 , n20657 , n20658 , n20659 , n20660 , n20661 , n20662 , n20663 , n20664 , n20665 , n20666 , n20667 , n20668 , n20669 , n20670 , n20671 , n20672 , n20673 , n20674 , n20675 , n20676 , n20677 , n20678 , n20679 , n20680 , n20681 , n20682 , n20683 , n20684 , n20685 , n20686 , n20687 , n20688 , n20689 , n20690 , n20691 , n20692 , n20693 , n20694 , n20695 , n20696 , n20697 , n20698 , n20699 , n20700 , n20701 , n20702 , n20703 , n20704 , n20705 , n20706 , n20707 , n20708 , n20709 , n20710 , n20711 , n20712 , n20713 , n20714 , n20715 , n20716 , n20717 , n20718 , n20719 , n20720 , n20721 , n20722 , n20723 , n20724 , n20725 , n20726 , n20727 , n20728 , n20729 , n20730 , n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , n20737 , n20738 , n20739 , n20740 , n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , n20747 , n20748 , n20749 , n20750 , n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , n20757 , n20758 , n20759 , n20760 , n20761 , n20762 , n20763 , n20764 , n20765 , n20766 , n20767 , n20768 , n20769 , n20770 , n20771 , n20772 , n20773 , n20774 , n20775 , n20776 , n20777 , n20778 , n20779 , n20780 , n20781 , n20782 , n20783 , n20784 , n20785 , n20786 , n20787 , n20788 , n20789 , n20790 , n20791 , n20792 , n20793 , n20794 , n20795 , n20796 , n20797 , n20798 , n20799 , n20800 , n20801 , n20802 , n20803 , n20804 , n20805 , n20806 , n20807 , n20808 , n20809 , n20810 , n20811 , n20812 , n20813 , n20814 , n20815 , n20816 , n20817 , n20818 , n20819 , n20820 , n20821 , n20822 , n20823 , n20824 , n20825 , n20826 , n20827 , n20828 , n20829 , n20830 , n20831 , n20832 , n20833 , n20834 , n20835 , n20836 , n20837 , n20838 , n20839 , n20840 , n20841 , n20842 , n20843 , n20844 , n20845 , n20846 , n20847 , n20848 , n20849 , n20850 , n20851 , n20852 , n20853 , n20854 , n20855 , n20856 , n20857 , n20858 , n20859 , n20860 , n20861 , n20862 , n20863 , n20864 , n20865 , n20866 , n20867 , n20868 , n20869 , n20870 , n20871 , n20872 , n20873 , n20874 , n20875 , n20876 , n20877 , n20878 , n20879 , n20880 , n20881 , n20882 , n20883 , n20884 , n20885 , n20886 , n20887 , n20888 , n20889 , n20890 , n20891 , n20892 , n20893 , n20894 , n20895 , n20896 , n20897 , n20898 , n20899 , n20900 , n20901 , n20902 , n20903 , n20904 , n20905 , n20906 , n20907 , n20908 , n20909 , n20910 , n20911 , n20912 , n20913 , n20914 , n20915 , n20916 , n20917 , n20918 , n20919 , n20920 , n20921 , n20922 , n20923 , n20924 , n20925 , n20926 , n20927 , n20928 , n20929 , n20930 , n20931 , n20932 , n20933 , n20934 , n20935 , n20936 , n20937 , n20938 , n20939 , n20940 , n20941 , n20942 , n20943 , n20944 , n20945 , n20946 , n20947 , n20948 , n20949 , n20950 , n20951 , n20952 , n20953 , n20954 , n20955 , n20956 , n20957 , n20958 , n20959 , n20960 , n20961 , n20962 , n20963 , n20964 , n20965 , n20966 , n20967 , n20968 , n20969 , n20970 , n20971 , n20972 , n20973 , n20974 , n20975 , n20976 , n20977 , n20978 , n20979 , n20980 , n20981 , n20982 , n20983 , n20984 , n20985 , n20986 , n20987 , n20988 , n20989 , n20990 , n20991 , n20992 , n20993 , n20994 , n20995 , n20996 , n20997 , n20998 , n20999 , n21000 , n21001 , n21002 , n21003 , n21004 , n21005 , n21006 , n21007 , n21008 , n21009 , n21010 , n21011 , n21012 , n21013 , n21014 , n21015 , n21016 , n21017 , n21018 , n21019 , n21020 , n21021 , n21022 , n21023 , n21024 , n21025 , n21026 , n21027 , n21028 , n21029 , n21030 , n21031 , n21032 , n21033 , n21034 , n21035 , n21036 , n21037 , n21038 , n21039 , n21040 , n21041 , n21042 , n21043 , n21044 , n21045 , n21046 , n21047 , n21048 , n21049 , n21050 , n21051 , n21052 , n21053 , n21054 , n21055 , n21056 , n21057 , n21058 , n21059 , n21060 , n21061 , n21062 , n21063 , n21064 , n21065 , n21066 , n21067 , n21068 , n21069 , n21070 , n21071 , n21072 , n21073 , n21074 , n21075 , n21076 , n21077 , n21078 , n21079 , n21080 , n21081 , n21082 , n21083 , n21084 , n21085 , n21086 , n21087 , n21088 , n21089 , n21090 , n21091 , n21092 , n21093 , n21094 , n21095 , n21096 , n21097 , n21098 , n21099 , n21100 , n21101 , n21102 , n21103 , n21104 , n21105 , n21106 , n21107 , n21108 , n21109 , n21110 , n21111 , n21112 , n21113 , n21114 , n21115 , n21116 , n21117 , n21118 , n21119 , n21120 , n21121 , n21122 , n21123 , n21124 , n21125 , n21126 , n21127 , n21128 , n21129 , n21130 , n21131 , n21132 , n21133 , n21134 , n21135 , n21136 , n21137 , n21138 , n21139 , n21140 , n21141 , n21142 , n21143 , n21144 , n21145 , n21146 , n21147 , n21148 , n21149 , n21150 , n21151 , n21152 , n21153 , n21154 , n21155 , n21156 , n21157 , n21158 , n21159 , n21160 , n21161 , n21162 , n21163 , n21164 , n21165 , n21166 , n21167 , n21168 , n21169 , n21170 , n21171 , n21172 , n21173 , n21174 , n21175 , n21176 , n21177 , n21178 , n21179 , n21180 , n21181 , n21182 , n21183 , n21184 , n21185 , n21186 , n21187 , n21188 , n21189 , n21190 , n21191 , n21192 , n21193 , n21194 , n21195 , n21196 , n21197 , n21198 , n21199 , n21200 , n21201 , n21202 , n21203 , n21204 , n21205 , n21206 , n21207 , n21208 , n21209 , n21210 , n21211 , n21212 , n21213 , n21214 , n21215 , n21216 , n21217 , n21218 , n21219 , n21220 , n21221 , n21222 , n21223 , n21224 , n21225 , n21226 , n21227 , n21228 , n21229 , n21230 , n21231 , n21232 , n21233 , n21234 , n21235 , n21236 , n21237 , n21238 , n21239 , n21240 , n21241 , n21242 , n21243 , n21244 , n21245 , n21246 , n21247 , n21248 , n21249 , n21250 , n21251 , n21252 , n21253 , n21254 , n21255 , n21256 , n21257 , n21258 , n21259 , n21260 , n21261 , n21262 , n21263 , n21264 , n21265 , n21266 , n21267 , n21268 , n21269 , n21270 , n21271 , n21272 , n21273 , n21274 , n21275 , n21276 , n21277 , n21278 , n21279 , n21280 , n21281 , n21282 , n21283 , n21284 , n21285 , n21286 , n21287 , n21288 , n21289 , n21290 , n21291 , n21292 , n21293 , n21294 , n21295 , n21296 , n21297 , n21298 , n21299 , n21300 , n21301 , n21302 , n21303 , n21304 , n21305 , n21306 , n21307 , n21308 , n21309 , n21310 , n21311 , n21312 , n21313 , n21314 , n21315 , n21316 , n21317 , n21318 , n21319 , n21320 , n21321 , n21322 , n21323 , n21324 , n21325 , n21326 , n21327 , n21328 , n21329 , n21330 , n21331 , n21332 , n21333 , n21334 , n21335 , n21336 , n21337 , n21338 , n21339 , n21340 , n21341 , n21342 , n21343 , n21344 , n21345 , n21346 , n21347 , n21348 , n21349 , n21350 , n21351 , n21352 , n21353 , n21354 , n21355 , n21356 , n21357 , n21358 , n21359 , n21360 , n21361 , n21362 , n21363 , n21364 , n21365 , n21366 , n21367 , n21368 , n21369 , n21370 , n21371 , n21372 , n21373 , n21374 , n21375 , n21376 , n21377 , n21378 , n21379 , n21380 , n21381 , n21382 , n21383 , n21384 , n21385 , n21386 , n21387 , n21388 , n21389 , n21390 , n21391 , n21392 , n21393 , n21394 , n21395 , n21396 , n21397 , n21398 , n21399 , n21400 , n21401 , n21402 , n21403 , n21404 , n21405 , n21406 , n21407 , n21408 , n21409 , n21410 , n21411 , n21412 , n21413 , n21414 , n21415 , n21416 , n21417 , n21418 , n21419 , n21420 , n21421 , n21422 , n21423 , n21424 , n21425 , n21426 , n21427 , n21428 , n21429 , n21430 , n21431 , n21432 , n21433 , n21434 , n21435 , n21436 , n21437 , n21438 , n21439 , n21440 , n21441 , n21442 , n21443 , n21444 , n21445 , n21446 , n21447 , n21448 , n21449 , n21450 , n21451 , n21452 , n21453 , n21454 , n21455 , n21456 , n21457 , n21458 , n21459 , n21460 , n21461 , n21462 , n21463 , n21464 , n21465 , n21466 , n21467 , n21468 , n21469 , n21470 , n21471 , n21472 , n21473 , n21474 , n21475 , n21476 , n21477 , n21478 , n21479 , n21480 , n21481 , n21482 , n21483 , n21484 , n21485 , n21486 , n21487 , n21488 , n21489 , n21490 , n21491 , n21492 , n21493 , n21494 , n21495 , n21496 , n21497 , n21498 , n21499 , n21500 , n21501 , n21502 , n21503 , n21504 , n21505 , n21506 , n21507 , n21508 , n21509 , n21510 , n21511 , n21512 , n21513 , n21514 , n21515 , n21516 , n21517 , n21518 , n21519 , n21520 , n21521 , n21522 , n21523 , n21524 , n21525 , n21526 , n21527 , n21528 , n21529 , n21530 , n21531 , n21532 , n21533 , n21534 , n21535 , n21536 , n21537 , n21538 , n21539 , n21540 , n21541 , n21542 , n21543 , n21544 , n21545 , n21546 , n21547 , n21548 , n21549 , n21550 , n21551 , n21552 , n21553 , n21554 , n21555 , n21556 , n21557 , n21558 , n21559 , n21560 , n21561 , n21562 , n21563 , n21564 , n21565 , n21566 , n21567 , n21568 , n21569 , n21570 , n21571 , n21572 , n21573 , n21574 , n21575 , n21576 , n21577 , n21578 , n21579 , n21580 , n21581 , n21582 , n21583 , n21584 , n21585 , n21586 , n21587 , n21588 , n21589 , n21590 , n21591 , n21592 , n21593 , n21594 , n21595 , n21596 , n21597 , n21598 , n21599 , n21600 , n21601 , n21602 , n21603 , n21604 , n21605 , n21606 , n21607 , n21608 , n21609 , n21610 , n21611 , n21612 , n21613 , n21614 , n21615 , n21616 , n21617 , n21618 , n21619 , n21620 , n21621 , n21622 , n21623 , n21624 , n21625 , n21626 , n21627 , n21628 , n21629 , n21630 , n21631 , n21632 , n21633 , n21634 , n21635 , n21636 , n21637 , n21638 , n21639 , n21640 , n21641 , n21642 , n21643 , n21644 , n21645 , n21646 , n21647 , n21648 , n21649 , n21650 , n21651 , n21652 , n21653 , n21654 , n21655 , n21656 , n21657 , n21658 , n21659 , n21660 , n21661 , n21662 , n21663 , n21664 , n21665 , n21666 , n21667 , n21668 , n21669 , n21670 , n21671 , n21672 , n21673 , n21674 , n21675 , n21676 , n21677 , n21678 , n21679 , n21680 , n21681 , n21682 , n21683 , n21684 , n21685 , n21686 , n21687 , n21688 , n21689 , n21690 , n21691 , n21692 , n21693 , n21694 , n21695 , n21696 , n21697 , n21698 , n21699 , n21700 , n21701 , n21702 , n21703 , n21704 , n21705 , n21706 , n21707 , n21708 , n21709 , n21710 , n21711 , n21712 , n21713 , n21714 , n21715 , n21716 , n21717 , n21718 , n21719 , n21720 , n21721 , n21722 , n21723 , n21724 , n21725 , n21726 , n21727 , n21728 , n21729 , n21730 , n21731 , n21732 , n21733 , n21734 , n21735 , n21736 , n21737 , n21738 , n21739 , n21740 , n21741 , n21742 , n21743 , n21744 , n21745 , n21746 , n21747 , n21748 , n21749 , n21750 , n21751 , n21752 , n21753 , n21754 , n21755 , n21756 , n21757 , n21758 , n21759 , n21760 , n21761 , n21762 , n21763 , n21764 , n21765 , n21766 , n21767 , n21768 , n21769 , n21770 , n21771 , n21772 , n21773 , n21774 , n21775 , n21776 , n21777 , n21778 , n21779 , n21780 , n21781 , n21782 , n21783 , n21784 , n21785 , n21786 , n21787 , n21788 , n21789 , n21790 , n21791 , n21792 , n21793 , n21794 , n21795 , n21796 , n21797 , n21798 , n21799 , n21800 , n21801 , n21802 , n21803 , n21804 , n21805 , n21806 , n21807 , n21808 , n21809 , n21810 , n21811 , n21812 , n21813 , n21814 , n21815 , n21816 , n21817 , n21818 , n21819 , n21820 , n21821 , n21822 , n21823 , n21824 , n21825 , n21826 , n21827 , n21828 , n21829 , n21830 , n21831 , n21832 , n21833 , n21834 , n21835 , n21836 , n21837 , n21838 , n21839 , n21840 , n21841 , n21842 , n21843 , n21844 , n21845 , n21846 , n21847 , n21848 , n21849 , n21850 , n21851 , n21852 , n21853 , n21854 , n21855 , n21856 , n21857 , n21858 , n21859 , n21860 , n21861 , n21862 , n21863 , n21864 , n21865 , n21866 , n21867 , n21868 , n21869 , n21870 , n21871 , n21872 , n21873 , n21874 , n21875 , n21876 , n21877 , n21878 , n21879 , n21880 , n21881 , n21882 , n21883 , n21884 , n21885 , n21886 , n21887 , n21888 , n21889 , n21890 , n21891 , n21892 , n21893 , n21894 , n21895 , n21896 , n21897 , n21898 , n21899 , n21900 , n21901 , n21902 , n21903 , n21904 , n21905 , n21906 , n21907 , n21908 , n21909 , n21910 , n21911 , n21912 , n21913 , n21914 , n21915 , n21916 , n21917 , n21918 , n21919 , n21920 , n21921 , n21922 , n21923 , n21924 , n21925 , n21926 , n21927 , n21928 , n21929 , n21930 , n21931 , n21932 , n21933 , n21934 , n21935 , n21936 , n21937 , n21938 , n21939 , n21940 , n21941 , n21942 , n21943 , n21944 , n21945 , n21946 , n21947 , n21948 , n21949 , n21950 , n21951 , n21952 , n21953 , n21954 , n21955 , n21956 , n21957 , n21958 , n21959 , n21960 , n21961 , n21962 , n21963 , n21964 , n21965 , n21966 , n21967 , n21968 , n21969 , n21970 , n21971 , n21972 , n21973 , n21974 , n21975 , n21976 , n21977 , n21978 , n21979 , n21980 , n21981 , n21982 , n21983 , n21984 , n21985 , n21986 , n21987 , n21988 , n21989 , n21990 , n21991 , n21992 , n21993 , n21994 , n21995 , n21996 , n21997 , n21998 , n21999 , n22000 , n22001 , n22002 , n22003 , n22004 , n22005 , n22006 , n22007 , n22008 , n22009 , n22010 , n22011 , n22012 , n22013 , n22014 , n22015 , n22016 , n22017 , n22018 , n22019 , n22020 , n22021 , n22022 , n22023 , n22024 , n22025 , n22026 , n22027 , n22028 , n22029 , n22030 , n22031 , n22032 , n22033 , n22034 , n22035 , n22036 , n22037 , n22038 , n22039 , n22040 , n22041 , n22042 , n22043 , n22044 , n22045 , n22046 , n22047 , n22048 , n22049 , n22050 , n22051 , n22052 , n22053 , n22054 , n22055 , n22056 , n22057 , n22058 , n22059 , n22060 , n22061 , n22062 , n22063 , n22064 , n22065 , n22066 , n22067 , n22068 , n22069 , n22070 , n22071 , n22072 , n22073 , n22074 , n22075 , n22076 , n22077 , n22078 , n22079 , n22080 , n22081 , n22082 , n22083 , n22084 , n22085 , n22086 , n22087 , n22088 , n22089 , n22090 , n22091 , n22092 , n22093 , n22094 , n22095 , n22096 , n22097 , n22098 , n22099 , n22100 , n22101 , n22102 , n22103 , n22104 , n22105 , n22106 , n22107 , n22108 , n22109 , n22110 , n22111 , n22112 , n22113 , n22114 , n22115 , n22116 , n22117 , n22118 , n22119 , n22120 , n22121 , n22122 , n22123 , n22124 , n22125 , n22126 , n22127 , n22128 , n22129 , n22130 , n22131 , n22132 , n22133 , n22134 , n22135 , n22136 , n22137 , n22138 , n22139 , n22140 , n22141 , n22142 , n22143 , n22144 , n22145 , n22146 , n22147 , n22148 , n22149 , n22150 , n22151 , n22152 , n22153 , n22154 , n22155 , n22156 , n22157 , n22158 , n22159 , n22160 , n22161 , n22162 , n22163 , n22164 , n22165 , n22166 , n22167 , n22168 , n22169 , n22170 , n22171 , n22172 , n22173 , n22174 , n22175 , n22176 , n22177 , n22178 , n22179 , n22180 , n22181 , n22182 , n22183 , n22184 , n22185 , n22186 , n22187 , n22188 , n22189 , n22190 , n22191 , n22192 , n22193 , n22194 , n22195 , n22196 , n22197 , n22198 , n22199 , n22200 , n22201 , n22202 , n22203 , n22204 , n22205 , n22206 , n22207 , n22208 , n22209 , n22210 , n22211 , n22212 , n22213 , n22214 , n22215 , n22216 , n22217 , n22218 , n22219 , n22220 , n22221 , n22222 , n22223 , n22224 , n22225 , n22226 , n22227 , n22228 , n22229 , n22230 , n22231 , n22232 , n22233 , n22234 , n22235 , n22236 , n22237 , n22238 , n22239 , n22240 , n22241 , n22242 , n22243 , n22244 , n22245 , n22246 , n22247 , n22248 , n22249 , n22250 , n22251 , n22252 , n22253 , n22254 , n22255 , n22256 , n22257 , n22258 , n22259 , n22260 , n22261 , n22262 , n22263 , n22264 , n22265 , n22266 , n22267 , n22268 , n22269 , n22270 , n22271 , n22272 , n22273 , n22274 , n22275 , n22276 , n22277 , n22278 , n22279 , n22280 , n22281 , n22282 , n22283 , n22284 , n22285 , n22286 , n22287 , n22288 , n22289 , n22290 , n22291 , n22292 , n22293 , n22294 , n22295 , n22296 , n22297 , n22298 , n22299 , n22300 , n22301 , n22302 , n22303 , n22304 , n22305 , n22306 , n22307 , n22308 , n22309 , n22310 , n22311 , n22312 , n22313 , n22314 , n22315 , n22316 , n22317 , n22318 , n22319 , n22320 , n22321 , n22322 , n22323 , n22324 , n22325 , n22326 , n22327 , n22328 , n22329 , n22330 , n22331 , n22332 , n22333 , n22334 , n22335 , n22336 , n22337 , n22338 , n22339 , n22340 , n22341 , n22342 , n22343 , n22344 , n22345 , n22346 , n22347 , n22348 , n22349 , n22350 , n22351 , n22352 , n22353 , n22354 , n22355 , n22356 , n22357 , n22358 , n22359 , n22360 , n22361 , n22362 , n22363 , n22364 , n22365 , n22366 , n22367 , n22368 , n22369 , n22370 , n22371 , n22372 , n22373 , n22374 , n22375 , n22376 , n22377 , n22378 , n22379 , n22380 , n22381 , n22382 , n22383 , n22384 , n22385 , n22386 , n22387 , n22388 , n22389 , n22390 , n22391 , n22392 , n22393 , n22394 , n22395 , n22396 , n22397 , n22398 , n22399 , n22400 , n22401 , n22402 , n22403 , n22404 , n22405 , n22406 , n22407 , n22408 , n22409 , n22410 , n22411 , n22412 , n22413 , n22414 , n22415 , n22416 , n22417 , n22418 , n22419 , n22420 , n22421 , n22422 , n22423 , n22424 , n22425 , n22426 , n22427 , n22428 , n22429 , n22430 , n22431 , n22432 , n22433 , n22434 , n22435 , n22436 , n22437 , n22438 , n22439 , n22440 , n22441 , n22442 , n22443 , n22444 , n22445 , n22446 , n22447 , n22448 , n22449 , n22450 , n22451 , n22452 , n22453 , n22454 , n22455 , n22456 , n22457 , n22458 , n22459 , n22460 , n22461 , n22462 , n22463 , n22464 , n22465 , n22466 , n22467 , n22468 , n22469 , n22470 , n22471 , n22472 , n22473 , n22474 , n22475 , n22476 , n22477 , n22478 , n22479 , n22480 , n22481 , n22482 , n22483 , n22484 , n22485 , n22486 , n22487 , n22488 , n22489 , n22490 , n22491 , n22492 , n22493 , n22494 , n22495 , n22496 , n22497 , n22498 , n22499 , n22500 , n22501 , n22502 , n22503 , n22504 , n22505 , n22506 , n22507 , n22508 , n22509 , n22510 , n22511 , n22512 , n22513 , n22514 , n22515 , n22516 , n22517 , n22518 , n22519 , n22520 , n22521 , n22522 , n22523 , n22524 , n22525 , n22526 , n22527 , n22528 , n22529 , n22530 , n22531 , n22532 , n22533 , n22534 , n22535 , n22536 , n22537 , n22538 , n22539 , n22540 , n22541 , n22542 , n22543 , n22544 , n22545 , n22546 , n22547 , n22548 , n22549 , n22550 , n22551 , n22552 , n22553 , n22554 , n22555 , n22556 , n22557 , n22558 , n22559 , n22560 , n22561 , n22562 , n22563 , n22564 , n22565 , n22566 , n22567 , n22568 , n22569 , n22570 , n22571 , n22572 , n22573 , n22574 , n22575 , n22576 , n22577 , n22578 , n22579 , n22580 , n22581 , n22582 , n22583 , n22584 , n22585 , n22586 , n22587 , n22588 , n22589 , n22590 , n22591 , n22592 , n22593 , n22594 , n22595 , n22596 , n22597 , n22598 , n22599 , n22600 , n22601 , n22602 , n22603 , n22604 , n22605 , n22606 , n22607 , n22608 , n22609 , n22610 , n22611 , n22612 , n22613 , n22614 , n22615 , n22616 , n22617 , n22618 , n22619 , n22620 , n22621 , n22622 , n22623 , n22624 , n22625 , n22626 , n22627 , n22628 , n22629 , n22630 , n22631 , n22632 , n22633 , n22634 , n22635 , n22636 , n22637 , n22638 , n22639 , n22640 , n22641 , n22642 , n22643 , n22644 , n22645 , n22646 , n22647 , n22648 , n22649 , n22650 , n22651 , n22652 , n22653 , n22654 , n22655 , n22656 , n22657 , n22658 , n22659 , n22660 , n22661 , n22662 , n22663 , n22664 , n22665 , n22666 , n22667 , n22668 , n22669 , n22670 , n22671 , n22672 , n22673 , n22674 , n22675 , n22676 , n22677 , n22678 , n22679 , n22680 , n22681 , n22682 , n22683 , n22684 , n22685 , n22686 , n22687 , n22688 , n22689 , n22690 , n22691 , n22692 , n22693 , n22694 , n22695 , n22696 , n22697 , n22698 , n22699 , n22700 , n22701 , n22702 , n22703 , n22704 , n22705 , n22706 , n22707 , n22708 , n22709 , n22710 , n22711 , n22712 , n22713 , n22714 , n22715 , n22716 , n22717 , n22718 , n22719 , n22720 , n22721 , n22722 , n22723 , n22724 , n22725 , n22726 , n22727 , n22728 , n22729 , n22730 , n22731 , n22732 , n22733 , n22734 , n22735 , n22736 , n22737 , n22738 , n22739 , n22740 , n22741 , n22742 , n22743 , n22744 , n22745 , n22746 , n22747 , n22748 , n22749 , n22750 , n22751 , n22752 , n22753 , n22754 , n22755 , n22756 , n22757 , n22758 , n22759 , n22760 , n22761 , n22762 , n22763 , n22764 , n22765 , n22766 , n22767 , n22768 , n22769 , n22770 , n22771 , n22772 , n22773 , n22774 , n22775 , n22776 , n22777 , n22778 , n22779 , n22780 , n22781 , n22782 , n22783 , n22784 , n22785 , n22786 , n22787 , n22788 , n22789 , n22790 , n22791 , n22792 , n22793 , n22794 , n22795 , n22796 , n22797 , n22798 , n22799 , n22800 , n22801 , n22802 , n22803 , n22804 , n22805 , n22806 , n22807 , n22808 , n22809 , n22810 , n22811 , n22812 , n22813 , n22814 , n22815 , n22816 , n22817 , n22818 , n22819 , n22820 , n22821 , n22822 , n22823 , n22824 , n22825 , n22826 , n22827 , n22828 , n22829 , n22830 , n22831 , n22832 , n22833 , n22834 , n22835 , n22836 , n22837 , n22838 , n22839 , n22840 , n22841 , n22842 , n22843 , n22844 , n22845 , n22846 , n22847 , n22848 , n22849 , n22850 , n22851 , n22852 , n22853 , n22854 , n22855 , n22856 , n22857 , n22858 , n22859 , n22860 , n22861 , n22862 , n22863 , n22864 , n22865 , n22866 , n22867 , n22868 , n22869 , n22870 , n22871 , n22872 , n22873 , n22874 , n22875 , n22876 , n22877 , n22878 , n22879 , n22880 , n22881 , n22882 , n22883 , n22884 , n22885 , n22886 , n22887 , n22888 , n22889 , n22890 , n22891 , n22892 , n22893 , n22894 , n22895 , n22896 , n22897 , n22898 , n22899 , n22900 , n22901 , n22902 , n22903 , n22904 , n22905 , n22906 , n22907 , n22908 , n22909 , n22910 , n22911 , n22912 , n22913 , n22914 , n22915 , n22916 , n22917 , n22918 , n22919 , n22920 , n22921 , n22922 , n22923 , n22924 , n22925 , n22926 , n22927 , n22928 , n22929 , n22930 , n22931 , n22932 , n22933 , n22934 , n22935 , n22936 , n22937 , n22938 , n22939 , n22940 , n22941 , n22942 , n22943 , n22944 , n22945 , n22946 , n22947 , n22948 , n22949 , n22950 , n22951 , n22952 , n22953 , n22954 , n22955 , n22956 , n22957 , n22958 , n22959 , n22960 , n22961 , n22962 , n22963 , n22964 , n22965 , n22966 , n22967 , n22968 , n22969 , n22970 , n22971 , n22972 , n22973 , n22974 , n22975 , n22976 , n22977 , n22978 , n22979 , n22980 , n22981 , n22982 , n22983 , n22984 , n22985 , n22986 , n22987 , n22988 , n22989 , n22990 , n22991 , n22992 , n22993 , n22994 , n22995 , n22996 , n22997 , n22998 , n22999 , n23000 , n23001 , n23002 , n23003 , n23004 , n23005 , n23006 , n23007 , n23008 , n23009 , n23010 , n23011 , n23012 , n23013 , n23014 , n23015 , n23016 , n23017 , n23018 , n23019 , n23020 , n23021 , n23022 , n23023 , n23024 , n23025 , n23026 , n23027 , n23028 , n23029 , n23030 , n23031 , n23032 , n23033 , n23034 , n23035 , n23036 , n23037 , n23038 , n23039 , n23040 , n23041 , n23042 , n23043 , n23044 , n23045 , n23046 , n23047 , n23048 , n23049 , n23050 , n23051 , n23052 , n23053 , n23054 , n23055 , n23056 , n23057 , n23058 , n23059 , n23060 , n23061 , n23062 , n23063 , n23064 , n23065 , n23066 , n23067 , n23068 , n23069 , n23070 , n23071 , n23072 , n23073 , n23074 , n23075 , n23076 , n23077 , n23078 , n23079 , n23080 , n23081 , n23082 , n23083 , n23084 , n23085 , n23086 , n23087 , n23088 , n23089 , n23090 , n23091 , n23092 , n23093 , n23094 , n23095 , n23096 , n23097 , n23098 , n23099 , n23100 , n23101 , n23102 , n23103 , n23104 , n23105 , n23106 , n23107 , n23108 , n23109 , n23110 , n23111 , n23112 , n23113 , n23114 , n23115 , n23116 , n23117 , n23118 , n23119 , n23120 , n23121 , n23122 , n23123 , n23124 , n23125 , n23126 , n23127 , n23128 , n23129 , n23130 , n23131 , n23132 , n23133 , n23134 , n23135 , n23136 , n23137 , n23138 , n23139 , n23140 , n23141 , n23142 , n23143 , n23144 , n23145 , n23146 , n23147 , n23148 , n23149 , n23150 , n23151 , n23152 , n23153 , n23154 , n23155 , n23156 , n23157 , n23158 , n23159 , n23160 , n23161 , n23162 , n23163 , n23164 , n23165 , n23166 , n23167 , n23168 , n23169 , n23170 , n23171 , n23172 , n23173 , n23174 , n23175 , n23176 , n23177 , n23178 , n23179 , n23180 , n23181 , n23182 , n23183 , n23184 , n23185 , n23186 , n23187 , n23188 , n23189 , n23190 , n23191 , n23192 , n23193 , n23194 , n23195 , n23196 , n23197 , n23198 , n23199 , n23200 , n23201 , n23202 , n23203 , n23204 , n23205 , n23206 , n23207 , n23208 , n23209 , n23210 , n23211 , n23212 , n23213 , n23214 , n23215 , n23216 , n23217 , n23218 , n23219 , n23220 , n23221 , n23222 , n23223 , n23224 , n23225 , n23226 , n23227 , n23228 , n23229 , n23230 , n23231 , n23232 , n23233 , n23234 , n23235 , n23236 , n23237 , n23238 , n23239 , n23240 , n23241 , n23242 , n23243 , n23244 , n23245 , n23246 , n23247 , n23248 , n23249 , n23250 , n23251 , n23252 , n23253 , n23254 , n23255 , n23256 , n23257 , n23258 , n23259 , n23260 , n23261 , n23262 , n23263 , n23264 , n23265 , n23266 , n23267 , n23268 , n23269 , n23270 , n23271 , n23272 , n23273 , n23274 , n23275 , n23276 , n23277 , n23278 , n23279 , n23280 , n23281 , n23282 , n23283 , n23284 , n23285 , n23286 , n23287 , n23288 , n23289 , n23290 , n23291 , n23292 , n23293 , n23294 , n23295 , n23296 , n23297 , n23298 , n23299 , n23300 , n23301 , n23302 , n23303 , n23304 , n23305 , n23306 , n23307 , n23308 , n23309 , n23310 , n23311 , n23312 , n23313 , n23314 , n23315 , n23316 , n23317 , n23318 , n23319 , n23320 , n23321 , n23322 , n23323 , n23324 , n23325 , n23326 , n23327 , n23328 , n23329 , n23330 , n23331 , n23332 , n23333 , n23334 , n23335 , n23336 , n23337 , n23338 , n23339 , n23340 , n23341 , n23342 , n23343 , n23344 , n23345 , n23346 , n23347 , n23348 , n23349 , n23350 , n23351 , n23352 , n23353 , n23354 , n23355 , n23356 , n23357 , n23358 , n23359 , n23360 , n23361 , n23362 , n23363 , n23364 , n23365 , n23366 , n23367 , n23368 , n23369 , n23370 , n23371 , n23372 , n23373 , n23374 , n23375 , n23376 , n23377 , n23378 , n23379 , n23380 , n23381 , n23382 , n23383 , n23384 , n23385 , n23386 , n23387 , n23388 , n23389 , n23390 , n23391 , n23392 , n23393 , n23394 , n23395 , n23396 , n23397 , n23398 , n23399 , n23400 , n23401 , n23402 , n23403 , n23404 , n23405 , n23406 , n23407 , n23408 , n23409 , n23410 , n23411 , n23412 , n23413 , n23414 , n23415 , n23416 , n23417 , n23418 , n23419 , n23420 , n23421 , n23422 , n23423 , n23424 , n23425 , n23426 , n23427 , n23428 , n23429 , n23430 , n23431 , n23432 , n23433 , n23434 , n23435 , n23436 , n23437 , n23438 , n23439 , n23440 , n23441 , n23442 , n23443 , n23444 , n23445 , n23446 , n23447 , n23448 , n23449 , n23450 , n23451 , n23452 , n23453 , n23454 , n23455 , n23456 , n23457 , n23458 , n23459 , n23460 , n23461 , n23462 , n23463 , n23464 , n23465 , n23466 , n23467 , n23468 , n23469 , n23470 , n23471 , n23472 , n23473 , n23474 , n23475 , n23476 , n23477 , n23478 , n23479 , n23480 , n23481 , n23482 , n23483 , n23484 , n23485 , n23486 , n23487 , n23488 , n23489 , n23490 , n23491 , n23492 , n23493 , n23494 , n23495 , n23496 , n23497 , n23498 , n23499 , n23500 , n23501 , n23502 , n23503 , n23504 , n23505 , n23506 , n23507 , n23508 , n23509 , n23510 , n23511 , n23512 , n23513 , n23514 , n23515 , n23516 , n23517 , n23518 , n23519 , n23520 , n23521 , n23522 , n23523 , n23524 , n23525 , n23526 , n23527 , n23528 , n23529 , n23530 , n23531 , n23532 , n23533 , n23534 , n23535 , n23536 , n23537 , n23538 , n23539 , n23540 , n23541 , n23542 , n23543 , n23544 , n23545 , n23546 , n23547 , n23548 , n23549 , n23550 , n23551 , n23552 , n23553 , n23554 , n23555 , n23556 , n23557 , n23558 , n23559 , n23560 , n23561 , n23562 , n23563 , n23564 , n23565 , n23566 , n23567 , n23568 , n23569 , n23570 , n23571 , n23572 , n23573 , n23574 , n23575 , n23576 , n23577 , n23578 , n23579 , n23580 , n23581 , n23582 , n23583 , n23584 , n23585 , n23586 , n23587 , n23588 , n23589 , n23590 , n23591 , n23592 , n23593 , n23594 , n23595 , n23596 , n23597 , n23598 , n23599 , n23600 , n23601 , n23602 , n23603 , n23604 , n23605 , n23606 , n23607 , n23608 , n23609 , n23610 , n23611 , n23612 , n23613 , n23614 , n23615 , n23616 , n23617 , n23618 , n23619 , n23620 , n23621 , n23622 , n23623 , n23624 , n23625 , n23626 , n23627 , n23628 , n23629 , n23630 , n23631 , n23632 , n23633 , n23634 , n23635 , n23636 , n23637 , n23638 , n23639 , n23640 , n23641 , n23642 , n23643 , n23644 , n23645 , n23646 , n23647 , n23648 , n23649 , n23650 , n23651 , n23652 , n23653 , n23654 , n23655 , n23656 , n23657 , n23658 , n23659 , n23660 , n23661 , n23662 , n23663 , n23664 , n23665 , n23666 , n23667 , n23668 , n23669 , n23670 , n23671 , n23672 , n23673 , n23674 , n23675 , n23676 , n23677 , n23678 , n23679 , n23680 , n23681 , n23682 , n23683 , n23684 , n23685 , n23686 , n23687 , n23688 , n23689 , n23690 , n23691 , n23692 , n23693 , n23694 , n23695 , n23696 , n23697 , n23698 , n23699 , n23700 , n23701 , n23702 , n23703 , n23704 , n23705 , n23706 , n23707 , n23708 , n23709 , n23710 , n23711 , n23712 , n23713 , n23714 , n23715 , n23716 , n23717 , n23718 , n23719 , n23720 , n23721 , n23722 , n23723 , n23724 , n23725 , n23726 , n23727 , n23728 , n23729 , n23730 , n23731 , n23732 , n23733 , n23734 , n23735 , n23736 , n23737 , n23738 , n23739 , n23740 , n23741 , n23742 , n23743 , n23744 , n23745 , n23746 , n23747 , n23748 , n23749 , n23750 , n23751 , n23752 , n23753 , n23754 , n23755 , n23756 , n23757 , n23758 , n23759 , n23760 , n23761 , n23762 , n23763 , n23764 , n23765 , n23766 , n23767 , n23768 , n23769 , n23770 , n23771 , n23772 , n23773 , n23774 , n23775 , n23776 , n23777 , n23778 , n23779 , n23780 , n23781 , n23782 , n23783 , n23784 , n23785 , n23786 , n23787 , n23788 , n23789 , n23790 , n23791 , n23792 , n23793 , n23794 , n23795 , n23796 , n23797 , n23798 , n23799 , n23800 , n23801 , n23802 , n23803 , n23804 , n23805 , n23806 , n23807 , n23808 , n23809 , n23810 , n23811 , n23812 , n23813 , n23814 , n23815 , n23816 , n23817 , n23818 , n23819 , n23820 , n23821 , n23822 , n23823 , n23824 , n23825 , n23826 , n23827 , n23828 , n23829 , n23830 , n23831 , n23832 , n23833 , n23834 , n23835 , n23836 , n23837 , n23838 , n23839 , n23840 , n23841 , n23842 , n23843 , n23844 , n23845 , n23846 , n23847 , n23848 , n23849 , n23850 , n23851 , n23852 , n23853 , n23854 , n23855 , n23856 , n23857 , n23858 , n23859 , n23860 , n23861 , n23862 , n23863 , n23864 , n23865 , n23866 , n23867 , n23868 , n23869 , n23870 , n23871 , n23872 , n23873 , n23874 , n23875 , n23876 , n23877 , n23878 , n23879 , n23880 , n23881 , n23882 , n23883 , n23884 , n23885 , n23886 , n23887 , n23888 , n23889 , n23890 , n23891 , n23892 , n23893 , n23894 , n23895 , n23896 , n23897 , n23898 , n23899 , n23900 , n23901 , n23902 , n23903 , n23904 , n23905 , n23906 , n23907 , n23908 , n23909 , n23910 , n23911 , n23912 , n23913 , n23914 , n23915 , n23916 , n23917 , n23918 , n23919 , n23920 , n23921 , n23922 , n23923 , n23924 , n23925 , n23926 , n23927 , n23928 , n23929 , n23930 , n23931 , n23932 , n23933 , n23934 , n23935 , n23936 , n23937 , n23938 , n23939 , n23940 , n23941 , n23942 , n23943 , n23944 , n23945 , n23946 , n23947 , n23948 , n23949 , n23950 , n23951 , n23952 , n23953 , n23954 , n23955 , n23956 , n23957 , n23958 , n23959 , n23960 , n23961 , n23962 , n23963 , n23964 , n23965 , n23966 , n23967 , n23968 , n23969 , n23970 , n23971 , n23972 , n23973 , n23974 , n23975 , n23976 , n23977 , n23978 , n23979 , n23980 , n23981 , n23982 , n23983 , n23984 , n23985 , n23986 , n23987 , n23988 , n23989 , n23990 , n23991 , n23992 , n23993 , n23994 , n23995 , n23996 , n23997 , n23998 , n23999 , n24000 , n24001 , n24002 , n24003 , n24004 , n24005 , n24006 , n24007 , n24008 , n24009 , n24010 , n24011 , n24012 , n24013 , n24014 , n24015 , n24016 , n24017 , n24018 , n24019 , n24020 , n24021 , n24022 , n24023 , n24024 , n24025 , n24026 , n24027 , n24028 , n24029 , n24030 , n24031 , n24032 , n24033 , n24034 , n24035 , n24036 , n24037 , n24038 , n24039 , n24040 , n24041 , n24042 , n24043 , n24044 , n24045 , n24046 , n24047 , n24048 , n24049 , n24050 , n24051 , n24052 , n24053 , n24054 , n24055 , n24056 , n24057 , n24058 , n24059 , n24060 , n24061 , n24062 , n24063 , n24064 , n24065 , n24066 , n24067 , n24068 , n24069 , n24070 , n24071 , n24072 , n24073 , n24074 , n24075 , n24076 , n24077 , n24078 , n24079 , n24080 , n24081 , n24082 , n24083 , n24084 , n24085 , n24086 , n24087 , n24088 , n24089 , n24090 , n24091 , n24092 , n24093 , n24094 , n24095 , n24096 , n24097 , n24098 , n24099 , n24100 , n24101 , n24102 , n24103 , n24104 , n24105 , n24106 , n24107 , n24108 , n24109 , n24110 , n24111 , n24112 , n24113 , n24114 , n24115 , n24116 , n24117 , n24118 , n24119 , n24120 , n24121 , n24122 , n24123 , n24124 , n24125 , n24126 , n24127 , n24128 , n24129 , n24130 , n24131 , n24132 , n24133 , n24134 , n24135 , n24136 , n24137 , n24138 , n24139 , n24140 , n24141 , n24142 , n24143 , n24144 , n24145 , n24146 , n24147 , n24148 , n24149 , n24150 , n24151 , n24152 , n24153 , n24154 , n24155 , n24156 , n24157 , n24158 , n24159 , n24160 , n24161 , n24162 , n24163 , n24164 , n24165 , n24166 , n24167 , n24168 , n24169 , n24170 , n24171 , n24172 , n24173 , n24174 , n24175 , n24176 , n24177 , n24178 , n24179 , n24180 , n24181 , n24182 , n24183 , n24184 , n24185 , n24186 , n24187 , n24188 , n24189 , n24190 , n24191 , n24192 , n24193 , n24194 , n24195 , n24196 , n24197 , n24198 , n24199 , n24200 , n24201 , n24202 , n24203 , n24204 , n24205 , n24206 , n24207 , n24208 , n24209 , n24210 , n24211 , n24212 , n24213 , n24214 , n24215 , n24216 , n24217 , n24218 , n24219 , n24220 , n24221 , n24222 , n24223 , n24224 , n24225 , n24226 , n24227 , n24228 , n24229 , n24230 , n24231 , n24232 , n24233 , n24234 , n24235 , n24236 , n24237 , n24238 , n24239 , n24240 , n24241 , n24242 , n24243 , n24244 , n24245 , n24246 , n24247 , n24248 , n24249 , n24250 , n24251 , n24252 , n24253 , n24254 , n24255 , n24256 , n24257 , n24258 , n24259 , n24260 , n24261 , n24262 , n24263 , n24264 , n24265 , n24266 , n24267 , n24268 , n24269 , n24270 , n24271 , n24272 , n24273 , n24274 , n24275 , n24276 , n24277 , n24278 , n24279 , n24280 , n24281 , n24282 , n24283 , n24284 , n24285 , n24286 , n24287 , n24288 , n24289 , n24290 , n24291 , n24292 , n24293 , n24294 , n24295 , n24296 , n24297 , n24298 , n24299 , n24300 , n24301 , n24302 , n24303 , n24304 , n24305 , n24306 , n24307 , n24308 , n24309 , n24310 , n24311 , n24312 , n24313 , n24314 , n24315 , n24316 , n24317 , n24318 , n24319 , n24320 , n24321 , n24322 , n24323 , n24324 , n24325 , n24326 , n24327 , n24328 , n24329 , n24330 , n24331 , n24332 , n24333 , n24334 , n24335 , n24336 , n24337 , n24338 , n24339 , n24340 , n24341 , n24342 , n24343 , n24344 , n24345 , n24346 , n24347 , n24348 , n24349 , n24350 , n24351 , n24352 , n24353 , n24354 , n24355 , n24356 , n24357 , n24358 , n24359 , n24360 , n24361 , n24362 , n24363 , n24364 , n24365 , n24366 , n24367 , n24368 , n24369 , n24370 , n24371 , n24372 , n24373 , n24374 , n24375 , n24376 , n24377 , n24378 , n24379 , n24380 , n24381 , n24382 , n24383 , n24384 , n24385 , n24386 , n24387 , n24388 , n24389 , n24390 , n24391 , n24392 , n24393 , n24394 , n24395 , n24396 , n24397 , n24398 , n24399 , n24400 , n24401 , n24402 , n24403 , n24404 , n24405 , n24406 , n24407 , n24408 , n24409 , n24410 , n24411 , n24412 , n24413 , n24414 , n24415 , n24416 , n24417 , n24418 , n24419 , n24420 , n24421 , n24422 , n24423 , n24424 , n24425 , n24426 , n24427 , n24428 , n24429 , n24430 , n24431 , n24432 , n24433 , n24434 , n24435 , n24436 , n24437 , n24438 , n24439 , n24440 , n24441 , n24442 , n24443 , n24444 , n24445 , n24446 , n24447 , n24448 , n24449 , n24450 , n24451 , n24452 , n24453 , n24454 , n24455 , n24456 , n24457 , n24458 , n24459 , n24460 , n24461 , n24462 , n24463 , n24464 , n24465 , n24466 , n24467 , n24468 , n24469 , n24470 , n24471 , n24472 , n24473 , n24474 , n24475 , n24476 , n24477 , n24478 , n24479 , n24480 , n24481 , n24482 , n24483 , n24484 , n24485 , n24486 , n24487 , n24488 , n24489 , n24490 , n24491 , n24492 , n24493 , n24494 , n24495 , n24496 , n24497 , n24498 , n24499 , n24500 , n24501 , n24502 , n24503 , n24504 , n24505 , n24506 , n24507 , n24508 , n24509 , n24510 , n24511 , n24512 , n24513 , n24514 , n24515 , n24516 , n24517 , n24518 , n24519 , n24520 , n24521 , n24522 , n24523 , n24524 , n24525 , n24526 , n24527 , n24528 , n24529 , n24530 , n24531 , n24532 , n24533 , n24534 , n24535 , n24536 , n24537 , n24538 , n24539 , n24540 , n24541 , n24542 , n24543 , n24544 , n24545 , n24546 , n24547 , n24548 , n24549 , n24550 , n24551 , n24552 , n24553 , n24554 , n24555 , n24556 , n24557 , n24558 , n24559 , n24560 , n24561 , n24562 , n24563 , n24564 , n24565 , n24566 , n24567 , n24568 , n24569 , n24570 , n24571 , n24572 , n24573 , n24574 , n24575 , n24576 , n24577 , n24578 , n24579 , n24580 , n24581 , n24582 , n24583 , n24584 , n24585 , n24586 , n24587 , n24588 , n24589 , n24590 , n24591 , n24592 , n24593 , n24594 , n24595 , n24596 , n24597 , n24598 , n24599 , n24600 , n24601 , n24602 , n24603 , n24604 , n24605 , n24606 , n24607 , n24608 , n24609 , n24610 , n24611 , n24612 , n24613 , n24614 , n24615 , n24616 , n24617 , n24618 , n24619 , n24620 , n24621 , n24622 , n24623 , n24624 , n24625 , n24626 , n24627 , n24628 , n24629 , n24630 , n24631 , n24632 , n24633 , n24634 , n24635 , n24636 , n24637 , n24638 , n24639 , n24640 , n24641 , n24642 , n24643 , n24644 , n24645 , n24646 , n24647 , n24648 , n24649 , n24650 , n24651 , n24652 , n24653 , n24654 , n24655 , n24656 , n24657 , n24658 , n24659 , n24660 , n24661 , n24662 , n24663 , n24664 , n24665 , n24666 , n24667 , n24668 , n24669 , n24670 , n24671 , n24672 , n24673 , n24674 , n24675 , n24676 , n24677 , n24678 , n24679 , n24680 , n24681 , n24682 , n24683 , n24684 , n24685 , n24686 , n24687 , n24688 , n24689 , n24690 , n24691 , n24692 , n24693 , n24694 , n24695 , n24696 , n24697 , n24698 , n24699 , n24700 , n24701 , n24702 , n24703 , n24704 , n24705 , n24706 , n24707 , n24708 , n24709 , n24710 , n24711 , n24712 , n24713 , n24714 , n24715 , n24716 , n24717 , n24718 , n24719 , n24720 , n24721 , n24722 , n24723 , n24724 , n24725 , n24726 , n24727 , n24728 , n24729 , n24730 , n24731 , n24732 , n24733 , n24734 , n24735 , n24736 , n24737 , n24738 , n24739 , n24740 , n24741 , n24742 , n24743 , n24744 , n24745 , n24746 , n24747 , n24748 , n24749 , n24750 , n24751 , n24752 , n24753 , n24754 , n24755 , n24756 , n24757 , n24758 , n24759 , n24760 , n24761 , n24762 , n24763 , n24764 , n24765 , n24766 , n24767 , n24768 , n24769 , n24770 , n24771 , n24772 , n24773 , n24774 , n24775 , n24776 , n24777 , n24778 , n24779 , n24780 , n24781 , n24782 , n24783 , n24784 , n24785 , n24786 , n24787 , n24788 , n24789 , n24790 , n24791 , n24792 , n24793 , n24794 , n24795 , n24796 , n24797 , n24798 , n24799 , n24800 , n24801 , n24802 , n24803 , n24804 , n24805 , n24806 , n24807 , n24808 , n24809 , n24810 , n24811 , n24812 , n24813 , n24814 , n24815 , n24816 , n24817 , n24818 , n24819 , n24820 , n24821 , n24822 , n24823 , n24824 , n24825 , n24826 , n24827 , n24828 , n24829 , n24830 , n24831 , n24832 , n24833 , n24834 , n24835 , n24836 , n24837 , n24838 , n24839 , n24840 , n24841 , n24842 , n24843 , n24844 , n24845 , n24846 , n24847 , n24848 , n24849 , n24850 , n24851 , n24852 , n24853 , n24854 , n24855 , n24856 , n24857 , n24858 , n24859 , n24860 , n24861 , n24862 , n24863 , n24864 , n24865 , n24866 , n24867 , n24868 , n24869 , n24870 , n24871 , n24872 , n24873 , n24874 , n24875 , n24876 , n24877 , n24878 , n24879 , n24880 , n24881 , n24882 , n24883 , n24884 , n24885 , n24886 , n24887 , n24888 , n24889 , n24890 , n24891 , n24892 , n24893 , n24894 , n24895 , n24896 , n24897 , n24898 , n24899 , n24900 , n24901 , n24902 , n24903 , n24904 , n24905 , n24906 , n24907 , n24908 , n24909 , n24910 , n24911 , n24912 , n24913 , n24914 , n24915 , n24916 , n24917 , n24918 , n24919 , n24920 , n24921 , n24922 , n24923 , n24924 , n24925 , n24926 , n24927 , n24928 , n24929 , n24930 , n24931 , n24932 , n24933 , n24934 , n24935 , n24936 , n24937 , n24938 , n24939 , n24940 , n24941 , n24942 , n24943 , n24944 , n24945 , n24946 , n24947 , n24948 , n24949 , n24950 , n24951 , n24952 , n24953 , n24954 , n24955 , n24956 , n24957 , n24958 , n24959 , n24960 , n24961 , n24962 , n24963 , n24964 , n24965 , n24966 , n24967 , n24968 , n24969 , n24970 , n24971 , n24972 , n24973 , n24974 , n24975 , n24976 , n24977 , n24978 , n24979 , n24980 , n24981 , n24982 , n24983 , n24984 , n24985 , n24986 , n24987 , n24988 , n24989 , n24990 , n24991 , n24992 , n24993 , n24994 , n24995 , n24996 , n24997 , n24998 , n24999 , n25000 , n25001 , n25002 , n25003 , n25004 , n25005 , n25006 , n25007 , n25008 , n25009 , n25010 , n25011 , n25012 , n25013 , n25014 , n25015 , n25016 , n25017 , n25018 , n25019 , n25020 , n25021 , n25022 , n25023 , n25024 , n25025 , n25026 , n25027 , n25028 , n25029 , n25030 , n25031 , n25032 , n25033 , n25034 , n25035 , n25036 , n25037 , n25038 , n25039 , n25040 , n25041 , n25042 , n25043 , n25044 , n25045 , n25046 , n25047 , n25048 , n25049 , n25050 , n25051 , n25052 , n25053 , n25054 , n25055 , n25056 , n25057 , n25058 , n25059 , n25060 , n25061 , n25062 , n25063 , n25064 , n25065 , n25066 , n25067 , n25068 , n25069 , n25070 , n25071 , n25072 , n25073 , n25074 , n25075 , n25076 , n25077 , n25078 , n25079 , n25080 , n25081 , n25082 , n25083 , n25084 , n25085 , n25086 , n25087 , n25088 , n25089 , n25090 , n25091 , n25092 , n25093 , n25094 , n25095 , n25096 , n25097 , n25098 , n25099 , n25100 , n25101 , n25102 , n25103 , n25104 , n25105 , n25106 , n25107 , n25108 , n25109 , n25110 , n25111 , n25112 , n25113 , n25114 , n25115 , n25116 , n25117 , n25118 , n25119 , n25120 , n25121 , n25122 , n25123 , n25124 , n25125 , n25126 , n25127 , n25128 , n25129 , n25130 , n25131 , n25132 , n25133 , n25134 , n25135 , n25136 , n25137 , n25138 , n25139 , n25140 , n25141 , n25142 , n25143 , n25144 , n25145 , n25146 , n25147 , n25148 , n25149 , n25150 , n25151 , n25152 , n25153 , n25154 , n25155 , n25156 , n25157 , n25158 , n25159 , n25160 , n25161 , n25162 , n25163 , n25164 , n25165 , n25166 , n25167 , n25168 , n25169 , n25170 , n25171 , n25172 , n25173 , n25174 , n25175 , n25176 , n25177 , n25178 , n25179 , n25180 , n25181 , n25182 , n25183 , n25184 , n25185 , n25186 , n25187 , n25188 , n25189 , n25190 , n25191 , n25192 , n25193 , n25194 , n25195 , n25196 , n25197 , n25198 , n25199 , n25200 , n25201 , n25202 , n25203 , n25204 , n25205 , n25206 , n25207 , n25208 , n25209 , n25210 , n25211 , n25212 , n25213 , n25214 , n25215 , n25216 , n25217 , n25218 , n25219 , n25220 , n25221 , n25222 , n25223 , n25224 , n25225 , n25226 , n25227 , n25228 , n25229 , n25230 , n25231 , n25232 , n25233 , n25234 , n25235 , n25236 , n25237 , n25238 , n25239 , n25240 , n25241 , n25242 , n25243 , n25244 , n25245 , n25246 , n25247 , n25248 , n25249 , n25250 , n25251 , n25252 , n25253 , n25254 , n25255 , n25256 , n25257 , n25258 , n25259 , n25260 , n25261 , n25262 , n25263 , n25264 , n25265 , n25266 , n25267 , n25268 , n25269 , n25270 , n25271 , n25272 , n25273 , n25274 , n25275 , n25276 , n25277 , n25278 , n25279 , n25280 , n25281 , n25282 , n25283 , n25284 , n25285 , n25286 , n25287 , n25288 , n25289 , n25290 , n25291 , n25292 , n25293 , n25294 , n25295 , n25296 , n25297 , n25298 , n25299 , n25300 , n25301 , n25302 , n25303 , n25304 , n25305 , n25306 , n25307 , n25308 , n25309 , n25310 , n25311 , n25312 , n25313 , n25314 , n25315 , n25316 , n25317 , n25318 , n25319 , n25320 , n25321 , n25322 , n25323 , n25324 , n25325 , n25326 , n25327 , n25328 , n25329 , n25330 , n25331 , n25332 , n25333 , n25334 , n25335 , n25336 , n25337 , n25338 , n25339 , n25340 , n25341 , n25342 , n25343 , n25344 , n25345 , n25346 , n25347 , n25348 , n25349 , n25350 , n25351 , n25352 , n25353 , n25354 , n25355 , n25356 , n25357 , n25358 , n25359 , n25360 , n25361 , n25362 , n25363 , n25364 , n25365 , n25366 , n25367 , n25368 , n25369 , n25370 , n25371 , n25372 , n25373 , n25374 , n25375 , n25376 , n25377 , n25378 , n25379 , n25380 , n25381 , n25382 , n25383 , n25384 , n25385 , n25386 , n25387 , n25388 , n25389 , n25390 , n25391 , n25392 , n25393 , n25394 , n25395 , n25396 , n25397 , n25398 , n25399 , n25400 , n25401 , n25402 , n25403 , n25404 , n25405 , n25406 , n25407 , n25408 , n25409 , n25410 , n25411 , n25412 , n25413 , n25414 , n25415 , n25416 , n25417 , n25418 , n25419 , n25420 , n25421 , n25422 , n25423 , n25424 , n25425 , n25426 , n25427 , n25428 , n25429 , n25430 , n25431 , n25432 , n25433 , n25434 , n25435 , n25436 , n25437 , n25438 , n25439 , n25440 , n25441 , n25442 , n25443 , n25444 , n25445 , n25446 , n25447 , n25448 , n25449 , n25450 , n25451 , n25452 , n25453 , n25454 , n25455 , n25456 , n25457 , n25458 , n25459 , n25460 , n25461 , n25462 , n25463 , n25464 , n25465 , n25466 , n25467 , n25468 , n25469 , n25470 , n25471 , n25472 , n25473 , n25474 , n25475 , n25476 , n25477 , n25478 , n25479 , n25480 , n25481 , n25482 , n25483 , n25484 , n25485 , n25486 , n25487 , n25488 , n25489 , n25490 , n25491 , n25492 , n25493 , n25494 , n25495 , n25496 , n25497 , n25498 , n25499 , n25500 , n25501 , n25502 , n25503 , n25504 , n25505 , n25506 , n25507 , n25508 , n25509 , n25510 , n25511 , n25512 , n25513 , n25514 , n25515 , n25516 , n25517 , n25518 , n25519 , n25520 , n25521 , n25522 , n25523 , n25524 , n25525 , n25526 , n25527 , n25528 , n25529 , n25530 , n25531 , n25532 , n25533 , n25534 , n25535 , n25536 , n25537 , n25538 , n25539 , n25540 , n25541 , n25542 , n25543 , n25544 , n25545 , n25546 , n25547 , n25548 , n25549 , n25550 , n25551 , n25552 , n25553 , n25554 , n25555 , n25556 , n25557 , n25558 , n25559 , n25560 , n25561 , n25562 , n25563 , n25564 , n25565 , n25566 , n25567 , n25568 , n25569 , n25570 , n25571 , n25572 , n25573 , n25574 , n25575 , n25576 , n25577 , n25578 , n25579 , n25580 , n25581 , n25582 , n25583 , n25584 , n25585 , n25586 , n25587 , n25588 , n25589 , n25590 , n25591 , n25592 , n25593 , n25594 , n25595 , n25596 , n25597 , n25598 , n25599 , n25600 , n25601 , n25602 , n25603 , n25604 , n25605 , n25606 , n25607 , n25608 , n25609 , n25610 , n25611 , n25612 , n25613 , n25614 , n25615 , n25616 , n25617 , n25618 , n25619 , n25620 , n25621 , n25622 , n25623 , n25624 , n25625 , n25626 , n25627 , n25628 , n25629 , n25630 , n25631 , n25632 , n25633 , n25634 , n25635 , n25636 , n25637 , n25638 , n25639 , n25640 , n25641 , n25642 , n25643 , n25644 , n25645 , n25646 , n25647 , n25648 , n25649 , n25650 , n25651 , n25652 , n25653 , n25654 , n25655 , n25656 , n25657 , n25658 , n25659 , n25660 , n25661 , n25662 , n25663 , n25664 , n25665 , n25666 , n25667 , n25668 , n25669 , n25670 , n25671 , n25672 , n25673 , n25674 , n25675 , n25676 , n25677 , n25678 , n25679 , n25680 , n25681 , n25682 , n25683 , n25684 , n25685 , n25686 , n25687 , n25688 , n25689 , n25690 , n25691 , n25692 , n25693 , n25694 , n25695 , n25696 , n25697 , n25698 , n25699 , n25700 , n25701 , n25702 , n25703 , n25704 , n25705 , n25706 , n25707 , n25708 , n25709 , n25710 , n25711 , n25712 , n25713 , n25714 , n25715 , n25716 , n25717 , n25718 , n25719 , n25720 , n25721 , n25722 , n25723 , n25724 , n25725 , n25726 , n25727 , n25728 , n25729 , n25730 , n25731 , n25732 , n25733 , n25734 , n25735 , n25736 , n25737 , n25738 , n25739 , n25740 , n25741 , n25742 , n25743 , n25744 , n25745 , n25746 , n25747 , n25748 , n25749 , n25750 , n25751 , n25752 , n25753 , n25754 , n25755 , n25756 , n25757 , n25758 , n25759 , n25760 , n25761 , n25762 , n25763 , n25764 , n25765 , n25766 , n25767 , n25768 , n25769 , n25770 , n25771 , n25772 , n25773 , n25774 , n25775 , n25776 , n25777 , n25778 , n25779 , n25780 , n25781 , n25782 , n25783 , n25784 , n25785 , n25786 , n25787 , n25788 , n25789 , n25790 , n25791 , n25792 , n25793 , n25794 , n25795 , n25796 , n25797 , n25798 , n25799 , n25800 , n25801 , n25802 , n25803 , n25804 , n25805 , n25806 , n25807 , n25808 , n25809 , n25810 , n25811 , n25812 , n25813 , n25814 , n25815 , n25816 , n25817 , n25818 , n25819 , n25820 , n25821 , n25822 , n25823 , n25824 , n25825 , n25826 , n25827 , n25828 , n25829 , n25830 , n25831 , n25832 , n25833 , n25834 , n25835 , n25836 , n25837 , n25838 , n25839 , n25840 , n25841 , n25842 , n25843 , n25844 , n25845 , n25846 , n25847 , n25848 , n25849 , n25850 , n25851 , n25852 , n25853 , n25854 , n25855 , n25856 , n25857 , n25858 , n25859 , n25860 , n25861 , n25862 , n25863 , n25864 , n25865 , n25866 , n25867 , n25868 , n25869 , n25870 , n25871 , n25872 , n25873 , n25874 , n25875 , n25876 , n25877 , n25878 , n25879 , n25880 , n25881 , n25882 , n25883 , n25884 , n25885 , n25886 , n25887 , n25888 , n25889 , n25890 , n25891 , n25892 , n25893 , n25894 , n25895 , n25896 , n25897 , n25898 , n25899 , n25900 , n25901 , n25902 , n25903 , n25904 , n25905 , n25906 , n25907 , n25908 , n25909 , n25910 , n25911 , n25912 , n25913 , n25914 , n25915 , n25916 , n25917 , n25918 , n25919 , n25920 , n25921 , n25922 , n25923 , n25924 , n25925 , n25926 , n25927 , n25928 , n25929 , n25930 , n25931 , n25932 , n25933 , n25934 , n25935 , n25936 , n25937 , n25938 , n25939 , n25940 , n25941 , n25942 , n25943 , n25944 , n25945 , n25946 , n25947 , n25948 , n25949 , n25950 , n25951 , n25952 , n25953 , n25954 , n25955 , n25956 , n25957 , n25958 , n25959 , n25960 , n25961 , n25962 , n25963 , n25964 , n25965 , n25966 , n25967 , n25968 , n25969 , n25970 , n25971 , n25972 , n25973 , n25974 , n25975 , n25976 , n25977 , n25978 , n25979 , n25980 , n25981 , n25982 , n25983 , n25984 , n25985 , n25986 , n25987 , n25988 , n25989 , n25990 , n25991 , n25992 , n25993 , n25994 , n25995 , n25996 , n25997 , n25998 , n25999 , n26000 , n26001 , n26002 , n26003 , n26004 , n26005 , n26006 , n26007 , n26008 , n26009 , n26010 , n26011 , n26012 , n26013 , n26014 , n26015 , n26016 , n26017 , n26018 , n26019 , n26020 , n26021 , n26022 , n26023 , n26024 , n26025 , n26026 , n26027 , n26028 , n26029 , n26030 , n26031 , n26032 , n26033 , n26034 , n26035 , n26036 , n26037 , n26038 , n26039 , n26040 , n26041 , n26042 , n26043 , n26044 , n26045 , n26046 , n26047 , n26048 , n26049 , n26050 , n26051 , n26052 , n26053 , n26054 , n26055 , n26056 , n26057 , n26058 , n26059 , n26060 , n26061 , n26062 , n26063 , n26064 , n26065 , n26066 , n26067 , n26068 , n26069 , n26070 , n26071 , n26072 , n26073 , n26074 , n26075 , n26076 , n26077 , n26078 , n26079 , n26080 , n26081 , n26082 , n26083 , n26084 , n26085 , n26086 , n26087 , n26088 , n26089 , n26090 , n26091 , n26092 , n26093 , n26094 , n26095 , n26096 , n26097 , n26098 , n26099 , n26100 , n26101 , n26102 , n26103 , n26104 , n26105 , n26106 , n26107 , n26108 , n26109 , n26110 , n26111 , n26112 , n26113 , n26114 , n26115 , n26116 , n26117 , n26118 , n26119 , n26120 , n26121 , n26122 , n26123 , n26124 , n26125 , n26126 , n26127 , n26128 , n26129 , n26130 , n26131 , n26132 , n26133 , n26134 , n26135 , n26136 , n26137 , n26138 , n26139 , n26140 , n26141 , n26142 , n26143 , n26144 , n26145 , n26146 , n26147 , n26148 , n26149 , n26150 , n26151 , n26152 , n26153 , n26154 , n26155 , n26156 , n26157 , n26158 , n26159 , n26160 , n26161 , n26162 , n26163 , n26164 , n26165 , n26166 , n26167 , n26168 , n26169 , n26170 , n26171 , n26172 , n26173 , n26174 , n26175 , n26176 , n26177 , n26178 , n26179 , n26180 , n26181 , n26182 , n26183 , n26184 , n26185 , n26186 , n26187 , n26188 , n26189 , n26190 , n26191 , n26192 , n26193 , n26194 , n26195 , n26196 , n26197 , n26198 , n26199 , n26200 , n26201 , n26202 , n26203 , n26204 , n26205 , n26206 , n26207 , n26208 , n26209 , n26210 , n26211 , n26212 , n26213 , n26214 , n26215 , n26216 , n26217 , n26218 , n26219 , n26220 , n26221 , n26222 , n26223 , n26224 , n26225 , n26226 , n26227 , n26228 , n26229 , n26230 , n26231 , n26232 , n26233 , n26234 , n26235 , n26236 , n26237 , n26238 , n26239 , n26240 , n26241 , n26242 , n26243 , n26244 , n26245 , n26246 , n26247 , n26248 , n26249 , n26250 , n26251 , n26252 , n26253 , n26254 , n26255 , n26256 , n26257 , n26258 , n26259 , n26260 , n26261 , n26262 , n26263 , n26264 , n26265 , n26266 , n26267 , n26268 , n26269 , n26270 , n26271 , n26272 , n26273 , n26274 , n26275 , n26276 , n26277 , n26278 , n26279 , n26280 , n26281 , n26282 , n26283 , n26284 , n26285 , n26286 , n26287 , n26288 , n26289 , n26290 , n26291 , n26292 , n26293 , n26294 , n26295 , n26296 , n26297 , n26298 , n26299 , n26300 , n26301 , n26302 , n26303 , n26304 , n26305 , n26306 , n26307 , n26308 , n26309 , n26310 , n26311 , n26312 , n26313 , n26314 , n26315 , n26316 , n26317 , n26318 , n26319 , n26320 , n26321 , n26322 , n26323 , n26324 , n26325 , n26326 , n26327 , n26328 , n26329 , n26330 , n26331 , n26332 , n26333 , n26334 , n26335 , n26336 , n26337 , n26338 , n26339 , n26340 , n26341 , n26342 , n26343 , n26344 , n26345 , n26346 , n26347 , n26348 , n26349 , n26350 , n26351 , n26352 , n26353 , n26354 , n26355 , n26356 , n26357 , n26358 , n26359 , n26360 , n26361 , n26362 , n26363 , n26364 , n26365 , n26366 , n26367 , n26368 , n26369 , n26370 , n26371 , n26372 , n26373 , n26374 , n26375 , n26376 , n26377 , n26378 , n26379 , n26380 , n26381 , n26382 , n26383 , n26384 , n26385 , n26386 , n26387 , n26388 , n26389 , n26390 , n26391 , n26392 , n26393 , n26394 , n26395 , n26396 , n26397 , n26398 , n26399 , n26400 , n26401 , n26402 , n26403 , n26404 , n26405 , n26406 , n26407 , n26408 , n26409 , n26410 , n26411 , n26412 , n26413 , n26414 , n26415 , n26416 , n26417 , n26418 , n26419 , n26420 , n26421 , n26422 , n26423 , n26424 , n26425 , n26426 , n26427 , n26428 , n26429 , n26430 , n26431 , n26432 , n26433 , n26434 , n26435 , n26436 , n26437 , n26438 , n26439 , n26440 , n26441 , n26442 , n26443 , n26444 , n26445 , n26446 , n26447 , n26448 , n26449 , n26450 , n26451 , n26452 , n26453 , n26454 , n26455 , n26456 , n26457 , n26458 , n26459 , n26460 , n26461 , n26462 , n26463 , n26464 , n26465 , n26466 , n26467 , n26468 , n26469 , n26470 , n26471 , n26472 , n26473 , n26474 , n26475 , n26476 , n26477 , n26478 , n26479 , n26480 , n26481 , n26482 , n26483 , n26484 , n26485 , n26486 , n26487 , n26488 , n26489 , n26490 , n26491 , n26492 , n26493 , n26494 , n26495 , n26496 , n26497 , n26498 , n26499 , n26500 , n26501 , n26502 , n26503 , n26504 , n26505 , n26506 , n26507 , n26508 , n26509 , n26510 , n26511 , n26512 , n26513 , n26514 , n26515 , n26516 , n26517 , n26518 , n26519 , n26520 , n26521 , n26522 , n26523 , n26524 , n26525 , n26526 , n26527 , n26528 , n26529 , n26530 , n26531 , n26532 , n26533 , n26534 , n26535 , n26536 , n26537 , n26538 , n26539 , n26540 , n26541 , n26542 , n26543 , n26544 , n26545 , n26546 , n26547 , n26548 , n26549 , n26550 , n26551 , n26552 , n26553 , n26554 , n26555 , n26556 , n26557 , n26558 , n26559 , n26560 , n26561 , n26562 , n26563 , n26564 , n26565 , n26566 , n26567 , n26568 , n26569 , n26570 , n26571 , n26572 , n26573 , n26574 , n26575 , n26576 , n26577 , n26578 , n26579 , n26580 , n26581 , n26582 , n26583 , n26584 , n26585 , n26586 , n26587 , n26588 , n26589 , n26590 , n26591 , n26592 , n26593 , n26594 , n26595 , n26596 , n26597 , n26598 , n26599 , n26600 , n26601 , n26602 , n26603 , n26604 , n26605 , n26606 , n26607 , n26608 , n26609 , n26610 , n26611 , n26612 , n26613 , n26614 , n26615 , n26616 , n26617 , n26618 , n26619 , n26620 , n26621 , n26622 , n26623 , n26624 , n26625 , n26626 , n26627 , n26628 , n26629 , n26630 , n26631 , n26632 , n26633 , n26634 , n26635 , n26636 , n26637 , n26638 , n26639 , n26640 , n26641 , n26642 , n26643 , n26644 , n26645 , n26646 , n26647 , n26648 , n26649 , n26650 , n26651 , n26652 , n26653 , n26654 , n26655 , n26656 , n26657 , n26658 , n26659 , n26660 , n26661 , n26662 , n26663 , n26664 , n26665 , n26666 , n26667 , n26668 , n26669 , n26670 , n26671 , n26672 , n26673 , n26674 , n26675 , n26676 , n26677 , n26678 , n26679 , n26680 , n26681 , n26682 , n26683 , n26684 , n26685 , n26686 , n26687 , n26688 , n26689 , n26690 , n26691 , n26692 , n26693 , n26694 , n26695 , n26696 , n26697 , n26698 , n26699 , n26700 , n26701 , n26702 , n26703 , n26704 , n26705 , n26706 , n26707 , n26708 , n26709 , n26710 , n26711 , n26712 , n26713 , n26714 , n26715 , n26716 , n26717 , n26718 , n26719 , n26720 , n26721 , n26722 , n26723 , n26724 , n26725 , n26726 , n26727 , n26728 , n26729 , n26730 , n26731 , n26732 , n26733 , n26734 , n26735 , n26736 , n26737 , n26738 , n26739 , n26740 , n26741 , n26742 , n26743 , n26744 , n26745 , n26746 , n26747 , n26748 , n26749 , n26750 , n26751 , n26752 , n26753 , n26754 , n26755 , n26756 , n26757 , n26758 , n26759 , n26760 , n26761 , n26762 , n26763 , n26764 , n26765 , n26766 , n26767 , n26768 , n26769 , n26770 , n26771 , n26772 , n26773 , n26774 , n26775 , n26776 , n26777 , n26778 , n26779 , n26780 , n26781 , n26782 , n26783 , n26784 , n26785 , n26786 , n26787 , n26788 , n26789 , n26790 , n26791 , n26792 , n26793 , n26794 , n26795 , n26796 , n26797 , n26798 , n26799 , n26800 , n26801 , n26802 , n26803 , n26804 , n26805 , n26806 , n26807 , n26808 , n26809 , n26810 , n26811 , n26812 , n26813 , n26814 , n26815 , n26816 , n26817 , n26818 , n26819 , n26820 , n26821 , n26822 , n26823 , n26824 , n26825 , n26826 , n26827 , n26828 , n26829 , n26830 , n26831 , n26832 , n26833 , n26834 , n26835 , n26836 , n26837 , n26838 , n26839 , n26840 , n26841 , n26842 , n26843 , n26844 , n26845 , n26846 , n26847 , n26848 , n26849 , n26850 , n26851 , n26852 , n26853 , n26854 , n26855 , n26856 , n26857 , n26858 , n26859 , n26860 , n26861 , n26862 , n26863 , n26864 , n26865 , n26866 , n26867 , n26868 , n26869 , n26870 , n26871 , n26872 , n26873 , n26874 , n26875 , n26876 , n26877 , n26878 , n26879 , n26880 , n26881 , n26882 , n26883 , n26884 , n26885 , n26886 , n26887 , n26888 , n26889 , n26890 , n26891 , n26892 , n26893 , n26894 , n26895 , n26896 , n26897 , n26898 , n26899 , n26900 , n26901 , n26902 , n26903 , n26904 , n26905 , n26906 , n26907 , n26908 , n26909 , n26910 , n26911 , n26912 , n26913 , n26914 , n26915 , n26916 , n26917 , n26918 , n26919 , n26920 , n26921 , n26922 , n26923 , n26924 , n26925 , n26926 , n26927 , n26928 , n26929 , n26930 , n26931 , n26932 , n26933 , n26934 , n26935 , n26936 , n26937 , n26938 , n26939 , n26940 , n26941 , n26942 , n26943 , n26944 , n26945 , n26946 , n26947 , n26948 , n26949 , n26950 , n26951 , n26952 , n26953 , n26954 , n26955 , n26956 , n26957 , n26958 , n26959 , n26960 , n26961 , n26962 , n26963 , n26964 , n26965 , n26966 , n26967 , n26968 , n26969 , n26970 , n26971 , n26972 , n26973 , n26974 , n26975 , n26976 , n26977 , n26978 , n26979 , n26980 , n26981 , n26982 , n26983 , n26984 , n26985 , n26986 , n26987 , n26988 , n26989 , n26990 , n26991 , n26992 , n26993 , n26994 , n26995 , n26996 , n26997 , n26998 , n26999 , n27000 , n27001 , n27002 , n27003 , n27004 , n27005 , n27006 , n27007 , n27008 , n27009 , n27010 , n27011 , n27012 , n27013 , n27014 , n27015 , n27016 , n27017 , n27018 , n27019 , n27020 , n27021 , n27022 , n27023 , n27024 , n27025 , n27026 , n27027 , n27028 , n27029 , n27030 , n27031 , n27032 , n27033 , n27034 , n27035 , n27036 , n27037 , n27038 , n27039 , n27040 , n27041 , n27042 , n27043 , n27044 , n27045 , n27046 , n27047 , n27048 , n27049 , n27050 , n27051 , n27052 , n27053 , n27054 , n27055 , n27056 , n27057 , n27058 , n27059 , n27060 , n27061 , n27062 , n27063 , n27064 , n27065 , n27066 , n27067 , n27068 , n27069 , n27070 , n27071 , n27072 , n27073 , n27074 , n27075 , n27076 , n27077 , n27078 , n27079 , n27080 , n27081 , n27082 , n27083 , n27084 , n27085 , n27086 , n27087 , n27088 , n27089 , n27090 , n27091 , n27092 , n27093 , n27094 , n27095 , n27096 , n27097 , n27098 , n27099 , n27100 , n27101 , n27102 , n27103 , n27104 , n27105 , n27106 , n27107 , n27108 , n27109 , n27110 , n27111 , n27112 , n27113 , n27114 , n27115 , n27116 , n27117 , n27118 , n27119 , n27120 , n27121 , n27122 , n27123 , n27124 , n27125 , n27126 , n27127 , n27128 , n27129 , n27130 , n27131 , n27132 , n27133 , n27134 , n27135 , n27136 , n27137 , n27138 , n27139 , n27140 , n27141 , n27142 , n27143 , n27144 , n27145 , n27146 , n27147 , n27148 , n27149 , n27150 , n27151 , n27152 , n27153 , n27154 , n27155 , n27156 , n27157 , n27158 , n27159 , n27160 , n27161 , n27162 , n27163 , n27164 , n27165 , n27166 , n27167 , n27168 , n27169 , n27170 , n27171 , n27172 , n27173 , n27174 , n27175 , n27176 , n27177 , n27178 , n27179 , n27180 , n27181 , n27182 , n27183 , n27184 , n27185 , n27186 , n27187 , n27188 , n27189 , n27190 , n27191 , n27192 , n27193 , n27194 , n27195 , n27196 , n27197 , n27198 , n27199 , n27200 , n27201 , n27202 , n27203 , n27204 , n27205 , n27206 , n27207 , n27208 , n27209 , n27210 , n27211 , n27212 , n27213 , n27214 , n27215 , n27216 , n27217 , n27218 , n27219 , n27220 , n27221 , n27222 , n27223 , n27224 , n27225 , n27226 , n27227 , n27228 , n27229 , n27230 , n27231 , n27232 , n27233 , n27234 , n27235 , n27236 , n27237 , n27238 , n27239 , n27240 , n27241 , n27242 , n27243 , n27244 , n27245 , n27246 , n27247 , n27248 , n27249 , n27250 , n27251 , n27252 , n27253 , n27254 , n27255 , n27256 , n27257 , n27258 , n27259 , n27260 , n27261 , n27262 , n27263 , n27264 , n27265 , n27266 , n27267 , n27268 , n27269 , n27270 , n27271 , n27272 , n27273 , n27274 , n27275 , n27276 , n27277 , n27278 , n27279 , n27280 , n27281 , n27282 , n27283 , n27284 , n27285 , n27286 , n27287 , n27288 , n27289 , n27290 , n27291 , n27292 , n27293 , n27294 , n27295 , n27296 , n27297 , n27298 , n27299 , n27300 , n27301 , n27302 , n27303 , n27304 , n27305 , n27306 , n27307 , n27308 , n27309 , n27310 , n27311 , n27312 , n27313 , n27314 , n27315 , n27316 , n27317 , n27318 , n27319 , n27320 , n27321 , n27322 , n27323 , n27324 , n27325 , n27326 , n27327 , n27328 , n27329 , n27330 , n27331 , n27332 , n27333 , n27334 , n27335 , n27336 , n27337 , n27338 , n27339 , n27340 , n27341 , n27342 , n27343 , n27344 , n27345 , n27346 , n27347 , n27348 , n27349 , n27350 , n27351 , n27352 , n27353 , n27354 , n27355 , n27356 , n27357 , n27358 , n27359 , n27360 , n27361 , n27362 , n27363 , n27364 , n27365 , n27366 , n27367 , n27368 , n27369 , n27370 , n27371 , n27372 , n27373 , n27374 , n27375 , n27376 , n27377 , n27378 , n27379 , n27380 , n27381 , n27382 , n27383 , n27384 , n27385 , n27386 , n27387 , n27388 , n27389 , n27390 , n27391 , n27392 , n27393 , n27394 , n27395 , n27396 , n27397 , n27398 , n27399 , n27400 , n27401 , n27402 , n27403 , n27404 , n27405 , n27406 , n27407 , n27408 , n27409 , n27410 , n27411 , n27412 , n27413 , n27414 , n27415 , n27416 , n27417 , n27418 , n27419 , n27420 , n27421 , n27422 , n27423 , n27424 , n27425 , n27426 , n27427 , n27428 , n27429 , n27430 , n27431 , n27432 , n27433 , n27434 , n27435 , n27436 , n27437 , n27438 , n27439 , n27440 , n27441 , n27442 , n27443 , n27444 , n27445 , n27446 , n27447 , n27448 , n27449 , n27450 , n27451 , n27452 , n27453 , n27454 , n27455 , n27456 , n27457 , n27458 , n27459 , n27460 , n27461 , n27462 , n27463 , n27464 , n27465 , n27466 , n27467 , n27468 , n27469 , n27470 , n27471 , n27472 , n27473 , n27474 , n27475 , n27476 , n27477 , n27478 , n27479 , n27480 , n27481 , n27482 , n27483 , n27484 , n27485 , n27486 , n27487 , n27488 , n27489 , n27490 , n27491 , n27492 , n27493 , n27494 , n27495 , n27496 , n27497 , n27498 , n27499 , n27500 , n27501 , n27502 , n27503 , n27504 , n27505 , n27506 , n27507 , n27508 , n27509 , n27510 , n27511 , n27512 , n27513 , n27514 , n27515 , n27516 , n27517 , n27518 , n27519 , n27520 , n27521 , n27522 , n27523 , n27524 , n27525 , n27526 , n27527 , n27528 , n27529 , n27530 , n27531 , n27532 , n27533 , n27534 , n27535 , n27536 , n27537 , n27538 , n27539 , n27540 , n27541 , n27542 , n27543 , n27544 , n27545 , n27546 , n27547 , n27548 , n27549 , n27550 , n27551 , n27552 , n27553 , n27554 , n27555 , n27556 , n27557 , n27558 , n27559 , n27560 , n27561 , n27562 , n27563 , n27564 , n27565 , n27566 , n27567 , n27568 , n27569 , n27570 , n27571 , n27572 , n27573 , n27574 , n27575 , n27576 , n27577 , n27578 , n27579 , n27580 , n27581 , n27582 , n27583 , n27584 , n27585 , n27586 , n27587 , n27588 , n27589 , n27590 , n27591 , n27592 , n27593 , n27594 , n27595 , n27596 , n27597 , n27598 , n27599 , n27600 , n27601 , n27602 , n27603 , n27604 , n27605 , n27606 , n27607 , n27608 , n27609 , n27610 , n27611 , n27612 , n27613 , n27614 , n27615 , n27616 , n27617 , n27618 , n27619 , n27620 , n27621 , n27622 , n27623 , n27624 , n27625 , n27626 , n27627 , n27628 , n27629 , n27630 , n27631 , n27632 , n27633 , n27634 , n27635 , n27636 , n27637 , n27638 , n27639 , n27640 , n27641 , n27642 , n27643 , n27644 , n27645 , n27646 , n27647 , n27648 , n27649 , n27650 , n27651 , n27652 , n27653 , n27654 , n27655 , n27656 , n27657 , n27658 , n27659 , n27660 , n27661 , n27662 , n27663 , n27664 , n27665 , n27666 , n27667 , n27668 , n27669 , n27670 , n27671 , n27672 , n27673 , n27674 , n27675 , n27676 , n27677 , n27678 , n27679 , n27680 , n27681 , n27682 , n27683 , n27684 , n27685 , n27686 , n27687 , n27688 , n27689 , n27690 , n27691 , n27692 , n27693 , n27694 , n27695 , n27696 , n27697 , n27698 , n27699 , n27700 , n27701 , n27702 , n27703 , n27704 , n27705 , n27706 , n27707 , n27708 , n27709 , n27710 , n27711 , n27712 , n27713 , n27714 , n27715 , n27716 , n27717 , n27718 , n27719 , n27720 , n27721 , n27722 , n27723 , n27724 , n27725 , n27726 , n27727 , n27728 , n27729 , n27730 , n27731 , n27732 , n27733 , n27734 , n27735 , n27736 , n27737 , n27738 , n27739 , n27740 , n27741 , n27742 , n27743 , n27744 , n27745 , n27746 , n27747 , n27748 , n27749 , n27750 , n27751 , n27752 , n27753 , n27754 , n27755 , n27756 , n27757 , n27758 , n27759 , n27760 , n27761 , n27762 , n27763 , n27764 , n27765 , n27766 , n27767 , n27768 , n27769 , n27770 , n27771 , n27772 , n27773 , n27774 , n27775 , n27776 , n27777 , n27778 , n27779 , n27780 , n27781 , n27782 , n27783 , n27784 , n27785 , n27786 , n27787 , n27788 , n27789 , n27790 , n27791 , n27792 , n27793 , n27794 , n27795 , n27796 , n27797 , n27798 , n27799 , n27800 , n27801 , n27802 , n27803 , n27804 , n27805 , n27806 , n27807 , n27808 , n27809 , n27810 , n27811 , n27812 , n27813 , n27814 , n27815 , n27816 , n27817 , n27818 , n27819 , n27820 , n27821 , n27822 , n27823 , n27824 , n27825 , n27826 , n27827 , n27828 , n27829 , n27830 , n27831 , n27832 , n27833 , n27834 , n27835 , n27836 , n27837 , n27838 , n27839 , n27840 , n27841 , n27842 , n27843 , n27844 , n27845 , n27846 , n27847 , n27848 , n27849 , n27850 , n27851 , n27852 , n27853 , n27854 , n27855 , n27856 , n27857 , n27858 , n27859 , n27860 , n27861 , n27862 , n27863 , n27864 , n27865 , n27866 , n27867 , n27868 , n27869 , n27870 , n27871 , n27872 , n27873 , n27874 , n27875 , n27876 , n27877 , n27878 , n27879 , n27880 , n27881 , n27882 , n27883 , n27884 , n27885 , n27886 , n27887 , n27888 , n27889 , n27890 , n27891 , n27892 , n27893 , n27894 , n27895 , n27896 , n27897 , n27898 , n27899 , n27900 , n27901 , n27902 , n27903 , n27904 , n27905 , n27906 , n27907 , n27908 , n27909 , n27910 , n27911 , n27912 , n27913 , n27914 , n27915 , n27916 , n27917 , n27918 , n27919 , n27920 , n27921 , n27922 , n27923 , n27924 , n27925 , n27926 , n27927 , n27928 , n27929 , n27930 , n27931 , n27932 , n27933 , n27934 , n27935 , n27936 , n27937 , n27938 , n27939 , n27940 , n27941 , n27942 , n27943 , n27944 , n27945 , n27946 , n27947 , n27948 , n27949 , n27950 , n27951 , n27952 , n27953 , n27954 , n27955 , n27956 , n27957 , n27958 , n27959 , n27960 , n27961 , n27962 , n27963 , n27964 , n27965 , n27966 , n27967 , n27968 , n27969 , n27970 , n27971 , n27972 , n27973 , n27974 , n27975 , n27976 , n27977 , n27978 , n27979 , n27980 , n27981 , n27982 , n27983 , n27984 , n27985 , n27986 , n27987 , n27988 , n27989 , n27990 , n27991 , n27992 , n27993 , n27994 , n27995 , n27996 , n27997 , n27998 , n27999 , n28000 , n28001 , n28002 , n28003 , n28004 , n28005 , n28006 , n28007 , n28008 , n28009 , n28010 , n28011 , n28012 , n28013 , n28014 , n28015 , n28016 , n28017 , n28018 , n28019 , n28020 , n28021 , n28022 , n28023 , n28024 , n28025 , n28026 , n28027 , n28028 , n28029 , n28030 , n28031 , n28032 , n28033 , n28034 , n28035 , n28036 , n28037 , n28038 , n28039 , n28040 , n28041 , n28042 , n28043 , n28044 , n28045 , n28046 , n28047 , n28048 , n28049 , n28050 , n28051 , n28052 , n28053 , n28054 , n28055 , n28056 , n28057 , n28058 , n28059 , n28060 , n28061 , n28062 , n28063 , n28064 , n28065 , n28066 , n28067 , n28068 , n28069 , n28070 , n28071 , n28072 , n28073 , n28074 , n28075 , n28076 , n28077 , n28078 , n28079 , n28080 , n28081 , n28082 , n28083 , n28084 , n28085 , n28086 , n28087 , n28088 , n28089 , n28090 , n28091 , n28092 , n28093 , n28094 , n28095 , n28096 , n28097 , n28098 , n28099 , n28100 , n28101 , n28102 , n28103 , n28104 , n28105 , n28106 , n28107 , n28108 , n28109 , n28110 , n28111 , n28112 , n28113 , n28114 , n28115 , n28116 , n28117 , n28118 , n28119 , n28120 , n28121 , n28122 , n28123 , n28124 , n28125 , n28126 , n28127 , n28128 , n28129 , n28130 , n28131 , n28132 , n28133 , n28134 , n28135 , n28136 , n28137 , n28138 , n28139 , n28140 , n28141 , n28142 , n28143 , n28144 , n28145 , n28146 , n28147 , n28148 , n28149 , n28150 , n28151 , n28152 , n28153 , n28154 , n28155 , n28156 , n28157 , n28158 , n28159 , n28160 , n28161 , n28162 , n28163 , n28164 , n28165 , n28166 , n28167 , n28168 , n28169 , n28170 , n28171 , n28172 , n28173 , n28174 , n28175 , n28176 , n28177 , n28178 , n28179 , n28180 , n28181 , n28182 , n28183 , n28184 , n28185 , n28186 , n28187 , n28188 , n28189 , n28190 , n28191 , n28192 , n28193 , n28194 , n28195 , n28196 , n28197 , n28198 , n28199 , n28200 , n28201 , n28202 , n28203 , n28204 , n28205 , n28206 , n28207 , n28208 , n28209 , n28210 , n28211 , n28212 , n28213 , n28214 , n28215 , n28216 , n28217 , n28218 , n28219 , n28220 , n28221 , n28222 , n28223 , n28224 , n28225 , n28226 , n28227 , n28228 , n28229 , n28230 , n28231 , n28232 , n28233 , n28234 , n28235 , n28236 , n28237 , n28238 , n28239 , n28240 , n28241 , n28242 , n28243 , n28244 , n28245 , n28246 , n28247 , n28248 , n28249 , n28250 , n28251 , n28252 , n28253 , n28254 , n28255 , n28256 , n28257 , n28258 , n28259 , n28260 , n28261 , n28262 , n28263 , n28264 , n28265 , n28266 , n28267 , n28268 , n28269 , n28270 , n28271 , n28272 , n28273 , n28274 , n28275 , n28276 , n28277 , n28278 , n28279 , n28280 , n28281 , n28282 , n28283 , n28284 , n28285 , n28286 , n28287 , n28288 , n28289 , n28290 , n28291 , n28292 , n28293 , n28294 , n28295 , n28296 , n28297 , n28298 , n28299 , n28300 , n28301 , n28302 , n28303 , n28304 , n28305 , n28306 , n28307 , n28308 , n28309 , n28310 , n28311 , n28312 , n28313 , n28314 , n28315 , n28316 , n28317 , n28318 , n28319 , n28320 , n28321 , n28322 , n28323 , n28324 , n28325 , n28326 , n28327 , n28328 , n28329 , n28330 , n28331 , n28332 , n28333 , n28334 , n28335 , n28336 , n28337 , n28338 , n28339 , n28340 , n28341 , n28342 , n28343 , n28344 , n28345 , n28346 , n28347 , n28348 , n28349 , n28350 , n28351 , n28352 , n28353 , n28354 , n28355 , n28356 , n28357 , n28358 , n28359 , n28360 , n28361 , n28362 , n28363 , n28364 , n28365 , n28366 , n28367 , n28368 , n28369 , n28370 , n28371 , n28372 , n28373 , n28374 , n28375 , n28376 , n28377 , n28378 , n28379 , n28380 , n28381 , n28382 , n28383 , n28384 , n28385 , n28386 , n28387 , n28388 , n28389 , n28390 , n28391 , n28392 , n28393 , n28394 , n28395 , n28396 , n28397 , n28398 , n28399 , n28400 , n28401 , n28402 , n28403 , n28404 , n28405 , n28406 , n28407 , n28408 , n28409 , n28410 , n28411 , n28412 , n28413 , n28414 , n28415 , n28416 , n28417 , n28418 , n28419 , n28420 , n28421 , n28422 , n28423 , n28424 , n28425 , n28426 , n28427 , n28428 , n28429 , n28430 , n28431 , n28432 , n28433 , n28434 , n28435 , n28436 , n28437 , n28438 , n28439 , n28440 , n28441 , n28442 , n28443 , n28444 , n28445 , n28446 , n28447 , n28448 , n28449 , n28450 , n28451 , n28452 , n28453 , n28454 , n28455 , n28456 , n28457 , n28458 , n28459 , n28460 , n28461 , n28462 , n28463 , n28464 , n28465 , n28466 , n28467 , n28468 , n28469 , n28470 , n28471 , n28472 , n28473 , n28474 , n28475 , n28476 , n28477 , n28478 , n28479 , n28480 , n28481 , n28482 , n28483 , n28484 , n28485 , n28486 , n28487 , n28488 , n28489 , n28490 , n28491 , n28492 , n28493 , n28494 , n28495 , n28496 , n28497 , n28498 , n28499 , n28500 , n28501 , n28502 , n28503 , n28504 , n28505 , n28506 , n28507 , n28508 , n28509 , n28510 , n28511 , n28512 , n28513 , n28514 , n28515 , n28516 , n28517 , n28518 , n28519 , n28520 , n28521 , n28522 , n28523 , n28524 , n28525 , n28526 , n28527 , n28528 , n28529 , n28530 , n28531 , n28532 , n28533 , n28534 , n28535 , n28536 , n28537 , n28538 , n28539 , n28540 , n28541 , n28542 , n28543 , n28544 , n28545 , n28546 , n28547 , n28548 , n28549 , n28550 , n28551 , n28552 , n28553 , n28554 , n28555 , n28556 , n28557 , n28558 , n28559 , n28560 , n28561 , n28562 , n28563 , n28564 , n28565 , n28566 , n28567 , n28568 , n28569 , n28570 , n28571 , n28572 , n28573 , n28574 , n28575 , n28576 , n28577 , n28578 , n28579 , n28580 , n28581 , n28582 , n28583 , n28584 , n28585 , n28586 , n28587 , n28588 , n28589 , n28590 , n28591 , n28592 , n28593 , n28594 , n28595 , n28596 , n28597 , n28598 , n28599 , n28600 , n28601 , n28602 , n28603 , n28604 , n28605 , n28606 , n28607 , n28608 , n28609 , n28610 , n28611 , n28612 , n28613 , n28614 , n28615 , n28616 , n28617 , n28618 , n28619 , n28620 , n28621 , n28622 , n28623 , n28624 , n28625 , n28626 , n28627 , n28628 , n28629 , n28630 , n28631 , n28632 , n28633 , n28634 , n28635 , n28636 , n28637 , n28638 , n28639 , n28640 , n28641 , n28642 , n28643 , n28644 , n28645 , n28646 , n28647 , n28648 , n28649 , n28650 , n28651 , n28652 , n28653 , n28654 , n28655 , n28656 , n28657 , n28658 , n28659 , n28660 , n28661 , n28662 , n28663 , n28664 , n28665 , n28666 , n28667 , n28668 , n28669 , n28670 , n28671 , n28672 , n28673 , n28674 , n28675 , n28676 , n28677 , n28678 , n28679 , n28680 , n28681 , n28682 , n28683 , n28684 , n28685 , n28686 , n28687 , n28688 , n28689 , n28690 , n28691 , n28692 , n28693 , n28694 , n28695 , n28696 , n28697 , n28698 , n28699 , n28700 , n28701 , n28702 , n28703 , n28704 , n28705 , n28706 , n28707 , n28708 , n28709 , n28710 , n28711 , n28712 , n28713 , n28714 , n28715 , n28716 , n28717 , n28718 , n28719 , n28720 , n28721 , n28722 , n28723 , n28724 , n28725 , n28726 , n28727 , n28728 , n28729 , n28730 , n28731 , n28732 , n28733 , n28734 , n28735 , n28736 , n28737 , n28738 , n28739 , n28740 , n28741 , n28742 , n28743 , n28744 , n28745 , n28746 , n28747 , n28748 , n28749 , n28750 , n28751 , n28752 , n28753 , n28754 , n28755 , n28756 , n28757 , n28758 , n28759 , n28760 , n28761 , n28762 , n28763 , n28764 , n28765 , n28766 , n28767 , n28768 , n28769 , n28770 , n28771 , n28772 , n28773 , n28774 , n28775 , n28776 , n28777 , n28778 , n28779 , n28780 , n28781 , n28782 , n28783 , n28784 , n28785 , n28786 , n28787 , n28788 , n28789 , n28790 , n28791 , n28792 , n28793 , n28794 , n28795 , n28796 , n28797 , n28798 , n28799 , n28800 , n28801 , n28802 , n28803 , n28804 , n28805 , n28806 , n28807 , n28808 , n28809 , n28810 , n28811 , n28812 , n28813 , n28814 , n28815 , n28816 , n28817 , n28818 , n28819 , n28820 , n28821 , n28822 , n28823 , n28824 , n28825 , n28826 , n28827 , n28828 , n28829 , n28830 , n28831 , n28832 , n28833 , n28834 , n28835 , n28836 , n28837 , n28838 , n28839 , n28840 , n28841 , n28842 , n28843 , n28844 , n28845 , n28846 , n28847 , n28848 , n28849 , n28850 , n28851 , n28852 , n28853 , n28854 , n28855 , n28856 , n28857 , n28858 , n28859 , n28860 , n28861 , n28862 , n28863 , n28864 , n28865 , n28866 , n28867 , n28868 , n28869 , n28870 , n28871 , n28872 , n28873 , n28874 , n28875 , n28876 , n28877 , n28878 , n28879 , n28880 , n28881 , n28882 , n28883 , n28884 , n28885 , n28886 , n28887 , n28888 , n28889 , n28890 , n28891 , n28892 , n28893 , n28894 , n28895 , n28896 , n28897 , n28898 , n28899 , n28900 , n28901 , n28902 , n28903 , n28904 , n28905 , n28906 , n28907 , n28908 , n28909 , n28910 , n28911 , n28912 , n28913 , n28914 , n28915 , n28916 , n28917 , n28918 , n28919 , n28920 , n28921 , n28922 , n28923 , n28924 , n28925 , n28926 , n28927 , n28928 , n28929 , n28930 , n28931 , n28932 , n28933 , n28934 , n28935 , n28936 , n28937 , n28938 , n28939 , n28940 , n28941 , n28942 , n28943 , n28944 , n28945 , n28946 , n28947 , n28948 , n28949 , n28950 , n28951 , n28952 , n28953 , n28954 , n28955 , n28956 , n28957 , n28958 , n28959 , n28960 , n28961 , n28962 , n28963 , n28964 , n28965 , n28966 , n28967 , n28968 , n28969 , n28970 , n28971 , n28972 , n28973 , n28974 , n28975 , n28976 , n28977 , n28978 , n28979 , n28980 , n28981 , n28982 , n28983 , n28984 , n28985 , n28986 , n28987 , n28988 , n28989 , n28990 , n28991 , n28992 , n28993 , n28994 , n28995 , n28996 , n28997 , n28998 , n28999 , n29000 , n29001 , n29002 , n29003 , n29004 , n29005 , n29006 , n29007 , n29008 , n29009 , n29010 , n29011 , n29012 , n29013 , n29014 , n29015 , n29016 , n29017 , n29018 , n29019 , n29020 , n29021 , n29022 , n29023 , n29024 , n29025 , n29026 , n29027 , n29028 , n29029 , n29030 , n29031 , n29032 , n29033 , n29034 , n29035 , n29036 , n29037 , n29038 , n29039 , n29040 , n29041 , n29042 , n29043 , n29044 , n29045 , n29046 , n29047 , n29048 , n29049 , n29050 , n29051 , n29052 , n29053 , n29054 , n29055 , n29056 , n29057 , n29058 , n29059 , n29060 , n29061 , n29062 , n29063 , n29064 , n29065 , n29066 , n29067 , n29068 , n29069 , n29070 , n29071 , n29072 , n29073 , n29074 , n29075 , n29076 , n29077 , n29078 , n29079 , n29080 , n29081 , n29082 , n29083 , n29084 , n29085 , n29086 , n29087 , n29088 , n29089 , n29090 , n29091 , n29092 , n29093 , n29094 , n29095 , n29096 , n29097 , n29098 , n29099 , n29100 , n29101 , n29102 , n29103 , n29104 , n29105 , n29106 , n29107 , n29108 , n29109 , n29110 , n29111 , n29112 , n29113 , n29114 , n29115 , n29116 , n29117 , n29118 , n29119 , n29120 , n29121 , n29122 , n29123 , n29124 , n29125 , n29126 , n29127 , n29128 , n29129 , n29130 , n29131 , n29132 , n29133 , n29134 , n29135 , n29136 , n29137 , n29138 , n29139 , n29140 , n29141 , n29142 , n29143 , n29144 , n29145 , n29146 , n29147 , n29148 , n29149 , n29150 , n29151 , n29152 , n29153 , n29154 , n29155 , n29156 , n29157 , n29158 , n29159 , n29160 , n29161 , n29162 , n29163 , n29164 , n29165 , n29166 , n29167 , n29168 , n29169 , n29170 , n29171 , n29172 , n29173 , n29174 , n29175 , n29176 , n29177 , n29178 , n29179 , n29180 , n29181 , n29182 , n29183 , n29184 , n29185 , n29186 , n29187 , n29188 , n29189 , n29190 , n29191 , n29192 , n29193 , n29194 , n29195 , n29196 , n29197 , n29198 , n29199 , n29200 , n29201 , n29202 , n29203 , n29204 , n29205 , n29206 , n29207 , n29208 , n29209 , n29210 , n29211 , n29212 , n29213 , n29214 , n29215 , n29216 , n29217 , n29218 , n29219 , n29220 , n29221 , n29222 , n29223 , n29224 , n29225 , n29226 , n29227 , n29228 , n29229 , n29230 , n29231 , n29232 , n29233 , n29234 , n29235 , n29236 , n29237 , n29238 , n29239 , n29240 , n29241 , n29242 , n29243 , n29244 , n29245 , n29246 , n29247 , n29248 , n29249 , n29250 , n29251 , n29252 , n29253 , n29254 , n29255 , n29256 , n29257 , n29258 , n29259 , n29260 , n29261 , n29262 , n29263 , n29264 , n29265 , n29266 , n29267 , n29268 , n29269 , n29270 , n29271 , n29272 , n29273 , n29274 , n29275 , n29276 , n29277 , n29278 , n29279 , n29280 , n29281 , n29282 , n29283 , n29284 , n29285 , n29286 , n29287 , n29288 , n29289 , n29290 , n29291 , n29292 , n29293 , n29294 , n29295 , n29296 , n29297 , n29298 , n29299 , n29300 , n29301 , n29302 , n29303 , n29304 , n29305 , n29306 , n29307 , n29308 , n29309 , n29310 , n29311 , n29312 , n29313 , n29314 , n29315 , n29316 , n29317 , n29318 , n29319 , n29320 , n29321 , n29322 , n29323 , n29324 , n29325 , n29326 , n29327 , n29328 , n29329 , n29330 , n29331 , n29332 , n29333 , n29334 , n29335 , n29336 , n29337 , n29338 , n29339 , n29340 , n29341 , n29342 , n29343 , n29344 , n29345 , n29346 , n29347 , n29348 , n29349 , n29350 , n29351 , n29352 , n29353 , n29354 , n29355 , n29356 , n29357 , n29358 , n29359 , n29360 , n29361 , n29362 , n29363 , n29364 , n29365 , n29366 , n29367 , n29368 , n29369 , n29370 , n29371 , n29372 , n29373 , n29374 , n29375 , n29376 , n29377 , n29378 , n29379 , n29380 , n29381 , n29382 , n29383 , n29384 , n29385 , n29386 , n29387 , n29388 , n29389 , n29390 , n29391 , n29392 , n29393 , n29394 , n29395 , n29396 , n29397 , n29398 , n29399 , n29400 , n29401 , n29402 , n29403 , n29404 , n29405 , n29406 , n29407 , n29408 , n29409 , n29410 , n29411 , n29412 , n29413 , n29414 , n29415 , n29416 , n29417 , n29418 , n29419 , n29420 , n29421 , n29422 , n29423 , n29424 , n29425 , n29426 , n29427 , n29428 , n29429 , n29430 , n29431 , n29432 , n29433 , n29434 , n29435 , n29436 , n29437 , n29438 , n29439 , n29440 , n29441 , n29442 , n29443 , n29444 , n29445 , n29446 , n29447 , n29448 , n29449 , n29450 , n29451 , n29452 , n29453 , n29454 , n29455 , n29456 , n29457 , n29458 , n29459 , n29460 , n29461 , n29462 , n29463 , n29464 , n29465 , n29466 , n29467 , n29468 , n29469 , n29470 , n29471 , n29472 , n29473 , n29474 , n29475 , n29476 , n29477 , n29478 , n29479 , n29480 , n29481 , n29482 , n29483 , n29484 , n29485 , n29486 , n29487 , n29488 , n29489 , n29490 , n29491 , n29492 , n29493 , n29494 , n29495 , n29496 , n29497 , n29498 , n29499 , n29500 , n29501 , n29502 , n29503 , n29504 , n29505 , n29506 , n29507 , n29508 , n29509 , n29510 , n29511 , n29512 , n29513 , n29514 , n29515 , n29516 , n29517 , n29518 , n29519 , n29520 , n29521 , n29522 , n29523 , n29524 , n29525 , n29526 , n29527 , n29528 , n29529 , n29530 , n29531 , n29532 , n29533 , n29534 , n29535 , n29536 , n29537 , n29538 , n29539 , n29540 , n29541 , n29542 , n29543 , n29544 , n29545 , n29546 , n29547 , n29548 , n29549 , n29550 , n29551 , n29552 , n29553 , n29554 , n29555 , n29556 , n29557 , n29558 , n29559 , n29560 , n29561 , n29562 , n29563 , n29564 , n29565 , n29566 , n29567 , n29568 , n29569 , n29570 , n29571 , n29572 , n29573 , n29574 , n29575 , n29576 , n29577 , n29578 , n29579 , n29580 , n29581 , n29582 , n29583 , n29584 , n29585 , n29586 , n29587 , n29588 , n29589 , n29590 , n29591 , n29592 , n29593 , n29594 , n29595 , n29596 , n29597 , n29598 , n29599 , n29600 , n29601 , n29602 , n29603 , n29604 , n29605 , n29606 , n29607 , n29608 , n29609 , n29610 , n29611 , n29612 , n29613 , n29614 , n29615 , n29616 , n29617 , n29618 , n29619 , n29620 , n29621 , n29622 , n29623 , n29624 , n29625 , n29626 , n29627 , n29628 , n29629 , n29630 , n29631 , n29632 , n29633 , n29634 , n29635 , n29636 , n29637 , n29638 , n29639 , n29640 , n29641 , n29642 , n29643 , n29644 , n29645 , n29646 , n29647 , n29648 , n29649 , n29650 , n29651 , n29652 , n29653 , n29654 , n29655 , n29656 , n29657 , n29658 , n29659 , n29660 , n29661 , n29662 , n29663 , n29664 , n29665 , n29666 , n29667 , n29668 , n29669 , n29670 , n29671 , n29672 , n29673 , n29674 , n29675 , n29676 , n29677 , n29678 , n29679 , n29680 , n29681 , n29682 , n29683 , n29684 , n29685 , n29686 , n29687 , n29688 , n29689 , n29690 , n29691 , n29692 , n29693 , n29694 , n29695 , n29696 , n29697 , n29698 , n29699 , n29700 , n29701 , n29702 , n29703 , n29704 , n29705 , n29706 , n29707 , n29708 , n29709 , n29710 , n29711 , n29712 , n29713 , n29714 , n29715 , n29716 , n29717 , n29718 , n29719 , n29720 , n29721 , n29722 , n29723 , n29724 , n29725 , n29726 , n29727 , n29728 , n29729 , n29730 , n29731 , n29732 , n29733 , n29734 , n29735 , n29736 , n29737 , n29738 , n29739 , n29740 , n29741 , n29742 , n29743 , n29744 , n29745 , n29746 , n29747 , n29748 , n29749 , n29750 , n29751 , n29752 , n29753 , n29754 , n29755 , n29756 , n29757 , n29758 , n29759 , n29760 , n29761 , n29762 , n29763 , n29764 , n29765 , n29766 , n29767 , n29768 , n29769 , n29770 , n29771 , n29772 , n29773 , n29774 , n29775 , n29776 , n29777 , n29778 , n29779 , n29780 , n29781 , n29782 , n29783 , n29784 , n29785 , n29786 , n29787 , n29788 , n29789 , n29790 , n29791 , n29792 , n29793 , n29794 , n29795 , n29796 , n29797 , n29798 , n29799 , n29800 , n29801 , n29802 , n29803 , n29804 , n29805 , n29806 , n29807 , n29808 , n29809 , n29810 , n29811 , n29812 , n29813 , n29814 , n29815 , n29816 , n29817 , n29818 , n29819 , n29820 , n29821 , n29822 , n29823 , n29824 , n29825 , n29826 , n29827 , n29828 , n29829 , n29830 , n29831 , n29832 , n29833 , n29834 , n29835 , n29836 , n29837 , n29838 , n29839 , n29840 , n29841 , n29842 , n29843 , n29844 , n29845 , n29846 , n29847 , n29848 , n29849 , n29850 , n29851 , n29852 , n29853 , n29854 , n29855 , n29856 , n29857 , n29858 , n29859 , n29860 , n29861 , n29862 , n29863 , n29864 , n29865 , n29866 , n29867 , n29868 , n29869 , n29870 , n29871 , n29872 , n29873 , n29874 , n29875 , n29876 , n29877 , n29878 , n29879 , n29880 , n29881 , n29882 , n29883 , n29884 , n29885 , n29886 , n29887 , n29888 , n29889 , n29890 , n29891 , n29892 , n29893 , n29894 , n29895 , n29896 , n29897 , n29898 , n29899 , n29900 , n29901 , n29902 , n29903 , n29904 , n29905 , n29906 , n29907 , n29908 , n29909 , n29910 , n29911 , n29912 , n29913 , n29914 , n29915 , n29916 , n29917 , n29918 , n29919 , n29920 , n29921 , n29922 , n29923 , n29924 , n29925 , n29926 , n29927 , n29928 , n29929 , n29930 , n29931 , n29932 , n29933 , n29934 , n29935 , n29936 , n29937 , n29938 , n29939 , n29940 , n29941 , n29942 , n29943 , n29944 , n29945 , n29946 , n29947 , n29948 , n29949 , n29950 , n29951 , n29952 , n29953 , n29954 , n29955 , n29956 , n29957 , n29958 , n29959 , n29960 , n29961 , n29962 , n29963 , n29964 , n29965 , n29966 , n29967 , n29968 , n29969 , n29970 , n29971 , n29972 , n29973 , n29974 , n29975 , n29976 , n29977 , n29978 , n29979 , n29980 , n29981 , n29982 , n29983 , n29984 , n29985 , n29986 , n29987 , n29988 , n29989 , n29990 , n29991 , n29992 , n29993 , n29994 , n29995 , n29996 , n29997 , n29998 , n29999 , n30000 , n30001 , n30002 , n30003 , n30004 , n30005 , n30006 , n30007 , n30008 , n30009 , n30010 , n30011 , n30012 , n30013 , n30014 , n30015 , n30016 , n30017 , n30018 , n30019 , n30020 , n30021 , n30022 , n30023 , n30024 , n30025 , n30026 , n30027 , n30028 , n30029 , n30030 , n30031 , n30032 , n30033 , n30034 , n30035 , n30036 , n30037 , n30038 , n30039 , n30040 , n30041 , n30042 , n30043 , n30044 , n30045 , n30046 , n30047 , n30048 , n30049 , n30050 , n30051 , n30052 , n30053 , n30054 , n30055 , n30056 , n30057 , n30058 , n30059 , n30060 , n30061 , n30062 , n30063 , n30064 , n30065 , n30066 , n30067 , n30068 , n30069 , n30070 , n30071 , n30072 , n30073 , n30074 , n30075 , n30076 , n30077 , n30078 , n30079 , n30080 , n30081 , n30082 , n30083 , n30084 , n30085 , n30086 , n30087 , n30088 , n30089 , n30090 , n30091 , n30092 , n30093 , n30094 , n30095 , n30096 , n30097 , n30098 , n30099 , n30100 , n30101 , n30102 , n30103 , n30104 , n30105 , n30106 , n30107 , n30108 , n30109 , n30110 , n30111 , n30112 , n30113 , n30114 , n30115 , n30116 , n30117 , n30118 , n30119 , n30120 , n30121 , n30122 , n30123 , n30124 , n30125 , n30126 , n30127 , n30128 , n30129 , n30130 , n30131 , n30132 , n30133 , n30134 , n30135 , n30136 , n30137 , n30138 , n30139 , n30140 , n30141 , n30142 , n30143 , n30144 , n30145 , n30146 , n30147 , n30148 , n30149 , n30150 , n30151 , n30152 , n30153 , n30154 , n30155 , n30156 , n30157 , n30158 , n30159 , n30160 , n30161 , n30162 , n30163 , n30164 , n30165 , n30166 , n30167 , n30168 , n30169 , n30170 , n30171 , n30172 , n30173 , n30174 , n30175 , n30176 , n30177 , n30178 , n30179 , n30180 , n30181 , n30182 , n30183 , n30184 , n30185 , n30186 , n30187 , n30188 , n30189 , n30190 , n30191 , n30192 , n30193 , n30194 , n30195 , n30196 , n30197 , n30198 , n30199 , n30200 , n30201 , n30202 , n30203 , n30204 , n30205 , n30206 , n30207 , n30208 , n30209 , n30210 , n30211 , n30212 , n30213 , n30214 , n30215 , n30216 , n30217 , n30218 , n30219 , n30220 , n30221 , n30222 , n30223 , n30224 , n30225 , n30226 , n30227 , n30228 , n30229 , n30230 , n30231 , n30232 , n30233 , n30234 , n30235 , n30236 , n30237 , n30238 , n30239 , n30240 , n30241 , n30242 , n30243 , n30244 , n30245 , n30246 , n30247 , n30248 , n30249 , n30250 , n30251 , n30252 , n30253 , n30254 , n30255 , n30256 , n30257 , n30258 , n30259 , n30260 , n30261 , n30262 , n30263 , n30264 , n30265 , n30266 , n30267 , n30268 , n30269 , n30270 , n30271 , n30272 , n30273 , n30274 , n30275 , n30276 , n30277 , n30278 , n30279 , n30280 , n30281 , n30282 , n30283 , n30284 , n30285 , n30286 , n30287 , n30288 , n30289 , n30290 , n30291 , n30292 , n30293 , n30294 , n30295 , n30296 , n30297 , n30298 , n30299 , n30300 , n30301 , n30302 , n30303 , n30304 , n30305 , n30306 , n30307 , n30308 , n30309 , n30310 , n30311 , n30312 , n30313 , n30314 , n30315 , n30316 , n30317 , n30318 , n30319 , n30320 , n30321 , n30322 , n30323 , n30324 , n30325 , n30326 , n30327 , n30328 , n30329 , n30330 , n30331 , n30332 , n30333 , n30334 , n30335 , n30336 , n30337 , n30338 , n30339 , n30340 , n30341 , n30342 , n30343 , n30344 , n30345 , n30346 , n30347 , n30348 , n30349 , n30350 , n30351 , n30352 , n30353 , n30354 , n30355 , n30356 , n30357 , n30358 , n30359 , n30360 , n30361 , n30362 , n30363 , n30364 , n30365 , n30366 , n30367 , n30368 , n30369 , n30370 , n30371 , n30372 , n30373 , n30374 , n30375 , n30376 , n30377 , n30378 , n30379 , n30380 , n30381 , n30382 , n30383 , n30384 , n30385 , n30386 , n30387 , n30388 , n30389 , n30390 , n30391 , n30392 , n30393 , n30394 , n30395 , n30396 , n30397 , n30398 , n30399 , n30400 , n30401 , n30402 , n30403 , n30404 , n30405 , n30406 , n30407 , n30408 , n30409 , n30410 , n30411 , n30412 , n30413 , n30414 , n30415 , n30416 , n30417 , n30418 , n30419 , n30420 , n30421 , n30422 , n30423 , n30424 , n30425 , n30426 , n30427 , n30428 , n30429 , n30430 , n30431 , n30432 , n30433 , n30434 , n30435 , n30436 , n30437 , n30438 , n30439 , n30440 , n30441 , n30442 , n30443 , n30444 , n30445 , n30446 , n30447 , n30448 , n30449 , n30450 , n30451 , n30452 , n30453 , n30454 , n30455 , n30456 , n30457 , n30458 , n30459 , n30460 , n30461 , n30462 , n30463 , n30464 , n30465 , n30466 , n30467 , n30468 , n30469 , n30470 , n30471 , n30472 , n30473 , n30474 , n30475 , n30476 , n30477 , n30478 , n30479 , n30480 , n30481 , n30482 , n30483 , n30484 , n30485 , n30486 , n30487 , n30488 , n30489 , n30490 , n30491 , n30492 , n30493 , n30494 , n30495 , n30496 , n30497 , n30498 , n30499 , n30500 , n30501 , n30502 , n30503 , n30504 , n30505 , n30506 , n30507 , n30508 , n30509 , n30510 , n30511 , n30512 , n30513 , n30514 , n30515 , n30516 , n30517 , n30518 , n30519 , n30520 , n30521 , n30522 , n30523 , n30524 , n30525 , n30526 , n30527 , n30528 , n30529 , n30530 , n30531 , n30532 , n30533 , n30534 , n30535 , n30536 , n30537 , n30538 , n30539 , n30540 , n30541 , n30542 , n30543 , n30544 , n30545 , n30546 , n30547 , n30548 , n30549 , n30550 , n30551 , n30552 , n30553 , n30554 , n30555 , n30556 , n30557 , n30558 , n30559 , n30560 , n30561 , n30562 , n30563 , n30564 , n30565 , n30566 , n30567 , n30568 , n30569 , n30570 , n30571 , n30572 , n30573 , n30574 , n30575 , n30576 , n30577 , n30578 , n30579 , n30580 , n30581 , n30582 , n30583 , n30584 , n30585 , n30586 , n30587 , n30588 , n30589 , n30590 , n30591 , n30592 , n30593 , n30594 , n30595 , n30596 , n30597 , n30598 , n30599 , n30600 , n30601 , n30602 , n30603 , n30604 , n30605 , n30606 , n30607 , n30608 , n30609 , n30610 , n30611 , n30612 , n30613 , n30614 , n30615 , n30616 , n30617 , n30618 , n30619 , n30620 , n30621 , n30622 , n30623 , n30624 , n30625 , n30626 , n30627 , n30628 , n30629 , n30630 , n30631 , n30632 , n30633 , n30634 , n30635 , n30636 , n30637 , n30638 , n30639 , n30640 , n30641 , n30642 , n30643 , n30644 , n30645 , n30646 , n30647 , n30648 , n30649 , n30650 , n30651 , n30652 , n30653 , n30654 , n30655 , n30656 , n30657 , n30658 , n30659 , n30660 , n30661 , n30662 , n30663 , n30664 , n30665 , n30666 , n30667 , n30668 , n30669 , n30670 , n30671 , n30672 , n30673 , n30674 , n30675 , n30676 , n30677 , n30678 , n30679 , n30680 , n30681 , n30682 , n30683 , n30684 , n30685 , n30686 , n30687 , n30688 , n30689 , n30690 , n30691 , n30692 , n30693 , n30694 , n30695 , n30696 , n30697 , n30698 , n30699 , n30700 , n30701 , n30702 , n30703 , n30704 , n30705 , n30706 , n30707 , n30708 , n30709 , n30710 , n30711 , n30712 , n30713 , n30714 , n30715 , n30716 , n30717 , n30718 , n30719 , n30720 , n30721 , n30722 , n30723 , n30724 , n30725 , n30726 , n30727 , n30728 , n30729 , n30730 , n30731 , n30732 , n30733 , n30734 , n30735 , n30736 , n30737 , n30738 , n30739 , n30740 , n30741 , n30742 , n30743 , n30744 , n30745 , n30746 , n30747 , n30748 , n30749 , n30750 , n30751 , n30752 , n30753 , n30754 , n30755 , n30756 , n30757 , n30758 , n30759 , n30760 , n30761 , n30762 , n30763 , n30764 , n30765 , n30766 , n30767 , n30768 , n30769 , n30770 , n30771 , n30772 , n30773 , n30774 , n30775 , n30776 , n30777 , n30778 , n30779 , n30780 , n30781 , n30782 , n30783 , n30784 , n30785 , n30786 , n30787 , n30788 , n30789 , n30790 , n30791 , n30792 , n30793 , n30794 , n30795 , n30796 , n30797 , n30798 , n30799 , n30800 , n30801 , n30802 , n30803 , n30804 , n30805 , n30806 , n30807 , n30808 , n30809 , n30810 , n30811 , n30812 , n30813 , n30814 , n30815 , n30816 , n30817 , n30818 , n30819 , n30820 , n30821 , n30822 , n30823 , n30824 , n30825 , n30826 , n30827 , n30828 , n30829 , n30830 , n30831 , n30832 , n30833 , n30834 , n30835 , n30836 , n30837 , n30838 , n30839 , n30840 , n30841 , n30842 , n30843 , n30844 , n30845 , n30846 , n30847 , n30848 , n30849 , n30850 , n30851 , n30852 , n30853 , n30854 , n30855 , n30856 , n30857 , n30858 , n30859 , n30860 , n30861 , n30862 , n30863 , n30864 , n30865 , n30866 , n30867 , n30868 , n30869 , n30870 , n30871 , n30872 , n30873 , n30874 , n30875 , n30876 , n30877 , n30878 , n30879 , n30880 , n30881 , n30882 , n30883 , n30884 , n30885 , n30886 , n30887 , n30888 , n30889 , n30890 , n30891 , n30892 , n30893 , n30894 , n30895 , n30896 , n30897 , n30898 , n30899 , n30900 , n30901 , n30902 , n30903 , n30904 , n30905 , n30906 , n30907 , n30908 , n30909 , n30910 , n30911 , n30912 , n30913 , n30914 , n30915 , n30916 , n30917 , n30918 , n30919 , n30920 , n30921 , n30922 , n30923 , n30924 , n30925 , n30926 , n30927 , n30928 , n30929 , n30930 , n30931 , n30932 , n30933 , n30934 , n30935 , n30936 , n30937 , n30938 , n30939 , n30940 , n30941 , n30942 , n30943 , n30944 , n30945 , n30946 , n30947 , n30948 , n30949 , n30950 , n30951 , n30952 , n30953 , n30954 , n30955 , n30956 , n30957 , n30958 , n30959 , n30960 , n30961 , n30962 , n30963 , n30964 , n30965 , n30966 , n30967 , n30968 , n30969 , n30970 , n30971 , n30972 , n30973 , n30974 , n30975 , n30976 , n30977 , n30978 , n30979 , n30980 , n30981 , n30982 , n30983 , n30984 , n30985 , n30986 , n30987 , n30988 , n30989 , n30990 , n30991 , n30992 , n30993 , n30994 , n30995 , n30996 , n30997 , n30998 , n30999 , n31000 , n31001 , n31002 , n31003 , n31004 , n31005 , n31006 , n31007 , n31008 , n31009 , n31010 , n31011 , n31012 , n31013 , n31014 , n31015 , n31016 , n31017 , n31018 , n31019 , n31020 , n31021 , n31022 , n31023 , n31024 , n31025 , n31026 , n31027 , n31028 , n31029 , n31030 , n31031 , n31032 , n31033 , n31034 , n31035 , n31036 , n31037 , n31038 , n31039 , n31040 , n31041 , n31042 , n31043 , n31044 , n31045 , n31046 , n31047 , n31048 , n31049 , n31050 , n31051 , n31052 , n31053 , n31054 , n31055 , n31056 , n31057 , n31058 , n31059 , n31060 , n31061 , n31062 , n31063 , n31064 , n31065 , n31066 , n31067 , n31068 , n31069 , n31070 , n31071 , n31072 , n31073 , n31074 , n31075 , n31076 , n31077 , n31078 , n31079 , n31080 , n31081 , n31082 , n31083 , n31084 , n31085 , n31086 , n31087 , n31088 , n31089 , n31090 , n31091 , n31092 , n31093 , n31094 , n31095 , n31096 , n31097 , n31098 , n31099 , n31100 , n31101 , n31102 , n31103 , n31104 , n31105 , n31106 , n31107 , n31108 , n31109 , n31110 , n31111 , n31112 , n31113 , n31114 , n31115 , n31116 , n31117 , n31118 , n31119 , n31120 , n31121 , n31122 , n31123 , n31124 , n31125 , n31126 , n31127 , n31128 , n31129 , n31130 , n31131 , n31132 , n31133 , n31134 , n31135 , n31136 , n31137 , n31138 , n31139 , n31140 , n31141 , n31142 , n31143 , n31144 , n31145 , n31146 , n31147 , n31148 , n31149 , n31150 , n31151 , n31152 , n31153 , n31154 , n31155 , n31156 , n31157 , n31158 , n31159 , n31160 , n31161 , n31162 , n31163 , n31164 , n31165 , n31166 , n31167 , n31168 , n31169 , n31170 , n31171 , n31172 , n31173 , n31174 , n31175 , n31176 , n31177 , n31178 , n31179 , n31180 , n31181 , n31182 , n31183 , n31184 , n31185 , n31186 , n31187 , n31188 , n31189 , n31190 , n31191 , n31192 , n31193 , n31194 , n31195 , n31196 , n31197 , n31198 , n31199 , n31200 , n31201 , n31202 , n31203 , n31204 , n31205 , n31206 , n31207 , n31208 , n31209 , n31210 , n31211 , n31212 , n31213 , n31214 , n31215 , n31216 , n31217 , n31218 , n31219 , n31220 , n31221 , n31222 , n31223 , n31224 , n31225 , n31226 , n31227 , n31228 , n31229 , n31230 , n31231 , n31232 , n31233 , n31234 , n31235 , n31236 , n31237 , n31238 , n31239 , n31240 , n31241 , n31242 , n31243 , n31244 , n31245 , n31246 , n31247 , n31248 , n31249 , n31250 , n31251 , n31252 , n31253 , n31254 , n31255 , n31256 , n31257 , n31258 , n31259 , n31260 , n31261 , n31262 , n31263 , n31264 , n31265 , n31266 , n31267 , n31268 , n31269 , n31270 , n31271 , n31272 , n31273 , n31274 , n31275 , n31276 , n31277 , n31278 , n31279 , n31280 , n31281 , n31282 , n31283 , n31284 , n31285 , n31286 , n31287 , n31288 , n31289 , n31290 , n31291 , n31292 , n31293 , n31294 , n31295 , n31296 , n31297 , n31298 , n31299 , n31300 , n31301 , n31302 , n31303 , n31304 , n31305 , n31306 , n31307 , n31308 , n31309 , n31310 , n31311 , n31312 , n31313 , n31314 , n31315 , n31316 , n31317 , n31318 , n31319 , n31320 , n31321 , n31322 , n31323 , n31324 , n31325 , n31326 , n31327 , n31328 , n31329 , n31330 , n31331 , n31332 , n31333 , n31334 , n31335 , n31336 , n31337 , n31338 , n31339 , n31340 , n31341 , n31342 , n31343 , n31344 , n31345 , n31346 , n31347 , n31348 , n31349 , n31350 , n31351 , n31352 , n31353 , n31354 , n31355 , n31356 , n31357 , n31358 , n31359 , n31360 , n31361 , n31362 , n31363 , n31364 , n31365 , n31366 , n31367 , n31368 , n31369 , n31370 , n31371 , n31372 , n31373 , n31374 , n31375 , n31376 , n31377 , n31378 , n31379 , n31380 , n31381 , n31382 , n31383 , n31384 , n31385 , n31386 , n31387 , n31388 , n31389 , n31390 , n31391 , n31392 , n31393 , n31394 , n31395 , n31396 , n31397 , n31398 , n31399 , n31400 , n31401 , n31402 , n31403 , n31404 , n31405 , n31406 , n31407 , n31408 , n31409 , n31410 , n31411 , n31412 , n31413 , n31414 , n31415 , n31416 , n31417 , n31418 , n31419 , n31420 , n31421 , n31422 , n31423 , n31424 , n31425 , n31426 , n31427 , n31428 , n31429 , n31430 , n31431 , n31432 , n31433 , n31434 , n31435 , n31436 , n31437 , n31438 , n31439 , n31440 , n31441 , n31442 , n31443 , n31444 , n31445 , n31446 , n31447 , n31448 , n31449 , n31450 , n31451 , n31452 , n31453 , n31454 , n31455 , n31456 , n31457 , n31458 , n31459 , n31460 , n31461 , n31462 , n31463 , n31464 , n31465 , n31466 , n31467 , n31468 , n31469 , n31470 , n31471 , n31472 , n31473 ;
  assign n129 = ( ~x56 & x108 ) | ( ~x56 & x119 ) | ( x108 & x119 ) ;
  assign n130 = x114 ^ x102 ^ x26 ;
  assign n131 = x62 ^ x42 ^ x23 ;
  assign n132 = x57 & x112 ;
  assign n133 = n132 ^ x70 ^ 1'b0 ;
  assign n134 = n129 ^ x97 ^ x87 ;
  assign n135 = x41 & x55 ;
  assign n136 = ~x44 & n135 ;
  assign n137 = ( x5 & x45 ) | ( x5 & n136 ) | ( x45 & n136 ) ;
  assign n138 = x70 ^ x22 ^ x3 ;
  assign n140 = x26 ^ x2 ^ 1'b0 ;
  assign n141 = x7 & n140 ;
  assign n139 = x39 & x82 ;
  assign n142 = n141 ^ n139 ^ 1'b0 ;
  assign n143 = ( x36 & x63 ) | ( x36 & n142 ) | ( x63 & n142 ) ;
  assign n144 = x115 ^ x18 ^ 1'b0 ;
  assign n145 = x107 & n144 ;
  assign n146 = n145 ^ x106 ^ x78 ;
  assign n147 = ( x20 & x71 ) | ( x20 & ~x112 ) | ( x71 & ~x112 ) ;
  assign n148 = n147 ^ x70 ^ x34 ;
  assign n149 = n148 ^ x27 ^ x21 ;
  assign n150 = n149 ^ x63 ^ x58 ;
  assign n151 = x127 ^ x69 ^ 1'b0 ;
  assign n154 = x53 ^ x7 ^ 1'b0 ;
  assign n155 = x16 & n154 ;
  assign n156 = n155 ^ n142 ^ x42 ;
  assign n152 = x65 & ~n148 ;
  assign n153 = ~x112 & n152 ;
  assign n157 = n156 ^ n153 ^ 1'b0 ;
  assign n158 = ( x13 & ~x43 ) | ( x13 & x92 ) | ( ~x43 & x92 ) ;
  assign n159 = n158 ^ x87 ^ x9 ;
  assign n160 = n131 | n159 ;
  assign n163 = x117 ^ x111 ^ x69 ;
  assign n161 = ( ~x53 & x59 ) | ( ~x53 & x81 ) | ( x59 & x81 ) ;
  assign n162 = ~x0 & n161 ;
  assign n164 = n163 ^ n162 ^ 1'b0 ;
  assign n167 = ( x49 & x52 ) | ( x49 & ~x92 ) | ( x52 & ~x92 ) ;
  assign n165 = x118 ^ x85 ^ x40 ;
  assign n166 = n165 ^ x53 ^ x25 ;
  assign n168 = n167 ^ n166 ^ x53 ;
  assign n169 = ( ~x65 & x66 ) | ( ~x65 & n168 ) | ( x66 & n168 ) ;
  assign n170 = x56 & n160 ;
  assign n171 = x53 ^ x39 ^ x33 ;
  assign n173 = x35 & ~n171 ;
  assign n174 = ~x32 & n173 ;
  assign n172 = ( x1 & ~n133 ) | ( x1 & n171 ) | ( ~n133 & n171 ) ;
  assign n175 = n174 ^ n172 ^ 1'b0 ;
  assign n176 = x30 & ~n175 ;
  assign n177 = x101 ^ x17 ^ x4 ;
  assign n178 = n177 ^ n141 ^ x8 ;
  assign n179 = ( x59 & ~x90 ) | ( x59 & n169 ) | ( ~x90 & n169 ) ;
  assign n180 = x126 ^ x106 ^ x70 ;
  assign n181 = n180 ^ x124 ^ x32 ;
  assign n182 = x27 & x73 ;
  assign n183 = ( ~x18 & x32 ) | ( ~x18 & x125 ) | ( x32 & x125 ) ;
  assign n184 = ( x3 & ~x66 ) | ( x3 & n183 ) | ( ~x66 & n183 ) ;
  assign n185 = x117 ^ x37 ^ x30 ;
  assign n186 = n185 ^ n165 ^ x9 ;
  assign n187 = x78 ^ x27 ^ 1'b0 ;
  assign n188 = ~n186 & n187 ;
  assign n189 = n188 ^ x86 ^ 1'b0 ;
  assign n190 = ( ~n182 & n184 ) | ( ~n182 & n189 ) | ( n184 & n189 ) ;
  assign n191 = x63 & x73 ;
  assign n192 = n191 ^ x118 ^ 1'b0 ;
  assign n193 = n192 ^ n129 ^ 1'b0 ;
  assign n194 = x30 & ~n193 ;
  assign n195 = ( x46 & n145 ) | ( x46 & n170 ) | ( n145 & n170 ) ;
  assign n198 = ( x64 & ~x100 ) | ( x64 & n147 ) | ( ~x100 & n147 ) ;
  assign n196 = x35 & x122 ;
  assign n197 = ~n155 & n196 ;
  assign n199 = n198 ^ n197 ^ x108 ;
  assign n200 = ( x1 & x7 ) | ( x1 & ~x28 ) | ( x7 & ~x28 ) ;
  assign n201 = ( x124 & n161 ) | ( x124 & ~n200 ) | ( n161 & ~n200 ) ;
  assign n206 = n183 ^ x75 ^ x52 ;
  assign n202 = x50 & ~n163 ;
  assign n203 = n202 ^ x3 ^ 1'b0 ;
  assign n204 = ( ~x66 & x97 ) | ( ~x66 & n203 ) | ( x97 & n203 ) ;
  assign n205 = n204 ^ x105 ^ x15 ;
  assign n207 = n206 ^ n205 ^ x113 ;
  assign n210 = x90 ^ x66 ^ 1'b0 ;
  assign n211 = x90 & n210 ;
  assign n212 = x13 & x89 ;
  assign n213 = ~n211 & n212 ;
  assign n214 = n213 ^ n134 ^ x55 ;
  assign n208 = x33 & ~n206 ;
  assign n209 = ~x24 & n208 ;
  assign n215 = n214 ^ n209 ^ 1'b0 ;
  assign n216 = x71 & ~n171 ;
  assign n217 = ~x35 & n216 ;
  assign n218 = n217 ^ n185 ^ x51 ;
  assign n219 = ( ~x100 & n183 ) | ( ~x100 & n213 ) | ( n183 & n213 ) ;
  assign n220 = n159 ^ n151 ^ x35 ;
  assign n221 = n220 ^ x6 ^ 1'b0 ;
  assign n222 = x59 & n221 ;
  assign n223 = n198 ^ x91 ^ 1'b0 ;
  assign n224 = ~n131 & n155 ;
  assign n225 = ~x105 & n224 ;
  assign n226 = x74 | n225 ;
  assign n227 = ( ~x84 & n223 ) | ( ~x84 & n226 ) | ( n223 & n226 ) ;
  assign n228 = x95 ^ x45 ^ 1'b0 ;
  assign n229 = x105 & n228 ;
  assign n230 = n229 ^ x100 ^ x18 ;
  assign n236 = n159 ^ n147 ^ n130 ;
  assign n237 = x23 & ~n236 ;
  assign n238 = n237 ^ x17 ^ 1'b0 ;
  assign n239 = ( x49 & ~n168 ) | ( x49 & n238 ) | ( ~n168 & n238 ) ;
  assign n240 = n179 ^ x127 ^ x36 ;
  assign n241 = n240 ^ x110 ^ 1'b0 ;
  assign n242 = n239 & n241 ;
  assign n243 = n242 ^ x77 ^ x2 ;
  assign n234 = n229 ^ x60 ^ x24 ;
  assign n231 = ( ~x57 & x60 ) | ( ~x57 & x67 ) | ( x60 & x67 ) ;
  assign n232 = n141 & n231 ;
  assign n233 = n232 ^ x126 ^ 1'b0 ;
  assign n235 = n234 ^ n233 ^ x26 ;
  assign n244 = n243 ^ n235 ^ 1'b0 ;
  assign n245 = ~x73 & n211 ;
  assign n246 = n245 ^ n147 ^ x95 ;
  assign n247 = ( x106 & n192 ) | ( x106 & n246 ) | ( n192 & n246 ) ;
  assign n248 = x24 & ~x53 ;
  assign n249 = n183 ^ n163 ^ 1'b0 ;
  assign n250 = x111 ^ x78 ^ x17 ;
  assign n251 = n171 | n250 ;
  assign n252 = n251 ^ x33 ^ 1'b0 ;
  assign n253 = ( x123 & n148 ) | ( x123 & ~n194 ) | ( n148 & ~n194 ) ;
  assign n254 = ( x65 & n252 ) | ( x65 & n253 ) | ( n252 & n253 ) ;
  assign n255 = x5 & x97 ;
  assign n256 = ~x32 & n255 ;
  assign n257 = ( x9 & x11 ) | ( x9 & n256 ) | ( x11 & n256 ) ;
  assign n258 = n257 ^ n235 ^ 1'b0 ;
  assign n259 = n254 & ~n258 ;
  assign n260 = x76 & ~n158 ;
  assign n262 = x16 & x113 ;
  assign n263 = n262 ^ x121 ^ 1'b0 ;
  assign n264 = n181 & n263 ;
  assign n265 = x56 & n264 ;
  assign n261 = n182 & ~n238 ;
  assign n266 = n265 ^ n261 ^ 1'b0 ;
  assign n267 = n138 ^ x17 ^ 1'b0 ;
  assign n271 = x59 & ~x84 ;
  assign n272 = n271 ^ x26 ^ x9 ;
  assign n268 = x86 ^ x46 ^ x37 ;
  assign n269 = x49 & ~n168 ;
  assign n270 = n268 & n269 ;
  assign n273 = n272 ^ n270 ^ x127 ;
  assign n274 = x94 & ~n138 ;
  assign n275 = ~n273 & n274 ;
  assign n276 = n182 & ~n275 ;
  assign n277 = ~x88 & n276 ;
  assign n281 = x105 ^ x21 ^ x15 ;
  assign n278 = x51 & ~n136 ;
  assign n279 = ~x43 & n278 ;
  assign n280 = x81 & ~n279 ;
  assign n282 = n281 ^ n280 ^ 1'b0 ;
  assign n283 = x103 & x114 ;
  assign n284 = n283 ^ n178 ^ 1'b0 ;
  assign n285 = ( n263 & n282 ) | ( n263 & ~n284 ) | ( n282 & ~n284 ) ;
  assign n286 = ( x87 & ~x106 ) | ( x87 & n253 ) | ( ~x106 & n253 ) ;
  assign n287 = n236 ^ n172 ^ x4 ;
  assign n299 = n161 & n198 ;
  assign n300 = ~x7 & n299 ;
  assign n298 = n133 ^ x51 ^ x17 ;
  assign n301 = n300 ^ n298 ^ 1'b0 ;
  assign n302 = n159 | n301 ;
  assign n296 = x20 & x126 ;
  assign n297 = n296 ^ x69 ^ 1'b0 ;
  assign n303 = n302 ^ n297 ^ 1'b0 ;
  assign n304 = x60 & n303 ;
  assign n288 = ( x82 & x127 ) | ( x82 & ~n149 ) | ( x127 & ~n149 ) ;
  assign n289 = n288 ^ n133 ^ x90 ;
  assign n293 = n271 ^ n148 ^ 1'b0 ;
  assign n290 = ~n142 & n172 ;
  assign n291 = n256 & n290 ;
  assign n292 = n291 ^ x120 ^ x16 ;
  assign n294 = n293 ^ n292 ^ n155 ;
  assign n295 = ( x14 & n289 ) | ( x14 & n294 ) | ( n289 & n294 ) ;
  assign n305 = n304 ^ n295 ^ x26 ;
  assign n309 = n279 ^ x16 ^ 1'b0 ;
  assign n306 = x5 & x88 ;
  assign n307 = n306 ^ x73 ^ 1'b0 ;
  assign n308 = n307 ^ n167 ^ x115 ;
  assign n310 = n309 ^ n308 ^ n148 ;
  assign n311 = n310 ^ x2 ^ 1'b0 ;
  assign n312 = n311 ^ n219 ^ x72 ;
  assign n313 = n164 ^ x83 ^ x45 ;
  assign n314 = x109 & n313 ;
  assign n321 = x54 & x100 ;
  assign n322 = n177 & n321 ;
  assign n318 = x88 & x96 ;
  assign n319 = n318 ^ x6 ^ 1'b0 ;
  assign n320 = n194 & ~n319 ;
  assign n323 = n322 ^ n320 ^ 1'b0 ;
  assign n316 = x72 & ~x89 ;
  assign n315 = x85 ^ x71 ^ 1'b0 ;
  assign n317 = n316 ^ n315 ^ n223 ;
  assign n324 = n323 ^ n317 ^ n150 ;
  assign n325 = n270 & n324 ;
  assign n328 = n158 ^ x94 ^ x55 ;
  assign n327 = x37 & ~n203 ;
  assign n329 = n328 ^ n327 ^ 1'b0 ;
  assign n326 = x101 ^ x40 ^ x28 ;
  assign n330 = n329 ^ n326 ^ x23 ;
  assign n331 = x5 & x27 ;
  assign n332 = ~x6 & n331 ;
  assign n333 = x97 & ~n332 ;
  assign n334 = ~x13 & n333 ;
  assign n335 = ( x114 & ~n153 ) | ( x114 & n300 ) | ( ~n153 & n300 ) ;
  assign n336 = n305 ^ x79 ^ 1'b0 ;
  assign n337 = n335 & ~n336 ;
  assign n338 = ( x40 & x120 ) | ( x40 & n294 ) | ( x120 & n294 ) ;
  assign n339 = x92 & ~n227 ;
  assign n340 = n339 ^ n178 ^ 1'b0 ;
  assign n341 = n340 ^ x56 ^ 1'b0 ;
  assign n342 = n338 & ~n341 ;
  assign n343 = n198 | n203 ;
  assign n344 = ~n192 & n343 ;
  assign n345 = n344 ^ x87 ^ 1'b0 ;
  assign n346 = n345 ^ n141 ^ x57 ;
  assign n358 = x71 ^ x45 ^ 1'b0 ;
  assign n359 = x41 & n358 ;
  assign n360 = ( ~x82 & n279 ) | ( ~x82 & n359 ) | ( n279 & n359 ) ;
  assign n361 = n360 ^ n195 ^ 1'b0 ;
  assign n362 = n328 | n361 ;
  assign n347 = n180 ^ n146 ^ 1'b0 ;
  assign n348 = x115 & n347 ;
  assign n349 = x71 & n348 ;
  assign n350 = ~x109 & n349 ;
  assign n351 = n350 ^ x0 ^ 1'b0 ;
  assign n353 = ( x84 & x107 ) | ( x84 & n236 ) | ( x107 & n236 ) ;
  assign n354 = ~n351 & n353 ;
  assign n355 = n354 ^ n153 ^ 1'b0 ;
  assign n356 = n355 ^ n263 ^ x94 ;
  assign n352 = n351 ^ n281 ^ n206 ;
  assign n357 = n356 ^ n352 ^ n131 ;
  assign n363 = n362 ^ n357 ^ 1'b0 ;
  assign n364 = n230 | n363 ;
  assign n365 = n257 ^ x5 ^ 1'b0 ;
  assign n366 = x124 ^ x56 ^ x39 ;
  assign n367 = n366 ^ n293 ^ 1'b0 ;
  assign n368 = n360 ^ x117 ^ x99 ;
  assign n369 = ( x49 & n231 ) | ( x49 & ~n368 ) | ( n231 & ~n368 ) ;
  assign n370 = n369 ^ n225 ^ x13 ;
  assign n371 = n166 ^ x120 ^ 1'b0 ;
  assign n372 = x97 & n371 ;
  assign n373 = x60 & ~x123 ;
  assign n374 = n373 ^ n142 ^ x5 ;
  assign n375 = ( n307 & n372 ) | ( n307 & ~n374 ) | ( n372 & ~n374 ) ;
  assign n382 = x117 ^ x13 ^ 1'b0 ;
  assign n383 = ~n271 & n382 ;
  assign n384 = ~n245 & n383 ;
  assign n385 = ~n156 & n384 ;
  assign n386 = n199 & ~n385 ;
  assign n387 = x120 & n386 ;
  assign n380 = n257 ^ n240 ^ x58 ;
  assign n376 = n155 ^ x93 ^ x26 ;
  assign n377 = n226 ^ x2 ^ 1'b0 ;
  assign n378 = n377 ^ n348 ^ x5 ;
  assign n379 = ( x26 & n376 ) | ( x26 & ~n378 ) | ( n376 & ~n378 ) ;
  assign n381 = n380 ^ n379 ^ x19 ;
  assign n388 = n387 ^ n381 ^ x44 ;
  assign n389 = ~n375 & n388 ;
  assign n390 = n389 ^ x4 ^ 1'b0 ;
  assign n392 = x79 & ~x90 ;
  assign n391 = x61 & ~n219 ;
  assign n393 = n392 ^ n391 ^ x94 ;
  assign n394 = ( x37 & x55 ) | ( x37 & ~x91 ) | ( x55 & ~x91 ) ;
  assign n395 = n394 ^ n159 ^ x18 ;
  assign n396 = n395 ^ x28 ^ 1'b0 ;
  assign n397 = n229 & n396 ;
  assign n398 = x57 & n397 ;
  assign n399 = n238 & n398 ;
  assign n403 = x14 & x99 ;
  assign n404 = n403 ^ x11 ^ 1'b0 ;
  assign n405 = n315 & n404 ;
  assign n401 = x60 ^ x5 ^ 1'b0 ;
  assign n400 = n166 & n369 ;
  assign n402 = n401 ^ n400 ^ 1'b0 ;
  assign n406 = n405 ^ n402 ^ x48 ;
  assign n407 = n366 ^ x87 ^ x42 ;
  assign n408 = n171 & n407 ;
  assign n411 = x127 ^ x10 ^ 1'b0 ;
  assign n412 = x119 & n411 ;
  assign n413 = ( x99 & ~n373 ) | ( x99 & n412 ) | ( ~n373 & n412 ) ;
  assign n414 = n413 ^ x108 ^ x90 ;
  assign n415 = ( ~x18 & n323 ) | ( ~x18 & n414 ) | ( n323 & n414 ) ;
  assign n410 = n171 ^ x45 ^ x14 ;
  assign n409 = n227 ^ n204 ^ n169 ;
  assign n416 = n415 ^ n410 ^ n409 ;
  assign n417 = n137 & ~n250 ;
  assign n418 = n197 & n417 ;
  assign n419 = x54 & x103 ;
  assign n420 = n419 ^ x39 ^ 1'b0 ;
  assign n421 = ( n151 & n231 ) | ( n151 & n420 ) | ( n231 & n420 ) ;
  assign n422 = n226 ^ n201 ^ 1'b0 ;
  assign n423 = x85 & x87 ;
  assign n424 = n423 ^ x57 ^ 1'b0 ;
  assign n425 = n424 ^ x108 ^ 1'b0 ;
  assign n426 = n422 | n425 ;
  assign n427 = x123 & n185 ;
  assign n428 = n160 ^ x27 ^ 1'b0 ;
  assign n429 = ( x18 & ~x24 ) | ( x18 & n302 ) | ( ~x24 & n302 ) ;
  assign n430 = n429 ^ n133 ^ 1'b0 ;
  assign n431 = n428 & n430 ;
  assign n432 = x61 ^ x17 ^ 1'b0 ;
  assign n433 = ( n427 & ~n431 ) | ( n427 & n432 ) | ( ~n431 & n432 ) ;
  assign n434 = x47 & ~n145 ;
  assign n435 = ( n305 & n433 ) | ( n305 & n434 ) | ( n433 & n434 ) ;
  assign n436 = ~x120 & n343 ;
  assign n437 = n436 ^ n148 ^ 1'b0 ;
  assign n438 = n315 ^ x94 ^ 1'b0 ;
  assign n440 = ( ~x58 & x117 ) | ( ~x58 & n134 ) | ( x117 & n134 ) ;
  assign n439 = x71 & n205 ;
  assign n441 = n440 ^ n439 ^ 1'b0 ;
  assign n442 = n359 ^ x43 ^ 1'b0 ;
  assign n443 = ( n131 & n142 ) | ( n131 & ~n165 ) | ( n142 & ~n165 ) ;
  assign n444 = n443 ^ x23 ^ x2 ;
  assign n445 = ( n365 & n442 ) | ( n365 & ~n444 ) | ( n442 & ~n444 ) ;
  assign n446 = n441 & n445 ;
  assign n447 = n169 & n446 ;
  assign n448 = ~n169 & n359 ;
  assign n449 = ~n394 & n448 ;
  assign n450 = n413 & n449 ;
  assign n451 = ( x33 & x115 ) | ( x33 & n169 ) | ( x115 & n169 ) ;
  assign n452 = ( ~x38 & x114 ) | ( ~x38 & n153 ) | ( x114 & n153 ) ;
  assign n453 = ~n256 & n452 ;
  assign n454 = ( x74 & ~x78 ) | ( x74 & n453 ) | ( ~x78 & n453 ) ;
  assign n455 = x18 & n454 ;
  assign n456 = ~n451 & n455 ;
  assign n460 = n443 ^ x30 ^ 1'b0 ;
  assign n461 = x116 & ~n460 ;
  assign n457 = ( x78 & x122 ) | ( x78 & n319 ) | ( x122 & n319 ) ;
  assign n458 = x100 & n457 ;
  assign n459 = n163 & n458 ;
  assign n462 = n461 ^ n459 ^ 1'b0 ;
  assign n463 = n223 & ~n279 ;
  assign n464 = n463 ^ n207 ^ 1'b0 ;
  assign n465 = ( n192 & ~n462 ) | ( n192 & n464 ) | ( ~n462 & n464 ) ;
  assign n466 = n159 ^ n143 ^ x102 ;
  assign n467 = n394 & n466 ;
  assign n468 = n467 ^ x108 ^ 1'b0 ;
  assign n469 = n468 ^ n201 ^ 1'b0 ;
  assign n470 = n421 & ~n469 ;
  assign n471 = ~n145 & n470 ;
  assign n472 = n397 ^ n272 ^ n145 ;
  assign n473 = n350 ^ x72 ^ 1'b0 ;
  assign n474 = n322 | n473 ;
  assign n475 = n474 ^ x94 ^ 1'b0 ;
  assign n476 = n472 | n475 ;
  assign n477 = n316 ^ x93 ^ 1'b0 ;
  assign n478 = n477 ^ n284 ^ x97 ;
  assign n479 = ( x96 & n214 ) | ( x96 & ~n431 ) | ( n214 & ~n431 ) ;
  assign n480 = n479 ^ n353 ^ x100 ;
  assign n481 = x57 & n345 ;
  assign n482 = n220 & ~n481 ;
  assign n483 = ~n386 & n482 ;
  assign n484 = x0 | n483 ;
  assign n485 = ( x30 & ~n151 ) | ( x30 & n211 ) | ( ~n151 & n211 ) ;
  assign n486 = n485 ^ n366 ^ 1'b0 ;
  assign n487 = n309 & n317 ;
  assign n488 = ~n167 & n487 ;
  assign n489 = n488 ^ n445 ^ n405 ;
  assign n490 = n308 ^ n153 ^ 1'b0 ;
  assign n491 = n203 | n452 ;
  assign n492 = x12 | n491 ;
  assign n493 = n492 ^ x93 ^ x57 ;
  assign n494 = n133 | n493 ;
  assign n495 = n490 | n494 ;
  assign n496 = n492 ^ n186 ^ 1'b0 ;
  assign n497 = n129 & ~n496 ;
  assign n498 = n141 & n497 ;
  assign n499 = ~x52 & n498 ;
  assign n500 = n307 ^ x115 ^ x85 ;
  assign n501 = n500 ^ n256 ^ 1'b0 ;
  assign n502 = n415 ^ n220 ^ 1'b0 ;
  assign n503 = n380 | n502 ;
  assign n507 = x46 & x51 ;
  assign n508 = n507 ^ n273 ^ 1'b0 ;
  assign n504 = n214 ^ x60 ^ 1'b0 ;
  assign n505 = n288 & n504 ;
  assign n506 = n505 ^ n170 ^ 1'b0 ;
  assign n509 = n508 ^ n506 ^ x126 ;
  assign n510 = ~x53 & n201 ;
  assign n511 = n510 ^ n447 ^ n434 ;
  assign n512 = n511 ^ n369 ^ x52 ;
  assign n513 = x59 ^ x10 ^ 1'b0 ;
  assign n514 = x24 & n513 ;
  assign n515 = n514 ^ n225 ^ 1'b0 ;
  assign n516 = x95 & n147 ;
  assign n517 = n345 & n516 ;
  assign n518 = n517 ^ n259 ^ n249 ;
  assign n519 = n518 ^ n445 ^ n338 ;
  assign n520 = n414 ^ n236 ^ x118 ;
  assign n521 = n427 & ~n520 ;
  assign n522 = n521 ^ n300 ^ 1'b0 ;
  assign n523 = ( x80 & n345 ) | ( x80 & ~n522 ) | ( n345 & ~n522 ) ;
  assign n524 = n523 ^ n142 ^ x65 ;
  assign n525 = n148 ^ x54 ^ x4 ;
  assign n526 = n525 ^ n523 ^ n172 ;
  assign n527 = ( n158 & n179 ) | ( n158 & ~n342 ) | ( n179 & ~n342 ) ;
  assign n530 = n293 ^ x114 ^ x112 ;
  assign n528 = n195 & ~n345 ;
  assign n529 = n449 & n528 ;
  assign n531 = n530 ^ n529 ^ 1'b0 ;
  assign n532 = ( x75 & ~n231 ) | ( x75 & n531 ) | ( ~n231 & n531 ) ;
  assign n533 = n532 ^ n145 ^ 1'b0 ;
  assign n540 = n198 ^ x100 ^ x14 ;
  assign n535 = n271 ^ x86 ^ 1'b0 ;
  assign n536 = n146 | n535 ;
  assign n537 = ( x27 & x127 ) | ( x27 & n530 ) | ( x127 & n530 ) ;
  assign n538 = x76 & ~n537 ;
  assign n539 = ( ~n385 & n536 ) | ( ~n385 & n538 ) | ( n536 & n538 ) ;
  assign n541 = n540 ^ n539 ^ n375 ;
  assign n534 = ~n263 & n356 ;
  assign n542 = n541 ^ n534 ^ 1'b0 ;
  assign n543 = ( x69 & n366 ) | ( x69 & ~n420 ) | ( n366 & ~n420 ) ;
  assign n544 = ( x45 & n529 ) | ( x45 & ~n543 ) | ( n529 & ~n543 ) ;
  assign n545 = n256 ^ x112 ^ x48 ;
  assign n546 = ~n197 & n545 ;
  assign n547 = n544 & n546 ;
  assign n548 = x73 & n393 ;
  assign n549 = n548 ^ n523 ^ 1'b0 ;
  assign n554 = x114 & ~n130 ;
  assign n555 = n554 ^ x57 ^ 1'b0 ;
  assign n551 = n164 & ~n394 ;
  assign n550 = n449 ^ n284 ^ n174 ;
  assign n552 = n551 ^ n550 ^ 1'b0 ;
  assign n553 = n381 | n552 ;
  assign n556 = n555 ^ n553 ^ n434 ;
  assign n557 = ( n547 & n549 ) | ( n547 & n556 ) | ( n549 & n556 ) ;
  assign n561 = x43 ^ x42 ^ 1'b0 ;
  assign n562 = ( ~n388 & n529 ) | ( ~n388 & n561 ) | ( n529 & n561 ) ;
  assign n558 = x81 ^ x72 ^ 1'b0 ;
  assign n559 = x61 & n558 ;
  assign n560 = n497 & n559 ;
  assign n563 = n562 ^ n560 ^ 1'b0 ;
  assign n564 = x95 & ~n180 ;
  assign n565 = n564 ^ x8 ^ 1'b0 ;
  assign n566 = n429 ^ n372 ^ 1'b0 ;
  assign n567 = n565 | n566 ;
  assign n568 = n567 ^ n203 ^ 1'b0 ;
  assign n569 = x18 & n407 ;
  assign n570 = ( n536 & ~n568 ) | ( n536 & n569 ) | ( ~n568 & n569 ) ;
  assign n572 = x91 ^ x28 ^ x13 ;
  assign n573 = n572 ^ n407 ^ n279 ;
  assign n574 = n573 ^ n366 ^ 1'b0 ;
  assign n575 = n231 & n574 ;
  assign n571 = x113 & ~n379 ;
  assign n576 = n575 ^ n571 ^ 1'b0 ;
  assign n577 = n527 ^ n401 ^ 1'b0 ;
  assign n578 = x20 & n156 ;
  assign n579 = n578 ^ n198 ^ 1'b0 ;
  assign n580 = ( ~x112 & n171 ) | ( ~x112 & n393 ) | ( n171 & n393 ) ;
  assign n581 = n580 ^ n568 ^ 1'b0 ;
  assign n582 = n272 ^ n233 ^ n226 ;
  assign n583 = ( x2 & ~n293 ) | ( x2 & n582 ) | ( ~n293 & n582 ) ;
  assign n584 = n493 ^ n360 ^ x38 ;
  assign n585 = n352 & ~n584 ;
  assign n586 = ~n353 & n585 ;
  assign n587 = n364 | n586 ;
  assign n588 = n587 ^ n519 ^ 1'b0 ;
  assign n589 = ( n313 & n420 ) | ( n313 & ~n530 ) | ( n420 & ~n530 ) ;
  assign n597 = ( x31 & ~n429 ) | ( x31 & n449 ) | ( ~n429 & n449 ) ;
  assign n590 = ( x122 & n244 ) | ( x122 & ~n395 ) | ( n244 & ~n395 ) ;
  assign n591 = n590 ^ n134 ^ x61 ;
  assign n592 = ( x65 & n157 ) | ( x65 & n591 ) | ( n157 & n591 ) ;
  assign n593 = n178 & n179 ;
  assign n594 = n353 & ~n593 ;
  assign n595 = n429 & n594 ;
  assign n596 = n592 | n595 ;
  assign n598 = n597 ^ n596 ^ 1'b0 ;
  assign n599 = ( ~x36 & x57 ) | ( ~x36 & n526 ) | ( x57 & n526 ) ;
  assign n600 = n599 ^ n593 ^ 1'b0 ;
  assign n601 = ( n141 & n245 ) | ( n141 & ~n275 ) | ( n245 & ~n275 ) ;
  assign n602 = n181 ^ x99 ^ 1'b0 ;
  assign n604 = ( x0 & n167 ) | ( x0 & n234 ) | ( n167 & n234 ) ;
  assign n605 = n604 ^ n209 ^ 1'b0 ;
  assign n603 = n260 & n372 ;
  assign n606 = n605 ^ n603 ^ 1'b0 ;
  assign n609 = n544 ^ n462 ^ 1'b0 ;
  assign n607 = n273 ^ n180 ^ x32 ;
  assign n608 = ~n190 & n607 ;
  assign n610 = n609 ^ n608 ^ 1'b0 ;
  assign n611 = ( n138 & n231 ) | ( n138 & ~n385 ) | ( n231 & ~n385 ) ;
  assign n612 = ( x60 & n138 ) | ( x60 & ~n316 ) | ( n138 & ~n316 ) ;
  assign n613 = ~n153 & n612 ;
  assign n614 = ~n611 & n613 ;
  assign n615 = ( x20 & ~n316 ) | ( x20 & n614 ) | ( ~n316 & n614 ) ;
  assign n616 = n129 ^ x37 ^ 1'b0 ;
  assign n617 = n616 ^ n213 ^ 1'b0 ;
  assign n618 = ( ~n142 & n615 ) | ( ~n142 & n617 ) | ( n615 & n617 ) ;
  assign n619 = n618 ^ x90 ^ x15 ;
  assign n620 = n289 ^ n192 ^ x20 ;
  assign n621 = n620 ^ n532 ^ x35 ;
  assign n624 = n449 ^ n240 ^ x127 ;
  assign n625 = n624 ^ n172 ^ n145 ;
  assign n622 = n368 & n555 ;
  assign n623 = ~n350 & n622 ;
  assign n626 = n625 ^ n623 ^ 1'b0 ;
  assign n627 = n305 ^ n246 ^ 1'b0 ;
  assign n628 = n330 & ~n627 ;
  assign n629 = n149 ^ n133 ^ 1'b0 ;
  assign n630 = n604 ^ n158 ^ 1'b0 ;
  assign n631 = n629 & n630 ;
  assign n632 = n198 ^ x109 ^ x26 ;
  assign n633 = n201 & n632 ;
  assign n635 = x93 ^ x85 ^ 1'b0 ;
  assign n634 = n195 & n461 ;
  assign n636 = n635 ^ n634 ^ 1'b0 ;
  assign n637 = n636 ^ n415 ^ n309 ;
  assign n638 = x63 & ~n637 ;
  assign n639 = n633 & n638 ;
  assign n642 = x115 ^ x89 ^ 1'b0 ;
  assign n643 = n642 ^ n394 ^ n322 ;
  assign n640 = n297 ^ x101 ^ 1'b0 ;
  assign n641 = x93 & ~n640 ;
  assign n644 = n643 ^ n641 ^ n364 ;
  assign n645 = ( x91 & ~x100 ) | ( x91 & n130 ) | ( ~x100 & n130 ) ;
  assign n646 = x8 & ~x45 ;
  assign n647 = n646 ^ x126 ^ 1'b0 ;
  assign n648 = n645 | n647 ;
  assign n649 = n526 | n648 ;
  assign n650 = ( n267 & ~n644 ) | ( n267 & n649 ) | ( ~n644 & n649 ) ;
  assign n651 = n300 | n350 ;
  assign n652 = n651 ^ x68 ^ 1'b0 ;
  assign n653 = n215 ^ n209 ^ x73 ;
  assign n654 = ( n300 & n368 ) | ( n300 & n653 ) | ( n368 & n653 ) ;
  assign n655 = n654 ^ n397 ^ 1'b0 ;
  assign n656 = ~n652 & n655 ;
  assign n657 = n656 ^ n639 ^ n606 ;
  assign n658 = n291 | n429 ;
  assign n659 = n436 & ~n658 ;
  assign n660 = ( x60 & ~x97 ) | ( x60 & x122 ) | ( ~x97 & x122 ) ;
  assign n669 = n359 ^ x94 ^ 1'b0 ;
  assign n670 = x44 & n669 ;
  assign n671 = n243 ^ x92 ^ 1'b0 ;
  assign n672 = n670 & ~n671 ;
  assign n673 = n672 ^ x107 ^ x66 ;
  assign n668 = x73 & ~n420 ;
  assign n674 = n673 ^ n668 ^ 1'b0 ;
  assign n664 = n457 ^ n309 ^ x50 ;
  assign n665 = n664 ^ n412 ^ x123 ;
  assign n666 = x105 & n665 ;
  assign n667 = ~n272 & n666 ;
  assign n675 = n674 ^ n667 ^ 1'b0 ;
  assign n676 = n265 | n675 ;
  assign n680 = n537 ^ n231 ^ x4 ;
  assign n681 = n680 ^ n230 ^ n187 ;
  assign n682 = n136 | n681 ;
  assign n683 = n246 | n682 ;
  assign n684 = n683 ^ n137 ^ n133 ;
  assign n677 = n648 ^ n544 ^ x70 ;
  assign n678 = ( x72 & n323 ) | ( x72 & n677 ) | ( n323 & n677 ) ;
  assign n679 = n607 & n678 ;
  assign n685 = n684 ^ n679 ^ 1'b0 ;
  assign n686 = n676 & ~n685 ;
  assign n661 = n319 ^ n150 ^ 1'b0 ;
  assign n662 = ~n530 & n661 ;
  assign n663 = n662 ^ x76 ^ 1'b0 ;
  assign n687 = n686 ^ n663 ^ 1'b0 ;
  assign n688 = n660 & ~n687 ;
  assign n689 = x40 & n394 ;
  assign n690 = ~n156 & n689 ;
  assign n691 = n690 ^ n207 ^ 1'b0 ;
  assign n692 = n691 ^ n194 ^ 1'b0 ;
  assign n693 = x98 & n324 ;
  assign n694 = n693 ^ x43 ^ 1'b0 ;
  assign n695 = x90 ^ x70 ^ x18 ;
  assign n696 = ( n688 & n694 ) | ( n688 & ~n695 ) | ( n694 & ~n695 ) ;
  assign n697 = n600 ^ x121 ^ x59 ;
  assign n698 = n158 | n270 ;
  assign n699 = n660 ^ n504 ^ n420 ;
  assign n700 = ( x34 & ~n698 ) | ( x34 & n699 ) | ( ~n698 & n699 ) ;
  assign n701 = x91 & n166 ;
  assign n702 = n701 ^ n654 ^ 1'b0 ;
  assign n703 = n462 ^ x120 ^ x73 ;
  assign n704 = n203 | n551 ;
  assign n705 = n704 ^ n394 ^ 1'b0 ;
  assign n706 = ( x25 & n149 ) | ( x25 & ~n705 ) | ( n149 & ~n705 ) ;
  assign n707 = n161 & ~n582 ;
  assign n708 = n707 ^ x69 ^ 1'b0 ;
  assign n709 = ( ~n300 & n392 ) | ( ~n300 & n708 ) | ( n392 & n708 ) ;
  assign n712 = ( ~x78 & x118 ) | ( ~x78 & n236 ) | ( x118 & n236 ) ;
  assign n713 = ( x58 & n165 ) | ( x58 & ~n712 ) | ( n165 & ~n712 ) ;
  assign n710 = ( x43 & ~x49 ) | ( x43 & x125 ) | ( ~x49 & x125 ) ;
  assign n711 = ( x96 & n636 ) | ( x96 & ~n710 ) | ( n636 & ~n710 ) ;
  assign n714 = n713 ^ n711 ^ n383 ;
  assign n715 = ~n219 & n714 ;
  assign n716 = n709 & n715 ;
  assign n717 = ( n703 & n706 ) | ( n703 & n716 ) | ( n706 & n716 ) ;
  assign n718 = ~n214 & n717 ;
  assign n719 = n702 & n718 ;
  assign n720 = n719 ^ n386 ^ n285 ;
  assign n721 = n380 ^ n217 ^ 1'b0 ;
  assign n722 = ~n319 & n721 ;
  assign n723 = x111 & n532 ;
  assign n724 = ~x106 & n723 ;
  assign n725 = n531 ^ n492 ^ n441 ;
  assign n726 = n710 ^ n635 ^ 1'b0 ;
  assign n727 = ~n725 & n726 ;
  assign n728 = ~x13 & n727 ;
  assign n729 = n691 ^ n680 ^ n142 ;
  assign n730 = ( ~x46 & x95 ) | ( ~x46 & n146 ) | ( x95 & n146 ) ;
  assign n731 = ( n259 & n329 ) | ( n259 & n730 ) | ( n329 & n730 ) ;
  assign n732 = n512 & n731 ;
  assign n733 = ( ~n165 & n205 ) | ( ~n165 & n226 ) | ( n205 & n226 ) ;
  assign n734 = n733 ^ n428 ^ n248 ;
  assign n735 = n579 ^ n203 ^ 1'b0 ;
  assign n736 = ~n573 & n735 ;
  assign n737 = ~n579 & n736 ;
  assign n738 = ~n304 & n737 ;
  assign n739 = x84 & ~n738 ;
  assign n740 = ~n734 & n739 ;
  assign n741 = ( x60 & x91 ) | ( x60 & n447 ) | ( x91 & n447 ) ;
  assign n742 = x82 & n231 ;
  assign n743 = ~n466 & n742 ;
  assign n744 = ( x114 & ~n184 ) | ( x114 & n743 ) | ( ~n184 & n743 ) ;
  assign n745 = n744 ^ n495 ^ 1'b0 ;
  assign n746 = x66 | n745 ;
  assign n750 = n443 ^ n137 ^ x60 ;
  assign n749 = n263 | n582 ;
  assign n751 = n750 ^ n749 ^ 1'b0 ;
  assign n747 = n366 ^ n335 ^ 1'b0 ;
  assign n748 = ( n708 & n711 ) | ( n708 & ~n747 ) | ( n711 & ~n747 ) ;
  assign n752 = n751 ^ n748 ^ n379 ;
  assign n753 = n199 ^ x100 ^ x31 ;
  assign n755 = n543 ^ n186 ^ 1'b0 ;
  assign n756 = x33 & ~n755 ;
  assign n754 = n377 ^ n272 ^ n240 ;
  assign n757 = n756 ^ n754 ^ x27 ;
  assign n758 = n416 ^ n197 ^ x17 ;
  assign n759 = n254 ^ x71 ^ 1'b0 ;
  assign n760 = n414 ^ n178 ^ n161 ;
  assign n761 = n760 ^ x70 ^ 1'b0 ;
  assign n762 = n759 & n761 ;
  assign n763 = ( x96 & x101 ) | ( x96 & ~n762 ) | ( x101 & ~n762 ) ;
  assign n764 = ( n625 & ~n758 ) | ( n625 & n763 ) | ( ~n758 & n763 ) ;
  assign n765 = ( x9 & ~n298 ) | ( x9 & n436 ) | ( ~n298 & n436 ) ;
  assign n766 = n765 ^ n751 ^ n162 ;
  assign n767 = n424 ^ n319 ^ x103 ;
  assign n768 = n767 ^ n346 ^ x41 ;
  assign n769 = n353 ^ x65 ^ 1'b0 ;
  assign n770 = x23 & n769 ;
  assign n771 = n770 ^ n531 ^ n360 ;
  assign n772 = n771 ^ n372 ^ x42 ;
  assign n773 = ( n766 & n768 ) | ( n766 & n772 ) | ( n768 & n772 ) ;
  assign n774 = ( x25 & ~x62 ) | ( x25 & n168 ) | ( ~x62 & n168 ) ;
  assign n775 = n568 ^ n474 ^ n307 ;
  assign n776 = ~n774 & n775 ;
  assign n777 = n773 & n776 ;
  assign n778 = n167 ^ n138 ^ n130 ;
  assign n779 = n778 ^ n291 ^ 1'b0 ;
  assign n780 = n373 & n779 ;
  assign n781 = n543 & ~n606 ;
  assign n782 = n781 ^ n597 ^ 1'b0 ;
  assign n783 = n530 ^ n201 ^ 1'b0 ;
  assign n784 = x126 & ~n268 ;
  assign n785 = ~n654 & n784 ;
  assign n786 = n138 ^ x75 ^ 1'b0 ;
  assign n787 = ( x79 & n186 ) | ( x79 & n256 ) | ( n186 & n256 ) ;
  assign n788 = ( n765 & n786 ) | ( n765 & ~n787 ) | ( n786 & ~n787 ) ;
  assign n789 = n369 & n401 ;
  assign n790 = ~n674 & n789 ;
  assign n791 = n691 | n790 ;
  assign n792 = n416 | n791 ;
  assign n793 = n454 ^ n319 ^ 1'b0 ;
  assign n794 = n711 | n793 ;
  assign n795 = n794 ^ n537 ^ n170 ;
  assign n796 = ( n352 & ~n508 ) | ( n352 & n795 ) | ( ~n508 & n795 ) ;
  assign n797 = x16 & ~n190 ;
  assign n798 = n797 ^ x77 ^ 1'b0 ;
  assign n799 = n798 ^ x62 ^ 1'b0 ;
  assign n800 = x61 & ~n799 ;
  assign n801 = n279 ^ n270 ^ x90 ;
  assign n802 = ( ~x25 & n415 ) | ( ~x25 & n434 ) | ( n415 & n434 ) ;
  assign n803 = ~n801 & n802 ;
  assign n804 = n744 | n803 ;
  assign n805 = n804 ^ n159 ^ 1'b0 ;
  assign n806 = n805 ^ n654 ^ x117 ;
  assign n807 = n227 ^ n217 ^ x68 ;
  assign n808 = n807 ^ n479 ^ n177 ;
  assign n809 = x20 & ~n163 ;
  assign n810 = n364 & n809 ;
  assign n811 = n628 | n810 ;
  assign n812 = n355 & ~n478 ;
  assign n813 = ~x52 & n812 ;
  assign n814 = n813 ^ n312 ^ n131 ;
  assign n815 = n257 ^ n185 ^ x127 ;
  assign n816 = ( x3 & ~x29 ) | ( x3 & n815 ) | ( ~x29 & n815 ) ;
  assign n817 = n654 ^ n355 ^ 1'b0 ;
  assign n818 = n394 & n726 ;
  assign n819 = n818 ^ n334 ^ 1'b0 ;
  assign n821 = ( n272 & n298 ) | ( n272 & ~n525 ) | ( n298 & ~n525 ) ;
  assign n820 = ~n267 & n346 ;
  assign n822 = n821 ^ n820 ^ 1'b0 ;
  assign n823 = ( n616 & n819 ) | ( n616 & n822 ) | ( n819 & n822 ) ;
  assign n824 = n823 ^ x70 ^ 1'b0 ;
  assign n825 = n824 ^ n672 ^ n295 ;
  assign n826 = n825 ^ n158 ^ n130 ;
  assign n827 = n509 & n644 ;
  assign n828 = ~n317 & n827 ;
  assign n829 = n828 ^ n264 ^ n155 ;
  assign n830 = n829 ^ n307 ^ 1'b0 ;
  assign n831 = n614 ^ n383 ^ n293 ;
  assign n832 = ( n147 & n441 ) | ( n147 & ~n831 ) | ( n441 & ~n831 ) ;
  assign n833 = ~n190 & n665 ;
  assign n834 = n833 ^ x74 ^ 1'b0 ;
  assign n835 = ( ~n367 & n734 ) | ( ~n367 & n834 ) | ( n734 & n834 ) ;
  assign n837 = ~n377 & n444 ;
  assign n838 = n837 ^ n319 ^ 1'b0 ;
  assign n836 = ( x29 & ~x54 ) | ( x29 & x121 ) | ( ~x54 & x121 ) ;
  assign n839 = n838 ^ n836 ^ 1'b0 ;
  assign n840 = n839 ^ n462 ^ 1'b0 ;
  assign n845 = n229 & n324 ;
  assign n846 = n845 ^ n156 ^ 1'b0 ;
  assign n841 = x30 & n575 ;
  assign n842 = n841 ^ n289 ^ 1'b0 ;
  assign n843 = x77 & ~n842 ;
  assign n844 = n843 ^ n422 ^ 1'b0 ;
  assign n847 = n846 ^ n844 ^ n775 ;
  assign n852 = x19 & n756 ;
  assign n853 = n138 & n852 ;
  assign n854 = n252 & n853 ;
  assign n855 = n705 ^ x109 ^ 1'b0 ;
  assign n856 = n607 & n855 ;
  assign n857 = ( x10 & ~n854 ) | ( x10 & n856 ) | ( ~n854 & n856 ) ;
  assign n848 = n177 | n591 ;
  assign n849 = n848 ^ n268 ^ 1'b0 ;
  assign n850 = n580 ^ n468 ^ n260 ;
  assign n851 = n849 | n850 ;
  assign n858 = n857 ^ n851 ^ 1'b0 ;
  assign n859 = n489 ^ n459 ^ 1'b0 ;
  assign n860 = x50 & n684 ;
  assign n861 = n860 ^ x84 ^ 1'b0 ;
  assign n862 = n518 | n849 ;
  assign n863 = n862 ^ x109 ^ 1'b0 ;
  assign n864 = x33 & n863 ;
  assign n865 = n864 ^ n415 ^ 1'b0 ;
  assign n866 = ( n267 & n637 ) | ( n267 & n865 ) | ( n637 & n865 ) ;
  assign n867 = ( n525 & n861 ) | ( n525 & n866 ) | ( n861 & n866 ) ;
  assign n868 = n461 ^ n259 ^ 1'b0 ;
  assign n869 = n660 & n868 ;
  assign n870 = n869 ^ n780 ^ 1'b0 ;
  assign n871 = ~n853 & n870 ;
  assign n872 = ( x6 & n267 ) | ( x6 & n710 ) | ( n267 & n710 ) ;
  assign n873 = ~n681 & n872 ;
  assign n874 = ~n356 & n873 ;
  assign n875 = ( n338 & n694 ) | ( n338 & ~n713 ) | ( n694 & ~n713 ) ;
  assign n876 = n738 ^ n377 ^ 1'b0 ;
  assign n877 = ~n875 & n876 ;
  assign n878 = n874 & n877 ;
  assign n883 = ( ~x3 & x66 ) | ( ~x3 & n615 ) | ( x66 & n615 ) ;
  assign n884 = n883 ^ n357 ^ x36 ;
  assign n882 = x79 & n674 ;
  assign n885 = n884 ^ n882 ^ 1'b0 ;
  assign n880 = n169 ^ x68 ^ 1'b0 ;
  assign n879 = ( x119 & n211 ) | ( x119 & ~n819 ) | ( n211 & ~n819 ) ;
  assign n881 = n880 ^ n879 ^ n743 ;
  assign n886 = n885 ^ n881 ^ n747 ;
  assign n887 = n176 ^ x124 ^ 1'b0 ;
  assign n888 = ( n390 & ~n418 ) | ( n390 & n887 ) | ( ~n418 & n887 ) ;
  assign n889 = x87 & x107 ;
  assign n890 = n236 & n889 ;
  assign n891 = n890 ^ n831 ^ n223 ;
  assign n892 = n888 & n891 ;
  assign n893 = x117 & n190 ;
  assign n894 = n796 & n893 ;
  assign n895 = ( ~x102 & n656 ) | ( ~x102 & n674 ) | ( n656 & n674 ) ;
  assign n896 = ~n568 & n895 ;
  assign n897 = n359 ^ x72 ^ x47 ;
  assign n898 = ( x124 & ~n200 ) | ( x124 & n897 ) | ( ~n200 & n897 ) ;
  assign n899 = n898 ^ x38 ^ 1'b0 ;
  assign n900 = n317 & ~n899 ;
  assign n901 = n624 ^ x81 ^ 1'b0 ;
  assign n902 = n293 & n410 ;
  assign n903 = n901 & n902 ;
  assign n904 = x73 ^ x48 ^ 1'b0 ;
  assign n905 = n903 | n904 ;
  assign n906 = ( n265 & ~n418 ) | ( n265 & n471 ) | ( ~n418 & n471 ) ;
  assign n907 = ( x58 & n646 ) | ( x58 & n906 ) | ( n646 & n906 ) ;
  assign n909 = ( x72 & ~n313 ) | ( x72 & n322 ) | ( ~n313 & n322 ) ;
  assign n908 = x67 & n808 ;
  assign n910 = n909 ^ n908 ^ 1'b0 ;
  assign n911 = n849 ^ n264 ^ x2 ;
  assign n912 = ( n240 & n298 ) | ( n240 & n911 ) | ( n298 & n911 ) ;
  assign n913 = n509 ^ n377 ^ n182 ;
  assign n914 = n913 ^ n839 ^ 1'b0 ;
  assign n915 = n760 & n914 ;
  assign n916 = n242 ^ n205 ^ x46 ;
  assign n917 = n656 ^ n319 ^ 1'b0 ;
  assign n918 = n813 | n917 ;
  assign n919 = x72 & n918 ;
  assign n920 = n919 ^ x99 ^ 1'b0 ;
  assign n921 = n866 | n920 ;
  assign n923 = x10 & x65 ;
  assign n924 = n242 ^ x43 ^ x14 ;
  assign n925 = ( n334 & n923 ) | ( n334 & n924 ) | ( n923 & n924 ) ;
  assign n926 = n925 ^ n242 ^ x16 ;
  assign n922 = n253 | n621 ;
  assign n927 = n926 ^ n922 ^ 1'b0 ;
  assign n928 = n611 & n750 ;
  assign n929 = ~n760 & n928 ;
  assign n930 = x90 & ~n890 ;
  assign n931 = ~n821 & n930 ;
  assign n932 = n931 ^ n345 ^ 1'b0 ;
  assign n933 = ~n929 & n932 ;
  assign n935 = x36 | n136 ;
  assign n934 = n683 ^ n397 ^ n292 ;
  assign n936 = n935 ^ n934 ^ 1'b0 ;
  assign n937 = n163 | n936 ;
  assign n938 = n328 ^ n136 ^ 1'b0 ;
  assign n939 = ~n937 & n938 ;
  assign n940 = n939 ^ n728 ^ 1'b0 ;
  assign n941 = n933 & ~n940 ;
  assign n942 = x38 ^ x17 ^ 1'b0 ;
  assign n943 = n201 & n942 ;
  assign n944 = n187 ^ n142 ^ 1'b0 ;
  assign n945 = n943 & ~n944 ;
  assign n946 = n444 & n945 ;
  assign n947 = n946 ^ n839 ^ 1'b0 ;
  assign n948 = n133 | n947 ;
  assign n953 = ( n227 & ~n557 ) | ( n227 & n676 ) | ( ~n557 & n676 ) ;
  assign n949 = x110 ^ x100 ^ x62 ;
  assign n950 = n949 ^ n582 ^ 1'b0 ;
  assign n951 = n523 ^ n338 ^ 1'b0 ;
  assign n952 = n950 & ~n951 ;
  assign n954 = n953 ^ n952 ^ 1'b0 ;
  assign n955 = ~n711 & n954 ;
  assign n956 = n650 ^ n222 ^ x125 ;
  assign n957 = x82 & ~n183 ;
  assign n958 = ~x3 & x102 ;
  assign n959 = n958 ^ n340 ^ 1'b0 ;
  assign n960 = ~n957 & n959 ;
  assign n961 = x0 & n960 ;
  assign n962 = ( ~n165 & n328 ) | ( ~n165 & n383 ) | ( n328 & n383 ) ;
  assign n963 = ~n281 & n962 ;
  assign n964 = n963 ^ n148 ^ 1'b0 ;
  assign n965 = ( n415 & ~n593 ) | ( n415 & n964 ) | ( ~n593 & n964 ) ;
  assign n966 = n591 | n622 ;
  assign n967 = n966 ^ n527 ^ 1'b0 ;
  assign n970 = n380 | n637 ;
  assign n968 = x47 & ~n591 ;
  assign n969 = n968 ^ n759 ^ 1'b0 ;
  assign n971 = n970 ^ n969 ^ x50 ;
  assign n972 = n872 ^ n395 ^ x66 ;
  assign n973 = n378 ^ n323 ^ n150 ;
  assign n974 = n972 | n973 ;
  assign n975 = n230 ^ n148 ^ x38 ;
  assign n976 = n975 ^ n890 ^ 1'b0 ;
  assign n977 = x27 & x31 ;
  assign n978 = n977 ^ n164 ^ 1'b0 ;
  assign n979 = n764 ^ n292 ^ 1'b0 ;
  assign n980 = n978 | n979 ;
  assign n981 = n545 ^ n248 ^ 1'b0 ;
  assign n982 = n187 ^ n171 ^ 1'b0 ;
  assign n983 = n981 | n982 ;
  assign n984 = n427 ^ n206 ^ 1'b0 ;
  assign n985 = n984 ^ n861 ^ n297 ;
  assign n986 = ( ~n345 & n983 ) | ( ~n345 & n985 ) | ( n983 & n985 ) ;
  assign n987 = n323 ^ n163 ^ 1'b0 ;
  assign n988 = n180 | n987 ;
  assign n989 = n988 ^ n636 ^ 1'b0 ;
  assign n990 = n524 | n989 ;
  assign n991 = n667 ^ n279 ^ n141 ;
  assign n992 = ( x81 & ~n407 ) | ( x81 & n695 ) | ( ~n407 & n695 ) ;
  assign n993 = n991 | n992 ;
  assign n994 = n367 & ~n993 ;
  assign n995 = ( x23 & n657 ) | ( x23 & ~n994 ) | ( n657 & ~n994 ) ;
  assign n996 = n995 ^ n273 ^ 1'b0 ;
  assign n997 = n996 ^ n754 ^ n680 ;
  assign n998 = n985 ^ n219 ^ 1'b0 ;
  assign n999 = n589 ^ n323 ^ 1'b0 ;
  assign n1000 = n259 & ~n999 ;
  assign n1001 = n1000 ^ n973 ^ 1'b0 ;
  assign n1002 = n293 ^ n236 ^ n218 ;
  assign n1003 = ( ~n466 & n525 ) | ( ~n466 & n1002 ) | ( n525 & n1002 ) ;
  assign n1004 = ( ~n750 & n974 ) | ( ~n750 & n1003 ) | ( n974 & n1003 ) ;
  assign n1005 = n350 ^ x106 ^ 1'b0 ;
  assign n1009 = n145 & n239 ;
  assign n1010 = n1009 ^ x94 ^ 1'b0 ;
  assign n1006 = x86 ^ x16 ^ 1'b0 ;
  assign n1007 = ( n395 & n504 ) | ( n395 & ~n599 ) | ( n504 & ~n599 ) ;
  assign n1008 = ( n168 & n1006 ) | ( n168 & n1007 ) | ( n1006 & n1007 ) ;
  assign n1011 = n1010 ^ n1008 ^ 1'b0 ;
  assign n1012 = n493 & ~n590 ;
  assign n1013 = ~n757 & n1012 ;
  assign n1014 = ~n1011 & n1013 ;
  assign n1015 = ( x123 & n270 ) | ( x123 & ~n1014 ) | ( n270 & ~n1014 ) ;
  assign n1016 = ( n486 & n519 ) | ( n486 & n680 ) | ( n519 & n680 ) ;
  assign n1017 = ( n374 & ~n595 ) | ( n374 & n1016 ) | ( ~n595 & n1016 ) ;
  assign n1018 = n934 ^ n316 ^ x110 ;
  assign n1019 = n1018 ^ n947 ^ x14 ;
  assign n1020 = n1019 ^ n1018 ^ n654 ;
  assign n1021 = ( n442 & n1017 ) | ( n442 & n1020 ) | ( n1017 & n1020 ) ;
  assign n1029 = n597 ^ n485 ^ n420 ;
  assign n1022 = ( ~x65 & x109 ) | ( ~x65 & n198 ) | ( x109 & n198 ) ;
  assign n1023 = ( x68 & n756 ) | ( x68 & ~n1022 ) | ( n756 & ~n1022 ) ;
  assign n1024 = n1023 ^ n322 ^ x17 ;
  assign n1025 = n1024 ^ n264 ^ x95 ;
  assign n1026 = ( n273 & ~n480 ) | ( n273 & n1025 ) | ( ~n480 & n1025 ) ;
  assign n1027 = n1026 ^ n901 ^ 1'b0 ;
  assign n1028 = x39 & ~n1027 ;
  assign n1030 = n1029 ^ n1028 ^ x43 ;
  assign n1031 = n182 & n490 ;
  assign n1032 = n1031 ^ n624 ^ 1'b0 ;
  assign n1033 = n370 & ~n520 ;
  assign n1034 = ~n758 & n1033 ;
  assign n1035 = x24 & ~n1034 ;
  assign n1036 = n1035 ^ n452 ^ 1'b0 ;
  assign n1037 = x10 & ~n414 ;
  assign n1038 = n203 & n1037 ;
  assign n1039 = n1036 & ~n1038 ;
  assign n1040 = x68 & n1039 ;
  assign n1041 = ( x60 & n182 ) | ( x60 & ~n880 ) | ( n182 & ~n880 ) ;
  assign n1042 = ~n743 & n1041 ;
  assign n1043 = n312 & n1042 ;
  assign n1044 = ( n198 & n888 ) | ( n198 & n1043 ) | ( n888 & n1043 ) ;
  assign n1045 = ~x121 & n317 ;
  assign n1046 = x85 & ~n1045 ;
  assign n1047 = n1046 ^ n359 ^ 1'b0 ;
  assign n1048 = x48 & n1047 ;
  assign n1049 = n1046 & n1048 ;
  assign n1050 = ( x37 & x110 ) | ( x37 & n853 ) | ( x110 & n853 ) ;
  assign n1051 = n1050 ^ n129 ^ x85 ;
  assign n1052 = n1051 ^ x112 ^ 1'b0 ;
  assign n1053 = n1052 ^ n733 ^ n525 ;
  assign n1054 = ~n540 & n1053 ;
  assign n1055 = n1054 ^ n787 ^ 1'b0 ;
  assign n1056 = n706 & n1055 ;
  assign n1057 = n850 & n1056 ;
  assign n1062 = n929 ^ n834 ^ 1'b0 ;
  assign n1058 = n989 ^ x102 ^ 1'b0 ;
  assign n1059 = ~n499 & n1058 ;
  assign n1060 = n542 & n1059 ;
  assign n1061 = n1060 ^ n307 ^ 1'b0 ;
  assign n1063 = n1062 ^ n1061 ^ n1059 ;
  assign n1069 = n978 ^ x50 ^ 1'b0 ;
  assign n1064 = x22 & n298 ;
  assign n1065 = n1064 ^ n172 ^ 1'b0 ;
  assign n1066 = n703 ^ n436 ^ x2 ;
  assign n1067 = ~x68 & n1066 ;
  assign n1068 = n1065 & n1067 ;
  assign n1070 = n1069 ^ n1068 ^ n549 ;
  assign n1071 = n1070 ^ n903 ^ n711 ;
  assign n1075 = x4 & ~n162 ;
  assign n1076 = ~n670 & n1075 ;
  assign n1077 = n300 | n1076 ;
  assign n1078 = x24 | n1077 ;
  assign n1072 = x101 & n223 ;
  assign n1073 = n1072 ^ n223 ^ 1'b0 ;
  assign n1074 = ( n348 & ~n540 ) | ( n348 & n1073 ) | ( ~n540 & n1073 ) ;
  assign n1079 = n1078 ^ n1074 ^ n991 ;
  assign n1080 = ~n402 & n1079 ;
  assign n1081 = n1080 ^ n342 ^ 1'b0 ;
  assign n1082 = ( ~x52 & n254 ) | ( ~x52 & n277 ) | ( n254 & n277 ) ;
  assign n1083 = n436 ^ n319 ^ x67 ;
  assign n1084 = n492 ^ x82 ^ 1'b0 ;
  assign n1085 = ( n307 & n324 ) | ( n307 & n1084 ) | ( n324 & n1084 ) ;
  assign n1086 = ( n539 & n1083 ) | ( n539 & n1085 ) | ( n1083 & n1085 ) ;
  assign n1087 = n890 ^ n165 ^ 1'b0 ;
  assign n1088 = ~n170 & n1087 ;
  assign n1089 = ~n981 & n1088 ;
  assign n1090 = ~n1086 & n1089 ;
  assign n1091 = ( n780 & n1082 ) | ( n780 & n1090 ) | ( n1082 & n1090 ) ;
  assign n1092 = x37 & ~n1091 ;
  assign n1093 = n1081 & n1092 ;
  assign n1094 = n236 | n1093 ;
  assign n1095 = n1050 | n1094 ;
  assign n1096 = n713 ^ n302 ^ x76 ;
  assign n1097 = n178 & ~n565 ;
  assign n1098 = n1097 ^ n413 ^ n233 ;
  assign n1099 = ( n786 & ~n1096 ) | ( n786 & n1098 ) | ( ~n1096 & n1098 ) ;
  assign n1100 = ( x53 & n412 ) | ( x53 & ~n806 ) | ( n412 & ~n806 ) ;
  assign n1101 = n923 ^ n215 ^ 1'b0 ;
  assign n1102 = x73 & n1101 ;
  assign n1103 = n984 ^ n956 ^ 1'b0 ;
  assign n1104 = n1102 & ~n1103 ;
  assign n1105 = x60 & n414 ;
  assign n1106 = n1105 ^ n187 ^ 1'b0 ;
  assign n1107 = ( x7 & n764 ) | ( x7 & n866 ) | ( n764 & n866 ) ;
  assign n1108 = ~n391 & n750 ;
  assign n1109 = x65 & n1108 ;
  assign n1110 = n788 | n1109 ;
  assign n1111 = n1107 & ~n1110 ;
  assign n1112 = n466 | n794 ;
  assign n1113 = ( n716 & n1079 ) | ( n716 & n1112 ) | ( n1079 & n1112 ) ;
  assign n1114 = ( ~n197 & n1093 ) | ( ~n197 & n1113 ) | ( n1093 & n1113 ) ;
  assign n1115 = n635 ^ n580 ^ n134 ;
  assign n1118 = ( x37 & n265 ) | ( x37 & ~n285 ) | ( n265 & ~n285 ) ;
  assign n1116 = x74 & x77 ;
  assign n1117 = n1116 ^ n326 ^ 1'b0 ;
  assign n1119 = n1118 ^ n1117 ^ n545 ;
  assign n1120 = n1119 ^ n217 ^ 1'b0 ;
  assign n1125 = ~n165 & n350 ;
  assign n1121 = n198 & n394 ;
  assign n1122 = n1121 ^ x114 ^ 1'b0 ;
  assign n1123 = ( ~x10 & n141 ) | ( ~x10 & n1122 ) | ( n141 & n1122 ) ;
  assign n1124 = n1123 ^ n337 ^ 1'b0 ;
  assign n1126 = n1125 ^ n1124 ^ n194 ;
  assign n1127 = n1036 ^ n802 ^ n360 ;
  assign n1128 = n133 & ~n436 ;
  assign n1129 = ( x23 & x66 ) | ( x23 & ~n1128 ) | ( x66 & ~n1128 ) ;
  assign n1130 = ( ~n239 & n253 ) | ( ~n239 & n1129 ) | ( n253 & n1129 ) ;
  assign n1132 = ( n142 & ~n265 ) | ( n142 & n291 ) | ( ~n265 & n291 ) ;
  assign n1133 = x9 & ~n325 ;
  assign n1134 = n235 & n1133 ;
  assign n1135 = ~n1083 & n1134 ;
  assign n1136 = n1132 & n1135 ;
  assign n1131 = n194 & ~n544 ;
  assign n1137 = n1136 ^ n1131 ^ 1'b0 ;
  assign n1138 = n1066 & n1137 ;
  assign n1139 = ~x39 & n1138 ;
  assign n1140 = x126 & ~n1118 ;
  assign n1141 = ~n242 & n1140 ;
  assign n1142 = n1141 ^ n859 ^ x108 ;
  assign n1147 = n490 & ~n500 ;
  assign n1145 = n1045 ^ n242 ^ n141 ;
  assign n1146 = n1145 ^ n145 ^ 1'b0 ;
  assign n1143 = n1023 ^ n978 ^ n690 ;
  assign n1144 = n1143 ^ n673 ^ 1'b0 ;
  assign n1148 = n1147 ^ n1146 ^ n1144 ;
  assign n1149 = ( n912 & ~n1017 ) | ( n912 & n1124 ) | ( ~n1017 & n1124 ) ;
  assign n1150 = n1149 ^ n1002 ^ x54 ;
  assign n1152 = n662 ^ n595 ^ n315 ;
  assign n1151 = n617 | n931 ;
  assign n1153 = n1152 ^ n1151 ^ n599 ;
  assign n1154 = n225 ^ n156 ^ x23 ;
  assign n1155 = n1154 ^ n573 ^ x127 ;
  assign n1156 = n643 & n1155 ;
  assign n1157 = n699 & n1156 ;
  assign n1158 = ( ~x123 & n380 ) | ( ~x123 & n1088 ) | ( n380 & n1088 ) ;
  assign n1159 = ( n316 & ~n730 ) | ( n316 & n1006 ) | ( ~n730 & n1006 ) ;
  assign n1160 = n213 & n1159 ;
  assign n1162 = n167 & n653 ;
  assign n1163 = n1162 ^ x113 ^ 1'b0 ;
  assign n1161 = n183 & ~n302 ;
  assign n1164 = n1163 ^ n1161 ^ 1'b0 ;
  assign n1165 = ~n591 & n1164 ;
  assign n1166 = n1160 & n1165 ;
  assign n1167 = n1158 | n1166 ;
  assign n1168 = n509 | n1167 ;
  assign n1171 = n1016 ^ x28 ^ x13 ;
  assign n1169 = ( n330 & ~n395 ) | ( n330 & n407 ) | ( ~n395 & n407 ) ;
  assign n1170 = n579 & n1169 ;
  assign n1172 = n1171 ^ n1170 ^ n759 ;
  assign n1173 = n158 & n1172 ;
  assign n1174 = n1020 & n1173 ;
  assign n1175 = n166 ^ n153 ^ x26 ;
  assign n1176 = n1175 ^ n1068 ^ n597 ;
  assign n1177 = n1176 ^ n839 ^ x57 ;
  assign n1182 = ( ~x74 & n229 ) | ( ~x74 & n750 ) | ( n229 & n750 ) ;
  assign n1178 = n869 & ~n1065 ;
  assign n1179 = n1178 ^ n1074 ^ 1'b0 ;
  assign n1180 = n429 & n943 ;
  assign n1181 = ~n1179 & n1180 ;
  assign n1183 = n1182 ^ n1181 ^ 1'b0 ;
  assign n1190 = ( x87 & ~n171 ) | ( x87 & n385 ) | ( ~n171 & n385 ) ;
  assign n1188 = ( ~n547 & n561 ) | ( ~n547 & n911 ) | ( n561 & n911 ) ;
  assign n1184 = ~n597 & n706 ;
  assign n1185 = n816 ^ n155 ^ 1'b0 ;
  assign n1186 = n717 & n1185 ;
  assign n1187 = ~n1184 & n1186 ;
  assign n1189 = n1188 ^ n1187 ^ 1'b0 ;
  assign n1191 = n1190 ^ n1189 ^ n1182 ;
  assign n1192 = ( x23 & n236 ) | ( x23 & n550 ) | ( n236 & n550 ) ;
  assign n1193 = n1192 ^ n184 ^ 1'b0 ;
  assign n1202 = n719 ^ n626 ^ 1'b0 ;
  assign n1203 = n449 | n1202 ;
  assign n1204 = n884 & ~n1203 ;
  assign n1194 = ( n242 & n437 ) | ( n242 & ~n492 ) | ( n437 & ~n492 ) ;
  assign n1195 = ~n477 & n1194 ;
  assign n1196 = n1043 & n1195 ;
  assign n1197 = ( ~n555 & n823 ) | ( ~n555 & n898 ) | ( n823 & n898 ) ;
  assign n1198 = n1197 ^ n1171 ^ 1'b0 ;
  assign n1199 = n1006 & n1198 ;
  assign n1200 = ( n376 & n481 ) | ( n376 & n1199 ) | ( n481 & n1199 ) ;
  assign n1201 = n1196 | n1200 ;
  assign n1205 = n1204 ^ n1201 ^ 1'b0 ;
  assign n1206 = n1154 ^ n340 ^ x61 ;
  assign n1207 = n667 ^ n601 ^ 1'b0 ;
  assign n1208 = x89 & ~n1207 ;
  assign n1209 = n732 & ~n1208 ;
  assign n1210 = ( ~n207 & n270 ) | ( ~n207 & n292 ) | ( n270 & n292 ) ;
  assign n1211 = n421 & ~n590 ;
  assign n1212 = n1211 ^ n973 ^ 1'b0 ;
  assign n1213 = ( n1169 & n1210 ) | ( n1169 & ~n1212 ) | ( n1210 & ~n1212 ) ;
  assign n1214 = ( ~n1203 & n1209 ) | ( ~n1203 & n1213 ) | ( n1209 & n1213 ) ;
  assign n1218 = n863 ^ n512 ^ 1'b0 ;
  assign n1219 = n856 & n1218 ;
  assign n1215 = n397 & n628 ;
  assign n1216 = n270 & n1215 ;
  assign n1217 = ~n375 & n1216 ;
  assign n1220 = n1219 ^ n1217 ^ n390 ;
  assign n1221 = n1220 ^ n1049 ^ 1'b0 ;
  assign n1224 = n134 | n592 ;
  assign n1225 = n1224 ^ x108 ^ 1'b0 ;
  assign n1223 = x81 & ~n180 ;
  assign n1226 = n1225 ^ n1223 ^ 1'b0 ;
  assign n1222 = n381 | n1020 ;
  assign n1227 = n1226 ^ n1222 ^ 1'b0 ;
  assign n1228 = ( x24 & n174 ) | ( x24 & ~n607 ) | ( n174 & ~n607 ) ;
  assign n1230 = x80 & n960 ;
  assign n1231 = n1230 ^ n295 ^ 1'b0 ;
  assign n1229 = x97 & n1149 ;
  assign n1232 = n1231 ^ n1229 ^ 1'b0 ;
  assign n1233 = ( n298 & n1228 ) | ( n298 & n1232 ) | ( n1228 & n1232 ) ;
  assign n1234 = n145 & n302 ;
  assign n1235 = ( x86 & ~n1216 ) | ( x86 & n1234 ) | ( ~n1216 & n1234 ) ;
  assign n1236 = n401 & ~n1068 ;
  assign n1237 = n1236 ^ n583 ^ 1'b0 ;
  assign n1238 = n453 & n1219 ;
  assign n1239 = n1203 & n1238 ;
  assign n1240 = n215 & ~n713 ;
  assign n1241 = n1240 ^ n252 ^ 1'b0 ;
  assign n1242 = n556 | n1241 ;
  assign n1243 = n934 ^ n445 ^ 1'b0 ;
  assign n1247 = n846 ^ n375 ^ 1'b0 ;
  assign n1248 = ( ~n186 & n646 ) | ( ~n186 & n1247 ) | ( n646 & n1247 ) ;
  assign n1244 = ( n315 & n360 ) | ( n315 & ~n853 ) | ( n360 & ~n853 ) ;
  assign n1245 = n921 ^ n847 ^ 1'b0 ;
  assign n1246 = n1244 & ~n1245 ;
  assign n1249 = n1248 ^ n1246 ^ 1'b0 ;
  assign n1250 = ~n849 & n1249 ;
  assign n1251 = n1250 ^ n1005 ^ n984 ;
  assign n1252 = ~n270 & n1247 ;
  assign n1253 = ~n1251 & n1252 ;
  assign n1254 = n166 ^ x47 ^ 1'b0 ;
  assign n1255 = x15 & n1254 ;
  assign n1256 = n883 ^ n520 ^ 1'b0 ;
  assign n1257 = n434 & ~n1256 ;
  assign n1258 = ~n1212 & n1257 ;
  assign n1259 = ~n1255 & n1258 ;
  assign n1260 = n549 ^ x64 ^ 1'b0 ;
  assign n1261 = n1260 ^ n317 ^ x124 ;
  assign n1262 = ( ~n307 & n1259 ) | ( ~n307 & n1261 ) | ( n1259 & n1261 ) ;
  assign n1263 = ( n145 & n304 ) | ( n145 & ~n355 ) | ( n304 & ~n355 ) ;
  assign n1264 = ( x64 & ~n741 ) | ( x64 & n1263 ) | ( ~n741 & n1263 ) ;
  assign n1265 = ~x3 & n720 ;
  assign n1266 = ( n288 & ~n1095 ) | ( n288 & n1265 ) | ( ~n1095 & n1265 ) ;
  assign n1267 = ~n508 & n751 ;
  assign n1268 = n1267 ^ n434 ^ 1'b0 ;
  assign n1269 = ( n189 & n370 ) | ( n189 & ~n474 ) | ( n370 & ~n474 ) ;
  assign n1270 = ( n195 & n645 ) | ( n195 & ~n786 ) | ( n645 & ~n786 ) ;
  assign n1271 = ~n471 & n1145 ;
  assign n1272 = n426 & n1271 ;
  assign n1273 = ( n492 & n1270 ) | ( n492 & n1272 ) | ( n1270 & n1272 ) ;
  assign n1274 = n1273 ^ n1008 ^ 1'b0 ;
  assign n1275 = n1269 & ~n1274 ;
  assign n1276 = ( n1150 & n1268 ) | ( n1150 & n1275 ) | ( n1268 & n1275 ) ;
  assign n1279 = ( n263 & ~n284 ) | ( n263 & n604 ) | ( ~n284 & n604 ) ;
  assign n1280 = x66 ^ x23 ^ 1'b0 ;
  assign n1281 = ( n782 & n1279 ) | ( n782 & ~n1280 ) | ( n1279 & ~n1280 ) ;
  assign n1282 = n1281 ^ n503 ^ x17 ;
  assign n1277 = n632 ^ n500 ^ 1'b0 ;
  assign n1278 = n445 & ~n1277 ;
  assign n1283 = n1282 ^ n1278 ^ 1'b0 ;
  assign n1284 = n806 & n975 ;
  assign n1287 = n207 & ~n551 ;
  assign n1285 = ( x73 & x88 ) | ( x73 & ~n607 ) | ( x88 & ~n607 ) ;
  assign n1286 = n1285 ^ n738 ^ n432 ;
  assign n1288 = n1287 ^ n1286 ^ 1'b0 ;
  assign n1289 = n1106 ^ n876 ^ n433 ;
  assign n1292 = x32 & n748 ;
  assign n1290 = ( x40 & ~x58 ) | ( x40 & n1002 ) | ( ~x58 & n1002 ) ;
  assign n1291 = n598 & n1290 ;
  assign n1293 = n1292 ^ n1291 ^ n643 ;
  assign n1294 = ~n203 & n445 ;
  assign n1295 = ( n160 & n185 ) | ( n160 & n1294 ) | ( n185 & n1294 ) ;
  assign n1296 = ( ~n730 & n1293 ) | ( ~n730 & n1295 ) | ( n1293 & n1295 ) ;
  assign n1297 = x124 & ~n129 ;
  assign n1298 = ( ~n831 & n1025 ) | ( ~n831 & n1297 ) | ( n1025 & n1297 ) ;
  assign n1299 = n1298 ^ n1036 ^ x51 ;
  assign n1300 = n145 & n206 ;
  assign n1301 = n555 ^ n214 ^ x39 ;
  assign n1302 = n1300 | n1301 ;
  assign n1303 = n1299 | n1302 ;
  assign n1304 = ( x49 & n573 ) | ( x49 & ~n1303 ) | ( n573 & ~n1303 ) ;
  assign n1305 = ( x56 & n1117 ) | ( x56 & n1304 ) | ( n1117 & n1304 ) ;
  assign n1306 = n1305 ^ n1242 ^ 1'b0 ;
  assign n1309 = n1123 ^ n176 ^ 1'b0 ;
  assign n1310 = n834 | n1309 ;
  assign n1311 = ( x33 & n236 ) | ( x33 & ~n1310 ) | ( n236 & ~n1310 ) ;
  assign n1307 = n951 ^ n787 ^ n179 ;
  assign n1308 = n1307 ^ n1108 ^ 1'b0 ;
  assign n1312 = n1311 ^ n1308 ^ n1065 ;
  assign n1313 = n1312 ^ n916 ^ n298 ;
  assign n1314 = n1284 ^ n991 ^ x116 ;
  assign n1315 = n1034 ^ n892 ^ n725 ;
  assign n1316 = n531 ^ n309 ^ 1'b0 ;
  assign n1317 = ( n568 & n653 ) | ( n568 & n1316 ) | ( n653 & n1316 ) ;
  assign n1318 = ( x9 & n1315 ) | ( x9 & n1317 ) | ( n1315 & n1317 ) ;
  assign n1323 = n719 ^ n656 ^ 1'b0 ;
  assign n1319 = n854 ^ n590 ^ 1'b0 ;
  assign n1320 = x57 & ~n1319 ;
  assign n1321 = n1320 ^ n485 ^ 1'b0 ;
  assign n1322 = n892 & n1321 ;
  assign n1324 = n1323 ^ n1322 ^ n234 ;
  assign n1325 = n732 ^ n238 ^ 1'b0 ;
  assign n1326 = n673 | n1325 ;
  assign n1338 = n989 ^ n988 ^ n359 ;
  assign n1337 = n369 & ~n1228 ;
  assign n1339 = n1338 ^ n1337 ^ 1'b0 ;
  assign n1333 = n170 ^ n161 ^ 1'b0 ;
  assign n1334 = n130 & ~n1333 ;
  assign n1332 = n277 & ~n486 ;
  assign n1335 = n1334 ^ n1332 ^ n716 ;
  assign n1336 = ( n757 & n1074 ) | ( n757 & n1335 ) | ( n1074 & n1335 ) ;
  assign n1327 = ( x2 & n717 ) | ( x2 & ~n863 ) | ( n717 & ~n863 ) ;
  assign n1328 = ~n505 & n1327 ;
  assign n1329 = n1328 ^ n782 ^ 1'b0 ;
  assign n1330 = n1329 ^ n1084 ^ n1069 ;
  assign n1331 = n167 & n1330 ;
  assign n1340 = n1339 ^ n1336 ^ n1331 ;
  assign n1341 = n366 ^ x68 ^ 1'b0 ;
  assign n1343 = x39 | n813 ;
  assign n1342 = n771 ^ n265 ^ 1'b0 ;
  assign n1344 = n1343 ^ n1342 ^ n178 ;
  assign n1345 = n1012 & n1344 ;
  assign n1346 = n1345 ^ n836 ^ 1'b0 ;
  assign n1348 = n1041 ^ n159 ^ x75 ;
  assign n1347 = ~n359 & n437 ;
  assign n1349 = n1348 ^ n1347 ^ n179 ;
  assign n1350 = n385 ^ n310 ^ n213 ;
  assign n1351 = n1350 ^ n633 ^ 1'b0 ;
  assign n1352 = n222 & n1322 ;
  assign n1353 = ~n1351 & n1352 ;
  assign n1354 = x2 & ~x88 ;
  assign n1355 = n359 ^ x115 ^ 1'b0 ;
  assign n1356 = n1355 ^ n207 ^ n143 ;
  assign n1357 = n1356 ^ n1297 ^ n957 ;
  assign n1358 = n853 & n1357 ;
  assign n1359 = n1358 ^ n1297 ^ n335 ;
  assign n1368 = ( x52 & ~n256 ) | ( x52 & n435 ) | ( ~n256 & n435 ) ;
  assign n1360 = ( ~x4 & n220 ) | ( ~x4 & n432 ) | ( n220 & n432 ) ;
  assign n1361 = n1360 ^ n821 ^ n142 ;
  assign n1362 = ( n166 & n330 ) | ( n166 & n1361 ) | ( n330 & n1361 ) ;
  assign n1363 = x3 & n166 ;
  assign n1364 = n1363 ^ n709 ^ 1'b0 ;
  assign n1365 = x63 & n1364 ;
  assign n1366 = ~n1362 & n1365 ;
  assign n1367 = n1076 | n1366 ;
  assign n1369 = n1368 ^ n1367 ^ 1'b0 ;
  assign n1370 = ~x10 & x33 ;
  assign n1371 = n1123 & ~n1370 ;
  assign n1372 = n1371 ^ n949 ^ 1'b0 ;
  assign n1373 = ~n743 & n1372 ;
  assign n1374 = x120 | n673 ;
  assign n1375 = n972 ^ n178 ^ x53 ;
  assign n1376 = ( n305 & ~n1374 ) | ( n305 & n1375 ) | ( ~n1374 & n1375 ) ;
  assign n1377 = n408 ^ x90 ^ 1'b0 ;
  assign n1378 = n1376 | n1377 ;
  assign n1379 = ( ~n503 & n648 ) | ( ~n503 & n842 ) | ( n648 & n842 ) ;
  assign n1380 = ( n500 & ~n974 ) | ( n500 & n1379 ) | ( ~n974 & n1379 ) ;
  assign n1381 = n853 ^ n492 ^ x101 ;
  assign n1382 = n595 | n1381 ;
  assign n1383 = n568 ^ n429 ^ 1'b0 ;
  assign n1384 = n1287 & n1383 ;
  assign n1385 = n1384 ^ n242 ^ 1'b0 ;
  assign n1386 = ~n226 & n1385 ;
  assign n1387 = ( x67 & n375 ) | ( x67 & n663 ) | ( n375 & n663 ) ;
  assign n1388 = n1387 ^ n1017 ^ n732 ;
  assign n1389 = n1349 & ~n1388 ;
  assign n1390 = ~n1386 & n1389 ;
  assign n1391 = ( x24 & n295 ) | ( x24 & ~n1006 ) | ( n295 & ~n1006 ) ;
  assign n1392 = ( n1192 & n1197 ) | ( n1192 & ~n1391 ) | ( n1197 & ~n1391 ) ;
  assign n1393 = ( x123 & n367 ) | ( x123 & n1392 ) | ( n367 & n1392 ) ;
  assign n1394 = n1393 ^ n863 ^ 1'b0 ;
  assign n1395 = n1247 ^ n366 ^ 1'b0 ;
  assign n1396 = n884 ^ n513 ^ 1'b0 ;
  assign n1397 = x50 & n840 ;
  assign n1398 = n168 ^ x50 ^ 1'b0 ;
  assign n1399 = x42 & ~n1398 ;
  assign n1400 = n1399 ^ x123 ^ 1'b0 ;
  assign n1401 = n328 | n1400 ;
  assign n1402 = n184 & n372 ;
  assign n1403 = n1402 ^ n217 ^ 1'b0 ;
  assign n1404 = ( n1297 & n1316 ) | ( n1297 & ~n1403 ) | ( n1316 & ~n1403 ) ;
  assign n1405 = n525 & ~n1404 ;
  assign n1406 = n1108 ^ n519 ^ n190 ;
  assign n1407 = n1066 ^ n620 ^ n259 ;
  assign n1410 = n1096 ^ n415 ^ 1'b0 ;
  assign n1411 = n266 & ~n1410 ;
  assign n1408 = ( x25 & ~x77 ) | ( x25 & n706 ) | ( ~x77 & n706 ) ;
  assign n1409 = ( n166 & ~n257 ) | ( n166 & n1408 ) | ( ~n257 & n1408 ) ;
  assign n1412 = n1411 ^ n1409 ^ n1265 ;
  assign n1413 = ~n1407 & n1412 ;
  assign n1414 = n1413 ^ n287 ^ 1'b0 ;
  assign n1415 = n1112 ^ n181 ^ 1'b0 ;
  assign n1416 = n1392 | n1415 ;
  assign n1417 = n1357 & ~n1416 ;
  assign n1418 = n846 & n1417 ;
  assign n1419 = n674 ^ n428 ^ 1'b0 ;
  assign n1420 = n572 | n1419 ;
  assign n1421 = n1420 ^ n145 ^ 1'b0 ;
  assign n1422 = n1421 ^ n692 ^ n298 ;
  assign n1423 = n615 & n1299 ;
  assign n1424 = n1109 & n1423 ;
  assign n1425 = ( n943 & ~n1422 ) | ( n943 & n1424 ) | ( ~n1422 & n1424 ) ;
  assign n1426 = n1303 ^ n765 ^ n565 ;
  assign n1427 = ( n408 & ~n676 ) | ( n408 & n879 ) | ( ~n676 & n879 ) ;
  assign n1428 = n722 & n1427 ;
  assign n1429 = n1428 ^ x46 ^ 1'b0 ;
  assign n1430 = ~n937 & n1429 ;
  assign n1431 = ( n131 & n407 ) | ( n131 & ~n506 ) | ( n407 & ~n506 ) ;
  assign n1432 = ~n695 & n1147 ;
  assign n1433 = ( n697 & n1431 ) | ( n697 & n1432 ) | ( n1431 & n1432 ) ;
  assign n1434 = n282 ^ x37 ^ x21 ;
  assign n1435 = n409 & ~n517 ;
  assign n1436 = n1435 ^ x23 ^ 1'b0 ;
  assign n1437 = n441 ^ n143 ^ 1'b0 ;
  assign n1438 = n1436 | n1437 ;
  assign n1439 = n1438 ^ n849 ^ 1'b0 ;
  assign n1440 = n1434 | n1439 ;
  assign n1441 = n1440 ^ n998 ^ 1'b0 ;
  assign n1442 = ( ~n160 & n572 ) | ( ~n160 & n981 ) | ( n572 & n981 ) ;
  assign n1443 = n1184 ^ n874 ^ 1'b0 ;
  assign n1444 = n1443 ^ n130 ^ 1'b0 ;
  assign n1445 = n1130 ^ n677 ^ x6 ;
  assign n1446 = n1445 ^ n931 ^ 1'b0 ;
  assign n1447 = n1444 & n1446 ;
  assign n1448 = n786 ^ n456 ^ x125 ;
  assign n1449 = x41 & ~n1448 ;
  assign n1450 = ~n1050 & n1449 ;
  assign n1451 = n653 ^ x17 ^ x7 ;
  assign n1452 = n1451 ^ n322 ^ n201 ;
  assign n1453 = n792 ^ n137 ^ 1'b0 ;
  assign n1454 = ~n1452 & n1453 ;
  assign n1455 = ( n311 & ~n360 ) | ( n311 & n824 ) | ( ~n360 & n824 ) ;
  assign n1456 = n543 ^ n479 ^ n377 ;
  assign n1457 = ( n796 & ~n1455 ) | ( n796 & n1456 ) | ( ~n1455 & n1456 ) ;
  assign n1458 = n195 ^ x6 ^ 1'b0 ;
  assign n1459 = ~n142 & n1458 ;
  assign n1462 = n337 & n1022 ;
  assign n1463 = n1462 ^ n264 ^ 1'b0 ;
  assign n1464 = x123 & ~n131 ;
  assign n1465 = ~n1463 & n1464 ;
  assign n1460 = ( n896 & n996 ) | ( n896 & n1136 ) | ( n996 & n1136 ) ;
  assign n1461 = x103 & n1460 ;
  assign n1466 = n1465 ^ n1461 ^ 1'b0 ;
  assign n1467 = n853 | n1111 ;
  assign n1468 = n1467 ^ n345 ^ 1'b0 ;
  assign n1469 = n260 ^ x121 ^ 1'b0 ;
  assign n1470 = n654 & n1469 ;
  assign n1471 = n1470 ^ n1053 ^ x72 ;
  assign n1472 = ( ~x11 & n392 ) | ( ~x11 & n413 ) | ( n392 & n413 ) ;
  assign n1473 = x26 & ~n1472 ;
  assign n1474 = ( x121 & n775 ) | ( x121 & ~n1473 ) | ( n775 & ~n1473 ) ;
  assign n1475 = ( n610 & ~n1471 ) | ( n610 & n1474 ) | ( ~n1471 & n1474 ) ;
  assign n1476 = ( n223 & n555 ) | ( n223 & n1475 ) | ( n555 & n1475 ) ;
  assign n1477 = n240 ^ x59 ^ x14 ;
  assign n1478 = n949 | n1477 ;
  assign n1479 = n1478 ^ n428 ^ 1'b0 ;
  assign n1482 = n758 ^ x72 ^ 1'b0 ;
  assign n1483 = n1046 & n1482 ;
  assign n1480 = n543 ^ n438 ^ x92 ;
  assign n1481 = n513 & n1480 ;
  assign n1484 = n1483 ^ n1481 ^ 1'b0 ;
  assign n1485 = n916 | n1484 ;
  assign n1488 = n1065 ^ n159 ^ x8 ;
  assign n1489 = ( x10 & ~n1403 ) | ( x10 & n1488 ) | ( ~n1403 & n1488 ) ;
  assign n1490 = n272 & ~n1489 ;
  assign n1491 = n688 & n1490 ;
  assign n1492 = n1491 ^ n499 ^ 1'b0 ;
  assign n1486 = ( n345 & n575 ) | ( n345 & ~n612 ) | ( n575 & ~n612 ) ;
  assign n1487 = n694 | n1486 ;
  assign n1493 = n1492 ^ n1487 ^ 1'b0 ;
  assign n1494 = n1022 ^ n184 ^ 1'b0 ;
  assign n1495 = n881 ^ n858 ^ 1'b0 ;
  assign n1496 = n1494 & n1495 ;
  assign n1497 = n1496 ^ n912 ^ n248 ;
  assign n1498 = ( ~n703 & n1052 ) | ( ~n703 & n1497 ) | ( n1052 & n1497 ) ;
  assign n1499 = n975 | n1498 ;
  assign n1500 = n1499 ^ n909 ^ 1'b0 ;
  assign n1501 = n1068 ^ n437 ^ x99 ;
  assign n1502 = ~n162 & n1403 ;
  assign n1503 = ~n1501 & n1502 ;
  assign n1504 = ~n719 & n1068 ;
  assign n1505 = n549 & ~n765 ;
  assign n1506 = n1505 ^ n846 ^ 1'b0 ;
  assign n1507 = ( n757 & n1504 ) | ( n757 & n1506 ) | ( n1504 & n1506 ) ;
  assign n1508 = ( n412 & n1503 ) | ( n412 & n1507 ) | ( n1503 & n1507 ) ;
  assign n1513 = n901 ^ n665 ^ n294 ;
  assign n1514 = n1513 ^ n155 ^ 1'b0 ;
  assign n1510 = x17 & n279 ;
  assign n1509 = ( ~n370 & n506 ) | ( ~n370 & n962 ) | ( n506 & n962 ) ;
  assign n1511 = n1510 ^ n1509 ^ n527 ;
  assign n1512 = x71 & n1511 ;
  assign n1515 = n1514 ^ n1512 ^ 1'b0 ;
  assign n1516 = ( n166 & n213 ) | ( n166 & ~n978 ) | ( n213 & ~n978 ) ;
  assign n1517 = n744 ^ n685 ^ x36 ;
  assign n1518 = ( ~n1048 & n1516 ) | ( ~n1048 & n1517 ) | ( n1516 & n1517 ) ;
  assign n1519 = x87 & ~n1096 ;
  assign n1520 = n836 & ~n1519 ;
  assign n1521 = n1520 ^ n522 ^ 1'b0 ;
  assign n1522 = n1521 ^ n248 ^ x97 ;
  assign n1523 = n831 ^ n493 ^ n324 ;
  assign n1524 = n1523 ^ x2 ^ 1'b0 ;
  assign n1525 = n644 | n712 ;
  assign n1526 = n1525 ^ n1448 ^ n385 ;
  assign n1527 = n1526 ^ n1370 ^ 1'b0 ;
  assign n1528 = ~n1286 & n1527 ;
  assign n1529 = n1528 ^ n427 ^ n312 ;
  assign n1530 = n218 ^ x120 ^ x21 ;
  assign n1531 = n1530 ^ n844 ^ n626 ;
  assign n1532 = n1219 ^ n499 ^ 1'b0 ;
  assign n1533 = n1531 | n1532 ;
  assign n1534 = ( n711 & n863 ) | ( n711 & n1533 ) | ( n863 & n1533 ) ;
  assign n1540 = x34 & ~n680 ;
  assign n1541 = ~n292 & n1540 ;
  assign n1537 = n575 ^ n559 ^ 1'b0 ;
  assign n1538 = n391 & n1537 ;
  assign n1539 = ( x97 & n706 ) | ( x97 & ~n1538 ) | ( n706 & ~n1538 ) ;
  assign n1542 = n1541 ^ n1539 ^ 1'b0 ;
  assign n1543 = n338 & ~n1542 ;
  assign n1535 = n893 ^ n418 ^ 1'b0 ;
  assign n1536 = n760 & ~n1535 ;
  assign n1544 = n1543 ^ n1536 ^ n853 ;
  assign n1546 = n744 ^ n376 ^ 1'b0 ;
  assign n1547 = ~n162 & n1546 ;
  assign n1545 = x100 & ~n970 ;
  assign n1548 = n1547 ^ n1545 ^ 1'b0 ;
  assign n1549 = n1548 ^ x44 ^ 1'b0 ;
  assign n1550 = n700 & ~n1549 ;
  assign n1551 = ( n1154 & ~n1273 ) | ( n1154 & n1550 ) | ( ~n1273 & n1550 ) ;
  assign n1554 = n316 ^ x70 ^ x37 ;
  assign n1553 = n399 & n413 ;
  assign n1552 = ~n130 & n295 ;
  assign n1555 = n1554 ^ n1553 ^ n1552 ;
  assign n1557 = ( n375 & n665 ) | ( n375 & n1066 ) | ( n665 & n1066 ) ;
  assign n1556 = n903 | n1366 ;
  assign n1558 = n1557 ^ n1556 ^ 1'b0 ;
  assign n1559 = ( x117 & n1171 ) | ( x117 & ~n1558 ) | ( n1171 & ~n1558 ) ;
  assign n1560 = n466 ^ n143 ^ 1'b0 ;
  assign n1561 = x109 & n1560 ;
  assign n1562 = n1561 ^ n513 ^ 1'b0 ;
  assign n1563 = ~n1452 & n1562 ;
  assign n1564 = x55 & n509 ;
  assign n1565 = n465 & n1564 ;
  assign n1566 = n1565 ^ n646 ^ 1'b0 ;
  assign n1567 = n1371 ^ n1257 ^ n754 ;
  assign n1568 = n373 & ~n1007 ;
  assign n1569 = n695 | n1515 ;
  assign n1570 = n1568 | n1569 ;
  assign n1571 = n1280 ^ n1171 ^ n481 ;
  assign n1572 = n1117 ^ n602 ^ x82 ;
  assign n1574 = n1297 ^ n667 ^ n572 ;
  assign n1573 = ( ~x65 & n223 ) | ( ~x65 & n1279 ) | ( n223 & n1279 ) ;
  assign n1575 = n1574 ^ n1573 ^ n570 ;
  assign n1576 = n295 & ~n553 ;
  assign n1577 = n1575 & n1576 ;
  assign n1578 = ( n248 & ~n1572 ) | ( n248 & n1577 ) | ( ~n1572 & n1577 ) ;
  assign n1579 = n611 ^ x71 ^ 1'b0 ;
  assign n1580 = ~n1578 & n1579 ;
  assign n1581 = n512 & n1580 ;
  assign n1582 = ~x20 & n1581 ;
  assign n1583 = n1403 ^ n643 ^ n307 ;
  assign n1584 = ( ~n217 & n1068 ) | ( ~n217 & n1496 ) | ( n1068 & n1496 ) ;
  assign n1585 = ( x110 & n1055 ) | ( x110 & n1174 ) | ( n1055 & n1174 ) ;
  assign n1586 = ( n1583 & ~n1584 ) | ( n1583 & n1585 ) | ( ~n1584 & n1585 ) ;
  assign n1587 = n215 | n582 ;
  assign n1588 = n1587 ^ n1005 ^ 1'b0 ;
  assign n1589 = ( n670 & n1132 ) | ( n670 & n1588 ) | ( n1132 & n1588 ) ;
  assign n1590 = n273 & ~n1083 ;
  assign n1591 = n420 ^ n192 ^ 1'b0 ;
  assign n1592 = ~n230 & n1591 ;
  assign n1593 = ( ~n771 & n900 ) | ( ~n771 & n1592 ) | ( n900 & n1592 ) ;
  assign n1594 = n633 ^ n616 ^ n479 ;
  assign n1595 = x20 & n1594 ;
  assign n1596 = n1199 & ~n1595 ;
  assign n1597 = n822 & n1596 ;
  assign n1599 = n1347 ^ n617 ^ 1'b0 ;
  assign n1598 = n620 & n880 ;
  assign n1600 = n1599 ^ n1598 ^ 1'b0 ;
  assign n1607 = n1279 ^ n1016 ^ 1'b0 ;
  assign n1608 = n151 & ~n1607 ;
  assign n1609 = n740 ^ n432 ^ 1'b0 ;
  assign n1610 = ( n726 & n1608 ) | ( n726 & n1609 ) | ( n1608 & n1609 ) ;
  assign n1606 = ( ~n158 & n775 ) | ( ~n158 & n811 ) | ( n775 & n811 ) ;
  assign n1611 = n1610 ^ n1606 ^ n814 ;
  assign n1612 = n1611 ^ n831 ^ n163 ;
  assign n1601 = ( x116 & n488 ) | ( x116 & ~n1279 ) | ( n488 & ~n1279 ) ;
  assign n1602 = n1125 ^ n713 ^ 1'b0 ;
  assign n1603 = n1602 ^ n923 ^ 1'b0 ;
  assign n1604 = ~n1601 & n1603 ;
  assign n1605 = n1604 ^ n844 ^ 1'b0 ;
  assign n1613 = n1612 ^ n1605 ^ n570 ;
  assign n1614 = n1216 ^ n1129 ^ n794 ;
  assign n1615 = n1614 ^ x46 ^ 1'b0 ;
  assign n1616 = n415 | n1615 ;
  assign n1617 = n828 ^ n500 ^ n495 ;
  assign n1618 = n839 ^ n270 ^ x95 ;
  assign n1619 = n412 ^ n153 ^ x119 ;
  assign n1620 = ( n185 & n1583 ) | ( n185 & n1619 ) | ( n1583 & n1619 ) ;
  assign n1621 = ( ~x49 & n166 ) | ( ~x49 & n911 ) | ( n166 & n911 ) ;
  assign n1622 = ( n169 & n346 ) | ( n169 & n1621 ) | ( n346 & n1621 ) ;
  assign n1623 = ( n131 & n1620 ) | ( n131 & ~n1622 ) | ( n1620 & ~n1622 ) ;
  assign n1624 = ( x7 & n681 ) | ( x7 & ~n733 ) | ( n681 & ~n733 ) ;
  assign n1625 = n590 | n1624 ;
  assign n1626 = n1625 ^ n215 ^ 1'b0 ;
  assign n1627 = n1626 ^ n1160 ^ 1'b0 ;
  assign n1628 = n688 & ~n1627 ;
  assign n1629 = ( ~n169 & n1038 ) | ( ~n169 & n1244 ) | ( n1038 & n1244 ) ;
  assign n1630 = n1629 ^ n1017 ^ n810 ;
  assign n1631 = ( n1623 & n1628 ) | ( n1623 & ~n1630 ) | ( n1628 & ~n1630 ) ;
  assign n1632 = n220 ^ x9 ^ 1'b0 ;
  assign n1633 = x57 & n1632 ;
  assign n1634 = ~n1029 & n1633 ;
  assign n1635 = n1081 ^ n373 ^ x64 ;
  assign n1636 = n1635 ^ n401 ^ n217 ;
  assign n1637 = x107 & n683 ;
  assign n1638 = ~n428 & n1637 ;
  assign n1639 = n1638 ^ n1619 ^ n950 ;
  assign n1640 = n1639 ^ n1381 ^ 1'b0 ;
  assign n1641 = n1563 & n1640 ;
  assign n1646 = n343 ^ n236 ^ x92 ;
  assign n1644 = n1160 ^ n909 ^ 1'b0 ;
  assign n1642 = n506 & n611 ;
  assign n1643 = ~x86 & n1642 ;
  assign n1645 = n1644 ^ n1643 ^ x85 ;
  assign n1647 = n1646 ^ n1645 ^ n829 ;
  assign n1648 = n1647 ^ n612 ^ n431 ;
  assign n1649 = n490 & n508 ;
  assign n1650 = n1649 ^ n966 ^ n282 ;
  assign n1651 = n1650 ^ x60 ^ 1'b0 ;
  assign n1652 = n1102 ^ n479 ^ 1'b0 ;
  assign n1653 = x98 & ~n1652 ;
  assign n1654 = ( x65 & ~n1096 ) | ( x65 & n1653 ) | ( ~n1096 & n1653 ) ;
  assign n1655 = n1654 ^ n1053 ^ n978 ;
  assign n1656 = n1655 ^ n568 ^ n499 ;
  assign n1657 = ~n1651 & n1656 ;
  assign n1660 = ( x3 & x54 ) | ( x3 & ~n346 ) | ( x54 & ~n346 ) ;
  assign n1658 = n885 & n1610 ;
  assign n1659 = n1658 ^ n854 ^ 1'b0 ;
  assign n1661 = n1660 ^ n1659 ^ 1'b0 ;
  assign n1662 = n1480 | n1661 ;
  assign n1663 = x47 | n1662 ;
  assign n1664 = ( n219 & n374 ) | ( n219 & ~n642 ) | ( n374 & ~n642 ) ;
  assign n1665 = ( n653 & n1300 ) | ( n653 & n1664 ) | ( n1300 & n1664 ) ;
  assign n1666 = n1018 ^ n828 ^ n711 ;
  assign n1667 = ~n351 & n815 ;
  assign n1668 = ~n1074 & n1667 ;
  assign n1669 = x19 & n1668 ;
  assign n1670 = n1669 ^ n803 ^ 1'b0 ;
  assign n1671 = n1097 & ~n1670 ;
  assign n1672 = n1463 & n1671 ;
  assign n1674 = n246 ^ x2 ^ 1'b0 ;
  assign n1673 = n145 & ~n568 ;
  assign n1675 = n1674 ^ n1673 ^ 1'b0 ;
  assign n1676 = n434 ^ n156 ^ 1'b0 ;
  assign n1677 = ~n1675 & n1676 ;
  assign n1678 = n381 ^ n286 ^ 1'b0 ;
  assign n1679 = n1677 & n1678 ;
  assign n1680 = n1679 ^ n644 ^ 1'b0 ;
  assign n1681 = n1672 & n1680 ;
  assign n1682 = x125 & ~n1437 ;
  assign n1683 = ~n819 & n1682 ;
  assign n1684 = n1010 ^ x65 ^ 1'b0 ;
  assign n1685 = n1684 ^ n288 ^ 1'b0 ;
  assign n1686 = ~n1683 & n1685 ;
  assign n1687 = n1686 ^ x50 ^ 1'b0 ;
  assign n1688 = n292 & n935 ;
  assign n1689 = n1688 ^ n581 ^ 1'b0 ;
  assign n1690 = ~n1439 & n1689 ;
  assign n1691 = n1122 ^ n1036 ^ n230 ;
  assign n1692 = n393 & n996 ;
  assign n1693 = n1691 & n1692 ;
  assign n1694 = ( ~x61 & n1690 ) | ( ~x61 & n1693 ) | ( n1690 & n1693 ) ;
  assign n1695 = n512 & ~n1694 ;
  assign n1696 = x76 & n844 ;
  assign n1697 = ~n1695 & n1696 ;
  assign n1698 = ( x56 & ~x120 ) | ( x56 & n484 ) | ( ~x120 & n484 ) ;
  assign n1699 = ( x21 & n500 ) | ( x21 & ~n1698 ) | ( n500 & ~n1698 ) ;
  assign n1700 = ( x80 & ~n636 ) | ( x80 & n1062 ) | ( ~n636 & n1062 ) ;
  assign n1701 = n1643 ^ n641 ^ 1'b0 ;
  assign n1702 = x18 & ~n1701 ;
  assign n1703 = n1702 ^ n1674 ^ 1'b0 ;
  assign n1704 = ( ~x70 & n165 ) | ( ~x70 & n401 ) | ( n165 & n401 ) ;
  assign n1705 = n717 & ~n929 ;
  assign n1706 = n1705 ^ n748 ^ 1'b0 ;
  assign n1707 = n1706 ^ n869 ^ 1'b0 ;
  assign n1708 = n1707 ^ n1567 ^ n1565 ;
  assign n1709 = ( n374 & ~n615 ) | ( n374 & n621 ) | ( ~n615 & n621 ) ;
  assign n1710 = n1709 ^ n1362 ^ 1'b0 ;
  assign n1711 = n1532 | n1710 ;
  assign n1712 = n246 & n570 ;
  assign n1713 = n136 & n1712 ;
  assign n1714 = n1636 & ~n1713 ;
  assign n1715 = ( ~n187 & n450 ) | ( ~n187 & n905 ) | ( n450 & n905 ) ;
  assign n1716 = n1584 ^ n1129 ^ x102 ;
  assign n1717 = n1716 ^ n1384 ^ n897 ;
  assign n1718 = x117 | n1717 ;
  assign n1719 = n1644 ^ n994 ^ 1'b0 ;
  assign n1720 = n1719 ^ n1148 ^ n145 ;
  assign n1721 = n766 | n1070 ;
  assign n1722 = n1629 | n1721 ;
  assign n1723 = ~n802 & n1722 ;
  assign n1724 = n1723 ^ n1390 ^ 1'b0 ;
  assign n1725 = n654 ^ n223 ^ x67 ;
  assign n1726 = n1079 & ~n1725 ;
  assign n1727 = n541 & n1726 ;
  assign n1728 = ( ~x45 & x121 ) | ( ~x45 & n1727 ) | ( x121 & n1727 ) ;
  assign n1729 = ( n579 & ~n1616 ) | ( n579 & n1728 ) | ( ~n1616 & n1728 ) ;
  assign n1731 = n147 & ~n238 ;
  assign n1730 = ~n520 & n896 ;
  assign n1732 = n1731 ^ n1730 ^ 1'b0 ;
  assign n1733 = x116 & n1466 ;
  assign n1734 = ~x96 & n1733 ;
  assign n1735 = ~n159 & n357 ;
  assign n1736 = n235 & n1735 ;
  assign n1737 = n1379 ^ n610 ^ n510 ;
  assign n1738 = ( ~n760 & n1736 ) | ( ~n760 & n1737 ) | ( n1736 & n1737 ) ;
  assign n1739 = n1716 ^ n716 ^ 1'b0 ;
  assign n1740 = n764 ^ n625 ^ n505 ;
  assign n1741 = n1740 ^ n1548 ^ 1'b0 ;
  assign n1742 = n1741 ^ n1196 ^ 1'b0 ;
  assign n1743 = n418 ^ x23 ^ 1'b0 ;
  assign n1744 = x109 & ~n1743 ;
  assign n1745 = ( n167 & ~n365 ) | ( n167 & n465 ) | ( ~n365 & n465 ) ;
  assign n1746 = n1744 & ~n1745 ;
  assign n1747 = n265 & n1746 ;
  assign n1748 = n1213 ^ n857 ^ n788 ;
  assign n1749 = n609 ^ n325 ^ x75 ;
  assign n1750 = n1749 ^ n401 ^ x47 ;
  assign n1751 = ~n478 & n1550 ;
  assign n1752 = n1751 ^ n524 ^ 1'b0 ;
  assign n1753 = ~n362 & n1752 ;
  assign n1754 = n1750 & n1753 ;
  assign n1755 = ( x120 & ~n141 ) | ( x120 & n1436 ) | ( ~n141 & n1436 ) ;
  assign n1756 = n1755 ^ n1380 ^ 1'b0 ;
  assign n1757 = n978 ^ n803 ^ n453 ;
  assign n1758 = ( ~n515 & n1539 ) | ( ~n515 & n1757 ) | ( n1539 & n1757 ) ;
  assign n1759 = n547 ^ x46 ^ 1'b0 ;
  assign n1760 = n1759 ^ n1618 ^ 1'b0 ;
  assign n1761 = n1758 | n1760 ;
  assign n1762 = ( n1515 & n1756 ) | ( n1515 & ~n1761 ) | ( n1756 & ~n1761 ) ;
  assign n1763 = ( n847 & n1132 ) | ( n847 & n1534 ) | ( n1132 & n1534 ) ;
  assign n1764 = ( x107 & n1091 ) | ( x107 & ~n1264 ) | ( n1091 & ~n1264 ) ;
  assign n1765 = ~n136 & n999 ;
  assign n1777 = n167 & n1633 ;
  assign n1778 = n1777 ^ n1664 ^ n352 ;
  assign n1766 = n198 ^ n129 ^ 1'b0 ;
  assign n1767 = ~n131 & n1766 ;
  assign n1768 = n838 & n1767 ;
  assign n1769 = n1768 ^ n1514 ^ 1'b0 ;
  assign n1770 = n904 & ~n1769 ;
  assign n1771 = n1770 ^ n309 ^ 1'b0 ;
  assign n1772 = n234 | n1079 ;
  assign n1773 = n1391 ^ n1085 ^ 1'b0 ;
  assign n1774 = ~n1772 & n1773 ;
  assign n1775 = n1774 ^ n360 ^ 1'b0 ;
  assign n1776 = ~n1771 & n1775 ;
  assign n1779 = n1778 ^ n1776 ^ 1'b0 ;
  assign n1780 = n1779 ^ n1070 ^ n569 ;
  assign n1786 = ( n180 & ~n252 ) | ( n180 & n537 ) | ( ~n252 & n537 ) ;
  assign n1787 = n338 & ~n1786 ;
  assign n1788 = n399 & n1787 ;
  assign n1781 = n243 | n667 ;
  assign n1782 = n143 | n1781 ;
  assign n1783 = n1782 ^ n451 ^ n130 ;
  assign n1784 = ( n497 & n1066 ) | ( n497 & ~n1783 ) | ( n1066 & ~n1783 ) ;
  assign n1785 = ( n645 & ~n1285 ) | ( n645 & n1784 ) | ( ~n1285 & n1784 ) ;
  assign n1789 = n1788 ^ n1785 ^ n808 ;
  assign n1790 = n1595 | n1789 ;
  assign n1791 = ( x10 & n162 ) | ( x10 & n673 ) | ( n162 & n673 ) ;
  assign n1792 = n483 | n1531 ;
  assign n1793 = n1792 ^ n1531 ^ 1'b0 ;
  assign n1794 = ( n147 & n685 ) | ( n147 & ~n1793 ) | ( n685 & ~n1793 ) ;
  assign n1795 = ( n808 & n1791 ) | ( n808 & n1794 ) | ( n1791 & n1794 ) ;
  assign n1796 = ( n253 & n971 ) | ( n253 & n1795 ) | ( n971 & n1795 ) ;
  assign n1798 = n476 ^ n133 ^ 1'b0 ;
  assign n1799 = n1798 ^ n850 ^ 1'b0 ;
  assign n1800 = n235 | n1799 ;
  assign n1801 = n633 | n911 ;
  assign n1802 = n1800 & ~n1801 ;
  assign n1797 = n654 ^ n643 ^ n489 ;
  assign n1803 = n1802 ^ n1797 ^ n620 ;
  assign n1804 = n335 & ~n1803 ;
  assign n1805 = n1331 & ~n1804 ;
  assign n1806 = ( x106 & ~n484 ) | ( x106 & n572 ) | ( ~n484 & n572 ) ;
  assign n1807 = n437 & ~n1806 ;
  assign n1808 = ~n1026 & n1807 ;
  assign n1809 = ( ~n244 & n1127 ) | ( ~n244 & n1808 ) | ( n1127 & n1808 ) ;
  assign n1818 = n597 ^ n392 ^ n145 ;
  assign n1819 = ( n317 & n366 ) | ( n317 & n1818 ) | ( n366 & n1818 ) ;
  assign n1817 = n264 | n314 ;
  assign n1820 = n1819 ^ n1817 ^ n1431 ;
  assign n1810 = n298 & ~n747 ;
  assign n1811 = n177 & n1810 ;
  assign n1812 = n169 | n1811 ;
  assign n1813 = n414 & ~n1812 ;
  assign n1814 = ( n641 & n714 ) | ( n641 & n1813 ) | ( n714 & n1813 ) ;
  assign n1815 = n1814 ^ n180 ^ x70 ;
  assign n1816 = n1815 ^ n253 ^ n250 ;
  assign n1821 = n1820 ^ n1816 ^ n1120 ;
  assign n1822 = x45 & ~n566 ;
  assign n1823 = n1822 ^ n1279 ^ 1'b0 ;
  assign n1824 = n366 | n1823 ;
  assign n1825 = n157 | n1824 ;
  assign n1826 = n1825 ^ n916 ^ 1'b0 ;
  assign n1827 = x43 & ~n872 ;
  assign n1828 = n584 & n1827 ;
  assign n1829 = n1828 ^ n1097 ^ n614 ;
  assign n1830 = ( ~x42 & x91 ) | ( ~x42 & n136 ) | ( x91 & n136 ) ;
  assign n1831 = ( n1194 & ~n1336 ) | ( n1194 & n1830 ) | ( ~n1336 & n1830 ) ;
  assign n1832 = ~n1028 & n1341 ;
  assign n1833 = ( n179 & n643 ) | ( n179 & n1832 ) | ( n643 & n1832 ) ;
  assign n1837 = n364 & n570 ;
  assign n1838 = ( x66 & ~n1473 ) | ( x66 & n1837 ) | ( ~n1473 & n1837 ) ;
  assign n1834 = ( x32 & n364 ) | ( x32 & n524 ) | ( n364 & n524 ) ;
  assign n1835 = n1834 ^ n1550 ^ n896 ;
  assign n1836 = n978 & n1835 ;
  assign n1839 = n1838 ^ n1836 ^ 1'b0 ;
  assign n1840 = n1839 ^ n1189 ^ 1'b0 ;
  assign n1841 = n1343 & ~n1840 ;
  assign n1842 = n1659 ^ n802 ^ 1'b0 ;
  assign n1843 = n1752 & n1842 ;
  assign n1844 = n1841 & n1843 ;
  assign n1847 = n768 ^ n436 ^ x64 ;
  assign n1848 = ( n272 & n1090 ) | ( n272 & ~n1847 ) | ( n1090 & ~n1847 ) ;
  assign n1846 = ( x116 & n1489 ) | ( x116 & ~n1553 ) | ( n1489 & ~n1553 ) ;
  assign n1845 = n1684 ^ n213 ^ 1'b0 ;
  assign n1849 = n1848 ^ n1846 ^ n1845 ;
  assign n1850 = n756 ^ n247 ^ n131 ;
  assign n1851 = ~n648 & n1850 ;
  assign n1852 = n1851 ^ n849 ^ 1'b0 ;
  assign n1853 = n1852 ^ n550 ^ n315 ;
  assign n1854 = ( x23 & ~n1357 ) | ( x23 & n1853 ) | ( ~n1357 & n1853 ) ;
  assign n1855 = ( x107 & n169 ) | ( x107 & n451 ) | ( n169 & n451 ) ;
  assign n1856 = n981 ^ n803 ^ x45 ;
  assign n1857 = ( ~n1451 & n1855 ) | ( ~n1451 & n1856 ) | ( n1855 & n1856 ) ;
  assign n1858 = n1795 ^ n1316 ^ n748 ;
  assign n1859 = ( n146 & ~n294 ) | ( n146 & n421 ) | ( ~n294 & n421 ) ;
  assign n1860 = n1102 ^ n1046 ^ n273 ;
  assign n1861 = n782 | n1860 ;
  assign n1862 = n1859 | n1861 ;
  assign n1863 = n1862 ^ n1830 ^ n676 ;
  assign n1864 = n1317 & n1364 ;
  assign n1865 = n1864 ^ n270 ^ 1'b0 ;
  assign n1866 = n1299 ^ n1154 ^ 1'b0 ;
  assign n1867 = n1865 & n1866 ;
  assign n1868 = n393 ^ n182 ^ 1'b0 ;
  assign n1869 = n1868 ^ n836 ^ 1'b0 ;
  assign n1870 = ~n568 & n1869 ;
  assign n1871 = n1084 ^ n523 ^ n414 ;
  assign n1872 = n1871 ^ x63 ^ 1'b0 ;
  assign n1873 = ( x83 & n1870 ) | ( x83 & ~n1872 ) | ( n1870 & ~n1872 ) ;
  assign n1874 = n876 ^ n706 ^ 1'b0 ;
  assign n1875 = ( n950 & ~n1193 ) | ( n950 & n1874 ) | ( ~n1193 & n1874 ) ;
  assign n1878 = n1244 ^ n250 ^ x14 ;
  assign n1879 = n1878 ^ n422 ^ x2 ;
  assign n1880 = ( n176 & n264 ) | ( n176 & n1879 ) | ( n264 & n1879 ) ;
  assign n1881 = ( ~n378 & n539 ) | ( ~n378 & n1880 ) | ( n539 & n1880 ) ;
  assign n1876 = ~x117 & n490 ;
  assign n1877 = n986 & n1876 ;
  assign n1882 = n1881 ^ n1877 ^ 1'b0 ;
  assign n1883 = n1882 ^ n1824 ^ 1'b0 ;
  assign n1884 = n288 & ~n544 ;
  assign n1885 = n1883 & n1884 ;
  assign n1886 = n1516 ^ n356 ^ n242 ;
  assign n1887 = ( n165 & n698 ) | ( n165 & ~n1886 ) | ( n698 & ~n1886 ) ;
  assign n1888 = n1778 ^ n1504 ^ n310 ;
  assign n1889 = n375 | n517 ;
  assign n1890 = x12 | n1889 ;
  assign n1891 = ( n497 & ~n901 ) | ( n497 & n1361 ) | ( ~n901 & n1361 ) ;
  assign n1892 = n1890 & n1891 ;
  assign n1893 = n1892 ^ n1376 ^ 1'b0 ;
  assign n1894 = n961 ^ n703 ^ x15 ;
  assign n1895 = ( n316 & ~n375 ) | ( n316 & n1894 ) | ( ~n375 & n1894 ) ;
  assign n1896 = ( n442 & ~n813 ) | ( n442 & n1073 ) | ( ~n813 & n1073 ) ;
  assign n1897 = n293 & n1896 ;
  assign n1898 = ( n253 & ~n1176 ) | ( n253 & n1897 ) | ( ~n1176 & n1897 ) ;
  assign n1899 = ~n511 & n1062 ;
  assign n1900 = n1454 & n1885 ;
  assign n1901 = ( ~x8 & n1305 ) | ( ~x8 & n1355 ) | ( n1305 & n1355 ) ;
  assign n1902 = n1901 ^ n1429 ^ n1145 ;
  assign n1903 = ( n454 & ~n472 ) | ( n454 & n667 ) | ( ~n472 & n667 ) ;
  assign n1904 = n372 & ~n1903 ;
  assign n1905 = n1904 ^ n1878 ^ n1727 ;
  assign n1908 = ( n483 & n1188 ) | ( n483 & ~n1879 ) | ( n1188 & ~n1879 ) ;
  assign n1906 = n895 & n1815 ;
  assign n1907 = ~n1847 & n1906 ;
  assign n1909 = n1908 ^ n1907 ^ n1603 ;
  assign n1910 = n1112 ^ n272 ^ n254 ;
  assign n1911 = n1910 ^ n1664 ^ n426 ;
  assign n1912 = n1132 ^ x89 ^ 1'b0 ;
  assign n1913 = n1912 ^ n1227 ^ 1'b0 ;
  assign n1914 = ( ~n1115 & n1911 ) | ( ~n1115 & n1913 ) | ( n1911 & n1913 ) ;
  assign n1915 = n964 ^ n530 ^ x112 ;
  assign n1916 = x114 & ~n1915 ;
  assign n1917 = ( x68 & ~n1043 ) | ( x68 & n1916 ) | ( ~n1043 & n1916 ) ;
  assign n1918 = n1303 & ~n1755 ;
  assign n1919 = ( x94 & n471 ) | ( x94 & n1233 ) | ( n471 & n1233 ) ;
  assign n1920 = n1919 ^ n1148 ^ n279 ;
  assign n1921 = n486 | n568 ;
  assign n1922 = n1672 | n1921 ;
  assign n1923 = n1922 ^ n670 ^ 1'b0 ;
  assign n1924 = ( n295 & ~n1616 ) | ( n295 & n1728 ) | ( ~n1616 & n1728 ) ;
  assign n1925 = ~n1575 & n1626 ;
  assign n1926 = n1924 & ~n1925 ;
  assign n1927 = n830 ^ x95 ^ 1'b0 ;
  assign n1928 = n1927 ^ n130 ^ x112 ;
  assign n1929 = n1619 ^ n1609 ^ n553 ;
  assign n1930 = n380 | n1929 ;
  assign n1931 = n1699 | n1930 ;
  assign n1932 = n1744 ^ x38 ^ x12 ;
  assign n1933 = n1932 ^ n1541 ^ n770 ;
  assign n1934 = x119 & ~n1203 ;
  assign n1935 = n1933 & n1934 ;
  assign n1936 = n297 | n1500 ;
  assign n1937 = n1638 ^ n180 ^ 1'b0 ;
  assign n1938 = ~n256 & n1937 ;
  assign n1939 = ~n621 & n1938 ;
  assign n1940 = n1939 ^ n153 ^ 1'b0 ;
  assign n1941 = n990 & n1940 ;
  assign n1942 = n1941 ^ n961 ^ 1'b0 ;
  assign n1943 = n1942 ^ n1586 ^ n422 ;
  assign n1944 = n582 | n1036 ;
  assign n1945 = x110 ^ x87 ^ x30 ;
  assign n1946 = n1945 ^ n988 ^ n880 ;
  assign n1947 = n1944 & ~n1946 ;
  assign n1952 = n1406 ^ n788 ^ n267 ;
  assign n1948 = x99 & ~n1123 ;
  assign n1949 = ~n713 & n1948 ;
  assign n1950 = n1189 ^ n1149 ^ 1'b0 ;
  assign n1951 = n1949 | n1950 ;
  assign n1953 = n1952 ^ n1951 ^ 1'b0 ;
  assign n1954 = n532 & n869 ;
  assign n1955 = n1954 ^ x100 ^ 1'b0 ;
  assign n1956 = ( n611 & n1519 ) | ( n611 & ~n1903 ) | ( n1519 & ~n1903 ) ;
  assign n1957 = ( ~x111 & n288 ) | ( ~x111 & n664 ) | ( n288 & n664 ) ;
  assign n1958 = ( n179 & n569 ) | ( n179 & ~n1370 ) | ( n569 & ~n1370 ) ;
  assign n1959 = n436 & n1958 ;
  assign n1960 = ( n1956 & n1957 ) | ( n1956 & ~n1959 ) | ( n1957 & ~n1959 ) ;
  assign n1961 = n1955 | n1960 ;
  assign n1962 = x86 | n1961 ;
  assign n1963 = n544 ^ x37 ^ 1'b0 ;
  assign n1964 = n1868 & ~n1963 ;
  assign n1965 = n1964 ^ n1197 ^ 1'b0 ;
  assign n1966 = ~n1765 & n1965 ;
  assign n1967 = n1966 ^ n1175 ^ 1'b0 ;
  assign n1968 = n1374 ^ n1104 ^ x2 ;
  assign n1969 = ( n986 & ~n1444 ) | ( n986 & n1968 ) | ( ~n1444 & n1968 ) ;
  assign n1987 = ( n186 & ~n236 ) | ( n186 & n1020 ) | ( ~n236 & n1020 ) ;
  assign n1985 = n1059 ^ n1015 ^ 1'b0 ;
  assign n1986 = n1795 & n1985 ;
  assign n1970 = n267 & ~n1073 ;
  assign n1971 = n1970 ^ n1206 ^ 1'b0 ;
  assign n1979 = n724 | n934 ;
  assign n1980 = n1979 ^ n1783 ^ 1'b0 ;
  assign n1981 = ~n1782 & n1980 ;
  assign n1977 = n326 ^ n302 ^ x29 ;
  assign n1972 = ( n397 & ~n601 ) | ( n397 & n615 ) | ( ~n601 & n615 ) ;
  assign n1973 = ( ~x14 & x17 ) | ( ~x14 & n1972 ) | ( x17 & n1972 ) ;
  assign n1974 = x39 ^ x34 ^ 1'b0 ;
  assign n1975 = n1973 & n1974 ;
  assign n1976 = ~n485 & n1975 ;
  assign n1978 = n1977 ^ n1976 ^ n1397 ;
  assign n1982 = n1981 ^ n1978 ^ n1647 ;
  assign n1983 = ~n1971 & n1982 ;
  assign n1984 = n1983 ^ n1785 ^ 1'b0 ;
  assign n1988 = n1987 ^ n1986 ^ n1984 ;
  assign n1989 = n1306 ^ n595 ^ n182 ;
  assign n1990 = n160 | n1727 ;
  assign n1991 = n1332 | n1990 ;
  assign n1992 = n1991 ^ n981 ^ 1'b0 ;
  assign n1993 = n500 & ~n619 ;
  assign n1994 = n1993 ^ n297 ^ 1'b0 ;
  assign n1995 = n1994 ^ x53 ^ 1'b0 ;
  assign n1996 = ~n1992 & n1995 ;
  assign n1997 = ~n1970 & n1996 ;
  assign n1998 = x11 & n1248 ;
  assign n1999 = ~n1466 & n1998 ;
  assign n2000 = n1999 ^ n561 ^ n179 ;
  assign n2013 = n1159 ^ x110 ^ x21 ;
  assign n2009 = n563 ^ n434 ^ n426 ;
  assign n2010 = n2009 ^ n164 ^ x42 ;
  assign n2011 = n1084 | n2010 ;
  assign n2012 = ( x80 & ~x111 ) | ( x80 & n2011 ) | ( ~x111 & n2011 ) ;
  assign n2001 = n485 & ~n1860 ;
  assign n2002 = n2001 ^ n217 ^ 1'b0 ;
  assign n2003 = n839 & ~n1456 ;
  assign n2004 = n2003 ^ n1656 ^ 1'b0 ;
  assign n2005 = n2004 ^ x114 ^ 1'b0 ;
  assign n2006 = n2002 & n2005 ;
  assign n2007 = n895 ^ n383 ^ 1'b0 ;
  assign n2008 = n2006 & n2007 ;
  assign n2014 = n2013 ^ n2012 ^ n2008 ;
  assign n2015 = n538 & n1525 ;
  assign n2016 = n1800 & n2015 ;
  assign n2017 = n1846 ^ x51 ^ 1'b0 ;
  assign n2018 = ~n2016 & n2017 ;
  assign n2020 = n943 ^ n353 ^ 1'b0 ;
  assign n2019 = n659 | n911 ;
  assign n2021 = n2020 ^ n2019 ^ 1'b0 ;
  assign n2022 = ~n523 & n2021 ;
  assign n2023 = ~n2018 & n2022 ;
  assign n2024 = n413 & n933 ;
  assign n2025 = ~n1671 & n2024 ;
  assign n2027 = n1915 ^ n629 ^ n271 ;
  assign n2026 = n1297 ^ n750 ^ 1'b0 ;
  assign n2028 = n2027 ^ n2026 ^ 1'b0 ;
  assign n2029 = x54 & ~n2028 ;
  assign n2030 = n561 & ~n1069 ;
  assign n2031 = n1639 & n2030 ;
  assign n2032 = n2031 ^ x79 ^ 1'b0 ;
  assign n2033 = ( n1912 & n2029 ) | ( n1912 & ~n2032 ) | ( n2029 & ~n2032 ) ;
  assign n2034 = x59 & n961 ;
  assign n2035 = ~n2033 & n2034 ;
  assign n2036 = x63 & ~n263 ;
  assign n2037 = n2036 ^ n632 ^ 1'b0 ;
  assign n2038 = ( ~n250 & n1082 ) | ( ~n250 & n1132 ) | ( n1082 & n1132 ) ;
  assign n2039 = n1412 & ~n2038 ;
  assign n2040 = n2039 ^ n656 ^ 1'b0 ;
  assign n2041 = x30 & ~n1122 ;
  assign n2042 = n213 & n2041 ;
  assign n2043 = n1472 ^ n572 ^ 1'b0 ;
  assign n2044 = ~n2042 & n2043 ;
  assign n2045 = ~n713 & n2044 ;
  assign n2046 = n1543 ^ n1025 ^ n438 ;
  assign n2047 = n828 & ~n2046 ;
  assign n2048 = ( x107 & ~n431 ) | ( x107 & n1213 ) | ( ~n431 & n1213 ) ;
  assign n2049 = n167 & ~n292 ;
  assign n2050 = ( ~n786 & n2048 ) | ( ~n786 & n2049 ) | ( n2048 & n2049 ) ;
  assign n2051 = ( n924 & n2047 ) | ( n924 & ~n2050 ) | ( n2047 & ~n2050 ) ;
  assign n2053 = x2 & x98 ;
  assign n2054 = n964 & n2053 ;
  assign n2055 = ~n198 & n2054 ;
  assign n2052 = ( x3 & ~n1095 ) | ( x3 & n1246 ) | ( ~n1095 & n1246 ) ;
  assign n2056 = n2055 ^ n2052 ^ x108 ;
  assign n2057 = ( x84 & n1084 ) | ( x84 & ~n1558 ) | ( n1084 & ~n1558 ) ;
  assign n2058 = n633 ^ n399 ^ x112 ;
  assign n2059 = ( x101 & ~n166 ) | ( x101 & n2058 ) | ( ~n166 & n2058 ) ;
  assign n2060 = ( n2056 & n2057 ) | ( n2056 & ~n2059 ) | ( n2057 & ~n2059 ) ;
  assign n2061 = n1531 | n1997 ;
  assign n2069 = n1728 ^ n1490 ^ n360 ;
  assign n2070 = ( n1533 & n1539 ) | ( n1533 & n2069 ) | ( n1539 & n2069 ) ;
  assign n2062 = n691 ^ n227 ^ x1 ;
  assign n2063 = ( n744 & n805 ) | ( n744 & ~n1431 ) | ( n805 & ~n1431 ) ;
  assign n2064 = n1541 ^ n426 ^ 1'b0 ;
  assign n2065 = ~n2063 & n2064 ;
  assign n2066 = ~x102 & n1155 ;
  assign n2067 = n2065 & n2066 ;
  assign n2068 = n2062 | n2067 ;
  assign n2071 = n2070 ^ n2068 ^ 1'b0 ;
  assign n2072 = ( x5 & ~n883 ) | ( x5 & n996 ) | ( ~n883 & n996 ) ;
  assign n2073 = n1769 ^ n1510 ^ n1183 ;
  assign n2074 = n1793 ^ n994 ^ 1'b0 ;
  assign n2075 = ~n2073 & n2074 ;
  assign n2076 = n1026 & ~n1806 ;
  assign n2077 = n2076 ^ n814 ^ n273 ;
  assign n2078 = n429 & ~n766 ;
  assign n2079 = ( n1323 & ~n2077 ) | ( n1323 & n2078 ) | ( ~n2077 & n2078 ) ;
  assign n2082 = x23 & ~n351 ;
  assign n2080 = n214 ^ x85 ^ 1'b0 ;
  assign n2081 = x37 & ~n2080 ;
  assign n2083 = n2082 ^ n2081 ^ n814 ;
  assign n2084 = n2083 ^ n1152 ^ 1'b0 ;
  assign n2085 = n1529 & ~n2084 ;
  assign n2086 = n772 ^ n195 ^ 1'b0 ;
  assign n2087 = n1847 ^ n1171 ^ n250 ;
  assign n2088 = n1530 ^ n639 ^ 1'b0 ;
  assign n2089 = ( n1870 & ~n2087 ) | ( n1870 & n2088 ) | ( ~n2087 & n2088 ) ;
  assign n2090 = n1022 & ~n2089 ;
  assign n2091 = n773 | n1656 ;
  assign n2092 = n725 | n2091 ;
  assign n2093 = n2090 | n2092 ;
  assign n2094 = n1725 ^ n435 ^ 1'b0 ;
  assign n2095 = n2094 ^ n1977 ^ n1483 ;
  assign n2096 = n366 & n1324 ;
  assign n2097 = ( n298 & n315 ) | ( n298 & ~n2082 ) | ( n315 & ~n2082 ) ;
  assign n2098 = n1547 & n2097 ;
  assign n2099 = ~n226 & n451 ;
  assign n2100 = n981 & n2099 ;
  assign n2101 = n1339 ^ n312 ^ 1'b0 ;
  assign n2102 = ~n250 & n2101 ;
  assign n2104 = x33 & ~n204 ;
  assign n2105 = n2104 ^ n1002 ^ 1'b0 ;
  assign n2103 = n1797 ^ n1736 ^ n880 ;
  assign n2106 = n2105 ^ n2103 ^ n404 ;
  assign n2107 = n244 | n2106 ;
  assign n2109 = n148 | n1053 ;
  assign n2108 = n391 & n484 ;
  assign n2110 = n2109 ^ n2108 ^ n315 ;
  assign n2112 = ( n172 & n759 ) | ( n172 & n937 ) | ( n759 & n937 ) ;
  assign n2111 = n972 ^ n615 ^ n512 ;
  assign n2113 = n2112 ^ n2111 ^ n918 ;
  assign n2114 = ( n1011 & n1470 ) | ( n1011 & ~n2113 ) | ( n1470 & ~n2113 ) ;
  assign n2115 = ~n462 & n2114 ;
  assign n2116 = ~n2110 & n2115 ;
  assign n2117 = ( n635 & ~n2107 ) | ( n635 & n2116 ) | ( ~n2107 & n2116 ) ;
  assign n2118 = n1426 ^ n240 ^ x74 ;
  assign n2119 = n1977 ^ n433 ^ x22 ;
  assign n2120 = ( ~n544 & n1353 ) | ( ~n544 & n1541 ) | ( n1353 & n1541 ) ;
  assign n2121 = ( ~x59 & n1285 ) | ( ~x59 & n2120 ) | ( n1285 & n2120 ) ;
  assign n2122 = ~n279 & n1360 ;
  assign n2123 = x115 & ~n2122 ;
  assign n2124 = n2121 & n2123 ;
  assign n2125 = n2124 ^ n798 ^ 1'b0 ;
  assign n2126 = x101 & n2125 ;
  assign n2132 = n688 ^ n676 ^ n392 ;
  assign n2127 = n617 ^ n530 ^ 1'b0 ;
  assign n2128 = n304 & n2127 ;
  assign n2129 = n1023 ^ n667 ^ 1'b0 ;
  assign n2130 = n2128 & ~n2129 ;
  assign n2131 = ( n145 & n2089 ) | ( n145 & ~n2130 ) | ( n2089 & ~n2130 ) ;
  assign n2133 = n2132 ^ n2131 ^ 1'b0 ;
  assign n2134 = n945 & n2133 ;
  assign n2135 = n1584 ^ n156 ^ x117 ;
  assign n2136 = n2135 ^ n1947 ^ n513 ;
  assign n2137 = n1732 ^ n572 ^ n447 ;
  assign n2138 = ( ~x99 & n814 ) | ( ~x99 & n1155 ) | ( n814 & n1155 ) ;
  assign n2139 = ~n1602 & n2138 ;
  assign n2140 = n2139 ^ n1149 ^ 1'b0 ;
  assign n2141 = ( n1010 & n1068 ) | ( n1010 & ~n1437 ) | ( n1068 & ~n1437 ) ;
  assign n2142 = n2141 ^ n622 ^ n522 ;
  assign n2143 = n1269 ^ n826 ^ 1'b0 ;
  assign n2144 = n2143 ^ n620 ^ 1'b0 ;
  assign n2145 = n2142 & ~n2144 ;
  assign n2146 = ~n924 & n2145 ;
  assign n2147 = n1159 ^ n625 ^ n616 ;
  assign n2148 = x116 & n2147 ;
  assign n2149 = n2148 ^ n426 ^ 1'b0 ;
  assign n2150 = n444 & ~n2149 ;
  assign n2151 = ( n394 & n1675 ) | ( n394 & n2150 ) | ( n1675 & n2150 ) ;
  assign n2152 = n2151 ^ n1582 ^ n1558 ;
  assign n2153 = ~n279 & n1813 ;
  assign n2154 = n2153 ^ n890 ^ 1'b0 ;
  assign n2155 = n323 & ~n1133 ;
  assign n2156 = ~n1360 & n2155 ;
  assign n2157 = ~n259 & n2156 ;
  assign n2160 = n2130 ^ n1220 ^ n147 ;
  assign n2158 = n834 ^ x50 ^ 1'b0 ;
  assign n2159 = n242 & ~n2158 ;
  assign n2161 = n2160 ^ n2159 ^ n555 ;
  assign n2162 = n2161 ^ n933 ^ 1'b0 ;
  assign n2163 = ~n2157 & n2162 ;
  assign n2164 = n311 ^ n272 ^ 1'b0 ;
  assign n2165 = n380 | n2164 ;
  assign n2166 = n2165 ^ n497 ^ 1'b0 ;
  assign n2167 = n1051 | n2166 ;
  assign n2168 = n2167 ^ n2066 ^ n1289 ;
  assign n2169 = n1057 ^ n588 ^ 1'b0 ;
  assign n2170 = ( n309 & n326 ) | ( n309 & n657 ) | ( n326 & n657 ) ;
  assign n2171 = n1870 ^ n1536 ^ n1477 ;
  assign n2172 = ( n1338 & n2170 ) | ( n1338 & n2171 ) | ( n2170 & n2171 ) ;
  assign n2176 = n2082 ^ n1419 ^ n1129 ;
  assign n2177 = n512 ^ n275 ^ 1'b0 ;
  assign n2178 = n2176 & ~n2177 ;
  assign n2173 = n716 ^ n636 ^ 1'b0 ;
  assign n2174 = x16 & n2173 ;
  assign n2175 = n2174 ^ n633 ^ n205 ;
  assign n2179 = n2178 ^ n2175 ^ n878 ;
  assign n2180 = n2179 ^ n949 ^ 1'b0 ;
  assign n2181 = n2172 & ~n2180 ;
  assign n2182 = ~n367 & n674 ;
  assign n2183 = ~n532 & n2182 ;
  assign n2184 = ( ~n279 & n1189 ) | ( ~n279 & n2183 ) | ( n1189 & n2183 ) ;
  assign n2185 = ( ~n1463 & n1876 ) | ( ~n1463 & n2184 ) | ( n1876 & n2184 ) ;
  assign n2186 = n1143 ^ n437 ^ 1'b0 ;
  assign n2187 = ( n1247 & n2185 ) | ( n1247 & n2186 ) | ( n2185 & n2186 ) ;
  assign n2188 = ( n145 & ~n172 ) | ( n145 & n1045 ) | ( ~n172 & n1045 ) ;
  assign n2189 = ( ~n767 & n1573 ) | ( ~n767 & n2188 ) | ( n1573 & n2188 ) ;
  assign n2190 = n935 ^ n211 ^ 1'b0 ;
  assign n2191 = n2190 ^ n762 ^ 1'b0 ;
  assign n2192 = n710 & n2191 ;
  assign n2193 = ( n890 & ~n2189 ) | ( n890 & n2192 ) | ( ~n2189 & n2192 ) ;
  assign n2194 = n2193 ^ n1711 ^ n322 ;
  assign n2195 = n2116 ^ n1943 ^ n1411 ;
  assign n2196 = n1509 ^ n1332 ^ n387 ;
  assign n2197 = n1899 ^ n1314 ^ n1108 ;
  assign n2198 = n2197 ^ n1424 ^ n295 ;
  assign n2199 = n1978 ^ n1476 ^ x53 ;
  assign n2200 = n1880 ^ n1348 ^ n180 ;
  assign n2201 = n2200 ^ n775 ^ 1'b0 ;
  assign n2203 = ( ~n151 & n826 ) | ( ~n151 & n832 ) | ( n826 & n832 ) ;
  assign n2202 = n756 & n1475 ;
  assign n2204 = n2203 ^ n2202 ^ 1'b0 ;
  assign n2205 = ( n270 & ~n1234 ) | ( n270 & n2204 ) | ( ~n1234 & n2204 ) ;
  assign n2206 = n2205 ^ n1441 ^ n386 ;
  assign n2207 = n1511 ^ n1234 ^ 1'b0 ;
  assign n2208 = n2207 ^ n948 ^ 1'b0 ;
  assign n2209 = n2206 & n2208 ;
  assign n2210 = n1134 ^ n378 ^ n263 ;
  assign n2211 = n2210 ^ n518 ^ 1'b0 ;
  assign n2212 = n1285 ^ n1273 ^ 1'b0 ;
  assign n2213 = n2212 ^ n1629 ^ 1'b0 ;
  assign n2214 = n880 ^ n190 ^ x25 ;
  assign n2215 = ( n1628 & n1767 ) | ( n1628 & ~n2214 ) | ( n1767 & ~n2214 ) ;
  assign n2216 = n1052 ^ n1026 ^ 1'b0 ;
  assign n2219 = ~n399 & n724 ;
  assign n2218 = n512 & ~n872 ;
  assign n2220 = n2219 ^ n2218 ^ n1280 ;
  assign n2221 = n285 & n896 ;
  assign n2222 = ~n2220 & n2221 ;
  assign n2217 = n1322 & ~n2006 ;
  assign n2223 = n2222 ^ n2217 ^ 1'b0 ;
  assign n2224 = ( n315 & ~n1273 ) | ( n315 & n1511 ) | ( ~n1273 & n1511 ) ;
  assign n2225 = n472 ^ x109 ^ 1'b0 ;
  assign n2226 = n981 | n2225 ;
  assign n2227 = n2226 ^ x120 ^ x27 ;
  assign n2230 = ~n217 & n501 ;
  assign n2228 = n956 ^ n553 ^ 1'b0 ;
  assign n2229 = n1559 & ~n2228 ;
  assign n2231 = n2230 ^ n2229 ^ 1'b0 ;
  assign n2232 = n2227 & n2231 ;
  assign n2240 = n645 | n828 ;
  assign n2241 = n1874 & ~n2240 ;
  assign n2233 = n988 | n1277 ;
  assign n2234 = n2233 ^ n695 ^ 1'b0 ;
  assign n2235 = n2234 ^ n1320 ^ 1'b0 ;
  assign n2236 = n138 | n2235 ;
  assign n2237 = ( n584 & n794 ) | ( n584 & ~n2236 ) | ( n794 & ~n2236 ) ;
  assign n2238 = n2237 ^ n1668 ^ 1'b0 ;
  assign n2239 = n1891 & n2238 ;
  assign n2242 = n2241 ^ n2239 ^ n927 ;
  assign n2243 = ( n444 & ~n1437 ) | ( n444 & n2042 ) | ( ~n1437 & n2042 ) ;
  assign n2244 = ~n593 & n1314 ;
  assign n2245 = ~n412 & n2244 ;
  assign n2246 = n2245 ^ n1905 ^ n550 ;
  assign n2247 = ( n450 & ~n2243 ) | ( n450 & n2246 ) | ( ~n2243 & n2246 ) ;
  assign n2248 = n1994 & n2020 ;
  assign n2249 = n2170 & n2248 ;
  assign n2250 = n1636 & n1740 ;
  assign n2251 = n2249 & n2250 ;
  assign n2252 = ( n513 & n1439 ) | ( n513 & ~n2251 ) | ( n1439 & ~n2251 ) ;
  assign n2253 = n1282 ^ n387 ^ 1'b0 ;
  assign n2254 = n2253 ^ n1795 ^ 1'b0 ;
  assign n2255 = n1506 ^ n219 ^ x63 ;
  assign n2256 = ~n526 & n750 ;
  assign n2257 = ( n984 & n1882 ) | ( n984 & ~n2256 ) | ( n1882 & ~n2256 ) ;
  assign n2258 = n1359 ^ n513 ^ 1'b0 ;
  assign n2259 = n2258 ^ n937 ^ n291 ;
  assign n2260 = ( x2 & ~n149 ) | ( x2 & n1175 ) | ( ~n149 & n1175 ) ;
  assign n2261 = n762 & n2260 ;
  assign n2267 = n2002 ^ n1531 ^ 1'b0 ;
  assign n2268 = n2267 ^ n1688 ^ 1'b0 ;
  assign n2269 = n950 & ~n2268 ;
  assign n2270 = n621 ^ n185 ^ x71 ;
  assign n2271 = n1008 | n2270 ;
  assign n2272 = n2269 | n2271 ;
  assign n2273 = n2272 ^ n1083 ^ 1'b0 ;
  assign n2262 = n143 & ~n1273 ;
  assign n2263 = n577 | n948 ;
  assign n2264 = n2263 ^ n702 ^ 1'b0 ;
  assign n2265 = n2264 ^ n1329 ^ n897 ;
  assign n2266 = n2262 & ~n2265 ;
  assign n2274 = n2273 ^ n2266 ^ 1'b0 ;
  assign n2275 = n2105 ^ n1109 ^ n600 ;
  assign n2276 = n2275 ^ n378 ^ 1'b0 ;
  assign n2277 = n1021 ^ n151 ^ 1'b0 ;
  assign n2278 = ( n811 & n1590 ) | ( n811 & ~n2111 ) | ( n1590 & ~n2111 ) ;
  assign n2279 = n2278 ^ n1334 ^ x73 ;
  assign n2280 = n2279 ^ n2026 ^ 1'b0 ;
  assign n2281 = n230 | n2280 ;
  assign n2283 = ( x121 & ~n474 ) | ( x121 & n476 ) | ( ~n474 & n476 ) ;
  assign n2284 = n844 ^ x84 ^ 1'b0 ;
  assign n2285 = n2284 ^ n218 ^ 1'b0 ;
  assign n2286 = n2283 & n2285 ;
  assign n2287 = n2286 ^ n644 ^ 1'b0 ;
  assign n2288 = n164 & n2287 ;
  assign n2282 = n1633 ^ n1049 ^ n790 ;
  assign n2289 = n2288 ^ n2282 ^ 1'b0 ;
  assign n2290 = n1006 ^ x37 ^ x34 ;
  assign n2291 = ( ~n665 & n773 ) | ( ~n665 & n1281 ) | ( n773 & n1281 ) ;
  assign n2293 = ( n367 & n412 ) | ( n367 & n1944 ) | ( n412 & n1944 ) ;
  assign n2292 = ( ~n517 & n866 ) | ( ~n517 & n1074 ) | ( n866 & n1074 ) ;
  assign n2294 = n2293 ^ n2292 ^ n1357 ;
  assign n2295 = ( ~n2290 & n2291 ) | ( ~n2290 & n2294 ) | ( n2291 & n2294 ) ;
  assign n2296 = ( ~x46 & n215 ) | ( ~x46 & n493 ) | ( n215 & n493 ) ;
  assign n2297 = n438 & ~n2296 ;
  assign n2298 = ~n763 & n2297 ;
  assign n2299 = n2298 ^ n1785 ^ n615 ;
  assign n2300 = n490 ^ n461 ^ 1'b0 ;
  assign n2301 = ~n1040 & n2300 ;
  assign n2302 = ~n1471 & n2301 ;
  assign n2303 = n2299 & n2302 ;
  assign n2304 = n2303 ^ n1888 ^ n941 ;
  assign n2305 = ~n867 & n1749 ;
  assign n2306 = n2305 ^ x82 ^ 1'b0 ;
  assign n2307 = n1797 ^ n244 ^ 1'b0 ;
  assign n2308 = ~n912 & n1818 ;
  assign n2309 = x118 & ~n2308 ;
  assign n2310 = ~n2307 & n2309 ;
  assign n2311 = n1828 | n2310 ;
  assign n2312 = n2306 & ~n2311 ;
  assign n2313 = ( n294 & ~n1788 ) | ( n294 & n1827 ) | ( ~n1788 & n1827 ) ;
  assign n2314 = n2313 ^ n2135 ^ n418 ;
  assign n2315 = ~n765 & n2314 ;
  assign n2316 = n169 | n901 ;
  assign n2317 = n550 & ~n2316 ;
  assign n2322 = n2029 ^ n1391 ^ 1'b0 ;
  assign n2323 = x3 & n2322 ;
  assign n2324 = n414 & n2323 ;
  assign n2318 = ( x104 & n184 ) | ( x104 & n798 ) | ( n184 & n798 ) ;
  assign n2319 = ( ~n368 & n1755 ) | ( ~n368 & n2318 ) | ( n1755 & n2318 ) ;
  assign n2320 = n989 & ~n2319 ;
  assign n2321 = n2320 ^ n621 ^ 1'b0 ;
  assign n2325 = n2324 ^ n2321 ^ 1'b0 ;
  assign n2326 = ~n660 & n2325 ;
  assign n2327 = n1835 ^ n1752 ^ n519 ;
  assign n2328 = n541 | n614 ;
  assign n2329 = n2328 ^ n835 ^ 1'b0 ;
  assign n2334 = ( n832 & ~n1272 ) | ( n832 & n1621 ) | ( ~n1272 & n1621 ) ;
  assign n2330 = n570 & n663 ;
  assign n2331 = n2330 ^ n1539 ^ 1'b0 ;
  assign n2332 = n2331 ^ n948 ^ 1'b0 ;
  assign n2333 = ~n305 & n2332 ;
  assign n2335 = n2334 ^ n2333 ^ 1'b0 ;
  assign n2336 = ( n1528 & n2329 ) | ( n1528 & n2335 ) | ( n2329 & n2335 ) ;
  assign n2337 = n2327 & n2336 ;
  assign n2338 = ( n457 & ~n599 ) | ( n457 & n674 ) | ( ~n599 & n674 ) ;
  assign n2339 = ~n1804 & n2338 ;
  assign n2340 = n388 & ~n1526 ;
  assign n2341 = ~n1858 & n2340 ;
  assign n2342 = ( ~n697 & n1096 ) | ( ~n697 & n1380 ) | ( n1096 & n1380 ) ;
  assign n2343 = ( n145 & ~n657 ) | ( n145 & n685 ) | ( ~n657 & n685 ) ;
  assign n2344 = n160 | n2343 ;
  assign n2345 = n699 | n724 ;
  assign n2346 = n2345 ^ n478 ^ 1'b0 ;
  assign n2347 = ( n2160 & n2290 ) | ( n2160 & ~n2346 ) | ( n2290 & ~n2346 ) ;
  assign n2348 = ( ~n1208 & n2344 ) | ( ~n1208 & n2347 ) | ( n2344 & n2347 ) ;
  assign n2349 = x94 & ~n598 ;
  assign n2350 = n2349 ^ n155 ^ 1'b0 ;
  assign n2351 = n2350 ^ x74 ^ 1'b0 ;
  assign n2352 = n2348 & ~n2351 ;
  assign n2353 = n2352 ^ n1899 ^ n1621 ;
  assign n2361 = n1977 ^ n484 ^ n410 ;
  assign n2362 = n2361 ^ n886 ^ 1'b0 ;
  assign n2363 = x1 & n2362 ;
  assign n2358 = n680 ^ n392 ^ n168 ;
  assign n2359 = n2358 ^ n896 ^ 1'b0 ;
  assign n2360 = ~n1929 & n2359 ;
  assign n2356 = n484 & ~n694 ;
  assign n2354 = n1419 ^ n468 ^ 1'b0 ;
  assign n2355 = n1913 & n2354 ;
  assign n2357 = n2356 ^ n2355 ^ n1259 ;
  assign n2364 = n2363 ^ n2360 ^ n2357 ;
  assign n2368 = n235 | n488 ;
  assign n2369 = n2368 ^ n432 ^ 1'b0 ;
  assign n2370 = ( x55 & n801 ) | ( x55 & n2369 ) | ( n801 & n2369 ) ;
  assign n2371 = n2370 ^ n1606 ^ 1'b0 ;
  assign n2365 = ( x69 & n298 ) | ( x69 & ~n512 ) | ( n298 & ~n512 ) ;
  assign n2366 = ~n146 & n2365 ;
  assign n2367 = ~n1506 & n2366 ;
  assign n2372 = n2371 ^ n2367 ^ 1'b0 ;
  assign n2373 = n421 & ~n2372 ;
  assign n2374 = n2373 ^ n189 ^ 1'b0 ;
  assign n2375 = n665 | n1313 ;
  assign n2376 = n2375 ^ n2088 ^ 1'b0 ;
  assign n2377 = n133 & ~n1517 ;
  assign n2378 = n1774 ^ n656 ^ 1'b0 ;
  assign n2384 = ( ~n1011 & n1248 ) | ( ~n1011 & n1583 ) | ( n1248 & n1583 ) ;
  assign n2382 = n878 | n1073 ;
  assign n2383 = n2382 ^ x44 ^ 1'b0 ;
  assign n2380 = x102 & n1065 ;
  assign n2379 = ( n1548 & ~n1638 ) | ( n1548 & n1769 ) | ( ~n1638 & n1769 ) ;
  assign n2381 = n2380 ^ n2379 ^ 1'b0 ;
  assign n2385 = n2384 ^ n2383 ^ n2381 ;
  assign n2386 = n1852 ^ n1052 ^ 1'b0 ;
  assign n2387 = n1533 | n2306 ;
  assign n2388 = n2386 & ~n2387 ;
  assign n2390 = ( n1411 & ~n1608 ) | ( n1411 & n1653 ) | ( ~n1608 & n1653 ) ;
  assign n2389 = n992 ^ n915 ^ n337 ;
  assign n2391 = n2390 ^ n2389 ^ n538 ;
  assign n2392 = ( n2197 & ~n2388 ) | ( n2197 & n2391 ) | ( ~n2388 & n2391 ) ;
  assign n2393 = n1217 ^ n807 ^ n315 ;
  assign n2394 = ( n931 & n1282 ) | ( n931 & ~n2393 ) | ( n1282 & ~n2393 ) ;
  assign n2395 = n346 ^ x18 ^ 1'b0 ;
  assign n2396 = n2395 ^ n294 ^ 1'b0 ;
  assign n2397 = n2394 & n2396 ;
  assign n2398 = n2397 ^ n926 ^ 1'b0 ;
  assign n2399 = n1525 ^ n1307 ^ n1298 ;
  assign n2400 = n2399 ^ n625 ^ 1'b0 ;
  assign n2401 = n633 | n2400 ;
  assign n2402 = ( n1573 & n1650 ) | ( n1573 & n2290 ) | ( n1650 & n2290 ) ;
  assign n2404 = n295 ^ x25 ^ 1'b0 ;
  assign n2405 = ~n648 & n2404 ;
  assign n2403 = x123 | n2321 ;
  assign n2406 = n2405 ^ n2403 ^ 1'b0 ;
  assign n2407 = n876 & ~n2406 ;
  assign n2408 = n2407 ^ n1192 ^ 1'b0 ;
  assign n2409 = ~n2402 & n2408 ;
  assign n2410 = ( n374 & n450 ) | ( n374 & n1269 ) | ( n450 & n1269 ) ;
  assign n2411 = n1151 ^ n945 ^ n702 ;
  assign n2412 = n2286 ^ x50 ^ 1'b0 ;
  assign n2413 = ~n2411 & n2412 ;
  assign n2414 = n2410 & n2413 ;
  assign n2415 = ( x121 & ~n441 ) | ( x121 & n1182 ) | ( ~n441 & n1182 ) ;
  assign n2416 = n2415 ^ n1654 ^ 1'b0 ;
  assign n2417 = ( n725 & ~n734 ) | ( n725 & n1171 ) | ( ~n734 & n1171 ) ;
  assign n2418 = ( n760 & n900 ) | ( n760 & n1480 ) | ( n900 & n1480 ) ;
  assign n2419 = n2418 ^ n588 ^ x76 ;
  assign n2420 = ( n1657 & n2417 ) | ( n1657 & ~n2419 ) | ( n2417 & ~n2419 ) ;
  assign n2421 = ( ~n1018 & n2416 ) | ( ~n1018 & n2420 ) | ( n2416 & n2420 ) ;
  assign n2422 = n1046 ^ n865 ^ n788 ;
  assign n2423 = n2422 ^ n1918 ^ 1'b0 ;
  assign n2424 = ( ~n187 & n429 ) | ( ~n187 & n995 ) | ( n429 & n995 ) ;
  assign n2425 = n2424 ^ n408 ^ 1'b0 ;
  assign n2426 = n1466 & n2425 ;
  assign n2427 = n2426 ^ n1266 ^ n353 ;
  assign n2428 = n436 ^ x33 ^ x15 ;
  assign n2429 = ( n256 & n1981 ) | ( n256 & n2428 ) | ( n1981 & n2428 ) ;
  assign n2430 = n199 & ~n1001 ;
  assign n2431 = n2430 ^ n464 ^ 1'b0 ;
  assign n2432 = n2431 ^ x70 ^ x33 ;
  assign n2433 = ( n2072 & n2429 ) | ( n2072 & n2432 ) | ( n2429 & n2432 ) ;
  assign n2434 = n1005 ^ n695 ^ 1'b0 ;
  assign n2435 = n2434 ^ n2267 ^ n1045 ;
  assign n2436 = n181 | n2135 ;
  assign n2437 = ~n1127 & n2436 ;
  assign n2438 = n2434 & n2437 ;
  assign n2439 = n226 | n245 ;
  assign n2440 = n677 & ~n2439 ;
  assign n2441 = n2440 ^ n1081 ^ n962 ;
  assign n2443 = ( n248 & n688 ) | ( n248 & ~n760 ) | ( n688 & ~n760 ) ;
  assign n2442 = n386 & ~n2170 ;
  assign n2444 = n2443 ^ n2442 ^ 1'b0 ;
  assign n2445 = n1225 & ~n1320 ;
  assign n2446 = ( n903 & n1124 ) | ( n903 & ~n2445 ) | ( n1124 & ~n2445 ) ;
  assign n2447 = n2444 & n2446 ;
  assign n2448 = n2441 & n2447 ;
  assign n2449 = n2448 ^ n1316 ^ 1'b0 ;
  assign n2450 = ( ~n272 & n684 ) | ( ~n272 & n1068 ) | ( n684 & n1068 ) ;
  assign n2451 = n2450 ^ n2370 ^ n2055 ;
  assign n2452 = n972 & n1074 ;
  assign n2453 = ~n131 & n2452 ;
  assign n2454 = n2086 | n2453 ;
  assign n2455 = n2454 ^ n2436 ^ 1'b0 ;
  assign n2456 = ( n590 & ~n1806 ) | ( n590 & n1896 ) | ( ~n1806 & n1896 ) ;
  assign n2457 = ~n157 & n863 ;
  assign n2458 = n2457 ^ n281 ^ 1'b0 ;
  assign n2459 = ( ~n1134 & n2456 ) | ( ~n1134 & n2458 ) | ( n2456 & n2458 ) ;
  assign n2460 = ~n351 & n2459 ;
  assign n2461 = n2460 ^ n416 ^ 1'b0 ;
  assign n2462 = n770 & ~n1217 ;
  assign n2463 = x102 & ~n1915 ;
  assign n2464 = n2171 ^ n816 ^ 1'b0 ;
  assign n2465 = ~n719 & n2110 ;
  assign n2466 = ~n1146 & n2465 ;
  assign n2467 = n277 | n2390 ;
  assign n2468 = n2467 ^ n1977 ^ n1621 ;
  assign n2469 = ~n566 & n1194 ;
  assign n2470 = ~n830 & n2469 ;
  assign n2471 = n2470 ^ n1144 ^ n532 ;
  assign n2472 = ( x46 & ~n223 ) | ( x46 & n2471 ) | ( ~n223 & n2471 ) ;
  assign n2473 = x55 & ~n551 ;
  assign n2474 = ~n289 & n2473 ;
  assign n2475 = ( n730 & n2012 ) | ( n730 & ~n2020 ) | ( n2012 & ~n2020 ) ;
  assign n2476 = n2474 | n2475 ;
  assign n2477 = n2476 ^ n1729 ^ 1'b0 ;
  assign n2478 = n1534 ^ n1353 ^ n489 ;
  assign n2479 = ( n289 & ~n610 ) | ( n289 & n2245 ) | ( ~n610 & n2245 ) ;
  assign n2480 = n519 & ~n1683 ;
  assign n2481 = n2480 ^ n783 ^ 1'b0 ;
  assign n2482 = n2481 ^ n910 ^ n515 ;
  assign n2483 = ~n541 & n2482 ;
  assign n2484 = ~n1881 & n2483 ;
  assign n2485 = ( x14 & n1847 ) | ( x14 & ~n2160 ) | ( n1847 & ~n2160 ) ;
  assign n2486 = ( n489 & n2484 ) | ( n489 & ~n2485 ) | ( n2484 & ~n2485 ) ;
  assign n2490 = ~x36 & n461 ;
  assign n2487 = n1959 ^ n1722 ^ n1375 ;
  assign n2488 = n2487 ^ n649 ^ n285 ;
  assign n2489 = ( ~n1048 & n1798 ) | ( ~n1048 & n2488 ) | ( n1798 & n2488 ) ;
  assign n2491 = n2490 ^ n2489 ^ 1'b0 ;
  assign n2492 = ( ~x38 & n598 ) | ( ~x38 & n998 ) | ( n598 & n998 ) ;
  assign n2493 = n2071 & ~n2492 ;
  assign n2494 = n1828 & n1873 ;
  assign n2495 = n2283 ^ n236 ^ n177 ;
  assign n2496 = n1731 | n2495 ;
  assign n2497 = ~n264 & n2496 ;
  assign n2498 = n1261 & n2497 ;
  assign n2499 = ( n203 & n2494 ) | ( n203 & n2498 ) | ( n2494 & n2498 ) ;
  assign n2500 = n1076 ^ n834 ^ n635 ;
  assign n2501 = n2500 ^ n1036 ^ 1'b0 ;
  assign n2502 = n2501 ^ n1468 ^ 1'b0 ;
  assign n2503 = n1838 | n2502 ;
  assign n2504 = n1007 & ~n2503 ;
  assign n2509 = n2176 ^ n834 ^ n395 ;
  assign n2510 = n2509 ^ n1030 ^ n323 ;
  assign n2511 = n2510 ^ n1082 ^ n929 ;
  assign n2505 = x126 & ~n1220 ;
  assign n2506 = ~n512 & n2505 ;
  assign n2507 = n2506 ^ n1706 ^ n865 ;
  assign n2508 = ~n2411 & n2507 ;
  assign n2512 = n2511 ^ n2508 ^ 1'b0 ;
  assign n2521 = n2452 ^ n1023 ^ x52 ;
  assign n2522 = n2521 ^ n826 ^ 1'b0 ;
  assign n2523 = n2236 | n2522 ;
  assign n2524 = n2523 ^ n2292 ^ n1550 ;
  assign n2530 = n530 & n1176 ;
  assign n2525 = n705 ^ n643 ^ 1'b0 ;
  assign n2526 = ~n163 & n2525 ;
  assign n2527 = n2526 ^ n1749 ^ n629 ;
  assign n2528 = n2527 ^ n2090 ^ 1'b0 ;
  assign n2529 = n750 & ~n2528 ;
  assign n2531 = n2530 ^ n2529 ^ 1'b0 ;
  assign n2532 = n2524 & n2531 ;
  assign n2518 = n1473 & ~n1788 ;
  assign n2519 = n2518 ^ n599 ^ 1'b0 ;
  assign n2516 = n1050 ^ n442 ^ 1'b0 ;
  assign n2517 = n2448 & n2516 ;
  assign n2513 = n1818 ^ n971 ^ 1'b0 ;
  assign n2514 = ( n291 & n526 ) | ( n291 & ~n2513 ) | ( n526 & ~n2513 ) ;
  assign n2515 = n2514 ^ n2360 ^ x100 ;
  assign n2520 = n2519 ^ n2517 ^ n2515 ;
  assign n2533 = n2532 ^ n2520 ^ 1'b0 ;
  assign n2534 = n1364 & ~n2533 ;
  assign n2535 = ( n130 & ~n1104 ) | ( n130 & n2149 ) | ( ~n1104 & n2149 ) ;
  assign n2536 = n2535 ^ x75 ^ 1'b0 ;
  assign n2537 = n916 | n2536 ;
  assign n2538 = x64 & n1159 ;
  assign n2539 = n2538 ^ n404 ^ 1'b0 ;
  assign n2540 = ~n1118 & n2539 ;
  assign n2541 = n2540 ^ n1525 ^ 1'b0 ;
  assign n2542 = n1503 ^ n1132 ^ n414 ;
  assign n2543 = ( n490 & ~n615 ) | ( n490 & n2542 ) | ( ~n615 & n2542 ) ;
  assign n2544 = n2541 & n2543 ;
  assign n2545 = ( ~n919 & n1234 ) | ( ~n919 & n2544 ) | ( n1234 & n2544 ) ;
  assign n2546 = ( n629 & n710 ) | ( n629 & n2545 ) | ( n710 & n2545 ) ;
  assign n2547 = n1090 | n2546 ;
  assign n2548 = ( n227 & n939 ) | ( n227 & ~n1066 ) | ( n939 & ~n1066 ) ;
  assign n2549 = n2548 ^ n2016 ^ n752 ;
  assign n2550 = n853 ^ n695 ^ n156 ;
  assign n2551 = x67 & ~n667 ;
  assign n2552 = n2551 ^ n550 ^ 1'b0 ;
  assign n2553 = n380 | n2552 ;
  assign n2554 = ( n525 & n2550 ) | ( n525 & n2553 ) | ( n2550 & n2553 ) ;
  assign n2556 = n2038 ^ n1386 ^ 1'b0 ;
  assign n2555 = n1182 ^ n743 ^ 1'b0 ;
  assign n2557 = n2556 ^ n2555 ^ 1'b0 ;
  assign n2558 = x108 ^ x88 ^ 1'b0 ;
  assign n2559 = n343 & n2558 ;
  assign n2560 = ( n1903 & ~n2013 ) | ( n1903 & n2544 ) | ( ~n2013 & n2544 ) ;
  assign n2561 = n1708 & n2560 ;
  assign n2562 = ~n2559 & n2561 ;
  assign n2563 = n1633 ^ n421 ^ n346 ;
  assign n2564 = ( ~n508 & n590 ) | ( ~n508 & n1088 ) | ( n590 & n1088 ) ;
  assign n2565 = n2563 | n2564 ;
  assign n2566 = n246 & n2565 ;
  assign n2567 = n2566 ^ n2114 ^ 1'b0 ;
  assign n2570 = n2405 ^ n1972 ^ 1'b0 ;
  assign n2571 = n2570 ^ n2029 ^ n501 ;
  assign n2568 = n1782 ^ n1608 ^ n543 ;
  assign n2569 = n814 & n2568 ;
  assign n2572 = n2571 ^ n2569 ^ 1'b0 ;
  assign n2573 = ~n169 & n2572 ;
  assign n2574 = ~n2461 & n2573 ;
  assign n2575 = n2574 ^ n171 ^ 1'b0 ;
  assign n2576 = ( x117 & n753 ) | ( x117 & ~n1471 ) | ( n753 & ~n1471 ) ;
  assign n2577 = n2004 & ~n2053 ;
  assign n2578 = x75 & ~n2174 ;
  assign n2579 = ( n1188 & n2319 ) | ( n1188 & n2578 ) | ( n2319 & n2578 ) ;
  assign n2580 = ( n2576 & n2577 ) | ( n2576 & n2579 ) | ( n2577 & n2579 ) ;
  assign n2581 = n1611 ^ n510 ^ n464 ;
  assign n2582 = ( ~n501 & n2580 ) | ( ~n501 & n2581 ) | ( n2580 & n2581 ) ;
  assign n2585 = x24 | n637 ;
  assign n2586 = n2585 ^ n1466 ^ 1'b0 ;
  assign n2587 = n1096 & n2586 ;
  assign n2583 = ( n300 & n2109 ) | ( n300 & ~n2519 ) | ( n2109 & ~n2519 ) ;
  assign n2584 = n2583 ^ n2361 ^ 1'b0 ;
  assign n2588 = n2587 ^ n2584 ^ n1517 ;
  assign n2589 = n1947 ^ n315 ^ 1'b0 ;
  assign n2595 = n1316 ^ n792 ^ n472 ;
  assign n2594 = n631 & n1124 ;
  assign n2596 = n2595 ^ n2594 ^ 1'b0 ;
  assign n2597 = n1677 & ~n2596 ;
  assign n2598 = n2597 ^ n476 ^ 1'b0 ;
  assign n2599 = ( ~n869 & n911 ) | ( ~n869 & n2598 ) | ( n911 & n2598 ) ;
  assign n2591 = x15 & n1427 ;
  assign n2592 = n2591 ^ n474 ^ 1'b0 ;
  assign n2593 = n2592 ^ n1868 ^ n839 ;
  assign n2590 = ( x81 & n1492 ) | ( x81 & ~n1559 ) | ( n1492 & ~n1559 ) ;
  assign n2600 = n2599 ^ n2593 ^ n2590 ;
  assign n2601 = ( n434 & n2589 ) | ( n434 & ~n2600 ) | ( n2589 & ~n2600 ) ;
  assign n2602 = ( n2420 & ~n2588 ) | ( n2420 & n2601 ) | ( ~n2588 & n2601 ) ;
  assign n2603 = ( ~n933 & n1880 ) | ( ~n933 & n2405 ) | ( n1880 & n2405 ) ;
  assign n2604 = n1831 ^ n1448 ^ n738 ;
  assign n2605 = n2603 & n2604 ;
  assign n2606 = n2605 ^ n1005 ^ 1'b0 ;
  assign n2607 = ( n644 & ~n1003 ) | ( n644 & n2606 ) | ( ~n1003 & n2606 ) ;
  assign n2613 = n1455 & ~n2058 ;
  assign n2614 = n2613 ^ n1040 ^ 1'b0 ;
  assign n2612 = ( ~n659 & n1782 ) | ( ~n659 & n2107 ) | ( n1782 & n2107 ) ;
  assign n2608 = n148 ^ x100 ^ 1'b0 ;
  assign n2609 = n1005 ^ n986 ^ 1'b0 ;
  assign n2610 = ~n2608 & n2609 ;
  assign n2611 = n2353 & n2610 ;
  assign n2615 = n2614 ^ n2612 ^ n2611 ;
  assign n2616 = ( ~n857 & n1399 ) | ( ~n857 & n1972 ) | ( n1399 & n1972 ) ;
  assign n2617 = n1838 ^ n785 ^ 1'b0 ;
  assign n2618 = ~n518 & n2617 ;
  assign n2619 = n2010 ^ x34 ^ 1'b0 ;
  assign n2620 = ~n885 & n1322 ;
  assign n2621 = n466 & n2620 ;
  assign n2622 = n2621 ^ n1221 ^ 1'b0 ;
  assign n2623 = n2319 ^ n1916 ^ n1525 ;
  assign n2624 = ( n1050 & n1471 ) | ( n1050 & ~n2623 ) | ( n1471 & ~n2623 ) ;
  assign n2625 = ( n712 & n1654 ) | ( n712 & ~n2624 ) | ( n1654 & ~n2624 ) ;
  assign n2626 = ~n2059 & n2432 ;
  assign n2630 = n480 ^ n472 ^ 1'b0 ;
  assign n2631 = n600 | n2630 ;
  assign n2632 = n2631 ^ n2138 ^ n500 ;
  assign n2633 = n2632 ^ n1595 ^ n1557 ;
  assign n2628 = n1437 ^ n437 ^ x10 ;
  assign n2627 = n901 | n2013 ;
  assign n2629 = n2628 ^ n2627 ^ 1'b0 ;
  assign n2634 = n2633 ^ n2629 ^ n1237 ;
  assign n2635 = n2634 ^ n2061 ^ n223 ;
  assign n2636 = n2290 ^ n1122 ^ 1'b0 ;
  assign n2637 = x0 & ~n505 ;
  assign n2638 = ( n185 & ~n1004 ) | ( n185 & n2637 ) | ( ~n1004 & n2637 ) ;
  assign n2639 = n1620 & n2638 ;
  assign n2640 = ~n2636 & n2639 ;
  assign n2641 = n1144 ^ n542 ^ 1'b0 ;
  assign n2642 = ( n1132 & ~n1594 ) | ( n1132 & n1728 ) | ( ~n1594 & n1728 ) ;
  assign n2643 = n2642 ^ n2014 ^ n1694 ;
  assign n2644 = ( ~n667 & n2232 ) | ( ~n667 & n2643 ) | ( n2232 & n2643 ) ;
  assign n2645 = x21 & n2128 ;
  assign n2646 = n2645 ^ n1489 ^ 1'b0 ;
  assign n2647 = n2646 ^ x3 ^ 1'b0 ;
  assign n2648 = n2647 ^ n1862 ^ n1194 ;
  assign n2649 = n2648 ^ n1451 ^ 1'b0 ;
  assign n2658 = n2361 ^ n1051 ^ n566 ;
  assign n2651 = n2027 ^ x30 ^ 1'b0 ;
  assign n2652 = ~n230 & n2651 ;
  assign n2650 = n1303 & ~n1308 ;
  assign n2653 = n2652 ^ n2650 ^ 1'b0 ;
  assign n2654 = n907 | n2234 ;
  assign n2655 = n986 | n2654 ;
  assign n2656 = n710 & ~n2655 ;
  assign n2657 = ( ~n1196 & n2653 ) | ( ~n1196 & n2656 ) | ( n2653 & n2656 ) ;
  assign n2659 = n2658 ^ n2657 ^ 1'b0 ;
  assign n2660 = n557 | n2144 ;
  assign n2661 = n969 & n1474 ;
  assign n2662 = ( n348 & n1999 ) | ( n348 & n2138 ) | ( n1999 & n2138 ) ;
  assign n2663 = ( n808 & n2661 ) | ( n808 & ~n2662 ) | ( n2661 & ~n2662 ) ;
  assign n2664 = n1119 & n2663 ;
  assign n2665 = n2664 ^ n1789 ^ 1'b0 ;
  assign n2666 = ( ~n642 & n662 ) | ( ~n642 & n694 ) | ( n662 & n694 ) ;
  assign n2667 = n2666 ^ n2570 ^ n1395 ;
  assign n2668 = ~n973 & n1539 ;
  assign n2669 = ~x66 & n894 ;
  assign n2670 = n2669 ^ n1775 ^ 1'b0 ;
  assign n2671 = n200 | n787 ;
  assign n2672 = n1145 & n2671 ;
  assign n2673 = n2672 ^ n2336 ^ 1'b0 ;
  assign n2674 = n2334 ^ n1672 ^ 1'b0 ;
  assign n2675 = n821 & ~n1361 ;
  assign n2676 = n2675 ^ n667 ^ 1'b0 ;
  assign n2677 = ( n875 & ~n885 ) | ( n875 & n2676 ) | ( ~n885 & n2676 ) ;
  assign n2678 = ( ~n685 & n1221 ) | ( ~n685 & n2677 ) | ( n1221 & n2677 ) ;
  assign n2679 = n2678 ^ n561 ^ n242 ;
  assign n2680 = n454 ^ n335 ^ n314 ;
  assign n2681 = n2458 ^ n2241 ^ n1860 ;
  assign n2682 = ~n2680 & n2681 ;
  assign n2683 = ( n272 & n422 ) | ( n272 & ~n1353 ) | ( n422 & ~n1353 ) ;
  assign n2684 = n1717 ^ n626 ^ 1'b0 ;
  assign n2685 = n622 ^ n390 ^ 1'b0 ;
  assign n2686 = n501 & n2685 ;
  assign n2687 = ~x18 & n2686 ;
  assign n2697 = ( n244 & ~n790 ) | ( n244 & n846 ) | ( ~n790 & n846 ) ;
  assign n2698 = ( n151 & n346 ) | ( n151 & n2697 ) | ( n346 & n2697 ) ;
  assign n2696 = n1868 ^ n298 ^ n297 ;
  assign n2695 = n1503 ^ n129 ^ 1'b0 ;
  assign n2699 = n2698 ^ n2696 ^ n2695 ;
  assign n2700 = n2699 ^ n1647 ^ n1025 ;
  assign n2690 = ~n1143 & n2637 ;
  assign n2691 = n2690 ^ x123 ^ 1'b0 ;
  assign n2688 = n1348 ^ n929 ^ n168 ;
  assign n2689 = n2688 ^ n1401 ^ 1'b0 ;
  assign n2692 = n2691 ^ n2689 ^ n2184 ;
  assign n2693 = n786 | n2692 ;
  assign n2694 = n1099 & ~n2693 ;
  assign n2701 = n2700 ^ n2694 ^ n2467 ;
  assign n2702 = n1330 & n2701 ;
  assign n2703 = ( ~n1533 & n2687 ) | ( ~n1533 & n2702 ) | ( n2687 & n2702 ) ;
  assign n2706 = n1045 ^ n916 ^ 1'b0 ;
  assign n2704 = n291 | n697 ;
  assign n2705 = n1244 & ~n2704 ;
  assign n2707 = n2706 ^ n2705 ^ n1641 ;
  assign n2708 = ( ~n1407 & n1575 ) | ( ~n1407 & n2234 ) | ( n1575 & n2234 ) ;
  assign n2709 = ~n462 & n2708 ;
  assign n2710 = n2709 ^ n2390 ^ x55 ;
  assign n2711 = n2414 ^ n1454 ^ 1'b0 ;
  assign n2712 = ( n853 & n1079 ) | ( n853 & ~n2088 ) | ( n1079 & ~n2088 ) ;
  assign n2713 = n2712 ^ n1081 ^ 1'b0 ;
  assign n2714 = n2713 ^ n2048 ^ 1'b0 ;
  assign n2715 = n2086 ^ x56 ^ 1'b0 ;
  assign n2716 = n298 & n2715 ;
  assign n2725 = n1360 ^ n884 ^ n565 ;
  assign n2722 = n1316 ^ n372 ^ 1'b0 ;
  assign n2723 = n2722 ^ n2456 ^ n1190 ;
  assign n2724 = ( n1069 & n2509 ) | ( n1069 & n2723 ) | ( n2509 & n2723 ) ;
  assign n2719 = n1399 ^ n1184 ^ 1'b0 ;
  assign n2720 = n1706 & ~n2719 ;
  assign n2717 = n1531 ^ n729 ^ n162 ;
  assign n2718 = ( ~n206 & n568 ) | ( ~n206 & n2717 ) | ( n568 & n2717 ) ;
  assign n2721 = n2720 ^ n2718 ^ 1'b0 ;
  assign n2726 = n2725 ^ n2724 ^ n2721 ;
  assign n2727 = n368 & ~n1375 ;
  assign n2728 = ~n1902 & n2727 ;
  assign n2729 = n2535 | n2568 ;
  assign n2730 = n2729 ^ n1034 ^ 1'b0 ;
  assign n2731 = ( ~n559 & n2079 ) | ( ~n559 & n2730 ) | ( n2079 & n2730 ) ;
  assign n2732 = n2097 ^ n644 ^ 1'b0 ;
  assign n2733 = ~n1727 & n2732 ;
  assign n2734 = n1806 ^ n765 ^ n635 ;
  assign n2735 = n1288 | n2734 ;
  assign n2736 = n1040 & ~n2735 ;
  assign n2737 = n1404 | n2736 ;
  assign n2738 = n563 | n2737 ;
  assign n2739 = ( n1539 & n2560 ) | ( n1539 & ~n2738 ) | ( n2560 & ~n2738 ) ;
  assign n2740 = n1883 ^ n740 ^ n733 ;
  assign n2741 = n566 ^ x69 ^ x49 ;
  assign n2742 = n1903 ^ n1755 ^ 1'b0 ;
  assign n2743 = n2030 ^ n773 ^ n764 ;
  assign n2744 = n2743 ^ n1375 ^ n672 ;
  assign n2745 = ( ~n159 & n875 ) | ( ~n159 & n1041 ) | ( n875 & n1041 ) ;
  assign n2746 = ( n565 & n2009 ) | ( n565 & ~n2745 ) | ( n2009 & ~n2745 ) ;
  assign n2747 = ~n639 & n2418 ;
  assign n2748 = n2747 ^ n1375 ^ 1'b0 ;
  assign n2749 = ~n2746 & n2748 ;
  assign n2750 = ~n1677 & n2749 ;
  assign n2751 = n2744 & n2750 ;
  assign n2752 = ~n1221 & n1671 ;
  assign n2753 = n2752 ^ n673 ^ 1'b0 ;
  assign n2754 = ~n2751 & n2753 ;
  assign n2755 = x40 & n485 ;
  assign n2756 = n2755 ^ n551 ^ 1'b0 ;
  assign n2757 = ( ~n418 & n2275 ) | ( ~n418 & n2756 ) | ( n2275 & n2756 ) ;
  assign n2758 = n2361 ^ n360 ^ 1'b0 ;
  assign n2759 = n1470 & ~n2758 ;
  assign n2760 = n1785 ^ x101 ^ 1'b0 ;
  assign n2770 = n829 | n1972 ;
  assign n2761 = n1855 ^ n1285 ^ n435 ;
  assign n2762 = n466 & n2761 ;
  assign n2763 = n2762 ^ n1755 ^ 1'b0 ;
  assign n2764 = x109 & n2763 ;
  assign n2765 = n919 & n2764 ;
  assign n2766 = n1357 ^ n706 ^ 1'b0 ;
  assign n2767 = ~n2765 & n2766 ;
  assign n2768 = ~n2089 & n2767 ;
  assign n2769 = n2768 ^ n1068 ^ 1'b0 ;
  assign n2771 = n2770 ^ n2769 ^ n1862 ;
  assign n2772 = n2178 & n2771 ;
  assign n2773 = ( ~n1014 & n2760 ) | ( ~n1014 & n2772 ) | ( n2760 & n2772 ) ;
  assign n2774 = n788 | n1636 ;
  assign n2775 = n2774 ^ n1049 ^ 1'b0 ;
  assign n2776 = ( ~x34 & x72 ) | ( ~x34 & n1848 ) | ( x72 & n1848 ) ;
  assign n2777 = n1247 & n2776 ;
  assign n2778 = ( n1697 & n2775 ) | ( n1697 & n2777 ) | ( n2775 & n2777 ) ;
  assign n2779 = n756 ^ n142 ^ 1'b0 ;
  assign n2780 = n1791 | n2779 ;
  assign n2781 = n1286 & ~n2780 ;
  assign n2782 = n2209 | n2781 ;
  assign n2783 = ~n520 & n2782 ;
  assign n2784 = n795 ^ n469 ^ x59 ;
  assign n2785 = ( ~n1348 & n1847 ) | ( ~n1348 & n2784 ) | ( n1847 & n2784 ) ;
  assign n2786 = ( n372 & n730 ) | ( n372 & ~n2785 ) | ( n730 & ~n2785 ) ;
  assign n2787 = n2786 ^ n1373 ^ n1030 ;
  assign n2788 = n1393 ^ n692 ^ n501 ;
  assign n2789 = n2787 | n2788 ;
  assign n2790 = n1297 | n2789 ;
  assign n2791 = n2226 & ~n2790 ;
  assign n2792 = n2544 ^ n2172 ^ 1'b0 ;
  assign n2793 = n2109 | n2792 ;
  assign n2794 = n642 | n702 ;
  assign n2795 = n2794 ^ n2390 ^ n219 ;
  assign n2796 = ( n1928 & n2624 ) | ( n1928 & n2795 ) | ( n2624 & n2795 ) ;
  assign n2797 = ( x5 & x38 ) | ( x5 & ~n545 ) | ( x38 & ~n545 ) ;
  assign n2798 = n2797 ^ n1463 ^ n539 ;
  assign n2799 = n1182 | n2798 ;
  assign n2800 = n520 ^ n459 ^ 1'b0 ;
  assign n2801 = ~n275 & n2800 ;
  assign n2802 = ( n1119 & n2013 ) | ( n1119 & n2801 ) | ( n2013 & n2801 ) ;
  assign n2803 = ( n223 & n1268 ) | ( n223 & n2802 ) | ( n1268 & n2802 ) ;
  assign n2804 = n2803 ^ n2211 ^ n1442 ;
  assign n2805 = n849 ^ n505 ^ x72 ;
  assign n2806 = n1480 | n2805 ;
  assign n2807 = n1041 | n2806 ;
  assign n2813 = n1850 ^ n798 ^ n418 ;
  assign n2808 = ( ~n162 & n919 ) | ( ~n162 & n1043 ) | ( n919 & n1043 ) ;
  assign n2809 = n1550 ^ n1285 ^ 1'b0 ;
  assign n2810 = ~n2808 & n2809 ;
  assign n2811 = n2450 & n2810 ;
  assign n2812 = n2811 ^ n2398 ^ n1784 ;
  assign n2814 = n2813 ^ n2812 ^ 1'b0 ;
  assign n2815 = n2023 | n2814 ;
  assign n2816 = n1595 ^ n1034 ^ n830 ;
  assign n2817 = n2816 ^ n2624 ^ n150 ;
  assign n2818 = n1622 ^ x125 ^ 1'b0 ;
  assign n2819 = ~n362 & n2070 ;
  assign n2820 = n2819 ^ n2756 ^ n741 ;
  assign n2821 = n692 ^ n674 ^ 1'b0 ;
  assign n2822 = n155 & ~n2821 ;
  assign n2823 = ( x26 & n151 ) | ( x26 & ~n2822 ) | ( n151 & ~n2822 ) ;
  assign n2824 = n760 ^ n580 ^ 1'b0 ;
  assign n2831 = n243 | n510 ;
  assign n2832 = n2831 ^ n719 ^ 1'b0 ;
  assign n2833 = ( n1465 & n1620 ) | ( n1465 & ~n2832 ) | ( n1620 & ~n2832 ) ;
  assign n2828 = n1096 & ~n1304 ;
  assign n2825 = n198 & n1364 ;
  assign n2826 = n2825 ^ n680 ^ 1'b0 ;
  assign n2827 = n2826 ^ n2801 ^ n367 ;
  assign n2829 = n2828 ^ n2827 ^ 1'b0 ;
  assign n2830 = ~n2226 & n2829 ;
  assign n2834 = n2833 ^ n2830 ^ n265 ;
  assign n2836 = n441 & n815 ;
  assign n2837 = ~x66 & n2836 ;
  assign n2835 = n2446 ^ n1085 ^ n291 ;
  assign n2838 = n2837 ^ n2835 ^ n1081 ;
  assign n2839 = ( n2000 & ~n2834 ) | ( n2000 & n2838 ) | ( ~n2834 & n2838 ) ;
  assign n2840 = ( x44 & n633 ) | ( x44 & n1316 ) | ( n633 & n1316 ) ;
  assign n2841 = n2840 ^ n1593 ^ 1'b0 ;
  assign n2842 = ~n249 & n2841 ;
  assign n2843 = n2842 ^ n1870 ^ n1408 ;
  assign n2844 = ~n381 & n2631 ;
  assign n2845 = ( n1066 & ~n1526 ) | ( n1066 & n2844 ) | ( ~n1526 & n2844 ) ;
  assign n2846 = n2539 ^ x3 ^ 1'b0 ;
  assign n2847 = ~n646 & n2846 ;
  assign n2848 = n2847 ^ n810 ^ n288 ;
  assign n2849 = n2848 ^ n2446 ^ n2169 ;
  assign n2850 = ( ~n2570 & n2845 ) | ( ~n2570 & n2849 ) | ( n2845 & n2849 ) ;
  assign n2851 = n2850 ^ n1356 ^ x75 ;
  assign n2852 = x123 & n1269 ;
  assign n2853 = n2851 & n2852 ;
  assign n2854 = ~n1528 & n1782 ;
  assign n2855 = n747 & n2712 ;
  assign n2856 = n1619 & ~n2855 ;
  assign n2857 = n499 & n2856 ;
  assign n2858 = n147 & n2799 ;
  assign n2859 = n2857 & n2858 ;
  assign n2860 = ~n642 & n1188 ;
  assign n2866 = ( n591 & ~n1498 ) | ( n591 & n1543 ) | ( ~n1498 & n1543 ) ;
  assign n2862 = n1494 ^ n1066 ^ n570 ;
  assign n2863 = n2862 ^ n1143 ^ n950 ;
  assign n2861 = n1973 ^ n263 ^ 1'b0 ;
  assign n2864 = n2863 ^ n2861 ^ n2389 ;
  assign n2865 = n2864 ^ n1387 ^ 1'b0 ;
  assign n2867 = n2866 ^ n2865 ^ n1827 ;
  assign n2868 = n2734 ^ x39 ^ 1'b0 ;
  assign n2869 = n1045 | n2868 ;
  assign n2870 = n957 ^ n945 ^ 1'b0 ;
  assign n2871 = n2360 ^ n1624 ^ n880 ;
  assign n2872 = n2871 ^ n1281 ^ 1'b0 ;
  assign n2873 = ~n2870 & n2872 ;
  assign n2874 = n1209 | n2832 ;
  assign n2875 = n2874 ^ n1727 ^ 1'b0 ;
  assign n2876 = n1126 ^ n957 ^ n607 ;
  assign n2877 = n2876 ^ n2441 ^ 1'b0 ;
  assign n2878 = n2877 ^ n1391 ^ 1'b0 ;
  assign n2879 = n1011 ^ x36 ^ 1'b0 ;
  assign n2880 = ~n2331 & n2879 ;
  assign n2881 = n2880 ^ n641 ^ n145 ;
  assign n2882 = ( n527 & ~n1507 ) | ( n527 & n2490 ) | ( ~n1507 & n2490 ) ;
  assign n2883 = ~n2881 & n2882 ;
  assign n2891 = n1742 ^ n540 ^ x121 ;
  assign n2884 = n945 ^ n597 ^ n424 ;
  assign n2885 = n505 ^ n182 ^ 1'b0 ;
  assign n2886 = n1996 & ~n2885 ;
  assign n2887 = n2886 ^ n484 ^ 1'b0 ;
  assign n2888 = x73 & n2887 ;
  assign n2889 = ~n2884 & n2888 ;
  assign n2890 = n2889 ^ n1693 ^ n1034 ;
  assign n2892 = n2891 ^ n2890 ^ n824 ;
  assign n2893 = n2273 ^ n933 ^ 1'b0 ;
  assign n2894 = n203 | n248 ;
  assign n2895 = n2894 ^ n2880 ^ n957 ;
  assign n2896 = n2076 & n2712 ;
  assign n2897 = ~n1327 & n2896 ;
  assign n2898 = ( n1122 & n2405 ) | ( n1122 & n2541 ) | ( n2405 & n2541 ) ;
  assign n2899 = n1388 | n2898 ;
  assign n2900 = n2899 ^ n421 ^ 1'b0 ;
  assign n2901 = n244 & n653 ;
  assign n2902 = n2901 ^ n1683 ^ 1'b0 ;
  assign n2903 = n2902 ^ n1460 ^ n943 ;
  assign n2904 = n1450 ^ n1441 ^ n245 ;
  assign n2905 = n1247 ^ x64 ^ 1'b0 ;
  assign n2906 = n2905 ^ n1460 ^ n309 ;
  assign n2907 = n2745 ^ n1544 ^ n631 ;
  assign n2908 = ( n2904 & ~n2906 ) | ( n2904 & n2907 ) | ( ~n2906 & n2907 ) ;
  assign n2909 = n2680 ^ n933 ^ n292 ;
  assign n2910 = n1555 ^ n1288 ^ n189 ;
  assign n2911 = n2910 ^ n390 ^ 1'b0 ;
  assign n2912 = ( x30 & n2909 ) | ( x30 & n2911 ) | ( n2909 & n2911 ) ;
  assign n2913 = ( n197 & n763 ) | ( n197 & n1933 ) | ( n763 & n1933 ) ;
  assign n2914 = n2331 ^ n1914 ^ n1788 ;
  assign n2915 = n2914 ^ n2676 ^ n2373 ;
  assign n2916 = n1859 ^ n375 ^ 1'b0 ;
  assign n2917 = n291 ^ n185 ^ 1'b0 ;
  assign n2918 = n2917 ^ n1483 ^ 1'b0 ;
  assign n2919 = ( n849 & n1106 ) | ( n849 & ~n2744 ) | ( n1106 & ~n2744 ) ;
  assign n2920 = n428 & n611 ;
  assign n2921 = n2920 ^ n1839 ^ 1'b0 ;
  assign n2922 = n2921 ^ n898 ^ 1'b0 ;
  assign n2923 = x16 & n2922 ;
  assign n2924 = n2310 ^ n1859 ^ 1'b0 ;
  assign n2927 = ~n918 & n1074 ;
  assign n2928 = n2927 ^ n1225 ^ 1'b0 ;
  assign n2929 = n2928 ^ n2021 ^ n1600 ;
  assign n2925 = n159 | n2440 ;
  assign n2926 = n1742 & ~n2925 ;
  assign n2930 = n2929 ^ n2926 ^ n960 ;
  assign n2933 = n1475 ^ n131 ^ 1'b0 ;
  assign n2934 = n401 & ~n2933 ;
  assign n2931 = n530 ^ n324 ^ n264 ;
  assign n2932 = ( n356 & ~n606 ) | ( n356 & n2931 ) | ( ~n606 & n2931 ) ;
  assign n2935 = n2934 ^ n2932 ^ n2161 ;
  assign n2936 = x18 & n1391 ;
  assign n2937 = n2936 ^ n2197 ^ 1'b0 ;
  assign n2942 = n1610 ^ n436 ^ 1'b0 ;
  assign n2943 = n2510 | n2942 ;
  assign n2944 = ( ~n788 & n2056 ) | ( ~n788 & n2943 ) | ( n2056 & n2943 ) ;
  assign n2945 = n2944 ^ n678 ^ 1'b0 ;
  assign n2946 = n670 & n2945 ;
  assign n2947 = n2008 ^ n268 ^ 1'b0 ;
  assign n2948 = n2946 & ~n2947 ;
  assign n2938 = n527 ^ x93 ^ 1'b0 ;
  assign n2939 = n1346 | n2938 ;
  assign n2940 = n1151 & ~n2939 ;
  assign n2941 = ~n2584 & n2940 ;
  assign n2949 = n2948 ^ n2941 ^ 1'b0 ;
  assign n2950 = ( n484 & n577 ) | ( n484 & n763 ) | ( n577 & n763 ) ;
  assign n2951 = n2950 ^ n1157 ^ 1'b0 ;
  assign n2952 = ( n1763 & ~n2548 ) | ( n1763 & n2951 ) | ( ~n2548 & n2951 ) ;
  assign n2953 = n2641 & ~n2952 ;
  assign n2954 = n2953 ^ n1129 ^ 1'b0 ;
  assign n2955 = ( n934 & n1123 ) | ( n934 & n1654 ) | ( n1123 & n1654 ) ;
  assign n2956 = n1828 ^ n1313 ^ 1'b0 ;
  assign n2957 = ~n2955 & n2956 ;
  assign n2958 = n1134 & ~n1785 ;
  assign n2959 = ~n2957 & n2958 ;
  assign n2964 = ~n588 & n887 ;
  assign n2960 = n1908 ^ n1226 ^ n1219 ;
  assign n2961 = n2960 ^ n2634 ^ n757 ;
  assign n2962 = n2782 ^ n746 ^ 1'b0 ;
  assign n2963 = ( ~n2569 & n2961 ) | ( ~n2569 & n2962 ) | ( n2961 & n2962 ) ;
  assign n2965 = n2964 ^ n2963 ^ n2628 ;
  assign n2966 = n1282 ^ n1008 ^ 1'b0 ;
  assign n2967 = n999 | n2966 ;
  assign n2968 = n645 | n1144 ;
  assign n2969 = ( ~n610 & n1212 ) | ( ~n610 & n2968 ) | ( n1212 & n2968 ) ;
  assign n2970 = ( n179 & ~n890 ) | ( n179 & n1644 ) | ( ~n890 & n1644 ) ;
  assign n2971 = x30 & ~n1370 ;
  assign n2972 = n1132 & n2971 ;
  assign n2973 = ( ~x24 & n1749 ) | ( ~x24 & n2972 ) | ( n1749 & n2972 ) ;
  assign n2974 = n1174 ^ n412 ^ 1'b0 ;
  assign n2975 = n796 & ~n2974 ;
  assign n2976 = n2973 & n2975 ;
  assign n2977 = n2976 ^ n2833 ^ 1'b0 ;
  assign n2978 = n2970 & ~n2977 ;
  assign n2979 = n2969 & n2978 ;
  assign n2980 = n2967 & n2979 ;
  assign n2981 = n2980 ^ n2010 ^ n1015 ;
  assign n2982 = ( n442 & n2144 ) | ( n442 & ~n2917 ) | ( n2144 & ~n2917 ) ;
  assign n2983 = ( x35 & ~n187 ) | ( x35 & n265 ) | ( ~n187 & n265 ) ;
  assign n2984 = n519 & ~n551 ;
  assign n2985 = ~n282 & n2984 ;
  assign n2986 = x116 & ~n2985 ;
  assign n2987 = n2983 & n2986 ;
  assign n2988 = n2472 & ~n2987 ;
  assign n2989 = n2982 & n2988 ;
  assign n2990 = ~n265 & n883 ;
  assign n2991 = n2990 ^ x53 ^ 1'b0 ;
  assign n2992 = n2991 ^ n919 ^ 1'b0 ;
  assign n2993 = ( n969 & n2020 ) | ( n969 & n2313 ) | ( n2020 & n2313 ) ;
  assign n2994 = n2993 ^ n1547 ^ n700 ;
  assign n2995 = x39 & ~n2994 ;
  assign n2996 = n2995 ^ n1329 ^ 1'b0 ;
  assign n2997 = ~n294 & n2283 ;
  assign n2998 = n2997 ^ n1786 ^ 1'b0 ;
  assign n2999 = n637 | n2998 ;
  assign n3000 = ~n2475 & n2999 ;
  assign n3001 = n1286 & n3000 ;
  assign n3002 = ( n1612 & n1697 ) | ( n1612 & ~n2299 ) | ( n1697 & ~n2299 ) ;
  assign n3003 = n368 & ~n2527 ;
  assign n3004 = n3003 ^ n1709 ^ 1'b0 ;
  assign n3005 = n1960 | n2069 ;
  assign n3006 = n3004 | n3005 ;
  assign n3007 = n2087 & ~n2468 ;
  assign n3008 = ( n3002 & ~n3006 ) | ( n3002 & n3007 ) | ( ~n3006 & n3007 ) ;
  assign n3009 = n245 | n2027 ;
  assign n3010 = ~n2070 & n3009 ;
  assign n3011 = n3010 ^ n2926 ^ 1'b0 ;
  assign n3012 = ( n185 & ~n189 ) | ( n185 & n284 ) | ( ~n189 & n284 ) ;
  assign n3013 = n3012 ^ x61 ^ 1'b0 ;
  assign n3014 = n1603 ^ n1513 ^ n1275 ;
  assign n3015 = n3014 ^ n2793 ^ 1'b0 ;
  assign n3016 = n1311 & ~n1901 ;
  assign n3017 = n512 & ~n1856 ;
  assign n3018 = n3017 ^ n746 ^ 1'b0 ;
  assign n3019 = ( n1841 & n3016 ) | ( n1841 & ~n3018 ) | ( n3016 & ~n3018 ) ;
  assign n3020 = n252 ^ x84 ^ 1'b0 ;
  assign n3021 = n740 | n3020 ;
  assign n3022 = ( ~n270 & n2692 ) | ( ~n270 & n3021 ) | ( n2692 & n3021 ) ;
  assign n3026 = ( n177 & n493 ) | ( n177 & n2763 ) | ( n493 & n2763 ) ;
  assign n3027 = ~n1648 & n2230 ;
  assign n3028 = ( ~n1192 & n3026 ) | ( ~n1192 & n3027 ) | ( n3026 & n3027 ) ;
  assign n3023 = ( n1441 & ~n1964 ) | ( n1441 & n2756 ) | ( ~n1964 & n2756 ) ;
  assign n3024 = ( n951 & ~n960 ) | ( n951 & n2526 ) | ( ~n960 & n2526 ) ;
  assign n3025 = n3023 | n3024 ;
  assign n3029 = n3028 ^ n3025 ^ 1'b0 ;
  assign n3030 = n2112 ^ n1609 ^ 1'b0 ;
  assign n3031 = ( x32 & n620 ) | ( x32 & ~n2418 ) | ( n620 & ~n2418 ) ;
  assign n3032 = ~n3030 & n3031 ;
  assign n3033 = n3032 ^ n2470 ^ 1'b0 ;
  assign n3034 = n1585 & n3033 ;
  assign n3035 = n3034 ^ n1808 ^ 1'b0 ;
  assign n3036 = n1960 ^ n468 ^ x98 ;
  assign n3037 = n598 & ~n3036 ;
  assign n3038 = n3037 ^ x117 ^ 1'b0 ;
  assign n3039 = n3035 & n3038 ;
  assign n3040 = n1226 ^ n854 ^ 1'b0 ;
  assign n3041 = n2063 | n3040 ;
  assign n3042 = ~n800 & n2767 ;
  assign n3043 = ( n138 & ~n3041 ) | ( n138 & n3042 ) | ( ~n3041 & n3042 ) ;
  assign n3044 = n2053 ^ n368 ^ n286 ;
  assign n3045 = n3044 ^ n2769 ^ n375 ;
  assign n3046 = n2490 ^ n878 ^ n248 ;
  assign n3047 = n3046 ^ n1725 ^ n288 ;
  assign n3053 = ( ~n226 & n933 ) | ( ~n226 & n1376 ) | ( n933 & n1376 ) ;
  assign n3054 = n3053 ^ n1257 ^ n378 ;
  assign n3048 = n1225 ^ n297 ^ n215 ;
  assign n3049 = ( ~n302 & n934 ) | ( ~n302 & n2176 ) | ( n934 & n2176 ) ;
  assign n3050 = n3049 ^ n2485 ^ n2179 ;
  assign n3051 = n3050 ^ n927 ^ n162 ;
  assign n3052 = n3048 & n3051 ;
  assign n3055 = n3054 ^ n3052 ^ 1'b0 ;
  assign n3056 = n3055 ^ n967 ^ 1'b0 ;
  assign n3057 = ~n849 & n3056 ;
  assign n3058 = ~n1024 & n1554 ;
  assign n3059 = n3058 ^ n531 ^ 1'b0 ;
  assign n3061 = n2239 ^ n1629 ^ n710 ;
  assign n3062 = ( n976 & ~n1129 ) | ( n976 & n3061 ) | ( ~n1129 & n3061 ) ;
  assign n3060 = n1091 | n2066 ;
  assign n3063 = n3062 ^ n3060 ^ 1'b0 ;
  assign n3064 = n3063 ^ n2520 ^ n1657 ;
  assign n3069 = n378 & ~n2541 ;
  assign n3070 = n3069 ^ n777 ^ 1'b0 ;
  assign n3066 = n489 & ~n884 ;
  assign n3067 = ~n383 & n3066 ;
  assign n3068 = n3067 ^ n2013 ^ n1601 ;
  assign n3071 = n3070 ^ n3068 ^ n512 ;
  assign n3065 = n553 | n584 ;
  assign n3072 = n3071 ^ n3065 ^ n2847 ;
  assign n3073 = n2736 ^ n553 ^ x119 ;
  assign n3074 = n3073 ^ n230 ^ 1'b0 ;
  assign n3075 = ( ~n874 & n1050 ) | ( ~n874 & n1949 ) | ( n1050 & n1949 ) ;
  assign n3076 = n1247 & n2411 ;
  assign n3077 = n3076 ^ n2418 ^ n591 ;
  assign n3078 = ( n408 & n3075 ) | ( n408 & n3077 ) | ( n3075 & n3077 ) ;
  assign n3079 = n281 | n3078 ;
  assign n3080 = n1674 ^ x66 ^ x24 ;
  assign n3081 = n200 & ~n988 ;
  assign n3082 = n1688 ^ n1122 ^ n1104 ;
  assign n3083 = ( n1361 & n3081 ) | ( n1361 & ~n3082 ) | ( n3081 & ~n3082 ) ;
  assign n3084 = ( ~x40 & n3080 ) | ( ~x40 & n3083 ) | ( n3080 & n3083 ) ;
  assign n3085 = n2428 ^ n1749 ^ n672 ;
  assign n3086 = n1649 ^ n1049 ^ n605 ;
  assign n3087 = n3085 & n3086 ;
  assign n3088 = n461 & n1203 ;
  assign n3089 = n2179 ^ n1997 ^ n1050 ;
  assign n3090 = n2392 | n3089 ;
  assign n3091 = n2930 | n3090 ;
  assign n3092 = n1451 ^ n624 ^ 1'b0 ;
  assign n3093 = ~n541 & n1021 ;
  assign n3094 = n3093 ^ x33 ^ 1'b0 ;
  assign n3095 = n973 & ~n1090 ;
  assign n3096 = ~x46 & n3095 ;
  assign n3097 = ( n1530 & n2415 ) | ( n1530 & n3096 ) | ( n2415 & n3096 ) ;
  assign n3098 = ( n1606 & n1612 ) | ( n1606 & n3097 ) | ( n1612 & n3097 ) ;
  assign n3099 = n3098 ^ n2620 ^ n766 ;
  assign n3100 = ~n230 & n705 ;
  assign n3101 = n366 & n3100 ;
  assign n3102 = n3101 ^ n2760 ^ 1'b0 ;
  assign n3103 = n3102 ^ n1287 ^ 1'b0 ;
  assign n3106 = ( n415 & n1355 ) | ( n415 & n2577 ) | ( n1355 & n2577 ) ;
  assign n3107 = n3106 ^ n2411 ^ 1'b0 ;
  assign n3104 = x100 & ~n438 ;
  assign n3105 = n3104 ^ n964 ^ 1'b0 ;
  assign n3108 = n3107 ^ n3105 ^ n305 ;
  assign n3116 = n1955 | n2296 ;
  assign n3117 = n3116 ^ n612 ^ 1'b0 ;
  assign n3111 = ( x18 & n390 ) | ( x18 & ~n1327 ) | ( n390 & ~n1327 ) ;
  assign n3112 = n3111 ^ n886 ^ 1'b0 ;
  assign n3113 = n2609 & ~n3112 ;
  assign n3109 = ( ~n896 & n2184 ) | ( ~n896 & n2402 ) | ( n2184 & n2402 ) ;
  assign n3110 = n3109 ^ n2147 ^ x19 ;
  assign n3114 = n3113 ^ n3110 ^ n1774 ;
  assign n3115 = ( ~n461 & n644 ) | ( ~n461 & n3114 ) | ( n644 & n3114 ) ;
  assign n3118 = n3117 ^ n3115 ^ 1'b0 ;
  assign n3119 = n1777 & n1955 ;
  assign n3120 = ~x80 & n1050 ;
  assign n3121 = n2519 | n3023 ;
  assign n3124 = ( ~n438 & n1514 ) | ( ~n438 & n1706 ) | ( n1514 & n1706 ) ;
  assign n3125 = ( n245 & ~n2122 ) | ( n245 & n3124 ) | ( ~n2122 & n3124 ) ;
  assign n3122 = n1978 ^ n1050 ^ x10 ;
  assign n3123 = n3122 ^ n1958 ^ n440 ;
  assign n3126 = n3125 ^ n3123 ^ n894 ;
  assign n3127 = n1123 & ~n1788 ;
  assign n3128 = n3127 ^ x19 ^ 1'b0 ;
  assign n3129 = n2313 & ~n3128 ;
  assign n3130 = n1334 & ~n1894 ;
  assign n3131 = ~n151 & n3130 ;
  assign n3132 = n2553 | n3131 ;
  assign n3133 = n3132 ^ n2060 ^ 1'b0 ;
  assign n3134 = ( x121 & ~n351 ) | ( x121 & n2440 ) | ( ~n351 & n2440 ) ;
  assign n3135 = n3134 ^ n543 ^ 1'b0 ;
  assign n3136 = n1832 | n2603 ;
  assign n3137 = ( n2931 & ~n3135 ) | ( n2931 & n3136 ) | ( ~n3135 & n3136 ) ;
  assign n3141 = n2301 ^ n1199 ^ n230 ;
  assign n3138 = n692 | n2677 ;
  assign n3139 = n376 | n3138 ;
  assign n3140 = n166 | n3139 ;
  assign n3142 = n3141 ^ n3140 ^ 1'b0 ;
  assign n3147 = ( x32 & n1090 ) | ( x32 & n2390 ) | ( n1090 & n2390 ) ;
  assign n3148 = ( n179 & n1655 ) | ( n179 & ~n3147 ) | ( n1655 & ~n3147 ) ;
  assign n3146 = n1592 & ~n1758 ;
  assign n3149 = n3148 ^ n3146 ^ n2689 ;
  assign n3143 = n246 & ~n813 ;
  assign n3144 = ~n2006 & n3143 ;
  assign n3145 = n3144 ^ n3122 ^ n1424 ;
  assign n3150 = n3149 ^ n3145 ^ n677 ;
  assign n3151 = ( n279 & ~n1307 ) | ( n279 & n2604 ) | ( ~n1307 & n2604 ) ;
  assign n3152 = n1713 ^ n1114 ^ 1'b0 ;
  assign n3153 = ~n3151 & n3152 ;
  assign n3154 = ~n3150 & n3153 ;
  assign n3155 = n429 ^ x68 ^ 1'b0 ;
  assign n3156 = ~n508 & n3155 ;
  assign n3157 = n3156 ^ n891 ^ n375 ;
  assign n3160 = n1958 ^ x93 ^ x65 ;
  assign n3158 = ~n1139 & n1619 ;
  assign n3159 = ~n550 & n3158 ;
  assign n3161 = n3160 ^ n3159 ^ n2564 ;
  assign n3162 = n728 & ~n1720 ;
  assign n3163 = n177 | n533 ;
  assign n3164 = x50 & ~n973 ;
  assign n3165 = n3164 ^ n3086 ^ n2996 ;
  assign n3166 = n3058 ^ n2398 ^ 1'b0 ;
  assign n3167 = ( n887 & n2349 ) | ( n887 & ~n3166 ) | ( n2349 & ~n3166 ) ;
  assign n3181 = x78 & n1749 ;
  assign n3182 = n1179 & n3181 ;
  assign n3168 = ~n1755 & n2114 ;
  assign n3169 = n3168 ^ n282 ^ 1'b0 ;
  assign n3174 = ( n1059 & n1090 ) | ( n1059 & n1316 ) | ( n1090 & n1316 ) ;
  assign n3170 = n1369 & n1719 ;
  assign n3171 = n3170 ^ n1015 ^ 1'b0 ;
  assign n3172 = n484 & ~n3171 ;
  assign n3173 = n3172 ^ n1126 ^ 1'b0 ;
  assign n3175 = n3174 ^ n3173 ^ n413 ;
  assign n3176 = n3175 ^ n2582 ^ n2048 ;
  assign n3177 = n2025 ^ n1662 ^ n752 ;
  assign n3178 = ~n1432 & n3177 ;
  assign n3179 = n3178 ^ n609 ^ 1'b0 ;
  assign n3180 = ( n3169 & n3176 ) | ( n3169 & ~n3179 ) | ( n3176 & ~n3179 ) ;
  assign n3183 = n3182 ^ n3180 ^ n332 ;
  assign n3184 = n526 & ~n970 ;
  assign n3185 = ~n767 & n2934 ;
  assign n3186 = ~n3184 & n3185 ;
  assign n3187 = n1791 ^ n1463 ^ n531 ;
  assign n3188 = n576 | n1555 ;
  assign n3189 = n703 & n1901 ;
  assign n3190 = ( n3187 & n3188 ) | ( n3187 & n3189 ) | ( n3188 & n3189 ) ;
  assign n3191 = n481 ^ n257 ^ 1'b0 ;
  assign n3192 = n2635 & n3191 ;
  assign n3193 = ~n199 & n3192 ;
  assign n3194 = n1439 & n1554 ;
  assign n3195 = n3194 ^ n2431 ^ n1239 ;
  assign n3196 = n2006 & ~n2612 ;
  assign n3198 = n1752 ^ n1706 ^ x100 ;
  assign n3197 = ( n999 & n1164 ) | ( n999 & ~n1301 ) | ( n1164 & ~n1301 ) ;
  assign n3199 = n3198 ^ n3197 ^ 1'b0 ;
  assign n3200 = n683 | n3199 ;
  assign n3201 = ( n3195 & n3196 ) | ( n3195 & ~n3200 ) | ( n3196 & ~n3200 ) ;
  assign n3202 = ( n1603 & n3193 ) | ( n1603 & ~n3201 ) | ( n3193 & ~n3201 ) ;
  assign n3203 = ( ~n322 & n426 ) | ( ~n322 & n612 ) | ( n426 & n612 ) ;
  assign n3204 = n1865 & n3203 ;
  assign n3205 = n3020 ^ n2168 ^ n330 ;
  assign n3206 = n1991 ^ n1697 ^ n584 ;
  assign n3207 = ( x103 & n964 ) | ( x103 & ~n1731 ) | ( n964 & ~n1731 ) ;
  assign n3208 = n1394 ^ n343 ^ 1'b0 ;
  assign n3209 = n1665 | n3208 ;
  assign n3210 = n3209 ^ n2772 ^ n731 ;
  assign n3211 = ~n786 & n2661 ;
  assign n3212 = n399 & n3211 ;
  assign n3213 = n2570 ^ n770 ^ 1'b0 ;
  assign n3214 = n1108 & n3213 ;
  assign n3215 = ~n3212 & n3214 ;
  assign n3216 = ( ~n1741 & n3007 ) | ( ~n1741 & n3215 ) | ( n3007 & n3215 ) ;
  assign n3217 = n414 ^ n259 ^ 1'b0 ;
  assign n3219 = n824 & n1294 ;
  assign n3220 = n3219 ^ n1251 ^ 1'b0 ;
  assign n3218 = n2298 ^ n2284 ^ n1908 ;
  assign n3221 = n3220 ^ n3218 ^ n1555 ;
  assign n3222 = ( ~n541 & n3217 ) | ( ~n541 & n3221 ) | ( n3217 & n3221 ) ;
  assign n3235 = n2249 ^ n2012 ^ n1959 ;
  assign n3236 = n3235 ^ n2863 ^ 1'b0 ;
  assign n3224 = n264 ^ x102 ^ 1'b0 ;
  assign n3225 = n1151 | n3224 ;
  assign n3226 = n1034 | n1823 ;
  assign n3227 = n1179 & ~n3226 ;
  assign n3228 = n1871 | n3227 ;
  assign n3229 = n2329 | n3228 ;
  assign n3230 = ( n1308 & ~n2355 ) | ( n1308 & n3113 ) | ( ~n2355 & n3113 ) ;
  assign n3231 = n3229 & n3230 ;
  assign n3232 = n3225 | n3231 ;
  assign n3233 = n2071 | n3232 ;
  assign n3234 = n509 | n3233 ;
  assign n3237 = n3236 ^ n3234 ^ 1'b0 ;
  assign n3223 = n2360 & n2459 ;
  assign n3238 = n3237 ^ n3223 ^ 1'b0 ;
  assign n3239 = n145 & ~n730 ;
  assign n3240 = n3239 ^ n854 ^ 1'b0 ;
  assign n3241 = n3240 ^ n2317 ^ 1'b0 ;
  assign n3242 = n2087 ^ n2052 ^ n1800 ;
  assign n3243 = ~n673 & n1434 ;
  assign n3244 = n625 | n3243 ;
  assign n3245 = n3244 ^ n636 ^ 1'b0 ;
  assign n3246 = n3240 ^ n1814 ^ 1'b0 ;
  assign n3247 = n291 | n3246 ;
  assign n3250 = x126 & n1483 ;
  assign n3251 = n3250 ^ n1133 ^ 1'b0 ;
  assign n3252 = ( n187 & ~n2258 ) | ( n187 & n3251 ) | ( ~n2258 & n3251 ) ;
  assign n3248 = x21 & x85 ;
  assign n3249 = n2150 | n3248 ;
  assign n3253 = n3252 ^ n3249 ^ n1646 ;
  assign n3254 = ( n285 & n3247 ) | ( n285 & n3253 ) | ( n3247 & n3253 ) ;
  assign n3255 = ( n243 & n786 ) | ( n243 & n1547 ) | ( n786 & n1547 ) ;
  assign n3256 = ( n1164 & n2940 ) | ( n1164 & n3255 ) | ( n2940 & n3255 ) ;
  assign n3257 = n2314 ^ n2283 ^ 1'b0 ;
  assign n3258 = n3161 ^ n2542 ^ x13 ;
  assign n3260 = n3124 ^ n1837 ^ n376 ;
  assign n3259 = n998 | n1816 ;
  assign n3261 = n3260 ^ n3259 ^ 1'b0 ;
  assign n3262 = n2809 ^ n996 ^ 1'b0 ;
  assign n3263 = n1180 & ~n1917 ;
  assign n3264 = n2481 ^ n2468 ^ n1594 ;
  assign n3265 = ( ~n778 & n1638 ) | ( ~n778 & n1699 ) | ( n1638 & n1699 ) ;
  assign n3266 = n1106 & n3265 ;
  assign n3267 = n3266 ^ n3041 ^ 1'b0 ;
  assign n3268 = n201 & ~n2808 ;
  assign n3269 = ( n620 & n1715 ) | ( n620 & n3268 ) | ( n1715 & n3268 ) ;
  assign n3270 = ( n2413 & ~n3081 ) | ( n2413 & n3269 ) | ( ~n3081 & n3269 ) ;
  assign n3271 = ~n849 & n945 ;
  assign n3272 = n3271 ^ n1025 ^ 1'b0 ;
  assign n3273 = n3272 ^ n480 ^ n220 ;
  assign n3274 = n3273 ^ n164 ^ 1'b0 ;
  assign n3279 = n1674 & ~n3272 ;
  assign n3280 = n529 & n3279 ;
  assign n3278 = n2446 ^ n2370 ^ 1'b0 ;
  assign n3275 = n1548 ^ n775 ^ n565 ;
  assign n3276 = n407 & ~n3275 ;
  assign n3277 = ~n2105 & n3276 ;
  assign n3281 = n3280 ^ n3278 ^ n3277 ;
  assign n3282 = n2747 ^ n2356 ^ n1677 ;
  assign n3283 = n3282 ^ n1507 ^ 1'b0 ;
  assign n3284 = n3281 & n3283 ;
  assign n3285 = ( n177 & ~n3274 ) | ( n177 & n3284 ) | ( ~n3274 & n3284 ) ;
  assign n3286 = n2940 ^ n1970 ^ n377 ;
  assign n3287 = n3286 ^ n3217 ^ 1'b0 ;
  assign n3288 = ~n624 & n1674 ;
  assign n3289 = ( n974 & ~n1068 ) | ( n974 & n3288 ) | ( ~n1068 & n3288 ) ;
  assign n3290 = n2723 ^ n1517 ^ 1'b0 ;
  assign n3291 = n3289 & n3290 ;
  assign n3292 = ( n2805 & ~n3179 ) | ( n2805 & n3291 ) | ( ~n3179 & n3291 ) ;
  assign n3296 = n220 & ~n302 ;
  assign n3297 = n1945 & n3296 ;
  assign n3295 = n2902 ^ n1429 ^ 1'b0 ;
  assign n3293 = n2948 ^ n840 ^ n536 ;
  assign n3294 = n3293 ^ n2267 ^ n2030 ;
  assign n3298 = n3297 ^ n3295 ^ n3294 ;
  assign n3299 = n3169 ^ n2532 ^ 1'b0 ;
  assign n3300 = ~n657 & n3175 ;
  assign n3301 = ~n770 & n3300 ;
  assign n3302 = n288 & ~n813 ;
  assign n3303 = ~n2289 & n3302 ;
  assign n3304 = n3171 ^ n1448 ^ 1'b0 ;
  assign n3305 = n2283 & n3304 ;
  assign n3306 = n1219 & n3305 ;
  assign n3307 = n3306 ^ n2635 ^ 1'b0 ;
  assign n3308 = n1741 ^ x36 ^ 1'b0 ;
  assign n3309 = n1541 | n3308 ;
  assign n3310 = n717 & ~n3309 ;
  assign n3311 = ~n3099 & n3310 ;
  assign n3312 = ( n169 & n1288 ) | ( n169 & n1399 ) | ( n1288 & n1399 ) ;
  assign n3313 = n3312 ^ n380 ^ 1'b0 ;
  assign n3314 = ~n3311 & n3313 ;
  assign n3315 = n710 ^ n264 ^ 1'b0 ;
  assign n3316 = n659 | n3315 ;
  assign n3317 = ~x68 & n3316 ;
  assign n3318 = n3317 ^ n1666 ^ n1306 ;
  assign n3319 = ( x25 & ~n2655 ) | ( x25 & n3318 ) | ( ~n2655 & n3318 ) ;
  assign n3320 = ( ~n1764 & n2043 ) | ( ~n1764 & n3319 ) | ( n2043 & n3319 ) ;
  assign n3321 = ~n1001 & n1263 ;
  assign n3322 = n774 | n3321 ;
  assign n3323 = n2167 & n3322 ;
  assign n3325 = n2197 ^ n1409 ^ n441 ;
  assign n3324 = n624 & n1459 ;
  assign n3326 = n3325 ^ n3324 ^ 1'b0 ;
  assign n3327 = n903 | n3326 ;
  assign n3328 = n1902 | n3327 ;
  assign n3329 = ( x2 & ~n1030 ) | ( x2 & n2197 ) | ( ~n1030 & n2197 ) ;
  assign n3330 = n3329 ^ n1636 ^ n1048 ;
  assign n3331 = n3319 ^ n3118 ^ 1'b0 ;
  assign n3332 = n887 & ~n1816 ;
  assign n3333 = n3332 ^ n388 ^ 1'b0 ;
  assign n3334 = ( ~n2279 & n2614 ) | ( ~n2279 & n3333 ) | ( n2614 & n3333 ) ;
  assign n3335 = n1193 | n3334 ;
  assign n3336 = ( n213 & ~n980 ) | ( n213 & n2324 ) | ( ~n980 & n2324 ) ;
  assign n3337 = n3336 ^ n1407 ^ 1'b0 ;
  assign n3338 = ( n391 & n891 ) | ( n391 & n1018 ) | ( n891 & n1018 ) ;
  assign n3339 = n1624 ^ n1477 ^ n203 ;
  assign n3340 = n607 & n1653 ;
  assign n3341 = n1725 & n3340 ;
  assign n3342 = n3339 & ~n3341 ;
  assign n3343 = ~n3338 & n3342 ;
  assign n3344 = ( n2397 & ~n3249 ) | ( n2397 & n3343 ) | ( ~n3249 & n3343 ) ;
  assign n3345 = ( x42 & n465 ) | ( x42 & ~n1950 ) | ( n465 & ~n1950 ) ;
  assign n3346 = n3345 ^ n2763 ^ n198 ;
  assign n3347 = n302 & ~n673 ;
  assign n3348 = n3346 | n3347 ;
  assign n3349 = n2772 | n3348 ;
  assign n3350 = n2521 & n3349 ;
  assign n3351 = n3344 & n3350 ;
  assign n3352 = ( x80 & n712 ) | ( x80 & n3234 ) | ( n712 & n3234 ) ;
  assign n3353 = n2628 ^ n1136 ^ 1'b0 ;
  assign n3354 = n1481 | n3353 ;
  assign n3355 = n839 & ~n1234 ;
  assign n3356 = n3354 & n3355 ;
  assign n3357 = n1946 | n3059 ;
  assign n3358 = n2315 ^ n2307 ^ n2183 ;
  assign n3359 = n1841 | n1976 ;
  assign n3360 = n3359 ^ n2967 ^ n271 ;
  assign n3361 = n3360 ^ n1119 ^ 1'b0 ;
  assign n3362 = n3358 | n3361 ;
  assign n3367 = n954 & n2576 ;
  assign n3368 = n345 & n3367 ;
  assign n3369 = n3068 & n3368 ;
  assign n3364 = n1752 ^ n1403 ^ 1'b0 ;
  assign n3365 = n1005 & ~n3364 ;
  assign n3363 = n1180 ^ n551 ^ n302 ;
  assign n3366 = n3365 ^ n3363 ^ n2056 ;
  assign n3370 = n3369 ^ n3366 ^ n1968 ;
  assign n3371 = n3141 ^ x4 ^ 1'b0 ;
  assign n3372 = n2150 ^ n1010 ^ n536 ;
  assign n3373 = n240 & n3372 ;
  assign n3374 = n3373 ^ n1068 ^ 1'b0 ;
  assign n3375 = n3374 ^ n3297 ^ 1'b0 ;
  assign n3376 = n1225 & n2611 ;
  assign n3377 = n1788 | n3376 ;
  assign n3378 = n2176 ^ n1610 ^ n631 ;
  assign n3379 = ( ~n259 & n672 ) | ( ~n259 & n3378 ) | ( n672 & n3378 ) ;
  assign n3380 = n1450 ^ n1357 ^ 1'b0 ;
  assign n3381 = n3379 | n3380 ;
  assign n3382 = n673 | n3030 ;
  assign n3383 = n234 & ~n1076 ;
  assign n3384 = n3382 & ~n3383 ;
  assign n3385 = n1020 & ~n3384 ;
  assign n3386 = ( n3377 & n3381 ) | ( n3377 & ~n3385 ) | ( n3381 & ~n3385 ) ;
  assign n3388 = n924 & ~n2955 ;
  assign n3389 = n3388 ^ n829 ^ 1'b0 ;
  assign n3387 = n2131 | n2749 ;
  assign n3390 = n3389 ^ n3387 ^ 1'b0 ;
  assign n3391 = n3389 ^ n1362 ^ x89 ;
  assign n3392 = n3107 ^ n562 ^ 1'b0 ;
  assign n3393 = ( n1977 & ~n3031 ) | ( n1977 & n3392 ) | ( ~n3031 & n3392 ) ;
  assign n3397 = n244 | n300 ;
  assign n3398 = n3397 ^ x84 ^ 1'b0 ;
  assign n3396 = x122 & n823 ;
  assign n3399 = n3398 ^ n3396 ^ 1'b0 ;
  assign n3394 = ~n972 & n1844 ;
  assign n3395 = n639 & n3394 ;
  assign n3400 = n3399 ^ n3395 ^ n1962 ;
  assign n3401 = n3400 ^ n2402 ^ n1393 ;
  assign n3403 = ~n994 & n1006 ;
  assign n3404 = n3403 ^ n2151 ^ 1'b0 ;
  assign n3402 = n1976 ^ n822 ^ 1'b0 ;
  assign n3405 = n3404 ^ n3402 ^ n2106 ;
  assign n3406 = n3405 ^ n2306 ^ n879 ;
  assign n3407 = ( n3321 & n3401 ) | ( n3321 & ~n3406 ) | ( n3401 & ~n3406 ) ;
  assign n3408 = n1547 ^ n438 ^ n364 ;
  assign n3409 = ~n973 & n3408 ;
  assign n3410 = n3409 ^ n1340 ^ x41 ;
  assign n3411 = ( n1364 & ~n2542 ) | ( n1364 & n2855 ) | ( ~n2542 & n2855 ) ;
  assign n3412 = n3411 ^ n974 ^ n223 ;
  assign n3413 = ( n1489 & n1684 ) | ( n1489 & n3412 ) | ( n1684 & n3412 ) ;
  assign n3414 = ( x125 & n2183 ) | ( x125 & ~n3413 ) | ( n2183 & ~n3413 ) ;
  assign n3415 = n3410 | n3414 ;
  assign n3416 = x64 & ~n2485 ;
  assign n3424 = ( x75 & ~n2498 ) | ( x75 & n3212 ) | ( ~n2498 & n3212 ) ;
  assign n3417 = ~n265 & n2178 ;
  assign n3418 = n3417 ^ x2 ^ 1'b0 ;
  assign n3419 = ( ~n1720 & n1967 ) | ( ~n1720 & n3321 ) | ( n1967 & n3321 ) ;
  assign n3420 = n3419 ^ n2541 ^ n639 ;
  assign n3421 = n1244 & ~n3420 ;
  assign n3422 = n3421 ^ n542 ^ 1'b0 ;
  assign n3423 = ( ~n1210 & n3418 ) | ( ~n1210 & n3422 ) | ( n3418 & n3422 ) ;
  assign n3425 = n3424 ^ n3423 ^ 1'b0 ;
  assign n3426 = n3058 & ~n3425 ;
  assign n3436 = n1011 ^ n847 ^ n181 ;
  assign n3434 = n654 & n1506 ;
  assign n3435 = n3434 ^ n620 ^ 1'b0 ;
  assign n3437 = n3436 ^ n3435 ^ n1539 ;
  assign n3431 = n378 ^ x21 ^ 1'b0 ;
  assign n3432 = ~n472 & n3431 ;
  assign n3427 = n499 ^ n387 ^ 1'b0 ;
  assign n3428 = n168 | n3427 ;
  assign n3429 = n949 ^ n692 ^ n450 ;
  assign n3430 = n3428 | n3429 ;
  assign n3433 = n3432 ^ n3430 ^ 1'b0 ;
  assign n3438 = n3437 ^ n3433 ^ n2376 ;
  assign n3440 = x35 & n1973 ;
  assign n3441 = n3440 ^ n181 ^ 1'b0 ;
  assign n3442 = n3441 ^ n1665 ^ x50 ;
  assign n3443 = n2519 ^ n2144 ^ n253 ;
  assign n3444 = ( n1890 & ~n3442 ) | ( n1890 & n3443 ) | ( ~n3442 & n3443 ) ;
  assign n3439 = n894 ^ n777 ^ n443 ;
  assign n3445 = n3444 ^ n3439 ^ n1909 ;
  assign n3446 = n1848 | n2588 ;
  assign n3447 = n3446 ^ n2788 ^ 1'b0 ;
  assign n3448 = ( n814 & n1558 ) | ( n814 & n3447 ) | ( n1558 & n3447 ) ;
  assign n3449 = n1315 ^ n381 ^ 1'b0 ;
  assign n3450 = n1044 & n3449 ;
  assign n3451 = ( n1125 & n2076 ) | ( n1125 & ~n3450 ) | ( n2076 & ~n3450 ) ;
  assign n3452 = n915 ^ n404 ^ x8 ;
  assign n3453 = ( x92 & n1456 ) | ( x92 & ~n3452 ) | ( n1456 & ~n3452 ) ;
  assign n3454 = n1341 & n2184 ;
  assign n3455 = ~n316 & n3454 ;
  assign n3456 = n3455 ^ n1895 ^ 1'b0 ;
  assign n3457 = n3364 ^ n3061 ^ n777 ;
  assign n3458 = n3457 ^ n1683 ^ n167 ;
  assign n3460 = n956 ^ n456 ^ 1'b0 ;
  assign n3461 = n3441 | n3460 ;
  assign n3459 = n1246 ^ n786 ^ 1'b0 ;
  assign n3462 = n3461 ^ n3459 ^ n1221 ;
  assign n3463 = x9 & ~n1513 ;
  assign n3464 = n3463 ^ n1756 ^ 1'b0 ;
  assign n3465 = ~n1755 & n3057 ;
  assign n3466 = n3465 ^ n2938 ^ 1'b0 ;
  assign n3467 = n3392 ^ n663 ^ 1'b0 ;
  assign n3468 = n1575 & n1654 ;
  assign n3469 = n3119 ^ n1559 ^ 1'b0 ;
  assign n3470 = ( n376 & n3468 ) | ( n376 & n3469 ) | ( n3468 & n3469 ) ;
  assign n3471 = n1051 & n1568 ;
  assign n3472 = n3471 ^ n1137 ^ 1'b0 ;
  assign n3473 = n3447 | n3472 ;
  assign n3474 = n3473 ^ n2106 ^ n1547 ;
  assign n3475 = n645 & n2175 ;
  assign n3476 = n2085 ^ n1498 ^ n447 ;
  assign n3477 = n2976 | n3476 ;
  assign n3478 = n3475 & ~n3477 ;
  assign n3479 = ~n524 & n2601 ;
  assign n3480 = n3479 ^ n2338 ^ 1'b0 ;
  assign n3481 = n2329 ^ n1896 ^ n236 ;
  assign n3482 = ( x16 & n355 ) | ( x16 & n3481 ) | ( n355 & n3481 ) ;
  assign n3483 = ( x79 & ~n697 ) | ( x79 & n1626 ) | ( ~n697 & n1626 ) ;
  assign n3484 = ( ~n129 & n605 ) | ( ~n129 & n1421 ) | ( n605 & n1421 ) ;
  assign n3485 = ( n2870 & n3483 ) | ( n2870 & ~n3484 ) | ( n3483 & ~n3484 ) ;
  assign n3486 = ( n314 & ~n2608 ) | ( n314 & n3485 ) | ( ~n2608 & n3485 ) ;
  assign n3487 = ( ~n1044 & n2700 ) | ( ~n1044 & n3486 ) | ( n2700 & n3486 ) ;
  assign n3488 = ( n1882 & n3482 ) | ( n1882 & ~n3487 ) | ( n3482 & ~n3487 ) ;
  assign n3489 = n620 & n2332 ;
  assign n3490 = n1736 & n3489 ;
  assign n3491 = n729 & n3490 ;
  assign n3492 = n2165 ^ n1182 ^ 1'b0 ;
  assign n3493 = n250 | n3492 ;
  assign n3494 = ~n233 & n2082 ;
  assign n3495 = n3493 & n3494 ;
  assign n3496 = ( n1405 & n2237 ) | ( n1405 & ~n3495 ) | ( n2237 & ~n3495 ) ;
  assign n3497 = n2358 ^ n1489 ^ 1'b0 ;
  assign n3498 = n758 & ~n3497 ;
  assign n3499 = n1525 & ~n3498 ;
  assign n3503 = n253 & ~n1268 ;
  assign n3504 = n3503 ^ n2371 ^ 1'b0 ;
  assign n3505 = n2759 ^ n955 ^ 1'b0 ;
  assign n3506 = ~n3504 & n3505 ;
  assign n3500 = n130 ^ x111 ^ 1'b0 ;
  assign n3501 = n537 & ~n3500 ;
  assign n3502 = n1896 & n3501 ;
  assign n3507 = n3506 ^ n3502 ^ 1'b0 ;
  assign n3508 = n3499 | n3507 ;
  assign n3509 = n3496 | n3508 ;
  assign n3511 = n2519 ^ n1397 ^ x70 ;
  assign n3510 = n3471 ^ n2687 ^ 1'b0 ;
  assign n3512 = n3511 ^ n3510 ^ n1580 ;
  assign n3513 = x20 | n3512 ;
  assign n3514 = n1952 ^ n1757 ^ n709 ;
  assign n3515 = n429 ^ n394 ^ 1'b0 ;
  assign n3516 = ( n1706 & ~n3097 ) | ( n1706 & n3359 ) | ( ~n3097 & n3359 ) ;
  assign n3517 = ( ~x24 & n3515 ) | ( ~x24 & n3516 ) | ( n3515 & n3516 ) ;
  assign n3519 = ( n282 & n2046 ) | ( n282 & ~n3461 ) | ( n2046 & ~n3461 ) ;
  assign n3518 = x87 & ~n3103 ;
  assign n3520 = n3519 ^ n3518 ^ 1'b0 ;
  assign n3521 = n3520 ^ n3401 ^ 1'b0 ;
  assign n3522 = n1964 ^ n1448 ^ n148 ;
  assign n3523 = ~n1578 & n2501 ;
  assign n3524 = n1578 & n3523 ;
  assign n3525 = n3524 ^ n2016 ^ 1'b0 ;
  assign n3526 = ~n3522 & n3525 ;
  assign n3527 = n762 ^ n300 ^ 1'b0 ;
  assign n3528 = n2070 | n3527 ;
  assign n3529 = n3528 ^ n934 ^ 1'b0 ;
  assign n3530 = n1847 ^ n1188 ^ n847 ;
  assign n3531 = n3530 ^ n1486 ^ n1360 ;
  assign n3536 = n2585 ^ n2185 ^ n205 ;
  assign n3537 = n924 | n1380 ;
  assign n3538 = n3536 & ~n3537 ;
  assign n3539 = ~n933 & n3538 ;
  assign n3533 = ( n969 & n1819 ) | ( n969 & n2521 ) | ( n1819 & n2521 ) ;
  assign n3532 = n159 | n268 ;
  assign n3534 = n3533 ^ n3532 ^ 1'b0 ;
  assign n3535 = ~n1976 & n3534 ;
  assign n3540 = n3539 ^ n3535 ^ 1'b0 ;
  assign n3541 = n3540 ^ n890 ^ 1'b0 ;
  assign n3543 = ( n129 & n330 ) | ( n129 & ~n2551 ) | ( n330 & ~n2551 ) ;
  assign n3542 = n179 | n2544 ;
  assign n3544 = n3543 ^ n3542 ^ 1'b0 ;
  assign n3548 = ( n642 & n772 ) | ( n642 & n904 ) | ( n772 & n904 ) ;
  assign n3549 = ( ~n520 & n1111 ) | ( ~n520 & n3548 ) | ( n1111 & n3548 ) ;
  assign n3545 = n1208 ^ n559 ^ n550 ;
  assign n3546 = n1217 | n3545 ;
  assign n3547 = n1280 | n3546 ;
  assign n3550 = n3549 ^ n3547 ^ 1'b0 ;
  assign n3551 = ( ~n1176 & n3544 ) | ( ~n1176 & n3550 ) | ( n3544 & n3550 ) ;
  assign n3552 = ~n259 & n3551 ;
  assign n3553 = ( x119 & n1235 ) | ( x119 & ~n1978 ) | ( n1235 & ~n1978 ) ;
  assign n3554 = n153 | n1227 ;
  assign n3555 = n2314 & ~n3554 ;
  assign n3556 = n3555 ^ n2167 ^ 1'b0 ;
  assign n3557 = x66 ^ x10 ^ 1'b0 ;
  assign n3558 = ~n366 & n3557 ;
  assign n3559 = n1356 ^ n186 ^ 1'b0 ;
  assign n3560 = n3558 & n3559 ;
  assign n3561 = n1852 & ~n3560 ;
  assign n3564 = ~n2596 & n2798 ;
  assign n3562 = ( n332 & n2090 ) | ( n332 & ~n2481 ) | ( n2090 & ~n2481 ) ;
  assign n3563 = n186 | n3562 ;
  assign n3565 = n3564 ^ n3563 ^ 1'b0 ;
  assign n3573 = ( n696 & n1356 ) | ( n696 & n2141 ) | ( n1356 & n2141 ) ;
  assign n3574 = n816 & ~n3573 ;
  assign n3575 = n1533 & n3574 ;
  assign n3566 = n918 ^ n607 ^ 1'b0 ;
  assign n3567 = n2785 | n3566 ;
  assign n3568 = n1650 | n3567 ;
  assign n3569 = n884 & ~n3568 ;
  assign n3570 = n1394 | n3569 ;
  assign n3571 = n3570 ^ n1045 ^ 1'b0 ;
  assign n3572 = n657 | n3571 ;
  assign n3576 = n3575 ^ n3572 ^ 1'b0 ;
  assign n3577 = n629 & ~n1096 ;
  assign n3580 = n1660 & ~n2844 ;
  assign n3581 = n3580 ^ x72 ^ 1'b0 ;
  assign n3578 = n3016 ^ n2570 ^ n835 ;
  assign n3579 = x56 & n3578 ;
  assign n3582 = n3581 ^ n3579 ^ 1'b0 ;
  assign n3583 = n3536 ^ n2343 ^ n1493 ;
  assign n3584 = x29 & ~n3583 ;
  assign n3585 = ~n2564 & n3584 ;
  assign n3599 = n1327 | n2136 ;
  assign n3586 = n1594 ^ n670 ^ 1'b0 ;
  assign n3588 = n2065 ^ x23 ^ 1'b0 ;
  assign n3587 = n3221 ^ n2985 ^ n1811 ;
  assign n3589 = n3588 ^ n3587 ^ n1051 ;
  assign n3590 = ~n897 & n2429 ;
  assign n3591 = ~n1847 & n3590 ;
  assign n3592 = n3591 ^ n2914 ^ n1718 ;
  assign n3593 = n3592 ^ n1452 ^ x75 ;
  assign n3594 = n2545 | n3593 ;
  assign n3595 = n2509 | n3594 ;
  assign n3596 = ( n2349 & n3589 ) | ( n2349 & n3595 ) | ( n3589 & n3595 ) ;
  assign n3597 = ( ~n1186 & n3586 ) | ( ~n1186 & n3596 ) | ( n3586 & n3596 ) ;
  assign n3598 = n3597 ^ n1390 ^ n524 ;
  assign n3600 = n3599 ^ n3598 ^ n1099 ;
  assign n3601 = ~n748 & n1154 ;
  assign n3602 = n1007 & n3601 ;
  assign n3604 = n1335 ^ n580 ^ n184 ;
  assign n3605 = ( n1316 & n1747 ) | ( n1316 & ~n3604 ) | ( n1747 & ~n3604 ) ;
  assign n3603 = n1762 | n3436 ;
  assign n3606 = n3605 ^ n3603 ^ 1'b0 ;
  assign n3607 = n3602 | n3606 ;
  assign n3608 = ( x28 & ~n740 ) | ( x28 & n1160 ) | ( ~n740 & n1160 ) ;
  assign n3609 = ~x79 & n3608 ;
  assign n3610 = n1470 & n3609 ;
  assign n3611 = n3269 & ~n3610 ;
  assign n3612 = n3611 ^ n1911 ^ 1'b0 ;
  assign n3613 = n416 & n2628 ;
  assign n3614 = n3613 ^ n206 ^ 1'b0 ;
  assign n3615 = ( x92 & ~n1164 ) | ( x92 & n3614 ) | ( ~n1164 & n3614 ) ;
  assign n3616 = n1050 & n3615 ;
  assign n3617 = n2788 & n3616 ;
  assign n3618 = x1 & ~n1896 ;
  assign n3619 = n2315 & n3618 ;
  assign n3620 = ( x5 & ~n915 ) | ( x5 & n2427 ) | ( ~n915 & n2427 ) ;
  assign n3621 = n1820 & n3620 ;
  assign n3622 = ~n3097 & n3621 ;
  assign n3623 = n130 & n1188 ;
  assign n3624 = n1282 & n3623 ;
  assign n3625 = n3624 ^ n1437 ^ 1'b0 ;
  assign n3626 = n1184 ^ n847 ^ 1'b0 ;
  assign n3627 = n330 & n3626 ;
  assign n3628 = ( n2488 & n2974 ) | ( n2488 & ~n3627 ) | ( n2974 & ~n3627 ) ;
  assign n3629 = ( n2062 & n2724 ) | ( n2062 & ~n3628 ) | ( n2724 & ~n3628 ) ;
  assign n3630 = n3629 ^ n412 ^ 1'b0 ;
  assign n3631 = n911 | n3630 ;
  assign n3632 = n2815 ^ n1436 ^ n839 ;
  assign n3633 = x4 & ~n2176 ;
  assign n3634 = ( n1220 & n3048 ) | ( n1220 & ~n3633 ) | ( n3048 & ~n3633 ) ;
  assign n3635 = n2130 ^ n1690 ^ 1'b0 ;
  assign n3640 = ~n756 & n887 ;
  assign n3636 = n3280 ^ n834 ^ n414 ;
  assign n3637 = n3636 ^ n2344 ^ 1'b0 ;
  assign n3638 = x66 & n3637 ;
  assign n3639 = n3638 ^ n3062 ^ n183 ;
  assign n3641 = n3640 ^ n3639 ^ n2257 ;
  assign n3642 = n3641 ^ n3359 ^ 1'b0 ;
  assign n3643 = n1977 & ~n3642 ;
  assign n3644 = n978 & n3643 ;
  assign n3645 = n3341 ^ n1012 ^ 1'b0 ;
  assign n3646 = n3645 ^ n3610 ^ n660 ;
  assign n3647 = n1290 ^ n1255 ^ n1065 ;
  assign n3648 = n3647 ^ n394 ^ x6 ;
  assign n3649 = n3646 & n3648 ;
  assign n3650 = n133 & ~n3649 ;
  assign n3657 = n512 & n3183 ;
  assign n3651 = n1071 ^ n1016 ^ n1011 ;
  assign n3652 = ( ~x75 & n2670 ) | ( ~x75 & n3651 ) | ( n2670 & n3651 ) ;
  assign n3653 = ( ~n481 & n1210 ) | ( ~n481 & n1431 ) | ( n1210 & n1431 ) ;
  assign n3654 = n3653 ^ n2657 ^ 1'b0 ;
  assign n3655 = n3522 | n3654 ;
  assign n3656 = n3652 & ~n3655 ;
  assign n3658 = n3657 ^ n3656 ^ 1'b0 ;
  assign n3659 = n1918 & n3658 ;
  assign n3660 = n1485 | n2914 ;
  assign n3661 = n3660 ^ n1828 ^ 1'b0 ;
  assign n3662 = n3661 ^ n1899 ^ 1'b0 ;
  assign n3663 = n2478 ^ x38 ^ 1'b0 ;
  assign n3664 = n1235 & ~n3663 ;
  assign n3665 = n1459 ^ n214 ^ 1'b0 ;
  assign n3666 = n3665 ^ n2776 ^ n698 ;
  assign n3667 = n2576 ^ n2436 ^ 1'b0 ;
  assign n3668 = n3667 ^ n526 ^ n503 ;
  assign n3669 = n714 & n3668 ;
  assign n3670 = n3669 ^ n2109 ^ 1'b0 ;
  assign n3671 = n2539 ^ n1952 ^ 1'b0 ;
  assign n3672 = n3671 ^ n652 ^ 1'b0 ;
  assign n3673 = n3672 ^ n3173 ^ n3037 ;
  assign n3674 = n2379 ^ n310 ^ 1'b0 ;
  assign n3685 = n1551 & ~n1738 ;
  assign n3686 = ~x34 & n3685 ;
  assign n3687 = ( x38 & n547 ) | ( x38 & n2428 ) | ( n547 & n2428 ) ;
  assign n3688 = ( n1136 & ~n2797 ) | ( n1136 & n3687 ) | ( ~n2797 & n3687 ) ;
  assign n3689 = n3688 ^ n2256 ^ n1886 ;
  assign n3690 = ( n2590 & n3686 ) | ( n2590 & ~n3689 ) | ( n3686 & ~n3689 ) ;
  assign n3691 = n3690 ^ n2682 ^ x89 ;
  assign n3678 = n2227 ^ n1548 ^ n134 ;
  assign n3677 = ( n1160 & n1422 ) | ( n1160 & ~n2405 ) | ( n1422 & ~n2405 ) ;
  assign n3679 = n3678 ^ n3677 ^ n1360 ;
  assign n3675 = n2256 ^ n1957 ^ n1422 ;
  assign n3676 = ( n1725 & n1831 ) | ( n1725 & ~n3675 ) | ( n1831 & ~n3675 ) ;
  assign n3680 = n3679 ^ n3676 ^ 1'b0 ;
  assign n3681 = n2405 ^ n2360 ^ n332 ;
  assign n3682 = ~n3063 & n3681 ;
  assign n3683 = n2474 & n3682 ;
  assign n3684 = ( n1239 & ~n3680 ) | ( n1239 & n3683 ) | ( ~n3680 & n3683 ) ;
  assign n3692 = n3691 ^ n3684 ^ 1'b0 ;
  assign n3693 = ~n3674 & n3692 ;
  assign n3696 = n3012 ^ n520 ^ 1'b0 ;
  assign n3697 = ( ~x123 & n319 ) | ( ~x123 & n3696 ) | ( n319 & n3696 ) ;
  assign n3694 = ~n999 & n2175 ;
  assign n3695 = n3694 ^ n1684 ^ 1'b0 ;
  assign n3698 = n3697 ^ n3695 ^ n1450 ;
  assign n3699 = n3379 & n3698 ;
  assign n3700 = n2471 ^ n1427 ^ n1315 ;
  assign n3701 = n2055 ^ n1755 ^ 1'b0 ;
  assign n3702 = n1176 ^ n356 ^ n246 ;
  assign n3703 = n3702 ^ x40 ^ 1'b0 ;
  assign n3704 = ( n2324 & n3701 ) | ( n2324 & n3703 ) | ( n3701 & n3703 ) ;
  assign n3705 = ( n369 & n1412 ) | ( n369 & ~n3498 ) | ( n1412 & ~n3498 ) ;
  assign n3706 = n2257 & n3705 ;
  assign n3707 = n3706 ^ n2822 ^ n1636 ;
  assign n3708 = n562 | n3437 ;
  assign n3709 = n3708 ^ n2972 ^ 1'b0 ;
  assign n3710 = ( n2090 & n2812 ) | ( n2090 & n3709 ) | ( n2812 & n3709 ) ;
  assign n3711 = ( n294 & n370 ) | ( n294 & n3710 ) | ( n370 & n3710 ) ;
  assign n3712 = n2486 ^ n1804 ^ n1683 ;
  assign n3713 = ( ~n205 & n3711 ) | ( ~n205 & n3712 ) | ( n3711 & n3712 ) ;
  assign n3714 = n3713 ^ n2076 ^ 1'b0 ;
  assign n3715 = n3707 | n3714 ;
  assign n3721 = n3452 ^ n1962 ^ n1019 ;
  assign n3717 = n1656 ^ n186 ^ 1'b0 ;
  assign n3718 = n2763 & n3717 ;
  assign n3719 = ( ~n1914 & n2344 ) | ( ~n1914 & n3718 ) | ( n2344 & n3718 ) ;
  assign n3720 = n3719 ^ x10 ^ 1'b0 ;
  assign n3716 = n1831 ^ n148 ^ 1'b0 ;
  assign n3722 = n3721 ^ n3720 ^ n3716 ;
  assign n3723 = n2718 ^ n951 ^ x50 ;
  assign n3724 = ( n150 & ~n2193 ) | ( n150 & n3723 ) | ( ~n2193 & n3723 ) ;
  assign n3725 = n3724 ^ n1808 ^ 1'b0 ;
  assign n3726 = ~n1947 & n3725 ;
  assign n3727 = n414 ^ n322 ^ 1'b0 ;
  assign n3728 = n2880 ^ n1030 ^ n849 ;
  assign n3729 = n3728 ^ n3336 ^ n1672 ;
  assign n3730 = ( n544 & ~n2579 ) | ( n544 & n3729 ) | ( ~n2579 & n3729 ) ;
  assign n3731 = n1296 ^ n1155 ^ 1'b0 ;
  assign n3732 = n1459 & ~n3731 ;
  assign n3733 = n3730 & ~n3732 ;
  assign n3734 = ( n1344 & n1894 ) | ( n1344 & n3195 ) | ( n1894 & n3195 ) ;
  assign n3735 = n1885 ^ n1318 ^ n332 ;
  assign n3736 = ( ~n611 & n3614 ) | ( ~n611 & n3735 ) | ( n3614 & n3735 ) ;
  assign n3737 = n1036 ^ n351 ^ 1'b0 ;
  assign n3738 = n2884 & ~n3737 ;
  assign n3739 = ( n375 & n2498 ) | ( n375 & n3738 ) | ( n2498 & n3738 ) ;
  assign n3741 = n219 & ~n772 ;
  assign n3740 = n2844 ^ n2696 ^ n619 ;
  assign n3742 = n3741 ^ n3740 ^ 1'b0 ;
  assign n3743 = ( x59 & x115 ) | ( x59 & ~n2178 ) | ( x115 & ~n2178 ) ;
  assign n3744 = n1497 ^ n656 ^ 1'b0 ;
  assign n3745 = n3744 ^ n3402 ^ n157 ;
  assign n3748 = ( n176 & n1838 ) | ( n176 & ~n2013 ) | ( n1838 & ~n2013 ) ;
  assign n3749 = ( ~x41 & n794 ) | ( ~x41 & n3748 ) | ( n794 & n3748 ) ;
  assign n3746 = n2772 ^ n1523 ^ 1'b0 ;
  assign n3747 = n3364 & n3746 ;
  assign n3750 = n3749 ^ n3747 ^ 1'b0 ;
  assign n3751 = n3750 ^ n1981 ^ 1'b0 ;
  assign n3752 = n549 & ~n3751 ;
  assign n3755 = n1391 ^ n598 ^ x67 ;
  assign n3756 = ( n469 & n2629 ) | ( n469 & n3755 ) | ( n2629 & n3755 ) ;
  assign n3753 = n1486 | n1933 ;
  assign n3754 = n3753 ^ n588 ^ 1'b0 ;
  assign n3757 = n3756 ^ n3754 ^ n1107 ;
  assign n3758 = n3247 ^ n3113 ^ n758 ;
  assign n3759 = ( n1622 & n1671 ) | ( n1622 & n3758 ) | ( n1671 & n3758 ) ;
  assign n3760 = n3759 ^ n3301 ^ 1'b0 ;
  assign n3761 = ( n472 & n770 ) | ( n472 & ~n796 ) | ( n770 & ~n796 ) ;
  assign n3762 = n2083 & n3761 ;
  assign n3763 = n3083 ^ n364 ^ 1'b0 ;
  assign n3764 = ( n839 & n3762 ) | ( n839 & ~n3763 ) | ( n3762 & ~n3763 ) ;
  assign n3765 = n2840 ^ n2224 ^ 1'b0 ;
  assign n3766 = n2288 & n3765 ;
  assign n3767 = ~n2335 & n2479 ;
  assign n3768 = ~n3766 & n3767 ;
  assign n3769 = ( n1912 & n3136 ) | ( n1912 & ~n3163 ) | ( n3136 & ~n3163 ) ;
  assign n3770 = n1269 ^ n445 ^ n244 ;
  assign n3771 = n3770 ^ n3689 ^ n1761 ;
  assign n3772 = n244 ^ n213 ^ 1'b0 ;
  assign n3773 = n2209 & n3772 ;
  assign n3774 = n3041 ^ n2121 ^ n1876 ;
  assign n3775 = n3774 ^ n3671 ^ 1'b0 ;
  assign n3776 = n2269 ^ n201 ^ 1'b0 ;
  assign n3777 = n3776 ^ n580 ^ 1'b0 ;
  assign n3778 = n310 & ~n3777 ;
  assign n3779 = ~n2559 & n3550 ;
  assign n3780 = n3779 ^ n3369 ^ 1'b0 ;
  assign n3781 = ( n1771 & ~n3778 ) | ( n1771 & n3780 ) | ( ~n3778 & n3780 ) ;
  assign n3782 = n2987 ^ n424 ^ 1'b0 ;
  assign n3783 = ~n3781 & n3782 ;
  assign n3784 = ( n415 & n1036 ) | ( n415 & n1269 ) | ( n1036 & n1269 ) ;
  assign n3785 = n3784 ^ n1987 ^ 1'b0 ;
  assign n3786 = n3785 ^ n1052 ^ 1'b0 ;
  assign n3787 = x42 & n3786 ;
  assign n3788 = n663 & n1714 ;
  assign n3789 = ~n3194 & n3788 ;
  assign n3790 = x70 & n2526 ;
  assign n3791 = n3790 ^ n706 ^ 1'b0 ;
  assign n3792 = n2301 ^ n626 ^ 1'b0 ;
  assign n3793 = n2972 | n3792 ;
  assign n3794 = n3791 & ~n3793 ;
  assign n3795 = ( n1008 & n1952 ) | ( n1008 & n3794 ) | ( n1952 & n3794 ) ;
  assign n3796 = n3009 ^ n2771 ^ n1346 ;
  assign n3798 = n155 ^ x84 ^ x58 ;
  assign n3799 = n3798 ^ n1136 ^ x2 ;
  assign n3797 = n3088 ^ n829 ^ x103 ;
  assign n3800 = n3799 ^ n3797 ^ n783 ;
  assign n3801 = n2216 | n3800 ;
  assign n3802 = n1097 | n3801 ;
  assign n3803 = n3149 ^ n790 ^ 1'b0 ;
  assign n3804 = n3802 & ~n3803 ;
  assign n3805 = n3622 ^ n2692 ^ n691 ;
  assign n3806 = n454 & ~n3409 ;
  assign n3809 = n1656 ^ n1391 ^ 1'b0 ;
  assign n3808 = n3260 ^ n1804 ^ n765 ;
  assign n3807 = n2883 ^ n1441 ^ x43 ;
  assign n3810 = n3809 ^ n3808 ^ n3807 ;
  assign n3811 = ( n1688 & n3806 ) | ( n1688 & ~n3810 ) | ( n3806 & ~n3810 ) ;
  assign n3812 = n538 ^ n266 ^ 1'b0 ;
  assign n3813 = ( n1152 & n1243 ) | ( n1152 & ~n3812 ) | ( n1243 & ~n3812 ) ;
  assign n3814 = n3813 ^ n2446 ^ n2264 ;
  assign n3815 = n3814 ^ n2237 ^ n888 ;
  assign n3816 = n2631 ^ x97 ^ x70 ;
  assign n3827 = n218 | n3187 ;
  assign n3826 = ( n584 & n1232 ) | ( n584 & n1919 ) | ( n1232 & n1919 ) ;
  assign n3828 = n3827 ^ n3826 ^ n1209 ;
  assign n3829 = n3828 ^ n1567 ^ x17 ;
  assign n3817 = x43 & n2833 ;
  assign n3818 = ( n324 & ~n2657 ) | ( n324 & n3817 ) | ( ~n2657 & n3817 ) ;
  assign n3819 = n2884 ^ n2713 ^ n2247 ;
  assign n3820 = n1978 ^ n533 ^ 1'b0 ;
  assign n3821 = n980 ^ x97 ^ 1'b0 ;
  assign n3822 = n3820 & ~n3821 ;
  assign n3823 = n3819 & n3822 ;
  assign n3824 = n3818 & ~n3823 ;
  assign n3825 = ~n2458 & n3824 ;
  assign n3830 = n3829 ^ n3825 ^ n483 ;
  assign n3831 = n3358 ^ n2778 ^ 1'b0 ;
  assign n3832 = n3831 ^ n2622 ^ n1737 ;
  assign n3833 = n2671 ^ n1294 ^ 1'b0 ;
  assign n3834 = ~n1894 & n3833 ;
  assign n3837 = x46 & n923 ;
  assign n3835 = n2203 ^ n1849 ^ n1117 ;
  assign n3836 = ( n2210 & ~n3207 ) | ( n2210 & n3835 ) | ( ~n3207 & n3835 ) ;
  assign n3838 = n3837 ^ n3836 ^ n1711 ;
  assign n3839 = n3838 ^ n1460 ^ n1084 ;
  assign n3840 = n3839 ^ n2993 ^ n1342 ;
  assign n3841 = n3382 ^ n3071 ^ n2443 ;
  assign n3842 = n2615 & n3841 ;
  assign n3843 = n3842 ^ n1999 ^ 1'b0 ;
  assign n3844 = n3240 ^ n662 ^ 1'b0 ;
  assign n3845 = n2210 & ~n3844 ;
  assign n3846 = n3845 ^ n850 ^ x29 ;
  assign n3847 = ( n748 & n2612 ) | ( n748 & n3846 ) | ( n2612 & n3846 ) ;
  assign n3848 = n2091 ^ x13 ^ 1'b0 ;
  assign n3849 = n1846 & ~n2046 ;
  assign n3850 = n3849 ^ n3379 ^ 1'b0 ;
  assign n3851 = n2599 & n3850 ;
  assign n3852 = ( n345 & n3406 ) | ( n345 & ~n3851 ) | ( n3406 & ~n3851 ) ;
  assign n3853 = ( n409 & ~n2249 ) | ( n409 & n2978 ) | ( ~n2249 & n2978 ) ;
  assign n3854 = x116 & ~n1740 ;
  assign n3855 = n2697 | n2863 ;
  assign n3856 = n3854 & ~n3855 ;
  assign n3857 = n3856 ^ n748 ^ 1'b0 ;
  assign n3858 = n879 & n3857 ;
  assign n3859 = n900 & ~n2697 ;
  assign n3860 = n3859 ^ n1343 ^ 1'b0 ;
  assign n3861 = n1685 & ~n3860 ;
  assign n3862 = ~n741 & n3861 ;
  assign n3863 = n764 | n3862 ;
  assign n3864 = n410 & ~n3863 ;
  assign n3871 = ( n998 & n3274 ) | ( n998 & ~n3385 ) | ( n3274 & ~n3385 ) ;
  assign n3868 = ~n2867 & n3050 ;
  assign n3865 = n1366 | n1555 ;
  assign n3866 = n3865 ^ n2347 ^ 1'b0 ;
  assign n3867 = ~n328 & n3866 ;
  assign n3869 = n3868 ^ n3867 ^ 1'b0 ;
  assign n3870 = n2970 & n3869 ;
  assign n3872 = n3871 ^ n3870 ^ 1'b0 ;
  assign n3873 = x96 & n2030 ;
  assign n3874 = ~x118 & n3873 ;
  assign n3875 = n1942 & ~n3874 ;
  assign n3876 = ( ~n1055 & n1828 ) | ( ~n1055 & n2307 ) | ( n1828 & n2307 ) ;
  assign n3877 = n1639 & n2893 ;
  assign n3878 = ~n3876 & n3877 ;
  assign n3879 = n3878 ^ n1645 ^ 1'b0 ;
  assign n3880 = ( n437 & n3875 ) | ( n437 & n3879 ) | ( n3875 & n3879 ) ;
  assign n3881 = n447 ^ n143 ^ 1'b0 ;
  assign n3882 = ( x6 & n3837 ) | ( x6 & n3881 ) | ( n3837 & n3881 ) ;
  assign n3883 = ( ~x56 & n2781 ) | ( ~x56 & n3882 ) | ( n2781 & n3882 ) ;
  assign n3884 = n1091 | n3883 ;
  assign n3885 = n476 & ~n3884 ;
  assign n3886 = n3468 ^ n3414 ^ n2633 ;
  assign n3887 = ( n2512 & ~n3885 ) | ( n2512 & n3886 ) | ( ~n3885 & n3886 ) ;
  assign n3888 = ( x4 & n1239 ) | ( x4 & ~n1358 ) | ( n1239 & ~n1358 ) ;
  assign n3889 = ( n1066 & ~n1316 ) | ( n1066 & n2132 ) | ( ~n1316 & n2132 ) ;
  assign n3890 = n408 | n1253 ;
  assign n3891 = x63 | n3890 ;
  assign n3892 = ( n2378 & n2464 ) | ( n2378 & ~n3891 ) | ( n2464 & ~n3891 ) ;
  assign n3893 = n3892 ^ n3544 ^ 1'b0 ;
  assign n3894 = n3889 | n3893 ;
  assign n3895 = n710 | n3894 ;
  assign n3896 = n1246 ^ n1085 ^ 1'b0 ;
  assign n3897 = n1113 ^ n762 ^ n434 ;
  assign n3898 = ( ~x68 & n2827 ) | ( ~x68 & n3897 ) | ( n2827 & n3897 ) ;
  assign n3899 = n3898 ^ x2 ^ 1'b0 ;
  assign n3900 = ( ~n901 & n2277 ) | ( ~n901 & n3169 ) | ( n2277 & n3169 ) ;
  assign n3901 = ( ~n1524 & n3341 ) | ( ~n1524 & n3900 ) | ( n3341 & n3900 ) ;
  assign n3902 = ( x112 & ~n1204 ) | ( x112 & n3901 ) | ( ~n1204 & n3901 ) ;
  assign n3913 = n1468 ^ n360 ^ 1'b0 ;
  assign n3903 = n792 & ~n1012 ;
  assign n3904 = n1518 ^ n1276 ^ 1'b0 ;
  assign n3907 = n697 & ~n801 ;
  assign n3908 = n206 & n3907 ;
  assign n3909 = ~n3282 & n3908 ;
  assign n3905 = n1717 ^ n653 ^ 1'b0 ;
  assign n3906 = n2012 & ~n3905 ;
  assign n3910 = n3909 ^ n3906 ^ 1'b0 ;
  assign n3911 = n3904 & n3910 ;
  assign n3912 = ~n3903 & n3911 ;
  assign n3914 = n3913 ^ n3912 ^ n302 ;
  assign n3916 = n2564 ^ n2269 ^ n2020 ;
  assign n3915 = ( n849 & n1296 ) | ( n849 & n1411 ) | ( n1296 & n1411 ) ;
  assign n3917 = n3916 ^ n3915 ^ n1534 ;
  assign n3918 = n602 & ~n892 ;
  assign n3919 = n2642 ^ x115 ^ 1'b0 ;
  assign n3920 = n2840 ^ n1090 ^ n420 ;
  assign n3921 = ( n3918 & n3919 ) | ( n3918 & ~n3920 ) | ( n3919 & ~n3920 ) ;
  assign n3925 = ( n777 & n794 ) | ( n777 & n1316 ) | ( n794 & n1316 ) ;
  assign n3922 = ( n493 & n678 ) | ( n493 & n2171 ) | ( n678 & n2171 ) ;
  assign n3923 = ~n1622 & n3922 ;
  assign n3924 = ~n2343 & n3923 ;
  assign n3926 = n3925 ^ n3924 ^ 1'b0 ;
  assign n3927 = n2847 ^ n2616 ^ n1158 ;
  assign n3928 = n2356 ^ n1361 ^ x2 ;
  assign n3929 = n3928 ^ n3544 ^ n174 ;
  assign n3930 = n3929 ^ n402 ^ 1'b0 ;
  assign n3931 = n1668 ^ n1500 ^ 1'b0 ;
  assign n3932 = n1796 & ~n3931 ;
  assign n3942 = n2159 ^ n2053 ^ 1'b0 ;
  assign n3940 = n3163 ^ n1769 ^ n531 ;
  assign n3933 = ~n426 & n656 ;
  assign n3934 = n3933 ^ n230 ^ 1'b0 ;
  assign n3935 = n3934 ^ n209 ^ 1'b0 ;
  assign n3937 = ~n1436 & n1911 ;
  assign n3936 = n1648 ^ n1429 ^ n874 ;
  assign n3938 = n3937 ^ n3936 ^ x5 ;
  assign n3939 = n3935 | n3938 ;
  assign n3941 = n3940 ^ n3939 ^ 1'b0 ;
  assign n3943 = n3942 ^ n3941 ^ n1722 ;
  assign n3944 = ( ~n480 & n3932 ) | ( ~n480 & n3943 ) | ( n3932 & n3943 ) ;
  assign n3945 = n256 | n1509 ;
  assign n3946 = n3945 ^ n145 ^ 1'b0 ;
  assign n3947 = n3944 & n3946 ;
  assign n3948 = ( n1914 & n2539 ) | ( n1914 & ~n3668 ) | ( n2539 & ~n3668 ) ;
  assign n3949 = n3834 & n3948 ;
  assign n3950 = n3949 ^ n2150 ^ 1'b0 ;
  assign n3952 = n1017 ^ n287 ^ 1'b0 ;
  assign n3953 = x83 & n3952 ;
  assign n3954 = n1188 & n3953 ;
  assign n3955 = ~n3146 & n3954 ;
  assign n3956 = ( n2365 & ~n3648 ) | ( n2365 & n3955 ) | ( ~n3648 & n3955 ) ;
  assign n3957 = n3956 ^ n2160 ^ 1'b0 ;
  assign n3958 = n3957 ^ n2513 ^ 1'b0 ;
  assign n3951 = n2663 & n3187 ;
  assign n3959 = n3958 ^ n3951 ^ 1'b0 ;
  assign n3963 = n2118 ^ n375 ^ x52 ;
  assign n3962 = n1646 ^ n199 ^ 1'b0 ;
  assign n3964 = n3963 ^ n3962 ^ 1'b0 ;
  assign n3960 = n3179 | n3255 ;
  assign n3961 = n3761 & ~n3960 ;
  assign n3965 = n3964 ^ n3961 ^ n1214 ;
  assign n3966 = ( ~n575 & n836 ) | ( ~n575 & n1100 ) | ( n836 & n1100 ) ;
  assign n3968 = ~n364 & n1373 ;
  assign n3969 = n903 & n3968 ;
  assign n3970 = n849 | n3969 ;
  assign n3971 = n3970 ^ n3461 ^ 1'b0 ;
  assign n3967 = n1025 ^ n497 ^ 1'b0 ;
  assign n3972 = n3971 ^ n3967 ^ 1'b0 ;
  assign n3973 = n754 & ~n3972 ;
  assign n3974 = ~n1468 & n3973 ;
  assign n3975 = n3521 & n3974 ;
  assign n3976 = n293 & ~n3936 ;
  assign n3977 = ~n1358 & n3976 ;
  assign n3978 = ( ~n561 & n2907 ) | ( ~n561 & n3977 ) | ( n2907 & n3977 ) ;
  assign n3979 = n3978 ^ n2955 ^ 1'b0 ;
  assign n3980 = n145 | n3282 ;
  assign n3981 = n3776 & ~n3980 ;
  assign n3982 = n814 & ~n1677 ;
  assign n3983 = n3982 ^ n2532 ^ 1'b0 ;
  assign n3984 = n374 & n3983 ;
  assign n3985 = n2587 ^ n2236 ^ n527 ;
  assign n3986 = n457 & ~n3985 ;
  assign n3987 = n2467 & n3986 ;
  assign n3988 = n3987 ^ n3759 ^ n2709 ;
  assign n3989 = n1873 ^ n690 ^ n562 ;
  assign n3990 = n1741 ^ n720 ^ 1'b0 ;
  assign n3991 = ( ~x36 & n3738 ) | ( ~x36 & n3990 ) | ( n3738 & n3990 ) ;
  assign n3992 = n1747 & n3991 ;
  assign n3993 = n309 & n2722 ;
  assign n3994 = ~n3198 & n3993 ;
  assign n3995 = n3994 ^ n1953 ^ 1'b0 ;
  assign n3996 = n2629 | n3704 ;
  assign n4003 = ( ~n158 & n714 ) | ( ~n158 & n1419 ) | ( n714 & n1419 ) ;
  assign n3997 = x97 & n1443 ;
  assign n3998 = ~x31 & n3997 ;
  assign n3999 = n2032 ^ n915 ^ 1'b0 ;
  assign n4000 = n3998 | n3999 ;
  assign n4001 = n2905 | n4000 ;
  assign n4002 = n1366 & ~n4001 ;
  assign n4004 = n4003 ^ n4002 ^ n2967 ;
  assign n4009 = n200 & n1427 ;
  assign n4010 = n4009 ^ n3319 ^ 1'b0 ;
  assign n4005 = n2826 ^ n2808 ^ n1018 ;
  assign n4006 = ( n1761 & n2624 ) | ( n1761 & ~n4005 ) | ( n2624 & ~n4005 ) ;
  assign n4007 = x105 & n4006 ;
  assign n4008 = n4007 ^ n481 ^ 1'b0 ;
  assign n4011 = n4010 ^ n4008 ^ n606 ;
  assign n4012 = ( n217 & ~n1756 ) | ( n217 & n3242 ) | ( ~n1756 & n3242 ) ;
  assign n4013 = ~n686 & n1476 ;
  assign n4014 = n4013 ^ n1335 ^ 1'b0 ;
  assign n4015 = n4011 ^ n3320 ^ 1'b0 ;
  assign n4016 = x87 & ~n309 ;
  assign n4019 = ( n1360 & n1479 ) | ( n1360 & n3341 ) | ( n1479 & n3341 ) ;
  assign n4017 = n1219 ^ n950 ^ n171 ;
  assign n4018 = ( n1695 & n2174 ) | ( n1695 & n4017 ) | ( n2174 & n4017 ) ;
  assign n4020 = n4019 ^ n4018 ^ n708 ;
  assign n4021 = n4020 ^ n270 ^ 1'b0 ;
  assign n4022 = ~n4016 & n4021 ;
  assign n4024 = n1553 ^ x115 ^ 1'b0 ;
  assign n4023 = n2004 ^ x110 ^ 1'b0 ;
  assign n4025 = n4024 ^ n4023 ^ 1'b0 ;
  assign n4026 = n2876 & n4025 ;
  assign n4027 = ~n248 & n4026 ;
  assign n4028 = ~n4022 & n4027 ;
  assign n4029 = n2141 ^ n925 ^ n459 ;
  assign n4030 = ( n380 & n1050 ) | ( n380 & n1558 ) | ( n1050 & n1558 ) ;
  assign n4031 = n4030 ^ n3007 ^ n725 ;
  assign n4032 = n3940 ^ n1411 ^ 1'b0 ;
  assign n4033 = n1620 & ~n4032 ;
  assign n4034 = n2827 ^ n736 ^ 1'b0 ;
  assign n4035 = ( n664 & n4033 ) | ( n664 & ~n4034 ) | ( n4033 & ~n4034 ) ;
  assign n4036 = ~n2379 & n3147 ;
  assign n4037 = ( n800 & n1139 ) | ( n800 & ~n4036 ) | ( n1139 & ~n4036 ) ;
  assign n4038 = n410 & n1026 ;
  assign n4039 = n4038 ^ n1237 ^ 1'b0 ;
  assign n4040 = ( n353 & ~n844 ) | ( n353 & n2585 ) | ( ~n844 & n2585 ) ;
  assign n4041 = ( n4037 & n4039 ) | ( n4037 & n4040 ) | ( n4039 & n4040 ) ;
  assign n4042 = n2599 | n4041 ;
  assign n4043 = n4042 ^ n1448 ^ 1'b0 ;
  assign n4044 = n1266 | n4043 ;
  assign n4045 = n1847 | n4044 ;
  assign n4046 = n2811 | n3096 ;
  assign n4047 = n4045 | n4046 ;
  assign n4049 = n2181 & n2489 ;
  assign n4048 = n3339 ^ n2056 ^ 1'b0 ;
  assign n4050 = n4049 ^ n4048 ^ n1891 ;
  assign n4051 = n4050 ^ n1266 ^ 1'b0 ;
  assign n4052 = ( ~n1633 & n1984 ) | ( ~n1633 & n3757 ) | ( n1984 & n3757 ) ;
  assign n4054 = n1100 & ~n1874 ;
  assign n4055 = ~x37 & n4054 ;
  assign n4053 = n1197 & ~n2151 ;
  assign n4056 = n4055 ^ n4053 ^ 1'b0 ;
  assign n4057 = n414 & ~n3586 ;
  assign n4058 = ~n1112 & n2685 ;
  assign n4059 = n4058 ^ n2629 ^ 1'b0 ;
  assign n4060 = ( n1147 & n2812 ) | ( n1147 & ~n3287 ) | ( n2812 & ~n3287 ) ;
  assign n4061 = ( n1970 & ~n4059 ) | ( n1970 & n4060 ) | ( ~n4059 & n4060 ) ;
  assign n4062 = n2720 ^ n527 ^ 1'b0 ;
  assign n4063 = ( n3551 & n4061 ) | ( n3551 & ~n4062 ) | ( n4061 & ~n4062 ) ;
  assign n4064 = n2020 ^ n1145 ^ 1'b0 ;
  assign n4065 = n3175 & n4064 ;
  assign n4066 = ( n1050 & n3344 ) | ( n1050 & ~n4065 ) | ( n3344 & ~n4065 ) ;
  assign n4067 = n1164 | n2256 ;
  assign n4068 = n2801 ^ n1351 ^ n540 ;
  assign n4069 = ( ~n1300 & n2571 ) | ( ~n1300 & n3238 ) | ( n2571 & n3238 ) ;
  assign n4073 = ( n350 & n454 ) | ( n350 & ~n555 ) | ( n454 & ~n555 ) ;
  assign n4074 = ( x93 & n736 ) | ( x93 & ~n2539 ) | ( n736 & ~n2539 ) ;
  assign n4075 = ( n883 & n4073 ) | ( n883 & ~n4074 ) | ( n4073 & ~n4074 ) ;
  assign n4070 = n1919 ^ n746 ^ n616 ;
  assign n4071 = ~n1090 & n4070 ;
  assign n4072 = n4071 ^ n3220 ^ 1'b0 ;
  assign n4076 = n4075 ^ n4072 ^ n1426 ;
  assign n4077 = n4076 ^ n3024 ^ x39 ;
  assign n4078 = ~n510 & n2279 ;
  assign n4079 = n4078 ^ n2242 ^ 1'b0 ;
  assign n4080 = n3969 ^ n3212 ^ 1'b0 ;
  assign n4081 = ( ~n3035 & n3273 ) | ( ~n3035 & n4080 ) | ( n3273 & n4080 ) ;
  assign n4082 = n4081 ^ n3898 ^ 1'b0 ;
  assign n4083 = n964 | n4082 ;
  assign n4084 = ( ~x0 & n2679 ) | ( ~x0 & n3510 ) | ( n2679 & n3510 ) ;
  assign n4085 = ~n878 & n2112 ;
  assign n4086 = n1755 & n4085 ;
  assign n4087 = ( n240 & ~n652 ) | ( n240 & n1394 ) | ( ~n652 & n1394 ) ;
  assign n4088 = ( x89 & n3109 ) | ( x89 & ~n4087 ) | ( n3109 & ~n4087 ) ;
  assign n4089 = ( n1106 & n4086 ) | ( n1106 & n4088 ) | ( n4086 & n4088 ) ;
  assign n4090 = n1118 & ~n1709 ;
  assign n4093 = n2622 ^ n1272 ^ 1'b0 ;
  assign n4091 = ~n907 & n3153 ;
  assign n4092 = n4091 ^ n3448 ^ 1'b0 ;
  assign n4094 = n4093 ^ n4092 ^ n2219 ;
  assign n4098 = n1602 & ~n4017 ;
  assign n4095 = x60 & ~n1424 ;
  assign n4096 = n4095 ^ n1119 ^ 1'b0 ;
  assign n4097 = n4096 ^ n1354 ^ 1'b0 ;
  assign n4099 = n4098 ^ n4097 ^ 1'b0 ;
  assign n4100 = n1736 | n4099 ;
  assign n4102 = n1643 ^ n842 ^ n168 ;
  assign n4101 = n1368 ^ n1234 ^ n730 ;
  assign n4103 = n4102 ^ n4101 ^ n1706 ;
  assign n4105 = n2506 ^ n2471 ^ n1098 ;
  assign n4104 = ~n253 & n2526 ;
  assign n4106 = n4105 ^ n4104 ^ 1'b0 ;
  assign n4107 = ( n744 & n4103 ) | ( n744 & n4106 ) | ( n4103 & n4106 ) ;
  assign n4108 = ( n1090 & ~n2470 ) | ( n1090 & n4107 ) | ( ~n2470 & n4107 ) ;
  assign n4113 = n1800 ^ n1361 ^ 1'b0 ;
  assign n4114 = n1386 & n4113 ;
  assign n4115 = ( n1335 & n3728 ) | ( n1335 & ~n4114 ) | ( n3728 & ~n4114 ) ;
  assign n4111 = ~n790 & n939 ;
  assign n4112 = ~x49 & n4111 ;
  assign n4109 = n1055 ^ n957 ^ n267 ;
  assign n4110 = n4109 ^ n3184 ^ n209 ;
  assign n4116 = n4115 ^ n4112 ^ n4110 ;
  assign n4117 = n738 | n2808 ;
  assign n4118 = n3115 & ~n4117 ;
  assign n4120 = ( n294 & n1244 ) | ( n294 & ~n1514 ) | ( n1244 & ~n1514 ) ;
  assign n4121 = ( ~x121 & x124 ) | ( ~x121 & n4120 ) | ( x124 & n4120 ) ;
  assign n4119 = n1307 & n2008 ;
  assign n4122 = n4121 ^ n4119 ^ 1'b0 ;
  assign n4123 = ( ~n204 & n974 ) | ( ~n204 & n1800 ) | ( n974 & n1800 ) ;
  assign n4124 = n3516 ^ n1974 ^ 1'b0 ;
  assign n4125 = n4123 & n4124 ;
  assign n4127 = n4041 ^ n1566 ^ 1'b0 ;
  assign n4126 = ~n225 & n2371 ;
  assign n4128 = n4127 ^ n4126 ^ 1'b0 ;
  assign n4129 = ( n1872 & ~n3068 ) | ( n1872 & n4128 ) | ( ~n3068 & n4128 ) ;
  assign n4130 = ( ~n1086 & n2812 ) | ( ~n1086 & n4129 ) | ( n2812 & n4129 ) ;
  assign n4131 = n1577 ^ n1565 ^ 1'b0 ;
  assign n4132 = x90 & n4131 ;
  assign n4133 = n3806 ^ n1394 ^ 1'b0 ;
  assign n4134 = ( n3356 & n4132 ) | ( n3356 & n4133 ) | ( n4132 & n4133 ) ;
  assign n4137 = n2643 ^ n1956 ^ n1498 ;
  assign n4135 = n536 & n1844 ;
  assign n4136 = n2765 | n4135 ;
  assign n4138 = n4137 ^ n4136 ^ 1'b0 ;
  assign n4144 = ( n413 & n1553 ) | ( n413 & n3744 ) | ( n1553 & n3744 ) ;
  assign n4141 = ~n364 & n746 ;
  assign n4142 = n4141 ^ n1823 ^ 1'b0 ;
  assign n4139 = n1388 ^ n815 ^ 1'b0 ;
  assign n4140 = n4139 ^ n1269 ^ 1'b0 ;
  assign n4143 = n4142 ^ n4140 ^ n1466 ;
  assign n4145 = n4144 ^ n4143 ^ n3312 ;
  assign n4146 = n253 ^ n236 ^ 1'b0 ;
  assign n4147 = n2681 ^ n512 ^ x44 ;
  assign n4148 = x0 & ~x6 ;
  assign n4149 = ( n2808 & n4147 ) | ( n2808 & ~n4148 ) | ( n4147 & ~n4148 ) ;
  assign n4150 = ( n1791 & n2736 ) | ( n1791 & n4149 ) | ( n2736 & n4149 ) ;
  assign n4151 = n650 | n1153 ;
  assign n4152 = ( n3220 & n4150 ) | ( n3220 & ~n4151 ) | ( n4150 & ~n4151 ) ;
  assign n4153 = n402 | n4152 ;
  assign n4154 = n1543 | n4153 ;
  assign n4155 = n822 & n4154 ;
  assign n4162 = n1777 ^ n300 ^ x31 ;
  assign n4163 = n2329 & n4162 ;
  assign n4156 = n3372 ^ n1146 ^ 1'b0 ;
  assign n4157 = n1708 & n4156 ;
  assign n4158 = ( n2301 & n2548 ) | ( n2301 & ~n4157 ) | ( n2548 & ~n4157 ) ;
  assign n4159 = ( n1344 & n1645 ) | ( n1344 & ~n4158 ) | ( n1645 & ~n4158 ) ;
  assign n4160 = ~n801 & n1255 ;
  assign n4161 = ~n4159 & n4160 ;
  assign n4164 = n4163 ^ n4161 ^ n2057 ;
  assign n4165 = ( n1083 & n3026 ) | ( n1083 & n4073 ) | ( n3026 & n4073 ) ;
  assign n4166 = n3410 & n4165 ;
  assign n4169 = n777 ^ n437 ^ n284 ;
  assign n4167 = ~n975 & n1570 ;
  assign n4168 = n586 & n4167 ;
  assign n4170 = n4169 ^ n4168 ^ 1'b0 ;
  assign n4171 = x2 & n1012 ;
  assign n4172 = n4171 ^ n815 ^ 1'b0 ;
  assign n4173 = n4172 ^ n4169 ^ 1'b0 ;
  assign n4174 = ( n522 & n3409 ) | ( n522 & ~n4173 ) | ( n3409 & ~n4173 ) ;
  assign n4175 = x55 & ~n2807 ;
  assign n4176 = ( ~n235 & n1455 ) | ( ~n235 & n3243 ) | ( n1455 & n3243 ) ;
  assign n4177 = n2553 | n2985 ;
  assign n4178 = n4177 ^ n2676 ^ 1'b0 ;
  assign n4179 = n428 & ~n4178 ;
  assign n4180 = ( ~n518 & n2438 ) | ( ~n518 & n4179 ) | ( n2438 & n4179 ) ;
  assign n4181 = ~n4176 & n4180 ;
  assign n4182 = n645 & ~n4181 ;
  assign n4183 = ( x88 & n2306 ) | ( x88 & n3812 ) | ( n2306 & n3812 ) ;
  assign n4184 = n1307 & n4183 ;
  assign n4185 = n2450 ^ n1633 ^ n787 ;
  assign n4186 = n1655 & ~n4185 ;
  assign n4187 = n3640 ^ n2725 ^ 1'b0 ;
  assign n4188 = n4187 ^ n1798 ^ n199 ;
  assign n4189 = n4186 & ~n4188 ;
  assign n4195 = n471 & n3037 ;
  assign n4190 = n1163 ^ n399 ^ 1'b0 ;
  assign n4191 = n4190 ^ n1758 ^ x59 ;
  assign n4192 = n4191 ^ n2634 ^ n1910 ;
  assign n4193 = n4192 ^ n136 ^ 1'b0 ;
  assign n4194 = n1715 | n4193 ;
  assign n4196 = n4195 ^ n4194 ^ 1'b0 ;
  assign n4197 = ( n1644 & ~n3909 ) | ( n1644 & n4196 ) | ( ~n3909 & n4196 ) ;
  assign n4198 = ( ~n1709 & n3169 ) | ( ~n1709 & n4197 ) | ( n3169 & n4197 ) ;
  assign n4199 = n3257 & ~n4198 ;
  assign n4200 = ~n4189 & n4199 ;
  assign n4202 = ~n413 & n865 ;
  assign n4201 = n2772 ^ n649 ^ 1'b0 ;
  assign n4203 = n4202 ^ n4201 ^ n2369 ;
  assign n4204 = n2827 ^ n2178 ^ 1'b0 ;
  assign n4206 = ~n392 & n1982 ;
  assign n4207 = ~n1506 & n4206 ;
  assign n4205 = n167 & n2122 ;
  assign n4208 = n4207 ^ n4205 ^ n3551 ;
  assign n4209 = ( n3464 & n4204 ) | ( n3464 & ~n4208 ) | ( n4204 & ~n4208 ) ;
  assign n4212 = ~n1004 & n3082 ;
  assign n4213 = ~n489 & n4212 ;
  assign n4214 = n1765 ^ x59 ^ 1'b0 ;
  assign n4215 = ( n1950 & n4213 ) | ( n1950 & n4214 ) | ( n4213 & n4214 ) ;
  assign n4216 = n4215 ^ n1341 ^ 1'b0 ;
  assign n4210 = n2144 | n3916 ;
  assign n4211 = n863 | n4210 ;
  assign n4217 = n4216 ^ n4211 ^ 1'b0 ;
  assign n4218 = ( n265 & n1129 ) | ( n265 & ~n1767 ) | ( n1129 & ~n1767 ) ;
  assign n4219 = n4218 ^ n1189 ^ 1'b0 ;
  assign n4220 = n189 | n3081 ;
  assign n4221 = ( ~n1310 & n1339 ) | ( ~n1310 & n3806 ) | ( n1339 & n3806 ) ;
  assign n4222 = ~n610 & n1046 ;
  assign n4223 = n1281 ^ n551 ^ 1'b0 ;
  assign n4224 = n4222 & ~n4223 ;
  assign n4225 = n1190 & n2509 ;
  assign n4226 = n4225 ^ n3668 ^ 1'b0 ;
  assign n4227 = n2695 | n4158 ;
  assign n4228 = n3395 & ~n4227 ;
  assign n4229 = ~n3940 & n4228 ;
  assign n4230 = ( ~x53 & n758 ) | ( ~x53 & n3645 ) | ( n758 & n3645 ) ;
  assign n4231 = n379 | n1431 ;
  assign n4232 = n1339 | n3626 ;
  assign n4233 = n4232 ^ n1122 ^ 1'b0 ;
  assign n4234 = n3339 ^ n1823 ^ n1623 ;
  assign n4235 = ( x120 & n337 ) | ( x120 & ~n4234 ) | ( n337 & ~n4234 ) ;
  assign n4236 = ( n3053 & n4233 ) | ( n3053 & ~n4235 ) | ( n4233 & ~n4235 ) ;
  assign n4237 = ( n2527 & n4231 ) | ( n2527 & ~n4236 ) | ( n4231 & ~n4236 ) ;
  assign n4238 = ( ~n512 & n1613 ) | ( ~n512 & n2934 ) | ( n1613 & n2934 ) ;
  assign n4239 = n2210 ^ n1700 ^ n1259 ;
  assign n4240 = n4239 ^ n692 ^ x95 ;
  assign n4241 = ~n4238 & n4240 ;
  assign n4242 = n2982 ^ n1483 ^ n1350 ;
  assign n4243 = n4242 ^ n4097 ^ 1'b0 ;
  assign n4244 = n660 & n1850 ;
  assign n4245 = n4244 ^ n999 ^ 1'b0 ;
  assign n4246 = ~n3209 & n4245 ;
  assign n4247 = ~n895 & n4246 ;
  assign n4249 = n1630 ^ n1336 ^ n1177 ;
  assign n4248 = n2838 ^ n926 ^ 1'b0 ;
  assign n4250 = n4249 ^ n4248 ^ n1871 ;
  assign n4251 = n881 & ~n4250 ;
  assign n4252 = n4247 & n4251 ;
  assign n4253 = ( x16 & x62 ) | ( x16 & n2218 ) | ( x62 & n2218 ) ;
  assign n4254 = n2684 & ~n4253 ;
  assign n4256 = n955 ^ n231 ^ 1'b0 ;
  assign n4255 = n1294 & ~n2306 ;
  assign n4257 = n4256 ^ n4255 ^ 1'b0 ;
  assign n4258 = n1426 | n4257 ;
  assign n4259 = n4258 ^ n2484 ^ 1'b0 ;
  assign n4260 = n549 & n2170 ;
  assign n4261 = n4260 ^ n3962 ^ 1'b0 ;
  assign n4262 = n1550 & ~n4261 ;
  assign n4263 = n762 & n891 ;
  assign n4264 = ~n806 & n4263 ;
  assign n4265 = ( ~n624 & n646 ) | ( ~n624 & n1847 ) | ( n646 & n1847 ) ;
  assign n4266 = n984 | n4265 ;
  assign n4267 = n4266 ^ n2331 ^ 1'b0 ;
  assign n4268 = n4267 ^ x30 ^ 1'b0 ;
  assign n4270 = ~n1020 & n2496 ;
  assign n4271 = n1304 & n4270 ;
  assign n4269 = ~n681 & n750 ;
  assign n4272 = n4271 ^ n4269 ^ 1'b0 ;
  assign n4273 = ( n951 & n2742 ) | ( n951 & n4272 ) | ( n2742 & n4272 ) ;
  assign n4274 = n4273 ^ n2081 ^ n392 ;
  assign n4275 = ( n214 & n1874 ) | ( n214 & ~n4274 ) | ( n1874 & ~n4274 ) ;
  assign n4276 = ( ~n4264 & n4268 ) | ( ~n4264 & n4275 ) | ( n4268 & n4275 ) ;
  assign n4277 = n4262 & n4276 ;
  assign n4278 = n4277 ^ n1656 ^ 1'b0 ;
  assign n4279 = ( ~n1707 & n4259 ) | ( ~n1707 & n4278 ) | ( n4259 & n4278 ) ;
  assign n4281 = ( n1069 & n1346 ) | ( n1069 & ~n2770 ) | ( n1346 & ~n2770 ) ;
  assign n4282 = ( n372 & ~n576 ) | ( n372 & n4281 ) | ( ~n576 & n4281 ) ;
  assign n4280 = n2855 ^ n1489 ^ n433 ;
  assign n4283 = n4282 ^ n4280 ^ n3018 ;
  assign n4284 = x81 & n2922 ;
  assign n4285 = ~n1409 & n4284 ;
  assign n4286 = n4285 ^ n3809 ^ n2488 ;
  assign n4289 = n2946 ^ n1405 ^ 1'b0 ;
  assign n4290 = n3817 & n4289 ;
  assign n4287 = n2832 ^ n2765 ^ n2475 ;
  assign n4288 = ( ~n561 & n1113 ) | ( ~n561 & n4287 ) | ( n1113 & n4287 ) ;
  assign n4291 = n4290 ^ n4288 ^ 1'b0 ;
  assign n4292 = n4052 | n4291 ;
  assign n4294 = ( n1977 & n2407 ) | ( n1977 & ~n3799 ) | ( n2407 & ~n3799 ) ;
  assign n4293 = n4267 ^ n1125 ^ n897 ;
  assign n4295 = n4294 ^ n4293 ^ 1'b0 ;
  assign n4296 = n709 | n4120 ;
  assign n4297 = n4296 ^ n2246 ^ 1'b0 ;
  assign n4298 = n2608 | n4297 ;
  assign n4299 = ~n2379 & n4298 ;
  assign n4300 = ~n2416 & n3832 ;
  assign n4301 = n4151 & n4300 ;
  assign n4302 = n3919 ^ n1597 ^ 1'b0 ;
  assign n4303 = n4302 ^ n3614 ^ 1'b0 ;
  assign n4304 = ( n253 & n706 ) | ( n253 & ~n1868 ) | ( n706 & ~n1868 ) ;
  assign n4305 = n990 | n4304 ;
  assign n4306 = n4305 ^ n2830 ^ n657 ;
  assign n4307 = n601 & n1621 ;
  assign n4311 = ( n203 & ~n878 ) | ( n203 & n2632 ) | ( ~n878 & n2632 ) ;
  assign n4309 = ~n659 & n3837 ;
  assign n4310 = ~n3993 & n4309 ;
  assign n4308 = n4239 ^ n1299 ^ n431 ;
  assign n4312 = n4311 ^ n4310 ^ n4308 ;
  assign n4313 = n846 | n4020 ;
  assign n4314 = n3157 | n4313 ;
  assign n4315 = n1804 ^ n748 ^ x102 ;
  assign n4316 = ~n2441 & n2704 ;
  assign n4317 = n4316 ^ n2276 ^ 1'b0 ;
  assign n4318 = x74 | n2392 ;
  assign n4319 = n3798 ^ n2042 ^ 1'b0 ;
  assign n4320 = ~n2723 & n4319 ;
  assign n4321 = ( n1149 & ~n1570 ) | ( n1149 & n4320 ) | ( ~n1570 & n4320 ) ;
  assign n4322 = ( ~n324 & n3214 ) | ( ~n324 & n4321 ) | ( n3214 & n4321 ) ;
  assign n4323 = n2527 ^ n2361 ^ 1'b0 ;
  assign n4324 = n1728 | n4323 ;
  assign n4325 = n2245 ^ n1964 ^ 1'b0 ;
  assign n4326 = ( n598 & n4324 ) | ( n598 & n4325 ) | ( n4324 & n4325 ) ;
  assign n4327 = ~n2520 & n4326 ;
  assign n4328 = n826 & n4327 ;
  assign n4329 = n4322 & ~n4328 ;
  assign n4330 = n4318 & ~n4329 ;
  assign n4331 = ~n4317 & n4330 ;
  assign n4332 = ( n1594 & n4315 ) | ( n1594 & n4331 ) | ( n4315 & n4331 ) ;
  assign n4333 = n3839 ^ n3199 ^ n773 ;
  assign n4334 = n4317 & n4333 ;
  assign n4335 = ( n696 & n1355 ) | ( n696 & n1736 ) | ( n1355 & n1736 ) ;
  assign n4336 = n1332 ^ n768 ^ n702 ;
  assign n4337 = ( n1268 & ~n2761 ) | ( n1268 & n4336 ) | ( ~n2761 & n4336 ) ;
  assign n4338 = ( n2543 & ~n4335 ) | ( n2543 & n4337 ) | ( ~n4335 & n4337 ) ;
  assign n4339 = n4338 ^ n2507 ^ n826 ;
  assign n4340 = n2378 & ~n2972 ;
  assign n4341 = n4340 ^ n2688 ^ 1'b0 ;
  assign n4342 = ( n954 & n2865 ) | ( n954 & n2914 ) | ( n2865 & n2914 ) ;
  assign n4343 = n4341 & n4342 ;
  assign n4344 = ( n1522 & n3099 ) | ( n1522 & ~n3488 ) | ( n3099 & ~n3488 ) ;
  assign n4345 = ( ~n962 & n4343 ) | ( ~n962 & n4344 ) | ( n4343 & n4344 ) ;
  assign n4346 = n171 | n2032 ;
  assign n4347 = n1068 & ~n4346 ;
  assign n4349 = n2535 ^ n2126 ^ n575 ;
  assign n4348 = n298 & ~n3735 ;
  assign n4350 = n4349 ^ n4348 ^ 1'b0 ;
  assign n4351 = ( n4275 & n4347 ) | ( n4275 & ~n4350 ) | ( n4347 & ~n4350 ) ;
  assign n4352 = x22 & ~x62 ;
  assign n4353 = n867 & n4352 ;
  assign n4354 = n3351 ^ n3231 ^ n179 ;
  assign n4355 = n1405 ^ n966 ^ 1'b0 ;
  assign n4356 = n2614 & ~n4355 ;
  assign n4357 = ( n857 & n1848 ) | ( n857 & n4356 ) | ( n1848 & n4356 ) ;
  assign n4358 = n1444 ^ n705 ^ 1'b0 ;
  assign n4359 = n4358 ^ n2703 ^ 1'b0 ;
  assign n4360 = n4357 & ~n4359 ;
  assign n4361 = ( n618 & n4354 ) | ( n618 & n4360 ) | ( n4354 & n4360 ) ;
  assign n4366 = n964 ^ n825 ^ n705 ;
  assign n4362 = n512 & n896 ;
  assign n4363 = n4362 ^ n906 ^ 1'b0 ;
  assign n4364 = n4363 ^ n2077 ^ 1'b0 ;
  assign n4365 = n2918 | n4364 ;
  assign n4367 = n4366 ^ n4365 ^ n4294 ;
  assign n4368 = n1609 | n1832 ;
  assign n4369 = n4368 ^ n3696 ^ 1'b0 ;
  assign n4371 = n631 & ~n794 ;
  assign n4372 = ~x22 & n4371 ;
  assign n4370 = n357 & n1419 ;
  assign n4373 = n4372 ^ n4370 ^ n2964 ;
  assign n4374 = ( n1573 & n3101 ) | ( n1573 & ~n3145 ) | ( n3101 & ~n3145 ) ;
  assign n4375 = ( ~n2713 & n2972 ) | ( ~n2713 & n3636 ) | ( n2972 & n3636 ) ;
  assign n4376 = ( n488 & n1212 ) | ( n488 & n4375 ) | ( n1212 & n4375 ) ;
  assign n4377 = ( ~n1082 & n3536 ) | ( ~n1082 & n4376 ) | ( n3536 & n4376 ) ;
  assign n4378 = n1422 & n4377 ;
  assign n4379 = n4374 | n4378 ;
  assign n4380 = n1427 | n4379 ;
  assign n4381 = ( n624 & ~n1364 ) | ( n624 & n1778 ) | ( ~n1364 & n1778 ) ;
  assign n4382 = n4381 ^ n3567 ^ x121 ;
  assign n4383 = ( n591 & n1099 ) | ( n591 & ~n1426 ) | ( n1099 & ~n1426 ) ;
  assign n4384 = ( n3755 & ~n3800 ) | ( n3755 & n4383 ) | ( ~n3800 & n4383 ) ;
  assign n4385 = n1683 & ~n4384 ;
  assign n4386 = n195 | n319 ;
  assign n4387 = n4386 ^ n1171 ^ 1'b0 ;
  assign n4388 = ~n2380 & n4387 ;
  assign n4389 = ~n1217 & n1847 ;
  assign n4390 = n4389 ^ n2308 ^ 1'b0 ;
  assign n4391 = n4390 ^ n2178 ^ n1794 ;
  assign n4392 = ( ~n2816 & n4388 ) | ( ~n2816 & n4391 ) | ( n4388 & n4391 ) ;
  assign n4393 = ~n157 & n2203 ;
  assign n4394 = n1026 & n4393 ;
  assign n4395 = n4201 ^ n1288 ^ 1'b0 ;
  assign n4396 = n3447 | n4395 ;
  assign n4397 = ( ~x65 & n788 ) | ( ~x65 & n4190 ) | ( n788 & n4190 ) ;
  assign n4398 = ~n1552 & n1844 ;
  assign n4399 = ~x53 & n4398 ;
  assign n4400 = n4399 ^ n1933 ^ 1'b0 ;
  assign n4401 = n474 | n4400 ;
  assign n4402 = ( x30 & ~n967 ) | ( x30 & n1524 ) | ( ~n967 & n1524 ) ;
  assign n4403 = n4402 ^ n1534 ^ n319 ;
  assign n4404 = ( n3435 & ~n4401 ) | ( n3435 & n4403 ) | ( ~n4401 & n4403 ) ;
  assign n4405 = n2014 ^ n1441 ^ 1'b0 ;
  assign n4406 = n1702 ^ n1286 ^ x35 ;
  assign n4407 = n445 & ~n2378 ;
  assign n4408 = ( n136 & n416 ) | ( n136 & n2712 ) | ( n416 & n2712 ) ;
  assign n4409 = ~n3004 & n4408 ;
  assign n4410 = ~n4250 & n4409 ;
  assign n4411 = n4407 & n4410 ;
  assign n4414 = n1395 ^ n1180 ^ n165 ;
  assign n4412 = ( n1269 & n1991 ) | ( n1269 & n2010 ) | ( n1991 & n2010 ) ;
  assign n4413 = n2105 & n4412 ;
  assign n4415 = n4414 ^ n4413 ^ 1'b0 ;
  assign n4416 = n433 | n1653 ;
  assign n4417 = ~n1719 & n4416 ;
  assign n4420 = n2944 ^ x33 ^ 1'b0 ;
  assign n4421 = n1051 | n4163 ;
  assign n4422 = n4421 ^ n1357 ^ 1'b0 ;
  assign n4423 = n4420 & n4422 ;
  assign n4424 = n2446 & n4423 ;
  assign n4425 = n4424 ^ n3385 ^ 1'b0 ;
  assign n4418 = n4304 ^ n1442 ^ 1'b0 ;
  assign n4419 = ~n1395 & n4418 ;
  assign n4426 = n4425 ^ n4419 ^ 1'b0 ;
  assign n4427 = n4426 ^ x114 ^ 1'b0 ;
  assign n4428 = n1496 & ~n4427 ;
  assign n4429 = n2171 ^ n1630 ^ n442 ;
  assign n4430 = ~n1378 & n4421 ;
  assign n4431 = n4430 ^ n2628 ^ 1'b0 ;
  assign n4446 = n607 & ~n2256 ;
  assign n4447 = ~n1554 & n4446 ;
  assign n4441 = n1355 ^ n1071 ^ 1'b0 ;
  assign n4442 = ~n593 & n4441 ;
  assign n4443 = n2978 ^ n1731 ^ n633 ;
  assign n4444 = n4442 & n4443 ;
  assign n4445 = n4444 ^ n3221 ^ 1'b0 ;
  assign n4448 = n4447 ^ n4445 ^ 1'b0 ;
  assign n4449 = n4448 ^ n2795 ^ n2323 ;
  assign n4432 = n1940 ^ n1647 ^ 1'b0 ;
  assign n4433 = n4432 ^ n3603 ^ 1'b0 ;
  assign n4434 = ~n1375 & n4433 ;
  assign n4435 = ~n168 & n4434 ;
  assign n4436 = n4435 ^ n3186 ^ 1'b0 ;
  assign n4437 = n1584 ^ n867 ^ 1'b0 ;
  assign n4438 = n468 | n4437 ;
  assign n4439 = n4436 & ~n4438 ;
  assign n4440 = n4439 ^ x61 ^ 1'b0 ;
  assign n4450 = n4449 ^ n4440 ^ 1'b0 ;
  assign n4451 = ~n1811 & n3243 ;
  assign n4452 = ( n410 & ~n1867 ) | ( n410 & n4451 ) | ( ~n1867 & n4451 ) ;
  assign n4453 = n3240 & n3827 ;
  assign n4454 = n4453 ^ n3187 ^ 1'b0 ;
  assign n4455 = n1040 & ~n4454 ;
  assign n4457 = n2237 ^ n378 ^ 1'b0 ;
  assign n4456 = n4162 ^ n1742 ^ n747 ;
  assign n4458 = n4457 ^ n4456 ^ n3998 ;
  assign n4459 = n3522 ^ n260 ^ 1'b0 ;
  assign n4460 = n720 & ~n4459 ;
  assign n4461 = ( n3261 & ~n4458 ) | ( n3261 & n4460 ) | ( ~n4458 & n4460 ) ;
  assign n4462 = n4461 ^ n1356 ^ 1'b0 ;
  assign n4463 = ( n2090 & ~n2260 ) | ( n2090 & n4462 ) | ( ~n2260 & n4462 ) ;
  assign n4464 = n1055 & n3209 ;
  assign n4465 = n155 & ~n1411 ;
  assign n4469 = ( n190 & ~n1375 ) | ( n190 & n1506 ) | ( ~n1375 & n1506 ) ;
  assign n4470 = n387 & n3263 ;
  assign n4471 = n4469 & n4470 ;
  assign n4466 = n3184 ^ n477 ^ 1'b0 ;
  assign n4467 = n854 & ~n4466 ;
  assign n4468 = n4467 ^ n3818 ^ n2026 ;
  assign n4472 = n4471 ^ n4468 ^ n355 ;
  assign n4473 = n2464 ^ n1734 ^ 1'b0 ;
  assign n4474 = x124 & ~n4473 ;
  assign n4475 = n4343 ^ n159 ^ 1'b0 ;
  assign n4477 = ( n1734 & n2207 ) | ( n1734 & ~n3312 ) | ( n2207 & ~n3312 ) ;
  assign n4476 = n2390 & n3074 ;
  assign n4478 = n4477 ^ n4476 ^ 1'b0 ;
  assign n4479 = ~n402 & n4164 ;
  assign n4480 = n416 | n2218 ;
  assign n4481 = ~n3365 & n4480 ;
  assign n4482 = n4481 ^ n611 ^ 1'b0 ;
  assign n4483 = n1697 | n4482 ;
  assign n4484 = n3709 & ~n4483 ;
  assign n4485 = n3678 ^ n453 ^ 1'b0 ;
  assign n4486 = n319 | n4485 ;
  assign n4487 = n1029 | n4486 ;
  assign n4488 = n4487 ^ n134 ^ 1'b0 ;
  assign n4489 = n4488 ^ n1901 ^ n1188 ;
  assign n4492 = ~n1093 & n1412 ;
  assign n4490 = ~n1912 & n2241 ;
  assign n4491 = n4490 ^ n1748 ^ n186 ;
  assign n4493 = n4492 ^ n4491 ^ x44 ;
  assign n4494 = n3013 ^ x113 ^ 1'b0 ;
  assign n4495 = n659 | n1433 ;
  assign n4496 = n4495 ^ n407 ^ 1'b0 ;
  assign n4497 = ~x17 & n4496 ;
  assign n4511 = n894 ^ n326 ^ n137 ;
  assign n4512 = n4511 ^ n3898 ^ n480 ;
  assign n4506 = n1758 ^ n1626 ^ n1106 ;
  assign n4507 = n2283 & n4506 ;
  assign n4508 = n4507 ^ n3217 ^ 1'b0 ;
  assign n4504 = n3636 ^ n773 ^ 1'b0 ;
  assign n4505 = n1772 | n4504 ;
  assign n4498 = n2347 ^ n311 ^ 1'b0 ;
  assign n4499 = n161 & ~n4498 ;
  assign n4500 = n385 & n4499 ;
  assign n4501 = ( n1573 & n3023 ) | ( n1573 & n4500 ) | ( n3023 & n4500 ) ;
  assign n4502 = n4501 ^ n562 ^ 1'b0 ;
  assign n4503 = ~n2236 & n4502 ;
  assign n4509 = n4508 ^ n4505 ^ n4503 ;
  assign n4510 = n1475 & n4509 ;
  assign n4513 = n4512 ^ n4510 ^ 1'b0 ;
  assign n4514 = ( ~n374 & n1528 ) | ( ~n374 & n1971 ) | ( n1528 & n1971 ) ;
  assign n4515 = ( x24 & n586 ) | ( x24 & ~n773 ) | ( n586 & ~n773 ) ;
  assign n4516 = ( n3473 & n3603 ) | ( n3473 & ~n4515 ) | ( n3603 & ~n4515 ) ;
  assign n4517 = n4514 | n4516 ;
  assign n4518 = n1875 | n4517 ;
  assign n4519 = n2058 & n2344 ;
  assign n4520 = n4519 ^ n586 ^ 1'b0 ;
  assign n4521 = n1050 & n4520 ;
  assign n4522 = ~n1720 & n4521 ;
  assign n4523 = ~n479 & n2375 ;
  assign n4524 = n4523 ^ n3880 ^ 1'b0 ;
  assign n4525 = ( x107 & n1488 ) | ( x107 & ~n1553 ) | ( n1488 & ~n1553 ) ;
  assign n4526 = n3721 ^ n1517 ^ 1'b0 ;
  assign n4527 = n4525 & ~n4526 ;
  assign n4528 = ( n1210 & n2482 ) | ( n1210 & ~n4500 ) | ( n2482 & ~n4500 ) ;
  assign n4529 = n243 | n468 ;
  assign n4530 = n4210 & ~n4529 ;
  assign n4531 = n4528 | n4530 ;
  assign n4532 = n2358 ^ n2046 ^ n802 ;
  assign n4533 = n2360 ^ n541 ^ 1'b0 ;
  assign n4534 = n3806 & ~n4533 ;
  assign n4535 = n2608 ^ n1010 ^ x63 ;
  assign n4536 = ( ~x117 & n2902 ) | ( ~x117 & n3697 ) | ( n2902 & n3697 ) ;
  assign n4537 = ( n1853 & n4535 ) | ( n1853 & n4536 ) | ( n4535 & n4536 ) ;
  assign n4538 = ( n2088 & ~n4491 ) | ( n2088 & n4537 ) | ( ~n4491 & n4537 ) ;
  assign n4539 = n4534 & n4538 ;
  assign n4540 = n4539 ^ n4224 ^ n249 ;
  assign n4541 = n2941 & n3668 ;
  assign n4542 = ( x68 & ~n1078 ) | ( x68 & n1268 ) | ( ~n1078 & n1268 ) ;
  assign n4543 = n1287 & n1828 ;
  assign n4544 = ( ~n3688 & n4542 ) | ( ~n3688 & n4543 ) | ( n4542 & n4543 ) ;
  assign n4545 = n1184 ^ n1176 ^ 1'b0 ;
  assign n4546 = n1068 ^ n557 ^ n159 ;
  assign n4547 = n2962 ^ n503 ^ 1'b0 ;
  assign n4548 = ~n4164 & n4547 ;
  assign n4549 = n4548 ^ n2684 ^ 1'b0 ;
  assign n4550 = ( n1894 & n4546 ) | ( n1894 & n4549 ) | ( n4546 & n4549 ) ;
  assign n4552 = ( n219 & ~n289 ) | ( n219 & n1443 ) | ( ~n289 & n1443 ) ;
  assign n4553 = ( n1021 & ~n2325 ) | ( n1021 & n4552 ) | ( ~n2325 & n4552 ) ;
  assign n4551 = n2146 & n3701 ;
  assign n4554 = n4553 ^ n4551 ^ n3973 ;
  assign n4555 = ( n170 & n1137 ) | ( n170 & n1989 ) | ( n1137 & n1989 ) ;
  assign n4556 = n4555 ^ n4544 ^ 1'b0 ;
  assign n4564 = n628 & ~n1794 ;
  assign n4565 = n2227 & ~n4564 ;
  assign n4566 = ~n1980 & n4565 ;
  assign n4557 = n329 & ~n1886 ;
  assign n4558 = n4557 ^ n741 ^ 1'b0 ;
  assign n4559 = n4558 ^ n2369 ^ 1'b0 ;
  assign n4560 = ( ~n215 & n760 ) | ( ~n215 & n4559 ) | ( n760 & n4559 ) ;
  assign n4561 = x123 & ~n3227 ;
  assign n4562 = ~n4560 & n4561 ;
  assign n4563 = n2165 | n4562 ;
  assign n4567 = n4566 ^ n4563 ^ 1'b0 ;
  assign n4568 = ( n310 & n1196 ) | ( n310 & n2245 ) | ( n1196 & n2245 ) ;
  assign n4569 = n4567 | n4568 ;
  assign n4570 = n4569 ^ n1403 ^ 1'b0 ;
  assign n4571 = ~n492 & n3322 ;
  assign n4581 = n551 | n720 ;
  assign n4572 = ( n2717 & ~n2746 ) | ( n2717 & n2855 ) | ( ~n2746 & n2855 ) ;
  assign n4573 = n924 ^ n582 ^ 1'b0 ;
  assign n4574 = n956 & n4573 ;
  assign n4575 = n4574 ^ n1580 ^ n348 ;
  assign n4576 = n2209 ^ n1141 ^ 1'b0 ;
  assign n4577 = n4575 | n4576 ;
  assign n4578 = n1865 & ~n4577 ;
  assign n4579 = n2912 & ~n4578 ;
  assign n4580 = n4572 & n4579 ;
  assign n4582 = n4581 ^ n4580 ^ 1'b0 ;
  assign n4583 = n824 & n4582 ;
  assign n4585 = n2282 ^ n1306 ^ 1'b0 ;
  assign n4586 = n2974 ^ n953 ^ 1'b0 ;
  assign n4587 = n4585 & n4586 ;
  assign n4584 = n4352 ^ n3896 ^ n1904 ;
  assign n4588 = n4587 ^ n4584 ^ n532 ;
  assign n4599 = n512 | n2488 ;
  assign n4595 = n3021 ^ n2832 ^ 1'b0 ;
  assign n4596 = n1603 & n4595 ;
  assign n4597 = n1301 ^ n1244 ^ 1'b0 ;
  assign n4598 = n4596 & ~n4597 ;
  assign n4600 = n4599 ^ n4598 ^ 1'b0 ;
  assign n4601 = n1036 & n4600 ;
  assign n4589 = n1073 ^ n725 ^ n346 ;
  assign n4590 = n762 & ~n4589 ;
  assign n4591 = n4590 ^ n600 ^ 1'b0 ;
  assign n4592 = n4591 ^ n1541 ^ x118 ;
  assign n4593 = n4592 ^ n1151 ^ 1'b0 ;
  assign n4594 = n4593 ^ n3628 ^ n1500 ;
  assign n4602 = n4601 ^ n4594 ^ 1'b0 ;
  assign n4606 = n1312 | n1366 ;
  assign n4607 = n3583 & ~n4606 ;
  assign n4603 = n343 & n696 ;
  assign n4604 = n4603 ^ n2283 ^ 1'b0 ;
  assign n4605 = n1967 | n4604 ;
  assign n4608 = n4607 ^ n4605 ^ 1'b0 ;
  assign n4609 = n3186 ^ n2649 ^ 1'b0 ;
  assign n4610 = n4608 | n4609 ;
  assign n4611 = n4610 ^ n2837 ^ 1'b0 ;
  assign n4612 = ( n1073 & n2021 ) | ( n1073 & n4229 ) | ( n2021 & n4229 ) ;
  assign n4618 = n4036 ^ x70 ^ 1'b0 ;
  assign n4619 = ~n1932 & n4618 ;
  assign n4617 = n3536 ^ n1606 ^ n992 ;
  assign n4616 = ( n2159 & n2370 ) | ( n2159 & ~n3482 ) | ( n2370 & ~n3482 ) ;
  assign n4620 = n4619 ^ n4617 ^ n4616 ;
  assign n4614 = n3341 ^ n2485 ^ n1159 ;
  assign n4613 = ~n757 & n1154 ;
  assign n4615 = n4614 ^ n4613 ^ 1'b0 ;
  assign n4621 = n4620 ^ n4615 ^ n768 ;
  assign n4622 = n1130 & ~n4581 ;
  assign n4623 = n4622 ^ n2016 ^ 1'b0 ;
  assign n4624 = n1419 ^ n268 ^ 1'b0 ;
  assign n4625 = n4624 ^ n3805 ^ 1'b0 ;
  assign n4626 = n4074 & n4625 ;
  assign n4627 = n3651 ^ n2194 ^ 1'b0 ;
  assign n4628 = n3334 ^ n2346 ^ 1'b0 ;
  assign n4629 = n1553 | n4628 ;
  assign n4630 = n4629 ^ n2813 ^ n2154 ;
  assign n4631 = n4630 ^ n254 ^ 1'b0 ;
  assign n4632 = n4627 & ~n4631 ;
  assign n4633 = n1522 | n2335 ;
  assign n4634 = n815 | n4633 ;
  assign n4635 = n4634 ^ n4510 ^ n1514 ;
  assign n4636 = ( n1965 & n4632 ) | ( n1965 & n4635 ) | ( n4632 & n4635 ) ;
  assign n4637 = ~n2931 & n3412 ;
  assign n4638 = n4637 ^ n4416 ^ 1'b0 ;
  assign n4639 = n2317 & n2607 ;
  assign n4640 = n1429 ^ n1155 ^ 1'b0 ;
  assign n4642 = ( n1136 & n1971 ) | ( n1136 & ~n3436 ) | ( n1971 & ~n3436 ) ;
  assign n4641 = ( n2291 & n2689 ) | ( n2291 & ~n4280 ) | ( n2689 & ~n4280 ) ;
  assign n4643 = n4642 ^ n4641 ^ 1'b0 ;
  assign n4644 = ( n1720 & n4640 ) | ( n1720 & n4643 ) | ( n4640 & n4643 ) ;
  assign n4645 = n3495 & ~n4644 ;
  assign n4646 = n2577 ^ n859 ^ 1'b0 ;
  assign n4647 = n3184 & ~n4646 ;
  assign n4648 = n1342 | n4647 ;
  assign n4649 = n3519 | n4648 ;
  assign n4650 = ~n275 & n953 ;
  assign n4651 = n913 & ~n4650 ;
  assign n4652 = n1486 & n4587 ;
  assign n4653 = n2399 & n2507 ;
  assign n4654 = n4653 ^ n3081 ^ 1'b0 ;
  assign n4655 = n4654 ^ n3062 ^ n2355 ;
  assign n4656 = n1225 & ~n3475 ;
  assign n4657 = n4656 ^ n3522 ^ 1'b0 ;
  assign n4658 = n399 & n4657 ;
  assign n4659 = ( n150 & n509 ) | ( n150 & ~n1082 ) | ( n509 & ~n1082 ) ;
  assign n4660 = ( n2539 & n4414 ) | ( n2539 & ~n4659 ) | ( n4414 & ~n4659 ) ;
  assign n4661 = ( x20 & n1393 ) | ( x20 & n3160 ) | ( n1393 & n3160 ) ;
  assign n4662 = x59 & n3195 ;
  assign n4663 = ~n3265 & n4662 ;
  assign n4664 = n3016 | n4663 ;
  assign n4665 = n4661 & ~n4664 ;
  assign n4669 = ( n2142 & n3579 ) | ( n2142 & n4036 ) | ( n3579 & n4036 ) ;
  assign n4666 = ( ~x47 & x99 ) | ( ~x47 & n263 ) | ( x99 & n263 ) ;
  assign n4667 = ( n249 & n3150 ) | ( n249 & n4666 ) | ( n3150 & n4666 ) ;
  assign n4668 = n1163 | n4667 ;
  assign n4670 = n4669 ^ n4668 ^ 1'b0 ;
  assign n4671 = ( ~n4503 & n4587 ) | ( ~n4503 & n4670 ) | ( n4587 & n4670 ) ;
  assign n4672 = ( n1259 & n1982 ) | ( n1259 & n4311 ) | ( n1982 & n4311 ) ;
  assign n4674 = ( ~n234 & n798 ) | ( ~n234 & n1406 ) | ( n798 & n1406 ) ;
  assign n4673 = n771 & ~n937 ;
  assign n4675 = n4674 ^ n4673 ^ 1'b0 ;
  assign n4676 = x25 & n4675 ;
  assign n4677 = n4676 ^ n1237 ^ 1'b0 ;
  assign n4679 = ( n836 & n1657 ) | ( n836 & ~n3812 ) | ( n1657 & ~n3812 ) ;
  assign n4680 = n1012 | n2743 ;
  assign n4681 = n4680 ^ n813 ^ 1'b0 ;
  assign n4682 = n4679 | n4681 ;
  assign n4683 = n1936 | n4682 ;
  assign n4678 = n4202 ^ n2394 ^ 1'b0 ;
  assign n4684 = n4683 ^ n4678 ^ n4629 ;
  assign n4685 = ( n4672 & n4677 ) | ( n4672 & ~n4684 ) | ( n4677 & ~n4684 ) ;
  assign n4686 = n3164 ^ n1117 ^ 1'b0 ;
  assign n4687 = n447 | n4686 ;
  assign n4688 = ( n1933 & n3882 ) | ( n1933 & ~n4163 ) | ( n3882 & ~n4163 ) ;
  assign n4690 = n589 | n1713 ;
  assign n4691 = ( n2030 & ~n4558 ) | ( n2030 & n4690 ) | ( ~n4558 & n4690 ) ;
  assign n4692 = n2301 & n4691 ;
  assign n4693 = n1128 & n4692 ;
  assign n4689 = ~n984 & n3111 ;
  assign n4694 = n4693 ^ n4689 ^ n747 ;
  assign n4695 = n2190 ^ n788 ^ n570 ;
  assign n4696 = n4695 ^ n4375 ^ n2963 ;
  assign n4697 = n4694 | n4696 ;
  assign n4698 = ( n4687 & ~n4688 ) | ( n4687 & n4697 ) | ( ~n4688 & n4697 ) ;
  assign n4699 = n645 | n2931 ;
  assign n4700 = ( ~n943 & n2051 ) | ( ~n943 & n4699 ) | ( n2051 & n4699 ) ;
  assign n4701 = ( ~n1203 & n1936 ) | ( ~n1203 & n4230 ) | ( n1936 & n4230 ) ;
  assign n4702 = n4701 ^ n4037 ^ n1291 ;
  assign n4703 = ( ~n1488 & n4700 ) | ( ~n1488 & n4702 ) | ( n4700 & n4702 ) ;
  assign n4704 = ( n1374 & ~n3333 ) | ( n1374 & n3622 ) | ( ~n3333 & n3622 ) ;
  assign n4705 = n1078 ^ n426 ^ 1'b0 ;
  assign n4706 = ( ~n319 & n894 ) | ( ~n319 & n2237 ) | ( n894 & n2237 ) ;
  assign n4707 = ( ~n2130 & n4705 ) | ( ~n2130 & n4706 ) | ( n4705 & n4706 ) ;
  assign n4708 = ~n2103 & n3377 ;
  assign n4709 = n783 & n4708 ;
  assign n4710 = ( n4704 & ~n4707 ) | ( n4704 & n4709 ) | ( ~n4707 & n4709 ) ;
  assign n4711 = ( ~n1622 & n3707 ) | ( ~n1622 & n3804 ) | ( n3707 & n3804 ) ;
  assign n4712 = n1617 & n2073 ;
  assign n4713 = n2383 ^ n1301 ^ 1'b0 ;
  assign n4714 = n4713 ^ n4068 ^ 1'b0 ;
  assign n4717 = n3891 ^ n2325 ^ 1'b0 ;
  assign n4718 = n4717 ^ n559 ^ n277 ;
  assign n4719 = ( n388 & n4666 ) | ( n388 & ~n4718 ) | ( n4666 & ~n4718 ) ;
  assign n4715 = ( n381 & n1029 ) | ( n381 & ~n1068 ) | ( n1029 & ~n1068 ) ;
  assign n4716 = n4715 ^ n3106 ^ n1088 ;
  assign n4720 = n4719 ^ n4716 ^ n3104 ;
  assign n4728 = x50 & ~n850 ;
  assign n4729 = n1431 & n4728 ;
  assign n4726 = ( n1717 & n1890 ) | ( n1717 & ~n3160 ) | ( n1890 & ~n3160 ) ;
  assign n4727 = ~n3389 & n4726 ;
  assign n4723 = ( ~n1022 & n1102 ) | ( ~n1022 & n1622 ) | ( n1102 & n1622 ) ;
  assign n4721 = n2527 ^ n183 ^ 1'b0 ;
  assign n4722 = ( n2876 & n4498 ) | ( n2876 & n4721 ) | ( n4498 & n4721 ) ;
  assign n4724 = n4723 ^ n4722 ^ n2960 ;
  assign n4725 = n4614 & n4724 ;
  assign n4730 = n4729 ^ n4727 ^ n4725 ;
  assign n4731 = n1806 | n4157 ;
  assign n4732 = n4114 & n4731 ;
  assign n4733 = n586 | n4264 ;
  assign n4734 = n4733 ^ n1391 ^ n1158 ;
  assign n4735 = n726 & ~n1228 ;
  assign n4736 = n4735 ^ n3272 ^ 1'b0 ;
  assign n4737 = ( ~n1235 & n3288 ) | ( ~n1235 & n4191 ) | ( n3288 & n4191 ) ;
  assign n4738 = ( ~n1706 & n4736 ) | ( ~n1706 & n4737 ) | ( n4736 & n4737 ) ;
  assign n4749 = n618 & n2637 ;
  assign n4750 = n2237 & n4749 ;
  assign n4746 = n3835 ^ n879 ^ 1'b0 ;
  assign n4747 = n1809 | n4746 ;
  assign n4748 = ( n765 & n970 ) | ( n765 & ~n4747 ) | ( n970 & ~n4747 ) ;
  assign n4739 = ~n923 & n2336 ;
  assign n4740 = n3243 ^ n2303 ^ 1'b0 ;
  assign n4741 = n3776 & n4740 ;
  assign n4742 = n4739 & n4741 ;
  assign n4743 = n183 & ~n2642 ;
  assign n4744 = n4743 ^ n1233 ^ 1'b0 ;
  assign n4745 = n4742 | n4744 ;
  assign n4751 = n4750 ^ n4748 ^ n4745 ;
  assign n4753 = n767 | n3070 ;
  assign n4754 = ( n2151 & n3308 ) | ( n2151 & n4753 ) | ( n3308 & n4753 ) ;
  assign n4752 = ~n3256 & n4352 ;
  assign n4755 = n4754 ^ n4752 ^ 1'b0 ;
  assign n4756 = n716 | n4376 ;
  assign n4757 = n4755 | n4756 ;
  assign n4758 = n557 & ~n903 ;
  assign n4759 = n2661 ^ n2655 ^ n1532 ;
  assign n4760 = n4759 ^ n3534 ^ 1'b0 ;
  assign n4761 = ~n4758 & n4760 ;
  assign n4762 = n4615 | n4761 ;
  assign n4763 = n3812 & ~n4497 ;
  assign n4764 = n4530 & n4763 ;
  assign n4766 = ( n484 & ~n906 ) | ( n484 & n975 ) | ( ~n906 & n975 ) ;
  assign n4767 = ( x54 & n831 ) | ( x54 & ~n4766 ) | ( n831 & ~n4766 ) ;
  assign n4765 = n3510 ^ n2843 ^ n960 ;
  assign n4768 = n4767 ^ n4765 ^ 1'b0 ;
  assign n4769 = n2332 & ~n4768 ;
  assign n4770 = ~n199 & n2902 ;
  assign n4771 = n4770 ^ n2393 ^ 1'b0 ;
  assign n4772 = ( n1665 & n2919 ) | ( n1665 & n4771 ) | ( n2919 & n4771 ) ;
  assign n4773 = n1247 | n4772 ;
  assign n4774 = n1378 ^ n440 ^ 1'b0 ;
  assign n4775 = ( ~n1169 & n1620 ) | ( ~n1169 & n3808 ) | ( n1620 & n3808 ) ;
  assign n4776 = n1912 & ~n4775 ;
  assign n4777 = n3811 ^ n1434 ^ 1'b0 ;
  assign n4778 = x89 & ~n4777 ;
  assign n4779 = n1521 ^ n1063 ^ 1'b0 ;
  assign n4780 = n1205 | n4779 ;
  assign n4781 = n4304 | n4780 ;
  assign n4782 = n4677 & ~n4781 ;
  assign n4783 = n601 & n4139 ;
  assign n4784 = n1772 & n4783 ;
  assign n4785 = n2976 | n4501 ;
  assign n4786 = n1899 & ~n4785 ;
  assign n4787 = ( n2559 & n4456 ) | ( n2559 & ~n4786 ) | ( n4456 & ~n4786 ) ;
  assign n4788 = n1587 ^ n1041 ^ 1'b0 ;
  assign n4789 = n4464 ^ n3412 ^ 1'b0 ;
  assign n4790 = ~n4788 & n4789 ;
  assign n4791 = n3075 & ~n3656 ;
  assign n4792 = n4791 ^ n1933 ^ 1'b0 ;
  assign n4793 = ( n369 & n766 ) | ( n369 & n3033 ) | ( n766 & n3033 ) ;
  assign n4794 = ( n272 & n4472 ) | ( n272 & n4793 ) | ( n4472 & n4793 ) ;
  assign n4795 = n2530 ^ n951 ^ 1'b0 ;
  assign n4796 = ( n164 & n3044 ) | ( n164 & n4795 ) | ( n3044 & n4795 ) ;
  assign n4797 = n4515 & ~n4796 ;
  assign n4798 = n918 & n4797 ;
  assign n4799 = ~n1526 & n4033 ;
  assign n4800 = n576 & n4799 ;
  assign n4801 = n4800 ^ n1663 ^ n540 ;
  assign n4802 = n665 & ~n4801 ;
  assign n4803 = n4798 & n4802 ;
  assign n4804 = n2570 ^ n690 ^ 1'b0 ;
  assign n4805 = n4287 & ~n4804 ;
  assign n4806 = n3773 ^ n2048 ^ 1'b0 ;
  assign n4807 = n215 & n4806 ;
  assign n4808 = n1656 ^ x93 ^ 1'b0 ;
  assign n4809 = n4161 | n4808 ;
  assign n4810 = n4809 ^ n1196 ^ 1'b0 ;
  assign n4811 = n4810 ^ n3262 ^ n2828 ;
  assign n4812 = n4811 ^ n1852 ^ 1'b0 ;
  assign n4813 = n4666 ^ n442 ^ 1'b0 ;
  assign n4814 = ( n1971 & n2602 ) | ( n1971 & n3971 ) | ( n2602 & n3971 ) ;
  assign n4815 = ( n1558 & n2256 ) | ( n1558 & n3124 ) | ( n2256 & n3124 ) ;
  assign n4816 = ( n4813 & n4814 ) | ( n4813 & n4815 ) | ( n4814 & n4815 ) ;
  assign n4819 = n497 ^ n465 ^ x79 ;
  assign n4817 = n896 ^ n777 ^ 1'b0 ;
  assign n4818 = x0 & ~n4817 ;
  assign n4820 = n4819 ^ n4818 ^ n4767 ;
  assign n4821 = n4599 | n4820 ;
  assign n4822 = n4821 ^ n2052 ^ n1239 ;
  assign n4824 = ( n179 & n1572 ) | ( n179 & ~n1957 ) | ( n1572 & ~n1957 ) ;
  assign n4825 = n3797 & ~n4824 ;
  assign n4823 = n2747 & n3778 ;
  assign n4826 = n4825 ^ n4823 ^ 1'b0 ;
  assign n4827 = n1024 | n4826 ;
  assign n4828 = n388 & n3044 ;
  assign n4829 = n4828 ^ n551 ^ 1'b0 ;
  assign n4830 = n4829 ^ n1314 ^ 1'b0 ;
  assign n4831 = n3088 & n4830 ;
  assign n4832 = n155 & ~n4138 ;
  assign n4833 = n1361 | n3285 ;
  assign n4834 = n3906 | n4833 ;
  assign n4835 = n4834 ^ n2274 ^ 1'b0 ;
  assign n4836 = n519 & n4070 ;
  assign n4837 = n4836 ^ n1494 ^ 1'b0 ;
  assign n4838 = n3553 ^ n3026 ^ n660 ;
  assign n4839 = ( n1183 & n4654 ) | ( n1183 & n4838 ) | ( n4654 & n4838 ) ;
  assign n4840 = ~n1376 & n4839 ;
  assign n4841 = n157 & ~n1949 ;
  assign n4842 = n4841 ^ n1967 ^ n1382 ;
  assign n4843 = n631 & n4754 ;
  assign n4844 = ( n387 & n4842 ) | ( n387 & ~n4843 ) | ( n4842 & ~n4843 ) ;
  assign n4845 = n4844 ^ n2196 ^ 1'b0 ;
  assign n4846 = ~n4840 & n4845 ;
  assign n4847 = n4846 ^ n462 ^ 1'b0 ;
  assign n4848 = n4825 & ~n4847 ;
  assign n4849 = n4191 ^ n2091 ^ n1808 ;
  assign n4850 = ~n465 & n2647 ;
  assign n4851 = ~n4280 & n4850 ;
  assign n4852 = n1976 ^ x5 ^ 1'b0 ;
  assign n4853 = ( n4849 & ~n4851 ) | ( n4849 & n4852 ) | ( ~n4851 & n4852 ) ;
  assign n4854 = ( ~n1944 & n3471 ) | ( ~n1944 & n4041 ) | ( n3471 & n4041 ) ;
  assign n4855 = n4101 ^ n3876 ^ 1'b0 ;
  assign n4856 = n4855 ^ n4815 ^ n386 ;
  assign n4861 = n933 & n2346 ;
  assign n4862 = ( n770 & ~n1186 ) | ( n770 & n2106 ) | ( ~n1186 & n2106 ) ;
  assign n4863 = ( n2279 & ~n2335 ) | ( n2279 & n4862 ) | ( ~n2335 & n4862 ) ;
  assign n4864 = ( n1827 & n4861 ) | ( n1827 & ~n4863 ) | ( n4861 & ~n4863 ) ;
  assign n4857 = n1609 ^ n1589 ^ n846 ;
  assign n4858 = ( n2717 & n2900 ) | ( n2717 & ~n4857 ) | ( n2900 & ~n4857 ) ;
  assign n4859 = n4858 ^ n3184 ^ n2089 ;
  assign n4860 = ( ~x60 & n1336 ) | ( ~x60 & n4859 ) | ( n1336 & n4859 ) ;
  assign n4865 = n4864 ^ n4860 ^ 1'b0 ;
  assign n4866 = n369 & ~n469 ;
  assign n4867 = n4866 ^ n159 ^ 1'b0 ;
  assign n4868 = n1614 & n4867 ;
  assign n4869 = ( ~n1629 & n1660 ) | ( ~n1629 & n4617 ) | ( n1660 & n4617 ) ;
  assign n4870 = n4869 ^ n1507 ^ 1'b0 ;
  assign n4874 = n3360 ^ n2526 ^ n1217 ;
  assign n4872 = ( n912 & ~n1199 ) | ( n912 & n3182 ) | ( ~n1199 & n3182 ) ;
  assign n4873 = n1062 | n4872 ;
  assign n4875 = n4874 ^ n4873 ^ 1'b0 ;
  assign n4871 = ~n1151 & n4559 ;
  assign n4876 = n4875 ^ n4871 ^ 1'b0 ;
  assign n4877 = n4876 ^ n1539 ^ n1406 ;
  assign n4879 = n3566 ^ n1373 ^ x118 ;
  assign n4878 = n2495 ^ n1451 ^ n586 ;
  assign n4880 = n4879 ^ n4878 ^ 1'b0 ;
  assign n4881 = ~n916 & n4880 ;
  assign n4882 = n4881 ^ n1158 ^ 1'b0 ;
  assign n4883 = n871 & ~n4882 ;
  assign n4884 = n4883 ^ n2200 ^ n440 ;
  assign n4885 = ( n2259 & ~n3218 ) | ( n2259 & n4884 ) | ( ~n3218 & n4884 ) ;
  assign n4886 = ~n765 & n891 ;
  assign n4887 = ~n872 & n4886 ;
  assign n4888 = n1761 & ~n4887 ;
  assign n4889 = n4888 ^ n3540 ^ 1'b0 ;
  assign n4890 = n4889 ^ n1910 ^ x55 ;
  assign n4891 = n4890 ^ n3273 ^ n1611 ;
  assign n4892 = n2745 ^ n506 ^ 1'b0 ;
  assign n4893 = n2081 & n4892 ;
  assign n4895 = n4358 ^ x81 ^ 1'b0 ;
  assign n4894 = n1269 & ~n1657 ;
  assign n4896 = n4895 ^ n4894 ^ 1'b0 ;
  assign n4897 = n1543 & n4896 ;
  assign n4898 = ~n3053 & n4897 ;
  assign n4899 = ( n2057 & ~n2833 ) | ( n2057 & n3639 ) | ( ~n2833 & n3639 ) ;
  assign n4900 = ( n1147 & ~n2638 ) | ( n1147 & n2978 ) | ( ~n2638 & n2978 ) ;
  assign n4901 = n3077 ^ n1573 ^ 1'b0 ;
  assign n4902 = n4900 | n4901 ;
  assign n4903 = ( n1755 & n3674 ) | ( n1755 & ~n4902 ) | ( n3674 & ~n4902 ) ;
  assign n4904 = n2906 & n3776 ;
  assign n4905 = n2444 & ~n4795 ;
  assign n4906 = ( n1439 & ~n4163 ) | ( n1439 & n4905 ) | ( ~n4163 & n4905 ) ;
  assign n4907 = n3024 | n4906 ;
  assign n4908 = n4907 ^ n2289 ^ 1'b0 ;
  assign n4909 = n4813 ^ n1707 ^ 1'b0 ;
  assign n4910 = n2021 & ~n4909 ;
  assign n4911 = ( n547 & n633 ) | ( n547 & n876 ) | ( n633 & n876 ) ;
  assign n4912 = n980 ^ n338 ^ 1'b0 ;
  assign n4913 = n2794 & ~n4912 ;
  assign n4914 = n4207 ^ n1841 ^ n141 ;
  assign n4915 = n4913 & n4914 ;
  assign n4916 = n4911 & n4915 ;
  assign n4917 = n4356 ^ n1220 ^ n260 ;
  assign n4918 = ( n177 & n2282 ) | ( n177 & ~n4917 ) | ( n2282 & ~n4917 ) ;
  assign n4919 = n4918 ^ n1650 ^ 1'b0 ;
  assign n4920 = n4919 ^ n3349 ^ 1'b0 ;
  assign n4921 = n2103 ^ n713 ^ 1'b0 ;
  assign n4922 = n4921 ^ n3252 ^ 1'b0 ;
  assign n4923 = x17 & n1659 ;
  assign n4924 = n4923 ^ n2388 ^ 1'b0 ;
  assign n4925 = n1380 & ~n3809 ;
  assign n4926 = n4925 ^ n3544 ^ 1'b0 ;
  assign n4927 = n4924 & ~n4926 ;
  assign n4928 = n4375 ^ n4144 ^ 1'b0 ;
  assign n4929 = n4927 & n4928 ;
  assign n4930 = ( n265 & n1220 ) | ( n265 & n1914 ) | ( n1220 & n1914 ) ;
  assign n4931 = n4930 ^ n2555 ^ n859 ;
  assign n4932 = n4931 ^ n3204 ^ n2075 ;
  assign n4933 = ( n1763 & ~n2840 ) | ( n1763 & n4669 ) | ( ~n2840 & n4669 ) ;
  assign n4934 = x2 | n4933 ;
  assign n4935 = n4059 ^ n1334 ^ 1'b0 ;
  assign n4936 = x72 & ~n4935 ;
  assign n4937 = n4936 ^ n3054 ^ 1'b0 ;
  assign n4938 = n4818 & ~n4937 ;
  assign n4939 = n1639 & n4938 ;
  assign n4940 = n4939 ^ n510 ^ 1'b0 ;
  assign n4941 = n4940 ^ n4065 ^ 1'b0 ;
  assign n4942 = n4934 & n4941 ;
  assign n4943 = n4942 ^ n1777 ^ 1'b0 ;
  assign n4944 = n4036 ^ n859 ^ 1'b0 ;
  assign n4945 = ~n2251 & n2946 ;
  assign n4946 = ~n2087 & n4945 ;
  assign n4947 = n2241 | n4946 ;
  assign n4948 = n2622 ^ n2523 ^ n1900 ;
  assign n4949 = n4948 ^ n4572 ^ 1'b0 ;
  assign n4950 = ( ~n531 & n2179 ) | ( ~n531 & n4229 ) | ( n2179 & n4229 ) ;
  assign n4951 = ( ~n1806 & n1978 ) | ( ~n1806 & n2837 ) | ( n1978 & n2837 ) ;
  assign n4952 = n2860 ^ n259 ^ 1'b0 ;
  assign n4953 = n4951 & ~n4952 ;
  assign n4954 = n4953 ^ n4734 ^ n3186 ;
  assign n4955 = n3142 & ~n4954 ;
  assign n4956 = n4955 ^ n2857 ^ 1'b0 ;
  assign n4957 = n1282 ^ n929 ^ n910 ;
  assign n4958 = n3800 | n4957 ;
  assign n4959 = n4958 ^ n1655 ^ 1'b0 ;
  assign n4960 = n1355 & n3589 ;
  assign n4961 = ( ~n729 & n1496 ) | ( ~n729 & n4766 ) | ( n1496 & n4766 ) ;
  assign n4962 = ( n4959 & ~n4960 ) | ( n4959 & n4961 ) | ( ~n4960 & n4961 ) ;
  assign n4963 = ~n1468 & n3200 ;
  assign n4964 = ~n4962 & n4963 ;
  assign n4965 = n4560 ^ n351 ^ 1'b0 ;
  assign n4966 = n2553 | n4965 ;
  assign n4967 = n4966 ^ n2523 ^ 1'b0 ;
  assign n4968 = n2273 & n2722 ;
  assign n4969 = ( n145 & n326 ) | ( n145 & ~n1334 ) | ( n326 & ~n1334 ) ;
  assign n4970 = ( n1299 & n2864 ) | ( n1299 & n4969 ) | ( n2864 & n4969 ) ;
  assign n4971 = ( n4967 & n4968 ) | ( n4967 & ~n4970 ) | ( n4968 & ~n4970 ) ;
  assign n4972 = n2994 ^ n579 ^ 1'b0 ;
  assign n4973 = ~n3712 & n4972 ;
  assign n4974 = n4207 ^ n2451 ^ 1'b0 ;
  assign n4975 = n2862 | n4974 ;
  assign n4982 = n913 | n3439 ;
  assign n4976 = ~n795 & n1405 ;
  assign n4977 = n3889 ^ n1286 ^ n315 ;
  assign n4978 = n980 | n4977 ;
  assign n4979 = n4978 ^ n4680 ^ 1'b0 ;
  assign n4980 = n4121 ^ n998 ^ n404 ;
  assign n4981 = ( n4976 & n4979 ) | ( n4976 & ~n4980 ) | ( n4979 & ~n4980 ) ;
  assign n4983 = n4982 ^ n4981 ^ 1'b0 ;
  assign n4984 = n3587 & n4983 ;
  assign n4985 = ( ~n282 & n1334 ) | ( ~n282 & n4589 ) | ( n1334 & n4589 ) ;
  assign n4986 = ( n1693 & n2756 ) | ( n1693 & n4985 ) | ( n2756 & n4985 ) ;
  assign n4987 = ( ~n822 & n3548 ) | ( ~n822 & n4986 ) | ( n3548 & n4986 ) ;
  assign n4988 = n1204 | n2466 ;
  assign n4989 = n4813 & ~n4988 ;
  assign n4990 = ( ~n939 & n1017 ) | ( ~n939 & n1114 ) | ( n1017 & n1114 ) ;
  assign n4991 = ( n2292 & n4989 ) | ( n2292 & n4990 ) | ( n4989 & n4990 ) ;
  assign n4992 = n4991 ^ n4482 ^ n4221 ;
  assign n4993 = n1684 ^ n1163 ^ n846 ;
  assign n4994 = n4993 ^ n3540 ^ 1'b0 ;
  assign n4995 = n4463 ^ n1169 ^ 1'b0 ;
  assign n4996 = n4994 | n4995 ;
  assign n4997 = ( ~n1196 & n3573 ) | ( ~n1196 & n4930 ) | ( n3573 & n4930 ) ;
  assign n4998 = n2325 ^ n1472 ^ 1'b0 ;
  assign n4999 = n3061 | n4998 ;
  assign n5000 = n401 & ~n452 ;
  assign n5001 = ~n4680 & n5000 ;
  assign n5002 = ( n572 & n1832 ) | ( n572 & n3947 ) | ( n1832 & n3947 ) ;
  assign n5003 = n4961 ^ n856 ^ 1'b0 ;
  assign n5007 = n2556 & ~n3530 ;
  assign n5008 = n3860 & n5007 ;
  assign n5004 = ~n1356 & n1997 ;
  assign n5005 = ~n656 & n5004 ;
  assign n5006 = n5005 ^ n2230 ^ n898 ;
  assign n5009 = n5008 ^ n5006 ^ n2426 ;
  assign n5010 = n5009 ^ n3880 ^ x95 ;
  assign n5011 = ~n1532 & n1597 ;
  assign n5012 = n5011 ^ n1045 ^ 1'b0 ;
  assign n5013 = n248 | n1830 ;
  assign n5014 = n5013 ^ n1695 ^ 1'b0 ;
  assign n5015 = n239 ^ x104 ^ x63 ;
  assign n5016 = n4132 ^ n4006 ^ n192 ;
  assign n5017 = ~n2411 & n5016 ;
  assign n5018 = n2251 & n5017 ;
  assign n5019 = n5015 & n5018 ;
  assign n5020 = n4997 ^ n2014 ^ 1'b0 ;
  assign n5021 = ( x80 & n1595 ) | ( x80 & n3272 ) | ( n1595 & n3272 ) ;
  assign n5022 = n2157 | n5021 ;
  assign n5023 = n612 | n5022 ;
  assign n5024 = n3013 ^ n264 ^ 1'b0 ;
  assign n5025 = n831 & n1102 ;
  assign n5026 = ( n179 & ~n1248 ) | ( n179 & n1346 ) | ( ~n1248 & n1346 ) ;
  assign n5027 = ( n3317 & n3435 ) | ( n3317 & ~n5026 ) | ( n3435 & ~n5026 ) ;
  assign n5028 = ~n1697 & n4381 ;
  assign n5029 = ~n5027 & n5028 ;
  assign n5030 = n293 & n3825 ;
  assign n5031 = ( n2239 & n2860 ) | ( n2239 & n3948 ) | ( n2860 & n3948 ) ;
  assign n5032 = n515 & n5031 ;
  assign n5033 = n2492 & n5032 ;
  assign n5034 = n4841 ^ n3843 ^ n2067 ;
  assign n5035 = n4508 & ~n5034 ;
  assign n5036 = ~n3841 & n5035 ;
  assign n5037 = n5036 ^ n998 ^ 1'b0 ;
  assign n5040 = n415 | n1917 ;
  assign n5041 = n5040 ^ n3229 ^ 1'b0 ;
  assign n5038 = n204 | n1308 ;
  assign n5039 = n5038 ^ n2215 ^ 1'b0 ;
  assign n5042 = n5041 ^ n5039 ^ n1702 ;
  assign n5043 = n5042 ^ n3564 ^ n3415 ;
  assign n5044 = ~n1003 & n4659 ;
  assign n5045 = n5044 ^ n612 ^ 1'b0 ;
  assign n5046 = n5045 ^ n3827 ^ 1'b0 ;
  assign n5047 = ( n1251 & n4721 ) | ( n1251 & n4837 ) | ( n4721 & n4837 ) ;
  assign n5051 = ( ~x12 & n2213 ) | ( ~x12 & n2798 ) | ( n2213 & n2798 ) ;
  assign n5048 = ( n454 & ~n2801 ) | ( n454 & n4218 ) | ( ~n2801 & n4218 ) ;
  assign n5049 = n5048 ^ n462 ^ 1'b0 ;
  assign n5050 = n2834 & n5049 ;
  assign n5052 = n5051 ^ n5050 ^ n743 ;
  assign n5053 = n4030 | n5052 ;
  assign n5054 = n3289 ^ n1144 ^ 1'b0 ;
  assign n5055 = ( ~x106 & n3519 ) | ( ~x106 & n3840 ) | ( n3519 & n3840 ) ;
  assign n5056 = n5055 ^ n3452 ^ n1330 ;
  assign n5057 = n2270 ^ n504 ^ 1'b0 ;
  assign n5058 = n1275 ^ n1117 ^ n254 ;
  assign n5059 = n5058 ^ n2199 ^ n1220 ;
  assign n5060 = ( n967 & n3650 ) | ( n967 & ~n4530 ) | ( n3650 & ~n4530 ) ;
  assign n5061 = ( n690 & n898 ) | ( n690 & ~n1601 ) | ( n898 & ~n1601 ) ;
  assign n5062 = n5061 ^ n4666 ^ n1767 ;
  assign n5063 = n3595 & ~n5062 ;
  assign n5064 = n5063 ^ n492 ^ 1'b0 ;
  assign n5065 = n2842 ^ n2352 ^ n1204 ;
  assign n5066 = n1353 | n5065 ;
  assign n5067 = n2763 ^ n1347 ^ 1'b0 ;
  assign n5068 = n3338 & n5067 ;
  assign n5069 = ( n162 & n2524 ) | ( n162 & ~n5068 ) | ( n2524 & ~n5068 ) ;
  assign n5070 = n5069 ^ n2501 ^ n1128 ;
  assign n5071 = n768 & ~n3047 ;
  assign n5072 = n5070 | n5071 ;
  assign n5073 = n5072 ^ n4860 ^ 1'b0 ;
  assign n5074 = n5073 ^ n4980 ^ n3428 ;
  assign n5075 = n1504 | n5073 ;
  assign n5076 = n3716 & ~n5075 ;
  assign n5077 = n3688 | n5076 ;
  assign n5078 = n5077 ^ n725 ^ 1'b0 ;
  assign n5079 = n1500 & n3272 ;
  assign n5080 = ( n242 & n4916 ) | ( n242 & ~n5015 ) | ( n4916 & ~n5015 ) ;
  assign n5081 = ~n524 & n3918 ;
  assign n5082 = n5081 ^ n3194 ^ 1'b0 ;
  assign n5083 = n1190 & n5082 ;
  assign n5084 = n5083 ^ n340 ^ 1'b0 ;
  assign n5085 = n2161 & ~n5084 ;
  assign n5086 = n2513 | n4691 ;
  assign n5087 = n2356 & ~n5086 ;
  assign n5088 = n5087 ^ n2963 ^ 1'b0 ;
  assign n5089 = n5088 ^ n4888 ^ x91 ;
  assign n5090 = ~n4488 & n5089 ;
  assign n5091 = n1016 & n5090 ;
  assign n5092 = ( ~n581 & n2880 ) | ( ~n581 & n4478 ) | ( n2880 & n4478 ) ;
  assign n5093 = n3227 ^ n2032 ^ n1280 ;
  assign n5094 = ~n2234 & n5093 ;
  assign n5095 = n5094 ^ n1901 ^ 1'b0 ;
  assign n5096 = ( n1285 & n3024 ) | ( n1285 & ~n5095 ) | ( n3024 & ~n5095 ) ;
  assign n5097 = ~n4101 & n5096 ;
  assign n5098 = n5097 ^ n4073 ^ 1'b0 ;
  assign n5099 = n1346 | n5098 ;
  assign n5100 = n5099 ^ n1295 ^ 1'b0 ;
  assign n5101 = n5100 ^ n2778 ^ n1910 ;
  assign n5102 = n5053 ^ n3918 ^ n265 ;
  assign n5103 = ( ~n164 & n832 ) | ( ~n164 & n4331 ) | ( n832 & n4331 ) ;
  assign n5104 = ( n2264 & n3868 ) | ( n2264 & ~n5103 ) | ( n3868 & ~n5103 ) ;
  assign n5105 = n2113 | n4841 ;
  assign n5106 = n774 & n5105 ;
  assign n5112 = x71 & n503 ;
  assign n5109 = n1553 ^ n315 ^ 1'b0 ;
  assign n5110 = n1347 & ~n5109 ;
  assign n5111 = n5110 ^ n352 ^ 1'b0 ;
  assign n5113 = n5112 ^ n5111 ^ 1'b0 ;
  assign n5114 = n457 & ~n5113 ;
  assign n5107 = n1628 ^ n1488 ^ 1'b0 ;
  assign n5108 = n2234 | n5107 ;
  assign n5115 = n5114 ^ n5108 ^ 1'b0 ;
  assign n5116 = n1919 ^ n178 ^ 1'b0 ;
  assign n5117 = ~n2728 & n3687 ;
  assign n5118 = n5116 & n5117 ;
  assign n5119 = n4596 ^ n1426 ^ 1'b0 ;
  assign n5120 = n5119 ^ n4786 ^ n2016 ;
  assign n5121 = ( n1651 & ~n2569 ) | ( n1651 & n5120 ) | ( ~n2569 & n5120 ) ;
  assign n5122 = ( n2262 & n3891 ) | ( n2262 & ~n5121 ) | ( n3891 & ~n5121 ) ;
  assign n5123 = n5122 ^ n3308 ^ n943 ;
  assign n5126 = ~n1553 & n2239 ;
  assign n5124 = n1197 & ~n2706 ;
  assign n5125 = n5124 ^ n656 ^ 1'b0 ;
  assign n5127 = n5126 ^ n5125 ^ 1'b0 ;
  assign n5128 = n5127 ^ n4855 ^ 1'b0 ;
  assign n5129 = n4500 ^ n3958 ^ n2682 ;
  assign n5130 = n239 & ~n1414 ;
  assign n5131 = n2067 & n5130 ;
  assign n5132 = n1170 & ~n5131 ;
  assign n5135 = ( x116 & ~n1052 ) | ( x116 & n4248 ) | ( ~n1052 & n4248 ) ;
  assign n5133 = n1220 ^ n1041 ^ n499 ;
  assign n5134 = n1820 & n5133 ;
  assign n5136 = n5135 ^ n5134 ^ n3061 ;
  assign n5137 = n5136 ^ n3900 ^ n3081 ;
  assign n5138 = n3798 ^ n716 ^ n540 ;
  assign n5139 = ( ~n4910 & n5137 ) | ( ~n4910 & n5138 ) | ( n5137 & n5138 ) ;
  assign n5140 = ( ~n1832 & n3309 ) | ( ~n1832 & n3436 ) | ( n3309 & n3436 ) ;
  assign n5141 = n5140 ^ n2178 ^ n1311 ;
  assign n5142 = ~n2915 & n3006 ;
  assign n5143 = n3583 ^ n513 ^ 1'b0 ;
  assign n5144 = n1620 & ~n5143 ;
  assign n5145 = n5144 ^ n1323 ^ 1'b0 ;
  assign n5146 = ~n1393 & n5145 ;
  assign n5147 = ( n4711 & ~n5142 ) | ( n4711 & n5146 ) | ( ~n5142 & n5146 ) ;
  assign n5153 = ( ~n445 & n2723 ) | ( ~n445 & n3125 ) | ( n2723 & n3125 ) ;
  assign n5148 = n3035 ^ n2057 ^ 1'b0 ;
  assign n5149 = n1348 & ~n5148 ;
  assign n5150 = n1806 ^ n1148 ^ n699 ;
  assign n5151 = n4163 ^ n3799 ^ n2236 ;
  assign n5152 = ( n5149 & n5150 ) | ( n5149 & n5151 ) | ( n5150 & n5151 ) ;
  assign n5154 = n5153 ^ n5152 ^ n708 ;
  assign n5155 = n4913 ^ n4596 ^ 1'b0 ;
  assign n5156 = n5155 ^ n515 ^ n207 ;
  assign n5157 = n5156 ^ n3404 ^ n2073 ;
  assign n5158 = n357 & ~n1693 ;
  assign n5159 = ( x64 & ~n240 ) | ( x64 & n1183 ) | ( ~n240 & n1183 ) ;
  assign n5160 = n5158 & ~n5159 ;
  assign n5161 = n5157 & n5160 ;
  assign n5162 = n935 ^ n657 ^ x27 ;
  assign n5163 = ~n424 & n5162 ;
  assign n5164 = n5163 ^ n1419 ^ 1'b0 ;
  assign n5165 = n5164 ^ n483 ^ n305 ;
  assign n5166 = ( n645 & n1351 ) | ( n645 & ~n2049 ) | ( n1351 & ~n2049 ) ;
  assign n5167 = n4292 ^ n4066 ^ n626 ;
  assign n5168 = n5166 & n5167 ;
  assign n5169 = n5168 ^ n3573 ^ 1'b0 ;
  assign n5170 = n357 & ~n2504 ;
  assign n5171 = n504 & n5170 ;
  assign n5172 = ( n1393 & ~n2010 ) | ( n1393 & n4889 ) | ( ~n2010 & n4889 ) ;
  assign n5173 = n1609 ^ n1460 ^ 1'b0 ;
  assign n5174 = n3891 & ~n5173 ;
  assign n5175 = n3485 ^ n1958 ^ n863 ;
  assign n5176 = n5175 ^ n3925 ^ n1347 ;
  assign n5177 = ( n1083 & n1380 ) | ( n1083 & ~n4049 ) | ( n1380 & ~n4049 ) ;
  assign n5178 = n1950 ^ n1638 ^ n1210 ;
  assign n5179 = n5178 ^ n643 ^ 1'b0 ;
  assign n5180 = ( ~n2239 & n5177 ) | ( ~n2239 & n5179 ) | ( n5177 & n5179 ) ;
  assign n5181 = ( ~n3904 & n3916 ) | ( ~n3904 & n4647 ) | ( n3916 & n4647 ) ;
  assign n5182 = n3188 ^ n2999 ^ n569 ;
  assign n5183 = n5182 ^ n4457 ^ 1'b0 ;
  assign n5184 = n3186 & n5183 ;
  assign n5185 = n501 & ~n1190 ;
  assign n5186 = ( n1364 & n1817 ) | ( n1364 & n5185 ) | ( n1817 & n5185 ) ;
  assign n5187 = ~n1578 & n2339 ;
  assign n5188 = n5187 ^ n618 ^ 1'b0 ;
  assign n5189 = n823 & ~n5188 ;
  assign n5190 = n3022 ^ n2815 ^ 1'b0 ;
  assign n5191 = n5189 & n5190 ;
  assign n5192 = ~n3054 & n5191 ;
  assign n5193 = ~n5186 & n5192 ;
  assign n5194 = n1109 | n1288 ;
  assign n5195 = n5194 ^ n4333 ^ 1'b0 ;
  assign n5196 = ( x7 & n5193 ) | ( x7 & n5195 ) | ( n5193 & n5195 ) ;
  assign n5197 = n5196 ^ n5062 ^ 1'b0 ;
  assign n5198 = n4559 ^ n1059 ^ x21 ;
  assign n5199 = n1944 & n2313 ;
  assign n5200 = n3701 ^ n1568 ^ 1'b0 ;
  assign n5201 = ( n5198 & n5199 ) | ( n5198 & n5200 ) | ( n5199 & n5200 ) ;
  assign n5210 = n2023 ^ n323 ^ n265 ;
  assign n5211 = n2350 | n3261 ;
  assign n5212 = n5210 & ~n5211 ;
  assign n5213 = ~n2723 & n2871 ;
  assign n5214 = n5212 & n5213 ;
  assign n5202 = n1817 ^ n958 ^ 1'b0 ;
  assign n5203 = n847 & ~n5202 ;
  assign n5204 = n5203 ^ n377 ^ 1'b0 ;
  assign n5205 = n927 | n5204 ;
  assign n5206 = n5205 ^ n3083 ^ 1'b0 ;
  assign n5207 = n5206 ^ n2243 ^ 1'b0 ;
  assign n5208 = n607 | n4052 ;
  assign n5209 = n5207 & n5208 ;
  assign n5215 = n5214 ^ n5209 ^ 1'b0 ;
  assign n5216 = n1507 ^ n542 ^ 1'b0 ;
  assign n5219 = ( n220 & ~n1017 ) | ( n220 & n1069 ) | ( ~n1017 & n1069 ) ;
  assign n5217 = n1808 ^ n883 ^ 1'b0 ;
  assign n5218 = n1833 & ~n5217 ;
  assign n5220 = n5219 ^ n5218 ^ n141 ;
  assign n5221 = ( n3318 & n5216 ) | ( n3318 & ~n5220 ) | ( n5216 & ~n5220 ) ;
  assign n5222 = n2016 ^ n1151 ^ 1'b0 ;
  assign n5227 = n1474 ^ x4 ^ 1'b0 ;
  assign n5225 = n2128 ^ n1609 ^ n1102 ;
  assign n5226 = ( ~x49 & n3058 ) | ( ~x49 & n5225 ) | ( n3058 & n5225 ) ;
  assign n5223 = n1863 | n2237 ;
  assign n5224 = n2045 & ~n5223 ;
  assign n5228 = n5227 ^ n5226 ^ n5224 ;
  assign n5229 = n5228 ^ n3673 ^ n3031 ;
  assign n5237 = x90 & ~n1239 ;
  assign n5238 = ~x35 & n5237 ;
  assign n5231 = ( n732 & n2057 ) | ( n732 & n2887 ) | ( n2057 & n2887 ) ;
  assign n5232 = ( n313 & n988 ) | ( n313 & n5231 ) | ( n988 & n5231 ) ;
  assign n5233 = ( x105 & ~n159 ) | ( x105 & n1170 ) | ( ~n159 & n1170 ) ;
  assign n5234 = n5233 ^ x15 ^ 1'b0 ;
  assign n5235 = ( n3560 & n5232 ) | ( n3560 & n5234 ) | ( n5232 & n5234 ) ;
  assign n5230 = n3817 ^ n1456 ^ 1'b0 ;
  assign n5236 = n5235 ^ n5230 ^ n3700 ;
  assign n5239 = n5238 ^ n5236 ^ n887 ;
  assign n5241 = n3023 | n4231 ;
  assign n5242 = n5241 ^ n1298 ^ 1'b0 ;
  assign n5240 = n4629 ^ n1806 ^ 1'b0 ;
  assign n5243 = n5242 ^ n5240 ^ n3829 ;
  assign n5244 = ( n1597 & n1900 ) | ( n1597 & ~n3334 ) | ( n1900 & ~n3334 ) ;
  assign n5245 = n1511 & n1977 ;
  assign n5246 = ( x105 & n3612 ) | ( x105 & n3926 ) | ( n3612 & n3926 ) ;
  assign n5247 = ( n165 & n5245 ) | ( n165 & ~n5246 ) | ( n5245 & ~n5246 ) ;
  assign n5248 = n2771 ^ n533 ^ 1'b0 ;
  assign n5249 = n1786 ^ n1506 ^ n1044 ;
  assign n5250 = n5249 ^ n3544 ^ n1826 ;
  assign n5251 = n3773 & n5250 ;
  assign n5252 = n5251 ^ n5062 ^ 1'b0 ;
  assign n5253 = ( n2959 & n5248 ) | ( n2959 & n5252 ) | ( n5248 & n5252 ) ;
  assign n5254 = n4947 ^ n2870 ^ n649 ;
  assign n5255 = n1725 | n4489 ;
  assign n5256 = n1293 & n2756 ;
  assign n5257 = n1176 ^ x89 ^ 1'b0 ;
  assign n5258 = ~n859 & n5257 ;
  assign n5259 = n4341 ^ n2288 ^ n1376 ;
  assign n5260 = ( n2590 & n5258 ) | ( n2590 & ~n5259 ) | ( n5258 & ~n5259 ) ;
  assign n5261 = ( n1093 & n1574 ) | ( n1093 & ~n2722 ) | ( n1574 & ~n2722 ) ;
  assign n5262 = ( ~x68 & n513 ) | ( ~x68 & n5261 ) | ( n513 & n5261 ) ;
  assign n5263 = n329 & ~n5262 ;
  assign n5264 = n748 & n5263 ;
  assign n5265 = n314 & n943 ;
  assign n5266 = n5265 ^ n2198 ^ 1'b0 ;
  assign n5267 = ( n1416 & n3950 ) | ( n1416 & ~n5266 ) | ( n3950 & ~n5266 ) ;
  assign n5268 = ( n2509 & ~n5264 ) | ( n2509 & n5267 ) | ( ~n5264 & n5267 ) ;
  assign n5270 = n1647 | n4679 ;
  assign n5271 = n1977 | n5270 ;
  assign n5269 = ( ~n129 & n1375 ) | ( ~n129 & n1685 ) | ( n1375 & n1685 ) ;
  assign n5272 = n5271 ^ n5269 ^ 1'b0 ;
  assign n5273 = n4465 & n5272 ;
  assign n5274 = n5261 ^ n2631 ^ 1'b0 ;
  assign n5275 = ~n3936 & n5274 ;
  assign n5277 = n3539 ^ n1779 ^ 1'b0 ;
  assign n5276 = n3774 ^ n1068 ^ 1'b0 ;
  assign n5278 = n5277 ^ n5276 ^ n5266 ;
  assign n5279 = ( n1339 & n5275 ) | ( n1339 & n5278 ) | ( n5275 & n5278 ) ;
  assign n5281 = ( x103 & ~n913 ) | ( x103 & n1959 ) | ( ~n913 & n1959 ) ;
  assign n5280 = n1641 & n1833 ;
  assign n5282 = n5281 ^ n5280 ^ 1'b0 ;
  assign n5283 = n1847 & ~n5282 ;
  assign n5284 = ~n1073 & n1679 ;
  assign n5285 = n5284 ^ n4938 ^ 1'b0 ;
  assign n5286 = n3892 ^ n2375 ^ n1481 ;
  assign n5296 = n609 | n1786 ;
  assign n5287 = n1023 ^ n620 ^ 1'b0 ;
  assign n5288 = ~n1565 & n5287 ;
  assign n5289 = n484 ^ x115 ^ 1'b0 ;
  assign n5290 = n2082 & n5289 ;
  assign n5291 = n2436 & n5290 ;
  assign n5292 = ~n5288 & n5291 ;
  assign n5293 = n5292 ^ n4770 ^ 1'b0 ;
  assign n5294 = ~n2489 & n5293 ;
  assign n5295 = ( n1671 & n3203 ) | ( n1671 & ~n5294 ) | ( n3203 & ~n5294 ) ;
  assign n5297 = n5296 ^ n5295 ^ n1059 ;
  assign n5298 = n4630 | n5297 ;
  assign n5299 = n5286 | n5298 ;
  assign n5300 = n3080 & n5080 ;
  assign n5301 = n5300 ^ n3147 ^ x19 ;
  assign n5302 = ( n805 & ~n4480 ) | ( n805 & n4878 ) | ( ~n4480 & n4878 ) ;
  assign n5303 = ( n3230 & n3305 ) | ( n3230 & n5302 ) | ( n3305 & n5302 ) ;
  assign n5304 = n5303 ^ n5175 ^ n958 ;
  assign n5305 = n5304 ^ n3028 ^ n2047 ;
  assign n5306 = n4356 | n4562 ;
  assign n5307 = ( n307 & n1599 ) | ( n307 & n2161 ) | ( n1599 & n2161 ) ;
  assign n5308 = ( n1199 & n4305 ) | ( n1199 & n5307 ) | ( n4305 & n5307 ) ;
  assign n5309 = n1558 | n5308 ;
  assign n5310 = n2272 ^ n1533 ^ 1'b0 ;
  assign n5313 = ~n199 & n857 ;
  assign n5314 = ~n907 & n4824 ;
  assign n5315 = x23 & ~n5314 ;
  assign n5316 = n5315 ^ n3364 ^ 1'b0 ;
  assign n5317 = n2479 & n4619 ;
  assign n5318 = n5317 ^ n4601 ^ 1'b0 ;
  assign n5319 = ( n5313 & ~n5316 ) | ( n5313 & n5318 ) | ( ~n5316 & n5318 ) ;
  assign n5311 = ( n187 & n2131 ) | ( n187 & n2150 ) | ( n2131 & n2150 ) ;
  assign n5312 = n1558 & ~n5311 ;
  assign n5320 = n5319 ^ n5312 ^ n1532 ;
  assign n5321 = ( n2887 & n5310 ) | ( n2887 & ~n5320 ) | ( n5310 & ~n5320 ) ;
  assign n5322 = n2149 ^ x43 ^ 1'b0 ;
  assign n5323 = n2671 & n5322 ;
  assign n5324 = ~n3987 & n5323 ;
  assign n5325 = ~n2141 & n2313 ;
  assign n5326 = n5325 ^ n305 ^ 1'b0 ;
  assign n5327 = n5324 & ~n5326 ;
  assign n5328 = ~n130 & n3404 ;
  assign n5329 = ( ~n1588 & n1664 ) | ( ~n1588 & n5328 ) | ( n1664 & n5328 ) ;
  assign n5330 = n3998 ^ n2798 ^ n1001 ;
  assign n5331 = n2055 & n3110 ;
  assign n5332 = ~n1647 & n2117 ;
  assign n5333 = n2653 | n3145 ;
  assign n5334 = ( n618 & n5332 ) | ( n618 & ~n5333 ) | ( n5332 & ~n5333 ) ;
  assign n5335 = ( n5330 & n5331 ) | ( n5330 & n5334 ) | ( n5331 & n5334 ) ;
  assign n5336 = ~n5329 & n5335 ;
  assign n5337 = ~n5327 & n5336 ;
  assign n5338 = n656 ^ n340 ^ x123 ;
  assign n5339 = n4864 & ~n5338 ;
  assign n5340 = ( n2680 & ~n4055 ) | ( n2680 & n5339 ) | ( ~n4055 & n5339 ) ;
  assign n5343 = n1677 | n2816 ;
  assign n5344 = n5343 ^ n1603 ^ 1'b0 ;
  assign n5345 = n3486 & ~n5344 ;
  assign n5341 = ( n884 & ~n4149 ) | ( n884 & n4766 ) | ( ~n4149 & n4766 ) ;
  assign n5342 = ( n1606 & n4690 ) | ( n1606 & ~n5341 ) | ( n4690 & ~n5341 ) ;
  assign n5346 = n5345 ^ n5342 ^ n454 ;
  assign n5347 = n5346 ^ n3098 ^ 1'b0 ;
  assign n5348 = ~n248 & n5347 ;
  assign n5349 = n2014 & n4770 ;
  assign n5350 = ( ~n767 & n3453 ) | ( ~n767 & n4230 ) | ( n3453 & n4230 ) ;
  assign n5351 = n5350 ^ n2199 ^ 1'b0 ;
  assign n5352 = n187 & n5351 ;
  assign n5353 = n582 ^ x79 ^ 1'b0 ;
  assign n5354 = ( n1493 & n4016 ) | ( n1493 & ~n5353 ) | ( n4016 & ~n5353 ) ;
  assign n5355 = n5354 ^ n2441 ^ 1'b0 ;
  assign n5356 = n335 & ~n5355 ;
  assign n5357 = n233 & n3338 ;
  assign n5358 = n5356 & n5357 ;
  assign n5359 = n4541 ^ n1978 ^ 1'b0 ;
  assign n5360 = n5358 & n5359 ;
  assign n5361 = n5356 ^ n1049 ^ n317 ;
  assign n5362 = ( ~n332 & n685 ) | ( ~n332 & n907 ) | ( n685 & n907 ) ;
  assign n5363 = ~n334 & n1134 ;
  assign n5364 = n5363 ^ x110 ^ 1'b0 ;
  assign n5365 = n2093 & ~n5364 ;
  assign n5366 = n5362 & n5365 ;
  assign n5367 = n2725 & ~n5366 ;
  assign n5368 = n5367 ^ x124 ^ 1'b0 ;
  assign n5369 = n2700 & ~n5368 ;
  assign n5373 = n1323 ^ n1034 ^ 1'b0 ;
  assign n5370 = n2157 | n2784 ;
  assign n5371 = n5370 ^ n1601 ^ 1'b0 ;
  assign n5372 = ( n427 & n2293 ) | ( n427 & ~n5371 ) | ( n2293 & ~n5371 ) ;
  assign n5374 = n5373 ^ n5372 ^ 1'b0 ;
  assign n5375 = n678 & ~n1809 ;
  assign n5376 = n5374 & n5375 ;
  assign n5377 = ( n765 & n2103 ) | ( n765 & ~n2226 ) | ( n2103 & ~n2226 ) ;
  assign n5378 = n351 | n2364 ;
  assign n5379 = n2089 | n5378 ;
  assign n5380 = n5379 ^ n2365 ^ n399 ;
  assign n5382 = n525 ^ n215 ^ x84 ;
  assign n5381 = n680 | n4862 ;
  assign n5383 = n5382 ^ n5381 ^ 1'b0 ;
  assign n5384 = n3357 | n3423 ;
  assign n5385 = ( n3120 & n5337 ) | ( n3120 & ~n5384 ) | ( n5337 & ~n5384 ) ;
  assign n5386 = ( n1119 & ~n2055 ) | ( n1119 & n5242 ) | ( ~n2055 & n5242 ) ;
  assign n5387 = n670 | n3023 ;
  assign n5388 = n1780 & n5387 ;
  assign n5389 = n5388 ^ n1107 ^ n418 ;
  assign n5390 = n5389 ^ n4500 ^ n3755 ;
  assign n5391 = n2253 | n2488 ;
  assign n5392 = n5391 ^ n3829 ^ 1'b0 ;
  assign n5393 = n1984 & ~n5392 ;
  assign n5394 = n3009 & n5393 ;
  assign n5395 = ~x59 & n5394 ;
  assign n5396 = n5395 ^ n4014 ^ n943 ;
  assign n5397 = n5396 ^ n1994 ^ n1020 ;
  assign n5398 = n5397 ^ n3625 ^ n1747 ;
  assign n5399 = n1332 | n3955 ;
  assign n5400 = n2598 & n5399 ;
  assign n5401 = ~n4515 & n5400 ;
  assign n5402 = n211 & n266 ;
  assign n5403 = n1424 & n5402 ;
  assign n5404 = n5403 ^ n1200 ^ 1'b0 ;
  assign n5405 = ~n2407 & n5404 ;
  assign n5407 = ~n1651 & n2050 ;
  assign n5408 = ~n4867 & n5407 ;
  assign n5406 = n2542 & n3963 ;
  assign n5409 = n5408 ^ n5406 ^ 1'b0 ;
  assign n5410 = ~n619 & n4249 ;
  assign n5411 = n5410 ^ n2560 ^ 1'b0 ;
  assign n5412 = n5411 ^ n4150 ^ 1'b0 ;
  assign n5413 = ( ~n4889 & n5409 ) | ( ~n4889 & n5412 ) | ( n5409 & n5412 ) ;
  assign n5414 = n981 | n1663 ;
  assign n5415 = n5414 ^ n4786 ^ n3352 ;
  assign n5416 = ( n1290 & n2974 ) | ( n1290 & ~n4264 ) | ( n2974 & ~n4264 ) ;
  assign n5417 = n3969 ^ n1444 ^ 1'b0 ;
  assign n5418 = n5416 | n5417 ;
  assign n5419 = n5418 ^ n3825 ^ n2653 ;
  assign n5420 = n2331 ^ n2150 ^ 1'b0 ;
  assign n5421 = ~n568 & n5420 ;
  assign n5422 = n2403 ^ n199 ^ 1'b0 ;
  assign n5423 = n5421 & n5422 ;
  assign n5424 = n5423 ^ n1057 ^ x84 ;
  assign n5425 = ( n545 & n1299 ) | ( n545 & ~n2676 ) | ( n1299 & ~n2676 ) ;
  assign n5426 = n5425 ^ n5162 ^ 1'b0 ;
  assign n5427 = ~n5424 & n5426 ;
  assign n5428 = n5419 & n5427 ;
  assign n5429 = n4096 & n5428 ;
  assign n5430 = n3835 ^ n1353 ^ 1'b0 ;
  assign n5431 = ~n1769 & n5430 ;
  assign n5432 = ( n690 & ~n2055 ) | ( n690 & n5431 ) | ( ~n2055 & n5431 ) ;
  assign n5433 = n730 | n3309 ;
  assign n5434 = n5432 | n5433 ;
  assign n5435 = n5115 & ~n5301 ;
  assign n5436 = ~n5434 & n5435 ;
  assign n5437 = n322 | n3442 ;
  assign n5438 = n5437 ^ n4461 ^ 1'b0 ;
  assign n5439 = n5438 ^ n4505 ^ 1'b0 ;
  assign n5440 = n5439 ^ n708 ^ n377 ;
  assign n5444 = ( n595 & n1137 ) | ( n595 & n2828 ) | ( n1137 & n2828 ) ;
  assign n5445 = ~n3409 & n5444 ;
  assign n5446 = ~x49 & n5445 ;
  assign n5447 = n5446 ^ x24 ^ 1'b0 ;
  assign n5441 = ~n226 & n1334 ;
  assign n5442 = n5441 ^ n1118 ^ n635 ;
  assign n5443 = n4848 & n5442 ;
  assign n5448 = n5447 ^ n5443 ^ 1'b0 ;
  assign n5449 = n3193 | n5306 ;
  assign n5452 = n2548 & n4335 ;
  assign n5450 = n3205 & n4843 ;
  assign n5451 = ~n1819 & n5450 ;
  assign n5453 = n5452 ^ n5451 ^ n199 ;
  assign n5454 = ( ~n2926 & n3451 ) | ( ~n2926 & n4701 ) | ( n3451 & n4701 ) ;
  assign n5455 = n5454 ^ n2915 ^ n2378 ;
  assign n5456 = n5455 ^ n5391 ^ n4036 ;
  assign n5461 = n4811 ^ n1706 ^ n1330 ;
  assign n5457 = ( n1076 & n1152 ) | ( n1076 & ~n1503 ) | ( n1152 & ~n1503 ) ;
  assign n5458 = n5457 ^ n3102 ^ n1823 ;
  assign n5459 = n5458 ^ n2884 ^ 1'b0 ;
  assign n5460 = n5459 ^ n2306 ^ 1'b0 ;
  assign n5462 = n5461 ^ n5460 ^ n3936 ;
  assign n5463 = n823 & ~n2247 ;
  assign n5464 = ~n2946 & n5463 ;
  assign n5465 = n3277 | n5464 ;
  assign n5466 = x28 | n5465 ;
  assign n5467 = n2599 ^ n1593 ^ 1'b0 ;
  assign n5468 = n5466 & ~n5467 ;
  assign n5469 = n5468 ^ n2710 ^ 1'b0 ;
  assign n5470 = ( ~n307 & n2109 ) | ( ~n307 & n4722 ) | ( n2109 & n4722 ) ;
  assign n5471 = n5470 ^ n4750 ^ 1'b0 ;
  assign n5472 = ( ~n159 & n787 ) | ( ~n159 & n5471 ) | ( n787 & n5471 ) ;
  assign n5473 = n1330 & n1393 ;
  assign n5474 = n5472 | n5473 ;
  assign n5475 = n2006 & ~n2688 ;
  assign n5476 = n692 ^ n293 ^ x98 ;
  assign n5477 = n1074 & n5476 ;
  assign n5478 = n5477 ^ n3202 ^ 1'b0 ;
  assign n5479 = n2413 | n5478 ;
  assign n5480 = ~n366 & n646 ;
  assign n5481 = x20 & ~n5480 ;
  assign n5482 = n5481 ^ n911 ^ 1'b0 ;
  assign n5483 = n1543 | n1943 ;
  assign n5484 = n2094 & n5483 ;
  assign n5485 = n5484 ^ n3620 ^ 1'b0 ;
  assign n5486 = n3117 ^ n2876 ^ n519 ;
  assign n5489 = n2329 ^ n844 ^ 1'b0 ;
  assign n5487 = n3379 & n4341 ;
  assign n5488 = n5288 & ~n5487 ;
  assign n5490 = n5489 ^ n5488 ^ 1'b0 ;
  assign n5491 = n338 | n919 ;
  assign n5492 = n5491 ^ n2226 ^ 1'b0 ;
  assign n5493 = n3220 ^ n2887 ^ 1'b0 ;
  assign n5494 = n5492 | n5493 ;
  assign n5495 = n3248 ^ n880 ^ 1'b0 ;
  assign n5496 = ~n4721 & n5495 ;
  assign n5497 = ( ~n1129 & n5494 ) | ( ~n1129 & n5496 ) | ( n5494 & n5496 ) ;
  assign n5498 = n3698 & ~n5497 ;
  assign n5499 = n5490 & n5498 ;
  assign n5500 = n4308 | n5499 ;
  assign n5501 = n3625 & ~n5500 ;
  assign n5502 = n5501 ^ n4624 ^ n1583 ;
  assign n5506 = ( n500 & n1106 ) | ( n500 & n1388 ) | ( n1106 & n1388 ) ;
  assign n5507 = ( ~n1048 & n1323 ) | ( ~n1048 & n5506 ) | ( n1323 & n5506 ) ;
  assign n5508 = ( n1475 & ~n2842 ) | ( n1475 & n5507 ) | ( ~n2842 & n5507 ) ;
  assign n5509 = n5508 ^ n4546 ^ 1'b0 ;
  assign n5503 = n783 | n3360 ;
  assign n5504 = n5503 ^ n190 ^ 1'b0 ;
  assign n5505 = n1729 & ~n5504 ;
  assign n5510 = n5509 ^ n5505 ^ 1'b0 ;
  assign n5512 = ( n1143 & n1243 ) | ( n1143 & n1322 ) | ( n1243 & n1322 ) ;
  assign n5511 = n171 | n1371 ;
  assign n5513 = n5512 ^ n5511 ^ 1'b0 ;
  assign n5514 = ( n343 & n1644 ) | ( n343 & ~n3137 ) | ( n1644 & ~n3137 ) ;
  assign n5515 = ( n4428 & n5513 ) | ( n4428 & ~n5514 ) | ( n5513 & ~n5514 ) ;
  assign n5522 = ( x90 & n194 ) | ( x90 & n3696 ) | ( n194 & n3696 ) ;
  assign n5523 = n5522 ^ n732 ^ x31 ;
  assign n5517 = n909 & ~n1109 ;
  assign n5518 = n5517 ^ n1501 ^ 1'b0 ;
  assign n5519 = n1879 & n5518 ;
  assign n5520 = ( n1589 & ~n1788 ) | ( n1589 & n5519 ) | ( ~n1788 & n5519 ) ;
  assign n5516 = ( n4648 & n4672 ) | ( n4648 & n4815 ) | ( n4672 & n4815 ) ;
  assign n5521 = n5520 ^ n5516 ^ n3447 ;
  assign n5524 = n5523 ^ n5521 ^ 1'b0 ;
  assign n5525 = ( x54 & ~n2624 ) | ( x54 & n2633 ) | ( ~n2624 & n2633 ) ;
  assign n5526 = ( n397 & ~n2683 ) | ( n397 & n5525 ) | ( ~n2683 & n5525 ) ;
  assign n5527 = ( n1477 & ~n2919 ) | ( n1477 & n5526 ) | ( ~n2919 & n5526 ) ;
  assign n5529 = n1595 ^ n605 ^ 1'b0 ;
  assign n5530 = ( n616 & n2699 ) | ( n616 & ~n5529 ) | ( n2699 & ~n5529 ) ;
  assign n5528 = n2383 & n3349 ;
  assign n5531 = n5530 ^ n5528 ^ 1'b0 ;
  assign n5532 = n5531 ^ n3305 ^ n1574 ;
  assign n5533 = ( n2272 & n2957 ) | ( n2272 & ~n4838 ) | ( n2957 & ~n4838 ) ;
  assign n5534 = n1504 ^ x43 ^ 1'b0 ;
  assign n5535 = ( n415 & n5533 ) | ( n415 & n5534 ) | ( n5533 & n5534 ) ;
  assign n5536 = n1690 | n5535 ;
  assign n5537 = n5536 ^ n3485 ^ 1'b0 ;
  assign n5538 = n2346 | n5537 ;
  assign n5539 = ( n935 & n2424 ) | ( n935 & n5538 ) | ( n2424 & n5538 ) ;
  assign n5540 = ( ~n2378 & n2638 ) | ( ~n2378 & n3033 ) | ( n2638 & n3033 ) ;
  assign n5541 = n1481 | n1926 ;
  assign n5542 = n5338 & ~n5541 ;
  assign n5543 = n3581 & ~n5542 ;
  assign n5544 = n3475 ^ n654 ^ 1'b0 ;
  assign n5545 = n4102 & ~n5544 ;
  assign n5546 = n5545 ^ n2217 ^ n1192 ;
  assign n5557 = n509 & ~n1407 ;
  assign n5558 = n5557 ^ n2349 ^ 1'b0 ;
  assign n5552 = n1623 ^ n1592 ^ n903 ;
  assign n5553 = ( n523 & n1496 ) | ( n523 & n5552 ) | ( n1496 & n5552 ) ;
  assign n5554 = n5553 ^ n3943 ^ 1'b0 ;
  assign n5555 = n335 & ~n5554 ;
  assign n5556 = n5555 ^ n620 ^ 1'b0 ;
  assign n5547 = n1572 | n4566 ;
  assign n5548 = n5547 ^ n238 ^ 1'b0 ;
  assign n5549 = n5548 ^ n2076 ^ n980 ;
  assign n5550 = n5549 ^ n4381 ^ 1'b0 ;
  assign n5551 = ( n1714 & ~n2365 ) | ( n1714 & n5550 ) | ( ~n2365 & n5550 ) ;
  assign n5559 = n5558 ^ n5556 ^ n5551 ;
  assign n5560 = n5559 ^ n4943 ^ n326 ;
  assign n5561 = ( n2262 & ~n5121 ) | ( n2262 & n5461 ) | ( ~n5121 & n5461 ) ;
  assign n5562 = ( n674 & n1450 ) | ( n674 & ~n1972 ) | ( n1450 & ~n1972 ) ;
  assign n5563 = n4620 ^ n4425 ^ n3724 ;
  assign n5564 = ~n199 & n4592 ;
  assign n5565 = ( ~n2912 & n5421 ) | ( ~n2912 & n5564 ) | ( n5421 & n5564 ) ;
  assign n5566 = ( ~n5562 & n5563 ) | ( ~n5562 & n5565 ) | ( n5563 & n5565 ) ;
  assign n5567 = n4849 ^ n390 ^ 1'b0 ;
  assign n5568 = ~n3001 & n5567 ;
  assign n5569 = ~n203 & n405 ;
  assign n5570 = n3595 | n5569 ;
  assign n5571 = n2819 & n5570 ;
  assign n5572 = n2692 & n5571 ;
  assign n5573 = n5568 | n5572 ;
  assign n5575 = n486 ^ n445 ^ 1'b0 ;
  assign n5574 = n1340 & ~n2069 ;
  assign n5576 = n5575 ^ n5574 ^ 1'b0 ;
  assign n5577 = ( ~n3825 & n5158 ) | ( ~n3825 & n5180 ) | ( n5158 & n5180 ) ;
  assign n5578 = n4412 ^ n1709 ^ n699 ;
  assign n5579 = ( n2272 & ~n3338 ) | ( n2272 & n5578 ) | ( ~n3338 & n5578 ) ;
  assign n5580 = n1821 | n5579 ;
  assign n5581 = n5580 ^ n1307 ^ 1'b0 ;
  assign n5582 = ( n308 & n2097 ) | ( n308 & ~n2163 ) | ( n2097 & ~n2163 ) ;
  assign n5586 = n2405 & n4115 ;
  assign n5587 = n5586 ^ n2079 ^ 1'b0 ;
  assign n5588 = x54 & ~n5587 ;
  assign n5589 = n499 & n5588 ;
  assign n5583 = n1896 ^ n1045 ^ n474 ;
  assign n5584 = n5583 ^ n2265 ^ 1'b0 ;
  assign n5585 = n3724 | n5584 ;
  assign n5590 = n5589 ^ n5585 ^ n3209 ;
  assign n5591 = n4575 | n5562 ;
  assign n5592 = n5591 ^ n2020 ^ 1'b0 ;
  assign n5593 = n5592 ^ n2405 ^ 1'b0 ;
  assign n5594 = ~n2339 & n5593 ;
  assign n5595 = ( n1063 & n2317 ) | ( n1063 & n5105 ) | ( n2317 & n5105 ) ;
  assign n5596 = n2329 & ~n5492 ;
  assign n5597 = n478 & n5596 ;
  assign n5598 = n239 | n3436 ;
  assign n5599 = n5179 & n5598 ;
  assign n5600 = n5597 & n5599 ;
  assign n5606 = n1503 & n5250 ;
  assign n5607 = n5606 ^ n1717 ^ n325 ;
  assign n5602 = n762 ^ n374 ^ x84 ;
  assign n5601 = n2237 & n3718 ;
  assign n5603 = n5602 ^ n5601 ^ 1'b0 ;
  assign n5604 = ~n1606 & n5603 ;
  assign n5605 = ( n844 & n5174 ) | ( n844 & ~n5604 ) | ( n5174 & ~n5604 ) ;
  assign n5608 = n5607 ^ n5605 ^ 1'b0 ;
  assign n5609 = n4840 | n5608 ;
  assign n5611 = n3701 | n5198 ;
  assign n5610 = ( n420 & ~n2219 ) | ( n420 & n3118 ) | ( ~n2219 & n3118 ) ;
  assign n5612 = n5611 ^ n5610 ^ n2579 ;
  assign n5618 = ~n795 & n4619 ;
  assign n5619 = n2983 & n5618 ;
  assign n5615 = x78 & n1819 ;
  assign n5616 = ~n531 & n5615 ;
  assign n5613 = n4072 ^ n3268 ^ n1146 ;
  assign n5614 = n3704 | n5613 ;
  assign n5617 = n5616 ^ n5614 ^ 1'b0 ;
  assign n5620 = n5619 ^ n5617 ^ n2973 ;
  assign n5621 = ~n686 & n2272 ;
  assign n5622 = n5621 ^ n2059 ^ 1'b0 ;
  assign n5623 = n677 & n1320 ;
  assign n5624 = ( ~n412 & n5622 ) | ( ~n412 & n5623 ) | ( n5622 & n5623 ) ;
  assign n5625 = n984 & n1618 ;
  assign n5626 = ~n1614 & n2884 ;
  assign n5627 = n5626 ^ n4642 ^ 1'b0 ;
  assign n5628 = n5627 ^ n3091 ^ n604 ;
  assign n5630 = ( n1036 & ~n2230 ) | ( n1036 & n2633 ) | ( ~n2230 & n2633 ) ;
  assign n5629 = n3334 & ~n4123 ;
  assign n5631 = n5630 ^ n5629 ^ 1'b0 ;
  assign n5632 = ~n5628 & n5631 ;
  assign n5633 = n3105 & n5632 ;
  assign n5634 = n4059 ^ n3207 ^ n1366 ;
  assign n5636 = n4158 ^ n1944 ^ n176 ;
  assign n5635 = ~n287 & n1270 ;
  assign n5637 = n5636 ^ n5635 ^ 1'b0 ;
  assign n5638 = n2682 ^ n2295 ^ 1'b0 ;
  assign n5639 = n5637 & ~n5638 ;
  assign n5640 = n1166 ^ n650 ^ 1'b0 ;
  assign n5641 = n4736 & n5640 ;
  assign n5642 = ( n3330 & n4075 ) | ( n3330 & n5641 ) | ( n4075 & n5641 ) ;
  assign n5643 = n1111 & n5642 ;
  assign n5646 = x124 & ~n810 ;
  assign n5647 = n160 & n5646 ;
  assign n5648 = ( n673 & ~n4257 ) | ( n673 & n5647 ) | ( ~n4257 & n5647 ) ;
  assign n5649 = n5648 ^ n3442 ^ 1'b0 ;
  assign n5650 = n3251 ^ n1411 ^ 1'b0 ;
  assign n5651 = ~n5021 & n5650 ;
  assign n5652 = n5651 ^ n2324 ^ n235 ;
  assign n5653 = n5649 & n5652 ;
  assign n5644 = n2734 ^ n2666 ^ n1388 ;
  assign n5645 = n5644 ^ n5036 ^ n5027 ;
  assign n5654 = n5653 ^ n5645 ^ n4107 ;
  assign n5655 = n1829 | n3441 ;
  assign n5656 = n786 & n830 ;
  assign n5658 = n5140 ^ n2730 ^ 1'b0 ;
  assign n5659 = n5658 ^ x1 ^ 1'b0 ;
  assign n5657 = n4175 | n5601 ;
  assign n5660 = n5659 ^ n5657 ^ 1'b0 ;
  assign n5661 = ( n2218 & n2390 ) | ( n2218 & ~n3096 ) | ( n2390 & ~n3096 ) ;
  assign n5662 = n5332 & n5661 ;
  assign n5663 = n5662 ^ n4148 ^ 1'b0 ;
  assign n5664 = n4055 ^ n1266 ^ 1'b0 ;
  assign n5665 = ~n422 & n5664 ;
  assign n5666 = n4648 ^ n575 ^ 1'b0 ;
  assign n5667 = n1331 & ~n5666 ;
  assign n5668 = ( n351 & ~n1018 ) | ( n351 & n3696 ) | ( ~n1018 & n3696 ) ;
  assign n5669 = n5668 ^ n5616 ^ n1148 ;
  assign n5670 = n5669 ^ n4977 ^ 1'b0 ;
  assign n5671 = ( n3443 & ~n4260 ) | ( n3443 & n5670 ) | ( ~n4260 & n5670 ) ;
  assign n5672 = n5159 ^ n3448 ^ n3146 ;
  assign n5677 = n5512 ^ n1468 ^ n1107 ;
  assign n5673 = n3761 ^ n328 ^ n160 ;
  assign n5674 = n4500 ^ n1999 ^ n1737 ;
  assign n5675 = n1843 & n5674 ;
  assign n5676 = ( n3159 & n5673 ) | ( n3159 & n5675 ) | ( n5673 & n5675 ) ;
  assign n5678 = n5677 ^ n5676 ^ 1'b0 ;
  assign n5679 = n5120 & ~n5678 ;
  assign n5680 = n4426 | n5679 ;
  assign n5681 = n5672 & n5680 ;
  assign n5682 = n5510 ^ n2441 ^ 1'b0 ;
  assign n5683 = n4729 | n5682 ;
  assign n5684 = n5081 ^ n2364 ^ 1'b0 ;
  assign n5685 = n1111 & n2394 ;
  assign n5686 = ( x27 & ~n364 ) | ( x27 & n5685 ) | ( ~n364 & n5685 ) ;
  assign n5687 = n5686 ^ n3006 ^ 1'b0 ;
  assign n5688 = n3134 & ~n5264 ;
  assign n5689 = ~n783 & n5688 ;
  assign n5699 = ( n282 & ~n512 ) | ( n282 & n1248 ) | ( ~n512 & n1248 ) ;
  assign n5700 = n451 & ~n5699 ;
  assign n5701 = n4214 & n5700 ;
  assign n5696 = x123 | n4112 ;
  assign n5692 = n2403 ^ n1483 ^ 1'b0 ;
  assign n5693 = x112 & n328 ;
  assign n5694 = ( n3012 & n5692 ) | ( n3012 & ~n5693 ) | ( n5692 & ~n5693 ) ;
  assign n5695 = ( n1666 & n2482 ) | ( n1666 & ~n5694 ) | ( n2482 & ~n5694 ) ;
  assign n5697 = n5696 ^ n5695 ^ 1'b0 ;
  assign n5698 = n3051 & n5697 ;
  assign n5690 = n3558 & ~n5242 ;
  assign n5691 = n199 & n5690 ;
  assign n5702 = n5701 ^ n5698 ^ n5691 ;
  assign n5703 = n5195 ^ n4108 ^ n2895 ;
  assign n5704 = n3134 ^ n2472 ^ n1338 ;
  assign n5705 = ( n2130 & n2251 ) | ( n2130 & ~n5552 ) | ( n2251 & ~n5552 ) ;
  assign n5706 = n941 ^ n238 ^ x39 ;
  assign n5707 = n2833 ^ n1445 ^ 1'b0 ;
  assign n5708 = x101 & ~n5707 ;
  assign n5709 = ( n5539 & ~n5706 ) | ( n5539 & n5708 ) | ( ~n5706 & n5708 ) ;
  assign n5710 = n367 & n1711 ;
  assign n5711 = n5710 ^ n4849 ^ n3164 ;
  assign n5712 = n2220 ^ n472 ^ 1'b0 ;
  assign n5713 = n5712 ^ n3312 ^ 1'b0 ;
  assign n5714 = n2451 & n5713 ;
  assign n5715 = n5714 ^ n264 ^ 1'b0 ;
  assign n5716 = ( n568 & n819 ) | ( n568 & n4570 ) | ( n819 & n4570 ) ;
  assign n5717 = n4947 ^ n357 ^ 1'b0 ;
  assign n5718 = n1886 | n5717 ;
  assign n5720 = ( n605 & n1152 ) | ( n605 & n1531 ) | ( n1152 & n1531 ) ;
  assign n5721 = ( n2243 & ~n5529 ) | ( n2243 & n5720 ) | ( ~n5529 & n5720 ) ;
  assign n5722 = n5721 ^ n1575 ^ 1'b0 ;
  assign n5719 = x79 & n4680 ;
  assign n5723 = n5722 ^ n5719 ^ 1'b0 ;
  assign n5724 = ~n1200 & n5723 ;
  assign n5727 = n199 | n773 ;
  assign n5728 = n2788 & ~n5727 ;
  assign n5725 = n2838 ^ n1111 ^ n926 ;
  assign n5726 = n5725 ^ n3147 ^ n2420 ;
  assign n5729 = n5728 ^ n5726 ^ 1'b0 ;
  assign n5730 = n5729 ^ n1341 ^ 1'b0 ;
  assign n5731 = n5730 ^ n3161 ^ n220 ;
  assign n5732 = n5731 ^ n5139 ^ n778 ;
  assign n5733 = n5732 ^ n4584 ^ n192 ;
  assign n5734 = n1306 & n3014 ;
  assign n5735 = ~n4614 & n5734 ;
  assign n5736 = ( n1370 & n1381 ) | ( n1370 & n3625 ) | ( n1381 & n3625 ) ;
  assign n5737 = n5735 | n5736 ;
  assign n5738 = ( n1724 & n1860 ) | ( n1724 & n2324 ) | ( n1860 & n2324 ) ;
  assign n5739 = n5738 ^ n4390 ^ n1644 ;
  assign n5740 = n477 ^ n268 ^ n248 ;
  assign n5741 = ( n1681 & n2530 ) | ( n1681 & ~n5740 ) | ( n2530 & ~n5740 ) ;
  assign n5742 = n5741 ^ n2040 ^ 1'b0 ;
  assign n5743 = n5739 | n5742 ;
  assign n5744 = n3235 & ~n4519 ;
  assign n5745 = n4903 ^ n2557 ^ n427 ;
  assign n5748 = n3144 ^ n1310 ^ 1'b0 ;
  assign n5746 = n3096 ^ n2770 ^ n2556 ;
  assign n5747 = n5746 ^ x61 ^ 1'b0 ;
  assign n5749 = n5748 ^ n5747 ^ n3035 ;
  assign n5750 = n5749 ^ n1153 ^ 1'b0 ;
  assign n5751 = n4145 ^ n1645 ^ x2 ;
  assign n5752 = ( x15 & ~n2413 ) | ( x15 & n5751 ) | ( ~n2413 & n5751 ) ;
  assign n5753 = n3825 ^ n3169 ^ 1'b0 ;
  assign n5754 = n4150 ^ n1832 ^ 1'b0 ;
  assign n5755 = ~n133 & n4293 ;
  assign n5756 = ~x29 & n5755 ;
  assign n5757 = n2378 | n5756 ;
  assign n5758 = n5757 ^ n4560 ^ 1'b0 ;
  assign n5759 = n5754 & n5758 ;
  assign n5760 = ( n3930 & ~n5753 ) | ( n3930 & n5759 ) | ( ~n5753 & n5759 ) ;
  assign n5761 = n4157 ^ n3675 ^ 1'b0 ;
  assign n5762 = ( ~n643 & n2149 ) | ( ~n643 & n2544 ) | ( n2149 & n2544 ) ;
  assign n5763 = ( n2445 & ~n2940 ) | ( n2445 & n5762 ) | ( ~n2940 & n5762 ) ;
  assign n5764 = n5245 ^ n136 ^ 1'b0 ;
  assign n5765 = n3409 ^ n3135 ^ 1'b0 ;
  assign n5766 = ( n973 & n5764 ) | ( n973 & n5765 ) | ( n5764 & n5765 ) ;
  assign n5767 = ~n1343 & n4623 ;
  assign n5768 = n2713 | n5497 ;
  assign n5769 = n5768 ^ x78 ^ 1'b0 ;
  assign n5770 = n5769 ^ n3039 ^ 1'b0 ;
  assign n5779 = n4114 ^ n896 ^ 1'b0 ;
  assign n5780 = ( n2227 & n3198 ) | ( n2227 & ~n5779 ) | ( n3198 & ~n5779 ) ;
  assign n5781 = n5780 ^ n298 ^ 1'b0 ;
  assign n5771 = ~n1946 & n2272 ;
  assign n5772 = n1959 & n5771 ;
  assign n5773 = n5772 ^ n469 ^ n257 ;
  assign n5774 = ( x84 & n1544 ) | ( x84 & n5773 ) | ( n1544 & n5773 ) ;
  assign n5775 = n5774 ^ n3924 ^ n162 ;
  assign n5776 = ( ~n420 & n3459 ) | ( ~n420 & n3461 ) | ( n3459 & n3461 ) ;
  assign n5777 = n5776 ^ n2455 ^ 1'b0 ;
  assign n5778 = n5775 & ~n5777 ;
  assign n5782 = n5781 ^ n5778 ^ 1'b0 ;
  assign n5783 = n260 & n3887 ;
  assign n5784 = n3541 & n5783 ;
  assign n5785 = n5784 ^ n2032 ^ 1'b0 ;
  assign n5786 = n5661 ^ n5174 ^ n3825 ;
  assign n5787 = n5512 ^ n1040 ^ 1'b0 ;
  assign n5788 = n2079 | n2750 ;
  assign n5791 = n792 | n1062 ;
  assign n5790 = n2745 ^ x52 ^ 1'b0 ;
  assign n5792 = n5791 ^ n5790 ^ n3193 ;
  assign n5793 = n1284 & n5792 ;
  assign n5789 = n5556 ^ n4094 ^ n3604 ;
  assign n5794 = n5793 ^ n5789 ^ 1'b0 ;
  assign n5795 = n4022 ^ n2109 ^ 1'b0 ;
  assign n5796 = n2207 | n5795 ;
  assign n5797 = n4030 & n5796 ;
  assign n5798 = n5797 ^ n4307 ^ n2426 ;
  assign n5799 = n1151 ^ n1062 ^ n268 ;
  assign n5800 = ( n1557 & ~n3902 ) | ( n1557 & n5799 ) | ( ~n3902 & n5799 ) ;
  assign n5801 = n3255 ^ n1012 ^ 1'b0 ;
  assign n5802 = n838 & ~n5801 ;
  assign n5803 = ~n3019 & n5802 ;
  assign n5804 = ~n5800 & n5803 ;
  assign n5805 = n2284 ^ n1565 ^ 1'b0 ;
  assign n5806 = ( n1915 & n4457 ) | ( n1915 & n5805 ) | ( n4457 & n5805 ) ;
  assign n5807 = n1052 ^ n270 ^ 1'b0 ;
  assign n5808 = n5807 ^ n1833 ^ 1'b0 ;
  assign n5809 = n5806 & n5808 ;
  assign n5810 = n406 & ~n2682 ;
  assign n5811 = x126 & n580 ;
  assign n5812 = n1767 & ~n5811 ;
  assign n5813 = n5812 ^ n1053 ^ 1'b0 ;
  assign n5814 = ( n254 & n1815 ) | ( n254 & ~n1819 ) | ( n1815 & ~n1819 ) ;
  assign n5815 = n3016 | n3443 ;
  assign n5816 = ( n1283 & n5814 ) | ( n1283 & n5815 ) | ( n5814 & n5815 ) ;
  assign n5817 = n2381 & n5816 ;
  assign n5818 = n2402 ^ n513 ^ 1'b0 ;
  assign n5819 = n5818 ^ n3471 ^ 1'b0 ;
  assign n5820 = ~n5817 & n5819 ;
  assign n5821 = ( ~n1174 & n2631 ) | ( ~n1174 & n5820 ) | ( n2631 & n5820 ) ;
  assign n5822 = ( x19 & n744 ) | ( x19 & ~n2016 ) | ( n744 & ~n2016 ) ;
  assign n5823 = n1436 | n1729 ;
  assign n5824 = n220 | n5823 ;
  assign n5825 = n905 & n4474 ;
  assign n5826 = ~n5824 & n5825 ;
  assign n5827 = ( n910 & n1147 ) | ( n910 & ~n5653 ) | ( n1147 & ~n5653 ) ;
  assign n5828 = ( n5822 & ~n5826 ) | ( n5822 & n5827 ) | ( ~n5826 & n5827 ) ;
  assign n5829 = ( n1777 & n4986 ) | ( n1777 & n5358 ) | ( n4986 & n5358 ) ;
  assign n5830 = n4846 ^ n4496 ^ 1'b0 ;
  assign n5831 = n1550 & n5830 ;
  assign n5832 = ~n2623 & n5016 ;
  assign n5833 = n1917 & n5832 ;
  assign n5834 = ( ~n1183 & n3895 ) | ( ~n1183 & n5833 ) | ( n3895 & n5833 ) ;
  assign n5835 = n3301 ^ n186 ^ 1'b0 ;
  assign n5836 = ~n5015 & n5835 ;
  assign n5837 = n2422 ^ n1725 ^ 1'b0 ;
  assign n5838 = n5837 ^ n1106 ^ n476 ;
  assign n5839 = ~n5268 & n5781 ;
  assign n5840 = n374 & ~n5816 ;
  assign n5841 = ~n4478 & n5840 ;
  assign n5851 = n1070 | n1841 ;
  assign n5852 = ~n3085 & n3615 ;
  assign n5853 = n5852 ^ n3230 ^ 1'b0 ;
  assign n5854 = ( ~n2501 & n2808 ) | ( ~n2501 & n4726 ) | ( n2808 & n4726 ) ;
  assign n5855 = n954 & n1387 ;
  assign n5856 = n5855 ^ n2830 ^ 1'b0 ;
  assign n5857 = ( n324 & n5854 ) | ( n324 & n5856 ) | ( n5854 & n5856 ) ;
  assign n5858 = n5853 & ~n5857 ;
  assign n5859 = ~n5851 & n5858 ;
  assign n5842 = n1225 ^ n1183 ^ 1'b0 ;
  assign n5843 = n380 | n5842 ;
  assign n5844 = n5843 ^ n2801 ^ n562 ;
  assign n5845 = n3080 ^ n2642 ^ 1'b0 ;
  assign n5846 = x18 & ~n5845 ;
  assign n5847 = ( n1139 & ~n5844 ) | ( n1139 & n5846 ) | ( ~n5844 & n5846 ) ;
  assign n5848 = ~n3674 & n5847 ;
  assign n5849 = ~n1547 & n5848 ;
  assign n5850 = n821 & ~n5849 ;
  assign n5860 = n5859 ^ n5850 ^ 1'b0 ;
  assign n5861 = n3080 ^ n2749 ^ 1'b0 ;
  assign n5862 = n4911 ^ n4875 ^ n2144 ;
  assign n5863 = n5862 ^ n2643 ^ n659 ;
  assign n5869 = ( n468 & n2526 ) | ( n468 & ~n4691 ) | ( n2526 & ~n4691 ) ;
  assign n5870 = n5869 ^ n2023 ^ n1217 ;
  assign n5871 = ( n1287 & n2678 ) | ( n1287 & ~n5870 ) | ( n2678 & ~n5870 ) ;
  assign n5864 = n1287 ^ n357 ^ 1'b0 ;
  assign n5865 = n5864 ^ n765 ^ 1'b0 ;
  assign n5866 = n5249 ^ n2067 ^ 1'b0 ;
  assign n5867 = n5865 | n5866 ;
  assign n5868 = n5867 ^ n1944 ^ 1'b0 ;
  assign n5872 = n5871 ^ n5868 ^ 1'b0 ;
  assign n5873 = n5863 & ~n5872 ;
  assign n5874 = x115 & n4045 ;
  assign n5875 = n2855 & n5874 ;
  assign n5876 = n3415 & ~n5036 ;
  assign n5877 = n2583 & n5876 ;
  assign n5878 = ~n4005 & n4336 ;
  assign n5879 = n829 & n5878 ;
  assign n5880 = n5879 ^ n510 ^ 1'b0 ;
  assign n5881 = n5860 & n5880 ;
  assign n5885 = n5814 ^ n4100 ^ n3485 ;
  assign n5882 = ~n2066 & n2726 ;
  assign n5883 = n5882 ^ n245 ^ 1'b0 ;
  assign n5884 = n4183 & n5883 ;
  assign n5886 = n5885 ^ n5884 ^ 1'b0 ;
  assign n5887 = ( ~n1232 & n4895 ) | ( ~n1232 & n5886 ) | ( n4895 & n5886 ) ;
  assign n5888 = n734 & n3959 ;
  assign n5889 = n297 & n5888 ;
  assign n5890 = n5526 ^ n1007 ^ n816 ;
  assign n5897 = ~n3344 & n5630 ;
  assign n5898 = ~n927 & n5897 ;
  assign n5899 = n2573 ^ n1240 ^ 1'b0 ;
  assign n5900 = n5898 | n5899 ;
  assign n5891 = n1455 ^ n983 ^ 1'b0 ;
  assign n5892 = ( n2214 & ~n2356 ) | ( n2214 & n5891 ) | ( ~n2356 & n5891 ) ;
  assign n5893 = n4824 ^ n2892 ^ 1'b0 ;
  assign n5894 = n5892 & ~n5893 ;
  assign n5895 = n5212 ^ n4197 ^ 1'b0 ;
  assign n5896 = n5894 & n5895 ;
  assign n5901 = n5900 ^ n5896 ^ x2 ;
  assign n5902 = n5901 ^ n3762 ^ 1'b0 ;
  assign n5903 = n881 & ~n3278 ;
  assign n5904 = n2736 & n5903 ;
  assign n5905 = n3585 ^ n194 ^ 1'b0 ;
  assign n5906 = ~n601 & n1237 ;
  assign n5907 = n1334 & ~n3191 ;
  assign n5908 = n5906 | n5907 ;
  assign n5909 = n5905 & ~n5908 ;
  assign n5910 = n5904 | n5909 ;
  assign n5911 = n1970 ^ n871 ^ 1'b0 ;
  assign n5912 = n1916 & n2336 ;
  assign n5913 = ( n5802 & n5911 ) | ( n5802 & n5912 ) | ( n5911 & n5912 ) ;
  assign n5914 = n1480 | n1496 ;
  assign n5915 = n1992 & n2137 ;
  assign n5916 = n5915 ^ n3903 ^ n2969 ;
  assign n5917 = ( n1550 & n5914 ) | ( n1550 & ~n5916 ) | ( n5914 & ~n5916 ) ;
  assign n5918 = n395 & n1514 ;
  assign n5919 = ~n5523 & n5918 ;
  assign n5920 = n5919 ^ n2759 ^ 1'b0 ;
  assign n5921 = n3889 ^ n1014 ^ n260 ;
  assign n5922 = n5921 ^ n225 ^ 1'b0 ;
  assign n5923 = n5920 | n5922 ;
  assign n5924 = n213 | n2160 ;
  assign n5925 = n5924 ^ n525 ^ 1'b0 ;
  assign n5926 = n575 & n5925 ;
  assign n5927 = n5926 ^ n4516 ^ 1'b0 ;
  assign n5928 = n246 & ~n2743 ;
  assign n5935 = ~n631 & n2797 ;
  assign n5930 = ~n619 & n815 ;
  assign n5931 = n5930 ^ n3678 ^ 1'b0 ;
  assign n5932 = ~n709 & n5931 ;
  assign n5933 = n5932 ^ n4024 ^ 1'b0 ;
  assign n5934 = n4426 | n5933 ;
  assign n5936 = n5935 ^ n5934 ^ n2815 ;
  assign n5929 = n1550 & n3806 ;
  assign n5937 = n5936 ^ n5929 ^ 1'b0 ;
  assign n5938 = n734 ^ n390 ^ 1'b0 ;
  assign n5939 = n1972 & ~n5938 ;
  assign n5940 = n2494 ^ n1450 ^ 1'b0 ;
  assign n5941 = n5939 & n5940 ;
  assign n5942 = n5941 ^ n999 ^ 1'b0 ;
  assign n5943 = n2205 & ~n4264 ;
  assign n5944 = ~n4697 & n5943 ;
  assign n5946 = ( ~n1083 & n2608 ) | ( ~n1083 & n3820 ) | ( n2608 & n3820 ) ;
  assign n5947 = n1530 ^ n177 ^ 1'b0 ;
  assign n5948 = n5947 ^ n3236 ^ n2077 ;
  assign n5949 = n5948 ^ n5473 ^ n2725 ;
  assign n5950 = n5949 ^ n1752 ^ 1'b0 ;
  assign n5951 = n5946 & ~n5950 ;
  assign n5945 = n2232 & ~n4793 ;
  assign n5952 = n5951 ^ n5945 ^ 1'b0 ;
  assign n5954 = n1552 | n3736 ;
  assign n5955 = n3615 | n5954 ;
  assign n5953 = n3047 & ~n4616 ;
  assign n5956 = n5955 ^ n5953 ^ 1'b0 ;
  assign n5957 = n5956 ^ n2014 ^ n686 ;
  assign n5958 = n2440 ^ n1336 ^ 1'b0 ;
  assign n5959 = n2395 | n5958 ;
  assign n5960 = n1613 & ~n2658 ;
  assign n5961 = n5960 ^ n1407 ^ 1'b0 ;
  assign n5962 = ( n5136 & n5959 ) | ( n5136 & ~n5961 ) | ( n5959 & ~n5961 ) ;
  assign n5963 = n4088 & ~n5962 ;
  assign n5964 = ~n948 & n2211 ;
  assign n5965 = n5964 ^ n2743 ^ 1'b0 ;
  assign n5966 = ( x107 & n757 ) | ( x107 & ~n5965 ) | ( n757 & ~n5965 ) ;
  assign n5967 = n5966 ^ n5478 ^ 1'b0 ;
  assign n5968 = n3016 ^ n2467 ^ n910 ;
  assign n5969 = n4271 ^ n1761 ^ n1095 ;
  assign n5970 = n2296 & n5969 ;
  assign n5971 = n5970 ^ n5065 ^ n686 ;
  assign n5972 = ~n5968 & n5971 ;
  assign n5973 = ~n5612 & n5972 ;
  assign n5974 = n3937 ^ n1468 ^ 1'b0 ;
  assign n5975 = ( n937 & n2149 ) | ( n937 & n2623 ) | ( n2149 & n2623 ) ;
  assign n5976 = ( n235 & n1879 ) | ( n235 & ~n2009 ) | ( n1879 & ~n2009 ) ;
  assign n5977 = ( ~n525 & n1859 ) | ( ~n525 & n5976 ) | ( n1859 & n5976 ) ;
  assign n5978 = ( n5974 & n5975 ) | ( n5974 & ~n5977 ) | ( n5975 & ~n5977 ) ;
  assign n5979 = ( n3597 & n4510 ) | ( n3597 & n5978 ) | ( n4510 & n5978 ) ;
  assign n5980 = n4864 & n5144 ;
  assign n5981 = n5980 ^ n3862 ^ n2694 ;
  assign n5982 = ~n1371 & n5529 ;
  assign n5983 = n5982 ^ n2468 ^ 1'b0 ;
  assign n5984 = n3101 | n5983 ;
  assign n5985 = n5984 ^ n1426 ^ 1'b0 ;
  assign n5986 = n1154 & ~n5985 ;
  assign n5987 = ~n5981 & n5986 ;
  assign n5988 = n3312 ^ n1841 ^ 1'b0 ;
  assign n5989 = ( n2426 & n3593 ) | ( n2426 & n5988 ) | ( n3593 & n5988 ) ;
  assign n5990 = n897 & n5457 ;
  assign n5991 = ( n3852 & ~n4163 ) | ( n3852 & n5990 ) | ( ~n4163 & n5990 ) ;
  assign n5992 = n2010 | n5373 ;
  assign n5993 = n5992 ^ n2691 ^ 1'b0 ;
  assign n5994 = ( n1761 & n2038 ) | ( n1761 & ~n5993 ) | ( n2038 & ~n5993 ) ;
  assign n5995 = ( n1774 & n2653 ) | ( n1774 & ~n5994 ) | ( n2653 & ~n5994 ) ;
  assign n5996 = n4260 ^ n2174 ^ 1'b0 ;
  assign n6000 = n1308 | n2623 ;
  assign n6001 = n6000 ^ n1703 ^ 1'b0 ;
  assign n5997 = n5569 ^ n1475 ^ 1'b0 ;
  assign n5998 = n1588 | n5997 ;
  assign n5999 = n728 | n5998 ;
  assign n6002 = n6001 ^ n5999 ^ 1'b0 ;
  assign n6003 = ( ~n3444 & n4541 ) | ( ~n3444 & n6002 ) | ( n4541 & n6002 ) ;
  assign n6005 = n2421 ^ n678 ^ x4 ;
  assign n6006 = n6005 ^ n5258 ^ n1790 ;
  assign n6004 = n4070 ^ n2397 ^ n1674 ;
  assign n6007 = n6006 ^ n6004 ^ n3797 ;
  assign n6008 = n2029 ^ n1472 ^ n699 ;
  assign n6009 = ( n1514 & ~n2950 ) | ( n1514 & n6008 ) | ( ~n2950 & n6008 ) ;
  assign n6010 = ( n4554 & n5460 ) | ( n4554 & n6009 ) | ( n5460 & n6009 ) ;
  assign n6011 = ( n1065 & n2246 ) | ( n1065 & ~n2786 ) | ( n2246 & ~n2786 ) ;
  assign n6013 = ~n2243 & n3070 ;
  assign n6012 = n2413 & n3784 ;
  assign n6014 = n6013 ^ n6012 ^ 1'b0 ;
  assign n6015 = n6014 ^ n4659 ^ n3021 ;
  assign n6016 = n4839 ^ n2110 ^ n1006 ;
  assign n6017 = n1002 ^ n892 ^ 1'b0 ;
  assign n6018 = ( ~n198 & n3562 ) | ( ~n198 & n3784 ) | ( n3562 & n3784 ) ;
  assign n6019 = n5693 ^ n148 ^ 1'b0 ;
  assign n6020 = ~n6018 & n6019 ;
  assign n6021 = n6017 & n6020 ;
  assign n6022 = ( ~n238 & n378 ) | ( ~n238 & n6021 ) | ( n378 & n6021 ) ;
  assign n6023 = n6016 & n6022 ;
  assign n6024 = n6023 ^ n2506 ^ 1'b0 ;
  assign n6025 = ( n5487 & n6015 ) | ( n5487 & ~n6024 ) | ( n6015 & ~n6024 ) ;
  assign n6026 = n6025 ^ n2929 ^ n1845 ;
  assign n6027 = ~n2293 & n3413 ;
  assign n6028 = n6027 ^ n3896 ^ 1'b0 ;
  assign n6029 = ( n4221 & n4541 ) | ( n4221 & ~n6028 ) | ( n4541 & ~n6028 ) ;
  assign n6030 = ( n3299 & ~n3383 ) | ( n3299 & n6029 ) | ( ~n3383 & n6029 ) ;
  assign n6031 = ~n1139 & n4868 ;
  assign n6032 = n1003 | n5981 ;
  assign n6033 = n4740 ^ n4598 ^ 1'b0 ;
  assign n6034 = n2464 & n6033 ;
  assign n6035 = n2337 & n6034 ;
  assign n6036 = n1945 ^ n1344 ^ 1'b0 ;
  assign n6037 = n2109 ^ n1141 ^ 1'b0 ;
  assign n6038 = n1399 & n6037 ;
  assign n6039 = n6038 ^ n2921 ^ n2843 ;
  assign n6040 = ~n2545 & n3623 ;
  assign n6041 = n6040 ^ n3475 ^ 1'b0 ;
  assign n6042 = n1818 & n6041 ;
  assign n6043 = ( n1981 & n3109 ) | ( n1981 & ~n6042 ) | ( n3109 & ~n6042 ) ;
  assign n6044 = ( ~n6036 & n6039 ) | ( ~n6036 & n6043 ) | ( n6039 & n6043 ) ;
  assign n6045 = ( n444 & ~n1657 ) | ( n444 & n2677 ) | ( ~n1657 & n2677 ) ;
  assign n6046 = n5837 & n6045 ;
  assign n6047 = ( n5385 & ~n5509 ) | ( n5385 & n6046 ) | ( ~n5509 & n6046 ) ;
  assign n6048 = n4421 ^ n2708 ^ n2695 ;
  assign n6049 = n6048 ^ n6030 ^ n1945 ;
  assign n6050 = ~n1439 & n1833 ;
  assign n6051 = ( x109 & ~n5566 ) | ( x109 & n6050 ) | ( ~n5566 & n6050 ) ;
  assign n6052 = n1144 & ~n3840 ;
  assign n6053 = ( ~n1782 & n3891 ) | ( ~n1782 & n4115 ) | ( n3891 & n4115 ) ;
  assign n6054 = n6039 | n6053 ;
  assign n6055 = n854 & ~n6054 ;
  assign n6056 = ( n1126 & ~n2301 ) | ( n1126 & n6055 ) | ( ~n2301 & n6055 ) ;
  assign n6057 = n3006 ^ n884 ^ 1'b0 ;
  assign n6058 = ~n3835 & n6057 ;
  assign n6059 = n148 | n2016 ;
  assign n6060 = x40 & ~n2130 ;
  assign n6061 = n1261 | n3024 ;
  assign n6062 = n6060 & ~n6061 ;
  assign n6063 = n6059 & ~n6062 ;
  assign n6064 = n6063 ^ n4588 ^ 1'b0 ;
  assign n6065 = n2559 ^ n559 ^ 1'b0 ;
  assign n6066 = ~n2954 & n6065 ;
  assign n6067 = ( n1128 & n1538 ) | ( n1128 & n1757 ) | ( n1538 & n1757 ) ;
  assign n6068 = ( n386 & ~n1376 ) | ( n386 & n6067 ) | ( ~n1376 & n6067 ) ;
  assign n6069 = n6059 ^ n360 ^ 1'b0 ;
  assign n6070 = n2131 & ~n3495 ;
  assign n6071 = ( n1073 & n1395 ) | ( n1073 & n1529 ) | ( n1395 & n1529 ) ;
  assign n6072 = ( ~n2440 & n6070 ) | ( ~n2440 & n6071 ) | ( n6070 & n6071 ) ;
  assign n6073 = n4598 & n6072 ;
  assign n6074 = n3562 | n6073 ;
  assign n6075 = n6069 & ~n6074 ;
  assign n6076 = n943 ^ x38 ^ 1'b0 ;
  assign n6077 = n550 | n6076 ;
  assign n6078 = n3586 & n6077 ;
  assign n6079 = n4479 ^ n4393 ^ 1'b0 ;
  assign n6080 = ( ~n1608 & n6078 ) | ( ~n1608 & n6079 ) | ( n6078 & n6079 ) ;
  assign n6081 = ( n1636 & n4177 ) | ( n1636 & n5469 ) | ( n4177 & n5469 ) ;
  assign n6083 = ~n1797 & n2415 ;
  assign n6084 = n6083 ^ n2967 ^ x45 ;
  assign n6082 = n3292 & n4755 ;
  assign n6085 = n6084 ^ n6082 ^ 1'b0 ;
  assign n6086 = n5724 & ~n6085 ;
  assign n6087 = n2105 & ~n3134 ;
  assign n6088 = n673 | n6087 ;
  assign n6089 = n6088 ^ n5820 ^ 1'b0 ;
  assign n6090 = n1920 & n6089 ;
  assign n6094 = ( n1369 & n3969 ) | ( n1369 & ~n5227 ) | ( n3969 & ~n5227 ) ;
  assign n6091 = n1475 | n5011 ;
  assign n6092 = n6091 ^ n2239 ^ n905 ;
  assign n6093 = ~n1578 & n6092 ;
  assign n6095 = n6094 ^ n6093 ^ n1137 ;
  assign n6096 = n3976 & ~n4524 ;
  assign n6097 = n6095 & n6096 ;
  assign n6098 = n1349 ^ n1251 ^ n1225 ;
  assign n6099 = n145 | n6098 ;
  assign n6100 = n3588 & n5507 ;
  assign n6101 = n725 & n6100 ;
  assign n6102 = n6101 ^ n3521 ^ 1'b0 ;
  assign n6103 = n1530 & n2553 ;
  assign n6104 = n6103 ^ n4222 ^ n3441 ;
  assign n6105 = n6104 ^ n4902 ^ n4185 ;
  assign n6106 = n2992 & n6105 ;
  assign n6107 = n6102 & ~n6106 ;
  assign n6108 = n6107 ^ n4927 ^ 1'b0 ;
  assign n6109 = n6108 ^ n3341 ^ 1'b0 ;
  assign n6110 = ~n2184 & n6109 ;
  assign n6111 = n6110 ^ n5606 ^ n2744 ;
  assign n6114 = n5961 ^ n4075 ^ 1'b0 ;
  assign n6115 = n4293 & n6114 ;
  assign n6112 = ~n2565 & n2801 ;
  assign n6113 = ~n3836 & n6112 ;
  assign n6116 = n6115 ^ n6113 ^ 1'b0 ;
  assign n6117 = ( ~n617 & n1804 ) | ( ~n617 & n2308 ) | ( n1804 & n2308 ) ;
  assign n6118 = ~n1572 & n6117 ;
  assign n6119 = ~n1996 & n6118 ;
  assign n6120 = n5846 ^ n5199 ^ 1'b0 ;
  assign n6121 = n2384 & n6120 ;
  assign n6122 = ( ~n1176 & n2668 ) | ( ~n1176 & n4675 ) | ( n2668 & n4675 ) ;
  assign n6123 = n5189 & n6094 ;
  assign n6124 = n6123 ^ n2662 ^ n677 ;
  assign n6125 = n5969 ^ n3236 ^ 1'b0 ;
  assign n6126 = ( ~x20 & n4660 ) | ( ~x20 & n6125 ) | ( n4660 & n6125 ) ;
  assign n6127 = n4180 ^ n4122 ^ n1772 ;
  assign n6128 = n3797 ^ n3571 ^ n1412 ;
  assign n6129 = n6128 ^ n3184 ^ 1'b0 ;
  assign n6130 = n6127 & n6129 ;
  assign n6131 = n2344 & n2509 ;
  assign n6132 = n5228 ^ n4253 ^ 1'b0 ;
  assign n6133 = ~n5647 & n6132 ;
  assign n6134 = n6133 ^ n4657 ^ n3058 ;
  assign n6137 = n624 & n3937 ;
  assign n6135 = n2973 | n3893 ;
  assign n6136 = n790 & ~n6135 ;
  assign n6138 = n6137 ^ n6136 ^ n1635 ;
  assign n6144 = n409 ^ n174 ^ 1'b0 ;
  assign n6145 = n3016 & ~n6144 ;
  assign n6146 = n6145 ^ n1588 ^ 1'b0 ;
  assign n6147 = n1891 & ~n6146 ;
  assign n6148 = n6147 ^ n3325 ^ 1'b0 ;
  assign n6149 = n3509 & n6148 ;
  assign n6139 = n1261 ^ x15 ^ 1'b0 ;
  assign n6140 = n2694 ^ n910 ^ n840 ;
  assign n6141 = n6140 ^ n656 ^ 1'b0 ;
  assign n6142 = ~n6139 & n6141 ;
  assign n6143 = ~n5034 & n6142 ;
  assign n6150 = n6149 ^ n6143 ^ 1'b0 ;
  assign n6153 = ( ~n391 & n1096 ) | ( ~n391 & n3160 ) | ( n1096 & n3160 ) ;
  assign n6151 = n1340 ^ n302 ^ n233 ;
  assign n6152 = n6151 ^ n2326 ^ n1704 ;
  assign n6154 = n6153 ^ n6152 ^ n5767 ;
  assign n6155 = ~x24 & n3967 ;
  assign n6156 = n3964 & n6155 ;
  assign n6157 = n6156 ^ n5399 ^ 1'b0 ;
  assign n6158 = n590 | n6157 ;
  assign n6159 = n544 | n1427 ;
  assign n6160 = n6159 ^ n1511 ^ 1'b0 ;
  assign n6161 = n2809 & ~n6160 ;
  assign n6162 = n6161 ^ n5225 ^ 1'b0 ;
  assign n6163 = ~n958 & n1629 ;
  assign n6164 = n6163 ^ n2067 ^ 1'b0 ;
  assign n6165 = n3903 ^ n2981 ^ n887 ;
  assign n6166 = ( n4358 & n6164 ) | ( n4358 & ~n6165 ) | ( n6164 & ~n6165 ) ;
  assign n6167 = n1580 & ~n4247 ;
  assign n6168 = ~n273 & n6167 ;
  assign n6169 = n6168 ^ n4805 ^ 1'b0 ;
  assign n6170 = n4665 ^ n753 ^ 1'b0 ;
  assign n6171 = ( ~n131 & n3129 ) | ( ~n131 & n6170 ) | ( n3129 & n6170 ) ;
  assign n6172 = n486 & ~n4660 ;
  assign n6173 = n1164 & n4311 ;
  assign n6174 = n6173 ^ n4253 ^ 1'b0 ;
  assign n6175 = n6174 ^ n3180 ^ 1'b0 ;
  assign n6176 = n1421 ^ n346 ^ x7 ;
  assign n6177 = n6176 ^ n4501 ^ n1439 ;
  assign n6178 = n2661 & n6177 ;
  assign n6179 = n6175 & n6178 ;
  assign n6180 = n2598 & n3328 ;
  assign n6181 = n6180 ^ n1880 ^ 1'b0 ;
  assign n6182 = ( n2429 & n4429 ) | ( n2429 & ~n6181 ) | ( n4429 & ~n6181 ) ;
  assign n6183 = ( n752 & n849 ) | ( n752 & n1700 ) | ( n849 & n1700 ) ;
  assign n6184 = n6183 ^ n2962 ^ 1'b0 ;
  assign n6185 = ~n4765 & n6184 ;
  assign n6190 = n3648 ^ n505 ^ n217 ;
  assign n6188 = n5865 ^ n504 ^ 1'b0 ;
  assign n6189 = ~n1638 & n6188 ;
  assign n6191 = n6190 ^ n6189 ^ n3163 ;
  assign n6192 = n4342 & ~n6191 ;
  assign n6193 = n6192 ^ n1729 ^ 1'b0 ;
  assign n6186 = n615 & n2876 ;
  assign n6187 = n6186 ^ n4841 ^ 1'b0 ;
  assign n6194 = n6193 ^ n6187 ^ 1'b0 ;
  assign n6197 = n1268 | n2198 ;
  assign n6198 = n1297 & ~n6197 ;
  assign n6199 = ~n1992 & n3551 ;
  assign n6200 = n6198 & n6199 ;
  assign n6201 = n4801 | n6200 ;
  assign n6202 = n2175 | n6201 ;
  assign n6195 = n2103 ^ n978 ^ n577 ;
  assign n6196 = n5598 & n6195 ;
  assign n6203 = n6202 ^ n6196 ^ 1'b0 ;
  assign n6204 = n1112 ^ n410 ^ 1'b0 ;
  assign n6205 = n5110 & ~n6204 ;
  assign n6206 = n6205 ^ n4968 ^ 1'b0 ;
  assign n6207 = ( x2 & x114 ) | ( x2 & n2452 ) | ( x114 & n2452 ) ;
  assign n6208 = n6207 ^ n2096 ^ n231 ;
  assign n6209 = ~n1927 & n2830 ;
  assign n6210 = ~n6208 & n6209 ;
  assign n6212 = x107 & n1523 ;
  assign n6213 = n6212 ^ n149 ^ 1'b0 ;
  assign n6214 = ~n4215 & n6213 ;
  assign n6211 = n5762 | n5776 ;
  assign n6215 = n6214 ^ n6211 ^ 1'b0 ;
  assign n6216 = ( ~n186 & n6210 ) | ( ~n186 & n6215 ) | ( n6210 & n6215 ) ;
  assign n6217 = n2555 ^ n381 ^ 1'b0 ;
  assign n6218 = ~n2857 & n6217 ;
  assign n6219 = ~n786 & n2699 ;
  assign n6220 = ( ~n576 & n859 ) | ( ~n576 & n1922 ) | ( n859 & n1922 ) ;
  assign n6221 = n1169 ^ n994 ^ 1'b0 ;
  assign n6222 = n6221 ^ n3408 ^ 1'b0 ;
  assign n6223 = n6220 & ~n6222 ;
  assign n6224 = ( n6218 & ~n6219 ) | ( n6218 & n6223 ) | ( ~n6219 & n6223 ) ;
  assign n6225 = ~n6043 & n6219 ;
  assign n6226 = ~n145 & n6225 ;
  assign n6227 = ( n2763 & ~n4542 ) | ( n2763 & n6226 ) | ( ~n4542 & n6226 ) ;
  assign n6228 = n6227 ^ n974 ^ n582 ;
  assign n6229 = n348 & ~n2688 ;
  assign n6230 = n6229 ^ n2105 ^ 1'b0 ;
  assign n6231 = n2185 | n6230 ;
  assign n6232 = n6231 ^ n3255 ^ 1'b0 ;
  assign n6239 = n2140 & ~n5512 ;
  assign n6240 = ( n2511 & ~n4723 ) | ( n2511 & n6239 ) | ( ~n4723 & n6239 ) ;
  assign n6241 = n3097 & n6240 ;
  assign n6233 = n1528 & n3733 ;
  assign n6234 = n2515 | n4458 ;
  assign n6235 = n5277 | n6234 ;
  assign n6236 = ( ~n970 & n1193 ) | ( ~n970 & n6235 ) | ( n1193 & n6235 ) ;
  assign n6237 = ( n4392 & n6226 ) | ( n4392 & n6236 ) | ( n6226 & n6236 ) ;
  assign n6238 = ( ~n5138 & n6233 ) | ( ~n5138 & n6237 ) | ( n6233 & n6237 ) ;
  assign n6242 = n6241 ^ n6238 ^ 1'b0 ;
  assign n6243 = ~n6232 & n6242 ;
  assign n6245 = n1066 & ~n3885 ;
  assign n6246 = n6245 ^ n2432 ^ 1'b0 ;
  assign n6247 = n2749 & ~n6246 ;
  assign n6248 = ( n190 & n2422 ) | ( n190 & n4329 ) | ( n2422 & n4329 ) ;
  assign n6249 = n6248 ^ n943 ^ 1'b0 ;
  assign n6250 = n6247 | n6249 ;
  assign n6244 = n5918 ^ n1691 ^ 1'b0 ;
  assign n6251 = n6250 ^ n6244 ^ 1'b0 ;
  assign n6252 = n4245 & n6251 ;
  assign n6253 = n6183 ^ x51 ^ 1'b0 ;
  assign n6254 = n6253 ^ n1208 ^ 1'b0 ;
  assign n6255 = n2644 & n6254 ;
  assign n6256 = n4939 | n6255 ;
  assign n6257 = n632 & n3877 ;
  assign n6258 = n4964 | n6257 ;
  assign n6259 = n6258 ^ n3920 ^ 1'b0 ;
  assign n6261 = n2264 ^ n372 ^ 1'b0 ;
  assign n6260 = n2994 ^ n2394 ^ n2098 ;
  assign n6262 = n6261 ^ n6260 ^ n542 ;
  assign n6263 = n481 | n6262 ;
  assign n6264 = n277 & ~n6263 ;
  assign n6265 = ( n490 & n676 ) | ( n490 & n1633 ) | ( n676 & n1633 ) ;
  assign n6266 = n6265 ^ n2983 ^ 1'b0 ;
  assign n6267 = n1119 & ~n6266 ;
  assign n6268 = n6267 ^ n4694 ^ 1'b0 ;
  assign n6269 = n3935 ^ n319 ^ 1'b0 ;
  assign n6270 = ~n2500 & n6269 ;
  assign n6271 = n6270 ^ n2159 ^ n1344 ;
  assign n6272 = n3156 & ~n6271 ;
  assign n6273 = n6268 & n6272 ;
  assign n6274 = n6273 ^ n5523 ^ n4055 ;
  assign n6275 = ~n828 & n5568 ;
  assign n6276 = n3378 ^ n545 ^ n388 ;
  assign n6277 = n6276 ^ n4568 ^ n1643 ;
  assign n6278 = ( n322 & n4357 ) | ( n322 & ~n6277 ) | ( n4357 & ~n6277 ) ;
  assign n6279 = n6278 ^ n2426 ^ 1'b0 ;
  assign n6280 = ~n1014 & n6279 ;
  assign n6281 = ( n480 & ~n1957 ) | ( n480 & n3400 ) | ( ~n1957 & n3400 ) ;
  assign n6282 = ( ~n2492 & n2604 ) | ( ~n2492 & n3586 ) | ( n2604 & n3586 ) ;
  assign n6283 = n1648 ^ n447 ^ 1'b0 ;
  assign n6284 = n6283 ^ n3323 ^ 1'b0 ;
  assign n6285 = n6282 & ~n6284 ;
  assign n6286 = n6285 ^ n892 ^ 1'b0 ;
  assign n6287 = ( n454 & ~n6281 ) | ( n454 & n6286 ) | ( ~n6281 & n6286 ) ;
  assign n6288 = n2229 ^ n1609 ^ 1'b0 ;
  assign n6289 = ~n3330 & n3836 ;
  assign n6301 = n4006 ^ n2890 ^ n1575 ;
  assign n6300 = n505 | n1246 ;
  assign n6295 = ( n500 & n724 ) | ( n500 & n1090 ) | ( n724 & n1090 ) ;
  assign n6296 = n2628 ^ n1697 ^ 1'b0 ;
  assign n6297 = n2805 | n6296 ;
  assign n6298 = n6295 | n6297 ;
  assign n6299 = n2455 | n6298 ;
  assign n6302 = n6301 ^ n6300 ^ n6299 ;
  assign n6303 = n6302 ^ n4493 ^ n4394 ;
  assign n6291 = n5108 ^ n3514 ^ n282 ;
  assign n6292 = n5178 & ~n6291 ;
  assign n6293 = n6292 ^ n3796 ^ 1'b0 ;
  assign n6290 = n4250 ^ n2086 ^ n1227 ;
  assign n6294 = n6293 ^ n6290 ^ n3698 ;
  assign n6304 = n6303 ^ n6294 ^ n4670 ;
  assign n6305 = n3450 ^ n2136 ^ 1'b0 ;
  assign n6306 = n4841 ^ n185 ^ 1'b0 ;
  assign n6307 = n1145 & n6306 ;
  assign n6308 = ( n2126 & ~n3651 ) | ( n2126 & n6307 ) | ( ~n3651 & n6307 ) ;
  assign n6309 = n3162 ^ n2403 ^ 1'b0 ;
  assign n6310 = n6308 & ~n6309 ;
  assign n6311 = ( ~n1989 & n6305 ) | ( ~n1989 & n6310 ) | ( n6305 & n6310 ) ;
  assign n6312 = n5150 ^ n1124 ^ x3 ;
  assign n6313 = n2785 | n5826 ;
  assign n6314 = n6312 & ~n6313 ;
  assign n6315 = n6314 ^ n3634 ^ 1'b0 ;
  assign n6316 = n4070 ^ n3471 ^ 1'b0 ;
  assign n6318 = n2427 & n3218 ;
  assign n6319 = ~n4511 & n6318 ;
  assign n6317 = n1873 & ~n2680 ;
  assign n6320 = n6319 ^ n6317 ^ n4329 ;
  assign n6321 = n6316 & ~n6320 ;
  assign n6322 = n5397 & n6321 ;
  assign n6323 = ~n1758 & n2346 ;
  assign n6324 = n5549 ^ n2232 ^ x3 ;
  assign n6325 = n6324 ^ n3990 ^ 1'b0 ;
  assign n6326 = n1052 ^ n459 ^ 1'b0 ;
  assign n6329 = n4010 ^ n1248 ^ 1'b0 ;
  assign n6330 = ~n1734 & n6329 ;
  assign n6327 = ( x107 & n1404 ) | ( x107 & ~n2688 ) | ( n1404 & ~n2688 ) ;
  assign n6328 = ( ~n1471 & n2341 ) | ( ~n1471 & n6327 ) | ( n2341 & n6327 ) ;
  assign n6331 = n6330 ^ n6328 ^ n1143 ;
  assign n6332 = ( n4004 & ~n6326 ) | ( n4004 & n6331 ) | ( ~n6326 & n6331 ) ;
  assign n6333 = n6332 ^ n3948 ^ 1'b0 ;
  assign n6334 = n6325 & n6333 ;
  assign n6335 = n5602 ^ n3072 ^ 1'b0 ;
  assign n6336 = ( n3358 & ~n4949 ) | ( n3358 & n6335 ) | ( ~n4949 & n6335 ) ;
  assign n6337 = n6336 ^ n5233 ^ n988 ;
  assign n6338 = ( ~n3641 & n4498 ) | ( ~n3641 & n6175 ) | ( n4498 & n6175 ) ;
  assign n6339 = n5083 ^ n1507 ^ n854 ;
  assign n6346 = n427 & n892 ;
  assign n6347 = n807 & n6346 ;
  assign n6348 = ( n253 & n768 ) | ( n253 & ~n6347 ) | ( n768 & ~n6347 ) ;
  assign n6349 = n6348 ^ n5095 ^ n171 ;
  assign n6340 = x68 & ~n3457 ;
  assign n6341 = n2659 & n6340 ;
  assign n6342 = n6341 ^ n3627 ^ 1'b0 ;
  assign n6343 = n601 & n6342 ;
  assign n6344 = n392 | n1447 ;
  assign n6345 = n6343 & n6344 ;
  assign n6350 = n6349 ^ n6345 ^ 1'b0 ;
  assign n6359 = n3019 ^ n2736 ^ n771 ;
  assign n6351 = n3412 ^ n1927 ^ 1'b0 ;
  assign n6352 = n2027 & ~n6351 ;
  assign n6353 = n6352 ^ n3723 ^ 1'b0 ;
  assign n6354 = n2964 | n3540 ;
  assign n6355 = n6354 ^ n2020 ^ 1'b0 ;
  assign n6356 = ~n3987 & n6355 ;
  assign n6357 = n6356 ^ n4279 ^ 1'b0 ;
  assign n6358 = n6353 | n6357 ;
  assign n6360 = n6359 ^ n6358 ^ n130 ;
  assign n6361 = n1784 ^ n616 ^ x127 ;
  assign n6362 = n575 & ~n1253 ;
  assign n6363 = n1759 & n6362 ;
  assign n6364 = ( n3452 & n5774 ) | ( n3452 & ~n6363 ) | ( n5774 & ~n6363 ) ;
  assign n6365 = n561 & n3726 ;
  assign n6366 = ~x55 & n6365 ;
  assign n6367 = n962 & n1530 ;
  assign n6368 = n6367 ^ x70 ^ 1'b0 ;
  assign n6369 = ( n2826 & n3757 ) | ( n2826 & ~n6368 ) | ( n3757 & ~n6368 ) ;
  assign n6370 = n6369 ^ n2989 ^ n253 ;
  assign n6371 = n2105 ^ n633 ^ n223 ;
  assign n6372 = ( ~n2152 & n2562 ) | ( ~n2152 & n6371 ) | ( n2562 & n6371 ) ;
  assign n6373 = n6372 ^ n3982 ^ n3087 ;
  assign n6374 = n6373 ^ n2580 ^ 1'b0 ;
  assign n6375 = x37 & n6374 ;
  assign n6385 = n5122 ^ n3716 ^ 1'b0 ;
  assign n6377 = ( n1190 & n3366 ) | ( n1190 & ~n3378 ) | ( n3366 & ~n3378 ) ;
  assign n6378 = ( n2193 & ~n3302 ) | ( n2193 & n6377 ) | ( ~n3302 & n6377 ) ;
  assign n6376 = x59 & ~n1500 ;
  assign n6379 = n6378 ^ n6376 ^ n4766 ;
  assign n6380 = n6379 ^ n3150 ^ 1'b0 ;
  assign n6381 = n1789 ^ n929 ^ 1'b0 ;
  assign n6382 = n6381 ^ n5585 ^ n1070 ;
  assign n6383 = ( n5905 & ~n6380 ) | ( n5905 & n6382 ) | ( ~n6380 & n6382 ) ;
  assign n6384 = n6383 ^ n2701 ^ 1'b0 ;
  assign n6386 = n6385 ^ n6384 ^ n4127 ;
  assign n6387 = n209 | n4295 ;
  assign n6388 = n6387 ^ n2369 ^ 1'b0 ;
  assign n6389 = n3009 | n6388 ;
  assign n6390 = n3177 & n5452 ;
  assign n6391 = ~x41 & n4465 ;
  assign n6392 = ( n1691 & n2259 ) | ( n1691 & ~n4923 ) | ( n2259 & ~n4923 ) ;
  assign n6393 = n6392 ^ n3516 ^ x12 ;
  assign n6394 = n6393 ^ n6338 ^ n2388 ;
  assign n6395 = n6182 ^ n4642 ^ n215 ;
  assign n6396 = ( n990 & n2549 ) | ( n990 & n3118 ) | ( n2549 & n3118 ) ;
  assign n6397 = ( x44 & n2798 ) | ( x44 & ~n4414 ) | ( n2798 & ~n4414 ) ;
  assign n6414 = ( n1681 & n2194 ) | ( n1681 & ~n6397 ) | ( n2194 & ~n6397 ) ;
  assign n6415 = n6414 ^ n2256 ^ 1'b0 ;
  assign n6413 = ~n2462 & n3328 ;
  assign n6398 = n286 ^ n164 ^ 1'b0 ;
  assign n6399 = n6398 ^ n1572 ^ n960 ;
  assign n6400 = n461 & ~n6399 ;
  assign n6401 = ~n6397 & n6400 ;
  assign n6404 = ( n169 & n2822 ) | ( n169 & n3639 ) | ( n2822 & n3639 ) ;
  assign n6402 = ~n906 & n4074 ;
  assign n6403 = n6402 ^ n162 ^ 1'b0 ;
  assign n6405 = n6404 ^ n6403 ^ 1'b0 ;
  assign n6406 = ~n3312 & n6405 ;
  assign n6407 = ( n1021 & n6401 ) | ( n1021 & ~n6406 ) | ( n6401 & ~n6406 ) ;
  assign n6408 = n6067 ^ n2171 ^ 1'b0 ;
  assign n6409 = n1451 | n6408 ;
  assign n6410 = n6409 ^ n4844 ^ 1'b0 ;
  assign n6411 = ~n6407 & n6410 ;
  assign n6412 = n6411 ^ n2310 ^ n2131 ;
  assign n6416 = n6415 ^ n6413 ^ n6412 ;
  assign n6417 = n3316 ^ n2260 ^ 1'b0 ;
  assign n6418 = n259 | n3043 ;
  assign n6419 = n6418 ^ n3936 ^ 1'b0 ;
  assign n6420 = n5243 & ~n6419 ;
  assign n6421 = ( n1304 & n1338 ) | ( n1304 & n1465 ) | ( n1338 & n1465 ) ;
  assign n6424 = n2699 ^ n1255 ^ n1163 ;
  assign n6422 = ~n1308 & n4560 ;
  assign n6423 = ~n1496 & n6422 ;
  assign n6425 = n6424 ^ n6423 ^ n1879 ;
  assign n6428 = x55 & n3766 ;
  assign n6429 = n6428 ^ n3964 ^ 1'b0 ;
  assign n6426 = n1912 | n4304 ;
  assign n6427 = n4780 & ~n6426 ;
  assign n6430 = n6429 ^ n6427 ^ 1'b0 ;
  assign n6431 = ( ~n6421 & n6425 ) | ( ~n6421 & n6430 ) | ( n6425 & n6430 ) ;
  assign n6434 = n4969 ^ n1106 ^ n367 ;
  assign n6432 = n1778 ^ n1248 ^ 1'b0 ;
  assign n6433 = ~n424 & n6432 ;
  assign n6435 = n6434 ^ n6433 ^ 1'b0 ;
  assign n6436 = n6435 ^ n2130 ^ 1'b0 ;
  assign n6437 = n2227 ^ n1085 ^ 1'b0 ;
  assign n6438 = n5548 ^ n1691 ^ 1'b0 ;
  assign n6439 = n1411 ^ n1221 ^ n885 ;
  assign n6440 = n5975 ^ n678 ^ 1'b0 ;
  assign n6441 = n133 | n6440 ;
  assign n6442 = ( n3490 & ~n6439 ) | ( n3490 & n6441 ) | ( ~n6439 & n6441 ) ;
  assign n6443 = n6442 ^ n3804 ^ n2951 ;
  assign n6444 = ( n1621 & n2030 ) | ( n1621 & ~n6443 ) | ( n2030 & ~n6443 ) ;
  assign n6445 = ( n6437 & ~n6438 ) | ( n6437 & n6444 ) | ( ~n6438 & n6444 ) ;
  assign n6447 = n934 ^ x38 ^ 1'b0 ;
  assign n6446 = ( x31 & n4312 ) | ( x31 & ~n5736 ) | ( n4312 & ~n5736 ) ;
  assign n6448 = n6447 ^ n6446 ^ 1'b0 ;
  assign n6449 = n2134 ^ n683 ^ 1'b0 ;
  assign n6450 = n1246 & n6449 ;
  assign n6451 = n6397 & n6450 ;
  assign n6452 = n6451 ^ n684 ^ 1'b0 ;
  assign n6453 = n6452 ^ n5789 ^ n5711 ;
  assign n6454 = n5792 ^ n618 ^ n268 ;
  assign n6455 = n6454 ^ n5977 ^ n1041 ;
  assign n6456 = n257 | n981 ;
  assign n6457 = n6455 & ~n6456 ;
  assign n6458 = n6457 ^ n4116 ^ 1'b0 ;
  assign n6461 = n915 ^ n478 ^ n234 ;
  assign n6459 = n644 & ~n2785 ;
  assign n6460 = n6459 ^ n665 ^ 1'b0 ;
  assign n6462 = n6461 ^ n6460 ^ n814 ;
  assign n6463 = n716 | n5974 ;
  assign n6464 = n390 & ~n6463 ;
  assign n6465 = n6462 | n6464 ;
  assign n6466 = n2236 & ~n6465 ;
  assign n6467 = n614 & ~n6466 ;
  assign n6473 = n1778 & n4381 ;
  assign n6474 = n6473 ^ n2255 ^ 1'b0 ;
  assign n6468 = n788 | n2380 ;
  assign n6469 = n773 & ~n6468 ;
  assign n6470 = n275 | n6469 ;
  assign n6471 = n6470 ^ n3106 ^ 1'b0 ;
  assign n6472 = n947 | n6471 ;
  assign n6475 = n6474 ^ n6472 ^ n356 ;
  assign n6477 = ( n568 & ~n1544 ) | ( n568 & n5225 ) | ( ~n1544 & n5225 ) ;
  assign n6476 = n4139 ^ n3374 ^ 1'b0 ;
  assign n6478 = n6477 ^ n6476 ^ n1867 ;
  assign n6487 = n4471 ^ n2159 ^ n1900 ;
  assign n6479 = x49 & n441 ;
  assign n6480 = n6479 ^ n286 ^ 1'b0 ;
  assign n6481 = ( n2411 & n5570 ) | ( n2411 & ~n6480 ) | ( n5570 & ~n6480 ) ;
  assign n6482 = n2043 & n4069 ;
  assign n6483 = n2278 ^ x18 ^ 1'b0 ;
  assign n6484 = n6483 ^ n5871 ^ 1'b0 ;
  assign n6485 = n6482 & n6484 ;
  assign n6486 = ~n6481 & n6485 ;
  assign n6488 = n6487 ^ n6486 ^ 1'b0 ;
  assign n6489 = n6409 ^ n3854 ^ 1'b0 ;
  assign n6490 = ( ~n1065 & n2924 ) | ( ~n1065 & n4182 ) | ( n2924 & n4182 ) ;
  assign n6491 = n5597 ^ n2290 ^ 1'b0 ;
  assign n6492 = ~n3083 & n6491 ;
  assign n6493 = ( ~n5340 & n6490 ) | ( ~n5340 & n6492 ) | ( n6490 & n6492 ) ;
  assign n6504 = n2347 & ~n2877 ;
  assign n6499 = ( n131 & n337 ) | ( n131 & n517 ) | ( n337 & n517 ) ;
  assign n6494 = n2299 ^ n130 ^ 1'b0 ;
  assign n6495 = n6494 ^ n4185 ^ n3176 ;
  assign n6496 = ~n2188 & n6495 ;
  assign n6497 = n1592 & ~n2379 ;
  assign n6498 = n6496 & n6497 ;
  assign n6500 = n6499 ^ n6498 ^ n2325 ;
  assign n6501 = n6500 ^ n3926 ^ n3305 ;
  assign n6502 = n1624 | n2278 ;
  assign n6503 = n6501 & ~n6502 ;
  assign n6505 = n6504 ^ n6503 ^ n3599 ;
  assign n6506 = n1194 | n5061 ;
  assign n6507 = n3976 ^ n2293 ^ n2016 ;
  assign n6508 = ( n2660 & n6506 ) | ( n2660 & ~n6507 ) | ( n6506 & ~n6507 ) ;
  assign n6509 = ( n710 & n1250 ) | ( n710 & n6508 ) | ( n1250 & n6508 ) ;
  assign n6510 = n6509 ^ n2490 ^ 1'b0 ;
  assign n6511 = x7 & ~n807 ;
  assign n6512 = n6510 & n6511 ;
  assign n6513 = n5052 & n5694 ;
  assign n6514 = n6265 ^ n822 ^ 1'b0 ;
  assign n6515 = n6513 | n6514 ;
  assign n6516 = n4393 ^ n2147 ^ 1'b0 ;
  assign n6517 = n6516 ^ n2580 ^ 1'b0 ;
  assign n6519 = n2612 ^ n2580 ^ 1'b0 ;
  assign n6518 = ~n5689 & n6283 ;
  assign n6520 = n6519 ^ n6518 ^ 1'b0 ;
  assign n6521 = n3614 & n5925 ;
  assign n6522 = n4862 & n6521 ;
  assign n6523 = n1079 & ~n6522 ;
  assign n6524 = n6523 ^ x67 ^ 1'b0 ;
  assign n6525 = ( n163 & ~n2446 ) | ( n163 & n2720 ) | ( ~n2446 & n2720 ) ;
  assign n6526 = n6525 ^ n2167 ^ 1'b0 ;
  assign n6527 = ~n6524 & n6526 ;
  assign n6528 = n1783 & n3114 ;
  assign n6529 = n4546 ^ n2935 ^ 1'b0 ;
  assign n6530 = n3586 | n5784 ;
  assign n6531 = n6529 & ~n6530 ;
  assign n6532 = n322 | n1472 ;
  assign n6533 = n3850 & n6532 ;
  assign n6534 = n6533 ^ n4094 ^ n1203 ;
  assign n6542 = n2239 & ~n4324 ;
  assign n6543 = n2599 & n6542 ;
  assign n6544 = ( n592 & n6404 ) | ( n592 & ~n6543 ) | ( n6404 & ~n6543 ) ;
  assign n6538 = n161 & ~n4957 ;
  assign n6539 = n2367 & n6538 ;
  assign n6540 = ( n2083 & n2761 ) | ( n2083 & n6539 ) | ( n2761 & n6539 ) ;
  assign n6541 = n6540 ^ n3636 ^ n1024 ;
  assign n6535 = ( x47 & n483 ) | ( x47 & n783 ) | ( n483 & n783 ) ;
  assign n6536 = n2539 & ~n6535 ;
  assign n6537 = n6536 ^ n2276 ^ 1'b0 ;
  assign n6545 = n6544 ^ n6541 ^ n6537 ;
  assign n6546 = n1470 & ~n1725 ;
  assign n6547 = n3686 ^ n2612 ^ 1'b0 ;
  assign n6548 = n6546 & ~n6547 ;
  assign n6549 = ~n811 & n880 ;
  assign n6550 = n6549 ^ n3316 ^ 1'b0 ;
  assign n6551 = n6550 ^ n5364 ^ n1693 ;
  assign n6552 = n4987 ^ n3395 ^ 1'b0 ;
  assign n6553 = n6551 | n6552 ;
  assign n6557 = n6005 ^ n440 ^ 1'b0 ;
  assign n6558 = n310 & ~n6557 ;
  assign n6554 = n1526 | n5597 ;
  assign n6555 = n533 & ~n6554 ;
  assign n6556 = n3063 & ~n6555 ;
  assign n6559 = n6558 ^ n6556 ^ 1'b0 ;
  assign n6560 = n3146 & ~n6559 ;
  assign n6561 = n1496 ^ n844 ^ 1'b0 ;
  assign n6565 = x105 & n1749 ;
  assign n6566 = n6565 ^ n691 ^ 1'b0 ;
  assign n6562 = n2994 ^ n2467 ^ 1'b0 ;
  assign n6563 = ~n5108 & n6562 ;
  assign n6564 = n6563 ^ n5936 ^ 1'b0 ;
  assign n6567 = n6566 ^ n6564 ^ 1'b0 ;
  assign n6569 = n1105 & n3213 ;
  assign n6570 = n6569 ^ n510 ^ 1'b0 ;
  assign n6568 = ( n1393 & n2706 ) | ( n1393 & ~n2808 ) | ( n2706 & ~n2808 ) ;
  assign n6571 = n6570 ^ n6568 ^ n1878 ;
  assign n6572 = n6571 ^ n5438 ^ 1'b0 ;
  assign n6573 = n6567 & n6572 ;
  assign n6574 = n6078 ^ n4442 ^ n2276 ;
  assign n6575 = n646 & n985 ;
  assign n6576 = n6575 ^ n6335 ^ n1847 ;
  assign n6577 = ( n3328 & n3938 ) | ( n3328 & n5677 ) | ( n3938 & n5677 ) ;
  assign n6578 = ~x98 & n6577 ;
  assign n6579 = n958 ^ n450 ^ 1'b0 ;
  assign n6580 = ~n399 & n6579 ;
  assign n6581 = ~n5103 & n6580 ;
  assign n6582 = ( n355 & n5342 ) | ( n355 & n6055 ) | ( n5342 & n6055 ) ;
  assign n6583 = n6582 ^ n3903 ^ 1'b0 ;
  assign n6584 = n3853 & ~n6583 ;
  assign n6598 = n5144 ^ n2637 ^ 1'b0 ;
  assign n6586 = ( n304 & n619 ) | ( n304 & n4824 ) | ( n619 & n4824 ) ;
  assign n6585 = n5070 ^ n4879 ^ 1'b0 ;
  assign n6587 = n6586 ^ n6585 ^ n867 ;
  assign n6594 = ( ~n1186 & n1847 ) | ( ~n1186 & n2171 ) | ( n1847 & n2171 ) ;
  assign n6595 = n6594 ^ n6223 ^ n1443 ;
  assign n6591 = n1991 & ~n2420 ;
  assign n6592 = ~n1570 & n6591 ;
  assign n6588 = n916 ^ x81 ^ 1'b0 ;
  assign n6589 = n6588 ^ n4815 ^ 1'b0 ;
  assign n6590 = n6589 ^ n2319 ^ n249 ;
  assign n6593 = n6592 ^ n6590 ^ n2251 ;
  assign n6596 = n6595 ^ n6593 ^ n5036 ;
  assign n6597 = n6587 & n6596 ;
  assign n6599 = n6598 ^ n6597 ^ 1'b0 ;
  assign n6600 = n3302 ^ n1443 ^ x123 ;
  assign n6601 = ( n733 & n990 ) | ( n733 & ~n1251 ) | ( n990 & ~n1251 ) ;
  assign n6602 = n1268 | n4562 ;
  assign n6603 = n5675 & ~n6602 ;
  assign n6604 = n418 | n6603 ;
  assign n6605 = n6604 ^ n1214 ^ 1'b0 ;
  assign n6606 = ( ~n2373 & n4353 ) | ( ~n2373 & n4891 ) | ( n4353 & n4891 ) ;
  assign n6607 = ~n6254 & n6606 ;
  assign n6608 = n1714 ^ n326 ^ 1'b0 ;
  assign n6609 = n3631 | n6608 ;
  assign n6610 = n6609 ^ n3671 ^ n970 ;
  assign n6611 = n1947 & n5271 ;
  assign n6612 = n2131 ^ n481 ^ 1'b0 ;
  assign n6613 = n3585 | n6612 ;
  assign n6614 = n6613 ^ n4639 ^ n1844 ;
  assign n6618 = n1264 & n2348 ;
  assign n6619 = ( n362 & ~n828 ) | ( n362 & n6618 ) | ( ~n828 & n6618 ) ;
  assign n6620 = ( n549 & ~n3153 ) | ( n549 & n6619 ) | ( ~n3153 & n6619 ) ;
  assign n6617 = ~n4333 & n6220 ;
  assign n6615 = n3383 ^ n2178 ^ 1'b0 ;
  assign n6616 = n3794 | n6615 ;
  assign n6621 = n6620 ^ n6617 ^ n6616 ;
  assign n6623 = ~n2376 & n2397 ;
  assign n6622 = n2075 & ~n2653 ;
  assign n6624 = n6623 ^ n6622 ^ 1'b0 ;
  assign n6625 = x83 & n887 ;
  assign n6626 = n6625 ^ n1977 ^ 1'b0 ;
  assign n6627 = n1820 | n2131 ;
  assign n6628 = ( n2057 & n6626 ) | ( n2057 & ~n6627 ) | ( n6626 & ~n6627 ) ;
  assign n6629 = n6628 ^ n4276 ^ 1'b0 ;
  assign n6630 = n302 | n6629 ;
  assign n6631 = n3736 ^ n1126 ^ 1'b0 ;
  assign n6632 = n338 & ~n6631 ;
  assign n6633 = ( ~n1714 & n6461 ) | ( ~n1714 & n6632 ) | ( n6461 & n6632 ) ;
  assign n6636 = n5864 ^ n4458 ^ n4039 ;
  assign n6634 = ( n1109 & ~n2086 ) | ( n1109 & n3596 ) | ( ~n2086 & n3596 ) ;
  assign n6635 = n6634 ^ n2588 ^ n393 ;
  assign n6637 = n6636 ^ n6635 ^ n4242 ;
  assign n6639 = ( n1355 & ~n1409 ) | ( n1355 & n1530 ) | ( ~n1409 & n1530 ) ;
  assign n6640 = ( n1022 & ~n2269 ) | ( n1022 & n6639 ) | ( ~n2269 & n6639 ) ;
  assign n6641 = n6640 ^ x113 ^ 1'b0 ;
  assign n6638 = ( ~n247 & n1630 ) | ( ~n247 & n4290 ) | ( n1630 & n4290 ) ;
  assign n6642 = n6641 ^ n6638 ^ n1091 ;
  assign n6643 = n2689 ^ n1911 ^ n1839 ;
  assign n6644 = n6643 ^ n2734 ^ n235 ;
  assign n6646 = ( ~n617 & n900 ) | ( ~n617 & n3447 ) | ( n900 & n3447 ) ;
  assign n6647 = n906 ^ n744 ^ 1'b0 ;
  assign n6648 = n1867 & n6647 ;
  assign n6649 = ( n1771 & n6646 ) | ( n1771 & n6648 ) | ( n6646 & n6648 ) ;
  assign n6645 = x99 & n1681 ;
  assign n6650 = n6649 ^ n6645 ^ 1'b0 ;
  assign n6651 = ( n1210 & n6644 ) | ( n1210 & ~n6650 ) | ( n6644 & ~n6650 ) ;
  assign n6652 = n6651 ^ n5076 ^ n4184 ;
  assign n6653 = ( n2781 & n2833 ) | ( n2781 & ~n2903 ) | ( n2833 & ~n2903 ) ;
  assign n6654 = n6570 ^ n3468 ^ n1419 ;
  assign n6655 = ( ~n1017 & n5539 ) | ( ~n1017 & n6654 ) | ( n5539 & n6654 ) ;
  assign n6656 = ( ~n2498 & n2770 ) | ( ~n2498 & n2982 ) | ( n2770 & n2982 ) ;
  assign n6657 = n6656 ^ n913 ^ 1'b0 ;
  assign n6658 = n3562 ^ n444 ^ 1'b0 ;
  assign n6659 = n6658 ^ n2126 ^ n247 ;
  assign n6660 = n4320 ^ n1153 ^ 1'b0 ;
  assign n6661 = ~n1043 & n6660 ;
  assign n6662 = ( n4224 & n6659 ) | ( n4224 & n6661 ) | ( n6659 & n6661 ) ;
  assign n6663 = n5549 ^ n5042 ^ n131 ;
  assign n6664 = n476 | n3956 ;
  assign n6665 = n6664 ^ n4824 ^ 1'b0 ;
  assign n6666 = n5469 | n6665 ;
  assign n6667 = n6666 ^ n3928 ^ 1'b0 ;
  assign n6668 = n2025 | n6667 ;
  assign n6674 = ( n988 & n1856 ) | ( n988 & ~n2124 ) | ( n1856 & ~n2124 ) ;
  assign n6675 = n6674 ^ n5865 ^ n1783 ;
  assign n6672 = ( n345 & n1628 ) | ( n345 & n2269 ) | ( n1628 & n2269 ) ;
  assign n6669 = ( ~n1166 & n2141 ) | ( ~n1166 & n2629 ) | ( n2141 & n2629 ) ;
  assign n6670 = ( x34 & n2928 ) | ( x34 & ~n3011 ) | ( n2928 & ~n3011 ) ;
  assign n6671 = ( n3898 & ~n6669 ) | ( n3898 & n6670 ) | ( ~n6669 & n6670 ) ;
  assign n6673 = n6672 ^ n6671 ^ n2777 ;
  assign n6676 = n6675 ^ n6673 ^ 1'b0 ;
  assign n6677 = n5775 & n6676 ;
  assign n6678 = n892 & ~n1143 ;
  assign n6679 = n6678 ^ n1518 ^ 1'b0 ;
  assign n6680 = n4888 ^ n1679 ^ 1'b0 ;
  assign n6681 = n6679 & n6680 ;
  assign n6682 = n6681 ^ n1747 ^ 1'b0 ;
  assign n6683 = n6682 ^ n1518 ^ 1'b0 ;
  assign n6684 = n6325 ^ n5756 ^ 1'b0 ;
  assign n6685 = n476 | n1316 ;
  assign n6686 = ( n3409 & ~n3919 ) | ( n3409 & n5955 ) | ( ~n3919 & n5955 ) ;
  assign n6687 = n5820 ^ n2446 ^ 1'b0 ;
  assign n6688 = ( n1541 & n3284 ) | ( n1541 & ~n3553 ) | ( n3284 & ~n3553 ) ;
  assign n6689 = n6688 ^ n1711 ^ 1'b0 ;
  assign n6694 = n895 & ~n4019 ;
  assign n6695 = n3308 & n6694 ;
  assign n6692 = n825 & n2909 ;
  assign n6693 = n6692 ^ n3794 ^ n1130 ;
  assign n6690 = ( n443 & n909 ) | ( n443 & n1782 ) | ( n909 & n1782 ) ;
  assign n6691 = n6690 ^ n2622 ^ n1587 ;
  assign n6696 = n6695 ^ n6693 ^ n6691 ;
  assign n6697 = ( ~n597 & n1021 ) | ( ~n597 & n5931 ) | ( n1021 & n5931 ) ;
  assign n6698 = ~n583 & n6697 ;
  assign n6699 = n155 & n287 ;
  assign n6700 = n2847 ^ n1430 ^ n1356 ;
  assign n6701 = ( n726 & n4098 ) | ( n726 & n6700 ) | ( n4098 & n6700 ) ;
  assign n6702 = n3451 | n6701 ;
  assign n6703 = n6702 ^ n3530 ^ 1'b0 ;
  assign n6704 = n6699 & ~n6703 ;
  assign n6705 = ~n4774 & n6704 ;
  assign n6706 = ( n996 & n5558 ) | ( n996 & ~n6639 ) | ( n5558 & ~n6639 ) ;
  assign n6707 = ( n2818 & ~n4043 ) | ( n2818 & n5587 ) | ( ~n4043 & n5587 ) ;
  assign n6708 = n6707 ^ n4813 ^ n1193 ;
  assign n6709 = n6708 ^ n2273 ^ 1'b0 ;
  assign n6710 = n5232 ^ n3499 ^ n2218 ;
  assign n6711 = ( n2081 & n3243 ) | ( n2081 & ~n6710 ) | ( n3243 & ~n6710 ) ;
  assign n6712 = n5490 ^ n2837 ^ x3 ;
  assign n6713 = n2151 | n2584 ;
  assign n6714 = n6713 ^ n2718 ^ 1'b0 ;
  assign n6715 = n6714 ^ n3956 ^ n691 ;
  assign n6716 = n6712 & n6715 ;
  assign n6717 = n6716 ^ n4288 ^ 1'b0 ;
  assign n6718 = ~n6705 & n6717 ;
  assign n6719 = ( ~n2197 & n2818 ) | ( ~n2197 & n4977 ) | ( n2818 & n4977 ) ;
  assign n6720 = ( n686 & ~n2515 ) | ( n686 & n6719 ) | ( ~n2515 & n6719 ) ;
  assign n6721 = ( n3193 & n3996 ) | ( n3193 & ~n6720 ) | ( n3996 & ~n6720 ) ;
  assign n6722 = n1664 ^ n1463 ^ 1'b0 ;
  assign n6725 = ~n483 & n2794 ;
  assign n6726 = n1533 & n6725 ;
  assign n6723 = n5587 ^ n5145 ^ 1'b0 ;
  assign n6724 = ~n1346 & n6723 ;
  assign n6727 = n6726 ^ n6724 ^ 1'b0 ;
  assign n6731 = ( n1005 & ~n2079 ) | ( n1005 & n4723 ) | ( ~n2079 & n4723 ) ;
  assign n6729 = n4986 ^ n418 ^ n275 ;
  assign n6730 = n6729 ^ n230 ^ 1'b0 ;
  assign n6728 = n4298 ^ n155 ^ 1'b0 ;
  assign n6732 = n6731 ^ n6730 ^ n6728 ;
  assign n6733 = n6732 ^ n5458 ^ n1870 ;
  assign n6737 = ( ~n1552 & n2393 ) | ( ~n1552 & n4855 ) | ( n2393 & n4855 ) ;
  assign n6734 = n909 & n1684 ;
  assign n6735 = n6734 ^ n2666 ^ 1'b0 ;
  assign n6736 = ~n1635 & n6735 ;
  assign n6738 = n6737 ^ n6736 ^ 1'b0 ;
  assign n6739 = n2611 | n3217 ;
  assign n6740 = n6739 ^ n974 ^ n795 ;
  assign n6741 = ( ~n1409 & n3834 ) | ( ~n1409 & n4287 ) | ( n3834 & n4287 ) ;
  assign n6742 = ( n5476 & ~n6213 ) | ( n5476 & n6741 ) | ( ~n6213 & n6741 ) ;
  assign n6743 = ( n1375 & n5229 ) | ( n1375 & n6742 ) | ( n5229 & n6742 ) ;
  assign n6744 = n2065 ^ n1910 ^ 1'b0 ;
  assign n6745 = n6744 ^ n2323 ^ 1'b0 ;
  assign n6746 = x32 & n6745 ;
  assign n6747 = n6746 ^ n3667 ^ n294 ;
  assign n6748 = n6747 ^ n5756 ^ n1504 ;
  assign n6749 = n2527 ^ n1392 ^ 1'b0 ;
  assign n6750 = n1949 ^ n1590 ^ n345 ;
  assign n6751 = ( x102 & n6270 ) | ( x102 & n6750 ) | ( n6270 & n6750 ) ;
  assign n6752 = n5609 | n6751 ;
  assign n6753 = n2760 | n5436 ;
  assign n6754 = n6753 ^ n3812 ^ 1'b0 ;
  assign n6755 = ~n4542 & n6754 ;
  assign n6756 = n6755 ^ n3289 ^ 1'b0 ;
  assign n6757 = ( ~n313 & n633 ) | ( ~n313 & n6756 ) | ( n633 & n6756 ) ;
  assign n6758 = n130 & n5859 ;
  assign n6759 = ~n4944 & n6299 ;
  assign n6760 = n6759 ^ n2120 ^ 1'b0 ;
  assign n6761 = ( n483 & ~n625 ) | ( n483 & n6760 ) | ( ~n625 & n6760 ) ;
  assign n6762 = n6356 ^ n3650 ^ 1'b0 ;
  assign n6763 = ( n1180 & n3280 ) | ( n1180 & ~n4304 ) | ( n3280 & ~n4304 ) ;
  assign n6765 = ( ~n424 & n1419 ) | ( ~n424 & n3990 ) | ( n1419 & n3990 ) ;
  assign n6764 = ~n1589 & n2487 ;
  assign n6766 = n6765 ^ n6764 ^ 1'b0 ;
  assign n6767 = ( n3212 & n6763 ) | ( n3212 & n6766 ) | ( n6763 & n6766 ) ;
  assign n6768 = ( n179 & n6762 ) | ( n179 & n6767 ) | ( n6762 & n6767 ) ;
  assign n6769 = n2174 & n2414 ;
  assign n6770 = ~n545 & n6769 ;
  assign n6771 = ( n3351 & n3433 ) | ( n3351 & ~n6770 ) | ( n3433 & ~n6770 ) ;
  assign n6772 = n990 & ~n4396 ;
  assign n6773 = n2070 & n6772 ;
  assign n6774 = n6773 ^ n2126 ^ n751 ;
  assign n6775 = n6039 ^ n2510 ^ n248 ;
  assign n6776 = ( n1283 & n2033 ) | ( n1283 & ~n4770 ) | ( n2033 & ~n4770 ) ;
  assign n6782 = n348 & ~n610 ;
  assign n6783 = n6782 ^ n1141 ^ 1'b0 ;
  assign n6781 = ( ~n719 & n934 ) | ( ~n719 & n2339 ) | ( n934 & n2339 ) ;
  assign n6777 = n4185 ^ n2348 ^ 1'b0 ;
  assign n6778 = n4222 & ~n6777 ;
  assign n6779 = n2175 ^ n1364 ^ 1'b0 ;
  assign n6780 = n6778 & n6779 ;
  assign n6784 = n6783 ^ n6781 ^ n6780 ;
  assign n6785 = n6776 & n6784 ;
  assign n6786 = n6785 ^ n2249 ^ 1'b0 ;
  assign n6787 = ( n3045 & n6775 ) | ( n3045 & ~n6786 ) | ( n6775 & ~n6786 ) ;
  assign n6788 = x108 & ~n4535 ;
  assign n6789 = n6788 ^ n2075 ^ 1'b0 ;
  assign n6790 = n6789 ^ n385 ^ 1'b0 ;
  assign n6791 = n1378 | n2494 ;
  assign n6792 = n6790 | n6791 ;
  assign n6795 = ( n368 & ~n438 ) | ( n368 & n1828 ) | ( ~n438 & n1828 ) ;
  assign n6796 = ( n1977 & ~n3134 ) | ( n1977 & n6795 ) | ( ~n3134 & n6795 ) ;
  assign n6793 = n1649 ^ n849 ^ 1'b0 ;
  assign n6794 = ( n1752 & n2116 ) | ( n1752 & ~n6793 ) | ( n2116 & ~n6793 ) ;
  assign n6797 = n6796 ^ n6794 ^ n6619 ;
  assign n6798 = n619 ^ x114 ^ 1'b0 ;
  assign n6799 = x39 & n3272 ;
  assign n6805 = n3023 ^ n1397 ^ n614 ;
  assign n6800 = ( n3376 & n4946 ) | ( n3376 & ~n5508 ) | ( n4946 & ~n5508 ) ;
  assign n6801 = ( ~n744 & n760 ) | ( ~n744 & n1183 ) | ( n760 & n1183 ) ;
  assign n6802 = n2623 ^ n1329 ^ 1'b0 ;
  assign n6803 = ( ~n2514 & n6801 ) | ( ~n2514 & n6802 ) | ( n6801 & n6802 ) ;
  assign n6804 = ~n6800 & n6803 ;
  assign n6806 = n6805 ^ n6804 ^ n1762 ;
  assign n6807 = n5454 ^ n1295 ^ 1'b0 ;
  assign n6808 = ( n3125 & ~n4493 ) | ( n3125 & n6807 ) | ( ~n4493 & n6807 ) ;
  assign n6809 = n2381 ^ n148 ^ 1'b0 ;
  assign n6810 = ~n270 & n1097 ;
  assign n6811 = ( n1940 & n3180 ) | ( n1940 & ~n6810 ) | ( n3180 & ~n6810 ) ;
  assign n6812 = ( ~n1583 & n6809 ) | ( ~n1583 & n6811 ) | ( n6809 & n6811 ) ;
  assign n6813 = n5093 ^ n1444 ^ 1'b0 ;
  assign n6814 = ~n3724 & n6813 ;
  assign n6815 = n6814 ^ n4767 ^ n2209 ;
  assign n6816 = ( ~n5025 & n6812 ) | ( ~n5025 & n6815 ) | ( n6812 & n6815 ) ;
  assign n6817 = ~n825 & n2797 ;
  assign n6818 = ~n356 & n6817 ;
  assign n6819 = n6818 ^ n5859 ^ n5178 ;
  assign n6820 = n3610 ^ n2773 ^ 1'b0 ;
  assign n6821 = n4274 & ~n6820 ;
  assign n6822 = n6821 ^ n3422 ^ 1'b0 ;
  assign n6823 = n6822 ^ n4087 ^ n3210 ;
  assign n6824 = ( n512 & n1247 ) | ( n512 & n3697 ) | ( n1247 & n3697 ) ;
  assign n6825 = n6824 ^ n2030 ^ 1'b0 ;
  assign n6830 = n3626 ^ n586 ^ 1'b0 ;
  assign n6826 = ( n2057 & ~n2419 ) | ( n2057 & n2745 ) | ( ~n2419 & n2745 ) ;
  assign n6827 = n6826 ^ n2895 ^ n2189 ;
  assign n6828 = n4036 ^ n2883 ^ n1034 ;
  assign n6829 = n6827 & ~n6828 ;
  assign n6831 = n6830 ^ n6829 ^ 1'b0 ;
  assign n6832 = n6831 ^ n2042 ^ n1427 ;
  assign n6833 = n6832 ^ n5534 ^ 1'b0 ;
  assign n6834 = ( n3632 & n6382 ) | ( n3632 & n6830 ) | ( n6382 & n6830 ) ;
  assign n6836 = ( n3205 & n4497 ) | ( n3205 & ~n5220 ) | ( n4497 & ~n5220 ) ;
  assign n6835 = n4370 ^ n1320 ^ n1240 ;
  assign n6837 = n6836 ^ n6835 ^ n1622 ;
  assign n6838 = n6283 ^ n2207 ^ n1875 ;
  assign n6839 = n6838 ^ n4450 ^ n2479 ;
  assign n6840 = n5286 ^ n1189 ^ n884 ;
  assign n6841 = n6840 ^ n5212 ^ 1'b0 ;
  assign n6842 = ~n1450 & n2102 ;
  assign n6843 = n1052 | n4616 ;
  assign n6844 = n6842 | n6843 ;
  assign n6850 = ( n1872 & n2754 ) | ( n1872 & n3732 ) | ( n2754 & n3732 ) ;
  assign n6845 = n1193 ^ n223 ^ 1'b0 ;
  assign n6846 = ~n5773 & n6845 ;
  assign n6847 = ~n4434 & n6846 ;
  assign n6848 = n6793 ^ n6198 ^ 1'b0 ;
  assign n6849 = n6847 | n6848 ;
  assign n6851 = n6850 ^ n6849 ^ n2206 ;
  assign n6852 = n399 ^ n305 ^ 1'b0 ;
  assign n6853 = ~n3151 & n6852 ;
  assign n6854 = n3030 ^ n1736 ^ 1'b0 ;
  assign n6855 = n6853 & n6854 ;
  assign n6856 = n6712 ^ n4612 ^ 1'b0 ;
  assign n6857 = ( n1668 & n3487 ) | ( n1668 & ~n4622 ) | ( n3487 & ~n4622 ) ;
  assign n6858 = n5587 & n6857 ;
  assign n6859 = n6858 ^ n832 ^ 1'b0 ;
  assign n6866 = n5364 ^ n1813 ^ 1'b0 ;
  assign n6860 = n4994 ^ n1132 ^ n760 ;
  assign n6861 = n5587 ^ n4698 ^ n520 ;
  assign n6862 = n1698 ^ n1296 ^ 1'b0 ;
  assign n6863 = n6862 ^ n6608 ^ n2584 ;
  assign n6864 = ( n1127 & n6861 ) | ( n1127 & ~n6863 ) | ( n6861 & ~n6863 ) ;
  assign n6865 = ( ~n1886 & n6860 ) | ( ~n1886 & n6864 ) | ( n6860 & n6864 ) ;
  assign n6867 = n6866 ^ n6865 ^ n5224 ;
  assign n6870 = n6480 ^ n2587 ^ n2253 ;
  assign n6871 = n905 & n6870 ;
  assign n6868 = n2086 ^ n1379 ^ 1'b0 ;
  assign n6869 = n4946 | n6868 ;
  assign n6872 = n6871 ^ n6869 ^ 1'b0 ;
  assign n6873 = n441 & n1166 ;
  assign n6874 = ( n509 & ~n754 ) | ( n509 & n3509 ) | ( ~n754 & n3509 ) ;
  assign n6875 = n6874 ^ n4910 ^ n4414 ;
  assign n6876 = n2012 & n3689 ;
  assign n6877 = ~n273 & n6876 ;
  assign n6878 = n199 & ~n6877 ;
  assign n6879 = n5568 ^ n3936 ^ 1'b0 ;
  assign n6880 = ( n3041 & n4705 ) | ( n3041 & ~n6879 ) | ( n4705 & ~n6879 ) ;
  assign n6881 = ( ~n2193 & n2474 ) | ( ~n2193 & n4911 ) | ( n2474 & n4911 ) ;
  assign n6882 = n2126 & ~n3640 ;
  assign n6883 = n6881 & n6882 ;
  assign n6884 = ( n1859 & n2547 ) | ( n1859 & n3762 ) | ( n2547 & n3762 ) ;
  assign n6885 = ( n1835 & ~n3088 ) | ( n1835 & n4447 ) | ( ~n3088 & n4447 ) ;
  assign n6886 = n3335 & ~n6885 ;
  assign n6887 = n6884 & n6886 ;
  assign n6888 = n6883 | n6887 ;
  assign n6889 = n4939 | n6888 ;
  assign n6893 = ( n288 & n2991 ) | ( n288 & n4120 ) | ( n2991 & n4120 ) ;
  assign n6894 = n316 | n1828 ;
  assign n6895 = n1118 & ~n6894 ;
  assign n6896 = x51 & ~n6895 ;
  assign n6897 = ( n3125 & n6893 ) | ( n3125 & ~n6896 ) | ( n6893 & ~n6896 ) ;
  assign n6890 = ~n566 & n1059 ;
  assign n6891 = n3114 & n6890 ;
  assign n6892 = n6112 | n6891 ;
  assign n6898 = n6897 ^ n6892 ^ 1'b0 ;
  assign n6899 = n6053 ^ n3633 ^ n1040 ;
  assign n6904 = x50 & n1798 ;
  assign n6905 = n6904 ^ n1261 ^ 1'b0 ;
  assign n6900 = ( x21 & ~n1955 ) | ( x21 & n2928 ) | ( ~n1955 & n2928 ) ;
  assign n6901 = ( n786 & n867 ) | ( n786 & n2294 ) | ( n867 & n2294 ) ;
  assign n6902 = n6900 & ~n6901 ;
  assign n6903 = ~n6219 & n6902 ;
  assign n6906 = n6905 ^ n6903 ^ n223 ;
  assign n6907 = ( n3101 & ~n6899 ) | ( n3101 & n6906 ) | ( ~n6899 & n6906 ) ;
  assign n6908 = n254 & ~n924 ;
  assign n6909 = n6908 ^ n2788 ^ 1'b0 ;
  assign n6910 = n1209 | n6909 ;
  assign n6911 = ( x41 & ~n5230 ) | ( x41 & n6286 ) | ( ~n5230 & n6286 ) ;
  assign n6912 = n3145 & n4114 ;
  assign n6913 = ~n6014 & n6912 ;
  assign n6914 = ( n989 & n3036 ) | ( n989 & n6913 ) | ( n3036 & n6913 ) ;
  assign n6915 = ( n2181 & n2611 ) | ( n2181 & ~n5844 ) | ( n2611 & ~n5844 ) ;
  assign n6916 = ( x2 & n1355 ) | ( x2 & ~n6915 ) | ( n1355 & ~n6915 ) ;
  assign n6917 = ~n6914 & n6916 ;
  assign n6918 = n4635 & n6917 ;
  assign n6919 = ( n4954 & n5947 ) | ( n4954 & ~n6918 ) | ( n5947 & ~n6918 ) ;
  assign n6920 = n645 | n1933 ;
  assign n6921 = ( n1359 & n5573 ) | ( n1359 & n6255 ) | ( n5573 & n6255 ) ;
  assign n6922 = n624 | n5371 ;
  assign n6923 = ~n3808 & n5483 ;
  assign n6924 = n6923 ^ n4023 ^ 1'b0 ;
  assign n6925 = ~n1142 & n3764 ;
  assign n6926 = n2883 & n6925 ;
  assign n6927 = n6926 ^ n3693 ^ 1'b0 ;
  assign n6928 = ( n598 & n3401 ) | ( n598 & ~n5891 ) | ( n3401 & ~n5891 ) ;
  assign n6929 = n2343 & n6928 ;
  assign n6930 = n586 ^ n297 ^ 1'b0 ;
  assign n6931 = n1059 & n6930 ;
  assign n6932 = n3237 | n6931 ;
  assign n6933 = n3693 & ~n6932 ;
  assign n6934 = ~n5706 & n6933 ;
  assign n6935 = n6929 & ~n6934 ;
  assign n6936 = n6935 ^ n1038 ^ 1'b0 ;
  assign n6937 = x23 & n1132 ;
  assign n6938 = n6937 ^ n6067 ^ n3402 ;
  assign n6939 = x101 & n6397 ;
  assign n6940 = ( ~n5023 & n6938 ) | ( ~n5023 & n6939 ) | ( n6938 & n6939 ) ;
  assign n6944 = n3955 ^ n2327 ^ 1'b0 ;
  assign n6945 = n750 & n6944 ;
  assign n6946 = ~n3330 & n6945 ;
  assign n6947 = n964 & n6946 ;
  assign n6941 = ( ~n872 & n2393 ) | ( ~n872 & n2969 ) | ( n2393 & n2969 ) ;
  assign n6942 = n6941 ^ n3915 ^ n696 ;
  assign n6943 = n1062 | n6942 ;
  assign n6948 = n6947 ^ n6943 ^ 1'b0 ;
  assign n6956 = n6555 ^ n4144 ^ 1'b0 ;
  assign n6957 = n2008 & ~n6956 ;
  assign n6958 = n6957 ^ n6181 ^ n4765 ;
  assign n6953 = ~n586 & n3892 ;
  assign n6954 = ~n665 & n6953 ;
  assign n6955 = n6954 ^ n6608 ^ 1'b0 ;
  assign n6952 = n6881 ^ n5977 ^ n5520 ;
  assign n6959 = n6958 ^ n6955 ^ n6952 ;
  assign n6949 = n1555 & n2224 ;
  assign n6950 = n563 & ~n6949 ;
  assign n6951 = n6950 ^ n1358 ^ 1'b0 ;
  assign n6960 = n6959 ^ n6951 ^ n5119 ;
  assign n6961 = ~n1038 & n4069 ;
  assign n6962 = n1192 ^ x76 ^ 1'b0 ;
  assign n6963 = n3365 | n6962 ;
  assign n6964 = ( n3906 & ~n6117 ) | ( n3906 & n6963 ) | ( ~n6117 & n6963 ) ;
  assign n6965 = n6964 ^ n2839 ^ n2785 ;
  assign n6966 = n2898 ^ n2392 ^ n1503 ;
  assign n6967 = ~n6965 & n6966 ;
  assign n6981 = ( ~n177 & n830 ) | ( ~n177 & n1401 ) | ( n830 & n1401 ) ;
  assign n6972 = ~n1318 & n2172 ;
  assign n6969 = n1137 & n1794 ;
  assign n6970 = n6969 ^ n5026 ^ 1'b0 ;
  assign n6971 = ( n2267 & n2468 ) | ( n2267 & ~n6970 ) | ( n2468 & ~n6970 ) ;
  assign n6973 = n6972 ^ n6971 ^ n4740 ;
  assign n6974 = n5203 & n6973 ;
  assign n6975 = n6974 ^ n6316 ^ n4443 ;
  assign n6976 = n2706 & n6975 ;
  assign n6977 = n6976 ^ n3511 ^ 1'b0 ;
  assign n6978 = x66 | n5739 ;
  assign n6979 = n3382 | n6978 ;
  assign n6980 = n6977 | n6979 ;
  assign n6968 = n1568 ^ n588 ^ 1'b0 ;
  assign n6982 = n6981 ^ n6980 ^ n6968 ;
  assign n6983 = ( ~n885 & n1350 ) | ( ~n885 & n2969 ) | ( n1350 & n2969 ) ;
  assign n6984 = ( n1614 & n5457 ) | ( n1614 & n5569 ) | ( n5457 & n5569 ) ;
  assign n6985 = ( n3107 & n6983 ) | ( n3107 & ~n6984 ) | ( n6983 & ~n6984 ) ;
  assign n6986 = n6985 ^ n4460 ^ 1'b0 ;
  assign n6987 = n6986 ^ n3161 ^ n2217 ;
  assign n6988 = n561 & n1626 ;
  assign n6989 = n6988 ^ n2822 ^ 1'b0 ;
  assign n6991 = n4245 ^ n1411 ^ n531 ;
  assign n6990 = n2239 & ~n3015 ;
  assign n6992 = n6991 ^ n6990 ^ n4005 ;
  assign n6993 = n6992 ^ n4322 ^ 1'b0 ;
  assign n6994 = n6989 | n6993 ;
  assign n6995 = n2429 & ~n6994 ;
  assign n6996 = n6995 ^ n3393 ^ 1'b0 ;
  assign n6999 = n3258 ^ n2427 ^ n1213 ;
  assign n6997 = n4875 ^ n2089 ^ 1'b0 ;
  assign n6998 = n1935 | n6997 ;
  assign n7000 = n6999 ^ n6998 ^ 1'b0 ;
  assign n7002 = ( ~n1430 & n2234 ) | ( ~n1430 & n2788 ) | ( n2234 & n2788 ) ;
  assign n7001 = n3664 ^ n1437 ^ 1'b0 ;
  assign n7003 = n7002 ^ n7001 ^ 1'b0 ;
  assign n7004 = n7003 ^ n4934 ^ 1'b0 ;
  assign n7013 = n445 & n6504 ;
  assign n7006 = n1883 & ~n4705 ;
  assign n7007 = n599 & n1078 ;
  assign n7008 = n7007 ^ n1809 ^ 1'b0 ;
  assign n7009 = ( n2788 & ~n2940 ) | ( n2788 & n7008 ) | ( ~n2940 & n7008 ) ;
  assign n7010 = n7006 & n7009 ;
  assign n7005 = x33 & ~n300 ;
  assign n7011 = n7010 ^ n7005 ^ 1'b0 ;
  assign n7012 = ~n4755 & n7011 ;
  assign n7014 = n7013 ^ n7012 ^ n218 ;
  assign n7015 = ~n714 & n4776 ;
  assign n7016 = n2256 ^ n1628 ^ 1'b0 ;
  assign n7017 = n5747 | n7016 ;
  assign n7018 = n6015 ^ n3990 ^ 1'b0 ;
  assign n7019 = n3519 & n7018 ;
  assign n7020 = n4820 & n7019 ;
  assign n7021 = n7020 ^ n566 ^ n209 ;
  assign n7022 = n4645 ^ n3401 ^ 1'b0 ;
  assign n7023 = n4353 ^ n2553 ^ 1'b0 ;
  assign n7024 = n7023 ^ n195 ^ 1'b0 ;
  assign n7025 = ( ~n2643 & n4887 ) | ( ~n2643 & n7024 ) | ( n4887 & n7024 ) ;
  assign n7026 = n7025 ^ n5227 ^ 1'b0 ;
  assign n7027 = n1911 | n7026 ;
  assign n7028 = ~n2895 & n3055 ;
  assign n7029 = n1778 & n2178 ;
  assign n7030 = n7029 ^ n1977 ^ 1'b0 ;
  assign n7031 = n3631 ^ n878 ^ n714 ;
  assign n7032 = n7031 ^ n4174 ^ x107 ;
  assign n7033 = ( n2548 & n7030 ) | ( n2548 & ~n7032 ) | ( n7030 & ~n7032 ) ;
  assign n7034 = n1539 | n6495 ;
  assign n7035 = ( ~n7028 & n7033 ) | ( ~n7028 & n7034 ) | ( n7033 & n7034 ) ;
  assign n7036 = n4701 ^ n2198 ^ 1'b0 ;
  assign n7037 = n3248 & ~n7036 ;
  assign n7038 = ( n374 & n4236 ) | ( n374 & ~n7037 ) | ( n4236 & ~n7037 ) ;
  assign n7039 = n663 | n7038 ;
  assign n7041 = n1081 ^ n733 ^ 1'b0 ;
  assign n7040 = n3030 | n3196 ;
  assign n7042 = n7041 ^ n7040 ^ 1'b0 ;
  assign n7043 = n6663 & ~n7042 ;
  assign n7044 = n1923 | n3356 ;
  assign n7045 = n7044 ^ n1452 ^ 1'b0 ;
  assign n7048 = n3011 & ~n3571 ;
  assign n7049 = n7048 ^ n3442 ^ 1'b0 ;
  assign n7047 = n772 | n1382 ;
  assign n7046 = ( n635 & n1298 ) | ( n635 & ~n2789 ) | ( n1298 & ~n2789 ) ;
  assign n7050 = n7049 ^ n7047 ^ n7046 ;
  assign n7051 = ( n1298 & n2206 ) | ( n1298 & n4729 ) | ( n2206 & n4729 ) ;
  assign n7052 = n7051 ^ n1695 ^ 1'b0 ;
  assign n7053 = n2163 & n6586 ;
  assign n7054 = n3947 ^ n1593 ^ 1'b0 ;
  assign n7055 = ~n7053 & n7054 ;
  assign n7056 = n2753 ^ n526 ^ 1'b0 ;
  assign n7057 = n7056 ^ n6241 ^ 1'b0 ;
  assign n7058 = n7055 & ~n7057 ;
  assign n7067 = x37 & n5391 ;
  assign n7059 = ( ~n1479 & n1590 ) | ( ~n1479 & n3428 ) | ( n1590 & n3428 ) ;
  assign n7060 = ( n3062 & n4574 ) | ( n3062 & ~n7059 ) | ( n4574 & ~n7059 ) ;
  assign n7061 = n7055 & ~n7060 ;
  assign n7062 = ( ~n825 & n1806 ) | ( ~n825 & n2200 ) | ( n1806 & n2200 ) ;
  assign n7063 = n6775 ^ n6156 ^ 1'b0 ;
  assign n7064 = n1643 | n7063 ;
  assign n7065 = ( n4773 & n7062 ) | ( n4773 & n7064 ) | ( n7062 & n7064 ) ;
  assign n7066 = n7061 & n7065 ;
  assign n7068 = n7067 ^ n7066 ^ 1'b0 ;
  assign n7069 = n7068 ^ n2847 ^ 1'b0 ;
  assign n7070 = n3007 ^ n2433 ^ 1'b0 ;
  assign n7071 = n2411 | n7070 ;
  assign n7072 = n1839 & n1982 ;
  assign n7073 = n1272 & n7072 ;
  assign n7074 = ( n1419 & n7071 ) | ( n1419 & ~n7073 ) | ( n7071 & ~n7073 ) ;
  assign n7075 = n7074 ^ n252 ^ 1'b0 ;
  assign n7076 = n2179 | n7075 ;
  assign n7078 = ( n2474 & n3882 ) | ( n2474 & ~n4974 ) | ( n3882 & ~n4974 ) ;
  assign n7079 = n346 & n7078 ;
  assign n7080 = n7079 ^ n5434 ^ 1'b0 ;
  assign n7077 = n2578 | n3288 ;
  assign n7081 = n7080 ^ n7077 ^ 1'b0 ;
  assign n7082 = n5647 ^ n4331 ^ n3871 ;
  assign n7083 = n7082 ^ n1146 ^ n947 ;
  assign n7084 = ~n716 & n2801 ;
  assign n7085 = n7084 ^ n2370 ^ 1'b0 ;
  assign n7086 = n7085 ^ n501 ^ 1'b0 ;
  assign n7087 = ~n3697 & n7086 ;
  assign n7088 = n5780 ^ n1942 ^ n509 ;
  assign n7089 = n6658 ^ n4643 ^ n2313 ;
  assign n7090 = ( n1797 & n7088 ) | ( n1797 & ~n7089 ) | ( n7088 & ~n7089 ) ;
  assign n7091 = ( n1886 & ~n4617 ) | ( n1886 & n7090 ) | ( ~n4617 & n7090 ) ;
  assign n7092 = n383 & n1620 ;
  assign n7093 = ( ~n1901 & n2699 ) | ( ~n1901 & n7092 ) | ( n2699 & n7092 ) ;
  assign n7094 = ( n2839 & ~n3971 ) | ( n2839 & n7093 ) | ( ~n3971 & n7093 ) ;
  assign n7099 = ~n1189 & n6715 ;
  assign n7100 = n7099 ^ n1128 ^ 1'b0 ;
  assign n7095 = n6053 ^ n1806 ^ n1384 ;
  assign n7096 = n7095 ^ n3896 ^ 1'b0 ;
  assign n7097 = n7096 ^ n1603 ^ x26 ;
  assign n7098 = n7097 ^ n2397 ^ n532 ;
  assign n7101 = n7100 ^ n7098 ^ n4118 ;
  assign n7105 = n6001 ^ n1761 ^ 1'b0 ;
  assign n7106 = x35 & n3389 ;
  assign n7107 = n7105 & n7106 ;
  assign n7108 = n7107 ^ n858 ^ 1'b0 ;
  assign n7103 = n4190 & ~n5048 ;
  assign n7104 = ~n1633 & n7103 ;
  assign n7102 = n2147 & n5034 ;
  assign n7109 = n7108 ^ n7104 ^ n7102 ;
  assign n7110 = ~n4876 & n7109 ;
  assign n7111 = n7101 & n7110 ;
  assign n7112 = n1105 ^ n722 ^ 1'b0 ;
  assign n7117 = n4185 ^ n1918 ^ 1'b0 ;
  assign n7114 = n2928 | n3510 ;
  assign n7115 = n6700 | n7114 ;
  assign n7116 = n6590 | n7115 ;
  assign n7118 = n7117 ^ n7116 ^ 1'b0 ;
  assign n7119 = n971 | n7118 ;
  assign n7113 = n5353 ^ n1086 ^ n652 ;
  assign n7120 = n7119 ^ n7113 ^ x52 ;
  assign n7124 = ~n297 & n3334 ;
  assign n7121 = n3537 ^ n3249 ^ 1'b0 ;
  assign n7122 = ~n2778 & n7121 ;
  assign n7123 = n7122 ^ n858 ^ n748 ;
  assign n7125 = n7124 ^ n7123 ^ n878 ;
  assign n7126 = ( n1347 & n4098 ) | ( n1347 & ~n7125 ) | ( n4098 & ~n7125 ) ;
  assign n7128 = ( n547 & ~n786 ) | ( n547 & n3316 ) | ( ~n786 & n3316 ) ;
  assign n7129 = n7128 ^ n4176 ^ n1914 ;
  assign n7127 = ( ~n3051 & n4147 ) | ( ~n3051 & n7121 ) | ( n4147 & n7121 ) ;
  assign n7130 = n7129 ^ n7127 ^ n5424 ;
  assign n7131 = x16 & n7130 ;
  assign n7132 = n7131 ^ n1548 ^ 1'b0 ;
  assign n7133 = n853 & n2111 ;
  assign n7134 = n7133 ^ n1324 ^ n731 ;
  assign n7135 = ( ~n909 & n3640 ) | ( ~n909 & n7134 ) | ( n3640 & n7134 ) ;
  assign n7136 = n7135 ^ n4959 ^ 1'b0 ;
  assign n7137 = n5904 | n7136 ;
  assign n7138 = ~n973 & n2807 ;
  assign n7139 = ~n376 & n2134 ;
  assign n7140 = n2555 & n7139 ;
  assign n7141 = ( n1279 & n2921 ) | ( n1279 & ~n7140 ) | ( n2921 & ~n7140 ) ;
  assign n7143 = ( ~n720 & n1561 ) | ( ~n720 & n3784 ) | ( n1561 & n3784 ) ;
  assign n7144 = n7143 ^ n5065 ^ n3298 ;
  assign n7145 = n7144 ^ n2210 ^ 1'b0 ;
  assign n7146 = ~n4127 & n7145 ;
  assign n7142 = ( n1886 & n2905 ) | ( n1886 & n4022 ) | ( n2905 & n4022 ) ;
  assign n7147 = n7146 ^ n7142 ^ n2253 ;
  assign n7148 = n7141 & n7147 ;
  assign n7149 = n7148 ^ n1300 ^ 1'b0 ;
  assign n7150 = n4598 ^ n1933 ^ n978 ;
  assign n7151 = n7150 ^ n5409 ^ n381 ;
  assign n7152 = n7151 ^ n2089 ^ x122 ;
  assign n7153 = n1597 ^ n511 ^ 1'b0 ;
  assign n7154 = n3934 & n7153 ;
  assign n7155 = n7154 ^ n4249 ^ x11 ;
  assign n7156 = n7155 ^ n5865 ^ n692 ;
  assign n7157 = ( n6915 & n7152 ) | ( n6915 & ~n7156 ) | ( n7152 & ~n7156 ) ;
  assign n7158 = n1159 | n2349 ;
  assign n7159 = n7158 ^ n2443 ^ 1'b0 ;
  assign n7160 = n1380 | n7159 ;
  assign n7161 = n4240 ^ n2048 ^ n1617 ;
  assign n7162 = n767 & ~n1471 ;
  assign n7163 = n2049 & n7162 ;
  assign n7168 = ~n637 & n6810 ;
  assign n7169 = n1992 & n7168 ;
  assign n7164 = x125 & n3016 ;
  assign n7165 = n811 & n7164 ;
  assign n7166 = n7165 ^ n584 ^ 1'b0 ;
  assign n7167 = ~n2880 & n7166 ;
  assign n7170 = n7169 ^ n7167 ^ 1'b0 ;
  assign n7171 = n7163 | n7170 ;
  assign n7172 = n187 & ~n7171 ;
  assign n7173 = n2203 & n7172 ;
  assign n7174 = n7173 ^ n696 ^ 1'b0 ;
  assign n7175 = n7161 | n7174 ;
  assign n7176 = n3944 ^ n2760 ^ n2179 ;
  assign n7177 = ( n329 & n1855 ) | ( n329 & n3318 ) | ( n1855 & n3318 ) ;
  assign n7178 = ~x23 & n7177 ;
  assign n7179 = n1053 & n6016 ;
  assign n7180 = n443 & n7179 ;
  assign n7181 = n2590 & ~n7180 ;
  assign n7182 = n7181 ^ n7012 ^ 1'b0 ;
  assign n7183 = ~n2091 & n2606 ;
  assign n7184 = ( ~n3679 & n5341 ) | ( ~n3679 & n6541 ) | ( n5341 & n6541 ) ;
  assign n7185 = ( n1498 & ~n7183 ) | ( n1498 & n7184 ) | ( ~n7183 & n7184 ) ;
  assign n7186 = n1559 & n2410 ;
  assign n7187 = n7186 ^ n3247 ^ 1'b0 ;
  assign n7188 = x8 & n412 ;
  assign n7189 = n1082 & n7188 ;
  assign n7190 = n7187 & n7189 ;
  assign n7193 = n6283 & ~n6783 ;
  assign n7191 = n1473 & n2644 ;
  assign n7192 = ~n4302 & n7191 ;
  assign n7194 = n7193 ^ n7192 ^ n315 ;
  assign n7197 = n6326 ^ n4139 ^ n3511 ;
  assign n7195 = ~n1297 & n1803 ;
  assign n7196 = n4384 | n7195 ;
  assign n7198 = n7197 ^ n7196 ^ 1'b0 ;
  assign n7199 = n7198 ^ n5738 ^ n1510 ;
  assign n7200 = n215 & n7199 ;
  assign n7201 = n4369 & n7200 ;
  assign n7202 = n1508 & n1814 ;
  assign n7203 = ( n372 & ~n6139 ) | ( n372 & n7202 ) | ( ~n6139 & n7202 ) ;
  assign n7204 = ~n1694 & n2301 ;
  assign n7205 = n1179 & n7204 ;
  assign n7207 = n4591 ^ n1336 ^ n746 ;
  assign n7208 = n7207 ^ n1500 ^ n562 ;
  assign n7209 = n4826 | n6781 ;
  assign n7210 = n176 | n7209 ;
  assign n7211 = n4353 & n7210 ;
  assign n7212 = ~n7208 & n7211 ;
  assign n7206 = n1550 & n1843 ;
  assign n7213 = n7212 ^ n7206 ^ 1'b0 ;
  assign n7214 = ~n3874 & n7213 ;
  assign n7215 = ~n2539 & n7214 ;
  assign n7216 = ( n350 & n7205 ) | ( n350 & ~n7215 ) | ( n7205 & ~n7215 ) ;
  assign n7217 = n553 | n3406 ;
  assign n7218 = n180 | n7217 ;
  assign n7219 = n7177 | n7218 ;
  assign n7220 = n5114 ^ n3026 ^ 1'b0 ;
  assign n7221 = n7219 & ~n7220 ;
  assign n7222 = n7221 ^ n5081 ^ 1'b0 ;
  assign n7227 = n2698 ^ n2213 ^ 1'b0 ;
  assign n7228 = n934 & ~n2889 ;
  assign n7229 = ( n2908 & n7227 ) | ( n2908 & ~n7228 ) | ( n7227 & ~n7228 ) ;
  assign n7224 = ( n1287 & n3374 ) | ( n1287 & n3640 ) | ( n3374 & n3640 ) ;
  assign n7225 = ( n2398 & n6845 ) | ( n2398 & ~n7224 ) | ( n6845 & ~n7224 ) ;
  assign n7223 = ( n1763 & ~n3457 ) | ( n1763 & n4679 ) | ( ~n3457 & n4679 ) ;
  assign n7226 = n7225 ^ n7223 ^ n3716 ;
  assign n7230 = n7229 ^ n7226 ^ 1'b0 ;
  assign n7232 = n1086 ^ n366 ^ 1'b0 ;
  assign n7231 = ~n2820 & n4851 ;
  assign n7233 = n7232 ^ n7231 ^ n362 ;
  assign n7234 = ( n1330 & n3272 ) | ( n1330 & ~n6864 ) | ( n3272 & ~n6864 ) ;
  assign n7235 = n2592 & ~n3850 ;
  assign n7236 = n7235 ^ n2941 ^ n2607 ;
  assign n7237 = ( ~n4729 & n5837 ) | ( ~n4729 & n7236 ) | ( n5837 & n7236 ) ;
  assign n7238 = n7237 ^ n5340 ^ n3761 ;
  assign n7239 = n7177 ^ x60 ^ 1'b0 ;
  assign n7240 = n6480 ^ n4726 ^ n1806 ;
  assign n7241 = n7240 ^ n6359 ^ n4443 ;
  assign n7242 = n7241 ^ n3261 ^ 1'b0 ;
  assign n7243 = n7239 & ~n7242 ;
  assign n7244 = n3993 ^ n1144 ^ n464 ;
  assign n7245 = n2027 | n6092 ;
  assign n7246 = n7245 ^ n4640 ^ 1'b0 ;
  assign n7247 = n7244 & ~n7246 ;
  assign n7248 = ~n2838 & n7247 ;
  assign n7249 = n7248 ^ n7123 ^ 1'b0 ;
  assign n7250 = ~n765 & n3605 ;
  assign n7258 = n200 & ~n719 ;
  assign n7259 = n7258 ^ n1654 ^ 1'b0 ;
  assign n7254 = n6368 ^ n2595 ^ n1105 ;
  assign n7255 = n3459 ^ n1382 ^ 1'b0 ;
  assign n7256 = n7254 & ~n7255 ;
  assign n7251 = n3148 ^ n1414 ^ 1'b0 ;
  assign n7252 = ~n1439 & n7251 ;
  assign n7253 = ~n1548 & n7252 ;
  assign n7257 = n7256 ^ n7253 ^ 1'b0 ;
  assign n7260 = n7259 ^ n7257 ^ n373 ;
  assign n7261 = n2390 & ~n6423 ;
  assign n7262 = n2291 & n7261 ;
  assign n7263 = n7260 | n7262 ;
  assign n7264 = n2809 ^ x48 ^ 1'b0 ;
  assign n7265 = ~n975 & n7264 ;
  assign n7266 = ( n806 & n7163 ) | ( n806 & n7265 ) | ( n7163 & n7265 ) ;
  assign n7267 = ~n1210 & n7266 ;
  assign n7268 = n7267 ^ n287 ^ 1'b0 ;
  assign n7269 = n2086 | n7268 ;
  assign n7270 = n7263 & ~n7269 ;
  assign n7271 = n7250 & ~n7270 ;
  assign n7272 = n4120 ^ n1793 ^ n1346 ;
  assign n7273 = ( n849 & ~n2443 ) | ( n849 & n7272 ) | ( ~n2443 & n7272 ) ;
  assign n7274 = ~n3082 & n4356 ;
  assign n7275 = n2832 ^ n1170 ^ n374 ;
  assign n7276 = ( ~x56 & n629 ) | ( ~x56 & n7275 ) | ( n629 & n7275 ) ;
  assign n7277 = n7276 ^ n1024 ^ n383 ;
  assign n7278 = n2094 & n7277 ;
  assign n7279 = ~n7274 & n7278 ;
  assign n7280 = n7279 ^ n315 ^ 1'b0 ;
  assign n7281 = n7273 & n7280 ;
  assign n7282 = ( n1308 & ~n4175 ) | ( n1308 & n4295 ) | ( ~n4175 & n4295 ) ;
  assign n7283 = n3197 ^ n356 ^ x29 ;
  assign n7284 = n7283 ^ n3917 ^ 1'b0 ;
  assign n7285 = n7282 | n7284 ;
  assign n7286 = n1536 & ~n6060 ;
  assign n7287 = n1681 & ~n4086 ;
  assign n7288 = ~n5975 & n7287 ;
  assign n7289 = n7288 ^ n4399 ^ n1299 ;
  assign n7290 = n461 & ~n3719 ;
  assign n7291 = ( n5306 & ~n7289 ) | ( n5306 & n7290 ) | ( ~n7289 & n7290 ) ;
  assign n7292 = n6810 ^ n2321 ^ n2165 ;
  assign n7293 = ~n1510 & n7292 ;
  assign n7294 = n2602 ^ n1964 ^ 1'b0 ;
  assign n7295 = n1049 & ~n1552 ;
  assign n7296 = ~n6223 & n7295 ;
  assign n7297 = n2167 | n6524 ;
  assign n7298 = n7297 ^ n450 ^ 1'b0 ;
  assign n7299 = n2847 ^ n1246 ^ x53 ;
  assign n7300 = n7299 ^ n2078 ^ n1306 ;
  assign n7301 = n3785 ^ n1504 ^ 1'b0 ;
  assign n7302 = n2381 & n7301 ;
  assign n7304 = n1919 ^ n1076 ^ n954 ;
  assign n7303 = n4320 & ~n5589 ;
  assign n7305 = n7304 ^ n7303 ^ 1'b0 ;
  assign n7306 = ( n5483 & ~n7302 ) | ( n5483 & n7305 ) | ( ~n7302 & n7305 ) ;
  assign n7307 = n3261 ^ n3074 ^ n2050 ;
  assign n7308 = n7307 ^ n2844 ^ 1'b0 ;
  assign n7309 = n7308 ^ n2169 ^ n876 ;
  assign n7323 = n6295 ^ n2219 ^ n236 ;
  assign n7320 = ( n309 & ~n570 ) | ( n309 & n3581 ) | ( ~n570 & n3581 ) ;
  assign n7321 = n5277 ^ n2058 ^ 1'b0 ;
  assign n7322 = n7320 | n7321 ;
  assign n7324 = n7323 ^ n7322 ^ n5645 ;
  assign n7325 = n7324 ^ n7195 ^ n3723 ;
  assign n7316 = n2147 ^ n748 ^ 1'b0 ;
  assign n7317 = n2292 & ~n7316 ;
  assign n7318 = ~n4993 & n7317 ;
  assign n7319 = ( n4560 & n5088 ) | ( n4560 & n7318 ) | ( n5088 & n7318 ) ;
  assign n7313 = ~n1038 & n1989 ;
  assign n7314 = ~n733 & n7313 ;
  assign n7310 = n819 & ~n910 ;
  assign n7311 = n7310 ^ x1 ^ 1'b0 ;
  assign n7312 = n597 & ~n7311 ;
  assign n7315 = n7314 ^ n7312 ^ 1'b0 ;
  assign n7326 = n7325 ^ n7319 ^ n7315 ;
  assign n7327 = n6670 ^ n5242 ^ 1'b0 ;
  assign n7328 = ~n2608 & n6592 ;
  assign n7329 = n4102 ^ n2422 ^ n1641 ;
  assign n7330 = n7329 ^ n2877 ^ 1'b0 ;
  assign n7331 = ~n7328 & n7330 ;
  assign n7332 = n7331 ^ n3462 ^ n1010 ;
  assign n7333 = n4672 ^ n619 ^ n383 ;
  assign n7334 = n6383 ^ n4181 ^ n1316 ;
  assign n7335 = ~n2805 & n5244 ;
  assign n7336 = n7335 ^ n2026 ^ 1'b0 ;
  assign n7337 = n4498 ^ n4141 ^ n1709 ;
  assign n7338 = ~n2046 & n2761 ;
  assign n7339 = n7337 & n7338 ;
  assign n7340 = n4650 ^ n4513 ^ n4034 ;
  assign n7341 = n2721 ^ n1099 ^ 1'b0 ;
  assign n7342 = n4969 | n7341 ;
  assign n7343 = n4247 ^ n1571 ^ n1061 ;
  assign n7344 = ( n1243 & n5295 ) | ( n1243 & n7343 ) | ( n5295 & n7343 ) ;
  assign n7345 = ( n7340 & ~n7342 ) | ( n7340 & n7344 ) | ( ~n7342 & n7344 ) ;
  assign n7347 = n2195 ^ n1264 ^ n759 ;
  assign n7348 = ~n1205 & n7347 ;
  assign n7349 = n7062 | n7348 ;
  assign n7346 = ~n131 & n1933 ;
  assign n7350 = n7349 ^ n7346 ^ 1'b0 ;
  assign n7355 = x93 & ~n429 ;
  assign n7356 = ~n1373 & n7355 ;
  assign n7357 = x40 & ~n1534 ;
  assign n7358 = n7357 ^ n364 ^ 1'b0 ;
  assign n7359 = ( x2 & n7356 ) | ( x2 & n7358 ) | ( n7356 & n7358 ) ;
  assign n7360 = n1875 & n7359 ;
  assign n7361 = ( x43 & n3336 ) | ( x43 & n7360 ) | ( n3336 & n7360 ) ;
  assign n7351 = n6397 ^ n1708 ^ n863 ;
  assign n7352 = n7351 ^ n4986 ^ n3546 ;
  assign n7353 = n7352 ^ n6413 ^ x123 ;
  assign n7354 = n4280 & ~n7353 ;
  assign n7362 = n7361 ^ n7354 ^ 1'b0 ;
  assign n7363 = ~n2490 & n4260 ;
  assign n7366 = n2475 & n2892 ;
  assign n7364 = ~n2284 & n6406 ;
  assign n7365 = ~n1525 & n7364 ;
  assign n7367 = n7366 ^ n7365 ^ n2511 ;
  assign n7368 = n7367 ^ n1732 ^ 1'b0 ;
  assign n7369 = ( n1141 & ~n3700 ) | ( n1141 & n3816 ) | ( ~n3700 & n3816 ) ;
  assign n7370 = n7369 ^ n3536 ^ n2998 ;
  assign n7371 = ( n1044 & n2542 ) | ( n1044 & n2903 ) | ( n2542 & n2903 ) ;
  assign n7372 = n5559 & ~n7371 ;
  assign n7373 = n7372 ^ n505 ^ 1'b0 ;
  assign n7374 = ~n4747 & n7373 ;
  assign n7375 = n4363 & ~n6067 ;
  assign n7376 = n138 | n1750 ;
  assign n7377 = n7376 ^ n461 ^ 1'b0 ;
  assign n7378 = n7377 ^ n6919 ^ n1713 ;
  assign n7379 = n2636 ^ n2067 ^ n1648 ;
  assign n7380 = ~n6564 & n7379 ;
  assign n7381 = ( n786 & n2456 ) | ( n786 & ~n3856 ) | ( n2456 & ~n3856 ) ;
  assign n7382 = n5851 ^ n3888 ^ 1'b0 ;
  assign n7383 = n7382 ^ n4759 ^ n1311 ;
  assign n7384 = n7381 & ~n7383 ;
  assign n7385 = n7384 ^ n227 ^ 1'b0 ;
  assign n7386 = ~n5393 & n7124 ;
  assign n7387 = n1336 & ~n3645 ;
  assign n7388 = n2694 & n7387 ;
  assign n7389 = n7388 ^ n6731 ^ n5689 ;
  assign n7390 = ~n130 & n1819 ;
  assign n7391 = ~n7389 & n7390 ;
  assign n7392 = n2260 & n3858 ;
  assign n7402 = n1919 ^ n1644 ^ 1'b0 ;
  assign n7399 = n3967 ^ n2424 ^ n1088 ;
  assign n7400 = n7399 ^ n1270 ^ 1'b0 ;
  assign n7401 = ~n2470 & n7400 ;
  assign n7396 = n4519 ^ n2093 ^ n716 ;
  assign n7397 = ( n1528 & n3443 ) | ( n1528 & n7396 ) | ( n3443 & n7396 ) ;
  assign n7395 = n1175 & ~n2417 ;
  assign n7398 = n7397 ^ n7395 ^ 1'b0 ;
  assign n7403 = n7402 ^ n7401 ^ n7398 ;
  assign n7393 = n4985 ^ n1871 ^ 1'b0 ;
  assign n7394 = n6392 & n7393 ;
  assign n7404 = n7403 ^ n7394 ^ 1'b0 ;
  assign n7405 = n5065 ^ n2477 ^ 1'b0 ;
  assign n7406 = ~n5058 & n6795 ;
  assign n7407 = ( n2290 & n7405 ) | ( n2290 & n7406 ) | ( n7405 & n7406 ) ;
  assign n7408 = n2418 & ~n7407 ;
  assign n7409 = ~n308 & n5234 ;
  assign n7410 = n6397 & n7409 ;
  assign n7411 = ( n2381 & n7408 ) | ( n2381 & n7410 ) | ( n7408 & n7410 ) ;
  assign n7412 = ( n1694 & n3115 ) | ( n1694 & n7411 ) | ( n3115 & n7411 ) ;
  assign n7413 = n3686 ^ x105 ^ 1'b0 ;
  assign n7414 = n4793 & ~n7413 ;
  assign n7415 = ( n1629 & n5983 ) | ( n1629 & n7414 ) | ( n5983 & n7414 ) ;
  assign n7416 = n3285 & n7415 ;
  assign n7417 = ( n1805 & n4924 ) | ( n1805 & n5118 ) | ( n4924 & n5118 ) ;
  assign n7418 = ( n929 & ~n1275 ) | ( n929 & n7219 ) | ( ~n1275 & n7219 ) ;
  assign n7419 = ( ~n1896 & n3354 ) | ( ~n1896 & n7151 ) | ( n3354 & n7151 ) ;
  assign n7420 = ( ~n541 & n1465 ) | ( ~n541 & n2725 ) | ( n1465 & n2725 ) ;
  assign n7421 = n1388 & n7420 ;
  assign n7422 = ( ~n3770 & n4747 ) | ( ~n3770 & n5431 ) | ( n4747 & n5431 ) ;
  assign n7423 = ~n7421 & n7422 ;
  assign n7427 = ( n178 & ~n2229 ) | ( n178 & n4051 ) | ( ~n2229 & n4051 ) ;
  assign n7425 = ( n409 & n3457 ) | ( n409 & n3482 ) | ( n3457 & n3482 ) ;
  assign n7424 = x94 & n170 ;
  assign n7426 = n7425 ^ n7424 ^ n5331 ;
  assign n7428 = n7427 ^ n7426 ^ n4240 ;
  assign n7429 = ~n142 & n492 ;
  assign n7430 = n1791 & n7429 ;
  assign n7431 = n7430 ^ n1091 ^ 1'b0 ;
  assign n7435 = n5961 ^ n958 ^ 1'b0 ;
  assign n7432 = n2644 & n3963 ;
  assign n7433 = n7432 ^ n2014 ^ 1'b0 ;
  assign n7434 = n1468 | n7433 ;
  assign n7436 = n7435 ^ n7434 ^ n949 ;
  assign n7443 = ~n1142 & n1795 ;
  assign n7444 = n2488 & n7443 ;
  assign n7445 = n6308 & ~n7444 ;
  assign n7446 = n7445 ^ n6268 ^ 1'b0 ;
  assign n7437 = n1394 | n1834 ;
  assign n7438 = n7437 ^ n6220 ^ n1859 ;
  assign n7439 = n1623 & ~n4491 ;
  assign n7440 = ~n7438 & n7439 ;
  assign n7441 = n872 | n7440 ;
  assign n7442 = ~n2918 & n7441 ;
  assign n7447 = n7446 ^ n7442 ^ 1'b0 ;
  assign n7448 = x79 | n3935 ;
  assign n7449 = ~n849 & n7448 ;
  assign n7450 = ~n370 & n7449 ;
  assign n7455 = n6480 ^ n2114 ^ 1'b0 ;
  assign n7456 = ~n5328 & n7455 ;
  assign n7451 = n3625 & n4599 ;
  assign n7452 = n1541 & n7451 ;
  assign n7453 = n2313 & ~n5070 ;
  assign n7454 = n7452 & n7453 ;
  assign n7457 = n7456 ^ n7454 ^ 1'b0 ;
  assign n7458 = n7450 | n7457 ;
  assign n7459 = n7458 ^ n5806 ^ n2426 ;
  assign n7460 = n3904 | n6081 ;
  assign n7468 = ( n803 & n2914 ) | ( n803 & ~n3645 ) | ( n2914 & ~n3645 ) ;
  assign n7462 = ~n459 & n6970 ;
  assign n7463 = n131 & n7462 ;
  assign n7464 = n6649 ^ n2321 ^ 1'b0 ;
  assign n7465 = ~n171 & n7464 ;
  assign n7466 = ~n7463 & n7465 ;
  assign n7467 = ~n4559 & n7466 ;
  assign n7469 = n7468 ^ n7467 ^ n4036 ;
  assign n7461 = ~n2488 & n3588 ;
  assign n7470 = n7469 ^ n7461 ^ 1'b0 ;
  assign n7473 = n1234 ^ n929 ^ x53 ;
  assign n7471 = n2886 & n6793 ;
  assign n7472 = n7471 ^ n5081 ^ 1'b0 ;
  assign n7474 = n7473 ^ n7472 ^ 1'b0 ;
  assign n7475 = n2999 & ~n7474 ;
  assign n7476 = n227 | n4788 ;
  assign n7477 = n2697 & ~n7476 ;
  assign n7478 = ( n1427 & ~n6008 ) | ( n1427 & n7477 ) | ( ~n6008 & n7477 ) ;
  assign n7487 = n1881 & n3899 ;
  assign n7488 = ~n626 & n7487 ;
  assign n7489 = n3316 | n7488 ;
  assign n7490 = n4350 & ~n7489 ;
  assign n7482 = ( n181 & n1675 ) | ( n181 & ~n3113 ) | ( n1675 & ~n3113 ) ;
  assign n7483 = n3703 | n7482 ;
  assign n7484 = n4593 | n7483 ;
  assign n7485 = n1894 | n7484 ;
  assign n7479 = ( ~n2560 & n4510 ) | ( ~n2560 & n5891 ) | ( n4510 & n5891 ) ;
  assign n7480 = ~n5436 & n7479 ;
  assign n7481 = n4715 & n7480 ;
  assign n7486 = n7485 ^ n7481 ^ 1'b0 ;
  assign n7491 = n7490 ^ n7486 ^ 1'b0 ;
  assign n7492 = n7478 & n7491 ;
  assign n7493 = ~n145 & n3364 ;
  assign n7494 = n5714 & ~n7493 ;
  assign n7495 = n7494 ^ n3349 ^ 1'b0 ;
  assign n7496 = ( n334 & n2803 ) | ( n334 & n5955 ) | ( n2803 & n5955 ) ;
  assign n7497 = n7244 ^ n3140 ^ n896 ;
  assign n7498 = n550 & n4460 ;
  assign n7499 = n7498 ^ n2272 ^ 1'b0 ;
  assign n7500 = n4482 | n7499 ;
  assign n7501 = n4230 & ~n7500 ;
  assign n7502 = ~n7222 & n7501 ;
  assign n7503 = n4786 & n7067 ;
  assign n7504 = ~n1513 & n7183 ;
  assign n7505 = n326 | n1082 ;
  assign n7506 = n7505 ^ n4220 ^ 1'b0 ;
  assign n7507 = n4030 ^ n2210 ^ n964 ;
  assign n7508 = ~n2598 & n4072 ;
  assign n7509 = n7507 & n7508 ;
  assign n7510 = ~n6489 & n7509 ;
  assign n7511 = ~n1873 & n7274 ;
  assign n7512 = n7511 ^ n3848 ^ n2534 ;
  assign n7513 = n3385 & n7512 ;
  assign n7514 = x87 & ~n1141 ;
  assign n7515 = n250 & n7514 ;
  assign n7516 = x9 & ~n2962 ;
  assign n7517 = n1210 & n7516 ;
  assign n7518 = ~n3028 & n3147 ;
  assign n7519 = n7518 ^ n7193 ^ n2830 ;
  assign n7520 = n759 & n7519 ;
  assign n7521 = n7520 ^ n7222 ^ 1'b0 ;
  assign n7522 = n7517 | n7521 ;
  assign n7523 = n5949 ^ n5060 ^ n3784 ;
  assign n7524 = n903 & ~n7523 ;
  assign n7525 = ( n294 & n1767 ) | ( n294 & ~n7199 ) | ( n1767 & ~n7199 ) ;
  assign n7526 = n2050 ^ n1349 ^ n418 ;
  assign n7527 = n7526 ^ n4581 ^ n256 ;
  assign n7528 = ( n1496 & n3062 ) | ( n1496 & n6568 ) | ( n3062 & n6568 ) ;
  assign n7529 = n7528 ^ n6057 ^ 1'b0 ;
  assign n7530 = ( n4451 & ~n6283 ) | ( n4451 & n7146 ) | ( ~n6283 & n7146 ) ;
  assign n7531 = ( n6368 & n7529 ) | ( n6368 & n7530 ) | ( n7529 & n7530 ) ;
  assign n7532 = n3541 | n7236 ;
  assign n7533 = n7532 ^ n646 ^ 1'b0 ;
  assign n7534 = ~n1107 & n5595 ;
  assign n7535 = ~n1015 & n7534 ;
  assign n7536 = n1285 & ~n3249 ;
  assign n7537 = n7536 ^ n492 ^ 1'b0 ;
  assign n7538 = n7535 | n7537 ;
  assign n7540 = ~n4393 & n6437 ;
  assign n7541 = n7540 ^ n6098 ^ 1'b0 ;
  assign n7542 = n7541 ^ n3109 ^ n1163 ;
  assign n7543 = n6200 | n7542 ;
  assign n7544 = n7543 ^ n4842 ^ 1'b0 ;
  assign n7539 = ~n2207 & n7407 ;
  assign n7545 = n7544 ^ n7539 ^ n3079 ;
  assign n7546 = n3483 ^ n1802 ^ n1088 ;
  assign n7547 = ~n698 & n7546 ;
  assign n7548 = ~n2700 & n7547 ;
  assign n7549 = n3061 ^ n2326 ^ x4 ;
  assign n7550 = ( ~n2583 & n4049 ) | ( ~n2583 & n7549 ) | ( n4049 & n7549 ) ;
  assign n7551 = ( n481 & n5617 ) | ( n481 & ~n7550 ) | ( n5617 & ~n7550 ) ;
  assign n7552 = ( n1817 & n7548 ) | ( n1817 & ~n7551 ) | ( n7548 & ~n7551 ) ;
  assign n7555 = n1477 | n3076 ;
  assign n7556 = n7165 | n7555 ;
  assign n7557 = n5779 & ~n7556 ;
  assign n7553 = n1809 ^ n601 ^ 1'b0 ;
  assign n7554 = ( ~n1698 & n4106 ) | ( ~n1698 & n7553 ) | ( n4106 & n7553 ) ;
  assign n7558 = n7557 ^ n7554 ^ n5843 ;
  assign n7559 = n2245 ^ n1956 ^ 1'b0 ;
  assign n7560 = n4671 & n7559 ;
  assign n7561 = x31 & ~n5210 ;
  assign n7562 = n7561 ^ n2738 ^ 1'b0 ;
  assign n7563 = n1592 & n3305 ;
  assign n7564 = ( ~n252 & n7562 ) | ( ~n252 & n7563 ) | ( n7562 & n7563 ) ;
  assign n7565 = n2904 ^ n512 ^ 1'b0 ;
  assign n7566 = ~n7564 & n7565 ;
  assign n7567 = n374 & n706 ;
  assign n7568 = n7567 ^ n1306 ^ 1'b0 ;
  assign n7569 = n7568 ^ n6439 ^ 1'b0 ;
  assign n7570 = n7566 & n7569 ;
  assign n7571 = n3295 ^ n2777 ^ 1'b0 ;
  assign n7572 = ( ~n2877 & n3016 ) | ( ~n2877 & n7571 ) | ( n3016 & n7571 ) ;
  assign n7585 = ~n680 & n3558 ;
  assign n7584 = ( n4098 & n6429 ) | ( n4098 & ~n7151 ) | ( n6429 & ~n7151 ) ;
  assign n7580 = n2519 & n6778 ;
  assign n7573 = n2209 ^ n918 ^ 1'b0 ;
  assign n7574 = n332 | n7573 ;
  assign n7575 = n4311 ^ n2209 ^ n1288 ;
  assign n7576 = n2358 & n7575 ;
  assign n7577 = n7574 & n7576 ;
  assign n7578 = ( ~n293 & n2420 ) | ( ~n293 & n7245 ) | ( n2420 & n7245 ) ;
  assign n7579 = n7577 | n7578 ;
  assign n7581 = n7580 ^ n7579 ^ 1'b0 ;
  assign n7582 = n2862 | n6098 ;
  assign n7583 = ( ~n5811 & n7581 ) | ( ~n5811 & n7582 ) | ( n7581 & n7582 ) ;
  assign n7586 = n7585 ^ n7584 ^ n7583 ;
  assign n7587 = ( n2247 & ~n7572 ) | ( n2247 & n7586 ) | ( ~n7572 & n7586 ) ;
  assign n7588 = n5822 ^ n5249 ^ n3115 ;
  assign n7589 = n5230 | n5368 ;
  assign n7590 = n7588 & n7589 ;
  assign n7591 = n7001 ^ n5672 ^ n1665 ;
  assign n7592 = n7591 ^ n6945 ^ n3791 ;
  assign n7593 = n5978 ^ n1606 ^ 1'b0 ;
  assign n7594 = ~n4793 & n7593 ;
  assign n7595 = n1529 & ~n2234 ;
  assign n7596 = n7595 ^ n1217 ^ 1'b0 ;
  assign n7597 = n7596 ^ n1387 ^ 1'b0 ;
  assign n7598 = ( x2 & n1477 ) | ( x2 & n7597 ) | ( n1477 & n7597 ) ;
  assign n7599 = ( n5419 & n6303 ) | ( n5419 & n7598 ) | ( n6303 & n7598 ) ;
  assign n7600 = n156 & ~n1234 ;
  assign n7601 = ( n1227 & n1901 ) | ( n1227 & ~n7600 ) | ( n1901 & ~n7600 ) ;
  assign n7602 = x52 & ~n895 ;
  assign n7603 = n3354 | n7602 ;
  assign n7604 = ( ~n447 & n7601 ) | ( ~n447 & n7603 ) | ( n7601 & n7603 ) ;
  assign n7605 = n7604 ^ n4604 ^ n2667 ;
  assign n7606 = ( n1684 & ~n2921 ) | ( n1684 & n4689 ) | ( ~n2921 & n4689 ) ;
  assign n7607 = n7606 ^ n1624 ^ n1357 ;
  assign n7608 = n5918 ^ n2553 ^ n1953 ;
  assign n7609 = n6458 & ~n7608 ;
  assign n7610 = n532 & ~n3022 ;
  assign n7611 = n3062 & n7610 ;
  assign n7612 = x23 & n824 ;
  assign n7613 = n7612 ^ n4589 ^ 1'b0 ;
  assign n7614 = n7613 ^ n2588 ^ n1277 ;
  assign n7615 = ( n1281 & ~n7611 ) | ( n1281 & n7614 ) | ( ~n7611 & n7614 ) ;
  assign n7616 = ~n387 & n7615 ;
  assign n7617 = n1679 & ~n4089 ;
  assign n7618 = ~n7616 & n7617 ;
  assign n7619 = n5610 ^ n2837 ^ n134 ;
  assign n7620 = n2414 ^ n1190 ^ 1'b0 ;
  assign n7621 = ~n3171 & n3841 ;
  assign n7622 = ~n7620 & n7621 ;
  assign n7623 = n7622 ^ n3896 ^ 1'b0 ;
  assign n7624 = n7619 & n7623 ;
  assign n7635 = n5411 ^ n2026 ^ 1'b0 ;
  assign n7636 = n2738 & n5558 ;
  assign n7637 = n7635 & n7636 ;
  assign n7625 = n1728 | n2143 ;
  assign n7626 = n7625 ^ n1310 ^ 1'b0 ;
  assign n7627 = n7626 ^ n3081 ^ n2335 ;
  assign n7628 = ( ~n1323 & n6261 ) | ( ~n1323 & n7627 ) | ( n6261 & n7627 ) ;
  assign n7629 = n3454 & ~n6983 ;
  assign n7630 = ~n1915 & n7629 ;
  assign n7631 = n170 | n7630 ;
  assign n7632 = n2862 & ~n7631 ;
  assign n7633 = ( n1583 & ~n7628 ) | ( n1583 & n7632 ) | ( ~n7628 & n7632 ) ;
  assign n7634 = ( n677 & n5818 ) | ( n677 & n7633 ) | ( n5818 & n7633 ) ;
  assign n7638 = n7637 ^ n7634 ^ 1'b0 ;
  assign n7644 = n7399 ^ n4176 ^ x11 ;
  assign n7639 = n3734 ^ n3016 ^ x88 ;
  assign n7640 = ~n3814 & n7639 ;
  assign n7641 = n1148 & n2343 ;
  assign n7642 = n1872 & ~n7641 ;
  assign n7643 = ( n4560 & n7640 ) | ( n4560 & ~n7642 ) | ( n7640 & ~n7642 ) ;
  assign n7645 = n7644 ^ n7643 ^ n7399 ;
  assign n7646 = n5922 ^ n2259 ^ 1'b0 ;
  assign n7647 = n2251 | n7646 ;
  assign n7648 = ~n2089 & n3273 ;
  assign n7650 = n3546 | n3704 ;
  assign n7651 = n7450 & ~n7650 ;
  assign n7649 = x18 & ~n6506 ;
  assign n7652 = n7651 ^ n7649 ^ 1'b0 ;
  assign n7653 = n7648 & ~n7652 ;
  assign n7654 = ( n937 & ~n2770 ) | ( n937 & n6690 ) | ( ~n2770 & n6690 ) ;
  assign n7655 = n4837 ^ n3789 ^ 1'b0 ;
  assign n7656 = n2002 & n7655 ;
  assign n7657 = ~n7654 & n7656 ;
  assign n7658 = ( x101 & n1108 ) | ( x101 & n1903 ) | ( n1108 & n1903 ) ;
  assign n7659 = n7658 ^ n1004 ^ 1'b0 ;
  assign n7660 = n2575 & ~n7659 ;
  assign n7661 = ( n4560 & n4910 ) | ( n4560 & ~n7660 ) | ( n4910 & ~n7660 ) ;
  assign n7662 = n972 & n1041 ;
  assign n7663 = n7662 ^ n1659 ^ 1'b0 ;
  assign n7664 = n7661 & ~n7663 ;
  assign n7665 = ( n1986 & ~n6243 ) | ( n1986 & n7307 ) | ( ~n6243 & n7307 ) ;
  assign n7666 = n4888 ^ n2175 ^ 1'b0 ;
  assign n7667 = n1403 & n7666 ;
  assign n7668 = n5118 & n7667 ;
  assign n7669 = ~n652 & n6919 ;
  assign n7670 = ( ~n4341 & n6668 ) | ( ~n4341 & n7240 ) | ( n6668 & n7240 ) ;
  assign n7671 = ( n2464 & ~n3300 ) | ( n2464 & n5575 ) | ( ~n3300 & n5575 ) ;
  assign n7672 = n6640 ^ n6131 ^ 1'b0 ;
  assign n7673 = n7671 | n7672 ;
  assign n7679 = n2608 ^ n696 ^ 1'b0 ;
  assign n7680 = n738 ^ n334 ^ 1'b0 ;
  assign n7681 = ( n3826 & n7679 ) | ( n3826 & n7680 ) | ( n7679 & n7680 ) ;
  assign n7677 = ( ~x121 & n330 ) | ( ~x121 & n3061 ) | ( n330 & n3061 ) ;
  assign n7674 = ( n182 & ~n3882 ) | ( n182 & n4213 ) | ( ~n3882 & n4213 ) ;
  assign n7675 = n7674 ^ n6398 ^ n474 ;
  assign n7676 = ( n374 & ~n3727 ) | ( n374 & n7675 ) | ( ~n3727 & n7675 ) ;
  assign n7678 = n7677 ^ n7676 ^ 1'b0 ;
  assign n7682 = n7681 ^ n7678 ^ n1820 ;
  assign n7683 = n1748 ^ n529 ^ 1'b0 ;
  assign n7684 = n4506 & ~n7683 ;
  assign n7685 = n1107 | n1904 ;
  assign n7686 = n7684 & n7685 ;
  assign n7687 = n4469 & n7686 ;
  assign n7688 = n1107 & n2371 ;
  assign n7689 = n4432 ^ n844 ^ 1'b0 ;
  assign n7690 = n7689 ^ n3565 ^ 1'b0 ;
  assign n7691 = n7073 ^ n4310 ^ n2894 ;
  assign n7696 = n5262 ^ n3756 ^ n1301 ;
  assign n7693 = ( n659 & n1017 ) | ( n659 & n2422 ) | ( n1017 & n2422 ) ;
  assign n7692 = ( x93 & ~n2477 ) | ( x93 & n5779 ) | ( ~n2477 & n5779 ) ;
  assign n7694 = n7693 ^ n7692 ^ 1'b0 ;
  assign n7695 = n7694 ^ n3602 ^ 1'b0 ;
  assign n7697 = n7696 ^ n7695 ^ n2374 ;
  assign n7698 = ~n7691 & n7697 ;
  assign n7699 = n1082 & n7698 ;
  assign n7700 = ( n4434 & ~n5747 ) | ( n4434 & n7424 ) | ( ~n5747 & n7424 ) ;
  assign n7701 = n7620 & n7700 ;
  assign n7702 = n5598 & n5641 ;
  assign n7703 = n7702 ^ n4862 ^ 1'b0 ;
  assign n7704 = x23 & n7703 ;
  assign n7705 = ~n7701 & n7704 ;
  assign n7706 = n6123 ^ n4407 ^ 1'b0 ;
  assign n7707 = ~n5772 & n7411 ;
  assign n7708 = n7706 & n7707 ;
  assign n7709 = n3608 ^ n1898 ^ 1'b0 ;
  assign n7710 = n1772 | n7709 ;
  assign n7711 = n7710 ^ n4408 ^ 1'b0 ;
  assign n7712 = x58 & ~n7711 ;
  assign n7713 = ~n3137 & n7712 ;
  assign n7714 = ~n1196 & n3934 ;
  assign n7715 = n7714 ^ n6261 ^ x30 ;
  assign n7716 = n7715 ^ n1422 ^ n1206 ;
  assign n7717 = n3229 & n7716 ;
  assign n7718 = n7717 ^ n798 ^ 1'b0 ;
  assign n7719 = n7352 & n7718 ;
  assign n7720 = n6644 ^ n2779 ^ 1'b0 ;
  assign n7730 = n2383 ^ n1107 ^ 1'b0 ;
  assign n7724 = n5685 | n7600 ;
  assign n7725 = ~n3998 & n7724 ;
  assign n7726 = ~n3452 & n7725 ;
  assign n7721 = n2475 | n2648 ;
  assign n7722 = n7721 ^ n5290 ^ 1'b0 ;
  assign n7723 = n664 | n7722 ;
  assign n7727 = n7726 ^ n7723 ^ 1'b0 ;
  assign n7728 = n7727 ^ n1331 ^ 1'b0 ;
  assign n7729 = ~n6214 & n7728 ;
  assign n7731 = n7730 ^ n7729 ^ n1115 ;
  assign n7732 = ( x11 & ~n3674 ) | ( x11 & n4354 ) | ( ~n3674 & n4354 ) ;
  assign n7733 = n4278 & ~n4904 ;
  assign n7734 = n7733 ^ n4696 ^ n1798 ;
  assign n7737 = n4795 ^ n2072 ^ n1649 ;
  assign n7735 = n4040 ^ n2652 ^ n2176 ;
  assign n7736 = n7735 ^ n3668 ^ n1734 ;
  assign n7738 = n7737 ^ n7736 ^ n4412 ;
  assign n7739 = n7734 & n7738 ;
  assign n7740 = ~n3550 & n7739 ;
  assign n7741 = n4341 ^ n2253 ^ 1'b0 ;
  assign n7742 = ( ~n1145 & n5276 ) | ( ~n1145 & n7741 ) | ( n5276 & n7741 ) ;
  assign n7743 = ( n4336 & ~n5810 ) | ( n4336 & n7742 ) | ( ~n5810 & n7742 ) ;
  assign n7744 = ~n300 & n945 ;
  assign n7745 = n4169 ^ n2062 ^ 1'b0 ;
  assign n7746 = n1154 & n7745 ;
  assign n7747 = n7746 ^ n298 ^ 1'b0 ;
  assign n7748 = n7747 ^ n7438 ^ 1'b0 ;
  assign n7749 = ~n5390 & n7748 ;
  assign n7750 = n7749 ^ n697 ^ 1'b0 ;
  assign n7756 = n7680 ^ n3498 ^ 1'b0 ;
  assign n7757 = n2699 & n7756 ;
  assign n7751 = n6516 ^ n3036 ^ 1'b0 ;
  assign n7752 = n4896 & n7751 ;
  assign n7753 = ( n2509 & n3493 ) | ( n2509 & ~n5110 ) | ( n3493 & ~n5110 ) ;
  assign n7754 = ( n931 & n5114 ) | ( n931 & n7753 ) | ( n5114 & n7753 ) ;
  assign n7755 = ( n1153 & n7752 ) | ( n1153 & n7754 ) | ( n7752 & n7754 ) ;
  assign n7758 = n7757 ^ n7755 ^ n6281 ;
  assign n7759 = n4273 ^ n2573 ^ n1876 ;
  assign n7760 = n7759 ^ n3603 ^ n268 ;
  assign n7761 = ~n1184 & n1387 ;
  assign n7762 = n7761 ^ n5961 ^ 1'b0 ;
  assign n7763 = n561 & n607 ;
  assign n7764 = n2550 ^ n1403 ^ x69 ;
  assign n7765 = ( n452 & n1783 ) | ( n452 & ~n6941 ) | ( n1783 & ~n6941 ) ;
  assign n7766 = x111 & n3236 ;
  assign n7767 = n7765 & n7766 ;
  assign n7768 = ~n7764 & n7767 ;
  assign n7773 = x82 & n1005 ;
  assign n7774 = n7773 ^ n2481 ^ 1'b0 ;
  assign n7769 = n2291 ^ n1590 ^ n702 ;
  assign n7770 = n2291 ^ n1331 ^ n537 ;
  assign n7771 = n7770 ^ n6024 ^ n3154 ;
  assign n7772 = ( n6556 & ~n7769 ) | ( n6556 & n7771 ) | ( ~n7769 & n7771 ) ;
  assign n7775 = n7774 ^ n7772 ^ 1'b0 ;
  assign n7776 = ( ~n285 & n2026 ) | ( ~n285 & n4325 ) | ( n2026 & n4325 ) ;
  assign n7777 = ~n7147 & n7765 ;
  assign n7778 = ( n592 & ~n7776 ) | ( n592 & n7777 ) | ( ~n7776 & n7777 ) ;
  assign n7780 = n413 ^ n362 ^ 1'b0 ;
  assign n7781 = ( ~n3813 & n6658 ) | ( ~n3813 & n7780 ) | ( n6658 & n7780 ) ;
  assign n7779 = n1128 | n3674 ;
  assign n7782 = n7781 ^ n7779 ^ 1'b0 ;
  assign n7783 = n7782 ^ n5092 ^ n2588 ;
  assign n7784 = n3347 ^ n775 ^ 1'b0 ;
  assign n7785 = n1756 & ~n7784 ;
  assign n7786 = n1344 & ~n4501 ;
  assign n7787 = n7786 ^ n680 ^ 1'b0 ;
  assign n7788 = n7787 ^ n3991 ^ 1'b0 ;
  assign n7789 = n7785 & n7788 ;
  assign n7790 = ( n2699 & ~n2991 ) | ( n2699 & n4456 ) | ( ~n2991 & n4456 ) ;
  assign n7791 = ( n1507 & n6128 ) | ( n1507 & ~n7790 ) | ( n6128 & ~n7790 ) ;
  assign n7792 = ( ~n421 & n6260 ) | ( ~n421 & n6870 ) | ( n6260 & n6870 ) ;
  assign n7793 = n7792 ^ n4087 ^ n2682 ;
  assign n7794 = ( n4350 & n7791 ) | ( n4350 & ~n7793 ) | ( n7791 & ~n7793 ) ;
  assign n7795 = ( n7783 & ~n7789 ) | ( n7783 & n7794 ) | ( ~n7789 & n7794 ) ;
  assign n7796 = n7194 ^ n5514 ^ 1'b0 ;
  assign n7797 = n886 & n7796 ;
  assign n7799 = n1126 & n3305 ;
  assign n7800 = n7799 ^ n3336 ^ 1'b0 ;
  assign n7798 = ( ~x21 & n559 ) | ( ~x21 & n5189 ) | ( n559 & n5189 ) ;
  assign n7801 = n7800 ^ n7798 ^ 1'b0 ;
  assign n7802 = ~n5653 & n7801 ;
  assign n7804 = n624 & n629 ;
  assign n7805 = n7804 ^ n2738 ^ 1'b0 ;
  assign n7803 = n1401 | n7793 ;
  assign n7806 = n7805 ^ n7803 ^ 1'b0 ;
  assign n7809 = n1186 & n1406 ;
  assign n7810 = n7809 ^ n5562 ^ 1'b0 ;
  assign n7811 = ~n540 & n7810 ;
  assign n7812 = ~n1097 & n7811 ;
  assign n7807 = n6693 ^ n4677 ^ 1'b0 ;
  assign n7808 = n4959 | n7807 ;
  assign n7813 = n7812 ^ n7808 ^ x32 ;
  assign n7824 = n1623 & ~n4066 ;
  assign n7825 = n7824 ^ n4306 ^ 1'b0 ;
  assign n7823 = n4249 ^ n3031 ^ n788 ;
  assign n7815 = ( x38 & n743 ) | ( x38 & ~n1439 ) | ( n743 & ~n1439 ) ;
  assign n7816 = ( n181 & n2109 ) | ( n181 & ~n7815 ) | ( n2109 & ~n7815 ) ;
  assign n7817 = n948 | n4666 ;
  assign n7818 = n7817 ^ x125 ^ 1'b0 ;
  assign n7819 = ( n6810 & n7816 ) | ( n6810 & n7818 ) | ( n7816 & n7818 ) ;
  assign n7820 = ~n1456 & n7819 ;
  assign n7814 = ( ~n442 & n1509 ) | ( ~n442 & n5507 ) | ( n1509 & n5507 ) ;
  assign n7821 = n7820 ^ n7814 ^ n1577 ;
  assign n7822 = n7821 ^ n6640 ^ n3710 ;
  assign n7826 = n7825 ^ n7823 ^ n7822 ;
  assign n7827 = ~n667 & n6480 ;
  assign n7828 = n486 & n7827 ;
  assign n7829 = n7828 ^ n1450 ^ 1'b0 ;
  assign n7830 = ~n4629 & n4888 ;
  assign n7831 = n7830 ^ x66 ^ 1'b0 ;
  assign n7832 = n7831 ^ n5278 ^ n1636 ;
  assign n7833 = x32 & ~n7832 ;
  assign n7834 = n7833 ^ n243 ^ 1'b0 ;
  assign n7836 = n1736 ^ n832 ^ 1'b0 ;
  assign n7837 = n7836 ^ n3467 ^ 1'b0 ;
  assign n7838 = n7195 ^ n3813 ^ n1473 ;
  assign n7839 = ( n5096 & n7837 ) | ( n5096 & n7838 ) | ( n7837 & n7838 ) ;
  assign n7835 = ~n2492 & n7210 ;
  assign n7840 = n7839 ^ n7835 ^ 1'b0 ;
  assign n7841 = n1996 & ~n2520 ;
  assign n7842 = ~n819 & n7841 ;
  assign n7843 = ( n2511 & ~n5518 ) | ( n2511 & n6477 ) | ( ~n5518 & n6477 ) ;
  assign n7844 = n7843 ^ n2081 ^ 1'b0 ;
  assign n7845 = ~n7842 & n7844 ;
  assign n7846 = n7845 ^ n4571 ^ 1'b0 ;
  assign n7847 = n7207 ^ n6447 ^ n5311 ;
  assign n7848 = ( n541 & ~n5857 ) | ( n541 & n7847 ) | ( ~n5857 & n7847 ) ;
  assign n7849 = n7848 ^ n839 ^ 1'b0 ;
  assign n7850 = n7176 | n7849 ;
  assign n7851 = ( n376 & ~n6414 ) | ( n376 & n7850 ) | ( ~n6414 & n7850 ) ;
  assign n7852 = n5228 & ~n6368 ;
  assign n7853 = n5131 ^ n2765 ^ n379 ;
  assign n7854 = ~n4128 & n4361 ;
  assign n7855 = n5671 ^ n2581 ^ 1'b0 ;
  assign n7856 = n738 | n7855 ;
  assign n7857 = n4970 & ~n7856 ;
  assign n7863 = ~n1147 & n5001 ;
  assign n7858 = n4189 ^ n2241 ^ 1'b0 ;
  assign n7859 = ( ~n606 & n894 ) | ( ~n606 & n1763 ) | ( n894 & n1763 ) ;
  assign n7860 = n4200 ^ n984 ^ 1'b0 ;
  assign n7861 = n7859 & n7860 ;
  assign n7862 = n7858 & n7861 ;
  assign n7864 = n7863 ^ n7862 ^ 1'b0 ;
  assign n7865 = ~n619 & n2678 ;
  assign n7866 = n3163 & n7865 ;
  assign n7867 = n5299 ^ n4571 ^ n337 ;
  assign n7868 = n7867 ^ n3193 ^ 1'b0 ;
  assign n7869 = n5438 & n7868 ;
  assign n7870 = ~n805 & n1654 ;
  assign n7871 = n7870 ^ n7056 ^ 1'b0 ;
  assign n7872 = x65 & ~n894 ;
  assign n7873 = n7872 ^ n2295 ^ 1'b0 ;
  assign n7874 = n7873 ^ n2364 ^ 1'b0 ;
  assign n7875 = x15 & ~n6348 ;
  assign n7876 = n7441 ^ n3549 ^ 1'b0 ;
  assign n7877 = n7876 ^ n7073 ^ 1'b0 ;
  assign n7878 = ( ~n5607 & n5777 ) | ( ~n5607 & n7877 ) | ( n5777 & n7877 ) ;
  assign n7881 = n4525 & ~n6847 ;
  assign n7882 = n7881 ^ n909 ^ 1'b0 ;
  assign n7880 = n5366 ^ n616 ^ x66 ;
  assign n7879 = n2029 ^ n652 ^ 1'b0 ;
  assign n7883 = n7882 ^ n7880 ^ n7879 ;
  assign n7884 = n7677 ^ n4593 ^ n3979 ;
  assign n7885 = n5243 & ~n7884 ;
  assign n7886 = n214 & n1168 ;
  assign n7887 = x15 & n965 ;
  assign n7888 = n7887 ^ n1404 ^ 1'b0 ;
  assign n7889 = ( n2922 & ~n3534 ) | ( n2922 & n7888 ) | ( ~n3534 & n7888 ) ;
  assign n7890 = ( n401 & n664 ) | ( n401 & ~n1422 ) | ( n664 & ~n1422 ) ;
  assign n7897 = n3628 ^ n2415 ^ 1'b0 ;
  assign n7898 = ( n393 & n2960 ) | ( n393 & n7897 ) | ( n2960 & n7897 ) ;
  assign n7892 = n3588 & n6352 ;
  assign n7893 = n7892 ^ n1330 ^ 1'b0 ;
  assign n7894 = n7893 ^ n4512 ^ 1'b0 ;
  assign n7895 = ~n925 & n7894 ;
  assign n7891 = n1648 ^ n1366 ^ 1'b0 ;
  assign n7896 = n7895 ^ n7891 ^ 1'b0 ;
  assign n7899 = n7898 ^ n7896 ^ 1'b0 ;
  assign n7900 = ( n3883 & ~n7890 ) | ( n3883 & n7899 ) | ( ~n7890 & n7899 ) ;
  assign n7901 = ( ~n176 & n1270 ) | ( ~n176 & n2103 ) | ( n1270 & n2103 ) ;
  assign n7902 = ( n4932 & n7189 ) | ( n4932 & ~n7901 ) | ( n7189 & ~n7901 ) ;
  assign n7906 = n3922 ^ n1918 ^ n586 ;
  assign n7904 = n3674 ^ n1704 ^ 1'b0 ;
  assign n7905 = ~n6156 & n7904 ;
  assign n7907 = n7906 ^ n7905 ^ 1'b0 ;
  assign n7908 = n6716 | n7907 ;
  assign n7909 = n7528 & ~n7908 ;
  assign n7903 = ~n2670 & n3262 ;
  assign n7910 = n7909 ^ n7903 ^ 1'b0 ;
  assign n7913 = n4559 ^ n1002 ^ n683 ;
  assign n7911 = n1217 & ~n2135 ;
  assign n7912 = n7911 ^ n3188 ^ n842 ;
  assign n7914 = n7913 ^ n7912 ^ n4644 ;
  assign n7915 = n1374 & ~n1977 ;
  assign n7916 = n7915 ^ n2970 ^ 1'b0 ;
  assign n7917 = x68 ^ x38 ^ 1'b0 ;
  assign n7918 = ( n3528 & n7916 ) | ( n3528 & ~n7917 ) | ( n7916 & ~n7917 ) ;
  assign n7919 = ( ~n1819 & n3237 ) | ( ~n1819 & n5216 ) | ( n3237 & n5216 ) ;
  assign n7920 = n6532 ^ x48 ^ 1'b0 ;
  assign n7921 = ( ~n7918 & n7919 ) | ( ~n7918 & n7920 ) | ( n7919 & n7920 ) ;
  assign n7922 = ~n1388 & n5630 ;
  assign n7923 = ~n3487 & n7922 ;
  assign n7924 = ~n3085 & n6908 ;
  assign n7925 = n7924 ^ n449 ^ 1'b0 ;
  assign n7928 = ( ~n583 & n5071 ) | ( ~n583 & n5871 ) | ( n5071 & n5871 ) ;
  assign n7926 = n1379 | n3515 ;
  assign n7927 = n7926 ^ n3957 ^ 1'b0 ;
  assign n7929 = n7928 ^ n7927 ^ n6046 ;
  assign n7931 = n1148 & n2894 ;
  assign n7932 = ~n179 & n7931 ;
  assign n7933 = n1711 | n7932 ;
  assign n7934 = n4659 | n7933 ;
  assign n7930 = n5343 ^ n3597 ^ n562 ;
  assign n7935 = n7934 ^ n7930 ^ n945 ;
  assign n7936 = n1226 | n7935 ;
  assign n7937 = n7929 | n7936 ;
  assign n7938 = n7356 ^ n7133 ^ 1'b0 ;
  assign n7939 = ( n2887 & n4689 ) | ( n2887 & ~n7938 ) | ( n4689 & ~n7938 ) ;
  assign n7940 = n1797 ^ n1312 ^ n1203 ;
  assign n7941 = n7939 | n7940 ;
  assign n7942 = n7941 ^ n1563 ^ 1'b0 ;
  assign n7943 = n7942 ^ n1854 ^ n1653 ;
  assign n7944 = n7943 ^ n5824 ^ n828 ;
  assign n7945 = ~n367 & n1782 ;
  assign n7946 = ~n7944 & n7945 ;
  assign n7947 = n2178 & ~n3045 ;
  assign n7948 = ~n3292 & n7947 ;
  assign n7949 = n5616 ^ n279 ^ 1'b0 ;
  assign n7950 = n2464 & n2900 ;
  assign n7951 = ~n7949 & n7950 ;
  assign n7952 = n3769 ^ n3035 ^ n1592 ;
  assign n7953 = ( n2506 & n2830 ) | ( n2506 & ~n4101 ) | ( n2830 & ~n4101 ) ;
  assign n7954 = n5891 ^ n934 ^ x110 ;
  assign n7955 = ( ~n2334 & n7953 ) | ( ~n2334 & n7954 ) | ( n7953 & n7954 ) ;
  assign n7956 = n2601 & n7955 ;
  assign n7957 = ~n7952 & n7956 ;
  assign n7958 = n7957 ^ n6325 ^ 1'b0 ;
  assign n7959 = n7951 | n7958 ;
  assign n7963 = n4132 ^ n1646 ^ n505 ;
  assign n7964 = ( n2414 & n2569 ) | ( n2414 & ~n5483 ) | ( n2569 & ~n5483 ) ;
  assign n7965 = ( n5597 & n7963 ) | ( n5597 & n7964 ) | ( n7963 & n7964 ) ;
  assign n7966 = n7965 ^ n4867 ^ 1'b0 ;
  assign n7967 = n6535 | n7966 ;
  assign n7960 = n3409 ^ n263 ^ 1'b0 ;
  assign n7961 = n2102 & n7960 ;
  assign n7962 = n7961 ^ n4305 ^ n3625 ;
  assign n7968 = n7967 ^ n7962 ^ n6064 ;
  assign n7969 = n1902 & ~n2905 ;
  assign n7970 = n7969 ^ n3915 ^ 1'b0 ;
  assign n7971 = ( n1611 & ~n7067 ) | ( n1611 & n7970 ) | ( ~n7067 & n7970 ) ;
  assign n7972 = n7971 ^ n4254 ^ 1'b0 ;
  assign n7973 = n2530 & ~n7972 ;
  assign n7974 = n5353 ^ n915 ^ 1'b0 ;
  assign n7975 = n7957 | n7974 ;
  assign n7976 = n3124 & n3732 ;
  assign n7977 = n5103 & n7976 ;
  assign n7978 = n1553 ^ n1355 ^ 1'b0 ;
  assign n7979 = ( n635 & ~n2172 ) | ( n635 & n7978 ) | ( ~n2172 & n7978 ) ;
  assign n7980 = n7979 ^ n6686 ^ n6244 ;
  assign n7981 = n7317 ^ n6737 ^ n3150 ;
  assign n7982 = n5494 ^ n3007 ^ 1'b0 ;
  assign n7983 = n880 & n6957 ;
  assign n7984 = n5650 & n7983 ;
  assign n7985 = ~n7982 & n7984 ;
  assign n7986 = n5649 & n7985 ;
  assign n7987 = ( n388 & n694 ) | ( n388 & ~n1357 ) | ( n694 & ~n1357 ) ;
  assign n7989 = n1273 & ~n3998 ;
  assign n7990 = n2523 & n7989 ;
  assign n7991 = n3147 & ~n4780 ;
  assign n7992 = ~n1767 & n7991 ;
  assign n7993 = ( n172 & ~n7990 ) | ( n172 & n7992 ) | ( ~n7990 & n7992 ) ;
  assign n7988 = n1732 | n3979 ;
  assign n7994 = n7993 ^ n7988 ^ 1'b0 ;
  assign n7995 = ( ~n2295 & n7987 ) | ( ~n2295 & n7994 ) | ( n7987 & n7994 ) ;
  assign n7996 = n1052 & n3091 ;
  assign n8005 = ~n4840 & n7667 ;
  assign n8000 = ~n3297 & n7187 ;
  assign n8001 = n8000 ^ n2523 ^ 1'b0 ;
  assign n8002 = n8001 ^ n2643 ^ n2116 ;
  assign n7997 = x122 & n2749 ;
  assign n7998 = n7997 ^ n6093 ^ 1'b0 ;
  assign n7999 = n4087 & n7998 ;
  assign n8003 = n8002 ^ n7999 ^ 1'b0 ;
  assign n8004 = ( n1133 & n1645 ) | ( n1133 & ~n8003 ) | ( n1645 & ~n8003 ) ;
  assign n8006 = n8005 ^ n8004 ^ n4657 ;
  assign n8014 = n2466 & ~n7405 ;
  assign n8015 = n8014 ^ n7542 ^ n2077 ;
  assign n8007 = n6368 ^ n879 ^ n211 ;
  assign n8008 = n8007 ^ n7651 ^ n5286 ;
  assign n8009 = n1514 & n4924 ;
  assign n8010 = ~n401 & n8009 ;
  assign n8011 = n4028 ^ n2232 ^ 1'b0 ;
  assign n8012 = n8010 | n8011 ;
  assign n8013 = n8008 & n8012 ;
  assign n8016 = n8015 ^ n8013 ^ n4360 ;
  assign n8017 = n3092 ^ n3026 ^ n1888 ;
  assign n8018 = n915 & ~n8017 ;
  assign n8019 = n3186 & n8018 ;
  assign n8020 = n5356 ^ n2951 ^ 1'b0 ;
  assign n8021 = ~n503 & n3014 ;
  assign n8022 = n8020 & n8021 ;
  assign n8026 = ( n1434 & n3442 ) | ( n1434 & n3963 ) | ( n3442 & n3963 ) ;
  assign n8027 = n8026 ^ n6300 ^ 1'b0 ;
  assign n8028 = n233 | n8027 ;
  assign n8023 = ( ~n225 & n268 ) | ( ~n225 & n2519 ) | ( n268 & n2519 ) ;
  assign n8024 = n8023 ^ n5296 ^ 1'b0 ;
  assign n8025 = n1172 | n8024 ;
  assign n8029 = n8028 ^ n8025 ^ 1'b0 ;
  assign n8030 = n4983 & n8029 ;
  assign n8032 = n6378 ^ n4090 ^ n654 ;
  assign n8031 = ~n834 & n5413 ;
  assign n8033 = n8032 ^ n8031 ^ 1'b0 ;
  assign n8034 = n6758 ^ n510 ^ 1'b0 ;
  assign n8040 = n1026 & n1639 ;
  assign n8041 = ~n1639 & n8040 ;
  assign n8042 = n136 | n186 ;
  assign n8043 = n8041 & ~n8042 ;
  assign n8044 = n6795 ^ n277 ^ x49 ;
  assign n8045 = n1913 & ~n8044 ;
  assign n8046 = n8044 & n8045 ;
  assign n8047 = n4036 & ~n8046 ;
  assign n8048 = n8043 & n8047 ;
  assign n8049 = n649 & ~n3680 ;
  assign n8050 = n8048 & n8049 ;
  assign n8037 = n5120 ^ n2584 ^ n2338 ;
  assign n8035 = n426 ^ n377 ^ 1'b0 ;
  assign n8036 = ~n7151 & n8035 ;
  assign n8038 = n8037 ^ n8036 ^ 1'b0 ;
  assign n8039 = n3627 | n8038 ;
  assign n8051 = n8050 ^ n8039 ^ 1'b0 ;
  assign n8052 = n3677 ^ n2293 ^ 1'b0 ;
  assign n8053 = ~n3451 & n8052 ;
  assign n8054 = n795 & n8053 ;
  assign n8055 = n6191 | n8054 ;
  assign n8056 = n8055 ^ n4758 ^ 1'b0 ;
  assign n8057 = n4641 ^ n4189 ^ 1'b0 ;
  assign n8058 = n8056 | n8057 ;
  assign n8061 = n1125 | n4535 ;
  assign n8062 = n1616 & ~n8061 ;
  assign n8063 = n7691 | n8062 ;
  assign n8064 = n4016 & ~n8063 ;
  assign n8059 = n3317 ^ n1196 ^ n611 ;
  assign n8060 = ~n1114 & n8059 ;
  assign n8065 = n8064 ^ n8060 ^ 1'b0 ;
  assign n8066 = n8065 ^ n4276 ^ n2994 ;
  assign n8067 = n8058 & n8066 ;
  assign n8068 = n1876 & ~n5469 ;
  assign n8069 = n8067 & n8068 ;
  assign n8070 = n1504 | n2593 ;
  assign n8071 = n8070 ^ n1648 ^ 1'b0 ;
  assign n8072 = n8071 ^ n3567 ^ 1'b0 ;
  assign n8073 = n2288 & n6282 ;
  assign n8074 = n1481 & n8073 ;
  assign n8075 = n8074 ^ n6472 ^ n5531 ;
  assign n8076 = n8075 ^ n5182 ^ 1'b0 ;
  assign n8077 = n1516 & ~n2151 ;
  assign n8078 = n8076 & n8077 ;
  assign n8079 = ( ~n362 & n8072 ) | ( ~n362 & n8078 ) | ( n8072 & n8078 ) ;
  assign n8080 = n1828 | n6454 ;
  assign n8081 = n2691 & ~n8080 ;
  assign n8082 = ~n6633 & n7272 ;
  assign n8083 = n3726 & n4497 ;
  assign n8084 = ( n846 & n1320 ) | ( n846 & n2557 ) | ( n1320 & n2557 ) ;
  assign n8085 = n8084 ^ n1874 ^ 1'b0 ;
  assign n8086 = n2665 & n8085 ;
  assign n8087 = n8086 ^ n1620 ^ n284 ;
  assign n8088 = n2573 & n8087 ;
  assign n8089 = n4383 & n8088 ;
  assign n8090 = ~n958 & n5496 ;
  assign n8091 = ~n4320 & n8090 ;
  assign n8092 = n8091 ^ n7654 ^ 1'b0 ;
  assign n8102 = ~n3749 & n3891 ;
  assign n8103 = n8102 ^ n7602 ^ 1'b0 ;
  assign n8099 = n1095 & ~n7468 ;
  assign n8100 = n8099 ^ n844 ^ 1'b0 ;
  assign n8093 = n6226 ^ n663 ^ 1'b0 ;
  assign n8094 = n3898 & n6123 ;
  assign n8095 = n7821 & n8094 ;
  assign n8096 = n3085 & n8095 ;
  assign n8097 = n4240 ^ n1706 ^ x49 ;
  assign n8098 = ( n8093 & ~n8096 ) | ( n8093 & n8097 ) | ( ~n8096 & n8097 ) ;
  assign n8101 = n8100 ^ n8098 ^ n7302 ;
  assign n8104 = n8103 ^ n8101 ^ n7657 ;
  assign n8105 = n7317 ^ n5168 ^ n233 ;
  assign n8106 = n1270 & ~n6964 ;
  assign n8107 = n8106 ^ n568 ^ 1'b0 ;
  assign n8108 = n8107 ^ n3469 ^ 1'b0 ;
  assign n8109 = n501 & ~n8108 ;
  assign n8110 = n8109 ^ n2816 ^ 1'b0 ;
  assign n8111 = n2026 & ~n2303 ;
  assign n8112 = n8111 ^ n4004 ^ n702 ;
  assign n8113 = ( n4867 & ~n5393 ) | ( n4867 & n8112 ) | ( ~n5393 & n8112 ) ;
  assign n8114 = ( n253 & n5229 ) | ( n253 & n5789 ) | ( n5229 & n5789 ) ;
  assign n8116 = n4864 ^ n3317 ^ 1'b0 ;
  assign n8117 = n2837 | n8116 ;
  assign n8118 = n8117 ^ n6836 ^ n1973 ;
  assign n8119 = ( ~n265 & n6735 ) | ( ~n265 & n8118 ) | ( n6735 & n8118 ) ;
  assign n8120 = n8119 ^ n5913 ^ 1'b0 ;
  assign n8121 = n2710 & ~n8120 ;
  assign n8122 = n8121 ^ n7085 ^ n4151 ;
  assign n8115 = n1999 | n2649 ;
  assign n8123 = n8122 ^ n8115 ^ 1'b0 ;
  assign n8129 = n1898 ^ n947 ^ n649 ;
  assign n8124 = ~n456 & n800 ;
  assign n8125 = ~n167 & n8124 ;
  assign n8126 = n8125 ^ n2557 ^ x55 ;
  assign n8127 = n8126 ^ n3569 ^ n697 ;
  assign n8128 = n8127 ^ n2583 ^ n2523 ;
  assign n8130 = n8129 ^ n8128 ^ n4528 ;
  assign n8131 = ( x96 & ~n714 ) | ( x96 & n8130 ) | ( ~n714 & n8130 ) ;
  assign n8132 = n5391 ^ n219 ^ 1'b0 ;
  assign n8133 = ~n698 & n816 ;
  assign n8134 = n5843 & n8133 ;
  assign n8135 = ( n2304 & n8132 ) | ( n2304 & n8134 ) | ( n8132 & n8134 ) ;
  assign n8136 = ~n1093 & n3295 ;
  assign n8138 = ( n1808 & n2523 ) | ( n1808 & ~n3382 ) | ( n2523 & ~n3382 ) ;
  assign n8139 = ( ~n281 & n971 ) | ( ~n281 & n8138 ) | ( n971 & n8138 ) ;
  assign n8137 = n2625 | n2754 ;
  assign n8140 = n8139 ^ n8137 ^ 1'b0 ;
  assign n8141 = ~n8136 & n8140 ;
  assign n8142 = ( n6317 & n8135 ) | ( n6317 & ~n8141 ) | ( n8135 & ~n8141 ) ;
  assign n8143 = n1368 & ~n2667 ;
  assign n8144 = n5585 & n8143 ;
  assign n8145 = n2832 ^ n2815 ^ n1099 ;
  assign n8146 = n828 ^ n767 ^ n677 ;
  assign n8147 = n8145 | n8146 ;
  assign n8148 = n2914 ^ n1454 ^ 1'b0 ;
  assign n8149 = n5679 ^ n1794 ^ 1'b0 ;
  assign n8150 = n1611 & n2174 ;
  assign n8151 = n8150 ^ n434 ^ 1'b0 ;
  assign n8152 = x127 & ~n8151 ;
  assign n8153 = n8152 ^ n4394 ^ 1'b0 ;
  assign n8154 = n5809 & ~n8153 ;
  assign n8156 = n7405 ^ n2046 ^ n1166 ;
  assign n8155 = n2331 | n7306 ;
  assign n8157 = n8156 ^ n8155 ^ 1'b0 ;
  assign n8158 = n141 & n3553 ;
  assign n8159 = n5589 ^ n3631 ^ n1330 ;
  assign n8162 = ( ~n691 & n751 ) | ( ~n691 & n2615 ) | ( n751 & n2615 ) ;
  assign n8160 = n2461 | n4580 ;
  assign n8161 = n2557 & ~n8160 ;
  assign n8163 = n8162 ^ n8161 ^ n7109 ;
  assign n8164 = n3626 ^ n1392 ^ 1'b0 ;
  assign n8165 = n8164 ^ n7092 ^ n4744 ;
  assign n8166 = n1374 ^ n811 ^ 1'b0 ;
  assign n8167 = ( n550 & n1575 ) | ( n550 & ~n2067 ) | ( n1575 & ~n2067 ) ;
  assign n8168 = ~n5331 & n8167 ;
  assign n8169 = n8168 ^ n7511 ^ 1'b0 ;
  assign n8170 = ( ~x19 & n2374 ) | ( ~x19 & n7181 ) | ( n2374 & n7181 ) ;
  assign n8171 = n595 | n8170 ;
  assign n8175 = ( ~n974 & n1674 ) | ( ~n974 & n3033 ) | ( n1674 & n3033 ) ;
  assign n8172 = ( n374 & n1837 ) | ( n374 & ~n3705 ) | ( n1837 & ~n3705 ) ;
  assign n8173 = ( ~n2021 & n5807 ) | ( ~n2021 & n8172 ) | ( n5807 & n8172 ) ;
  assign n8174 = n3347 | n8173 ;
  assign n8176 = n8175 ^ n8174 ^ 1'b0 ;
  assign n8177 = n6800 ^ n6579 ^ 1'b0 ;
  assign n8178 = n3603 & ~n8177 ;
  assign n8179 = n6964 ^ n6735 ^ n1612 ;
  assign n8180 = ( ~n1922 & n3539 ) | ( ~n1922 & n8179 ) | ( n3539 & n8179 ) ;
  assign n8181 = n2491 | n3741 ;
  assign n8183 = n6690 ^ n1859 ^ n184 ;
  assign n8184 = ~n530 & n8183 ;
  assign n8185 = n2598 & n8184 ;
  assign n8186 = ~n2390 & n8185 ;
  assign n8182 = n4377 & ~n5464 ;
  assign n8187 = n8186 ^ n8182 ^ n8147 ;
  assign n8188 = n345 | n3012 ;
  assign n8189 = n4498 & ~n8188 ;
  assign n8190 = n8189 ^ n5780 ^ n3925 ;
  assign n8191 = n3690 ^ n2583 ^ n575 ;
  assign n8192 = ~n4305 & n6354 ;
  assign n8193 = n8191 & n8192 ;
  assign n8194 = n8193 ^ n1149 ^ 1'b0 ;
  assign n8195 = n8190 | n8194 ;
  assign n8196 = n2847 & n3205 ;
  assign n8197 = n8195 & n8196 ;
  assign n8198 = n4882 & n5650 ;
  assign n8199 = n8198 ^ n3703 ^ 1'b0 ;
  assign n8200 = n6046 | n8199 ;
  assign n8201 = n2596 ^ n2293 ^ n443 ;
  assign n8202 = n8201 ^ n2021 ^ n1865 ;
  assign n8203 = ( ~n2781 & n6218 ) | ( ~n2781 & n8202 ) | ( n6218 & n8202 ) ;
  assign n8204 = n8203 ^ n8059 ^ n1744 ;
  assign n8205 = n1073 | n8204 ;
  assign n8206 = n8205 ^ x99 ^ 1'b0 ;
  assign n8207 = n3582 | n8206 ;
  assign n8208 = ( n1298 & ~n2682 ) | ( n1298 & n6980 ) | ( ~n2682 & n6980 ) ;
  assign n8209 = n8208 ^ n7113 ^ n6002 ;
  assign n8210 = n8209 ^ n1268 ^ 1'b0 ;
  assign n8211 = ( n3785 & ~n5655 ) | ( n3785 & n5740 ) | ( ~n5655 & n5740 ) ;
  assign n8212 = n4961 & ~n6636 ;
  assign n8213 = n8212 ^ n7660 ^ n2667 ;
  assign n8214 = ( ~n3157 & n3657 ) | ( ~n3157 & n8213 ) | ( n3657 & n8213 ) ;
  assign n8215 = n1479 & n2985 ;
  assign n8216 = n8215 ^ n5530 ^ n929 ;
  assign n8217 = n8216 ^ n4279 ^ n3593 ;
  assign n8218 = x35 & ~n4948 ;
  assign n8219 = n8218 ^ n6247 ^ 1'b0 ;
  assign n8220 = n8219 ^ n2657 ^ 1'b0 ;
  assign n8221 = ~n1926 & n8220 ;
  assign n8222 = n8221 ^ n5438 ^ 1'b0 ;
  assign n8224 = ~n2383 & n2679 ;
  assign n8223 = ( ~n667 & n834 ) | ( ~n667 & n3662 ) | ( n834 & n3662 ) ;
  assign n8225 = n8224 ^ n8223 ^ 1'b0 ;
  assign n8226 = n580 ^ x83 ^ 1'b0 ;
  assign n8227 = n1507 | n8226 ;
  assign n8229 = n207 & ~n399 ;
  assign n8230 = n8229 ^ n2349 ^ 1'b0 ;
  assign n8228 = ( n1332 & n4682 ) | ( n1332 & n7691 ) | ( n4682 & n7691 ) ;
  assign n8231 = n8230 ^ n8228 ^ 1'b0 ;
  assign n8232 = n8227 | n8231 ;
  assign n8233 = n7232 | n8232 ;
  assign n8234 = ( n2334 & ~n5041 ) | ( n2334 & n5199 ) | ( ~n5041 & n5199 ) ;
  assign n8235 = n8234 ^ n3432 ^ 1'b0 ;
  assign n8236 = n8235 ^ n5862 ^ 1'b0 ;
  assign n8237 = n950 & ~n8236 ;
  assign n8238 = n2970 & n4412 ;
  assign n8239 = n3814 & n8238 ;
  assign n8240 = ~n1358 & n8239 ;
  assign n8241 = n8240 ^ n7850 ^ n1304 ;
  assign n8242 = n6230 ^ n2789 ^ n1593 ;
  assign n8243 = n3909 ^ n1639 ^ 1'b0 ;
  assign n8244 = ( n1411 & n6582 ) | ( n1411 & ~n8243 ) | ( n6582 & ~n8243 ) ;
  assign n8245 = ( n2541 & n7583 ) | ( n2541 & ~n8244 ) | ( n7583 & ~n8244 ) ;
  assign n8246 = ~n8242 & n8245 ;
  assign n8255 = n3943 ^ n386 ^ 1'b0 ;
  assign n8256 = n8255 ^ n731 ^ n453 ;
  assign n8253 = n5725 & ~n5837 ;
  assign n8249 = n2424 & ~n3769 ;
  assign n8250 = ~n3267 & n8249 ;
  assign n8251 = n8250 ^ n2012 ^ 1'b0 ;
  assign n8247 = n1969 & n2405 ;
  assign n8248 = n3733 & ~n8247 ;
  assign n8252 = n8251 ^ n8248 ^ 1'b0 ;
  assign n8254 = n8253 ^ n8252 ^ 1'b0 ;
  assign n8257 = n8256 ^ n8254 ^ 1'b0 ;
  assign n8258 = n2815 ^ n2229 ^ 1'b0 ;
  assign n8259 = n7828 & n8258 ;
  assign n8260 = ( n2179 & n4145 ) | ( n2179 & n8259 ) | ( n4145 & n8259 ) ;
  assign n8268 = ( ~n1388 & n2079 ) | ( ~n1388 & n6284 ) | ( n2079 & n6284 ) ;
  assign n8267 = n4159 & ~n7584 ;
  assign n8269 = n8268 ^ n8267 ^ 1'b0 ;
  assign n8270 = n4591 ^ n1391 ^ 1'b0 ;
  assign n8271 = ~n7736 & n8270 ;
  assign n8272 = n8269 & n8271 ;
  assign n8262 = n3942 ^ n1213 ^ x124 ;
  assign n8263 = ( n4076 & n5674 ) | ( n4076 & n8262 ) | ( n5674 & n8262 ) ;
  assign n8261 = n8094 ^ n7549 ^ n4353 ;
  assign n8264 = n8263 ^ n8261 ^ 1'b0 ;
  assign n8265 = n2399 | n8264 ;
  assign n8266 = n8227 | n8265 ;
  assign n8273 = n8272 ^ n8266 ^ 1'b0 ;
  assign n8274 = n4033 & ~n4121 ;
  assign n8275 = n8274 ^ n1899 ^ 1'b0 ;
  assign n8276 = n6690 ^ n2781 ^ n1123 ;
  assign n8277 = n8276 ^ n259 ^ 1'b0 ;
  assign n8278 = n5865 ^ n3471 ^ 1'b0 ;
  assign n8279 = n3511 | n8278 ;
  assign n8280 = n437 & n4320 ;
  assign n8281 = n8279 & n8280 ;
  assign n8282 = ~n8277 & n8281 ;
  assign n8283 = n8282 ^ n337 ^ 1'b0 ;
  assign n8284 = ( ~x97 & n1707 ) | ( ~x97 & n6220 ) | ( n1707 & n6220 ) ;
  assign n8285 = n956 & n8284 ;
  assign n8286 = n4438 ^ n1320 ^ 1'b0 ;
  assign n8291 = n379 | n6870 ;
  assign n8292 = n3620 | n8291 ;
  assign n8287 = n986 ^ n964 ^ 1'b0 ;
  assign n8288 = n7626 ^ n4016 ^ n3561 ;
  assign n8289 = n8288 ^ n6371 ^ 1'b0 ;
  assign n8290 = n8287 & ~n8289 ;
  assign n8293 = n8292 ^ n8290 ^ 1'b0 ;
  assign n8294 = n2283 & n8293 ;
  assign n8295 = n8294 ^ n1656 ^ n190 ;
  assign n8296 = n8026 | n8295 ;
  assign n8301 = ( n1011 & n2802 ) | ( n1011 & n6160 ) | ( n2802 & n6160 ) ;
  assign n8297 = n3163 ^ n3027 ^ 1'b0 ;
  assign n8298 = ~n5871 & n8297 ;
  assign n8299 = n2113 ^ n1534 ^ 1'b0 ;
  assign n8300 = n8298 & ~n8299 ;
  assign n8302 = n8301 ^ n8300 ^ n7675 ;
  assign n8303 = n8302 ^ n4918 ^ n2738 ;
  assign n8304 = n3071 | n6270 ;
  assign n8305 = ( ~n3926 & n8303 ) | ( ~n3926 & n8304 ) | ( n8303 & n8304 ) ;
  assign n8306 = n8305 ^ n7680 ^ 1'b0 ;
  assign n8307 = n5060 & n8306 ;
  assign n8308 = n8307 ^ n5460 ^ n4865 ;
  assign n8309 = n4137 ^ n719 ^ 1'b0 ;
  assign n8310 = x41 & ~n8309 ;
  assign n8311 = ( n1343 & n2089 ) | ( n1343 & n6845 ) | ( n2089 & n6845 ) ;
  assign n8312 = n8311 ^ n4249 ^ n2089 ;
  assign n8314 = ( n575 & ~n5096 ) | ( n575 & n5680 ) | ( ~n5096 & n5680 ) ;
  assign n8313 = n5337 ^ n3377 ^ n275 ;
  assign n8315 = n8314 ^ n8313 ^ 1'b0 ;
  assign n8316 = ~n2310 & n8315 ;
  assign n8317 = n1470 & n5121 ;
  assign n8318 = n8317 ^ n4450 ^ 1'b0 ;
  assign n8319 = n8318 ^ n2002 ^ n1452 ;
  assign n8320 = n4895 ^ n1997 ^ 1'b0 ;
  assign n8321 = n8320 ^ n1444 ^ 1'b0 ;
  assign n8322 = n5715 & ~n7508 ;
  assign n8323 = n8322 ^ n6707 ^ 1'b0 ;
  assign n8324 = ~n3640 & n8323 ;
  assign n8325 = n3845 ^ n3262 ^ 1'b0 ;
  assign n8326 = ( n2475 & ~n6672 ) | ( n2475 & n8325 ) | ( ~n6672 & n8325 ) ;
  assign n8327 = n8247 & ~n8326 ;
  assign n8335 = ( n1929 & n2329 ) | ( n1929 & ~n6159 ) | ( n2329 & ~n6159 ) ;
  assign n8336 = n1633 & ~n4016 ;
  assign n8337 = ~n602 & n8336 ;
  assign n8338 = ( ~n5776 & n8335 ) | ( ~n5776 & n8337 ) | ( n8335 & n8337 ) ;
  assign n8334 = n4202 ^ n2787 ^ 1'b0 ;
  assign n8328 = n2798 | n6796 ;
  assign n8329 = n4705 & ~n8328 ;
  assign n8330 = n5150 ^ n481 ^ 1'b0 ;
  assign n8331 = n8330 ^ n8156 ^ n1450 ;
  assign n8332 = n8331 ^ n4043 ^ n915 ;
  assign n8333 = n8329 & n8332 ;
  assign n8339 = n8338 ^ n8334 ^ n8333 ;
  assign n8340 = n6665 ^ n955 ^ 1'b0 ;
  assign n8341 = n377 | n8340 ;
  assign n8342 = n945 & n3371 ;
  assign n8343 = ~n5706 & n8342 ;
  assign n8344 = ( n162 & n6997 ) | ( n162 & ~n8343 ) | ( n6997 & ~n8343 ) ;
  assign n8345 = n5656 ^ n1409 ^ 1'b0 ;
  assign n8346 = ( ~n8341 & n8344 ) | ( ~n8341 & n8345 ) | ( n8344 & n8345 ) ;
  assign n8347 = ~n2863 & n4521 ;
  assign n8348 = n8347 ^ n1798 ^ 1'b0 ;
  assign n8349 = n8348 ^ n8255 ^ n3953 ;
  assign n8350 = ( n872 & n1531 ) | ( n872 & ~n8349 ) | ( n1531 & ~n8349 ) ;
  assign n8351 = n3839 ^ n468 ^ 1'b0 ;
  assign n8354 = n162 & ~n712 ;
  assign n8352 = ( n1394 & ~n4665 ) | ( n1394 & n5261 ) | ( ~n4665 & n5261 ) ;
  assign n8353 = n6324 & ~n8352 ;
  assign n8355 = n8354 ^ n8353 ^ 1'b0 ;
  assign n8356 = n3077 & ~n4098 ;
  assign n8357 = n8355 & ~n8356 ;
  assign n8358 = ~n1904 & n8357 ;
  assign n8359 = n7415 & ~n8358 ;
  assign n8360 = n8359 ^ x17 ^ 1'b0 ;
  assign n8361 = ( n4022 & n5034 ) | ( n4022 & ~n5566 ) | ( n5034 & ~n5566 ) ;
  assign n8362 = n8361 ^ n6570 ^ n2826 ;
  assign n8363 = n8007 ^ n1235 ^ n1109 ;
  assign n8364 = ( ~n729 & n2909 ) | ( ~n729 & n8363 ) | ( n2909 & n8363 ) ;
  assign n8366 = ( x51 & ~n4163 ) | ( x51 & n5870 ) | ( ~n4163 & n5870 ) ;
  assign n8367 = ( n570 & n1524 ) | ( n570 & n4864 ) | ( n1524 & n4864 ) ;
  assign n8368 = n8367 ^ n2428 ^ 1'b0 ;
  assign n8369 = ( n5294 & ~n8366 ) | ( n5294 & n8368 ) | ( ~n8366 & n8368 ) ;
  assign n8370 = ( n7256 & n7322 ) | ( n7256 & n8369 ) | ( n7322 & n8369 ) ;
  assign n8365 = ~n1802 & n5831 ;
  assign n8371 = n8370 ^ n8365 ^ 1'b0 ;
  assign n8374 = n7250 ^ n6067 ^ 1'b0 ;
  assign n8372 = n2105 ^ n466 ^ 1'b0 ;
  assign n8373 = x51 & n8372 ;
  assign n8375 = n8374 ^ n8373 ^ 1'b0 ;
  assign n8376 = n6752 & ~n8375 ;
  assign n8377 = n8376 ^ n3428 ^ 1'b0 ;
  assign n8378 = n8377 ^ n6187 ^ n1643 ;
  assign n8379 = ( n136 & ~n511 ) | ( n136 & n1104 ) | ( ~n511 & n1104 ) ;
  assign n8380 = ( n485 & n802 ) | ( n485 & ~n7970 ) | ( n802 & ~n7970 ) ;
  assign n8381 = n8380 ^ n5770 ^ 1'b0 ;
  assign n8382 = ( n6812 & n8379 ) | ( n6812 & n8381 ) | ( n8379 & n8381 ) ;
  assign n8383 = n879 ^ n875 ^ n692 ;
  assign n8384 = n2388 | n7236 ;
  assign n8385 = n6262 & ~n8384 ;
  assign n8386 = ( n7614 & n8383 ) | ( n7614 & ~n8385 ) | ( n8383 & ~n8385 ) ;
  assign n8387 = ( n880 & ~n3028 ) | ( n880 & n4140 ) | ( ~n3028 & n4140 ) ;
  assign n8388 = n876 & n7665 ;
  assign n8389 = ( n1561 & n4407 ) | ( n1561 & n5330 ) | ( n4407 & n5330 ) ;
  assign n8390 = ( n910 & ~n4786 ) | ( n910 & n8007 ) | ( ~n4786 & n8007 ) ;
  assign n8391 = n2589 ^ n424 ^ 1'b0 ;
  assign n8392 = ~n2185 & n2277 ;
  assign n8393 = ~n8391 & n8392 ;
  assign n8394 = n5915 | n8393 ;
  assign n8395 = n8390 | n8394 ;
  assign n8396 = ~n2090 & n3364 ;
  assign n8397 = n783 | n8396 ;
  assign n8398 = n8397 ^ n5449 ^ 1'b0 ;
  assign n8399 = n8395 & ~n8398 ;
  assign n8400 = n2631 ^ n990 ^ 1'b0 ;
  assign n8401 = ( n483 & ~n1036 ) | ( n483 & n1859 ) | ( ~n1036 & n1859 ) ;
  assign n8402 = n8401 ^ n4592 ^ 1'b0 ;
  assign n8403 = n8400 | n8402 ;
  assign n8404 = n1399 | n8403 ;
  assign n8408 = n153 | n3079 ;
  assign n8405 = x22 & n1324 ;
  assign n8406 = n1881 ^ x68 ^ 1'b0 ;
  assign n8407 = ( ~n6305 & n8405 ) | ( ~n6305 & n8406 ) | ( n8405 & n8406 ) ;
  assign n8409 = n8408 ^ n8407 ^ n6073 ;
  assign n8410 = n1291 ^ x99 ^ 1'b0 ;
  assign n8411 = n3919 | n8410 ;
  assign n8412 = n8411 ^ n2374 ^ 1'b0 ;
  assign n8413 = ~n568 & n8412 ;
  assign n8414 = n1514 ^ n298 ^ 1'b0 ;
  assign n8415 = n8413 & ~n8414 ;
  assign n8416 = ( n5624 & n8409 ) | ( n5624 & ~n8415 ) | ( n8409 & ~n8415 ) ;
  assign n8417 = n8416 ^ n1694 ^ n468 ;
  assign n8424 = n5062 | n5597 ;
  assign n8425 = n7420 ^ n2537 ^ 1'b0 ;
  assign n8426 = n8424 | n8425 ;
  assign n8427 = n2318 | n8426 ;
  assign n8418 = n253 & n3248 ;
  assign n8419 = ~n615 & n8418 ;
  assign n8420 = n4016 ^ n2093 ^ 1'b0 ;
  assign n8421 = n8420 ^ n3186 ^ 1'b0 ;
  assign n8422 = n8421 ^ n7648 ^ n1177 ;
  assign n8423 = ( ~n7819 & n8419 ) | ( ~n7819 & n8422 ) | ( n8419 & n8422 ) ;
  assign n8428 = n8427 ^ n8423 ^ 1'b0 ;
  assign n8429 = n5797 | n8428 ;
  assign n8432 = n2859 ^ n2590 ^ n226 ;
  assign n8433 = n5210 | n8432 ;
  assign n8434 = n7716 | n8433 ;
  assign n8430 = ~n131 & n489 ;
  assign n8431 = n8430 ^ n5472 ^ 1'b0 ;
  assign n8435 = n8434 ^ n8431 ^ n1084 ;
  assign n8436 = ( n7208 & n8429 ) | ( n7208 & ~n8435 ) | ( n8429 & ~n8435 ) ;
  assign n8438 = x19 & n257 ;
  assign n8439 = ~n6679 & n8438 ;
  assign n8440 = ( n3065 & n6751 ) | ( n3065 & ~n8439 ) | ( n6751 & ~n8439 ) ;
  assign n8437 = ( x121 & ~n4207 ) | ( x121 & n5201 ) | ( ~n4207 & n5201 ) ;
  assign n8441 = n8440 ^ n8437 ^ n3119 ;
  assign n8443 = n5791 ^ n4913 ^ 1'b0 ;
  assign n8442 = n5054 ^ n1859 ^ 1'b0 ;
  assign n8444 = n8443 ^ n8442 ^ n670 ;
  assign n8445 = n4409 | n6954 ;
  assign n8446 = n8445 ^ n1150 ^ 1'b0 ;
  assign n8447 = n8446 ^ n2299 ^ 1'b0 ;
  assign n8448 = ~n451 & n2274 ;
  assign n8449 = ~n6976 & n8448 ;
  assign n8450 = n2647 ^ n569 ^ 1'b0 ;
  assign n8451 = n5532 ^ n4793 ^ 1'b0 ;
  assign n8454 = ( ~n466 & n4158 ) | ( ~n466 & n4904 ) | ( n4158 & n4904 ) ;
  assign n8452 = n5542 ^ n1811 ^ n625 ;
  assign n8453 = ~x40 & n8452 ;
  assign n8455 = n8454 ^ n8453 ^ n6659 ;
  assign n8456 = n622 & n2840 ;
  assign n8457 = ~n8455 & n8456 ;
  assign n8458 = n214 & n1024 ;
  assign n8459 = n8458 ^ n2887 ^ 1'b0 ;
  assign n8460 = n8459 ^ n5513 ^ 1'b0 ;
  assign n8461 = ~n1691 & n2061 ;
  assign n8462 = ( ~n763 & n1022 ) | ( ~n763 & n8461 ) | ( n1022 & n8461 ) ;
  assign n8463 = n7198 ^ n5414 ^ n1310 ;
  assign n8464 = n388 & n8463 ;
  assign n8465 = n8464 ^ n6265 ^ 1'b0 ;
  assign n8466 = n8462 & n8465 ;
  assign n8467 = n2000 & n2786 ;
  assign n8468 = n4404 & n8467 ;
  assign n8469 = n5281 | n8468 ;
  assign n8470 = n2827 | n8469 ;
  assign n8471 = ( n1404 & n8466 ) | ( n1404 & ~n8470 ) | ( n8466 & ~n8470 ) ;
  assign n8472 = n5350 ^ n4811 ^ n2646 ;
  assign n8473 = ( n2537 & n2554 ) | ( n2537 & n8472 ) | ( n2554 & n8472 ) ;
  assign n8474 = n8272 ^ n5248 ^ n4479 ;
  assign n8477 = n5613 ^ n4462 ^ 1'b0 ;
  assign n8475 = n2535 ^ n1641 ^ 1'b0 ;
  assign n8476 = n8475 ^ n8228 ^ n5549 ;
  assign n8478 = n8477 ^ n8476 ^ n285 ;
  assign n8479 = ( n617 & n662 ) | ( n617 & ~n1108 ) | ( n662 & ~n1108 ) ;
  assign n8480 = n2542 & n8479 ;
  assign n8481 = n2541 & n8480 ;
  assign n8482 = ( ~n1100 & n2060 ) | ( ~n1100 & n4158 ) | ( n2060 & n4158 ) ;
  assign n8483 = n8482 ^ n5796 ^ n2449 ;
  assign n8484 = n1789 | n5364 ;
  assign n8485 = n2416 & ~n8484 ;
  assign n8486 = n2458 ^ n1903 ^ n394 ;
  assign n8487 = n1588 | n4447 ;
  assign n8488 = n1634 & ~n8487 ;
  assign n8489 = ( n5981 & n8486 ) | ( n5981 & ~n8488 ) | ( n8486 & ~n8488 ) ;
  assign n8490 = n801 | n4726 ;
  assign n8491 = ( n378 & n783 ) | ( n378 & ~n8490 ) | ( n783 & ~n8490 ) ;
  assign n8492 = n4347 ^ n1450 ^ 1'b0 ;
  assign n8493 = n1617 & n8492 ;
  assign n8494 = n8493 ^ n5219 ^ n614 ;
  assign n8495 = ( ~n6071 & n8491 ) | ( ~n6071 & n8494 ) | ( n8491 & n8494 ) ;
  assign n8496 = n1644 | n2931 ;
  assign n8497 = n8496 ^ n1630 ^ 1'b0 ;
  assign n8498 = ( ~x45 & n2569 ) | ( ~x45 & n8497 ) | ( n2569 & n8497 ) ;
  assign n8499 = n203 & ~n8498 ;
  assign n8500 = n2860 & n8499 ;
  assign n8501 = n8500 ^ n6942 ^ 1'b0 ;
  assign n8502 = n8495 & n8501 ;
  assign n8504 = n3418 ^ n1368 ^ n190 ;
  assign n8505 = ( n259 & n4666 ) | ( n259 & ~n8504 ) | ( n4666 & ~n8504 ) ;
  assign n8506 = n7680 ^ n2486 ^ 1'b0 ;
  assign n8507 = n1331 & ~n8506 ;
  assign n8508 = ( n1718 & n5751 ) | ( n1718 & n8507 ) | ( n5751 & n8507 ) ;
  assign n8509 = ~n130 & n8508 ;
  assign n8510 = ~n8505 & n8509 ;
  assign n8503 = ~n5255 & n5454 ;
  assign n8511 = n8510 ^ n8503 ^ 1'b0 ;
  assign n8512 = n850 ^ n829 ^ 1'b0 ;
  assign n8513 = n8512 ^ n3302 ^ n3021 ;
  assign n8514 = n3131 | n7113 ;
  assign n8515 = n1929 | n5844 ;
  assign n8516 = n8515 ^ x12 ^ 1'b0 ;
  assign n8517 = n8516 ^ n4622 ^ 1'b0 ;
  assign n8518 = n8517 ^ n5469 ^ n4331 ;
  assign n8519 = n1430 & ~n5116 ;
  assign n8520 = ( ~n4329 & n5706 ) | ( ~n4329 & n8519 ) | ( n5706 & n8519 ) ;
  assign n8521 = ( n1255 & n3071 ) | ( n1255 & ~n3371 ) | ( n3071 & ~n3371 ) ;
  assign n8522 = n8521 ^ n7861 ^ 1'b0 ;
  assign n8523 = n3016 | n8522 ;
  assign n8528 = n6626 ^ n1152 ^ x88 ;
  assign n8529 = n5628 & ~n8528 ;
  assign n8524 = n2343 ^ n599 ^ 1'b0 ;
  assign n8525 = x25 & n8524 ;
  assign n8526 = n8525 ^ n3176 ^ 1'b0 ;
  assign n8527 = n1867 & n8526 ;
  assign n8530 = n8529 ^ n8527 ^ n8494 ;
  assign n8531 = n4065 ^ n2972 ^ 1'b0 ;
  assign n8532 = ( n4878 & ~n5578 ) | ( n4878 & n8531 ) | ( ~n5578 & n8531 ) ;
  assign n8533 = n3496 ^ n1265 ^ 1'b0 ;
  assign n8534 = n3011 & ~n8533 ;
  assign n8535 = n8534 ^ n2178 ^ 1'b0 ;
  assign n8536 = n1133 & ~n3383 ;
  assign n8537 = n8536 ^ n5296 ^ 1'b0 ;
  assign n8538 = n8537 ^ n2510 ^ n248 ;
  assign n8539 = n6731 | n7735 ;
  assign n8540 = n8539 ^ n3019 ^ 1'b0 ;
  assign n8544 = ( ~n468 & n4365 ) | ( ~n468 & n7381 ) | ( n4365 & n7381 ) ;
  assign n8545 = n8544 ^ n5153 ^ n4960 ;
  assign n8541 = n253 | n3942 ;
  assign n8542 = ~n4524 & n8541 ;
  assign n8543 = n8542 ^ n3191 ^ 1'b0 ;
  assign n8546 = n8545 ^ n8543 ^ n6241 ;
  assign n8547 = ( ~n8538 & n8540 ) | ( ~n8538 & n8546 ) | ( n8540 & n8546 ) ;
  assign n8548 = n3321 ^ n1086 ^ n1034 ;
  assign n8549 = n8300 & n8548 ;
  assign n8550 = n8549 ^ n8247 ^ 1'b0 ;
  assign n8551 = ( x1 & n5487 ) | ( x1 & ~n5714 ) | ( n5487 & ~n5714 ) ;
  assign n8552 = n2795 ^ n780 ^ 1'b0 ;
  assign n8553 = n750 & n8552 ;
  assign n8554 = ( ~n8550 & n8551 ) | ( ~n8550 & n8553 ) | ( n8551 & n8553 ) ;
  assign n8558 = n1515 ^ n734 ^ 1'b0 ;
  assign n8559 = ( n2282 & ~n6594 ) | ( n2282 & n8558 ) | ( ~n6594 & n8558 ) ;
  assign n8555 = n5294 ^ n4726 ^ n595 ;
  assign n8556 = ( n859 & ~n2697 ) | ( n859 & n5974 ) | ( ~n2697 & n5974 ) ;
  assign n8557 = ( n4496 & n8555 ) | ( n4496 & n8556 ) | ( n8555 & n8556 ) ;
  assign n8560 = n8559 ^ n8557 ^ n2689 ;
  assign n8566 = n1994 & ~n4137 ;
  assign n8561 = ~n2478 & n8452 ;
  assign n8562 = n8561 ^ n3851 ^ 1'b0 ;
  assign n8563 = n5387 ^ n4049 ^ 1'b0 ;
  assign n8564 = n8562 & ~n8563 ;
  assign n8565 = n7243 & n8564 ;
  assign n8567 = n8566 ^ n8565 ^ 1'b0 ;
  assign n8568 = n2723 ^ n1294 ^ 1'b0 ;
  assign n8569 = n582 | n8568 ;
  assign n8570 = n8569 ^ n5773 ^ n1953 ;
  assign n8571 = n8570 ^ n464 ^ 1'b0 ;
  assign n8572 = x31 & n8571 ;
  assign n8573 = ~n2834 & n8572 ;
  assign n8574 = n6989 ^ n4365 ^ 1'b0 ;
  assign n8575 = n5513 | n8574 ;
  assign n8576 = n5299 ^ n3273 ^ n711 ;
  assign n8577 = ( n1051 & n2091 ) | ( n1051 & n6261 ) | ( n2091 & n6261 ) ;
  assign n8578 = n8577 ^ n6807 ^ 1'b0 ;
  assign n8579 = n4555 & ~n8578 ;
  assign n8580 = n8579 ^ n1553 ^ 1'b0 ;
  assign n8584 = n2631 ^ n1327 ^ x88 ;
  assign n8581 = n2745 & ~n3299 ;
  assign n8582 = ~n3745 & n8581 ;
  assign n8583 = n8582 ^ n8505 ^ n3085 ;
  assign n8585 = n8584 ^ n8583 ^ 1'b0 ;
  assign n8586 = ( n6965 & ~n7285 ) | ( n6965 & n8585 ) | ( ~n7285 & n8585 ) ;
  assign n8587 = n5645 ^ n3724 ^ 1'b0 ;
  assign n8588 = n421 & ~n8587 ;
  assign n8589 = n8588 ^ n4712 ^ n4674 ;
  assign n8590 = n3924 & ~n3961 ;
  assign n8591 = n5962 ^ n1081 ^ 1'b0 ;
  assign n8592 = n3115 ^ n2745 ^ n160 ;
  assign n8593 = n3064 & n8592 ;
  assign n8594 = n8593 ^ n2819 ^ 1'b0 ;
  assign n8595 = n6918 | n8594 ;
  assign n8596 = n2843 ^ n1490 ^ 1'b0 ;
  assign n8597 = ( n966 & ~n1095 ) | ( n966 & n2423 ) | ( ~n1095 & n2423 ) ;
  assign n8598 = n8597 ^ n6648 ^ 1'b0 ;
  assign n8599 = n1514 & ~n8598 ;
  assign n8600 = n5807 & n8599 ;
  assign n8601 = ( n648 & n3433 ) | ( n648 & ~n3681 ) | ( n3433 & ~n3681 ) ;
  assign n8602 = n8389 & ~n8601 ;
  assign n8603 = n8602 ^ n6790 ^ n5269 ;
  assign n8604 = n4544 ^ n484 ^ 1'b0 ;
  assign n8605 = n4867 & ~n8604 ;
  assign n8606 = x57 & ~n8605 ;
  assign n8607 = n2615 ^ n531 ^ n235 ;
  assign n8608 = n8607 ^ n5177 ^ 1'b0 ;
  assign n8609 = n8606 | n8608 ;
  assign n8610 = ~n1430 & n7716 ;
  assign n8611 = n4652 & n8610 ;
  assign n8612 = n831 & ~n8611 ;
  assign n8613 = n610 & n8612 ;
  assign n8618 = ~n159 & n5696 ;
  assign n8619 = n8618 ^ n3961 ^ 1'b0 ;
  assign n8614 = n702 | n2746 ;
  assign n8615 = n2883 & ~n8614 ;
  assign n8616 = n8615 ^ n1096 ^ 1'b0 ;
  assign n8617 = n8616 ^ n2471 ^ n532 ;
  assign n8620 = n8619 ^ n8617 ^ 1'b0 ;
  assign n8621 = n2462 & n8620 ;
  assign n8623 = ( ~n1952 & n2492 ) | ( ~n1952 & n3826 ) | ( n2492 & n3826 ) ;
  assign n8622 = n214 & ~n238 ;
  assign n8624 = n8623 ^ n8622 ^ 1'b0 ;
  assign n8625 = n3409 ^ n2638 ^ n2441 ;
  assign n8626 = n6630 ^ n5262 ^ 1'b0 ;
  assign n8627 = ~n8625 & n8626 ;
  assign n8628 = ( n1247 & n2464 ) | ( n1247 & ~n2786 ) | ( n2464 & ~n2786 ) ;
  assign n8629 = n5748 ^ n5319 ^ 1'b0 ;
  assign n8630 = ( ~n380 & n4039 ) | ( ~n380 & n8629 ) | ( n4039 & n8629 ) ;
  assign n8631 = n4884 & ~n8630 ;
  assign n8632 = n7135 ^ n6626 ^ n628 ;
  assign n8633 = n6378 ^ n5507 ^ 1'b0 ;
  assign n8634 = n1859 ^ n1326 ^ 1'b0 ;
  assign n8635 = n962 & ~n8634 ;
  assign n8636 = ( n5563 & n8633 ) | ( n5563 & n8635 ) | ( n8633 & n8635 ) ;
  assign n8637 = ~n8632 & n8636 ;
  assign n8638 = ( n3088 & n4539 ) | ( n3088 & ~n6104 ) | ( n4539 & ~n6104 ) ;
  assign n8639 = n8139 ^ n5589 ^ n2978 ;
  assign n8640 = n380 & ~n7574 ;
  assign n8641 = n2346 ^ x13 ^ 1'b0 ;
  assign n8642 = n2220 & ~n8641 ;
  assign n8643 = n8640 | n8642 ;
  assign n8644 = ( n238 & ~n568 ) | ( n238 & n3443 ) | ( ~n568 & n3443 ) ;
  assign n8645 = n8644 ^ n2304 ^ 1'b0 ;
  assign n8646 = n5782 & ~n8645 ;
  assign n8648 = ( ~n1928 & n5900 ) | ( ~n1928 & n6008 ) | ( n5900 & n6008 ) ;
  assign n8647 = ( n4339 & n4985 ) | ( n4339 & n6319 ) | ( n4985 & n6319 ) ;
  assign n8649 = n8648 ^ n8647 ^ n3302 ;
  assign n8650 = n6837 ^ n2955 ^ 1'b0 ;
  assign n8651 = ~n441 & n3599 ;
  assign n8652 = n2644 ^ n309 ^ 1'b0 ;
  assign n8653 = n5165 ^ n2957 ^ n1882 ;
  assign n8654 = n8652 & ~n8653 ;
  assign n8655 = n8651 & n8654 ;
  assign n8656 = n200 & ~n1808 ;
  assign n8657 = ~n2994 & n8656 ;
  assign n8662 = n3289 ^ n887 ^ x28 ;
  assign n8663 = n8662 ^ n5262 ^ n3499 ;
  assign n8664 = n7732 & ~n8663 ;
  assign n8658 = n3653 ^ n2524 ^ n393 ;
  assign n8659 = ( n2510 & n6038 ) | ( n2510 & n8658 ) | ( n6038 & n8658 ) ;
  assign n8660 = ( n2985 & n4243 ) | ( n2985 & n8659 ) | ( n4243 & n8659 ) ;
  assign n8661 = n2564 & ~n8660 ;
  assign n8665 = n8664 ^ n8661 ^ 1'b0 ;
  assign n8666 = n2922 ^ n667 ^ n176 ;
  assign n8667 = n6643 ^ n5981 ^ 1'b0 ;
  assign n8668 = n8667 ^ n6354 ^ n2319 ;
  assign n8669 = n6695 ^ n2402 ^ 1'b0 ;
  assign n8670 = n386 & n8669 ;
  assign n8671 = n976 & ~n8118 ;
  assign n8672 = ~n8670 & n8671 ;
  assign n8673 = n2701 ^ n2213 ^ 1'b0 ;
  assign n8674 = n8673 ^ n5050 ^ n3299 ;
  assign n8675 = ~n418 & n8674 ;
  assign n8676 = ~n1016 & n4917 ;
  assign n8677 = n8676 ^ n244 ^ 1'b0 ;
  assign n8678 = n7402 ^ n6008 ^ n1079 ;
  assign n8679 = n8677 & ~n8678 ;
  assign n8680 = n8679 ^ n3167 ^ 1'b0 ;
  assign n8681 = n8680 ^ n4250 ^ n3207 ;
  assign n8682 = x1 & ~n8681 ;
  assign n8683 = n8682 ^ n5253 ^ 1'b0 ;
  assign n8684 = ( n3272 & ~n4976 ) | ( n3272 & n8491 ) | ( ~n4976 & n8491 ) ;
  assign n8685 = ( n7714 & n7921 ) | ( n7714 & n8684 ) | ( n7921 & n8684 ) ;
  assign n8686 = n2227 ^ n346 ^ 1'b0 ;
  assign n8687 = ( n2178 & ~n5516 ) | ( n2178 & n8135 ) | ( ~n5516 & n8135 ) ;
  assign n8688 = ( n4197 & n6802 ) | ( n4197 & ~n8687 ) | ( n6802 & ~n8687 ) ;
  assign n8689 = n8686 | n8688 ;
  assign n8690 = n7105 ^ n2210 ^ 1'b0 ;
  assign n8691 = n8690 ^ n2809 ^ 1'b0 ;
  assign n8692 = n8691 ^ n3742 ^ 1'b0 ;
  assign n8693 = n8692 ^ n5357 ^ n1791 ;
  assign n8694 = n8015 ^ n3161 ^ 1'b0 ;
  assign n8695 = n8693 | n8694 ;
  assign n8696 = ~n3362 & n5868 ;
  assign n8697 = n536 & n8696 ;
  assign n8698 = ( n205 & n3368 ) | ( n205 & ~n8697 ) | ( n3368 & ~n8697 ) ;
  assign n8699 = n3745 ^ n1154 ^ n376 ;
  assign n8700 = n8699 ^ n7518 ^ n4457 ;
  assign n8701 = n4721 ^ n1411 ^ n316 ;
  assign n8702 = n593 | n730 ;
  assign n8703 = n4045 | n8702 ;
  assign n8704 = ( n1407 & ~n8701 ) | ( n1407 & n8703 ) | ( ~n8701 & n8703 ) ;
  assign n8705 = n8704 ^ n8186 ^ n1501 ;
  assign n8707 = ( n1050 & n1750 ) | ( n1050 & ~n3297 ) | ( n1750 & ~n3297 ) ;
  assign n8706 = n5329 ^ n4265 ^ 1'b0 ;
  assign n8708 = n8707 ^ n8706 ^ n7498 ;
  assign n8714 = ( ~n1085 & n1510 ) | ( ~n1085 & n2301 ) | ( n1510 & n2301 ) ;
  assign n8710 = n1853 ^ n1208 ^ x67 ;
  assign n8711 = ( n235 & ~n1533 ) | ( n235 & n8710 ) | ( ~n1533 & n8710 ) ;
  assign n8712 = n2360 & n8711 ;
  assign n8709 = ( ~n3162 & n6160 ) | ( ~n3162 & n6893 ) | ( n6160 & n6893 ) ;
  assign n8713 = n8712 ^ n8709 ^ n6756 ;
  assign n8715 = n8714 ^ n8713 ^ 1'b0 ;
  assign n8716 = n8715 ^ n5292 ^ 1'b0 ;
  assign n8721 = n227 & ~n4440 ;
  assign n8718 = n3400 ^ n857 ^ 1'b0 ;
  assign n8719 = n5126 ^ n2284 ^ 1'b0 ;
  assign n8720 = ~n8718 & n8719 ;
  assign n8717 = n8395 ^ n3359 ^ n1343 ;
  assign n8722 = n8721 ^ n8720 ^ n8717 ;
  assign n8723 = n7394 ^ n5008 ^ n415 ;
  assign n8724 = n8723 ^ n3985 ^ n3681 ;
  assign n8725 = n8619 ^ n6827 ^ 1'b0 ;
  assign n8726 = n2968 & ~n3212 ;
  assign n8727 = n2286 & n8726 ;
  assign n8728 = n8725 & n8727 ;
  assign n8729 = ( n2455 & ~n3273 ) | ( n2455 & n8138 ) | ( ~n3273 & n8138 ) ;
  assign n8730 = ( n2195 & ~n4287 ) | ( n2195 & n5920 ) | ( ~n4287 & n5920 ) ;
  assign n8731 = n8729 | n8730 ;
  assign n8732 = n8731 ^ n6136 ^ 1'b0 ;
  assign n8733 = n1295 | n8732 ;
  assign n8734 = n7585 ^ n1411 ^ 1'b0 ;
  assign n8735 = n8734 ^ n3337 ^ n690 ;
  assign n8742 = n3016 | n4098 ;
  assign n8743 = n8742 ^ n4157 ^ 1'b0 ;
  assign n8736 = ~n966 & n2607 ;
  assign n8737 = n8736 ^ n6939 ^ 1'b0 ;
  assign n8738 = ( n2703 & n3068 ) | ( n2703 & ~n4196 ) | ( n3068 & ~n4196 ) ;
  assign n8739 = ~n8737 & n8738 ;
  assign n8740 = n8739 ^ n459 ^ 1'b0 ;
  assign n8741 = n427 & n8740 ;
  assign n8744 = n8743 ^ n8741 ^ 1'b0 ;
  assign n8745 = n4337 ^ n4334 ^ n3726 ;
  assign n8746 = n8745 ^ n6992 ^ 1'b0 ;
  assign n8747 = ~n362 & n2804 ;
  assign n8748 = n8747 ^ n3689 ^ 1'b0 ;
  assign n8749 = n8748 ^ n5161 ^ 1'b0 ;
  assign n8750 = n8749 ^ n5751 ^ n5296 ;
  assign n8751 = ( n620 & ~n1084 ) | ( n620 & n8427 ) | ( ~n1084 & n8427 ) ;
  assign n8752 = n2100 & n8751 ;
  assign n8753 = ( n1431 & n3408 ) | ( n1431 & n8407 ) | ( n3408 & n8407 ) ;
  assign n8754 = n8753 ^ n3579 ^ n3058 ;
  assign n8755 = n8754 ^ n5668 ^ n4098 ;
  assign n8756 = n6508 ^ n5116 ^ 1'b0 ;
  assign n8758 = n4230 & ~n8139 ;
  assign n8757 = n8109 ^ n5197 ^ 1'b0 ;
  assign n8759 = n8758 ^ n8757 ^ n4003 ;
  assign n8760 = ( n3593 & ~n8091 ) | ( n3593 & n8759 ) | ( ~n8091 & n8759 ) ;
  assign n8761 = ~n3345 & n4286 ;
  assign n8762 = ( n5408 & ~n5464 ) | ( n5408 & n8761 ) | ( ~n5464 & n8761 ) ;
  assign n8763 = n4440 ^ n3816 ^ 1'b0 ;
  assign n8764 = ( n4717 & ~n6218 ) | ( n4717 & n8763 ) | ( ~n6218 & n8763 ) ;
  assign n8765 = n6891 ^ n6487 ^ 1'b0 ;
  assign n8766 = ( n1228 & n1331 ) | ( n1228 & ~n8765 ) | ( n1331 & ~n8765 ) ;
  assign n8767 = n3629 ^ n1876 ^ n422 ;
  assign n8768 = n8767 ^ n7747 ^ 1'b0 ;
  assign n8769 = n8766 & ~n8768 ;
  assign n8770 = ( n3206 & n3764 ) | ( n3206 & n6472 ) | ( n3764 & n6472 ) ;
  assign n8771 = n7780 ^ n6978 ^ n746 ;
  assign n8772 = ( ~n386 & n7551 ) | ( ~n386 & n8771 ) | ( n7551 & n8771 ) ;
  assign n8773 = n8772 ^ n2242 ^ n1856 ;
  assign n8774 = n8773 ^ n6983 ^ n4822 ;
  assign n8775 = n3227 ^ n792 ^ 1'b0 ;
  assign n8776 = n8775 ^ n5142 ^ n1895 ;
  assign n8777 = n8776 ^ n7596 ^ 1'b0 ;
  assign n8778 = n7356 ^ n4039 ^ n1789 ;
  assign n8779 = ( x72 & ~n821 ) | ( x72 & n4736 ) | ( ~n821 & n4736 ) ;
  assign n8780 = n8779 ^ n1371 ^ 1'b0 ;
  assign n8781 = ( n7780 & n8778 ) | ( n7780 & ~n8780 ) | ( n8778 & ~n8780 ) ;
  assign n8782 = n7411 & n8781 ;
  assign n8793 = n3678 ^ n1460 ^ 1'b0 ;
  assign n8794 = n8793 ^ n456 ^ 1'b0 ;
  assign n8791 = n156 & ~n2904 ;
  assign n8792 = ( n1164 & n7637 ) | ( n1164 & ~n8791 ) | ( n7637 & ~n8791 ) ;
  assign n8795 = n8794 ^ n8792 ^ n5225 ;
  assign n8787 = ~n2440 & n6001 ;
  assign n8788 = n8787 ^ x121 ^ 1'b0 ;
  assign n8789 = n3245 & n7911 ;
  assign n8790 = n8788 & ~n8789 ;
  assign n8783 = ( n442 & n760 ) | ( n442 & n1366 ) | ( n760 & n1366 ) ;
  assign n8784 = n264 | n5728 ;
  assign n8785 = n8783 & ~n8784 ;
  assign n8786 = ~n7599 & n8785 ;
  assign n8796 = n8795 ^ n8790 ^ n8786 ;
  assign n8797 = n376 & n3264 ;
  assign n8798 = n8797 ^ n2218 ^ 1'b0 ;
  assign n8799 = n8592 ^ n8443 ^ n2429 ;
  assign n8800 = n4445 & n6703 ;
  assign n8801 = n2058 ^ n131 ^ 1'b0 ;
  assign n8802 = ( n1145 & n2935 ) | ( n1145 & n5602 ) | ( n2935 & n5602 ) ;
  assign n8803 = ~n5247 & n8683 ;
  assign n8804 = n8802 & n8803 ;
  assign n8805 = n3362 | n4000 ;
  assign n8806 = n1063 & ~n8805 ;
  assign n8807 = n1356 & n8806 ;
  assign n8808 = n8807 ^ n964 ^ 1'b0 ;
  assign n8809 = n6763 ^ n2950 ^ n1463 ;
  assign n8810 = ( n3263 & n6580 ) | ( n3263 & ~n8809 ) | ( n6580 & ~n8809 ) ;
  assign n8811 = n1809 ^ n1523 ^ 1'b0 ;
  assign n8812 = n8811 ^ x99 ^ 1'b0 ;
  assign n8813 = ( n1022 & n2567 ) | ( n1022 & ~n8812 ) | ( n2567 & ~n8812 ) ;
  assign n8816 = n926 & ~n2515 ;
  assign n8815 = n4287 & n4559 ;
  assign n8817 = n8816 ^ n8815 ^ 1'b0 ;
  assign n8814 = n8301 ^ n5487 ^ n3647 ;
  assign n8818 = n8817 ^ n8814 ^ n3653 ;
  assign n8819 = n3513 & n7663 ;
  assign n8820 = ( n4831 & ~n5637 ) | ( n4831 & n7146 ) | ( ~n5637 & n7146 ) ;
  assign n8821 = n1190 & ~n7023 ;
  assign n8822 = ~n2638 & n8821 ;
  assign n8823 = ( ~n886 & n8820 ) | ( ~n886 & n8822 ) | ( n8820 & n8822 ) ;
  assign n8824 = ~n263 & n6123 ;
  assign n8825 = n8824 ^ n413 ^ 1'b0 ;
  assign n8827 = n6116 ^ n4040 ^ n2633 ;
  assign n8826 = n629 & n6842 ;
  assign n8828 = n8827 ^ n8826 ^ 1'b0 ;
  assign n8829 = n8828 ^ n5981 ^ n3598 ;
  assign n8830 = ( n8476 & ~n8825 ) | ( n8476 & n8829 ) | ( ~n8825 & n8829 ) ;
  assign n8831 = n8096 ^ n6105 ^ n4943 ;
  assign n8834 = n2513 ^ n1146 ^ n828 ;
  assign n8832 = n4045 ^ n3203 ^ 1'b0 ;
  assign n8833 = ~n2982 & n8832 ;
  assign n8835 = n8834 ^ n8833 ^ n1790 ;
  assign n8836 = n4497 | n8835 ;
  assign n8837 = n8831 | n8836 ;
  assign n8838 = n5686 ^ n3602 ^ n3089 ;
  assign n8839 = ( ~n6383 & n8037 ) | ( ~n6383 & n8283 ) | ( n8037 & n8283 ) ;
  assign n8840 = n1912 | n5470 ;
  assign n8841 = n6510 & ~n8840 ;
  assign n8842 = n5145 & ~n7396 ;
  assign n8843 = n8842 ^ n6409 ^ n915 ;
  assign n8844 = ( n3386 & n6881 ) | ( n3386 & ~n8843 ) | ( n6881 & ~n8843 ) ;
  assign n8845 = n6891 ^ n3622 ^ 1'b0 ;
  assign n8846 = n8844 & ~n8845 ;
  assign n8847 = ~n2026 & n4423 ;
  assign n8848 = n1828 | n2578 ;
  assign n8849 = n3743 | n8848 ;
  assign n8850 = ( ~n2117 & n3115 ) | ( ~n2117 & n8849 ) | ( n3115 & n8849 ) ;
  assign n8851 = ( ~n3605 & n8847 ) | ( ~n3605 & n8850 ) | ( n8847 & n8850 ) ;
  assign n8854 = n3272 ^ n1169 ^ n1034 ;
  assign n8852 = n7753 ^ n2393 ^ 1'b0 ;
  assign n8853 = n8852 ^ n5607 ^ n2611 ;
  assign n8855 = n8854 ^ n8853 ^ 1'b0 ;
  assign n8856 = ( n636 & n2980 ) | ( n636 & n8855 ) | ( n2980 & n8855 ) ;
  assign n8858 = n253 & ~n4109 ;
  assign n8859 = n8858 ^ n4951 ^ 1'b0 ;
  assign n8857 = n8183 ^ n4276 ^ n1718 ;
  assign n8860 = n8859 ^ n8857 ^ n5105 ;
  assign n8861 = n3020 ^ n294 ^ 1'b0 ;
  assign n8862 = n8861 ^ n5695 ^ 1'b0 ;
  assign n8863 = ( n734 & n6812 ) | ( n734 & n7064 ) | ( n6812 & n7064 ) ;
  assign n8864 = n1699 & n8656 ;
  assign n8865 = n8370 & n8864 ;
  assign n8866 = ( ~n165 & n1011 ) | ( ~n165 & n4644 ) | ( n1011 & n4644 ) ;
  assign n8867 = n5686 ^ n3413 ^ 1'b0 ;
  assign n8868 = n1069 | n3122 ;
  assign n8869 = n8868 ^ n7420 ^ n2799 ;
  assign n8870 = ( n1232 & n3395 ) | ( n1232 & n3762 ) | ( n3395 & n3762 ) ;
  assign n8871 = n8870 ^ n5385 ^ 1'b0 ;
  assign n8872 = n8869 & n8871 ;
  assign n8873 = n572 & n1459 ;
  assign n8877 = n2726 ^ n1375 ^ 1'b0 ;
  assign n8874 = n5487 | n7816 ;
  assign n8875 = n8874 ^ x106 ^ 1'b0 ;
  assign n8876 = n8875 ^ n2893 ^ n1343 ;
  assign n8878 = n8877 ^ n8876 ^ 1'b0 ;
  assign n8879 = n8878 ^ n2435 ^ 1'b0 ;
  assign n8880 = ~n1003 & n8879 ;
  assign n8881 = n6393 ^ n3577 ^ 1'b0 ;
  assign n8882 = n8448 ^ n4500 ^ n1262 ;
  assign n8883 = n8882 ^ n5595 ^ n698 ;
  assign n8884 = ( n3872 & n4960 ) | ( n3872 & n8883 ) | ( n4960 & n8883 ) ;
  assign n8885 = n5476 & n7326 ;
  assign n8886 = n2150 ^ n951 ^ n760 ;
  assign n8887 = n8886 ^ n3230 ^ 1'b0 ;
  assign n8888 = ~n1946 & n8887 ;
  assign n8889 = ( n1239 & ~n1650 ) | ( n1239 & n8888 ) | ( ~n1650 & n8888 ) ;
  assign n8890 = n4070 & n8889 ;
  assign n8891 = ~n5384 & n8890 ;
  assign n8892 = n8713 ^ n5836 ^ n5006 ;
  assign n8893 = n5419 ^ n2499 ^ 1'b0 ;
  assign n8894 = n4132 & ~n8893 ;
  assign n8895 = ( n3791 & ~n8247 ) | ( n3791 & n8894 ) | ( ~n8247 & n8894 ) ;
  assign n8898 = n3882 ^ n576 ^ 1'b0 ;
  assign n8899 = n3980 & ~n8898 ;
  assign n8900 = n8899 ^ n1823 ^ 1'b0 ;
  assign n8896 = n5356 ^ n2922 ^ n1346 ;
  assign n8897 = ~n1301 & n8896 ;
  assign n8901 = n8900 ^ n8897 ^ 1'b0 ;
  assign n8902 = ( n985 & n8895 ) | ( n985 & n8901 ) | ( n8895 & n8901 ) ;
  assign n8903 = n4170 ^ n490 ^ 1'b0 ;
  assign n8904 = n8902 & n8903 ;
  assign n8905 = n2616 & ~n7130 ;
  assign n8906 = ~x122 & n4882 ;
  assign n8909 = n1800 ^ n955 ^ 1'b0 ;
  assign n8910 = n1294 & ~n8909 ;
  assign n8911 = ( n1834 & n4213 ) | ( n1834 & n8910 ) | ( n4213 & n8910 ) ;
  assign n8907 = n3858 & ~n4918 ;
  assign n8908 = n8907 ^ n6495 ^ 1'b0 ;
  assign n8912 = n8911 ^ n8908 ^ 1'b0 ;
  assign n8913 = n6650 & ~n8912 ;
  assign n8916 = x40 & n4820 ;
  assign n8914 = n6780 ^ n236 ^ 1'b0 ;
  assign n8915 = n8914 ^ n4571 ^ n3179 ;
  assign n8917 = n8916 ^ n8915 ^ n3947 ;
  assign n8920 = n7828 ^ n3363 ^ 1'b0 ;
  assign n8918 = n2907 ^ x3 ^ 1'b0 ;
  assign n8919 = n8918 ^ n3722 ^ n1683 ;
  assign n8921 = n8920 ^ n8919 ^ n2255 ;
  assign n8922 = n1046 | n3819 ;
  assign n8923 = n8922 ^ n2481 ^ n2069 ;
  assign n8924 = n3329 | n8923 ;
  assign n8925 = n8924 ^ n7274 ^ 1'b0 ;
  assign n8926 = n7715 ^ n3491 ^ n2713 ;
  assign n8927 = n4404 & n8926 ;
  assign n8928 = ( ~n8921 & n8925 ) | ( ~n8921 & n8927 ) | ( n8925 & n8927 ) ;
  assign n8929 = n7806 | n8746 ;
  assign n8930 = n4351 ^ n4070 ^ n3742 ;
  assign n8931 = n6981 ^ n2998 ^ n499 ;
  assign n8932 = n3201 ^ n3084 ^ 1'b0 ;
  assign n8933 = n7134 & n8932 ;
  assign n8934 = n8933 ^ n1203 ^ 1'b0 ;
  assign n8935 = n8934 ^ n6992 ^ 1'b0 ;
  assign n8936 = n8931 & n8935 ;
  assign n8937 = n1791 & n3064 ;
  assign n8938 = n8936 & n8937 ;
  assign n8940 = n4693 ^ n3125 ^ 1'b0 ;
  assign n8941 = n990 & ~n8940 ;
  assign n8939 = n796 & n5932 ;
  assign n8942 = n8941 ^ n8939 ^ 1'b0 ;
  assign n8943 = ( n504 & n6404 ) | ( n504 & n8635 ) | ( n6404 & n8635 ) ;
  assign n8944 = n8943 ^ n3564 ^ n2887 ;
  assign n8959 = n2576 | n6739 ;
  assign n8960 = ( n1578 & ~n4114 ) | ( n1578 & n8959 ) | ( ~n4114 & n8959 ) ;
  assign n8954 = n7180 ^ n2234 ^ 1'b0 ;
  assign n8955 = n5186 & n8954 ;
  assign n8956 = ~n2062 & n8955 ;
  assign n8957 = n8956 ^ n1373 ^ 1'b0 ;
  assign n8953 = n4272 & n5105 ;
  assign n8958 = n8957 ^ n8953 ^ 1'b0 ;
  assign n8945 = n1558 | n2495 ;
  assign n8946 = n2059 ^ n1272 ^ n575 ;
  assign n8947 = ( ~n3571 & n7107 ) | ( ~n3571 & n8946 ) | ( n7107 & n8946 ) ;
  assign n8948 = n4017 ^ n1445 ^ 1'b0 ;
  assign n8949 = ~x68 & n3349 ;
  assign n8950 = ~n8948 & n8949 ;
  assign n8951 = ( ~n1697 & n4402 ) | ( ~n1697 & n8950 ) | ( n4402 & n8950 ) ;
  assign n8952 = ( n8945 & n8947 ) | ( n8945 & ~n8951 ) | ( n8947 & ~n8951 ) ;
  assign n8961 = n8960 ^ n8958 ^ n8952 ;
  assign n8962 = ( n1411 & n8944 ) | ( n1411 & n8961 ) | ( n8944 & n8961 ) ;
  assign n8963 = n3280 & n6113 ;
  assign n8964 = n5699 & n7396 ;
  assign n8965 = x9 & n6397 ;
  assign n8966 = n8964 & n8965 ;
  assign n8967 = n1036 & ~n3917 ;
  assign n8968 = ( n1243 & ~n5486 ) | ( n1243 & n8967 ) | ( ~n5486 & n8967 ) ;
  assign n8972 = n2494 | n5494 ;
  assign n8973 = n8972 ^ n6750 ^ 1'b0 ;
  assign n8969 = n2906 & ~n4405 ;
  assign n8970 = n3975 & n8969 ;
  assign n8971 = ( n831 & n971 ) | ( n831 & ~n8970 ) | ( n971 & ~n8970 ) ;
  assign n8974 = n8973 ^ n8971 ^ n399 ;
  assign n8975 = n4075 ^ n1393 ^ n999 ;
  assign n8976 = n6053 ^ n4408 ^ 1'b0 ;
  assign n8977 = n8975 & n8976 ;
  assign n8978 = n8977 ^ n7180 ^ n722 ;
  assign n8979 = n8978 ^ n6089 ^ n1483 ;
  assign n8982 = ~n691 & n1447 ;
  assign n8983 = n8982 ^ n665 ^ 1'b0 ;
  assign n8984 = n2638 & ~n8983 ;
  assign n8985 = n1220 & n8984 ;
  assign n8980 = n4191 ^ n1706 ^ n1247 ;
  assign n8981 = n6282 | n8980 ;
  assign n8986 = n8985 ^ n8981 ^ 1'b0 ;
  assign n8987 = n4715 | n8986 ;
  assign n8988 = ( n4719 & n6693 ) | ( n4719 & n7286 ) | ( n6693 & n7286 ) ;
  assign n8991 = n2843 ^ n2498 ^ 1'b0 ;
  assign n8992 = n2612 & n8991 ;
  assign n8989 = ( x85 & ~n3981 ) | ( x85 & n8973 ) | ( ~n3981 & n8973 ) ;
  assign n8990 = n2911 | n8989 ;
  assign n8993 = n8992 ^ n8990 ^ 1'b0 ;
  assign n8994 = n322 & ~n7183 ;
  assign n8995 = ( n1439 & ~n4202 ) | ( n1439 & n8994 ) | ( ~n4202 & n8994 ) ;
  assign n8996 = n2234 ^ n2081 ^ 1'b0 ;
  assign n8997 = n2181 ^ n1136 ^ 1'b0 ;
  assign n8998 = n368 & ~n8997 ;
  assign n8999 = n8996 | n8998 ;
  assign n9000 = ( n875 & ~n1695 ) | ( n875 & n2428 ) | ( ~n1695 & n2428 ) ;
  assign n9001 = ( n3092 & n8334 ) | ( n3092 & ~n9000 ) | ( n8334 & ~n9000 ) ;
  assign n9002 = ( n4467 & n6883 ) | ( n4467 & ~n9001 ) | ( n6883 & ~n9001 ) ;
  assign n9004 = n6128 ^ n5308 ^ 1'b0 ;
  assign n9005 = x126 & ~n9004 ;
  assign n9006 = n2553 ^ n927 ^ 1'b0 ;
  assign n9007 = n500 & ~n9006 ;
  assign n9008 = ~n9005 & n9007 ;
  assign n9003 = n7141 ^ n3151 ^ 1'b0 ;
  assign n9009 = n9008 ^ n9003 ^ n1269 ;
  assign n9010 = ( ~n1599 & n2111 ) | ( ~n1599 & n3958 ) | ( n2111 & n3958 ) ;
  assign n9011 = n3115 ^ n2346 ^ 1'b0 ;
  assign n9012 = n9010 & n9011 ;
  assign n9013 = n3312 ^ n1989 ^ 1'b0 ;
  assign n9014 = n5024 | n9013 ;
  assign n9015 = n7780 ^ n7425 ^ n2911 ;
  assign n9016 = x79 | n9015 ;
  assign n9017 = n5358 | n9016 ;
  assign n9018 = n3588 & n9017 ;
  assign n9019 = n9018 ^ n4190 ^ 1'b0 ;
  assign n9020 = n2043 & n3341 ;
  assign n9023 = n896 & n2445 ;
  assign n9021 = x120 & ~n302 ;
  assign n9022 = n9021 ^ n1364 ^ 1'b0 ;
  assign n9024 = n9023 ^ n9022 ^ n6675 ;
  assign n9025 = ( ~n4451 & n9020 ) | ( ~n4451 & n9024 ) | ( n9020 & n9024 ) ;
  assign n9026 = ( ~n2837 & n5447 ) | ( ~n2837 & n8097 ) | ( n5447 & n8097 ) ;
  assign n9027 = n6366 ^ n1182 ^ 1'b0 ;
  assign n9028 = n2312 | n4026 ;
  assign n9029 = n9028 ^ n8642 ^ 1'b0 ;
  assign n9030 = ~n2461 & n5116 ;
  assign n9031 = n9030 ^ n2539 ^ n894 ;
  assign n9032 = n4491 ^ n2065 ^ 1'b0 ;
  assign n9033 = n3407 & ~n9032 ;
  assign n9034 = ~n9031 & n9033 ;
  assign n9035 = x18 & ~n379 ;
  assign n9036 = n9035 ^ n2120 ^ 1'b0 ;
  assign n9037 = n2498 ^ n1707 ^ 1'b0 ;
  assign n9038 = n5542 | n9037 ;
  assign n9039 = n5922 & ~n9038 ;
  assign n9040 = n9036 & ~n9039 ;
  assign n9041 = ~n9034 & n9040 ;
  assign n9042 = n5059 ^ n542 ^ 1'b0 ;
  assign n9043 = n7454 ^ n5380 ^ n2718 ;
  assign n9044 = n6792 & ~n9043 ;
  assign n9045 = n9044 ^ n183 ^ 1'b0 ;
  assign n9046 = ( n7325 & n9042 ) | ( n7325 & ~n9045 ) | ( n9042 & ~n9045 ) ;
  assign n9047 = ~n6289 & n7733 ;
  assign n9048 = n9046 & n9047 ;
  assign n9049 = n4033 ^ n2291 ^ n388 ;
  assign n9050 = n234 & n9049 ;
  assign n9051 = ( x46 & ~n199 ) | ( x46 & n4363 ) | ( ~n199 & n4363 ) ;
  assign n9052 = ~n1053 & n6121 ;
  assign n9053 = n6828 ^ n5969 ^ 1'b0 ;
  assign n9054 = n1294 & n5881 ;
  assign n9055 = ~n2160 & n9054 ;
  assign n9065 = n8996 ^ n5607 ^ 1'b0 ;
  assign n9066 = n9065 ^ n620 ^ 1'b0 ;
  assign n9067 = ~n555 & n9066 ;
  assign n9057 = ( n2272 & n6504 ) | ( n2272 & ~n6765 ) | ( n6504 & ~n6765 ) ;
  assign n9056 = n6124 & ~n7038 ;
  assign n9058 = n9057 ^ n9056 ^ 1'b0 ;
  assign n9059 = n635 & ~n6543 ;
  assign n9060 = ~n378 & n9059 ;
  assign n9061 = n9060 ^ n3031 ^ 1'b0 ;
  assign n9062 = n9061 ^ n1720 ^ x124 ;
  assign n9063 = n601 & ~n9062 ;
  assign n9064 = n9058 & n9063 ;
  assign n9068 = n9067 ^ n9064 ^ 1'b0 ;
  assign n9069 = n2304 ^ n1758 ^ n386 ;
  assign n9070 = ( x5 & n424 ) | ( x5 & ~n9069 ) | ( n424 & ~n9069 ) ;
  assign n9071 = ( ~x0 & n1375 ) | ( ~x0 & n9070 ) | ( n1375 & n9070 ) ;
  assign n9072 = ( ~n1452 & n8759 ) | ( ~n1452 & n9071 ) | ( n8759 & n9071 ) ;
  assign n9073 = n6481 ^ n4028 ^ 1'b0 ;
  assign n9074 = ~n4677 & n9073 ;
  assign n9075 = n2178 & ~n3645 ;
  assign n9076 = n6506 & n9075 ;
  assign n9077 = ~n2167 & n9076 ;
  assign n9078 = ( ~n2964 & n9074 ) | ( ~n2964 & n9077 ) | ( n9074 & n9077 ) ;
  assign n9082 = ( n2135 & n3291 ) | ( n2135 & n4128 ) | ( n3291 & n4128 ) ;
  assign n9079 = ~n6586 & n8461 ;
  assign n9080 = ( n5377 & n6541 ) | ( n5377 & ~n8439 ) | ( n6541 & ~n8439 ) ;
  assign n9081 = ( n7793 & ~n9079 ) | ( n7793 & n9080 ) | ( ~n9079 & n9080 ) ;
  assign n9083 = n9082 ^ n9081 ^ 1'b0 ;
  assign n9084 = n9078 & ~n9083 ;
  assign n9085 = x14 & n654 ;
  assign n9086 = n9085 ^ n2289 ^ 1'b0 ;
  assign n9087 = ( ~n2293 & n8507 ) | ( ~n2293 & n9086 ) | ( n8507 & n9086 ) ;
  assign n9088 = ( n4572 & n8164 ) | ( n4572 & ~n9087 ) | ( n8164 & ~n9087 ) ;
  assign n9089 = n5335 & ~n9088 ;
  assign n9090 = n9089 ^ n7948 ^ 1'b0 ;
  assign n9091 = ~n1517 & n5421 ;
  assign n9092 = n9091 ^ n1621 ^ 1'b0 ;
  assign n9093 = ~n2291 & n4535 ;
  assign n9094 = ( ~n2844 & n3451 ) | ( ~n2844 & n9093 ) | ( n3451 & n9093 ) ;
  assign n9095 = n1451 | n2568 ;
  assign n9096 = n9095 ^ n2256 ^ 1'b0 ;
  assign n9097 = n2252 & n6307 ;
  assign n9098 = n1291 & n9097 ;
  assign n9099 = n9098 ^ n2196 ^ 1'b0 ;
  assign n9100 = ~n9096 & n9099 ;
  assign n9101 = n9100 ^ n8420 ^ 1'b0 ;
  assign n9102 = ~n7454 & n9101 ;
  assign n9103 = ( n9092 & ~n9094 ) | ( n9092 & n9102 ) | ( ~n9094 & n9102 ) ;
  assign n9104 = ( n2598 & n3541 ) | ( n2598 & ~n3886 ) | ( n3541 & ~n3886 ) ;
  assign n9105 = n8300 ^ n2842 ^ x49 ;
  assign n9106 = n9105 ^ n4414 ^ n209 ;
  assign n9107 = ( n705 & ~n4158 ) | ( n705 & n5198 ) | ( ~n4158 & n5198 ) ;
  assign n9108 = n6937 ^ n2867 ^ x101 ;
  assign n9109 = ( n4059 & n9107 ) | ( n4059 & n9108 ) | ( n9107 & n9108 ) ;
  assign n9110 = n9109 ^ n7847 ^ n6312 ;
  assign n9111 = ( n9104 & ~n9106 ) | ( n9104 & n9110 ) | ( ~n9106 & n9110 ) ;
  assign n9112 = n3864 | n9111 ;
  assign n9128 = n6312 ^ n1418 ^ n1294 ;
  assign n9129 = n9128 ^ n1126 ^ x66 ;
  assign n9124 = ( n6236 & n6460 ) | ( n6236 & n7433 ) | ( n6460 & n7433 ) ;
  assign n9122 = n3814 ^ n3499 ^ 1'b0 ;
  assign n9123 = ~n4974 & n9122 ;
  assign n9125 = n9124 ^ n9123 ^ 1'b0 ;
  assign n9113 = n586 | n1394 ;
  assign n9114 = n357 | n9113 ;
  assign n9115 = n9114 ^ n4734 ^ 1'b0 ;
  assign n9119 = ( n1474 & n2866 ) | ( n1474 & ~n6937 ) | ( n2866 & ~n6937 ) ;
  assign n9116 = n5045 ^ n4727 ^ n3339 ;
  assign n9117 = ( n646 & ~n1577 ) | ( n646 & n9116 ) | ( ~n1577 & n9116 ) ;
  assign n9118 = ( n1419 & ~n1945 ) | ( n1419 & n9117 ) | ( ~n1945 & n9117 ) ;
  assign n9120 = n9119 ^ n9118 ^ 1'b0 ;
  assign n9121 = n9115 | n9120 ;
  assign n9126 = n9125 ^ n9121 ^ n2753 ;
  assign n9127 = n5790 & ~n9126 ;
  assign n9130 = n9129 ^ n9127 ^ 1'b0 ;
  assign n9131 = ( n3920 & n4188 ) | ( n3920 & n8475 ) | ( n4188 & n8475 ) ;
  assign n9132 = n5624 & n6638 ;
  assign n9133 = ~n9131 & n9132 ;
  assign n9134 = n1362 ^ n829 ^ n549 ;
  assign n9135 = n9134 ^ n5526 ^ n3987 ;
  assign n9136 = ~n6624 & n9135 ;
  assign n9137 = n9136 ^ n372 ^ 1'b0 ;
  assign n9139 = n1688 & ~n3115 ;
  assign n9140 = n9139 ^ n6354 ^ 1'b0 ;
  assign n9138 = ( n2692 & n4176 ) | ( n2692 & n6671 ) | ( n4176 & n6671 ) ;
  assign n9141 = n9140 ^ n9138 ^ n3541 ;
  assign n9142 = ( n326 & n7167 ) | ( n326 & ~n9141 ) | ( n7167 & ~n9141 ) ;
  assign n9150 = n2789 | n8424 ;
  assign n9151 = n5121 | n9150 ;
  assign n9152 = n4574 & n9151 ;
  assign n9153 = n9152 ^ n1608 ^ 1'b0 ;
  assign n9143 = ~n2445 & n2772 ;
  assign n9144 = n9143 ^ n5145 ^ 1'b0 ;
  assign n9145 = n832 & n6495 ;
  assign n9146 = ( n4694 & ~n9144 ) | ( n4694 & n9145 ) | ( ~n9144 & n9145 ) ;
  assign n9147 = n9146 ^ n2116 ^ 1'b0 ;
  assign n9148 = n9147 ^ n6149 ^ n2314 ;
  assign n9149 = ~n7274 & n9148 ;
  assign n9154 = n9153 ^ n9149 ^ 1'b0 ;
  assign n9161 = ~n3275 & n3964 ;
  assign n9162 = n9161 ^ n1073 ^ 1'b0 ;
  assign n9163 = n9162 ^ n6729 ^ n1899 ;
  assign n9160 = n2426 | n3858 ;
  assign n9156 = n7254 ^ n5364 ^ 1'b0 ;
  assign n9157 = n762 & ~n9156 ;
  assign n9155 = n7680 ^ n6606 ^ n2142 ;
  assign n9158 = n9157 ^ n9155 ^ n2703 ;
  assign n9159 = ( ~n2982 & n7074 ) | ( ~n2982 & n9158 ) | ( n7074 & n9158 ) ;
  assign n9164 = n9163 ^ n9160 ^ n9159 ;
  assign n9173 = ( n1943 & n2847 ) | ( n1943 & ~n8183 ) | ( n2847 & ~n8183 ) ;
  assign n9174 = n275 | n1118 ;
  assign n9175 = n9173 | n9174 ;
  assign n9176 = ~n4375 & n9175 ;
  assign n9177 = ( n1132 & n3688 ) | ( n1132 & n9176 ) | ( n3688 & n9176 ) ;
  assign n9166 = n2020 ^ n222 ^ 1'b0 ;
  assign n9167 = n1320 & n9166 ;
  assign n9165 = ( ~n2500 & n3188 ) | ( ~n2500 & n4390 ) | ( n3188 & n4390 ) ;
  assign n9168 = n9167 ^ n9165 ^ n1513 ;
  assign n9169 = n314 & ~n3336 ;
  assign n9170 = ( n449 & ~n2418 ) | ( n449 & n9169 ) | ( ~n2418 & n9169 ) ;
  assign n9171 = ( n4281 & n9168 ) | ( n4281 & n9170 ) | ( n9168 & n9170 ) ;
  assign n9172 = n9171 ^ n6976 ^ 1'b0 ;
  assign n9178 = n9177 ^ n9172 ^ 1'b0 ;
  assign n9179 = n5175 | n9178 ;
  assign n9180 = n4650 & ~n6766 ;
  assign n9181 = ~n2507 & n9180 ;
  assign n9182 = n5545 & n6424 ;
  assign n9183 = ~n4970 & n9182 ;
  assign n9184 = n9181 | n9183 ;
  assign n9188 = n3552 & n3698 ;
  assign n9189 = n9188 ^ n4384 ^ 1'b0 ;
  assign n9185 = n6814 ^ n2342 ^ 1'b0 ;
  assign n9186 = n6236 & ~n9185 ;
  assign n9187 = n9186 ^ n4511 ^ 1'b0 ;
  assign n9190 = n9189 ^ n9187 ^ n1307 ;
  assign n9191 = n2747 ^ n2323 ^ x76 ;
  assign n9192 = n6999 | n9191 ;
  assign n9193 = n1318 | n9192 ;
  assign n9194 = n728 | n4500 ;
  assign n9195 = n9194 ^ n3461 ^ 1'b0 ;
  assign n9196 = n2992 & ~n9195 ;
  assign n9197 = n9196 ^ n2081 ^ 1'b0 ;
  assign n9198 = n9197 ^ n3740 ^ n1197 ;
  assign n9199 = n9193 & ~n9198 ;
  assign n9200 = n821 & ~n4019 ;
  assign n9201 = n3830 & n9200 ;
  assign n9202 = n9201 ^ n8964 ^ 1'b0 ;
  assign n9203 = n1894 ^ x19 ^ 1'b0 ;
  assign n9204 = n266 & ~n9203 ;
  assign n9205 = n4896 & n9204 ;
  assign n9206 = n2381 ^ n2023 ^ n1326 ;
  assign n9207 = n8619 | n9206 ;
  assign n9208 = ( n6505 & n7311 ) | ( n6505 & ~n9207 ) | ( n7311 & ~n9207 ) ;
  assign n9209 = ( ~n4601 & n9205 ) | ( ~n4601 & n9208 ) | ( n9205 & n9208 ) ;
  assign n9210 = n6957 ^ n1775 ^ n1725 ;
  assign n9211 = n9210 ^ n4522 ^ 1'b0 ;
  assign n9212 = n4115 & n9211 ;
  assign n9213 = ( ~n7227 & n8202 ) | ( ~n7227 & n9212 ) | ( n8202 & n9212 ) ;
  assign n9214 = n2636 & ~n9031 ;
  assign n9215 = ~n4501 & n8716 ;
  assign n9216 = ~n5894 & n9215 ;
  assign n9223 = n3687 ^ n2954 ^ n1208 ;
  assign n9224 = n9223 ^ n4445 ^ n1266 ;
  assign n9218 = x103 & ~n6862 ;
  assign n9219 = n9218 ^ n2795 ^ 1'b0 ;
  assign n9220 = n9219 ^ n5151 ^ n729 ;
  assign n9221 = n9220 ^ n4793 ^ n171 ;
  assign n9217 = n5464 ^ n2219 ^ n1856 ;
  assign n9222 = n9221 ^ n9217 ^ 1'b0 ;
  assign n9225 = n9224 ^ n9222 ^ 1'b0 ;
  assign n9226 = n1308 & n4235 ;
  assign n9227 = n9226 ^ n7382 ^ 1'b0 ;
  assign n9228 = n2175 & ~n3784 ;
  assign n9229 = ~n5102 & n9228 ;
  assign n9230 = n505 & ~n9229 ;
  assign n9231 = n4511 ^ n3877 ^ n2016 ;
  assign n9232 = ( n3138 & n5486 ) | ( n3138 & ~n8054 ) | ( n5486 & ~n8054 ) ;
  assign n9233 = n2198 | n8659 ;
  assign n9235 = n1257 & n2721 ;
  assign n9236 = n9235 ^ n1049 ^ 1'b0 ;
  assign n9237 = n9236 ^ n4905 ^ n1280 ;
  assign n9234 = x65 & n7641 ;
  assign n9238 = n9237 ^ n9234 ^ 1'b0 ;
  assign n9239 = n7362 ^ n4846 ^ n559 ;
  assign n9240 = ( n1702 & n5010 ) | ( n1702 & n5196 ) | ( n5010 & n5196 ) ;
  assign n9241 = n9240 ^ n9045 ^ n6706 ;
  assign n9242 = ( ~n2949 & n3589 ) | ( ~n2949 & n4538 ) | ( n3589 & n4538 ) ;
  assign n9243 = n9242 ^ n906 ^ 1'b0 ;
  assign n9244 = n2922 ^ n2739 ^ 1'b0 ;
  assign n9245 = n4002 ^ n2109 ^ n838 ;
  assign n9246 = ( n2823 & ~n4594 ) | ( n2823 & n9245 ) | ( ~n4594 & n9245 ) ;
  assign n9247 = n734 ^ n197 ^ 1'b0 ;
  assign n9248 = n2029 & n9247 ;
  assign n9249 = ~n2638 & n9248 ;
  assign n9250 = ( n1854 & n4020 ) | ( n1854 & n4429 ) | ( n4020 & n4429 ) ;
  assign n9251 = ( n3706 & n7144 ) | ( n3706 & n9250 ) | ( n7144 & n9250 ) ;
  assign n9252 = n2674 ^ n595 ^ 1'b0 ;
  assign n9258 = ( n130 & n481 ) | ( n130 & ~n1693 ) | ( n481 & ~n1693 ) ;
  assign n9259 = n9258 ^ n871 ^ 1'b0 ;
  assign n9260 = ( n2470 & ~n3312 ) | ( n2470 & n9259 ) | ( ~n3312 & n9259 ) ;
  assign n9257 = ~n765 & n1191 ;
  assign n9261 = n9260 ^ n9257 ^ n582 ;
  assign n9262 = n9261 ^ n5548 ^ x39 ;
  assign n9253 = ( ~n447 & n2314 ) | ( ~n447 & n3407 ) | ( n2314 & n3407 ) ;
  assign n9254 = ~n3329 & n9253 ;
  assign n9255 = n3610 & n9254 ;
  assign n9256 = n5139 | n9255 ;
  assign n9263 = n9262 ^ n9256 ^ 1'b0 ;
  assign n9264 = n5127 ^ n3912 ^ n504 ;
  assign n9265 = n9264 ^ n7108 ^ n4550 ;
  assign n9269 = n5522 ^ n872 ^ 1'b0 ;
  assign n9270 = ~n2631 & n9269 ;
  assign n9266 = ~n1424 & n4643 ;
  assign n9267 = ~x73 & n9266 ;
  assign n9268 = n7743 | n9267 ;
  assign n9271 = n9270 ^ n9268 ^ 1'b0 ;
  assign n9272 = n5054 ^ n1659 ^ x82 ;
  assign n9273 = n1281 & n9272 ;
  assign n9274 = ( n2167 & n8605 ) | ( n2167 & n9273 ) | ( n8605 & n9273 ) ;
  assign n9275 = ( n1989 & n3016 ) | ( n1989 & ~n4134 ) | ( n3016 & ~n4134 ) ;
  assign n9277 = n7107 ^ n2037 ^ n1456 ;
  assign n9278 = n6409 ^ n4098 ^ 1'b0 ;
  assign n9279 = ~n9277 & n9278 ;
  assign n9276 = n5698 ^ n3269 ^ x47 ;
  assign n9280 = n9279 ^ n9276 ^ n4250 ;
  assign n9281 = n1843 & ~n2513 ;
  assign n9282 = ~n5931 & n9281 ;
  assign n9283 = n9282 ^ n6818 ^ 1'b0 ;
  assign n9285 = ( ~n2259 & n2738 ) | ( ~n2259 & n4271 ) | ( n2738 & n4271 ) ;
  assign n9284 = n9141 ^ n5674 ^ x80 ;
  assign n9286 = n9285 ^ n9284 ^ n7100 ;
  assign n9287 = n9286 ^ n6021 ^ 1'b0 ;
  assign n9288 = n9283 | n9287 ;
  assign n9289 = n5166 ^ n3491 ^ 1'b0 ;
  assign n9290 = n7814 & ~n9289 ;
  assign n9291 = n4180 & ~n9290 ;
  assign n9292 = n4408 ^ n880 ^ 1'b0 ;
  assign n9293 = n4207 ^ n698 ^ 1'b0 ;
  assign n9294 = n2094 & n9293 ;
  assign n9295 = ~n4084 & n9294 ;
  assign n9296 = n9295 ^ n8473 ^ 1'b0 ;
  assign n9297 = n8320 ^ n7734 ^ n2549 ;
  assign n9298 = ( ~n2671 & n8926 ) | ( ~n2671 & n9297 ) | ( n8926 & n9297 ) ;
  assign n9299 = n7798 ^ n3378 ^ 1'b0 ;
  assign n9300 = n3977 ^ n652 ^ 1'b0 ;
  assign n9301 = n5595 & ~n9300 ;
  assign n9302 = n4282 ^ n275 ^ 1'b0 ;
  assign n9303 = n626 & n4278 ;
  assign n9304 = n9303 ^ n9073 ^ n7876 ;
  assign n9305 = n2307 | n4288 ;
  assign n9306 = n9305 ^ n1226 ^ n976 ;
  assign n9307 = ( n5605 & n8028 ) | ( n5605 & n9306 ) | ( n8028 & n9306 ) ;
  assign n9308 = ~n275 & n648 ;
  assign n9309 = n9308 ^ n8689 ^ 1'b0 ;
  assign n9310 = n4712 | n5018 ;
  assign n9311 = n9310 ^ n4213 ^ 1'b0 ;
  assign n9313 = n1539 ^ n814 ^ n187 ;
  assign n9312 = n7049 ^ n3083 ^ n2765 ;
  assign n9314 = n9313 ^ n9312 ^ 1'b0 ;
  assign n9315 = ~n8111 & n9314 ;
  assign n9316 = ~n360 & n6265 ;
  assign n9317 = n4140 & n9316 ;
  assign n9318 = n5277 & n9317 ;
  assign n9319 = n1149 & n2403 ;
  assign n9320 = ~n5279 & n9319 ;
  assign n9324 = n1452 ^ n878 ^ 1'b0 ;
  assign n9321 = n1826 ^ n1344 ^ 1'b0 ;
  assign n9322 = n1687 | n9321 ;
  assign n9323 = n9322 ^ n7008 ^ n646 ;
  assign n9325 = n9324 ^ n9323 ^ n4198 ;
  assign n9326 = n9259 & ~n9325 ;
  assign n9327 = n9326 ^ n8406 ^ 1'b0 ;
  assign n9328 = n1986 & ~n9327 ;
  assign n9329 = n7173 ^ n6955 ^ 1'b0 ;
  assign n9330 = n8955 & n9329 ;
  assign n9331 = n1839 ^ n1171 ^ 1'b0 ;
  assign n9332 = n9331 ^ n1982 ^ n1636 ;
  assign n9333 = n5592 ^ n5411 ^ 1'b0 ;
  assign n9334 = n9332 | n9333 ;
  assign n9342 = n6690 ^ n2795 ^ n984 ;
  assign n9339 = n4971 ^ n431 ^ 1'b0 ;
  assign n9340 = n2861 & ~n9339 ;
  assign n9341 = n9340 ^ n223 ^ 1'b0 ;
  assign n9335 = n5323 ^ n1025 ^ 1'b0 ;
  assign n9336 = n9335 ^ n4813 ^ n3493 ;
  assign n9337 = n5529 & ~n9336 ;
  assign n9338 = n9337 ^ n8716 ^ 1'b0 ;
  assign n9343 = n9342 ^ n9341 ^ n9338 ;
  assign n9346 = ( n1828 & ~n3077 ) | ( n1828 & n3268 ) | ( ~n3077 & n3268 ) ;
  assign n9347 = ( n1339 & n6624 ) | ( n1339 & ~n9346 ) | ( n6624 & ~n9346 ) ;
  assign n9344 = n2094 | n3087 ;
  assign n9345 = n9344 ^ n5178 ^ n4636 ;
  assign n9348 = n9347 ^ n9345 ^ n3213 ;
  assign n9350 = n5965 ^ n5095 ^ n2175 ;
  assign n9349 = ( n1095 & ~n1456 ) | ( n1095 & n2045 ) | ( ~n1456 & n2045 ) ;
  assign n9351 = n9350 ^ n9349 ^ n2016 ;
  assign n9352 = n6551 ^ n1803 ^ n989 ;
  assign n9353 = n9352 ^ n8379 ^ 1'b0 ;
  assign n9354 = n9353 ^ n4162 ^ 1'b0 ;
  assign n9355 = n3370 | n9354 ;
  assign n9356 = n3887 ^ n1580 ^ n1232 ;
  assign n9357 = n9356 ^ n7114 ^ 1'b0 ;
  assign n9358 = ( n2595 & n3695 ) | ( n2595 & ~n9357 ) | ( n3695 & ~n9357 ) ;
  assign n9359 = n9358 ^ n2845 ^ 1'b0 ;
  assign n9360 = ( ~n1533 & n3123 ) | ( ~n1533 & n9359 ) | ( n3123 & n9359 ) ;
  assign n9362 = n7722 ^ n5158 ^ n731 ;
  assign n9363 = n9362 ^ n635 ^ 1'b0 ;
  assign n9364 = n9363 ^ n5558 ^ n1666 ;
  assign n9361 = n5332 ^ n4016 ^ n2495 ;
  assign n9365 = n9364 ^ n9361 ^ n2682 ;
  assign n9366 = ( ~n1903 & n3044 ) | ( ~n1903 & n7399 ) | ( n3044 & n7399 ) ;
  assign n9367 = n9366 ^ n6038 ^ 1'b0 ;
  assign n9368 = n9367 ^ n4414 ^ 1'b0 ;
  assign n9369 = n967 & n6735 ;
  assign n9370 = n9369 ^ n1025 ^ 1'b0 ;
  assign n9371 = n4479 | n7848 ;
  assign n9372 = n9371 ^ n7596 ^ 1'b0 ;
  assign n9373 = n9370 | n9372 ;
  assign n9374 = n3322 & n5346 ;
  assign n9375 = n6885 ^ n6363 ^ n454 ;
  assign n9376 = n3595 ^ n3289 ^ 1'b0 ;
  assign n9377 = n1332 & n9376 ;
  assign n9378 = n8783 ^ n2787 ^ n1168 ;
  assign n9379 = n3326 ^ n1380 ^ n1078 ;
  assign n9380 = n9378 & ~n9379 ;
  assign n9381 = n9377 & n9380 ;
  assign n9382 = n2983 ^ n674 ^ n622 ;
  assign n9383 = n5552 & n9382 ;
  assign n9384 = n7712 ^ n3370 ^ n2582 ;
  assign n9385 = n3858 ^ x98 ^ 1'b0 ;
  assign n9386 = n8758 | n9385 ;
  assign n9387 = ( n2837 & n4458 ) | ( n2837 & ~n9098 ) | ( n4458 & ~n9098 ) ;
  assign n9388 = n9387 ^ n618 ^ 1'b0 ;
  assign n9389 = n4377 & ~n9388 ;
  assign n9390 = n8888 ^ n8415 ^ n2685 ;
  assign n9391 = ( n1145 & n7897 ) | ( n1145 & ~n8219 ) | ( n7897 & ~n8219 ) ;
  assign n9392 = n9391 ^ n1711 ^ 1'b0 ;
  assign n9393 = n717 & ~n4644 ;
  assign n9394 = n9393 ^ n923 ^ 1'b0 ;
  assign n9395 = ~n2245 & n9394 ;
  assign n9396 = ( ~n667 & n5799 ) | ( ~n667 & n9395 ) | ( n5799 & n9395 ) ;
  assign n9398 = n5934 ^ n5357 ^ 1'b0 ;
  assign n9399 = n1457 | n9398 ;
  assign n9397 = ( ~n2276 & n2911 ) | ( ~n2276 & n4578 ) | ( n2911 & n4578 ) ;
  assign n9400 = n9399 ^ n9397 ^ n1421 ;
  assign n9401 = n3263 & n9263 ;
  assign n9402 = n9401 ^ n8672 ^ 1'b0 ;
  assign n9403 = n8172 ^ n4307 ^ n2478 ;
  assign n9404 = ~n927 & n9403 ;
  assign n9405 = ( n1583 & ~n3300 ) | ( n1583 & n5660 ) | ( ~n3300 & n5660 ) ;
  assign n9413 = ( n2277 & ~n3227 ) | ( n2277 & n4946 ) | ( ~n3227 & n4946 ) ;
  assign n9406 = n1093 | n1312 ;
  assign n9407 = n1602 & ~n9406 ;
  assign n9408 = ( n3070 & ~n9021 ) | ( n3070 & n9407 ) | ( ~n9021 & n9407 ) ;
  assign n9409 = ( n2606 & n2847 ) | ( n2606 & n9408 ) | ( n2847 & n9408 ) ;
  assign n9410 = ~n2310 & n5870 ;
  assign n9411 = n9410 ^ n4702 ^ 1'b0 ;
  assign n9412 = ( ~n6161 & n9409 ) | ( ~n6161 & n9411 ) | ( n9409 & n9411 ) ;
  assign n9414 = n9413 ^ n9412 ^ n8983 ;
  assign n9415 = ( n9404 & n9405 ) | ( n9404 & n9414 ) | ( n9405 & n9414 ) ;
  assign n9417 = ( n2349 & n2706 ) | ( n2349 & n3484 ) | ( n2706 & n3484 ) ;
  assign n9416 = n1741 | n3698 ;
  assign n9418 = n9417 ^ n9416 ^ n1664 ;
  assign n9419 = n6747 ^ n4900 ^ 1'b0 ;
  assign n9420 = n8389 & ~n9419 ;
  assign n9421 = ~n645 & n3747 ;
  assign n9422 = ~n3710 & n9421 ;
  assign n9423 = n2547 | n9422 ;
  assign n9424 = n2063 & ~n9423 ;
  assign n9425 = n7928 ^ n1865 ^ 1'b0 ;
  assign n9426 = n1871 ^ n1567 ^ 1'b0 ;
  assign n9427 = n883 & ~n9426 ;
  assign n9428 = n5579 | n9427 ;
  assign n9429 = n5425 & ~n7584 ;
  assign n9430 = n7288 & n9429 ;
  assign n9431 = ( ~n271 & n1737 ) | ( ~n271 & n7276 ) | ( n1737 & n7276 ) ;
  assign n9432 = n9431 ^ n8861 ^ 1'b0 ;
  assign n9433 = ( n1304 & n2808 ) | ( n1304 & n9432 ) | ( n2808 & n9432 ) ;
  assign n9434 = n3889 ^ n903 ^ n466 ;
  assign n9435 = ( n1828 & ~n2157 ) | ( n1828 & n4677 ) | ( ~n2157 & n4677 ) ;
  assign n9436 = n6957 ^ n2249 ^ n435 ;
  assign n9437 = ( n4065 & n9435 ) | ( n4065 & n9436 ) | ( n9435 & n9436 ) ;
  assign n9438 = ( n3716 & ~n9434 ) | ( n3716 & n9437 ) | ( ~n9434 & n9437 ) ;
  assign n9439 = n2746 ^ n1797 ^ 1'b0 ;
  assign n9440 = n5120 & n9439 ;
  assign n9441 = n3457 | n9440 ;
  assign n9442 = n1050 ^ n490 ^ 1'b0 ;
  assign n9443 = n1038 | n4721 ;
  assign n9444 = n340 & ~n9443 ;
  assign n9445 = n3619 | n9444 ;
  assign n9446 = n9445 ^ n6404 ^ 1'b0 ;
  assign n9447 = ~n1268 & n6091 ;
  assign n9448 = ~x119 & n9447 ;
  assign n9449 = ( n5105 & n9446 ) | ( n5105 & n9448 ) | ( n9446 & n9448 ) ;
  assign n9450 = ~n2038 & n3648 ;
  assign n9451 = ~n9449 & n9450 ;
  assign n9452 = n1012 ^ n865 ^ 1'b0 ;
  assign n9453 = n4834 & n9452 ;
  assign n9454 = n9451 & n9453 ;
  assign n9455 = n9260 ^ n3405 ^ n2723 ;
  assign n9456 = n6277 ^ n1818 ^ 1'b0 ;
  assign n9457 = n1994 ^ n197 ^ 1'b0 ;
  assign n9458 = n420 | n9457 ;
  assign n9459 = n5627 & ~n9458 ;
  assign n9460 = n9459 ^ n8582 ^ 1'b0 ;
  assign n9461 = n538 & ~n2247 ;
  assign n9462 = ( n307 & n3534 ) | ( n307 & ~n8151 ) | ( n3534 & ~n8151 ) ;
  assign n9463 = n9461 & n9462 ;
  assign n9464 = n8523 & n9463 ;
  assign n9465 = ( n991 & n3335 ) | ( n991 & ~n3720 ) | ( n3335 & ~n3720 ) ;
  assign n9466 = ( n3272 & n4077 ) | ( n3272 & n9465 ) | ( n4077 & n9465 ) ;
  assign n9467 = ~n8343 & n9466 ;
  assign n9468 = n9467 ^ n4555 ^ n244 ;
  assign n9469 = n2543 ^ n2422 ^ 1'b0 ;
  assign n9470 = ( ~n2620 & n3379 ) | ( ~n2620 & n9469 ) | ( n3379 & n9469 ) ;
  assign n9471 = n9470 ^ n5702 ^ n2397 ;
  assign n9472 = n3031 & n3963 ;
  assign n9473 = n931 & n9472 ;
  assign n9474 = n9473 ^ n5770 ^ 1'b0 ;
  assign n9475 = ( ~n7249 & n9471 ) | ( ~n7249 & n9474 ) | ( n9471 & n9474 ) ;
  assign n9478 = ~n2837 & n7714 ;
  assign n9479 = n9478 ^ n4640 ^ n481 ;
  assign n9476 = n8421 ^ n2105 ^ 1'b0 ;
  assign n9477 = n5709 & n9476 ;
  assign n9480 = n9479 ^ n9477 ^ n6889 ;
  assign n9481 = n7121 & n9409 ;
  assign n9482 = n7272 & ~n9481 ;
  assign n9483 = n9482 ^ x23 ^ 1'b0 ;
  assign n9484 = n759 | n4407 ;
  assign n9485 = ( n2787 & n6187 ) | ( n2787 & n9205 ) | ( n6187 & n9205 ) ;
  assign n9486 = n9485 ^ n705 ^ 1'b0 ;
  assign n9487 = n7126 & ~n7348 ;
  assign n9488 = x12 & ~n1914 ;
  assign n9491 = ( n476 & n1592 ) | ( n476 & ~n2710 ) | ( n1592 & ~n2710 ) ;
  assign n9489 = n2131 ^ x118 ^ 1'b0 ;
  assign n9490 = n3232 | n9489 ;
  assign n9492 = n9491 ^ n9490 ^ n6055 ;
  assign n9493 = n5011 ^ n2932 ^ n2641 ;
  assign n9494 = n3816 & n4956 ;
  assign n9495 = ~n9493 & n9494 ;
  assign n9496 = ( n1228 & n7608 ) | ( n1228 & n9495 ) | ( n7608 & n9495 ) ;
  assign n9497 = n5589 ^ n2314 ^ n2021 ;
  assign n9498 = n8444 & ~n9361 ;
  assign n9499 = n9497 & n9498 ;
  assign n9500 = ( n712 & n2108 ) | ( n712 & ~n5288 ) | ( n2108 & ~n5288 ) ;
  assign n9501 = n9134 ^ n6385 ^ 1'b0 ;
  assign n9505 = ~n404 & n1409 ;
  assign n9506 = n9505 ^ n2165 ^ 1'b0 ;
  assign n9507 = n9506 ^ n2051 ^ n593 ;
  assign n9503 = n964 ^ n931 ^ 1'b0 ;
  assign n9502 = n1475 & n3981 ;
  assign n9504 = n9503 ^ n9502 ^ 1'b0 ;
  assign n9508 = n9507 ^ n9504 ^ n5249 ;
  assign n9509 = n1805 | n2337 ;
  assign n9511 = n4228 ^ n3044 ^ n2470 ;
  assign n9512 = n3163 & n9511 ;
  assign n9513 = n9512 ^ n4230 ^ 1'b0 ;
  assign n9510 = n4997 | n8465 ;
  assign n9514 = n9513 ^ n9510 ^ 1'b0 ;
  assign n9515 = ~n790 & n3047 ;
  assign n9516 = ( n971 & n8711 ) | ( n971 & n9515 ) | ( n8711 & n9515 ) ;
  assign n9517 = n9516 ^ n2777 ^ 1'b0 ;
  assign n9518 = ~n3381 & n9517 ;
  assign n9519 = ~n6716 & n9518 ;
  assign n9520 = ( n330 & n8331 ) | ( n330 & ~n9519 ) | ( n8331 & ~n9519 ) ;
  assign n9521 = ( ~n1677 & n3402 ) | ( ~n1677 & n5352 ) | ( n3402 & n5352 ) ;
  assign n9522 = n763 & n2819 ;
  assign n9523 = n9522 ^ n4682 ^ 1'b0 ;
  assign n9524 = n8635 ^ n6092 ^ n477 ;
  assign n9527 = n1483 ^ x23 ^ 1'b0 ;
  assign n9528 = ~n131 & n9527 ;
  assign n9529 = n863 & ~n3799 ;
  assign n9530 = ~n9528 & n9529 ;
  assign n9525 = n227 | n7223 ;
  assign n9526 = n9525 ^ n6025 ^ 1'b0 ;
  assign n9531 = n9530 ^ n9526 ^ n7633 ;
  assign n9532 = n4695 ^ n3190 ^ 1'b0 ;
  assign n9533 = ( n429 & n605 ) | ( n429 & ~n9532 ) | ( n605 & ~n9532 ) ;
  assign n9534 = n9533 ^ n4283 ^ n2745 ;
  assign n9535 = n9534 ^ n6992 ^ n6046 ;
  assign n9536 = ( n4846 & n5320 ) | ( n4846 & ~n6718 ) | ( n5320 & ~n6718 ) ;
  assign n9537 = n9536 ^ n760 ^ 1'b0 ;
  assign n9538 = n3234 ^ n3160 ^ n2798 ;
  assign n9539 = n5757 & n9538 ;
  assign n9540 = ( ~x31 & n223 ) | ( ~x31 & n9539 ) | ( n223 & n9539 ) ;
  assign n9541 = n9540 ^ n8164 ^ 1'b0 ;
  assign n9542 = ~n311 & n2242 ;
  assign n9543 = ( n5681 & n5708 ) | ( n5681 & ~n6001 ) | ( n5708 & ~n6001 ) ;
  assign n9544 = ~n1285 & n9543 ;
  assign n9545 = n3011 ^ x17 ^ 1'b0 ;
  assign n9546 = n1759 | n1907 ;
  assign n9547 = n9546 ^ n2077 ^ 1'b0 ;
  assign n9548 = n4739 | n9547 ;
  assign n9549 = n9548 ^ n561 ^ 1'b0 ;
  assign n9550 = n4011 & n9549 ;
  assign n9551 = ~n9545 & n9550 ;
  assign n9552 = n492 & ~n2109 ;
  assign n9553 = n9552 ^ n1859 ^ 1'b0 ;
  assign n9554 = ( n2842 & n7001 ) | ( n2842 & ~n9553 ) | ( n7001 & ~n9553 ) ;
  assign n9555 = n7233 & n9554 ;
  assign n9556 = n9555 ^ n8175 ^ 1'b0 ;
  assign n9561 = ~n136 & n6369 ;
  assign n9562 = ( n1388 & ~n4666 ) | ( n1388 & n6690 ) | ( ~n4666 & n6690 ) ;
  assign n9563 = ( ~n929 & n3379 ) | ( ~n929 & n9562 ) | ( n3379 & n9562 ) ;
  assign n9564 = n9563 ^ n1442 ^ 1'b0 ;
  assign n9565 = n9561 & ~n9564 ;
  assign n9566 = ~n6304 & n9565 ;
  assign n9567 = ~n3359 & n9566 ;
  assign n9558 = n1107 | n7107 ;
  assign n9557 = n3377 & n8175 ;
  assign n9559 = n9558 ^ n9557 ^ 1'b0 ;
  assign n9560 = ( n1419 & n9466 ) | ( n1419 & n9559 ) | ( n9466 & n9559 ) ;
  assign n9568 = n9567 ^ n9560 ^ n1899 ;
  assign n9569 = ~n8303 & n9568 ;
  assign n9571 = n7680 ^ n4294 ^ 1'b0 ;
  assign n9570 = ( ~x15 & n2163 ) | ( ~x15 & n5324 ) | ( n2163 & n5324 ) ;
  assign n9572 = n9571 ^ n9570 ^ n4404 ;
  assign n9573 = ( n198 & n743 ) | ( n198 & n2506 ) | ( n743 & n2506 ) ;
  assign n9574 = n9573 ^ n2527 ^ 1'b0 ;
  assign n9575 = ~n5150 & n9574 ;
  assign n9576 = n3269 & n9575 ;
  assign n9577 = ~n3317 & n9576 ;
  assign n9578 = n9577 ^ n7074 ^ 1'b0 ;
  assign n9579 = n2805 & n3846 ;
  assign n9580 = n9413 ^ n3882 ^ 1'b0 ;
  assign n9581 = ( ~n1472 & n5021 ) | ( ~n1472 & n9580 ) | ( n5021 & n9580 ) ;
  assign n9582 = ( ~n9339 & n9579 ) | ( ~n9339 & n9581 ) | ( n9579 & n9581 ) ;
  assign n9583 = ( n4924 & ~n7789 ) | ( n4924 & n9039 ) | ( ~n7789 & n9039 ) ;
  assign n9588 = n2334 ^ n954 ^ 1'b0 ;
  assign n9589 = n1018 | n1521 ;
  assign n9590 = n9588 & ~n9589 ;
  assign n9591 = n9590 ^ n3303 ^ n2281 ;
  assign n9586 = n2902 & n7596 ;
  assign n9587 = n9586 ^ n8644 ^ 1'b0 ;
  assign n9592 = n9591 ^ n9587 ^ 1'b0 ;
  assign n9593 = n4691 & ~n9592 ;
  assign n9594 = n1788 & n1915 ;
  assign n9595 = ( n1369 & n3920 ) | ( n1369 & ~n9594 ) | ( n3920 & ~n9594 ) ;
  assign n9596 = n8668 & n9595 ;
  assign n9597 = ~n9593 & n9596 ;
  assign n9584 = ( n2212 & n3705 ) | ( n2212 & ~n3820 ) | ( n3705 & ~n3820 ) ;
  assign n9585 = ( n7441 & n7776 ) | ( n7441 & n9584 ) | ( n7776 & n9584 ) ;
  assign n9598 = n9597 ^ n9585 ^ n4096 ;
  assign n9599 = ( n2679 & n3815 ) | ( n2679 & ~n9515 ) | ( n3815 & ~n9515 ) ;
  assign n9600 = n3706 ^ n2827 ^ 1'b0 ;
  assign n9601 = n1493 & ~n5157 ;
  assign n9602 = n9601 ^ n1107 ^ 1'b0 ;
  assign n9603 = n1516 & n9602 ;
  assign n9604 = n9600 & n9603 ;
  assign n9605 = n1557 ^ n1317 ^ n508 ;
  assign n9606 = ~n7858 & n9605 ;
  assign n9610 = n7229 ^ n3804 ^ 1'b0 ;
  assign n9611 = ~n3084 & n9610 ;
  assign n9607 = n1568 ^ n1399 ^ n162 ;
  assign n9608 = n3412 & n9607 ;
  assign n9609 = ~n6128 & n9608 ;
  assign n9612 = n9611 ^ n9609 ^ n6140 ;
  assign n9613 = n9612 ^ n729 ^ 1'b0 ;
  assign n9614 = n4956 & n9613 ;
  assign n9615 = n9614 ^ n5460 ^ 1'b0 ;
  assign n9616 = ( n5066 & ~n6510 ) | ( n5066 & n6731 ) | ( ~n6510 & n6731 ) ;
  assign n9617 = n4882 | n8640 ;
  assign n9618 = n9617 ^ n2337 ^ n1427 ;
  assign n9619 = ~n9616 & n9618 ;
  assign n9621 = n543 ^ n157 ^ 1'b0 ;
  assign n9622 = n2179 & ~n9621 ;
  assign n9623 = n9622 ^ n2247 ^ n265 ;
  assign n9620 = ~n4152 & n8199 ;
  assign n9624 = n9623 ^ n9620 ^ 1'b0 ;
  assign n9625 = n1984 & n3217 ;
  assign n9626 = n9625 ^ n7003 ^ 1'b0 ;
  assign n9627 = ( n2691 & ~n4629 ) | ( n2691 & n4684 ) | ( ~n4629 & n4684 ) ;
  assign n9628 = n9627 ^ n3640 ^ n2596 ;
  assign n9629 = ( ~n3098 & n9561 ) | ( ~n3098 & n9628 ) | ( n9561 & n9628 ) ;
  assign n9630 = n6159 ^ n2002 ^ n866 ;
  assign n9631 = ( n1767 & n1917 ) | ( n1767 & ~n9630 ) | ( n1917 & ~n9630 ) ;
  assign n9632 = ( n1955 & n2754 ) | ( n1955 & ~n9631 ) | ( n2754 & ~n9631 ) ;
  assign n9633 = n9632 ^ n6862 ^ 1'b0 ;
  assign n9634 = n9629 & n9633 ;
  assign n9635 = ( ~n3414 & n9626 ) | ( ~n3414 & n9634 ) | ( n9626 & n9634 ) ;
  assign n9636 = n3579 ^ n1361 ^ 1'b0 ;
  assign n9642 = ( n450 & ~n3565 ) | ( n450 & n7639 ) | ( ~n3565 & n7639 ) ;
  assign n9640 = n4729 ^ n2615 ^ n1143 ;
  assign n9641 = n9640 ^ n6066 ^ 1'b0 ;
  assign n9637 = n7425 ^ n4544 ^ n2901 ;
  assign n9638 = n9637 ^ n2967 ^ n1346 ;
  assign n9639 = n9638 ^ n4271 ^ 1'b0 ;
  assign n9643 = n9642 ^ n9641 ^ n9639 ;
  assign n9649 = n1748 ^ n1191 ^ 1'b0 ;
  assign n9650 = ~n4107 & n9649 ;
  assign n9647 = n2571 ^ n1284 ^ 1'b0 ;
  assign n9648 = n2413 & n9647 ;
  assign n9651 = n9650 ^ n9648 ^ 1'b0 ;
  assign n9645 = ( n4616 & n4837 ) | ( n4616 & n5969 ) | ( n4837 & n5969 ) ;
  assign n9644 = ~n772 & n4363 ;
  assign n9646 = n9645 ^ n9644 ^ 1'b0 ;
  assign n9652 = n9651 ^ n9646 ^ 1'b0 ;
  assign n9653 = n5932 & ~n9652 ;
  assign n9654 = n1918 & n3433 ;
  assign n9655 = n9654 ^ n2289 ^ 1'b0 ;
  assign n9656 = n6207 & n9655 ;
  assign n9657 = n7427 ^ n3065 ^ 1'b0 ;
  assign n9658 = ( ~n8997 & n9656 ) | ( ~n8997 & n9657 ) | ( n9656 & n9657 ) ;
  assign n9659 = ( n4103 & n4535 ) | ( n4103 & ~n7006 ) | ( n4535 & ~n7006 ) ;
  assign n9660 = n6257 ^ n3522 ^ 1'b0 ;
  assign n9661 = n7564 ^ n6482 ^ n3138 ;
  assign n9662 = ( ~n6765 & n9660 ) | ( ~n6765 & n9661 ) | ( n9660 & n9661 ) ;
  assign n9663 = ( n5108 & n9659 ) | ( n5108 & n9662 ) | ( n9659 & n9662 ) ;
  assign n9664 = n9098 ^ n5854 ^ n4148 ;
  assign n9665 = ~n8272 & n9664 ;
  assign n9666 = n9665 ^ n1633 ^ 1'b0 ;
  assign n9667 = n9204 ^ n4701 ^ n1100 ;
  assign n9671 = n6989 ^ n1668 ^ 1'b0 ;
  assign n9672 = ~n2919 & n9671 ;
  assign n9673 = n6057 ^ n5686 ^ 1'b0 ;
  assign n9674 = n9672 & ~n9673 ;
  assign n9668 = ( n1210 & ~n4815 ) | ( n1210 & n8931 ) | ( ~n4815 & n8931 ) ;
  assign n9669 = ( n1418 & ~n9016 ) | ( n1418 & n9668 ) | ( ~n9016 & n9668 ) ;
  assign n9670 = n5395 | n9669 ;
  assign n9675 = n9674 ^ n9670 ^ 1'b0 ;
  assign n9676 = n9667 & n9675 ;
  assign n9677 = n6471 ^ n6195 ^ n2120 ;
  assign n9682 = ( n7314 & ~n8084 ) | ( n7314 & n9335 ) | ( ~n8084 & n9335 ) ;
  assign n9678 = ( n606 & ~n1685 ) | ( n606 & n4281 ) | ( ~n1685 & n4281 ) ;
  assign n9679 = n7828 | n9678 ;
  assign n9680 = n9679 ^ n8017 ^ 1'b0 ;
  assign n9681 = n2622 & n9680 ;
  assign n9683 = n9682 ^ n9681 ^ n736 ;
  assign n9684 = n9683 ^ n4040 ^ 1'b0 ;
  assign n9685 = n2170 | n9684 ;
  assign n9686 = n9685 ^ n7281 ^ 1'b0 ;
  assign n9687 = n9677 & n9686 ;
  assign n9688 = ( n311 & ~n3030 ) | ( n311 & n9687 ) | ( ~n3030 & n9687 ) ;
  assign n9689 = n6646 & ~n7022 ;
  assign n9690 = n4610 ^ n4057 ^ n3750 ;
  assign n9691 = n9690 ^ n7288 ^ n3697 ;
  assign n9696 = n416 & n2332 ;
  assign n9697 = n9696 ^ n4233 ^ 1'b0 ;
  assign n9698 = n9697 ^ n6210 ^ n422 ;
  assign n9692 = n6326 ^ n407 ^ n378 ;
  assign n9693 = n2633 & ~n9692 ;
  assign n9694 = n9693 ^ n5891 ^ 1'b0 ;
  assign n9695 = n9694 ^ n9481 ^ n731 ;
  assign n9699 = n9698 ^ n9695 ^ 1'b0 ;
  assign n9700 = n9691 & n9699 ;
  assign n9701 = ~n9689 & n9700 ;
  assign n9702 = n2911 ^ n2905 ^ 1'b0 ;
  assign n9703 = ~n8403 & n9702 ;
  assign n9708 = ( ~n1915 & n4144 ) | ( ~n1915 & n4399 ) | ( n4144 & n4399 ) ;
  assign n9704 = ~n1486 & n5354 ;
  assign n9705 = n9704 ^ n5687 ^ 1'b0 ;
  assign n9706 = n3593 & n9705 ;
  assign n9707 = n9706 ^ n8354 ^ n1371 ;
  assign n9709 = n9708 ^ n9707 ^ n1228 ;
  assign n9710 = x15 | n5619 ;
  assign n9712 = n2222 ^ n2070 ^ n348 ;
  assign n9711 = n5598 ^ n3583 ^ n2296 ;
  assign n9713 = n9712 ^ n9711 ^ n7769 ;
  assign n9714 = n9710 & ~n9713 ;
  assign n9715 = ( n456 & n956 ) | ( n456 & n1587 ) | ( n956 & n1587 ) ;
  assign n9716 = ( x6 & n4552 ) | ( x6 & ~n8732 ) | ( n4552 & ~n8732 ) ;
  assign n9717 = ~n6026 & n6090 ;
  assign n9718 = n9717 ^ n1300 ^ 1'b0 ;
  assign n9719 = ~n4860 & n7010 ;
  assign n9720 = n5904 ^ n3278 ^ 1'b0 ;
  assign n9721 = n9720 ^ n1649 ^ 1'b0 ;
  assign n9722 = n9719 | n9721 ;
  assign n9723 = n9722 ^ n3023 ^ 1'b0 ;
  assign n9724 = n1015 & n9723 ;
  assign n9725 = ( n2739 & ~n7441 ) | ( n2739 & n9724 ) | ( ~n7441 & n9724 ) ;
  assign n9726 = n2160 & n7970 ;
  assign n9727 = n9726 ^ n2395 ^ 1'b0 ;
  assign n9728 = n2799 ^ n1671 ^ 1'b0 ;
  assign n9729 = n2286 ^ n1119 ^ 1'b0 ;
  assign n9730 = n4022 & n9729 ;
  assign n9731 = n9730 ^ n4666 ^ 1'b0 ;
  assign n9732 = ( ~n5939 & n9728 ) | ( ~n5939 & n9731 ) | ( n9728 & n9731 ) ;
  assign n9733 = n9732 ^ n9554 ^ n3678 ;
  assign n9735 = n422 ^ x72 ^ 1'b0 ;
  assign n9736 = n168 | n9735 ;
  assign n9737 = n9736 ^ x28 ^ 1'b0 ;
  assign n9734 = n5123 & ~n7853 ;
  assign n9738 = n9737 ^ n9734 ^ 1'b0 ;
  assign n9739 = ( n631 & ~n4736 ) | ( n631 & n6319 ) | ( ~n4736 & n6319 ) ;
  assign n9740 = x30 & n9739 ;
  assign n9741 = n9740 ^ n8896 ^ 1'b0 ;
  assign n9742 = ( ~n462 & n2175 ) | ( ~n462 & n6984 ) | ( n2175 & n6984 ) ;
  assign n9743 = n3471 ^ x54 ^ 1'b0 ;
  assign n9744 = ( ~n4622 & n9742 ) | ( ~n4622 & n9743 ) | ( n9742 & n9743 ) ;
  assign n9745 = n3548 ^ n1295 ^ 1'b0 ;
  assign n9753 = ( ~n1984 & n3759 ) | ( ~n1984 & n4634 ) | ( n3759 & n4634 ) ;
  assign n9746 = n5492 ^ n910 ^ 1'b0 ;
  assign n9747 = ~n1732 & n9746 ;
  assign n9748 = n8778 ^ n7107 ^ n2562 ;
  assign n9749 = n1200 | n9748 ;
  assign n9750 = n2934 | n9749 ;
  assign n9751 = ( n2448 & n9747 ) | ( n2448 & n9750 ) | ( n9747 & n9750 ) ;
  assign n9752 = ~n7690 & n9751 ;
  assign n9754 = n9753 ^ n9752 ^ 1'b0 ;
  assign n9756 = n1836 | n8311 ;
  assign n9755 = ( n1674 & ~n7377 ) | ( n1674 & n8674 ) | ( ~n7377 & n8674 ) ;
  assign n9757 = n9756 ^ n9755 ^ n2609 ;
  assign n9758 = n1316 & n1793 ;
  assign n9759 = n9758 ^ n5606 ^ 1'b0 ;
  assign n9760 = ( ~n1292 & n4649 ) | ( ~n1292 & n9759 ) | ( n4649 & n9759 ) ;
  assign n9761 = n3770 | n6288 ;
  assign n9762 = ~n8136 & n9761 ;
  assign n9763 = ~n5743 & n8382 ;
  assign n9764 = ~n7713 & n9763 ;
  assign n9768 = n3213 & ~n6048 ;
  assign n9769 = n9768 ^ n2071 ^ 1'b0 ;
  assign n9770 = ( n1568 & n6913 ) | ( n1568 & ~n9769 ) | ( n6913 & ~n9769 ) ;
  assign n9771 = n9770 ^ n2663 ^ n1675 ;
  assign n9766 = ~n3835 & n6159 ;
  assign n9767 = ~n7252 & n9766 ;
  assign n9765 = n3423 & ~n7421 ;
  assign n9772 = n9771 ^ n9767 ^ n9765 ;
  assign n9773 = n9772 ^ n2835 ^ n1276 ;
  assign n9774 = ( x121 & n2475 ) | ( x121 & n8383 ) | ( n2475 & n8383 ) ;
  assign n9775 = n8126 & ~n9774 ;
  assign n9776 = n3723 ^ n3061 ^ x42 ;
  assign n9777 = n7825 & n9776 ;
  assign n9778 = ( n472 & n2527 ) | ( n472 & ~n9777 ) | ( n2527 & ~n9777 ) ;
  assign n9782 = n1553 & ~n5546 ;
  assign n9779 = n5138 ^ n5058 ^ 1'b0 ;
  assign n9780 = n4096 | n9779 ;
  assign n9781 = n9780 ^ n7425 ^ 1'b0 ;
  assign n9783 = n9782 ^ n9781 ^ 1'b0 ;
  assign n9784 = n5749 & ~n9783 ;
  assign n9785 = n8844 & ~n9233 ;
  assign n9786 = ~n3091 & n9785 ;
  assign n9787 = n8146 ^ n6057 ^ 1'b0 ;
  assign n9788 = ( n3581 & ~n8920 ) | ( n3581 & n9787 ) | ( ~n8920 & n9787 ) ;
  assign n9789 = n4249 & ~n8835 ;
  assign n9790 = n9789 ^ n2418 ^ 1'b0 ;
  assign n9791 = n3577 & ~n9790 ;
  assign n9792 = n9791 ^ n2993 ^ 1'b0 ;
  assign n9793 = ( n231 & n1955 ) | ( n231 & n6399 ) | ( n1955 & n6399 ) ;
  assign n9794 = n9793 ^ n8010 ^ n6281 ;
  assign n9795 = ( n348 & n9792 ) | ( n348 & n9794 ) | ( n9792 & n9794 ) ;
  assign n9796 = ( n1157 & n6927 ) | ( n1157 & ~n9795 ) | ( n6927 & ~n9795 ) ;
  assign n9797 = ~n256 & n5133 ;
  assign n9798 = ~n5413 & n5489 ;
  assign n9799 = n5174 ^ n3117 ^ 1'b0 ;
  assign n9800 = ~n9798 & n9799 ;
  assign n9801 = ~n846 & n1279 ;
  assign n9802 = ~n7898 & n9801 ;
  assign n9803 = n9802 ^ n2088 ^ 1'b0 ;
  assign n9804 = n9803 ^ n9607 ^ 1'b0 ;
  assign n9805 = n9800 & n9804 ;
  assign n9806 = n9797 | n9805 ;
  assign n9807 = n9796 | n9806 ;
  assign n9808 = n4352 | n9807 ;
  assign n9809 = n4608 | n7217 ;
  assign n9811 = n4401 ^ n395 ^ 1'b0 ;
  assign n9812 = n7121 & ~n9811 ;
  assign n9813 = n2230 ^ n561 ^ 1'b0 ;
  assign n9814 = n9812 & n9813 ;
  assign n9815 = ( ~n808 & n4165 ) | ( ~n808 & n9814 ) | ( n4165 & n9814 ) ;
  assign n9810 = n6541 ^ n5885 ^ n4996 ;
  assign n9816 = n9815 ^ n9810 ^ 1'b0 ;
  assign n9817 = ~n1091 & n7790 ;
  assign n9818 = n2783 & n9817 ;
  assign n9819 = ( x30 & ~n5959 ) | ( x30 & n9818 ) | ( ~n5959 & n9818 ) ;
  assign n9820 = n1953 & ~n7113 ;
  assign n9821 = ~n2033 & n9820 ;
  assign n9822 = ( n1631 & n9819 ) | ( n1631 & n9821 ) | ( n9819 & n9821 ) ;
  assign n9823 = n9822 ^ n1342 ^ 1'b0 ;
  assign n9824 = n6579 ^ n3697 ^ 1'b0 ;
  assign n9825 = n9823 & n9824 ;
  assign n9826 = x110 & ~n4453 ;
  assign n9827 = n7059 ^ n4879 ^ 1'b0 ;
  assign n9828 = n4311 ^ n2648 ^ 1'b0 ;
  assign n9833 = ~n875 & n1629 ;
  assign n9834 = n9833 ^ n933 ^ 1'b0 ;
  assign n9835 = ( ~n861 & n2347 ) | ( ~n861 & n9834 ) | ( n2347 & n9834 ) ;
  assign n9836 = n9835 ^ n8455 ^ n6833 ;
  assign n9829 = n4076 ^ n1765 ^ 1'b0 ;
  assign n9830 = n9829 ^ n1828 ^ n1246 ;
  assign n9831 = n3934 & n4107 ;
  assign n9832 = ~n9830 & n9831 ;
  assign n9837 = n9836 ^ n9832 ^ 1'b0 ;
  assign n9838 = n9828 | n9837 ;
  assign n9839 = n3016 ^ n1688 ^ 1'b0 ;
  assign n9840 = n1616 & n5864 ;
  assign n9841 = n8204 | n9840 ;
  assign n9842 = n3683 & ~n9841 ;
  assign n9843 = n1862 | n9842 ;
  assign n9844 = n5807 ^ n1457 ^ 1'b0 ;
  assign n9845 = n7396 | n9844 ;
  assign n9846 = n9845 ^ n4045 ^ 1'b0 ;
  assign n9851 = n4753 ^ n3260 ^ n1043 ;
  assign n9849 = n660 & ~n6008 ;
  assign n9850 = n9849 ^ n1085 ^ 1'b0 ;
  assign n9847 = ( n4512 & ~n5542 ) | ( n4512 & n7641 ) | ( ~n5542 & n7641 ) ;
  assign n9848 = ( ~n2938 & n9771 ) | ( ~n2938 & n9847 ) | ( n9771 & n9847 ) ;
  assign n9852 = n9851 ^ n9850 ^ n9848 ;
  assign n9853 = n9846 & ~n9852 ;
  assign n9854 = ~n766 & n9043 ;
  assign n9855 = n2109 ^ n2030 ^ n1636 ;
  assign n9856 = n857 | n9774 ;
  assign n9857 = ~n9855 & n9856 ;
  assign n9858 = n3657 & n9857 ;
  assign n9859 = n203 & ~n4977 ;
  assign n9860 = n9859 ^ n2332 ^ 1'b0 ;
  assign n9861 = ( n2325 & n9858 ) | ( n2325 & n9860 ) | ( n9858 & n9860 ) ;
  assign n9862 = ~n1480 & n5282 ;
  assign n9863 = n4260 & n9862 ;
  assign n9864 = n8128 ^ n2521 ^ 1'b0 ;
  assign n9865 = ~n4562 & n9864 ;
  assign n9866 = n9865 ^ n3928 ^ n3847 ;
  assign n9867 = ( n9229 & ~n9682 ) | ( n9229 & n9866 ) | ( ~n9682 & n9866 ) ;
  assign n9868 = ~n3622 & n5383 ;
  assign n9869 = n9868 ^ n3495 ^ 1'b0 ;
  assign n9870 = n2823 & ~n3138 ;
  assign n9871 = n307 & n9870 ;
  assign n9874 = n5647 | n8136 ;
  assign n9875 = n2394 | n9874 ;
  assign n9876 = n9875 ^ n1590 ^ x43 ;
  assign n9872 = n6299 ^ n2773 ^ 1'b0 ;
  assign n9873 = ( n1006 & n3654 ) | ( n1006 & ~n9872 ) | ( n3654 & ~n9872 ) ;
  assign n9877 = n9876 ^ n9873 ^ 1'b0 ;
  assign n9878 = n2527 & ~n5373 ;
  assign n9880 = n2397 & ~n5712 ;
  assign n9881 = n9880 ^ n5918 ^ 1'b0 ;
  assign n9879 = ~n3785 & n8398 ;
  assign n9882 = n9881 ^ n9879 ^ 1'b0 ;
  assign n9883 = n9793 ^ n1488 ^ 1'b0 ;
  assign n9884 = n9883 ^ x15 ^ 1'b0 ;
  assign n9885 = n3444 & n9884 ;
  assign n9886 = n5421 | n7754 ;
  assign n9887 = ~n275 & n9886 ;
  assign n9888 = n3743 & n9887 ;
  assign n9890 = n6818 ^ n3690 ^ n1763 ;
  assign n9891 = n9890 ^ n5576 ^ 1'b0 ;
  assign n9892 = ~n6705 & n9891 ;
  assign n9889 = n6553 ^ n4803 ^ 1'b0 ;
  assign n9893 = n9892 ^ n9889 ^ 1'b0 ;
  assign n9896 = ~n2299 & n4528 ;
  assign n9897 = n9896 ^ n990 ^ 1'b0 ;
  assign n9898 = n9897 ^ n4933 ^ n2712 ;
  assign n9894 = n3779 ^ n2102 ^ 1'b0 ;
  assign n9895 = ~n6860 & n9894 ;
  assign n9899 = n9898 ^ n9895 ^ 1'b0 ;
  assign n9900 = n1928 & n2638 ;
  assign n9901 = n9900 ^ n5065 ^ 1'b0 ;
  assign n9902 = n9901 ^ n5031 ^ x81 ;
  assign n9903 = ( n4598 & n5539 ) | ( n4598 & n9533 ) | ( n5539 & n9533 ) ;
  assign n9904 = ~n1283 & n3991 ;
  assign n9905 = n9904 ^ n2700 ^ 1'b0 ;
  assign n9906 = n9905 ^ n872 ^ n744 ;
  assign n9907 = n8804 ^ n8646 ^ n6807 ;
  assign n9908 = n7613 ^ x7 ^ 1'b0 ;
  assign n9909 = ~n8482 & n9908 ;
  assign n9910 = ~n3303 & n9909 ;
  assign n9911 = ( n1603 & n2851 ) | ( n1603 & ~n6824 ) | ( n2851 & ~n6824 ) ;
  assign n9912 = ( n1628 & n9910 ) | ( n1628 & ~n9911 ) | ( n9910 & ~n9911 ) ;
  assign n9913 = n2487 ^ n2170 ^ n1500 ;
  assign n9914 = n6662 ^ n726 ^ 1'b0 ;
  assign n9915 = n7247 ^ n7117 ^ 1'b0 ;
  assign n9916 = n1969 | n7419 ;
  assign n9917 = n9915 & ~n9916 ;
  assign n9918 = ~n6427 & n9917 ;
  assign n9919 = n4727 ^ n3977 ^ n2866 ;
  assign n9920 = n9919 ^ n4230 ^ n610 ;
  assign n9921 = n2279 & ~n3295 ;
  assign n9922 = ~n9920 & n9921 ;
  assign n9923 = n9774 ^ n2637 ^ n461 ;
  assign n9924 = n9923 ^ n226 ^ 1'b0 ;
  assign n9925 = x34 & ~n9924 ;
  assign n9926 = n1575 | n9925 ;
  assign n9927 = ( n8688 & ~n9922 ) | ( n8688 & n9926 ) | ( ~n9922 & n9926 ) ;
  assign n9928 = n6145 ^ n4911 ^ 1'b0 ;
  assign n9929 = n7221 & ~n9928 ;
  assign n9930 = n8265 ^ n6376 ^ 1'b0 ;
  assign n9931 = n2197 | n2256 ;
  assign n9932 = n9931 ^ n253 ^ 1'b0 ;
  assign n9933 = n5296 ^ n965 ^ 1'b0 ;
  assign n9934 = n5441 & n9933 ;
  assign n9935 = n6746 ^ n5083 ^ n1283 ;
  assign n9936 = n2964 | n9935 ;
  assign n9937 = n9936 ^ n6363 ^ n3825 ;
  assign n9938 = ( n2200 & n5146 ) | ( n2200 & n9937 ) | ( n5146 & n9937 ) ;
  assign n9939 = n9934 & ~n9938 ;
  assign n9940 = n9932 & n9939 ;
  assign n9941 = n8870 ^ n5313 ^ n4591 ;
  assign n9942 = n4048 & ~n7180 ;
  assign n9943 = ~n9941 & n9942 ;
  assign n9949 = n1062 | n1745 ;
  assign n9950 = n9949 ^ n5327 ^ 1'b0 ;
  assign n9947 = ~n767 & n4445 ;
  assign n9948 = n6588 & n9947 ;
  assign n9944 = n8843 ^ n8010 ^ n4403 ;
  assign n9945 = ~n1163 & n9944 ;
  assign n9946 = n9945 ^ n5054 ^ 1'b0 ;
  assign n9951 = n9950 ^ n9948 ^ n9946 ;
  assign n9952 = n7542 ^ n2905 ^ 1'b0 ;
  assign n9953 = ( n557 & n4832 ) | ( n557 & ~n6113 ) | ( n4832 & ~n6113 ) ;
  assign n9954 = n9952 & ~n9953 ;
  assign n9955 = n6438 & n9954 ;
  assign n9956 = ( n332 & n3200 ) | ( n332 & n4281 ) | ( n3200 & n4281 ) ;
  assign n9957 = n2802 ^ n2544 ^ n1368 ;
  assign n9958 = n9957 ^ n7769 ^ n785 ;
  assign n9959 = n9958 ^ n1008 ^ 1'b0 ;
  assign n9960 = x54 & ~n9959 ;
  assign n9961 = n7102 ^ n5538 ^ 1'b0 ;
  assign n9962 = ~n1450 & n2094 ;
  assign n9963 = ~n176 & n9962 ;
  assign n9964 = n2237 | n9963 ;
  assign n9965 = n9964 ^ n3103 ^ 1'b0 ;
  assign n9966 = ( ~n7759 & n7990 ) | ( ~n7759 & n9000 ) | ( n7990 & n9000 ) ;
  assign n9967 = n9965 & n9966 ;
  assign n9968 = ( n1757 & ~n6030 ) | ( n1757 & n7265 ) | ( ~n6030 & n7265 ) ;
  assign n9969 = ~n9967 & n9968 ;
  assign n9970 = n9969 ^ n2210 ^ 1'b0 ;
  assign n9971 = n9970 ^ n9294 ^ 1'b0 ;
  assign n9972 = n9971 ^ n4888 ^ 1'b0 ;
  assign n9973 = n9961 & ~n9972 ;
  assign n9974 = n6267 ^ n3028 ^ n890 ;
  assign n9975 = n9974 ^ n6324 ^ 1'b0 ;
  assign n9976 = x94 & ~n3482 ;
  assign n9979 = n549 & n6693 ;
  assign n9980 = n8348 & n9979 ;
  assign n9977 = ~n2105 & n8811 ;
  assign n9978 = n9977 ^ n4239 ^ 1'b0 ;
  assign n9981 = n9980 ^ n9978 ^ 1'b0 ;
  assign n9982 = n5894 & n9981 ;
  assign n9983 = n9982 ^ n8636 ^ n6274 ;
  assign n9984 = n8599 ^ n393 ^ x25 ;
  assign n9985 = n7539 | n7848 ;
  assign n9986 = x12 | n9985 ;
  assign n9987 = n9986 ^ n1802 ^ n242 ;
  assign n9988 = ( n6406 & n7391 ) | ( n6406 & ~n9339 ) | ( n7391 & ~n9339 ) ;
  assign n9989 = ( n1085 & n7146 ) | ( n1085 & ~n9988 ) | ( n7146 & ~n9988 ) ;
  assign n9993 = ( n3156 & n3221 ) | ( n3156 & ~n4726 ) | ( n3221 & ~n4726 ) ;
  assign n9990 = ~n4187 & n5096 ;
  assign n9991 = n9990 ^ n5790 ^ 1'b0 ;
  assign n9992 = n9991 ^ n7911 ^ n4695 ;
  assign n9994 = n9993 ^ n9992 ^ n714 ;
  assign n9998 = ( x3 & n242 ) | ( x3 & n4758 ) | ( n242 & n4758 ) ;
  assign n9999 = n9998 ^ n3702 ^ n1427 ;
  assign n9995 = n3904 & ~n4017 ;
  assign n9996 = n9995 ^ n1164 ^ 1'b0 ;
  assign n9997 = ( n7769 & n8368 ) | ( n7769 & ~n9996 ) | ( n8368 & ~n9996 ) ;
  assign n10000 = n9999 ^ n9997 ^ n5692 ;
  assign n10003 = n1373 | n1727 ;
  assign n10001 = ~n5625 & n7456 ;
  assign n10002 = n10001 ^ n1987 ^ 1'b0 ;
  assign n10004 = n10003 ^ n10002 ^ n3891 ;
  assign n10005 = n5562 | n9440 ;
  assign n10006 = n10005 ^ n2040 ^ n1504 ;
  assign n10007 = n4161 ^ n2835 ^ n1288 ;
  assign n10008 = n2753 & n10007 ;
  assign n10009 = ~n592 & n2392 ;
  assign n10010 = n10009 ^ n4748 ^ n1685 ;
  assign n10011 = ( n2094 & ~n9298 ) | ( n2094 & n10010 ) | ( ~n9298 & n10010 ) ;
  assign n10013 = n536 | n1436 ;
  assign n10014 = n10013 ^ n1473 ^ 1'b0 ;
  assign n10015 = n10014 ^ n493 ^ 1'b0 ;
  assign n10012 = n2138 & ~n6091 ;
  assign n10016 = n10015 ^ n10012 ^ 1'b0 ;
  assign n10017 = n4304 ^ n4245 ^ 1'b0 ;
  assign n10018 = n2406 & ~n10017 ;
  assign n10019 = n10018 ^ n7166 ^ n893 ;
  assign n10020 = ( n1838 & n2812 ) | ( n1838 & n8959 ) | ( n2812 & n8959 ) ;
  assign n10021 = ( n3164 & n3679 ) | ( n3164 & ~n10020 ) | ( n3679 & ~n10020 ) ;
  assign n10022 = ( ~n6123 & n6164 ) | ( ~n6123 & n10021 ) | ( n6164 & n10021 ) ;
  assign n10023 = n8681 ^ n6616 ^ 1'b0 ;
  assign n10024 = ~n10022 & n10023 ;
  assign n10025 = ~n9656 & n10024 ;
  assign n10026 = n10019 & n10025 ;
  assign n10027 = n9157 ^ n1513 ^ 1'b0 ;
  assign n10028 = n1727 | n10027 ;
  assign n10029 = ( ~x61 & n5300 ) | ( ~x61 & n10028 ) | ( n5300 & n10028 ) ;
  assign n10030 = n281 | n308 ;
  assign n10031 = n10030 ^ n1984 ^ 1'b0 ;
  assign n10032 = n10031 ^ n1466 ^ 1'b0 ;
  assign n10033 = n3886 & n10032 ;
  assign n10034 = n4967 ^ n2292 ^ 1'b0 ;
  assign n10035 = n706 & n10034 ;
  assign n10036 = n10035 ^ n611 ^ 1'b0 ;
  assign n10037 = ( ~n7035 & n8211 ) | ( ~n7035 & n8636 ) | ( n8211 & n8636 ) ;
  assign n10043 = n2924 | n8504 ;
  assign n10044 = n4545 | n10043 ;
  assign n10039 = n966 | n4705 ;
  assign n10040 = n10039 ^ n3716 ^ 1'b0 ;
  assign n10038 = n1933 & n5564 ;
  assign n10041 = n10040 ^ n10038 ^ 1'b0 ;
  assign n10042 = n3174 & n10041 ;
  assign n10045 = n10044 ^ n10042 ^ 1'b0 ;
  assign n10046 = ( ~n326 & n3491 ) | ( ~n326 & n3519 ) | ( n3491 & n3519 ) ;
  assign n10047 = n1551 & n7895 ;
  assign n10048 = ~n4658 & n10047 ;
  assign n10049 = ( n1456 & n5259 ) | ( n1456 & n10048 ) | ( n5259 & n10048 ) ;
  assign n10050 = n10046 & ~n10049 ;
  assign n10051 = n10050 ^ n7291 ^ 1'b0 ;
  assign n10052 = n7925 ^ n1098 ^ n136 ;
  assign n10053 = n10052 ^ n579 ^ n240 ;
  assign n10056 = ~n8854 & n9173 ;
  assign n10057 = n350 & n10056 ;
  assign n10058 = n4691 ^ n1762 ^ 1'b0 ;
  assign n10059 = ~n3710 & n10058 ;
  assign n10060 = ( n3343 & n10057 ) | ( n3343 & ~n10059 ) | ( n10057 & ~n10059 ) ;
  assign n10054 = n8724 ^ n2443 ^ 1'b0 ;
  assign n10055 = n7028 & ~n10054 ;
  assign n10061 = n10060 ^ n10055 ^ 1'b0 ;
  assign n10062 = n7283 & ~n7550 ;
  assign n10063 = n10062 ^ n5761 ^ n1268 ;
  assign n10064 = ( ~n257 & n771 ) | ( ~n257 & n2120 ) | ( n771 & n2120 ) ;
  assign n10065 = ( n308 & n606 ) | ( n308 & n10064 ) | ( n606 & n10064 ) ;
  assign n10066 = ( n885 & n4298 ) | ( n885 & n10065 ) | ( n4298 & n10065 ) ;
  assign n10067 = n10066 ^ n5542 ^ n1563 ;
  assign n10068 = x112 | n4514 ;
  assign n10069 = n6847 ^ n988 ^ 1'b0 ;
  assign n10070 = n2269 & n10069 ;
  assign n10071 = n10070 ^ n1320 ^ 1'b0 ;
  assign n10072 = n4377 & n10071 ;
  assign n10073 = ~n3012 & n10072 ;
  assign n10074 = ~n3113 & n10073 ;
  assign n10075 = n10068 | n10074 ;
  assign n10076 = n7574 ^ n4057 ^ n2388 ;
  assign n10077 = n10076 ^ n5199 ^ 1'b0 ;
  assign n10078 = ( n7772 & n8792 ) | ( n7772 & n10077 ) | ( n8792 & n10077 ) ;
  assign n10081 = n2569 | n5540 ;
  assign n10079 = ( ~n1097 & n2086 ) | ( ~n1097 & n3432 ) | ( n2086 & n3432 ) ;
  assign n10080 = n10079 ^ n6728 ^ n3641 ;
  assign n10082 = n10081 ^ n10080 ^ n1454 ;
  assign n10083 = n4162 & ~n7426 ;
  assign n10090 = n3741 ^ n3636 ^ n1290 ;
  assign n10091 = n624 & n1679 ;
  assign n10092 = n10090 & n10091 ;
  assign n10089 = ( n376 & n7469 ) | ( n376 & n8816 ) | ( n7469 & n8816 ) ;
  assign n10093 = n10092 ^ n10089 ^ n3551 ;
  assign n10084 = ( n3212 & n4453 ) | ( n3212 & ~n8202 ) | ( n4453 & ~n8202 ) ;
  assign n10085 = n10084 ^ n9322 ^ n2060 ;
  assign n10086 = n4305 | n10085 ;
  assign n10087 = n7897 & ~n10086 ;
  assign n10088 = n10087 ^ n7611 ^ n1846 ;
  assign n10094 = n10093 ^ n10088 ^ n7696 ;
  assign n10095 = n7192 ^ n5831 ^ n170 ;
  assign n10096 = n3935 ^ n3887 ^ n495 ;
  assign n10097 = ~n4399 & n10096 ;
  assign n10098 = n10095 & n10097 ;
  assign n10099 = ( n1327 & ~n3452 ) | ( n1327 & n3993 ) | ( ~n3452 & n3993 ) ;
  assign n10101 = n5475 ^ n1814 ^ n1014 ;
  assign n10100 = n8740 ^ n6359 ^ n2646 ;
  assign n10102 = n10101 ^ n10100 ^ 1'b0 ;
  assign n10103 = n5851 ^ n414 ^ x22 ;
  assign n10104 = ( n2336 & n6316 ) | ( n2336 & n6593 ) | ( n6316 & n6593 ) ;
  assign n10105 = n4821 ^ n242 ^ 1'b0 ;
  assign n10109 = ~n376 & n3820 ;
  assign n10110 = n5157 & n10109 ;
  assign n10106 = n8559 ^ n662 ^ 1'b0 ;
  assign n10107 = ~n3198 & n10106 ;
  assign n10108 = n10107 ^ n9704 ^ n2002 ;
  assign n10111 = n10110 ^ n10108 ^ 1'b0 ;
  assign n10112 = ( n10104 & n10105 ) | ( n10104 & ~n10111 ) | ( n10105 & ~n10111 ) ;
  assign n10113 = n4695 ^ n677 ^ 1'b0 ;
  assign n10114 = ( n242 & n2171 ) | ( n242 & n5774 ) | ( n2171 & n5774 ) ;
  assign n10115 = n8084 | n10114 ;
  assign n10116 = n3202 & ~n8195 ;
  assign n10117 = n10116 ^ n1633 ^ 1'b0 ;
  assign n10118 = ( n10113 & n10115 ) | ( n10113 & n10117 ) | ( n10115 & n10117 ) ;
  assign n10119 = ( n1675 & n4500 ) | ( n1675 & ~n7535 ) | ( n4500 & ~n7535 ) ;
  assign n10120 = ( n1105 & n9815 ) | ( n1105 & ~n10119 ) | ( n9815 & ~n10119 ) ;
  assign n10123 = n510 | n1353 ;
  assign n10124 = n2779 & ~n10123 ;
  assign n10125 = ( n1263 & ~n1880 ) | ( n1263 & n10124 ) | ( ~n1880 & n10124 ) ;
  assign n10126 = n10125 ^ n5746 ^ n3813 ;
  assign n10121 = n1122 | n6029 ;
  assign n10122 = n10121 ^ n7684 ^ 1'b0 ;
  assign n10127 = n10126 ^ n10122 ^ n1024 ;
  assign n10128 = n4936 ^ n3718 ^ n939 ;
  assign n10129 = n10128 ^ n8662 ^ n5915 ;
  assign n10130 = n4468 & ~n7152 ;
  assign n10131 = ~n10129 & n10130 ;
  assign n10138 = ~n192 & n1437 ;
  assign n10132 = ( ~n1644 & n1955 ) | ( ~n1644 & n6423 ) | ( n1955 & n6423 ) ;
  assign n10134 = n3780 ^ n916 ^ n732 ;
  assign n10133 = n1282 & n1570 ;
  assign n10135 = n10134 ^ n10133 ^ 1'b0 ;
  assign n10136 = ( ~n8970 & n10132 ) | ( ~n8970 & n10135 ) | ( n10132 & n10135 ) ;
  assign n10137 = n9759 | n10136 ;
  assign n10139 = n10138 ^ n10137 ^ 1'b0 ;
  assign n10140 = n10139 ^ n4344 ^ 1'b0 ;
  assign n10141 = n1739 | n5112 ;
  assign n10142 = n10141 ^ n7008 ^ n3092 ;
  assign n10143 = ( ~n7273 & n7420 ) | ( ~n7273 & n10142 ) | ( n7420 & n10142 ) ;
  assign n10144 = n4983 ^ n4629 ^ 1'b0 ;
  assign n10145 = n352 & ~n10144 ;
  assign n10146 = n8779 & n10145 ;
  assign n10147 = n10146 ^ n8355 ^ 1'b0 ;
  assign n10148 = x67 & n5249 ;
  assign n10149 = n10148 ^ n6160 ^ 1'b0 ;
  assign n10150 = n7694 ^ n672 ^ 1'b0 ;
  assign n10151 = n3205 ^ n3138 ^ n861 ;
  assign n10152 = n6919 ^ n6170 ^ n760 ;
  assign n10154 = n3015 ^ n2489 ^ 1'b0 ;
  assign n10155 = n6448 & ~n10154 ;
  assign n10153 = n2186 & ~n3096 ;
  assign n10156 = n10155 ^ n10153 ^ 1'b0 ;
  assign n10157 = ( n5151 & n8240 ) | ( n5151 & ~n10156 ) | ( n8240 & ~n10156 ) ;
  assign n10158 = n2728 | n5776 ;
  assign n10159 = n10158 ^ n3882 ^ 1'b0 ;
  assign n10161 = n2744 ^ n1580 ^ n1268 ;
  assign n10162 = n10161 ^ n5279 ^ n894 ;
  assign n10163 = n10162 ^ n2411 ^ 1'b0 ;
  assign n10160 = n4887 ^ n4298 ^ 1'b0 ;
  assign n10164 = n10163 ^ n10160 ^ n8776 ;
  assign n10165 = ( n215 & n249 ) | ( n215 & ~n1647 ) | ( n249 & ~n1647 ) ;
  assign n10166 = ( n5177 & ~n6672 ) | ( n5177 & n10165 ) | ( ~n6672 & n10165 ) ;
  assign n10167 = ( n3216 & n4250 ) | ( n3216 & n4581 ) | ( n4250 & n4581 ) ;
  assign n10168 = ( n2347 & ~n10166 ) | ( n2347 & n10167 ) | ( ~n10166 & n10167 ) ;
  assign n10169 = n8244 ^ n1744 ^ 1'b0 ;
  assign n10170 = n2684 | n10169 ;
  assign n10171 = n7134 & ~n10170 ;
  assign n10172 = n10171 ^ n8022 ^ 1'b0 ;
  assign n10173 = n9206 ^ n1452 ^ 1'b0 ;
  assign n10174 = ~n4002 & n10173 ;
  assign n10175 = ( ~n3540 & n6327 ) | ( ~n3540 & n6406 ) | ( n6327 & n6406 ) ;
  assign n10176 = ( n3800 & ~n9323 ) | ( n3800 & n10175 ) | ( ~n9323 & n10175 ) ;
  assign n10177 = n2081 & n10176 ;
  assign n10178 = ~n10174 & n10177 ;
  assign n10179 = n5434 ^ n4570 ^ 1'b0 ;
  assign n10180 = n1168 & ~n8423 ;
  assign n10181 = n8389 ^ n563 ^ 1'b0 ;
  assign n10182 = n7265 ^ n3581 ^ 1'b0 ;
  assign n10183 = ( x79 & ~n325 ) | ( x79 & n3220 ) | ( ~n325 & n3220 ) ;
  assign n10184 = ( n732 & n4780 ) | ( n732 & n10183 ) | ( n4780 & n10183 ) ;
  assign n10187 = n1832 & ~n4572 ;
  assign n10185 = n8084 ^ n4122 ^ n503 ;
  assign n10186 = n6070 | n10185 ;
  assign n10188 = n10187 ^ n10186 ^ 1'b0 ;
  assign n10189 = ( n10182 & n10184 ) | ( n10182 & n10188 ) | ( n10184 & n10188 ) ;
  assign n10190 = n7235 ^ n4509 ^ 1'b0 ;
  assign n10191 = n3174 & ~n10190 ;
  assign n10192 = ~n1301 & n10191 ;
  assign n10193 = n10192 ^ n3499 ^ 1'b0 ;
  assign n10194 = ( ~n2242 & n9540 ) | ( ~n2242 & n10134 ) | ( n9540 & n10134 ) ;
  assign n10195 = ( n4216 & n10193 ) | ( n4216 & ~n10194 ) | ( n10193 & ~n10194 ) ;
  assign n10196 = n10108 ^ n3054 ^ 1'b0 ;
  assign n10197 = n3895 ^ n1700 ^ 1'b0 ;
  assign n10198 = ~n7320 & n10197 ;
  assign n10199 = ~n2153 & n10198 ;
  assign n10200 = ~n10196 & n10199 ;
  assign n10202 = ~n1899 & n6359 ;
  assign n10203 = n5847 & n10202 ;
  assign n10201 = n9255 ^ n8443 ^ n8250 ;
  assign n10204 = n10203 ^ n10201 ^ 1'b0 ;
  assign n10205 = n7747 & n10204 ;
  assign n10206 = n3649 | n9037 ;
  assign n10207 = n10206 ^ n2944 ^ 1'b0 ;
  assign n10208 = ~n6299 & n10207 ;
  assign n10209 = n3042 ^ n1455 ^ 1'b0 ;
  assign n10210 = n4761 & n10209 ;
  assign n10211 = ~n3851 & n7318 ;
  assign n10212 = n5520 & n10211 ;
  assign n10213 = n10212 ^ n980 ^ 1'b0 ;
  assign n10214 = ( ~n6385 & n10210 ) | ( ~n6385 & n10213 ) | ( n10210 & n10213 ) ;
  assign n10215 = x28 & n3990 ;
  assign n10216 = n3504 & n10215 ;
  assign n10217 = ( n664 & n5108 ) | ( n664 & ~n10216 ) | ( n5108 & ~n10216 ) ;
  assign n10218 = n2187 & n10217 ;
  assign n10219 = x116 & ~n2731 ;
  assign n10220 = n10219 ^ n6710 ^ n5941 ;
  assign n10222 = n756 & n2602 ;
  assign n10223 = ~n5814 & n10222 ;
  assign n10224 = ( n2230 & n2472 ) | ( n2230 & n10223 ) | ( n2472 & n10223 ) ;
  assign n10225 = n10224 ^ n2282 ^ 1'b0 ;
  assign n10221 = x119 | n5791 ;
  assign n10226 = n10225 ^ n10221 ^ n4479 ;
  assign n10227 = n1628 ^ n527 ^ 1'b0 ;
  assign n10228 = n10227 ^ n8916 ^ n2383 ;
  assign n10229 = n10228 ^ n9710 ^ 1'b0 ;
  assign n10230 = n4197 | n10229 ;
  assign n10231 = n969 | n5994 ;
  assign n10232 = n1752 | n10231 ;
  assign n10233 = n10232 ^ n7418 ^ n7280 ;
  assign n10234 = n985 & n6712 ;
  assign n10235 = ( n10230 & ~n10233 ) | ( n10230 & n10234 ) | ( ~n10233 & n10234 ) ;
  assign n10236 = n5070 ^ n4172 ^ 1'b0 ;
  assign n10237 = ~n170 & n10236 ;
  assign n10238 = n10237 ^ n7265 ^ 1'b0 ;
  assign n10239 = ( n136 & ~n4546 ) | ( n136 & n9756 ) | ( ~n4546 & n9756 ) ;
  assign n10240 = ~n4049 & n7667 ;
  assign n10241 = ~x41 & n10240 ;
  assign n10242 = n10241 ^ n2629 ^ n1977 ;
  assign n10243 = ( n4215 & n9315 ) | ( n4215 & n9462 ) | ( n9315 & n9462 ) ;
  assign n10244 = n6501 | n9925 ;
  assign n10245 = n3475 | n3626 ;
  assign n10246 = n3068 | n10245 ;
  assign n10247 = ( ~n1522 & n9900 ) | ( ~n1522 & n10246 ) | ( n9900 & n10246 ) ;
  assign n10248 = ( ~n3530 & n6198 ) | ( ~n3530 & n10247 ) | ( n6198 & n10247 ) ;
  assign n10249 = ( n7379 & ~n9286 ) | ( n7379 & n10248 ) | ( ~n9286 & n10248 ) ;
  assign n10250 = ( n2461 & n4305 ) | ( n2461 & n10249 ) | ( n4305 & n10249 ) ;
  assign n10251 = n3135 & ~n5578 ;
  assign n10252 = n171 & n10251 ;
  assign n10253 = n1664 & ~n2217 ;
  assign n10254 = n10253 ^ n6068 ^ 1'b0 ;
  assign n10255 = n10252 | n10254 ;
  assign n10256 = x118 & n4242 ;
  assign n10257 = n9079 & ~n10256 ;
  assign n10258 = n2665 & n5788 ;
  assign n10259 = ~n6639 & n10258 ;
  assign n10260 = ( n880 & ~n10257 ) | ( n880 & n10259 ) | ( ~n10257 & n10259 ) ;
  assign n10261 = ~n9530 & n10260 ;
  assign n10262 = n6627 & ~n6984 ;
  assign n10263 = n10262 ^ n1503 ^ 1'b0 ;
  assign n10264 = n10263 ^ n8595 ^ 1'b0 ;
  assign n10265 = n2839 ^ x61 ^ 1'b0 ;
  assign n10266 = n10265 ^ n3344 ^ 1'b0 ;
  assign n10267 = ( ~n4101 & n9313 ) | ( ~n4101 & n10266 ) | ( n9313 & n10266 ) ;
  assign n10268 = n4971 ^ n4515 ^ n353 ;
  assign n10269 = n10268 ^ x36 ^ 1'b0 ;
  assign n10270 = n8307 | n10269 ;
  assign n10271 = n10270 ^ n4061 ^ 1'b0 ;
  assign n10272 = ~n2116 & n10271 ;
  assign n10274 = x84 & ~n4861 ;
  assign n10275 = n6766 & ~n10274 ;
  assign n10273 = ( ~n1548 & n5579 ) | ( ~n1548 & n8475 ) | ( n5579 & n8475 ) ;
  assign n10276 = n10275 ^ n10273 ^ n7435 ;
  assign n10280 = n5712 ^ n3157 ^ n1533 ;
  assign n10281 = n759 & ~n10280 ;
  assign n10282 = n7917 & n10281 ;
  assign n10277 = ( n2312 & n3891 ) | ( n2312 & n9627 ) | ( n3891 & n9627 ) ;
  assign n10278 = ( n2364 & n4034 ) | ( n2364 & ~n10277 ) | ( n4034 & ~n10277 ) ;
  assign n10279 = ~n4657 & n10278 ;
  assign n10283 = n10282 ^ n10279 ^ n2884 ;
  assign n10284 = ( n2584 & n4017 ) | ( n2584 & ~n10283 ) | ( n4017 & ~n10283 ) ;
  assign n10285 = n7755 ^ n374 ^ 1'b0 ;
  assign n10286 = ~n5816 & n10285 ;
  assign n10287 = ( n971 & ~n4583 ) | ( n971 & n10286 ) | ( ~n4583 & n10286 ) ;
  assign n10288 = ( ~n559 & n1790 ) | ( ~n559 & n2803 ) | ( n1790 & n2803 ) ;
  assign n10289 = n7058 | n10288 ;
  assign n10296 = ( n1605 & n1920 ) | ( n1605 & n5550 ) | ( n1920 & n5550 ) ;
  assign n10290 = n233 | n1943 ;
  assign n10291 = n10290 ^ n440 ^ 1'b0 ;
  assign n10292 = n813 | n7409 ;
  assign n10293 = n8584 | n10292 ;
  assign n10294 = ~n3312 & n10293 ;
  assign n10295 = n10291 & n10294 ;
  assign n10297 = n10296 ^ n10295 ^ 1'b0 ;
  assign n10299 = ( n157 & n1024 ) | ( n157 & n4835 ) | ( n1024 & n4835 ) ;
  assign n10298 = n3776 & ~n7901 ;
  assign n10300 = n10299 ^ n10298 ^ 1'b0 ;
  assign n10301 = n1431 ^ n1182 ^ 1'b0 ;
  assign n10302 = ( n1900 & ~n4188 ) | ( n1900 & n10301 ) | ( ~n4188 & n10301 ) ;
  assign n10303 = ( n874 & n4500 ) | ( n874 & n10302 ) | ( n4500 & n10302 ) ;
  assign n10304 = n5525 & n5724 ;
  assign n10305 = ~n724 & n10304 ;
  assign n10306 = n10305 ^ n6985 ^ 1'b0 ;
  assign n10307 = n10306 ^ n9197 ^ n1952 ;
  assign n10313 = n9399 ^ n5513 ^ n4273 ;
  assign n10308 = ( n1436 & n1584 ) | ( n1436 & ~n2763 ) | ( n1584 & ~n2763 ) ;
  assign n10309 = n6618 ^ n3667 ^ n2943 ;
  assign n10310 = ~n7926 & n10309 ;
  assign n10311 = n10308 & n10310 ;
  assign n10312 = n7587 | n10311 ;
  assign n10314 = n10313 ^ n10312 ^ 1'b0 ;
  assign n10315 = n2249 & ~n3399 ;
  assign n10316 = n751 & ~n8288 ;
  assign n10317 = ( ~n4097 & n7987 ) | ( ~n4097 & n10316 ) | ( n7987 & n10316 ) ;
  assign n10318 = n10317 ^ n763 ^ 1'b0 ;
  assign n10319 = n2941 & ~n9491 ;
  assign n10320 = ~n3209 & n6182 ;
  assign n10330 = n5059 ^ n3985 ^ n2923 ;
  assign n10327 = ( n1164 & ~n1301 ) | ( n1164 & n1326 ) | ( ~n1301 & n1326 ) ;
  assign n10328 = ( ~n5641 & n6381 ) | ( ~n5641 & n10327 ) | ( n6381 & n10327 ) ;
  assign n10321 = n2694 ^ n1408 ^ 1'b0 ;
  assign n10322 = n2873 & n5965 ;
  assign n10323 = n1439 & n10322 ;
  assign n10324 = n1767 & ~n8761 ;
  assign n10325 = n10323 & ~n10324 ;
  assign n10326 = n10321 & ~n10325 ;
  assign n10329 = n10328 ^ n10326 ^ 1'b0 ;
  assign n10331 = n10330 ^ n10329 ^ n3243 ;
  assign n10332 = n4293 & n4829 ;
  assign n10333 = n10332 ^ n5470 ^ 1'b0 ;
  assign n10341 = x30 & n7272 ;
  assign n10342 = n1694 & n10341 ;
  assign n10334 = ( ~n4954 & n5565 ) | ( ~n4954 & n6847 ) | ( n5565 & n6847 ) ;
  assign n10335 = ( n800 & n3323 ) | ( n800 & ~n4636 ) | ( n3323 & ~n4636 ) ;
  assign n10336 = ( n509 & n7388 ) | ( n509 & ~n10335 ) | ( n7388 & ~n10335 ) ;
  assign n10337 = n7891 & n10336 ;
  assign n10338 = n2218 & n10337 ;
  assign n10339 = n10334 | n10338 ;
  assign n10340 = n913 & n10339 ;
  assign n10343 = n10342 ^ n10340 ^ 1'b0 ;
  assign n10344 = ( n1114 & n2655 ) | ( n1114 & ~n4304 ) | ( n2655 & ~n4304 ) ;
  assign n10345 = n10344 ^ n4347 ^ n973 ;
  assign n10346 = n450 | n1518 ;
  assign n10347 = n6300 | n10346 ;
  assign n10348 = n10347 ^ n3992 ^ 1'b0 ;
  assign n10349 = ( ~n279 & n897 ) | ( ~n279 & n10348 ) | ( n897 & n10348 ) ;
  assign n10350 = ( n3764 & n3768 ) | ( n3764 & ~n3958 ) | ( n3768 & ~n3958 ) ;
  assign n10351 = n395 & ~n8423 ;
  assign n10352 = ~n10350 & n10351 ;
  assign n10353 = n10352 ^ n3334 ^ n3247 ;
  assign n10354 = ( n1838 & n2624 ) | ( n1838 & ~n8184 ) | ( n2624 & ~n8184 ) ;
  assign n10355 = n9255 ^ n2857 ^ n1714 ;
  assign n10356 = ( ~n6675 & n6963 ) | ( ~n6675 & n10355 ) | ( n6963 & n10355 ) ;
  assign n10357 = n9701 ^ n6004 ^ 1'b0 ;
  assign n10358 = n9827 & n10357 ;
  assign n10359 = n2692 ^ n1183 ^ 1'b0 ;
  assign n10360 = n10359 ^ x83 ^ 1'b0 ;
  assign n10361 = ~n4793 & n10360 ;
  assign n10362 = n1186 & n9941 ;
  assign n10363 = ~n10361 & n10362 ;
  assign n10364 = ~n170 & n3264 ;
  assign n10365 = n5837 ^ n4948 ^ 1'b0 ;
  assign n10366 = n2332 & n10365 ;
  assign n10367 = n10366 ^ n1706 ^ 1'b0 ;
  assign n10368 = n10364 & ~n10367 ;
  assign n10369 = ( n6413 & n7195 ) | ( n6413 & n10368 ) | ( n7195 & n10368 ) ;
  assign n10370 = n9732 ^ n8270 ^ n7971 ;
  assign n10371 = n7046 & n10370 ;
  assign n10372 = n2030 & ~n4611 ;
  assign n10377 = ( ~n3514 & n5029 ) | ( ~n3514 & n9043 ) | ( n5029 & n9043 ) ;
  assign n10374 = n2968 ^ x70 ^ 1'b0 ;
  assign n10375 = n10374 ^ n6427 ^ n5833 ;
  assign n10373 = n1199 & ~n4454 ;
  assign n10376 = n10375 ^ n10373 ^ 1'b0 ;
  assign n10378 = n10377 ^ n10376 ^ n8490 ;
  assign n10379 = n6564 | n10082 ;
  assign n10380 = n10379 ^ n3688 ^ 1'b0 ;
  assign n10381 = n1199 & n3792 ;
  assign n10382 = n3263 ^ n909 ^ 1'b0 ;
  assign n10383 = n4761 & n10382 ;
  assign n10384 = n8934 ^ n6320 ^ 1'b0 ;
  assign n10385 = ( n7963 & ~n10383 ) | ( n7963 & n10384 ) | ( ~n10383 & n10384 ) ;
  assign n10386 = n440 & ~n1313 ;
  assign n10387 = ~n3125 & n10386 ;
  assign n10388 = n10387 ^ n10080 ^ n5108 ;
  assign n10389 = ( n1384 & n5875 ) | ( n1384 & n10029 ) | ( n5875 & n10029 ) ;
  assign n10390 = n3220 & ~n4447 ;
  assign n10391 = n1994 & n10390 ;
  assign n10392 = n10391 ^ n1182 ^ 1'b0 ;
  assign n10393 = ( ~n1817 & n2159 ) | ( ~n1817 & n7926 ) | ( n2159 & n7926 ) ;
  assign n10394 = ~n542 & n7504 ;
  assign n10395 = n3213 & ~n3752 ;
  assign n10396 = n9452 ^ n4508 ^ n943 ;
  assign n10397 = ( n2045 & ~n6718 ) | ( n2045 & n10396 ) | ( ~n6718 & n10396 ) ;
  assign n10398 = n10397 ^ n1908 ^ 1'b0 ;
  assign n10399 = n4157 | n5560 ;
  assign n10400 = n3468 ^ n645 ^ 1'b0 ;
  assign n10401 = n6972 | n10400 ;
  assign n10402 = n10401 ^ n7662 ^ 1'b0 ;
  assign n10403 = ~n783 & n10402 ;
  assign n10404 = ( ~n4030 & n8970 ) | ( ~n4030 & n10403 ) | ( n8970 & n10403 ) ;
  assign n10405 = ~n4089 & n10404 ;
  assign n10406 = ( n1008 & ~n1578 ) | ( n1008 & n2837 ) | ( ~n1578 & n2837 ) ;
  assign n10407 = n8738 | n10406 ;
  assign n10408 = ~x105 & n10407 ;
  assign n10409 = ( n201 & n4770 ) | ( n201 & ~n10408 ) | ( n4770 & ~n10408 ) ;
  assign n10410 = n2008 ^ n609 ^ n352 ;
  assign n10411 = ~n1380 & n2661 ;
  assign n10412 = n10411 ^ n2967 ^ 1'b0 ;
  assign n10413 = ( n8807 & ~n10410 ) | ( n8807 & n10412 ) | ( ~n10410 & n10412 ) ;
  assign n10414 = n10413 ^ n4081 ^ 1'b0 ;
  assign n10415 = n10409 & ~n10414 ;
  assign n10416 = ( ~n5155 & n5746 ) | ( ~n5155 & n6640 ) | ( n5746 & n6640 ) ;
  assign n10417 = ( n1821 & ~n5487 ) | ( n1821 & n10416 ) | ( ~n5487 & n10416 ) ;
  assign n10418 = n10417 ^ n5299 ^ 1'b0 ;
  assign n10419 = n10415 & ~n10418 ;
  assign n10420 = n9350 ^ n432 ^ 1'b0 ;
  assign n10421 = ( x10 & n2716 ) | ( x10 & ~n8934 ) | ( n2716 & ~n8934 ) ;
  assign n10422 = ~n9043 & n10166 ;
  assign n10423 = ~n2057 & n6091 ;
  assign n10424 = n10423 ^ n1266 ^ 1'b0 ;
  assign n10425 = ( ~n8125 & n10422 ) | ( ~n8125 & n10424 ) | ( n10422 & n10424 ) ;
  assign n10426 = n7405 ^ n3362 ^ 1'b0 ;
  assign n10427 = n2950 & n10426 ;
  assign n10439 = n6695 ^ n5635 ^ n4860 ;
  assign n10437 = n1668 ^ n716 ^ 1'b0 ;
  assign n10435 = n1012 | n3924 ;
  assign n10436 = ~n3385 & n10435 ;
  assign n10438 = n10437 ^ n10436 ^ 1'b0 ;
  assign n10440 = n10439 ^ n10438 ^ 1'b0 ;
  assign n10441 = n1955 | n10440 ;
  assign n10433 = n10359 ^ n5396 ^ 1'b0 ;
  assign n10434 = n4420 & ~n10433 ;
  assign n10428 = ( n1275 & n4684 ) | ( n1275 & ~n9905 ) | ( n4684 & ~n9905 ) ;
  assign n10429 = n4691 ^ n3953 ^ n1714 ;
  assign n10430 = ( n3827 & n10428 ) | ( n3827 & n10429 ) | ( n10428 & n10429 ) ;
  assign n10431 = x100 & n10430 ;
  assign n10432 = ~x106 & n10431 ;
  assign n10442 = n10441 ^ n10434 ^ n10432 ;
  assign n10443 = n2171 & ~n5482 ;
  assign n10444 = n7414 ^ n1583 ^ 1'b0 ;
  assign n10445 = n1529 & ~n10444 ;
  assign n10446 = n10445 ^ n9547 ^ 1'b0 ;
  assign n10451 = n1141 | n1720 ;
  assign n10447 = n4033 ^ n2712 ^ n181 ;
  assign n10448 = n6881 ^ n3145 ^ x31 ;
  assign n10449 = ( ~n3118 & n10447 ) | ( ~n3118 & n10448 ) | ( n10447 & n10448 ) ;
  assign n10450 = ~n8685 & n10449 ;
  assign n10452 = n10451 ^ n10450 ^ 1'b0 ;
  assign n10453 = ( n786 & n871 ) | ( n786 & ~n1378 ) | ( n871 & ~n1378 ) ;
  assign n10454 = n464 | n3747 ;
  assign n10455 = n3744 & n6381 ;
  assign n10456 = n10087 & n10455 ;
  assign n10457 = ( ~n308 & n4055 ) | ( ~n308 & n4196 ) | ( n4055 & n4196 ) ;
  assign n10458 = ~n10456 & n10457 ;
  assign n10459 = n10458 ^ n437 ^ 1'b0 ;
  assign n10460 = n3501 & ~n10459 ;
  assign n10461 = n10460 ^ n8760 ^ 1'b0 ;
  assign n10462 = n6262 & n8087 ;
  assign n10463 = ( n156 & n2938 ) | ( n156 & n7944 ) | ( n2938 & n7944 ) ;
  assign n10464 = n615 ^ n337 ^ 1'b0 ;
  assign n10465 = ~n4795 & n10464 ;
  assign n10466 = n10465 ^ n3398 ^ n3196 ;
  assign n10467 = n1374 & n10466 ;
  assign n10468 = n10467 ^ n6822 ^ 1'b0 ;
  assign n10469 = x61 & n2943 ;
  assign n10470 = n5957 & n7938 ;
  assign n10471 = ( ~n7644 & n10469 ) | ( ~n7644 & n10470 ) | ( n10469 & n10470 ) ;
  assign n10472 = ( n3536 & n6914 ) | ( n3536 & n8014 ) | ( n6914 & n8014 ) ;
  assign n10473 = n10022 ^ n2448 ^ 1'b0 ;
  assign n10474 = ~n9828 & n10473 ;
  assign n10475 = n6453 & ~n10474 ;
  assign n10476 = ( ~n3963 & n10472 ) | ( ~n3963 & n10475 ) | ( n10472 & n10475 ) ;
  assign n10477 = n10476 ^ n3105 ^ 1'b0 ;
  assign n10478 = n10471 & n10477 ;
  assign n10479 = n6730 ^ n3488 ^ 1'b0 ;
  assign n10480 = n10479 ^ n4739 ^ 1'b0 ;
  assign n10484 = n1291 & ~n4354 ;
  assign n10481 = n2568 ^ n1656 ^ n1052 ;
  assign n10482 = n10481 ^ n3696 ^ n3148 ;
  assign n10483 = n568 | n10482 ;
  assign n10485 = n10484 ^ n10483 ^ 1'b0 ;
  assign n10486 = n990 ^ n418 ^ 1'b0 ;
  assign n10487 = n8477 ^ n3742 ^ 1'b0 ;
  assign n10488 = n10486 & n10487 ;
  assign n10489 = ( n1911 & ~n2073 ) | ( n1911 & n10488 ) | ( ~n2073 & n10488 ) ;
  assign n10490 = n2581 | n10489 ;
  assign n10491 = n10490 ^ n6300 ^ 1'b0 ;
  assign n10497 = n5158 ^ n3703 ^ n1553 ;
  assign n10492 = n367 | n878 ;
  assign n10493 = n2226 & ~n10492 ;
  assign n10494 = ~n2542 & n9015 ;
  assign n10495 = n1896 | n10494 ;
  assign n10496 = n10493 & ~n10495 ;
  assign n10498 = n10497 ^ n10496 ^ n1152 ;
  assign n10499 = ( n3420 & ~n3647 ) | ( n3420 & n4440 ) | ( ~n3647 & n4440 ) ;
  assign n10500 = n6533 ^ n6324 ^ 1'b0 ;
  assign n10501 = n1204 & n2661 ;
  assign n10502 = n3748 & n10501 ;
  assign n10503 = n5611 & n10502 ;
  assign n10504 = ( n834 & ~n1210 ) | ( n834 & n4750 ) | ( ~n1210 & n4750 ) ;
  assign n10505 = n10504 ^ n8633 ^ n5411 ;
  assign n10506 = n10505 ^ n6686 ^ 1'b0 ;
  assign n10507 = n10503 | n10506 ;
  assign n10508 = n10507 ^ n5536 ^ n1847 ;
  assign n10518 = n1219 & n1732 ;
  assign n10509 = n906 | n2165 ;
  assign n10510 = x80 | n10509 ;
  assign n10512 = n3269 ^ n2033 ^ 1'b0 ;
  assign n10513 = n8677 & n10512 ;
  assign n10514 = n10513 ^ n9440 ^ 1'b0 ;
  assign n10515 = n4320 & n10514 ;
  assign n10511 = n6802 | n8368 ;
  assign n10516 = n10515 ^ n10511 ^ 1'b0 ;
  assign n10517 = n10510 & n10516 ;
  assign n10519 = n10518 ^ n10517 ^ 1'b0 ;
  assign n10520 = n5080 & n10519 ;
  assign n10521 = ~n6420 & n10520 ;
  assign n10522 = n2021 & n4492 ;
  assign n10523 = n7497 & n10522 ;
  assign n10526 = n4957 ^ n2275 ^ n1192 ;
  assign n10524 = n569 | n2073 ;
  assign n10525 = n10524 ^ n9165 ^ 1'b0 ;
  assign n10527 = n10526 ^ n10525 ^ n2089 ;
  assign n10528 = n6693 ^ n5166 ^ n3164 ;
  assign n10529 = n9558 ^ n7488 ^ 1'b0 ;
  assign n10530 = ~n2217 & n10529 ;
  assign n10531 = n10528 & n10530 ;
  assign n10532 = n10531 ^ n9905 ^ 1'b0 ;
  assign n10533 = ( n1750 & n1929 ) | ( n1750 & ~n2989 ) | ( n1929 & ~n2989 ) ;
  assign n10534 = n3334 & n5031 ;
  assign n10535 = ~n3704 & n10534 ;
  assign n10536 = n6831 & n10535 ;
  assign n10537 = n10536 ^ n4322 ^ 1'b0 ;
  assign n10538 = n999 | n10537 ;
  assign n10539 = n10533 & ~n10538 ;
  assign n10540 = ( n1183 & n5612 ) | ( n1183 & ~n7062 ) | ( n5612 & ~n7062 ) ;
  assign n10541 = n7088 ^ n2713 ^ 1'b0 ;
  assign n10542 = n8406 & ~n10541 ;
  assign n10543 = n10542 ^ n6992 ^ n4651 ;
  assign n10544 = n3647 & n10543 ;
  assign n10545 = n5978 ^ n2446 ^ n1465 ;
  assign n10546 = n10545 ^ n6677 ^ n1265 ;
  assign n10547 = n10546 ^ n1305 ^ 1'b0 ;
  assign n10548 = ( ~n6445 & n10544 ) | ( ~n6445 & n10547 ) | ( n10544 & n10547 ) ;
  assign n10549 = ~n1694 & n8201 ;
  assign n10550 = n10549 ^ n2488 ^ 1'b0 ;
  assign n10551 = ( n1298 & n3892 ) | ( n1298 & n5773 ) | ( n3892 & n5773 ) ;
  assign n10552 = n10551 ^ n8812 ^ 1'b0 ;
  assign n10553 = n9575 & ~n10552 ;
  assign n10554 = n1148 & n6612 ;
  assign n10555 = n3061 & n10554 ;
  assign n10556 = n4966 | n7848 ;
  assign n10557 = n10555 & ~n10556 ;
  assign n10558 = n282 & ~n2802 ;
  assign n10559 = ~n6989 & n10558 ;
  assign n10560 = n6508 & n10559 ;
  assign n10564 = n6881 ^ n1443 ^ 1'b0 ;
  assign n10565 = ( ~n550 & n780 ) | ( ~n550 & n10564 ) | ( n780 & n10564 ) ;
  assign n10566 = n10565 ^ n5616 ^ 1'b0 ;
  assign n10567 = n5661 ^ n2264 ^ n1841 ;
  assign n10568 = n10567 ^ n5126 ^ n1666 ;
  assign n10569 = n10568 ^ n2581 ^ 1'b0 ;
  assign n10570 = ( ~n1468 & n3540 ) | ( ~n1468 & n10569 ) | ( n3540 & n10569 ) ;
  assign n10571 = ( ~n2456 & n10566 ) | ( ~n2456 & n10570 ) | ( n10566 & n10570 ) ;
  assign n10563 = ( ~n2419 & n4843 ) | ( ~n2419 & n10022 ) | ( n4843 & n10022 ) ;
  assign n10561 = n7323 ^ n825 ^ 1'b0 ;
  assign n10562 = n3967 & ~n10561 ;
  assign n10572 = n10571 ^ n10563 ^ n10562 ;
  assign n10573 = ( n5057 & n6519 ) | ( n5057 & n10572 ) | ( n6519 & n10572 ) ;
  assign n10574 = ~n1317 & n10573 ;
  assign n10576 = n9818 ^ n8761 ^ 1'b0 ;
  assign n10577 = n1455 & ~n10576 ;
  assign n10575 = n1016 ^ n800 ^ 1'b0 ;
  assign n10578 = n10577 ^ n10575 ^ n9477 ;
  assign n10579 = n7982 & n10578 ;
  assign n10580 = n10579 ^ n5439 ^ 1'b0 ;
  assign n10581 = n4880 ^ n4280 ^ 1'b0 ;
  assign n10582 = n10581 ^ n6152 ^ 1'b0 ;
  assign n10583 = ~n652 & n10582 ;
  assign n10584 = n6705 ^ n3021 ^ 1'b0 ;
  assign n10585 = n10584 ^ n7888 ^ 1'b0 ;
  assign n10586 = n2339 | n10585 ;
  assign n10587 = n5314 ^ n2485 ^ n861 ;
  assign n10588 = n10587 ^ n10194 ^ 1'b0 ;
  assign n10589 = ~n195 & n1494 ;
  assign n10590 = ( n1533 & n5670 ) | ( n1533 & n10589 ) | ( n5670 & n10589 ) ;
  assign n10591 = n9118 ^ n4547 ^ n395 ;
  assign n10595 = ( ~n1248 & n3932 ) | ( ~n1248 & n4819 ) | ( n3932 & n4819 ) ;
  assign n10592 = n4208 | n8721 ;
  assign n10593 = n1285 ^ n376 ^ 1'b0 ;
  assign n10594 = ( n4960 & n10592 ) | ( n4960 & ~n10593 ) | ( n10592 & ~n10593 ) ;
  assign n10596 = n10595 ^ n10594 ^ n7883 ;
  assign n10598 = n6460 ^ n143 ^ 1'b0 ;
  assign n10599 = ( n888 & n7932 ) | ( n888 & n10598 ) | ( n7932 & n10598 ) ;
  assign n10597 = ~n1361 & n8927 ;
  assign n10600 = n10599 ^ n10597 ^ n7648 ;
  assign n10601 = n6832 ^ n6094 ^ 1'b0 ;
  assign n10602 = n1690 & n10601 ;
  assign n10603 = n1346 ^ n897 ^ 1'b0 ;
  assign n10604 = n8962 & ~n10603 ;
  assign n10605 = n10057 ^ n6313 ^ x62 ;
  assign n10606 = ( ~n1369 & n4457 ) | ( ~n1369 & n10605 ) | ( n4457 & n10605 ) ;
  assign n10608 = n3442 ^ n3045 ^ n2898 ;
  assign n10609 = n10608 ^ n6297 ^ n1719 ;
  assign n10607 = n2734 | n7250 ;
  assign n10610 = n10609 ^ n10607 ^ 1'b0 ;
  assign n10611 = ( ~n763 & n7661 ) | ( ~n763 & n10610 ) | ( n7661 & n10610 ) ;
  assign n10612 = n911 | n4088 ;
  assign n10613 = n10612 ^ n9545 ^ 1'b0 ;
  assign n10614 = ( n1342 & ~n7419 ) | ( n1342 & n9627 ) | ( ~n7419 & n9627 ) ;
  assign n10615 = n7122 ^ n5749 ^ n5466 ;
  assign n10616 = x106 & n397 ;
  assign n10617 = ~n2021 & n10616 ;
  assign n10618 = n1313 & n8390 ;
  assign n10619 = n2900 & n10618 ;
  assign n10620 = n1475 ^ x15 ^ 1'b0 ;
  assign n10621 = ~n1315 & n8753 ;
  assign n10622 = ~n10620 & n10621 ;
  assign n10623 = n10482 ^ n3176 ^ n2514 ;
  assign n10624 = ( n3201 & n5641 ) | ( n3201 & n6403 ) | ( n5641 & n6403 ) ;
  assign n10625 = n6255 ^ n5011 ^ n1473 ;
  assign n10626 = ( ~n5723 & n10624 ) | ( ~n5723 & n10625 ) | ( n10624 & n10625 ) ;
  assign n10627 = ( n8004 & n8343 ) | ( n8004 & n8658 ) | ( n8343 & n8658 ) ;
  assign n10628 = n10626 & ~n10627 ;
  assign n10629 = ~n10623 & n10628 ;
  assign n10630 = n8324 & n8922 ;
  assign n10636 = ( x105 & ~n5854 ) | ( x105 & n8127 ) | ( ~n5854 & n8127 ) ;
  assign n10637 = n815 ^ n690 ^ 1'b0 ;
  assign n10638 = n10636 & ~n10637 ;
  assign n10634 = ( n1023 & ~n4018 ) | ( n1023 & n7397 ) | ( ~n4018 & n7397 ) ;
  assign n10631 = n847 & ~n2363 ;
  assign n10632 = ( n1850 & n5650 ) | ( n1850 & n7282 ) | ( n5650 & n7282 ) ;
  assign n10633 = ( n3716 & n10631 ) | ( n3716 & n10632 ) | ( n10631 & n10632 ) ;
  assign n10635 = n10634 ^ n10633 ^ 1'b0 ;
  assign n10639 = n10638 ^ n10635 ^ 1'b0 ;
  assign n10640 = n1095 & ~n3745 ;
  assign n10641 = n2411 | n4954 ;
  assign n10642 = n10641 ^ n4245 ^ 1'b0 ;
  assign n10643 = ~n8151 & n10642 ;
  assign n10644 = n10640 & n10643 ;
  assign n10645 = n6513 ^ n857 ^ 1'b0 ;
  assign n10646 = n10644 | n10645 ;
  assign n10647 = n10646 ^ n2807 ^ 1'b0 ;
  assign n10648 = n10647 ^ n3070 ^ 1'b0 ;
  assign n10650 = n2815 ^ n581 ^ n572 ;
  assign n10649 = n2293 | n5597 ;
  assign n10651 = n10650 ^ n10649 ^ n6663 ;
  assign n10652 = n9003 ^ n3452 ^ 1'b0 ;
  assign n10653 = ~n8383 & n10652 ;
  assign n10659 = n192 & n1590 ;
  assign n10654 = n540 | n8625 ;
  assign n10655 = n2247 & ~n10654 ;
  assign n10656 = n10655 ^ n4259 ^ n1448 ;
  assign n10657 = ~n2714 & n10656 ;
  assign n10658 = ~n5023 & n10657 ;
  assign n10660 = n10659 ^ n10658 ^ 1'b0 ;
  assign n10661 = ( n2269 & n2905 ) | ( n2269 & ~n4200 ) | ( n2905 & ~n4200 ) ;
  assign n10662 = ( n409 & ~n2778 ) | ( n409 & n5362 ) | ( ~n2778 & n5362 ) ;
  assign n10663 = ( ~n6369 & n10661 ) | ( ~n6369 & n10662 ) | ( n10661 & n10662 ) ;
  assign n10664 = n3207 ^ n2724 ^ 1'b0 ;
  assign n10665 = n5471 ^ n3360 ^ 1'b0 ;
  assign n10666 = n3106 & ~n10665 ;
  assign n10667 = n10666 ^ n386 ^ 1'b0 ;
  assign n10668 = ~n5775 & n10667 ;
  assign n10669 = n10668 ^ n9238 ^ n2255 ;
  assign n10670 = ( ~n4385 & n5324 ) | ( ~n4385 & n6425 ) | ( n5324 & n6425 ) ;
  assign n10671 = n10202 ^ n7549 ^ 1'b0 ;
  assign n10672 = n3028 | n10671 ;
  assign n10673 = n7776 ^ n4146 ^ n1277 ;
  assign n10674 = ~n8915 & n10673 ;
  assign n10675 = n1900 & ~n2959 ;
  assign n10676 = n1863 & n10675 ;
  assign n10677 = ( x26 & n2323 ) | ( x26 & n10676 ) | ( n2323 & n10676 ) ;
  assign n10678 = n10677 ^ n7712 ^ n3461 ;
  assign n10679 = n2258 & n10678 ;
  assign n10680 = n1646 & ~n7337 ;
  assign n10681 = ~n10679 & n10680 ;
  assign n10682 = n926 & ~n4865 ;
  assign n10683 = ( n519 & n2957 ) | ( n519 & n5587 ) | ( n2957 & n5587 ) ;
  assign n10684 = n2698 ^ n304 ^ 1'b0 ;
  assign n10685 = n10684 ^ n1515 ^ 1'b0 ;
  assign n10690 = n10493 ^ n9259 ^ x121 ;
  assign n10691 = n1029 | n10690 ;
  assign n10686 = ~n972 & n7008 ;
  assign n10687 = ~n3795 & n10686 ;
  assign n10688 = n10687 ^ n7224 ^ 1'b0 ;
  assign n10689 = ( ~n1958 & n3398 ) | ( ~n1958 & n10688 ) | ( n3398 & n10688 ) ;
  assign n10692 = n10691 ^ n10689 ^ n6392 ;
  assign n10693 = n9781 ^ n650 ^ 1'b0 ;
  assign n10694 = n6624 | n10693 ;
  assign n10695 = n1220 ^ n260 ^ 1'b0 ;
  assign n10696 = n2991 | n6750 ;
  assign n10697 = n3886 | n10696 ;
  assign n10698 = n6238 ^ n3272 ^ n2484 ;
  assign n10699 = ( ~n10695 & n10697 ) | ( ~n10695 & n10698 ) | ( n10697 & n10698 ) ;
  assign n10700 = ( ~n965 & n4875 ) | ( ~n965 & n6659 ) | ( n4875 & n6659 ) ;
  assign n10701 = n401 & n10700 ;
  assign n10710 = n353 & ~n934 ;
  assign n10711 = n810 & n10710 ;
  assign n10705 = n950 & ~n3144 ;
  assign n10706 = ~n3404 & n10705 ;
  assign n10707 = n9892 & ~n10706 ;
  assign n10708 = n10707 ^ n5519 ^ 1'b0 ;
  assign n10709 = ~n2524 & n10708 ;
  assign n10702 = ( n1208 & n4103 ) | ( n1208 & ~n8916 ) | ( n4103 & ~n8916 ) ;
  assign n10703 = n6617 ^ n2057 ^ n853 ;
  assign n10704 = ( n1926 & n10702 ) | ( n1926 & n10703 ) | ( n10702 & n10703 ) ;
  assign n10712 = n10711 ^ n10709 ^ n10704 ;
  assign n10713 = n2088 ^ n1500 ^ n1292 ;
  assign n10714 = n2459 & ~n10713 ;
  assign n10715 = n6860 & n10714 ;
  assign n10716 = n6481 ^ n1065 ^ 1'b0 ;
  assign n10717 = n10715 | n10716 ;
  assign n10718 = n4888 | n10717 ;
  assign n10719 = ~n7180 & n10718 ;
  assign n10720 = n3364 ^ n532 ^ 1'b0 ;
  assign n10721 = ~n934 & n10720 ;
  assign n10722 = n10721 ^ n7847 ^ 1'b0 ;
  assign n10723 = n3819 | n10722 ;
  assign n10724 = n10723 ^ n9876 ^ 1'b0 ;
  assign n10725 = ~n3749 & n10724 ;
  assign n10726 = ( n1308 & n2399 ) | ( n1308 & n3562 ) | ( n2399 & n3562 ) ;
  assign n10727 = ( n201 & n1251 ) | ( n201 & n3740 ) | ( n1251 & n3740 ) ;
  assign n10728 = ~n2541 & n2559 ;
  assign n10729 = ~n10727 & n10728 ;
  assign n10730 = n10726 | n10729 ;
  assign n10731 = n10725 | n10730 ;
  assign n10732 = ~n489 & n10731 ;
  assign n10733 = n10356 ^ n8673 ^ 1'b0 ;
  assign n10734 = n2526 & ~n4971 ;
  assign n10735 = n551 & n10734 ;
  assign n10736 = ~n10235 & n10735 ;
  assign n10737 = ( n3602 & n4761 ) | ( n3602 & n5172 ) | ( n4761 & n5172 ) ;
  assign n10738 = ( x106 & n6880 ) | ( x106 & n10737 ) | ( n6880 & n10737 ) ;
  assign n10739 = ( n181 & n778 ) | ( n181 & ~n6093 ) | ( n778 & ~n6093 ) ;
  assign n10740 = n1915 ^ n1169 ^ n606 ;
  assign n10741 = n6914 ^ n2089 ^ 1'b0 ;
  assign n10742 = n10740 & ~n10741 ;
  assign n10743 = ( x56 & n573 ) | ( x56 & ~n6970 ) | ( n573 & ~n6970 ) ;
  assign n10744 = n10743 ^ n8381 ^ n3196 ;
  assign n10745 = ( n4215 & n5849 ) | ( n4215 & ~n10744 ) | ( n5849 & ~n10744 ) ;
  assign n10746 = n10309 ^ n509 ^ 1'b0 ;
  assign n10747 = n10746 ^ n4464 ^ 1'b0 ;
  assign n10748 = ( ~n10742 & n10745 ) | ( ~n10742 & n10747 ) | ( n10745 & n10747 ) ;
  assign n10753 = ( n273 & n3450 ) | ( n273 & ~n5627 ) | ( n3450 & ~n5627 ) ;
  assign n10754 = n10753 ^ n2083 ^ 1'b0 ;
  assign n10755 = ( x107 & n1557 ) | ( x107 & n6460 ) | ( n1557 & n6460 ) ;
  assign n10756 = n10755 ^ n7302 ^ n1026 ;
  assign n10757 = n10756 ^ n7058 ^ 1'b0 ;
  assign n10758 = n10754 | n10757 ;
  assign n10749 = n8854 ^ n2181 ^ 1'b0 ;
  assign n10750 = n10749 ^ n5516 ^ n5139 ;
  assign n10751 = n10750 ^ n5624 ^ 1'b0 ;
  assign n10752 = n6232 | n10751 ;
  assign n10759 = n10758 ^ n10752 ^ n604 ;
  assign n10760 = n10748 | n10759 ;
  assign n10761 = n10739 | n10760 ;
  assign n10762 = ( n378 & n1960 ) | ( n378 & ~n3595 ) | ( n1960 & ~n3595 ) ;
  assign n10763 = n10762 ^ n234 ^ 1'b0 ;
  assign n10764 = n605 & n10763 ;
  assign n10768 = n6564 ^ n3300 ^ 1'b0 ;
  assign n10769 = n6507 | n10768 ;
  assign n10765 = ( ~n3922 & n4240 ) | ( ~n3922 & n7665 ) | ( n4240 & n7665 ) ;
  assign n10766 = ~n1824 & n1896 ;
  assign n10767 = ~n10765 & n10766 ;
  assign n10770 = n10769 ^ n10767 ^ n8754 ;
  assign n10771 = n8592 ^ n3298 ^ 1'b0 ;
  assign n10774 = ( ~x37 & n133 ) | ( ~x37 & n839 ) | ( n133 & n839 ) ;
  assign n10773 = n8597 ^ n6644 ^ 1'b0 ;
  assign n10775 = n10774 ^ n10773 ^ n189 ;
  assign n10772 = n8781 ^ n2159 ^ 1'b0 ;
  assign n10776 = n10775 ^ n10772 ^ n10534 ;
  assign n10777 = ( n8117 & n10771 ) | ( n8117 & ~n10776 ) | ( n10771 & ~n10776 ) ;
  assign n10778 = n5224 & n6669 ;
  assign n10779 = ( ~n1015 & n1829 ) | ( ~n1015 & n2602 ) | ( n1829 & n2602 ) ;
  assign n10780 = ( n4905 & ~n5669 ) | ( n4905 & n10779 ) | ( ~n5669 & n10779 ) ;
  assign n10783 = n1085 & ~n9821 ;
  assign n10784 = n10783 ^ n2634 ^ 1'b0 ;
  assign n10785 = ( n6519 & ~n7277 ) | ( n6519 & n10784 ) | ( ~n7277 & n10784 ) ;
  assign n10781 = n4647 & n7177 ;
  assign n10782 = n6883 & n10781 ;
  assign n10786 = n10785 ^ n10782 ^ n6747 ;
  assign n10787 = n9889 ^ n5155 ^ n3776 ;
  assign n10788 = ~n9146 & n10787 ;
  assign n10789 = ( n4544 & ~n4825 ) | ( n4544 & n8833 ) | ( ~n4825 & n8833 ) ;
  assign n10790 = ( n4758 & n6371 ) | ( n4758 & n9506 ) | ( n6371 & n9506 ) ;
  assign n10791 = ~n2869 & n10790 ;
  assign n10792 = ( n275 & n5165 ) | ( n275 & ~n8997 ) | ( n5165 & ~n8997 ) ;
  assign n10793 = n8465 | n10792 ;
  assign n10794 = n8443 & ~n10793 ;
  assign n10795 = ~x30 & n1248 ;
  assign n10796 = n4386 ^ x42 ^ 1'b0 ;
  assign n10797 = n5135 & n10796 ;
  assign n10798 = n10459 ^ n10223 ^ 1'b0 ;
  assign n10799 = n1084 & n10798 ;
  assign n10800 = n489 & n1443 ;
  assign n10801 = n3528 & n10800 ;
  assign n10802 = n2060 & ~n9735 ;
  assign n10803 = n10802 ^ n3344 ^ 1'b0 ;
  assign n10804 = n10125 ^ n6250 ^ 1'b0 ;
  assign n10805 = n2716 & n10804 ;
  assign n10806 = n10805 ^ n2072 ^ 1'b0 ;
  assign n10807 = n4453 | n10806 ;
  assign n10808 = n10807 ^ n712 ^ 1'b0 ;
  assign n10809 = ~n184 & n5558 ;
  assign n10810 = n6290 & n10809 ;
  assign n10811 = n10810 ^ n5550 ^ 1'b0 ;
  assign n10812 = ~n10808 & n10811 ;
  assign n10813 = n10812 ^ n3357 ^ 1'b0 ;
  assign n10817 = ( ~x34 & n1989 ) | ( ~x34 & n9847 ) | ( n1989 & n9847 ) ;
  assign n10818 = n10347 ^ n2256 ^ 1'b0 ;
  assign n10819 = n3667 ^ n1929 ^ n625 ;
  assign n10820 = n10819 ^ n10057 ^ 1'b0 ;
  assign n10821 = n8422 & n10820 ;
  assign n10822 = ( n10817 & n10818 ) | ( n10817 & ~n10821 ) | ( n10818 & ~n10821 ) ;
  assign n10814 = n499 & ~n5156 ;
  assign n10815 = n9845 ^ n5471 ^ 1'b0 ;
  assign n10816 = ( n8559 & n10814 ) | ( n8559 & ~n10815 ) | ( n10814 & ~n10815 ) ;
  assign n10823 = n10822 ^ n10816 ^ n9772 ;
  assign n10829 = n632 | n2402 ;
  assign n10830 = n10829 ^ n8505 ^ 1'b0 ;
  assign n10831 = n9378 & n10830 ;
  assign n10832 = n10831 ^ n2118 ^ 1'b0 ;
  assign n10827 = n5076 ^ n4953 ^ 1'b0 ;
  assign n10824 = ( n297 & n370 ) | ( n297 & ~n3676 ) | ( n370 & ~n3676 ) ;
  assign n10825 = n3148 ^ n609 ^ 1'b0 ;
  assign n10826 = ( n6742 & n10824 ) | ( n6742 & ~n10825 ) | ( n10824 & ~n10825 ) ;
  assign n10828 = n10827 ^ n10826 ^ n4096 ;
  assign n10833 = n10832 ^ n10828 ^ n4815 ;
  assign n10834 = n2976 | n8943 ;
  assign n10835 = n7992 ^ n7041 ^ n1378 ;
  assign n10836 = ( n4614 & ~n7042 ) | ( n4614 & n10835 ) | ( ~n7042 & n10835 ) ;
  assign n10837 = n1010 | n2625 ;
  assign n10838 = n10837 ^ n1061 ^ 1'b0 ;
  assign n10839 = x74 & ~n2402 ;
  assign n10840 = n10839 ^ n317 ^ 1'b0 ;
  assign n10841 = n10840 ^ n6934 ^ 1'b0 ;
  assign n10842 = n4043 ^ n948 ^ 1'b0 ;
  assign n10843 = n10842 ^ n9835 ^ n635 ;
  assign n10845 = ( n1780 & n2338 ) | ( n1780 & n2943 ) | ( n2338 & n2943 ) ;
  assign n10846 = n2757 & ~n10845 ;
  assign n10847 = ~x29 & n10846 ;
  assign n10848 = n9366 ^ n7518 ^ n2114 ;
  assign n10849 = ( n4208 & ~n10847 ) | ( n4208 & n10848 ) | ( ~n10847 & n10848 ) ;
  assign n10844 = n6140 & ~n10397 ;
  assign n10850 = n10849 ^ n10844 ^ 1'b0 ;
  assign n10851 = n4226 ^ n592 ^ 1'b0 ;
  assign n10852 = n2016 & n10851 ;
  assign n10853 = n10852 ^ n4238 ^ n1193 ;
  assign n10854 = n9282 ^ n853 ^ 1'b0 ;
  assign n10855 = n10853 & n10854 ;
  assign n10856 = n2227 ^ n310 ^ n240 ;
  assign n10857 = n5304 | n5948 ;
  assign n10858 = ~n10856 & n10857 ;
  assign n10859 = ~n10449 & n10858 ;
  assign n10860 = n1147 | n10859 ;
  assign n10861 = n9335 | n10860 ;
  assign n10862 = n10861 ^ n5123 ^ 1'b0 ;
  assign n10863 = n10862 ^ n9890 ^ n2471 ;
  assign n10864 = n1838 ^ n990 ^ 1'b0 ;
  assign n10865 = n8013 ^ n285 ^ x116 ;
  assign n10866 = n10864 | n10865 ;
  assign n10867 = ( n9297 & n10863 ) | ( n9297 & n10866 ) | ( n10863 & n10866 ) ;
  assign n10868 = n8658 ^ n4024 ^ n757 ;
  assign n10869 = n10868 ^ n3054 ^ 1'b0 ;
  assign n10873 = ( ~n674 & n2456 ) | ( ~n674 & n5164 ) | ( n2456 & n5164 ) ;
  assign n10870 = n8391 ^ n5021 ^ n915 ;
  assign n10871 = ( n1898 & ~n2583 ) | ( n1898 & n10870 ) | ( ~n2583 & n10870 ) ;
  assign n10872 = ~n8729 & n10871 ;
  assign n10874 = n10873 ^ n10872 ^ 1'b0 ;
  assign n10875 = ( n1566 & n2778 ) | ( n1566 & n10874 ) | ( n2778 & n10874 ) ;
  assign n10876 = n4010 ^ n2264 ^ 1'b0 ;
  assign n10877 = ( n1240 & ~n7757 ) | ( n1240 & n10876 ) | ( ~n7757 & n10876 ) ;
  assign n10878 = n10877 ^ n4864 ^ n3127 ;
  assign n10880 = n6015 ^ n5757 ^ n949 ;
  assign n10879 = n9584 ^ n1304 ^ 1'b0 ;
  assign n10881 = n10880 ^ n10879 ^ 1'b0 ;
  assign n10882 = n10878 & n10881 ;
  assign n10883 = n2840 & n5785 ;
  assign n10884 = ~n5539 & n10883 ;
  assign n10885 = n10884 ^ n8157 ^ 1'b0 ;
  assign n10886 = n1572 | n2954 ;
  assign n10887 = n334 ^ n166 ^ 1'b0 ;
  assign n10888 = n3188 & ~n10887 ;
  assign n10892 = n9835 ^ n5429 ^ n5129 ;
  assign n10889 = n758 & ~n2118 ;
  assign n10890 = ( n4237 & n5706 ) | ( n4237 & ~n10277 ) | ( n5706 & ~n10277 ) ;
  assign n10891 = ~n10889 & n10890 ;
  assign n10893 = n10892 ^ n10891 ^ 1'b0 ;
  assign n10894 = n4453 ^ n1030 ^ 1'b0 ;
  assign n10895 = n5356 & ~n10894 ;
  assign n10896 = ~n4757 & n10895 ;
  assign n10897 = n10896 ^ n3080 ^ 1'b0 ;
  assign n10898 = n7101 ^ n4105 ^ n1048 ;
  assign n10899 = n6814 & n10898 ;
  assign n10900 = ~n10897 & n10899 ;
  assign n10905 = n7667 ^ n3344 ^ n2982 ;
  assign n10906 = n433 | n2417 ;
  assign n10907 = n10906 ^ n6516 ^ 1'b0 ;
  assign n10908 = n8215 | n10907 ;
  assign n10909 = n372 | n10908 ;
  assign n10911 = ( n450 & n1623 ) | ( n450 & ~n2312 ) | ( n1623 & ~n2312 ) ;
  assign n10910 = ( ~n748 & n3443 ) | ( ~n748 & n4911 ) | ( n3443 & n4911 ) ;
  assign n10912 = n10911 ^ n10910 ^ n883 ;
  assign n10913 = ( ~x97 & n10482 ) | ( ~x97 & n10912 ) | ( n10482 & n10912 ) ;
  assign n10914 = n10909 & ~n10913 ;
  assign n10915 = n10905 & n10914 ;
  assign n10901 = n5965 ^ n1836 ^ n1641 ;
  assign n10902 = ( n1903 & n6703 ) | ( n1903 & n7691 ) | ( n6703 & n7691 ) ;
  assign n10903 = n10902 ^ n7890 ^ n5732 ;
  assign n10904 = ( ~x92 & n10901 ) | ( ~x92 & n10903 ) | ( n10901 & n10903 ) ;
  assign n10916 = n10915 ^ n10904 ^ x104 ;
  assign n10917 = ( n244 & n954 ) | ( n244 & n2097 ) | ( n954 & n2097 ) ;
  assign n10918 = ( ~n4511 & n8630 ) | ( ~n4511 & n10917 ) | ( n8630 & n10917 ) ;
  assign n10930 = n2681 ^ n1956 ^ x87 ;
  assign n10931 = ( n4081 & n6283 ) | ( n4081 & ~n10930 ) | ( n6283 & ~n10930 ) ;
  assign n10927 = n6103 ^ n4612 ^ n4602 ;
  assign n10928 = ~n7216 & n10927 ;
  assign n10921 = n3945 & ~n7165 ;
  assign n10922 = n10921 ^ n4443 ^ 1'b0 ;
  assign n10923 = n1154 & ~n10922 ;
  assign n10924 = n6017 & n10923 ;
  assign n10919 = n7187 ^ n249 ^ 1'b0 ;
  assign n10920 = n10919 ^ n6071 ^ n5079 ;
  assign n10925 = n10924 ^ n10920 ^ n2636 ;
  assign n10926 = ( ~n4706 & n10335 ) | ( ~n4706 & n10925 ) | ( n10335 & n10925 ) ;
  assign n10929 = n10928 ^ n10926 ^ n1575 ;
  assign n10932 = n10931 ^ n10929 ^ 1'b0 ;
  assign n10933 = n7964 ^ n2167 ^ 1'b0 ;
  assign n10934 = n1674 & n10933 ;
  assign n10935 = n294 | n1874 ;
  assign n10936 = n10934 | n10935 ;
  assign n10940 = n9114 ^ n3808 ^ n1082 ;
  assign n10938 = ~n5781 & n6045 ;
  assign n10939 = n10938 ^ n8960 ^ 1'b0 ;
  assign n10937 = n4096 | n4142 ;
  assign n10941 = n10940 ^ n10939 ^ n10937 ;
  assign n10942 = n5277 ^ n1393 ^ 1'b0 ;
  assign n10943 = n222 & n10942 ;
  assign n10944 = n10943 ^ n10266 ^ 1'b0 ;
  assign n10945 = ( n1285 & n7197 ) | ( n1285 & n9020 ) | ( n7197 & n9020 ) ;
  assign n10946 = n10945 ^ n6766 ^ n2395 ;
  assign n10959 = ~n690 & n6733 ;
  assign n10947 = ( n2083 & ~n2875 ) | ( n2083 & n5980 ) | ( ~n2875 & n5980 ) ;
  assign n10948 = n5892 ^ n3027 ^ n740 ;
  assign n10949 = ~n4755 & n6649 ;
  assign n10950 = ( n1946 & ~n3592 ) | ( n1946 & n7685 ) | ( ~n3592 & n7685 ) ;
  assign n10951 = ~n10949 & n10950 ;
  assign n10952 = n10948 & n10951 ;
  assign n10953 = ( n9000 & ~n10947 ) | ( n9000 & n10952 ) | ( ~n10947 & n10952 ) ;
  assign n10954 = n8424 | n10953 ;
  assign n10955 = n6347 & ~n10954 ;
  assign n10956 = n5026 ^ n4852 ^ 1'b0 ;
  assign n10957 = ~n10955 & n10956 ;
  assign n10958 = n4636 & n10957 ;
  assign n10960 = n10959 ^ n10958 ^ 1'b0 ;
  assign n10961 = n7193 & ~n10960 ;
  assign n10962 = n1907 & ~n10961 ;
  assign n10965 = n957 ^ n624 ^ n203 ;
  assign n10964 = ( ~n570 & n6783 ) | ( ~n570 & n7274 ) | ( n6783 & n7274 ) ;
  assign n10963 = ( n3837 & n6305 ) | ( n3837 & n10308 ) | ( n6305 & n10308 ) ;
  assign n10966 = n10965 ^ n10964 ^ n10963 ;
  assign n10967 = ~n1969 & n10396 ;
  assign n10968 = ~n522 & n10967 ;
  assign n10969 = n10968 ^ n8054 ^ n3700 ;
  assign n10970 = n129 & n7454 ;
  assign n10973 = n8341 ^ n1885 ^ 1'b0 ;
  assign n10971 = n4162 ^ n1130 ^ 1'b0 ;
  assign n10972 = n456 | n10971 ;
  assign n10974 = n10973 ^ n10972 ^ n1959 ;
  assign n10975 = n10974 ^ n6501 ^ n3544 ;
  assign n10976 = ( n7735 & n10970 ) | ( n7735 & ~n10975 ) | ( n10970 & ~n10975 ) ;
  assign n10977 = n10861 ^ n1353 ^ 1'b0 ;
  assign n10978 = n4110 ^ n3412 ^ 1'b0 ;
  assign n10979 = n545 & ~n10978 ;
  assign n10980 = ( ~n1331 & n7302 ) | ( ~n1331 & n10979 ) | ( n7302 & n10979 ) ;
  assign n10981 = n1081 | n7107 ;
  assign n10982 = n10981 ^ n5735 ^ 1'b0 ;
  assign n10983 = ( ~n1158 & n4960 ) | ( ~n1158 & n7898 ) | ( n4960 & n7898 ) ;
  assign n10984 = n10983 ^ n6373 ^ n3511 ;
  assign n10985 = ~n7482 & n10984 ;
  assign n10986 = n7176 & n10985 ;
  assign n10987 = ( n9490 & n9742 ) | ( n9490 & n10986 ) | ( n9742 & n10986 ) ;
  assign n10995 = n4472 & ~n8691 ;
  assign n10990 = ( n1339 & ~n1926 ) | ( n1339 & n3445 ) | ( ~n1926 & n3445 ) ;
  assign n10991 = ( ~n949 & n5776 ) | ( ~n949 & n10990 ) | ( n5776 & n10990 ) ;
  assign n10992 = n3241 ^ n2750 ^ 1'b0 ;
  assign n10993 = ~n10991 & n10992 ;
  assign n10989 = ( ~n927 & n7062 ) | ( ~n927 & n8282 ) | ( n7062 & n8282 ) ;
  assign n10988 = n5039 ^ n1725 ^ 1'b0 ;
  assign n10994 = n10993 ^ n10989 ^ n10988 ;
  assign n10996 = n10995 ^ n10994 ^ 1'b0 ;
  assign n10998 = n2550 | n9125 ;
  assign n10997 = n1465 | n2049 ;
  assign n10999 = n10998 ^ n10997 ^ 1'b0 ;
  assign n11000 = n3292 ^ n2643 ^ n1633 ;
  assign n11001 = ~n10441 & n11000 ;
  assign n11002 = ~x8 & n11001 ;
  assign n11003 = n313 | n6017 ;
  assign n11004 = ( n6984 & n7121 ) | ( n6984 & ~n11003 ) | ( n7121 & ~n11003 ) ;
  assign n11005 = n11004 ^ n7116 ^ n2267 ;
  assign n11006 = n3530 ^ n3021 ^ 1'b0 ;
  assign n11008 = ( n4140 & ~n5342 ) | ( n4140 & n5644 ) | ( ~n5342 & n5644 ) ;
  assign n11007 = n6414 & n8994 ;
  assign n11009 = n11008 ^ n11007 ^ 1'b0 ;
  assign n11010 = n11009 ^ n5185 ^ 1'b0 ;
  assign n11011 = n9082 ^ n8455 ^ n7298 ;
  assign n11012 = n5569 ^ n3280 ^ 1'b0 ;
  assign n11013 = ~n10682 & n11012 ;
  assign n11014 = n4968 ^ n1681 ^ 1'b0 ;
  assign n11015 = n11014 ^ n5320 ^ 1'b0 ;
  assign n11018 = ( ~n4016 & n4514 ) | ( ~n4016 & n4738 ) | ( n4514 & n4738 ) ;
  assign n11016 = ( n129 & n2776 ) | ( n129 & n3940 ) | ( n2776 & n3940 ) ;
  assign n11017 = n11016 ^ n5968 ^ n3771 ;
  assign n11019 = n11018 ^ n11017 ^ n4380 ;
  assign n11020 = n1418 & n4129 ;
  assign n11022 = n2435 & n7665 ;
  assign n11021 = n259 & ~n5256 ;
  assign n11023 = n11022 ^ n11021 ^ n10740 ;
  assign n11024 = n11023 ^ n5366 ^ n4298 ;
  assign n11032 = n1280 ^ n348 ^ 1'b0 ;
  assign n11033 = n6659 | n11032 ;
  assign n11034 = ( n142 & n5408 ) | ( n142 & ~n11033 ) | ( n5408 & ~n11033 ) ;
  assign n11031 = ( ~n2635 & n3925 ) | ( ~n2635 & n5419 ) | ( n3925 & n5419 ) ;
  assign n11035 = n11034 ^ n11031 ^ n2869 ;
  assign n11025 = ~n1219 & n1374 ;
  assign n11026 = ~n673 & n1024 ;
  assign n11027 = n136 & n11026 ;
  assign n11028 = n7241 & n10673 ;
  assign n11029 = n11027 | n11028 ;
  assign n11030 = n11025 | n11029 ;
  assign n11036 = n11035 ^ n11030 ^ 1'b0 ;
  assign n11037 = n1153 & n2904 ;
  assign n11038 = n11037 ^ n313 ^ 1'b0 ;
  assign n11039 = n5731 ^ n5543 ^ 1'b0 ;
  assign n11040 = ~n9086 & n11039 ;
  assign n11041 = ( n6221 & ~n11038 ) | ( n6221 & n11040 ) | ( ~n11038 & n11040 ) ;
  assign n11042 = n3742 & ~n9571 ;
  assign n11043 = n11042 ^ n4629 ^ 1'b0 ;
  assign n11044 = n9706 ^ n7679 ^ n2471 ;
  assign n11053 = ~n381 & n966 ;
  assign n11054 = n11053 ^ n2721 ^ n674 ;
  assign n11055 = n3379 & ~n11054 ;
  assign n11049 = n6437 ^ n4726 ^ n508 ;
  assign n11050 = n1817 ^ x66 ^ 1'b0 ;
  assign n11051 = n11049 & ~n11050 ;
  assign n11045 = n1368 & n8491 ;
  assign n11046 = ~n7654 & n11045 ;
  assign n11047 = n2573 & n8548 ;
  assign n11048 = n11046 & n11047 ;
  assign n11052 = n11051 ^ n11048 ^ n7358 ;
  assign n11056 = n11055 ^ n11052 ^ 1'b0 ;
  assign n11057 = n11044 & n11056 ;
  assign n11058 = n7571 ^ n6662 ^ 1'b0 ;
  assign n11059 = ~n2078 & n10740 ;
  assign n11060 = n424 & n11059 ;
  assign n11064 = n3747 ^ n1117 ^ 1'b0 ;
  assign n11061 = ~n4844 & n4889 ;
  assign n11062 = n11061 ^ n6580 ^ 1'b0 ;
  assign n11063 = ( n1226 & n4257 ) | ( n1226 & n11062 ) | ( n4257 & n11062 ) ;
  assign n11065 = n11064 ^ n11063 ^ 1'b0 ;
  assign n11066 = ~n11060 & n11065 ;
  assign n11068 = n4665 ^ n1960 ^ 1'b0 ;
  assign n11067 = ( n1026 & ~n5807 ) | ( n1026 & n6683 ) | ( ~n5807 & n6683 ) ;
  assign n11069 = n11068 ^ n11067 ^ n8546 ;
  assign n11070 = n8476 ^ n5088 ^ 1'b0 ;
  assign n11071 = ~n3582 & n11070 ;
  assign n11074 = n6675 ^ n2210 ^ n1108 ;
  assign n11073 = ( n1944 & n2046 ) | ( n1944 & n6735 ) | ( n2046 & n6735 ) ;
  assign n11075 = n11074 ^ n11073 ^ n4571 ;
  assign n11076 = n11075 ^ n10238 ^ n4008 ;
  assign n11072 = n1896 & n7998 ;
  assign n11077 = n11076 ^ n11072 ^ 1'b0 ;
  assign n11078 = ( ~n3645 & n4947 ) | ( ~n3645 & n10897 ) | ( n4947 & n10897 ) ;
  assign n11079 = n11078 ^ n3483 ^ x120 ;
  assign n11080 = ( n635 & n4337 ) | ( n635 & n4946 ) | ( n4337 & n4946 ) ;
  assign n11081 = n1371 | n1608 ;
  assign n11084 = n7047 ^ n3636 ^ n3285 ;
  assign n11085 = n1364 & ~n2893 ;
  assign n11086 = ~n11084 & n11085 ;
  assign n11082 = ~n1599 & n7379 ;
  assign n11083 = n11082 ^ n9875 ^ 1'b0 ;
  assign n11087 = n11086 ^ n11083 ^ n836 ;
  assign n11091 = n3249 ^ n2720 ^ n1707 ;
  assign n11088 = ( n1346 & n1775 ) | ( n1346 & ~n5607 ) | ( n1775 & ~n5607 ) ;
  assign n11089 = n8477 & n9729 ;
  assign n11090 = ~n11088 & n11089 ;
  assign n11092 = n11091 ^ n11090 ^ n6127 ;
  assign n11093 = n1285 & n3816 ;
  assign n11094 = n10110 & n11093 ;
  assign n11095 = n2519 & ~n11094 ;
  assign n11098 = n5058 | n6441 ;
  assign n11099 = n879 | n11098 ;
  assign n11100 = ~n8224 & n11099 ;
  assign n11101 = n11100 ^ n4678 ^ 1'b0 ;
  assign n11096 = n5756 & n7963 ;
  assign n11097 = ( n2100 & n10871 ) | ( n2100 & n11096 ) | ( n10871 & n11096 ) ;
  assign n11102 = n11101 ^ n11097 ^ n6469 ;
  assign n11103 = ~n1517 & n6418 ;
  assign n11104 = n590 & n11103 ;
  assign n11105 = n2560 & ~n11104 ;
  assign n11106 = n2157 & n11105 ;
  assign n11107 = n3035 ^ n1153 ^ 1'b0 ;
  assign n11108 = n5637 | n10523 ;
  assign n11109 = n5366 ^ n4351 ^ 1'b0 ;
  assign n11110 = n1436 | n7970 ;
  assign n11111 = n1915 & ~n2046 ;
  assign n11112 = n11111 ^ n215 ^ 1'b0 ;
  assign n11113 = n9535 | n10750 ;
  assign n11114 = n11112 & ~n11113 ;
  assign n11115 = ~n1526 & n9906 ;
  assign n11117 = n1839 & ~n11074 ;
  assign n11118 = n6353 & n11117 ;
  assign n11116 = n7602 ^ n4268 ^ n161 ;
  assign n11119 = n11118 ^ n11116 ^ 1'b0 ;
  assign n11120 = n11119 ^ n5708 ^ n2061 ;
  assign n11121 = ~n2714 & n2895 ;
  assign n11122 = n11121 ^ n6824 ^ 1'b0 ;
  assign n11123 = n11122 ^ n5556 ^ n2000 ;
  assign n11124 = ~n5705 & n11123 ;
  assign n11125 = n5112 ^ n2661 ^ n1007 ;
  assign n11126 = n7309 ^ n6733 ^ 1'b0 ;
  assign n11127 = n11125 | n11126 ;
  assign n11128 = n3438 ^ n1778 ^ n1738 ;
  assign n11129 = n11128 ^ n1507 ^ 1'b0 ;
  assign n11130 = n8585 ^ n4500 ^ n4431 ;
  assign n11131 = n7770 & n11130 ;
  assign n11132 = ~n828 & n1208 ;
  assign n11133 = n1290 & n11132 ;
  assign n11134 = ( n5285 & ~n10998 ) | ( n5285 & n11133 ) | ( ~n10998 & n11133 ) ;
  assign n11135 = n6991 ^ n4224 ^ 1'b0 ;
  assign n11136 = n11135 ^ n6181 ^ n1348 ;
  assign n11137 = n5177 ^ n4960 ^ n3020 ;
  assign n11138 = n11137 ^ n1456 ^ 1'b0 ;
  assign n11139 = n10260 ^ n7759 ^ 1'b0 ;
  assign n11140 = n8745 ^ n7361 ^ n1272 ;
  assign n11141 = ( n3272 & n7752 ) | ( n3272 & ~n11140 ) | ( n7752 & ~n11140 ) ;
  assign n11142 = ( n1088 & n2900 ) | ( n1088 & ~n11141 ) | ( n2900 & ~n11141 ) ;
  assign n11143 = ( n1796 & n7518 ) | ( n1796 & n9399 ) | ( n7518 & n9399 ) ;
  assign n11144 = ( n643 & n2960 ) | ( n643 & ~n11143 ) | ( n2960 & ~n11143 ) ;
  assign n11145 = n8282 | n11144 ;
  assign n11146 = n7930 | n11145 ;
  assign n11147 = n10172 ^ n9351 ^ 1'b0 ;
  assign n11148 = n8128 & n11147 ;
  assign n11149 = n7302 ^ n2207 ^ n1612 ;
  assign n11150 = ~n1212 & n11149 ;
  assign n11151 = n2155 & ~n4164 ;
  assign n11152 = ( n2237 & ~n10686 ) | ( n2237 & n11151 ) | ( ~n10686 & n11151 ) ;
  assign n11153 = ~n657 & n3934 ;
  assign n11154 = ~n7240 & n11153 ;
  assign n11159 = n3650 & ~n5843 ;
  assign n11160 = n11159 ^ n5710 ^ 1'b0 ;
  assign n11161 = n11160 ^ n5516 ^ 1'b0 ;
  assign n11155 = n8262 ^ n3452 ^ n1719 ;
  assign n11156 = n11155 ^ n6945 ^ n6786 ;
  assign n11157 = n3975 | n11156 ;
  assign n11158 = n11157 ^ n8324 ^ 1'b0 ;
  assign n11162 = n11161 ^ n11158 ^ n10323 ;
  assign n11166 = n645 & n6742 ;
  assign n11167 = n11166 ^ n5619 ^ 1'b0 ;
  assign n11163 = n3636 & ~n4324 ;
  assign n11164 = n11163 ^ n9664 ^ 1'b0 ;
  assign n11165 = n11164 ^ n2754 ^ 1'b0 ;
  assign n11168 = n11167 ^ n11165 ^ n7572 ;
  assign n11169 = n1955 | n4663 ;
  assign n11170 = n11169 ^ n6543 ^ 1'b0 ;
  assign n11171 = n6253 ^ n6207 ^ n6042 ;
  assign n11172 = ( n5331 & n6648 ) | ( n5331 & n11171 ) | ( n6648 & n11171 ) ;
  assign n11173 = ~n4049 & n11172 ;
  assign n11174 = n9524 | n11011 ;
  assign n11175 = n3899 | n11174 ;
  assign n11176 = n10877 ^ n9291 ^ n2438 ;
  assign n11177 = ( n900 & ~n6406 ) | ( n900 & n7815 ) | ( ~n6406 & n7815 ) ;
  assign n11178 = n2819 & n11177 ;
  assign n11179 = n9579 & n11178 ;
  assign n11180 = n11179 ^ n4501 ^ n3886 ;
  assign n11181 = ~n5701 & n7776 ;
  assign n11182 = ( ~n990 & n1871 ) | ( ~n990 & n2053 ) | ( n1871 & n2053 ) ;
  assign n11183 = ( n2922 & ~n6461 ) | ( n2922 & n11182 ) | ( ~n6461 & n11182 ) ;
  assign n11184 = n11183 ^ n10934 ^ n3115 ;
  assign n11185 = ( ~n8870 & n8910 ) | ( ~n8870 & n11184 ) | ( n8910 & n11184 ) ;
  assign n11186 = n4748 ^ n4005 ^ 1'b0 ;
  assign n11187 = n11185 & n11186 ;
  assign n11188 = ~n136 & n575 ;
  assign n11189 = n11188 ^ n762 ^ 1'b0 ;
  assign n11190 = n11189 ^ n5829 ^ 1'b0 ;
  assign n11191 = n3577 & ~n11190 ;
  assign n11192 = n814 & n6377 ;
  assign n11193 = n11192 ^ n4183 ^ 1'b0 ;
  assign n11194 = ( x48 & n6300 ) | ( x48 & n11193 ) | ( n6300 & n11193 ) ;
  assign n11195 = n8876 ^ n5122 ^ 1'b0 ;
  assign n11196 = n11195 ^ n9327 ^ n2058 ;
  assign n11197 = n11115 ^ n10165 ^ 1'b0 ;
  assign n11198 = ~n7185 & n10006 ;
  assign n11199 = ( n6202 & ~n9078 ) | ( n6202 & n11198 ) | ( ~n9078 & n11198 ) ;
  assign n11200 = n2666 ^ n2549 ^ n825 ;
  assign n11201 = n4767 & n11200 ;
  assign n11202 = n11201 ^ n8470 ^ n468 ;
  assign n11203 = ( ~n1117 & n2595 ) | ( ~n1117 & n9119 ) | ( n2595 & n9119 ) ;
  assign n11204 = ( n700 & n3647 ) | ( n700 & ~n11203 ) | ( n3647 & ~n11203 ) ;
  assign n11205 = x80 & ~n11204 ;
  assign n11206 = n11202 & n11205 ;
  assign n11207 = n166 & n4353 ;
  assign n11208 = n11207 ^ n5033 ^ 1'b0 ;
  assign n11209 = ( n3955 & n4004 ) | ( n3955 & n8656 ) | ( n4004 & n8656 ) ;
  assign n11213 = ( n1566 & n1953 ) | ( n1566 & n2448 ) | ( n1953 & n2448 ) ;
  assign n11214 = x101 & n8201 ;
  assign n11215 = ~n11213 & n11214 ;
  assign n11210 = n8370 | n9414 ;
  assign n11211 = n11210 ^ n1044 ^ 1'b0 ;
  assign n11212 = n11211 ^ n10811 ^ n3265 ;
  assign n11216 = n11215 ^ n11212 ^ n9518 ;
  assign n11217 = n5152 ^ n4793 ^ 1'b0 ;
  assign n11218 = ~n3105 & n11217 ;
  assign n11219 = ( ~n867 & n2124 ) | ( ~n867 & n11218 ) | ( n2124 & n11218 ) ;
  assign n11220 = n7468 ^ n531 ^ 1'b0 ;
  assign n11221 = n4596 & ~n11220 ;
  assign n11222 = n4925 ^ n3987 ^ n1844 ;
  assign n11223 = ( n3103 & ~n3836 ) | ( n3103 & n11222 ) | ( ~n3836 & n11222 ) ;
  assign n11224 = n11223 ^ n2431 ^ n1255 ;
  assign n11225 = ( n885 & ~n11221 ) | ( n885 & n11224 ) | ( ~n11221 & n11224 ) ;
  assign n11226 = n2871 & n11225 ;
  assign n11227 = n8375 & n11226 ;
  assign n11228 = n11227 ^ n1602 ^ 1'b0 ;
  assign n11229 = ~n3107 & n11228 ;
  assign n11230 = n6832 ^ n6452 ^ 1'b0 ;
  assign n11231 = n11230 ^ n8971 ^ 1'b0 ;
  assign n11232 = ~n9974 & n11231 ;
  assign n11233 = n10845 ^ n8239 ^ n2167 ;
  assign n11234 = n11233 ^ n9630 ^ n5441 ;
  assign n11235 = n11234 ^ n4770 ^ 1'b0 ;
  assign n11236 = ( n5288 & n5675 ) | ( n5288 & ~n11235 ) | ( n5675 & ~n11235 ) ;
  assign n11237 = ( ~n808 & n2410 ) | ( ~n808 & n5329 ) | ( n2410 & n5329 ) ;
  assign n11243 = n646 | n3007 ;
  assign n11244 = n11243 ^ n3334 ^ 1'b0 ;
  assign n11245 = ( ~n1228 & n5622 ) | ( ~n1228 & n11244 ) | ( n5622 & n11244 ) ;
  assign n11238 = n6746 ^ n1062 ^ 1'b0 ;
  assign n11239 = n1513 | n11238 ;
  assign n11240 = n11239 ^ x7 ^ 1'b0 ;
  assign n11241 = n5592 ^ n4748 ^ 1'b0 ;
  assign n11242 = n11240 | n11241 ;
  assign n11246 = n11245 ^ n11242 ^ 1'b0 ;
  assign n11247 = ( n2864 & ~n10505 ) | ( n2864 & n11246 ) | ( ~n10505 & n11246 ) ;
  assign n11248 = ( ~n3605 & n11237 ) | ( ~n3605 & n11247 ) | ( n11237 & n11247 ) ;
  assign n11249 = n6885 ^ n3798 ^ n995 ;
  assign n11250 = n11249 ^ n8583 ^ 1'b0 ;
  assign n11251 = ~n3565 & n11250 ;
  assign n11252 = ~n7108 & n11251 ;
  assign n11253 = n10555 & n11252 ;
  assign n11254 = n5033 | n7644 ;
  assign n11255 = n11254 ^ n7508 ^ 1'b0 ;
  assign n11257 = n421 & n2210 ;
  assign n11258 = n5773 & n11257 ;
  assign n11259 = n6794 | n11258 ;
  assign n11260 = n11259 ^ n1614 ^ 1'b0 ;
  assign n11256 = ~n1977 & n9801 ;
  assign n11261 = n11260 ^ n11256 ^ n9052 ;
  assign n11262 = ( n1913 & ~n4385 ) | ( n1913 & n5146 ) | ( ~n4385 & n5146 ) ;
  assign n11266 = n4989 ^ n1592 ^ n206 ;
  assign n11263 = n3071 & n4315 ;
  assign n11264 = ~n3513 & n11263 ;
  assign n11265 = n11264 ^ n4975 ^ 1'b0 ;
  assign n11267 = n11266 ^ n11265 ^ n1833 ;
  assign n11268 = ( ~n2521 & n2556 ) | ( ~n2521 & n3823 ) | ( n2556 & n3823 ) ;
  assign n11269 = ( n2898 & n4325 ) | ( n2898 & ~n11268 ) | ( n4325 & ~n11268 ) ;
  assign n11270 = n11269 ^ x80 ^ 1'b0 ;
  assign n11271 = ~n10970 & n11270 ;
  assign n11272 = n9923 ^ n9682 ^ n310 ;
  assign n11273 = n7571 | n11272 ;
  assign n11274 = n11273 ^ n6683 ^ 1'b0 ;
  assign n11275 = n6094 ^ n2484 ^ 1'b0 ;
  assign n11276 = ( n1929 & ~n3779 ) | ( n1929 & n11275 ) | ( ~n3779 & n11275 ) ;
  assign n11277 = n11276 ^ n7129 ^ n2045 ;
  assign n11278 = n3785 ^ n3671 ^ n656 ;
  assign n11279 = ~n7311 & n11278 ;
  assign n11280 = n11277 & n11279 ;
  assign n11281 = n7490 ^ n2967 ^ n2917 ;
  assign n11282 = ~n2392 & n11281 ;
  assign n11283 = ~n2112 & n11282 ;
  assign n11284 = ~n7402 & n7917 ;
  assign n11288 = n1133 & ~n3436 ;
  assign n11289 = n11288 ^ n1269 ^ 1'b0 ;
  assign n11290 = ( ~n1217 & n3334 ) | ( ~n1217 & n11289 ) | ( n3334 & n11289 ) ;
  assign n11285 = n4030 & ~n10021 ;
  assign n11286 = n11285 ^ n2435 ^ 1'b0 ;
  assign n11287 = n11286 ^ n5811 ^ 1'b0 ;
  assign n11291 = n11290 ^ n11287 ^ n3386 ;
  assign n11292 = ( n653 & ~n11284 ) | ( n653 & n11291 ) | ( ~n11284 & n11291 ) ;
  assign n11293 = n7472 ^ n1524 ^ 1'b0 ;
  assign n11294 = n2882 ^ n672 ^ n616 ;
  assign n11295 = n6195 & ~n11294 ;
  assign n11296 = ( n726 & n1691 ) | ( n726 & ~n11295 ) | ( n1691 & ~n11295 ) ;
  assign n11297 = n11296 ^ n8754 ^ n4509 ;
  assign n11298 = n5700 ^ n4754 ^ n3092 ;
  assign n11299 = n11298 ^ n4188 ^ n3146 ;
  assign n11300 = ( n7142 & ~n9008 ) | ( n7142 & n9774 ) | ( ~n9008 & n9774 ) ;
  assign n11301 = n11300 ^ n10194 ^ 1'b0 ;
  assign n11302 = n5879 | n11301 ;
  assign n11303 = n6612 ^ n3868 ^ 1'b0 ;
  assign n11304 = n4157 & ~n11303 ;
  assign n11305 = n11304 ^ n5233 ^ 1'b0 ;
  assign n11306 = n11305 ^ n1154 ^ n342 ;
  assign n11307 = n4553 & n10912 ;
  assign n11308 = n8241 ^ n1619 ^ 1'b0 ;
  assign n11309 = n337 & n620 ;
  assign n11310 = n11309 ^ n1297 ^ 1'b0 ;
  assign n11311 = n11310 ^ n5969 ^ 1'b0 ;
  assign n11312 = ~n4795 & n11311 ;
  assign n11313 = ( ~n6820 & n10313 ) | ( ~n6820 & n11312 ) | ( n10313 & n11312 ) ;
  assign n11314 = n2897 ^ n2529 ^ 1'b0 ;
  assign n11315 = n6104 & ~n11314 ;
  assign n11316 = ( ~n1996 & n4275 ) | ( ~n1996 & n11315 ) | ( n4275 & n11315 ) ;
  assign n11317 = n11316 ^ n6700 ^ 1'b0 ;
  assign n11318 = n11317 ^ n1065 ^ 1'b0 ;
  assign n11324 = n317 & ~n6112 ;
  assign n11325 = ~n6775 & n11324 ;
  assign n11319 = n3759 ^ n2327 ^ 1'b0 ;
  assign n11320 = n9577 ^ n2206 ^ 1'b0 ;
  assign n11321 = n5106 | n11320 ;
  assign n11322 = n11319 | n11321 ;
  assign n11323 = n1260 | n11322 ;
  assign n11326 = n11325 ^ n11323 ^ n6580 ;
  assign n11327 = n7615 & ~n11326 ;
  assign n11328 = ~n3184 & n11327 ;
  assign n11329 = n8516 ^ n6635 ^ n526 ;
  assign n11330 = n11329 ^ n2463 ^ 1'b0 ;
  assign n11331 = n6972 ^ n3928 ^ 1'b0 ;
  assign n11332 = ( ~n8100 & n11330 ) | ( ~n8100 & n11331 ) | ( n11330 & n11331 ) ;
  assign n11333 = n11332 ^ n9356 ^ 1'b0 ;
  assign n11334 = ~n3936 & n6667 ;
  assign n11335 = ~n5829 & n11334 ;
  assign n11336 = n11335 ^ n5987 ^ 1'b0 ;
  assign n11337 = n6938 ^ n2152 ^ n949 ;
  assign n11338 = n8774 ^ n1633 ^ 1'b0 ;
  assign n11339 = ~n11337 & n11338 ;
  assign n11340 = ( n348 & n1118 ) | ( n348 & ~n3965 ) | ( n1118 & ~n3965 ) ;
  assign n11341 = n11340 ^ n5949 ^ 1'b0 ;
  assign n11342 = ~n866 & n11341 ;
  assign n11345 = x106 & n2113 ;
  assign n11343 = n3217 ^ x2 ^ 1'b0 ;
  assign n11344 = n11343 ^ n8833 ^ 1'b0 ;
  assign n11346 = n11345 ^ n11344 ^ 1'b0 ;
  assign n11347 = n11346 ^ n4803 ^ n819 ;
  assign n11348 = n8707 ^ n2395 ^ 1'b0 ;
  assign n11349 = n7403 & ~n11348 ;
  assign n11350 = ( ~n664 & n2974 ) | ( ~n664 & n4737 ) | ( n2974 & n4737 ) ;
  assign n11351 = n1199 ^ n385 ^ 1'b0 ;
  assign n11352 = ~n7017 & n11351 ;
  assign n11353 = ( ~n754 & n11350 ) | ( ~n754 & n11352 ) | ( n11350 & n11352 ) ;
  assign n11354 = n10697 ^ n2443 ^ 1'b0 ;
  assign n11355 = n10686 & ~n11354 ;
  assign n11356 = ( n4827 & n5120 ) | ( n4827 & ~n11355 ) | ( n5120 & ~n11355 ) ;
  assign n11357 = n7435 ^ n1107 ^ 1'b0 ;
  assign n11358 = ~n4974 & n11357 ;
  assign n11359 = n11358 ^ n3874 ^ n3509 ;
  assign n11360 = n2833 & n11359 ;
  assign n11361 = ~n10198 & n11360 ;
  assign n11363 = n1709 | n7318 ;
  assign n11362 = n3501 & ~n11319 ;
  assign n11364 = n11363 ^ n11362 ^ 1'b0 ;
  assign n11365 = n2272 ^ n176 ^ 1'b0 ;
  assign n11366 = n1827 & n11365 ;
  assign n11367 = n11366 ^ n5923 ^ n5255 ;
  assign n11368 = n6617 ^ n4105 ^ 1'b0 ;
  assign n11374 = n672 & n4543 ;
  assign n11369 = n8145 ^ n3345 ^ 1'b0 ;
  assign n11370 = ~n3791 & n11369 ;
  assign n11371 = ~n4002 & n11370 ;
  assign n11372 = n11371 ^ n6490 ^ 1'b0 ;
  assign n11373 = n11372 ^ n2209 ^ 1'b0 ;
  assign n11375 = n11374 ^ n11373 ^ n2603 ;
  assign n11376 = n11375 ^ n5121 ^ 1'b0 ;
  assign n11377 = ( ~x37 & x43 ) | ( ~x37 & n9761 ) | ( x43 & n9761 ) ;
  assign n11378 = n3712 ^ n3107 ^ n1244 ;
  assign n11379 = n4440 ^ n4365 ^ n142 ;
  assign n11380 = n11379 ^ n5757 ^ n5551 ;
  assign n11381 = ( ~n652 & n2834 ) | ( ~n652 & n11380 ) | ( n2834 & n11380 ) ;
  assign n11382 = ( ~n300 & n4869 ) | ( ~n300 & n9358 ) | ( n4869 & n9358 ) ;
  assign n11383 = ( ~n7759 & n11381 ) | ( ~n7759 & n11382 ) | ( n11381 & n11382 ) ;
  assign n11384 = ~n3193 & n11383 ;
  assign n11385 = n11378 & n11384 ;
  assign n11386 = n9795 ^ n8017 ^ n7142 ;
  assign n11387 = n11386 ^ n7727 ^ n7358 ;
  assign n11388 = n5027 & ~n5575 ;
  assign n11389 = ~n2056 & n11388 ;
  assign n11390 = n2687 | n5385 ;
  assign n11391 = n11390 ^ n5373 ^ 1'b0 ;
  assign n11392 = ( n11387 & n11389 ) | ( n11387 & ~n11391 ) | ( n11389 & ~n11391 ) ;
  assign n11393 = n1977 ^ n880 ^ 1'b0 ;
  assign n11394 = n11393 ^ n4198 ^ 1'b0 ;
  assign n11395 = ( n4567 & n5497 ) | ( n4567 & ~n11394 ) | ( n5497 & ~n11394 ) ;
  assign n11396 = n11395 ^ n6659 ^ n3990 ;
  assign n11397 = n11396 ^ n5665 ^ n2081 ;
  assign n11398 = n11022 ^ n6053 ^ 1'b0 ;
  assign n11399 = n11398 ^ n4816 ^ 1'b0 ;
  assign n11406 = n7307 ^ n6001 ^ n2905 ;
  assign n11407 = ~n133 & n11406 ;
  assign n11408 = n4612 & n11407 ;
  assign n11409 = ~n7305 & n11408 ;
  assign n11400 = n3325 ^ n2428 ^ n1935 ;
  assign n11401 = n11400 ^ n5234 ^ 1'b0 ;
  assign n11402 = n11401 ^ n7001 ^ n631 ;
  assign n11403 = ~n7386 & n11402 ;
  assign n11404 = n3877 & ~n8566 ;
  assign n11405 = n11403 & n11404 ;
  assign n11410 = n11409 ^ n11405 ^ 1'b0 ;
  assign n11411 = ( ~n1761 & n3442 ) | ( ~n1761 & n9141 ) | ( n3442 & n9141 ) ;
  assign n11412 = n6630 ^ n4023 ^ n648 ;
  assign n11413 = ( ~n11076 & n11411 ) | ( ~n11076 & n11412 ) | ( n11411 & n11412 ) ;
  assign n11415 = ( n3593 & n5133 ) | ( n3593 & n11303 ) | ( n5133 & n11303 ) ;
  assign n11414 = n1899 | n7096 ;
  assign n11416 = n11415 ^ n11414 ^ n365 ;
  assign n11418 = ( n2835 & n3201 ) | ( n2835 & n7585 ) | ( n3201 & n7585 ) ;
  assign n11419 = n11418 ^ n3436 ^ 1'b0 ;
  assign n11420 = n3424 & n7116 ;
  assign n11421 = n11419 & n11420 ;
  assign n11417 = ( ~n888 & n9069 ) | ( ~n888 & n9131 ) | ( n9069 & n9131 ) ;
  assign n11422 = n11421 ^ n11417 ^ 1'b0 ;
  assign n11423 = n3468 ^ n2828 ^ n1717 ;
  assign n11424 = ( n10774 & n11422 ) | ( n10774 & ~n11423 ) | ( n11422 & ~n11423 ) ;
  assign n11425 = n8450 ^ n4572 ^ n2418 ;
  assign n11426 = n9422 ^ n8008 ^ n6123 ;
  assign n11427 = n11426 ^ n2946 ^ 1'b0 ;
  assign n11432 = n8816 ^ x122 ^ 1'b0 ;
  assign n11431 = n4477 ^ n3556 ^ n1255 ;
  assign n11433 = n11432 ^ n11431 ^ n5487 ;
  assign n11429 = ( n1510 & n3919 ) | ( n1510 & n10469 ) | ( n3919 & n10469 ) ;
  assign n11428 = n1665 | n3906 ;
  assign n11430 = n11429 ^ n11428 ^ 1'b0 ;
  assign n11434 = n11433 ^ n11430 ^ 1'b0 ;
  assign n11435 = ( n2424 & n3166 ) | ( n2424 & ~n9448 ) | ( n3166 & ~n9448 ) ;
  assign n11436 = n11435 ^ n6454 ^ 1'b0 ;
  assign n11437 = n11436 ^ n11249 ^ 1'b0 ;
  assign n11438 = n11052 & n11437 ;
  assign n11439 = ( ~n2245 & n5802 ) | ( ~n2245 & n6650 ) | ( n5802 & n6650 ) ;
  assign n11440 = n2623 | n6022 ;
  assign n11441 = n4766 ^ n4378 ^ n3169 ;
  assign n11442 = n11441 ^ n6627 ^ n4383 ;
  assign n11443 = ( n10666 & ~n11440 ) | ( n10666 & n11442 ) | ( ~n11440 & n11442 ) ;
  assign n11444 = ( n724 & ~n2844 ) | ( n724 & n11443 ) | ( ~n2844 & n11443 ) ;
  assign n11445 = n11108 ^ n1425 ^ 1'b0 ;
  assign n11446 = n9629 & ~n11445 ;
  assign n11447 = n6420 & n7890 ;
  assign n11453 = n6068 ^ n2541 ^ n490 ;
  assign n11448 = ~n1468 & n8008 ;
  assign n11449 = ~n7765 & n11448 ;
  assign n11450 = n11449 ^ n5664 ^ n3202 ;
  assign n11451 = ~n1533 & n11450 ;
  assign n11452 = n11451 ^ n609 ^ 1'b0 ;
  assign n11454 = n11453 ^ n11452 ^ 1'b0 ;
  assign n11455 = ( n8517 & n11447 ) | ( n8517 & ~n11454 ) | ( n11447 & ~n11454 ) ;
  assign n11456 = ~x87 & n10176 ;
  assign n11457 = n11456 ^ n7440 ^ n6095 ;
  assign n11458 = ( n6999 & n8992 ) | ( n6999 & ~n9411 ) | ( n8992 & ~n9411 ) ;
  assign n11459 = n1532 ^ n1359 ^ 1'b0 ;
  assign n11460 = n4289 & n11459 ;
  assign n11461 = n11460 ^ n9155 ^ n7008 ;
  assign n11462 = n4369 | n11461 ;
  assign n11463 = n11462 ^ n9631 ^ 1'b0 ;
  assign n11464 = n3814 ^ n2544 ^ 1'b0 ;
  assign n11465 = ~n1003 & n11464 ;
  assign n11466 = n11465 ^ n8584 ^ 1'b0 ;
  assign n11472 = ( ~n3996 & n6805 ) | ( ~n3996 & n8507 ) | ( n6805 & n8507 ) ;
  assign n11467 = ( n2612 & n5559 ) | ( n2612 & n6380 ) | ( n5559 & n6380 ) ;
  assign n11468 = n1592 ^ n699 ^ n229 ;
  assign n11469 = n11468 ^ n10873 ^ n524 ;
  assign n11470 = ~n3795 & n11469 ;
  assign n11471 = ~n11467 & n11470 ;
  assign n11473 = n11472 ^ n11471 ^ n1454 ;
  assign n11474 = n442 & ~n6267 ;
  assign n11475 = ( n1470 & n5490 ) | ( n1470 & n7792 ) | ( n5490 & n7792 ) ;
  assign n11476 = n2061 & n7606 ;
  assign n11477 = n11475 & n11476 ;
  assign n11478 = n1314 & n1561 ;
  assign n11479 = n11478 ^ n6198 ^ 1'b0 ;
  assign n11480 = ( n1936 & ~n3847 ) | ( n1936 & n11479 ) | ( ~n3847 & n11479 ) ;
  assign n11481 = n11480 ^ n383 ^ 1'b0 ;
  assign n11482 = n4132 & n11481 ;
  assign n11483 = n11482 ^ n10677 ^ n6435 ;
  assign n11484 = n794 | n8732 ;
  assign n11485 = n6709 & ~n11484 ;
  assign n11486 = n231 & n4448 ;
  assign n11487 = n3044 & n4810 ;
  assign n11488 = ( ~n4608 & n8151 ) | ( ~n4608 & n11487 ) | ( n8151 & n11487 ) ;
  assign n11489 = n11488 ^ n8316 ^ n3309 ;
  assign n11490 = n4363 ^ n1273 ^ 1'b0 ;
  assign n11491 = ~n6887 & n11490 ;
  assign n11492 = ~n9014 & n11491 ;
  assign n11493 = n7416 & n11492 ;
  assign n11497 = ( ~n3676 & n4620 ) | ( ~n3676 & n6297 ) | ( n4620 & n6297 ) ;
  assign n11495 = ( n659 & n2289 ) | ( n659 & n6628 ) | ( n2289 & n6628 ) ;
  assign n11496 = n11495 ^ n9349 ^ 1'b0 ;
  assign n11494 = n10061 ^ n7667 ^ n249 ;
  assign n11498 = n11497 ^ n11496 ^ n11494 ;
  assign n11499 = ~n2151 & n2828 ;
  assign n11500 = n11499 ^ n724 ^ 1'b0 ;
  assign n11501 = n2020 & ~n11500 ;
  assign n11502 = ( n1034 & n9306 ) | ( n1034 & ~n11501 ) | ( n9306 & ~n11501 ) ;
  assign n11503 = n563 & ~n11502 ;
  assign n11504 = ( ~n3372 & n3609 ) | ( ~n3372 & n9659 ) | ( n3609 & n9659 ) ;
  assign n11505 = n11504 ^ n8831 ^ n1566 ;
  assign n11512 = ~n1117 & n2086 ;
  assign n11509 = n2724 | n9118 ;
  assign n11510 = n11509 ^ n4189 ^ 1'b0 ;
  assign n11511 = n5514 & ~n11510 ;
  assign n11506 = n5413 ^ n3996 ^ n2132 ;
  assign n11507 = n11506 ^ n9588 ^ 1'b0 ;
  assign n11508 = ( n4452 & n8631 ) | ( n4452 & ~n11507 ) | ( n8631 & ~n11507 ) ;
  assign n11513 = n11512 ^ n11511 ^ n11508 ;
  assign n11514 = n5088 ^ n3995 ^ n901 ;
  assign n11515 = n8262 ^ n7651 ^ n338 ;
  assign n11516 = n765 | n11515 ;
  assign n11517 = n11516 ^ n1957 ^ 1'b0 ;
  assign n11518 = n4452 | n11517 ;
  assign n11519 = n5390 & ~n11518 ;
  assign n11526 = n3058 ^ n850 ^ x118 ;
  assign n11523 = n9176 | n10819 ;
  assign n11521 = n4414 ^ n569 ^ 1'b0 ;
  assign n11522 = n1209 | n11521 ;
  assign n11520 = n1977 ^ n584 ^ 1'b0 ;
  assign n11524 = n11523 ^ n11522 ^ n11520 ;
  assign n11525 = ~n5693 & n11524 ;
  assign n11527 = n11526 ^ n11525 ^ 1'b0 ;
  assign n11528 = n9322 ^ n1834 ^ 1'b0 ;
  assign n11529 = n11528 ^ n10750 ^ 1'b0 ;
  assign n11530 = n1159 & ~n11529 ;
  assign n11531 = n11527 | n11530 ;
  assign n11532 = ~n8921 & n11531 ;
  assign n11533 = n11519 & n11532 ;
  assign n11534 = ( n3628 & ~n6741 ) | ( n3628 & n8126 ) | ( ~n6741 & n8126 ) ;
  assign n11535 = n9925 ^ n7013 ^ 1'b0 ;
  assign n11536 = ~n6363 & n11535 ;
  assign n11537 = n11534 | n11536 ;
  assign n11538 = ( n3513 & ~n4183 ) | ( n3513 & n4793 ) | ( ~n4183 & n4793 ) ;
  assign n11539 = ( n4554 & ~n9708 ) | ( n4554 & n9994 ) | ( ~n9708 & n9994 ) ;
  assign n11540 = ~x56 & n324 ;
  assign n11541 = n1759 ^ n559 ^ n529 ;
  assign n11542 = n11541 ^ n3602 ^ 1'b0 ;
  assign n11543 = n7954 & n11542 ;
  assign n11544 = ( n3695 & n3962 ) | ( n3695 & ~n11543 ) | ( n3962 & ~n11543 ) ;
  assign n11545 = ( n3634 & n7667 ) | ( n3634 & n11544 ) | ( n7667 & n11544 ) ;
  assign n11546 = ( n6799 & n7781 ) | ( n6799 & n11545 ) | ( n7781 & n11545 ) ;
  assign n11547 = ( n7107 & ~n11540 ) | ( n7107 & n11546 ) | ( ~n11540 & n11546 ) ;
  assign n11548 = ( n3368 & n11539 ) | ( n3368 & n11547 ) | ( n11539 & n11547 ) ;
  assign n11549 = ( n1636 & n8324 ) | ( n1636 & n11548 ) | ( n8324 & n11548 ) ;
  assign n11550 = ( n7598 & n11538 ) | ( n7598 & ~n11549 ) | ( n11538 & ~n11549 ) ;
  assign n11555 = n808 & n3442 ;
  assign n11551 = n532 & n1583 ;
  assign n11552 = n11551 ^ n10990 ^ n6916 ;
  assign n11553 = n7854 ^ n6035 ^ 1'b0 ;
  assign n11554 = n11552 & n11553 ;
  assign n11556 = n11555 ^ n11554 ^ 1'b0 ;
  assign n11557 = ( n1419 & ~n2584 ) | ( n1419 & n8235 ) | ( ~n2584 & n8235 ) ;
  assign n11558 = ( n5011 & n5461 ) | ( n5011 & n11557 ) | ( n5461 & n11557 ) ;
  assign n11564 = n6371 ^ n1243 ^ n426 ;
  assign n11563 = ( n3334 & ~n3936 ) | ( n3334 & n9366 ) | ( ~n3936 & n9366 ) ;
  assign n11559 = n2502 ^ n410 ^ 1'b0 ;
  assign n11560 = n1782 & ~n11559 ;
  assign n11561 = n600 | n5867 ;
  assign n11562 = n11560 | n11561 ;
  assign n11565 = n11564 ^ n11563 ^ n11562 ;
  assign n11566 = ( n5142 & ~n7712 ) | ( n5142 & n11565 ) | ( ~n7712 & n11565 ) ;
  assign n11567 = n11566 ^ n697 ^ 1'b0 ;
  assign n11568 = n1490 & n11567 ;
  assign n11569 = ( n492 & n1163 ) | ( n492 & ~n5175 ) | ( n1163 & ~n5175 ) ;
  assign n11570 = ( n5556 & n6418 ) | ( n5556 & ~n11569 ) | ( n6418 & ~n11569 ) ;
  assign n11571 = n9853 ^ n9573 ^ 1'b0 ;
  assign n11572 = n11570 | n11571 ;
  assign n11573 = ~n4065 & n9102 ;
  assign n11574 = n11573 ^ n8284 ^ 1'b0 ;
  assign n11578 = n2718 ^ n2611 ^ 1'b0 ;
  assign n11579 = n5491 & n11578 ;
  assign n11580 = n7640 ^ n2273 ^ 1'b0 ;
  assign n11581 = n11579 & ~n11580 ;
  assign n11575 = x30 & n2603 ;
  assign n11576 = ~n3075 & n11575 ;
  assign n11577 = n9753 & ~n11576 ;
  assign n11582 = n11581 ^ n11577 ^ 1'b0 ;
  assign n11583 = ( n7977 & ~n11574 ) | ( n7977 & n11582 ) | ( ~n11574 & n11582 ) ;
  assign n11584 = n1146 & n2405 ;
  assign n11585 = n11584 ^ n1323 ^ 1'b0 ;
  assign n11586 = n11585 ^ n3935 ^ 1'b0 ;
  assign n11587 = ( n504 & n7766 ) | ( n504 & n11586 ) | ( n7766 & n11586 ) ;
  assign n11588 = n11587 ^ n508 ^ 1'b0 ;
  assign n11589 = n8486 | n9656 ;
  assign n11590 = n11588 & ~n11589 ;
  assign n11591 = n5512 ^ n1243 ^ n726 ;
  assign n11592 = n11591 ^ n5616 ^ n2930 ;
  assign n11593 = n11352 & ~n11592 ;
  assign n11604 = ( n1160 & n2507 ) | ( n1160 & ~n2870 ) | ( n2507 & ~n2870 ) ;
  assign n11594 = ( n1898 & n3785 ) | ( n1898 & ~n9711 ) | ( n3785 & ~n9711 ) ;
  assign n11595 = n4098 | n5648 ;
  assign n11596 = n7940 | n11595 ;
  assign n11597 = ( ~n9221 & n9397 ) | ( ~n9221 & n11596 ) | ( n9397 & n11596 ) ;
  assign n11598 = ( x114 & n5756 ) | ( x114 & n5863 ) | ( n5756 & n5863 ) ;
  assign n11599 = n2999 & n3779 ;
  assign n11600 = n6999 & n11599 ;
  assign n11601 = ( n518 & n11598 ) | ( n518 & ~n11600 ) | ( n11598 & ~n11600 ) ;
  assign n11602 = ( n7644 & n11597 ) | ( n7644 & ~n11601 ) | ( n11597 & ~n11601 ) ;
  assign n11603 = ( n6436 & n11594 ) | ( n6436 & ~n11602 ) | ( n11594 & ~n11602 ) ;
  assign n11605 = n11604 ^ n11603 ^ n2804 ;
  assign n11614 = n4187 ^ n1451 ^ 1'b0 ;
  assign n11606 = ( ~n2050 & n3971 ) | ( ~n2050 & n7265 ) | ( n3971 & n7265 ) ;
  assign n11607 = n1916 | n11606 ;
  assign n11608 = n2256 & ~n11607 ;
  assign n11609 = n11469 & ~n11608 ;
  assign n11611 = ( n225 & n2932 ) | ( n225 & ~n9267 ) | ( n2932 & ~n9267 ) ;
  assign n11610 = n3339 & n7919 ;
  assign n11612 = n11611 ^ n11610 ^ 1'b0 ;
  assign n11613 = n11609 & ~n11612 ;
  assign n11615 = n11614 ^ n11613 ^ 1'b0 ;
  assign n11616 = ( n3413 & n4989 ) | ( n3413 & ~n9057 ) | ( n4989 & ~n9057 ) ;
  assign n11617 = n11616 ^ n11500 ^ 1'b0 ;
  assign n11618 = n6441 | n11617 ;
  assign n11619 = ( n4562 & n5455 ) | ( n4562 & ~n11618 ) | ( n5455 & ~n11618 ) ;
  assign n11620 = ~n2742 & n6780 ;
  assign n11621 = n2968 & ~n5104 ;
  assign n11622 = n11621 ^ n1675 ^ 1'b0 ;
  assign n11623 = ~n11620 & n11622 ;
  assign n11624 = n5629 & n11623 ;
  assign n11625 = n2622 & ~n3445 ;
  assign n11626 = ~n3163 & n11625 ;
  assign n11627 = ( ~n6566 & n8707 ) | ( ~n6566 & n11626 ) | ( n8707 & n11626 ) ;
  assign n11628 = n2242 ^ n2217 ^ n1829 ;
  assign n11630 = ( n2494 & n7154 ) | ( n2494 & n8886 ) | ( n7154 & n8886 ) ;
  assign n11631 = n11630 ^ n5676 ^ 1'b0 ;
  assign n11632 = ~n5499 & n11631 ;
  assign n11633 = n11632 ^ n6477 ^ n3967 ;
  assign n11629 = n3016 ^ n2495 ^ 1'b0 ;
  assign n11634 = n11633 ^ n11629 ^ 1'b0 ;
  assign n11635 = ( ~n7130 & n11628 ) | ( ~n7130 & n11634 ) | ( n11628 & n11634 ) ;
  assign n11636 = n1714 & ~n2680 ;
  assign n11637 = ~n10143 & n11636 ;
  assign n11638 = n11637 ^ n7701 ^ 1'b0 ;
  assign n11641 = n523 & ~n5221 ;
  assign n11639 = n2295 & n6742 ;
  assign n11640 = n6789 & n11639 ;
  assign n11642 = n11641 ^ n11640 ^ 1'b0 ;
  assign n11643 = ( n5928 & n9115 ) | ( n5928 & ~n9283 ) | ( n9115 & ~n9283 ) ;
  assign n11644 = n11643 ^ n7907 ^ n2580 ;
  assign n11645 = n10605 ^ n834 ^ 1'b0 ;
  assign n11646 = n7940 ^ n4449 ^ n767 ;
  assign n11647 = n3291 & ~n8348 ;
  assign n11648 = n11647 ^ n2512 ^ 1'b0 ;
  assign n11649 = n3268 ^ n2667 ^ 1'b0 ;
  assign n11650 = n9532 & ~n11649 ;
  assign n11651 = ( n11646 & ~n11648 ) | ( n11646 & n11650 ) | ( ~n11648 & n11650 ) ;
  assign n11652 = ~n7300 & n11651 ;
  assign n11653 = n10650 ^ n5976 ^ 1'b0 ;
  assign n11654 = ( n1330 & ~n4084 ) | ( n1330 & n11653 ) | ( ~n4084 & n11653 ) ;
  assign n11655 = n11654 ^ n2661 ^ n575 ;
  assign n11658 = n4150 | n8644 ;
  assign n11659 = n1029 | n11658 ;
  assign n11660 = ( n1933 & n2317 ) | ( n1933 & n11659 ) | ( n2317 & n11659 ) ;
  assign n11657 = ( n2461 & n2585 ) | ( n2461 & ~n8372 ) | ( n2585 & ~n8372 ) ;
  assign n11661 = n11660 ^ n11657 ^ n5546 ;
  assign n11656 = n368 & n2590 ;
  assign n11662 = n11661 ^ n11656 ^ 1'b0 ;
  assign n11663 = n11662 ^ n9240 ^ n2433 ;
  assign n11664 = n10871 ^ n4540 ^ 1'b0 ;
  assign n11665 = ( n1835 & n3442 ) | ( n1835 & ~n5738 ) | ( n3442 & ~n5738 ) ;
  assign n11666 = n11665 ^ n10220 ^ n7020 ;
  assign n11667 = ( n3739 & n8145 ) | ( n3739 & ~n9469 ) | ( n8145 & ~n9469 ) ;
  assign n11668 = n2128 & ~n11667 ;
  assign n11669 = n11668 ^ n4634 ^ 1'b0 ;
  assign n11670 = ( n1664 & n9226 ) | ( n1664 & ~n10859 ) | ( n9226 & ~n10859 ) ;
  assign n11671 = n4712 | n8757 ;
  assign n11672 = n11670 & ~n11671 ;
  assign n11673 = n10762 ^ n5821 ^ n916 ;
  assign n11674 = n11673 ^ n11355 ^ n3288 ;
  assign n11681 = n5921 ^ n5694 ^ 1'b0 ;
  assign n11682 = n6540 | n11681 ;
  assign n11683 = ( n376 & ~n2312 ) | ( n376 & n11682 ) | ( ~n2312 & n11682 ) ;
  assign n11684 = n11683 ^ n4550 ^ 1'b0 ;
  assign n11685 = n2564 & ~n3541 ;
  assign n11686 = n765 & n11685 ;
  assign n11688 = n6450 & ~n8276 ;
  assign n11687 = n10505 ^ n3645 ^ n896 ;
  assign n11689 = n11688 ^ n11687 ^ 1'b0 ;
  assign n11690 = n11686 | n11689 ;
  assign n11691 = ~n11684 & n11690 ;
  assign n11675 = n3541 ^ n1895 ^ 1'b0 ;
  assign n11676 = ~n11616 & n11675 ;
  assign n11677 = ( n4632 & n8096 ) | ( n4632 & ~n11128 ) | ( n8096 & ~n11128 ) ;
  assign n11678 = n8700 ^ n7038 ^ 1'b0 ;
  assign n11679 = n11677 | n11678 ;
  assign n11680 = ( n9006 & n11676 ) | ( n9006 & n11679 ) | ( n11676 & n11679 ) ;
  assign n11692 = n11691 ^ n11680 ^ n5634 ;
  assign n11693 = ( ~x74 & n1565 ) | ( ~x74 & n5313 ) | ( n1565 & n5313 ) ;
  assign n11694 = n506 & ~n3792 ;
  assign n11695 = n11694 ^ n5153 ^ n434 ;
  assign n11696 = ( n5577 & n11693 ) | ( n5577 & ~n11695 ) | ( n11693 & ~n11695 ) ;
  assign n11697 = n11696 ^ n9691 ^ 1'b0 ;
  assign n11698 = n11692 & ~n11697 ;
  assign n11699 = n9207 ^ n7195 ^ n1493 ;
  assign n11700 = n11699 ^ n3014 ^ 1'b0 ;
  assign n11701 = ~n629 & n4953 ;
  assign n11702 = ( n582 & n2954 ) | ( n582 & ~n10682 ) | ( n2954 & ~n10682 ) ;
  assign n11703 = ( n5813 & n7467 ) | ( n5813 & ~n8583 ) | ( n7467 & ~n8583 ) ;
  assign n11704 = n10334 & ~n11703 ;
  assign n11705 = n6244 & n11704 ;
  assign n11706 = n2585 ^ x43 ^ 1'b0 ;
  assign n11707 = n10481 ^ n6877 ^ 1'b0 ;
  assign n11708 = n7901 | n11707 ;
  assign n11709 = n11708 ^ n8666 ^ 1'b0 ;
  assign n11710 = n10534 & n11709 ;
  assign n11714 = n11686 ^ n6293 ^ n4982 ;
  assign n11711 = n7307 ^ n702 ^ n150 ;
  assign n11712 = n7729 ^ n4670 ^ n1709 ;
  assign n11713 = ( n11585 & n11711 ) | ( n11585 & ~n11712 ) | ( n11711 & ~n11712 ) ;
  assign n11715 = n11714 ^ n11713 ^ 1'b0 ;
  assign n11716 = n5965 ^ n2592 ^ n189 ;
  assign n11717 = n5134 & ~n5554 ;
  assign n11718 = ~n2930 & n11717 ;
  assign n11719 = n11716 & ~n11718 ;
  assign n11720 = n11719 ^ n3756 ^ 1'b0 ;
  assign n11721 = ( n6508 & n11546 ) | ( n6508 & n11720 ) | ( n11546 & n11720 ) ;
  assign n11722 = ~n1862 & n8955 ;
  assign n11723 = n11722 ^ n8297 ^ n5663 ;
  assign n11724 = n6247 ^ n1666 ^ 1'b0 ;
  assign n11725 = n563 & ~n11724 ;
  assign n11726 = n11725 ^ n9500 ^ n3998 ;
  assign n11727 = n964 & ~n3558 ;
  assign n11728 = n8709 ^ n4861 ^ 1'b0 ;
  assign n11729 = ~n11727 & n11728 ;
  assign n11730 = n4975 ^ n3775 ^ n1018 ;
  assign n11731 = ( n1488 & ~n1594 ) | ( n1488 & n3260 ) | ( ~n1594 & n3260 ) ;
  assign n11732 = n8809 | n11731 ;
  assign n11733 = ~n980 & n11732 ;
  assign n11734 = n1327 | n11733 ;
  assign n11735 = n3706 | n6435 ;
  assign n11736 = n11735 ^ n2843 ^ 1'b0 ;
  assign n11737 = n11736 ^ n7583 ^ n2863 ;
  assign n11738 = n501 & n4279 ;
  assign n11739 = n9835 & ~n11660 ;
  assign n11740 = n11738 & n11739 ;
  assign n11741 = ( n1359 & n1508 ) | ( n1359 & ~n11740 ) | ( n1508 & ~n11740 ) ;
  assign n11742 = n6941 | n11741 ;
  assign n11743 = n11742 ^ n716 ^ 1'b0 ;
  assign n11744 = ~n11737 & n11743 ;
  assign n11745 = ( n10194 & n11003 ) | ( n10194 & n11440 ) | ( n11003 & n11440 ) ;
  assign n11746 = n6900 & n8486 ;
  assign n11747 = n2802 ^ n1843 ^ n1612 ;
  assign n11748 = n1804 & n5981 ;
  assign n11749 = n11748 ^ n1601 ^ 1'b0 ;
  assign n11750 = ( n1175 & ~n8103 ) | ( n1175 & n11749 ) | ( ~n8103 & n11749 ) ;
  assign n11751 = ~n11747 & n11750 ;
  assign n11752 = n11746 & n11751 ;
  assign n11753 = n1318 & ~n6029 ;
  assign n11754 = ~n2286 & n11753 ;
  assign n11755 = n7671 | n11754 ;
  assign n11756 = n2474 | n3678 ;
  assign n11757 = n1881 | n11756 ;
  assign n11758 = n11757 ^ n2157 ^ n698 ;
  assign n11759 = n11758 ^ n10963 ^ n1283 ;
  assign n11760 = ~n4784 & n10052 ;
  assign n11761 = n11760 ^ x84 ^ 1'b0 ;
  assign n11762 = n7676 ^ n1899 ^ n619 ;
  assign n11764 = n6013 ^ n4393 ^ 1'b0 ;
  assign n11763 = n2523 | n4350 ;
  assign n11765 = n11764 ^ n11763 ^ 1'b0 ;
  assign n11766 = n11765 ^ n3407 ^ 1'b0 ;
  assign n11767 = n11766 ^ n8276 ^ 1'b0 ;
  assign n11768 = n2993 & ~n11767 ;
  assign n11769 = n515 & ~n3969 ;
  assign n11770 = ~n9943 & n11769 ;
  assign n11771 = ( n2526 & ~n6223 ) | ( n2526 & n7107 ) | ( ~n6223 & n7107 ) ;
  assign n11772 = n4776 ^ n4500 ^ n1301 ;
  assign n11773 = n11772 ^ n4118 ^ 1'b0 ;
  assign n11774 = ( n926 & n9846 ) | ( n926 & n11773 ) | ( n9846 & n11773 ) ;
  assign n11775 = ( n2213 & n2269 ) | ( n2213 & ~n2773 ) | ( n2269 & ~n2773 ) ;
  assign n11776 = n7407 ^ n5003 ^ n3582 ;
  assign n11777 = n10912 & ~n11776 ;
  assign n11778 = ~n6601 & n11777 ;
  assign n11779 = n6119 | n11778 ;
  assign n11784 = n288 & n3345 ;
  assign n11785 = n11784 ^ n3379 ^ 1'b0 ;
  assign n11781 = n2950 & ~n6991 ;
  assign n11782 = ~n5345 & n11781 ;
  assign n11780 = n1933 & n10257 ;
  assign n11783 = n11782 ^ n11780 ^ 1'b0 ;
  assign n11786 = n11785 ^ n11783 ^ n6628 ;
  assign n11787 = n7329 ^ n624 ^ n324 ;
  assign n11788 = ( n7446 & n11651 ) | ( n7446 & ~n11787 ) | ( n11651 & ~n11787 ) ;
  assign n11789 = n6588 ^ n2153 ^ n1744 ;
  assign n11790 = n11789 ^ n9704 ^ n7008 ;
  assign n11792 = ( n910 & n2307 ) | ( n910 & n7828 ) | ( n2307 & n7828 ) ;
  assign n11793 = n3057 | n11792 ;
  assign n11791 = n5354 & ~n5683 ;
  assign n11794 = n11793 ^ n11791 ^ 1'b0 ;
  assign n11795 = n3189 ^ n1933 ^ 1'b0 ;
  assign n11796 = n11795 ^ n8476 ^ n3084 ;
  assign n11797 = n1798 & ~n11796 ;
  assign n11803 = n2138 | n4135 ;
  assign n11804 = n11803 ^ n6025 ^ n2026 ;
  assign n11805 = n10344 & n11804 ;
  assign n11806 = n11259 & n11805 ;
  assign n11798 = n2420 | n5674 ;
  assign n11799 = n11798 ^ n183 ^ 1'b0 ;
  assign n11800 = n4713 & n11646 ;
  assign n11801 = ~n11799 & n11800 ;
  assign n11802 = n600 | n11801 ;
  assign n11807 = n11806 ^ n11802 ^ 1'b0 ;
  assign n11808 = n11807 ^ n9840 ^ n5641 ;
  assign n11809 = n3522 ^ n2134 ^ 1'b0 ;
  assign n11810 = n646 | n11809 ;
  assign n11811 = n6506 ^ n3418 ^ n2378 ;
  assign n11812 = n11811 ^ n753 ^ 1'b0 ;
  assign n11813 = n986 & n11812 ;
  assign n11814 = n6203 ^ n2493 ^ n1659 ;
  assign n11815 = n10018 ^ n904 ^ 1'b0 ;
  assign n11816 = ~n1308 & n11815 ;
  assign n11817 = n11814 & n11816 ;
  assign n11821 = n6019 ^ n4733 ^ 1'b0 ;
  assign n11822 = n11821 ^ n9647 ^ n7957 ;
  assign n11819 = n249 & n1299 ;
  assign n11818 = ~n577 & n1240 ;
  assign n11820 = n11819 ^ n11818 ^ 1'b0 ;
  assign n11823 = n11822 ^ n11820 ^ 1'b0 ;
  assign n11824 = ~n8964 & n11216 ;
  assign n11825 = n9135 ^ n6087 ^ 1'b0 ;
  assign n11826 = n5891 & ~n11825 ;
  assign n11827 = ( ~n289 & n859 ) | ( ~n289 & n7600 ) | ( n859 & n7600 ) ;
  assign n11828 = n11827 ^ n8129 ^ n4271 ;
  assign n11829 = ( n3733 & n9257 ) | ( n3733 & ~n11828 ) | ( n9257 & ~n11828 ) ;
  assign n11830 = n7257 ^ n3299 ^ 1'b0 ;
  assign n11831 = ~n3272 & n11830 ;
  assign n11832 = n3985 & n11831 ;
  assign n11833 = ( n11038 & n11829 ) | ( n11038 & n11832 ) | ( n11829 & n11832 ) ;
  assign n11834 = ~n910 & n7934 ;
  assign n11835 = n5911 & n11834 ;
  assign n11836 = n11835 ^ n6600 ^ n4281 ;
  assign n11837 = x68 & ~n2421 ;
  assign n11838 = n11837 ^ n6042 ^ 1'b0 ;
  assign n11839 = n11838 ^ n4884 ^ 1'b0 ;
  assign n11840 = n10172 | n11839 ;
  assign n11841 = n11840 ^ n3024 ^ n2604 ;
  assign n11842 = n7401 ^ n2551 ^ n2426 ;
  assign n11843 = n11842 ^ n4325 ^ 1'b0 ;
  assign n11844 = n8904 ^ n5814 ^ n2198 ;
  assign n11849 = n6330 & n7127 ;
  assign n11850 = n9378 & n11849 ;
  assign n11851 = n11850 ^ n4680 ^ 1'b0 ;
  assign n11852 = n11851 ^ n9612 ^ n9261 ;
  assign n11845 = n231 & n6679 ;
  assign n11846 = n11845 ^ n4159 ^ 1'b0 ;
  assign n11847 = n5507 & ~n11846 ;
  assign n11848 = n11847 ^ n2004 ^ 1'b0 ;
  assign n11853 = n11852 ^ n11848 ^ n1134 ;
  assign n11854 = n6291 ^ n2614 ^ n1395 ;
  assign n11858 = n4918 ^ n2622 ^ n2403 ;
  assign n11857 = n10740 ^ n1403 ^ n1146 ;
  assign n11859 = n11858 ^ n11857 ^ 1'b0 ;
  assign n11855 = n4268 ^ n1226 ^ n495 ;
  assign n11856 = n3487 & n11855 ;
  assign n11860 = n11859 ^ n11856 ^ 1'b0 ;
  assign n11861 = n3918 & ~n11860 ;
  assign n11862 = n11861 ^ n2811 ^ 1'b0 ;
  assign n11863 = ~n788 & n1338 ;
  assign n11864 = ~n166 & n11863 ;
  assign n11865 = n10207 ^ n3232 ^ 1'b0 ;
  assign n11866 = n3959 & ~n11865 ;
  assign n11867 = n3906 ^ n2435 ^ n2255 ;
  assign n11868 = n11867 ^ n4518 ^ 1'b0 ;
  assign n11869 = n11866 & ~n11868 ;
  assign n11870 = n11869 ^ n4385 ^ 1'b0 ;
  assign n11871 = n11864 | n11870 ;
  assign n11872 = n5732 & ~n11303 ;
  assign n11873 = n9171 ^ n3218 ^ n2782 ;
  assign n11874 = n11872 & n11873 ;
  assign n11875 = n11874 ^ n8023 ^ 1'b0 ;
  assign n11877 = n2121 ^ n1049 ^ n921 ;
  assign n11876 = ( ~n1129 & n3749 ) | ( ~n1129 & n7594 ) | ( n3749 & n7594 ) ;
  assign n11878 = n11877 ^ n11876 ^ 1'b0 ;
  assign n11879 = ~n6674 & n11878 ;
  assign n11880 = n3134 ^ n1010 ^ n913 ;
  assign n11881 = n10889 ^ n4688 ^ n4426 ;
  assign n11882 = n11881 ^ n1019 ^ n264 ;
  assign n11883 = n9712 ^ n1608 ^ 1'b0 ;
  assign n11884 = n6776 & ~n11883 ;
  assign n11885 = n11884 ^ n4989 ^ n1511 ;
  assign n11892 = n2795 ^ n2377 ^ 1'b0 ;
  assign n11890 = n10356 & n10578 ;
  assign n11891 = n849 & n11890 ;
  assign n11886 = ( n3061 & n3862 ) | ( n3061 & n4555 ) | ( n3862 & n4555 ) ;
  assign n11887 = n2842 & ~n11886 ;
  assign n11888 = n2449 & n11887 ;
  assign n11889 = n9131 & ~n11888 ;
  assign n11893 = n11892 ^ n11891 ^ n11889 ;
  assign n11894 = ( ~n6127 & n6254 ) | ( ~n6127 & n7930 ) | ( n6254 & n7930 ) ;
  assign n11895 = n11894 ^ n7268 ^ 1'b0 ;
  assign n11896 = n7992 & n11895 ;
  assign n11898 = ( n796 & ~n4511 ) | ( n796 & n5332 ) | ( ~n4511 & n5332 ) ;
  assign n11897 = ~n2567 & n5816 ;
  assign n11899 = n11898 ^ n11897 ^ 1'b0 ;
  assign n11900 = n5449 & ~n11899 ;
  assign n11901 = n11900 ^ n6262 ^ 1'b0 ;
  assign n11902 = n700 & ~n10212 ;
  assign n11903 = ~n11901 & n11902 ;
  assign n11904 = ~n2660 & n11456 ;
  assign n11905 = n8674 & n11904 ;
  assign n11906 = ~n874 & n6544 ;
  assign n11907 = n11906 ^ n7644 ^ 1'b0 ;
  assign n11908 = n11907 ^ n1475 ^ n859 ;
  assign n11909 = n9165 & n11908 ;
  assign n11910 = n11909 ^ n4778 ^ 1'b0 ;
  assign n11911 = n11910 ^ n5859 ^ 1'b0 ;
  assign n11912 = n1522 ^ n148 ^ 1'b0 ;
  assign n11913 = n11912 ^ n6761 ^ n2851 ;
  assign n11914 = n2209 & n2726 ;
  assign n11915 = n1677 & n7484 ;
  assign n11916 = ~n9605 & n11915 ;
  assign n11917 = n4094 & ~n11916 ;
  assign n11918 = ( n7100 & ~n11914 ) | ( n7100 & n11917 ) | ( ~n11914 & n11917 ) ;
  assign n11919 = n10317 & n11918 ;
  assign n11920 = n960 & ~n9444 ;
  assign n11921 = n7690 & n11920 ;
  assign n11922 = n7911 ^ n3769 ^ n3555 ;
  assign n11923 = n7546 & ~n11922 ;
  assign n11924 = n11923 ^ n3242 ^ 1'b0 ;
  assign n11925 = n11924 ^ n3569 ^ n2179 ;
  assign n11926 = n11925 ^ n4525 ^ n366 ;
  assign n11931 = n1273 & n1815 ;
  assign n11932 = n11931 ^ n9167 ^ 1'b0 ;
  assign n11927 = ~n5937 & n7065 ;
  assign n11928 = n11927 ^ n2938 ^ 1'b0 ;
  assign n11929 = n10043 | n11928 ;
  assign n11930 = ( n2773 & ~n6019 ) | ( n2773 & n11929 ) | ( ~n6019 & n11929 ) ;
  assign n11933 = n11932 ^ n11930 ^ 1'b0 ;
  assign n11934 = n3101 | n10441 ;
  assign n11935 = n11934 ^ n4205 ^ 1'b0 ;
  assign n11936 = ~n561 & n1737 ;
  assign n11937 = ( n7130 & n11049 ) | ( n7130 & n11936 ) | ( n11049 & n11936 ) ;
  assign n11938 = ( ~n7065 & n11935 ) | ( ~n7065 & n11937 ) | ( n11935 & n11937 ) ;
  assign n11939 = ~n863 & n4961 ;
  assign n11940 = n2894 & n10703 ;
  assign n11941 = n11940 ^ n9331 ^ n6506 ;
  assign n11942 = ~n8847 & n11941 ;
  assign n11943 = n3461 | n11942 ;
  assign n11949 = n11140 ^ n10459 ^ n865 ;
  assign n11950 = n11949 ^ n6344 ^ 1'b0 ;
  assign n11944 = n2147 | n5187 ;
  assign n11945 = n8297 | n11944 ;
  assign n11946 = n5906 ^ n3147 ^ 1'b0 ;
  assign n11947 = n1244 & ~n11946 ;
  assign n11948 = n11945 & n11947 ;
  assign n11951 = n11950 ^ n11948 ^ 1'b0 ;
  assign n11952 = ~n2420 & n3586 ;
  assign n11953 = n8281 | n11952 ;
  assign n11954 = n10172 ^ n3123 ^ n2760 ;
  assign n11955 = n7193 ^ n5554 ^ 1'b0 ;
  assign n11956 = ( ~n6871 & n9108 ) | ( ~n6871 & n11955 ) | ( n9108 & n11955 ) ;
  assign n11957 = n343 & n11956 ;
  assign n11958 = n11957 ^ n11337 ^ 1'b0 ;
  assign n11959 = n5342 ^ n2398 ^ n1356 ;
  assign n11960 = ~n6913 & n11959 ;
  assign n11961 = n1022 | n11696 ;
  assign n11962 = n11961 ^ n9358 ^ n738 ;
  assign n11963 = n10213 ^ n4954 ^ 1'b0 ;
  assign n11964 = n11786 & ~n11963 ;
  assign n11965 = ~n332 & n8379 ;
  assign n11966 = n4471 & n11965 ;
  assign n11967 = n247 & n5052 ;
  assign n11968 = ( n10639 & n11687 ) | ( n10639 & ~n11967 ) | ( n11687 & ~n11967 ) ;
  assign n11969 = n4641 ^ n141 ^ 1'b0 ;
  assign n11970 = n11246 ^ n10942 ^ n4771 ;
  assign n11974 = x112 & ~n3193 ;
  assign n11975 = n11974 ^ n1830 ^ 1'b0 ;
  assign n11971 = n9223 ^ n3110 ^ 1'b0 ;
  assign n11972 = x98 & n11971 ;
  assign n11973 = n11972 ^ n11428 ^ n3186 ;
  assign n11976 = n11975 ^ n11973 ^ n10301 ;
  assign n11977 = ( n2459 & n3346 ) | ( n2459 & n7762 ) | ( n3346 & n7762 ) ;
  assign n11978 = n6639 ^ n4765 ^ n253 ;
  assign n11979 = n11978 ^ n10950 ^ n9236 ;
  assign n11980 = n4306 ^ n179 ^ 1'b0 ;
  assign n11981 = n11980 ^ n656 ^ 1'b0 ;
  assign n11982 = n11725 & ~n11981 ;
  assign n11983 = ~n1636 & n8948 ;
  assign n11984 = n11983 ^ n7633 ^ n7585 ;
  assign n11985 = n11984 ^ n589 ^ 1'b0 ;
  assign n11986 = n1447 ^ n1405 ^ 1'b0 ;
  assign n11987 = n11986 ^ n4248 ^ 1'b0 ;
  assign n11988 = n3379 | n11987 ;
  assign n11989 = n11988 ^ n5813 ^ n2660 ;
  assign n11990 = ( ~n1005 & n3914 ) | ( ~n1005 & n11989 ) | ( n3914 & n11989 ) ;
  assign n11991 = n6690 ^ n2418 ^ n592 ;
  assign n11992 = ( n3696 & ~n6500 ) | ( n3696 & n11991 ) | ( ~n6500 & n11991 ) ;
  assign n11993 = n11992 ^ n11938 ^ 1'b0 ;
  assign n11994 = n4447 ^ n2197 ^ n2110 ;
  assign n11995 = n10739 ^ n5058 ^ 1'b0 ;
  assign n11996 = ( n7926 & n11994 ) | ( n7926 & ~n11995 ) | ( n11994 & ~n11995 ) ;
  assign n11997 = n5320 & n11996 ;
  assign n11998 = n11997 ^ n4951 ^ n766 ;
  assign n11999 = n5382 ^ n3212 ^ 1'b0 ;
  assign n12000 = ( n686 & ~n9905 ) | ( n686 & n11999 ) | ( ~n9905 & n11999 ) ;
  assign n12001 = n6756 ^ n151 ^ 1'b0 ;
  assign n12002 = ( n6010 & n12000 ) | ( n6010 & ~n12001 ) | ( n12000 & ~n12001 ) ;
  assign n12003 = ( n4415 & n5249 ) | ( n4415 & ~n6639 ) | ( n5249 & ~n6639 ) ;
  assign n12004 = ( ~n6182 & n7692 ) | ( ~n6182 & n12003 ) | ( n7692 & n12003 ) ;
  assign n12008 = n6399 ^ n4957 ^ n3364 ;
  assign n12009 = ( n376 & n6159 ) | ( n376 & n12008 ) | ( n6159 & n12008 ) ;
  assign n12010 = ( n1486 & n4257 ) | ( n1486 & n12009 ) | ( n4257 & n12009 ) ;
  assign n12005 = ~n3450 & n4262 ;
  assign n12006 = n12005 ^ n5747 ^ 1'b0 ;
  assign n12007 = n2775 & n12006 ;
  assign n12011 = n12010 ^ n12007 ^ 1'b0 ;
  assign n12012 = n10845 & n12011 ;
  assign n12013 = n9473 ^ n6454 ^ 1'b0 ;
  assign n12014 = n1717 & n12013 ;
  assign n12015 = n11038 ^ n2865 ^ 1'b0 ;
  assign n12016 = ( ~n5956 & n11881 ) | ( ~n5956 & n12015 ) | ( n11881 & n12015 ) ;
  assign n12017 = n12016 ^ n2616 ^ n2013 ;
  assign n12018 = ( n969 & ~n2380 ) | ( n969 & n5909 ) | ( ~n2380 & n5909 ) ;
  assign n12019 = ( n6090 & n11867 ) | ( n6090 & ~n12018 ) | ( n11867 & ~n12018 ) ;
  assign n12022 = n10784 ^ n1437 ^ n187 ;
  assign n12020 = n884 & n5313 ;
  assign n12021 = ( n1477 & n6015 ) | ( n1477 & ~n12020 ) | ( n6015 & ~n12020 ) ;
  assign n12023 = n12022 ^ n12021 ^ n4562 ;
  assign n12024 = n8454 ^ n4715 ^ n1933 ;
  assign n12025 = ( n4859 & n6136 ) | ( n4859 & n12024 ) | ( n6136 & n12024 ) ;
  assign n12033 = n7718 ^ n7414 ^ n6151 ;
  assign n12026 = n2468 & ~n3385 ;
  assign n12027 = n9553 & n12026 ;
  assign n12028 = n12027 ^ n11562 ^ n1991 ;
  assign n12029 = n6703 ^ n4614 ^ n2435 ;
  assign n12030 = ~n4142 & n12029 ;
  assign n12031 = n12030 ^ n8583 ^ 1'b0 ;
  assign n12032 = ( ~n6406 & n12028 ) | ( ~n6406 & n12031 ) | ( n12028 & n12031 ) ;
  assign n12034 = n12033 ^ n12032 ^ n392 ;
  assign n12035 = n3548 ^ n275 ^ 1'b0 ;
  assign n12036 = ( n4274 & n8439 ) | ( n4274 & ~n12035 ) | ( n8439 & ~n12035 ) ;
  assign n12037 = n9797 | n12036 ;
  assign n12038 = n1856 & n2733 ;
  assign n12039 = ( n4048 & n8701 ) | ( n4048 & n12038 ) | ( n8701 & n12038 ) ;
  assign n12044 = ( n192 & n4571 ) | ( n192 & n7671 ) | ( n4571 & n7671 ) ;
  assign n12045 = n12044 ^ n2293 ^ n253 ;
  assign n12041 = n6354 ^ n374 ^ 1'b0 ;
  assign n12042 = n3944 & n12041 ;
  assign n12040 = n6081 | n9852 ;
  assign n12043 = n12042 ^ n12040 ^ 1'b0 ;
  assign n12046 = n12045 ^ n12043 ^ n6991 ;
  assign n12047 = ~n5554 & n6373 ;
  assign n12048 = ~n10876 & n12047 ;
  assign n12051 = ( ~n4208 & n8125 ) | ( ~n4208 & n8389 ) | ( n8125 & n8389 ) ;
  assign n12049 = n1312 & ~n3041 ;
  assign n12050 = n9485 & ~n12049 ;
  assign n12052 = n12051 ^ n12050 ^ 1'b0 ;
  assign n12053 = n11329 ^ n2596 ^ 1'b0 ;
  assign n12054 = n6677 ^ x13 ^ 1'b0 ;
  assign n12055 = ( n4980 & ~n12053 ) | ( n4980 & n12054 ) | ( ~n12053 & n12054 ) ;
  assign n12056 = n5476 ^ n3661 ^ n2282 ;
  assign n12057 = n12056 ^ n11468 ^ n4162 ;
  assign n12058 = n3337 & n4716 ;
  assign n12059 = n6827 | n12058 ;
  assign n12060 = n6183 ^ n5252 ^ n342 ;
  assign n12061 = ( ~x1 & n1748 ) | ( ~x1 & n4976 ) | ( n1748 & n4976 ) ;
  assign n12062 = ~n6310 & n12061 ;
  assign n12063 = ( ~n315 & n7124 ) | ( ~n315 & n11160 ) | ( n7124 & n11160 ) ;
  assign n12064 = ( n1684 & ~n2255 ) | ( n1684 & n12063 ) | ( ~n2255 & n12063 ) ;
  assign n12068 = n9737 ^ n710 ^ n575 ;
  assign n12065 = n1144 & ~n7053 ;
  assign n12066 = ~n3553 & n12065 ;
  assign n12067 = n12066 ^ n3707 ^ n3638 ;
  assign n12069 = n12068 ^ n12067 ^ n10815 ;
  assign n12070 = ( n665 & n1827 ) | ( n665 & ~n7889 ) | ( n1827 & ~n7889 ) ;
  assign n12071 = n12070 ^ n4388 ^ 1'b0 ;
  assign n12072 = ( n5550 & n10302 ) | ( n5550 & n10963 ) | ( n10302 & n10963 ) ;
  assign n12073 = ( n4282 & ~n7358 ) | ( n4282 & n8550 ) | ( ~n7358 & n8550 ) ;
  assign n12074 = ~n486 & n12073 ;
  assign n12075 = n12074 ^ n6977 ^ 1'b0 ;
  assign n12076 = n7775 | n12075 ;
  assign n12077 = n12072 & ~n12076 ;
  assign n12078 = n12071 & ~n12077 ;
  assign n12079 = n12078 ^ n1583 ^ 1'b0 ;
  assign n12080 = n4407 & n10934 ;
  assign n12081 = n569 & ~n9163 ;
  assign n12082 = ~n1184 & n3811 ;
  assign n12083 = n12082 ^ n3316 ^ 1'b0 ;
  assign n12084 = n9288 & n10100 ;
  assign n12085 = ~n12083 & n12084 ;
  assign n12095 = n2409 ^ n2353 ^ 1'b0 ;
  assign n12086 = n5703 ^ n4019 ^ 1'b0 ;
  assign n12087 = n1126 & n12086 ;
  assign n12088 = ( n1049 & n1503 ) | ( n1049 & ~n3077 ) | ( n1503 & ~n3077 ) ;
  assign n12089 = ( n471 & ~n12087 ) | ( n471 & n12088 ) | ( ~n12087 & n12088 ) ;
  assign n12090 = n656 & ~n1785 ;
  assign n12091 = ~n731 & n12090 ;
  assign n12092 = n5177 | n12091 ;
  assign n12093 = n9675 | n12092 ;
  assign n12094 = ( n1905 & n12089 ) | ( n1905 & n12093 ) | ( n12089 & n12093 ) ;
  assign n12096 = n12095 ^ n12094 ^ 1'b0 ;
  assign n12097 = n7630 | n12096 ;
  assign n12098 = ( n136 & ~n1300 ) | ( n136 & n2695 ) | ( ~n1300 & n2695 ) ;
  assign n12099 = n12098 ^ n2864 ^ n1956 ;
  assign n12100 = ( n2077 & n3718 ) | ( n2077 & n5055 ) | ( n3718 & n5055 ) ;
  assign n12101 = ( x27 & n9629 ) | ( x27 & ~n10058 ) | ( n9629 & ~n10058 ) ;
  assign n12102 = n6655 & n8908 ;
  assign n12103 = n12102 ^ n7254 ^ 1'b0 ;
  assign n12104 = n9570 | n12103 ;
  assign n12105 = n10079 & ~n12104 ;
  assign n12106 = n6407 & n12105 ;
  assign n12107 = n3914 & ~n5185 ;
  assign n12108 = n225 | n2077 ;
  assign n12109 = n12108 ^ n5048 ^ 1'b0 ;
  assign n12110 = ( n6663 & n6910 ) | ( n6663 & n12109 ) | ( n6910 & n12109 ) ;
  assign n12114 = n3818 & n7859 ;
  assign n12115 = n1791 & n12114 ;
  assign n12116 = ( ~n2695 & n3409 ) | ( ~n2695 & n12115 ) | ( n3409 & n12115 ) ;
  assign n12112 = n3815 | n8263 ;
  assign n12113 = n12112 ^ n4112 ^ 1'b0 ;
  assign n12111 = ( n2834 & n7278 ) | ( n2834 & n10270 ) | ( n7278 & n10270 ) ;
  assign n12117 = n12116 ^ n12113 ^ n12111 ;
  assign n12118 = n9444 ^ n3836 ^ n1928 ;
  assign n12119 = n12118 ^ n8649 ^ n1422 ;
  assign n12120 = n2784 ^ n2126 ^ 1'b0 ;
  assign n12121 = ~n1977 & n12120 ;
  assign n12122 = n1034 | n3724 ;
  assign n12123 = n12122 ^ n4555 ^ 1'b0 ;
  assign n12124 = n12123 ^ n696 ^ 1'b0 ;
  assign n12125 = ~n12121 & n12124 ;
  assign n12128 = n3036 ^ n1124 ^ 1'b0 ;
  assign n12129 = n10301 | n12128 ;
  assign n12130 = n12129 ^ n7551 ^ n7143 ;
  assign n12126 = n5553 ^ n3293 ^ n2676 ;
  assign n12127 = ( n325 & ~n1160 ) | ( n325 & n12126 ) | ( ~n1160 & n12126 ) ;
  assign n12131 = n12130 ^ n12127 ^ n751 ;
  assign n12132 = ( n1819 & n5264 ) | ( n1819 & ~n10430 ) | ( n5264 & ~n10430 ) ;
  assign n12133 = n3643 ^ n2863 ^ 1'b0 ;
  assign n12134 = n1659 | n12133 ;
  assign n12139 = ~n405 & n4949 ;
  assign n12137 = n4969 ^ n2785 ^ n1953 ;
  assign n12135 = n572 | n1107 ;
  assign n12136 = n12135 ^ n1068 ^ 1'b0 ;
  assign n12138 = n12137 ^ n12136 ^ n8161 ;
  assign n12140 = n12139 ^ n12138 ^ 1'b0 ;
  assign n12141 = n12134 | n12140 ;
  assign n12142 = n3197 ^ n1953 ^ n1590 ;
  assign n12143 = n8766 & ~n12142 ;
  assign n12144 = n12143 ^ n197 ^ 1'b0 ;
  assign n12145 = n5804 | n10671 ;
  assign n12146 = ~n7481 & n12145 ;
  assign n12147 = ~n12144 & n12146 ;
  assign n12148 = n4515 ^ n1798 ^ n325 ;
  assign n12149 = ( n5206 & ~n8764 ) | ( n5206 & n12148 ) | ( ~n8764 & n12148 ) ;
  assign n12150 = n478 | n11950 ;
  assign n12151 = n12149 | n12150 ;
  assign n12155 = ( n2580 & n3253 ) | ( n2580 & ~n3882 ) | ( n3253 & ~n3882 ) ;
  assign n12152 = ( n4285 & ~n6657 ) | ( n4285 & n10887 ) | ( ~n6657 & n10887 ) ;
  assign n12153 = n9012 & ~n9838 ;
  assign n12154 = n12152 & n12153 ;
  assign n12156 = n12155 ^ n12154 ^ n565 ;
  assign n12161 = ~n4287 & n7925 ;
  assign n12162 = ~n6855 & n12161 ;
  assign n12159 = ~x66 & n10577 ;
  assign n12160 = n12159 ^ n2023 ^ 1'b0 ;
  assign n12157 = ( n179 & ~n5301 ) | ( n179 & n7917 ) | ( ~n5301 & n7917 ) ;
  assign n12158 = n1629 & n12157 ;
  assign n12163 = n12162 ^ n12160 ^ n12158 ;
  assign n12164 = x12 & ~n4412 ;
  assign n12165 = n8996 | n12164 ;
  assign n12166 = n11633 ^ n1277 ^ 1'b0 ;
  assign n12167 = n3467 & ~n12166 ;
  assign n12168 = ~n1200 & n3659 ;
  assign n12169 = n12168 ^ n1532 ^ 1'b0 ;
  assign n12170 = n6067 ^ n5027 ^ n3586 ;
  assign n12171 = ~n11916 & n12170 ;
  assign n12172 = ~n12169 & n12171 ;
  assign n12173 = n11530 ^ n5631 ^ 1'b0 ;
  assign n12174 = ~n6716 & n12173 ;
  assign n12175 = ~n7105 & n12174 ;
  assign n12176 = n12175 ^ n5725 ^ 1'b0 ;
  assign n12177 = ( n1672 & n5186 ) | ( n1672 & ~n9093 ) | ( n5186 & ~n9093 ) ;
  assign n12178 = ~n3166 & n12177 ;
  assign n12179 = n8247 | n12178 ;
  assign n12180 = n12179 ^ n1572 ^ 1'b0 ;
  assign n12181 = n6480 ^ n568 ^ n405 ;
  assign n12182 = ~n6881 & n12181 ;
  assign n12183 = n12182 ^ n5605 ^ 1'b0 ;
  assign n12184 = ( x81 & n1639 ) | ( x81 & ~n2232 ) | ( n1639 & ~n2232 ) ;
  assign n12185 = n12184 ^ n716 ^ 1'b0 ;
  assign n12186 = n4471 | n12185 ;
  assign n12187 = ( n3875 & n7030 ) | ( n3875 & n12186 ) | ( n7030 & n12186 ) ;
  assign n12188 = ( n12180 & n12183 ) | ( n12180 & ~n12187 ) | ( n12183 & ~n12187 ) ;
  assign n12189 = ~n1589 & n10432 ;
  assign n12190 = n12189 ^ n5165 ^ 1'b0 ;
  assign n12191 = ( ~n2718 & n3207 ) | ( ~n2718 & n5408 ) | ( n3207 & n5408 ) ;
  assign n12192 = n12191 ^ n7679 ^ n2555 ;
  assign n12193 = n10719 ^ n9296 ^ n6396 ;
  assign n12194 = n724 | n12193 ;
  assign n12197 = ~n4354 & n7904 ;
  assign n12198 = ~n2683 & n12197 ;
  assign n12195 = x100 & ~n4205 ;
  assign n12196 = ~x32 & n12195 ;
  assign n12199 = n12198 ^ n12196 ^ 1'b0 ;
  assign n12200 = ~n5390 & n12199 ;
  assign n12201 = n3562 ^ n365 ^ 1'b0 ;
  assign n12202 = ( n1894 & n1952 ) | ( n1894 & n4607 ) | ( n1952 & n4607 ) ;
  assign n12203 = n12202 ^ n5673 ^ n4795 ;
  assign n12204 = n12203 ^ n8216 ^ 1'b0 ;
  assign n12205 = n12201 & n12204 ;
  assign n12206 = ( ~n3253 & n4812 ) | ( ~n3253 & n6153 ) | ( n4812 & n6153 ) ;
  assign n12207 = ( n584 & n5898 ) | ( n584 & n12206 ) | ( n5898 & n12206 ) ;
  assign n12208 = ( n4702 & ~n10113 ) | ( n4702 & n12207 ) | ( ~n10113 & n12207 ) ;
  assign n12209 = n218 | n10961 ;
  assign n12210 = n12209 ^ n11315 ^ 1'b0 ;
  assign n12220 = n2946 & n11235 ;
  assign n12221 = n12220 ^ n582 ^ 1'b0 ;
  assign n12222 = n12221 ^ n7132 ^ x107 ;
  assign n12215 = n3316 ^ n2839 ^ 1'b0 ;
  assign n12216 = n2622 & n12215 ;
  assign n12217 = n4531 & n12216 ;
  assign n12218 = n12217 ^ n5728 ^ n2103 ;
  assign n12211 = n3160 | n9793 ;
  assign n12212 = n12211 ^ n5079 ^ 1'b0 ;
  assign n12213 = n3481 | n12212 ;
  assign n12214 = n9444 & ~n12213 ;
  assign n12219 = n12218 ^ n12214 ^ n7377 ;
  assign n12223 = n12222 ^ n12219 ^ n9756 ;
  assign n12224 = n2484 ^ n2171 ^ n1316 ;
  assign n12225 = n12224 ^ n7728 ^ n5080 ;
  assign n12226 = n12225 ^ n10636 ^ 1'b0 ;
  assign n12227 = n1447 & ~n10277 ;
  assign n12228 = n6665 & n12227 ;
  assign n12229 = ~n243 & n2253 ;
  assign n12230 = n12229 ^ n2209 ^ 1'b0 ;
  assign n12231 = ~n11215 & n12230 ;
  assign n12232 = n12231 ^ n5005 ^ n3063 ;
  assign n12233 = ( x2 & n1429 ) | ( x2 & ~n2433 ) | ( n1429 & ~n2433 ) ;
  assign n12234 = ( n7328 & n12232 ) | ( n7328 & ~n12233 ) | ( n12232 & ~n12233 ) ;
  assign n12235 = n5788 ^ n4555 ^ 1'b0 ;
  assign n12236 = n12235 ^ n2257 ^ n1174 ;
  assign n12237 = n9017 & n12236 ;
  assign n12238 = n2805 ^ n1283 ^ 1'b0 ;
  assign n12239 = n12238 ^ n4700 ^ n393 ;
  assign n12240 = n6889 & n9595 ;
  assign n12241 = ~n10942 & n12240 ;
  assign n12242 = n2601 & n7673 ;
  assign n12243 = ( n12239 & n12241 ) | ( n12239 & ~n12242 ) | ( n12241 & ~n12242 ) ;
  assign n12244 = n10526 ^ n4112 ^ n3596 ;
  assign n12245 = n1595 & n12244 ;
  assign n12246 = n4959 & ~n12245 ;
  assign n12247 = n12246 ^ n2308 ^ 1'b0 ;
  assign n12248 = n12247 ^ n6358 ^ n2607 ;
  assign n12249 = n5473 & ~n5987 ;
  assign n12250 = ~n1300 & n4492 ;
  assign n12251 = n12250 ^ n7482 ^ 1'b0 ;
  assign n12252 = n12251 ^ n11239 ^ n5150 ;
  assign n12253 = n2900 & n12252 ;
  assign n12254 = ( n6392 & n6858 ) | ( n6392 & n12228 ) | ( n6858 & n12228 ) ;
  assign n12255 = ( n1468 & n2943 ) | ( n1468 & n5335 ) | ( n2943 & n5335 ) ;
  assign n12256 = ( ~x94 & n7030 ) | ( ~x94 & n12255 ) | ( n7030 & n12255 ) ;
  assign n12258 = n8383 ^ n1005 ^ 1'b0 ;
  assign n12259 = n1111 | n12258 ;
  assign n12257 = n895 & ~n4687 ;
  assign n12260 = n12259 ^ n12257 ^ 1'b0 ;
  assign n12261 = n1924 & ~n2555 ;
  assign n12262 = ~n1905 & n12261 ;
  assign n12263 = n12262 ^ n5149 ^ n850 ;
  assign n12264 = n12263 ^ n11506 ^ 1'b0 ;
  assign n12265 = n12070 & ~n12264 ;
  assign n12266 = n12260 & n12265 ;
  assign n12267 = n12256 & n12266 ;
  assign n12271 = ~n6215 & n8570 ;
  assign n12268 = n166 & ~n1253 ;
  assign n12269 = ( n3830 & n11683 ) | ( n3830 & n12268 ) | ( n11683 & n12268 ) ;
  assign n12270 = n12269 ^ n10589 ^ 1'b0 ;
  assign n12272 = n12271 ^ n12270 ^ x30 ;
  assign n12273 = ( n335 & n3347 ) | ( n335 & ~n4310 ) | ( n3347 & ~n4310 ) ;
  assign n12274 = n3485 | n12273 ;
  assign n12275 = n12274 ^ n10979 ^ n8559 ;
  assign n12276 = ( n2291 & n11313 ) | ( n2291 & n12275 ) | ( n11313 & n12275 ) ;
  assign n12277 = n5383 & n7772 ;
  assign n12278 = n12277 ^ n4220 ^ 1'b0 ;
  assign n12279 = n6179 ^ n6112 ^ n4192 ;
  assign n12280 = ~n284 & n12279 ;
  assign n12281 = ~n12278 & n12280 ;
  assign n12282 = n7753 ^ n6891 ^ 1'b0 ;
  assign n12283 = ( n814 & ~n1105 ) | ( n814 & n11034 ) | ( ~n1105 & n11034 ) ;
  assign n12284 = n12283 ^ x123 ^ 1'b0 ;
  assign n12285 = n6608 ^ n2137 ^ 1'b0 ;
  assign n12286 = ( n2212 & ~n4856 ) | ( n2212 & n12285 ) | ( ~n4856 & n12285 ) ;
  assign n12287 = n12286 ^ n10507 ^ 1'b0 ;
  assign n12288 = n858 & ~n12287 ;
  assign n12289 = n9677 ^ n665 ^ 1'b0 ;
  assign n12290 = n10167 ^ n1967 ^ n568 ;
  assign n12291 = n2795 & n7370 ;
  assign n12292 = n12291 ^ n8615 ^ 1'b0 ;
  assign n12293 = ( n1660 & n4670 ) | ( n1660 & n9397 ) | ( n4670 & n9397 ) ;
  assign n12294 = n12293 ^ n8010 ^ 1'b0 ;
  assign n12299 = ~n990 & n4221 ;
  assign n12297 = n8505 ^ n3828 ^ n1599 ;
  assign n12298 = n6973 & n12297 ;
  assign n12295 = n8389 ^ n7667 ^ n7318 ;
  assign n12296 = n12295 ^ n8173 ^ n6985 ;
  assign n12300 = n12299 ^ n12298 ^ n12296 ;
  assign n12301 = ( n7935 & n10415 ) | ( n7935 & n12148 ) | ( n10415 & n12148 ) ;
  assign n12302 = n8352 & n10918 ;
  assign n12303 = n2700 & n8779 ;
  assign n12304 = n12303 ^ n10934 ^ 1'b0 ;
  assign n12305 = n2385 & ~n2553 ;
  assign n12306 = ( n4745 & ~n7288 ) | ( n4745 & n12305 ) | ( ~n7288 & n12305 ) ;
  assign n12307 = n7187 ^ n5773 ^ n2615 ;
  assign n12308 = n12307 ^ n374 ^ 1'b0 ;
  assign n12309 = n12043 | n12308 ;
  assign n12310 = n12306 & ~n12309 ;
  assign n12311 = x32 & n1481 ;
  assign n12312 = n4581 | n12311 ;
  assign n12313 = n12312 ^ n6596 ^ 1'b0 ;
  assign n12315 = ( n6980 & n8224 ) | ( n6980 & n11818 ) | ( n8224 & n11818 ) ;
  assign n12316 = n10930 | n12315 ;
  assign n12314 = n2504 | n8709 ;
  assign n12317 = n12316 ^ n12314 ^ 1'b0 ;
  assign n12318 = n1142 | n2713 ;
  assign n12319 = n714 | n12318 ;
  assign n12320 = n6319 ^ n1375 ^ n572 ;
  assign n12321 = n12320 ^ n1375 ^ n1041 ;
  assign n12322 = ( ~n10324 & n12319 ) | ( ~n10324 & n12321 ) | ( n12319 & n12321 ) ;
  assign n12323 = n12322 ^ n2751 ^ 1'b0 ;
  assign n12324 = n12323 ^ n7398 ^ 1'b0 ;
  assign n12325 = n2272 & n2834 ;
  assign n12326 = n12325 ^ n2495 ^ 1'b0 ;
  assign n12327 = n12326 ^ n4093 ^ 1'b0 ;
  assign n12328 = n4521 ^ n3225 ^ 1'b0 ;
  assign n12329 = n12327 & ~n12328 ;
  assign n12330 = n2049 | n5978 ;
  assign n12331 = n2468 | n12330 ;
  assign n12332 = n9866 & n12331 ;
  assign n12333 = ~n12329 & n12332 ;
  assign n12334 = n10532 ^ n6373 ^ 1'b0 ;
  assign n12335 = ( n1896 & n8286 ) | ( n1896 & ~n11400 ) | ( n8286 & ~n11400 ) ;
  assign n12336 = n1275 | n9793 ;
  assign n12337 = n7448 ^ n3195 ^ 1'b0 ;
  assign n12338 = n614 | n3875 ;
  assign n12339 = n9528 | n12338 ;
  assign n12340 = ~n6927 & n12339 ;
  assign n12341 = n12340 ^ n6867 ^ 1'b0 ;
  assign n12342 = ( ~n520 & n11682 ) | ( ~n520 & n12341 ) | ( n11682 & n12341 ) ;
  assign n12343 = ( n5159 & n11511 ) | ( n5159 & ~n12188 ) | ( n11511 & ~n12188 ) ;
  assign n12344 = n4436 ^ n3930 ^ n3816 ;
  assign n12345 = n12344 ^ n7679 ^ n5268 ;
  assign n12346 = n12345 ^ n3886 ^ 1'b0 ;
  assign n12347 = n1899 | n12346 ;
  assign n12352 = ( n1740 & n1808 ) | ( n1740 & n4879 ) | ( n1808 & n4879 ) ;
  assign n12353 = n796 & ~n12352 ;
  assign n12348 = n4390 & ~n4620 ;
  assign n12349 = n12348 ^ n4363 ^ 1'b0 ;
  assign n12350 = ( n4298 & n4795 ) | ( n4298 & n12349 ) | ( n4795 & n12349 ) ;
  assign n12351 = ( n2743 & n6354 ) | ( n2743 & n12350 ) | ( n6354 & n12350 ) ;
  assign n12354 = n12353 ^ n12351 ^ n3337 ;
  assign n12355 = n12354 ^ n11758 ^ n2485 ;
  assign n12356 = ~n2265 & n4150 ;
  assign n12358 = ( ~n4202 & n4407 ) | ( ~n4202 & n5288 ) | ( n4407 & n5288 ) ;
  assign n12357 = n5523 ^ n3231 ^ n539 ;
  assign n12359 = n12358 ^ n12357 ^ n579 ;
  assign n12360 = ( ~n7231 & n12356 ) | ( ~n7231 & n12359 ) | ( n12356 & n12359 ) ;
  assign n12361 = n4943 | n8424 ;
  assign n12362 = n7888 | n12361 ;
  assign n12363 = n10195 ^ n6287 ^ n6142 ;
  assign n12364 = ~n5108 & n7090 ;
  assign n12365 = n12364 ^ n976 ^ 1'b0 ;
  assign n12366 = ~n1956 & n7452 ;
  assign n12367 = ( n697 & ~n7477 ) | ( n697 & n12366 ) | ( ~n7477 & n12366 ) ;
  assign n12368 = n12367 ^ n4930 ^ n4024 ;
  assign n12369 = ~n4307 & n12368 ;
  assign n12370 = n5834 & n7816 ;
  assign n12371 = ( n2839 & ~n2904 ) | ( n2839 & n11986 ) | ( ~n2904 & n11986 ) ;
  assign n12372 = n770 & ~n1609 ;
  assign n12373 = n12372 ^ n4429 ^ 1'b0 ;
  assign n12374 = n5560 & n12373 ;
  assign n12375 = n12058 ^ n10432 ^ n7230 ;
  assign n12376 = ( x6 & n12374 ) | ( x6 & n12375 ) | ( n12374 & n12375 ) ;
  assign n12379 = ~n5535 & n8585 ;
  assign n12377 = n9609 ^ n5665 ^ 1'b0 ;
  assign n12378 = n9190 & ~n12377 ;
  assign n12380 = n12379 ^ n12378 ^ 1'b0 ;
  assign n12381 = n4129 & ~n6392 ;
  assign n12383 = n2324 | n4116 ;
  assign n12384 = n5959 & ~n12383 ;
  assign n12382 = ~n3650 & n3758 ;
  assign n12385 = n12384 ^ n12382 ^ 1'b0 ;
  assign n12386 = n4468 & ~n8788 ;
  assign n12387 = ~n6830 & n12386 ;
  assign n12388 = n8369 | n12387 ;
  assign n12389 = n12388 ^ n5034 ^ 1'b0 ;
  assign n12390 = n2444 & n12389 ;
  assign n12391 = n12343 ^ n5226 ^ n1068 ;
  assign n12392 = n7847 ^ n4337 ^ 1'b0 ;
  assign n12393 = n12392 ^ n9070 ^ n6768 ;
  assign n12394 = n1233 & n10096 ;
  assign n12395 = n12394 ^ n3713 ^ 1'b0 ;
  assign n12396 = n12395 ^ n385 ^ 1'b0 ;
  assign n12397 = n12396 ^ n2138 ^ 1'b0 ;
  assign n12398 = ~n8288 & n12397 ;
  assign n12399 = n12398 ^ n8401 ^ 1'b0 ;
  assign n12400 = n515 & ~n2767 ;
  assign n12401 = n12400 ^ n2410 ^ n1029 ;
  assign n12402 = ( n926 & ~n5153 ) | ( n926 & n12401 ) | ( ~n5153 & n12401 ) ;
  assign n12403 = ~n9407 & n12402 ;
  assign n12404 = n12403 ^ n12103 ^ n4074 ;
  assign n12405 = ( n1597 & n7351 ) | ( n1597 & ~n10659 ) | ( n7351 & ~n10659 ) ;
  assign n12406 = ~n4638 & n6951 ;
  assign n12411 = ( n2701 & n3481 ) | ( n2701 & ~n6398 ) | ( n3481 & ~n6398 ) ;
  assign n12412 = ~n2718 & n12411 ;
  assign n12408 = n4851 ^ n4784 ^ n1082 ;
  assign n12409 = n12408 ^ n1158 ^ 1'b0 ;
  assign n12407 = n9096 ^ n9077 ^ n7222 ;
  assign n12410 = n12409 ^ n12407 ^ n1316 ;
  assign n12413 = n12412 ^ n12410 ^ 1'b0 ;
  assign n12414 = n7373 & ~n8037 ;
  assign n12415 = n206 & n12414 ;
  assign n12416 = n12415 ^ n7426 ^ n4805 ;
  assign n12417 = n969 | n12416 ;
  assign n12418 = n10910 ^ n1911 ^ n1605 ;
  assign n12419 = n12418 ^ n1817 ^ n156 ;
  assign n12420 = n1935 ^ n1572 ^ 1'b0 ;
  assign n12421 = n2206 & n12420 ;
  assign n12422 = n4751 & ~n11903 ;
  assign n12423 = ~n12421 & n12422 ;
  assign n12424 = n3871 ^ n1659 ^ 1'b0 ;
  assign n12425 = ( ~n1510 & n7438 ) | ( ~n1510 & n12424 ) | ( n7438 & n12424 ) ;
  assign n12426 = n12425 ^ n3151 ^ 1'b0 ;
  assign n12427 = n12426 ^ n5627 ^ n323 ;
  assign n12428 = ( ~n1001 & n3482 ) | ( ~n1001 & n6651 ) | ( n3482 & n6651 ) ;
  assign n12429 = n12428 ^ n4024 ^ 1'b0 ;
  assign n12430 = ( n983 & n2277 ) | ( n983 & n2789 ) | ( n2277 & n2789 ) ;
  assign n12431 = n12430 ^ n2434 ^ 1'b0 ;
  assign n12432 = n10087 ^ n3317 ^ 1'b0 ;
  assign n12433 = ( n3383 & n3826 ) | ( n3383 & ~n6080 ) | ( n3826 & ~n6080 ) ;
  assign n12434 = ( n5786 & n6741 ) | ( n5786 & n12433 ) | ( n6741 & n12433 ) ;
  assign n12435 = n5102 & n12424 ;
  assign n12436 = ~n2365 & n12435 ;
  assign n12437 = n12436 ^ n4711 ^ 1'b0 ;
  assign n12438 = n7649 & ~n12437 ;
  assign n12439 = n1391 & ~n2433 ;
  assign n12440 = n7690 & n12439 ;
  assign n12441 = ( n3088 & n6213 ) | ( n3088 & n9612 ) | ( n6213 & n9612 ) ;
  assign n12442 = ( n6155 & n9364 ) | ( n6155 & ~n12441 ) | ( n9364 & ~n12441 ) ;
  assign n12443 = n6879 ^ n2652 ^ n2176 ;
  assign n12444 = n12443 ^ n4426 ^ n4036 ;
  assign n12445 = ( n5051 & n5333 ) | ( n5051 & ~n9347 ) | ( n5333 & ~n9347 ) ;
  assign n12446 = n12445 ^ n4694 ^ 1'b0 ;
  assign n12447 = ~n11474 & n12446 ;
  assign n12448 = ~n4744 & n5271 ;
  assign n12449 = n7964 & n12448 ;
  assign n12451 = ( n187 & ~n229 ) | ( n187 & n10084 ) | ( ~n229 & n10084 ) ;
  assign n12452 = n12451 ^ n4264 ^ n2529 ;
  assign n12450 = n2502 | n4185 ;
  assign n12453 = n12452 ^ n12450 ^ 1'b0 ;
  assign n12454 = ( n11602 & ~n12449 ) | ( n11602 & n12453 ) | ( ~n12449 & n12453 ) ;
  assign n12455 = ( n2844 & n12447 ) | ( n2844 & n12454 ) | ( n12447 & n12454 ) ;
  assign n12456 = n8936 & n11052 ;
  assign n12457 = n7663 ^ n6634 ^ 1'b0 ;
  assign n12458 = n12281 & ~n12457 ;
  assign n12459 = n325 & n1991 ;
  assign n12460 = n12459 ^ n5811 ^ 1'b0 ;
  assign n12461 = ( n5098 & n6931 ) | ( n5098 & ~n8415 ) | ( n6931 & ~n8415 ) ;
  assign n12462 = ( n3386 & n4501 ) | ( n3386 & n10973 ) | ( n4501 & n10973 ) ;
  assign n12463 = n4075 & ~n11033 ;
  assign n12464 = ~n3203 & n12463 ;
  assign n12465 = n4383 ^ n3196 ^ 1'b0 ;
  assign n12466 = n12465 ^ n1651 ^ 1'b0 ;
  assign n12467 = n12464 | n12466 ;
  assign n12468 = n3904 | n12467 ;
  assign n12469 = ( n12461 & n12462 ) | ( n12461 & ~n12468 ) | ( n12462 & ~n12468 ) ;
  assign n12470 = n12307 ^ n12299 ^ n7971 ;
  assign n12471 = n3487 & n4776 ;
  assign n12472 = ~n4249 & n12471 ;
  assign n12473 = n5031 & n6324 ;
  assign n12474 = ~x95 & n12473 ;
  assign n12475 = n7694 & ~n12474 ;
  assign n12476 = n12472 & n12475 ;
  assign n12477 = n8380 ^ n5606 ^ 1'b0 ;
  assign n12478 = n12476 | n12477 ;
  assign n12479 = n2724 & ~n12478 ;
  assign n12480 = ( n238 & n395 ) | ( n238 & ~n2047 ) | ( n395 & ~n2047 ) ;
  assign n12481 = ( n1344 & ~n11815 ) | ( n1344 & n12480 ) | ( ~n11815 & n12480 ) ;
  assign n12485 = ~n743 & n1843 ;
  assign n12486 = n6073 | n12485 ;
  assign n12487 = n3387 & n6270 ;
  assign n12488 = ~n12486 & n12487 ;
  assign n12482 = ~n5276 & n10609 ;
  assign n12483 = n10952 & n12482 ;
  assign n12484 = n12483 ^ n10145 ^ n5600 ;
  assign n12489 = n12488 ^ n12484 ^ 1'b0 ;
  assign n12490 = n3115 ^ n1199 ^ 1'b0 ;
  assign n12491 = n7322 | n12490 ;
  assign n12492 = n12491 ^ n8459 ^ 1'b0 ;
  assign n12494 = ( n2168 & n3083 ) | ( n2168 & ~n3207 ) | ( n3083 & ~n3207 ) ;
  assign n12493 = n9660 ^ n3443 ^ x11 ;
  assign n12495 = n12494 ^ n12493 ^ n2169 ;
  assign n12496 = n12495 ^ n6022 ^ n1550 ;
  assign n12497 = n1225 ^ n1115 ^ 1'b0 ;
  assign n12498 = n10114 & ~n12497 ;
  assign n12499 = n813 ^ n628 ^ 1'b0 ;
  assign n12500 = n12498 & ~n12499 ;
  assign n12503 = n2962 & n5136 ;
  assign n12504 = n5775 ^ n4610 ^ n4148 ;
  assign n12505 = ( n4267 & n12503 ) | ( n4267 & ~n12504 ) | ( n12503 & ~n12504 ) ;
  assign n12501 = ( x120 & n286 ) | ( x120 & n733 ) | ( n286 & n733 ) ;
  assign n12502 = n12501 ^ n6095 ^ n2472 ;
  assign n12506 = n12505 ^ n12502 ^ 1'b0 ;
  assign n12507 = n9653 ^ n2367 ^ 1'b0 ;
  assign n12508 = n3195 & ~n12507 ;
  assign n12509 = n12472 ^ n9399 ^ n1940 ;
  assign n12510 = n5371 | n12509 ;
  assign n12511 = n5947 & ~n12510 ;
  assign n12512 = n2356 & ~n2360 ;
  assign n12513 = n12512 ^ n413 ^ 1'b0 ;
  assign n12514 = n12513 ^ n9306 ^ n8680 ;
  assign n12515 = n4135 & ~n12311 ;
  assign n12516 = n4758 ^ n3976 ^ n2306 ;
  assign n12517 = n5625 & ~n8886 ;
  assign n12518 = n12253 & ~n12517 ;
  assign n12519 = n12516 & n12518 ;
  assign n12520 = n4256 & n5477 ;
  assign n12521 = ~n6751 & n12520 ;
  assign n12522 = ( n7791 & n12379 ) | ( n7791 & ~n12521 ) | ( n12379 & ~n12521 ) ;
  assign n12523 = n11545 ^ n3374 ^ n378 ;
  assign n12524 = n6842 ^ n6819 ^ x24 ;
  assign n12529 = n9872 ^ n6183 ^ n5111 ;
  assign n12530 = ( n5786 & n9197 ) | ( n5786 & ~n12529 ) | ( n9197 & ~n12529 ) ;
  assign n12525 = ~n311 & n5319 ;
  assign n12526 = ~n4927 & n12525 ;
  assign n12527 = n5319 & ~n12526 ;
  assign n12528 = n7030 & n12527 ;
  assign n12531 = n12530 ^ n12528 ^ n4236 ;
  assign n12532 = n8658 & n11049 ;
  assign n12533 = n9840 & n12532 ;
  assign n12534 = ( ~n1019 & n1624 ) | ( ~n1019 & n12533 ) | ( n1624 & n12533 ) ;
  assign n12535 = n12534 ^ n9738 ^ n3294 ;
  assign n12541 = ( n5862 & ~n5912 ) | ( n5862 & n6303 ) | ( ~n5912 & n6303 ) ;
  assign n12540 = n11141 ^ n10809 ^ 1'b0 ;
  assign n12536 = n4726 & n5545 ;
  assign n12537 = ~n1817 & n12536 ;
  assign n12538 = ( n703 & ~n7562 ) | ( n703 & n12537 ) | ( ~n7562 & n12537 ) ;
  assign n12539 = ( ~n7994 & n9071 ) | ( ~n7994 & n12538 ) | ( n9071 & n12538 ) ;
  assign n12542 = n12541 ^ n12540 ^ n12539 ;
  assign n12543 = n8779 ^ n6703 ^ n4474 ;
  assign n12544 = n12543 ^ n1145 ^ 1'b0 ;
  assign n12545 = ~n1572 & n12544 ;
  assign n12546 = ( ~n3453 & n8465 ) | ( ~n3453 & n11510 ) | ( n8465 & n11510 ) ;
  assign n12547 = n12546 ^ n2424 ^ n642 ;
  assign n12548 = n12547 ^ n12008 ^ n6966 ;
  assign n12549 = n1860 | n4172 ;
  assign n12550 = n12549 ^ n3659 ^ 1'b0 ;
  assign n12551 = n4981 & ~n12550 ;
  assign n12552 = ~n2267 & n7720 ;
  assign n12553 = ~n12465 & n12552 ;
  assign n12554 = n10661 | n12553 ;
  assign n12555 = ( n5542 & n11830 ) | ( n5542 & n12554 ) | ( n11830 & n12554 ) ;
  assign n12556 = ~n6545 & n12059 ;
  assign n12557 = ~n12555 & n12556 ;
  assign n12558 = n3814 | n12557 ;
  assign n12559 = n12558 ^ n10909 ^ 1'b0 ;
  assign n12560 = n2919 | n11683 ;
  assign n12561 = n12560 ^ n5059 ^ 1'b0 ;
  assign n12562 = ( n2236 & n10327 ) | ( n2236 & ~n12561 ) | ( n10327 & ~n12561 ) ;
  assign n12564 = ~n1992 & n4472 ;
  assign n12565 = n12564 ^ n3678 ^ 1'b0 ;
  assign n12563 = n9193 ^ n7056 ^ n1344 ;
  assign n12566 = n12565 ^ n12563 ^ 1'b0 ;
  assign n12567 = n5900 & ~n8653 ;
  assign n12568 = n6047 ^ n5749 ^ n4723 ;
  assign n12569 = n9518 | n12568 ;
  assign n12570 = n453 ^ n244 ^ 1'b0 ;
  assign n12571 = n886 & ~n12570 ;
  assign n12572 = n12571 ^ n12222 ^ 1'b0 ;
  assign n12573 = n11063 | n12572 ;
  assign n12574 = ( n3995 & n5115 ) | ( n3995 & ~n12573 ) | ( n5115 & ~n12573 ) ;
  assign n12575 = ~n9146 & n12574 ;
  assign n12576 = ~n5220 & n9108 ;
  assign n12578 = n1655 ^ n1105 ^ 1'b0 ;
  assign n12579 = ( n2432 & ~n3909 ) | ( n2432 & n12578 ) | ( ~n3909 & n12578 ) ;
  assign n12577 = ( n581 & n2397 ) | ( n581 & ~n6874 ) | ( n2397 & ~n6874 ) ;
  assign n12580 = n12579 ^ n12577 ^ 1'b0 ;
  assign n12581 = ( n7918 & n12576 ) | ( n7918 & n12580 ) | ( n12576 & n12580 ) ;
  assign n12582 = n11995 ^ n8078 ^ 1'b0 ;
  assign n12583 = n5554 | n6820 ;
  assign n12584 = n5250 ^ n2745 ^ 1'b0 ;
  assign n12585 = n2338 & n12584 ;
  assign n12586 = n3856 ^ n931 ^ 1'b0 ;
  assign n12587 = n12229 ^ n9394 ^ n5023 ;
  assign n12588 = ( n12585 & ~n12586 ) | ( n12585 & n12587 ) | ( ~n12586 & n12587 ) ;
  assign n12594 = n1336 & n11222 ;
  assign n12595 = ( n6446 & n8398 ) | ( n6446 & n12594 ) | ( n8398 & n12594 ) ;
  assign n12589 = n1270 & n3018 ;
  assign n12590 = n12589 ^ n1982 ^ 1'b0 ;
  assign n12591 = n9659 & ~n12590 ;
  assign n12592 = n12591 ^ n3007 ^ 1'b0 ;
  assign n12593 = n7981 & n12592 ;
  assign n12596 = n12595 ^ n12593 ^ 1'b0 ;
  assign n12597 = ( n866 & n5218 ) | ( n866 & ~n8725 ) | ( n5218 & ~n8725 ) ;
  assign n12598 = n1393 ^ n1132 ^ 1'b0 ;
  assign n12599 = ~n2247 & n12598 ;
  assign n12600 = n12599 ^ n943 ^ 1'b0 ;
  assign n12601 = n1474 & n3603 ;
  assign n12602 = n5068 & n12601 ;
  assign n12603 = ( n1088 & n5957 ) | ( n1088 & ~n12602 ) | ( n5957 & ~n12602 ) ;
  assign n12604 = n1358 | n9850 ;
  assign n12605 = n6415 & ~n12604 ;
  assign n12606 = n12605 ^ n10963 ^ n8235 ;
  assign n12607 = n1018 & n3826 ;
  assign n12608 = n12607 ^ n2308 ^ n2267 ;
  assign n12609 = ~n11846 & n12608 ;
  assign n12610 = n11408 & n12609 ;
  assign n12611 = n12610 ^ n6524 ^ 1'b0 ;
  assign n12612 = ~n2593 & n12611 ;
  assign n12613 = n10983 & n12612 ;
  assign n12614 = ~n3548 & n12613 ;
  assign n12615 = n1832 ^ n598 ^ 1'b0 ;
  assign n12616 = n9659 & ~n12615 ;
  assign n12617 = n760 & n4356 ;
  assign n12618 = n12617 ^ x118 ^ 1'b0 ;
  assign n12619 = n12618 ^ n6371 ^ 1'b0 ;
  assign n12620 = n12616 & ~n12619 ;
  assign n12621 = n10772 ^ n9543 ^ 1'b0 ;
  assign n12622 = n4347 ^ n401 ^ n286 ;
  assign n12623 = ~n6490 & n9975 ;
  assign n12624 = n9479 & n12623 ;
  assign n12625 = n5971 & n12624 ;
  assign n12626 = n8528 ^ n572 ^ 1'b0 ;
  assign n12627 = n2600 | n12005 ;
  assign n12628 = n6442 & ~n12627 ;
  assign n12629 = n11501 | n12628 ;
  assign n12630 = n12629 ^ n8074 ^ 1'b0 ;
  assign n12631 = ( n5446 & n12626 ) | ( n5446 & n12630 ) | ( n12626 & n12630 ) ;
  assign n12632 = x17 & ~n7478 ;
  assign n12633 = ( ~n6286 & n10703 ) | ( ~n6286 & n12632 ) | ( n10703 & n12632 ) ;
  assign n12634 = ( n11358 & n12008 ) | ( n11358 & ~n12633 ) | ( n12008 & ~n12633 ) ;
  assign n12635 = ~n6644 & n6710 ;
  assign n12636 = n12635 ^ n6706 ^ 1'b0 ;
  assign n12637 = n12636 ^ n8545 ^ n7482 ;
  assign n12638 = n12637 ^ n4479 ^ 1'b0 ;
  assign n12639 = ( ~n12353 & n12634 ) | ( ~n12353 & n12638 ) | ( n12634 & n12638 ) ;
  assign n12640 = n11204 ^ n9110 ^ n6185 ;
  assign n12641 = n12640 ^ n6972 ^ n1749 ;
  assign n12642 = n8833 ^ n1942 ^ 1'b0 ;
  assign n12645 = ( ~n2869 & n4902 ) | ( ~n2869 & n5409 ) | ( n4902 & n5409 ) ;
  assign n12643 = n956 ^ n503 ^ 1'b0 ;
  assign n12644 = n8072 | n12643 ;
  assign n12646 = n12645 ^ n12644 ^ 1'b0 ;
  assign n12647 = n10099 & ~n12646 ;
  assign n12648 = ~n3761 & n10917 ;
  assign n12649 = n12648 ^ n2413 ^ 1'b0 ;
  assign n12650 = n1859 & n12649 ;
  assign n12651 = n142 | n3610 ;
  assign n12652 = n2277 | n12651 ;
  assign n12653 = n12652 ^ n249 ^ 1'b0 ;
  assign n12654 = n8184 & n9647 ;
  assign n12655 = ( n2436 & n12653 ) | ( n2436 & n12654 ) | ( n12653 & n12654 ) ;
  assign n12660 = n5552 ^ n4542 ^ 1'b0 ;
  assign n12661 = n8103 & ~n12660 ;
  assign n12657 = n2969 & n3543 ;
  assign n12658 = ~n7800 & n12657 ;
  assign n12656 = ~n223 & n5216 ;
  assign n12659 = n12658 ^ n12656 ^ n8435 ;
  assign n12662 = n12661 ^ n12659 ^ n6519 ;
  assign n12663 = n4973 ^ n2423 ^ n639 ;
  assign n12664 = n3586 ^ n2807 ^ n1108 ;
  assign n12665 = ( n6204 & n12663 ) | ( n6204 & ~n12664 ) | ( n12663 & ~n12664 ) ;
  assign n12678 = n3989 & n7994 ;
  assign n12679 = ~n5491 & n12678 ;
  assign n12673 = n2704 & n7811 ;
  assign n12674 = ~n7675 & n12673 ;
  assign n12668 = x19 | n148 ;
  assign n12669 = n1368 ^ n665 ^ 1'b0 ;
  assign n12670 = n3687 & n12669 ;
  assign n12671 = n9220 & n12670 ;
  assign n12672 = n12668 & ~n12671 ;
  assign n12675 = n12674 ^ n12672 ^ 1'b0 ;
  assign n12676 = n6905 & n12675 ;
  assign n12677 = n12676 ^ n6335 ^ 1'b0 ;
  assign n12680 = n12679 ^ n12677 ^ 1'b0 ;
  assign n12681 = n12680 ^ n4678 ^ x89 ;
  assign n12666 = n3295 & ~n6359 ;
  assign n12667 = n7568 | n12666 ;
  assign n12682 = n12681 ^ n12667 ^ 1'b0 ;
  assign n12683 = ( ~n1909 & n2880 ) | ( ~n1909 & n9507 ) | ( n2880 & n9507 ) ;
  assign n12684 = n7011 ^ n6446 ^ n2822 ;
  assign n12685 = n3743 | n7388 ;
  assign n12686 = n12685 ^ n8234 ^ 1'b0 ;
  assign n12687 = n10737 & n12686 ;
  assign n12688 = ~n12684 & n12687 ;
  assign n12689 = n207 & ~n8950 ;
  assign n12690 = n5723 & n12689 ;
  assign n12691 = n5540 & ~n12690 ;
  assign n12692 = n7848 ^ n6815 ^ n2107 ;
  assign n12693 = n12692 ^ n1247 ^ 1'b0 ;
  assign n12694 = n12693 ^ n12225 ^ 1'b0 ;
  assign n12695 = n6970 ^ n6949 ^ 1'b0 ;
  assign n12697 = ~n1228 & n6881 ;
  assign n12696 = ~n1716 & n4496 ;
  assign n12698 = n12697 ^ n12696 ^ 1'b0 ;
  assign n12699 = n4522 & ~n11564 ;
  assign n12700 = ~n182 & n12699 ;
  assign n12701 = ( n1501 & ~n6626 ) | ( n1501 & n12700 ) | ( ~n6626 & n12700 ) ;
  assign n12702 = n12701 ^ n8770 ^ 1'b0 ;
  assign n12705 = n6013 ^ n4133 ^ 1'b0 ;
  assign n12706 = n9206 | n12705 ;
  assign n12703 = n12495 ^ n1717 ^ 1'b0 ;
  assign n12704 = n2828 & ~n12703 ;
  assign n12707 = n12706 ^ n12704 ^ n12181 ;
  assign n12708 = n5227 & ~n12707 ;
  assign n12715 = n2876 ^ n2138 ^ n886 ;
  assign n12709 = ~n1315 & n5639 ;
  assign n12710 = ~n6453 & n12709 ;
  assign n12711 = ( ~n3314 & n3916 ) | ( ~n3314 & n4412 ) | ( n3916 & n4412 ) ;
  assign n12712 = ( n223 & n3214 ) | ( n223 & n12711 ) | ( n3214 & n12711 ) ;
  assign n12713 = n12712 ^ n5425 ^ n5224 ;
  assign n12714 = ~n12710 & n12713 ;
  assign n12716 = n12715 ^ n12714 ^ n2797 ;
  assign n12717 = n9079 ^ n5283 ^ 1'b0 ;
  assign n12718 = ( ~n3993 & n4438 ) | ( ~n3993 & n7054 ) | ( n4438 & n7054 ) ;
  assign n12719 = n2705 | n12718 ;
  assign n12720 = n12719 ^ n3543 ^ 1'b0 ;
  assign n12721 = n9031 ^ n3854 ^ 1'b0 ;
  assign n12722 = n10268 ^ n462 ^ 1'b0 ;
  assign n12723 = n3339 & n3387 ;
  assign n12724 = n12723 ^ n2839 ^ 1'b0 ;
  assign n12725 = n12722 | n12724 ;
  assign n12726 = n12725 ^ n6584 ^ 1'b0 ;
  assign n12727 = n3280 | n12726 ;
  assign n12730 = n3480 ^ n2884 ^ n1800 ;
  assign n12728 = ~n1085 & n10469 ;
  assign n12729 = ( n2794 & ~n8261 ) | ( n2794 & n12728 ) | ( ~n8261 & n12728 ) ;
  assign n12731 = n12730 ^ n12729 ^ n8625 ;
  assign n12732 = n8686 ^ n3054 ^ n2970 ;
  assign n12733 = n12732 ^ n9440 ^ 1'b0 ;
  assign n12734 = ~n12731 & n12733 ;
  assign n12735 = n6671 & ~n12534 ;
  assign n12736 = n9325 ^ n7589 ^ 1'b0 ;
  assign n12737 = ( n4366 & n6827 ) | ( n4366 & ~n12736 ) | ( n6827 & ~n12736 ) ;
  assign n12738 = n10335 ^ n5200 ^ n1518 ;
  assign n12739 = ( ~n2496 & n6123 ) | ( ~n2496 & n12738 ) | ( n6123 & n12738 ) ;
  assign n12740 = n6532 | n12739 ;
  assign n12741 = n12740 ^ x48 ^ 1'b0 ;
  assign n12742 = n8483 & ~n9352 ;
  assign n12743 = n6450 ^ n5479 ^ n414 ;
  assign n12744 = n12743 ^ n10999 ^ n7333 ;
  assign n12745 = ( n2091 & ~n8162 ) | ( n2091 & n8599 ) | ( ~n8162 & n8599 ) ;
  assign n12746 = n12745 ^ n5005 ^ 1'b0 ;
  assign n12747 = n1674 ^ n981 ^ 1'b0 ;
  assign n12748 = n9286 ^ n2959 ^ 1'b0 ;
  assign n12749 = ( n12746 & ~n12747 ) | ( n12746 & n12748 ) | ( ~n12747 & n12748 ) ;
  assign n12750 = ( n356 & ~n927 ) | ( n356 & n3103 ) | ( ~n927 & n3103 ) ;
  assign n12751 = ~n9631 & n12750 ;
  assign n12752 = n8611 & n12751 ;
  assign n12753 = n10586 ^ n6243 ^ 1'b0 ;
  assign n12754 = n11370 & ~n12753 ;
  assign n12755 = ( ~n1063 & n3339 ) | ( ~n1063 & n7954 ) | ( n3339 & n7954 ) ;
  assign n12756 = n6501 | n12755 ;
  assign n12757 = n2873 & ~n5103 ;
  assign n12758 = n11975 ^ n10963 ^ n7408 ;
  assign n12759 = n12757 | n12758 ;
  assign n12761 = n1896 ^ n599 ^ 1'b0 ;
  assign n12762 = n330 & n12761 ;
  assign n12760 = n2038 | n3785 ;
  assign n12763 = n12762 ^ n12760 ^ 1'b0 ;
  assign n12764 = ~n1346 & n12763 ;
  assign n12765 = ~n7042 & n12764 ;
  assign n12766 = n12765 ^ n2232 ^ 1'b0 ;
  assign n12767 = n1566 ^ n884 ^ 1'b0 ;
  assign n12768 = n9823 ^ n7848 ^ 1'b0 ;
  assign n12769 = n12768 ^ n1095 ^ 1'b0 ;
  assign n12770 = n8529 ^ n3227 ^ n1635 ;
  assign n12771 = ( ~n1836 & n3608 ) | ( ~n1836 & n3702 ) | ( n3608 & n3702 ) ;
  assign n12772 = n8559 ^ n7724 ^ n7662 ;
  assign n12773 = n6102 ^ n4000 ^ 1'b0 ;
  assign n12774 = x96 & ~n12773 ;
  assign n12775 = n12772 & n12774 ;
  assign n12776 = n12775 ^ n1227 ^ 1'b0 ;
  assign n12777 = ( ~n10424 & n12771 ) | ( ~n10424 & n12776 ) | ( n12771 & n12776 ) ;
  assign n12778 = ( n2798 & n6433 ) | ( n2798 & ~n9336 ) | ( n6433 & ~n9336 ) ;
  assign n12779 = n12778 ^ n8403 ^ n3798 ;
  assign n12780 = n9640 ^ n8596 ^ 1'b0 ;
  assign n12781 = ( n1809 & ~n6543 ) | ( n1809 & n7436 ) | ( ~n6543 & n7436 ) ;
  assign n12783 = n6300 & n11524 ;
  assign n12784 = ~n1654 & n12783 ;
  assign n12782 = n4691 & n6686 ;
  assign n12785 = n12784 ^ n12782 ^ 1'b0 ;
  assign n12786 = n12785 ^ n9146 ^ 1'b0 ;
  assign n12787 = n12781 & ~n12786 ;
  assign n12788 = n1651 | n7757 ;
  assign n12789 = n12788 ^ n10256 ^ 1'b0 ;
  assign n12790 = n12789 ^ n1943 ^ 1'b0 ;
  assign n12791 = n11988 ^ n5847 ^ n4702 ;
  assign n12792 = n815 | n12791 ;
  assign n12793 = ( n599 & n896 ) | ( n599 & ~n11676 ) | ( n896 & ~n11676 ) ;
  assign n12794 = n12793 ^ n9562 ^ n5861 ;
  assign n12795 = ~n214 & n12794 ;
  assign n12796 = ~n12792 & n12795 ;
  assign n12797 = ( n444 & n11378 ) | ( n444 & ~n12796 ) | ( n11378 & ~n12796 ) ;
  assign n12798 = ( ~n5634 & n6349 ) | ( ~n5634 & n10096 ) | ( n6349 & n10096 ) ;
  assign n12799 = n11317 & ~n12798 ;
  assign n12800 = ~n600 & n1199 ;
  assign n12801 = n11727 & n12800 ;
  assign n12802 = ( ~n4953 & n7596 ) | ( ~n4953 & n7891 ) | ( n7596 & n7891 ) ;
  assign n12803 = ~n4281 & n5679 ;
  assign n12804 = n12803 ^ n11799 ^ 1'b0 ;
  assign n12805 = n12804 ^ n8326 ^ 1'b0 ;
  assign n12806 = n12802 & n12805 ;
  assign n12807 = n7874 ^ n3930 ^ 1'b0 ;
  assign n12808 = n5635 ^ n2643 ^ 1'b0 ;
  assign n12809 = n6663 & n7722 ;
  assign n12810 = ~n526 & n12809 ;
  assign n12811 = ( ~x116 & n8653 ) | ( ~x116 & n9856 ) | ( n8653 & n9856 ) ;
  assign n12812 = n12811 ^ n10663 ^ 1'b0 ;
  assign n12813 = n722 & ~n12812 ;
  assign n12814 = n10070 & ~n10284 ;
  assign n12815 = n12814 ^ n7818 ^ 1'b0 ;
  assign n12816 = ( ~n5442 & n6002 ) | ( ~n5442 & n7288 ) | ( n6002 & n7288 ) ;
  assign n12817 = n12816 ^ n12397 ^ n10413 ;
  assign n12820 = n3048 ^ n785 ^ 1'b0 ;
  assign n12818 = ( n2216 & n4048 ) | ( n2216 & ~n9553 ) | ( n4048 & ~n9553 ) ;
  assign n12819 = ( n6737 & n10565 ) | ( n6737 & n12818 ) | ( n10565 & n12818 ) ;
  assign n12821 = n12820 ^ n12819 ^ n11412 ;
  assign n12822 = ~n3252 & n6838 ;
  assign n12823 = n10114 & ~n12822 ;
  assign n12824 = n9798 & n12823 ;
  assign n12825 = ( n1376 & ~n3529 ) | ( n1376 & n9920 ) | ( ~n3529 & n9920 ) ;
  assign n12826 = n9697 ^ n3153 ^ 1'b0 ;
  assign n12827 = ( n177 & n207 ) | ( n177 & ~n3249 ) | ( n207 & ~n3249 ) ;
  assign n12828 = n12826 & ~n12827 ;
  assign n12829 = n6445 ^ n5312 ^ n4320 ;
  assign n12830 = ( n1102 & n1456 ) | ( n1102 & n12829 ) | ( n1456 & n12829 ) ;
  assign n12831 = n9964 ^ n9534 ^ n8261 ;
  assign n12832 = ( n5554 & n9067 ) | ( n5554 & n9929 ) | ( n9067 & n9929 ) ;
  assign n12833 = n3177 & n12245 ;
  assign n12834 = n12638 ^ n4879 ^ n167 ;
  assign n12835 = n2835 & n5329 ;
  assign n12836 = n12835 ^ n6013 ^ 1'b0 ;
  assign n12837 = n709 | n2183 ;
  assign n12838 = n5145 & ~n12837 ;
  assign n12839 = ( n4545 & n8465 ) | ( n4545 & n12838 ) | ( n8465 & n12838 ) ;
  assign n12840 = ~n12836 & n12839 ;
  assign n12841 = n1326 | n12706 ;
  assign n12845 = n9515 ^ n2612 ^ n373 ;
  assign n12842 = n300 | n2587 ;
  assign n12843 = n12842 ^ n3106 ^ 1'b0 ;
  assign n12844 = n3110 & n12843 ;
  assign n12846 = n12845 ^ n12844 ^ n7648 ;
  assign n12847 = n1370 & n9087 ;
  assign n12848 = n2648 ^ n2159 ^ 1'b0 ;
  assign n12849 = n12848 ^ n7758 ^ 1'b0 ;
  assign n12850 = n2241 | n12849 ;
  assign n12851 = n12847 & ~n12850 ;
  assign n12852 = n11289 ^ n3020 ^ 1'b0 ;
  assign n12853 = n1621 | n11932 ;
  assign n12854 = n12853 ^ n168 ^ 1'b0 ;
  assign n12855 = ( ~n2544 & n4088 ) | ( ~n2544 & n12854 ) | ( n4088 & n12854 ) ;
  assign n12856 = n298 & n4987 ;
  assign n12857 = n2103 ^ n1174 ^ 1'b0 ;
  assign n12858 = ~n1401 & n12857 ;
  assign n12859 = n12858 ^ n3354 ^ 1'b0 ;
  assign n12860 = n12859 ^ n2491 ^ n2288 ;
  assign n12861 = n12822 ^ n12731 ^ n6334 ;
  assign n12862 = ( n12856 & n12860 ) | ( n12856 & n12861 ) | ( n12860 & n12861 ) ;
  assign n12863 = ( ~n478 & n1532 ) | ( ~n478 & n3723 ) | ( n1532 & n3723 ) ;
  assign n12864 = n2820 | n6836 ;
  assign n12865 = n3265 | n12864 ;
  assign n12866 = n5345 & ~n9116 ;
  assign n12867 = n12866 ^ n1046 ^ 1'b0 ;
  assign n12868 = ~n12865 & n12867 ;
  assign n12873 = ( x114 & n1719 ) | ( x114 & ~n5105 ) | ( n1719 & ~n5105 ) ;
  assign n12874 = n12873 ^ n6735 ^ 1'b0 ;
  assign n12875 = ~n11273 & n12874 ;
  assign n12869 = n705 & n3064 ;
  assign n12870 = ~x76 & n12869 ;
  assign n12871 = n5306 & n8378 ;
  assign n12872 = ( ~n483 & n12870 ) | ( ~n483 & n12871 ) | ( n12870 & n12871 ) ;
  assign n12876 = n12875 ^ n12872 ^ 1'b0 ;
  assign n12877 = ( n3111 & n5036 ) | ( n3111 & ~n9332 ) | ( n5036 & ~n9332 ) ;
  assign n12878 = n12877 ^ n2950 ^ 1'b0 ;
  assign n12879 = n199 & n9205 ;
  assign n12880 = ~n3254 & n12879 ;
  assign n12881 = n12880 ^ n4375 ^ 1'b0 ;
  assign n12882 = n8460 ^ n6156 ^ 1'b0 ;
  assign n12883 = n5207 ^ n4488 ^ 1'b0 ;
  assign n12884 = n5058 | n12883 ;
  assign n12885 = n12884 ^ n10325 ^ 1'b0 ;
  assign n12886 = n8126 ^ n7790 ^ n3891 ;
  assign n12887 = n10589 ^ n4084 ^ 1'b0 ;
  assign n12888 = ( n4152 & n12068 ) | ( n4152 & ~n12887 ) | ( n12068 & ~n12887 ) ;
  assign n12889 = n12888 ^ n10472 ^ 1'b0 ;
  assign n12890 = n12889 ^ n3947 ^ n1929 ;
  assign n12891 = n1237 & ~n8738 ;
  assign n12892 = ( n1020 & n2889 ) | ( n1020 & ~n12891 ) | ( n2889 & ~n12891 ) ;
  assign n12893 = n5604 ^ n3841 ^ 1'b0 ;
  assign n12894 = ~n1813 & n3899 ;
  assign n12895 = n12894 ^ n4217 ^ 1'b0 ;
  assign n12896 = n12895 ^ n1279 ^ 1'b0 ;
  assign n12897 = n5867 | n12896 ;
  assign n12898 = ( ~n3799 & n12893 ) | ( ~n3799 & n12897 ) | ( n12893 & n12897 ) ;
  assign n12899 = n12892 | n12898 ;
  assign n12900 = n12890 | n12899 ;
  assign n12901 = n4727 ^ n3282 ^ 1'b0 ;
  assign n12902 = ( ~n204 & n464 ) | ( ~n204 & n2577 ) | ( n464 & n2577 ) ;
  assign n12903 = n12902 ^ n11393 ^ n1175 ;
  assign n12904 = n12903 ^ n3839 ^ 1'b0 ;
  assign n12905 = n6805 & n12904 ;
  assign n12906 = n12905 ^ n10434 ^ 1'b0 ;
  assign n12908 = n2661 & ~n11932 ;
  assign n12909 = n12908 ^ n2962 ^ 1'b0 ;
  assign n12910 = n12909 ^ n5047 ^ 1'b0 ;
  assign n12911 = n1115 | n12910 ;
  assign n12912 = n12911 ^ n9473 ^ 1'b0 ;
  assign n12907 = n1873 | n5723 ;
  assign n12913 = n12912 ^ n12907 ^ n7328 ;
  assign n12915 = n3984 & n11086 ;
  assign n12914 = n8093 ^ n4458 ^ n2776 ;
  assign n12916 = n12915 ^ n12914 ^ n2910 ;
  assign n12917 = ~n4501 & n12916 ;
  assign n12918 = n12917 ^ n2445 ^ 1'b0 ;
  assign n12919 = n5195 ^ n4612 ^ n450 ;
  assign n12920 = n3531 & ~n6624 ;
  assign n12921 = ~n12919 & n12920 ;
  assign n12922 = n9812 ^ n6238 ^ n5164 ;
  assign n12923 = n9193 ^ n6710 ^ n4372 ;
  assign n12924 = n12791 ^ n5669 ^ n3713 ;
  assign n12928 = ( n7703 & ~n8550 ) | ( n7703 & n10754 ) | ( ~n8550 & n10754 ) ;
  assign n12925 = n4852 | n11620 ;
  assign n12926 = n2530 | n12925 ;
  assign n12927 = ( n878 & n9630 ) | ( n878 & ~n12926 ) | ( n9630 & ~n12926 ) ;
  assign n12929 = n12928 ^ n12927 ^ 1'b0 ;
  assign n12930 = n12924 & n12929 ;
  assign n12933 = n11799 ^ n698 ^ 1'b0 ;
  assign n12934 = n8875 & ~n12933 ;
  assign n12931 = ( ~n4528 & n6128 ) | ( ~n4528 & n8441 ) | ( n6128 & n8441 ) ;
  assign n12932 = n12931 ^ n8703 ^ n5349 ;
  assign n12935 = n12934 ^ n12932 ^ n4040 ;
  assign n12936 = ~n7205 & n9165 ;
  assign n12937 = n12935 & n12936 ;
  assign n12938 = n1729 | n8625 ;
  assign n12939 = n5382 | n12938 ;
  assign n12940 = n6006 & ~n12939 ;
  assign n12941 = n12005 | n12940 ;
  assign n12942 = n12941 ^ n8341 ^ 1'b0 ;
  assign n12943 = n3742 & ~n12942 ;
  assign n12944 = n12943 ^ n5587 ^ 1'b0 ;
  assign n12945 = n12944 ^ n7241 ^ n1902 ;
  assign n12946 = n6320 ^ n2794 ^ 1'b0 ;
  assign n12947 = x114 & ~n12946 ;
  assign n12948 = n12947 ^ n1532 ^ 1'b0 ;
  assign n12949 = n12948 ^ n2149 ^ 1'b0 ;
  assign n12950 = ~n2107 & n3150 ;
  assign n12953 = n1411 & n12778 ;
  assign n12954 = ~n2436 & n12953 ;
  assign n12955 = n12954 ^ n598 ^ 1'b0 ;
  assign n12951 = n3242 & ~n4108 ;
  assign n12952 = n12951 ^ n5650 ^ 1'b0 ;
  assign n12956 = n12955 ^ n12952 ^ n11453 ;
  assign n12957 = n12412 ^ n5865 ^ n5288 ;
  assign n12958 = n10994 ^ n10480 ^ n3078 ;
  assign n12959 = n3075 & n12958 ;
  assign n12960 = ( n6605 & ~n7460 ) | ( n6605 & n12819 ) | ( ~n7460 & n12819 ) ;
  assign n12961 = n9104 ^ n3115 ^ n2025 ;
  assign n12962 = n12961 ^ n9297 ^ x29 ;
  assign n12963 = n6075 ^ n201 ^ 1'b0 ;
  assign n12964 = n12962 | n12963 ;
  assign n12965 = n7575 & ~n12964 ;
  assign n12966 = n12275 & n12965 ;
  assign n12967 = n12966 ^ n2346 ^ 1'b0 ;
  assign n12968 = n12960 & n12967 ;
  assign n12969 = ( n2027 & n2648 ) | ( n2027 & ~n10979 ) | ( n2648 & ~n10979 ) ;
  assign n12978 = n8783 ^ n8497 ^ n8129 ;
  assign n12979 = n12978 ^ n4254 ^ 1'b0 ;
  assign n12980 = n2757 & ~n12979 ;
  assign n12981 = n12980 ^ n8933 ^ n2016 ;
  assign n12970 = ( ~n1403 & n3046 ) | ( ~n1403 & n6239 ) | ( n3046 & n6239 ) ;
  assign n12971 = n12970 ^ n5921 ^ n1777 ;
  assign n12972 = n3085 ^ n2203 ^ 1'b0 ;
  assign n12973 = n6377 ^ n2689 ^ n1553 ;
  assign n12974 = n11435 & n12973 ;
  assign n12975 = ~n1074 & n12974 ;
  assign n12976 = n12972 | n12975 ;
  assign n12977 = n12971 & ~n12976 ;
  assign n12982 = n12981 ^ n12977 ^ n815 ;
  assign n12983 = ( n695 & n12969 ) | ( n695 & n12982 ) | ( n12969 & n12982 ) ;
  assign n12990 = ~n2579 & n9157 ;
  assign n12984 = n557 | n2848 ;
  assign n12985 = ~n3769 & n8455 ;
  assign n12986 = ~n11565 & n12985 ;
  assign n12987 = ( n2749 & n12984 ) | ( n2749 & n12986 ) | ( n12984 & n12986 ) ;
  assign n12988 = n7792 ^ n757 ^ 1'b0 ;
  assign n12989 = ( n2681 & n12987 ) | ( n2681 & ~n12988 ) | ( n12987 & ~n12988 ) ;
  assign n12991 = n12990 ^ n12989 ^ n10937 ;
  assign n12992 = n3754 ^ n2830 ^ n767 ;
  assign n12993 = ( n3838 & n4108 ) | ( n3838 & n12992 ) | ( n4108 & n12992 ) ;
  assign n12994 = ~n1295 & n8812 ;
  assign n12995 = n10913 & n12994 ;
  assign n12996 = ( n6116 & ~n9795 ) | ( n6116 & n12562 ) | ( ~n9795 & n12562 ) ;
  assign n12997 = n12996 ^ n8923 ^ n5302 ;
  assign n12998 = ( n4149 & n4918 ) | ( n4149 & ~n5460 ) | ( n4918 & ~n5460 ) ;
  assign n12999 = n5743 ^ n3697 ^ 1'b0 ;
  assign n13000 = ~n12998 & n12999 ;
  assign n13001 = ~n6522 & n10742 ;
  assign n13002 = n459 & n13001 ;
  assign n13003 = n6872 | n10401 ;
  assign n13004 = n8529 & ~n13003 ;
  assign n13005 = ~n6999 & n13004 ;
  assign n13006 = ( n6106 & n13002 ) | ( n6106 & ~n13005 ) | ( n13002 & ~n13005 ) ;
  assign n13007 = n13006 ^ n9081 ^ n8375 ;
  assign n13008 = ( n2934 & n3551 ) | ( n2934 & n6155 ) | ( n3551 & n6155 ) ;
  assign n13009 = ~n2981 & n13008 ;
  assign n13010 = ( n7667 & n7932 ) | ( n7667 & ~n8703 ) | ( n7932 & ~n8703 ) ;
  assign n13011 = ( n3138 & n6238 ) | ( n3138 & n13010 ) | ( n6238 & n13010 ) ;
  assign n13012 = n7065 & ~n10174 ;
  assign n13013 = n13004 ^ n2587 ^ 1'b0 ;
  assign n13014 = n13013 ^ n11718 ^ 1'b0 ;
  assign n13015 = ~n13012 & n13014 ;
  assign n13016 = ~n4196 & n6325 ;
  assign n13017 = n13016 ^ n11183 ^ 1'b0 ;
  assign n13018 = n7925 ^ n4546 ^ n853 ;
  assign n13019 = ~n4344 & n13018 ;
  assign n13020 = n13019 ^ n7173 ^ 1'b0 ;
  assign n13021 = ( n3971 & n13017 ) | ( n3971 & n13020 ) | ( n13017 & n13020 ) ;
  assign n13022 = ~n10131 & n13021 ;
  assign n13023 = n6010 & n13022 ;
  assign n13024 = n9352 ^ n4452 ^ 1'b0 ;
  assign n13025 = n11959 ^ n10006 ^ n8525 ;
  assign n13026 = n5829 & ~n7221 ;
  assign n13027 = n6723 ^ n5989 ^ n1486 ;
  assign n13028 = n13027 ^ n10397 ^ 1'b0 ;
  assign n13029 = n13026 | n13028 ;
  assign n13030 = ( x21 & n5108 ) | ( x21 & ~n7089 ) | ( n5108 & ~n7089 ) ;
  assign n13031 = n6243 ^ n6104 ^ n3485 ;
  assign n13032 = n4858 & ~n5756 ;
  assign n13034 = n3631 | n5685 ;
  assign n13035 = n7615 | n13034 ;
  assign n13036 = n7158 ^ n3919 ^ n1943 ;
  assign n13037 = n6908 & ~n13036 ;
  assign n13038 = ~n13035 & n13037 ;
  assign n13033 = n10011 | n10089 ;
  assign n13039 = n13038 ^ n13033 ^ 1'b0 ;
  assign n13041 = ( n3407 & n4674 ) | ( n3407 & n9953 ) | ( n4674 & n9953 ) ;
  assign n13040 = n10606 ^ n9159 ^ n4248 ;
  assign n13042 = n13041 ^ n13040 ^ n1126 ;
  assign n13043 = ~n4519 & n7208 ;
  assign n13044 = x65 & ~n5030 ;
  assign n13045 = ~n6747 & n13044 ;
  assign n13046 = n8658 ^ n6784 ^ n2135 ;
  assign n13048 = n4345 ^ n3631 ^ n2788 ;
  assign n13047 = n5356 & ~n7809 ;
  assign n13049 = n13048 ^ n13047 ^ 1'b0 ;
  assign n13050 = n4326 & n13049 ;
  assign n13051 = ( x30 & n7092 ) | ( x30 & n11394 ) | ( n7092 & n11394 ) ;
  assign n13052 = ( ~n13046 & n13050 ) | ( ~n13046 & n13051 ) | ( n13050 & n13051 ) ;
  assign n13053 = ( n1097 & ~n1629 ) | ( n1097 & n3922 ) | ( ~n1629 & n3922 ) ;
  assign n13054 = ( n4294 & ~n11746 ) | ( n4294 & n13053 ) | ( ~n11746 & n13053 ) ;
  assign n13055 = n1899 & ~n3439 ;
  assign n13056 = n5477 & n9448 ;
  assign n13057 = n13055 | n13056 ;
  assign n13058 = n13057 ^ n8349 ^ 1'b0 ;
  assign n13059 = ~n10174 & n13058 ;
  assign n13060 = n1833 | n5073 ;
  assign n13061 = ( n1455 & n5674 ) | ( n1455 & ~n6661 ) | ( n5674 & ~n6661 ) ;
  assign n13062 = ( n2253 & ~n4396 ) | ( n2253 & n6539 ) | ( ~n4396 & n6539 ) ;
  assign n13063 = n3730 & n13062 ;
  assign n13064 = ~n11400 & n13063 ;
  assign n13065 = ( n8685 & ~n13061 ) | ( n8685 & n13064 ) | ( ~n13061 & n13064 ) ;
  assign n13066 = n3346 ^ n808 ^ n454 ;
  assign n13070 = n4819 ^ n2949 ^ 1'b0 ;
  assign n13071 = n2346 | n13070 ;
  assign n13072 = n11143 & ~n13071 ;
  assign n13073 = n2638 | n10441 ;
  assign n13074 = ~n13072 & n13073 ;
  assign n13067 = n7437 ^ n6060 ^ 1'b0 ;
  assign n13068 = ~n2448 & n13067 ;
  assign n13069 = ( n1827 & n2726 ) | ( n1827 & ~n13068 ) | ( n2726 & ~n13068 ) ;
  assign n13075 = n13074 ^ n13069 ^ 1'b0 ;
  assign n13076 = n13066 & ~n13075 ;
  assign n13077 = n4837 | n8720 ;
  assign n13088 = n1818 | n4687 ;
  assign n13080 = ( n2692 & n4585 ) | ( n2692 & n9435 ) | ( n4585 & n9435 ) ;
  assign n13081 = n13080 ^ n3274 ^ 1'b0 ;
  assign n13082 = ( ~n680 & n10014 ) | ( ~n680 & n13081 ) | ( n10014 & n13081 ) ;
  assign n13083 = n13082 ^ n10949 ^ 1'b0 ;
  assign n13079 = n2812 ^ n956 ^ 1'b0 ;
  assign n13084 = n13083 ^ n13079 ^ n7591 ;
  assign n13085 = n13084 ^ n7082 ^ n6154 ;
  assign n13086 = n7787 & n13085 ;
  assign n13087 = n13086 ^ n9324 ^ 1'b0 ;
  assign n13078 = n5249 ^ n3147 ^ 1'b0 ;
  assign n13089 = n13088 ^ n13087 ^ n13078 ;
  assign n13090 = ( n2249 & ~n8239 ) | ( n2249 & n9814 ) | ( ~n8239 & n9814 ) ;
  assign n13091 = n7677 ^ n393 ^ 1'b0 ;
  assign n13092 = n2037 & ~n13091 ;
  assign n13093 = ( n620 & n5911 ) | ( n620 & ~n13092 ) | ( n5911 & ~n13092 ) ;
  assign n13094 = n13093 ^ n3487 ^ 1'b0 ;
  assign n13095 = n13090 & ~n13094 ;
  assign n13096 = n13095 ^ n3006 ^ n1159 ;
  assign n13097 = n3555 & n6312 ;
  assign n13098 = ( x33 & n2176 ) | ( x33 & n13097 ) | ( n2176 & n13097 ) ;
  assign n13099 = n12512 ^ n2393 ^ n2334 ;
  assign n13100 = ( n3586 & n11053 ) | ( n3586 & n13099 ) | ( n11053 & n13099 ) ;
  assign n13101 = n13100 ^ n12219 ^ n4534 ;
  assign n13102 = n12009 ^ n2303 ^ 1'b0 ;
  assign n13103 = n13102 ^ n7981 ^ n4215 ;
  assign n13104 = n2163 & ~n4989 ;
  assign n13105 = ( n618 & ~n1528 ) | ( n618 & n13104 ) | ( ~n1528 & n13104 ) ;
  assign n13106 = n6693 ^ n3851 ^ 1'b0 ;
  assign n13107 = n13105 | n13106 ;
  assign n13108 = n711 & n12029 ;
  assign n13109 = n7694 ^ n4084 ^ n4003 ;
  assign n13110 = n13109 ^ n10965 ^ 1'b0 ;
  assign n13111 = ( n13107 & n13108 ) | ( n13107 & ~n13110 ) | ( n13108 & ~n13110 ) ;
  assign n13112 = n3537 & ~n3666 ;
  assign n13113 = ( n1999 & ~n6085 ) | ( n1999 & n13112 ) | ( ~n6085 & n13112 ) ;
  assign n13114 = ( n5294 & n9774 ) | ( n5294 & ~n13113 ) | ( n9774 & ~n13113 ) ;
  assign n13119 = n2563 & ~n6101 ;
  assign n13120 = n7143 | n13119 ;
  assign n13121 = n13120 ^ n7604 ^ n881 ;
  assign n13115 = n12152 ^ n4069 ^ 1'b0 ;
  assign n13116 = n13008 & ~n13115 ;
  assign n13117 = ~n380 & n5671 ;
  assign n13118 = ~n13116 & n13117 ;
  assign n13122 = n13121 ^ n13118 ^ 1'b0 ;
  assign n13123 = n183 | n12098 ;
  assign n13124 = n6316 & n13054 ;
  assign n13125 = ~n9493 & n13124 ;
  assign n13126 = n4670 & ~n5214 ;
  assign n13127 = ~x116 & n13126 ;
  assign n13128 = n13127 ^ n5068 ^ n3263 ;
  assign n13129 = ~n6510 & n7091 ;
  assign n13130 = ~n7519 & n13129 ;
  assign n13131 = ~n13128 & n13130 ;
  assign n13132 = n12235 ^ n9538 ^ n1525 ;
  assign n13133 = n8481 ^ n1648 ^ 1'b0 ;
  assign n13134 = n13132 & ~n13133 ;
  assign n13135 = n13134 ^ n11618 ^ 1'b0 ;
  assign n13136 = n11807 | n13135 ;
  assign n13144 = n6789 & ~n8337 ;
  assign n13137 = ~n2349 & n5323 ;
  assign n13138 = n2206 & n5444 ;
  assign n13139 = n13138 ^ n1833 ^ 1'b0 ;
  assign n13140 = n7919 | n13139 ;
  assign n13141 = n10605 & ~n13140 ;
  assign n13142 = n3818 & ~n13141 ;
  assign n13143 = ~n13137 & n13142 ;
  assign n13145 = n13144 ^ n13143 ^ n3727 ;
  assign n13146 = n207 & ~n2709 ;
  assign n13147 = n13146 ^ n3364 ^ n2498 ;
  assign n13148 = n13147 ^ n6055 ^ 1'b0 ;
  assign n13149 = ( n1659 & ~n3981 ) | ( n1659 & n4008 ) | ( ~n3981 & n4008 ) ;
  assign n13150 = n5968 | n13149 ;
  assign n13151 = n13150 ^ n1739 ^ 1'b0 ;
  assign n13155 = n5526 ^ n3732 ^ n3595 ;
  assign n13152 = n4500 ^ n3033 ^ n1217 ;
  assign n13153 = n10166 & n13152 ;
  assign n13154 = n12436 | n13153 ;
  assign n13156 = n13155 ^ n13154 ^ 1'b0 ;
  assign n13157 = ~n4005 & n6596 ;
  assign n13158 = n11544 & n13157 ;
  assign n13159 = ( n6138 & n6376 ) | ( n6138 & ~n13158 ) | ( n6376 & ~n13158 ) ;
  assign n13163 = n2279 & n3482 ;
  assign n13164 = n13163 ^ n12009 ^ 1'b0 ;
  assign n13160 = n4198 | n8251 ;
  assign n13161 = n4130 & ~n13160 ;
  assign n13162 = n13161 ^ n2360 ^ 1'b0 ;
  assign n13165 = n13164 ^ n13162 ^ n2521 ;
  assign n13166 = n12344 ^ n10065 ^ n5951 ;
  assign n13171 = n5864 ^ n3471 ^ 1'b0 ;
  assign n13172 = n3530 | n13171 ;
  assign n13173 = n2131 | n13172 ;
  assign n13174 = n717 | n13173 ;
  assign n13169 = ( ~n2254 & n3252 ) | ( ~n2254 & n4391 ) | ( n3252 & n4391 ) ;
  assign n13170 = n13169 ^ n10697 ^ 1'b0 ;
  assign n13175 = n13174 ^ n13170 ^ n8615 ;
  assign n13167 = n3888 & ~n11016 ;
  assign n13168 = n13167 ^ n9287 ^ 1'b0 ;
  assign n13176 = n13175 ^ n13168 ^ n11633 ;
  assign n13177 = n9639 ^ n5622 ^ n268 ;
  assign n13178 = n13177 ^ n4772 ^ 1'b0 ;
  assign n13179 = n10057 ^ n8712 ^ 1'b0 ;
  assign n13180 = n13179 ^ n6162 ^ 1'b0 ;
  assign n13181 = ~n861 & n10915 ;
  assign n13182 = n7146 ^ n1429 ^ n660 ;
  assign n13183 = n13182 ^ n2502 ^ 1'b0 ;
  assign n13184 = n8973 | n13183 ;
  assign n13185 = ~n2914 & n4024 ;
  assign n13186 = n13185 ^ n6336 ^ n2197 ;
  assign n13187 = ( ~n4059 & n12534 ) | ( ~n4059 & n13186 ) | ( n12534 & n13186 ) ;
  assign n13188 = n6198 ^ n3216 ^ 1'b0 ;
  assign n13189 = n5134 & ~n13188 ;
  assign n13190 = n13189 ^ n7006 ^ n3048 ;
  assign n13191 = n3769 ^ n2371 ^ n2365 ;
  assign n13192 = n1994 & n5201 ;
  assign n13193 = n2526 & ~n9323 ;
  assign n13194 = n13192 & n13193 ;
  assign n13195 = ( ~n4233 & n5457 ) | ( ~n4233 & n13194 ) | ( n5457 & n13194 ) ;
  assign n13196 = n2138 & ~n9255 ;
  assign n13197 = n5913 ^ n5108 ^ n2604 ;
  assign n13198 = ( n1481 & ~n1946 ) | ( n1481 & n13197 ) | ( ~n1946 & n13197 ) ;
  assign n13199 = ( ~n1285 & n13196 ) | ( ~n1285 & n13198 ) | ( n13196 & n13198 ) ;
  assign n13200 = n11110 ^ n10205 ^ n2910 ;
  assign n13201 = n2094 & n10489 ;
  assign n13202 = n3097 & n7712 ;
  assign n13203 = n13202 ^ n1719 ^ 1'b0 ;
  assign n13204 = ( n4559 & n5617 ) | ( n4559 & ~n13203 ) | ( n5617 & ~n13203 ) ;
  assign n13205 = n13201 | n13204 ;
  assign n13216 = n6121 ^ n1645 ^ n260 ;
  assign n13223 = ( n2170 & ~n5951 ) | ( n2170 & n7712 ) | ( ~n5951 & n7712 ) ;
  assign n13221 = ~n7010 & n11064 ;
  assign n13220 = ~n4295 & n5927 ;
  assign n13222 = n13221 ^ n13220 ^ 1'b0 ;
  assign n13224 = n13223 ^ n13222 ^ n7987 ;
  assign n13225 = n3452 & ~n13224 ;
  assign n13217 = ( n6617 & n7708 ) | ( n6617 & ~n9070 ) | ( n7708 & ~n9070 ) ;
  assign n13218 = ( n6276 & n8559 ) | ( n6276 & ~n10577 ) | ( n8559 & ~n10577 ) ;
  assign n13219 = n13217 & ~n13218 ;
  assign n13226 = n13225 ^ n13219 ^ 1'b0 ;
  assign n13227 = n13216 & ~n13226 ;
  assign n13206 = n6748 ^ n3904 ^ x36 ;
  assign n13207 = n1134 & ~n2789 ;
  assign n13208 = n13207 ^ n9016 ^ 1'b0 ;
  assign n13209 = ~n3821 & n13208 ;
  assign n13210 = n13209 ^ n6054 ^ 1'b0 ;
  assign n13211 = n10081 & ~n13210 ;
  assign n13212 = n13211 ^ n9413 ^ 1'b0 ;
  assign n13213 = n11229 & ~n13212 ;
  assign n13214 = ~n13206 & n13213 ;
  assign n13215 = n8170 | n13214 ;
  assign n13228 = n13227 ^ n13215 ^ 1'b0 ;
  assign n13234 = n1353 | n11233 ;
  assign n13229 = n4701 & ~n11546 ;
  assign n13230 = n6398 ^ n1798 ^ n1045 ;
  assign n13231 = n13230 ^ n5136 ^ 1'b0 ;
  assign n13232 = n13231 ^ n7544 ^ n5576 ;
  assign n13233 = n13229 | n13232 ;
  assign n13235 = n13234 ^ n13233 ^ 1'b0 ;
  assign n13236 = n4627 & ~n11408 ;
  assign n13237 = n12942 ^ n2976 ^ n2355 ;
  assign n13238 = n2894 ^ n2135 ^ n231 ;
  assign n13239 = n2075 & n13238 ;
  assign n13240 = n13239 ^ n4118 ^ 1'b0 ;
  assign n13241 = n5644 & n13240 ;
  assign n13242 = ~n282 & n13241 ;
  assign n13243 = n2602 & ~n2805 ;
  assign n13244 = n13243 ^ n12214 ^ 1'b0 ;
  assign n13245 = ( n863 & n13242 ) | ( n863 & n13244 ) | ( n13242 & n13244 ) ;
  assign n13246 = n13245 ^ n7388 ^ 1'b0 ;
  assign n13247 = n2130 & ~n2341 ;
  assign n13248 = n13247 ^ n2880 ^ 1'b0 ;
  assign n13249 = n12126 ^ n7073 ^ n5809 ;
  assign n13250 = n13249 ^ n7021 ^ n2753 ;
  assign n13251 = x50 & ~n13250 ;
  assign n13252 = n13251 ^ n479 ^ 1'b0 ;
  assign n13253 = ( ~n1143 & n2955 ) | ( ~n1143 & n6091 ) | ( n2955 & n6091 ) ;
  assign n13254 = n13253 ^ n10478 ^ 1'b0 ;
  assign n13255 = n4101 ^ n2527 ^ n985 ;
  assign n13256 = ( n1113 & n2609 ) | ( n1113 & n13255 ) | ( n2609 & n13255 ) ;
  assign n13257 = n8636 | n10202 ;
  assign n13258 = ( n1970 & n13256 ) | ( n1970 & n13257 ) | ( n13256 & n13257 ) ;
  assign n13259 = ( n2370 & ~n3662 ) | ( n2370 & n3668 ) | ( ~n3662 & n3668 ) ;
  assign n13260 = n4331 & ~n13259 ;
  assign n13261 = n13260 ^ n1697 ^ 1'b0 ;
  assign n13262 = ( n12914 & n13258 ) | ( n12914 & ~n13261 ) | ( n13258 & ~n13261 ) ;
  assign n13265 = ~n1901 & n8779 ;
  assign n13266 = n6471 ^ n2930 ^ 1'b0 ;
  assign n13267 = n2763 & n13266 ;
  assign n13268 = n5409 & ~n13267 ;
  assign n13269 = n5354 & ~n13268 ;
  assign n13270 = ~n13265 & n13269 ;
  assign n13263 = n3375 | n13173 ;
  assign n13264 = n13263 ^ n7128 ^ n4393 ;
  assign n13271 = n13270 ^ n13264 ^ n3831 ;
  assign n13275 = n1338 | n4578 ;
  assign n13272 = n300 | n7463 ;
  assign n13273 = n13272 ^ n7454 ^ 1'b0 ;
  assign n13274 = n1561 & ~n13273 ;
  assign n13276 = n13275 ^ n13274 ^ 1'b0 ;
  assign n13277 = n13276 ^ n2570 ^ 1'b0 ;
  assign n13278 = n13071 | n13277 ;
  assign n13279 = n10194 & n12337 ;
  assign n13280 = ~n5216 & n13279 ;
  assign n13281 = n8331 ^ n6271 ^ n1624 ;
  assign n13282 = n3436 | n13281 ;
  assign n13283 = n13282 ^ n2521 ^ 1'b0 ;
  assign n13284 = ( n2788 & ~n3950 ) | ( n2788 & n13283 ) | ( ~n3950 & n13283 ) ;
  assign n13285 = n1873 & n2205 ;
  assign n13286 = n2723 & n9753 ;
  assign n13287 = ( n5531 & n13285 ) | ( n5531 & ~n13286 ) | ( n13285 & ~n13286 ) ;
  assign n13290 = n1927 | n3709 ;
  assign n13291 = n13290 ^ n2901 ^ 1'b0 ;
  assign n13288 = ( n1805 & n6276 ) | ( n1805 & n9427 ) | ( n6276 & n9427 ) ;
  assign n13289 = n247 & n13288 ;
  assign n13292 = n13291 ^ n13289 ^ 1'b0 ;
  assign n13293 = n2620 & ~n5091 ;
  assign n13294 = n13293 ^ n6317 ^ 1'b0 ;
  assign n13295 = n3466 ^ n3341 ^ 1'b0 ;
  assign n13296 = ( ~n7733 & n13294 ) | ( ~n7733 & n13295 ) | ( n13294 & n13295 ) ;
  assign n13298 = ( n3740 & n3804 ) | ( n3740 & n7942 ) | ( n3804 & n7942 ) ;
  assign n13297 = n2433 & n5397 ;
  assign n13299 = n13298 ^ n13297 ^ 1'b0 ;
  assign n13300 = n5012 & n13299 ;
  assign n13301 = ~n13296 & n13300 ;
  assign n13302 = ~n9286 & n13301 ;
  assign n13303 = n2710 & n3359 ;
  assign n13304 = ~n1873 & n13303 ;
  assign n13305 = n1629 & n1915 ;
  assign n13306 = n2107 & n13305 ;
  assign n13307 = ( ~n2567 & n4000 ) | ( ~n2567 & n13306 ) | ( n4000 & n13306 ) ;
  assign n13308 = n4994 | n13307 ;
  assign n13309 = n13308 ^ n12848 ^ 1'b0 ;
  assign n13310 = ( n8292 & n13304 ) | ( n8292 & ~n13309 ) | ( n13304 & ~n13309 ) ;
  assign n13311 = n1795 | n12109 ;
  assign n13312 = ~n3926 & n9250 ;
  assign n13313 = n13312 ^ n3826 ^ 1'b0 ;
  assign n13314 = n9625 ^ n4356 ^ 1'b0 ;
  assign n13315 = ~n10758 & n13314 ;
  assign n13316 = n12804 ^ n8538 ^ n8014 ;
  assign n13317 = ( n2006 & n5409 ) | ( n2006 & n13316 ) | ( n5409 & n13316 ) ;
  assign n13318 = ( n13313 & ~n13315 ) | ( n13313 & n13317 ) | ( ~n13315 & n13317 ) ;
  assign n13319 = n13311 & ~n13318 ;
  assign n13320 = ~n13310 & n13319 ;
  assign n13321 = n1832 & n5230 ;
  assign n13322 = n13321 ^ n7651 ^ n6133 ;
  assign n13323 = n12644 ^ n12296 ^ 1'b0 ;
  assign n13324 = n13323 ^ n10776 ^ 1'b0 ;
  assign n13325 = n3912 & ~n5922 ;
  assign n13326 = n2526 ^ n1728 ^ n1382 ;
  assign n13327 = n2157 & n13326 ;
  assign n13328 = ( n1310 & n4050 ) | ( n1310 & n13327 ) | ( n4050 & n13327 ) ;
  assign n13329 = n340 | n2754 ;
  assign n13330 = n1740 | n13329 ;
  assign n13331 = n13330 ^ n10198 ^ n8491 ;
  assign n13332 = ( n1093 & n2358 ) | ( n1093 & n6774 ) | ( n2358 & n6774 ) ;
  assign n13333 = n1343 & ~n4234 ;
  assign n13334 = n1285 ^ n316 ^ 1'b0 ;
  assign n13335 = ( ~n2932 & n6103 ) | ( ~n2932 & n13334 ) | ( n6103 & n13334 ) ;
  assign n13336 = ( ~n2588 & n7193 ) | ( ~n2588 & n13335 ) | ( n7193 & n13335 ) ;
  assign n13337 = n5995 & n13336 ;
  assign n13338 = n13333 & n13337 ;
  assign n13339 = ~n319 & n4546 ;
  assign n13340 = n2609 & ~n3362 ;
  assign n13341 = ~n13339 & n13340 ;
  assign n13342 = ( ~n3678 & n11428 ) | ( ~n3678 & n13341 ) | ( n11428 & n13341 ) ;
  assign n13347 = ( n7943 & n8200 ) | ( n7943 & n8828 ) | ( n8200 & n8828 ) ;
  assign n13343 = n7528 ^ n3666 ^ 1'b0 ;
  assign n13344 = ( ~n1850 & n5507 ) | ( ~n1850 & n13343 ) | ( n5507 & n13343 ) ;
  assign n13345 = n10383 ^ n8978 ^ n2178 ;
  assign n13346 = n13344 | n13345 ;
  assign n13348 = n13347 ^ n13346 ^ 1'b0 ;
  assign n13353 = ( n1999 & n6115 ) | ( n1999 & ~n6750 ) | ( n6115 & ~n6750 ) ;
  assign n13349 = ( n2834 & n3644 ) | ( n2834 & n10484 ) | ( n3644 & n10484 ) ;
  assign n13350 = ~n4231 & n8636 ;
  assign n13351 = n13350 ^ n2048 ^ 1'b0 ;
  assign n13352 = n13349 & ~n13351 ;
  assign n13354 = n13353 ^ n13352 ^ 1'b0 ;
  assign n13355 = n5546 ^ n5457 ^ 1'b0 ;
  assign n13356 = n4880 & ~n13355 ;
  assign n13357 = ( n5854 & n9225 ) | ( n5854 & ~n10940 ) | ( n9225 & ~n10940 ) ;
  assign n13358 = n13357 ^ n8302 ^ n6700 ;
  assign n13359 = n1547 & ~n6112 ;
  assign n13360 = n2523 & n13359 ;
  assign n13361 = n298 | n13360 ;
  assign n13362 = n7185 & ~n13361 ;
  assign n13363 = n13362 ^ n9829 ^ n8269 ;
  assign n13364 = x26 & ~n8870 ;
  assign n13365 = n2579 & n13364 ;
  assign n13366 = n3690 ^ n2370 ^ n1062 ;
  assign n13367 = n3085 | n13366 ;
  assign n13368 = n13367 ^ n2209 ^ 1'b0 ;
  assign n13370 = n11027 ^ n415 ^ 1'b0 ;
  assign n13371 = n13370 ^ n4468 ^ x70 ;
  assign n13369 = n8475 & ~n11246 ;
  assign n13372 = n13371 ^ n13369 ^ 1'b0 ;
  assign n13373 = n1179 ^ n788 ^ 1'b0 ;
  assign n13374 = n4186 & n13373 ;
  assign n13375 = n13374 ^ n1962 ^ 1'b0 ;
  assign n13376 = ~n219 & n13375 ;
  assign n13377 = n5061 | n13222 ;
  assign n13378 = n13376 | n13377 ;
  assign n13379 = n13378 ^ n10390 ^ n4226 ;
  assign n13380 = n13379 ^ n13253 ^ 1'b0 ;
  assign n13381 = n4944 & n13380 ;
  assign n13382 = n2414 & ~n3763 ;
  assign n13383 = ( n5759 & ~n12273 ) | ( n5759 & n13382 ) | ( ~n12273 & n13382 ) ;
  assign n13384 = n13383 ^ n8582 ^ 1'b0 ;
  assign n13385 = n13384 ^ n13024 ^ 1'b0 ;
  assign n13386 = ~n3957 & n5409 ;
  assign n13387 = ( n2507 & ~n2913 ) | ( n2507 & n13386 ) | ( ~n2913 & n13386 ) ;
  assign n13388 = n13387 ^ n1786 ^ 1'b0 ;
  assign n13389 = n12207 ^ n6937 ^ 1'b0 ;
  assign n13390 = n2911 | n13389 ;
  assign n13391 = ( n1244 & n3292 ) | ( n1244 & n3941 ) | ( n3292 & n3941 ) ;
  assign n13392 = ~n9198 & n13391 ;
  assign n13393 = n13392 ^ n5076 ^ 1'b0 ;
  assign n13397 = n905 & ~n5397 ;
  assign n13398 = n13397 ^ n11249 ^ 1'b0 ;
  assign n13399 = n941 & n13398 ;
  assign n13400 = ~n7141 & n13399 ;
  assign n13394 = n5623 & n6770 ;
  assign n13395 = ~n828 & n9941 ;
  assign n13396 = n13394 & n13395 ;
  assign n13401 = n13400 ^ n13396 ^ n10463 ;
  assign n13408 = n1813 ^ n1356 ^ 1'b0 ;
  assign n13409 = n2334 & n13408 ;
  assign n13402 = ( n2458 & n2801 ) | ( n2458 & n5048 ) | ( n2801 & n5048 ) ;
  assign n13403 = n13402 ^ n438 ^ 1'b0 ;
  assign n13404 = n10041 & n13403 ;
  assign n13405 = n13404 ^ n12178 ^ n699 ;
  assign n13406 = n13405 ^ n13035 ^ 1'b0 ;
  assign n13407 = ( n6430 & n9819 ) | ( n6430 & ~n13406 ) | ( n9819 & ~n13406 ) ;
  assign n13410 = n13409 ^ n13407 ^ 1'b0 ;
  assign n13414 = n4477 ^ n3985 ^ 1'b0 ;
  assign n13411 = n8281 ^ n7825 ^ n3053 ;
  assign n13412 = ~n5477 & n13411 ;
  assign n13413 = n3218 & n13412 ;
  assign n13415 = n13414 ^ n13413 ^ 1'b0 ;
  assign n13416 = ( ~n1260 & n3558 ) | ( ~n1260 & n3577 ) | ( n3558 & n3577 ) ;
  assign n13417 = n13416 ^ n5600 ^ 1'b0 ;
  assign n13418 = n6815 & ~n13417 ;
  assign n13421 = ( n821 & ~n3798 ) | ( n821 & n6441 ) | ( ~n3798 & n6441 ) ;
  assign n13422 = n13421 ^ n1494 ^ 1'b0 ;
  assign n13423 = n2021 & n13422 ;
  assign n13424 = n8037 & n13423 ;
  assign n13425 = n13424 ^ n6308 ^ 1'b0 ;
  assign n13419 = ~n1431 & n3850 ;
  assign n13420 = n13419 ^ n2973 ^ 1'b0 ;
  assign n13426 = n13425 ^ n13420 ^ n7549 ;
  assign n13427 = n5998 ^ n422 ^ 1'b0 ;
  assign n13428 = ~n3393 & n13427 ;
  assign n13429 = n13428 ^ n5048 ^ 1'b0 ;
  assign n13430 = n13429 ^ n6868 ^ x32 ;
  assign n13431 = n13430 ^ n13032 ^ n11083 ;
  assign n13432 = n3002 & ~n9041 ;
  assign n13433 = n13432 ^ n3063 ^ 1'b0 ;
  assign n13434 = ( n6715 & n7616 ) | ( n6715 & n11166 ) | ( n7616 & n11166 ) ;
  assign n13435 = ~n9088 & n12307 ;
  assign n13436 = ~x26 & n13435 ;
  assign n13437 = ( n3841 & n5068 ) | ( n3841 & n13436 ) | ( n5068 & n13436 ) ;
  assign n13438 = ( n4342 & n4923 ) | ( n4342 & ~n10286 ) | ( n4923 & ~n10286 ) ;
  assign n13439 = n13438 ^ n2494 ^ 1'b0 ;
  assign n13440 = n13439 ^ n10503 ^ n10413 ;
  assign n13441 = ( n778 & n924 ) | ( n778 & ~n11585 ) | ( n924 & ~n11585 ) ;
  assign n13442 = ( n8360 & n9966 ) | ( n8360 & n13441 ) | ( n9966 & n13441 ) ;
  assign n13443 = n2634 | n13442 ;
  assign n13444 = n11125 ^ n8127 ^ n386 ;
  assign n13445 = ( n5865 & n9260 ) | ( n5865 & n13444 ) | ( n9260 & n13444 ) ;
  assign n13446 = n4162 ^ n642 ^ 1'b0 ;
  assign n13447 = n8686 & n13446 ;
  assign n13448 = ( n5721 & n10166 ) | ( n5721 & n13447 ) | ( n10166 & n13447 ) ;
  assign n13449 = n1123 ^ n674 ^ 1'b0 ;
  assign n13450 = ( n2390 & ~n13448 ) | ( n2390 & n13449 ) | ( ~n13448 & n13449 ) ;
  assign n13452 = n1783 & ~n6901 ;
  assign n13453 = n3475 & n13452 ;
  assign n13454 = ( n6115 & n8465 ) | ( n6115 & n13453 ) | ( n8465 & n13453 ) ;
  assign n13451 = n1893 & n6239 ;
  assign n13455 = n13454 ^ n13451 ^ n6627 ;
  assign n13458 = n6937 ^ n1095 ^ n836 ;
  assign n13459 = ( n4940 & n5568 ) | ( n4940 & ~n13458 ) | ( n5568 & ~n13458 ) ;
  assign n13456 = n1341 & n2414 ;
  assign n13457 = n5947 & n13456 ;
  assign n13460 = n13459 ^ n13457 ^ n8338 ;
  assign n13461 = n2274 & ~n13460 ;
  assign n13462 = n13461 ^ n5031 ^ 1'b0 ;
  assign n13463 = ( n1744 & n7342 ) | ( n1744 & n10344 ) | ( n7342 & n10344 ) ;
  assign n13464 = ~n1166 & n13463 ;
  assign n13465 = ~n9265 & n13464 ;
  assign n13466 = ( ~n10618 & n13462 ) | ( ~n10618 & n13465 ) | ( n13462 & n13465 ) ;
  assign n13467 = n12715 ^ n6619 ^ 1'b0 ;
  assign n13468 = n5193 ^ n4739 ^ n2818 ;
  assign n13469 = ~n7927 & n11426 ;
  assign n13470 = ~n13468 & n13469 ;
  assign n13471 = n1528 & ~n2713 ;
  assign n13472 = ~n8204 & n9890 ;
  assign n13473 = n13472 ^ n10753 ^ 1'b0 ;
  assign n13474 = n13473 ^ n8792 ^ n5310 ;
  assign n13475 = n13474 ^ n9190 ^ n2834 ;
  assign n13477 = n1262 | n1926 ;
  assign n13478 = n13477 ^ n2633 ^ 1'b0 ;
  assign n13479 = ( n6579 & ~n7845 ) | ( n6579 & n13478 ) | ( ~n7845 & n13478 ) ;
  assign n13476 = ~n4150 & n8591 ;
  assign n13480 = n13479 ^ n13476 ^ 1'b0 ;
  assign n13485 = n1651 | n10533 ;
  assign n13486 = n13485 ^ n3484 ^ 1'b0 ;
  assign n13487 = n7141 & n13486 ;
  assign n13481 = n5622 & ~n13460 ;
  assign n13482 = n5139 & n13481 ;
  assign n13483 = n13482 ^ n9617 ^ n1270 ;
  assign n13484 = ~n1359 & n13483 ;
  assign n13488 = n13487 ^ n13484 ^ n1871 ;
  assign n13489 = ( n2851 & n8849 ) | ( n2851 & n12178 ) | ( n8849 & n12178 ) ;
  assign n13490 = n12626 ^ n8703 ^ 1'b0 ;
  assign n13491 = n5598 & ~n8559 ;
  assign n13492 = n957 ^ n539 ^ 1'b0 ;
  assign n13493 = ( n2116 & n5060 ) | ( n2116 & ~n8258 ) | ( n5060 & ~n8258 ) ;
  assign n13494 = n7765 ^ n5431 ^ 1'b0 ;
  assign n13495 = n13493 & n13494 ;
  assign n13496 = n1448 ^ n602 ^ 1'b0 ;
  assign n13497 = n4521 ^ n2938 ^ 1'b0 ;
  assign n13498 = n601 & ~n13497 ;
  assign n13499 = n13498 ^ n8367 ^ 1'b0 ;
  assign n13500 = n2029 & n13499 ;
  assign n13501 = n2419 & n13500 ;
  assign n13502 = n13501 ^ n7789 ^ n6378 ;
  assign n13503 = n4688 & n4761 ;
  assign n13504 = n3285 & n13503 ;
  assign n13505 = n7560 ^ n4145 ^ n1916 ;
  assign n13506 = n13504 & ~n13505 ;
  assign n13507 = n8482 ^ n8431 ^ n219 ;
  assign n13508 = ( n4282 & ~n7275 ) | ( n4282 & n12279 ) | ( ~n7275 & n12279 ) ;
  assign n13509 = n13508 ^ n5327 ^ 1'b0 ;
  assign n13510 = n13479 ^ n8825 ^ n7276 ;
  assign n13511 = ( ~n476 & n1038 ) | ( ~n476 & n13510 ) | ( n1038 & n13510 ) ;
  assign n13512 = n4834 & n13511 ;
  assign n13513 = n13509 & n13512 ;
  assign n13514 = x93 & ~n8814 ;
  assign n13515 = n13513 & n13514 ;
  assign n13518 = ( n312 & n2356 ) | ( n312 & ~n2541 ) | ( n2356 & ~n2541 ) ;
  assign n13519 = n13518 ^ n8834 ^ n4010 ;
  assign n13516 = ( n3062 & ~n3627 ) | ( n3062 & n3834 ) | ( ~n3627 & n3834 ) ;
  assign n13517 = n7192 | n13516 ;
  assign n13520 = n13519 ^ n13517 ^ n4363 ;
  assign n13521 = ( n747 & n6307 ) | ( n747 & n13520 ) | ( n6307 & n13520 ) ;
  assign n13522 = n2674 ^ n405 ^ 1'b0 ;
  assign n13523 = ~n7274 & n13522 ;
  assign n13524 = n7893 & n13523 ;
  assign n13525 = n13524 ^ n13265 ^ n12958 ;
  assign n13526 = n5357 & n10957 ;
  assign n13527 = n13526 ^ n783 ^ 1'b0 ;
  assign n13528 = n4372 & ~n9370 ;
  assign n13530 = n1953 ^ n1672 ^ n527 ;
  assign n13529 = n6361 ^ n5127 ^ x96 ;
  assign n13531 = n13530 ^ n13529 ^ n1118 ;
  assign n13532 = ( ~n2698 & n3291 ) | ( ~n2698 & n12826 ) | ( n3291 & n12826 ) ;
  assign n13533 = n13532 ^ n11686 ^ n4148 ;
  assign n13534 = n1945 | n10416 ;
  assign n13535 = n13534 ^ n4758 ^ 1'b0 ;
  assign n13536 = ( n309 & n4848 ) | ( n309 & n7627 ) | ( n4848 & n7627 ) ;
  assign n13537 = ~n4265 & n13536 ;
  assign n13538 = n13537 ^ n11248 ^ 1'b0 ;
  assign n13539 = ( ~n10260 & n13535 ) | ( ~n10260 & n13538 ) | ( n13535 & n13538 ) ;
  assign n13540 = n10480 ^ x36 ^ 1'b0 ;
  assign n13541 = n12268 ^ n10947 ^ n3035 ;
  assign n13542 = ~n8180 & n13541 ;
  assign n13543 = ( n1477 & n3510 ) | ( n1477 & n13542 ) | ( n3510 & n13542 ) ;
  assign n13544 = n7281 | n13543 ;
  assign n13545 = n13544 ^ n2991 ^ 1'b0 ;
  assign n13546 = n5466 | n12449 ;
  assign n13547 = n3210 & ~n4248 ;
  assign n13548 = n13547 ^ n7770 ^ 1'b0 ;
  assign n13549 = n12585 ^ n1996 ^ n971 ;
  assign n13550 = n13549 ^ n12228 ^ n5550 ;
  assign n13551 = n4704 ^ n2486 ^ 1'b0 ;
  assign n13552 = n13551 ^ n10325 ^ n6343 ;
  assign n13553 = ( n9835 & n12653 ) | ( n9835 & n13552 ) | ( n12653 & n13552 ) ;
  assign n13554 = ( n1567 & ~n3248 ) | ( n1567 & n11523 ) | ( ~n3248 & n11523 ) ;
  assign n13555 = ( n6452 & n9079 ) | ( n6452 & n13554 ) | ( n9079 & n13554 ) ;
  assign n13556 = n10701 ^ n9297 ^ 1'b0 ;
  assign n13557 = n12305 ^ n6835 ^ 1'b0 ;
  assign n13558 = n2072 & n13557 ;
  assign n13559 = ( n10185 & n13326 ) | ( n10185 & n13558 ) | ( n13326 & n13558 ) ;
  assign n13561 = ( n8322 & n9397 ) | ( n8322 & ~n10701 ) | ( n9397 & ~n10701 ) ;
  assign n13560 = ( n577 & n1335 ) | ( n577 & n12339 ) | ( n1335 & n12339 ) ;
  assign n13562 = n13561 ^ n13560 ^ n6880 ;
  assign n13563 = n5384 & n5904 ;
  assign n13564 = n13563 ^ n2026 ^ 1'b0 ;
  assign n13565 = n2999 & ~n13564 ;
  assign n13566 = ( n9344 & n10438 ) | ( n9344 & n12268 ) | ( n10438 & n12268 ) ;
  assign n13567 = n9214 ^ n8660 ^ 1'b0 ;
  assign n13568 = x38 & ~n7334 ;
  assign n13569 = ( ~n5041 & n5959 ) | ( ~n5041 & n13568 ) | ( n5959 & n13568 ) ;
  assign n13570 = n6522 ^ n294 ^ 1'b0 ;
  assign n13571 = ~n5264 & n13570 ;
  assign n13572 = ~n13569 & n13571 ;
  assign n13573 = n13572 ^ n10575 ^ 1'b0 ;
  assign n13574 = n13573 ^ n8722 ^ 1'b0 ;
  assign n13575 = ~n11395 & n13574 ;
  assign n13576 = ( n517 & n13567 ) | ( n517 & n13575 ) | ( n13567 & n13575 ) ;
  assign n13577 = n10599 ^ n8635 ^ n3439 ;
  assign n13578 = ( n298 & n8118 ) | ( n298 & ~n13577 ) | ( n8118 & ~n13577 ) ;
  assign n13579 = n13578 ^ n10227 ^ n9291 ;
  assign n13580 = ( x48 & n3619 ) | ( x48 & ~n4906 ) | ( n3619 & ~n4906 ) ;
  assign n13581 = n5732 ^ n4759 ^ n967 ;
  assign n13582 = ( n4072 & ~n13189 ) | ( n4072 & n13581 ) | ( ~n13189 & n13581 ) ;
  assign n13584 = n11528 ^ n7243 ^ n3925 ;
  assign n13583 = n9319 & n10785 ;
  assign n13585 = n13584 ^ n13583 ^ 1'b0 ;
  assign n13586 = n4010 & ~n13585 ;
  assign n13587 = n11783 & ~n12827 ;
  assign n13588 = n13587 ^ n11764 ^ 1'b0 ;
  assign n13589 = n897 ^ n450 ^ 1'b0 ;
  assign n13590 = n10930 | n13589 ;
  assign n13591 = n7033 ^ n4220 ^ 1'b0 ;
  assign n13592 = ( n6992 & n12028 ) | ( n6992 & ~n13591 ) | ( n12028 & ~n13591 ) ;
  assign n13595 = n9563 ^ n1154 ^ n1127 ;
  assign n13596 = ~n983 & n13595 ;
  assign n13597 = n5436 & n13596 ;
  assign n13593 = n2435 & n6334 ;
  assign n13594 = n13593 ^ n8119 ^ 1'b0 ;
  assign n13598 = n13597 ^ n13594 ^ n4108 ;
  assign n13599 = ( ~n1994 & n4063 ) | ( ~n1994 & n5023 ) | ( n4063 & n5023 ) ;
  assign n13600 = ( ~n10982 & n13173 ) | ( ~n10982 & n13599 ) | ( n13173 & n13599 ) ;
  assign n13601 = ( ~n6504 & n13598 ) | ( ~n6504 & n13600 ) | ( n13598 & n13600 ) ;
  assign n13602 = n7904 | n8132 ;
  assign n13603 = n2106 & n8211 ;
  assign n13604 = n1783 & ~n4084 ;
  assign n13605 = n13603 & n13604 ;
  assign n13606 = n12587 ^ n2432 ^ 1'b0 ;
  assign n13607 = n3892 & n13206 ;
  assign n13608 = n413 & n1275 ;
  assign n13609 = ~n8559 & n13608 ;
  assign n13610 = n13609 ^ n6708 ^ n4453 ;
  assign n13611 = ~n6300 & n7401 ;
  assign n13612 = n13611 ^ n810 ^ 1'b0 ;
  assign n13613 = n570 & n2481 ;
  assign n13614 = ~n4801 & n13613 ;
  assign n13615 = n12336 & ~n13338 ;
  assign n13616 = n13615 ^ x19 ^ 1'b0 ;
  assign n13618 = ( n7288 & n12059 ) | ( n7288 & ~n12541 ) | ( n12059 & ~n12541 ) ;
  assign n13617 = n8994 & ~n10157 ;
  assign n13619 = n13618 ^ n13617 ^ 1'b0 ;
  assign n13620 = x8 & ~n2502 ;
  assign n13621 = n13620 ^ n1259 ^ 1'b0 ;
  assign n13622 = ( n1654 & ~n10035 ) | ( n1654 & n13621 ) | ( ~n10035 & n13621 ) ;
  assign n13623 = ~n6610 & n13622 ;
  assign n13624 = n13482 ^ n10930 ^ 1'b0 ;
  assign n13625 = ( ~n3335 & n6013 ) | ( ~n3335 & n13624 ) | ( n6013 & n13624 ) ;
  assign n13627 = n1656 | n7135 ;
  assign n13628 = n13627 ^ n5936 ^ 1'b0 ;
  assign n13626 = n3408 & ~n7468 ;
  assign n13629 = n13628 ^ n13626 ^ 1'b0 ;
  assign n13630 = n13629 ^ n4074 ^ 1'b0 ;
  assign n13631 = n8372 & ~n13630 ;
  assign n13632 = x86 & ~n1738 ;
  assign n13633 = n13632 ^ n5282 ^ 1'b0 ;
  assign n13634 = n12449 | n13633 ;
  assign n13635 = n13634 ^ n11978 ^ 1'b0 ;
  assign n13636 = n1775 ^ n976 ^ 1'b0 ;
  assign n13637 = n13635 | n13636 ;
  assign n13638 = n13637 ^ n4953 ^ 1'b0 ;
  assign n13639 = n11405 | n13638 ;
  assign n13646 = n5149 & ~n6024 ;
  assign n13643 = n7611 ^ n4077 ^ 1'b0 ;
  assign n13644 = n7893 | n13643 ;
  assign n13645 = ( n1767 & n8302 ) | ( n1767 & n13644 ) | ( n8302 & n13644 ) ;
  assign n13640 = ( ~n1765 & n6822 ) | ( ~n1765 & n9655 ) | ( n6822 & n9655 ) ;
  assign n13641 = n13640 ^ n3602 ^ 1'b0 ;
  assign n13642 = n5769 & ~n13641 ;
  assign n13647 = n13646 ^ n13645 ^ n13642 ;
  assign n13648 = n4373 ^ n1744 ^ n733 ;
  assign n13649 = ( x26 & n323 ) | ( x26 & n13648 ) | ( n323 & n13648 ) ;
  assign n13650 = ( n6576 & n7241 ) | ( n6576 & n9748 ) | ( n7241 & n9748 ) ;
  assign n13651 = ( n11515 & ~n13649 ) | ( n11515 & n13650 ) | ( ~n13649 & n13650 ) ;
  assign n13652 = n7225 ^ n2965 ^ 1'b0 ;
  assign n13653 = ~n9943 & n13652 ;
  assign n13654 = ( n5269 & n8172 ) | ( n5269 & ~n13653 ) | ( n8172 & ~n13653 ) ;
  assign n13655 = ~n3019 & n6090 ;
  assign n13656 = n3346 & n13655 ;
  assign n13657 = n7210 ^ n5562 ^ n1583 ;
  assign n13658 = n1418 & n13657 ;
  assign n13659 = n6016 ^ n3205 ^ 1'b0 ;
  assign n13660 = ~n13658 & n13659 ;
  assign n13661 = ( x20 & ~n1180 ) | ( x20 & n8026 ) | ( ~n1180 & n8026 ) ;
  assign n13662 = n8147 & n13661 ;
  assign n13663 = n13662 ^ n10100 ^ 1'b0 ;
  assign n13664 = n13663 ^ n5250 ^ n1426 ;
  assign n13665 = ~n4462 & n13664 ;
  assign n13670 = n6741 ^ n3474 ^ 1'b0 ;
  assign n13666 = n11305 ^ x7 ^ 1'b0 ;
  assign n13667 = n7309 & ~n13666 ;
  assign n13668 = n1999 ^ n1636 ^ 1'b0 ;
  assign n13669 = n13667 & n13668 ;
  assign n13671 = n13670 ^ n13669 ^ 1'b0 ;
  assign n13672 = ( n1334 & n7347 ) | ( n1334 & ~n8877 ) | ( n7347 & ~n8877 ) ;
  assign n13673 = ( n3785 & ~n7091 ) | ( n3785 & n13672 ) | ( ~n7091 & n13672 ) ;
  assign n13674 = n6067 ^ n2794 ^ 1'b0 ;
  assign n13675 = ( n5123 & ~n6607 ) | ( n5123 & n7180 ) | ( ~n6607 & n7180 ) ;
  assign n13676 = n13675 ^ n9677 ^ 1'b0 ;
  assign n13677 = ( n1053 & n4576 ) | ( n1053 & n13676 ) | ( n4576 & n13676 ) ;
  assign n13678 = n1543 ^ n1474 ^ 1'b0 ;
  assign n13679 = n11028 ^ n3364 ^ 1'b0 ;
  assign n13680 = n2209 & ~n13679 ;
  assign n13681 = ( n6265 & n13678 ) | ( n6265 & ~n13680 ) | ( n13678 & ~n13680 ) ;
  assign n13682 = ~n5634 & n7895 ;
  assign n13683 = n13682 ^ n7820 ^ 1'b0 ;
  assign n13684 = n10960 ^ n6736 ^ n4575 ;
  assign n13686 = n1284 & n6455 ;
  assign n13687 = n11488 & n13686 ;
  assign n13688 = n13687 ^ n9646 ^ n9016 ;
  assign n13685 = n4620 ^ n3593 ^ n1509 ;
  assign n13689 = n13688 ^ n13685 ^ n9577 ;
  assign n13692 = ~n10167 & n12871 ;
  assign n13693 = n3969 & n13692 ;
  assign n13694 = ( n625 & n3374 ) | ( n625 & ~n3441 ) | ( n3374 & ~n3441 ) ;
  assign n13695 = ~n8757 & n13694 ;
  assign n13696 = n13693 & n13695 ;
  assign n13690 = n12893 ^ n6190 ^ n3819 ;
  assign n13691 = n3976 & ~n13690 ;
  assign n13697 = n13696 ^ n13691 ^ 1'b0 ;
  assign n13698 = n13697 ^ n2789 ^ 1'b0 ;
  assign n13699 = n12071 ^ n10994 ^ n5641 ;
  assign n13700 = ( n263 & n495 ) | ( n263 & ~n1137 ) | ( n495 & ~n1137 ) ;
  assign n13701 = n2930 & ~n13700 ;
  assign n13702 = ( n5205 & n7566 ) | ( n5205 & ~n7882 ) | ( n7566 & ~n7882 ) ;
  assign n13703 = ( n2584 & n13701 ) | ( n2584 & n13702 ) | ( n13701 & n13702 ) ;
  assign n13709 = ~n199 & n4220 ;
  assign n13710 = ~n5770 & n13709 ;
  assign n13711 = n13710 ^ n983 ^ 1'b0 ;
  assign n13707 = ~n3706 & n7315 ;
  assign n13708 = n4514 & n13707 ;
  assign n13712 = n13711 ^ n13708 ^ n5489 ;
  assign n13704 = ( ~n2865 & n3386 ) | ( ~n2865 & n12298 ) | ( n3386 & n12298 ) ;
  assign n13705 = ( n1714 & n3383 ) | ( n1714 & n13704 ) | ( n3383 & n13704 ) ;
  assign n13706 = n13705 ^ n9236 ^ n6193 ;
  assign n13713 = n13712 ^ n13706 ^ n7640 ;
  assign n13714 = n2405 & n13713 ;
  assign n13715 = ~n1364 & n13714 ;
  assign n13716 = n8037 ^ n7299 ^ 1'b0 ;
  assign n13717 = n529 | n13716 ;
  assign n13718 = n1964 | n6741 ;
  assign n13719 = ~n13717 & n13718 ;
  assign n13720 = ( ~x62 & n4209 ) | ( ~x62 & n10697 ) | ( n4209 & n10697 ) ;
  assign n13721 = ( n289 & ~n334 ) | ( n289 & n840 ) | ( ~n334 & n840 ) ;
  assign n13722 = n13721 ^ n189 ^ 1'b0 ;
  assign n13723 = n13722 ^ n1588 ^ n1277 ;
  assign n13724 = n13723 ^ n10548 ^ 1'b0 ;
  assign n13725 = x51 & ~n1180 ;
  assign n13726 = n13725 ^ n8978 ^ 1'b0 ;
  assign n13727 = n3330 ^ n2169 ^ n2067 ;
  assign n13728 = n13727 ^ n12662 ^ n2243 ;
  assign n13729 = n13172 ^ n3829 ^ 1'b0 ;
  assign n13730 = n7859 ^ n1460 ^ 1'b0 ;
  assign n13731 = ( ~n444 & n924 ) | ( ~n444 & n6187 ) | ( n924 & n6187 ) ;
  assign n13732 = n2681 & ~n13731 ;
  assign n13733 = ~n2875 & n13732 ;
  assign n13734 = n4538 & n13733 ;
  assign n13741 = n7104 ^ n3595 ^ n1490 ;
  assign n13738 = ( n1292 & n2431 ) | ( n1292 & ~n2761 ) | ( n2431 & ~n2761 ) ;
  assign n13739 = n13738 ^ n5977 ^ n3516 ;
  assign n13736 = n7018 ^ n5806 ^ n1911 ;
  assign n13735 = ( n5564 & n6671 ) | ( n5564 & ~n8633 ) | ( n6671 & ~n8633 ) ;
  assign n13737 = n13736 ^ n13735 ^ 1'b0 ;
  assign n13740 = n13739 ^ n13737 ^ 1'b0 ;
  assign n13742 = n13741 ^ n13740 ^ n2254 ;
  assign n13743 = ( n3213 & n4788 ) | ( n3213 & ~n8419 ) | ( n4788 & ~n8419 ) ;
  assign n13744 = ( n4566 & ~n7167 ) | ( n4566 & n13743 ) | ( ~n7167 & n13743 ) ;
  assign n13745 = n13744 ^ n4860 ^ x92 ;
  assign n13746 = n3160 & ~n8329 ;
  assign n13747 = n5149 ^ n4482 ^ n2487 ;
  assign n13748 = ~n8582 & n13747 ;
  assign n13749 = n7643 & n13748 ;
  assign n13753 = ~n8678 & n9461 ;
  assign n13754 = n8577 & n13753 ;
  assign n13750 = n8783 ^ n2983 ^ n2622 ;
  assign n13751 = ( n2470 & ~n10090 ) | ( n2470 & n12129 ) | ( ~n10090 & n12129 ) ;
  assign n13752 = ( n461 & n13750 ) | ( n461 & n13751 ) | ( n13750 & n13751 ) ;
  assign n13755 = n13754 ^ n13752 ^ n10608 ;
  assign n13756 = n13755 ^ n7929 ^ n7781 ;
  assign n13757 = n2136 & ~n6168 ;
  assign n13758 = ~n10235 & n11622 ;
  assign n13759 = n8450 & n13758 ;
  assign n13760 = n4022 & ~n4208 ;
  assign n13761 = ~n1586 & n13760 ;
  assign n13762 = ( ~n4411 & n10774 ) | ( ~n4411 & n13761 ) | ( n10774 & n13761 ) ;
  assign n13763 = n6715 ^ n5804 ^ n617 ;
  assign n13764 = n13763 ^ n5046 ^ 1'b0 ;
  assign n13765 = ~n7344 & n13764 ;
  assign n13766 = n13765 ^ n8743 ^ 1'b0 ;
  assign n13767 = n13423 ^ n256 ^ 1'b0 ;
  assign n13768 = n13767 ^ n472 ^ 1'b0 ;
  assign n13769 = n1940 ^ n391 ^ 1'b0 ;
  assign n13770 = n9403 ^ n7627 ^ 1'b0 ;
  assign n13771 = n13769 & ~n13770 ;
  assign n13772 = ~n2859 & n9941 ;
  assign n13773 = ~n3664 & n13772 ;
  assign n13774 = ~n3150 & n7952 ;
  assign n13776 = n12349 ^ n1444 ^ 1'b0 ;
  assign n13775 = n5125 ^ n3269 ^ n624 ;
  assign n13777 = n13776 ^ n13775 ^ n6064 ;
  assign n13778 = n5331 | n10922 ;
  assign n13779 = n13747 | n13778 ;
  assign n13780 = n13779 ^ n825 ^ 1'b0 ;
  assign n13781 = n9843 ^ n7951 ^ n6057 ;
  assign n13782 = ( ~n1426 & n4870 ) | ( ~n1426 & n13781 ) | ( n4870 & n13781 ) ;
  assign n13783 = ( ~n2035 & n13780 ) | ( ~n2035 & n13782 ) | ( n13780 & n13782 ) ;
  assign n13784 = ( n4956 & n9739 ) | ( n4956 & n12283 ) | ( n9739 & n12283 ) ;
  assign n13785 = ~n1964 & n5114 ;
  assign n13786 = ( n1205 & n5891 ) | ( n1205 & ~n13785 ) | ( n5891 & ~n13785 ) ;
  assign n13787 = n580 | n6610 ;
  assign n13788 = n13787 ^ n6714 ^ 1'b0 ;
  assign n13789 = ( n8566 & ~n11677 ) | ( n8566 & n13788 ) | ( ~n11677 & n13788 ) ;
  assign n13790 = n13789 ^ n11515 ^ 1'b0 ;
  assign n13791 = ~n5784 & n8955 ;
  assign n13792 = n7270 & n13791 ;
  assign n13793 = n13792 ^ n4376 ^ 1'b0 ;
  assign n13794 = n2346 & n12668 ;
  assign n13795 = n13605 ^ n2347 ^ n1259 ;
  assign n13796 = n12691 ^ n9528 ^ n4824 ;
  assign n13799 = ( n2880 & n3354 ) | ( n2880 & n5735 ) | ( n3354 & n5735 ) ;
  assign n13800 = ~n709 & n13799 ;
  assign n13797 = ( ~n5425 & n11632 ) | ( ~n5425 & n13529 ) | ( n11632 & n13529 ) ;
  assign n13798 = n551 | n13797 ;
  assign n13801 = n13800 ^ n13798 ^ 1'b0 ;
  assign n13802 = n1547 ^ n1498 ^ 1'b0 ;
  assign n13803 = ( n8371 & ~n10740 ) | ( n8371 & n12595 ) | ( ~n10740 & n12595 ) ;
  assign n13804 = n13802 & n13803 ;
  assign n13805 = n13804 ^ n8987 ^ 1'b0 ;
  assign n13806 = n13801 | n13805 ;
  assign n13807 = n4818 ^ n1925 ^ 1'b0 ;
  assign n13808 = n999 | n5613 ;
  assign n13809 = n13807 | n13808 ;
  assign n13810 = ( n547 & ~n6787 ) | ( n547 & n13809 ) | ( ~n6787 & n13809 ) ;
  assign n13815 = n5333 ^ n1608 ^ 1'b0 ;
  assign n13816 = ~n2548 & n13815 ;
  assign n13811 = n1299 | n8718 ;
  assign n13812 = n13811 ^ n4674 ^ 1'b0 ;
  assign n13813 = n12201 | n13812 ;
  assign n13814 = n410 & ~n13813 ;
  assign n13817 = n13816 ^ n13814 ^ 1'b0 ;
  assign n13818 = ( n2459 & n6532 ) | ( n2459 & ~n13817 ) | ( n6532 & ~n13817 ) ;
  assign n13819 = n3188 | n7724 ;
  assign n13820 = n3969 ^ n1334 ^ 1'b0 ;
  assign n13821 = n13820 ^ n12785 ^ 1'b0 ;
  assign n13822 = ( n1662 & n2549 ) | ( n1662 & n8352 ) | ( n2549 & n8352 ) ;
  assign n13823 = n13822 ^ n654 ^ 1'b0 ;
  assign n13824 = ~n2417 & n10267 ;
  assign n13825 = n4989 & n13824 ;
  assign n13827 = n9015 & ~n13504 ;
  assign n13828 = n4974 ^ n2906 ^ n2341 ;
  assign n13829 = ~n11344 & n13828 ;
  assign n13830 = n13827 & n13829 ;
  assign n13826 = n5729 & ~n9245 ;
  assign n13831 = n13830 ^ n13826 ^ 1'b0 ;
  assign n13833 = n5981 ^ n5928 ^ 1'b0 ;
  assign n13834 = ~n10949 & n13833 ;
  assign n13835 = ( n1900 & n5883 ) | ( n1900 & ~n13834 ) | ( n5883 & ~n13834 ) ;
  assign n13832 = ~n4639 & n8252 ;
  assign n13836 = n13835 ^ n13832 ^ 1'b0 ;
  assign n13837 = ~n1887 & n12044 ;
  assign n13838 = n4496 & n5065 ;
  assign n13839 = n3579 & n13838 ;
  assign n13840 = n13839 ^ n452 ^ 1'b0 ;
  assign n13841 = ~n829 & n13840 ;
  assign n13842 = ( n9822 & n13837 ) | ( n9822 & n13841 ) | ( n13837 & n13841 ) ;
  assign n13843 = n13842 ^ n9387 ^ n5446 ;
  assign n13844 = n4541 | n9116 ;
  assign n13845 = ~n2440 & n13844 ;
  assign n13846 = n13845 ^ n8570 ^ n8534 ;
  assign n13847 = n13846 ^ n7330 ^ n2053 ;
  assign n13848 = ( n9342 & n10151 ) | ( n9342 & n11343 ) | ( n10151 & n11343 ) ;
  assign n13849 = n13848 ^ n5086 ^ 1'b0 ;
  assign n13850 = n8662 ^ n1887 ^ 1'b0 ;
  assign n13851 = ~n7836 & n13850 ;
  assign n13852 = n13851 ^ n5865 ^ n488 ;
  assign n13853 = n4370 | n5248 ;
  assign n13854 = n13853 ^ n5205 ^ 1'b0 ;
  assign n13855 = n13854 ^ n3706 ^ 1'b0 ;
  assign n13856 = ~n5464 & n12443 ;
  assign n13857 = n13856 ^ n13449 ^ n9651 ;
  assign n13858 = n10459 & ~n13835 ;
  assign n13859 = n1369 & n2363 ;
  assign n13860 = ~n2357 & n13859 ;
  assign n13861 = ~n2226 & n5963 ;
  assign n13862 = n13860 & n13861 ;
  assign n13863 = ( ~n2658 & n11872 ) | ( ~n2658 & n13862 ) | ( n11872 & n13862 ) ;
  assign n13864 = ( ~n3274 & n11774 ) | ( ~n3274 & n13863 ) | ( n11774 & n13863 ) ;
  assign n13865 = n8711 ^ n4773 ^ n3683 ;
  assign n13866 = n6198 ^ n1324 ^ 1'b0 ;
  assign n13867 = n2045 | n13866 ;
  assign n13868 = n4697 ^ n4172 ^ 1'b0 ;
  assign n13869 = ( n6142 & n13867 ) | ( n6142 & n13868 ) | ( n13867 & n13868 ) ;
  assign n13871 = n2799 ^ n2553 ^ n2102 ;
  assign n13870 = ~n1519 & n3745 ;
  assign n13872 = n13871 ^ n13870 ^ 1'b0 ;
  assign n13873 = ( n1421 & n6929 ) | ( n1421 & ~n9677 ) | ( n6929 & ~n9677 ) ;
  assign n13874 = n13873 ^ n2834 ^ 1'b0 ;
  assign n13875 = ~n6274 & n13874 ;
  assign n13876 = n13875 ^ n6320 ^ 1'b0 ;
  assign n13877 = n2593 | n10301 ;
  assign n13878 = n13877 ^ n2108 ^ 1'b0 ;
  assign n13879 = n13296 ^ n10811 ^ n6858 ;
  assign n13880 = ( ~n5853 & n13878 ) | ( ~n5853 & n13879 ) | ( n13878 & n13879 ) ;
  assign n13881 = n738 | n2606 ;
  assign n13882 = n2826 | n13881 ;
  assign n13883 = n2089 & n13882 ;
  assign n13884 = n13883 ^ n7156 ^ 1'b0 ;
  assign n13885 = n8790 & ~n9966 ;
  assign n13886 = n13885 ^ n13321 ^ 1'b0 ;
  assign n13887 = ~n10667 & n13886 ;
  assign n13888 = n8688 ^ n5472 ^ 1'b0 ;
  assign n13889 = n8416 | n13888 ;
  assign n13890 = n7780 | n9851 ;
  assign n13891 = ( n9319 & n13194 ) | ( n9319 & ~n13890 ) | ( n13194 & ~n13890 ) ;
  assign n13892 = n8915 ^ n5409 ^ 1'b0 ;
  assign n13896 = n4688 ^ n4294 ^ n2733 ;
  assign n13897 = n13896 ^ n957 ^ 1'b0 ;
  assign n13898 = n2902 & ~n13897 ;
  assign n13893 = n3804 ^ n1149 ^ n1024 ;
  assign n13894 = ( n2212 & ~n11908 ) | ( n2212 & n13893 ) | ( ~n11908 & n13893 ) ;
  assign n13895 = n13894 ^ n4811 ^ n2864 ;
  assign n13899 = n13898 ^ n13895 ^ n10645 ;
  assign n13900 = ( ~n4408 & n4751 ) | ( ~n4408 & n5695 ) | ( n4751 & n5695 ) ;
  assign n13901 = ~n4805 & n13900 ;
  assign n13902 = n1500 & ~n12598 ;
  assign n13903 = ( n12035 & ~n13901 ) | ( n12035 & n13902 ) | ( ~n13901 & n13902 ) ;
  assign n13904 = n969 & ~n4202 ;
  assign n13905 = n7015 | n13904 ;
  assign n13906 = n12750 ^ n7655 ^ n7010 ;
  assign n13907 = n13906 ^ n11794 ^ n7024 ;
  assign n13908 = n12768 ^ n6008 ^ 1'b0 ;
  assign n13909 = ~n2245 & n13908 ;
  assign n13911 = n9452 ^ x113 ^ 1'b0 ;
  assign n13912 = ~n10947 & n13911 ;
  assign n13910 = n2357 ^ n2128 ^ 1'b0 ;
  assign n13913 = n13912 ^ n13910 ^ n11534 ;
  assign n13914 = n5335 | n10634 ;
  assign n13916 = ( n3278 & n3925 ) | ( n3278 & n13554 ) | ( n3925 & n13554 ) ;
  assign n13915 = ~n1750 & n11040 ;
  assign n13917 = n13916 ^ n13915 ^ 1'b0 ;
  assign n13918 = ( n5675 & n13914 ) | ( n5675 & n13917 ) | ( n13914 & n13917 ) ;
  assign n13919 = n4793 ^ n4134 ^ n553 ;
  assign n13920 = ( n5763 & ~n9627 ) | ( n5763 & n13919 ) | ( ~n9627 & n13919 ) ;
  assign n13921 = n5144 & n9856 ;
  assign n13922 = n13921 ^ n233 ^ 1'b0 ;
  assign n13923 = ( n7789 & n13920 ) | ( n7789 & n13922 ) | ( n13920 & n13922 ) ;
  assign n13924 = n6842 ^ n3649 ^ n1828 ;
  assign n13925 = n8680 ^ n5863 ^ 1'b0 ;
  assign n13926 = n4092 ^ n2900 ^ n2037 ;
  assign n13927 = ( ~n6881 & n8802 ) | ( ~n6881 & n13926 ) | ( n8802 & n13926 ) ;
  assign n13928 = n13927 ^ n6575 ^ n6235 ;
  assign n13929 = ( n4713 & ~n13925 ) | ( n4713 & n13928 ) | ( ~n13925 & n13928 ) ;
  assign n13930 = n10220 ^ n8001 ^ 1'b0 ;
  assign n13934 = n13327 ^ n359 ^ 1'b0 ;
  assign n13931 = n13708 ^ x70 ^ 1'b0 ;
  assign n13932 = n13931 ^ n12895 ^ 1'b0 ;
  assign n13933 = n6899 & n13932 ;
  assign n13935 = n13934 ^ n13933 ^ 1'b0 ;
  assign n13936 = n1793 & ~n9125 ;
  assign n13937 = n2147 | n2799 ;
  assign n13938 = n6646 ^ n1188 ^ 1'b0 ;
  assign n13939 = ( n3965 & ~n11947 ) | ( n3965 & n13938 ) | ( ~n11947 & n13938 ) ;
  assign n13940 = ~n13937 & n13939 ;
  assign n13941 = ~n3049 & n13940 ;
  assign n13942 = n2159 & ~n8592 ;
  assign n13943 = n13942 ^ n5562 ^ 1'b0 ;
  assign n13944 = ( ~n4849 & n7270 ) | ( ~n4849 & n7471 ) | ( n7270 & n7471 ) ;
  assign n13945 = ( ~n5312 & n13146 ) | ( ~n5312 & n13944 ) | ( n13146 & n13944 ) ;
  assign n13946 = ( ~n2122 & n6945 ) | ( ~n2122 & n11239 ) | ( n6945 & n11239 ) ;
  assign n13947 = n13206 & n13946 ;
  assign n13948 = ( ~n7478 & n8697 ) | ( ~n7478 & n13947 ) | ( n8697 & n13947 ) ;
  assign n13949 = n13948 ^ n7529 ^ n4861 ;
  assign n13950 = n12693 ^ n783 ^ n323 ;
  assign n13951 = n13950 ^ n2583 ^ 1'b0 ;
  assign n13952 = n2042 | n7423 ;
  assign n13953 = n2534 | n13952 ;
  assign n13954 = ( x101 & n242 ) | ( x101 & ~n10742 ) | ( n242 & ~n10742 ) ;
  assign n13955 = ( n9219 & ~n13953 ) | ( n9219 & n13954 ) | ( ~n13953 & n13954 ) ;
  assign n13956 = ~n2198 & n12914 ;
  assign n13957 = ~n11961 & n13956 ;
  assign n13958 = ( n1394 & n7553 ) | ( n1394 & n9741 ) | ( n7553 & n9741 ) ;
  assign n13959 = ( n1834 & n3770 ) | ( n1834 & ~n5689 ) | ( n3770 & ~n5689 ) ;
  assign n13960 = n2603 & n7880 ;
  assign n13961 = ~n13959 & n13960 ;
  assign n13966 = n7046 ^ n6646 ^ n1648 ;
  assign n13967 = ( n7897 & ~n10301 ) | ( n7897 & n13966 ) | ( ~n10301 & n13966 ) ;
  assign n13962 = n1704 ^ n576 ^ 1'b0 ;
  assign n13963 = n10061 & n12255 ;
  assign n13964 = ( n6938 & ~n13962 ) | ( n6938 & n13963 ) | ( ~n13962 & n13963 ) ;
  assign n13965 = ~n10489 & n13964 ;
  assign n13968 = n13967 ^ n13965 ^ 1'b0 ;
  assign n13969 = n7583 & n13968 ;
  assign n13970 = n13969 ^ n7550 ^ 1'b0 ;
  assign n13971 = n13961 | n13970 ;
  assign n13972 = n7116 & ~n9042 ;
  assign n13973 = n13972 ^ n6017 ^ 1'b0 ;
  assign n13976 = n5030 ^ n4426 ^ n3877 ;
  assign n13974 = ( n5867 & ~n11300 ) | ( n5867 & n12186 ) | ( ~n11300 & n12186 ) ;
  assign n13975 = n11669 | n13974 ;
  assign n13977 = n13976 ^ n13975 ^ 1'b0 ;
  assign n13978 = n7082 ^ n6004 ^ n4353 ;
  assign n13979 = x27 & ~n5669 ;
  assign n13980 = n13979 ^ n2580 ^ 1'b0 ;
  assign n13981 = n171 | n1381 ;
  assign n13982 = ( n11396 & n13980 ) | ( n11396 & n13981 ) | ( n13980 & n13981 ) ;
  assign n13989 = n12585 ^ n4235 ^ 1'b0 ;
  assign n13990 = ( n6546 & n8132 ) | ( n6546 & n13989 ) | ( n8132 & n13989 ) ;
  assign n13985 = x23 & ~n4712 ;
  assign n13986 = ~n3720 & n13985 ;
  assign n13983 = ~n263 & n803 ;
  assign n13984 = ( n523 & ~n7320 ) | ( n523 & n13983 ) | ( ~n7320 & n13983 ) ;
  assign n13987 = n13986 ^ n13984 ^ n8553 ;
  assign n13988 = n12374 & n13987 ;
  assign n13991 = n13990 ^ n13988 ^ 1'b0 ;
  assign n13992 = n1943 ^ n731 ^ 1'b0 ;
  assign n13993 = n13992 ^ n11429 ^ n3450 ;
  assign n13994 = n13993 ^ n6093 ^ n5865 ;
  assign n13995 = n440 & n854 ;
  assign n13996 = n13994 | n13995 ;
  assign n13997 = n2931 ^ n1860 ^ 1'b0 ;
  assign n13998 = n153 & n13997 ;
  assign n13999 = n3716 & n4737 ;
  assign n14000 = n9409 ^ n8260 ^ n6208 ;
  assign n14001 = ( n4555 & ~n5917 ) | ( n4555 & n8998 ) | ( ~n5917 & n8998 ) ;
  assign n14006 = n3318 ^ n3045 ^ 1'b0 ;
  assign n14007 = ~n2100 & n14006 ;
  assign n14002 = ( n239 & n2696 ) | ( n239 & ~n3284 ) | ( n2696 & ~n3284 ) ;
  assign n14003 = n10459 | n14002 ;
  assign n14004 = n14003 ^ n1387 ^ 1'b0 ;
  assign n14005 = n6039 | n14004 ;
  assign n14008 = n14007 ^ n14005 ^ 1'b0 ;
  assign n14009 = n7477 | n14008 ;
  assign n14010 = n863 ^ n664 ^ n185 ;
  assign n14011 = ( n5983 & ~n12279 ) | ( n5983 & n14010 ) | ( ~n12279 & n14010 ) ;
  assign n14012 = n14011 ^ n4128 ^ n141 ;
  assign n14013 = n8693 ^ n8096 ^ n3481 ;
  assign n14014 = ( n9369 & n9695 ) | ( n9369 & n14013 ) | ( n9695 & n14013 ) ;
  assign n14015 = n8065 ^ n6738 ^ 1'b0 ;
  assign n14016 = n2026 | n14015 ;
  assign n14017 = n14016 ^ n4567 ^ n2171 ;
  assign n14018 = ( n6172 & n8424 ) | ( n6172 & ~n14017 ) | ( n8424 & ~n14017 ) ;
  assign n14019 = n14018 ^ n7581 ^ 1'b0 ;
  assign n14020 = ~n433 & n969 ;
  assign n14021 = ~n11024 & n14020 ;
  assign n14022 = n10216 ^ n5147 ^ 1'b0 ;
  assign n14023 = ~n14021 & n14022 ;
  assign n14024 = ( n730 & n6176 ) | ( n730 & n7588 ) | ( n6176 & n7588 ) ;
  assign n14025 = ( n5661 & n13210 ) | ( n5661 & ~n14024 ) | ( n13210 & ~n14024 ) ;
  assign n14026 = n792 & n14025 ;
  assign n14027 = n13197 & n14026 ;
  assign n14028 = ~n4578 & n6049 ;
  assign n14029 = n2926 & n14028 ;
  assign n14030 = n11958 & n12738 ;
  assign n14031 = ( n5011 & n14029 ) | ( n5011 & n14030 ) | ( n14029 & n14030 ) ;
  assign n14032 = ( ~n6881 & n7890 ) | ( ~n6881 & n8947 ) | ( n7890 & n8947 ) ;
  assign n14033 = n14032 ^ n6466 ^ 1'b0 ;
  assign n14034 = ~n4334 & n14033 ;
  assign n14035 = n5281 & ~n13259 ;
  assign n14036 = n14035 ^ n6814 ^ 1'b0 ;
  assign n14037 = ~n14034 & n14036 ;
  assign n14038 = n995 ^ n490 ^ 1'b0 ;
  assign n14039 = n14038 ^ n7676 ^ 1'b0 ;
  assign n14040 = ~n1926 & n14039 ;
  assign n14041 = n9080 & n14040 ;
  assign n14042 = n14041 ^ n7425 ^ 1'b0 ;
  assign n14045 = n3964 ^ n3750 ^ n3385 ;
  assign n14046 = ( n3716 & n4931 ) | ( n3716 & n14045 ) | ( n4931 & n14045 ) ;
  assign n14043 = ( ~n3240 & n7215 ) | ( ~n3240 & n9451 ) | ( n7215 & n9451 ) ;
  assign n14044 = ( ~n8161 & n10895 ) | ( ~n8161 & n14043 ) | ( n10895 & n14043 ) ;
  assign n14047 = n14046 ^ n14044 ^ 1'b0 ;
  assign n14049 = n13708 ^ n11091 ^ 1'b0 ;
  assign n14050 = ~n1802 & n14049 ;
  assign n14051 = ( ~n5792 & n5889 ) | ( ~n5792 & n14050 ) | ( n5889 & n14050 ) ;
  assign n14048 = n9067 & n13802 ;
  assign n14052 = n14051 ^ n14048 ^ 1'b0 ;
  assign n14053 = n9125 ^ n3666 ^ 1'b0 ;
  assign n14054 = ( n943 & n13240 ) | ( n943 & n14053 ) | ( n13240 & n14053 ) ;
  assign n14055 = n4290 ^ x32 ^ 1'b0 ;
  assign n14056 = n1663 & n14055 ;
  assign n14057 = n14056 ^ n5542 ^ 1'b0 ;
  assign n14058 = n14057 ^ n3088 ^ 1'b0 ;
  assign n14059 = n12856 & ~n14058 ;
  assign n14060 = n5166 | n6160 ;
  assign n14061 = n886 | n12130 ;
  assign n14062 = n14061 ^ n9588 ^ 1'b0 ;
  assign n14063 = ~n14060 & n14062 ;
  assign n14072 = n12502 ^ n7096 ^ n2399 ;
  assign n14073 = n14072 ^ n2216 ^ 1'b0 ;
  assign n14070 = n444 & n5738 ;
  assign n14064 = ( n265 & n7580 ) | ( n265 & ~n7765 ) | ( n7580 & ~n7765 ) ;
  assign n14065 = ( n598 & n11703 ) | ( n598 & n14064 ) | ( n11703 & n14064 ) ;
  assign n14066 = n203 & ~n6927 ;
  assign n14067 = ( n6941 & ~n14065 ) | ( n6941 & n14066 ) | ( ~n14065 & n14066 ) ;
  assign n14068 = n14067 ^ n5915 ^ 1'b0 ;
  assign n14069 = n8334 & ~n14068 ;
  assign n14071 = n14070 ^ n14069 ^ n10518 ;
  assign n14074 = n14073 ^ n14071 ^ 1'b0 ;
  assign n14075 = n3645 | n14074 ;
  assign n14076 = n6580 ^ n1757 ^ 1'b0 ;
  assign n14077 = n9246 ^ n6910 ^ n961 ;
  assign n14078 = n10359 ^ n2862 ^ 1'b0 ;
  assign n14080 = ( n6494 & ~n7961 ) | ( n6494 & n8103 ) | ( ~n7961 & n8103 ) ;
  assign n14079 = ~n4453 & n9660 ;
  assign n14081 = n14080 ^ n14079 ^ 1'b0 ;
  assign n14082 = ( n2582 & ~n14078 ) | ( n2582 & n14081 ) | ( ~n14078 & n14081 ) ;
  assign n14083 = ~n14077 & n14082 ;
  assign n14084 = n4568 & n14083 ;
  assign n14085 = n5469 & ~n8915 ;
  assign n14086 = n8730 | n8957 ;
  assign n14096 = ( n2378 & n2911 ) | ( n2378 & ~n5461 ) | ( n2911 & ~n5461 ) ;
  assign n14087 = n8281 & ~n10367 ;
  assign n14090 = n2500 ^ n550 ^ n428 ;
  assign n14091 = n4188 & n14090 ;
  assign n14092 = ~n9446 & n14091 ;
  assign n14088 = n10237 & ~n13105 ;
  assign n14089 = n14088 ^ n6320 ^ 1'b0 ;
  assign n14093 = n14092 ^ n14089 ^ n7705 ;
  assign n14094 = n14093 ^ n5385 ^ n1908 ;
  assign n14095 = ~n14087 & n14094 ;
  assign n14097 = n14096 ^ n14095 ^ 1'b0 ;
  assign n14098 = ( n824 & n1146 ) | ( n824 & ~n6805 ) | ( n1146 & ~n6805 ) ;
  assign n14099 = n14097 & n14098 ;
  assign n14100 = n14099 ^ n8584 ^ 1'b0 ;
  assign n14101 = n2860 ^ n577 ^ 1'b0 ;
  assign n14102 = n8902 & n14101 ;
  assign n14103 = n14102 ^ n11609 ^ 1'b0 ;
  assign n14104 = n5867 | n9183 ;
  assign n14105 = n5594 | n14104 ;
  assign n14106 = n1243 | n4747 ;
  assign n14107 = n14106 ^ n4189 ^ 1'b0 ;
  assign n14108 = ~n9567 & n14107 ;
  assign n14109 = n14108 ^ n5010 ^ 1'b0 ;
  assign n14110 = n14109 ^ n9866 ^ n6644 ;
  assign n14111 = ( n1594 & ~n8157 ) | ( n1594 & n14110 ) | ( ~n8157 & n14110 ) ;
  assign n14113 = n1867 & ~n2625 ;
  assign n14114 = n14113 ^ n4887 ^ 1'b0 ;
  assign n14112 = n1991 & n7770 ;
  assign n14115 = n14114 ^ n14112 ^ 1'b0 ;
  assign n14116 = ( ~n9679 & n10132 ) | ( ~n9679 & n14115 ) | ( n10132 & n14115 ) ;
  assign n14117 = n12739 & ~n14116 ;
  assign n14118 = n14117 ^ n8791 ^ 1'b0 ;
  assign n14119 = ( n7032 & ~n14111 ) | ( n7032 & n14118 ) | ( ~n14111 & n14118 ) ;
  assign n14120 = n14119 ^ n2700 ^ 1'b0 ;
  assign n14121 = n8783 & ~n12343 ;
  assign n14122 = n4588 & n14121 ;
  assign n14123 = n1055 & ~n11731 ;
  assign n14124 = ~n13599 & n14123 ;
  assign n14125 = ( n8881 & n9267 ) | ( n8881 & ~n14124 ) | ( n9267 & ~n14124 ) ;
  assign n14126 = n2772 & ~n3243 ;
  assign n14127 = n5765 & n14126 ;
  assign n14128 = ~n365 & n7465 ;
  assign n14129 = n10809 ^ n1184 ^ 1'b0 ;
  assign n14130 = n1303 & ~n14129 ;
  assign n14131 = ~n10142 & n10663 ;
  assign n14132 = ~n14130 & n14131 ;
  assign n14133 = n9567 | n14132 ;
  assign n14134 = n10309 ^ x75 ^ 1'b0 ;
  assign n14135 = n14134 ^ n4280 ^ 1'b0 ;
  assign n14136 = ~n5776 & n14135 ;
  assign n14137 = ( ~n5051 & n13563 ) | ( ~n5051 & n14136 ) | ( n13563 & n14136 ) ;
  assign n14138 = n6793 ^ n5364 ^ 1'b0 ;
  assign n14139 = ( n760 & ~n811 ) | ( n760 & n14138 ) | ( ~n811 & n14138 ) ;
  assign n14140 = ( n4022 & n11852 ) | ( n4022 & n14139 ) | ( n11852 & n14139 ) ;
  assign n14141 = n3389 & ~n10228 ;
  assign n14142 = ( ~n1647 & n4640 ) | ( ~n1647 & n5102 ) | ( n4640 & n5102 ) ;
  assign n14143 = ( n969 & n8885 ) | ( n969 & ~n14142 ) | ( n8885 & ~n14142 ) ;
  assign n14144 = n11628 ^ n1619 ^ 1'b0 ;
  assign n14145 = n3193 & ~n5248 ;
  assign n14146 = n5011 ^ n4052 ^ n284 ;
  assign n14147 = n6863 & n13530 ;
  assign n14148 = n7884 & n14147 ;
  assign n14149 = n8677 & n14148 ;
  assign n14150 = ( n4889 & ~n14146 ) | ( n4889 & n14149 ) | ( ~n14146 & n14149 ) ;
  assign n14151 = n250 | n8975 ;
  assign n14152 = ( n3929 & n5691 ) | ( n3929 & n12739 ) | ( n5691 & n12739 ) ;
  assign n14153 = n14152 ^ n1717 ^ 1'b0 ;
  assign n14154 = n2880 & ~n14153 ;
  assign n14155 = n9860 & n14154 ;
  assign n14156 = ~n1955 & n6014 ;
  assign n14157 = ~n3531 & n14156 ;
  assign n14158 = n10348 ^ n2509 ^ 1'b0 ;
  assign n14159 = ( ~n243 & n3688 ) | ( ~n243 & n14158 ) | ( n3688 & n14158 ) ;
  assign n14160 = n14159 ^ n12031 ^ 1'b0 ;
  assign n14161 = ~n14157 & n14160 ;
  assign n14162 = ( ~x45 & n3183 ) | ( ~x45 & n3673 ) | ( n3183 & n3673 ) ;
  assign n14163 = n14162 ^ n7412 ^ n325 ;
  assign n14164 = n6261 ^ n4652 ^ n1911 ;
  assign n14165 = n13552 ^ n3377 ^ 1'b0 ;
  assign n14166 = n7378 ^ n2750 ^ 1'b0 ;
  assign n14167 = ( n2673 & n2731 ) | ( n2673 & ~n6595 ) | ( n2731 & ~n6595 ) ;
  assign n14168 = n13036 ^ n5988 ^ n4196 ;
  assign n14169 = n14168 ^ n13459 ^ n9674 ;
  assign n14170 = ( n12895 & n13891 ) | ( n12895 & n14169 ) | ( n13891 & n14169 ) ;
  assign n14171 = ( n1629 & n6881 ) | ( n1629 & n12155 ) | ( n6881 & n12155 ) ;
  assign n14172 = n6005 & n14171 ;
  assign n14173 = n14172 ^ n11828 ^ n3180 ;
  assign n14174 = ( ~n6937 & n9138 ) | ( ~n6937 & n14173 ) | ( n9138 & n14173 ) ;
  assign n14175 = n13212 ^ n2959 ^ x103 ;
  assign n14176 = n14175 ^ n9958 ^ 1'b0 ;
  assign n14177 = ( n967 & ~n5238 ) | ( n967 & n12847 ) | ( ~n5238 & n12847 ) ;
  assign n14178 = n9790 ^ n7741 ^ n7408 ;
  assign n14179 = n14178 ^ n9020 ^ 1'b0 ;
  assign n14180 = n8495 & ~n14179 ;
  assign n14181 = ( n9758 & n12121 ) | ( n9758 & n14180 ) | ( n12121 & n14180 ) ;
  assign n14182 = n7006 ^ n6102 ^ 1'b0 ;
  assign n14183 = n12512 | n14182 ;
  assign n14184 = n14183 ^ n14063 ^ n5059 ;
  assign n14185 = ~n184 & n4560 ;
  assign n14186 = n6984 ^ n6691 ^ n1442 ;
  assign n14187 = ~n14185 & n14186 ;
  assign n14188 = n14187 ^ n2802 ^ 1'b0 ;
  assign n14189 = ( n11118 & n13676 ) | ( n11118 & ~n14188 ) | ( n13676 & ~n14188 ) ;
  assign n14190 = n6558 ^ x47 ^ 1'b0 ;
  assign n14191 = ~n483 & n14190 ;
  assign n14192 = n6920 & n10368 ;
  assign n14193 = n14192 ^ n4822 ^ 1'b0 ;
  assign n14194 = n14191 & ~n14193 ;
  assign n14195 = n14194 ^ n2539 ^ 1'b0 ;
  assign n14196 = ( ~n6257 & n13841 ) | ( ~n6257 & n14195 ) | ( n13841 & n14195 ) ;
  assign n14198 = n1900 ^ n1395 ^ 1'b0 ;
  assign n14197 = ( ~n150 & n2866 ) | ( ~n150 & n5815 ) | ( n2866 & n5815 ) ;
  assign n14199 = n14198 ^ n14197 ^ 1'b0 ;
  assign n14200 = n14199 ^ n11771 ^ n1984 ;
  assign n14201 = n2378 & ~n14200 ;
  assign n14202 = n14201 ^ n13737 ^ 1'b0 ;
  assign n14203 = n9786 ^ n8186 ^ n2638 ;
  assign n14204 = n8219 ^ n2820 ^ 1'b0 ;
  assign n14211 = n7932 ^ n311 ^ 1'b0 ;
  assign n14209 = n7665 ^ n2082 ^ 1'b0 ;
  assign n14210 = ~n2226 & n14209 ;
  assign n14205 = ( ~n2911 & n8239 ) | ( ~n2911 & n8459 ) | ( n8239 & n8459 ) ;
  assign n14206 = ( ~n4553 & n8268 ) | ( ~n4553 & n14205 ) | ( n8268 & n14205 ) ;
  assign n14207 = n10218 ^ n2346 ^ 1'b0 ;
  assign n14208 = n14206 & n14207 ;
  assign n14212 = n14211 ^ n14210 ^ n14208 ;
  assign n14213 = n270 | n10655 ;
  assign n14214 = n14213 ^ n2530 ^ 1'b0 ;
  assign n14215 = n14214 ^ n9691 ^ n7929 ;
  assign n14216 = n2016 & ~n7176 ;
  assign n14217 = n14216 ^ x12 ^ 1'b0 ;
  assign n14218 = n7067 ^ n3561 ^ n1391 ;
  assign n14219 = n1565 & n8562 ;
  assign n14220 = n11630 ^ n3628 ^ 1'b0 ;
  assign n14223 = n2112 & n5324 ;
  assign n14224 = n14223 ^ n3044 ^ 1'b0 ;
  assign n14225 = n1722 & n14224 ;
  assign n14226 = ( n1739 & n3131 ) | ( n1739 & ~n14225 ) | ( n3131 & ~n14225 ) ;
  assign n14227 = ~n5301 & n14226 ;
  assign n14221 = ( ~n1434 & n4497 ) | ( ~n1434 & n6746 ) | ( n4497 & n6746 ) ;
  assign n14222 = n14221 ^ n7361 ^ 1'b0 ;
  assign n14228 = n14227 ^ n14222 ^ n6781 ;
  assign n14229 = ~n308 & n14228 ;
  assign n14233 = n5602 ^ n2291 ^ 1'b0 ;
  assign n14234 = n14233 ^ n5374 ^ 1'b0 ;
  assign n14235 = n7729 | n14234 ;
  assign n14230 = n4289 ^ n1980 ^ 1'b0 ;
  assign n14231 = ~n3061 & n14230 ;
  assign n14232 = ( n3253 & n7278 ) | ( n3253 & ~n14231 ) | ( n7278 & ~n14231 ) ;
  assign n14236 = n14235 ^ n14232 ^ n12202 ;
  assign n14237 = n6612 ^ n4331 ^ 1'b0 ;
  assign n14238 = n12571 ^ n8426 ^ n5419 ;
  assign n14239 = ( n767 & n3275 ) | ( n767 & n14238 ) | ( n3275 & n14238 ) ;
  assign n14240 = ( n538 & n2120 ) | ( n538 & ~n9082 ) | ( n2120 & ~n9082 ) ;
  assign n14241 = n14240 ^ n12071 ^ 1'b0 ;
  assign n14242 = n4438 | n14241 ;
  assign n14243 = ( ~n420 & n3227 ) | ( ~n420 & n12827 ) | ( n3227 & n12827 ) ;
  assign n14244 = n10991 ^ n4500 ^ 1'b0 ;
  assign n14245 = n14244 ^ n2544 ^ 1'b0 ;
  assign n14246 = ~n14243 & n14245 ;
  assign n14247 = n5507 ^ n2914 ^ 1'b0 ;
  assign n14248 = n14247 ^ n7930 ^ 1'b0 ;
  assign n14249 = n2230 & n14248 ;
  assign n14250 = n14249 ^ n10965 ^ 1'b0 ;
  assign n14251 = ( n3654 & n8604 ) | ( n3654 & ~n10323 ) | ( n8604 & ~n10323 ) ;
  assign n14252 = n14251 ^ n9793 ^ 1'b0 ;
  assign n14253 = n14250 & ~n14252 ;
  assign n14254 = n7024 ^ n4248 ^ n3787 ;
  assign n14255 = ~n3051 & n4036 ;
  assign n14256 = n9238 & ~n14255 ;
  assign n14257 = ~n8546 & n14256 ;
  assign n14258 = n2199 | n13517 ;
  assign n14259 = n14258 ^ n4146 ^ 1'b0 ;
  assign n14260 = n9544 ^ n6462 ^ 1'b0 ;
  assign n14261 = ( n969 & ~n6840 ) | ( n969 & n12914 ) | ( ~n6840 & n12914 ) ;
  assign n14262 = ( n2002 & ~n12093 ) | ( n2002 & n14261 ) | ( ~n12093 & n14261 ) ;
  assign n14263 = ~n8749 & n14262 ;
  assign n14264 = n3135 ^ x27 ^ 1'b0 ;
  assign n14265 = ~n3232 & n14264 ;
  assign n14266 = n5947 & n14265 ;
  assign n14267 = ~n4292 & n14266 ;
  assign n14268 = ~n607 & n14267 ;
  assign n14269 = ( n7785 & n8649 ) | ( n7785 & n14268 ) | ( n8649 & n14268 ) ;
  assign n14271 = n11268 ^ n8729 ^ 1'b0 ;
  assign n14270 = ~n9048 & n9134 ;
  assign n14272 = n14271 ^ n14270 ^ 1'b0 ;
  assign n14273 = n5911 | n13845 ;
  assign n14274 = n6072 & ~n14273 ;
  assign n14275 = n3490 ^ n1967 ^ 1'b0 ;
  assign n14276 = n12954 & n14275 ;
  assign n14277 = n14276 ^ n9890 ^ 1'b0 ;
  assign n14278 = ~n3416 & n13008 ;
  assign n14279 = ~n12669 & n14278 ;
  assign n14280 = n14279 ^ n9567 ^ n1655 ;
  assign n14281 = ( n3420 & n9251 ) | ( n3420 & n12907 ) | ( n9251 & n12907 ) ;
  assign n14282 = n194 & n4527 ;
  assign n14283 = ~x108 & n14282 ;
  assign n14284 = ( n11249 & n12053 ) | ( n11249 & n14283 ) | ( n12053 & n14283 ) ;
  assign n14285 = n4576 & n14284 ;
  assign n14286 = n10119 & n14285 ;
  assign n14287 = ~n2067 & n3776 ;
  assign n14288 = n14287 ^ n5259 ^ 1'b0 ;
  assign n14290 = n5865 & ~n9006 ;
  assign n14291 = n2011 ^ n500 ^ x33 ;
  assign n14292 = n14291 ^ n1285 ^ 1'b0 ;
  assign n14293 = n14290 | n14292 ;
  assign n14289 = n6965 & n9865 ;
  assign n14294 = n14293 ^ n14289 ^ 1'b0 ;
  assign n14295 = ~n325 & n14294 ;
  assign n14296 = n14295 ^ n4017 ^ 1'b0 ;
  assign n14297 = ( n3898 & n7073 ) | ( n3898 & n12811 ) | ( n7073 & n12811 ) ;
  assign n14298 = n8028 ^ n5934 ^ n203 ;
  assign n14299 = ( n1519 & n1920 ) | ( n1519 & n14298 ) | ( n1920 & n14298 ) ;
  assign n14300 = n12273 ^ n11682 ^ n6638 ;
  assign n14301 = n14300 ^ n896 ^ 1'b0 ;
  assign n14302 = ( n4868 & ~n8577 ) | ( n4868 & n14193 ) | ( ~n8577 & n14193 ) ;
  assign n14303 = n14302 ^ n10429 ^ 1'b0 ;
  assign n14304 = n14301 & ~n14303 ;
  assign n14305 = n8822 ^ n3706 ^ n2241 ;
  assign n14306 = n13896 & n14305 ;
  assign n14307 = n14306 ^ n13129 ^ 1'b0 ;
  assign n14308 = n8153 | n14307 ;
  assign n14309 = n1671 | n14308 ;
  assign n14310 = ( n14299 & n14304 ) | ( n14299 & ~n14309 ) | ( n14304 & ~n14309 ) ;
  assign n14311 = n7589 & ~n9679 ;
  assign n14312 = ~n1049 & n14311 ;
  assign n14313 = ( n1441 & ~n6710 ) | ( n1441 & n10481 ) | ( ~n6710 & n10481 ) ;
  assign n14314 = n5668 | n14313 ;
  assign n14315 = n12285 & ~n14314 ;
  assign n14316 = n10634 ^ n8129 ^ 1'b0 ;
  assign n14317 = n14316 ^ n8680 ^ 1'b0 ;
  assign n14318 = n5509 | n14317 ;
  assign n14319 = n760 & ~n3163 ;
  assign n14320 = n3599 & n7586 ;
  assign n14321 = n14320 ^ n12633 ^ 1'b0 ;
  assign n14327 = n4865 & n8003 ;
  assign n14328 = n14327 ^ n6240 ^ 1'b0 ;
  assign n14329 = n3607 | n14328 ;
  assign n14330 = n11055 & ~n14329 ;
  assign n14322 = n2950 ^ n1953 ^ 1'b0 ;
  assign n14323 = ~n3627 & n14322 ;
  assign n14324 = ( ~n831 & n5568 ) | ( ~n831 & n7774 ) | ( n5568 & n7774 ) ;
  assign n14325 = ( n445 & n13155 ) | ( n445 & n14324 ) | ( n13155 & n14324 ) ;
  assign n14326 = n14323 & ~n14325 ;
  assign n14331 = n14330 ^ n14326 ^ 1'b0 ;
  assign n14332 = n7116 ^ n4910 ^ n1649 ;
  assign n14333 = n13962 ^ n4639 ^ 1'b0 ;
  assign n14334 = n3819 | n14333 ;
  assign n14335 = n3789 & ~n14334 ;
  assign n14336 = ( ~x25 & n3354 ) | ( ~x25 & n14335 ) | ( n3354 & n14335 ) ;
  assign n14337 = n7020 ^ n433 ^ 1'b0 ;
  assign n14338 = n5699 ^ n2154 ^ 1'b0 ;
  assign n14339 = n641 & n14338 ;
  assign n14340 = n14339 ^ n5312 ^ n2562 ;
  assign n14341 = n2018 & ~n6230 ;
  assign n14342 = n14341 ^ n3004 ^ 1'b0 ;
  assign n14343 = n6372 ^ n664 ^ 1'b0 ;
  assign n14344 = n14343 ^ n11654 ^ n4863 ;
  assign n14345 = n14344 ^ n1724 ^ n214 ;
  assign n14346 = n14342 & ~n14345 ;
  assign n14356 = n3218 & n7889 ;
  assign n14357 = ~n5598 & n14356 ;
  assign n14358 = n14357 ^ n4650 ^ 1'b0 ;
  assign n14347 = n2161 ^ n2159 ^ n691 ;
  assign n14353 = ( ~n730 & n3369 ) | ( ~n730 & n3447 ) | ( n3369 & n3447 ) ;
  assign n14348 = n4086 ^ n691 ^ n174 ;
  assign n14349 = n7087 & ~n14348 ;
  assign n14350 = n14349 ^ n5238 ^ 1'b0 ;
  assign n14351 = n6373 & n10979 ;
  assign n14352 = ~n14350 & n14351 ;
  assign n14354 = n14353 ^ n14352 ^ 1'b0 ;
  assign n14355 = n14347 | n14354 ;
  assign n14359 = n14358 ^ n14355 ^ 1'b0 ;
  assign n14360 = n1154 ^ n263 ^ 1'b0 ;
  assign n14361 = n14360 ^ n1473 ^ n488 ;
  assign n14362 = ( n4568 & n7906 ) | ( n4568 & ~n14361 ) | ( n7906 & ~n14361 ) ;
  assign n14363 = n5454 ^ n2684 ^ 1'b0 ;
  assign n14364 = n3321 & ~n14363 ;
  assign n14365 = n14364 ^ n10287 ^ n4882 ;
  assign n14366 = ( n4214 & n12592 ) | ( n4214 & ~n14365 ) | ( n12592 & ~n14365 ) ;
  assign n14367 = n14366 ^ n4070 ^ 1'b0 ;
  assign n14368 = n13479 ^ n9695 ^ n888 ;
  assign n14369 = n13664 ^ n9411 ^ n3507 ;
  assign n14370 = n13755 ^ n10279 ^ n2077 ;
  assign n14371 = n6905 & ~n14370 ;
  assign n14372 = n14371 ^ n10051 ^ 1'b0 ;
  assign n14373 = n4486 | n12430 ;
  assign n14374 = n2811 & ~n14373 ;
  assign n14375 = n7001 & ~n14374 ;
  assign n14376 = n4773 ^ n1817 ^ 1'b0 ;
  assign n14377 = ~n5112 & n14376 ;
  assign n14378 = n5198 | n14377 ;
  assign n14379 = n14375 & ~n14378 ;
  assign n14380 = x86 & n956 ;
  assign n14381 = n9223 ^ n8207 ^ n2940 ;
  assign n14382 = ( n13986 & n14380 ) | ( n13986 & ~n14381 ) | ( n14380 & ~n14381 ) ;
  assign n14383 = ~n2726 & n4838 ;
  assign n14384 = ( n1698 & ~n11794 ) | ( n1698 & n14383 ) | ( ~n11794 & n14383 ) ;
  assign n14385 = n2323 | n9371 ;
  assign n14386 = n11524 & n14385 ;
  assign n14387 = n14386 ^ n2350 ^ 1'b0 ;
  assign n14388 = ( ~n8176 & n9704 ) | ( ~n8176 & n14387 ) | ( n9704 & n14387 ) ;
  assign n14389 = ( n964 & n4125 ) | ( n964 & ~n7166 ) | ( n4125 & ~n7166 ) ;
  assign n14390 = n4870 & n12051 ;
  assign n14391 = n14389 & n14390 ;
  assign n14392 = n14391 ^ n7780 ^ 1'b0 ;
  assign n14393 = ( ~n3236 & n14388 ) | ( ~n3236 & n14392 ) | ( n14388 & n14392 ) ;
  assign n14394 = n8204 ^ n5125 ^ 1'b0 ;
  assign n14395 = n2239 & n6790 ;
  assign n14396 = n14395 ^ n3402 ^ 1'b0 ;
  assign n14397 = n6476 ^ n1369 ^ n703 ;
  assign n14398 = ( n4701 & ~n14396 ) | ( n4701 & n14397 ) | ( ~n14396 & n14397 ) ;
  assign n14399 = n14398 ^ n13886 ^ n6945 ;
  assign n14400 = n3419 & n9843 ;
  assign n14401 = n14400 ^ n12010 ^ 1'b0 ;
  assign n14402 = n9584 ^ n8262 ^ n5513 ;
  assign n14403 = ( n678 & ~n2491 ) | ( n678 & n12715 ) | ( ~n2491 & n12715 ) ;
  assign n14404 = ( n2765 & n14402 ) | ( n2765 & ~n14403 ) | ( n14402 & ~n14403 ) ;
  assign n14405 = n14404 ^ n9112 ^ 1'b0 ;
  assign n14406 = n1232 & n14405 ;
  assign n14407 = n158 & ~n9440 ;
  assign n14408 = n2640 | n14407 ;
  assign n14409 = n6415 & ~n14408 ;
  assign n14410 = n3184 & n7256 ;
  assign n14411 = n14410 ^ n9186 ^ 1'b0 ;
  assign n14412 = n10565 ^ n4287 ^ 1'b0 ;
  assign n14413 = ( n11355 & n14411 ) | ( n11355 & ~n14412 ) | ( n14411 & ~n14412 ) ;
  assign n14414 = n1567 & ~n9935 ;
  assign n14415 = ( n3195 & n7927 ) | ( n3195 & ~n14414 ) | ( n7927 & ~n14414 ) ;
  assign n14416 = n14415 ^ n12436 ^ 1'b0 ;
  assign n14417 = n14413 & ~n14416 ;
  assign n14418 = ( ~n4065 & n5357 ) | ( ~n4065 & n8017 ) | ( n5357 & n8017 ) ;
  assign n14419 = n14418 ^ n6086 ^ n3591 ;
  assign n14420 = n566 | n3908 ;
  assign n14421 = n5253 & ~n14420 ;
  assign n14422 = n14419 & ~n14421 ;
  assign n14427 = n11830 ^ n10924 ^ 1'b0 ;
  assign n14428 = ( n9591 & n10084 ) | ( n9591 & ~n14427 ) | ( n10084 & ~n14427 ) ;
  assign n14423 = ( n4740 & ~n5055 ) | ( n4740 & n6019 ) | ( ~n5055 & n6019 ) ;
  assign n14424 = ( n3912 & n4130 ) | ( n3912 & ~n14423 ) | ( n4130 & ~n14423 ) ;
  assign n14425 = n14424 ^ n11409 ^ n2930 ;
  assign n14426 = n12684 | n14425 ;
  assign n14429 = n14428 ^ n14426 ^ 1'b0 ;
  assign n14430 = n9005 ^ n6010 ^ 1'b0 ;
  assign n14431 = n8690 ^ n5133 ^ n4878 ;
  assign n14432 = n8037 & ~n14431 ;
  assign n14433 = n4081 ^ n1191 ^ 1'b0 ;
  assign n14434 = n14433 ^ n11591 ^ 1'b0 ;
  assign n14435 = ~n5836 & n10230 ;
  assign n14436 = n7863 | n9499 ;
  assign n14437 = n3710 | n14436 ;
  assign n14438 = n14437 ^ n14174 ^ n3978 ;
  assign n14439 = n8855 ^ n8729 ^ n3104 ;
  assign n14440 = n8529 ^ n4713 ^ 1'b0 ;
  assign n14441 = n7371 | n14440 ;
  assign n14442 = n11942 ^ n2619 ^ x14 ;
  assign n14443 = ( n4450 & ~n14441 ) | ( n4450 & n14442 ) | ( ~n14441 & n14442 ) ;
  assign n14444 = n12847 ^ n7054 ^ 1'b0 ;
  assign n14446 = ( n8379 & n10567 ) | ( n8379 & ~n10911 ) | ( n10567 & ~n10911 ) ;
  assign n14445 = n11323 ^ n8191 ^ n6294 ;
  assign n14447 = n14446 ^ n14445 ^ 1'b0 ;
  assign n14448 = ~n8915 & n14447 ;
  assign n14449 = n159 & ~n14376 ;
  assign n14450 = n11839 | n12008 ;
  assign n14451 = n14450 ^ n11659 ^ 1'b0 ;
  assign n14452 = ( n3014 & n14449 ) | ( n3014 & ~n14451 ) | ( n14449 & ~n14451 ) ;
  assign n14453 = n7874 & ~n14452 ;
  assign n14454 = n14453 ^ n4948 ^ 1'b0 ;
  assign n14455 = n14454 ^ n8199 ^ n5920 ;
  assign n14456 = ( n1170 & ~n3924 ) | ( n1170 & n14455 ) | ( ~n3924 & n14455 ) ;
  assign n14457 = n13782 ^ n3111 ^ 1'b0 ;
  assign n14458 = n14457 ^ n11540 ^ n698 ;
  assign n14459 = n4730 | n13983 ;
  assign n14460 = n14459 ^ n10868 ^ 1'b0 ;
  assign n14461 = n6016 & n13554 ;
  assign n14462 = n14460 & n14461 ;
  assign n14463 = n3636 & ~n14462 ;
  assign n14464 = ~n3197 & n14463 ;
  assign n14465 = n3671 & ~n5461 ;
  assign n14466 = n14465 ^ n6112 ^ 1'b0 ;
  assign n14467 = n12366 | n14466 ;
  assign n14468 = n2373 & n13735 ;
  assign n14469 = n14468 ^ n7602 ^ 1'b0 ;
  assign n14470 = n14469 ^ n4455 ^ n1329 ;
  assign n14471 = n5785 ^ n3639 ^ 1'b0 ;
  assign n14472 = ~n5977 & n14471 ;
  assign n14473 = n14472 ^ n3354 ^ n3269 ;
  assign n14474 = ( n1019 & n7319 ) | ( n1019 & ~n14473 ) | ( n7319 & ~n14473 ) ;
  assign n14475 = n2319 | n11048 ;
  assign n14476 = n14475 ^ n3780 ^ 1'b0 ;
  assign n14477 = n14476 ^ n6594 ^ 1'b0 ;
  assign n14478 = n14477 ^ n7256 ^ 1'b0 ;
  assign n14479 = ~n5711 & n8981 ;
  assign n14480 = ( n10706 & n14478 ) | ( n10706 & n14479 ) | ( n14478 & n14479 ) ;
  assign n14482 = ( n641 & ~n1894 ) | ( n641 & n2955 ) | ( ~n1894 & n2955 ) ;
  assign n14483 = n6090 ^ n5462 ^ n2883 ;
  assign n14484 = ( n5802 & ~n14482 ) | ( n5802 & n14483 ) | ( ~n14482 & n14483 ) ;
  assign n14481 = ( ~n1605 & n2112 ) | ( ~n1605 & n4453 ) | ( n2112 & n4453 ) ;
  assign n14485 = n14484 ^ n14481 ^ n5740 ;
  assign n14486 = n10443 & n14485 ;
  assign n14487 = ~n2822 & n14486 ;
  assign n14488 = n7446 | n8672 ;
  assign n14489 = n7898 & ~n14488 ;
  assign n14492 = n6233 & n10678 ;
  assign n14493 = n14492 ^ n11400 ^ 1'b0 ;
  assign n14490 = n13248 ^ n10150 ^ 1'b0 ;
  assign n14491 = n3666 & ~n14490 ;
  assign n14494 = n14493 ^ n14491 ^ n13344 ;
  assign n14495 = n9195 ^ n2284 ^ n1814 ;
  assign n14496 = n14495 ^ n12582 ^ n9948 ;
  assign n14497 = n9518 ^ n1788 ^ 1'b0 ;
  assign n14498 = n3991 ^ n1411 ^ 1'b0 ;
  assign n14499 = x10 & ~n10568 ;
  assign n14500 = ( n7011 & n14498 ) | ( n7011 & n14499 ) | ( n14498 & n14499 ) ;
  assign n14503 = n4574 ^ n3823 ^ n3748 ;
  assign n14501 = ( n1071 & ~n3258 ) | ( n1071 & n5297 ) | ( ~n3258 & n5297 ) ;
  assign n14502 = n10513 & ~n14501 ;
  assign n14504 = n14503 ^ n14502 ^ 1'b0 ;
  assign n14505 = ( n4158 & n9010 ) | ( n4158 & ~n14504 ) | ( n9010 & ~n14504 ) ;
  assign n14506 = n14505 ^ n1896 ^ 1'b0 ;
  assign n14507 = n1192 | n13738 ;
  assign n14508 = n14418 & ~n14507 ;
  assign n14509 = n14508 ^ n13981 ^ n3212 ;
  assign n14510 = n3490 ^ n3203 ^ n379 ;
  assign n14511 = ( n1923 & ~n7628 ) | ( n1923 & n14510 ) | ( ~n7628 & n14510 ) ;
  assign n14512 = n3967 & n5389 ;
  assign n14513 = ~n14511 & n14512 ;
  assign n14514 = n5193 | n13127 ;
  assign n14515 = n14513 & ~n14514 ;
  assign n14516 = ( n1010 & n7087 ) | ( n1010 & ~n14515 ) | ( n7087 & ~n14515 ) ;
  assign n14517 = n3820 & ~n9364 ;
  assign n14518 = n9436 ^ n4150 ^ 1'b0 ;
  assign n14520 = n4556 ^ n3747 ^ n1468 ;
  assign n14521 = ( n170 & n981 ) | ( n170 & ~n14520 ) | ( n981 & ~n14520 ) ;
  assign n14519 = n10907 | n11596 ;
  assign n14522 = n14521 ^ n14519 ^ n13412 ;
  assign n14523 = ( ~n11213 & n12322 ) | ( ~n11213 & n14522 ) | ( n12322 & n14522 ) ;
  assign n14524 = n5669 & n13459 ;
  assign n14525 = n14078 ^ n2085 ^ 1'b0 ;
  assign n14526 = n14525 ^ n6596 ^ n2242 ;
  assign n14527 = ( n1785 & n8947 ) | ( n1785 & n10150 ) | ( n8947 & n10150 ) ;
  assign n14528 = n9925 ^ n4159 ^ n1364 ;
  assign n14531 = ~n2775 & n9033 ;
  assign n14529 = ~n5915 & n10114 ;
  assign n14530 = n821 & n14529 ;
  assign n14532 = n14531 ^ n14530 ^ n4539 ;
  assign n14533 = ~n450 & n5946 ;
  assign n14534 = n3629 | n14533 ;
  assign n14535 = n14534 ^ n11182 ^ 1'b0 ;
  assign n14536 = ~n2728 & n5890 ;
  assign n14537 = n5504 & n14536 ;
  assign n14538 = n14537 ^ n14220 ^ n12860 ;
  assign n14539 = ( ~n9364 & n10434 ) | ( ~n9364 & n13304 ) | ( n10434 & n13304 ) ;
  assign n14540 = n14539 ^ n11165 ^ n10699 ;
  assign n14541 = n14540 ^ n10569 ^ n2573 ;
  assign n14542 = n5297 ^ n3908 ^ x30 ;
  assign n14543 = n12650 & ~n14542 ;
  assign n14544 = n14543 ^ n760 ^ 1'b0 ;
  assign n14545 = ( n1002 & n1112 ) | ( n1002 & ~n4660 ) | ( n1112 & ~n4660 ) ;
  assign n14546 = n14545 ^ n8002 ^ 1'b0 ;
  assign n14547 = ~n14544 & n14546 ;
  assign n14548 = n5726 ^ n1561 ^ 1'b0 ;
  assign n14549 = ( n1160 & n3748 ) | ( n1160 & ~n14548 ) | ( n3748 & ~n14548 ) ;
  assign n14550 = n11052 | n14549 ;
  assign n14551 = n4249 & n10965 ;
  assign n14552 = n2881 & n14551 ;
  assign n14553 = n14552 ^ n9261 ^ 1'b0 ;
  assign n14554 = ( n2452 & n2589 ) | ( n2452 & ~n3481 ) | ( n2589 & ~n3481 ) ;
  assign n14555 = n14554 ^ n4943 ^ n1339 ;
  assign n14556 = n14555 ^ n11291 ^ n6865 ;
  assign n14565 = n2646 ^ n197 ^ 1'b0 ;
  assign n14557 = n5330 ^ n2935 ^ n1032 ;
  assign n14558 = n14557 ^ n9848 ^ n5765 ;
  assign n14559 = ( n5911 & n13755 ) | ( n5911 & n14558 ) | ( n13755 & n14558 ) ;
  assign n14560 = n7178 ^ n243 ^ 1'b0 ;
  assign n14561 = n7222 & n14560 ;
  assign n14562 = n14483 ^ n13739 ^ n9964 ;
  assign n14563 = ( ~n14559 & n14561 ) | ( ~n14559 & n14562 ) | ( n14561 & n14562 ) ;
  assign n14564 = n164 & n14563 ;
  assign n14566 = n14565 ^ n14564 ^ 1'b0 ;
  assign n14567 = n1316 | n3995 ;
  assign n14568 = n374 | n14567 ;
  assign n14569 = n10884 ^ n9173 ^ n3678 ;
  assign n14570 = n9902 | n14569 ;
  assign n14571 = n14568 & ~n14570 ;
  assign n14572 = n12329 ^ n9361 ^ n3609 ;
  assign n14573 = ( n3345 & n5691 ) | ( n3345 & n10344 ) | ( n5691 & n10344 ) ;
  assign n14574 = ( ~n533 & n11936 ) | ( ~n533 & n14573 ) | ( n11936 & n14573 ) ;
  assign n14575 = n14574 ^ n4475 ^ 1'b0 ;
  assign n14576 = n13933 ^ n8753 ^ n7765 ;
  assign n14577 = n1266 & n3973 ;
  assign n14578 = ( n2576 & ~n5179 ) | ( n2576 & n14577 ) | ( ~n5179 & n14577 ) ;
  assign n14579 = n14578 ^ n9000 ^ n1541 ;
  assign n14580 = n11500 ^ n1026 ^ 1'b0 ;
  assign n14581 = ( n3186 & n3381 ) | ( n3186 & n5242 ) | ( n3381 & n5242 ) ;
  assign n14582 = n14581 ^ n11396 ^ n7837 ;
  assign n14583 = n14582 ^ n10627 ^ 1'b0 ;
  assign n14584 = n14580 & ~n14583 ;
  assign n14585 = ( ~n6948 & n10974 ) | ( ~n6948 & n14584 ) | ( n10974 & n14584 ) ;
  assign n14586 = n5651 ^ n3488 ^ 1'b0 ;
  assign n14587 = ( n6221 & ~n8719 ) | ( n6221 & n14586 ) | ( ~n8719 & n14586 ) ;
  assign n14588 = n316 | n14587 ;
  assign n14589 = n8269 & ~n14588 ;
  assign n14590 = ~n3562 & n6537 ;
  assign n14591 = n6663 & ~n14590 ;
  assign n14592 = n14591 ^ n9322 ^ n8314 ;
  assign n14593 = n1668 | n13345 ;
  assign n14594 = n14592 | n14593 ;
  assign n14595 = n2365 | n14594 ;
  assign n14596 = n2204 | n10587 ;
  assign n14597 = ~n3965 & n14596 ;
  assign n14598 = n5225 & n13546 ;
  assign n14599 = n14598 ^ n10505 ^ 1'b0 ;
  assign n14600 = n2734 ^ n1903 ^ 1'b0 ;
  assign n14601 = n5680 ^ n5175 ^ n3207 ;
  assign n14602 = n3690 & n14601 ;
  assign n14603 = ( n5048 & n9582 ) | ( n5048 & ~n14602 ) | ( n9582 & ~n14602 ) ;
  assign n14604 = n4739 | n10963 ;
  assign n14605 = n14604 ^ n5308 ^ 1'b0 ;
  assign n14606 = n2537 | n14605 ;
  assign n14607 = n6656 ^ n4374 ^ 1'b0 ;
  assign n14608 = ( ~n217 & n14292 ) | ( ~n217 & n14607 ) | ( n14292 & n14607 ) ;
  assign n14609 = ~n2889 & n8553 ;
  assign n14610 = ~n10911 & n14609 ;
  assign n14611 = ( n4870 & n7626 ) | ( n4870 & ~n13974 ) | ( n7626 & ~n13974 ) ;
  assign n14613 = n3303 ^ n1783 ^ 1'b0 ;
  assign n14614 = ~n11276 & n14613 ;
  assign n14615 = n14614 ^ n7046 ^ n6134 ;
  assign n14616 = ( n1515 & ~n11433 ) | ( n1515 & n14615 ) | ( ~n11433 & n14615 ) ;
  assign n14612 = n11264 ^ n10110 ^ n1639 ;
  assign n14617 = n14616 ^ n14612 ^ 1'b0 ;
  assign n14618 = ( n365 & ~n5501 ) | ( n365 & n7792 ) | ( ~n5501 & n7792 ) ;
  assign n14619 = ( n3944 & ~n8728 ) | ( n3944 & n14618 ) | ( ~n8728 & n14618 ) ;
  assign n14620 = n5864 ^ n3826 ^ 1'b0 ;
  assign n14621 = n9155 & ~n9313 ;
  assign n14622 = n4247 & n14621 ;
  assign n14623 = n14622 ^ n8816 ^ 1'b0 ;
  assign n14624 = ( n392 & ~n2323 ) | ( n392 & n7843 ) | ( ~n2323 & n7843 ) ;
  assign n14625 = ~n600 & n12898 ;
  assign n14628 = n3991 & n8331 ;
  assign n14629 = ( n7337 & ~n11027 ) | ( n7337 & n14628 ) | ( ~n11027 & n14628 ) ;
  assign n14626 = ~n7067 & n10510 ;
  assign n14627 = n6215 & n14626 ;
  assign n14630 = n14629 ^ n14627 ^ n8772 ;
  assign n14632 = n3031 & ~n5634 ;
  assign n14633 = n14632 ^ n3386 ^ 1'b0 ;
  assign n14631 = ~n1899 & n4848 ;
  assign n14634 = n14633 ^ n14631 ^ 1'b0 ;
  assign n14635 = ~n7618 & n10939 ;
  assign n14636 = n7774 & n14635 ;
  assign n14637 = ( ~n632 & n14634 ) | ( ~n632 & n14636 ) | ( n14634 & n14636 ) ;
  assign n14638 = ~n2736 & n4574 ;
  assign n14639 = n14638 ^ n8432 ^ 1'b0 ;
  assign n14641 = n10481 ^ n5674 ^ n263 ;
  assign n14640 = ( ~n4386 & n5401 ) | ( ~n4386 & n10224 ) | ( n5401 & n10224 ) ;
  assign n14642 = n14641 ^ n14640 ^ 1'b0 ;
  assign n14643 = n5969 & n14642 ;
  assign n14644 = ( n10762 & n14639 ) | ( n10762 & n14643 ) | ( n14639 & n14643 ) ;
  assign n14645 = n2662 & ~n14644 ;
  assign n14646 = ( n717 & n2010 ) | ( n717 & ~n9957 ) | ( n2010 & ~n9957 ) ;
  assign n14647 = n5477 & n10564 ;
  assign n14649 = n1270 ^ n260 ^ 1'b0 ;
  assign n14648 = n3122 | n4041 ;
  assign n14650 = n14649 ^ n14648 ^ 1'b0 ;
  assign n14651 = n1114 ^ n522 ^ 1'b0 ;
  assign n14652 = n14650 & ~n14651 ;
  assign n14653 = n1220 | n14652 ;
  assign n14654 = n4989 ^ n1401 ^ 1'b0 ;
  assign n14655 = ~n6535 & n10309 ;
  assign n14656 = n5147 & n14655 ;
  assign n14657 = ( n972 & n13026 ) | ( n972 & ~n14656 ) | ( n13026 & ~n14656 ) ;
  assign n14658 = n14657 ^ n14569 ^ n12201 ;
  assign n14659 = ~n7212 & n14658 ;
  assign n14660 = ~n14654 & n14659 ;
  assign n14661 = n9258 ^ n8010 ^ 1'b0 ;
  assign n14662 = n8504 ^ n4761 ^ 1'b0 ;
  assign n14663 = n1150 & ~n14662 ;
  assign n14664 = ( n4796 & ~n10664 ) | ( n4796 & n14663 ) | ( ~n10664 & n14663 ) ;
  assign n14665 = ( ~n6847 & n7911 ) | ( ~n6847 & n8326 ) | ( n7911 & n8326 ) ;
  assign n14666 = n14665 ^ n2668 ^ 1'b0 ;
  assign n14667 = n5726 ^ n424 ^ 1'b0 ;
  assign n14668 = n14667 ^ n1684 ^ n595 ;
  assign n14669 = n2269 & ~n11877 ;
  assign n14670 = ~n14668 & n14669 ;
  assign n14674 = n4018 & n6165 ;
  assign n14671 = n867 ^ n316 ^ 1'b0 ;
  assign n14672 = n5687 & n14671 ;
  assign n14673 = n14672 ^ n1447 ^ 1'b0 ;
  assign n14675 = n14674 ^ n14673 ^ n7517 ;
  assign n14676 = n6954 ^ n3896 ^ 1'b0 ;
  assign n14677 = n253 & n14676 ;
  assign n14678 = n11606 ^ n5642 ^ 1'b0 ;
  assign n14679 = n4914 & ~n14678 ;
  assign n14680 = ( n4215 & ~n7423 ) | ( n4215 & n8262 ) | ( ~n7423 & n8262 ) ;
  assign n14681 = n14679 | n14680 ;
  assign n14686 = n4511 & n5088 ;
  assign n14687 = n14686 ^ n14554 ^ n9623 ;
  assign n14683 = n7517 ^ n1474 ^ n149 ;
  assign n14684 = ( n11184 & ~n13868 ) | ( n11184 & n14683 ) | ( ~n13868 & n14683 ) ;
  assign n14685 = n14684 ^ n13416 ^ n3843 ;
  assign n14682 = n7446 ^ n3436 ^ 1'b0 ;
  assign n14688 = n14687 ^ n14685 ^ n14682 ;
  assign n14689 = ~n2153 & n6352 ;
  assign n14690 = n6155 & n14689 ;
  assign n14691 = n14690 ^ n11520 ^ n9251 ;
  assign n14693 = ( n3189 & ~n3659 ) | ( n3189 & n8541 ) | ( ~n3659 & n8541 ) ;
  assign n14692 = ( n1558 & ~n3149 ) | ( n1558 & n10666 ) | ( ~n3149 & n10666 ) ;
  assign n14694 = n14693 ^ n14692 ^ n13725 ;
  assign n14695 = n6434 ^ n1102 ^ 1'b0 ;
  assign n14696 = n6677 ^ n2705 ^ n597 ;
  assign n14697 = n5791 ^ n1700 ^ 1'b0 ;
  assign n14698 = n14697 ^ n10896 ^ n10119 ;
  assign n14699 = n14698 ^ n2458 ^ 1'b0 ;
  assign n14700 = n5288 & n14699 ;
  assign n14701 = n14700 ^ n5458 ^ 1'b0 ;
  assign n14702 = ( n1284 & n14696 ) | ( n1284 & n14701 ) | ( n14696 & n14701 ) ;
  assign n14703 = n7236 ^ n3047 ^ n1021 ;
  assign n14704 = ( n5193 & n13571 ) | ( n5193 & ~n14703 ) | ( n13571 & ~n14703 ) ;
  assign n14707 = n11064 ^ n7673 ^ n214 ;
  assign n14705 = n5868 & n6295 ;
  assign n14706 = ( ~n965 & n6735 ) | ( ~n965 & n14705 ) | ( n6735 & n14705 ) ;
  assign n14708 = n14707 ^ n14706 ^ n13384 ;
  assign n14709 = n9609 ^ n2455 ^ 1'b0 ;
  assign n14715 = n8324 | n8886 ;
  assign n14711 = ( n2761 & n5210 ) | ( n2761 & n10301 ) | ( n5210 & n10301 ) ;
  assign n14712 = ( n884 & ~n2991 ) | ( n884 & n8584 ) | ( ~n2991 & n8584 ) ;
  assign n14713 = ( ~n1538 & n5391 ) | ( ~n1538 & n14712 ) | ( n5391 & n14712 ) ;
  assign n14714 = ( n1183 & n14711 ) | ( n1183 & n14713 ) | ( n14711 & n14713 ) ;
  assign n14716 = n14715 ^ n14714 ^ n8759 ;
  assign n14710 = n9826 & ~n13093 ;
  assign n14717 = n14716 ^ n14710 ^ 1'b0 ;
  assign n14718 = n6607 & n7676 ;
  assign n14719 = ~n11648 & n14718 ;
  assign n14720 = n1314 & ~n3964 ;
  assign n14721 = ( n1817 & n9842 ) | ( n1817 & n14720 ) | ( n9842 & n14720 ) ;
  assign n14725 = ( ~n842 & n1216 ) | ( ~n842 & n2842 ) | ( n1216 & n2842 ) ;
  assign n14723 = ( n1199 & n1700 ) | ( n1199 & ~n8585 ) | ( n1700 & ~n8585 ) ;
  assign n14722 = ( n1386 & n3302 ) | ( n1386 & n7482 ) | ( n3302 & n7482 ) ;
  assign n14724 = n14723 ^ n14722 ^ n12441 ;
  assign n14726 = n14725 ^ n14724 ^ 1'b0 ;
  assign n14727 = n4187 | n11703 ;
  assign n14728 = n7082 | n14727 ;
  assign n14729 = ( n5123 & ~n7101 ) | ( n5123 & n14087 ) | ( ~n7101 & n14087 ) ;
  assign n14730 = ( ~n12636 & n13192 ) | ( ~n12636 & n14729 ) | ( n13192 & n14729 ) ;
  assign n14731 = n11086 ^ n5776 ^ n3579 ;
  assign n14732 = ( ~n316 & n10115 ) | ( ~n316 & n14276 ) | ( n10115 & n14276 ) ;
  assign n14748 = x15 & ~n4841 ;
  assign n14749 = n14748 ^ x7 ^ 1'b0 ;
  assign n14750 = n14749 ^ n5527 ^ 1'b0 ;
  assign n14751 = n4575 ^ n1635 ^ 1'b0 ;
  assign n14752 = n2728 | n14751 ;
  assign n14753 = ( n1968 & n4308 ) | ( n1968 & ~n14752 ) | ( n4308 & ~n14752 ) ;
  assign n14754 = ( n9357 & ~n14750 ) | ( n9357 & n14753 ) | ( ~n14750 & n14753 ) ;
  assign n14736 = n4679 ^ n3164 ^ 1'b0 ;
  assign n14737 = n11660 ^ n6165 ^ n880 ;
  assign n14738 = n4418 & n14737 ;
  assign n14739 = n14738 ^ n3671 ^ 1'b0 ;
  assign n14740 = n218 | n14739 ;
  assign n14741 = n2549 | n14740 ;
  assign n14742 = ~n3478 & n7811 ;
  assign n14743 = n2921 & n14742 ;
  assign n14744 = ( ~n1597 & n14741 ) | ( ~n1597 & n14743 ) | ( n14741 & n14743 ) ;
  assign n14745 = n14744 ^ n3365 ^ 1'b0 ;
  assign n14746 = n14736 | n14745 ;
  assign n14733 = ( n4059 & n5523 ) | ( n4059 & n6219 ) | ( n5523 & n6219 ) ;
  assign n14734 = n4445 & n4468 ;
  assign n14735 = n14733 & n14734 ;
  assign n14747 = n14746 ^ n14735 ^ n5197 ;
  assign n14755 = n14754 ^ n14747 ^ n4566 ;
  assign n14756 = n2211 & n6689 ;
  assign n14757 = x105 | n1160 ;
  assign n14758 = n11922 & n14757 ;
  assign n14759 = ~n6519 & n10232 ;
  assign n14760 = n14759 ^ n1434 ^ 1'b0 ;
  assign n14761 = n14758 & n14760 ;
  assign n14763 = ~n953 & n3875 ;
  assign n14764 = n14763 ^ n3836 ^ 1'b0 ;
  assign n14762 = n4501 ^ n770 ^ 1'b0 ;
  assign n14765 = n14764 ^ n14762 ^ n11603 ;
  assign n14766 = ( n1841 & ~n2406 ) | ( n1841 & n4295 ) | ( ~n2406 & n4295 ) ;
  assign n14767 = ( n3607 & n8490 ) | ( n3607 & ~n14766 ) | ( n8490 & ~n14766 ) ;
  assign n14769 = ( n5266 & n6075 ) | ( n5266 & ~n8440 ) | ( n6075 & ~n8440 ) ;
  assign n14770 = n14769 ^ n2981 ^ n381 ;
  assign n14768 = ~n4770 & n6638 ;
  assign n14771 = n14770 ^ n14768 ^ 1'b0 ;
  assign n14772 = ( n12469 & ~n14767 ) | ( n12469 & n14771 ) | ( ~n14767 & n14771 ) ;
  assign n14773 = n1850 & n12769 ;
  assign n14774 = n14773 ^ n13563 ^ 1'b0 ;
  assign n14775 = ~n7578 & n12659 ;
  assign n14776 = ~n7953 & n14775 ;
  assign n14777 = n5507 & n14649 ;
  assign n14778 = n14777 ^ n14148 ^ n1160 ;
  assign n14779 = n14778 ^ n9387 ^ 1'b0 ;
  assign n14780 = n14779 ^ n14656 ^ n1610 ;
  assign n14781 = ( n1896 & n5266 ) | ( n1896 & n10162 ) | ( n5266 & n10162 ) ;
  assign n14782 = n14781 ^ n3019 ^ 1'b0 ;
  assign n14783 = n519 & n12776 ;
  assign n14784 = ( n4201 & n12652 ) | ( n4201 & ~n14783 ) | ( n12652 & ~n14783 ) ;
  assign n14785 = n10489 ^ n8551 ^ x14 ;
  assign n14786 = ( n3841 & n12816 ) | ( n3841 & ~n14785 ) | ( n12816 & ~n14785 ) ;
  assign n14788 = n5071 ^ n2065 ^ 1'b0 ;
  assign n14789 = n3232 | n14788 ;
  assign n14787 = n246 & ~n7365 ;
  assign n14790 = n14789 ^ n14787 ^ 1'b0 ;
  assign n14791 = n14790 ^ n10438 ^ n6794 ;
  assign n14792 = n7961 ^ n1375 ^ 1'b0 ;
  assign n14793 = x81 | n7180 ;
  assign n14794 = ( ~n138 & n6101 ) | ( ~n138 & n14793 ) | ( n6101 & n14793 ) ;
  assign n14795 = n11793 & ~n14794 ;
  assign n14796 = ~n14792 & n14795 ;
  assign n14797 = n2500 & n7765 ;
  assign n14798 = n5725 ^ n3084 ^ 1'b0 ;
  assign n14799 = ~n404 & n14798 ;
  assign n14800 = ~n14797 & n14799 ;
  assign n14801 = ~n5379 & n14800 ;
  assign n14802 = n6730 | n14801 ;
  assign n14803 = n8507 | n14802 ;
  assign n14804 = ( n1761 & n10713 ) | ( n1761 & n14803 ) | ( n10713 & n14803 ) ;
  assign n14805 = n2181 & n2183 ;
  assign n14806 = n2785 & n3147 ;
  assign n14807 = ( n11264 & n14805 ) | ( n11264 & ~n14806 ) | ( n14805 & ~n14806 ) ;
  assign n14808 = n12549 ^ n5966 ^ n773 ;
  assign n14809 = ( ~n6102 & n14807 ) | ( ~n6102 & n14808 ) | ( n14807 & n14808 ) ;
  assign n14810 = n1732 & ~n14809 ;
  assign n14811 = n3871 & ~n10673 ;
  assign n14812 = n8180 | n14811 ;
  assign n14813 = n14812 ^ n8195 ^ n2900 ;
  assign n14814 = n9612 ^ n3926 ^ 1'b0 ;
  assign n14815 = n9656 ^ n4713 ^ 1'b0 ;
  assign n14819 = ~n1651 & n7679 ;
  assign n14820 = n6443 | n14819 ;
  assign n14821 = n14820 ^ n7102 ^ 1'b0 ;
  assign n14816 = n895 & ~n4135 ;
  assign n14817 = ~n206 & n14816 ;
  assign n14818 = n14817 ^ n1887 ^ 1'b0 ;
  assign n14822 = n14821 ^ n14818 ^ n7678 ;
  assign n14823 = n3981 & n14822 ;
  assign n14824 = n14823 ^ n11936 ^ 1'b0 ;
  assign n14825 = n4325 & n14824 ;
  assign n14826 = ( ~n645 & n2249 ) | ( ~n645 & n7348 ) | ( n2249 & n7348 ) ;
  assign n14827 = n14826 ^ n8793 ^ n4542 ;
  assign n14828 = ( n1312 & n4930 ) | ( n1312 & n14827 ) | ( n4930 & n14827 ) ;
  assign n14829 = ~n4107 & n14055 ;
  assign n14830 = ~n5452 & n14829 ;
  assign n14831 = ~n6887 & n14830 ;
  assign n14832 = n14831 ^ n4468 ^ 1'b0 ;
  assign n14833 = n14832 ^ n267 ^ 1'b0 ;
  assign n14834 = n3470 & n14833 ;
  assign n14835 = n14834 ^ n12924 ^ 1'b0 ;
  assign n14836 = ~n3221 & n14835 ;
  assign n14837 = n5024 ^ n285 ^ 1'b0 ;
  assign n14840 = n11660 ^ n10678 ^ n2904 ;
  assign n14838 = n8632 ^ n5384 ^ n5325 ;
  assign n14839 = n14838 ^ n5245 ^ n1688 ;
  assign n14841 = n14840 ^ n14839 ^ n2137 ;
  assign n14842 = n14837 | n14841 ;
  assign n14843 = x107 | n14842 ;
  assign n14844 = n10565 ^ n7920 ^ n2550 ;
  assign n14845 = ( n147 & n1829 ) | ( n147 & n7223 ) | ( n1829 & n7223 ) ;
  assign n14846 = n14845 ^ n5961 ^ 1'b0 ;
  assign n14847 = ( n489 & n9349 ) | ( n489 & n14846 ) | ( n9349 & n14846 ) ;
  assign n14848 = ( ~x125 & n14844 ) | ( ~x125 & n14847 ) | ( n14844 & n14847 ) ;
  assign n14849 = ( n5497 & n13552 ) | ( n5497 & ~n13954 ) | ( n13552 & ~n13954 ) ;
  assign n14850 = n14290 ^ n12549 ^ n4325 ;
  assign n14851 = n14850 ^ n11860 ^ n2154 ;
  assign n14852 = n5833 ^ n3077 ^ n1199 ;
  assign n14853 = n14852 ^ n13294 ^ n7472 ;
  assign n14854 = ~n2623 & n9843 ;
  assign n14855 = n14854 ^ n8958 ^ 1'b0 ;
  assign n14856 = n10272 & ~n12882 ;
  assign n14857 = n652 & n14856 ;
  assign n14858 = ( n1567 & n1997 ) | ( n1567 & ~n3184 ) | ( n1997 & ~n3184 ) ;
  assign n14859 = n14858 ^ n6462 ^ 1'b0 ;
  assign n14860 = n14859 ^ n4477 ^ n2917 ;
  assign n14861 = ( n3335 & n4819 ) | ( n3335 & ~n14860 ) | ( n4819 & ~n14860 ) ;
  assign n14862 = ~n219 & n14861 ;
  assign n14863 = n8593 & n14862 ;
  assign n14864 = n10386 ^ n4304 ^ 1'b0 ;
  assign n14865 = n7596 & ~n14864 ;
  assign n14866 = n7340 ^ n1769 ^ 1'b0 ;
  assign n14867 = n847 | n14866 ;
  assign n14868 = n14867 ^ n9866 ^ n1796 ;
  assign n14869 = n9364 ^ n1217 ^ 1'b0 ;
  assign n14870 = n9360 ^ n8942 ^ 1'b0 ;
  assign n14871 = ( n3007 & n14869 ) | ( n3007 & n14870 ) | ( n14869 & n14870 ) ;
  assign n14872 = ( ~n14865 & n14868 ) | ( ~n14865 & n14871 ) | ( n14868 & n14871 ) ;
  assign n14873 = n12293 | n12740 ;
  assign n14874 = ( ~n8930 & n10234 ) | ( ~n8930 & n14873 ) | ( n10234 & n14873 ) ;
  assign n14875 = ~n11344 & n14874 ;
  assign n14882 = n6472 ^ n2189 ^ 1'b0 ;
  assign n14883 = ~n3022 & n14882 ;
  assign n14884 = n14883 ^ n5525 ^ 1'b0 ;
  assign n14885 = n7858 & n14884 ;
  assign n14881 = n3597 | n14199 ;
  assign n14886 = n14885 ^ n14881 ^ 1'b0 ;
  assign n14876 = n5677 & n6970 ;
  assign n14877 = n14876 ^ n1504 ^ 1'b0 ;
  assign n14878 = n8573 ^ n3047 ^ 1'b0 ;
  assign n14879 = n14877 & ~n14878 ;
  assign n14880 = n10058 & n14879 ;
  assign n14887 = n14886 ^ n14880 ^ 1'b0 ;
  assign n14888 = ~n1780 & n5760 ;
  assign n14889 = ~n4180 & n14888 ;
  assign n14891 = n7282 | n7705 ;
  assign n14892 = n14891 ^ n9257 ^ 1'b0 ;
  assign n14893 = n14892 ^ n7446 ^ n134 ;
  assign n14890 = n6896 ^ n6029 ^ n5277 ;
  assign n14894 = n14893 ^ n14890 ^ 1'b0 ;
  assign n14895 = ~n14889 & n14894 ;
  assign n14896 = ( n11582 & ~n14146 ) | ( n11582 & n14895 ) | ( ~n14146 & n14895 ) ;
  assign n14899 = n2270 | n3381 ;
  assign n14900 = n5451 & ~n14899 ;
  assign n14897 = n4949 ^ n1314 ^ n374 ;
  assign n14898 = ( ~n270 & n5482 ) | ( ~n270 & n14897 ) | ( n5482 & n14897 ) ;
  assign n14901 = n14900 ^ n14898 ^ n8493 ;
  assign n14902 = ( n7715 & n10676 ) | ( n7715 & n14901 ) | ( n10676 & n14901 ) ;
  assign n14903 = n822 | n9062 ;
  assign n14904 = ( ~n215 & n5081 ) | ( ~n215 & n7025 ) | ( n5081 & n7025 ) ;
  assign n14905 = n14904 ^ n4067 ^ 1'b0 ;
  assign n14906 = n14903 | n14905 ;
  assign n14907 = ~n6425 & n6749 ;
  assign n14908 = n14907 ^ n1370 ^ 1'b0 ;
  assign n14909 = n12845 ^ n3787 ^ 1'b0 ;
  assign n14910 = ( n3213 & n10015 ) | ( n3213 & ~n14909 ) | ( n10015 & ~n14909 ) ;
  assign n14911 = ( n2785 & ~n4334 ) | ( n2785 & n4578 ) | ( ~n4334 & n4578 ) ;
  assign n14912 = n14911 ^ n13900 ^ n10953 ;
  assign n14913 = ( n4840 & ~n5342 ) | ( n4840 & n8877 ) | ( ~n5342 & n8877 ) ;
  assign n14920 = ( ~n1049 & n3550 ) | ( ~n1049 & n4578 ) | ( n3550 & n4578 ) ;
  assign n14914 = n3438 ^ n1261 ^ 1'b0 ;
  assign n14915 = n143 & ~n14914 ;
  assign n14916 = ( ~n1070 & n2042 ) | ( ~n1070 & n3076 ) | ( n2042 & n3076 ) ;
  assign n14917 = n4710 & ~n14916 ;
  assign n14918 = ~n3588 & n14917 ;
  assign n14919 = ( n10087 & n14915 ) | ( n10087 & ~n14918 ) | ( n14915 & ~n14918 ) ;
  assign n14921 = n14920 ^ n14919 ^ 1'b0 ;
  assign n14922 = ( n2087 & n8719 ) | ( n2087 & ~n14921 ) | ( n8719 & ~n14921 ) ;
  assign n14923 = n7333 ^ n1192 ^ 1'b0 ;
  assign n14924 = n13275 & n14923 ;
  assign n14925 = ~n998 & n1965 ;
  assign n14926 = n14925 ^ n6973 ^ 1'b0 ;
  assign n14927 = ( n6590 & ~n8706 ) | ( n6590 & n14926 ) | ( ~n8706 & n14926 ) ;
  assign n14932 = n665 & ~n1592 ;
  assign n14933 = n2450 | n14932 ;
  assign n14934 = n14933 ^ n7765 ^ 1'b0 ;
  assign n14928 = ( n1645 & n3045 ) | ( n1645 & n3390 ) | ( n3045 & n3390 ) ;
  assign n14929 = n14928 ^ n8809 ^ n4742 ;
  assign n14930 = n14929 ^ n5006 ^ n1531 ;
  assign n14931 = n13050 & ~n14930 ;
  assign n14935 = n14934 ^ n14931 ^ 1'b0 ;
  assign n14936 = ( n1016 & n14927 ) | ( n1016 & ~n14935 ) | ( n14927 & ~n14935 ) ;
  assign n14939 = n427 | n625 ;
  assign n14937 = n8877 ^ n1468 ^ 1'b0 ;
  assign n14938 = n3210 & n14937 ;
  assign n14940 = n14939 ^ n14938 ^ 1'b0 ;
  assign n14943 = n854 & ~n1790 ;
  assign n14944 = n14943 ^ x44 ^ 1'b0 ;
  assign n14941 = n13046 ^ n11394 ^ n3836 ;
  assign n14942 = ( n1052 & n11793 ) | ( n1052 & ~n14941 ) | ( n11793 & ~n14941 ) ;
  assign n14945 = n14944 ^ n14942 ^ 1'b0 ;
  assign n14946 = ( n147 & n3665 ) | ( n147 & ~n11885 ) | ( n3665 & ~n11885 ) ;
  assign n14953 = n3234 ^ n2793 ^ n2004 ;
  assign n14950 = ( n1688 & n7478 ) | ( n1688 & ~n9173 ) | ( n7478 & ~n9173 ) ;
  assign n14948 = ( n1589 & ~n7747 ) | ( n1589 & n11263 ) | ( ~n7747 & n11263 ) ;
  assign n14949 = n5563 | n14948 ;
  assign n14951 = n14950 ^ n14949 ^ 1'b0 ;
  assign n14952 = ~n3016 & n14951 ;
  assign n14954 = n14953 ^ n14952 ^ 1'b0 ;
  assign n14947 = n7620 ^ n1750 ^ n748 ;
  assign n14955 = n14954 ^ n14947 ^ 1'b0 ;
  assign n14956 = ~n1788 & n14955 ;
  assign n14957 = n2541 | n14956 ;
  assign n14958 = n10065 ^ n3073 ^ 1'b0 ;
  assign n14959 = ~n11732 & n14958 ;
  assign n14960 = ( ~n4564 & n5329 ) | ( ~n4564 & n14959 ) | ( n5329 & n14959 ) ;
  assign n14961 = ~x32 & n14960 ;
  assign n14963 = n4260 | n10165 ;
  assign n14964 = n1382 & n2575 ;
  assign n14965 = n14964 ^ n2438 ^ 1'b0 ;
  assign n14966 = n14963 & ~n14965 ;
  assign n14962 = n4946 ^ n3540 ^ 1'b0 ;
  assign n14967 = n14966 ^ n14962 ^ n1594 ;
  assign n14968 = n885 & n11627 ;
  assign n14969 = n14968 ^ n397 ^ 1'b0 ;
  assign n14970 = n10625 ^ n884 ^ 1'b0 ;
  assign n14971 = n3922 & n14970 ;
  assign n14972 = ~n2475 & n3636 ;
  assign n14973 = ~n2155 & n14972 ;
  assign n14974 = n1935 | n14973 ;
  assign n14975 = n14971 | n14974 ;
  assign n14976 = ( n1294 & n4386 ) | ( n1294 & n5147 ) | ( n4386 & n5147 ) ;
  assign n14977 = n14976 ^ n5078 ^ 1'b0 ;
  assign n14978 = n1982 ^ n1763 ^ 1'b0 ;
  assign n14979 = ( ~n282 & n1318 ) | ( ~n282 & n4973 ) | ( n1318 & n4973 ) ;
  assign n14980 = n9294 & n14979 ;
  assign n14981 = ( n871 & n924 ) | ( n871 & n1388 ) | ( n924 & n1388 ) ;
  assign n14982 = ~n4704 & n14981 ;
  assign n14983 = n14221 ^ n3328 ^ 1'b0 ;
  assign n14984 = ~n5849 & n14983 ;
  assign n14985 = ( n7811 & n10910 ) | ( n7811 & ~n14984 ) | ( n10910 & ~n14984 ) ;
  assign n14986 = n14985 ^ n7694 ^ 1'b0 ;
  assign n14988 = ~n2603 & n11406 ;
  assign n14987 = n12020 ^ n1025 ^ 1'b0 ;
  assign n14989 = n14988 ^ n14987 ^ n10704 ;
  assign n14990 = n9796 ^ n9397 ^ n8224 ;
  assign n14991 = ~n1996 & n14990 ;
  assign n14992 = n6579 ^ n5754 ^ 1'b0 ;
  assign n14993 = n4697 & ~n14992 ;
  assign n14994 = n5906 ^ n2769 ^ 1'b0 ;
  assign n14995 = n14994 ^ n10202 ^ n4425 ;
  assign n14996 = n14995 ^ n13890 ^ 1'b0 ;
  assign n14997 = ( n1436 & n14993 ) | ( n1436 & n14996 ) | ( n14993 & n14996 ) ;
  assign n14998 = n6344 & n10925 ;
  assign n14999 = n2734 ^ n2720 ^ n2517 ;
  assign n15000 = ( n803 & n11636 ) | ( n803 & ~n14999 ) | ( n11636 & ~n14999 ) ;
  assign n15001 = n12365 ^ n10824 ^ n1335 ;
  assign n15002 = ( n4921 & ~n14979 ) | ( n4921 & n15001 ) | ( ~n14979 & n15001 ) ;
  assign n15003 = n13084 ^ n10599 ^ n2946 ;
  assign n15005 = n976 & ~n4842 ;
  assign n15006 = n5904 & n15005 ;
  assign n15004 = n5714 & n5761 ;
  assign n15007 = n15006 ^ n15004 ^ 1'b0 ;
  assign n15008 = ( n7254 & n10871 ) | ( n7254 & n14845 ) | ( n10871 & n14845 ) ;
  assign n15009 = ( n593 & ~n5405 ) | ( n593 & n15008 ) | ( ~n5405 & n15008 ) ;
  assign n15010 = ( n4820 & n11534 ) | ( n4820 & n13847 ) | ( n11534 & n13847 ) ;
  assign n15012 = n8967 ^ n7615 ^ 1'b0 ;
  assign n15013 = n3182 | n15012 ;
  assign n15011 = ~n677 & n11573 ;
  assign n15014 = n15013 ^ n15011 ^ 1'b0 ;
  assign n15015 = n3880 & n4496 ;
  assign n15016 = n3646 & n15015 ;
  assign n15017 = ( n6371 & n9698 ) | ( n6371 & ~n15016 ) | ( n9698 & ~n15016 ) ;
  assign n15018 = n15017 ^ n11159 ^ 1'b0 ;
  assign n15019 = ~n4990 & n15018 ;
  assign n15020 = n15019 ^ n1470 ^ 1'b0 ;
  assign n15021 = ( n5304 & ~n15014 ) | ( n5304 & n15020 ) | ( ~n15014 & n15020 ) ;
  assign n15022 = ( n2453 & n6537 ) | ( n2453 & ~n9205 ) | ( n6537 & ~n9205 ) ;
  assign n15023 = n1289 | n5705 ;
  assign n15024 = n15023 ^ n12178 ^ n4341 ;
  assign n15025 = n15024 ^ n2709 ^ n1143 ;
  assign n15026 = ( n195 & ~n15022 ) | ( n195 & n15025 ) | ( ~n15022 & n15025 ) ;
  assign n15027 = ( n5692 & ~n7560 ) | ( n5692 & n13073 ) | ( ~n7560 & n13073 ) ;
  assign n15030 = n3667 | n8648 ;
  assign n15029 = n3325 ^ n2827 ^ n2331 ;
  assign n15031 = n15030 ^ n15029 ^ n7502 ;
  assign n15028 = ( n5331 & ~n10459 ) | ( n5331 & n10948 ) | ( ~n10459 & n10948 ) ;
  assign n15032 = n15031 ^ n15028 ^ n14206 ;
  assign n15033 = ~n15027 & n15032 ;
  assign n15034 = n8239 ^ n5338 ^ 1'b0 ;
  assign n15035 = n15034 ^ n10376 ^ n2916 ;
  assign n15045 = n4301 ^ n3652 ^ 1'b0 ;
  assign n15036 = n7961 ^ n7352 ^ n2889 ;
  assign n15037 = ~n2141 & n15036 ;
  assign n15038 = n8082 & n15037 ;
  assign n15039 = n10524 ^ n4747 ^ n2544 ;
  assign n15040 = ( ~n4048 & n5699 ) | ( ~n4048 & n7283 ) | ( n5699 & n7283 ) ;
  assign n15041 = ( n5491 & ~n15039 ) | ( n5491 & n15040 ) | ( ~n15039 & n15040 ) ;
  assign n15042 = ( ~n8602 & n9597 ) | ( ~n8602 & n15041 ) | ( n9597 & n15041 ) ;
  assign n15043 = n15042 ^ n4149 ^ 1'b0 ;
  assign n15044 = n15038 | n15043 ;
  assign n15046 = n15045 ^ n15044 ^ 1'b0 ;
  assign n15047 = ( ~n1578 & n15035 ) | ( ~n1578 & n15046 ) | ( n15035 & n15046 ) ;
  assign n15048 = n14628 ^ n5288 ^ n422 ;
  assign n15049 = n8212 ^ n2143 ^ n894 ;
  assign n15050 = n15049 ^ n9160 ^ 1'b0 ;
  assign n15051 = n8330 & ~n15050 ;
  assign n15052 = n15051 ^ n11230 ^ n9711 ;
  assign n15053 = ( n2416 & n4862 ) | ( n2416 & ~n5703 ) | ( n4862 & ~n5703 ) ;
  assign n15054 = n15053 ^ n3825 ^ n2051 ;
  assign n15055 = n13704 | n15054 ;
  assign n15056 = n14641 ^ n12236 ^ 1'b0 ;
  assign n15057 = ~n15055 & n15056 ;
  assign n15058 = n14437 ^ n8977 ^ n431 ;
  assign n15059 = ( ~n1865 & n7929 ) | ( ~n1865 & n11556 ) | ( n7929 & n11556 ) ;
  assign n15060 = ~n1821 & n3314 ;
  assign n15061 = n15060 ^ n12960 ^ 1'b0 ;
  assign n15062 = n14017 ^ n6688 ^ 1'b0 ;
  assign n15063 = ~n15061 & n15062 ;
  assign n15072 = n9539 ^ n3981 ^ 1'b0 ;
  assign n15073 = n7421 | n15072 ;
  assign n15074 = n3802 & ~n15073 ;
  assign n15075 = n15074 ^ n6598 ^ n386 ;
  assign n15070 = n2414 & n3643 ;
  assign n15071 = n14065 & n15070 ;
  assign n15076 = n15075 ^ n15071 ^ n6377 ;
  assign n15065 = ~n3785 & n7121 ;
  assign n15066 = n15065 ^ n3578 ^ 1'b0 ;
  assign n15067 = ~n5201 & n15066 ;
  assign n15068 = n9980 & n15067 ;
  assign n15069 = n15068 ^ n3577 ^ 1'b0 ;
  assign n15077 = n15076 ^ n15069 ^ 1'b0 ;
  assign n15064 = n6887 | n10131 ;
  assign n15078 = n15077 ^ n15064 ^ n1978 ;
  assign n15079 = ( ~n2186 & n7342 ) | ( ~n2186 & n8003 ) | ( n7342 & n8003 ) ;
  assign n15080 = n357 | n1883 ;
  assign n15081 = ( n6142 & n10927 ) | ( n6142 & ~n15080 ) | ( n10927 & ~n15080 ) ;
  assign n15082 = ( ~n577 & n8918 ) | ( ~n577 & n15081 ) | ( n8918 & n15081 ) ;
  assign n15083 = ~n6652 & n15082 ;
  assign n15084 = n15083 ^ n14472 ^ 1'b0 ;
  assign n15085 = ( n598 & n624 ) | ( n598 & n2319 ) | ( n624 & n2319 ) ;
  assign n15086 = ( n3969 & n9953 ) | ( n3969 & n15085 ) | ( n9953 & n15085 ) ;
  assign n15087 = n3506 & ~n10270 ;
  assign n15088 = n4295 & n15087 ;
  assign n15089 = n15086 & ~n15088 ;
  assign n15090 = n834 | n13066 ;
  assign n15092 = n8132 ^ n8023 ^ n867 ;
  assign n15093 = n2663 ^ n1360 ^ 1'b0 ;
  assign n15094 = n15092 & ~n15093 ;
  assign n15095 = n11283 ^ n6692 ^ 1'b0 ;
  assign n15096 = n15094 & n15095 ;
  assign n15091 = n3899 & n4751 ;
  assign n15097 = n15096 ^ n15091 ^ n7555 ;
  assign n15098 = n12757 & n15097 ;
  assign n15099 = n15098 ^ n10703 ^ 1'b0 ;
  assign n15100 = n9506 ^ n1702 ^ 1'b0 ;
  assign n15101 = n2820 & n15100 ;
  assign n15103 = ( ~n2761 & n6649 ) | ( ~n2761 & n13648 ) | ( n6649 & n13648 ) ;
  assign n15104 = ( ~n12711 & n13685 ) | ( ~n12711 & n15103 ) | ( n13685 & n15103 ) ;
  assign n15102 = n3484 & n6315 ;
  assign n15105 = n15104 ^ n15102 ^ 1'b0 ;
  assign n15107 = ( ~n203 & n1669 ) | ( ~n203 & n9391 ) | ( n1669 & n9391 ) ;
  assign n15108 = n15107 ^ n7482 ^ n3862 ;
  assign n15106 = ( ~n2611 & n6160 ) | ( ~n2611 & n9503 ) | ( n6160 & n9503 ) ;
  assign n15109 = n15108 ^ n15106 ^ n6429 ;
  assign n15110 = n3774 | n8448 ;
  assign n15111 = n14090 | n15110 ;
  assign n15112 = n15111 ^ n9822 ^ 1'b0 ;
  assign n15113 = ( n2247 & ~n3678 ) | ( n2247 & n14233 ) | ( ~n3678 & n14233 ) ;
  assign n15114 = n15113 ^ n9096 ^ n5913 ;
  assign n15115 = n8652 ^ n2905 ^ 1'b0 ;
  assign n15116 = n13008 & ~n15115 ;
  assign n15117 = ~n452 & n15116 ;
  assign n15118 = ~n7688 & n15117 ;
  assign n15119 = n3344 & n15118 ;
  assign n15120 = ( n1736 & n3186 ) | ( n1736 & ~n5250 ) | ( n3186 & ~n5250 ) ;
  assign n15121 = n15120 ^ n3229 ^ 1'b0 ;
  assign n15123 = n6128 ^ n1740 ^ 1'b0 ;
  assign n15122 = n11653 ^ n9352 ^ n213 ;
  assign n15124 = n15123 ^ n15122 ^ n3051 ;
  assign n15132 = n12273 ^ n9105 ^ 1'b0 ;
  assign n15133 = n3359 & ~n15132 ;
  assign n15130 = n12217 ^ n4541 ^ n2301 ;
  assign n15131 = ( n6443 & n14557 ) | ( n6443 & n15130 ) | ( n14557 & n15130 ) ;
  assign n15134 = n15133 ^ n15131 ^ n7806 ;
  assign n15125 = n714 & n6820 ;
  assign n15126 = n15125 ^ n1329 ^ 1'b0 ;
  assign n15127 = n6659 ^ n2798 ^ n1697 ;
  assign n15128 = n15127 ^ n2835 ^ 1'b0 ;
  assign n15129 = n15126 & n15128 ;
  assign n15135 = n15134 ^ n15129 ^ n646 ;
  assign n15136 = n374 & ~n12528 ;
  assign n15137 = n10743 & n15136 ;
  assign n15138 = ( n2157 & ~n9285 ) | ( n2157 & n15137 ) | ( ~n9285 & n15137 ) ;
  assign n15139 = ( ~n1510 & n9313 ) | ( ~n1510 & n10070 ) | ( n9313 & n10070 ) ;
  assign n15140 = n15139 ^ n9292 ^ 1'b0 ;
  assign n15141 = n15140 ^ n7041 ^ n6029 ;
  assign n15142 = n15141 ^ n10533 ^ 1'b0 ;
  assign n15143 = n13893 & ~n15142 ;
  assign n15144 = ( n360 & n5912 ) | ( n360 & n15143 ) | ( n5912 & n15143 ) ;
  assign n15148 = n4189 & n11596 ;
  assign n15149 = n966 & n15148 ;
  assign n15150 = ( ~n9081 & n12186 ) | ( ~n9081 & n15149 ) | ( n12186 & n15149 ) ;
  assign n15145 = n6714 | n8242 ;
  assign n15146 = n15145 ^ n4505 ^ 1'b0 ;
  assign n15147 = n15146 ^ n5582 ^ n1239 ;
  assign n15151 = n15150 ^ n15147 ^ n4164 ;
  assign n15152 = n1001 & ~n1154 ;
  assign n15153 = n11234 ^ n2917 ^ 1'b0 ;
  assign n15154 = n5948 ^ n2954 ^ 1'b0 ;
  assign n15155 = ~n15153 & n15154 ;
  assign n15156 = n4338 | n7718 ;
  assign n15157 = ( ~n1153 & n2049 ) | ( ~n1153 & n15156 ) | ( n2049 & n15156 ) ;
  assign n15160 = n1335 & ~n4707 ;
  assign n15161 = n14766 & n15160 ;
  assign n15158 = n3083 | n6289 ;
  assign n15159 = n12419 & ~n15158 ;
  assign n15162 = n15161 ^ n15159 ^ n8286 ;
  assign n15163 = ( x68 & n15157 ) | ( x68 & n15162 ) | ( n15157 & n15162 ) ;
  assign n15164 = n3461 | n15163 ;
  assign n15166 = n442 & ~n3639 ;
  assign n15165 = n14146 ^ n2646 ^ n1172 ;
  assign n15167 = n15166 ^ n15165 ^ n3743 ;
  assign n15173 = n4576 ^ n4092 ^ 1'b0 ;
  assign n15174 = n3468 & n15173 ;
  assign n15169 = ~n1123 & n1244 ;
  assign n15170 = n1426 & n15169 ;
  assign n15168 = n4093 ^ n3131 ^ 1'b0 ;
  assign n15171 = n15170 ^ n15168 ^ n5453 ;
  assign n15172 = n563 & ~n15171 ;
  assign n15175 = n15174 ^ n15172 ^ 1'b0 ;
  assign n15176 = n413 & n9086 ;
  assign n15177 = ( n7580 & ~n7620 ) | ( n7580 & n11976 ) | ( ~n7620 & n11976 ) ;
  assign n15178 = n12259 ^ n3918 ^ 1'b0 ;
  assign n15179 = n6598 & ~n15178 ;
  assign n15183 = ( n145 & n3127 ) | ( n145 & ~n5135 ) | ( n3127 & ~n5135 ) ;
  assign n15180 = n5828 & ~n13517 ;
  assign n15181 = n15180 ^ n11135 ^ 1'b0 ;
  assign n15182 = n7692 & ~n15181 ;
  assign n15184 = n15183 ^ n15182 ^ 1'b0 ;
  assign n15185 = n2954 | n7013 ;
  assign n15186 = n11104 ^ n4249 ^ 1'b0 ;
  assign n15187 = n10694 | n15186 ;
  assign n15188 = n15185 | n15187 ;
  assign n15189 = n15188 ^ n5816 ^ n4098 ;
  assign n15190 = n3163 | n5156 ;
  assign n15191 = x106 | n15190 ;
  assign n15195 = n11239 ^ n8486 ^ n1151 ;
  assign n15196 = ( n10767 & n15071 ) | ( n10767 & n15195 ) | ( n15071 & n15195 ) ;
  assign n15193 = ( x2 & ~n3035 ) | ( x2 & n4725 ) | ( ~n3035 & n4725 ) ;
  assign n15192 = n729 & ~n11248 ;
  assign n15194 = n15193 ^ n15192 ^ 1'b0 ;
  assign n15197 = n15196 ^ n15194 ^ 1'b0 ;
  assign n15198 = ~n10974 & n15197 ;
  assign n15199 = n15198 ^ n5793 ^ 1'b0 ;
  assign n15200 = n15191 & ~n15199 ;
  assign n15201 = n3869 ^ n1012 ^ 1'b0 ;
  assign n15202 = n15201 ^ n1523 ^ n986 ;
  assign n15203 = n4155 & n10457 ;
  assign n15204 = ~n8914 & n12033 ;
  assign n15205 = n15204 ^ n6162 ^ 1'b0 ;
  assign n15206 = n6939 & ~n15205 ;
  assign n15207 = n9062 & n15206 ;
  assign n15208 = ( n10442 & n15203 ) | ( n10442 & ~n15207 ) | ( n15203 & ~n15207 ) ;
  assign n15209 = n10913 ^ n4030 ^ 1'b0 ;
  assign n15210 = n4793 | n15209 ;
  assign n15211 = n15210 ^ n3966 ^ n1836 ;
  assign n15212 = n6857 ^ n4944 ^ 1'b0 ;
  assign n15213 = n10449 & ~n15212 ;
  assign n15214 = n9583 ^ n4152 ^ 1'b0 ;
  assign n15215 = ~n2955 & n6404 ;
  assign n15216 = n15215 ^ n5353 ^ 1'b0 ;
  assign n15217 = n9408 ^ n8421 ^ n1378 ;
  assign n15218 = ( n2278 & n5740 ) | ( n2278 & n7893 ) | ( n5740 & n7893 ) ;
  assign n15219 = n6605 & n15218 ;
  assign n15220 = ( n705 & ~n15217 ) | ( n705 & n15219 ) | ( ~n15217 & n15219 ) ;
  assign n15221 = n15216 & n15220 ;
  assign n15222 = n15214 & n15221 ;
  assign n15223 = n12459 ^ n10939 ^ n4273 ;
  assign n15224 = ~n5921 & n15223 ;
  assign n15225 = ( x13 & n310 ) | ( x13 & ~n2661 ) | ( n310 & ~n2661 ) ;
  assign n15226 = n15225 ^ n11137 ^ 1'b0 ;
  assign n15227 = ~n11091 & n15226 ;
  assign n15228 = n12238 ^ n2494 ^ n1905 ;
  assign n15229 = n15228 ^ n527 ^ 1'b0 ;
  assign n15230 = n7377 & n7381 ;
  assign n15231 = n15230 ^ n3825 ^ 1'b0 ;
  assign n15232 = n427 & n13978 ;
  assign n15233 = n5310 & n8860 ;
  assign n15234 = n15233 ^ n12576 ^ 1'b0 ;
  assign n15235 = ~n15232 & n15234 ;
  assign n15240 = n11263 ^ n6805 ^ n720 ;
  assign n15236 = ( n2023 & n4736 ) | ( n2023 & ~n13678 ) | ( n4736 & ~n13678 ) ;
  assign n15237 = ( n685 & ~n7758 ) | ( n685 & n15236 ) | ( ~n7758 & n15236 ) ;
  assign n15238 = n15237 ^ n1452 ^ 1'b0 ;
  assign n15239 = n5198 | n15238 ;
  assign n15241 = n15240 ^ n15239 ^ 1'b0 ;
  assign n15242 = ( n3008 & ~n3023 ) | ( n3008 & n15241 ) | ( ~n3023 & n15241 ) ;
  assign n15247 = n4530 | n6358 ;
  assign n15243 = n14503 ^ n2234 ^ 1'b0 ;
  assign n15244 = n10610 & ~n15243 ;
  assign n15245 = n15244 ^ n519 ^ 1'b0 ;
  assign n15246 = n1497 & n15245 ;
  assign n15248 = n15247 ^ n15246 ^ 1'b0 ;
  assign n15249 = ( n2661 & ~n7125 ) | ( n2661 & n15248 ) | ( ~n7125 & n15248 ) ;
  assign n15250 = n15249 ^ n8916 ^ 1'b0 ;
  assign n15251 = ~n468 & n504 ;
  assign n15252 = n2227 & ~n15251 ;
  assign n15255 = n4538 ^ n1366 ^ 1'b0 ;
  assign n15256 = ~n2199 & n15255 ;
  assign n15257 = n15256 ^ n7805 ^ n1593 ;
  assign n15258 = ~n7562 & n15257 ;
  assign n15259 = n15258 ^ n5415 ^ 1'b0 ;
  assign n15253 = n11897 ^ n7720 ^ 1'b0 ;
  assign n15254 = n4190 & ~n15253 ;
  assign n15260 = n15259 ^ n15254 ^ n6768 ;
  assign n15261 = n7591 ^ n5672 ^ 1'b0 ;
  assign n15262 = n15260 | n15261 ;
  assign n15263 = n12996 | n15202 ;
  assign n15264 = n15263 ^ n9385 ^ 1'b0 ;
  assign n15265 = n14457 ^ n5519 ^ 1'b0 ;
  assign n15266 = ( n2426 & n3015 ) | ( n2426 & n3255 ) | ( n3015 & n3255 ) ;
  assign n15267 = n15266 ^ n2070 ^ 1'b0 ;
  assign n15268 = n3302 & n14271 ;
  assign n15269 = n15268 ^ n14687 ^ 1'b0 ;
  assign n15270 = ( n5152 & n5822 ) | ( n5152 & n8943 ) | ( n5822 & n8943 ) ;
  assign n15271 = n3924 | n9427 ;
  assign n15272 = n10755 ^ n4253 ^ n1405 ;
  assign n15273 = ( n1443 & n1662 ) | ( n1443 & n9186 ) | ( n1662 & n9186 ) ;
  assign n15274 = n15273 ^ n14510 ^ 1'b0 ;
  assign n15275 = n15272 | n15274 ;
  assign n15279 = n8134 ^ n4218 ^ 1'b0 ;
  assign n15276 = n5769 & n11003 ;
  assign n15277 = n6308 ^ x25 ^ 1'b0 ;
  assign n15278 = ~n15276 & n15277 ;
  assign n15280 = n15279 ^ n15278 ^ n14224 ;
  assign n15281 = n10947 ^ n3688 ^ n1645 ;
  assign n15282 = n15281 ^ n13720 ^ n8604 ;
  assign n15283 = n2381 & ~n5318 ;
  assign n15284 = n15283 ^ n1828 ^ 1'b0 ;
  assign n15285 = n12274 ^ n7989 ^ 1'b0 ;
  assign n15286 = n15284 & n15285 ;
  assign n15287 = ~n590 & n7359 ;
  assign n15288 = n14627 | n15287 ;
  assign n15289 = n3336 | n5977 ;
  assign n15290 = n15030 ^ n3215 ^ 1'b0 ;
  assign n15291 = n5780 & n15290 ;
  assign n15292 = ~n3830 & n13568 ;
  assign n15293 = n259 & n1875 ;
  assign n15294 = n15293 ^ n9094 ^ 1'b0 ;
  assign n15295 = ( n15291 & n15292 ) | ( n15291 & n15294 ) | ( n15292 & n15294 ) ;
  assign n15299 = n11596 ^ n5542 ^ n621 ;
  assign n15296 = n10759 ^ n1259 ^ 1'b0 ;
  assign n15297 = n1914 & n15296 ;
  assign n15298 = n15297 ^ n9558 ^ n6487 ;
  assign n15300 = n15299 ^ n15298 ^ n12794 ;
  assign n15301 = n15300 ^ n8943 ^ 1'b0 ;
  assign n15303 = n941 & n3456 ;
  assign n15304 = n15303 ^ n6750 ^ 1'b0 ;
  assign n15305 = n2720 & n15304 ;
  assign n15306 = ~n1865 & n15305 ;
  assign n15307 = ( n2631 & n6436 ) | ( n2631 & ~n15306 ) | ( n6436 & ~n15306 ) ;
  assign n15302 = n579 & ~n1883 ;
  assign n15308 = n15307 ^ n15302 ^ n6203 ;
  assign n15309 = n15308 ^ n14388 ^ n3716 ;
  assign n15310 = n15309 ^ n4393 ^ 1'b0 ;
  assign n15311 = n15310 ^ n9855 ^ n4268 ;
  assign n15312 = ( ~n9994 & n15301 ) | ( ~n9994 & n15311 ) | ( n15301 & n15311 ) ;
  assign n15313 = n3439 & ~n4745 ;
  assign n15314 = n15313 ^ n4663 ^ 1'b0 ;
  assign n15315 = ( n4436 & n5669 ) | ( n4436 & n14607 ) | ( n5669 & n14607 ) ;
  assign n15316 = n10058 & n15315 ;
  assign n15317 = n15316 ^ n8857 ^ n2991 ;
  assign n15318 = ( n315 & n9902 ) | ( n315 & ~n15317 ) | ( n9902 & ~n15317 ) ;
  assign n15319 = n8300 & ~n15318 ;
  assign n15320 = n15314 & n15319 ;
  assign n15321 = n11785 ^ n10862 ^ n183 ;
  assign n15322 = n1817 & n15321 ;
  assign n15323 = n8294 & ~n10618 ;
  assign n15324 = n15323 ^ n2488 ^ n1219 ;
  assign n15325 = n15324 ^ n5648 ^ 1'b0 ;
  assign n15326 = n1370 | n3620 ;
  assign n15327 = n15326 ^ n8510 ^ n5397 ;
  assign n15328 = ( n5311 & n12323 ) | ( n5311 & n14582 ) | ( n12323 & n14582 ) ;
  assign n15329 = n6013 ^ n2292 ^ n2014 ;
  assign n15330 = n15329 ^ n7236 ^ n4954 ;
  assign n15331 = n15330 ^ n5216 ^ 1'b0 ;
  assign n15332 = n3333 | n15331 ;
  assign n15333 = n10880 & n15332 ;
  assign n15334 = n5985 | n15333 ;
  assign n15335 = n15334 ^ n2113 ^ 1'b0 ;
  assign n15337 = n2073 ^ n1011 ^ 1'b0 ;
  assign n15338 = n7898 | n15337 ;
  assign n15336 = ~n1040 & n11034 ;
  assign n15339 = n15338 ^ n15336 ^ 1'b0 ;
  assign n15340 = ~n4103 & n15339 ;
  assign n15341 = n15340 ^ n1758 ^ 1'b0 ;
  assign n15342 = n2509 ^ n265 ^ 1'b0 ;
  assign n15343 = n2685 & n15342 ;
  assign n15344 = n15343 ^ n13611 ^ 1'b0 ;
  assign n15345 = n5959 | n15344 ;
  assign n15346 = n1794 & ~n15345 ;
  assign n15347 = n2983 & n15346 ;
  assign n15348 = n3016 & ~n15347 ;
  assign n15349 = n14134 & ~n15348 ;
  assign n15353 = ~n3469 & n13411 ;
  assign n15354 = n3067 & n15353 ;
  assign n15350 = ( n863 & ~n2707 ) | ( n863 & n12068 ) | ( ~n2707 & n12068 ) ;
  assign n15351 = n9975 & ~n15350 ;
  assign n15352 = ~n10449 & n15351 ;
  assign n15355 = n15354 ^ n15352 ^ n713 ;
  assign n15356 = ( n166 & ~n5248 ) | ( n166 & n11441 ) | ( ~n5248 & n11441 ) ;
  assign n15357 = n1470 & ~n3382 ;
  assign n15358 = n2495 & n15357 ;
  assign n15359 = n2886 & ~n15251 ;
  assign n15360 = n15359 ^ n2600 ^ 1'b0 ;
  assign n15361 = n15360 ^ n3234 ^ 1'b0 ;
  assign n15362 = n15358 & n15361 ;
  assign n15363 = n3758 ^ n1900 ^ n322 ;
  assign n15364 = n15363 ^ n11609 ^ n6316 ;
  assign n15367 = n756 & n3666 ;
  assign n15365 = ~n9640 & n14482 ;
  assign n15366 = n9237 & n15365 ;
  assign n15368 = n15367 ^ n15366 ^ n8802 ;
  assign n15369 = n1836 & n5491 ;
  assign n15370 = n15369 ^ n14226 ^ n2023 ;
  assign n15371 = n5415 & n15370 ;
  assign n15372 = n15371 ^ n8370 ^ 1'b0 ;
  assign n15373 = ( n5559 & n13723 ) | ( n5559 & ~n15372 ) | ( n13723 & ~n15372 ) ;
  assign n15376 = n4112 | n6378 ;
  assign n15377 = n15376 ^ n6874 ^ 1'b0 ;
  assign n15374 = n8167 ^ n6145 ^ n3372 ;
  assign n15375 = n1149 & n15374 ;
  assign n15378 = n15377 ^ n15375 ^ n9435 ;
  assign n15379 = n15378 ^ n5598 ^ n2569 ;
  assign n15386 = ( x36 & n4501 ) | ( x36 & n12626 ) | ( n4501 & n12626 ) ;
  assign n15380 = n4401 ^ n2759 ^ 1'b0 ;
  assign n15381 = ( n2257 & ~n5702 ) | ( n2257 & n15380 ) | ( ~n5702 & n15380 ) ;
  assign n15382 = n6705 & ~n15381 ;
  assign n15383 = ( n8710 & n10430 ) | ( n8710 & ~n15382 ) | ( n10430 & ~n15382 ) ;
  assign n15384 = n15383 ^ n13961 ^ n5438 ;
  assign n15385 = ~n10823 & n15384 ;
  assign n15387 = n15386 ^ n15385 ^ n1474 ;
  assign n15388 = n10428 ^ n7325 ^ 1'b0 ;
  assign n15389 = n9582 & ~n15388 ;
  assign n15390 = n15389 ^ n4033 ^ 1'b0 ;
  assign n15399 = n1100 & ~n3854 ;
  assign n15400 = n15399 ^ n4971 ^ 1'b0 ;
  assign n15391 = n2286 & n5772 ;
  assign n15392 = ( ~n7177 & n13649 ) | ( ~n7177 & n15391 ) | ( n13649 & n15391 ) ;
  assign n15393 = ( n4974 & ~n6913 ) | ( n4974 & n8094 ) | ( ~n6913 & n8094 ) ;
  assign n15394 = n1617 & ~n11391 ;
  assign n15395 = n15394 ^ n4059 ^ 1'b0 ;
  assign n15396 = n15393 & n15395 ;
  assign n15397 = ~n14010 & n15396 ;
  assign n15398 = n15392 | n15397 ;
  assign n15401 = n15400 ^ n15398 ^ 1'b0 ;
  assign n15402 = n3125 | n4080 ;
  assign n15403 = n5798 ^ n5523 ^ 1'b0 ;
  assign n15404 = n2900 & n15403 ;
  assign n15405 = ( n1531 & n4030 ) | ( n1531 & ~n15404 ) | ( n4030 & ~n15404 ) ;
  assign n15406 = n8926 ^ n8505 ^ 1'b0 ;
  assign n15407 = ( n1460 & n8337 ) | ( n1460 & n15406 ) | ( n8337 & n15406 ) ;
  assign n15410 = n9277 ^ n4825 ^ n410 ;
  assign n15411 = ( ~n451 & n4776 ) | ( ~n451 & n15410 ) | ( n4776 & n15410 ) ;
  assign n15408 = n5016 & n6855 ;
  assign n15409 = ( n1157 & ~n5129 ) | ( n1157 & n15408 ) | ( ~n5129 & n15408 ) ;
  assign n15412 = n15411 ^ n15409 ^ n10721 ;
  assign n15413 = n935 & ~n1290 ;
  assign n15414 = ~n3339 & n15413 ;
  assign n15415 = n15414 ^ n8367 ^ 1'b0 ;
  assign n15416 = n1862 & ~n14554 ;
  assign n15417 = n15034 & n15416 ;
  assign n15418 = n15417 ^ n950 ^ 1'b0 ;
  assign n15419 = n15415 | n15418 ;
  assign n15420 = ( n5525 & ~n13513 ) | ( n5525 & n15419 ) | ( ~n13513 & n15419 ) ;
  assign n15421 = ~n4501 & n14152 ;
  assign n15424 = n13423 ^ n11137 ^ n7378 ;
  assign n15422 = n4168 ^ n2549 ^ 1'b0 ;
  assign n15423 = n15422 ^ n7568 ^ n5187 ;
  assign n15425 = n15424 ^ n15423 ^ 1'b0 ;
  assign n15426 = n6741 | n15425 ;
  assign n15427 = n2623 | n8275 ;
  assign n15428 = n3646 ^ n3625 ^ 1'b0 ;
  assign n15429 = n2464 & n15428 ;
  assign n15430 = ~n4289 & n15429 ;
  assign n15431 = ( n4365 & n15107 ) | ( n4365 & ~n15430 ) | ( n15107 & ~n15430 ) ;
  assign n15432 = n15431 ^ n1055 ^ 1'b0 ;
  assign n15433 = ~n7548 & n15432 ;
  assign n15434 = ( n356 & n8921 ) | ( n356 & n15433 ) | ( n8921 & n15433 ) ;
  assign n15435 = n15434 ^ n4226 ^ 1'b0 ;
  assign n15436 = n2730 | n15435 ;
  assign n15442 = n7904 ^ n3838 ^ n314 ;
  assign n15443 = n1660 & n15442 ;
  assign n15444 = ~n6054 & n15443 ;
  assign n15440 = n259 & n5961 ;
  assign n15441 = n3493 & n15440 ;
  assign n15437 = n8423 ^ n2643 ^ 1'b0 ;
  assign n15438 = n15437 ^ n1164 ^ x87 ;
  assign n15439 = n15438 ^ n12529 ^ n11106 ;
  assign n15445 = n15444 ^ n15441 ^ n15439 ;
  assign n15447 = ( ~n6584 & n8203 ) | ( ~n6584 & n9889 ) | ( n8203 & n9889 ) ;
  assign n15446 = n14358 ^ n11379 ^ n8444 ;
  assign n15448 = n15447 ^ n15446 ^ n4585 ;
  assign n15456 = n6642 & ~n7274 ;
  assign n15457 = ~n10739 & n15456 ;
  assign n15449 = ( n2102 & ~n4880 ) | ( n2102 & n8684 ) | ( ~n4880 & n8684 ) ;
  assign n15450 = n8730 & ~n15449 ;
  assign n15451 = ~n6160 & n6494 ;
  assign n15452 = n15451 ^ n4540 ^ n767 ;
  assign n15453 = n15452 ^ n4460 ^ 1'b0 ;
  assign n15454 = n15450 & n15453 ;
  assign n15455 = ~n4971 & n15454 ;
  assign n15458 = n15457 ^ n15455 ^ 1'b0 ;
  assign n15459 = n706 & n14050 ;
  assign n15460 = x23 & n15459 ;
  assign n15461 = n15460 ^ n2840 ^ 1'b0 ;
  assign n15462 = n12977 ^ n2968 ^ 1'b0 ;
  assign n15463 = n4528 & ~n15462 ;
  assign n15464 = n15463 ^ n12201 ^ 1'b0 ;
  assign n15465 = n4412 ^ n4000 ^ x47 ;
  assign n15466 = n3274 ^ n3207 ^ 1'b0 ;
  assign n15472 = n7415 & n15361 ;
  assign n15473 = ~n945 & n15472 ;
  assign n15470 = n1654 & ~n6323 ;
  assign n15471 = n15470 ^ n11216 ^ 1'b0 ;
  assign n15467 = ( n412 & ~n967 ) | ( n412 & n6043 ) | ( ~n967 & n6043 ) ;
  assign n15468 = n13919 ^ n8781 ^ n3412 ;
  assign n15469 = ( n1828 & ~n15467 ) | ( n1828 & n15468 ) | ( ~n15467 & n15468 ) ;
  assign n15474 = n15473 ^ n15471 ^ n15469 ;
  assign n15475 = n2751 & ~n5824 ;
  assign n15476 = n168 | n4248 ;
  assign n15477 = n5630 | n15476 ;
  assign n15478 = n1483 & n3088 ;
  assign n15479 = ~n522 & n15478 ;
  assign n15480 = n15479 ^ n6731 ^ 1'b0 ;
  assign n15481 = ( n7551 & ~n15477 ) | ( n7551 & n15480 ) | ( ~n15477 & n15480 ) ;
  assign n15482 = n2760 | n11660 ;
  assign n15483 = n15481 & ~n15482 ;
  assign n15484 = n15483 ^ n413 ^ 1'b0 ;
  assign n15486 = ( n6057 & n7741 ) | ( n6057 & ~n11676 ) | ( n7741 & ~n11676 ) ;
  assign n15487 = ( n6364 & n7760 ) | ( n6364 & n15486 ) | ( n7760 & n15486 ) ;
  assign n15485 = n1248 & n13467 ;
  assign n15488 = n15487 ^ n15485 ^ 1'b0 ;
  assign n15491 = n6862 ^ n3145 ^ 1'b0 ;
  assign n15492 = n6517 | n15491 ;
  assign n15489 = n1795 & ~n3201 ;
  assign n15490 = ~n8232 & n15489 ;
  assign n15493 = n15492 ^ n15490 ^ 1'b0 ;
  assign n15494 = ( n9353 & ~n13530 ) | ( n9353 & n15493 ) | ( ~n13530 & n15493 ) ;
  assign n15495 = ( n2278 & n4315 ) | ( n2278 & n7747 ) | ( n4315 & n7747 ) ;
  assign n15496 = n15495 ^ n7165 ^ 1'b0 ;
  assign n15497 = n12365 ^ n3743 ^ 1'b0 ;
  assign n15498 = n6714 | n15497 ;
  assign n15499 = ( n2733 & ~n12836 ) | ( n2733 & n15498 ) | ( ~n12836 & n15498 ) ;
  assign n15500 = n15496 & n15499 ;
  assign n15501 = ( n3191 & ~n8707 ) | ( n3191 & n11393 ) | ( ~n8707 & n11393 ) ;
  assign n15502 = n15165 ^ n12167 ^ 1'b0 ;
  assign n15503 = n15501 | n15502 ;
  assign n15504 = n6991 ^ n6566 ^ n3869 ;
  assign n15505 = n4574 & n15504 ;
  assign n15506 = n11193 & n15505 ;
  assign n15507 = n2114 & n14644 ;
  assign n15508 = ~n8988 & n15507 ;
  assign n15509 = ( n10632 & ~n15506 ) | ( n10632 & n15508 ) | ( ~n15506 & n15508 ) ;
  assign n15510 = n12056 ^ n3885 ^ n2411 ;
  assign n15511 = n5403 ^ n2095 ^ n1299 ;
  assign n15512 = n15511 ^ n8472 ^ 1'b0 ;
  assign n15513 = ( ~n5408 & n15510 ) | ( ~n5408 & n15512 ) | ( n15510 & n15512 ) ;
  assign n15514 = ( n1577 & ~n6513 ) | ( n1577 & n8778 ) | ( ~n6513 & n8778 ) ;
  assign n15515 = n14711 ^ n2720 ^ 1'b0 ;
  assign n15516 = n15514 & ~n15515 ;
  assign n15517 = ~n11244 & n13406 ;
  assign n15518 = n15517 ^ n14293 ^ 1'b0 ;
  assign n15519 = ( ~n340 & n4534 ) | ( ~n340 & n6941 ) | ( n4534 & n6941 ) ;
  assign n15520 = n4245 & ~n7419 ;
  assign n15521 = n15520 ^ n1477 ^ 1'b0 ;
  assign n15522 = ( n1324 & ~n15519 ) | ( n1324 & n15521 ) | ( ~n15519 & n15521 ) ;
  assign n15523 = n6596 & n15522 ;
  assign n15524 = n3307 & n15523 ;
  assign n15525 = n15524 ^ n7753 ^ n5837 ;
  assign n15526 = n15525 ^ n10953 ^ n2723 ;
  assign n15527 = n7039 & n10634 ;
  assign n15528 = n15527 ^ n7419 ^ 1'b0 ;
  assign n15529 = n2625 | n6849 ;
  assign n15530 = n14029 & ~n15529 ;
  assign n15531 = ( n2847 & ~n7971 ) | ( n2847 & n15530 ) | ( ~n7971 & n15530 ) ;
  assign n15532 = ( n3234 & n8074 ) | ( n3234 & n15531 ) | ( n8074 & n15531 ) ;
  assign n15533 = n6302 & ~n15532 ;
  assign n15539 = n335 & n8550 ;
  assign n15540 = n9712 & n15539 ;
  assign n15535 = ( n1924 & ~n4546 ) | ( n1924 & n8408 ) | ( ~n4546 & n8408 ) ;
  assign n15536 = n15535 ^ n2154 ^ 1'b0 ;
  assign n15534 = ( n1711 & n5552 ) | ( n1711 & n8378 ) | ( n5552 & n8378 ) ;
  assign n15537 = n15536 ^ n15534 ^ 1'b0 ;
  assign n15538 = n1362 & ~n15537 ;
  assign n15541 = n15540 ^ n15538 ^ 1'b0 ;
  assign n15542 = ( n1001 & n6223 ) | ( n1001 & ~n7994 ) | ( n6223 & ~n7994 ) ;
  assign n15543 = n8129 ^ n863 ^ 1'b0 ;
  assign n15544 = n15542 | n15543 ;
  assign n15545 = n7651 ^ n3078 ^ 1'b0 ;
  assign n15546 = ( n1729 & ~n13010 ) | ( n1729 & n15545 ) | ( ~n13010 & n15545 ) ;
  assign n15547 = n6617 & n15546 ;
  assign n15548 = n8032 | n13966 ;
  assign n15549 = n6915 | n15548 ;
  assign n15550 = ( n3026 & n4640 ) | ( n3026 & ~n9105 ) | ( n4640 & ~n9105 ) ;
  assign n15551 = ( ~n2940 & n15549 ) | ( ~n2940 & n15550 ) | ( n15549 & n15550 ) ;
  assign n15552 = n8738 & n11142 ;
  assign n15553 = ~n14511 & n15552 ;
  assign n15554 = ( ~n652 & n2633 ) | ( ~n652 & n3207 ) | ( n2633 & n3207 ) ;
  assign n15555 = n7144 ^ n6164 ^ 1'b0 ;
  assign n15556 = n15555 ^ n3796 ^ x100 ;
  assign n15557 = n15556 ^ n890 ^ 1'b0 ;
  assign n15558 = ~n2537 & n15557 ;
  assign n15559 = n15554 & n15558 ;
  assign n15560 = n15559 ^ n15379 ^ 1'b0 ;
  assign n15561 = n11054 ^ n1583 ^ 1'b0 ;
  assign n15562 = ( x30 & n6215 ) | ( x30 & n11855 ) | ( n6215 & n11855 ) ;
  assign n15563 = n15562 ^ n11164 ^ 1'b0 ;
  assign n15564 = n13146 ^ n9915 ^ n2073 ;
  assign n15565 = n5864 ^ n1896 ^ n1315 ;
  assign n15566 = n3748 & ~n5718 ;
  assign n15567 = n15566 ^ n3157 ^ 1'b0 ;
  assign n15568 = n15565 & ~n15567 ;
  assign n15569 = n15568 ^ n5779 ^ 1'b0 ;
  assign n15570 = ~n11603 & n15569 ;
  assign n15571 = n15570 ^ n14197 ^ 1'b0 ;
  assign n15572 = n15571 ^ n2511 ^ n670 ;
  assign n15573 = n867 | n8153 ;
  assign n15574 = n2410 | n15573 ;
  assign n15575 = ~n7482 & n15574 ;
  assign n15576 = n15575 ^ n9646 ^ 1'b0 ;
  assign n15577 = ( ~n1870 & n3843 ) | ( ~n1870 & n15576 ) | ( n3843 & n15576 ) ;
  assign n15578 = n13914 ^ n8269 ^ n7378 ;
  assign n15579 = ~n3359 & n6235 ;
  assign n15580 = n570 & n1668 ;
  assign n15581 = ( n4332 & n4778 ) | ( n4332 & ~n15580 ) | ( n4778 & ~n15580 ) ;
  assign n15582 = n13055 & n15581 ;
  assign n15583 = ( ~n15578 & n15579 ) | ( ~n15578 & n15582 ) | ( n15579 & n15582 ) ;
  assign n15584 = n14080 ^ n6599 ^ n6053 ;
  assign n15585 = n7733 & ~n10020 ;
  assign n15586 = n1151 | n9793 ;
  assign n15587 = ~n1480 & n15586 ;
  assign n15588 = n6674 | n11182 ;
  assign n15589 = n15587 | n15588 ;
  assign n15590 = n15589 ^ n6066 ^ 1'b0 ;
  assign n15591 = n15585 & ~n15590 ;
  assign n15592 = n10824 ^ n10753 ^ n8577 ;
  assign n15593 = ( n2088 & ~n3209 ) | ( n2088 & n3297 ) | ( ~n3209 & n3297 ) ;
  assign n15594 = n15593 ^ n4638 ^ 1'b0 ;
  assign n15595 = n2120 & n14236 ;
  assign n15597 = n10413 & ~n13457 ;
  assign n15598 = n10484 & n15597 ;
  assign n15596 = n5680 ^ n4611 ^ 1'b0 ;
  assign n15599 = n15598 ^ n15596 ^ 1'b0 ;
  assign n15600 = ~n5587 & n15599 ;
  assign n15601 = n954 & n1276 ;
  assign n15602 = n15601 ^ n2323 ^ 1'b0 ;
  assign n15603 = n15600 & ~n15602 ;
  assign n15604 = n7814 ^ n1945 ^ 1'b0 ;
  assign n15605 = n15604 ^ n10847 ^ n7349 ;
  assign n15606 = n2501 & ~n15605 ;
  assign n15607 = n2365 & ~n11811 ;
  assign n15608 = n15607 ^ n5773 ^ 1'b0 ;
  assign n15609 = n15608 ^ n15222 ^ n7873 ;
  assign n15610 = n15510 ^ n4190 ^ 1'b0 ;
  assign n15611 = n15610 ^ n14582 ^ n6255 ;
  assign n15612 = n4280 | n6106 ;
  assign n15613 = n7452 ^ n3129 ^ n787 ;
  assign n15614 = n3724 | n15613 ;
  assign n15615 = n15614 ^ n5475 ^ 1'b0 ;
  assign n15619 = n3938 ^ n3461 ^ 1'b0 ;
  assign n15620 = ( ~n9590 & n12139 ) | ( ~n9590 & n15619 ) | ( n12139 & n15619 ) ;
  assign n15617 = n9339 ^ n897 ^ 1'b0 ;
  assign n15618 = ( n1070 & ~n9353 ) | ( n1070 & n15617 ) | ( ~n9353 & n15617 ) ;
  assign n15621 = n15620 ^ n15618 ^ n12530 ;
  assign n15616 = n5607 ^ n4267 ^ 1'b0 ;
  assign n15622 = n15621 ^ n15616 ^ 1'b0 ;
  assign n15623 = ~n9181 & n15622 ;
  assign n15624 = n4051 ^ n412 ^ 1'b0 ;
  assign n15625 = n2120 | n15624 ;
  assign n15626 = n3567 & n5551 ;
  assign n15627 = n11653 ^ n7909 ^ 1'b0 ;
  assign n15628 = n13891 & ~n15627 ;
  assign n15629 = n15628 ^ n12281 ^ 1'b0 ;
  assign n15630 = ~n15626 & n15629 ;
  assign n15631 = ~n3249 & n6038 ;
  assign n15632 = n13721 & ~n15631 ;
  assign n15633 = n15632 ^ n6553 ^ 1'b0 ;
  assign n15634 = n15633 ^ n6729 ^ n3439 ;
  assign n15635 = ( ~n557 & n3182 ) | ( ~n557 & n9076 ) | ( n3182 & n9076 ) ;
  assign n15636 = ( n4190 & ~n13430 ) | ( n4190 & n15635 ) | ( ~n13430 & n15635 ) ;
  assign n15637 = ( ~n850 & n13585 ) | ( ~n850 & n15636 ) | ( n13585 & n15636 ) ;
  assign n15638 = n5507 & n6414 ;
  assign n15639 = ( ~n179 & n8688 ) | ( ~n179 & n9611 ) | ( n8688 & n9611 ) ;
  assign n15640 = n11864 ^ n544 ^ 1'b0 ;
  assign n15641 = ~n9918 & n15640 ;
  assign n15642 = n15641 ^ n3657 ^ 1'b0 ;
  assign n15643 = n15639 | n15642 ;
  assign n15644 = ( n1316 & ~n9787 ) | ( n1316 & n15001 ) | ( ~n9787 & n15001 ) ;
  assign n15645 = n15644 ^ n11507 ^ 1'b0 ;
  assign n15646 = ( n6406 & ~n7158 ) | ( n6406 & n13367 ) | ( ~n7158 & n13367 ) ;
  assign n15647 = n5777 ^ n5455 ^ n2549 ;
  assign n15648 = n10656 | n15647 ;
  assign n15649 = ( n6108 & n15646 ) | ( n6108 & ~n15648 ) | ( n15646 & ~n15648 ) ;
  assign n15650 = n10107 ^ n7224 ^ n4538 ;
  assign n15651 = n13699 ^ n3830 ^ 1'b0 ;
  assign n15652 = ~n459 & n4273 ;
  assign n15653 = n15652 ^ n2882 ^ 1'b0 ;
  assign n15654 = n15653 ^ n12608 ^ n10374 ;
  assign n15655 = n5129 ^ n1432 ^ n1243 ;
  assign n15656 = n10449 ^ n8701 ^ 1'b0 ;
  assign n15657 = n10046 & n15656 ;
  assign n15658 = n10861 & ~n12411 ;
  assign n15659 = n15658 ^ n691 ^ 1'b0 ;
  assign n15660 = n15657 & n15659 ;
  assign n15661 = n15660 ^ n11986 ^ 1'b0 ;
  assign n15662 = n13482 ^ n4217 ^ 1'b0 ;
  assign n15663 = n15662 ^ n10742 ^ n9305 ;
  assign n15664 = ( n15655 & n15661 ) | ( n15655 & ~n15663 ) | ( n15661 & ~n15663 ) ;
  assign n15665 = n2929 | n14525 ;
  assign n15666 = ~n5538 & n15665 ;
  assign n15667 = n5297 ^ n3071 ^ 1'b0 ;
  assign n15668 = n15667 ^ n2573 ^ 1'b0 ;
  assign n15669 = n2704 & n15668 ;
  assign n15670 = n15669 ^ n7426 ^ n3352 ;
  assign n15671 = n15670 ^ n13121 ^ 1'b0 ;
  assign n15672 = n2051 & ~n15671 ;
  assign n15679 = ( n2295 & n4862 ) | ( n2295 & ~n9448 ) | ( n4862 & ~n9448 ) ;
  assign n15673 = n2853 | n5540 ;
  assign n15674 = n11000 & n15673 ;
  assign n15675 = ~n8541 & n15674 ;
  assign n15676 = n15675 ^ n2324 ^ 1'b0 ;
  assign n15677 = n1571 | n7202 ;
  assign n15678 = n15676 | n15677 ;
  assign n15680 = n15679 ^ n15678 ^ 1'b0 ;
  assign n15681 = n7651 ^ n3498 ^ 1'b0 ;
  assign n15682 = n887 & ~n7619 ;
  assign n15683 = n8251 ^ n4256 ^ 1'b0 ;
  assign n15684 = ( n9850 & ~n10136 ) | ( n9850 & n15683 ) | ( ~n10136 & n15683 ) ;
  assign n15685 = n15684 ^ n11332 ^ n2724 ;
  assign n15686 = ( n15681 & n15682 ) | ( n15681 & ~n15685 ) | ( n15682 & ~n15685 ) ;
  assign n15687 = n11512 ^ n6006 ^ 1'b0 ;
  assign n15688 = ( ~n2549 & n3336 ) | ( ~n2549 & n10487 ) | ( n3336 & n10487 ) ;
  assign n15689 = n4612 | n15688 ;
  assign n15690 = ( n2494 & n3286 ) | ( n2494 & n6754 ) | ( n3286 & n6754 ) ;
  assign n15691 = n15690 ^ n12396 ^ 1'b0 ;
  assign n15692 = n7205 | n15691 ;
  assign n15693 = ( n313 & n1933 ) | ( n313 & n3922 ) | ( n1933 & n3922 ) ;
  assign n15694 = ( n399 & ~n11123 ) | ( n399 & n15693 ) | ( ~n11123 & n15693 ) ;
  assign n15695 = n15694 ^ n4040 ^ 1'b0 ;
  assign n15696 = n9338 & ~n13532 ;
  assign n15697 = n1494 & ~n3150 ;
  assign n15698 = n1881 & n15697 ;
  assign n15699 = ( ~n409 & n3928 ) | ( ~n409 & n7842 ) | ( n3928 & n7842 ) ;
  assign n15700 = x95 & n10989 ;
  assign n15701 = n15700 ^ n5912 ^ 1'b0 ;
  assign n15702 = n9411 & n10403 ;
  assign n15703 = n15702 ^ n3255 ^ 1'b0 ;
  assign n15704 = n774 & n15703 ;
  assign n15705 = ~n3856 & n8534 ;
  assign n15706 = ( n440 & ~n2436 ) | ( n440 & n15705 ) | ( ~n2436 & n15705 ) ;
  assign n15707 = n15706 ^ n10864 ^ n3230 ;
  assign n15708 = ~n6429 & n15707 ;
  assign n15709 = ~n7858 & n15708 ;
  assign n15710 = n15709 ^ n8255 ^ n4103 ;
  assign n15711 = n15710 ^ n11922 ^ n11505 ;
  assign n15712 = n6551 ^ n5332 ^ 1'b0 ;
  assign n15713 = n11866 ^ n8497 ^ n325 ;
  assign n15714 = n15713 ^ n14818 ^ n9339 ;
  assign n15715 = n15712 & ~n15714 ;
  assign n15716 = n9765 ^ n8366 ^ n1330 ;
  assign n15717 = n13451 & ~n15716 ;
  assign n15718 = ~n13079 & n14385 ;
  assign n15719 = n14903 | n15718 ;
  assign n15720 = n15719 ^ n13179 ^ 1'b0 ;
  assign n15721 = n15273 ^ n7222 ^ 1'b0 ;
  assign n15722 = ~n13775 & n15721 ;
  assign n15723 = n12576 ^ n6919 ^ 1'b0 ;
  assign n15726 = ( n2256 & n11218 ) | ( n2256 & n13036 ) | ( n11218 & n13036 ) ;
  assign n15727 = n15726 ^ n3483 ^ n1907 ;
  assign n15724 = n9728 ^ n8792 ^ 1'b0 ;
  assign n15725 = ( x63 & n8862 ) | ( x63 & ~n15724 ) | ( n8862 & ~n15724 ) ;
  assign n15728 = n15727 ^ n15725 ^ n6773 ;
  assign n15729 = n1522 & n14364 ;
  assign n15730 = n1175 ^ x57 ^ 1'b0 ;
  assign n15731 = n2587 & ~n4409 ;
  assign n15732 = n15730 & n15731 ;
  assign n15733 = n6563 | n13457 ;
  assign n15734 = ( n4274 & ~n10530 ) | ( n4274 & n15733 ) | ( ~n10530 & n15733 ) ;
  assign n15735 = ~n11281 & n15734 ;
  assign n15736 = n4509 ^ n3245 ^ 1'b0 ;
  assign n15737 = n15735 | n15736 ;
  assign n15738 = n3943 & ~n13206 ;
  assign n15743 = n2643 | n3937 ;
  assign n15744 = n15743 ^ n3174 ^ 1'b0 ;
  assign n15739 = n7580 ^ n5031 ^ n4775 ;
  assign n15740 = ( x5 & ~x6 ) | ( x5 & n15739 ) | ( ~x6 & n15739 ) ;
  assign n15741 = ~n360 & n15740 ;
  assign n15742 = n15741 ^ n13498 ^ 1'b0 ;
  assign n15745 = n15744 ^ n15742 ^ n8621 ;
  assign n15746 = n2577 & ~n10764 ;
  assign n15747 = ( n5403 & n6838 ) | ( n5403 & ~n15746 ) | ( n6838 & ~n15746 ) ;
  assign n15748 = n15031 ^ n8849 ^ n2042 ;
  assign n15749 = ( ~n5505 & n9438 ) | ( ~n5505 & n9923 ) | ( n9438 & n9923 ) ;
  assign n15750 = n15749 ^ n11833 ^ n4305 ;
  assign n15751 = n5695 & n10818 ;
  assign n15752 = n15751 ^ n6395 ^ 1'b0 ;
  assign n15753 = ( n4282 & n15123 ) | ( n4282 & ~n15752 ) | ( n15123 & ~n15752 ) ;
  assign n15754 = n4501 | n6466 ;
  assign n15755 = n1923 | n15754 ;
  assign n15756 = n15755 ^ n1318 ^ 1'b0 ;
  assign n15757 = n15756 ^ n9437 ^ 1'b0 ;
  assign n15758 = n15757 ^ n6991 ^ 1'b0 ;
  assign n15759 = n8292 ^ n7205 ^ n2592 ;
  assign n15760 = n14591 ^ n5123 ^ n4396 ;
  assign n15761 = n621 | n15760 ;
  assign n15762 = n15761 ^ n1468 ^ 1'b0 ;
  assign n15763 = ( ~n4682 & n15759 ) | ( ~n4682 & n15762 ) | ( n15759 & n15762 ) ;
  assign n15764 = ~n15758 & n15763 ;
  assign n15765 = ~n4108 & n4651 ;
  assign n15766 = ~n15032 & n15765 ;
  assign n15767 = n2348 | n15766 ;
  assign n15768 = n5706 ^ n3175 ^ n2053 ;
  assign n15769 = n15768 ^ n2991 ^ 1'b0 ;
  assign n15770 = n12217 ^ n7790 ^ n7015 ;
  assign n15771 = ( n11398 & ~n15769 ) | ( n11398 & n15770 ) | ( ~n15769 & n15770 ) ;
  assign n15772 = n12231 ^ n2688 ^ n1878 ;
  assign n15773 = ( n5278 & n10442 ) | ( n5278 & ~n15772 ) | ( n10442 & ~n15772 ) ;
  assign n15774 = n10105 & ~n13944 ;
  assign n15775 = n15774 ^ n2700 ^ n2440 ;
  assign n15776 = n7780 ^ n2863 ^ 1'b0 ;
  assign n15777 = n15776 ^ n10947 ^ n4253 ;
  assign n15778 = n12914 ^ n11759 ^ n2557 ;
  assign n15779 = n2059 ^ n334 ^ 1'b0 ;
  assign n15780 = ~n15778 & n15779 ;
  assign n15781 = n4632 & n6543 ;
  assign n15782 = n3759 ^ n3124 ^ 1'b0 ;
  assign n15783 = n11585 ^ n9184 ^ 1'b0 ;
  assign n15784 = n5659 & n15783 ;
  assign n15785 = ( x110 & ~n1698 ) | ( x110 & n6475 ) | ( ~n1698 & n6475 ) ;
  assign n15786 = n3080 & ~n14971 ;
  assign n15791 = n7232 ^ n6043 ^ n4344 ;
  assign n15787 = n14115 ^ n11128 ^ 1'b0 ;
  assign n15788 = n4680 & ~n15787 ;
  assign n15789 = ~n13360 & n15788 ;
  assign n15790 = n15789 ^ n5661 ^ 1'b0 ;
  assign n15792 = n15791 ^ n15790 ^ 1'b0 ;
  assign n15793 = n1459 & ~n6741 ;
  assign n15794 = ( ~n7588 & n15792 ) | ( ~n7588 & n15793 ) | ( n15792 & n15793 ) ;
  assign n15795 = n10762 ^ n10407 ^ n4486 ;
  assign n15796 = n9229 | n15795 ;
  assign n15797 = ( n461 & n13687 ) | ( n461 & ~n15796 ) | ( n13687 & ~n15796 ) ;
  assign n15798 = n13745 ^ n2985 ^ 1'b0 ;
  assign n15799 = n12569 & n15798 ;
  assign n15800 = n900 ^ n250 ^ 1'b0 ;
  assign n15801 = n15800 ^ n980 ^ 1'b0 ;
  assign n15802 = ( n5167 & n13384 ) | ( n5167 & ~n15801 ) | ( n13384 & ~n15801 ) ;
  assign n15803 = n13231 ^ n11726 ^ 1'b0 ;
  assign n15805 = n1987 ^ n545 ^ 1'b0 ;
  assign n15804 = n924 & n14958 ;
  assign n15806 = n15805 ^ n15804 ^ 1'b0 ;
  assign n15807 = ( n1284 & n3284 ) | ( n1284 & ~n12774 ) | ( n3284 & ~n12774 ) ;
  assign n15808 = x91 & ~n15807 ;
  assign n15809 = ( ~x74 & n1118 ) | ( ~x74 & n13750 ) | ( n1118 & n13750 ) ;
  assign n15810 = n2978 & ~n15809 ;
  assign n15811 = n15810 ^ n4826 ^ 1'b0 ;
  assign n15812 = n3912 ^ n777 ^ 1'b0 ;
  assign n15813 = n15812 ^ n10656 ^ n234 ;
  assign n15814 = n15813 ^ n12356 ^ 1'b0 ;
  assign n15815 = n7620 & ~n15814 ;
  assign n15816 = ( n11573 & n13307 ) | ( n11573 & n15815 ) | ( n13307 & n15815 ) ;
  assign n15817 = ( n1732 & n7407 ) | ( n1732 & ~n15816 ) | ( n7407 & ~n15816 ) ;
  assign n15821 = n3671 ^ n2415 ^ x121 ;
  assign n15818 = n5419 ^ n557 ^ 1'b0 ;
  assign n15819 = ( n5504 & n9890 ) | ( n5504 & ~n13008 ) | ( n9890 & ~n13008 ) ;
  assign n15820 = n15818 & n15819 ;
  assign n15822 = n15821 ^ n15820 ^ n10291 ;
  assign n15823 = n13066 ^ n6456 ^ 1'b0 ;
  assign n15824 = ( n2771 & n5753 ) | ( n2771 & ~n15823 ) | ( n5753 & ~n15823 ) ;
  assign n15825 = n726 & n15824 ;
  assign n15826 = ~n9605 & n15825 ;
  assign n15827 = n14510 ^ n859 ^ 1'b0 ;
  assign n15828 = n15827 ^ n15404 ^ n1736 ;
  assign n15829 = n10365 & n15828 ;
  assign n15830 = n11052 ^ n7360 ^ n4537 ;
  assign n15831 = n12610 ^ n11112 ^ 1'b0 ;
  assign n15832 = n15028 ^ n2667 ^ 1'b0 ;
  assign n15833 = ~n12208 & n15832 ;
  assign n15834 = n10845 ^ n149 ^ 1'b0 ;
  assign n15835 = n12973 ^ n11693 ^ n10175 ;
  assign n15836 = ( ~n5302 & n9667 ) | ( ~n5302 & n15835 ) | ( n9667 & n15835 ) ;
  assign n15837 = n15836 ^ n13914 ^ n6166 ;
  assign n15838 = ( n3775 & n7674 ) | ( n3775 & n13240 ) | ( n7674 & n13240 ) ;
  assign n15839 = n2817 | n15838 ;
  assign n15840 = n15839 ^ n14412 ^ 1'b0 ;
  assign n15841 = n167 & n15840 ;
  assign n15842 = n15841 ^ n6391 ^ 1'b0 ;
  assign n15843 = n14634 ^ n14587 ^ n3512 ;
  assign n15844 = n1850 & n2485 ;
  assign n15845 = ~n7479 & n15844 ;
  assign n15846 = n180 | n15845 ;
  assign n15847 = n4320 & n14064 ;
  assign n15848 = ( n2045 & n15555 ) | ( n2045 & ~n15847 ) | ( n15555 & ~n15847 ) ;
  assign n15849 = n9679 ^ n5068 ^ 1'b0 ;
  assign n15850 = n1857 & ~n15849 ;
  assign n15851 = n5195 ^ n4405 ^ 1'b0 ;
  assign n15852 = n15850 & n15851 ;
  assign n15853 = n2873 & n15852 ;
  assign n15854 = ~n15848 & n15853 ;
  assign n15855 = ~n5448 & n12177 ;
  assign n15856 = ~n15854 & n15855 ;
  assign n15857 = n15856 ^ n11838 ^ 1'b0 ;
  assign n15858 = n3405 & n9344 ;
  assign n15859 = ~n6952 & n15858 ;
  assign n15860 = n8126 ^ n6399 ^ 1'b0 ;
  assign n15861 = n3091 & n15860 ;
  assign n15862 = n15861 ^ n9485 ^ 1'b0 ;
  assign n15863 = n10953 ^ n495 ^ 1'b0 ;
  assign n15864 = n15862 | n15863 ;
  assign n15865 = n10481 ^ n9144 ^ n406 ;
  assign n15867 = n9195 & n12297 ;
  assign n15866 = n15236 ^ n10861 ^ n6857 ;
  assign n15868 = n15867 ^ n15866 ^ 1'b0 ;
  assign n15869 = n5821 & n15868 ;
  assign n15870 = ( n12612 & n15865 ) | ( n12612 & n15869 ) | ( n15865 & n15869 ) ;
  assign n15871 = n3761 ^ n1261 ^ 1'b0 ;
  assign n15872 = n5670 ^ n1516 ^ 1'b0 ;
  assign n15873 = ~n15871 & n15872 ;
  assign n15874 = n5154 ^ n3984 ^ n2459 ;
  assign n15875 = n15874 ^ n13321 ^ n4404 ;
  assign n15876 = ( n4295 & ~n15873 ) | ( n4295 & n15875 ) | ( ~n15873 & n15875 ) ;
  assign n15877 = n15876 ^ n1216 ^ 1'b0 ;
  assign n15878 = n4128 & ~n13967 ;
  assign n15879 = n15878 ^ n2301 ^ 1'b0 ;
  assign n15880 = ( n2119 & ~n4715 ) | ( n2119 & n5224 ) | ( ~n4715 & n5224 ) ;
  assign n15881 = n15880 ^ n10930 ^ n633 ;
  assign n15882 = n10101 ^ n5670 ^ n1450 ;
  assign n15883 = n5664 ^ n1375 ^ 1'b0 ;
  assign n15884 = n2405 & n5965 ;
  assign n15885 = n15884 ^ n1654 ^ 1'b0 ;
  assign n15886 = ~n8149 & n13906 ;
  assign n15887 = n6202 & ~n7228 ;
  assign n15888 = n7627 ^ n5300 ^ n530 ;
  assign n15889 = n6002 & ~n10161 ;
  assign n15890 = ( n15887 & n15888 ) | ( n15887 & ~n15889 ) | ( n15888 & ~n15889 ) ;
  assign n15898 = ( n1809 & ~n5292 ) | ( n1809 & n10661 ) | ( ~n5292 & n10661 ) ;
  assign n15893 = n3012 ^ x23 ^ 1'b0 ;
  assign n15894 = ( n179 & ~n1122 ) | ( n179 & n15893 ) | ( ~n1122 & n15893 ) ;
  assign n15891 = ~n1111 & n12571 ;
  assign n15892 = ~n5266 & n15891 ;
  assign n15895 = n15894 ^ n15892 ^ n10122 ;
  assign n15896 = n3895 & ~n15895 ;
  assign n15897 = ~n3498 & n15896 ;
  assign n15899 = n15898 ^ n15897 ^ n238 ;
  assign n15902 = n13597 ^ n863 ^ 1'b0 ;
  assign n15903 = ~n3712 & n15902 ;
  assign n15900 = n12331 ^ n12056 ^ n179 ;
  assign n15901 = ( n7508 & ~n11749 ) | ( n7508 & n15900 ) | ( ~n11749 & n15900 ) ;
  assign n15904 = n15903 ^ n15901 ^ n4411 ;
  assign n15905 = n11139 & ~n15350 ;
  assign n15906 = n15905 ^ n12890 ^ 1'b0 ;
  assign n15911 = n2269 | n4017 ;
  assign n15912 = ~n991 & n10567 ;
  assign n15913 = ~n15911 & n15912 ;
  assign n15909 = ( n1146 & n3359 ) | ( n1146 & ~n10342 ) | ( n3359 & ~n10342 ) ;
  assign n15907 = n1800 | n13296 ;
  assign n15908 = n4713 | n15907 ;
  assign n15910 = n15909 ^ n15908 ^ n3118 ;
  assign n15914 = n15913 ^ n15910 ^ 1'b0 ;
  assign n15915 = n3543 & ~n15914 ;
  assign n15916 = n1049 & n3088 ;
  assign n15917 = n1933 & n15916 ;
  assign n15921 = ~n3037 & n6751 ;
  assign n15918 = n13532 ^ n8354 ^ n5037 ;
  assign n15919 = n3930 ^ n632 ^ 1'b0 ;
  assign n15920 = n15918 & n15919 ;
  assign n15922 = n15921 ^ n15920 ^ 1'b0 ;
  assign n15923 = n2205 & ~n15922 ;
  assign n15924 = ~n15917 & n15923 ;
  assign n15925 = n15924 ^ n9635 ^ 1'b0 ;
  assign n15926 = n5849 | n15925 ;
  assign n15927 = n15926 ^ n2957 ^ 1'b0 ;
  assign n15929 = n4842 | n5628 ;
  assign n15930 = n1332 | n15929 ;
  assign n15928 = ( n3027 & n3285 ) | ( n3027 & ~n8964 ) | ( n3285 & ~n8964 ) ;
  assign n15931 = n15930 ^ n15928 ^ n1313 ;
  assign n15932 = ( n6295 & ~n6588 ) | ( n6295 & n13036 ) | ( ~n6588 & n13036 ) ;
  assign n15933 = n15932 ^ n9208 ^ n3938 ;
  assign n15934 = n15933 ^ n15693 ^ 1'b0 ;
  assign n15935 = n7615 ^ n2653 ^ 1'b0 ;
  assign n15936 = n10919 ^ n5835 ^ n1388 ;
  assign n15937 = n9953 ^ n601 ^ 1'b0 ;
  assign n15938 = n9427 & ~n15937 ;
  assign n15939 = n15938 ^ n8087 ^ n1008 ;
  assign n15940 = ( ~n8172 & n8752 ) | ( ~n8172 & n14472 ) | ( n8752 & n14472 ) ;
  assign n15941 = ( ~n4293 & n8015 ) | ( ~n4293 & n10090 ) | ( n8015 & n10090 ) ;
  assign n15942 = ( ~n2132 & n5467 ) | ( ~n2132 & n7331 ) | ( n5467 & n7331 ) ;
  assign n15943 = n15574 & ~n15942 ;
  assign n15944 = n15943 ^ n11769 ^ n6973 ;
  assign n15945 = n15631 ^ n10636 ^ 1'b0 ;
  assign n15946 = n1199 & ~n15945 ;
  assign n15950 = n8959 ^ n2440 ^ 1'b0 ;
  assign n15951 = n311 | n15950 ;
  assign n15952 = n15951 ^ n7979 ^ n5031 ;
  assign n15948 = n6371 ^ n3794 ^ 1'b0 ;
  assign n15949 = n15948 ^ n15860 ^ n10903 ;
  assign n15953 = n15952 ^ n15949 ^ n14735 ;
  assign n15947 = n5106 | n10856 ;
  assign n15954 = n15953 ^ n15947 ^ 1'b0 ;
  assign n15955 = ( n6558 & n15946 ) | ( n6558 & ~n15954 ) | ( n15946 & ~n15954 ) ;
  assign n15956 = ( n7369 & n15944 ) | ( n7369 & n15955 ) | ( n15944 & n15955 ) ;
  assign n15957 = n4180 & n7531 ;
  assign n15958 = n5480 & n15957 ;
  assign n15959 = n14601 ^ n6274 ^ n3787 ;
  assign n15960 = n15959 ^ n3720 ^ 1'b0 ;
  assign n15961 = ( n4185 & n5050 ) | ( n4185 & n5705 ) | ( n5050 & n5705 ) ;
  assign n15962 = ( n14062 & n15149 ) | ( n14062 & ~n15961 ) | ( n15149 & ~n15961 ) ;
  assign n15963 = ( n3593 & n6588 ) | ( n3593 & ~n8889 ) | ( n6588 & ~n8889 ) ;
  assign n15964 = n10567 & ~n15963 ;
  assign n15965 = n15964 ^ n14965 ^ 1'b0 ;
  assign n15966 = n7697 ^ n5763 ^ 1'b0 ;
  assign n15967 = n15386 & ~n15966 ;
  assign n15968 = n7655 & n8272 ;
  assign n15969 = n11101 ^ n3643 ^ 1'b0 ;
  assign n15972 = n7735 ^ n7273 ^ 1'b0 ;
  assign n15970 = ~n1494 & n3294 ;
  assign n15971 = ~n14954 & n15970 ;
  assign n15973 = n15972 ^ n15971 ^ n2262 ;
  assign n15974 = ( n2614 & n9438 ) | ( n2614 & ~n11569 ) | ( n9438 & ~n11569 ) ;
  assign n15975 = n2204 & ~n5026 ;
  assign n15976 = ~n13591 & n15975 ;
  assign n15977 = n12410 ^ n5708 ^ 1'b0 ;
  assign n15978 = n6750 | n15977 ;
  assign n15984 = n1100 & ~n1522 ;
  assign n15985 = ~n780 & n15984 ;
  assign n15986 = n15985 ^ n3225 ^ 1'b0 ;
  assign n15979 = n7806 ^ n4450 ^ n3341 ;
  assign n15980 = n11295 ^ n7224 ^ n3569 ;
  assign n15981 = n11128 ^ n10216 ^ 1'b0 ;
  assign n15982 = n15980 & ~n15981 ;
  assign n15983 = ( n5691 & n15979 ) | ( n5691 & ~n15982 ) | ( n15979 & ~n15982 ) ;
  assign n15987 = n15986 ^ n15983 ^ n8253 ;
  assign n15988 = ( n6803 & n9631 ) | ( n6803 & ~n13800 ) | ( n9631 & ~n13800 ) ;
  assign n15989 = n4888 & ~n15639 ;
  assign n15990 = n15989 ^ n11038 ^ 1'b0 ;
  assign n15991 = n7194 ^ n254 ^ 1'b0 ;
  assign n15992 = ( ~n5116 & n5451 ) | ( ~n5116 & n15991 ) | ( n5451 & n15991 ) ;
  assign n15993 = ( ~n159 & n7748 ) | ( ~n159 & n10603 ) | ( n7748 & n10603 ) ;
  assign n15994 = n15993 ^ n13227 ^ n10920 ;
  assign n15995 = n8959 ^ n1299 ^ 1'b0 ;
  assign n15996 = n14038 & n15995 ;
  assign n15997 = n15996 ^ n667 ^ n360 ;
  assign n15998 = n7228 ^ n4645 ^ 1'b0 ;
  assign n15999 = ( n1519 & n2303 ) | ( n1519 & n15998 ) | ( n2303 & n15998 ) ;
  assign n16000 = n4889 & n13625 ;
  assign n16001 = n13914 ^ n6330 ^ n4033 ;
  assign n16002 = n16001 ^ n7618 ^ n286 ;
  assign n16003 = n15848 & n16002 ;
  assign n16004 = n2870 | n12337 ;
  assign n16005 = n282 & n3752 ;
  assign n16006 = n16005 ^ n3371 ^ 1'b0 ;
  assign n16007 = n16006 ^ n14950 ^ 1'b0 ;
  assign n16008 = n8556 ^ n5412 ^ 1'b0 ;
  assign n16009 = n8139 ^ n5522 ^ n3892 ;
  assign n16010 = ~n2257 & n2274 ;
  assign n16011 = n7562 & n16010 ;
  assign n16012 = n1049 & n3376 ;
  assign n16013 = n16012 ^ n1980 ^ 1'b0 ;
  assign n16014 = ( n16009 & n16011 ) | ( n16009 & n16013 ) | ( n16011 & n16013 ) ;
  assign n16015 = n16008 | n16014 ;
  assign n16016 = n1568 | n16015 ;
  assign n16017 = ( n5126 & n8186 ) | ( n5126 & n10203 ) | ( n8186 & n10203 ) ;
  assign n16018 = n3917 ^ n2253 ^ n397 ;
  assign n16019 = n16018 ^ n5515 ^ 1'b0 ;
  assign n16020 = n3307 & n16019 ;
  assign n16022 = n1703 & n13035 ;
  assign n16023 = n16022 ^ n11538 ^ 1'b0 ;
  assign n16021 = n6139 | n7031 ;
  assign n16024 = n16023 ^ n16021 ^ 1'b0 ;
  assign n16031 = n9584 ^ n8272 ^ n3468 ;
  assign n16025 = ( x52 & n1754 ) | ( x52 & ~n2254 ) | ( n1754 & ~n2254 ) ;
  assign n16026 = n16025 ^ n5702 ^ 1'b0 ;
  assign n16027 = n6155 ^ n5452 ^ 1'b0 ;
  assign n16028 = n16027 ^ n522 ^ x37 ;
  assign n16029 = n8460 & ~n16028 ;
  assign n16030 = n16026 & n16029 ;
  assign n16032 = n16031 ^ n16030 ^ 1'b0 ;
  assign n16033 = ~n5898 & n16032 ;
  assign n16034 = ~n5314 & n9167 ;
  assign n16035 = ~n3033 & n16034 ;
  assign n16036 = ( n652 & ~n3036 ) | ( n652 & n4617 ) | ( ~n3036 & n4617 ) ;
  assign n16037 = n16035 & ~n16036 ;
  assign n16038 = n16037 ^ n6895 ^ n3335 ;
  assign n16042 = ( n1865 & n12712 ) | ( n1865 & n13851 ) | ( n12712 & n13851 ) ;
  assign n16039 = n2061 & n7414 ;
  assign n16040 = n16039 ^ n12120 ^ 1'b0 ;
  assign n16041 = ( n4157 & ~n8175 ) | ( n4157 & n16040 ) | ( ~n8175 & n16040 ) ;
  assign n16043 = n16042 ^ n16041 ^ n4803 ;
  assign n16044 = n11259 ^ n7536 ^ n2539 ;
  assign n16045 = ( n6353 & ~n14868 ) | ( n6353 & n16044 ) | ( ~n14868 & n16044 ) ;
  assign n16046 = n16045 ^ n5694 ^ n3723 ;
  assign n16047 = n8461 ^ n3432 ^ 1'b0 ;
  assign n16048 = ~n5672 & n16047 ;
  assign n16049 = ( n2579 & n5277 ) | ( n2579 & ~n6221 ) | ( n5277 & ~n6221 ) ;
  assign n16050 = ( n14261 & ~n16048 ) | ( n14261 & n16049 ) | ( ~n16048 & n16049 ) ;
  assign n16051 = n6106 | n8660 ;
  assign n16052 = n4240 | n16051 ;
  assign n16053 = n1456 & n16052 ;
  assign n16054 = ~n2683 & n16053 ;
  assign n16055 = ( ~n6881 & n10625 ) | ( ~n6881 & n15120 ) | ( n10625 & n15120 ) ;
  assign n16056 = n16055 ^ n147 ^ 1'b0 ;
  assign n16057 = n16054 | n16056 ;
  assign n16058 = n8886 ^ n2716 ^ 1'b0 ;
  assign n16059 = n11975 ^ n8132 ^ n6733 ;
  assign n16060 = n7219 ^ n4759 ^ 1'b0 ;
  assign n16061 = ~n4534 & n16060 ;
  assign n16062 = n2361 & n14233 ;
  assign n16063 = n16062 ^ n14607 ^ 1'b0 ;
  assign n16064 = n5267 | n5602 ;
  assign n16065 = n16064 ^ n3650 ^ 1'b0 ;
  assign n16066 = n14766 ^ n9547 ^ 1'b0 ;
  assign n16067 = ~n16036 & n16066 ;
  assign n16068 = ~n366 & n16067 ;
  assign n16069 = n16065 & n16068 ;
  assign n16070 = n16069 ^ n15495 ^ n12164 ;
  assign n16071 = n8420 ^ n1444 ^ n1034 ;
  assign n16072 = n10702 ^ n685 ^ 1'b0 ;
  assign n16073 = ( n12882 & n16071 ) | ( n12882 & ~n16072 ) | ( n16071 & ~n16072 ) ;
  assign n16074 = ( n7845 & n9676 ) | ( n7845 & ~n13740 ) | ( n9676 & ~n13740 ) ;
  assign n16077 = n10501 ^ n8748 ^ 1'b0 ;
  assign n16075 = n7770 ^ n624 ^ 1'b0 ;
  assign n16076 = ~n8448 & n16075 ;
  assign n16078 = n16077 ^ n16076 ^ n222 ;
  assign n16079 = n9876 ^ n4562 ^ n621 ;
  assign n16080 = ~n7276 & n16079 ;
  assign n16081 = n16080 ^ n1443 ^ 1'b0 ;
  assign n16083 = ~n4307 & n8204 ;
  assign n16082 = n4706 & n9106 ;
  assign n16084 = n16083 ^ n16082 ^ 1'b0 ;
  assign n16085 = n6423 ^ n3253 ^ 1'b0 ;
  assign n16086 = n10910 | n16085 ;
  assign n16087 = n14484 ^ n5767 ^ 1'b0 ;
  assign n16088 = x91 & n16087 ;
  assign n16089 = n13224 ^ n5836 ^ 1'b0 ;
  assign n16090 = n16089 ^ n1083 ^ 1'b0 ;
  assign n16091 = n11053 ^ n5623 ^ 1'b0 ;
  assign n16092 = ( n9206 & n14754 ) | ( n9206 & ~n16091 ) | ( n14754 & ~n16091 ) ;
  assign n16093 = ( n10151 & n16090 ) | ( n10151 & n16092 ) | ( n16090 & n16092 ) ;
  assign n16094 = n342 & ~n3173 ;
  assign n16095 = n16094 ^ n2254 ^ 1'b0 ;
  assign n16096 = ( ~n3713 & n14034 ) | ( ~n3713 & n14941 ) | ( n14034 & n14941 ) ;
  assign n16097 = ( ~n1994 & n4859 ) | ( ~n1994 & n6219 ) | ( n4859 & n6219 ) ;
  assign n16098 = n16097 ^ n12056 ^ n3159 ;
  assign n16099 = ( n2319 & ~n7283 ) | ( n2319 & n13925 ) | ( ~n7283 & n13925 ) ;
  assign n16100 = n3148 ^ n1943 ^ 1'b0 ;
  assign n16101 = n254 & n16100 ;
  assign n16105 = ( n5905 & n6159 ) | ( n5905 & n9934 ) | ( n6159 & n9934 ) ;
  assign n16106 = n6503 | n16105 ;
  assign n16107 = n16106 ^ n4145 ^ n1548 ;
  assign n16102 = ( n1083 & ~n3334 ) | ( n1083 & n13073 ) | ( ~n3334 & n13073 ) ;
  assign n16103 = ( ~n367 & n1217 ) | ( ~n367 & n9487 ) | ( n1217 & n9487 ) ;
  assign n16104 = n16102 & ~n16103 ;
  assign n16108 = n16107 ^ n16104 ^ 1'b0 ;
  assign n16109 = n13234 ^ n3571 ^ n722 ;
  assign n16110 = ~n2079 & n11659 ;
  assign n16111 = ( n7856 & n9836 ) | ( n7856 & ~n16110 ) | ( n9836 & ~n16110 ) ;
  assign n16118 = n4179 ^ n892 ^ n579 ;
  assign n16119 = ~n1477 & n16118 ;
  assign n16112 = n416 & n1153 ;
  assign n16113 = n16112 ^ n5702 ^ 1'b0 ;
  assign n16114 = n11067 ^ n5054 ^ 1'b0 ;
  assign n16115 = n16113 & n16114 ;
  assign n16116 = n12873 ^ n12839 ^ n5592 ;
  assign n16117 = n16115 & n16116 ;
  assign n16120 = n16119 ^ n16117 ^ 1'b0 ;
  assign n16121 = n13764 ^ n9681 ^ n7049 ;
  assign n16122 = n16121 ^ n15788 ^ n14744 ;
  assign n16123 = n14302 & ~n16122 ;
  assign n16124 = ( x104 & ~n6237 ) | ( x104 & n10128 ) | ( ~n6237 & n10128 ) ;
  assign n16125 = n16124 ^ n4539 ^ 1'b0 ;
  assign n16126 = n12932 ^ n8177 ^ 1'b0 ;
  assign n16127 = ~n16125 & n16126 ;
  assign n16130 = ~n5698 & n6699 ;
  assign n16128 = ( ~n1574 & n4420 ) | ( ~n1574 & n5296 ) | ( n4420 & n5296 ) ;
  assign n16129 = n7684 & n16128 ;
  assign n16131 = n16130 ^ n16129 ^ 1'b0 ;
  assign n16132 = ( n1204 & ~n12344 ) | ( n1204 & n16131 ) | ( ~n12344 & n16131 ) ;
  assign n16133 = ~n2385 & n8367 ;
  assign n16134 = n16133 ^ n2798 ^ 1'b0 ;
  assign n16135 = n13777 & n16134 ;
  assign n16136 = ( n2642 & n9485 ) | ( n2642 & ~n13152 ) | ( n9485 & ~n13152 ) ;
  assign n16137 = n16136 ^ n15254 ^ n11958 ;
  assign n16142 = ~n4700 & n14712 ;
  assign n16143 = n16142 ^ n4421 ^ 1'b0 ;
  assign n16144 = n15183 & ~n16143 ;
  assign n16138 = n8180 | n10447 ;
  assign n16139 = n16138 ^ n6596 ^ 1'b0 ;
  assign n16140 = n16139 ^ n13445 ^ n472 ;
  assign n16141 = n15965 & ~n16140 ;
  assign n16145 = n16144 ^ n16141 ^ 1'b0 ;
  assign n16146 = ~n5535 & n9165 ;
  assign n16147 = n16146 ^ n6149 ^ 1'b0 ;
  assign n16148 = n16147 ^ n11846 ^ n10853 ;
  assign n16149 = n16148 ^ n6649 ^ 1'b0 ;
  assign n16150 = n16149 ^ n10401 ^ 1'b0 ;
  assign n16151 = n3121 | n16150 ;
  assign n16152 = n11992 ^ n5232 ^ 1'b0 ;
  assign n16153 = ( n3962 & n15549 ) | ( n3962 & n16152 ) | ( n15549 & n16152 ) ;
  assign n16154 = n5395 | n15604 ;
  assign n16155 = n16054 ^ n10819 ^ 1'b0 ;
  assign n16156 = n15778 ^ n10551 ^ 1'b0 ;
  assign n16157 = n3629 | n4028 ;
  assign n16158 = n16157 ^ n1707 ^ 1'b0 ;
  assign n16159 = ~n3835 & n16158 ;
  assign n16160 = x68 & n16159 ;
  assign n16161 = n5014 & n9989 ;
  assign n16162 = n13121 & n16161 ;
  assign n16163 = ( n1955 & ~n16160 ) | ( n1955 & n16162 ) | ( ~n16160 & n16162 ) ;
  assign n16164 = n16163 ^ n9405 ^ 1'b0 ;
  assign n16165 = n10263 & ~n16164 ;
  assign n16166 = n1724 | n4788 ;
  assign n16167 = n16165 & n16166 ;
  assign n16168 = ( ~n8121 & n11074 ) | ( ~n8121 & n14728 ) | ( n11074 & n14728 ) ;
  assign n16169 = n11972 ^ n7675 ^ n2484 ;
  assign n16170 = n16169 ^ n3832 ^ 1'b0 ;
  assign n16172 = n895 & n5144 ;
  assign n16173 = ~n2332 & n16172 ;
  assign n16171 = n11155 ^ n5203 ^ n3122 ;
  assign n16174 = n16173 ^ n16171 ^ 1'b0 ;
  assign n16175 = ( ~n2138 & n5384 ) | ( ~n2138 & n10691 ) | ( n5384 & n10691 ) ;
  assign n16176 = n11720 ^ n7648 ^ n5689 ;
  assign n16177 = ( x116 & n1789 ) | ( x116 & n3292 ) | ( n1789 & n3292 ) ;
  assign n16178 = n16177 ^ n13966 ^ 1'b0 ;
  assign n16179 = n13427 ^ n4936 ^ n3693 ;
  assign n16180 = n16179 ^ n1184 ^ 1'b0 ;
  assign n16181 = ~n4490 & n16180 ;
  assign n16182 = ( n3198 & ~n14343 ) | ( n3198 & n16181 ) | ( ~n14343 & n16181 ) ;
  assign n16183 = n8177 ^ n3665 ^ 1'b0 ;
  assign n16184 = n7893 | n11290 ;
  assign n16185 = n16184 ^ n5735 ^ 1'b0 ;
  assign n16186 = ( n1694 & n6356 ) | ( n1694 & ~n16185 ) | ( n6356 & ~n16185 ) ;
  assign n16187 = n16186 ^ n8621 ^ 1'b0 ;
  assign n16188 = ~n15233 & n16187 ;
  assign n16189 = n12095 & n12859 ;
  assign n16190 = n2813 ^ n2429 ^ n1357 ;
  assign n16191 = n2243 & n2378 ;
  assign n16192 = n6766 & n16191 ;
  assign n16193 = ( ~n426 & n5698 ) | ( ~n426 & n16192 ) | ( n5698 & n16192 ) ;
  assign n16194 = n16193 ^ n3141 ^ 1'b0 ;
  assign n16195 = n4125 & n16194 ;
  assign n16196 = ~n3103 & n16195 ;
  assign n16197 = n5934 & n16196 ;
  assign n16198 = ( n4726 & n6078 ) | ( n4726 & n9436 ) | ( n6078 & n9436 ) ;
  assign n16199 = ( n1711 & n8488 ) | ( n1711 & ~n16198 ) | ( n8488 & ~n16198 ) ;
  assign n16200 = n2154 & ~n16199 ;
  assign n16201 = n3567 & n16200 ;
  assign n16202 = ( n15279 & n16197 ) | ( n15279 & ~n16201 ) | ( n16197 & ~n16201 ) ;
  assign n16203 = n16190 & ~n16202 ;
  assign n16204 = n10125 ^ n3490 ^ 1'b0 ;
  assign n16205 = n1660 & n16204 ;
  assign n16206 = n16205 ^ n15146 ^ n4842 ;
  assign n16207 = n15074 ^ n5931 ^ 1'b0 ;
  assign n16208 = n447 | n5521 ;
  assign n16209 = n1991 | n16208 ;
  assign n16210 = ( ~n2706 & n8800 ) | ( ~n2706 & n15340 ) | ( n8800 & n15340 ) ;
  assign n16211 = n7071 | n16210 ;
  assign n16212 = n16209 | n16211 ;
  assign n16213 = n11298 ^ n10216 ^ 1'b0 ;
  assign n16214 = n5391 & ~n16213 ;
  assign n16215 = n4154 & ~n4947 ;
  assign n16216 = n8500 & n16215 ;
  assign n16217 = n10084 ^ n9261 ^ 1'b0 ;
  assign n16218 = n612 & n2409 ;
  assign n16219 = n10288 & n16218 ;
  assign n16220 = n16219 ^ n5181 ^ 1'b0 ;
  assign n16221 = n16220 ^ n14549 ^ n2289 ;
  assign n16222 = n16221 ^ n7104 ^ 1'b0 ;
  assign n16223 = n531 & n16222 ;
  assign n16224 = n16223 ^ n5634 ^ 1'b0 ;
  assign n16225 = n5654 ^ n5285 ^ 1'b0 ;
  assign n16226 = n3932 & n16225 ;
  assign n16227 = ( n16217 & ~n16224 ) | ( n16217 & n16226 ) | ( ~n16224 & n16226 ) ;
  assign n16228 = ( n16214 & n16216 ) | ( n16214 & ~n16227 ) | ( n16216 & ~n16227 ) ;
  assign n16232 = n11400 ^ n3883 ^ 1'b0 ;
  assign n16233 = n10516 & ~n16232 ;
  assign n16234 = ( n13169 & n15850 ) | ( n13169 & ~n16233 ) | ( n15850 & ~n16233 ) ;
  assign n16230 = n12305 ^ n7642 ^ n1205 ;
  assign n16229 = n2484 | n8557 ;
  assign n16231 = n16230 ^ n16229 ^ 1'b0 ;
  assign n16235 = n16234 ^ n16231 ^ n16030 ;
  assign n16236 = n2254 ^ n1500 ^ 1'b0 ;
  assign n16237 = n16236 ^ n9323 ^ 1'b0 ;
  assign n16238 = n3675 & n5651 ;
  assign n16239 = ( ~n943 & n14703 ) | ( ~n943 & n16055 ) | ( n14703 & n16055 ) ;
  assign n16240 = n2914 | n10603 ;
  assign n16241 = n8925 & ~n16240 ;
  assign n16242 = n16239 | n16241 ;
  assign n16243 = n16238 | n16242 ;
  assign n16244 = n4980 & ~n13229 ;
  assign n16245 = ~n13313 & n16244 ;
  assign n16246 = n16245 ^ n15402 ^ 1'b0 ;
  assign n16247 = n4511 & n10368 ;
  assign n16248 = ~n13468 & n16247 ;
  assign n16249 = n12148 | n16248 ;
  assign n16250 = n16249 ^ n12271 ^ 1'b0 ;
  assign n16251 = ~n7155 & n16250 ;
  assign n16252 = ~n753 & n2149 ;
  assign n16253 = n16252 ^ n2826 ^ 1'b0 ;
  assign n16254 = ( n2625 & ~n3293 ) | ( n2625 & n16253 ) | ( ~n3293 & n16253 ) ;
  assign n16255 = n4562 ^ n2289 ^ 1'b0 ;
  assign n16256 = n16254 | n16255 ;
  assign n16257 = n16256 ^ n11648 ^ n2216 ;
  assign n16259 = ( n1349 & ~n3887 ) | ( n1349 & n12181 ) | ( ~n3887 & n12181 ) ;
  assign n16258 = n3602 | n11303 ;
  assign n16260 = n16259 ^ n16258 ^ 1'b0 ;
  assign n16261 = n12452 ^ n1441 ^ n356 ;
  assign n16262 = n16261 ^ n13650 ^ n8448 ;
  assign n16264 = ( n3164 & ~n11519 ) | ( n3164 & n11876 ) | ( ~n11519 & n11876 ) ;
  assign n16263 = ~n7275 & n11651 ;
  assign n16265 = n16264 ^ n16263 ^ 1'b0 ;
  assign n16266 = n6578 ^ n3055 ^ 1'b0 ;
  assign n16267 = n16265 & ~n16266 ;
  assign n16268 = n5034 ^ n1879 ^ 1'b0 ;
  assign n16269 = n8409 ^ n3614 ^ n1332 ;
  assign n16270 = n16269 ^ n5702 ^ n4066 ;
  assign n16271 = n6256 ^ n3934 ^ 1'b0 ;
  assign n16272 = ~n16270 & n16271 ;
  assign n16273 = n13898 & ~n16272 ;
  assign n16274 = n16273 ^ n14682 ^ n2137 ;
  assign n16275 = ( ~n10176 & n16268 ) | ( ~n10176 & n16274 ) | ( n16268 & n16274 ) ;
  assign n16276 = n7383 & n12924 ;
  assign n16277 = n5057 & ~n16276 ;
  assign n16278 = n16277 ^ n2671 ^ 1'b0 ;
  assign n16279 = ~n7043 & n15129 ;
  assign n16280 = ~n12429 & n16279 ;
  assign n16281 = n4448 & n9869 ;
  assign n16282 = n4088 | n16281 ;
  assign n16283 = n16280 & ~n16282 ;
  assign n16284 = n10901 ^ n6319 ^ n3123 ;
  assign n16285 = n7053 ^ n4385 ^ n3422 ;
  assign n16286 = ~n12634 & n16285 ;
  assign n16287 = n16284 & n16286 ;
  assign n16288 = n16287 ^ n13267 ^ 1'b0 ;
  assign n16289 = n4334 | n8354 ;
  assign n16290 = n16288 & ~n16289 ;
  assign n16291 = n7358 ^ n2058 ^ x115 ;
  assign n16292 = ~n740 & n16291 ;
  assign n16293 = ~n10046 & n16292 ;
  assign n16294 = n4505 ^ n1816 ^ 1'b0 ;
  assign n16295 = ~n2667 & n16294 ;
  assign n16296 = ( n3834 & n4370 ) | ( n3834 & ~n16295 ) | ( n4370 & ~n16295 ) ;
  assign n16297 = n16296 ^ n7187 ^ n1259 ;
  assign n16298 = ( n432 & n16293 ) | ( n432 & ~n16297 ) | ( n16293 & ~n16297 ) ;
  assign n16299 = ( n6293 & ~n9597 ) | ( n6293 & n16298 ) | ( ~n9597 & n16298 ) ;
  assign n16300 = n6974 ^ n5810 ^ 1'b0 ;
  assign n16301 = ( n3135 & n8320 ) | ( n3135 & ~n16300 ) | ( n8320 & ~n16300 ) ;
  assign n16302 = n5859 & n16301 ;
  assign n16303 = n3490 & n14261 ;
  assign n16305 = n13050 ^ n10704 ^ n6391 ;
  assign n16304 = n2289 | n3458 ;
  assign n16306 = n16305 ^ n16304 ^ 1'b0 ;
  assign n16307 = ( n518 & n2860 ) | ( n518 & ~n9542 ) | ( n2860 & ~n9542 ) ;
  assign n16308 = n13219 ^ n2338 ^ 1'b0 ;
  assign n16309 = n4281 & n16308 ;
  assign n16310 = n9487 ^ n1821 ^ 1'b0 ;
  assign n16311 = ~n12972 & n16310 ;
  assign n16312 = ( n1390 & ~n1957 ) | ( n1390 & n4127 ) | ( ~n1957 & n4127 ) ;
  assign n16313 = n16312 ^ n14765 ^ 1'b0 ;
  assign n16314 = n12852 & n16313 ;
  assign n16315 = ( n512 & n3519 ) | ( n512 & ~n16314 ) | ( n3519 & ~n16314 ) ;
  assign n16316 = ( n1904 & n4434 ) | ( n1904 & ~n16177 ) | ( n4434 & ~n16177 ) ;
  assign n16317 = ( n4500 & n5951 ) | ( n4500 & ~n16316 ) | ( n5951 & ~n16316 ) ;
  assign n16318 = n16317 ^ n15117 ^ 1'b0 ;
  assign n16320 = n6654 ^ n3779 ^ 1'b0 ;
  assign n16321 = n4510 & n16320 ;
  assign n16319 = ( n705 & ~n945 ) | ( n705 & n2867 ) | ( ~n945 & n2867 ) ;
  assign n16322 = n16321 ^ n16319 ^ 1'b0 ;
  assign n16323 = n8462 ^ n7584 ^ n6954 ;
  assign n16324 = n13112 ^ n7108 ^ 1'b0 ;
  assign n16325 = n8230 & ~n16324 ;
  assign n16326 = ( n1197 & ~n13752 ) | ( n1197 & n16325 ) | ( ~n13752 & n16325 ) ;
  assign n16329 = n10940 ^ n7909 ^ 1'b0 ;
  assign n16330 = ~n9138 & n16329 ;
  assign n16331 = ~n6093 & n16330 ;
  assign n16332 = n8780 & n16331 ;
  assign n16333 = ( n7068 & n15088 ) | ( n7068 & ~n16332 ) | ( n15088 & ~n16332 ) ;
  assign n16327 = n1872 & n15047 ;
  assign n16328 = n16327 ^ n12307 ^ 1'b0 ;
  assign n16334 = n16333 ^ n16328 ^ n5436 ;
  assign n16335 = n9801 & ~n13045 ;
  assign n16336 = ~n8904 & n16335 ;
  assign n16337 = n13627 & ~n16336 ;
  assign n16338 = ( n1747 & n3125 ) | ( n1747 & ~n6588 ) | ( n3125 & ~n6588 ) ;
  assign n16339 = ( ~n1118 & n10704 ) | ( ~n1118 & n16338 ) | ( n10704 & n16338 ) ;
  assign n16340 = n906 | n4041 ;
  assign n16341 = n16340 ^ n6383 ^ 1'b0 ;
  assign n16342 = n8971 ^ n3013 ^ n589 ;
  assign n16343 = ( n11115 & n16341 ) | ( n11115 & ~n16342 ) | ( n16341 & ~n16342 ) ;
  assign n16344 = n7414 ^ n6566 ^ n4913 ;
  assign n16345 = ( ~n6752 & n16066 ) | ( ~n6752 & n16344 ) | ( n16066 & n16344 ) ;
  assign n16346 = n13727 ^ n7604 ^ 1'b0 ;
  assign n16347 = ~n2284 & n16346 ;
  assign n16348 = n16347 ^ n12360 ^ n7589 ;
  assign n16349 = n9688 ^ n8511 ^ 1'b0 ;
  assign n16350 = n16349 ^ n11009 ^ n6330 ;
  assign n16351 = n6544 ^ n2295 ^ 1'b0 ;
  assign n16352 = n16350 & n16351 ;
  assign n16353 = n10386 ^ n9395 ^ 1'b0 ;
  assign n16354 = ( n8586 & n12000 ) | ( n8586 & ~n14596 ) | ( n12000 & ~n14596 ) ;
  assign n16355 = n16354 ^ n7604 ^ 1'b0 ;
  assign n16356 = ~n12700 & n16355 ;
  assign n16357 = n3008 & ~n9341 ;
  assign n16358 = ( ~n2492 & n3889 ) | ( ~n2492 & n4416 ) | ( n3889 & n4416 ) ;
  assign n16359 = n4409 & n16358 ;
  assign n16360 = n16359 ^ n15473 ^ 1'b0 ;
  assign n16361 = n16360 ^ n12104 ^ n3473 ;
  assign n16366 = ( n10889 & ~n11961 ) | ( n10889 & n14301 ) | ( ~n11961 & n14301 ) ;
  assign n16362 = ~n10386 & n11020 ;
  assign n16363 = ( n1226 & ~n4634 ) | ( n1226 & n16362 ) | ( ~n4634 & n16362 ) ;
  assign n16364 = ~n8032 & n10688 ;
  assign n16365 = n16363 | n16364 ;
  assign n16367 = n16366 ^ n16365 ^ 1'b0 ;
  assign n16368 = ( n7300 & n8275 ) | ( n7300 & ~n12202 ) | ( n8275 & ~n12202 ) ;
  assign n16369 = n16368 ^ n4559 ^ n1590 ;
  assign n16370 = n16369 ^ n4869 ^ 1'b0 ;
  assign n16371 = ( n15442 & n15887 ) | ( n15442 & ~n16370 ) | ( n15887 & ~n16370 ) ;
  assign n16372 = ~n12283 & n16371 ;
  assign n16373 = n9712 & n16372 ;
  assign n16374 = ( n1539 & ~n7598 ) | ( n1539 & n15532 ) | ( ~n7598 & n15532 ) ;
  assign n16375 = n11496 ^ n10054 ^ 1'b0 ;
  assign n16376 = n5059 ^ n4527 ^ 1'b0 ;
  assign n16377 = n16375 & n16376 ;
  assign n16378 = n579 | n6796 ;
  assign n16379 = n16378 ^ n2204 ^ 1'b0 ;
  assign n16380 = ~n6663 & n16379 ;
  assign n16381 = ( n499 & ~n1411 ) | ( n499 & n1714 ) | ( ~n1411 & n1714 ) ;
  assign n16382 = n16381 ^ n12009 ^ n4467 ;
  assign n16383 = n16382 ^ n15589 ^ 1'b0 ;
  assign n16384 = n11287 ^ n7978 ^ 1'b0 ;
  assign n16385 = n4101 ^ n2521 ^ 1'b0 ;
  assign n16386 = n1472 | n16385 ;
  assign n16387 = ( ~n2122 & n2847 ) | ( ~n2122 & n16386 ) | ( n2847 & n16386 ) ;
  assign n16388 = n16387 ^ n381 ^ 1'b0 ;
  assign n16389 = n2055 | n16388 ;
  assign n16390 = n16389 ^ n14966 ^ n6103 ;
  assign n16391 = n16390 ^ n15565 ^ n3787 ;
  assign n16392 = n182 & ~n1450 ;
  assign n16393 = ~n13914 & n16392 ;
  assign n16394 = n16393 ^ n9533 ^ n5582 ;
  assign n16395 = ( n7436 & ~n11429 ) | ( n7436 & n16394 ) | ( ~n11429 & n16394 ) ;
  assign n16396 = n8391 ^ n7133 ^ n2718 ;
  assign n16397 = ( n2428 & n7632 ) | ( n2428 & ~n16396 ) | ( n7632 & ~n16396 ) ;
  assign n16398 = n725 | n8523 ;
  assign n16399 = n16397 | n16398 ;
  assign n16400 = ( n4411 & n4769 ) | ( n4411 & n6425 ) | ( n4769 & n6425 ) ;
  assign n16401 = n10970 | n16400 ;
  assign n16402 = n5015 ^ n760 ^ 1'b0 ;
  assign n16403 = n4724 & ~n5549 ;
  assign n16404 = n16402 & n16403 ;
  assign n16405 = n16404 ^ n8305 ^ n3049 ;
  assign n16406 = n490 | n5585 ;
  assign n16407 = n16406 ^ n3135 ^ n2647 ;
  assign n16408 = n286 | n468 ;
  assign n16409 = n16408 ^ n3285 ^ 1'b0 ;
  assign n16410 = ( n657 & n7090 ) | ( n657 & n8482 ) | ( n7090 & n8482 ) ;
  assign n16411 = ( ~n11003 & n16409 ) | ( ~n11003 & n16410 ) | ( n16409 & n16410 ) ;
  assign n16412 = n16411 ^ n13591 ^ 1'b0 ;
  assign n16413 = n16412 ^ n14255 ^ 1'b0 ;
  assign n16414 = ~n16407 & n16413 ;
  assign n16415 = ( n1063 & ~n1802 ) | ( n1063 & n1992 ) | ( ~n1802 & n1992 ) ;
  assign n16416 = n12873 ^ n4506 ^ 1'b0 ;
  assign n16417 = n16394 & n16416 ;
  assign n16418 = n16417 ^ n8245 ^ n1886 ;
  assign n16419 = n6130 & n16418 ;
  assign n16420 = ~n16415 & n16419 ;
  assign n16421 = n6035 | n12033 ;
  assign n16422 = ( n7135 & n16027 ) | ( n7135 & n16421 ) | ( n16027 & n16421 ) ;
  assign n16423 = n16422 ^ n5705 ^ 1'b0 ;
  assign n16424 = ( n1170 & n2254 ) | ( n1170 & ~n15911 ) | ( n2254 & ~n15911 ) ;
  assign n16425 = ( n8814 & n9630 ) | ( n8814 & ~n13820 ) | ( n9630 & ~n13820 ) ;
  assign n16426 = n6793 & n15653 ;
  assign n16427 = n2808 | n7654 ;
  assign n16428 = n11063 ^ n5939 ^ n1204 ;
  assign n16429 = n6439 & ~n16428 ;
  assign n16430 = n7037 & ~n9468 ;
  assign n16431 = n16430 ^ n6856 ^ 1'b0 ;
  assign n16432 = n3099 & ~n11123 ;
  assign n16433 = n14826 & n16432 ;
  assign n16441 = n8697 | n8967 ;
  assign n16442 = n16441 ^ n2089 ^ 1'b0 ;
  assign n16443 = n7759 | n16442 ;
  assign n16444 = n13146 ^ n9154 ^ 1'b0 ;
  assign n16445 = ~n16443 & n16444 ;
  assign n16440 = ~n4906 & n8516 ;
  assign n16434 = ( x70 & n1519 ) | ( x70 & ~n1572 ) | ( n1519 & ~n1572 ) ;
  assign n16435 = n15604 & n16434 ;
  assign n16436 = n3294 & n16435 ;
  assign n16437 = n16436 ^ n8715 ^ n2557 ;
  assign n16438 = n16437 ^ n2210 ^ 1'b0 ;
  assign n16439 = n6492 & n16438 ;
  assign n16446 = n16445 ^ n16440 ^ n16439 ;
  assign n16448 = n14697 ^ n6522 ^ n1582 ;
  assign n16449 = ~n6190 & n6424 ;
  assign n16450 = n2527 & n16449 ;
  assign n16451 = n16448 & n16450 ;
  assign n16452 = ( ~n3111 & n3330 ) | ( ~n3111 & n16451 ) | ( n3330 & n16451 ) ;
  assign n16447 = ( ~n1472 & n7270 ) | ( ~n1472 & n14055 ) | ( n7270 & n14055 ) ;
  assign n16453 = n16452 ^ n16447 ^ n14045 ;
  assign n16454 = n12259 ^ n6584 ^ n4345 ;
  assign n16455 = ~n16143 & n16454 ;
  assign n16456 = ( n5726 & n14963 ) | ( n5726 & ~n15444 ) | ( n14963 & ~n15444 ) ;
  assign n16460 = n4528 ^ n2520 ^ n1917 ;
  assign n16457 = ( n1287 & n5395 ) | ( n1287 & ~n6978 ) | ( n5395 & ~n6978 ) ;
  assign n16458 = ~n2520 & n16457 ;
  assign n16459 = n16458 ^ n6801 ^ 1'b0 ;
  assign n16461 = n16460 ^ n16459 ^ n7511 ;
  assign n16462 = n9155 ^ n520 ^ 1'b0 ;
  assign n16463 = n1583 & ~n16462 ;
  assign n16464 = n2120 & n16463 ;
  assign n16465 = n16464 ^ n10052 ^ 1'b0 ;
  assign n16466 = ( n485 & n10064 ) | ( n485 & ~n16465 ) | ( n10064 & ~n16465 ) ;
  assign n16467 = n11096 ^ n6259 ^ 1'b0 ;
  assign n16468 = n7320 | n16467 ;
  assign n16469 = n4934 & n13774 ;
  assign n16470 = n3054 | n11687 ;
  assign n16471 = n16470 ^ n15330 ^ 1'b0 ;
  assign n16472 = n3320 | n16471 ;
  assign n16473 = n1804 & ~n4759 ;
  assign n16474 = n5679 & n7132 ;
  assign n16475 = n3263 ^ n653 ^ 1'b0 ;
  assign n16476 = n1143 & n5559 ;
  assign n16477 = n8427 ^ n7083 ^ 1'b0 ;
  assign n16478 = n11130 & ~n16477 ;
  assign n16479 = n16478 ^ n15191 ^ 1'b0 ;
  assign n16480 = n16479 ^ n9147 ^ 1'b0 ;
  assign n16481 = n15574 ^ n13584 ^ n11746 ;
  assign n16482 = ~n7366 & n16481 ;
  assign n16483 = n16482 ^ n10486 ^ n6358 ;
  assign n16484 = n16483 ^ n9509 ^ n3146 ;
  assign n16485 = n10217 ^ n7256 ^ n2620 ;
  assign n16486 = ( n4524 & n6906 ) | ( n4524 & n9516 ) | ( n6906 & n9516 ) ;
  assign n16487 = n15944 ^ n10288 ^ 1'b0 ;
  assign n16488 = n16486 | n16487 ;
  assign n16489 = n16488 ^ n5070 ^ 1'b0 ;
  assign n16490 = n2544 | n11457 ;
  assign n16491 = n7412 & ~n16490 ;
  assign n16492 = n5826 ^ n545 ^ 1'b0 ;
  assign n16493 = n4326 & ~n16492 ;
  assign n16494 = ~n2509 & n3743 ;
  assign n16495 = ( ~n1459 & n6877 ) | ( ~n1459 & n7745 ) | ( n6877 & n7745 ) ;
  assign n16496 = x5 & ~n3823 ;
  assign n16497 = n16496 ^ n1987 ^ 1'b0 ;
  assign n16498 = ( ~n16494 & n16495 ) | ( ~n16494 & n16497 ) | ( n16495 & n16497 ) ;
  assign n16499 = ( n3654 & n16493 ) | ( n3654 & ~n16498 ) | ( n16493 & ~n16498 ) ;
  assign n16501 = n4639 ^ n4416 ^ 1'b0 ;
  assign n16502 = x73 & ~n16501 ;
  assign n16500 = n4801 ^ n4510 ^ 1'b0 ;
  assign n16503 = n16502 ^ n16500 ^ n7060 ;
  assign n16504 = n9109 ^ n7328 ^ n537 ;
  assign n16505 = n4455 | n12180 ;
  assign n16506 = n16505 ^ n15733 ^ 1'b0 ;
  assign n16507 = ( n1012 & n16504 ) | ( n1012 & ~n16506 ) | ( n16504 & ~n16506 ) ;
  assign n16508 = ( n4084 & n13535 ) | ( n4084 & ~n16507 ) | ( n13535 & ~n16507 ) ;
  assign n16509 = n7916 ^ n6855 ^ n5915 ;
  assign n16510 = n16509 ^ n12011 ^ 1'b0 ;
  assign n16511 = n9835 ^ n7693 ^ 1'b0 ;
  assign n16512 = ~n7064 & n16511 ;
  assign n16519 = n4568 ^ n2671 ^ x85 ;
  assign n16520 = ( n310 & n663 ) | ( n310 & n10256 ) | ( n663 & n10256 ) ;
  assign n16521 = ( n11713 & ~n16519 ) | ( n11713 & n16520 ) | ( ~n16519 & n16520 ) ;
  assign n16513 = n14627 ^ n562 ^ 1'b0 ;
  assign n16514 = n10784 & n16513 ;
  assign n16515 = n863 ^ n663 ^ 1'b0 ;
  assign n16516 = n16515 ^ n161 ^ 1'b0 ;
  assign n16517 = n16514 & n16516 ;
  assign n16518 = n11701 & n16517 ;
  assign n16522 = n16521 ^ n16518 ^ n5073 ;
  assign n16530 = ( n1354 & ~n2132 ) | ( n1354 & n11936 ) | ( ~n2132 & n11936 ) ;
  assign n16528 = n3119 ^ n2402 ^ n1594 ;
  assign n16526 = n4295 | n4989 ;
  assign n16527 = n2985 & ~n16526 ;
  assign n16529 = n16528 ^ n16527 ^ 1'b0 ;
  assign n16523 = n3094 | n9414 ;
  assign n16524 = n4414 & ~n16523 ;
  assign n16525 = n16524 ^ n8038 ^ 1'b0 ;
  assign n16531 = n16530 ^ n16529 ^ n16525 ;
  assign n16532 = ( n1199 & n4587 ) | ( n1199 & n5869 ) | ( n4587 & n5869 ) ;
  assign n16533 = n8283 & n15703 ;
  assign n16534 = ~n4771 & n16533 ;
  assign n16535 = ~n9189 & n13640 ;
  assign n16536 = ( x47 & ~n16534 ) | ( x47 & n16535 ) | ( ~n16534 & n16535 ) ;
  assign n16537 = n2211 ^ n1887 ^ 1'b0 ;
  assign n16538 = n11955 | n16537 ;
  assign n16539 = n16536 | n16538 ;
  assign n16540 = ( ~n8201 & n14271 ) | ( ~n8201 & n14433 ) | ( n14271 & n14433 ) ;
  assign n16541 = n1663 & n16540 ;
  assign n16542 = n16541 ^ n7076 ^ n5781 ;
  assign n16543 = ( n243 & n7275 ) | ( n243 & ~n8653 ) | ( n7275 & ~n8653 ) ;
  assign n16545 = n7262 & n9607 ;
  assign n16546 = ( ~n1732 & n4338 ) | ( ~n1732 & n12356 ) | ( n4338 & n12356 ) ;
  assign n16547 = n16546 ^ n2539 ^ 1'b0 ;
  assign n16548 = ( ~n16462 & n16545 ) | ( ~n16462 & n16547 ) | ( n16545 & n16547 ) ;
  assign n16544 = n6215 | n12897 ;
  assign n16549 = n16548 ^ n16544 ^ 1'b0 ;
  assign n16551 = n12722 ^ n1514 ^ 1'b0 ;
  assign n16552 = ( n6887 & n8904 ) | ( n6887 & ~n16551 ) | ( n8904 & ~n16551 ) ;
  assign n16550 = n3119 | n5900 ;
  assign n16553 = n16552 ^ n16550 ^ 1'b0 ;
  assign n16554 = n7096 ^ n4182 ^ 1'b0 ;
  assign n16555 = n14859 & n16554 ;
  assign n16556 = ( n5314 & n10830 ) | ( n5314 & n16555 ) | ( n10830 & n16555 ) ;
  assign n16557 = n13036 ^ n8658 ^ n4744 ;
  assign n16558 = n10081 & ~n16557 ;
  assign n16561 = n10444 ^ n10132 ^ n5334 ;
  assign n16559 = n2292 & ~n8705 ;
  assign n16560 = n16559 ^ n2769 ^ 1'b0 ;
  assign n16562 = n16561 ^ n16560 ^ n10627 ;
  assign n16563 = n6438 ^ n4659 ^ n236 ;
  assign n16564 = ( ~n6433 & n8686 ) | ( ~n6433 & n16563 ) | ( n8686 & n16563 ) ;
  assign n16565 = ( n2194 & ~n3973 ) | ( n2194 & n8104 ) | ( ~n3973 & n8104 ) ;
  assign n16566 = n10704 ^ n9866 ^ n1815 ;
  assign n16567 = ( n10515 & n16565 ) | ( n10515 & ~n16566 ) | ( n16565 & ~n16566 ) ;
  assign n16568 = n12229 ^ n4522 ^ n757 ;
  assign n16569 = n9141 & n13420 ;
  assign n16570 = n6448 ^ n3009 ^ 1'b0 ;
  assign n16571 = n16570 ^ n15911 ^ 1'b0 ;
  assign n16572 = n858 & n16571 ;
  assign n16573 = n16149 ^ n1809 ^ 1'b0 ;
  assign n16574 = n4691 ^ n4249 ^ n2141 ;
  assign n16575 = n16574 ^ n12225 ^ n5572 ;
  assign n16576 = n11673 ^ n9532 ^ n1626 ;
  assign n16577 = n10982 ^ n10959 ^ n10842 ;
  assign n16578 = ( ~n15635 & n16576 ) | ( ~n15635 & n16577 ) | ( n16576 & n16577 ) ;
  assign n16579 = n7454 ^ n6270 ^ 1'b0 ;
  assign n16580 = ~n1004 & n1708 ;
  assign n16581 = n16579 & n16580 ;
  assign n16582 = ( n465 & n13595 ) | ( n465 & n16581 ) | ( n13595 & n16581 ) ;
  assign n16583 = n12123 | n14269 ;
  assign n16585 = n537 & ~n4923 ;
  assign n16584 = n832 & ~n15272 ;
  assign n16586 = n16585 ^ n16584 ^ 1'b0 ;
  assign n16587 = n16586 ^ n8389 ^ 1'b0 ;
  assign n16588 = n13567 | n16587 ;
  assign n16589 = ~n1132 & n1639 ;
  assign n16590 = ~n2415 & n16589 ;
  assign n16591 = n8148 | n16590 ;
  assign n16592 = n9049 | n16591 ;
  assign n16593 = ( n1257 & n6198 ) | ( n1257 & n10772 ) | ( n6198 & n10772 ) ;
  assign n16594 = n1126 & n6274 ;
  assign n16595 = n16594 ^ n14377 ^ n8316 ;
  assign n16596 = n16595 ^ n9958 ^ 1'b0 ;
  assign n16597 = ( ~n1719 & n9452 ) | ( ~n1719 & n15580 ) | ( n9452 & n15580 ) ;
  assign n16598 = n16597 ^ n15174 ^ 1'b0 ;
  assign n16599 = ( n6744 & ~n9563 ) | ( n6744 & n16598 ) | ( ~n9563 & n16598 ) ;
  assign n16600 = n10443 ^ n4770 ^ n1379 ;
  assign n16603 = ~n13749 & n15653 ;
  assign n16602 = n2680 | n15699 ;
  assign n16601 = ~n874 & n4353 ;
  assign n16604 = n16603 ^ n16602 ^ n16601 ;
  assign n16605 = ~n611 & n13736 ;
  assign n16606 = ~n3998 & n5917 ;
  assign n16607 = ~n16605 & n16606 ;
  assign n16608 = ~n15211 & n16607 ;
  assign n16609 = ~n10853 & n16608 ;
  assign n16610 = n12173 ^ n12018 ^ n4262 ;
  assign n16611 = ( n177 & ~n15679 ) | ( n177 & n16610 ) | ( ~n15679 & n16610 ) ;
  assign n16612 = n4961 & n8904 ;
  assign n16613 = ~n12987 & n16612 ;
  assign n16614 = n16613 ^ n12626 ^ n2713 ;
  assign n16615 = n16614 ^ n2176 ^ 1'b0 ;
  assign n16616 = ( n2113 & n5261 ) | ( n2113 & ~n9685 ) | ( n5261 & ~n9685 ) ;
  assign n16617 = n12875 ^ n8252 ^ n162 ;
  assign n16619 = n5548 ^ n4311 ^ 1'b0 ;
  assign n16618 = ~n1508 & n1586 ;
  assign n16620 = n16619 ^ n16618 ^ 1'b0 ;
  assign n16621 = n7512 ^ n5977 ^ 1'b0 ;
  assign n16625 = n3142 & ~n7502 ;
  assign n16626 = ~n6455 & n16625 ;
  assign n16627 = n16626 ^ n7575 ^ n2416 ;
  assign n16628 = ( n2085 & ~n3934 ) | ( n2085 & n16627 ) | ( ~n3934 & n16627 ) ;
  assign n16622 = n4608 ^ n3752 ^ 1'b0 ;
  assign n16623 = n597 & ~n6500 ;
  assign n16624 = n16622 & n16623 ;
  assign n16629 = n16628 ^ n16624 ^ n1805 ;
  assign n16630 = n12015 ^ n3740 ^ n239 ;
  assign n16631 = n760 & n7638 ;
  assign n16632 = n16631 ^ n909 ^ 1'b0 ;
  assign n16633 = n15952 ^ n14779 ^ 1'b0 ;
  assign n16634 = ~n8723 & n16633 ;
  assign n16635 = ~n6840 & n13809 ;
  assign n16636 = ~n12602 & n16635 ;
  assign n16637 = n12239 ^ n10636 ^ 1'b0 ;
  assign n16638 = ~n16636 & n16637 ;
  assign n16639 = n16638 ^ n15655 ^ n13345 ;
  assign n16640 = n8877 ^ n5212 ^ n1782 ;
  assign n16641 = n13095 | n16210 ;
  assign n16642 = n15585 ^ n13635 ^ n3476 ;
  assign n16643 = n4065 ^ n2710 ^ n1250 ;
  assign n16644 = n4403 | n11736 ;
  assign n16645 = n16644 ^ n3436 ^ 1'b0 ;
  assign n16646 = n16643 | n16645 ;
  assign n16647 = ( ~n1109 & n16642 ) | ( ~n1109 & n16646 ) | ( n16642 & n16646 ) ;
  assign n16651 = ( ~n1927 & n5655 ) | ( ~n1927 & n8121 ) | ( n5655 & n8121 ) ;
  assign n16652 = ( n823 & n4742 ) | ( n823 & ~n16651 ) | ( n4742 & ~n16651 ) ;
  assign n16653 = n16652 ^ n4093 ^ 1'b0 ;
  assign n16648 = n4344 ^ n3774 ^ n1554 ;
  assign n16649 = n12563 ^ n7001 ^ 1'b0 ;
  assign n16650 = n16648 | n16649 ;
  assign n16654 = n16653 ^ n16650 ^ n7181 ;
  assign n16655 = n2957 & n4072 ;
  assign n16656 = ~n8655 & n16655 ;
  assign n16657 = ~n1475 & n16656 ;
  assign n16658 = n688 & n5014 ;
  assign n16659 = ~n11725 & n16658 ;
  assign n16660 = ( n6742 & n9850 ) | ( n6742 & n16659 ) | ( n9850 & n16659 ) ;
  assign n16661 = ( n4946 & n12973 ) | ( n4946 & n16660 ) | ( n12973 & n16660 ) ;
  assign n16662 = n10090 ^ n7262 ^ n2267 ;
  assign n16663 = n16662 ^ n9710 ^ n8390 ;
  assign n16664 = ( n3674 & n5680 ) | ( n3674 & n5853 ) | ( n5680 & n5853 ) ;
  assign n16665 = ~n1441 & n11075 ;
  assign n16666 = ~n11838 & n16665 ;
  assign n16667 = n6939 ^ n5167 ^ 1'b0 ;
  assign n16668 = n1722 & ~n6919 ;
  assign n16669 = n16667 & n16668 ;
  assign n16670 = n9249 | n16669 ;
  assign n16671 = n7730 | n11819 ;
  assign n16672 = n16671 ^ n13816 ^ 1'b0 ;
  assign n16673 = n16672 ^ n16069 ^ 1'b0 ;
  assign n16674 = n12293 ^ n7876 ^ 1'b0 ;
  assign n16675 = n12337 & ~n16674 ;
  assign n16676 = ~n4726 & n16675 ;
  assign n16681 = ( ~n2698 & n2870 ) | ( ~n2698 & n6091 ) | ( n2870 & n6091 ) ;
  assign n16682 = n6662 ^ n3078 ^ 1'b0 ;
  assign n16683 = n1243 | n16682 ;
  assign n16684 = n16681 | n16683 ;
  assign n16685 = n11000 | n16684 ;
  assign n16679 = n12339 ^ n12293 ^ n8958 ;
  assign n16677 = ( n2549 & n8290 ) | ( n2549 & n10348 ) | ( n8290 & n10348 ) ;
  assign n16678 = ( n5539 & n6897 ) | ( n5539 & n16677 ) | ( n6897 & n16677 ) ;
  assign n16680 = n16679 ^ n16678 ^ n4486 ;
  assign n16686 = n16685 ^ n16680 ^ n3281 ;
  assign n16687 = ( ~n6281 & n16676 ) | ( ~n6281 & n16686 ) | ( n16676 & n16686 ) ;
  assign n16688 = n16687 ^ n14381 ^ 1'b0 ;
  assign n16689 = ( n3485 & n6344 ) | ( n3485 & ~n8300 ) | ( n6344 & ~n8300 ) ;
  assign n16690 = n7549 | n8699 ;
  assign n16691 = n4451 | n16690 ;
  assign n16692 = ( ~n6881 & n16689 ) | ( ~n6881 & n16691 ) | ( n16689 & n16691 ) ;
  assign n16693 = n3392 | n15898 ;
  assign n16696 = n11696 ^ n9842 ^ x41 ;
  assign n16694 = n3316 | n12863 ;
  assign n16695 = n8566 & ~n16694 ;
  assign n16697 = n16696 ^ n16695 ^ 1'b0 ;
  assign n16698 = n6113 & ~n7837 ;
  assign n16699 = n1811 & n16698 ;
  assign n16700 = n16699 ^ n15963 ^ 1'b0 ;
  assign n16701 = n16697 & n16700 ;
  assign n16702 = n10066 & n11557 ;
  assign n16708 = n8889 ^ n2512 ^ n393 ;
  assign n16706 = ( ~n3848 & n12058 ) | ( ~n3848 & n15272 ) | ( n12058 & n15272 ) ;
  assign n16705 = n4721 & n10278 ;
  assign n16707 = n16706 ^ n16705 ^ n3597 ;
  assign n16703 = ( n905 & n4729 ) | ( n905 & ~n9366 ) | ( n4729 & ~n9366 ) ;
  assign n16704 = ( ~n1976 & n12021 ) | ( ~n1976 & n16703 ) | ( n12021 & n16703 ) ;
  assign n16709 = n16708 ^ n16707 ^ n16704 ;
  assign n16710 = ( ~n8996 & n15886 ) | ( ~n8996 & n16709 ) | ( n15886 & n16709 ) ;
  assign n16711 = n15112 ^ n3898 ^ 1'b0 ;
  assign n16718 = ( n1597 & n2663 ) | ( n1597 & n6359 ) | ( n2663 & n6359 ) ;
  assign n16712 = n4920 ^ n3146 ^ n1239 ;
  assign n16713 = ( n909 & n4531 ) | ( n909 & n8725 ) | ( n4531 & n8725 ) ;
  assign n16714 = n16713 ^ n3289 ^ n1261 ;
  assign n16715 = n9876 ^ n4479 ^ 1'b0 ;
  assign n16716 = ( n16712 & n16714 ) | ( n16712 & ~n16715 ) | ( n16714 & ~n16715 ) ;
  assign n16717 = n16716 ^ n4841 ^ 1'b0 ;
  assign n16719 = n16718 ^ n16717 ^ n2860 ;
  assign n16720 = n3780 & ~n4991 ;
  assign n16721 = n16720 ^ n8348 ^ 1'b0 ;
  assign n16722 = ~n503 & n11783 ;
  assign n16723 = n16722 ^ n7217 ^ 1'b0 ;
  assign n16724 = ~n4118 & n8366 ;
  assign n16725 = ( n5905 & n9801 ) | ( n5905 & ~n16724 ) | ( n9801 & ~n16724 ) ;
  assign n16726 = ( ~n16721 & n16723 ) | ( ~n16721 & n16725 ) | ( n16723 & n16725 ) ;
  assign n16727 = n13315 ^ n9836 ^ n4391 ;
  assign n16728 = n14059 ^ n4816 ^ 1'b0 ;
  assign n16729 = x49 & ~n16728 ;
  assign n16730 = n15894 | n16729 ;
  assign n16732 = n12212 ^ n6475 ^ 1'b0 ;
  assign n16733 = n5103 | n16732 ;
  assign n16734 = n16733 ^ n3995 ^ n3014 ;
  assign n16731 = n5132 | n13687 ;
  assign n16735 = n16734 ^ n16731 ^ 1'b0 ;
  assign n16736 = n6060 | n13025 ;
  assign n16737 = n16736 ^ n9495 ^ 1'b0 ;
  assign n16738 = ~n4098 & n4843 ;
  assign n16739 = n16738 ^ x95 ^ 1'b0 ;
  assign n16740 = n13009 ^ n7300 ^ 1'b0 ;
  assign n16741 = n16740 ^ n12634 ^ 1'b0 ;
  assign n16742 = ( ~x59 & n242 ) | ( ~x59 & n591 ) | ( n242 & n591 ) ;
  assign n16743 = n1475 & ~n16742 ;
  assign n16744 = n11034 ^ n4210 ^ n2021 ;
  assign n16745 = n16743 & ~n16744 ;
  assign n16746 = ( x84 & n4904 ) | ( x84 & n5770 ) | ( n4904 & n5770 ) ;
  assign n16747 = n16746 ^ n8603 ^ n3837 ;
  assign n16748 = n14988 ^ n3486 ^ 1'b0 ;
  assign n16749 = n16748 ^ n13881 ^ n8109 ;
  assign n16750 = ( n925 & n2745 ) | ( n925 & ~n15873 ) | ( n2745 & ~n15873 ) ;
  assign n16751 = ( n5368 & n11988 ) | ( n5368 & ~n16750 ) | ( n11988 & ~n16750 ) ;
  assign n16752 = n10063 & n16751 ;
  assign n16753 = n16752 ^ n8422 ^ n7305 ;
  assign n16760 = n1636 ^ n410 ^ n197 ;
  assign n16757 = n9692 | n16011 ;
  assign n16758 = n16757 ^ n4821 ^ 1'b0 ;
  assign n16754 = ( n3374 & n5907 ) | ( n3374 & n12028 ) | ( n5907 & n12028 ) ;
  assign n16755 = n1292 & n16754 ;
  assign n16756 = n5233 & n16755 ;
  assign n16759 = n16758 ^ n16756 ^ n12201 ;
  assign n16761 = n16760 ^ n16759 ^ x2 ;
  assign n16767 = n2073 | n3988 ;
  assign n16768 = n6067 & ~n16767 ;
  assign n16769 = n3877 & ~n15254 ;
  assign n16770 = ( n2909 & ~n16768 ) | ( n2909 & n16769 ) | ( ~n16768 & n16769 ) ;
  assign n16762 = ( n1844 & ~n4530 ) | ( n1844 & n6895 ) | ( ~n4530 & n6895 ) ;
  assign n16763 = n9186 ^ n7147 ^ 1'b0 ;
  assign n16764 = n16762 & n16763 ;
  assign n16765 = n16764 ^ n14344 ^ n9259 ;
  assign n16766 = ( n8812 & ~n9661 ) | ( n8812 & n16765 ) | ( ~n9661 & n16765 ) ;
  assign n16771 = n16770 ^ n16766 ^ n12700 ;
  assign n16772 = n10725 ^ n5824 ^ 1'b0 ;
  assign n16773 = ( ~n3167 & n5236 ) | ( ~n3167 & n5977 ) | ( n5236 & n5977 ) ;
  assign n16774 = ( n7366 & n16772 ) | ( n7366 & n16773 ) | ( n16772 & n16773 ) ;
  assign n16775 = n9495 | n16774 ;
  assign n16776 = ( n7888 & n8553 ) | ( n7888 & ~n9889 ) | ( n8553 & ~n9889 ) ;
  assign n16777 = n3799 & n16776 ;
  assign n16778 = n16777 ^ n14883 ^ n7252 ;
  assign n16779 = n1777 & n9832 ;
  assign n16780 = n16779 ^ n2153 ^ 1'b0 ;
  assign n16781 = ( ~n4224 & n7840 ) | ( ~n4224 & n14930 ) | ( n7840 & n14930 ) ;
  assign n16782 = n16781 ^ n4957 ^ n2472 ;
  assign n16783 = n3088 & ~n8898 ;
  assign n16784 = n16783 ^ n10108 ^ n9937 ;
  assign n16785 = n5796 ^ n2803 ^ n1318 ;
  assign n16788 = ~n1430 & n13228 ;
  assign n16786 = ~n740 & n5981 ;
  assign n16787 = n16786 ^ n8923 ^ 1'b0 ;
  assign n16789 = n16788 ^ n16787 ^ n11984 ;
  assign n16797 = ( n2733 & ~n5877 ) | ( n2733 & n11112 ) | ( ~n5877 & n11112 ) ;
  assign n16796 = n16717 ^ n12718 ^ n422 ;
  assign n16798 = n16797 ^ n16796 ^ n3466 ;
  assign n16792 = n3880 & n8781 ;
  assign n16793 = ~n7800 & n16792 ;
  assign n16794 = n16793 ^ n16411 ^ n15705 ;
  assign n16795 = n8964 | n16794 ;
  assign n16799 = n16798 ^ n16795 ^ 1'b0 ;
  assign n16790 = ( n2517 & n9758 ) | ( n2517 & n11898 ) | ( n9758 & n11898 ) ;
  assign n16791 = ~n10972 & n16790 ;
  assign n16800 = n16799 ^ n16791 ^ 1'b0 ;
  assign n16801 = n10313 & n11538 ;
  assign n16802 = n13704 ^ n5786 ^ 1'b0 ;
  assign n16803 = n10416 ^ n5125 ^ n1791 ;
  assign n16804 = n16803 ^ n12777 ^ 1'b0 ;
  assign n16805 = ~n6018 & n16804 ;
  assign n16806 = ( n16801 & n16802 ) | ( n16801 & n16805 ) | ( n16802 & n16805 ) ;
  assign n16807 = n142 & n1217 ;
  assign n16808 = n1860 ^ n1511 ^ 1'b0 ;
  assign n16809 = n16808 ^ n7818 ^ 1'b0 ;
  assign n16810 = ( n8577 & n16807 ) | ( n8577 & ~n16809 ) | ( n16807 & ~n16809 ) ;
  assign n16811 = n5530 ^ n4418 ^ 1'b0 ;
  assign n16812 = n16811 ^ n12204 ^ n7684 ;
  assign n16813 = ( n3028 & n3405 ) | ( n3028 & n7668 ) | ( n3405 & n7668 ) ;
  assign n16814 = ~n10264 & n16813 ;
  assign n16815 = n15496 ^ n11913 ^ 1'b0 ;
  assign n16816 = n15983 | n16815 ;
  assign n16817 = n12229 ^ n6330 ^ n351 ;
  assign n16818 = n16817 ^ n14868 ^ 1'b0 ;
  assign n16819 = n1206 & n16209 ;
  assign n16820 = n16819 ^ n5694 ^ 1'b0 ;
  assign n16821 = n9204 & ~n16820 ;
  assign n16822 = n16821 ^ n3227 ^ 1'b0 ;
  assign n16823 = ( ~n4740 & n7030 ) | ( ~n4740 & n16822 ) | ( n7030 & n16822 ) ;
  assign n16824 = n13219 ^ n11201 ^ n3735 ;
  assign n16825 = n16824 ^ n3640 ^ 1'b0 ;
  assign n16826 = ~n499 & n16825 ;
  assign n16827 = n12826 & n16826 ;
  assign n16828 = n6609 | n12674 ;
  assign n16829 = n16828 ^ n9669 ^ 1'b0 ;
  assign n16830 = n14221 ^ n2931 ^ n590 ;
  assign n16831 = n10749 ^ n1631 ^ 1'b0 ;
  assign n16832 = n1778 & ~n16831 ;
  assign n16833 = n16832 ^ n6458 ^ n4149 ;
  assign n16834 = n8734 ^ n316 ^ 1'b0 ;
  assign n16835 = ~n6409 & n13890 ;
  assign n16836 = ( n4370 & n10304 ) | ( n4370 & n16835 ) | ( n10304 & n16835 ) ;
  assign n16837 = n10874 ^ n8403 ^ n3457 ;
  assign n16838 = n16837 ^ n11401 ^ 1'b0 ;
  assign n16839 = n13102 | n16838 ;
  assign n16840 = n11591 ^ n3390 ^ 1'b0 ;
  assign n16841 = n410 & ~n1205 ;
  assign n16842 = n16841 ^ n145 ^ 1'b0 ;
  assign n16843 = n9911 ^ n7745 ^ n401 ;
  assign n16844 = ( ~n12355 & n15972 ) | ( ~n12355 & n16843 ) | ( n15972 & n16843 ) ;
  assign n16845 = ~n8453 & n11159 ;
  assign n16846 = n12181 ^ n3886 ^ n989 ;
  assign n16847 = n2199 | n16846 ;
  assign n16848 = n305 & ~n16847 ;
  assign n16849 = n16848 ^ n11530 ^ n5881 ;
  assign n16850 = ( ~n1388 & n5911 ) | ( ~n1388 & n15404 ) | ( n5911 & n15404 ) ;
  assign n16851 = ~n4941 & n16850 ;
  assign n16852 = n15388 | n16851 ;
  assign n16856 = ( ~n492 & n1409 ) | ( ~n492 & n3169 ) | ( n1409 & n3169 ) ;
  assign n16853 = n5252 ^ n4521 ^ 1'b0 ;
  assign n16854 = x63 & n16853 ;
  assign n16855 = ~n8473 & n16854 ;
  assign n16857 = n16856 ^ n16855 ^ 1'b0 ;
  assign n16858 = n16857 ^ n11426 ^ 1'b0 ;
  assign n16859 = ( n4146 & n4630 ) | ( n4146 & ~n7793 ) | ( n4630 & ~n7793 ) ;
  assign n16860 = ( ~n2922 & n7838 ) | ( ~n2922 & n16859 ) | ( n7838 & n16859 ) ;
  assign n16861 = n14199 ^ n5946 ^ n1203 ;
  assign n16862 = n10094 | n14602 ;
  assign n16863 = n16862 ^ n6401 ^ 1'b0 ;
  assign n16864 = n1821 ^ n563 ^ x113 ;
  assign n16865 = ~n4884 & n16864 ;
  assign n16866 = n16863 & n16865 ;
  assign n16867 = n3343 | n10497 ;
  assign n16868 = n1772 | n16867 ;
  assign n16869 = n950 | n16868 ;
  assign n16870 = n15198 ^ n5250 ^ n1199 ;
  assign n16871 = n5534 | n8097 ;
  assign n16872 = n5102 ^ n1655 ^ 1'b0 ;
  assign n16873 = ~n11994 & n16872 ;
  assign n16874 = n16873 ^ n14249 ^ 1'b0 ;
  assign n16875 = n16874 ^ n15991 ^ n14343 ;
  assign n16883 = n10826 ^ n2122 ^ n692 ;
  assign n16876 = n15556 ^ n8519 ^ n5696 ;
  assign n16877 = ( n5039 & ~n6104 ) | ( n5039 & n6471 ) | ( ~n6104 & n6471 ) ;
  assign n16878 = n16877 ^ n3157 ^ n1817 ;
  assign n16879 = n10406 | n16410 ;
  assign n16880 = n2105 | n16879 ;
  assign n16881 = ( ~n16876 & n16878 ) | ( ~n16876 & n16880 ) | ( n16878 & n16880 ) ;
  assign n16882 = n1183 | n16881 ;
  assign n16884 = n16883 ^ n16882 ^ n6169 ;
  assign n16885 = ( n2027 & ~n2931 ) | ( n2027 & n2974 ) | ( ~n2931 & n2974 ) ;
  assign n16886 = ( n2862 & n12224 ) | ( n2862 & n16885 ) | ( n12224 & n16885 ) ;
  assign n16887 = n10663 & ~n16014 ;
  assign n16888 = n3579 & n16887 ;
  assign n16889 = n1466 & ~n6009 ;
  assign n16890 = n540 & n16889 ;
  assign n16891 = ( n678 & ~n3787 ) | ( n678 & n10031 ) | ( ~n3787 & n10031 ) ;
  assign n16892 = n14633 ^ n4497 ^ n4432 ;
  assign n16893 = ~n12308 & n16892 ;
  assign n16894 = n16893 ^ n6571 ^ 1'b0 ;
  assign n16895 = ( n16890 & n16891 ) | ( n16890 & ~n16894 ) | ( n16891 & ~n16894 ) ;
  assign n16896 = n12203 | n12706 ;
  assign n16897 = n16896 ^ n3467 ^ 1'b0 ;
  assign n16898 = n780 & ~n16897 ;
  assign n16899 = ( n5529 & n5827 ) | ( n5529 & ~n16898 ) | ( n5827 & ~n16898 ) ;
  assign n16900 = n2126 & n5474 ;
  assign n16901 = n2249 & n16900 ;
  assign n16902 = ( n4960 & n14251 ) | ( n4960 & n16901 ) | ( n14251 & n16901 ) ;
  assign n16903 = n3871 & n13776 ;
  assign n16904 = n2380 & n16903 ;
  assign n16905 = ( ~n1485 & n8472 ) | ( ~n1485 & n16904 ) | ( n8472 & n16904 ) ;
  assign n16906 = n16905 ^ n15685 ^ n5467 ;
  assign n16907 = n3709 ^ n1602 ^ 1'b0 ;
  assign n16909 = n7496 ^ n7128 ^ n1107 ;
  assign n16908 = n10065 | n15380 ;
  assign n16910 = n16909 ^ n16908 ^ 1'b0 ;
  assign n16913 = ~n2983 & n3928 ;
  assign n16914 = ~n2254 & n16913 ;
  assign n16911 = ~n4318 & n4934 ;
  assign n16912 = ~n975 & n16911 ;
  assign n16915 = n16914 ^ n16912 ^ n1750 ;
  assign n16916 = n8535 & n16915 ;
  assign n16917 = n6701 & n16916 ;
  assign n16918 = n7065 ^ x81 ^ 1'b0 ;
  assign n16919 = ( ~n1111 & n1136 ) | ( ~n1111 & n2283 ) | ( n1136 & n2283 ) ;
  assign n16920 = n11859 & ~n16919 ;
  assign n16921 = n1645 | n4867 ;
  assign n16924 = n14032 ^ n4259 ^ n3210 ;
  assign n16922 = n1018 | n13155 ;
  assign n16923 = n13809 | n16922 ;
  assign n16925 = n16924 ^ n16923 ^ 1'b0 ;
  assign n16926 = n6380 ^ n1270 ^ 1'b0 ;
  assign n16927 = ~n14418 & n16926 ;
  assign n16928 = ~n272 & n16927 ;
  assign n16929 = x84 | n16928 ;
  assign n16930 = n2954 | n4654 ;
  assign n16931 = n8497 | n16930 ;
  assign n16932 = ( n3377 & n11402 ) | ( n3377 & ~n16931 ) | ( n11402 & ~n16931 ) ;
  assign n16933 = n16932 ^ n6534 ^ 1'b0 ;
  assign n16934 = n16929 & ~n16933 ;
  assign n16935 = n7630 ^ n6123 ^ 1'b0 ;
  assign n16936 = n7847 | n16935 ;
  assign n16937 = n4875 ^ n4684 ^ 1'b0 ;
  assign n16938 = n533 | n16937 ;
  assign n16939 = n5362 ^ n367 ^ 1'b0 ;
  assign n16940 = ~n8870 & n16939 ;
  assign n16941 = ( ~n2772 & n3294 ) | ( ~n2772 & n11932 ) | ( n3294 & n11932 ) ;
  assign n16942 = ( n4286 & n15963 ) | ( n4286 & ~n16941 ) | ( n15963 & ~n16941 ) ;
  assign n16943 = ~n11624 & n16942 ;
  assign n16944 = n16943 ^ n7897 ^ 1'b0 ;
  assign n16945 = ( n16938 & n16940 ) | ( n16938 & n16944 ) | ( n16940 & n16944 ) ;
  assign n16946 = ( n129 & n1320 ) | ( n129 & ~n4326 ) | ( n1320 & ~n4326 ) ;
  assign n16947 = n16946 ^ n2353 ^ 1'b0 ;
  assign n16948 = n3917 & ~n16947 ;
  assign n16949 = n215 & ~n15330 ;
  assign n16950 = n16949 ^ n2643 ^ 1'b0 ;
  assign n16951 = n16950 ^ n12296 ^ 1'b0 ;
  assign n16952 = ~n3028 & n16951 ;
  assign n16953 = n16952 ^ n12027 ^ n8804 ;
  assign n16954 = n4843 & ~n8335 ;
  assign n16955 = n16954 ^ n4110 ^ 1'b0 ;
  assign n16956 = ~n3212 & n8959 ;
  assign n16957 = n16956 ^ n9828 ^ 1'b0 ;
  assign n16958 = n11060 ^ n10659 ^ 1'b0 ;
  assign n16959 = ~n7059 & n16958 ;
  assign n16960 = ~n16957 & n16959 ;
  assign n16961 = n16960 ^ n13038 ^ n1815 ;
  assign n16962 = n16955 & n16961 ;
  assign n16963 = ~n2830 & n16962 ;
  assign n16964 = n11818 ^ n2717 ^ n2475 ;
  assign n16965 = n664 | n6320 ;
  assign n16966 = n16412 ^ n12553 ^ 1'b0 ;
  assign n16967 = n407 & n16966 ;
  assign n16968 = n14783 ^ n13244 ^ 1'b0 ;
  assign n16969 = ~n5534 & n16968 ;
  assign n16970 = n14057 ^ n7239 ^ 1'b0 ;
  assign n16971 = n16970 ^ n11166 ^ 1'b0 ;
  assign n16972 = n16971 ^ n8406 ^ n1732 ;
  assign n16973 = n7435 ^ n1136 ^ 1'b0 ;
  assign n16974 = ~n3800 & n16973 ;
  assign n16975 = ( n748 & n4249 ) | ( n748 & ~n16974 ) | ( n4249 & ~n16974 ) ;
  assign n16979 = n3507 ^ n1310 ^ n681 ;
  assign n16976 = ( n1530 & ~n4127 ) | ( n1530 & n5854 ) | ( ~n4127 & n5854 ) ;
  assign n16977 = ( ~n4934 & n8084 ) | ( ~n4934 & n16976 ) | ( n8084 & n16976 ) ;
  assign n16978 = n16977 ^ n8978 ^ n7660 ;
  assign n16980 = n16979 ^ n16978 ^ 1'b0 ;
  assign n16981 = ~n9189 & n16980 ;
  assign n16982 = n11986 ^ n7934 ^ 1'b0 ;
  assign n16983 = ~n5987 & n16982 ;
  assign n16984 = n16983 ^ n9803 ^ n4489 ;
  assign n16985 = n13671 & ~n16984 ;
  assign n16986 = ~n5510 & n16985 ;
  assign n16987 = n1500 & ~n4089 ;
  assign n16988 = n16987 ^ n9296 ^ 1'b0 ;
  assign n16989 = ( n570 & n9379 ) | ( n570 & n16988 ) | ( n9379 & n16988 ) ;
  assign n16990 = ~n4331 & n5731 ;
  assign n16991 = n16990 ^ n13600 ^ n9661 ;
  assign n16992 = n4685 ^ n1719 ^ n131 ;
  assign n16993 = n3773 & ~n6574 ;
  assign n16994 = n589 & n16993 ;
  assign n16995 = ( n10141 & n16992 ) | ( n10141 & n16994 ) | ( n16992 & n16994 ) ;
  assign n16996 = ( n5133 & ~n12425 ) | ( n5133 & n16995 ) | ( ~n12425 & n16995 ) ;
  assign n16997 = n16091 ^ n6742 ^ n6221 ;
  assign n16998 = n16997 ^ n7798 ^ 1'b0 ;
  assign n16999 = ~n16996 & n16998 ;
  assign n17000 = ~n5920 & n9123 ;
  assign n17001 = n17000 ^ n13169 ^ 1'b0 ;
  assign n17002 = n4229 | n17001 ;
  assign n17003 = ( n6563 & n16999 ) | ( n6563 & n17002 ) | ( n16999 & n17002 ) ;
  assign n17004 = n5227 ^ n2906 ^ 1'b0 ;
  assign n17005 = n581 & n17004 ;
  assign n17006 = n17005 ^ n9221 ^ n4849 ;
  assign n17007 = n2176 & n13768 ;
  assign n17008 = n17006 & n17007 ;
  assign n17009 = n13249 ^ n9607 ^ x30 ;
  assign n17010 = n8349 ^ n523 ^ 1'b0 ;
  assign n17011 = n8408 | n17010 ;
  assign n17012 = n17009 | n17011 ;
  assign n17013 = n12049 & ~n17012 ;
  assign n17014 = n1722 & ~n4839 ;
  assign n17015 = ~n5438 & n17014 ;
  assign n17016 = ( ~n9772 & n16957 ) | ( ~n9772 & n17015 ) | ( n16957 & n17015 ) ;
  assign n17017 = n17016 ^ n11835 ^ n4858 ;
  assign n17018 = n5416 | n10301 ;
  assign n17019 = n14247 | n17018 ;
  assign n17020 = n17019 ^ n13667 ^ 1'b0 ;
  assign n17021 = ~n8752 & n14562 ;
  assign n17022 = ~n527 & n3030 ;
  assign n17023 = ~n1486 & n16506 ;
  assign n17024 = n10234 & n17023 ;
  assign n17025 = ( n3850 & n17022 ) | ( n3850 & ~n17024 ) | ( n17022 & ~n17024 ) ;
  assign n17026 = n17025 ^ n8765 ^ 1'b0 ;
  assign n17027 = n6555 ^ n5432 ^ n1823 ;
  assign n17028 = n17027 ^ n3734 ^ n3567 ;
  assign n17029 = n7755 | n17028 ;
  assign n17030 = n2878 | n16689 ;
  assign n17031 = n17030 ^ n4651 ^ 1'b0 ;
  assign n17032 = n13505 | n13830 ;
  assign n17033 = n2890 | n17032 ;
  assign n17034 = n15792 ^ n14345 ^ n13516 ;
  assign n17035 = n6850 ^ n4889 ^ n2708 ;
  assign n17036 = n9021 & n17035 ;
  assign n17037 = n8138 ^ n1349 ^ x78 ;
  assign n17038 = ( n8189 & n16546 ) | ( n8189 & n17037 ) | ( n16546 & n17037 ) ;
  assign n17039 = n1902 | n10422 ;
  assign n17040 = ( n3680 & ~n9501 ) | ( n3680 & n17039 ) | ( ~n9501 & n17039 ) ;
  assign n17041 = n4421 ^ n1597 ^ 1'b0 ;
  assign n17042 = n15276 | n17041 ;
  assign n17043 = n15722 ^ n4378 ^ n1672 ;
  assign n17044 = ~n209 & n2921 ;
  assign n17046 = ( n726 & ~n5545 ) | ( n726 & n6009 ) | ( ~n5545 & n6009 ) ;
  assign n17045 = n12292 ^ n2076 ^ 1'b0 ;
  assign n17047 = n17046 ^ n17045 ^ n12214 ;
  assign n17048 = n4011 & ~n5653 ;
  assign n17049 = n6934 & n17048 ;
  assign n17050 = n17049 ^ n16317 ^ n1368 ;
  assign n17051 = n10227 & ~n10754 ;
  assign n17052 = n17051 ^ n10280 ^ 1'b0 ;
  assign n17053 = n4061 ^ n2325 ^ 1'b0 ;
  assign n17054 = n5093 & ~n17053 ;
  assign n17055 = n17052 & n17054 ;
  assign n17056 = n9805 ^ n686 ^ 1'b0 ;
  assign n17057 = n5957 | n7899 ;
  assign n17058 = n1761 | n17057 ;
  assign n17059 = n9632 ^ n4913 ^ n1160 ;
  assign n17060 = ( ~n1791 & n13398 ) | ( ~n1791 & n13920 ) | ( n13398 & n13920 ) ;
  assign n17061 = n16797 & n17060 ;
  assign n17062 = n17059 & n17061 ;
  assign n17063 = n5187 ^ n2809 ^ 1'b0 ;
  assign n17064 = n17063 ^ n14173 ^ n767 ;
  assign n17065 = ~n2548 & n7585 ;
  assign n17066 = n17065 ^ n2358 ^ 1'b0 ;
  assign n17067 = ( n7627 & n11596 ) | ( n7627 & n13925 ) | ( n11596 & n13925 ) ;
  assign n17068 = n1872 & n17067 ;
  assign n17069 = n17066 & n17068 ;
  assign n17070 = n17069 ^ n8978 ^ 1'b0 ;
  assign n17071 = n13336 & n17070 ;
  assign n17072 = ( n7434 & n17064 ) | ( n7434 & n17071 ) | ( n17064 & n17071 ) ;
  assign n17073 = ~n437 & n12404 ;
  assign n17075 = ( n2111 & n3311 ) | ( n2111 & ~n7060 ) | ( n3311 & ~n7060 ) ;
  assign n17076 = n17075 ^ n3633 ^ n1541 ;
  assign n17077 = ~n660 & n5853 ;
  assign n17078 = n17077 ^ n6668 ^ 1'b0 ;
  assign n17079 = ( ~n3573 & n17076 ) | ( ~n3573 & n17078 ) | ( n17076 & n17078 ) ;
  assign n17074 = n1343 & n14186 ;
  assign n17080 = n17079 ^ n17074 ^ 1'b0 ;
  assign n17081 = n8311 & ~n17080 ;
  assign n17082 = n17081 ^ n7323 ^ 1'b0 ;
  assign n17083 = n10817 ^ n9843 ^ n1650 ;
  assign n17085 = n7399 ^ n291 ^ 1'b0 ;
  assign n17086 = n2952 | n17085 ;
  assign n17084 = n8103 & ~n8883 ;
  assign n17087 = n17086 ^ n17084 ^ 1'b0 ;
  assign n17088 = ( n17082 & n17083 ) | ( n17082 & ~n17087 ) | ( n17083 & ~n17087 ) ;
  assign n17089 = n7160 & ~n7774 ;
  assign n17090 = ~n10076 & n17089 ;
  assign n17091 = n17090 ^ n15462 ^ 1'b0 ;
  assign n17092 = ~n4168 & n15244 ;
  assign n17093 = n2584 & n17092 ;
  assign n17094 = n17093 ^ n5767 ^ n3892 ;
  assign n17095 = n11720 ^ n2578 ^ n1313 ;
  assign n17096 = ( n11382 & ~n17094 ) | ( n11382 & n17095 ) | ( ~n17094 & n17095 ) ;
  assign n17099 = n5134 & n7401 ;
  assign n17097 = n1663 & n10386 ;
  assign n17098 = ~n9010 & n17097 ;
  assign n17100 = n17099 ^ n17098 ^ n7992 ;
  assign n17101 = n6768 ^ n2293 ^ 1'b0 ;
  assign n17102 = n7664 & ~n7977 ;
  assign n17103 = n17102 ^ n7684 ^ 1'b0 ;
  assign n17104 = n3975 ^ n3610 ^ 1'b0 ;
  assign n17105 = ~n17103 & n17104 ;
  assign n17106 = n7207 ^ n6356 ^ 1'b0 ;
  assign n17107 = n17106 ^ n10416 ^ n7299 ;
  assign n17108 = ( n3691 & n10203 ) | ( n3691 & ~n17107 ) | ( n10203 & ~n17107 ) ;
  assign n17109 = n17108 ^ n12856 ^ n10494 ;
  assign n17112 = n4217 & ~n6215 ;
  assign n17113 = n13563 & n17112 ;
  assign n17110 = n6881 ^ n6822 ^ n1709 ;
  assign n17111 = n17110 ^ n8915 ^ n5140 ;
  assign n17114 = n17113 ^ n17111 ^ n10700 ;
  assign n17115 = ( n394 & ~n632 ) | ( n394 & n801 ) | ( ~n632 & n801 ) ;
  assign n17116 = ( n10401 & n11158 ) | ( n10401 & ~n17115 ) | ( n11158 & ~n17115 ) ;
  assign n17117 = ~n6004 & n12337 ;
  assign n17118 = ~n10286 & n17117 ;
  assign n17119 = n11793 & n17118 ;
  assign n17120 = n15039 ^ n15027 ^ 1'b0 ;
  assign n17121 = n4450 | n4505 ;
  assign n17122 = n17120 | n17121 ;
  assign n17123 = ( n5285 & n10815 ) | ( n5285 & ~n16689 ) | ( n10815 & ~n16689 ) ;
  assign n17124 = n17123 ^ n10060 ^ n6009 ;
  assign n17125 = n17124 ^ n13153 ^ n12242 ;
  assign n17126 = n10278 ^ n4192 ^ n1578 ;
  assign n17127 = ( n4899 & n14587 ) | ( n4899 & n17126 ) | ( n14587 & n17126 ) ;
  assign n17129 = n4252 | n4556 ;
  assign n17130 = n17129 ^ n8583 ^ 1'b0 ;
  assign n17128 = n11522 | n12822 ;
  assign n17131 = n17130 ^ n17128 ^ 1'b0 ;
  assign n17132 = n17131 ^ n10598 ^ n6598 ;
  assign n17136 = ( n447 & n457 ) | ( n447 & n6002 ) | ( n457 & n6002 ) ;
  assign n17137 = n17136 ^ n16001 ^ n11004 ;
  assign n17133 = ( n506 & n2042 ) | ( n506 & n9898 ) | ( n2042 & n9898 ) ;
  assign n17134 = n3247 ^ n912 ^ 1'b0 ;
  assign n17135 = n17133 & n17134 ;
  assign n17138 = n17137 ^ n17135 ^ 1'b0 ;
  assign n17139 = n5955 & n17138 ;
  assign n17140 = n10784 ^ n7777 ^ n2428 ;
  assign n17141 = ( n604 & n6608 ) | ( n604 & ~n7671 ) | ( n6608 & ~n7671 ) ;
  assign n17142 = n6840 & n17141 ;
  assign n17143 = ~n13081 & n17142 ;
  assign n17146 = n9908 ^ n3232 ^ n397 ;
  assign n17147 = n17146 ^ n12932 ^ n2527 ;
  assign n17144 = n4711 ^ n2881 ^ 1'b0 ;
  assign n17145 = n8869 & ~n17144 ;
  assign n17148 = n17147 ^ n17145 ^ n1774 ;
  assign n17149 = n16065 ^ n15657 ^ n8475 ;
  assign n17150 = n17149 ^ n5578 ^ 1'b0 ;
  assign n17151 = n4999 | n17150 ;
  assign n17152 = ( n8017 & n8413 ) | ( n8017 & n15800 ) | ( n8413 & n15800 ) ;
  assign n17153 = ~n2165 & n5981 ;
  assign n17154 = n17153 ^ x72 ^ 1'b0 ;
  assign n17155 = n1053 & n8784 ;
  assign n17156 = n8389 ^ n6826 ^ 1'b0 ;
  assign n17157 = x36 & n17156 ;
  assign n17158 = ( n3749 & n15667 ) | ( n3749 & ~n17157 ) | ( n15667 & ~n17157 ) ;
  assign n17159 = n8083 | n17158 ;
  assign n17160 = n17159 ^ n1986 ^ 1'b0 ;
  assign n17161 = ~n5470 & n13568 ;
  assign n17162 = n17161 ^ n4130 ^ 1'b0 ;
  assign n17163 = n17162 ^ n17054 ^ 1'b0 ;
  assign n17164 = ( ~n11538 & n17160 ) | ( ~n11538 & n17163 ) | ( n17160 & n17163 ) ;
  assign n17165 = n17155 | n17164 ;
  assign n17166 = n17154 & ~n17165 ;
  assign n17167 = ( n13685 & ~n17152 ) | ( n13685 & n17166 ) | ( ~n17152 & n17166 ) ;
  assign n17168 = x15 & n14867 ;
  assign n17169 = n17168 ^ n6112 ^ 1'b0 ;
  assign n17170 = n12977 ^ n7714 ^ 1'b0 ;
  assign n17171 = ( x106 & n506 ) | ( x106 & ~n2406 ) | ( n506 & ~n2406 ) ;
  assign n17172 = n17171 ^ n6750 ^ 1'b0 ;
  assign n17173 = n10608 ^ n8446 ^ n1651 ;
  assign n17174 = n17173 ^ n14545 ^ n12407 ;
  assign n17175 = n17174 ^ n8571 ^ n3091 ;
  assign n17176 = n14330 ^ n4253 ^ 1'b0 ;
  assign n17177 = ( n6240 & n9547 ) | ( n6240 & n10723 ) | ( n9547 & n10723 ) ;
  assign n17178 = n12265 | n17177 ;
  assign n17179 = n5444 & ~n15723 ;
  assign n17180 = n17179 ^ n3823 ^ 1'b0 ;
  assign n17181 = n8234 ^ n7119 ^ n1287 ;
  assign n17182 = n6442 ^ n3098 ^ n2093 ;
  assign n17183 = ( n9982 & n10808 ) | ( n9982 & ~n17182 ) | ( n10808 & ~n17182 ) ;
  assign n17184 = n9524 ^ n8664 ^ 1'b0 ;
  assign n17185 = ~n1210 & n17184 ;
  assign n17186 = ( ~n271 & n17183 ) | ( ~n271 & n17185 ) | ( n17183 & n17185 ) ;
  assign n17187 = ( n6939 & ~n7328 ) | ( n6939 & n9258 ) | ( ~n7328 & n9258 ) ;
  assign n17188 = ( n253 & n7472 ) | ( n253 & n17187 ) | ( n7472 & n17187 ) ;
  assign n17189 = ( n6378 & n15949 ) | ( n6378 & n17188 ) | ( n15949 & n17188 ) ;
  assign n17190 = ~n7758 & n9823 ;
  assign n17191 = ~n17189 & n17190 ;
  assign n17192 = ( n1465 & ~n3517 ) | ( n1465 & n11249 ) | ( ~n3517 & n11249 ) ;
  assign n17193 = n17192 ^ n14987 ^ n11842 ;
  assign n17194 = n4189 & ~n8980 ;
  assign n17195 = n17194 ^ n7628 ^ 1'b0 ;
  assign n17196 = n17195 ^ n9064 ^ 1'b0 ;
  assign n17197 = n8937 ^ n6708 ^ 1'b0 ;
  assign n17198 = ~n3151 & n9860 ;
  assign n17199 = ( ~n13102 & n17197 ) | ( ~n13102 & n17198 ) | ( n17197 & n17198 ) ;
  assign n17200 = ( n6335 & n16773 ) | ( n6335 & ~n17199 ) | ( n16773 & ~n17199 ) ;
  assign n17201 = n9600 ^ n6783 ^ n3144 ;
  assign n17202 = n11263 | n17201 ;
  assign n17203 = n11823 ^ n6506 ^ 1'b0 ;
  assign n17204 = n11996 | n17203 ;
  assign n17205 = n17202 & ~n17204 ;
  assign n17206 = n13425 ^ n9960 ^ 1'b0 ;
  assign n17207 = n17206 ^ n6429 ^ n3499 ;
  assign n17208 = n8786 ^ n6488 ^ 1'b0 ;
  assign n17209 = n4209 ^ n3030 ^ 1'b0 ;
  assign n17210 = n2769 & ~n17209 ;
  assign n17211 = n13423 ^ n7941 ^ n4288 ;
  assign n17213 = n5770 ^ n3880 ^ 1'b0 ;
  assign n17212 = n4094 & ~n11461 ;
  assign n17214 = n17213 ^ n17212 ^ 1'b0 ;
  assign n17215 = n17214 ^ n14762 ^ 1'b0 ;
  assign n17216 = n13888 ^ n11842 ^ n4694 ;
  assign n17217 = n8791 ^ n8707 ^ n1069 ;
  assign n17218 = n11820 & n15744 ;
  assign n17219 = n17217 | n17218 ;
  assign n17220 = ~n1020 & n3126 ;
  assign n17221 = n17220 ^ n11932 ^ 1'b0 ;
  assign n17222 = n11115 & n17221 ;
  assign n17223 = n17222 ^ n3389 ^ 1'b0 ;
  assign n17224 = n3569 | n4572 ;
  assign n17225 = n17224 ^ n7396 ^ 1'b0 ;
  assign n17226 = ( n15545 & ~n17042 ) | ( n15545 & n17225 ) | ( ~n17042 & n17225 ) ;
  assign n17227 = n10964 ^ n7061 ^ n625 ;
  assign n17228 = n15133 ^ n5268 ^ 1'b0 ;
  assign n17229 = n17227 & n17228 ;
  assign n17230 = n8140 ^ n883 ^ 1'b0 ;
  assign n17231 = ( ~n976 & n15562 ) | ( ~n976 & n17230 ) | ( n15562 & n17230 ) ;
  assign n17232 = n12968 ^ n10266 ^ 1'b0 ;
  assign n17233 = ~n8157 & n17232 ;
  assign n17234 = ~n11727 & n17233 ;
  assign n17235 = ~n9970 & n14993 ;
  assign n17236 = n17235 ^ n10214 ^ 1'b0 ;
  assign n17237 = ~n6748 & n7871 ;
  assign n17238 = n7775 & n17237 ;
  assign n17239 = n17238 ^ n8957 ^ 1'b0 ;
  assign n17240 = n1320 & n3408 ;
  assign n17241 = n5222 & n9777 ;
  assign n17242 = n9049 & ~n10401 ;
  assign n17243 = n17242 ^ n7598 ^ 1'b0 ;
  assign n17244 = n17038 ^ n15918 ^ n9123 ;
  assign n17245 = n15823 ^ n1434 ^ 1'b0 ;
  assign n17246 = n17245 ^ n4037 ^ x26 ;
  assign n17247 = n13092 ^ n12885 ^ 1'b0 ;
  assign n17248 = n11622 & n17247 ;
  assign n17249 = n4138 & ~n14959 ;
  assign n17250 = n644 | n4993 ;
  assign n17251 = n17250 ^ n10662 ^ n5255 ;
  assign n17252 = n3129 & ~n17251 ;
  assign n17253 = n17252 ^ n15247 ^ 1'b0 ;
  assign n17254 = ( n12490 & n12590 ) | ( n12490 & n16105 ) | ( n12590 & n16105 ) ;
  assign n17255 = n10068 ^ n4556 ^ 1'b0 ;
  assign n17256 = n8970 | n12396 ;
  assign n17257 = ( ~n6477 & n15043 ) | ( ~n6477 & n17256 ) | ( n15043 & n17256 ) ;
  assign n17258 = n13219 ^ n5369 ^ 1'b0 ;
  assign n17259 = n9078 & n12905 ;
  assign n17260 = n17259 ^ n12008 ^ 1'b0 ;
  assign n17261 = ~n8783 & n17260 ;
  assign n17262 = ~n9232 & n17261 ;
  assign n17263 = n7389 & ~n15454 ;
  assign n17266 = n7518 ^ n4198 ^ n2539 ;
  assign n17267 = n17266 ^ n10066 ^ 1'b0 ;
  assign n17264 = n878 ^ n876 ^ 1'b0 ;
  assign n17265 = n4711 & ~n17264 ;
  assign n17268 = n17267 ^ n17265 ^ n4293 ;
  assign n17269 = n17268 ^ n4758 ^ n2195 ;
  assign n17270 = ( n2620 & n9741 ) | ( n2620 & ~n15029 ) | ( n9741 & ~n15029 ) ;
  assign n17271 = n12659 & n17270 ;
  assign n17272 = n17271 ^ n11471 ^ 1'b0 ;
  assign n17273 = n15372 ^ n8387 ^ 1'b0 ;
  assign n17274 = ~n1445 & n17273 ;
  assign n17275 = ~n6254 & n6574 ;
  assign n17276 = n2546 | n17142 ;
  assign n17277 = ( ~n7155 & n13501 ) | ( ~n7155 & n17276 ) | ( n13501 & n17276 ) ;
  assign n17278 = n6560 & ~n14046 ;
  assign n17279 = n11033 & ~n17278 ;
  assign n17280 = n3203 & n4717 ;
  assign n17281 = n5796 & n17280 ;
  assign n17282 = ( n1672 & n10296 ) | ( n1672 & n17281 ) | ( n10296 & n17281 ) ;
  assign n17283 = n17279 | n17282 ;
  assign n17284 = n894 | n10181 ;
  assign n17285 = n17284 ^ n2042 ^ 1'b0 ;
  assign n17286 = n767 | n16835 ;
  assign n17287 = n17286 ^ n3238 ^ 1'b0 ;
  assign n17288 = n2314 | n3253 ;
  assign n17289 = ( n5137 & ~n12791 ) | ( n5137 & n17288 ) | ( ~n12791 & n17288 ) ;
  assign n17290 = n1999 | n4275 ;
  assign n17291 = n3109 & ~n17290 ;
  assign n17292 = n17291 ^ n7769 ^ n2835 ;
  assign n17293 = n2789 | n17292 ;
  assign n17294 = n11097 & n17293 ;
  assign n17295 = n8781 ^ n4020 ^ 1'b0 ;
  assign n17296 = n6239 ^ n4689 ^ 1'b0 ;
  assign n17297 = n17295 & n17296 ;
  assign n17298 = ~n7695 & n17297 ;
  assign n17299 = n9039 & ~n17298 ;
  assign n17304 = n11683 ^ n7143 ^ 1'b0 ;
  assign n17300 = n8193 ^ n6861 ^ 1'b0 ;
  assign n17301 = n2532 & ~n17300 ;
  assign n17302 = n17301 ^ n13334 ^ n11659 ;
  assign n17303 = n1369 & n17302 ;
  assign n17305 = n17304 ^ n17303 ^ 1'b0 ;
  assign n17306 = n5086 ^ n933 ^ n609 ;
  assign n17307 = n17306 ^ n3480 ^ n750 ;
  assign n17308 = n2857 & n14010 ;
  assign n17309 = n17307 & ~n17308 ;
  assign n17310 = n10090 & n17309 ;
  assign n17311 = ( x69 & n369 ) | ( x69 & n4213 ) | ( n369 & n4213 ) ;
  assign n17312 = n12488 ^ n5029 ^ 1'b0 ;
  assign n17313 = n9117 ^ n8559 ^ n2778 ;
  assign n17314 = n17313 ^ n13232 ^ 1'b0 ;
  assign n17315 = ( n1481 & ~n16389 ) | ( n1481 & n17314 ) | ( ~n16389 & n17314 ) ;
  assign n17316 = ( n6059 & n6903 ) | ( n6059 & n12345 ) | ( n6903 & n12345 ) ;
  assign n17317 = n13723 ^ n11003 ^ 1'b0 ;
  assign n17318 = n3054 | n17317 ;
  assign n17319 = n8781 & ~n16441 ;
  assign n17320 = n3326 ^ n831 ^ 1'b0 ;
  assign n17321 = n5483 ^ n3487 ^ n1612 ;
  assign n17322 = n4838 ^ n3610 ^ n1174 ;
  assign n17323 = n17322 ^ n11842 ^ n7836 ;
  assign n17324 = n17323 ^ n8684 ^ n6437 ;
  assign n17325 = ( ~n6474 & n17321 ) | ( ~n6474 & n17324 ) | ( n17321 & n17324 ) ;
  assign n17326 = ( n6966 & n17320 ) | ( n6966 & ~n17325 ) | ( n17320 & ~n17325 ) ;
  assign n17327 = n6507 | n17326 ;
  assign n17328 = n17319 | n17327 ;
  assign n17329 = n17328 ^ n10634 ^ n254 ;
  assign n17330 = n17318 | n17329 ;
  assign n17331 = n1500 & ~n10494 ;
  assign n17332 = n17331 ^ n7460 ^ 1'b0 ;
  assign n17338 = n14577 ^ n314 ^ 1'b0 ;
  assign n17333 = n10931 & ~n12887 ;
  assign n17334 = ~n1049 & n17333 ;
  assign n17335 = n2292 & n3359 ;
  assign n17336 = n17334 & n17335 ;
  assign n17337 = n5781 | n17336 ;
  assign n17339 = n17338 ^ n17337 ^ 1'b0 ;
  assign n17341 = n4164 ^ n1711 ^ 1'b0 ;
  assign n17342 = n4137 & n17341 ;
  assign n17340 = ~n5655 & n12616 ;
  assign n17343 = n17342 ^ n17340 ^ 1'b0 ;
  assign n17344 = n14753 & ~n17343 ;
  assign n17345 = n5356 ^ n4443 ^ n1315 ;
  assign n17346 = n17345 ^ n10973 ^ n10775 ;
  assign n17347 = n17346 ^ n2569 ^ 1'b0 ;
  assign n17348 = n17344 | n17347 ;
  assign n17349 = n12449 ^ n4546 ^ 1'b0 ;
  assign n17350 = n2989 | n17349 ;
  assign n17351 = n11346 & ~n17350 ;
  assign n17352 = ~n10740 & n17351 ;
  assign n17353 = n6524 | n8791 ;
  assign n17354 = n10922 & ~n17353 ;
  assign n17355 = ( n1323 & n6332 ) | ( n1323 & n17354 ) | ( n6332 & n17354 ) ;
  assign n17356 = ( n2306 & ~n2744 ) | ( n2306 & n17355 ) | ( ~n2744 & n17355 ) ;
  assign n17357 = ( n2743 & ~n3623 ) | ( n2743 & n12577 ) | ( ~n3623 & n12577 ) ;
  assign n17358 = ( n3490 & n3689 ) | ( n3490 & n17357 ) | ( n3689 & n17357 ) ;
  assign n17359 = n2747 | n8923 ;
  assign n17360 = n9801 | n17359 ;
  assign n17361 = ( n7208 & n8313 ) | ( n7208 & ~n16762 ) | ( n8313 & ~n16762 ) ;
  assign n17362 = ~n1655 & n5346 ;
  assign n17363 = n11278 & n15541 ;
  assign n17364 = n17362 & n17363 ;
  assign n17365 = n1703 ^ n785 ^ 1'b0 ;
  assign n17366 = n17365 ^ n4650 ^ 1'b0 ;
  assign n17367 = n2217 | n10059 ;
  assign n17369 = n12977 ^ n672 ^ 1'b0 ;
  assign n17368 = ~n4175 & n9484 ;
  assign n17370 = n17369 ^ n17368 ^ 1'b0 ;
  assign n17371 = ( n168 & n17367 ) | ( n168 & n17370 ) | ( n17367 & n17370 ) ;
  assign n17372 = ( n965 & n3566 ) | ( n965 & n14385 ) | ( n3566 & n14385 ) ;
  assign n17373 = n10012 ^ n6177 ^ 1'b0 ;
  assign n17374 = n5482 & ~n17373 ;
  assign n17375 = n11022 & ~n17374 ;
  assign n17376 = n10183 ^ n6786 ^ 1'b0 ;
  assign n17377 = n6906 & n17376 ;
  assign n17378 = n17377 ^ n323 ^ 1'b0 ;
  assign n17379 = n3410 & n17378 ;
  assign n17380 = n17375 & n17379 ;
  assign n17381 = n10742 ^ n7358 ^ 1'b0 ;
  assign n17382 = n8427 ^ n2343 ^ 1'b0 ;
  assign n17383 = n6699 ^ n2769 ^ n967 ;
  assign n17384 = n2707 ^ n253 ^ 1'b0 ;
  assign n17385 = n17384 ^ n8624 ^ 1'b0 ;
  assign n17386 = ( n17382 & n17383 ) | ( n17382 & n17385 ) | ( n17383 & n17385 ) ;
  assign n17387 = n8831 & n11604 ;
  assign n17388 = n17387 ^ n5889 ^ 1'b0 ;
  assign n17389 = n14358 ^ n13868 ^ n7212 ;
  assign n17390 = n12238 ^ n8059 ^ n2857 ;
  assign n17391 = ( ~n17388 & n17389 ) | ( ~n17388 & n17390 ) | ( n17389 & n17390 ) ;
  assign n17392 = ( n17381 & n17386 ) | ( n17381 & ~n17391 ) | ( n17386 & ~n17391 ) ;
  assign n17393 = n11370 ^ n4919 ^ 1'b0 ;
  assign n17394 = ~n11670 & n17393 ;
  assign n17395 = n3398 & ~n17394 ;
  assign n17396 = ~n1212 & n3596 ;
  assign n17397 = n17396 ^ n14132 ^ 1'b0 ;
  assign n17398 = n10776 & ~n17397 ;
  assign n17399 = n4004 & ~n5219 ;
  assign n17400 = n11860 & n17399 ;
  assign n17401 = n7962 ^ n4202 ^ n1566 ;
  assign n17402 = ( n6927 & ~n7490 ) | ( n6927 & n17401 ) | ( ~n7490 & n17401 ) ;
  assign n17403 = n17402 ^ n8204 ^ n6019 ;
  assign n17404 = ( n3302 & n4322 ) | ( n3302 & n7403 ) | ( n4322 & n7403 ) ;
  assign n17405 = n3930 | n12202 ;
  assign n17406 = n17405 ^ n10274 ^ 1'b0 ;
  assign n17407 = ~n13141 & n17406 ;
  assign n17408 = x38 & n17407 ;
  assign n17409 = ( ~n15762 & n17404 ) | ( ~n15762 & n17408 ) | ( n17404 & n17408 ) ;
  assign n17410 = n16436 ^ n9538 ^ 1'b0 ;
  assign n17411 = n17410 ^ n12711 ^ n7639 ;
  assign n17412 = n17411 ^ n9015 ^ n5405 ;
  assign n17413 = ( n2178 & n6104 ) | ( n2178 & ~n7620 ) | ( n6104 & ~n7620 ) ;
  assign n17414 = n10592 ^ n8980 ^ n8350 ;
  assign n17416 = n5681 & ~n6770 ;
  assign n17415 = n3877 & n5296 ;
  assign n17417 = n17416 ^ n17415 ^ 1'b0 ;
  assign n17418 = n2926 | n7083 ;
  assign n17419 = n17418 ^ n8098 ^ 1'b0 ;
  assign n17420 = n5397 ^ n2111 ^ n1414 ;
  assign n17421 = n7917 ^ n6598 ^ n4087 ;
  assign n17422 = ( n5844 & n16193 ) | ( n5844 & n17421 ) | ( n16193 & n17421 ) ;
  assign n17423 = ~n1830 & n3281 ;
  assign n17424 = ~n1490 & n17423 ;
  assign n17425 = ( ~n2611 & n12612 ) | ( ~n2611 & n17424 ) | ( n12612 & n17424 ) ;
  assign n17426 = ( ~n4878 & n9070 ) | ( ~n4878 & n12061 ) | ( n9070 & n12061 ) ;
  assign n17427 = n17426 ^ n10671 ^ 1'b0 ;
  assign n17428 = ( n2734 & n8718 ) | ( n2734 & ~n9731 ) | ( n8718 & ~n9731 ) ;
  assign n17429 = n14789 ^ n8443 ^ 1'b0 ;
  assign n17430 = ( n720 & n9416 ) | ( n720 & ~n16846 ) | ( n9416 & ~n16846 ) ;
  assign n17431 = n10092 ^ n5539 ^ n2510 ;
  assign n17432 = n9049 ^ n8066 ^ n4793 ;
  assign n17433 = n4990 ^ n2582 ^ 1'b0 ;
  assign n17434 = ( ~n2577 & n17432 ) | ( ~n2577 & n17433 ) | ( n17432 & n17433 ) ;
  assign n17435 = n17431 | n17434 ;
  assign n17436 = n17430 & n17435 ;
  assign n17437 = n17436 ^ n5121 ^ 1'b0 ;
  assign n17438 = n11278 ^ n2697 ^ 1'b0 ;
  assign n17439 = n1050 & ~n17438 ;
  assign n17442 = n10482 ^ n9347 ^ n7962 ;
  assign n17440 = n16091 ^ n9664 ^ n2026 ;
  assign n17441 = n17440 ^ n14627 ^ n1761 ;
  assign n17443 = n17442 ^ n17441 ^ n2211 ;
  assign n17444 = n17443 ^ n12521 ^ n5816 ;
  assign n17445 = n16931 ^ n4465 ^ 1'b0 ;
  assign n17446 = n11185 & n17445 ;
  assign n17447 = n2358 & n16864 ;
  assign n17448 = n1297 & n17447 ;
  assign n17449 = n17448 ^ n2521 ^ 1'b0 ;
  assign n17450 = n8933 & ~n17449 ;
  assign n17451 = n17450 ^ n15217 ^ n9553 ;
  assign n17452 = ( ~n4981 & n8734 ) | ( ~n4981 & n9642 ) | ( n8734 & n9642 ) ;
  assign n17453 = n5942 ^ n1145 ^ 1'b0 ;
  assign n17454 = ~n8673 & n17453 ;
  assign n17455 = n3595 & n3899 ;
  assign n17456 = ~n12669 & n17455 ;
  assign n17457 = n15244 ^ n9808 ^ n5645 ;
  assign n17458 = n12911 ^ n10854 ^ n9570 ;
  assign n17459 = n16769 | n17458 ;
  assign n17460 = n17459 ^ n1001 ^ 1'b0 ;
  assign n17461 = ( ~n4562 & n6588 ) | ( ~n4562 & n9001 ) | ( n6588 & n9001 ) ;
  assign n17462 = n17461 ^ n9355 ^ 1'b0 ;
  assign n17463 = n7286 ^ n6376 ^ 1'b0 ;
  assign n17464 = n12157 & ~n17463 ;
  assign n17465 = ( n629 & n1392 ) | ( n629 & n1803 ) | ( n1392 & n1803 ) ;
  assign n17466 = ( x123 & n3830 ) | ( x123 & ~n17465 ) | ( n3830 & ~n17465 ) ;
  assign n17467 = n9296 | n12098 ;
  assign n17468 = n2882 | n4408 ;
  assign n17469 = n7049 ^ n3269 ^ 1'b0 ;
  assign n17470 = ~n8643 & n10161 ;
  assign n17471 = n3513 & n17470 ;
  assign n17472 = n17471 ^ n2056 ^ 1'b0 ;
  assign n17473 = n14244 ^ n7363 ^ 1'b0 ;
  assign n17474 = n12351 | n17473 ;
  assign n17475 = ~n811 & n2847 ;
  assign n17476 = n17475 ^ n2295 ^ 1'b0 ;
  assign n17477 = n17476 ^ n10749 ^ n872 ;
  assign n17478 = n14554 ^ n3182 ^ n300 ;
  assign n17479 = n3840 & n17478 ;
  assign n17480 = n17477 & n17479 ;
  assign n17481 = ( n137 & n1347 ) | ( n137 & n10762 ) | ( n1347 & n10762 ) ;
  assign n17482 = ~n4016 & n12873 ;
  assign n17483 = n17482 ^ n8014 ^ 1'b0 ;
  assign n17484 = ~n17481 & n17483 ;
  assign n17485 = ~n919 & n17484 ;
  assign n17486 = n5980 ^ n1216 ^ 1'b0 ;
  assign n17487 = n2542 & n17486 ;
  assign n17488 = n17487 ^ n14238 ^ n7337 ;
  assign n17489 = n17488 ^ n12565 ^ n1561 ;
  assign n17490 = n1952 & ~n17489 ;
  assign n17491 = n311 & n17490 ;
  assign n17495 = ( n1972 & n2959 ) | ( n1972 & ~n6354 ) | ( n2959 & ~n6354 ) ;
  assign n17496 = n10311 ^ n7918 ^ n5564 ;
  assign n17497 = ( n3953 & ~n17495 ) | ( n3953 & n17496 ) | ( ~n17495 & n17496 ) ;
  assign n17492 = n4976 & n5083 ;
  assign n17493 = n17492 ^ n5754 ^ 1'b0 ;
  assign n17494 = n3253 & ~n17493 ;
  assign n17498 = n17497 ^ n17494 ^ 1'b0 ;
  assign n17499 = ( n13573 & n17491 ) | ( n13573 & ~n17498 ) | ( n17491 & ~n17498 ) ;
  assign n17500 = n6855 ^ n469 ^ 1'b0 ;
  assign n17501 = n1225 & ~n7598 ;
  assign n17502 = n4638 ^ n2880 ^ 1'b0 ;
  assign n17504 = n11694 ^ n429 ^ 1'b0 ;
  assign n17505 = n11119 | n17504 ;
  assign n17503 = n763 | n10503 ;
  assign n17506 = n17505 ^ n17503 ^ n13868 ;
  assign n17507 = n17506 ^ n11832 ^ n3800 ;
  assign n17508 = ( ~n2527 & n6427 ) | ( ~n2527 & n10825 ) | ( n6427 & n10825 ) ;
  assign n17509 = n1349 & n17508 ;
  assign n17510 = n17509 ^ n11523 ^ 1'b0 ;
  assign n17511 = n8916 ^ n6191 ^ n4344 ;
  assign n17512 = n6420 & n10633 ;
  assign n17513 = n17511 & n17512 ;
  assign n17514 = n17513 ^ n6802 ^ 1'b0 ;
  assign n17515 = n2098 & ~n7632 ;
  assign n17516 = ~n8316 & n17515 ;
  assign n17517 = n11225 & n12449 ;
  assign n17518 = n17517 ^ n14921 ^ n5751 ;
  assign n17519 = ( n5100 & n14947 ) | ( n5100 & n17518 ) | ( n14947 & n17518 ) ;
  assign n17520 = n3082 ^ n1895 ^ 1'b0 ;
  assign n17521 = ( n4181 & n4429 ) | ( n4181 & ~n17520 ) | ( n4429 & ~n17520 ) ;
  assign n17522 = n17354 ^ n16072 ^ n11394 ;
  assign n17523 = n9074 ^ n6319 ^ 1'b0 ;
  assign n17524 = ~n17522 & n17523 ;
  assign n17525 = ( n13221 & n17521 ) | ( n13221 & n17524 ) | ( n17521 & n17524 ) ;
  assign n17526 = n14890 ^ n3476 ^ n1606 ;
  assign n17527 = n14939 ^ n9609 ^ n676 ;
  assign n17528 = ( ~n1174 & n4310 ) | ( ~n1174 & n9828 ) | ( n4310 & n9828 ) ;
  assign n17529 = n17528 ^ n2915 ^ 1'b0 ;
  assign n17530 = ~n3467 & n6618 ;
  assign n17531 = n15477 ^ n4539 ^ n1406 ;
  assign n17532 = n13218 & n17531 ;
  assign n17533 = ~n4268 & n8607 ;
  assign n17535 = n7732 ^ n3779 ^ 1'b0 ;
  assign n17534 = ~n4020 & n6503 ;
  assign n17536 = n17535 ^ n17534 ^ n12446 ;
  assign n17537 = n11073 ^ n1411 ^ 1'b0 ;
  assign n17538 = n17537 ^ n14529 ^ n4129 ;
  assign n17540 = n4339 ^ n4161 ^ 1'b0 ;
  assign n17541 = n17540 ^ n8646 ^ 1'b0 ;
  assign n17539 = ~n1749 & n10273 ;
  assign n17542 = n17541 ^ n17539 ^ n12675 ;
  assign n17543 = n7074 ^ n5177 ^ 1'b0 ;
  assign n17544 = n2027 & n17543 ;
  assign n17545 = n13479 ^ n4846 ^ 1'b0 ;
  assign n17548 = n6033 ^ n1296 ^ n957 ;
  assign n17546 = n6783 ^ n6104 ^ n1338 ;
  assign n17547 = n17546 ^ n15801 ^ n4325 ;
  assign n17549 = n17548 ^ n17547 ^ n3689 ;
  assign n17550 = n6941 ^ n3614 ^ 1'b0 ;
  assign n17551 = n17550 ^ n8408 ^ n2236 ;
  assign n17552 = n17551 ^ n5849 ^ 1'b0 ;
  assign n17553 = n2321 & ~n2728 ;
  assign n17554 = ~n10667 & n17553 ;
  assign n17555 = ( ~n6352 & n10516 ) | ( ~n6352 & n16362 ) | ( n10516 & n16362 ) ;
  assign n17556 = n4486 | n4505 ;
  assign n17557 = n136 & ~n17556 ;
  assign n17558 = n17557 ^ n11596 ^ n3243 ;
  assign n17559 = n10808 | n17558 ;
  assign n17560 = n17559 ^ n13944 ^ n8265 ;
  assign n17561 = ~n5797 & n17560 ;
  assign n17562 = ( n9695 & ~n13061 ) | ( n9695 & n13203 ) | ( ~n13061 & n13203 ) ;
  assign n17563 = n7594 ^ n2643 ^ 1'b0 ;
  assign n17564 = n17563 ^ n5259 ^ 1'b0 ;
  assign n17565 = ( ~n2917 & n8003 ) | ( ~n2917 & n15450 ) | ( n8003 & n15450 ) ;
  assign n17566 = n14251 ^ n4179 ^ 1'b0 ;
  assign n17567 = n11698 & ~n17566 ;
  assign n17568 = n3131 & n6718 ;
  assign n17569 = ( n5216 & n12073 ) | ( n5216 & ~n13314 ) | ( n12073 & ~n13314 ) ;
  assign n17570 = n17569 ^ n7317 ^ n3916 ;
  assign n17573 = ( ~n3125 & n4094 ) | ( ~n3125 & n6815 ) | ( n4094 & n6815 ) ;
  assign n17571 = n6268 & ~n12077 ;
  assign n17572 = ~n16715 & n17571 ;
  assign n17574 = n17573 ^ n17572 ^ 1'b0 ;
  assign n17575 = n17574 ^ n5464 ^ n3071 ;
  assign n17576 = n9219 ^ n3077 ^ 1'b0 ;
  assign n17577 = n17576 ^ n4114 ^ n933 ;
  assign n17578 = n1280 & ~n7135 ;
  assign n17579 = ( n145 & ~n6913 ) | ( n145 & n17578 ) | ( ~n6913 & n17578 ) ;
  assign n17580 = ( n7838 & n17577 ) | ( n7838 & n17579 ) | ( n17577 & n17579 ) ;
  assign n17581 = n17580 ^ n8819 ^ 1'b0 ;
  assign n17582 = n4685 & ~n16030 ;
  assign n17583 = ~n7971 & n17582 ;
  assign n17584 = n17583 ^ n12728 ^ n5438 ;
  assign n17585 = ( n12594 & n17441 ) | ( n12594 & n17584 ) | ( n17441 & n17584 ) ;
  assign n17586 = ( n2107 & ~n4512 ) | ( n2107 & n6824 ) | ( ~n4512 & n6824 ) ;
  assign n17587 = ( ~n817 & n10323 ) | ( ~n817 & n11363 ) | ( n10323 & n11363 ) ;
  assign n17588 = n10152 & n17587 ;
  assign n17589 = n3588 & n13523 ;
  assign n17590 = n17589 ^ n5364 ^ 1'b0 ;
  assign n17591 = ( ~n7884 & n15492 ) | ( ~n7884 & n17590 ) | ( n15492 & n17590 ) ;
  assign n17592 = n5981 & n5990 ;
  assign n17593 = n7510 | n17592 ;
  assign n17594 = n6537 & ~n17593 ;
  assign n17595 = ~n17591 & n17594 ;
  assign n17596 = n4477 & n9157 ;
  assign n17597 = ( n559 & n8180 ) | ( n559 & ~n12024 ) | ( n8180 & ~n12024 ) ;
  assign n17598 = n1119 & n15848 ;
  assign n17599 = n17597 & n17598 ;
  assign n17600 = n17599 ^ n3702 ^ 1'b0 ;
  assign n17601 = ~n17596 & n17600 ;
  assign n17602 = ~n2157 & n4320 ;
  assign n17603 = ~n933 & n17602 ;
  assign n17604 = n8855 & n17603 ;
  assign n17605 = ( n1374 & n8703 ) | ( n1374 & n15511 ) | ( n8703 & n15511 ) ;
  assign n17606 = ( n2072 & n17604 ) | ( n2072 & n17605 ) | ( n17604 & n17605 ) ;
  assign n17607 = n17192 ^ n8577 ^ n903 ;
  assign n17608 = n17607 ^ n10484 ^ n1354 ;
  assign n17609 = n3374 & ~n16296 ;
  assign n17610 = n17609 ^ n9700 ^ 1'b0 ;
  assign n17611 = n5391 ^ n4190 ^ 1'b0 ;
  assign n17612 = n10913 ^ n2025 ^ 1'b0 ;
  assign n17613 = n17611 & n17612 ;
  assign n17614 = ( n4501 & ~n17610 ) | ( n4501 & n17613 ) | ( ~n17610 & n17613 ) ;
  assign n17615 = n7006 ^ n506 ^ 1'b0 ;
  assign n17616 = n17615 ^ n15665 ^ n8957 ;
  assign n17617 = ~x96 & n713 ;
  assign n17618 = n239 & n1018 ;
  assign n17619 = n17618 ^ n10564 ^ 1'b0 ;
  assign n17620 = ~n17617 & n17619 ;
  assign n17621 = n10182 & n17620 ;
  assign n17622 = n17621 ^ n17223 ^ 1'b0 ;
  assign n17623 = n7846 | n8580 ;
  assign n17624 = n13633 ^ n11432 ^ 1'b0 ;
  assign n17625 = n5073 | n11551 ;
  assign n17626 = ~n6579 & n7733 ;
  assign n17627 = n17626 ^ n2670 ^ 1'b0 ;
  assign n17628 = ( ~n9208 & n9897 ) | ( ~n9208 & n17627 ) | ( n9897 & n17627 ) ;
  assign n17629 = ( n9157 & n10566 ) | ( n9157 & ~n17628 ) | ( n10566 & ~n17628 ) ;
  assign n17630 = n10043 | n17629 ;
  assign n17631 = n2787 ^ n1636 ^ x90 ;
  assign n17632 = ( n10668 & n11769 ) | ( n10668 & n17631 ) | ( n11769 & n17631 ) ;
  assign n17633 = ( n978 & n11958 ) | ( n978 & ~n17632 ) | ( n11958 & ~n17632 ) ;
  assign n17636 = n9495 ^ n7478 ^ n5704 ;
  assign n17634 = ~n916 & n2301 ;
  assign n17635 = n17634 ^ n13993 ^ 1'b0 ;
  assign n17637 = n17636 ^ n17635 ^ n12879 ;
  assign n17638 = n3098 & ~n9306 ;
  assign n17639 = n6057 ^ x73 ^ 1'b0 ;
  assign n17640 = n12038 & ~n17639 ;
  assign n17641 = n2857 & ~n17640 ;
  assign n17642 = ( n12443 & n17638 ) | ( n12443 & n17641 ) | ( n17638 & n17641 ) ;
  assign n17643 = ( n2812 & n3462 ) | ( n2812 & n5546 ) | ( n3462 & n5546 ) ;
  assign n17644 = n11995 ^ n1887 ^ 1'b0 ;
  assign n17645 = n17643 & n17644 ;
  assign n17646 = n17645 ^ n5923 ^ 1'b0 ;
  assign n17647 = ( n645 & ~n8529 ) | ( n645 & n9086 ) | ( ~n8529 & n9086 ) ;
  assign n17648 = n11187 & ~n17647 ;
  assign n17649 = n17648 ^ n12327 ^ 1'b0 ;
  assign n17650 = n16627 ^ n13162 ^ 1'b0 ;
  assign n17651 = ~n10759 & n17650 ;
  assign n17652 = x2 & ~n17651 ;
  assign n17656 = n12404 & ~n14437 ;
  assign n17654 = ( n465 & n2565 ) | ( n465 & n11722 ) | ( n2565 & n11722 ) ;
  assign n17653 = ~n4448 & n5860 ;
  assign n17655 = n17654 ^ n17653 ^ 1'b0 ;
  assign n17657 = n17656 ^ n17655 ^ n15113 ;
  assign n17658 = n12101 & ~n17657 ;
  assign n17659 = ~n16316 & n17658 ;
  assign n17660 = n7718 | n17659 ;
  assign n17661 = n2255 & n17120 ;
  assign n17662 = n17661 ^ n13851 ^ 1'b0 ;
  assign n17663 = n17662 ^ n17213 ^ n16397 ;
  assign n17665 = n3363 ^ n3084 ^ 1'b0 ;
  assign n17666 = n4008 & n17665 ;
  assign n17664 = ( ~n2551 & n12286 ) | ( ~n2551 & n16347 ) | ( n12286 & n16347 ) ;
  assign n17667 = n17666 ^ n17664 ^ n6931 ;
  assign n17668 = n566 & ~n17667 ;
  assign n17669 = n763 & n835 ;
  assign n17670 = ~n763 & n17669 ;
  assign n17671 = n2567 | n17670 ;
  assign n17672 = n17670 & ~n17671 ;
  assign n17673 = ( n8475 & n9260 ) | ( n8475 & n17672 ) | ( n9260 & n17672 ) ;
  assign n17674 = ( ~n3126 & n4936 ) | ( ~n3126 & n17673 ) | ( n4936 & n17673 ) ;
  assign n17677 = ( ~n1645 & n11374 ) | ( ~n1645 & n13725 ) | ( n11374 & n13725 ) ;
  assign n17675 = n12897 ^ n4719 ^ 1'b0 ;
  assign n17676 = ( n4981 & ~n11972 ) | ( n4981 & n17675 ) | ( ~n11972 & n17675 ) ;
  assign n17678 = n17677 ^ n17676 ^ 1'b0 ;
  assign n17679 = n17174 | n17678 ;
  assign n17680 = ( n7256 & n7983 ) | ( n7256 & ~n8162 ) | ( n7983 & ~n8162 ) ;
  assign n17681 = n537 & ~n17680 ;
  assign n17682 = n17681 ^ n1816 ^ 1'b0 ;
  assign n17683 = ( n605 & ~n1465 ) | ( n605 & n11534 ) | ( ~n1465 & n11534 ) ;
  assign n17684 = n9310 ^ n5357 ^ n3928 ;
  assign n17686 = n5438 ^ n3766 ^ 1'b0 ;
  assign n17685 = n1815 & n2517 ;
  assign n17687 = n17686 ^ n17685 ^ 1'b0 ;
  assign n17688 = n10421 ^ n4059 ^ 1'b0 ;
  assign n17689 = n17687 | n17688 ;
  assign n17690 = n4366 ^ n2901 ^ 1'b0 ;
  assign n17691 = ( n876 & n7228 ) | ( n876 & ~n16877 ) | ( n7228 & ~n16877 ) ;
  assign n17692 = ( n1987 & n3976 ) | ( n1987 & n9258 ) | ( n3976 & n9258 ) ;
  assign n17693 = n7599 & ~n10769 ;
  assign n17694 = n17692 & n17693 ;
  assign n17695 = n16130 ^ n12859 ^ n7858 ;
  assign n17696 = n11008 ^ n1882 ^ 1'b0 ;
  assign n17697 = n2200 & ~n17696 ;
  assign n17698 = ~n17695 & n17697 ;
  assign n17699 = n513 & ~n2992 ;
  assign n17700 = n11053 & ~n17699 ;
  assign n17701 = n17700 ^ n4690 ^ 1'b0 ;
  assign n17702 = n10481 ^ n808 ^ 1'b0 ;
  assign n17703 = n17702 ^ n7762 ^ 1'b0 ;
  assign n17704 = n17701 & n17703 ;
  assign n17705 = n16203 & n17704 ;
  assign n17706 = n4826 & n17705 ;
  assign n17707 = n8002 ^ n5605 ^ n5065 ;
  assign n17708 = n17707 ^ n2556 ^ 1'b0 ;
  assign n17709 = n7938 & n17708 ;
  assign n17710 = n17709 ^ n3892 ^ n1929 ;
  assign n17711 = ( ~n4073 & n12865 ) | ( ~n4073 & n13164 ) | ( n12865 & n13164 ) ;
  assign n17712 = n1292 | n17711 ;
  assign n17713 = n15880 ^ n7213 ^ 1'b0 ;
  assign n17714 = n17402 ^ n11720 ^ n8543 ;
  assign n17715 = ( n1739 & n2955 ) | ( n1739 & n4879 ) | ( n2955 & n4879 ) ;
  assign n17716 = n17715 ^ n9322 ^ 1'b0 ;
  assign n17717 = n11341 & n17716 ;
  assign n17718 = n17717 ^ n12728 ^ 1'b0 ;
  assign n17719 = n17718 ^ n15216 ^ n7318 ;
  assign n17720 = n17719 ^ n16955 ^ 1'b0 ;
  assign n17721 = n3466 & ~n3548 ;
  assign n17722 = ( n2409 & n2728 ) | ( n2409 & ~n6121 ) | ( n2728 & ~n6121 ) ;
  assign n17723 = n2146 | n17722 ;
  assign n17724 = n17721 | n17723 ;
  assign n17725 = ( ~n1079 & n3466 ) | ( ~n1079 & n8983 ) | ( n3466 & n8983 ) ;
  assign n17726 = ( x52 & n16961 ) | ( x52 & n17725 ) | ( n16961 & n17725 ) ;
  assign n17727 = n15254 ^ n14046 ^ 1'b0 ;
  assign n17728 = n17727 ^ n14799 ^ n7780 ;
  assign n17729 = ( x89 & ~n314 ) | ( x89 & n1860 ) | ( ~n314 & n1860 ) ;
  assign n17730 = ( n1511 & n10085 ) | ( n1511 & n17729 ) | ( n10085 & n17729 ) ;
  assign n17731 = n16854 ^ n14932 ^ n7189 ;
  assign n17732 = n14244 ^ n459 ^ 1'b0 ;
  assign n17733 = n4018 & ~n15889 ;
  assign n17734 = n17733 ^ n10788 ^ 1'b0 ;
  assign n17735 = ( n2203 & ~n4403 ) | ( n2203 & n4674 ) | ( ~n4403 & n4674 ) ;
  assign n17736 = ( x69 & n1783 ) | ( x69 & n17735 ) | ( n1783 & n17735 ) ;
  assign n17741 = ( ~n824 & n1447 ) | ( ~n824 & n2042 ) | ( n1447 & n2042 ) ;
  assign n17742 = n17741 ^ n3666 ^ n1621 ;
  assign n17738 = n4654 ^ n243 ^ 1'b0 ;
  assign n17739 = n2292 & n17738 ;
  assign n17737 = n14788 ^ n9080 ^ n5256 ;
  assign n17740 = n17739 ^ n17737 ^ n677 ;
  assign n17743 = n17742 ^ n17740 ^ n2422 ;
  assign n17744 = n1832 & n6952 ;
  assign n17745 = n15219 ^ n14066 ^ 1'b0 ;
  assign n17746 = n16434 ^ n14034 ^ 1'b0 ;
  assign n17747 = n17746 ^ n3726 ^ 1'b0 ;
  assign n17748 = n1280 | n2661 ;
  assign n17749 = n14752 ^ n3591 ^ n197 ;
  assign n17750 = n2132 & n17749 ;
  assign n17751 = n9940 | n12860 ;
  assign n17752 = n8728 & ~n17751 ;
  assign n17753 = n17752 ^ n10909 ^ 1'b0 ;
  assign n17754 = n592 | n7492 ;
  assign n17755 = n5003 | n14690 ;
  assign n17756 = n1231 | n8820 ;
  assign n17757 = n9915 | n17756 ;
  assign n17758 = n17755 & ~n17757 ;
  assign n17759 = n9922 | n17758 ;
  assign n17760 = n3993 & n15514 ;
  assign n17761 = ( ~n3653 & n17759 ) | ( ~n3653 & n17760 ) | ( n17759 & n17760 ) ;
  assign n17764 = n4793 ^ n4695 ^ n2137 ;
  assign n17762 = n2471 & n8334 ;
  assign n17763 = n17762 ^ n10727 ^ 1'b0 ;
  assign n17765 = n17764 ^ n17763 ^ n15103 ;
  assign n17766 = n4704 & n10266 ;
  assign n17767 = n16864 ^ n12395 ^ n2472 ;
  assign n17768 = n17767 ^ n10300 ^ n8652 ;
  assign n17769 = n17766 & n17768 ;
  assign n17770 = n17769 ^ n12762 ^ 1'b0 ;
  assign n17771 = n5531 | n7281 ;
  assign n17772 = n17771 ^ n4471 ^ 1'b0 ;
  assign n17773 = n12772 | n17772 ;
  assign n17774 = ( n5524 & n10777 ) | ( n5524 & n17697 ) | ( n10777 & n17697 ) ;
  assign n17775 = ( n15041 & ~n17773 ) | ( n15041 & n17774 ) | ( ~n17773 & n17774 ) ;
  assign n17776 = n15035 ^ n10769 ^ n3938 ;
  assign n17777 = n14932 ^ n4718 ^ n3728 ;
  assign n17778 = n3174 & ~n8921 ;
  assign n17779 = ~n10677 & n17778 ;
  assign n17780 = ( n14590 & ~n17777 ) | ( n14590 & n17779 ) | ( ~n17777 & n17779 ) ;
  assign n17781 = n17780 ^ n2982 ^ n2907 ;
  assign n17786 = n15514 ^ n3836 ^ n1113 ;
  assign n17783 = n2030 ^ n1472 ^ 1'b0 ;
  assign n17784 = n1444 & ~n17783 ;
  assign n17785 = n17784 ^ n8337 ^ n3585 ;
  assign n17782 = n5025 & n17408 ;
  assign n17787 = n17786 ^ n17785 ^ n17782 ;
  assign n17788 = n11828 ^ n10187 ^ 1'b0 ;
  assign n17789 = ( ~n13706 & n13912 ) | ( ~n13706 & n15441 ) | ( n13912 & n15441 ) ;
  assign n17790 = n17789 ^ n2067 ^ 1'b0 ;
  assign n17791 = n15848 ^ n13230 ^ n11855 ;
  assign n17792 = ( ~n7322 & n7943 ) | ( ~n7322 & n11289 ) | ( n7943 & n11289 ) ;
  assign n17793 = ~n9371 & n12949 ;
  assign n17794 = n17793 ^ n11493 ^ 1'b0 ;
  assign n17795 = ~n12053 & n16502 ;
  assign n17796 = n8740 & n10605 ;
  assign n17797 = ~n3054 & n3953 ;
  assign n17798 = n17797 ^ n2492 ^ 1'b0 ;
  assign n17799 = n17798 ^ n4349 ^ 1'b0 ;
  assign n17804 = ( ~n5149 & n9581 ) | ( ~n5149 & n17120 ) | ( n9581 & n17120 ) ;
  assign n17805 = ( n863 & n10706 ) | ( n863 & n17804 ) | ( n10706 & n17804 ) ;
  assign n17800 = x23 & n1017 ;
  assign n17801 = ~n2876 & n17800 ;
  assign n17802 = n9747 | n17801 ;
  assign n17803 = ~n10218 & n17802 ;
  assign n17806 = n17805 ^ n17803 ^ 1'b0 ;
  assign n17807 = n1867 & n17806 ;
  assign n17808 = ~n1357 & n17807 ;
  assign n17811 = ~n823 & n12523 ;
  assign n17812 = n17811 ^ n9604 ^ 1'b0 ;
  assign n17813 = ~n11189 & n17812 ;
  assign n17809 = n14330 ^ n2898 ^ 1'b0 ;
  assign n17810 = n16475 | n17809 ;
  assign n17814 = n17813 ^ n17810 ^ 1'b0 ;
  assign n17815 = n17590 ^ n4699 ^ n4555 ;
  assign n17816 = n16894 ^ n12652 ^ 1'b0 ;
  assign n17817 = n17815 & n17816 ;
  assign n17818 = n7684 & ~n17596 ;
  assign n17819 = n17818 ^ n3023 ^ 1'b0 ;
  assign n17820 = ( n8962 & n15880 ) | ( n8962 & ~n17819 ) | ( n15880 & ~n17819 ) ;
  assign n17821 = n2485 & ~n7685 ;
  assign n17822 = n5108 | n11988 ;
  assign n17823 = n3352 | n17822 ;
  assign n17824 = n17823 ^ n2604 ^ 1'b0 ;
  assign n17825 = n16268 & n17824 ;
  assign n17826 = n17825 ^ n6461 ^ 1'b0 ;
  assign n17827 = n256 & ~n2970 ;
  assign n17828 = n11469 & ~n17827 ;
  assign n17829 = n17828 ^ n1251 ^ 1'b0 ;
  assign n17830 = x53 & ~n3971 ;
  assign n17831 = n17829 & n17830 ;
  assign n17834 = n7408 & n13173 ;
  assign n17832 = ( n4372 & n6862 ) | ( n4372 & ~n8372 ) | ( n6862 & ~n8372 ) ;
  assign n17833 = n17832 ^ n7884 ^ n6176 ;
  assign n17835 = n17834 ^ n17833 ^ n4770 ;
  assign n17836 = ( n9590 & n10743 ) | ( n9590 & ~n11021 ) | ( n10743 & ~n11021 ) ;
  assign n17837 = ( n17831 & n17835 ) | ( n17831 & ~n17836 ) | ( n17835 & ~n17836 ) ;
  assign n17838 = ( n10438 & ~n17826 ) | ( n10438 & n17837 ) | ( ~n17826 & n17837 ) ;
  assign n17839 = ( n610 & n14185 ) | ( n610 & ~n14782 ) | ( n14185 & ~n14782 ) ;
  assign n17840 = n5327 ^ n1143 ^ 1'b0 ;
  assign n17841 = ~n4257 & n17840 ;
  assign n17842 = n17841 ^ n10370 ^ 1'b0 ;
  assign n17843 = n9103 ^ n248 ^ 1'b0 ;
  assign n17844 = n4380 & ~n17559 ;
  assign n17845 = ~n2886 & n17844 ;
  assign n17846 = ( ~n4285 & n4982 ) | ( ~n4285 & n15157 ) | ( n4982 & n15157 ) ;
  assign n17847 = ( ~n12483 & n15278 ) | ( ~n12483 & n15838 ) | ( n15278 & n15838 ) ;
  assign n17848 = ( ~n3853 & n15343 ) | ( ~n3853 & n16071 ) | ( n15343 & n16071 ) ;
  assign n17849 = ( ~n9311 & n9638 ) | ( ~n9311 & n17848 ) | ( n9638 & n17848 ) ;
  assign n17850 = x127 & ~n981 ;
  assign n17851 = n17849 & n17850 ;
  assign n17852 = ( n4920 & n9416 ) | ( n4920 & ~n10503 ) | ( n9416 & ~n10503 ) ;
  assign n17853 = n17852 ^ n17615 ^ n4645 ;
  assign n17854 = n3320 ^ n1392 ^ 1'b0 ;
  assign n17855 = n6931 & ~n17854 ;
  assign n17856 = ( ~n6773 & n17853 ) | ( ~n6773 & n17855 ) | ( n17853 & n17855 ) ;
  assign n17857 = ( n872 & n1932 ) | ( n872 & n10095 ) | ( n1932 & n10095 ) ;
  assign n17858 = n8882 | n17857 ;
  assign n17859 = n17856 | n17858 ;
  assign n17860 = n8391 ^ n2067 ^ 1'b0 ;
  assign n17861 = n8748 ^ n7151 ^ n5105 ;
  assign n17862 = n17861 ^ n11204 ^ n5983 ;
  assign n17863 = ( n3346 & n8255 ) | ( n3346 & ~n9545 ) | ( n8255 & ~n9545 ) ;
  assign n17864 = n14895 ^ n12811 ^ n1280 ;
  assign n17865 = ( ~n10157 & n17863 ) | ( ~n10157 & n17864 ) | ( n17863 & n17864 ) ;
  assign n17866 = ( n2318 & n6675 ) | ( n2318 & ~n11109 ) | ( n6675 & ~n11109 ) ;
  assign n17867 = n2778 | n16650 ;
  assign n17868 = n17867 ^ n2455 ^ 1'b0 ;
  assign n17869 = n7989 ^ n5522 ^ n622 ;
  assign n17870 = n17869 ^ n8637 ^ 1'b0 ;
  assign n17871 = ~n17177 & n17870 ;
  assign n17872 = ~n468 & n17266 ;
  assign n17873 = n17872 ^ n9391 ^ 1'b0 ;
  assign n17874 = n14602 ^ n13160 ^ n12375 ;
  assign n17876 = n8550 ^ n6149 ^ 1'b0 ;
  assign n17877 = n17876 ^ n3985 ^ 1'b0 ;
  assign n17878 = x55 & n17877 ;
  assign n17875 = ( ~n6282 & n13600 ) | ( ~n6282 & n16665 ) | ( n13600 & n16665 ) ;
  assign n17879 = n17878 ^ n17875 ^ n5508 ;
  assign n17880 = n5837 ^ n5729 ^ n1073 ;
  assign n17881 = n12734 ^ n9569 ^ 1'b0 ;
  assign n17882 = ~n11583 & n17881 ;
  assign n17883 = ~n9481 & n17882 ;
  assign n17884 = ~n1112 & n17883 ;
  assign n17885 = n11793 ^ n182 ^ 1'b0 ;
  assign n17886 = n17885 ^ n13007 ^ 1'b0 ;
  assign n17887 = ~n11075 & n11563 ;
  assign n17888 = ~n3921 & n17887 ;
  assign n17889 = ( n688 & n771 ) | ( n688 & ~n12033 ) | ( n771 & ~n12033 ) ;
  assign n17890 = n16534 & n17889 ;
  assign n17891 = n3612 & n5777 ;
  assign n17895 = n1079 | n16197 ;
  assign n17892 = n4508 & ~n7965 ;
  assign n17893 = n17892 ^ n10010 ^ n10007 ;
  assign n17894 = n2187 & ~n17893 ;
  assign n17896 = n17895 ^ n17894 ^ 1'b0 ;
  assign n17897 = n6906 & ~n11712 ;
  assign n17898 = ~n10248 & n17897 ;
  assign n17899 = n17898 ^ n15273 ^ n11950 ;
  assign n17900 = n8346 ^ n3103 ^ n1489 ;
  assign n17901 = n5616 | n10982 ;
  assign n17902 = ( n405 & n5904 ) | ( n405 & n15731 ) | ( n5904 & n15731 ) ;
  assign n17903 = n2640 | n17902 ;
  assign n17904 = ~n16848 & n17903 ;
  assign n17905 = n17904 ^ n14151 ^ 1'b0 ;
  assign n17906 = ( x33 & ~n5916 ) | ( x33 & n7318 ) | ( ~n5916 & n7318 ) ;
  assign n17907 = ( n766 & n4514 ) | ( n766 & n9242 ) | ( n4514 & n9242 ) ;
  assign n17908 = n5405 ^ n2680 ^ 1'b0 ;
  assign n17909 = ( n10593 & n12353 ) | ( n10593 & n17908 ) | ( n12353 & n17908 ) ;
  assign n17910 = ( n4810 & ~n11452 ) | ( n4810 & n17909 ) | ( ~n11452 & n17909 ) ;
  assign n17911 = n14641 | n17910 ;
  assign n17912 = n17911 ^ n3164 ^ 1'b0 ;
  assign n17913 = n14415 ^ n9738 ^ n5235 ;
  assign n17914 = n3789 | n4477 ;
  assign n17915 = n17914 ^ n7687 ^ 1'b0 ;
  assign n17916 = n17915 ^ n6679 ^ n4040 ;
  assign n17917 = n3390 & n3992 ;
  assign n17918 = n15479 ^ n8389 ^ 1'b0 ;
  assign n17919 = ~n2571 & n17918 ;
  assign n17920 = n17919 ^ n1595 ^ n642 ;
  assign n17921 = n6594 & n12218 ;
  assign n17922 = n14797 ^ n2265 ^ 1'b0 ;
  assign n17923 = n11108 ^ n6986 ^ n1679 ;
  assign n17924 = ( n3996 & ~n11440 ) | ( n3996 & n16471 ) | ( ~n11440 & n16471 ) ;
  assign n17925 = ( n5844 & ~n8253 ) | ( n5844 & n10145 ) | ( ~n8253 & n10145 ) ;
  assign n17926 = ( n2849 & n7116 ) | ( n2849 & ~n17925 ) | ( n7116 & ~n17925 ) ;
  assign n17927 = n11440 | n13706 ;
  assign n17928 = n17927 ^ n7520 ^ 1'b0 ;
  assign n17929 = n10246 ^ n7286 ^ 1'b0 ;
  assign n17930 = n4654 | n17929 ;
  assign n17931 = n17930 ^ n9118 ^ 1'b0 ;
  assign n17932 = n10029 ^ n814 ^ 1'b0 ;
  assign n17933 = n12723 & n13402 ;
  assign n17934 = n17933 ^ n16036 ^ 1'b0 ;
  assign n17935 = n12902 ^ n11810 ^ n11298 ;
  assign n17936 = n14904 ^ n13771 ^ n3127 ;
  assign n17937 = n10029 ^ n1899 ^ n906 ;
  assign n17938 = n15467 ^ n5849 ^ n4230 ;
  assign n17941 = ~n753 & n3958 ;
  assign n17939 = n11469 ^ n3724 ^ n1022 ;
  assign n17940 = n9819 & n17939 ;
  assign n17942 = n17941 ^ n17940 ^ n9930 ;
  assign n17943 = ~n1442 & n5769 ;
  assign n17944 = n17943 ^ n16048 ^ 1'b0 ;
  assign n17945 = ~n1649 & n17944 ;
  assign n17946 = n4997 ^ n1488 ^ 1'b0 ;
  assign n17947 = n17946 ^ n17442 ^ n6972 ;
  assign n17948 = n17947 ^ n11487 ^ 1'b0 ;
  assign n17949 = n6987 & ~n17948 ;
  assign n17950 = n3665 ^ n673 ^ 1'b0 ;
  assign n17951 = ( n617 & ~n7482 ) | ( n617 & n17950 ) | ( ~n7482 & n17950 ) ;
  assign n17952 = n9731 ^ n9704 ^ n785 ;
  assign n17953 = n17952 ^ n7722 ^ n3756 ;
  assign n17956 = n4408 & ~n6183 ;
  assign n17957 = n17956 ^ n7651 ^ 1'b0 ;
  assign n17958 = n17001 & n17957 ;
  assign n17954 = ( n3242 & n9898 ) | ( n3242 & ~n14712 ) | ( n9898 & ~n14712 ) ;
  assign n17955 = n6928 & ~n17954 ;
  assign n17959 = n17958 ^ n17955 ^ 1'b0 ;
  assign n17960 = n17959 ^ n5369 ^ n3006 ;
  assign n17961 = n13657 ^ n13398 ^ n6628 ;
  assign n17969 = n13100 ^ n7961 ^ 1'b0 ;
  assign n17970 = n3702 | n17969 ;
  assign n17962 = n5817 | n12202 ;
  assign n17963 = n3035 | n17962 ;
  assign n17964 = n8975 ^ n2304 ^ 1'b0 ;
  assign n17965 = n10356 & n17964 ;
  assign n17966 = n17963 & n17965 ;
  assign n17967 = n17966 ^ n12011 ^ 1'b0 ;
  assign n17968 = n5915 | n17967 ;
  assign n17971 = n17970 ^ n17968 ^ 1'b0 ;
  assign n17972 = ~n975 & n17021 ;
  assign n17973 = n17972 ^ n14180 ^ 1'b0 ;
  assign n17974 = n9128 & n17540 ;
  assign n17975 = n17974 ^ n2839 ^ 1'b0 ;
  assign n17976 = n1967 | n8314 ;
  assign n17977 = n17976 ^ n1226 ^ 1'b0 ;
  assign n17978 = ( n8261 & n17448 ) | ( n8261 & n17977 ) | ( n17448 & n17977 ) ;
  assign n17979 = n3435 | n5232 ;
  assign n17980 = n12045 | n17979 ;
  assign n17981 = ~n13605 & n17980 ;
  assign n17982 = ~n10046 & n17981 ;
  assign n17983 = n10371 & n12740 ;
  assign n17984 = n10699 & n17983 ;
  assign n17985 = ~n17982 & n17984 ;
  assign n17986 = n17929 ^ n11372 ^ n7093 ;
  assign n17987 = n3406 | n17986 ;
  assign n17989 = n5348 ^ n405 ^ 1'b0 ;
  assign n17990 = ( n6853 & ~n12462 ) | ( n6853 & n17989 ) | ( ~n12462 & n17989 ) ;
  assign n17988 = n15104 ^ n4220 ^ 1'b0 ;
  assign n17991 = n17990 ^ n17988 ^ 1'b0 ;
  assign n17992 = n7257 ^ n2172 ^ 1'b0 ;
  assign n17993 = n6035 | n17992 ;
  assign n17994 = n17993 ^ n16115 ^ 1'b0 ;
  assign n17995 = n17292 ^ n8466 ^ n275 ;
  assign n17996 = ( x108 & n2916 ) | ( x108 & n17995 ) | ( n2916 & n17995 ) ;
  assign n17997 = ( n6050 & n14587 ) | ( n6050 & n17996 ) | ( n14587 & n17996 ) ;
  assign n17998 = n13881 | n17997 ;
  assign n17999 = n6766 & ~n17998 ;
  assign n18000 = ( n2529 & n5193 ) | ( n2529 & n10447 ) | ( n5193 & n10447 ) ;
  assign n18001 = n18000 ^ n7968 ^ 1'b0 ;
  assign n18002 = n4687 | n13627 ;
  assign n18003 = n12653 | n18002 ;
  assign n18004 = ( n4018 & n11300 ) | ( n4018 & n18003 ) | ( n11300 & n18003 ) ;
  assign n18005 = n5710 | n9758 ;
  assign n18006 = n18005 ^ n11769 ^ 1'b0 ;
  assign n18007 = n18006 ^ n11442 ^ n7943 ;
  assign n18008 = n4172 ^ n2096 ^ n1555 ;
  assign n18009 = ( n3483 & n3593 ) | ( n3483 & n18008 ) | ( n3593 & n18008 ) ;
  assign n18010 = ~n12424 & n18009 ;
  assign n18017 = n13551 ^ n6799 ^ n4521 ;
  assign n18011 = n12350 ^ n5052 ^ 1'b0 ;
  assign n18012 = n18011 ^ n12024 ^ n8122 ;
  assign n18013 = n1199 | n18012 ;
  assign n18014 = n10429 & ~n18013 ;
  assign n18015 = n5343 | n18014 ;
  assign n18016 = n18015 ^ n15159 ^ n13781 ;
  assign n18018 = n18017 ^ n18016 ^ n8950 ;
  assign n18019 = n9117 | n11815 ;
  assign n18023 = n1827 ^ n1239 ^ 1'b0 ;
  assign n18024 = n5014 & n7606 ;
  assign n18025 = ~n18023 & n18024 ;
  assign n18026 = n10762 & n18025 ;
  assign n18027 = n130 & ~n18026 ;
  assign n18028 = n18027 ^ n8503 ^ 1'b0 ;
  assign n18020 = ( ~n5178 & n6862 ) | ( ~n5178 & n7420 ) | ( n6862 & n7420 ) ;
  assign n18021 = ( ~n3123 & n14792 ) | ( ~n3123 & n18020 ) | ( n14792 & n18020 ) ;
  assign n18022 = n3035 & ~n18021 ;
  assign n18029 = n18028 ^ n18022 ^ 1'b0 ;
  assign n18031 = n5242 | n8757 ;
  assign n18030 = ~n2557 & n10266 ;
  assign n18032 = n18031 ^ n18030 ^ 1'b0 ;
  assign n18033 = ( n5869 & ~n6338 ) | ( n5869 & n14010 ) | ( ~n6338 & n14010 ) ;
  assign n18034 = ~n12835 & n18033 ;
  assign n18035 = ~n5098 & n7352 ;
  assign n18036 = n18034 & n18035 ;
  assign n18037 = ( ~n2053 & n7181 ) | ( ~n2053 & n17278 ) | ( n7181 & n17278 ) ;
  assign n18038 = n8793 ^ n1924 ^ 1'b0 ;
  assign n18039 = n787 | n18038 ;
  assign n18040 = ( n5489 & n7031 ) | ( n5489 & ~n18039 ) | ( n7031 & ~n18039 ) ;
  assign n18041 = n5660 & n18040 ;
  assign n18042 = n18041 ^ n17509 ^ 1'b0 ;
  assign n18043 = ( n1451 & n9539 ) | ( n1451 & ~n11616 ) | ( n9539 & ~n11616 ) ;
  assign n18044 = ( n905 & n2174 ) | ( n905 & n18043 ) | ( n2174 & n18043 ) ;
  assign n18045 = ( n8202 & n11256 ) | ( n8202 & n18044 ) | ( n11256 & n18044 ) ;
  assign n18046 = n14047 | n18045 ;
  assign n18047 = n18042 | n18046 ;
  assign n18048 = ~n4793 & n9860 ;
  assign n18049 = ( ~n10104 & n15266 ) | ( ~n10104 & n18048 ) | ( n15266 & n18048 ) ;
  assign n18050 = n934 | n18049 ;
  assign n18051 = n13082 | n18050 ;
  assign n18054 = n13249 ^ n235 ^ 1'b0 ;
  assign n18055 = n5496 & ~n18054 ;
  assign n18053 = n9627 ^ n6128 ^ n2350 ;
  assign n18052 = n10306 ^ n7208 ^ 1'b0 ;
  assign n18056 = n18055 ^ n18053 ^ n18052 ;
  assign n18060 = n2265 & ~n5316 ;
  assign n18057 = n510 | n13792 ;
  assign n18058 = n1859 | n18057 ;
  assign n18059 = ( n10022 & n15107 ) | ( n10022 & n18058 ) | ( n15107 & n18058 ) ;
  assign n18061 = n18060 ^ n18059 ^ n17241 ;
  assign n18062 = ( n2370 & n14302 ) | ( n2370 & ~n16368 ) | ( n14302 & ~n16368 ) ;
  assign n18063 = n18062 ^ n8406 ^ n5480 ;
  assign n18064 = ( ~n2615 & n5414 ) | ( ~n2615 & n18063 ) | ( n5414 & n18063 ) ;
  assign n18065 = ( ~n14087 & n14916 ) | ( ~n14087 & n18064 ) | ( n14916 & n18064 ) ;
  assign n18066 = n15830 & n16915 ;
  assign n18067 = n18066 ^ n8779 ^ 1'b0 ;
  assign n18068 = n6624 ^ n5395 ^ 1'b0 ;
  assign n18069 = ( n488 & n1989 ) | ( n488 & ~n7454 ) | ( n1989 & ~n7454 ) ;
  assign n18070 = ~n5582 & n18069 ;
  assign n18071 = n18070 ^ n2369 ^ 1'b0 ;
  assign n18072 = ( ~n227 & n345 ) | ( ~n227 & n12826 ) | ( n345 & n12826 ) ;
  assign n18073 = n18072 ^ n12327 ^ 1'b0 ;
  assign n18074 = ( n265 & n2970 ) | ( n265 & n18073 ) | ( n2970 & n18073 ) ;
  assign n18075 = ~n576 & n12865 ;
  assign n18076 = n18075 ^ n2837 ^ 1'b0 ;
  assign n18077 = ( n12661 & n18074 ) | ( n12661 & ~n18076 ) | ( n18074 & ~n18076 ) ;
  assign n18078 = n2853 & ~n8799 ;
  assign n18079 = n18078 ^ n8158 ^ 1'b0 ;
  assign n18080 = n18077 | n18079 ;
  assign n18081 = n17225 ^ n10688 ^ n3816 ;
  assign n18082 = n11160 & ~n18081 ;
  assign n18083 = n1738 & n18082 ;
  assign n18084 = ( n3456 & n14752 ) | ( n3456 & n18083 ) | ( n14752 & n18083 ) ;
  assign n18085 = ( n12919 & n14080 ) | ( n12919 & n18084 ) | ( n14080 & n18084 ) ;
  assign n18086 = ( n2445 & n11275 ) | ( n2445 & n17954 ) | ( n11275 & n17954 ) ;
  assign n18093 = n16219 ^ n5576 ^ 1'b0 ;
  assign n18094 = n1260 & ~n18093 ;
  assign n18091 = n14909 ^ n3995 ^ 1'b0 ;
  assign n18092 = n3908 | n18091 ;
  assign n18087 = ~n1771 & n16517 ;
  assign n18088 = ~n2178 & n18087 ;
  assign n18089 = n5266 ^ n5119 ^ n1381 ;
  assign n18090 = n18088 & n18089 ;
  assign n18095 = n18094 ^ n18092 ^ n18090 ;
  assign n18096 = ( n1862 & n1926 ) | ( n1862 & n9674 ) | ( n1926 & n9674 ) ;
  assign n18097 = x104 & ~n17618 ;
  assign n18098 = ~n1168 & n18097 ;
  assign n18099 = n18098 ^ n5692 ^ n2295 ;
  assign n18100 = ( n15963 & ~n18096 ) | ( n15963 & n18099 ) | ( ~n18096 & n18099 ) ;
  assign n18101 = n8553 & n9109 ;
  assign n18102 = n2777 & n18101 ;
  assign n18103 = n2517 & n7184 ;
  assign n18104 = ( n7551 & n10079 ) | ( n7551 & n17729 ) | ( n10079 & n17729 ) ;
  assign n18105 = n4303 ^ n984 ^ n404 ;
  assign n18106 = n18105 ^ n1669 ^ 1'b0 ;
  assign n18107 = n901 | n18106 ;
  assign n18108 = ( ~n10117 & n14799 ) | ( ~n10117 & n18107 ) | ( n14799 & n18107 ) ;
  assign n18109 = ~n18104 & n18108 ;
  assign n18110 = n18109 ^ n7583 ^ 1'b0 ;
  assign n18111 = ( ~n8437 & n10383 ) | ( ~n8437 & n11815 ) | ( n10383 & n11815 ) ;
  assign n18112 = ( n10198 & n10325 ) | ( n10198 & ~n12009 ) | ( n10325 & ~n12009 ) ;
  assign n18113 = ( n8553 & n12307 ) | ( n8553 & n18112 ) | ( n12307 & n18112 ) ;
  assign n18114 = ( ~n1919 & n3888 ) | ( ~n1919 & n6731 ) | ( n3888 & n6731 ) ;
  assign n18115 = n15486 | n18114 ;
  assign n18116 = n18115 ^ n8067 ^ 1'b0 ;
  assign n18117 = n387 | n18116 ;
  assign n18118 = n3345 & ~n15406 ;
  assign n18119 = n10986 ^ n2582 ^ 1'b0 ;
  assign n18120 = ~n9071 & n18119 ;
  assign n18121 = n5563 | n14358 ;
  assign n18122 = n5784 & ~n18121 ;
  assign n18123 = n18122 ^ n3816 ^ 1'b0 ;
  assign n18124 = n1144 | n3565 ;
  assign n18125 = n16239 ^ n10079 ^ 1'b0 ;
  assign n18128 = n6775 ^ n3758 ^ 1'b0 ;
  assign n18129 = n3755 | n18128 ;
  assign n18126 = n8202 ^ n1324 ^ 1'b0 ;
  assign n18127 = n6195 & ~n18126 ;
  assign n18130 = n18129 ^ n18127 ^ n3721 ;
  assign n18131 = n2710 & ~n8017 ;
  assign n18132 = n18131 ^ n10533 ^ 1'b0 ;
  assign n18135 = n11795 ^ n2915 ^ n1987 ;
  assign n18133 = ~n2791 & n3543 ;
  assign n18134 = n7452 & n18133 ;
  assign n18136 = n18135 ^ n18134 ^ n270 ;
  assign n18137 = n16298 ^ n8687 ^ n3567 ;
  assign n18138 = n9571 ^ n5225 ^ n3360 ;
  assign n18139 = ~n7853 & n18138 ;
  assign n18140 = ~n8766 & n18139 ;
  assign n18141 = ( n10635 & n11653 ) | ( n10635 & n18140 ) | ( n11653 & n18140 ) ;
  assign n18142 = n10581 ^ n8103 ^ n1977 ;
  assign n18143 = n1427 ^ n518 ^ 1'b0 ;
  assign n18144 = n10482 | n18143 ;
  assign n18145 = n18144 ^ n4023 ^ 1'b0 ;
  assign n18146 = n18145 ^ n15580 ^ n11545 ;
  assign n18147 = n2519 | n7927 ;
  assign n18148 = ( n2819 & ~n18146 ) | ( n2819 & n18147 ) | ( ~n18146 & n18147 ) ;
  assign n18149 = n18148 ^ n10063 ^ 1'b0 ;
  assign n18150 = n9221 ^ x23 ^ 1'b0 ;
  assign n18151 = n18149 | n18150 ;
  assign n18152 = n1878 & ~n7928 ;
  assign n18153 = n18152 ^ n7989 ^ 1'b0 ;
  assign n18154 = n3298 | n18153 ;
  assign n18155 = n18151 & ~n18154 ;
  assign n18156 = n13801 ^ n10767 ^ n8157 ;
  assign n18157 = n18156 ^ n14210 ^ n3485 ;
  assign n18158 = n15933 ^ n602 ^ 1'b0 ;
  assign n18159 = ( ~n243 & n2135 ) | ( ~n243 & n18158 ) | ( n2135 & n18158 ) ;
  assign n18163 = ( n6193 & n7052 ) | ( n6193 & ~n9297 ) | ( n7052 & ~n9297 ) ;
  assign n18161 = n5974 ^ n1097 ^ n1014 ;
  assign n18160 = n4585 ^ n1830 ^ x15 ;
  assign n18162 = n18161 ^ n18160 ^ n2827 ;
  assign n18164 = n18163 ^ n18162 ^ 1'b0 ;
  assign n18165 = n12594 ^ n3830 ^ n2326 ;
  assign n18166 = n18165 ^ n5910 ^ n3517 ;
  assign n18167 = n3055 ^ n2863 ^ n1605 ;
  assign n18168 = n18167 ^ n6746 ^ 1'b0 ;
  assign n18169 = n2183 | n18168 ;
  assign n18170 = n2037 & ~n6607 ;
  assign n18171 = n14545 ^ n10625 ^ 1'b0 ;
  assign n18172 = n18170 & ~n18171 ;
  assign n18173 = n18169 & n18172 ;
  assign n18174 = n17087 ^ n7020 ^ 1'b0 ;
  assign n18175 = n725 | n4826 ;
  assign n18176 = n3832 & ~n9310 ;
  assign n18177 = n7728 & n18176 ;
  assign n18178 = ( n13860 & ~n18175 ) | ( n13860 & n18177 ) | ( ~n18175 & n18177 ) ;
  assign n18179 = ( n856 & n1838 ) | ( n856 & n10065 ) | ( n1838 & n10065 ) ;
  assign n18180 = n8834 ^ n2053 ^ 1'b0 ;
  assign n18181 = n18180 ^ n11403 ^ n1263 ;
  assign n18182 = n18181 ^ n12369 ^ 1'b0 ;
  assign n18183 = ~n6442 & n18182 ;
  assign n18186 = n10827 ^ n10661 ^ n2750 ;
  assign n18184 = n14291 ^ n13155 ^ 1'b0 ;
  assign n18185 = ~n778 & n18184 ;
  assign n18187 = n18186 ^ n18185 ^ n5660 ;
  assign n18188 = n14094 | n18187 ;
  assign n18189 = n12960 ^ n8639 ^ 1'b0 ;
  assign n18191 = n6692 ^ n4461 ^ n2759 ;
  assign n18190 = ~n11495 & n13667 ;
  assign n18192 = n18191 ^ n18190 ^ n1068 ;
  assign n18193 = n12407 ^ n3031 ^ 1'b0 ;
  assign n18194 = n6177 & n10515 ;
  assign n18195 = n7250 & n18194 ;
  assign n18196 = ( n964 & n1679 ) | ( n964 & ~n7208 ) | ( n1679 & ~n7208 ) ;
  assign n18197 = n18196 ^ n7632 ^ 1'b0 ;
  assign n18198 = ( n292 & n2600 ) | ( n292 & ~n2949 ) | ( n2600 & ~n2949 ) ;
  assign n18199 = n18198 ^ n16031 ^ 1'b0 ;
  assign n18200 = ( ~n7017 & n18197 ) | ( ~n7017 & n18199 ) | ( n18197 & n18199 ) ;
  assign n18201 = ( n9607 & n12109 ) | ( n9607 & ~n14956 ) | ( n12109 & ~n14956 ) ;
  assign n18202 = n2959 ^ n1314 ^ 1'b0 ;
  assign n18203 = ( n2464 & n5772 ) | ( n2464 & ~n18202 ) | ( n5772 & ~n18202 ) ;
  assign n18204 = ( ~n3333 & n4226 ) | ( ~n3333 & n13858 ) | ( n4226 & n13858 ) ;
  assign n18205 = n6391 ^ n1497 ^ 1'b0 ;
  assign n18206 = n18204 | n18205 ;
  assign n18207 = n11940 ^ n11402 ^ n5659 ;
  assign n18208 = n18207 ^ n7622 ^ 1'b0 ;
  assign n18209 = n13529 ^ n2379 ^ n2147 ;
  assign n18210 = n16195 ^ n5696 ^ 1'b0 ;
  assign n18211 = n18210 ^ n12534 ^ n345 ;
  assign n18212 = n696 & n1133 ;
  assign n18213 = n18212 ^ n16333 ^ n3510 ;
  assign n18214 = n3138 ^ n1844 ^ 1'b0 ;
  assign n18215 = n12430 | n18214 ;
  assign n18216 = n10479 ^ n6080 ^ 1'b0 ;
  assign n18217 = n3019 | n18216 ;
  assign n18218 = n17721 & ~n18217 ;
  assign n18219 = n9744 & ~n12071 ;
  assign n18220 = n3756 | n18219 ;
  assign n18221 = n13781 & ~n18220 ;
  assign n18222 = n13735 ^ n4622 ^ n1664 ;
  assign n18223 = n7787 & n10740 ;
  assign n18224 = n18222 & n18223 ;
  assign n18225 = ( n7943 & ~n9661 ) | ( n7943 & n18224 ) | ( ~n9661 & n18224 ) ;
  assign n18226 = ( ~n11795 & n18221 ) | ( ~n11795 & n18225 ) | ( n18221 & n18225 ) ;
  assign n18227 = n15923 & ~n18226 ;
  assign n18228 = n17591 ^ n6274 ^ n2086 ;
  assign n18229 = n10361 & ~n18166 ;
  assign n18230 = n18229 ^ n3754 ^ 1'b0 ;
  assign n18231 = ~n1738 & n8372 ;
  assign n18232 = ~n3268 & n18231 ;
  assign n18233 = n447 | n18232 ;
  assign n18234 = n5837 & ~n18233 ;
  assign n18235 = n11659 ^ n5256 ^ 1'b0 ;
  assign n18236 = n14072 ^ n2254 ^ 1'b0 ;
  assign n18237 = n3063 | n18236 ;
  assign n18238 = ~n3795 & n10827 ;
  assign n18239 = n18238 ^ n7809 ^ 1'b0 ;
  assign n18240 = ~n5797 & n6673 ;
  assign n18241 = ~n589 & n5622 ;
  assign n18242 = n18240 & n18241 ;
  assign n18243 = n15419 ^ n11096 ^ 1'b0 ;
  assign n18244 = ~n1240 & n15123 ;
  assign n18245 = ~n13721 & n18244 ;
  assign n18246 = n6124 & ~n18245 ;
  assign n18247 = n18246 ^ n695 ^ 1'b0 ;
  assign n18248 = n5949 | n18247 ;
  assign n18252 = ~n4080 & n13306 ;
  assign n18253 = n10237 | n18252 ;
  assign n18254 = n18039 ^ n822 ^ 1'b0 ;
  assign n18255 = n7697 & n18254 ;
  assign n18256 = n18255 ^ n1956 ^ 1'b0 ;
  assign n18257 = n18253 & ~n18256 ;
  assign n18249 = n1530 | n9974 ;
  assign n18250 = n18249 ^ n9531 ^ n8177 ;
  assign n18251 = n18250 ^ n13131 ^ n10383 ;
  assign n18258 = n18257 ^ n18251 ^ n17768 ;
  assign n18259 = n7818 ^ n2467 ^ n2193 ;
  assign n18260 = n18259 ^ n17157 ^ n4216 ;
  assign n18261 = n18260 ^ n6580 ^ 1'b0 ;
  assign n18264 = n17523 ^ n13989 ^ n4448 ;
  assign n18265 = n1001 & n9251 ;
  assign n18266 = n18264 & ~n18265 ;
  assign n18262 = n2402 | n6802 ;
  assign n18263 = n5141 & ~n18262 ;
  assign n18267 = n18266 ^ n18263 ^ 1'b0 ;
  assign n18268 = ~n4542 & n4878 ;
  assign n18269 = ~n8268 & n18268 ;
  assign n18270 = n18269 ^ n5757 ^ n451 ;
  assign n18271 = n18270 ^ n11005 ^ 1'b0 ;
  assign n18272 = n2634 | n18271 ;
  assign n18273 = n13049 & ~n14927 ;
  assign n18275 = n8219 ^ n3955 ^ n1811 ;
  assign n18274 = n12486 ^ n10887 ^ n9104 ;
  assign n18276 = n18275 ^ n18274 ^ n10094 ;
  assign n18277 = n11792 ^ n2777 ^ 1'b0 ;
  assign n18278 = n10163 & n18277 ;
  assign n18279 = n18278 ^ n434 ^ 1'b0 ;
  assign n18280 = n18279 ^ n1282 ^ 1'b0 ;
  assign n18281 = n18280 ^ n7519 ^ n461 ;
  assign n18282 = n1477 ^ n410 ^ 1'b0 ;
  assign n18283 = ( n1145 & ~n18281 ) | ( n1145 & n18282 ) | ( ~n18281 & n18282 ) ;
  assign n18284 = n2030 & n11650 ;
  assign n18285 = n18284 ^ n13971 ^ 1'b0 ;
  assign n18288 = ( n4500 & n7780 ) | ( n4500 & n10437 ) | ( n7780 & n10437 ) ;
  assign n18286 = n14577 ^ n4429 ^ 1'b0 ;
  assign n18287 = n18286 ^ n1007 ^ x24 ;
  assign n18289 = n18288 ^ n18287 ^ 1'b0 ;
  assign n18290 = n18289 ^ n8389 ^ n3817 ;
  assign n18291 = n7034 & n18290 ;
  assign n18292 = ~n7883 & n17488 ;
  assign n18293 = n4784 & n18292 ;
  assign n18294 = n7416 ^ n5299 ^ 1'b0 ;
  assign n18295 = n2482 & ~n18294 ;
  assign n18296 = n14846 ^ n7073 ^ 1'b0 ;
  assign n18297 = n12390 & n17387 ;
  assign n18298 = n7002 & n18297 ;
  assign n18299 = n18298 ^ n5150 ^ 1'b0 ;
  assign n18300 = n10057 | n16749 ;
  assign n18301 = ( ~n10009 & n10620 ) | ( ~n10009 & n11544 ) | ( n10620 & n11544 ) ;
  assign n18302 = ( n5391 & n12505 ) | ( n5391 & ~n18301 ) | ( n12505 & ~n18301 ) ;
  assign n18303 = n18302 ^ n10911 ^ n2109 ;
  assign n18304 = ( n2063 & n6300 ) | ( n2063 & n8862 ) | ( n6300 & n8862 ) ;
  assign n18305 = ~n4140 & n16395 ;
  assign n18306 = n18305 ^ n413 ^ 1'b0 ;
  assign n18308 = ( ~x12 & n1186 ) | ( ~x12 & n1244 ) | ( n1186 & n1244 ) ;
  assign n18309 = ( n1761 & ~n6089 ) | ( n1761 & n18308 ) | ( ~n6089 & n18308 ) ;
  assign n18310 = ( ~n8295 & n11641 ) | ( ~n8295 & n18309 ) | ( n11641 & n18309 ) ;
  assign n18307 = n2554 | n11672 ;
  assign n18311 = n18310 ^ n18307 ^ 1'b0 ;
  assign n18313 = n1573 & ~n2955 ;
  assign n18314 = n4856 & n18313 ;
  assign n18312 = ( n3274 & n10755 ) | ( n3274 & n17401 ) | ( n10755 & n17401 ) ;
  assign n18315 = n18314 ^ n18312 ^ 1'b0 ;
  assign n18316 = x45 & ~n16319 ;
  assign n18317 = n14417 ^ n5920 ^ 1'b0 ;
  assign n18318 = ( ~n13179 & n18316 ) | ( ~n13179 & n18317 ) | ( n18316 & n18317 ) ;
  assign n18319 = n2867 & n5806 ;
  assign n18320 = ( n644 & n9153 ) | ( n644 & ~n18319 ) | ( n9153 & ~n18319 ) ;
  assign n18321 = n3561 | n13465 ;
  assign n18322 = n11913 | n13341 ;
  assign n18323 = ~n4333 & n12563 ;
  assign n18324 = ~n6729 & n18323 ;
  assign n18325 = n2731 | n18324 ;
  assign n18326 = n18322 | n18325 ;
  assign n18327 = n15982 ^ n13959 ^ n2741 ;
  assign n18328 = n5432 ^ n4819 ^ 1'b0 ;
  assign n18329 = n7097 & n18328 ;
  assign n18330 = n18329 ^ n2891 ^ 1'b0 ;
  assign n18331 = x21 & ~n18330 ;
  assign n18332 = ( ~n1424 & n15207 ) | ( ~n1424 & n18331 ) | ( n15207 & n18331 ) ;
  assign n18333 = n12785 | n13056 ;
  assign n18335 = n16755 ^ n8983 ^ 1'b0 ;
  assign n18334 = ~n1873 & n5299 ;
  assign n18336 = n18335 ^ n18334 ^ 1'b0 ;
  assign n18337 = n678 | n1193 ;
  assign n18338 = ( n1879 & n3945 ) | ( n1879 & ~n9965 ) | ( n3945 & ~n9965 ) ;
  assign n18339 = n15334 ^ n7971 ^ n7198 ;
  assign n18340 = n14361 ^ n11698 ^ 1'b0 ;
  assign n18341 = n2569 | n18340 ;
  assign n18342 = n5724 ^ n3698 ^ 1'b0 ;
  assign n18343 = n18342 ^ n3272 ^ n2913 ;
  assign n18344 = ~n493 & n6826 ;
  assign n18345 = n992 & n18344 ;
  assign n18346 = n6916 & ~n13121 ;
  assign n18347 = n18346 ^ n15302 ^ 1'b0 ;
  assign n18348 = ( ~n3389 & n4148 ) | ( ~n3389 & n6275 ) | ( n4148 & n6275 ) ;
  assign n18349 = n6472 & n18348 ;
  assign n18350 = ~n7064 & n18349 ;
  assign n18351 = ( n4088 & n5706 ) | ( n4088 & ~n10948 ) | ( n5706 & ~n10948 ) ;
  assign n18352 = n14169 & ~n18351 ;
  assign n18353 = n17629 ^ n17414 ^ n1519 ;
  assign n18354 = ( ~n2974 & n3586 ) | ( ~n2974 & n9226 ) | ( n3586 & n9226 ) ;
  assign n18355 = n406 & ~n8283 ;
  assign n18356 = n4549 & ~n18355 ;
  assign n18357 = n18356 ^ n13594 ^ n11386 ;
  assign n18358 = ~n1068 & n15918 ;
  assign n18359 = ~n8740 & n18358 ;
  assign n18360 = n752 | n1401 ;
  assign n18361 = n13498 | n18360 ;
  assign n18362 = n9657 & n10359 ;
  assign n18363 = n10569 & n18362 ;
  assign n18364 = ( n3648 & ~n18361 ) | ( n3648 & n18363 ) | ( ~n18361 & n18363 ) ;
  assign n18368 = n11522 ^ n2217 ^ 1'b0 ;
  assign n18369 = n6699 & n18368 ;
  assign n18370 = n14011 ^ n10220 ^ 1'b0 ;
  assign n18371 = n18369 & ~n18370 ;
  assign n18365 = n2668 & n6550 ;
  assign n18366 = ( ~n3125 & n9477 ) | ( ~n3125 & n15085 ) | ( n9477 & n15085 ) ;
  assign n18367 = ( ~n2190 & n18365 ) | ( ~n2190 & n18366 ) | ( n18365 & n18366 ) ;
  assign n18372 = n18371 ^ n18367 ^ n3956 ;
  assign n18373 = ~n8538 & n17195 ;
  assign n18374 = n16347 ^ n12722 ^ 1'b0 ;
  assign n18375 = ( n1493 & n1700 ) | ( n1493 & ~n4878 ) | ( n1700 & ~n4878 ) ;
  assign n18376 = ( n624 & n4813 ) | ( n624 & n18375 ) | ( n4813 & n18375 ) ;
  assign n18377 = ( n198 & n2547 ) | ( n198 & n18376 ) | ( n2547 & n18376 ) ;
  assign n18378 = n9147 & n18377 ;
  assign n18379 = n18378 ^ n7774 ^ 1'b0 ;
  assign n18380 = n5674 | n17901 ;
  assign n18381 = n18380 ^ n3298 ^ 1'b0 ;
  assign n18382 = n3134 & ~n13119 ;
  assign n18383 = n18382 ^ n10902 ^ 1'b0 ;
  assign n18384 = n4903 | n12228 ;
  assign n18385 = n18383 | n18384 ;
  assign n18386 = n7058 & n11653 ;
  assign n18387 = ~n5081 & n18386 ;
  assign n18388 = n18387 ^ n14423 ^ n8876 ;
  assign n18394 = ( n2911 & n2946 ) | ( n2911 & n17615 ) | ( n2946 & n17615 ) ;
  assign n18395 = n5206 & ~n18394 ;
  assign n18396 = n6081 & n18395 ;
  assign n18389 = n3626 ^ x30 ^ 1'b0 ;
  assign n18390 = n15703 & n18389 ;
  assign n18391 = ~n10011 & n18390 ;
  assign n18392 = n4045 & n8199 ;
  assign n18393 = n18391 & n18392 ;
  assign n18397 = n18396 ^ n18393 ^ n6356 ;
  assign n18398 = n18397 ^ n2151 ^ n1727 ;
  assign n18399 = n13777 & ~n18016 ;
  assign n18400 = n10821 & ~n11632 ;
  assign n18401 = n285 & n13092 ;
  assign n18402 = n18401 ^ n7363 ^ 1'b0 ;
  assign n18403 = n18402 ^ n1184 ^ 1'b0 ;
  assign n18404 = n18403 ^ n5429 ^ n2086 ;
  assign n18405 = ( n3360 & ~n18400 ) | ( n3360 & n18404 ) | ( ~n18400 & n18404 ) ;
  assign n18406 = n14544 ^ n1095 ^ 1'b0 ;
  assign n18407 = ~n1174 & n16131 ;
  assign n18408 = n18406 & n18407 ;
  assign n18409 = n16893 ^ n5389 ^ n424 ;
  assign n18410 = n12578 ^ n9661 ^ n1557 ;
  assign n18411 = ( ~n6786 & n16312 ) | ( ~n6786 & n18410 ) | ( n16312 & n18410 ) ;
  assign n18416 = ( n4127 & n13989 ) | ( n4127 & n17618 ) | ( n13989 & n17618 ) ;
  assign n18417 = n4596 | n18416 ;
  assign n18415 = n9208 ^ n6768 ^ 1'b0 ;
  assign n18412 = ~n4155 & n7722 ;
  assign n18413 = n18412 ^ n8689 ^ 1'b0 ;
  assign n18414 = n7459 & ~n18413 ;
  assign n18418 = n18417 ^ n18415 ^ n18414 ;
  assign n18419 = ( n2286 & n7458 ) | ( n2286 & ~n7832 ) | ( n7458 & ~n7832 ) ;
  assign n18420 = n4014 ^ n1648 ^ 1'b0 ;
  assign n18421 = ( n2543 & ~n16882 ) | ( n2543 & n18420 ) | ( ~n16882 & n18420 ) ;
  assign n18422 = n9105 | n9370 ;
  assign n18423 = ( n4503 & ~n17015 ) | ( n4503 & n18422 ) | ( ~n17015 & n18422 ) ;
  assign n18424 = n1714 & n18423 ;
  assign n18425 = n4471 & n18424 ;
  assign n18426 = ~n1090 & n6742 ;
  assign n18427 = ~n6005 & n18426 ;
  assign n18428 = n7375 | n18427 ;
  assign n18429 = n15580 & ~n18428 ;
  assign n18430 = ( n1679 & ~n2921 ) | ( n1679 & n18429 ) | ( ~n2921 & n18429 ) ;
  assign n18431 = n14779 ^ n13675 ^ n10002 ;
  assign n18439 = ( n2011 & n13273 ) | ( n2011 & n18308 ) | ( n13273 & n18308 ) ;
  assign n18440 = n18439 ^ n11417 ^ n8553 ;
  assign n18441 = ( n2623 & n4272 ) | ( n2623 & n8138 ) | ( n4272 & n8138 ) ;
  assign n18442 = n11398 & n13621 ;
  assign n18443 = n18441 & n18442 ;
  assign n18444 = ( n13721 & n18440 ) | ( n13721 & n18443 ) | ( n18440 & n18443 ) ;
  assign n18432 = ~n5245 & n15329 ;
  assign n18433 = n18432 ^ n16714 ^ 1'b0 ;
  assign n18436 = n6679 ^ n6535 ^ 1'b0 ;
  assign n18434 = n12992 ^ n364 ^ 1'b0 ;
  assign n18435 = n2086 | n18434 ;
  assign n18437 = n18436 ^ n18435 ^ n1911 ;
  assign n18438 = ~n18433 & n18437 ;
  assign n18445 = n18444 ^ n18438 ^ 1'b0 ;
  assign n18446 = n16125 ^ n4404 ^ 1'b0 ;
  assign n18447 = n6516 | n18446 ;
  assign n18448 = ( ~n5319 & n9159 ) | ( ~n5319 & n10955 ) | ( n9159 & n10955 ) ;
  assign n18449 = n2293 | n5693 ;
  assign n18450 = n18448 & ~n18449 ;
  assign n18451 = n5374 | n18450 ;
  assign n18452 = n6812 & ~n18451 ;
  assign n18453 = ~n351 & n7377 ;
  assign n18454 = ( n6409 & n18452 ) | ( n6409 & n18453 ) | ( n18452 & n18453 ) ;
  assign n18455 = n8298 ^ n3346 ^ n1880 ;
  assign n18456 = ( ~n6698 & n15900 ) | ( ~n6698 & n18455 ) | ( n15900 & n18455 ) ;
  assign n18457 = n9167 & ~n18456 ;
  assign n18458 = n18454 & n18457 ;
  assign n18459 = n5111 & n10577 ;
  assign n18460 = ( n10496 & ~n15903 ) | ( n10496 & n18459 ) | ( ~n15903 & n18459 ) ;
  assign n18462 = n13064 ^ n3711 ^ n2273 ;
  assign n18461 = n11265 ^ n2625 ^ n971 ;
  assign n18463 = n18462 ^ n18461 ^ n14313 ;
  assign n18464 = ( n7639 & n10469 ) | ( n7639 & ~n15724 ) | ( n10469 & ~n15724 ) ;
  assign n18465 = ~n673 & n6103 ;
  assign n18466 = n5745 & n18465 ;
  assign n18467 = n18466 ^ n15613 ^ 1'b0 ;
  assign n18468 = n15014 & ~n18467 ;
  assign n18469 = ~n5724 & n18468 ;
  assign n18470 = ( n16790 & n18464 ) | ( n16790 & n18469 ) | ( n18464 & n18469 ) ;
  assign n18471 = ~n1994 & n13917 ;
  assign n18472 = n3352 & ~n3912 ;
  assign n18473 = n18472 ^ n5092 ^ 1'b0 ;
  assign n18474 = n8946 ^ n5212 ^ 1'b0 ;
  assign n18475 = ( n1220 & ~n18473 ) | ( n1220 & n18474 ) | ( ~n18473 & n18474 ) ;
  assign n18476 = n1007 ^ n788 ^ 1'b0 ;
  assign n18477 = n1614 & ~n3896 ;
  assign n18478 = n9418 ^ n2835 ^ 1'b0 ;
  assign n18479 = n11382 | n16540 ;
  assign n18480 = n5979 & ~n18479 ;
  assign n18481 = ( ~n3061 & n3666 ) | ( ~n3061 & n6871 ) | ( n3666 & n6871 ) ;
  assign n18482 = n16076 & n18481 ;
  assign n18483 = n18480 & n18482 ;
  assign n18487 = n8082 & n12013 ;
  assign n18484 = n14053 ^ n9532 ^ n2467 ;
  assign n18485 = n18484 ^ n9902 ^ 1'b0 ;
  assign n18486 = n8221 & n18485 ;
  assign n18488 = n18487 ^ n18486 ^ n6260 ;
  assign n18491 = n13246 | n13754 ;
  assign n18492 = n6670 & ~n18491 ;
  assign n18489 = n16447 ^ n3593 ^ 1'b0 ;
  assign n18490 = n7583 & n18489 ;
  assign n18493 = n18492 ^ n18490 ^ 1'b0 ;
  assign n18494 = n3813 ^ n3447 ^ n1253 ;
  assign n18495 = ( n12307 & n15068 ) | ( n12307 & ~n18494 ) | ( n15068 & ~n18494 ) ;
  assign n18496 = ( n738 & n17188 ) | ( n738 & ~n18495 ) | ( n17188 & ~n18495 ) ;
  assign n18497 = ( ~n2048 & n4616 ) | ( ~n2048 & n18496 ) | ( n4616 & n18496 ) ;
  assign n18498 = n18497 ^ n2996 ^ 1'b0 ;
  assign n18499 = ~n1118 & n18498 ;
  assign n18500 = ( n368 & n5026 ) | ( n368 & n6828 ) | ( n5026 & n6828 ) ;
  assign n18501 = n2176 & ~n18500 ;
  assign n18502 = n6253 & n18501 ;
  assign n18503 = n10052 ^ n8405 ^ n549 ;
  assign n18504 = n5766 ^ n5380 ^ n5089 ;
  assign n18505 = ( n4150 & n18503 ) | ( n4150 & n18504 ) | ( n18503 & n18504 ) ;
  assign n18506 = n2364 | n18505 ;
  assign n18507 = n18371 | n18506 ;
  assign n18508 = n989 & n10476 ;
  assign n18509 = n13376 ^ n12099 ^ n9497 ;
  assign n18510 = n4793 & n4931 ;
  assign n18511 = ~n750 & n18510 ;
  assign n18512 = n3462 | n18511 ;
  assign n18513 = ( ~n7361 & n7871 ) | ( ~n7361 & n15900 ) | ( n7871 & n15900 ) ;
  assign n18514 = ( n4370 & ~n12049 ) | ( n4370 & n18513 ) | ( ~n12049 & n18513 ) ;
  assign n18515 = n18514 ^ n12729 ^ n1899 ;
  assign n18516 = n2085 & n3351 ;
  assign n18517 = n1340 & ~n2761 ;
  assign n18518 = n18517 ^ n1923 ^ n481 ;
  assign n18519 = n18518 ^ n11232 ^ 1'b0 ;
  assign n18520 = ( n2344 & n7056 ) | ( n2344 & ~n11183 ) | ( n7056 & ~n11183 ) ;
  assign n18521 = n9169 ^ n5449 ^ 1'b0 ;
  assign n18522 = n18521 ^ n561 ^ 1'b0 ;
  assign n18523 = n18522 ^ n16412 ^ n5627 ;
  assign n18524 = ( n5006 & n9169 ) | ( n5006 & ~n10031 ) | ( n9169 & ~n10031 ) ;
  assign n18525 = ~n8448 & n11078 ;
  assign n18526 = n18525 ^ n17915 ^ 1'b0 ;
  assign n18527 = n15139 ^ n4490 ^ n3661 ;
  assign n18528 = ( n7146 & n17662 ) | ( n7146 & ~n18527 ) | ( n17662 & ~n18527 ) ;
  assign n18529 = n8157 ^ n500 ^ 1'b0 ;
  assign n18530 = ~n18528 & n18529 ;
  assign n18531 = x32 | n13006 ;
  assign n18532 = n7800 & n14956 ;
  assign n18533 = ~n18531 & n18532 ;
  assign n18534 = n9549 ^ x76 ^ 1'b0 ;
  assign n18535 = ( n3330 & n5645 ) | ( n3330 & n18534 ) | ( n5645 & n18534 ) ;
  assign n18537 = n2154 ^ x92 ^ 1'b0 ;
  assign n18538 = n2424 & n18537 ;
  assign n18536 = n1858 & ~n5026 ;
  assign n18539 = n18538 ^ n18536 ^ n6845 ;
  assign n18541 = ~n1900 & n6746 ;
  assign n18540 = ~n2441 & n3079 ;
  assign n18542 = n18541 ^ n18540 ^ 1'b0 ;
  assign n18543 = n2254 & n11295 ;
  assign n18544 = ~n14385 & n18543 ;
  assign n18545 = n830 & n18042 ;
  assign n18546 = ~n11989 & n18545 ;
  assign n18547 = n18546 ^ n13706 ^ 1'b0 ;
  assign n18548 = n18547 ^ n2612 ^ 1'b0 ;
  assign n18549 = n3906 & ~n18548 ;
  assign n18554 = n9473 ^ n3436 ^ n1149 ;
  assign n18550 = n5133 ^ n3104 ^ 1'b0 ;
  assign n18551 = n7546 & ~n18550 ;
  assign n18552 = n3187 ^ n1253 ^ 1'b0 ;
  assign n18553 = n18551 & ~n18552 ;
  assign n18555 = n18554 ^ n18553 ^ n1539 ;
  assign n18556 = n12731 ^ n10762 ^ 1'b0 ;
  assign n18557 = ~n12075 & n17508 ;
  assign n18558 = n18557 ^ n12461 ^ n1777 ;
  assign n18559 = n15774 ^ n10818 ^ n9286 ;
  assign n18560 = ~n3042 & n3977 ;
  assign n18561 = n18560 ^ n2823 ^ 1'b0 ;
  assign n18562 = ( n2296 & n14424 ) | ( n2296 & ~n18561 ) | ( n14424 & ~n18561 ) ;
  assign n18563 = n1115 & ~n3280 ;
  assign n18564 = ( n4564 & ~n4733 ) | ( n4564 & n18563 ) | ( ~n4733 & n18563 ) ;
  assign n18565 = n8203 ^ n3608 ^ 1'b0 ;
  assign n18566 = ~n7205 & n18565 ;
  assign n18567 = n18564 | n18566 ;
  assign n18569 = n6261 ^ n825 ^ 1'b0 ;
  assign n18570 = n586 | n18569 ;
  assign n18571 = ( ~n8337 & n18107 ) | ( ~n8337 & n18570 ) | ( n18107 & n18570 ) ;
  assign n18568 = n10833 & ~n11358 ;
  assign n18572 = n18571 ^ n18568 ^ n13069 ;
  assign n18573 = n13111 ^ n1010 ^ n696 ;
  assign n18574 = n835 & n4672 ;
  assign n18575 = ~n5208 & n18574 ;
  assign n18576 = ( n2011 & n5196 ) | ( n2011 & n6778 ) | ( n5196 & n6778 ) ;
  assign n18577 = n5720 & ~n18576 ;
  assign n18578 = n18577 ^ n7638 ^ 1'b0 ;
  assign n18579 = ( n743 & ~n6866 ) | ( n743 & n13912 ) | ( ~n6866 & n13912 ) ;
  assign n18580 = ( n136 & n4172 ) | ( n136 & ~n18579 ) | ( n4172 & ~n18579 ) ;
  assign n18581 = n18580 ^ n2427 ^ 1'b0 ;
  assign n18582 = n18578 | n18581 ;
  assign n18583 = n17022 ^ n15027 ^ n11627 ;
  assign n18584 = ( n1268 & n15694 ) | ( n1268 & n18583 ) | ( n15694 & n18583 ) ;
  assign n18586 = n2378 ^ n1246 ^ 1'b0 ;
  assign n18587 = n3674 | n7435 ;
  assign n18588 = n2640 & ~n18587 ;
  assign n18589 = n18588 ^ n14714 ^ 1'b0 ;
  assign n18590 = n18586 & n18589 ;
  assign n18585 = ~n6501 & n10634 ;
  assign n18591 = n18590 ^ n18585 ^ 1'b0 ;
  assign n18592 = ( ~n312 & n14964 ) | ( ~n312 & n18591 ) | ( n14964 & n18591 ) ;
  assign n18593 = ( n924 & n2633 ) | ( n924 & ~n9422 ) | ( n2633 & ~n9422 ) ;
  assign n18594 = n11019 ^ n7067 ^ n4342 ;
  assign n18595 = n6006 ^ n2227 ^ 1'b0 ;
  assign n18596 = n18595 ^ n17138 ^ n410 ;
  assign n18597 = n16477 ^ n15447 ^ n2008 ;
  assign n18598 = n18562 ^ n11355 ^ n9344 ;
  assign n18599 = n12429 & n18598 ;
  assign n18600 = n8961 & n18599 ;
  assign n18603 = n7065 & n10112 ;
  assign n18604 = n2346 & n18603 ;
  assign n18601 = n9504 ^ n6931 ^ 1'b0 ;
  assign n18602 = n4962 & n18601 ;
  assign n18605 = n18604 ^ n18602 ^ 1'b0 ;
  assign n18606 = ~x23 & n1784 ;
  assign n18607 = ( n6042 & n8383 ) | ( n6042 & ~n18606 ) | ( n8383 & ~n18606 ) ;
  assign n18608 = ( n3107 & n6392 ) | ( n3107 & ~n12459 ) | ( n6392 & ~n12459 ) ;
  assign n18609 = ( n8711 & n10562 ) | ( n8711 & n16134 ) | ( n10562 & n16134 ) ;
  assign n18610 = ( n1375 & n5732 ) | ( n1375 & ~n18609 ) | ( n5732 & ~n18609 ) ;
  assign n18611 = n10321 ^ n9290 ^ n8434 ;
  assign n18612 = n2063 & n4105 ;
  assign n18613 = n18612 ^ n7486 ^ n2550 ;
  assign n18614 = n10950 ^ n10818 ^ x14 ;
  assign n18615 = n18614 ^ n17903 ^ n10504 ;
  assign n18616 = n7282 ^ n6116 ^ 1'b0 ;
  assign n18617 = ~n18615 & n18616 ;
  assign n18618 = n6845 ^ n4820 ^ n2016 ;
  assign n18619 = n5377 & n18618 ;
  assign n18620 = n18619 ^ n1583 ^ 1'b0 ;
  assign n18621 = n14945 | n18620 ;
  assign n18622 = ( n14381 & n16084 ) | ( n14381 & n18621 ) | ( n16084 & n18621 ) ;
  assign n18625 = n1022 & ~n4328 ;
  assign n18626 = ~n5706 & n18625 ;
  assign n18623 = n17954 ^ n15769 ^ n14964 ;
  assign n18624 = n18623 ^ n6776 ^ n2744 ;
  assign n18627 = n18626 ^ n18624 ^ n1403 ;
  assign n18628 = n14261 | n18627 ;
  assign n18629 = n3456 & ~n12237 ;
  assign n18630 = ~n3456 & n18629 ;
  assign n18631 = n9033 & ~n11517 ;
  assign n18632 = n18631 ^ n4885 ^ 1'b0 ;
  assign n18633 = n9131 & n18632 ;
  assign n18634 = n14769 ^ n13993 ^ n10659 ;
  assign n18635 = ~n4041 & n13267 ;
  assign n18636 = n18635 ^ n3666 ^ 1'b0 ;
  assign n18637 = ( n8695 & n11569 ) | ( n8695 & n18636 ) | ( n11569 & n18636 ) ;
  assign n18638 = n18637 ^ n3471 ^ n1412 ;
  assign n18639 = ( n1397 & n4164 ) | ( n1397 & ~n5408 ) | ( n4164 & ~n5408 ) ;
  assign n18640 = n18639 ^ n15646 ^ 1'b0 ;
  assign n18641 = n9536 ^ n2660 ^ 1'b0 ;
  assign n18642 = n10128 | n18641 ;
  assign n18643 = ( ~n6036 & n8140 ) | ( ~n6036 & n13761 ) | ( n8140 & n13761 ) ;
  assign n18646 = n16832 ^ n5656 ^ 1'b0 ;
  assign n18644 = ~n7133 & n9407 ;
  assign n18645 = n18644 ^ n11605 ^ 1'b0 ;
  assign n18647 = n18646 ^ n18645 ^ n7187 ;
  assign n18648 = n18647 ^ n5729 ^ n3668 ;
  assign n18652 = n5089 & n9395 ;
  assign n18649 = n12225 & n16457 ;
  assign n18650 = x48 & ~n8983 ;
  assign n18651 = ~n18649 & n18650 ;
  assign n18653 = n18652 ^ n18651 ^ n14024 ;
  assign n18654 = n4657 ^ n2051 ^ n1139 ;
  assign n18655 = n3910 ^ n3206 ^ n1945 ;
  assign n18656 = n18655 ^ n14557 ^ n8014 ;
  assign n18657 = n18656 ^ n15330 ^ n1797 ;
  assign n18659 = n13097 ^ n6589 ^ n402 ;
  assign n18658 = ~n4195 & n13847 ;
  assign n18660 = n18659 ^ n18658 ^ 1'b0 ;
  assign n18661 = n6844 & ~n18660 ;
  assign n18662 = n18661 ^ n3454 ^ 1'b0 ;
  assign n18664 = n10909 ^ n5460 ^ n1647 ;
  assign n18665 = ~n1442 & n18664 ;
  assign n18663 = n9405 & n16148 ;
  assign n18666 = n18665 ^ n18663 ^ 1'b0 ;
  assign n18667 = n13468 ^ n5767 ^ 1'b0 ;
  assign n18668 = n9385 | n18667 ;
  assign n18669 = n15534 ^ n14138 ^ n2875 ;
  assign n18670 = ( ~n720 & n7410 ) | ( ~n720 & n9004 ) | ( n7410 & n9004 ) ;
  assign n18671 = n5781 & n7843 ;
  assign n18672 = n1216 & ~n4923 ;
  assign n18673 = ( n4318 & ~n18671 ) | ( n4318 & n18672 ) | ( ~n18671 & n18672 ) ;
  assign n18674 = n1905 & n11786 ;
  assign n18675 = n18674 ^ x15 ^ 1'b0 ;
  assign n18676 = n4112 ^ n3345 ^ n431 ;
  assign n18677 = n18396 & n18676 ;
  assign n18678 = n12222 ^ n8434 ^ 1'b0 ;
  assign n18679 = n12206 & n18678 ;
  assign n18680 = n2741 | n3924 ;
  assign n18681 = ~n4092 & n18680 ;
  assign n18682 = ~n12912 & n18681 ;
  assign n18683 = n3452 & n13018 ;
  assign n18684 = ~n626 & n18683 ;
  assign n18685 = n11691 | n16045 ;
  assign n18686 = n18684 & ~n18685 ;
  assign n18687 = n2429 & n2711 ;
  assign n18690 = n8223 & n10870 ;
  assign n18691 = ( n4146 & n16319 ) | ( n4146 & ~n18690 ) | ( n16319 & ~n18690 ) ;
  assign n18692 = n18691 ^ n18319 ^ n15358 ;
  assign n18688 = n14714 ^ n7687 ^ 1'b0 ;
  assign n18689 = n15655 & ~n18688 ;
  assign n18693 = n18692 ^ n18689 ^ n14451 ;
  assign n18694 = n4574 & ~n13225 ;
  assign n18695 = n18694 ^ n5288 ^ 1'b0 ;
  assign n18699 = ( n3969 & n5681 ) | ( n3969 & n9989 ) | ( n5681 & n9989 ) ;
  assign n18696 = n1775 & n12576 ;
  assign n18697 = ~n11564 & n18696 ;
  assign n18698 = ( n12713 & n15107 ) | ( n12713 & ~n18697 ) | ( n15107 & ~n18697 ) ;
  assign n18700 = n18699 ^ n18698 ^ 1'b0 ;
  assign n18701 = n12577 ^ n3806 ^ 1'b0 ;
  assign n18702 = n18701 ^ n4048 ^ n3180 ;
  assign n18703 = ~n2545 & n8602 ;
  assign n18704 = ~n5915 & n17470 ;
  assign n18705 = n7851 & ~n17278 ;
  assign n18706 = n13247 ^ n5917 ^ 1'b0 ;
  assign n18707 = ( n1424 & n11583 ) | ( n1424 & ~n18706 ) | ( n11583 & ~n18706 ) ;
  assign n18708 = ( n18704 & n18705 ) | ( n18704 & ~n18707 ) | ( n18705 & ~n18707 ) ;
  assign n18709 = ( ~n1929 & n7228 ) | ( ~n1929 & n17802 ) | ( n7228 & n17802 ) ;
  assign n18710 = ( n3573 & n16622 ) | ( n3573 & n18709 ) | ( n16622 & n18709 ) ;
  assign n18714 = n10931 ^ n2181 ^ n1563 ;
  assign n18711 = ( n2119 & n5157 ) | ( n2119 & ~n6726 ) | ( n5157 & ~n6726 ) ;
  assign n18712 = n644 & n5399 ;
  assign n18713 = n18711 & n18712 ;
  assign n18715 = n18714 ^ n18713 ^ 1'b0 ;
  assign n18716 = n11088 ^ n6742 ^ n1419 ;
  assign n18717 = n13228 & n18716 ;
  assign n18718 = ~n179 & n18717 ;
  assign n18719 = n6833 & ~n18105 ;
  assign n18720 = n18719 ^ n13663 ^ 1'b0 ;
  assign n18721 = n18720 ^ n15845 ^ n1529 ;
  assign n18722 = ( ~n11067 & n12914 ) | ( ~n11067 & n16001 ) | ( n12914 & n16001 ) ;
  assign n18723 = n8540 ^ n5442 ^ n4436 ;
  assign n18724 = n5770 ^ n753 ^ 1'b0 ;
  assign n18725 = n18723 & n18724 ;
  assign n18726 = ( n1076 & ~n2281 ) | ( n1076 & n9157 ) | ( ~n2281 & n9157 ) ;
  assign n18727 = ( n10784 & n18725 ) | ( n10784 & ~n18726 ) | ( n18725 & ~n18726 ) ;
  assign n18728 = n7238 & ~n18727 ;
  assign n18729 = n6013 ^ n5934 ^ 1'b0 ;
  assign n18730 = n7298 & n18729 ;
  assign n18731 = n2072 & n7194 ;
  assign n18732 = n12713 & n18731 ;
  assign n18733 = n18732 ^ n6226 ^ 1'b0 ;
  assign n18734 = n3206 | n18733 ;
  assign n18735 = n11754 & ~n18734 ;
  assign n18739 = n9259 & n13816 ;
  assign n18740 = n9996 & n18739 ;
  assign n18741 = n18740 ^ n10991 ^ n4141 ;
  assign n18736 = ( ~n3153 & n3539 ) | ( ~n3153 & n9259 ) | ( n3539 & n9259 ) ;
  assign n18737 = n18736 ^ n11144 ^ n4016 ;
  assign n18738 = n18737 ^ n4925 ^ 1'b0 ;
  assign n18742 = n18741 ^ n18738 ^ n7163 ;
  assign n18743 = n8398 ^ n7907 ^ 1'b0 ;
  assign n18744 = ( ~n1023 & n4347 ) | ( ~n1023 & n10731 ) | ( n4347 & n10731 ) ;
  assign n18745 = ~n5019 & n17185 ;
  assign n18746 = n18745 ^ n18020 ^ 1'b0 ;
  assign n18747 = n8712 ^ n3254 ^ n346 ;
  assign n18748 = n18747 ^ n13700 ^ n5642 ;
  assign n18749 = n9168 ^ n4920 ^ n4658 ;
  assign n18750 = n18749 ^ n11952 ^ n10057 ;
  assign n18753 = n2444 & n5144 ;
  assign n18754 = n18753 ^ n9534 ^ 1'b0 ;
  assign n18755 = n11722 & ~n18754 ;
  assign n18756 = ( n2738 & n14939 ) | ( n2738 & ~n18755 ) | ( n14939 & ~n18755 ) ;
  assign n18751 = n13711 & n13771 ;
  assign n18752 = n2448 & n18751 ;
  assign n18757 = n18756 ^ n18752 ^ n9210 ;
  assign n18763 = ( n454 & n1897 ) | ( n454 & n4024 ) | ( n1897 & n4024 ) ;
  assign n18764 = ( n1583 & n5649 ) | ( n1583 & ~n18763 ) | ( n5649 & ~n18763 ) ;
  assign n18758 = n6101 | n9409 ;
  assign n18759 = n7049 | n18758 ;
  assign n18760 = n6986 | n10313 ;
  assign n18761 = n18760 ^ n4022 ^ 1'b0 ;
  assign n18762 = ( n6582 & n18759 ) | ( n6582 & n18761 ) | ( n18759 & n18761 ) ;
  assign n18765 = n18764 ^ n18762 ^ n4186 ;
  assign n18766 = n7201 & ~n17197 ;
  assign n18767 = n12723 ^ n10631 ^ 1'b0 ;
  assign n18768 = n12969 | n18767 ;
  assign n18769 = n18768 ^ n18659 ^ 1'b0 ;
  assign n18770 = ~n4107 & n18769 ;
  assign n18775 = n8505 ^ n4382 ^ n265 ;
  assign n18776 = n2550 | n18775 ;
  assign n18777 = n10792 & ~n18776 ;
  assign n18778 = ( ~n6723 & n15818 ) | ( ~n6723 & n18777 ) | ( n15818 & n18777 ) ;
  assign n18771 = n14423 ^ n12982 ^ n5948 ;
  assign n18772 = n18771 ^ n935 ^ n547 ;
  assign n18773 = n4345 & n18772 ;
  assign n18774 = n18773 ^ n14633 ^ 1'b0 ;
  assign n18779 = n18778 ^ n18774 ^ n4411 ;
  assign n18780 = n16301 ^ n9674 ^ n6814 ;
  assign n18781 = n6742 ^ n563 ^ 1'b0 ;
  assign n18782 = n1477 | n3711 ;
  assign n18783 = ( n604 & n8322 ) | ( n604 & n18782 ) | ( n8322 & n18782 ) ;
  assign n18784 = n3577 & n10443 ;
  assign n18785 = n18784 ^ n10041 ^ 1'b0 ;
  assign n18786 = n3510 | n8788 ;
  assign n18787 = n16926 ^ n13349 ^ 1'b0 ;
  assign n18788 = n5069 & ~n18787 ;
  assign n18789 = n4367 ^ n3459 ^ 1'b0 ;
  assign n18791 = n10524 ^ n2706 ^ n1086 ;
  assign n18790 = n2707 | n3582 ;
  assign n18792 = n18791 ^ n18790 ^ 1'b0 ;
  assign n18793 = n7594 & n18792 ;
  assign n18794 = ( n8345 & n10396 ) | ( n8345 & n18170 ) | ( n10396 & n18170 ) ;
  assign n18795 = n5054 & n10821 ;
  assign n18796 = n3365 | n18795 ;
  assign n18797 = ( ~n14657 & n17574 ) | ( ~n14657 & n18796 ) | ( n17574 & n18796 ) ;
  assign n18798 = n11842 | n13246 ;
  assign n18799 = n18798 ^ n7594 ^ 1'b0 ;
  assign n18800 = ~n6599 & n7465 ;
  assign n18801 = n18800 ^ n10818 ^ 1'b0 ;
  assign n18802 = n2616 ^ n1523 ^ 1'b0 ;
  assign n18803 = ~n468 & n18802 ;
  assign n18804 = n8015 ^ n3292 ^ n2786 ;
  assign n18805 = n4831 & ~n12089 ;
  assign n18806 = ~x96 & n18805 ;
  assign n18807 = n16451 ^ n7822 ^ 1'b0 ;
  assign n18808 = n14812 & ~n18807 ;
  assign n18809 = ( n12321 & n18806 ) | ( n12321 & n18808 ) | ( n18806 & n18808 ) ;
  assign n18812 = n4906 ^ n3150 ^ n1644 ;
  assign n18813 = ( n3589 & n5563 ) | ( n3589 & n8459 ) | ( n5563 & n8459 ) ;
  assign n18814 = n18813 ^ n4654 ^ n3652 ;
  assign n18815 = n18812 & n18814 ;
  assign n18810 = ( n1452 & ~n12410 ) | ( n1452 & n15847 ) | ( ~n12410 & n15847 ) ;
  assign n18811 = n16390 | n18810 ;
  assign n18816 = n18815 ^ n18811 ^ 1'b0 ;
  assign n18817 = n3169 | n4301 ;
  assign n18818 = n18817 ^ n14198 ^ 1'b0 ;
  assign n18819 = ( n6062 & ~n8261 ) | ( n6062 & n18818 ) | ( ~n8261 & n18818 ) ;
  assign n18820 = n5018 ^ n3810 ^ n2170 ;
  assign n18821 = n18820 ^ n1747 ^ 1'b0 ;
  assign n18822 = ( ~n5805 & n11460 ) | ( ~n5805 & n18821 ) | ( n11460 & n18821 ) ;
  assign n18823 = n3764 | n5813 ;
  assign n18824 = n18823 ^ n17084 ^ n2834 ;
  assign n18825 = n18824 ^ n17780 ^ n9701 ;
  assign n18827 = n5499 & ~n8793 ;
  assign n18826 = n1063 | n9698 ;
  assign n18828 = n18827 ^ n18826 ^ n13212 ;
  assign n18829 = ( n4713 & n5356 ) | ( n4713 & n18828 ) | ( n5356 & n18828 ) ;
  assign n18830 = n1459 & n14339 ;
  assign n18831 = ~n18829 & n18830 ;
  assign n18832 = n13328 ^ n604 ^ 1'b0 ;
  assign n18837 = n8227 | n10569 ;
  assign n18838 = n9144 | n18837 ;
  assign n18836 = n5286 & n13750 ;
  assign n18839 = n18838 ^ n18836 ^ n6127 ;
  assign n18834 = ( n3125 & n4152 ) | ( n3125 & ~n6409 ) | ( n4152 & ~n6409 ) ;
  assign n18833 = n14343 ^ n4695 ^ 1'b0 ;
  assign n18835 = n18834 ^ n18833 ^ n12595 ;
  assign n18840 = n18839 ^ n18835 ^ n633 ;
  assign n18841 = n8788 ^ n4190 ^ 1'b0 ;
  assign n18842 = n18841 ^ n9900 ^ n3428 ;
  assign n18843 = n12103 ^ n7078 ^ 1'b0 ;
  assign n18844 = n18842 & ~n18843 ;
  assign n18845 = ( x51 & n3928 ) | ( x51 & ~n18844 ) | ( n3928 & ~n18844 ) ;
  assign n18846 = n4443 & ~n15522 ;
  assign n18847 = ( ~n6517 & n7809 ) | ( ~n6517 & n9079 ) | ( n7809 & n9079 ) ;
  assign n18848 = n15107 ^ n6954 ^ n5767 ;
  assign n18849 = ( n18846 & n18847 ) | ( n18846 & n18848 ) | ( n18847 & n18848 ) ;
  assign n18850 = n2555 | n5239 ;
  assign n18851 = n8734 | n18850 ;
  assign n18852 = n6444 & ~n18851 ;
  assign n18853 = ( n4973 & ~n15675 ) | ( n4973 & n18852 ) | ( ~n15675 & n18852 ) ;
  assign n18854 = n18853 ^ n10157 ^ n8429 ;
  assign n18855 = ( x56 & ~n15620 ) | ( x56 & n16288 ) | ( ~n15620 & n16288 ) ;
  assign n18856 = n7274 ^ n912 ^ 1'b0 ;
  assign n18857 = n5369 & ~n18856 ;
  assign n18858 = n13259 & n18857 ;
  assign n18859 = ( ~n1086 & n10890 ) | ( ~n1086 & n18858 ) | ( n10890 & n18858 ) ;
  assign n18860 = n15796 ^ n7794 ^ n5142 ;
  assign n18862 = n10342 ^ n7712 ^ 1'b0 ;
  assign n18861 = n2259 ^ n1654 ^ n374 ;
  assign n18863 = n18862 ^ n18861 ^ n4914 ;
  assign n18864 = n5504 ^ n2381 ^ n1285 ;
  assign n18865 = n6482 & ~n18864 ;
  assign n18866 = n12762 ^ n8087 ^ 1'b0 ;
  assign n18867 = n683 & n18866 ;
  assign n18868 = ( n1409 & n1965 ) | ( n1409 & ~n18867 ) | ( n1965 & ~n18867 ) ;
  assign n18869 = ~n18865 & n18868 ;
  assign n18870 = ~n12320 & n17087 ;
  assign n18871 = ( ~n18045 & n18869 ) | ( ~n18045 & n18870 ) | ( n18869 & n18870 ) ;
  assign n18872 = n16067 ^ n12585 ^ n11988 ;
  assign n18873 = n18872 ^ n11221 ^ n7270 ;
  assign n18875 = n7687 ^ n4975 ^ 1'b0 ;
  assign n18876 = n7187 & ~n18875 ;
  assign n18874 = n15129 & ~n17965 ;
  assign n18877 = n18876 ^ n18874 ^ n18337 ;
  assign n18878 = n4010 & n6961 ;
  assign n18879 = n11687 & n18878 ;
  assign n18880 = ( ~n4267 & n7183 ) | ( ~n4267 & n11811 ) | ( n7183 & n11811 ) ;
  assign n18881 = n18880 ^ n8153 ^ n2038 ;
  assign n18882 = n14725 ^ n7192 ^ n5068 ;
  assign n18883 = ( ~n5162 & n14590 ) | ( ~n5162 & n18882 ) | ( n14590 & n18882 ) ;
  assign n18884 = ( ~n2026 & n6984 ) | ( ~n2026 & n18883 ) | ( n6984 & n18883 ) ;
  assign n18885 = n16961 ^ n10195 ^ n950 ;
  assign n18892 = n9167 ^ n2692 ^ 1'b0 ;
  assign n18887 = n11330 ^ n1450 ^ 1'b0 ;
  assign n18888 = n3856 & ~n18887 ;
  assign n18889 = n955 & ~n18888 ;
  assign n18890 = n18889 ^ n388 ^ 1'b0 ;
  assign n18886 = n1523 & ~n5519 ;
  assign n18891 = n18890 ^ n18886 ^ 1'b0 ;
  assign n18893 = n18892 ^ n18891 ^ 1'b0 ;
  assign n18894 = n18095 | n18893 ;
  assign n18895 = n544 | n1970 ;
  assign n18896 = ~n1283 & n18895 ;
  assign n18897 = ( n5258 & n6624 ) | ( n5258 & ~n15959 ) | ( n6624 & ~n15959 ) ;
  assign n18898 = n18085 | n18897 ;
  assign n18899 = n18898 ^ n3602 ^ 1'b0 ;
  assign n18900 = n8623 ^ n1330 ^ n529 ;
  assign n18902 = n1583 & n1737 ;
  assign n18901 = n13650 ^ n11894 ^ n5665 ;
  assign n18903 = n18902 ^ n18901 ^ n5648 ;
  assign n18904 = n6079 & n18903 ;
  assign n18905 = n18904 ^ n8511 ^ 1'b0 ;
  assign n18906 = ( n4982 & n18900 ) | ( n4982 & ~n18905 ) | ( n18900 & ~n18905 ) ;
  assign n18907 = n1242 ^ n602 ^ 1'b0 ;
  assign n18908 = ( ~n4295 & n5229 ) | ( ~n4295 & n6475 ) | ( n5229 & n6475 ) ;
  assign n18909 = ( n1707 & n12136 ) | ( n1707 & n18908 ) | ( n12136 & n18908 ) ;
  assign n18910 = ( ~n14715 & n18907 ) | ( ~n14715 & n18909 ) | ( n18907 & n18909 ) ;
  assign n18911 = n2787 ^ n1856 ^ 1'b0 ;
  assign n18912 = ~n18167 & n18911 ;
  assign n18913 = n5977 ^ n3953 ^ n3138 ;
  assign n18914 = ( ~n2170 & n18912 ) | ( ~n2170 & n18913 ) | ( n18912 & n18913 ) ;
  assign n18915 = n10485 ^ n2165 ^ 1'b0 ;
  assign n18916 = ~n8356 & n18915 ;
  assign n18917 = ( n522 & ~n7241 ) | ( n522 & n18474 ) | ( ~n7241 & n18474 ) ;
  assign n18918 = n2055 ^ n1902 ^ 1'b0 ;
  assign n18919 = n15952 & ~n18918 ;
  assign n18920 = n18919 ^ n6002 ^ n5864 ;
  assign n18921 = ( ~n17404 & n18917 ) | ( ~n17404 & n18920 ) | ( n18917 & n18920 ) ;
  assign n18922 = n18921 ^ n8896 ^ n6483 ;
  assign n18923 = n14821 ^ n10601 ^ 1'b0 ;
  assign n18924 = n18494 & ~n18923 ;
  assign n18925 = ( n18204 & n18783 ) | ( n18204 & n18924 ) | ( n18783 & n18924 ) ;
  assign n18926 = ( n1471 & n12882 ) | ( n1471 & ~n13895 ) | ( n12882 & ~n13895 ) ;
  assign n18927 = n15294 ^ n5894 ^ n5577 ;
  assign n18928 = n9863 | n18462 ;
  assign n18929 = n18928 ^ n315 ^ 1'b0 ;
  assign n18930 = n295 & n5060 ;
  assign n18931 = n18930 ^ n2089 ^ 1'b0 ;
  assign n18940 = n5401 & n7035 ;
  assign n18933 = n402 | n2275 ;
  assign n18934 = n18933 ^ n8431 ^ 1'b0 ;
  assign n18935 = n8915 | n18934 ;
  assign n18936 = n17365 & ~n18935 ;
  assign n18932 = n6424 ^ n2589 ^ 1'b0 ;
  assign n18937 = n18936 ^ n18932 ^ 1'b0 ;
  assign n18938 = n18937 ^ n7729 ^ 1'b0 ;
  assign n18939 = ~n18736 & n18938 ;
  assign n18941 = n18940 ^ n18939 ^ 1'b0 ;
  assign n18942 = n12978 ^ n12064 ^ 1'b0 ;
  assign n18943 = ~n1024 & n3191 ;
  assign n18944 = n2010 & n18943 ;
  assign n18945 = n6050 & n18944 ;
  assign n18946 = n3415 & n18747 ;
  assign n18947 = ~n18945 & n18946 ;
  assign n18948 = n8071 ^ n7876 ^ 1'b0 ;
  assign n18949 = n18948 ^ n12210 ^ 1'b0 ;
  assign n18950 = ~n11712 & n18949 ;
  assign n18951 = n15287 ^ n3896 ^ 1'b0 ;
  assign n18952 = ( n9126 & n14643 ) | ( n9126 & n15107 ) | ( n14643 & n15107 ) ;
  assign n18953 = ~n3631 & n18952 ;
  assign n18954 = ~n7843 & n18953 ;
  assign n18955 = ( n2546 & ~n5395 ) | ( n2546 & n7668 ) | ( ~n5395 & n7668 ) ;
  assign n18956 = ~n7867 & n18955 ;
  assign n18957 = ( n6712 & n9738 ) | ( n6712 & n18956 ) | ( n9738 & n18956 ) ;
  assign n18958 = n2405 & ~n17815 ;
  assign n18959 = ( n1711 & n6335 ) | ( n1711 & ~n18958 ) | ( n6335 & ~n18958 ) ;
  assign n18962 = n18944 ^ n3274 ^ n271 ;
  assign n18960 = n6110 ^ n3704 ^ 1'b0 ;
  assign n18961 = n4312 | n18960 ;
  assign n18963 = n18962 ^ n18961 ^ n7025 ;
  assign n18966 = n4077 ^ n3661 ^ n830 ;
  assign n18967 = ( n1336 & ~n3506 ) | ( n1336 & n18966 ) | ( ~n3506 & n18966 ) ;
  assign n18964 = n3016 ^ n1654 ^ 1'b0 ;
  assign n18965 = n8444 & ~n18964 ;
  assign n18968 = n18967 ^ n18965 ^ 1'b0 ;
  assign n18969 = ( n988 & n6796 ) | ( n988 & n7375 ) | ( n6796 & n7375 ) ;
  assign n18970 = ~n6174 & n6283 ;
  assign n18971 = n18970 ^ n7882 ^ 1'b0 ;
  assign n18972 = n18971 ^ n11519 ^ n6276 ;
  assign n18973 = n14956 ^ n2055 ^ 1'b0 ;
  assign n18974 = n18427 ^ n11811 ^ n449 ;
  assign n18975 = ( n2721 & n3411 ) | ( n2721 & ~n7373 ) | ( n3411 & ~n7373 ) ;
  assign n18976 = n18975 ^ n7512 ^ 1'b0 ;
  assign n18977 = ( x16 & n7907 ) | ( x16 & ~n14705 ) | ( n7907 & ~n14705 ) ;
  assign n18978 = n17339 ^ n6786 ^ 1'b0 ;
  assign n18979 = n3029 | n18978 ;
  assign n18980 = n2688 ^ n822 ^ 1'b0 ;
  assign n18981 = n11988 ^ n3932 ^ 1'b0 ;
  assign n18982 = n18981 ^ n9015 ^ n376 ;
  assign n18983 = ~n849 & n7670 ;
  assign n18984 = n18983 ^ n4522 ^ 1'b0 ;
  assign n18985 = ( n7528 & ~n14801 ) | ( n7528 & n18984 ) | ( ~n14801 & n18984 ) ;
  assign n18986 = n7169 ^ n2913 ^ 1'b0 ;
  assign n18987 = n3831 | n18986 ;
  assign n18988 = n11718 ^ n7926 ^ 1'b0 ;
  assign n18989 = n12474 & n18988 ;
  assign n18990 = n3628 & ~n18989 ;
  assign n18991 = n3360 | n12547 ;
  assign n18992 = n18991 ^ n13789 ^ 1'b0 ;
  assign n18993 = n18992 ^ n12587 ^ 1'b0 ;
  assign n18994 = n10826 ^ n9634 ^ n4993 ;
  assign n18995 = ( n13922 & n17848 ) | ( n13922 & ~n18994 ) | ( n17848 & ~n18994 ) ;
  assign n18996 = n18995 ^ n15576 ^ n4843 ;
  assign n18997 = n5681 & ~n8288 ;
  assign n18998 = n18997 ^ n6875 ^ 1'b0 ;
  assign n18999 = n2656 & ~n18998 ;
  assign n19000 = n17718 & n18999 ;
  assign n19001 = n18856 ^ n3339 ^ n1032 ;
  assign n19002 = n4226 | n12161 ;
  assign n19003 = n19001 & ~n19002 ;
  assign n19004 = n19003 ^ n18486 ^ n6860 ;
  assign n19006 = n364 & n792 ;
  assign n19005 = n12569 ^ n11102 ^ n3934 ;
  assign n19007 = n19006 ^ n19005 ^ 1'b0 ;
  assign n19008 = n10754 & ~n13131 ;
  assign n19009 = n7226 | n11587 ;
  assign n19010 = ( n2377 & n7785 ) | ( n2377 & ~n14698 ) | ( n7785 & ~n14698 ) ;
  assign n19011 = n19010 ^ n7011 ^ 1'b0 ;
  assign n19012 = n348 & ~n4943 ;
  assign n19013 = n19012 ^ n11062 ^ 1'b0 ;
  assign n19014 = n5210 | n19013 ;
  assign n19015 = n10005 & ~n11488 ;
  assign n19016 = ( n1946 & n6189 ) | ( n1946 & ~n6594 ) | ( n6189 & ~n6594 ) ;
  assign n19017 = n5847 & ~n19016 ;
  assign n19018 = ~n8167 & n19017 ;
  assign n19020 = n3743 & ~n4707 ;
  assign n19021 = ~n4344 & n19020 ;
  assign n19019 = n8380 ^ n2859 ^ 1'b0 ;
  assign n19022 = n19021 ^ n19019 ^ n352 ;
  assign n19023 = n11823 & n19022 ;
  assign n19024 = n19023 ^ n15310 ^ 1'b0 ;
  assign n19025 = ~n10759 & n13703 ;
  assign n19026 = n12476 & n19025 ;
  assign n19027 = ( n3940 & n9195 ) | ( n3940 & ~n19026 ) | ( n9195 & ~n19026 ) ;
  assign n19028 = ( n13447 & ~n19024 ) | ( n13447 & n19027 ) | ( ~n19024 & n19027 ) ;
  assign n19030 = n12402 ^ n7970 ^ n2342 ;
  assign n19031 = n457 & ~n8262 ;
  assign n19032 = ~n19030 & n19031 ;
  assign n19029 = n3540 ^ n1291 ^ 1'b0 ;
  assign n19033 = n19032 ^ n19029 ^ n10270 ;
  assign n19034 = ( n3654 & ~n9177 ) | ( n3654 & n18045 ) | ( ~n9177 & n18045 ) ;
  assign n19046 = ~n4190 & n7518 ;
  assign n19040 = n13589 ^ n9016 ^ n2703 ;
  assign n19041 = n6544 & ~n7836 ;
  assign n19042 = ~n4793 & n19041 ;
  assign n19043 = ( n3733 & n10176 ) | ( n3733 & n19042 ) | ( n10176 & n19042 ) ;
  assign n19044 = n16448 ^ n12000 ^ n10434 ;
  assign n19045 = ( n19040 & ~n19043 ) | ( n19040 & n19044 ) | ( ~n19043 & n19044 ) ;
  assign n19038 = n9611 & ~n13875 ;
  assign n19036 = n5285 ^ n3122 ^ 1'b0 ;
  assign n19035 = n18039 ^ n12541 ^ 1'b0 ;
  assign n19037 = n19036 ^ n19035 ^ n5053 ;
  assign n19039 = n19038 ^ n19037 ^ n4654 ;
  assign n19047 = n19046 ^ n19045 ^ n19039 ;
  assign n19048 = n18504 ^ n13779 ^ 1'b0 ;
  assign n19049 = n12612 & n19048 ;
  assign n19050 = n8521 ^ n1069 ^ n315 ;
  assign n19051 = n8660 ^ n7035 ^ 1'b0 ;
  assign n19052 = n19050 | n19051 ;
  assign n19053 = n19052 ^ n11585 ^ n10930 ;
  assign n19054 = n13648 ^ n360 ^ 1'b0 ;
  assign n19055 = ( n5598 & ~n10317 ) | ( n5598 & n14866 ) | ( ~n10317 & n14866 ) ;
  assign n19056 = ~n19054 & n19055 ;
  assign n19057 = ~n9053 & n10183 ;
  assign n19058 = n19057 ^ n7213 ^ n3665 ;
  assign n19059 = n7859 & ~n8898 ;
  assign n19060 = n5871 & n19059 ;
  assign n19061 = n15974 | n19060 ;
  assign n19062 = n10915 & ~n19061 ;
  assign n19063 = n8597 ^ n4036 ^ n3706 ;
  assign n19064 = ( n1330 & n3807 ) | ( n1330 & n4632 ) | ( n3807 & n4632 ) ;
  assign n19065 = n19064 ^ n17306 ^ n10723 ;
  assign n19066 = ( n4150 & n12691 ) | ( n4150 & ~n19065 ) | ( n12691 & ~n19065 ) ;
  assign n19067 = n19063 & ~n19066 ;
  assign n19068 = n18348 ^ n13048 ^ n2370 ;
  assign n19069 = n11346 ^ n7606 ^ 1'b0 ;
  assign n19070 = ( n11743 & n19068 ) | ( n11743 & n19069 ) | ( n19068 & n19069 ) ;
  assign n19071 = ( n2960 & ~n4149 ) | ( n2960 & n5295 ) | ( ~n4149 & n5295 ) ;
  assign n19072 = n2489 | n19071 ;
  assign n19073 = n2674 | n19072 ;
  assign n19074 = n19073 ^ n894 ^ 1'b0 ;
  assign n19075 = n18770 & ~n18937 ;
  assign n19076 = n7397 & n19075 ;
  assign n19077 = n12452 ^ n11159 ^ 1'b0 ;
  assign n19078 = n1587 & n14092 ;
  assign n19079 = n8403 | n19078 ;
  assign n19080 = n10815 & ~n19079 ;
  assign n19081 = n13991 ^ n9624 ^ 1'b0 ;
  assign n19082 = n19081 ^ n3205 ^ n1837 ;
  assign n19083 = n9028 | n15796 ;
  assign n19084 = n4114 & n4575 ;
  assign n19085 = n2091 & n5154 ;
  assign n19086 = n12093 & ~n14893 ;
  assign n19087 = n5604 ^ n2834 ^ 1'b0 ;
  assign n19088 = ~n18413 & n19087 ;
  assign n19092 = n4310 & ~n4351 ;
  assign n19089 = n201 & n6959 ;
  assign n19090 = n3900 ^ n3151 ^ n2587 ;
  assign n19091 = n19089 & n19090 ;
  assign n19093 = n19092 ^ n19091 ^ n11968 ;
  assign n19094 = n4951 ^ n151 ^ 1'b0 ;
  assign n19095 = n16574 ^ n15354 ^ n4475 ;
  assign n19096 = n18367 ^ n16036 ^ n15618 ;
  assign n19097 = ( n19094 & n19095 ) | ( n19094 & n19096 ) | ( n19095 & n19096 ) ;
  assign n19098 = n14335 ^ n9262 ^ 1'b0 ;
  assign n19099 = n8437 & ~n19098 ;
  assign n19100 = n19099 ^ n1577 ^ n149 ;
  assign n19101 = n18039 ^ n12730 ^ n505 ;
  assign n19102 = n19043 ^ n4500 ^ 1'b0 ;
  assign n19103 = n16362 & ~n18062 ;
  assign n19104 = n19103 ^ n888 ^ 1'b0 ;
  assign n19105 = n19104 ^ n17564 ^ 1'b0 ;
  assign n19106 = n17950 ^ n11720 ^ 1'b0 ;
  assign n19107 = n16590 | n17691 ;
  assign n19108 = n16048 | n19107 ;
  assign n19109 = ( n9977 & n10649 ) | ( n9977 & ~n12483 ) | ( n10649 & ~n12483 ) ;
  assign n19113 = n18521 ^ n8395 ^ n2537 ;
  assign n19110 = n9932 ^ n4531 ^ 1'b0 ;
  assign n19111 = ~n6474 & n10214 ;
  assign n19112 = n19110 & n19111 ;
  assign n19114 = n19113 ^ n19112 ^ n8360 ;
  assign n19115 = ~n4492 & n4726 ;
  assign n19116 = n19115 ^ n3720 ^ 1'b0 ;
  assign n19117 = n15690 ^ n12693 ^ 1'b0 ;
  assign n19118 = ( n690 & n7272 ) | ( n690 & n10407 ) | ( n7272 & n10407 ) ;
  assign n19119 = ~n19117 & n19118 ;
  assign n19120 = ~n17777 & n19119 ;
  assign n19121 = n16485 ^ n7102 ^ n5558 ;
  assign n19122 = ( n6415 & n7965 ) | ( n6415 & n15519 ) | ( n7965 & n15519 ) ;
  assign n19123 = n19122 ^ n17615 ^ n17160 ;
  assign n19125 = n2948 & ~n4414 ;
  assign n19124 = n9881 ^ n5236 ^ n3413 ;
  assign n19126 = n19125 ^ n19124 ^ n4761 ;
  assign n19127 = n6709 ^ n4035 ^ 1'b0 ;
  assign n19128 = ~n4581 & n19127 ;
  assign n19129 = n10915 ^ n4567 ^ 1'b0 ;
  assign n19130 = n11122 ^ n8258 ^ n6273 ;
  assign n19131 = n12097 ^ n8334 ^ 1'b0 ;
  assign n19132 = n19130 | n19131 ;
  assign n19133 = ( n3917 & n8531 ) | ( n3917 & n15125 ) | ( n8531 & n15125 ) ;
  assign n19134 = ( n6595 & n7456 ) | ( n6595 & n12049 ) | ( n7456 & n12049 ) ;
  assign n19135 = n19134 ^ n12045 ^ 1'b0 ;
  assign n19136 = n15648 ^ n7901 ^ n4902 ;
  assign n19137 = ( n13326 & ~n19135 ) | ( n13326 & n19136 ) | ( ~n19135 & n19136 ) ;
  assign n19138 = ~n4014 & n14693 ;
  assign n19139 = n19138 ^ n15375 ^ 1'b0 ;
  assign n19140 = n2667 | n4772 ;
  assign n19141 = n19140 ^ n1827 ^ 1'b0 ;
  assign n19142 = n14029 ^ n13251 ^ n5527 ;
  assign n19143 = ( ~n4073 & n14965 ) | ( ~n4073 & n19142 ) | ( n14965 & n19142 ) ;
  assign n19144 = n18287 ^ n4280 ^ n3990 ;
  assign n19145 = n19144 ^ n13333 ^ 1'b0 ;
  assign n19146 = n14063 | n19145 ;
  assign n19147 = ~n17498 & n19146 ;
  assign n19148 = n2169 & n10466 ;
  assign n19149 = n19148 ^ n19026 ^ 1'b0 ;
  assign n19150 = n15775 ^ n11796 ^ 1'b0 ;
  assign n19151 = n13685 & n19150 ;
  assign n19152 = n2357 | n13440 ;
  assign n19153 = ~n6429 & n14505 ;
  assign n19154 = n19153 ^ n15107 ^ 1'b0 ;
  assign n19155 = ( n9607 & n11110 ) | ( n9607 & n15307 ) | ( n11110 & n15307 ) ;
  assign n19156 = ( n11581 & n13792 ) | ( n11581 & ~n19155 ) | ( n13792 & ~n19155 ) ;
  assign n19158 = n3733 ^ n2033 ^ n1507 ;
  assign n19157 = n12916 | n15232 ;
  assign n19159 = n19158 ^ n19157 ^ 1'b0 ;
  assign n19160 = n16919 ^ n3677 ^ n2769 ;
  assign n19161 = ( n2974 & n7645 ) | ( n2974 & n8399 ) | ( n7645 & n8399 ) ;
  assign n19162 = n5230 & ~n19161 ;
  assign n19163 = n19162 ^ n1313 ^ 1'b0 ;
  assign n19169 = n2754 | n12666 ;
  assign n19170 = n7000 & ~n19169 ;
  assign n19168 = ( n1111 & n6783 ) | ( n1111 & n6913 ) | ( n6783 & n6913 ) ;
  assign n19164 = n750 & n1613 ;
  assign n19165 = n19164 ^ n2767 ^ 1'b0 ;
  assign n19166 = n19165 ^ n5536 ^ n4353 ;
  assign n19167 = n19166 ^ n8494 ^ 1'b0 ;
  assign n19171 = n19170 ^ n19168 ^ n19167 ;
  assign n19172 = n5752 | n11811 ;
  assign n19173 = n19172 ^ n3444 ^ 1'b0 ;
  assign n19174 = ~n11691 & n18763 ;
  assign n19176 = n10683 ^ n7660 ^ 1'b0 ;
  assign n19177 = n12750 & n19176 ;
  assign n19175 = n13698 & n18522 ;
  assign n19178 = n19177 ^ n19175 ^ 1'b0 ;
  assign n19179 = n4344 ^ n3284 ^ n695 ;
  assign n19180 = n19179 ^ n12505 ^ n6077 ;
  assign n19181 = n19180 ^ n4614 ^ n1434 ;
  assign n19182 = n905 & ~n19181 ;
  assign n19183 = n19178 & n19182 ;
  assign n19184 = n13253 & n14639 ;
  assign n19185 = ~n12508 & n19184 ;
  assign n19186 = n5772 & n6147 ;
  assign n19187 = n10589 & ~n19186 ;
  assign n19188 = n12207 ^ n1095 ^ 1'b0 ;
  assign n19189 = n18264 ^ n10061 ^ 1'b0 ;
  assign n19190 = n11303 | n17069 ;
  assign n19191 = n7604 & ~n19190 ;
  assign n19192 = ~n2504 & n12164 ;
  assign n19193 = n14292 & n19192 ;
  assign n19194 = n3591 | n17493 ;
  assign n19195 = n19194 ^ n10181 ^ 1'b0 ;
  assign n19196 = ( n966 & n6208 ) | ( n966 & n9270 ) | ( n6208 & n9270 ) ;
  assign n19197 = n19196 ^ n12909 ^ n878 ;
  assign n19198 = ( n2175 & n16102 ) | ( n2175 & ~n19197 ) | ( n16102 & ~n19197 ) ;
  assign n19199 = ( n9363 & ~n17039 ) | ( n9363 & n19198 ) | ( ~n17039 & n19198 ) ;
  assign n19200 = n2288 | n4679 ;
  assign n19201 = n19200 ^ n5478 ^ n3053 ;
  assign n19202 = n12543 ^ n4654 ^ n1534 ;
  assign n19203 = n10668 ^ n9425 ^ 1'b0 ;
  assign n19204 = n1197 & ~n19203 ;
  assign n19205 = n11833 & n19204 ;
  assign n19206 = n19205 ^ n9414 ^ 1'b0 ;
  assign n19207 = ( n2047 & ~n4876 ) | ( n2047 & n6750 ) | ( ~n4876 & n6750 ) ;
  assign n19208 = n19207 ^ n7504 ^ n3482 ;
  assign n19209 = n19208 ^ n7640 ^ 1'b0 ;
  assign n19210 = n15103 ^ n4157 ^ 1'b0 ;
  assign n19211 = ~n3441 & n12224 ;
  assign n19212 = n19211 ^ n3231 ^ 1'b0 ;
  assign n19213 = n19212 ^ n14863 ^ n14323 ;
  assign n19214 = n19213 ^ n1634 ^ 1'b0 ;
  assign n19215 = ~n2488 & n9131 ;
  assign n19216 = ~n1260 & n19215 ;
  assign n19217 = n2214 & ~n9385 ;
  assign n19218 = n19217 ^ n198 ^ 1'b0 ;
  assign n19219 = n1683 | n8138 ;
  assign n19220 = n19219 ^ n760 ^ 1'b0 ;
  assign n19221 = n19220 ^ n4425 ^ n2120 ;
  assign n19222 = ( n3762 & n19218 ) | ( n3762 & n19221 ) | ( n19218 & n19221 ) ;
  assign n19223 = ( n861 & n6487 ) | ( n861 & ~n7934 ) | ( n6487 & ~n7934 ) ;
  assign n19224 = n9102 & ~n14540 ;
  assign n19225 = ~n14832 & n19224 ;
  assign n19226 = n696 & ~n14100 ;
  assign n19227 = ~n4240 & n19226 ;
  assign n19228 = n6990 ^ n5373 ^ n1867 ;
  assign n19229 = n7899 & n19228 ;
  assign n19230 = n19229 ^ n14901 ^ 1'b0 ;
  assign n19231 = ~n9140 & n19230 ;
  assign n19232 = ( ~n8313 & n13709 ) | ( ~n8313 & n15276 ) | ( n13709 & n15276 ) ;
  assign n19233 = ~n8691 & n19232 ;
  assign n19234 = n16687 & n19233 ;
  assign n19235 = n6325 & n6997 ;
  assign n19236 = n7981 | n17174 ;
  assign n19237 = n19235 | n19236 ;
  assign n19241 = ~n5572 & n5914 ;
  assign n19239 = n12268 ^ n5201 ^ n1221 ;
  assign n19240 = n16703 | n19239 ;
  assign n19242 = n19241 ^ n19240 ^ 1'b0 ;
  assign n19238 = n5827 ^ n2548 ^ n302 ;
  assign n19243 = n19242 ^ n19238 ^ 1'b0 ;
  assign n19244 = n14993 & n19243 ;
  assign n19245 = n16035 ^ n4443 ^ n2554 ;
  assign n19246 = n6386 & ~n19245 ;
  assign n19247 = ~n13441 & n19246 ;
  assign n19248 = n4596 & ~n9655 ;
  assign n19249 = n19248 ^ n19016 ^ 1'b0 ;
  assign n19250 = ( n11699 & n13594 ) | ( n11699 & ~n14577 ) | ( n13594 & ~n14577 ) ;
  assign n19251 = ~n2555 & n2922 ;
  assign n19252 = n19251 ^ n11062 ^ 1'b0 ;
  assign n19253 = n19252 ^ n6414 ^ 1'b0 ;
  assign n19254 = n15147 & ~n19253 ;
  assign n19255 = n19254 ^ n9144 ^ n6824 ;
  assign n19256 = n6391 ^ n901 ^ n565 ;
  assign n19257 = ( n2258 & n18190 ) | ( n2258 & n19256 ) | ( n18190 & n19256 ) ;
  assign n19258 = ( n4647 & ~n9405 ) | ( n4647 & n13938 ) | ( ~n9405 & n13938 ) ;
  assign n19259 = n5545 & ~n7156 ;
  assign n19260 = n10564 ^ n4414 ^ 1'b0 ;
  assign n19261 = ~n6370 & n19260 ;
  assign n19262 = n12301 ^ n11693 ^ 1'b0 ;
  assign n19263 = n19261 & n19262 ;
  assign n19264 = ( ~n4461 & n15913 ) | ( ~n4461 & n18948 ) | ( n15913 & n18948 ) ;
  assign n19265 = n684 & ~n10840 ;
  assign n19266 = n2883 & n19265 ;
  assign n19267 = n6483 | n19266 ;
  assign n19268 = n19264 & ~n19267 ;
  assign n19269 = n10463 & ~n19268 ;
  assign n19270 = n17093 & n19269 ;
  assign n19271 = n580 | n6793 ;
  assign n19272 = n15620 ^ n4593 ^ 1'b0 ;
  assign n19273 = n19271 & n19272 ;
  assign n19274 = n8128 & n19273 ;
  assign n19275 = n19274 ^ n9134 ^ 1'b0 ;
  assign n19276 = n4315 ^ n1901 ^ 1'b0 ;
  assign n19277 = n19276 ^ n9327 ^ 1'b0 ;
  assign n19278 = n19277 ^ n6349 ^ 1'b0 ;
  assign n19279 = ~n14116 & n19278 ;
  assign n19280 = n12890 ^ n12793 ^ 1'b0 ;
  assign n19281 = n11033 & n19280 ;
  assign n19282 = ( n1795 & n19279 ) | ( n1795 & ~n19281 ) | ( n19279 & ~n19281 ) ;
  assign n19287 = n12927 ^ n4070 ^ 1'b0 ;
  assign n19283 = n7816 ^ n5252 ^ n3358 ;
  assign n19284 = n8125 | n19283 ;
  assign n19285 = n19284 ^ n3419 ^ 1'b0 ;
  assign n19286 = ( n9286 & n9639 ) | ( n9286 & ~n19285 ) | ( n9639 & ~n19285 ) ;
  assign n19288 = n19287 ^ n19286 ^ n7002 ;
  assign n19289 = ( ~n2909 & n6698 ) | ( ~n2909 & n8119 ) | ( n6698 & n8119 ) ;
  assign n19290 = n4306 | n17162 ;
  assign n19291 = n19290 ^ n4626 ^ n1182 ;
  assign n19292 = n372 & n4428 ;
  assign n19293 = n19292 ^ n7510 ^ 1'b0 ;
  assign n19298 = n4544 | n13366 ;
  assign n19297 = n7108 | n8672 ;
  assign n19299 = n19298 ^ n19297 ^ 1'b0 ;
  assign n19294 = n18563 ^ n6900 ^ 1'b0 ;
  assign n19295 = n3414 | n19294 ;
  assign n19296 = n10099 & ~n19295 ;
  assign n19300 = n19299 ^ n19296 ^ 1'b0 ;
  assign n19301 = n5096 | n9695 ;
  assign n19302 = ( n4028 & n5352 ) | ( n4028 & n9823 ) | ( n5352 & n9823 ) ;
  assign n19303 = n9158 ^ n260 ^ 1'b0 ;
  assign n19304 = n19302 & n19303 ;
  assign n19305 = ~n11738 & n19304 ;
  assign n19306 = ~n13020 & n19305 ;
  assign n19307 = n19306 ^ n16233 ^ n11804 ;
  assign n19308 = ~n7777 & n19307 ;
  assign n19309 = n19308 ^ n10519 ^ 1'b0 ;
  assign n19310 = ( n1074 & n1104 ) | ( n1074 & ~n17345 ) | ( n1104 & ~n17345 ) ;
  assign n19311 = ~n9795 & n16588 ;
  assign n19312 = x74 & n2318 ;
  assign n19313 = ~x74 & n19312 ;
  assign n19314 = ( n1127 & n8811 ) | ( n1127 & ~n19313 ) | ( n8811 & ~n19313 ) ;
  assign n19318 = n14858 ^ n4065 ^ 1'b0 ;
  assign n19316 = n7052 ^ n4335 ^ 1'b0 ;
  assign n19317 = ( n6445 & n11299 ) | ( n6445 & ~n19316 ) | ( n11299 & ~n19316 ) ;
  assign n19315 = ( ~n5356 & n7245 ) | ( ~n5356 & n14684 ) | ( n7245 & n14684 ) ;
  assign n19319 = n19318 ^ n19317 ^ n19315 ;
  assign n19320 = n19319 ^ n14347 ^ 1'b0 ;
  assign n19321 = n19314 & ~n19320 ;
  assign n19322 = ~n9347 & n12136 ;
  assign n19323 = n14977 ^ n13747 ^ 1'b0 ;
  assign n19324 = n11508 ^ n6937 ^ n5531 ;
  assign n19325 = n6364 & n14446 ;
  assign n19326 = n15888 & n19325 ;
  assign n19327 = n13121 | n14078 ;
  assign n19328 = n14455 | n19327 ;
  assign n19329 = n15888 & ~n18275 ;
  assign n19330 = n15222 ^ n10986 ^ 1'b0 ;
  assign n19331 = ~n3214 & n19330 ;
  assign n19332 = ( n10111 & ~n13616 ) | ( n10111 & n16699 ) | ( ~n13616 & n16699 ) ;
  assign n19334 = ( x63 & n4568 ) | ( x63 & n12911 ) | ( n4568 & n12911 ) ;
  assign n19333 = n11084 ^ n6877 ^ n6831 ;
  assign n19335 = n19334 ^ n19333 ^ n13959 ;
  assign n19336 = n1616 | n11540 ;
  assign n19337 = n19336 ^ n4163 ^ 1'b0 ;
  assign n19338 = n19337 ^ n7500 ^ n2065 ;
  assign n19339 = ( n1917 & n7781 ) | ( n1917 & ~n19338 ) | ( n7781 & ~n19338 ) ;
  assign n19340 = n11528 ^ n10879 ^ n3148 ;
  assign n19341 = n18913 ^ n11321 ^ n4648 ;
  assign n19342 = ( n2642 & n12648 ) | ( n2642 & n18749 ) | ( n12648 & n18749 ) ;
  assign n19343 = n5220 ^ n4568 ^ n1748 ;
  assign n19344 = n816 & ~n19343 ;
  assign n19345 = n18043 ^ n5144 ^ n2807 ;
  assign n19353 = n11991 ^ n6850 ^ n4550 ;
  assign n19354 = ( ~n5397 & n14963 ) | ( ~n5397 & n19353 ) | ( n14963 & n19353 ) ;
  assign n19350 = n14549 ^ n6729 ^ 1'b0 ;
  assign n19351 = n19350 ^ n15330 ^ 1'b0 ;
  assign n19347 = x63 | n3123 ;
  assign n19348 = n19347 ^ n15713 ^ 1'b0 ;
  assign n19349 = n19348 ^ n18232 ^ n206 ;
  assign n19346 = n2642 | n7381 ;
  assign n19352 = n19351 ^ n19349 ^ n19346 ;
  assign n19355 = n19354 ^ n19352 ^ n15311 ;
  assign n19356 = n18480 ^ n10437 ^ 1'b0 ;
  assign n19357 = n9744 & n19356 ;
  assign n19358 = ~n19355 & n19357 ;
  assign n19359 = n10584 | n13149 ;
  assign n19360 = n4537 & ~n19359 ;
  assign n19361 = ~n410 & n522 ;
  assign n19362 = n11555 ^ n6937 ^ 1'b0 ;
  assign n19363 = ( n1118 & n15923 ) | ( n1118 & n19362 ) | ( n15923 & n19362 ) ;
  assign n19364 = n18680 ^ n10494 ^ 1'b0 ;
  assign n19365 = n19038 ^ n2293 ^ 1'b0 ;
  assign n19366 = n13860 ^ n10232 ^ n8128 ;
  assign n19367 = n11479 & n18891 ;
  assign n19368 = ~n2580 & n19367 ;
  assign n19369 = n1414 | n4168 ;
  assign n19370 = n19369 ^ n3453 ^ 1'b0 ;
  assign n19372 = n2733 ^ n2462 ^ 1'b0 ;
  assign n19373 = ~n8010 & n19372 ;
  assign n19374 = ~n12852 & n19373 ;
  assign n19371 = ~n4383 & n13366 ;
  assign n19375 = n19374 ^ n19371 ^ 1'b0 ;
  assign n19376 = ( n2976 & n15774 ) | ( n2976 & ~n19375 ) | ( n15774 & ~n19375 ) ;
  assign n19379 = ( ~n2916 & n3105 ) | ( ~n2916 & n8583 ) | ( n3105 & n8583 ) ;
  assign n19380 = n5483 ^ n2418 ^ 1'b0 ;
  assign n19381 = ~n12829 & n19380 ;
  assign n19382 = ( n8037 & n12251 ) | ( n8037 & n19381 ) | ( n12251 & n19381 ) ;
  assign n19383 = ~n4696 & n16744 ;
  assign n19384 = ( n19379 & n19382 ) | ( n19379 & n19383 ) | ( n19382 & n19383 ) ;
  assign n19377 = n2789 | n14567 ;
  assign n19378 = n19377 ^ n16780 ^ 1'b0 ;
  assign n19385 = n19384 ^ n19378 ^ n11435 ;
  assign n19386 = n11994 ^ n3579 ^ 1'b0 ;
  assign n19387 = n19386 ^ n9591 ^ n1396 ;
  assign n19388 = ~n12690 & n19387 ;
  assign n19389 = n7032 ^ n2694 ^ 1'b0 ;
  assign n19390 = ~n6740 & n19389 ;
  assign n19391 = n18756 ^ n2554 ^ 1'b0 ;
  assign n19392 = ~n6723 & n15807 ;
  assign n19393 = n7456 & n19392 ;
  assign n19394 = n19393 ^ n9553 ^ n4657 ;
  assign n19395 = n1681 & ~n3422 ;
  assign n19396 = n19394 & n19395 ;
  assign n19397 = n4839 ^ n3595 ^ 1'b0 ;
  assign n19398 = n1295 | n6487 ;
  assign n19399 = n19398 ^ n13288 ^ n9286 ;
  assign n19402 = x37 & n324 ;
  assign n19403 = n19402 ^ n1290 ^ 1'b0 ;
  assign n19404 = n7613 ^ n2511 ^ 1'b0 ;
  assign n19405 = n19403 & ~n19404 ;
  assign n19400 = ( ~x59 & n5754 ) | ( ~x59 & n10421 ) | ( n5754 & n10421 ) ;
  assign n19401 = n8708 & n19400 ;
  assign n19406 = n19405 ^ n19401 ^ 1'b0 ;
  assign n19407 = n19406 ^ n19024 ^ n4983 ;
  assign n19408 = n14563 ^ n7755 ^ n3991 ;
  assign n19409 = n626 & ~n1010 ;
  assign n19410 = n19409 ^ n1023 ^ 1'b0 ;
  assign n19411 = n19410 ^ n13991 ^ 1'b0 ;
  assign n19412 = ~n9761 & n19411 ;
  assign n19419 = n10010 ^ n3129 ^ 1'b0 ;
  assign n19420 = n16994 | n19419 ;
  assign n19415 = ~n1662 & n3665 ;
  assign n19416 = n562 & n19415 ;
  assign n19417 = n19416 ^ n8023 ^ x72 ;
  assign n19413 = x76 & n17497 ;
  assign n19414 = ~n3189 & n19413 ;
  assign n19418 = n19417 ^ n19414 ^ 1'b0 ;
  assign n19421 = n19420 ^ n19418 ^ n4469 ;
  assign n19422 = ( n2785 & n12817 ) | ( n2785 & ~n19421 ) | ( n12817 & ~n19421 ) ;
  assign n19426 = n7639 ^ x75 ^ 1'b0 ;
  assign n19427 = ( n1742 & ~n7601 ) | ( n1742 & n19426 ) | ( ~n7601 & n19426 ) ;
  assign n19425 = ( n2040 & n6335 ) | ( n2040 & ~n16545 ) | ( n6335 & ~n16545 ) ;
  assign n19423 = ( ~n4402 & n5566 ) | ( ~n4402 & n16651 ) | ( n5566 & n16651 ) ;
  assign n19424 = ( n5266 & ~n11287 ) | ( n5266 & n19423 ) | ( ~n11287 & n19423 ) ;
  assign n19428 = n19427 ^ n19425 ^ n19424 ;
  assign n19429 = ~n1356 & n2338 ;
  assign n19430 = n14721 & ~n19429 ;
  assign n19434 = n8182 ^ n2342 ^ 1'b0 ;
  assign n19431 = n1797 | n10386 ;
  assign n19432 = n13752 | n19431 ;
  assign n19433 = n13248 & n19432 ;
  assign n19435 = n19434 ^ n19433 ^ 1'b0 ;
  assign n19436 = n10413 ^ n9998 ^ 1'b0 ;
  assign n19437 = ~n9409 & n9998 ;
  assign n19438 = ~n19436 & n19437 ;
  assign n19439 = ( ~n5076 & n9770 ) | ( ~n5076 & n18006 ) | ( n9770 & n18006 ) ;
  assign n19440 = ( n6331 & ~n12907 ) | ( n6331 & n19439 ) | ( ~n12907 & n19439 ) ;
  assign n19441 = n9838 ^ n8507 ^ 1'b0 ;
  assign n19442 = n6287 | n19441 ;
  assign n19443 = n7185 | n19442 ;
  assign n19444 = n19443 ^ n7274 ^ n7080 ;
  assign n19445 = ~n1879 & n16455 ;
  assign n19446 = n3766 & n14627 ;
  assign n19447 = n19446 ^ n12914 ^ 1'b0 ;
  assign n19448 = n9016 ^ n6226 ^ n3541 ;
  assign n19449 = ( ~n4543 & n8985 ) | ( ~n4543 & n19448 ) | ( n8985 & n19448 ) ;
  assign n19450 = ~n2326 & n19449 ;
  assign n19451 = ~n14043 & n19450 ;
  assign n19452 = n12849 | n19451 ;
  assign n19453 = n19452 ^ n3770 ^ 1'b0 ;
  assign n19454 = ( n1169 & n1611 ) | ( n1169 & ~n4879 ) | ( n1611 & ~n4879 ) ;
  assign n19455 = n2803 & ~n6673 ;
  assign n19456 = ~n4004 & n19455 ;
  assign n19457 = ( ~n3667 & n13267 ) | ( ~n3667 & n19456 ) | ( n13267 & n19456 ) ;
  assign n19458 = n19457 ^ n7450 ^ n6195 ;
  assign n19459 = n19458 ^ n17819 ^ n10367 ;
  assign n19460 = ( ~n19185 & n19454 ) | ( ~n19185 & n19459 ) | ( n19454 & n19459 ) ;
  assign n19461 = ( n568 & n7078 ) | ( n568 & ~n8406 ) | ( n7078 & ~n8406 ) ;
  assign n19462 = ( ~n741 & n1729 ) | ( ~n741 & n7660 ) | ( n1729 & n7660 ) ;
  assign n19463 = ( n6634 & ~n16506 ) | ( n6634 & n19462 ) | ( ~n16506 & n19462 ) ;
  assign n19464 = n19461 & ~n19463 ;
  assign n19465 = ~n8216 & n9259 ;
  assign n19466 = n2563 | n3307 ;
  assign n19467 = n19466 ^ n1913 ^ 1'b0 ;
  assign n19468 = n12885 ^ n2625 ^ 1'b0 ;
  assign n19469 = ( n12206 & n13688 ) | ( n12206 & n19468 ) | ( n13688 & n19468 ) ;
  assign n19470 = n3144 & n6899 ;
  assign n19471 = ( n3583 & n8543 ) | ( n3583 & ~n19470 ) | ( n8543 & ~n19470 ) ;
  assign n19472 = n19471 ^ n10309 ^ 1'b0 ;
  assign n19473 = n8398 ^ n7109 ^ 1'b0 ;
  assign n19474 = n8955 ^ n7857 ^ 1'b0 ;
  assign n19475 = ~n6606 & n19474 ;
  assign n19476 = n17640 ^ n10708 ^ n7780 ;
  assign n19480 = n3848 ^ n1360 ^ 1'b0 ;
  assign n19477 = n10407 ^ n7970 ^ 1'b0 ;
  assign n19478 = n11522 | n19477 ;
  assign n19479 = n16760 & ~n19478 ;
  assign n19481 = n19480 ^ n19479 ^ 1'b0 ;
  assign n19482 = n15441 | n19481 ;
  assign n19483 = ( ~n7733 & n19476 ) | ( ~n7733 & n19482 ) | ( n19476 & n19482 ) ;
  assign n19484 = n19475 & ~n19483 ;
  assign n19485 = n610 & n19484 ;
  assign n19489 = ( n4933 & n5205 ) | ( n4933 & ~n6739 ) | ( n5205 & ~n6739 ) ;
  assign n19490 = ( ~n863 & n7695 ) | ( ~n863 & n19489 ) | ( n7695 & n19489 ) ;
  assign n19491 = ~n3504 & n19490 ;
  assign n19492 = n4384 & n19491 ;
  assign n19486 = n9936 ^ n1248 ^ 1'b0 ;
  assign n19487 = ~n3677 & n19486 ;
  assign n19488 = n17243 & n19487 ;
  assign n19493 = n19492 ^ n19488 ^ 1'b0 ;
  assign n19494 = n1982 & n9157 ;
  assign n19495 = ~n431 & n19494 ;
  assign n19496 = n19495 ^ n5780 ^ 1'b0 ;
  assign n19497 = n11442 | n19496 ;
  assign n19499 = n2052 & ~n14205 ;
  assign n19500 = n12718 & n19499 ;
  assign n19498 = ( n530 & ~n4127 ) | ( n530 & n6609 ) | ( ~n4127 & n6609 ) ;
  assign n19501 = n19500 ^ n19498 ^ n5549 ;
  assign n19502 = n7639 & n14663 ;
  assign n19503 = ~n19501 & n19502 ;
  assign n19504 = ( n1050 & n11606 ) | ( n1050 & n12844 ) | ( n11606 & n12844 ) ;
  assign n19505 = n14757 ^ n1714 ^ 1'b0 ;
  assign n19506 = ( n7092 & n17407 ) | ( n7092 & n19505 ) | ( n17407 & n19505 ) ;
  assign n19511 = n18494 ^ n7317 ^ n2491 ;
  assign n19507 = n9118 & ~n10416 ;
  assign n19508 = n18936 ^ n14559 ^ 1'b0 ;
  assign n19509 = n12577 & ~n19508 ;
  assign n19510 = ~n19507 & n19509 ;
  assign n19512 = n19511 ^ n19510 ^ n6744 ;
  assign n19513 = n8548 ^ n3883 ^ 1'b0 ;
  assign n19514 = ( x29 & ~n8145 ) | ( x29 & n10765 ) | ( ~n8145 & n10765 ) ;
  assign n19515 = n16714 & n19514 ;
  assign n19516 = n19513 & n19515 ;
  assign n19517 = ~n2838 & n6661 ;
  assign n19518 = n1707 & ~n19517 ;
  assign n19519 = n19518 ^ n1695 ^ n428 ;
  assign n19520 = ( n19512 & ~n19516 ) | ( n19512 & n19519 ) | ( ~n19516 & n19519 ) ;
  assign n19521 = ( n3341 & n8288 ) | ( n3341 & n9411 ) | ( n8288 & n9411 ) ;
  assign n19522 = n19521 ^ n14109 ^ 1'b0 ;
  assign n19523 = n12740 ^ n12235 ^ 1'b0 ;
  assign n19524 = n14656 ^ n10062 ^ n3513 ;
  assign n19525 = n7408 | n12958 ;
  assign n19526 = n19524 & ~n19525 ;
  assign n19527 = n19523 & n19526 ;
  assign n19528 = n3292 & ~n4956 ;
  assign n19529 = n16704 ^ n11546 ^ 1'b0 ;
  assign n19530 = ~n19528 & n19529 ;
  assign n19531 = n18291 ^ n10481 ^ 1'b0 ;
  assign n19532 = n562 & ~n9071 ;
  assign n19533 = n15036 ^ n12523 ^ n7435 ;
  assign n19534 = ( n4403 & n19532 ) | ( n4403 & n19533 ) | ( n19532 & n19533 ) ;
  assign n19535 = n19534 ^ n8730 ^ 1'b0 ;
  assign n19536 = n6267 ^ n5187 ^ n4186 ;
  assign n19537 = ( ~n2258 & n2606 ) | ( ~n2258 & n19536 ) | ( n2606 & n19536 ) ;
  assign n19538 = n19537 ^ n13946 ^ 1'b0 ;
  assign n19539 = n2414 | n8403 ;
  assign n19540 = n19539 ^ n12061 ^ n7962 ;
  assign n19541 = n12341 & n13195 ;
  assign n19542 = n19541 ^ n14324 ^ 1'b0 ;
  assign n19544 = n19089 ^ n13174 ^ n4396 ;
  assign n19543 = n17430 ^ n7133 ^ n6600 ;
  assign n19545 = n19544 ^ n19543 ^ 1'b0 ;
  assign n19546 = n12990 & n19545 ;
  assign n19547 = n19546 ^ n9233 ^ n5266 ;
  assign n19548 = ( n2898 & ~n10608 ) | ( n2898 & n19547 ) | ( ~n10608 & n19547 ) ;
  assign n19549 = n19548 ^ n15077 ^ n9017 ;
  assign n19550 = ~n1143 & n5932 ;
  assign n19551 = n18092 & n19550 ;
  assign n19552 = n16650 ^ n4827 ^ 1'b0 ;
  assign n19553 = n19552 ^ n11867 ^ 1'b0 ;
  assign n19554 = ~n18081 & n19553 ;
  assign n19555 = n760 & n12062 ;
  assign n19558 = ~n2883 & n13700 ;
  assign n19557 = n19073 ^ n4980 ^ n177 ;
  assign n19556 = n7600 & ~n13898 ;
  assign n19559 = n19558 ^ n19557 ^ n19556 ;
  assign n19560 = ( ~n568 & n6014 ) | ( ~n568 & n16540 ) | ( n6014 & n16540 ) ;
  assign n19561 = n4976 & n9328 ;
  assign n19562 = ~n16167 & n19561 ;
  assign n19563 = n13530 ^ n2600 ^ 1'b0 ;
  assign n19564 = n5857 | n19563 ;
  assign n19565 = n317 & ~n5129 ;
  assign n19566 = n19565 ^ n1351 ^ 1'b0 ;
  assign n19567 = ( n10234 & ~n19564 ) | ( n10234 & n19566 ) | ( ~n19564 & n19566 ) ;
  assign n19568 = n7333 ^ n6017 ^ 1'b0 ;
  assign n19569 = n9919 & ~n19568 ;
  assign n19570 = n19569 ^ n10339 ^ n767 ;
  assign n19571 = n19570 ^ n11927 ^ 1'b0 ;
  assign n19572 = n10627 & ~n12049 ;
  assign n19573 = ( n9451 & n14692 ) | ( n9451 & ~n19572 ) | ( n14692 & ~n19572 ) ;
  assign n19574 = ( n1427 & n8602 ) | ( n1427 & ~n16832 ) | ( n8602 & ~n16832 ) ;
  assign n19575 = n5977 | n7538 ;
  assign n19576 = n19575 ^ n16891 ^ 1'b0 ;
  assign n19577 = x41 & n1857 ;
  assign n19578 = ~n7716 & n19577 ;
  assign n19579 = n19578 ^ n2210 ^ 1'b0 ;
  assign n19580 = n19579 ^ n10624 ^ n7877 ;
  assign n19581 = n19580 ^ n17784 ^ n13976 ;
  assign n19582 = ( n14866 & n19576 ) | ( n14866 & ~n19581 ) | ( n19576 & ~n19581 ) ;
  assign n19583 = n10397 ^ n4302 ^ 1'b0 ;
  assign n19584 = n19426 & ~n19583 ;
  assign n19585 = n9012 & ~n11737 ;
  assign n19586 = ~n19584 & n19585 ;
  assign n19587 = n3096 | n19586 ;
  assign n19588 = n2661 & ~n19587 ;
  assign n19589 = n19588 ^ n19221 ^ 1'b0 ;
  assign n19590 = ~n13351 & n17215 ;
  assign n19591 = n19590 ^ n5144 ^ 1'b0 ;
  assign n19592 = n4067 & n19276 ;
  assign n19593 = n1243 & n19592 ;
  assign n19594 = n19593 ^ n1659 ^ 1'b0 ;
  assign n19596 = n3213 & ~n4107 ;
  assign n19597 = ~n962 & n19596 ;
  assign n19598 = n6783 & ~n19597 ;
  assign n19599 = n19598 ^ n8882 ^ 1'b0 ;
  assign n19595 = ( n7634 & n11828 ) | ( n7634 & ~n19544 ) | ( n11828 & ~n19544 ) ;
  assign n19600 = n19599 ^ n19595 ^ n10746 ;
  assign n19601 = n9818 ^ n4654 ^ 1'b0 ;
  assign n19602 = n924 | n13238 ;
  assign n19603 = n5245 & ~n19602 ;
  assign n19604 = n5946 & ~n6814 ;
  assign n19605 = n8478 & n19604 ;
  assign n19606 = n11598 ^ n7008 ^ n5179 ;
  assign n19607 = n19606 ^ n4784 ^ 1'b0 ;
  assign n19608 = n3495 ^ n2661 ^ 1'b0 ;
  assign n19609 = ~n12411 & n19608 ;
  assign n19610 = ( n9167 & ~n18064 ) | ( n9167 & n19609 ) | ( ~n18064 & n19609 ) ;
  assign n19611 = ( ~n8926 & n13292 ) | ( ~n8926 & n18445 ) | ( n13292 & n18445 ) ;
  assign n19612 = n6770 ^ n5199 ^ 1'b0 ;
  assign n19613 = n2820 | n19612 ;
  assign n19614 = n2870 | n4519 ;
  assign n19615 = n19613 & ~n19614 ;
  assign n19616 = ( ~n3629 & n7553 ) | ( ~n3629 & n19615 ) | ( n7553 & n19615 ) ;
  assign n19617 = n19616 ^ n6973 ^ n392 ;
  assign n19619 = ~n2146 & n7140 ;
  assign n19618 = ( n8314 & n8623 ) | ( n8314 & ~n13577 ) | ( n8623 & ~n13577 ) ;
  assign n19620 = n19619 ^ n19618 ^ n12020 ;
  assign n19621 = n6187 ^ n5870 ^ 1'b0 ;
  assign n19622 = n19620 & n19621 ;
  assign n19623 = ~n7332 & n19622 ;
  assign n19624 = n19623 ^ n1926 ^ 1'b0 ;
  assign n19625 = n14240 ^ n8162 ^ 1'b0 ;
  assign n19626 = n19317 ^ n18530 ^ 1'b0 ;
  assign n19627 = ~n19625 & n19626 ;
  assign n19628 = n7993 ^ n1104 ^ 1'b0 ;
  assign n19634 = ~n5905 & n11053 ;
  assign n19635 = n19634 ^ n11479 ^ 1'b0 ;
  assign n19630 = n1059 & n4191 ;
  assign n19631 = ~n8301 & n19630 ;
  assign n19632 = n19631 ^ n15510 ^ n10526 ;
  assign n19629 = n14426 ^ n8660 ^ n2733 ;
  assign n19633 = n19632 ^ n19629 ^ n1083 ;
  assign n19636 = n19635 ^ n19633 ^ n13817 ;
  assign n19637 = ( n205 & n19628 ) | ( n205 & ~n19636 ) | ( n19628 & ~n19636 ) ;
  assign n19638 = ( n6388 & n14803 ) | ( n6388 & ~n19637 ) | ( n14803 & ~n19637 ) ;
  assign n19639 = ( n5685 & n9065 ) | ( n5685 & ~n17717 ) | ( n9065 & ~n17717 ) ;
  assign n19640 = n12849 ^ n9383 ^ n4002 ;
  assign n19641 = ~n8794 & n9666 ;
  assign n19645 = n2464 & n6395 ;
  assign n19646 = n19645 ^ n11491 ^ 1'b0 ;
  assign n19642 = n4005 | n7899 ;
  assign n19643 = n15449 & ~n19642 ;
  assign n19644 = n3092 | n19643 ;
  assign n19647 = n19646 ^ n19644 ^ 1'b0 ;
  assign n19648 = n13928 ^ n7867 ^ 1'b0 ;
  assign n19649 = ( n9978 & ~n19022 ) | ( n9978 & n19648 ) | ( ~n19022 & n19648 ) ;
  assign n19650 = ( ~n10219 & n12867 ) | ( ~n10219 & n14111 ) | ( n12867 & n14111 ) ;
  assign n19651 = ( n14499 & ~n19649 ) | ( n14499 & n19650 ) | ( ~n19649 & n19650 ) ;
  assign n19652 = ~n9543 & n10727 ;
  assign n19653 = ( ~n5306 & n11711 ) | ( ~n5306 & n19652 ) | ( n11711 & n19652 ) ;
  assign n19655 = n16459 ^ n6445 ^ n4535 ;
  assign n19654 = n13137 ^ n3638 ^ 1'b0 ;
  assign n19656 = n19655 ^ n19654 ^ n6133 ;
  assign n19657 = n9148 & n16941 ;
  assign n19658 = n13990 ^ n2632 ^ 1'b0 ;
  assign n19659 = ~n7539 & n19658 ;
  assign n19660 = ( n7932 & n8849 ) | ( n7932 & ~n19659 ) | ( n8849 & ~n19659 ) ;
  assign n19661 = n3097 & ~n5353 ;
  assign n19662 = ~n2016 & n19661 ;
  assign n19663 = ( n1416 & n4694 ) | ( n1416 & n19662 ) | ( n4694 & n19662 ) ;
  assign n19664 = ( ~n1621 & n6893 ) | ( ~n1621 & n19663 ) | ( n6893 & n19663 ) ;
  assign n19665 = ( ~n3810 & n5692 ) | ( ~n3810 & n15333 ) | ( n5692 & n15333 ) ;
  assign n19666 = ( n5865 & n11548 ) | ( n5865 & ~n19665 ) | ( n11548 & ~n19665 ) ;
  assign n19667 = ( n9100 & n19664 ) | ( n9100 & ~n19666 ) | ( n19664 & ~n19666 ) ;
  assign n19668 = n18237 ^ n11866 ^ 1'b0 ;
  assign n19669 = n12241 | n19668 ;
  assign n19670 = n9297 ^ n6489 ^ 1'b0 ;
  assign n19671 = ~n9043 & n19670 ;
  assign n19672 = ~n16986 & n19671 ;
  assign n19673 = n19672 ^ n1538 ^ 1'b0 ;
  assign n19674 = ( n5774 & n12578 ) | ( n5774 & ~n17041 ) | ( n12578 & ~n17041 ) ;
  assign n19675 = n19674 ^ n16092 ^ 1'b0 ;
  assign n19678 = n9779 ^ n4086 ^ 1'b0 ;
  assign n19679 = ~n6359 & n19678 ;
  assign n19676 = n3207 & ~n8400 ;
  assign n19677 = ( n9043 & n15273 ) | ( n9043 & n19676 ) | ( n15273 & n19676 ) ;
  assign n19680 = n19679 ^ n19677 ^ n6235 ;
  assign n19681 = n12186 ^ n10209 ^ 1'b0 ;
  assign n19682 = ~n5127 & n13194 ;
  assign n19686 = n18308 ^ n6289 ^ n6047 ;
  assign n19685 = ( n724 & n4123 ) | ( n724 & n16071 ) | ( n4123 & n16071 ) ;
  assign n19683 = n10713 ^ n8992 ^ n2820 ;
  assign n19684 = n19683 ^ n16645 ^ n8381 ;
  assign n19687 = n19686 ^ n19685 ^ n19684 ;
  assign n19688 = n8454 | n16983 ;
  assign n19689 = n4214 | n9363 ;
  assign n19691 = ( n3953 & n5490 ) | ( n3953 & ~n8775 ) | ( n5490 & ~n8775 ) ;
  assign n19692 = n8925 | n19691 ;
  assign n19693 = n15451 & ~n19692 ;
  assign n19690 = n1567 & ~n16464 ;
  assign n19694 = n19693 ^ n19690 ^ 1'b0 ;
  assign n19695 = n10606 ^ n8352 ^ 1'b0 ;
  assign n19697 = n7430 ^ n4404 ^ 1'b0 ;
  assign n19698 = n1305 & n19697 ;
  assign n19699 = n19698 ^ n5763 ^ n771 ;
  assign n19696 = n6706 & n8624 ;
  assign n19700 = n19699 ^ n19696 ^ 1'b0 ;
  assign n19701 = n19700 ^ n13871 ^ 1'b0 ;
  assign n19703 = n12684 | n16464 ;
  assign n19702 = n7985 ^ n493 ^ n242 ;
  assign n19704 = n19703 ^ n19702 ^ n13489 ;
  assign n19705 = n19054 ^ n8651 ^ n3220 ;
  assign n19707 = n10233 ^ n8699 ^ n2169 ;
  assign n19706 = n6784 & ~n15980 ;
  assign n19708 = n19707 ^ n19706 ^ n6495 ;
  assign n19709 = ~n2118 & n9155 ;
  assign n19710 = n19500 ^ n18554 ^ n9860 ;
  assign n19711 = ( ~n1316 & n2622 ) | ( ~n1316 & n19710 ) | ( n2622 & n19710 ) ;
  assign n19712 = ( ~n16081 & n19709 ) | ( ~n16081 & n19711 ) | ( n19709 & n19711 ) ;
  assign n19713 = n1756 & ~n8333 ;
  assign n19714 = n18002 ^ n2009 ^ 1'b0 ;
  assign n19715 = n2560 | n19714 ;
  assign n19716 = n5415 ^ n2647 ^ n941 ;
  assign n19717 = ( n2824 & n7689 ) | ( n2824 & n19716 ) | ( n7689 & n19716 ) ;
  assign n19718 = n19717 ^ n13270 ^ n1863 ;
  assign n19719 = n7473 ^ n3295 ^ 1'b0 ;
  assign n19720 = n18626 ^ n18563 ^ n7484 ;
  assign n19721 = n3448 ^ n1259 ^ 1'b0 ;
  assign n19722 = ( n7332 & n19720 ) | ( n7332 & ~n19721 ) | ( n19720 & ~n19721 ) ;
  assign n19723 = ~n19719 & n19722 ;
  assign n19724 = ( ~n3140 & n11149 ) | ( ~n3140 & n16457 ) | ( n11149 & n16457 ) ;
  assign n19725 = ~n1503 & n5016 ;
  assign n19726 = n19725 ^ n5535 ^ 1'b0 ;
  assign n19727 = n19726 ^ n16803 ^ n15889 ;
  assign n19728 = ( n1629 & n2184 ) | ( n1629 & n17590 ) | ( n2184 & n17590 ) ;
  assign n19729 = n12674 ^ n9298 ^ 1'b0 ;
  assign n19730 = n3147 & ~n19729 ;
  assign n19731 = n1124 & n19730 ;
  assign n19732 = ( n12830 & n19728 ) | ( n12830 & n19731 ) | ( n19728 & n19731 ) ;
  assign n19733 = n834 ^ n393 ^ 1'b0 ;
  assign n19734 = n10952 | n19733 ;
  assign n19735 = ~n11435 & n19734 ;
  assign n19737 = n5934 ^ n434 ^ x122 ;
  assign n19736 = ~n7957 & n13873 ;
  assign n19738 = n19737 ^ n19736 ^ 1'b0 ;
  assign n19739 = n19738 ^ n5785 ^ n875 ;
  assign n19740 = n19739 ^ n17667 ^ n730 ;
  assign n19741 = n10288 ^ n8352 ^ n6822 ;
  assign n19742 = n8241 & n19741 ;
  assign n19743 = n1146 & ~n9310 ;
  assign n19744 = ~n2172 & n19743 ;
  assign n19745 = ( n5518 & ~n12198 ) | ( n5518 & n14729 ) | ( ~n12198 & n14729 ) ;
  assign n19746 = n12321 ^ n11683 ^ 1'b0 ;
  assign n19747 = n6623 & n16919 ;
  assign n19748 = n12136 & n19747 ;
  assign n19749 = n6524 & ~n19748 ;
  assign n19750 = n16027 ^ n12704 ^ n5573 ;
  assign n19751 = ( n5780 & n7500 ) | ( n5780 & n19750 ) | ( n7500 & n19750 ) ;
  assign n19752 = n4690 | n12690 ;
  assign n19753 = n2537 & ~n19752 ;
  assign n19754 = n8364 & n19753 ;
  assign n19755 = n9927 ^ n8637 ^ n3352 ;
  assign n19756 = ( ~n5419 & n16689 ) | ( ~n5419 & n19755 ) | ( n16689 & n19755 ) ;
  assign n19757 = n1205 | n18936 ;
  assign n19758 = n19757 ^ n16827 ^ 1'b0 ;
  assign n19759 = n16534 ^ n6452 ^ 1'b0 ;
  assign n19760 = ( ~n834 & n3875 ) | ( ~n834 & n15555 ) | ( n3875 & n15555 ) ;
  assign n19761 = n19760 ^ n4558 ^ n1488 ;
  assign n19762 = n17293 | n19761 ;
  assign n19763 = n330 | n19762 ;
  assign n19764 = ~n12184 & n19763 ;
  assign n19765 = n3205 & n16856 ;
  assign n19766 = n5187 | n19765 ;
  assign n19767 = n180 & ~n19766 ;
  assign n19768 = ( n5711 & n11966 ) | ( n5711 & n18219 ) | ( n11966 & n18219 ) ;
  assign n19769 = n19768 ^ n7782 ^ 1'b0 ;
  assign n19770 = n11164 | n19769 ;
  assign n19771 = n194 & ~n635 ;
  assign n19772 = n1313 & ~n19771 ;
  assign n19773 = n13092 ^ n10268 ^ n4678 ;
  assign n19774 = n4844 | n18143 ;
  assign n19775 = n11866 | n19774 ;
  assign n19776 = n19775 ^ n11084 ^ 1'b0 ;
  assign n19777 = ~n8642 & n19776 ;
  assign n19778 = ( ~n12071 & n12923 ) | ( ~n12071 & n14482 ) | ( n12923 & n14482 ) ;
  assign n19779 = ~n13099 & n17130 ;
  assign n19780 = n6941 ^ n3903 ^ n1970 ;
  assign n19781 = n19780 ^ n1348 ^ 1'b0 ;
  assign n19782 = n7688 & ~n12680 ;
  assign n19783 = n11698 & n19782 ;
  assign n19784 = n5718 | n19783 ;
  assign n19785 = n19784 ^ n12875 ^ 1'b0 ;
  assign n19786 = n16074 ^ n8656 ^ n4081 ;
  assign n19787 = n691 & ~n1786 ;
  assign n19788 = n4250 & n19787 ;
  assign n19789 = n12674 | n19788 ;
  assign n19790 = n7847 ^ n4572 ^ 1'b0 ;
  assign n19791 = ( n2011 & ~n4342 ) | ( n2011 & n7564 ) | ( ~n4342 & n7564 ) ;
  assign n19792 = n1425 ^ n1260 ^ 1'b0 ;
  assign n19793 = n19792 ^ n12707 ^ 1'b0 ;
  assign n19794 = ~n19791 & n19793 ;
  assign n19795 = n12923 & n19794 ;
  assign n19796 = n11015 & n19795 ;
  assign n19797 = n19796 ^ n18127 ^ 1'b0 ;
  assign n19798 = ( n1754 & n2901 ) | ( n1754 & n13894 ) | ( n2901 & n13894 ) ;
  assign n19799 = ~n14254 & n19798 ;
  assign n19800 = n13321 ^ n11183 ^ n3024 ;
  assign n19801 = n19800 ^ n2181 ^ 1'b0 ;
  assign n19802 = n2809 & n19801 ;
  assign n19803 = n6553 | n12972 ;
  assign n19804 = n19803 ^ n1357 ^ 1'b0 ;
  assign n19805 = n3990 ^ n676 ^ 1'b0 ;
  assign n19806 = n19804 & ~n19805 ;
  assign n19807 = n8583 ^ n1069 ^ 1'b0 ;
  assign n19808 = n9173 ^ n1426 ^ n340 ;
  assign n19809 = ( n4158 & n19807 ) | ( n4158 & n19808 ) | ( n19807 & n19808 ) ;
  assign n19810 = n256 | n2100 ;
  assign n19811 = n3317 | n19810 ;
  assign n19812 = n19811 ^ n19204 ^ n6187 ;
  assign n19817 = ( n4209 & ~n6090 ) | ( n4209 & n13914 ) | ( ~n6090 & n13914 ) ;
  assign n19815 = n2733 & n8387 ;
  assign n19813 = n15188 ^ n7141 ^ n147 ;
  assign n19814 = ~n8636 & n19813 ;
  assign n19816 = n19815 ^ n19814 ^ n13987 ;
  assign n19818 = n19817 ^ n19816 ^ n686 ;
  assign n19819 = n9854 | n11496 ;
  assign n19820 = n19355 | n19819 ;
  assign n19821 = n409 | n2550 ;
  assign n19822 = n19821 ^ n7028 ^ 1'b0 ;
  assign n19823 = ( n2021 & ~n2894 ) | ( n2021 & n19822 ) | ( ~n2894 & n19822 ) ;
  assign n19824 = n19823 ^ n5870 ^ x38 ;
  assign n19825 = n9719 & ~n19824 ;
  assign n19826 = n6458 ^ n4587 ^ n840 ;
  assign n19827 = ~n3164 & n19826 ;
  assign n19828 = n19827 ^ n12654 ^ 1'b0 ;
  assign n19829 = n15973 | n19828 ;
  assign n19830 = n4535 & ~n19829 ;
  assign n19831 = ( n4123 & ~n4874 ) | ( n4123 & n16997 ) | ( ~n4874 & n16997 ) ;
  assign n19832 = ( n1614 & n11586 ) | ( n1614 & ~n19831 ) | ( n11586 & ~n19831 ) ;
  assign n19833 = n12634 ^ n11881 ^ n6380 ;
  assign n19834 = n19833 ^ n9772 ^ n7334 ;
  assign n19839 = n9345 ^ n5944 ^ 1'b0 ;
  assign n19840 = n17384 & n19839 ;
  assign n19835 = n14290 ^ n4377 ^ 1'b0 ;
  assign n19836 = n2968 & n19835 ;
  assign n19837 = n19836 ^ n6145 ^ n5230 ;
  assign n19838 = ( ~n1445 & n19245 ) | ( ~n1445 & n19837 ) | ( n19245 & n19837 ) ;
  assign n19841 = n19840 ^ n19838 ^ n7040 ;
  assign n19842 = n12728 ^ n12653 ^ n8970 ;
  assign n19843 = n6370 | n19211 ;
  assign n19848 = ( n725 & ~n1651 ) | ( n725 & n7710 ) | ( ~n1651 & n7710 ) ;
  assign n19844 = n3749 ^ n3297 ^ n222 ;
  assign n19845 = n8119 & n19844 ;
  assign n19846 = n19845 ^ n11046 ^ 1'b0 ;
  assign n19847 = n11079 | n19846 ;
  assign n19849 = n19848 ^ n19847 ^ 1'b0 ;
  assign n19850 = n12403 ^ n4775 ^ n1644 ;
  assign n19851 = n19850 ^ n15722 ^ n3976 ;
  assign n19852 = ~n5594 & n19851 ;
  assign n19853 = ( n2157 & n2511 ) | ( n2157 & ~n2657 ) | ( n2511 & ~n2657 ) ;
  assign n19854 = n3364 & ~n19853 ;
  assign n19855 = n17443 & ~n19854 ;
  assign n19856 = n9233 ^ n6975 ^ n2546 ;
  assign n19857 = n19026 ^ n5652 ^ 1'b0 ;
  assign n19862 = n6175 ^ n5774 ^ n1982 ;
  assign n19863 = n19862 ^ n17489 ^ n5922 ;
  assign n19858 = n7626 ^ n2422 ^ 1'b0 ;
  assign n19859 = n1300 | n19858 ;
  assign n19860 = n19859 ^ n15113 ^ n1982 ;
  assign n19861 = n19860 ^ n18480 ^ n7280 ;
  assign n19864 = n19863 ^ n19861 ^ n9417 ;
  assign n19865 = n12626 ^ n8015 ^ n4983 ;
  assign n19866 = ~n4660 & n19865 ;
  assign n19867 = n4776 ^ n2783 ^ 1'b0 ;
  assign n19868 = n3628 | n19867 ;
  assign n19869 = n619 | n19613 ;
  assign n19870 = n19868 & ~n19869 ;
  assign n19871 = n12508 & ~n19870 ;
  assign n19872 = ~n12367 & n19871 ;
  assign n19873 = n11912 & ~n18372 ;
  assign n19874 = ~n2782 & n19873 ;
  assign n19875 = n4271 | n7008 ;
  assign n19876 = n234 | n547 ;
  assign n19877 = n19875 & ~n19876 ;
  assign n19878 = ( n1021 & n5865 ) | ( n1021 & ~n6891 ) | ( n5865 & ~n6891 ) ;
  assign n19879 = n19878 ^ n19442 ^ n18870 ;
  assign n19880 = n2128 & ~n11471 ;
  assign n19881 = n17826 | n19880 ;
  assign n19882 = n5008 & n10072 ;
  assign n19883 = n4811 ^ n1909 ^ 1'b0 ;
  assign n19884 = n4948 | n19883 ;
  assign n19885 = n13961 ^ n4929 ^ 1'b0 ;
  assign n19886 = n231 & ~n6913 ;
  assign n19887 = ~x111 & n19886 ;
  assign n19888 = ( n2616 & ~n7479 ) | ( n2616 & n11897 ) | ( ~n7479 & n11897 ) ;
  assign n19889 = n19888 ^ n7228 ^ 1'b0 ;
  assign n19890 = ~n5784 & n19889 ;
  assign n19891 = ( ~n3713 & n19887 ) | ( ~n3713 & n19890 ) | ( n19887 & n19890 ) ;
  assign n19892 = ( n17123 & n19885 ) | ( n17123 & n19891 ) | ( n19885 & n19891 ) ;
  assign n19897 = n14036 ^ n7731 ^ 1'b0 ;
  assign n19898 = ~n9542 & n19897 ;
  assign n19893 = n3941 ^ n3238 ^ x65 ;
  assign n19894 = n7001 ^ n2035 ^ 1'b0 ;
  assign n19895 = n19893 & n19894 ;
  assign n19896 = ~n15997 & n19895 ;
  assign n19899 = n19898 ^ n19896 ^ 1'b0 ;
  assign n19901 = n2753 & n4848 ;
  assign n19902 = n19901 ^ n7675 ^ 1'b0 ;
  assign n19900 = ( n691 & n2695 ) | ( n691 & n4253 ) | ( n2695 & n4253 ) ;
  assign n19903 = n19902 ^ n19900 ^ 1'b0 ;
  assign n19904 = ( n607 & ~n8334 ) | ( n607 & n19903 ) | ( ~n8334 & n19903 ) ;
  assign n19905 = ( ~n157 & n6903 ) | ( ~n157 & n11543 ) | ( n6903 & n11543 ) ;
  assign n19906 = n19905 ^ n410 ^ 1'b0 ;
  assign n19907 = n18913 ^ n9872 ^ 1'b0 ;
  assign n19908 = ( n8366 & n19906 ) | ( n8366 & n19907 ) | ( n19906 & n19907 ) ;
  assign n19909 = ~n3436 & n4884 ;
  assign n19910 = n19909 ^ n2679 ^ 1'b0 ;
  assign n19911 = ~n11256 & n12186 ;
  assign n19912 = ( n14866 & n19910 ) | ( n14866 & ~n19911 ) | ( n19910 & ~n19911 ) ;
  assign n19913 = n3706 | n14424 ;
  assign n19914 = n14650 | n19913 ;
  assign n19915 = ~n2152 & n19914 ;
  assign n19916 = ~n12260 & n19915 ;
  assign n19917 = n19060 ^ n2422 ^ 1'b0 ;
  assign n19918 = n19917 ^ n16874 ^ 1'b0 ;
  assign n19919 = n2371 & n2632 ;
  assign n19920 = n8476 & n19919 ;
  assign n19921 = ( n3070 & n3650 ) | ( n3070 & n9666 ) | ( n3650 & n9666 ) ;
  assign n19922 = ( n16752 & ~n19920 ) | ( n16752 & n19921 ) | ( ~n19920 & n19921 ) ;
  assign n19924 = n4220 ^ n4066 ^ 1'b0 ;
  assign n19923 = n8371 & n10327 ;
  assign n19925 = n19924 ^ n19923 ^ 1'b0 ;
  assign n19926 = n579 & ~n5198 ;
  assign n19927 = n19926 ^ n15453 ^ n12075 ;
  assign n19928 = n14094 & ~n19060 ;
  assign n19929 = n19928 ^ n3941 ^ 1'b0 ;
  assign n19930 = n13206 ^ n9728 ^ n9100 ;
  assign n19931 = n11263 ^ n6663 ^ n519 ;
  assign n19932 = n6406 & ~n19931 ;
  assign n19933 = n19932 ^ n1848 ^ 1'b0 ;
  assign n19934 = n19933 ^ n15237 ^ n1584 ;
  assign n19935 = n6489 ^ n2086 ^ 1'b0 ;
  assign n19936 = n4478 & ~n19935 ;
  assign n19937 = ( ~n2817 & n5974 ) | ( ~n2817 & n16072 ) | ( n5974 & n16072 ) ;
  assign n19938 = ( n10664 & n14962 ) | ( n10664 & n19937 ) | ( n14962 & n19937 ) ;
  assign n19939 = n6747 ^ n474 ^ 1'b0 ;
  assign n19940 = n16846 & ~n18621 ;
  assign n19941 = n12914 & ~n13633 ;
  assign n19942 = n19941 ^ n5264 ^ 1'b0 ;
  assign n19943 = n11586 ^ n686 ^ 1'b0 ;
  assign n19944 = n15203 | n19943 ;
  assign n19945 = n15604 ^ n8882 ^ n7584 ;
  assign n19946 = ( n409 & ~n16717 ) | ( n409 & n19945 ) | ( ~n16717 & n19945 ) ;
  assign n19947 = ~n11556 & n16186 ;
  assign n19948 = n19946 & n19947 ;
  assign n19949 = n9797 ^ n6469 ^ 1'b0 ;
  assign n19950 = ~n3539 & n19949 ;
  assign n19951 = n19950 ^ n4185 ^ 1'b0 ;
  assign n19952 = n11215 ^ n1192 ^ 1'b0 ;
  assign n19953 = n19951 | n19952 ;
  assign n19954 = n5178 & n6729 ;
  assign n19955 = n19954 ^ n5325 ^ 1'b0 ;
  assign n19956 = ( n1828 & n2272 ) | ( n1828 & ~n19955 ) | ( n2272 & ~n19955 ) ;
  assign n19957 = n1585 & n19386 ;
  assign n19958 = ~n12177 & n19957 ;
  assign n19959 = ( n7594 & n10673 ) | ( n7594 & ~n19958 ) | ( n10673 & ~n19958 ) ;
  assign n19960 = n19439 & n19959 ;
  assign n19961 = ~n1011 & n19960 ;
  assign n19962 = n16409 ^ n9778 ^ 1'b0 ;
  assign n19963 = ~n5907 & n8778 ;
  assign n19964 = n3302 & n19963 ;
  assign n19965 = n9118 & n19964 ;
  assign n19966 = n3858 & n15094 ;
  assign n19967 = n19966 ^ n18259 ^ 1'b0 ;
  assign n19968 = n1748 & n19967 ;
  assign n19969 = n16333 & n19968 ;
  assign n19970 = n7158 ^ n4367 ^ 1'b0 ;
  assign n19971 = ( n5931 & n8896 ) | ( n5931 & n19970 ) | ( n8896 & n19970 ) ;
  assign n19972 = n19971 ^ n10203 ^ n8190 ;
  assign n19973 = ~n794 & n19972 ;
  assign n19974 = ( ~n4576 & n8781 ) | ( ~n4576 & n16402 ) | ( n8781 & n16402 ) ;
  assign n19975 = n19974 ^ n13835 ^ n6991 ;
  assign n19976 = n13421 | n16152 ;
  assign n19977 = n16606 ^ n8023 ^ n3384 ;
  assign n19978 = n935 & ~n11624 ;
  assign n19979 = n19978 ^ n11344 ^ 1'b0 ;
  assign n19980 = n11897 ^ n3864 ^ 1'b0 ;
  assign n19981 = n8869 & n19980 ;
  assign n19982 = n4068 & n19981 ;
  assign n19983 = ~n9501 & n19982 ;
  assign n19984 = ( n1601 & ~n4187 ) | ( n1601 & n19983 ) | ( ~n4187 & n19983 ) ;
  assign n19986 = n373 & ~n8537 ;
  assign n19987 = ~n11141 & n19986 ;
  assign n19985 = n8193 ^ n7332 ^ n7142 ;
  assign n19988 = n19987 ^ n19985 ^ n11741 ;
  assign n19989 = n3530 & ~n8937 ;
  assign n19990 = n7031 ^ n6696 ^ 1'b0 ;
  assign n19991 = n6699 & n19990 ;
  assign n19992 = n18827 ^ n14752 ^ n5957 ;
  assign n19993 = ( ~n9846 & n18202 ) | ( ~n9846 & n19992 ) | ( n18202 & n19992 ) ;
  assign n19994 = n260 & ~n1691 ;
  assign n19995 = n2666 & n19994 ;
  assign n19996 = n3776 ^ n744 ^ 1'b0 ;
  assign n19997 = n2599 ^ n839 ^ 1'b0 ;
  assign n19998 = n19996 | n19997 ;
  assign n19999 = ( n7722 & n19995 ) | ( n7722 & n19998 ) | ( n19995 & n19998 ) ;
  assign n20000 = ( n5304 & ~n11835 ) | ( n5304 & n19999 ) | ( ~n11835 & n19999 ) ;
  assign n20001 = ( ~n568 & n5655 ) | ( ~n568 & n13731 ) | ( n5655 & n13731 ) ;
  assign n20002 = n16923 ^ n9516 ^ 1'b0 ;
  assign n20003 = n20001 | n20002 ;
  assign n20004 = n6450 ^ n1814 ^ 1'b0 ;
  assign n20005 = n20004 ^ n11587 ^ n8355 ;
  assign n20006 = n10338 | n20005 ;
  assign n20007 = n3638 | n20006 ;
  assign n20008 = n20007 ^ n19537 ^ 1'b0 ;
  assign n20009 = n1007 | n7362 ;
  assign n20010 = n20008 & ~n20009 ;
  assign n20011 = n19944 ^ n17936 ^ 1'b0 ;
  assign n20014 = n11344 | n19489 ;
  assign n20015 = n20014 ^ n2815 ^ 1'b0 ;
  assign n20012 = n14053 ^ n5729 ^ n3036 ;
  assign n20013 = n20012 ^ n2206 ^ n910 ;
  assign n20016 = n20015 ^ n20013 ^ x108 ;
  assign n20017 = ( n5225 & n12940 ) | ( n5225 & ~n13314 ) | ( n12940 & ~n13314 ) ;
  assign n20018 = n4144 & n15797 ;
  assign n20019 = n19016 ^ n13110 ^ n5969 ;
  assign n20020 = ~n709 & n1876 ;
  assign n20021 = ~n5741 & n20020 ;
  assign n20022 = ( n702 & ~n10220 ) | ( n702 & n10983 ) | ( ~n10220 & n10983 ) ;
  assign n20023 = ~n20021 & n20022 ;
  assign n20024 = ~n7546 & n20023 ;
  assign n20025 = ( n513 & n4923 ) | ( n513 & n12161 ) | ( n4923 & n12161 ) ;
  assign n20026 = n508 | n1945 ;
  assign n20027 = n17130 & ~n20026 ;
  assign n20028 = ( n4500 & ~n9006 ) | ( n4500 & n10998 ) | ( ~n9006 & n10998 ) ;
  assign n20029 = ( n3009 & ~n20027 ) | ( n3009 & n20028 ) | ( ~n20027 & n20028 ) ;
  assign n20030 = n2142 & ~n2296 ;
  assign n20032 = ( ~n1522 & n2466 ) | ( ~n1522 & n2878 ) | ( n2466 & n2878 ) ;
  assign n20031 = n17411 ^ n16362 ^ n4803 ;
  assign n20033 = n20032 ^ n20031 ^ n4510 ;
  assign n20034 = n20033 ^ n7795 ^ n1795 ;
  assign n20035 = n18116 ^ n5740 ^ n2922 ;
  assign n20036 = n15430 ^ n533 ^ 1'b0 ;
  assign n20037 = n20036 ^ n14151 ^ 1'b0 ;
  assign n20038 = n20035 & n20037 ;
  assign n20039 = n4980 ^ n2403 ^ 1'b0 ;
  assign n20040 = n13642 & n20039 ;
  assign n20041 = ~n17875 & n20040 ;
  assign n20042 = n20041 ^ n10155 ^ 1'b0 ;
  assign n20043 = n15492 ^ n12056 ^ 1'b0 ;
  assign n20044 = ( n2321 & n5699 ) | ( n2321 & n20043 ) | ( n5699 & n20043 ) ;
  assign n20045 = n9344 ^ n2207 ^ 1'b0 ;
  assign n20046 = n4366 & n4373 ;
  assign n20047 = n3023 & n20046 ;
  assign n20048 = n7863 ^ n3424 ^ 1'b0 ;
  assign n20049 = n13561 | n20048 ;
  assign n20050 = ( n8800 & ~n20047 ) | ( n8800 & n20049 ) | ( ~n20047 & n20049 ) ;
  assign n20051 = ( n9008 & n20045 ) | ( n9008 & ~n20050 ) | ( n20045 & ~n20050 ) ;
  assign n20052 = n20051 ^ n4776 ^ 1'b0 ;
  assign n20053 = n20044 & ~n20052 ;
  assign n20054 = n2383 ^ n2073 ^ 1'b0 ;
  assign n20055 = ~n11952 & n15038 ;
  assign n20056 = n907 | n13105 ;
  assign n20057 = n8860 | n20056 ;
  assign n20058 = n2982 | n10884 ;
  assign n20059 = n20057 | n20058 ;
  assign n20060 = n20059 ^ n8334 ^ n2124 ;
  assign n20061 = n19946 ^ n4819 ^ n4611 ;
  assign n20062 = n5408 ^ n1575 ^ 1'b0 ;
  assign n20063 = ( n16027 & n20061 ) | ( n16027 & ~n20062 ) | ( n20061 & ~n20062 ) ;
  assign n20064 = n13963 & ~n20063 ;
  assign n20065 = ( ~n10201 & n10524 ) | ( ~n10201 & n20064 ) | ( n10524 & n20064 ) ;
  assign n20066 = ~n450 & n1403 ;
  assign n20067 = n4621 & n20066 ;
  assign n20068 = n20067 ^ n18842 ^ n12444 ;
  assign n20069 = ( ~n3661 & n4679 ) | ( ~n3661 & n4974 ) | ( n4679 & n4974 ) ;
  assign n20070 = n12046 & n20069 ;
  assign n20071 = n10416 & n20070 ;
  assign n20072 = n8693 & ~n20071 ;
  assign n20073 = n2407 | n9137 ;
  assign n20074 = n15923 | n20073 ;
  assign n20075 = x70 & n4217 ;
  assign n20076 = n20075 ^ n9946 ^ 1'b0 ;
  assign n20077 = n15400 ^ n7017 ^ n3127 ;
  assign n20078 = ~n7185 & n20077 ;
  assign n20079 = n16702 ^ n13722 ^ n9925 ;
  assign n20080 = ( n6316 & n10878 ) | ( n6316 & n20079 ) | ( n10878 & n20079 ) ;
  assign n20081 = n14889 ^ n14752 ^ n316 ;
  assign n20082 = n4342 & n18763 ;
  assign n20083 = n10063 ^ n8024 ^ 1'b0 ;
  assign n20084 = n5186 & ~n20083 ;
  assign n20085 = n20084 ^ n7840 ^ 1'b0 ;
  assign n20086 = n20082 & n20085 ;
  assign n20089 = n7942 ^ n5949 ^ 1'b0 ;
  assign n20090 = n1408 ^ n1284 ^ 1'b0 ;
  assign n20091 = n2211 & ~n20090 ;
  assign n20092 = ( n2963 & ~n20089 ) | ( n2963 & n20091 ) | ( ~n20089 & n20091 ) ;
  assign n20087 = ~n4193 & n6038 ;
  assign n20088 = n20087 ^ n1412 ^ 1'b0 ;
  assign n20093 = n20092 ^ n20088 ^ n493 ;
  assign n20094 = ( n4776 & ~n11230 ) | ( n4776 & n20093 ) | ( ~n11230 & n20093 ) ;
  assign n20097 = n11009 ^ n2184 ^ 1'b0 ;
  assign n20095 = n4503 & n8600 ;
  assign n20096 = n4231 & n20095 ;
  assign n20098 = n20097 ^ n20096 ^ 1'b0 ;
  assign n20103 = ( n7351 & ~n11579 ) | ( n7351 & n13621 ) | ( ~n11579 & n13621 ) ;
  assign n20101 = ~n764 & n3334 ;
  assign n20102 = ~n1566 & n20101 ;
  assign n20104 = n20103 ^ n20102 ^ n11292 ;
  assign n20099 = ( n1899 & n6319 ) | ( n1899 & n6633 ) | ( n6319 & n6633 ) ;
  assign n20100 = ( n1233 & n3242 ) | ( n1233 & n20099 ) | ( n3242 & n20099 ) ;
  assign n20105 = n20104 ^ n20100 ^ 1'b0 ;
  assign n20106 = n4813 ^ n2747 ^ 1'b0 ;
  assign n20107 = ( n14705 & n17654 ) | ( n14705 & n20106 ) | ( n17654 & n20106 ) ;
  assign n20109 = n12203 ^ n466 ^ 1'b0 ;
  assign n20108 = n10479 & n14070 ;
  assign n20110 = n20109 ^ n20108 ^ 1'b0 ;
  assign n20111 = n4321 & n7655 ;
  assign n20112 = n1261 & n20111 ;
  assign n20113 = n20112 ^ n4315 ^ 1'b0 ;
  assign n20114 = n11099 ^ n3925 ^ n247 ;
  assign n20115 = ( n3097 & n10569 ) | ( n3097 & ~n14173 ) | ( n10569 & ~n14173 ) ;
  assign n20116 = n20114 & ~n20115 ;
  assign n20117 = n20113 & n20116 ;
  assign n20118 = ( ~n1192 & n5745 ) | ( ~n1192 & n6060 ) | ( n5745 & n6060 ) ;
  assign n20119 = ( n397 & ~n2065 ) | ( n397 & n11222 ) | ( ~n2065 & n11222 ) ;
  assign n20120 = n2161 ^ n673 ^ 1'b0 ;
  assign n20121 = n1182 & ~n20120 ;
  assign n20122 = ~n20119 & n20121 ;
  assign n20123 = n20122 ^ n8170 ^ 1'b0 ;
  assign n20124 = ( ~n7813 & n9497 ) | ( ~n7813 & n20123 ) | ( n9497 & n20123 ) ;
  assign n20125 = n20124 ^ n6421 ^ 1'b0 ;
  assign n20126 = ( n3990 & n4918 ) | ( n3990 & n5268 ) | ( n4918 & n5268 ) ;
  assign n20127 = ( ~n1430 & n10852 ) | ( ~n1430 & n20126 ) | ( n10852 & n20126 ) ;
  assign n20128 = n20127 ^ n10048 ^ n947 ;
  assign n20129 = ~x84 & n7401 ;
  assign n20130 = n11125 & n20129 ;
  assign n20131 = ( n5723 & n20128 ) | ( n5723 & ~n20130 ) | ( n20128 & ~n20130 ) ;
  assign n20132 = n20131 ^ n19815 ^ n5753 ;
  assign n20133 = n20132 ^ n12233 ^ n10370 ;
  assign n20135 = n5036 ^ n1002 ^ 1'b0 ;
  assign n20136 = n20135 ^ n11694 ^ n1756 ;
  assign n20137 = n20136 ^ n17597 ^ n8695 ;
  assign n20134 = ~n4236 & n14729 ;
  assign n20138 = n20137 ^ n20134 ^ 1'b0 ;
  assign n20139 = n1923 & n10917 ;
  assign n20140 = n20139 ^ n5018 ^ 1'b0 ;
  assign n20141 = n20140 ^ n14441 ^ n9654 ;
  assign n20142 = ~n4519 & n20141 ;
  assign n20143 = ~n12781 & n20142 ;
  assign n20144 = n20143 ^ n11611 ^ 1'b0 ;
  assign n20145 = n19304 & ~n20144 ;
  assign n20146 = ( n1391 & n1853 ) | ( n1391 & n18561 ) | ( n1853 & n18561 ) ;
  assign n20151 = ( ~n1728 & n3433 ) | ( ~n1728 & n4727 ) | ( n3433 & n4727 ) ;
  assign n20149 = n13068 ^ n4767 ^ 1'b0 ;
  assign n20147 = n5796 | n8148 ;
  assign n20148 = n6883 & ~n20147 ;
  assign n20150 = n20149 ^ n20148 ^ n4513 ;
  assign n20152 = n20151 ^ n20150 ^ n7504 ;
  assign n20153 = n15423 ^ n6254 ^ 1'b0 ;
  assign n20154 = n20153 ^ n9867 ^ n4976 ;
  assign n20155 = n11750 ^ n9640 ^ n8337 ;
  assign n20156 = n16035 ^ n9994 ^ 1'b0 ;
  assign n20157 = n20155 | n20156 ;
  assign n20158 = n20157 ^ n18595 ^ 1'b0 ;
  assign n20165 = n3582 | n4344 ;
  assign n20166 = n20165 ^ n7964 ^ 1'b0 ;
  assign n20164 = n2894 & n19775 ;
  assign n20167 = n20166 ^ n20164 ^ 1'b0 ;
  assign n20168 = ( n8646 & n9792 ) | ( n8646 & n20167 ) | ( n9792 & n20167 ) ;
  assign n20160 = n7456 & ~n16941 ;
  assign n20161 = n20160 ^ n3351 ^ 1'b0 ;
  assign n20162 = n13058 & n20161 ;
  assign n20163 = n20162 ^ n2262 ^ 1'b0 ;
  assign n20159 = n10282 ^ n2833 ^ 1'b0 ;
  assign n20169 = n20168 ^ n20163 ^ n20159 ;
  assign n20170 = n20169 ^ n2684 ^ n1774 ;
  assign n20171 = ( n146 & n19525 ) | ( n146 & ~n20170 ) | ( n19525 & ~n20170 ) ;
  assign n20172 = n14542 ^ n14111 ^ 1'b0 ;
  assign n20175 = n10275 ^ n2415 ^ 1'b0 ;
  assign n20173 = ~n5764 & n20040 ;
  assign n20174 = n20173 ^ n4438 ^ 1'b0 ;
  assign n20176 = n20175 ^ n20174 ^ 1'b0 ;
  assign n20177 = n18764 ^ n12402 ^ 1'b0 ;
  assign n20178 = ( n1119 & n5198 ) | ( n1119 & ~n6102 ) | ( n5198 & ~n6102 ) ;
  assign n20179 = ( n6805 & n17889 ) | ( n6805 & ~n19319 ) | ( n17889 & ~n19319 ) ;
  assign n20180 = n12630 ^ n9978 ^ n757 ;
  assign n20181 = n20180 ^ n4273 ^ 1'b0 ;
  assign n20182 = ~n4409 & n20181 ;
  assign n20183 = n5818 ^ n939 ^ 1'b0 ;
  assign n20184 = ( n7677 & n20182 ) | ( n7677 & n20183 ) | ( n20182 & n20183 ) ;
  assign n20185 = n7266 ^ n3097 ^ n2682 ;
  assign n20186 = n20185 ^ n16499 ^ 1'b0 ;
  assign n20187 = ~n6244 & n20186 ;
  assign n20188 = n3784 ^ n2178 ^ 1'b0 ;
  assign n20189 = n16494 & ~n20188 ;
  assign n20190 = n14418 ^ n3779 ^ 1'b0 ;
  assign n20191 = n20190 ^ n10749 ^ n9927 ;
  assign n20192 = n965 & n20191 ;
  assign n20193 = ~n20189 & n20192 ;
  assign n20194 = n11508 ^ n4693 ^ 1'b0 ;
  assign n20195 = ( ~n12723 & n13678 ) | ( ~n12723 & n14067 ) | ( n13678 & n14067 ) ;
  assign n20197 = n4906 ^ n4505 ^ 1'b0 ;
  assign n20196 = n16126 ^ n3452 ^ 1'b0 ;
  assign n20198 = n20197 ^ n20196 ^ 1'b0 ;
  assign n20199 = n20198 ^ n12031 ^ 1'b0 ;
  assign n20200 = n1947 | n5473 ;
  assign n20201 = n4591 | n20200 ;
  assign n20202 = n15380 ^ n13141 ^ n8409 ;
  assign n20203 = ( n4259 & n5515 ) | ( n4259 & ~n17725 ) | ( n5515 & ~n17725 ) ;
  assign n20204 = n20202 & ~n20203 ;
  assign n20205 = n20204 ^ n5228 ^ 1'b0 ;
  assign n20213 = n3899 & ~n13104 ;
  assign n20214 = n20213 ^ n15236 ^ 1'b0 ;
  assign n20215 = ( n2677 & n7360 ) | ( n2677 & n20214 ) | ( n7360 & n20214 ) ;
  assign n20209 = n800 & ~n6095 ;
  assign n20210 = ~n3496 & n20209 ;
  assign n20206 = ( n5439 & ~n5757 ) | ( n5439 & n8497 ) | ( ~n5757 & n8497 ) ;
  assign n20207 = n20206 ^ n9905 ^ 1'b0 ;
  assign n20208 = n20207 ^ n13250 ^ 1'b0 ;
  assign n20211 = n20210 ^ n20208 ^ n3646 ;
  assign n20212 = ( n9840 & ~n19655 ) | ( n9840 & n20211 ) | ( ~n19655 & n20211 ) ;
  assign n20216 = n20215 ^ n20212 ^ 1'b0 ;
  assign n20218 = ~n1283 & n2037 ;
  assign n20219 = n20218 ^ n160 ^ 1'b0 ;
  assign n20217 = n3664 & n10770 ;
  assign n20220 = n20219 ^ n20217 ^ n2767 ;
  assign n20221 = n4808 | n11718 ;
  assign n20222 = n20221 ^ n17558 ^ 1'b0 ;
  assign n20223 = n18377 ^ n2209 ^ 1'b0 ;
  assign n20224 = ~n474 & n20223 ;
  assign n20225 = x87 & ~n7644 ;
  assign n20226 = n20225 ^ n189 ^ 1'b0 ;
  assign n20227 = n20226 ^ n10625 ^ 1'b0 ;
  assign n20228 = ~n9767 & n20227 ;
  assign n20229 = n1294 & ~n19040 ;
  assign n20230 = n777 & n20229 ;
  assign n20231 = n20230 ^ n5361 ^ 1'b0 ;
  assign n20232 = n1573 & n20231 ;
  assign n20233 = n20232 ^ n4588 ^ 1'b0 ;
  assign n20234 = n20233 ^ n3516 ^ 1'b0 ;
  assign n20235 = ( n8087 & n8415 ) | ( n8087 & n11159 ) | ( n8415 & n11159 ) ;
  assign n20236 = ( n17531 & n18814 ) | ( n17531 & n20235 ) | ( n18814 & n20235 ) ;
  assign n20239 = n622 & n7122 ;
  assign n20240 = ~n3322 & n20239 ;
  assign n20237 = n11340 ^ n6959 ^ 1'b0 ;
  assign n20238 = n10194 & n20237 ;
  assign n20241 = n20240 ^ n20238 ^ n2570 ;
  assign n20242 = ( n7486 & ~n8186 ) | ( n7486 & n20241 ) | ( ~n8186 & n20241 ) ;
  assign n20243 = n7452 | n18944 ;
  assign n20244 = n20243 ^ n14568 ^ 1'b0 ;
  assign n20245 = n3164 | n4701 ;
  assign n20246 = n20245 ^ n12776 ^ 1'b0 ;
  assign n20247 = n9473 ^ n8056 ^ 1'b0 ;
  assign n20252 = n1980 & ~n15174 ;
  assign n20253 = n20252 ^ n1614 ^ 1'b0 ;
  assign n20248 = ~n5011 & n8852 ;
  assign n20249 = n20248 ^ n9993 ^ 1'b0 ;
  assign n20250 = n3419 & n20249 ;
  assign n20251 = n6094 & n20250 ;
  assign n20254 = n20253 ^ n20251 ^ 1'b0 ;
  assign n20255 = n20247 | n20254 ;
  assign n20256 = n20255 ^ n9808 ^ n4402 ;
  assign n20257 = n14350 ^ n13198 ^ n4562 ;
  assign n20258 = n2743 | n14379 ;
  assign n20259 = n20258 ^ n7340 ^ 1'b0 ;
  assign n20260 = ( x77 & n10304 ) | ( x77 & n12259 ) | ( n10304 & n12259 ) ;
  assign n20261 = n13247 ^ n8525 ^ 1'b0 ;
  assign n20262 = ~n12223 & n20261 ;
  assign n20263 = ~n15643 & n20262 ;
  assign n20264 = ~n20260 & n20263 ;
  assign n20265 = n8510 | n13650 ;
  assign n20266 = ( ~n10124 & n10142 ) | ( ~n10124 & n20265 ) | ( n10142 & n20265 ) ;
  assign n20267 = n1488 | n20266 ;
  assign n20268 = ( n9530 & n11387 ) | ( n9530 & ~n13203 ) | ( n11387 & ~n13203 ) ;
  assign n20269 = ( n10715 & n15100 ) | ( n10715 & n15219 ) | ( n15100 & n15219 ) ;
  assign n20270 = n5431 & ~n20269 ;
  assign n20271 = n20268 & n20270 ;
  assign n20272 = ( n141 & ~n664 ) | ( n141 & n18768 ) | ( ~n664 & n18768 ) ;
  assign n20273 = n1871 ^ n1228 ^ 1'b0 ;
  assign n20274 = n20273 ^ n19629 ^ n8005 ;
  assign n20275 = n20274 ^ n15369 ^ n3044 ;
  assign n20276 = n4641 ^ n2560 ^ 1'b0 ;
  assign n20277 = n15769 & ~n20276 ;
  assign n20278 = n20277 ^ n17878 ^ 1'b0 ;
  assign n20279 = ( n6697 & n13104 ) | ( n6697 & n19860 ) | ( n13104 & n19860 ) ;
  assign n20280 = n11399 & n20279 ;
  assign n20282 = n1270 & n5814 ;
  assign n20281 = n5494 | n13317 ;
  assign n20283 = n20282 ^ n20281 ^ n16507 ;
  assign n20284 = n7955 & n20283 ;
  assign n20285 = n20284 ^ n19620 ^ 1'b0 ;
  assign n20286 = x40 & ~n1227 ;
  assign n20287 = n6017 & n20286 ;
  assign n20288 = ( n1216 & n1617 ) | ( n1216 & ~n1752 ) | ( n1617 & ~n1752 ) ;
  assign n20289 = n20287 | n20288 ;
  assign n20290 = n20210 ^ n16911 ^ 1'b0 ;
  assign n20291 = ( n265 & n413 ) | ( n265 & ~n1897 ) | ( n413 & ~n1897 ) ;
  assign n20292 = n7323 & ~n20291 ;
  assign n20293 = n20292 ^ n8861 ^ 1'b0 ;
  assign n20294 = ~n13141 & n20293 ;
  assign n20295 = n3092 & ~n9267 ;
  assign n20296 = n20295 ^ n5390 ^ 1'b0 ;
  assign n20297 = n3292 | n20296 ;
  assign n20298 = n20297 ^ n2683 ^ 1'b0 ;
  assign n20299 = n16301 & n20298 ;
  assign n20300 = n10575 ^ n8734 ^ 1'b0 ;
  assign n20301 = n8066 ^ n3759 ^ 1'b0 ;
  assign n20302 = n6681 ^ n6516 ^ 1'b0 ;
  assign n20303 = n18547 | n20302 ;
  assign n20304 = n9359 ^ n9210 ^ n4862 ;
  assign n20305 = n20304 ^ n5324 ^ 1'b0 ;
  assign n20306 = n10139 | n20305 ;
  assign n20308 = ( ~n1294 & n7288 ) | ( ~n1294 & n11381 ) | ( n7288 & n11381 ) ;
  assign n20309 = ( ~n3026 & n14698 ) | ( ~n3026 & n20308 ) | ( n14698 & n20308 ) ;
  assign n20307 = n2773 & n5081 ;
  assign n20310 = n20309 ^ n20307 ^ 1'b0 ;
  assign n20311 = n8728 & ~n17967 ;
  assign n20312 = n20311 ^ n4530 ^ 1'b0 ;
  assign n20313 = n18561 ^ n17488 ^ n2136 ;
  assign n20314 = n20313 ^ n16955 ^ n3699 ;
  assign n20315 = n20314 ^ n4041 ^ 1'b0 ;
  assign n20316 = n11418 ^ n9604 ^ n1989 ;
  assign n20317 = ( n992 & n11049 ) | ( n992 & ~n20316 ) | ( n11049 & ~n20316 ) ;
  assign n20318 = n20317 ^ n19537 ^ n5827 ;
  assign n20319 = n9352 ^ n7775 ^ 1'b0 ;
  assign n20320 = n8371 & n20319 ;
  assign n20321 = ( n16854 & n20103 ) | ( n16854 & n20320 ) | ( n20103 & n20320 ) ;
  assign n20322 = n19078 ^ n7598 ^ 1'b0 ;
  assign n20323 = ( ~n9687 & n20321 ) | ( ~n9687 & n20322 ) | ( n20321 & n20322 ) ;
  assign n20325 = n7158 ^ n1883 ^ 1'b0 ;
  assign n20326 = n3301 & ~n20325 ;
  assign n20327 = n20326 ^ n14629 ^ n2069 ;
  assign n20324 = n11341 ^ n8121 ^ 1'b0 ;
  assign n20328 = n20327 ^ n20324 ^ n14206 ;
  assign n20329 = n15542 ^ n5699 ^ n2502 ;
  assign n20330 = n13893 ^ n12652 ^ n9413 ;
  assign n20331 = ( n1038 & ~n3688 ) | ( n1038 & n13046 ) | ( ~n3688 & n13046 ) ;
  assign n20332 = n2342 | n5759 ;
  assign n20333 = n8722 & n20332 ;
  assign n20334 = n6515 & n20333 ;
  assign n20335 = n508 | n13989 ;
  assign n20336 = n11511 | n20335 ;
  assign n20337 = n20309 ^ n9815 ^ n201 ;
  assign n20339 = ( n1890 & n2869 ) | ( n1890 & n12358 ) | ( n2869 & n12358 ) ;
  assign n20338 = n1876 & n11862 ;
  assign n20340 = n20339 ^ n20338 ^ 1'b0 ;
  assign n20341 = n8481 & n9912 ;
  assign n20342 = n1029 & ~n4374 ;
  assign n20343 = n15439 & n20342 ;
  assign n20344 = n20109 ^ n1731 ^ 1'b0 ;
  assign n20345 = n8609 ^ n8389 ^ n256 ;
  assign n20346 = n20345 ^ n17375 ^ 1'b0 ;
  assign n20347 = ~n20344 & n20346 ;
  assign n20348 = n6226 & ~n11029 ;
  assign n20349 = ~n2153 & n3173 ;
  assign n20350 = ~n20348 & n20349 ;
  assign n20351 = ( ~n2607 & n4220 ) | ( ~n2607 & n7861 ) | ( n4220 & n7861 ) ;
  assign n20352 = n15583 ^ n14238 ^ n8151 ;
  assign n20357 = n16071 ^ n2212 ^ 1'b0 ;
  assign n20358 = ~n9631 & n20357 ;
  assign n20359 = ~n12847 & n20358 ;
  assign n20360 = n20359 ^ n1228 ^ 1'b0 ;
  assign n20354 = ( x91 & n2960 ) | ( x91 & ~n10028 ) | ( n2960 & ~n10028 ) ;
  assign n20353 = n8442 & ~n14493 ;
  assign n20355 = n20354 ^ n20353 ^ 1'b0 ;
  assign n20356 = n20355 ^ n14460 ^ n8961 ;
  assign n20361 = n20360 ^ n20356 ^ n15423 ;
  assign n20362 = n20361 ^ n7744 ^ n3724 ;
  assign n20363 = n11557 ^ n5730 ^ 1'b0 ;
  assign n20364 = n17099 ^ n10913 ^ n3962 ;
  assign n20365 = n6286 ^ n3150 ^ 1'b0 ;
  assign n20366 = n831 & ~n20365 ;
  assign n20367 = n632 & n20366 ;
  assign n20368 = n4209 & n4821 ;
  assign n20369 = ~n7302 & n20368 ;
  assign n20370 = n18787 | n20369 ;
  assign n20371 = n20370 ^ n12005 ^ 1'b0 ;
  assign n20372 = ( n14032 & n17711 ) | ( n14032 & ~n20371 ) | ( n17711 & ~n20371 ) ;
  assign n20373 = ( n909 & ~n20367 ) | ( n909 & n20372 ) | ( ~n20367 & n20372 ) ;
  assign n20374 = n17863 ^ n6301 ^ n572 ;
  assign n20375 = ( ~n557 & n3781 ) | ( ~n557 & n6013 ) | ( n3781 & n6013 ) ;
  assign n20376 = n203 & n8875 ;
  assign n20377 = n168 & n20376 ;
  assign n20378 = n20375 | n20377 ;
  assign n20379 = n20374 & ~n20378 ;
  assign n20380 = n15605 | n20208 ;
  assign n20381 = n9048 ^ n5008 ^ n4713 ;
  assign n20382 = n20381 ^ n11062 ^ 1'b0 ;
  assign n20383 = n20380 & n20382 ;
  assign n20384 = n5650 & n12361 ;
  assign n20385 = n20384 ^ n19904 ^ n3839 ;
  assign n20386 = ( n767 & ~n7953 ) | ( n767 & n10182 ) | ( ~n7953 & n10182 ) ;
  assign n20387 = n3337 & n8802 ;
  assign n20388 = ~n15442 & n20387 ;
  assign n20389 = ~n8957 & n20388 ;
  assign n20390 = ( n2057 & n20386 ) | ( n2057 & ~n20389 ) | ( n20386 & ~n20389 ) ;
  assign n20391 = n5444 & n6807 ;
  assign n20392 = n5302 ^ n1496 ^ n1260 ;
  assign n20393 = n15425 ^ n5139 ^ 1'b0 ;
  assign n20394 = n413 & ~n20393 ;
  assign n20395 = n20392 & n20394 ;
  assign n20396 = n20395 ^ n2652 ^ 1'b0 ;
  assign n20397 = ( n2011 & n4182 ) | ( n2011 & ~n4287 ) | ( n4182 & ~n4287 ) ;
  assign n20398 = n20397 ^ n6116 ^ n6056 ;
  assign n20399 = n14697 ^ n5186 ^ 1'b0 ;
  assign n20400 = n9086 & n10809 ;
  assign n20401 = n19537 & n20400 ;
  assign n20402 = n20401 ^ n2656 ^ 1'b0 ;
  assign n20403 = n9458 | n20402 ;
  assign n20404 = ~n6079 & n10058 ;
  assign n20405 = ( n3579 & n11512 ) | ( n3579 & ~n11600 ) | ( n11512 & ~n11600 ) ;
  assign n20407 = n1732 | n7498 ;
  assign n20408 = n6354 | n20407 ;
  assign n20406 = ( n4484 & ~n14706 ) | ( n4484 & n14796 ) | ( ~n14706 & n14796 ) ;
  assign n20409 = n20408 ^ n20406 ^ n12307 ;
  assign n20410 = n2009 & ~n5033 ;
  assign n20411 = n12354 ^ n8885 ^ 1'b0 ;
  assign n20412 = n8111 ^ n1539 ^ 1'b0 ;
  assign n20413 = n20411 | n20412 ;
  assign n20414 = n15414 ^ n2484 ^ 1'b0 ;
  assign n20415 = n1639 & n20414 ;
  assign n20416 = n20415 ^ n8243 ^ 1'b0 ;
  assign n20417 = n18580 | n20416 ;
  assign n20418 = n17498 ^ n11980 ^ 1'b0 ;
  assign n20419 = n20418 ^ n6548 ^ 1'b0 ;
  assign n20420 = n9167 & n20419 ;
  assign n20423 = n8603 ^ n646 ^ 1'b0 ;
  assign n20421 = ( n4482 & n9369 ) | ( n4482 & n16493 ) | ( n9369 & n16493 ) ;
  assign n20422 = n20421 ^ n14029 ^ n3597 ;
  assign n20424 = n20423 ^ n20422 ^ n6971 ;
  assign n20425 = n20424 ^ n17941 ^ 1'b0 ;
  assign n20426 = n1847 & n20425 ;
  assign n20427 = n2510 | n4748 ;
  assign n20428 = n20427 ^ n359 ^ 1'b0 ;
  assign n20429 = ( ~n8183 & n10065 ) | ( ~n8183 & n20428 ) | ( n10065 & n20428 ) ;
  assign n20430 = n20429 ^ n16144 ^ n3269 ;
  assign n20431 = ( ~n4599 & n7158 ) | ( ~n4599 & n10122 ) | ( n7158 & n10122 ) ;
  assign n20436 = ( x46 & ~n2687 ) | ( x46 & n18778 ) | ( ~n2687 & n18778 ) ;
  assign n20432 = n4202 | n6722 ;
  assign n20433 = n12513 & ~n20432 ;
  assign n20434 = n8888 & n15562 ;
  assign n20435 = n20433 & n20434 ;
  assign n20437 = n20436 ^ n20435 ^ n18852 ;
  assign n20438 = n19579 ^ n4146 ^ 1'b0 ;
  assign n20439 = n14454 & ~n20438 ;
  assign n20440 = n11020 ^ n9679 ^ 1'b0 ;
  assign n20441 = ~n1370 & n20440 ;
  assign n20442 = n6220 & ~n9971 ;
  assign n20443 = n18112 ^ n17935 ^ 1'b0 ;
  assign n20444 = n20442 & ~n20443 ;
  assign n20447 = ~n6363 & n12285 ;
  assign n20448 = n20447 ^ n7049 ^ n385 ;
  assign n20445 = n13174 | n16521 ;
  assign n20446 = n20445 ^ n13727 ^ 1'b0 ;
  assign n20449 = n20448 ^ n20446 ^ 1'b0 ;
  assign n20450 = n5530 & n20449 ;
  assign n20451 = n13326 ^ n12706 ^ n3009 ;
  assign n20452 = n14703 & ~n20451 ;
  assign n20453 = n20452 ^ n15998 ^ 1'b0 ;
  assign n20454 = n14526 ^ n8413 ^ n4616 ;
  assign n20455 = n20454 ^ n9719 ^ n1547 ;
  assign n20462 = n14449 ^ n11714 ^ n9191 ;
  assign n20456 = ( n315 & ~n4583 ) | ( n315 & n7347 ) | ( ~n4583 & n7347 ) ;
  assign n20457 = n20456 ^ n20175 ^ n6726 ;
  assign n20458 = n20457 ^ n16515 ^ n1731 ;
  assign n20459 = n6896 & n20458 ;
  assign n20460 = n10307 & ~n20459 ;
  assign n20461 = ~n10979 & n20460 ;
  assign n20463 = n20462 ^ n20461 ^ n4198 ;
  assign n20465 = n5146 | n13256 ;
  assign n20466 = n20465 ^ n840 ^ 1'b0 ;
  assign n20464 = n3007 ^ x115 ^ 1'b0 ;
  assign n20467 = n20466 ^ n20464 ^ n9413 ;
  assign n20468 = n14921 | n18623 ;
  assign n20469 = n4996 | n13255 ;
  assign n20470 = ( n5700 & n6871 ) | ( n5700 & n15041 ) | ( n6871 & n15041 ) ;
  assign n20471 = n1266 | n20470 ;
  assign n20472 = n20471 ^ n3571 ^ 1'b0 ;
  assign n20473 = ( n18676 & n20469 ) | ( n18676 & n20472 ) | ( n20469 & n20472 ) ;
  assign n20474 = n3948 ^ x101 ^ 1'b0 ;
  assign n20475 = ~n19210 & n20474 ;
  assign n20476 = n15865 & n20475 ;
  assign n20477 = ( n1536 & n5070 ) | ( n1536 & ~n11916 ) | ( n5070 & ~n11916 ) ;
  assign n20478 = ~n11905 & n20477 ;
  assign n20479 = ~n5892 & n20478 ;
  assign n20480 = n11430 ^ n1024 ^ 1'b0 ;
  assign n20481 = ~n9039 & n20480 ;
  assign n20482 = ~n6328 & n17035 ;
  assign n20483 = n3220 | n20482 ;
  assign n20484 = n20483 ^ n14412 ^ 1'b0 ;
  assign n20485 = ~n3163 & n16678 ;
  assign n20486 = ~n2801 & n20485 ;
  assign n20487 = ( n15437 & n20484 ) | ( n15437 & n20486 ) | ( n20484 & n20486 ) ;
  assign n20488 = n9834 ^ n243 ^ 1'b0 ;
  assign n20489 = n10024 & n20488 ;
  assign n20490 = n12739 ^ n8841 ^ 1'b0 ;
  assign n20491 = n6801 & ~n20490 ;
  assign n20492 = ( n2847 & n20489 ) | ( n2847 & ~n20491 ) | ( n20489 & ~n20491 ) ;
  assign n20493 = ( n10002 & n10922 ) | ( n10002 & n19625 ) | ( n10922 & n19625 ) ;
  assign n20495 = n2431 & n9709 ;
  assign n20494 = ~n5703 & n12750 ;
  assign n20496 = n20495 ^ n20494 ^ 1'b0 ;
  assign n20497 = n1806 | n20496 ;
  assign n20498 = n20497 ^ n17848 ^ 1'b0 ;
  assign n20499 = n3445 | n5923 ;
  assign n20500 = n3237 & ~n20499 ;
  assign n20501 = n20500 ^ n7073 ^ 1'b0 ;
  assign n20502 = n2546 & n20501 ;
  assign n20503 = n12003 & n20502 ;
  assign n20504 = n20503 ^ n16648 ^ 1'b0 ;
  assign n20513 = n4253 & n6534 ;
  assign n20508 = ~n6585 & n7655 ;
  assign n20509 = n20508 ^ n11475 ^ 1'b0 ;
  assign n20510 = n20509 ^ n9170 ^ n7856 ;
  assign n20511 = ( n324 & n3458 ) | ( n324 & n13486 ) | ( n3458 & n13486 ) ;
  assign n20512 = n20510 | n20511 ;
  assign n20505 = ( n1518 & n5570 ) | ( n1518 & ~n8172 ) | ( n5570 & ~n8172 ) ;
  assign n20506 = n20505 ^ n6670 ^ 1'b0 ;
  assign n20507 = n19906 & ~n20506 ;
  assign n20514 = n20513 ^ n20512 ^ n20507 ;
  assign n20515 = n8967 ^ n4665 ^ 1'b0 ;
  assign n20516 = n20515 ^ n11116 ^ n4361 ;
  assign n20517 = n14227 ^ n8025 ^ n4014 ;
  assign n20518 = n6219 ^ n401 ^ 1'b0 ;
  assign n20519 = ~n11519 & n20518 ;
  assign n20520 = ( n11980 & n20517 ) | ( n11980 & ~n20519 ) | ( n20517 & ~n20519 ) ;
  assign n20521 = n20516 | n20520 ;
  assign n20522 = n20313 ^ n9259 ^ n5112 ;
  assign n20523 = ( n214 & n1079 ) | ( n214 & ~n10361 ) | ( n1079 & ~n10361 ) ;
  assign n20524 = ( n6574 & ~n9304 ) | ( n6574 & n20523 ) | ( ~n9304 & n20523 ) ;
  assign n20525 = n11888 ^ n3528 ^ 1'b0 ;
  assign n20526 = ~n1715 & n20525 ;
  assign n20527 = n20526 ^ n12494 ^ 1'b0 ;
  assign n20528 = n10374 ^ n4920 ^ n1331 ;
  assign n20529 = n20528 ^ n14021 ^ 1'b0 ;
  assign n20530 = ( n5927 & n6579 ) | ( n5927 & n13318 ) | ( n6579 & n13318 ) ;
  assign n20532 = n11733 ^ n8284 ^ n7685 ;
  assign n20531 = ( n1958 & n4759 ) | ( n1958 & n5133 ) | ( n4759 & n5133 ) ;
  assign n20533 = n20532 ^ n20531 ^ n15913 ;
  assign n20534 = n3696 | n16941 ;
  assign n20535 = n370 | n20534 ;
  assign n20536 = ( n150 & ~n12334 ) | ( n150 & n20535 ) | ( ~n12334 & n20535 ) ;
  assign n20537 = n13739 ^ n8206 ^ 1'b0 ;
  assign n20538 = n20537 ^ n17717 ^ 1'b0 ;
  assign n20539 = n3807 | n20538 ;
  assign n20540 = n20536 | n20539 ;
  assign n20541 = ( n5111 & ~n14840 ) | ( n5111 & n20540 ) | ( ~n14840 & n20540 ) ;
  assign n20544 = n3647 | n8987 ;
  assign n20542 = n9832 & ~n16953 ;
  assign n20543 = n20542 ^ n12374 ^ 1'b0 ;
  assign n20545 = n20544 ^ n20543 ^ 1'b0 ;
  assign n20546 = n3496 & n6007 ;
  assign n20547 = n11747 & n20546 ;
  assign n20548 = ( n2218 & ~n9105 ) | ( n2218 & n20547 ) | ( ~n9105 & n20547 ) ;
  assign n20549 = n4973 & ~n20548 ;
  assign n20550 = n20549 ^ n2282 ^ 1'b0 ;
  assign n20551 = n9856 ^ n1563 ^ n566 ;
  assign n20552 = ~n9219 & n20551 ;
  assign n20553 = ~n19992 & n20552 ;
  assign n20554 = n368 & ~n9220 ;
  assign n20555 = ~n912 & n20554 ;
  assign n20556 = ~n1486 & n2884 ;
  assign n20557 = n20556 ^ n5390 ^ 1'b0 ;
  assign n20558 = n976 & n20557 ;
  assign n20559 = n18480 & n20558 ;
  assign n20560 = ~n503 & n10487 ;
  assign n20561 = n20560 ^ n16938 ^ 1'b0 ;
  assign n20562 = ( n2839 & n5011 ) | ( n2839 & n20561 ) | ( n5011 & n20561 ) ;
  assign n20563 = ( ~n20555 & n20559 ) | ( ~n20555 & n20562 ) | ( n20559 & n20562 ) ;
  assign n20564 = ( ~n6288 & n15140 ) | ( ~n6288 & n18251 ) | ( n15140 & n18251 ) ;
  assign n20565 = ( n2913 & n4159 ) | ( n2913 & ~n20564 ) | ( n4159 & ~n20564 ) ;
  assign n20566 = n17900 ^ n2174 ^ 1'b0 ;
  assign n20567 = n20484 ^ n6418 ^ n4409 ;
  assign n20568 = n20567 ^ n896 ^ 1'b0 ;
  assign n20569 = ~n15635 & n20568 ;
  assign n20570 = n5023 ^ n1029 ^ 1'b0 ;
  assign n20571 = n2089 | n20570 ;
  assign n20575 = ( n3681 & ~n3902 ) | ( n3681 & n10321 ) | ( ~n3902 & n10321 ) ;
  assign n20572 = n4377 & n5089 ;
  assign n20573 = n20572 ^ n17560 ^ 1'b0 ;
  assign n20574 = n20573 ^ n16300 ^ n6984 ;
  assign n20576 = n20575 ^ n20574 ^ n3537 ;
  assign n20577 = n20576 ^ n19750 ^ n3318 ;
  assign n20578 = n20577 ^ n16647 ^ 1'b0 ;
  assign n20579 = n9821 ^ n7402 ^ n1523 ;
  assign n20580 = n9577 ^ n6865 ^ n1758 ;
  assign n20582 = n5248 ^ n4333 ^ 1'b0 ;
  assign n20583 = ~n13055 & n20582 ;
  assign n20581 = n9781 & n12746 ;
  assign n20584 = n20583 ^ n20581 ^ 1'b0 ;
  assign n20585 = n10645 ^ n4322 ^ n1297 ;
  assign n20586 = n20585 ^ n4954 ^ n3356 ;
  assign n20587 = n20584 | n20586 ;
  assign n20588 = n13338 ^ n10709 ^ 1'b0 ;
  assign n20589 = ~n360 & n20588 ;
  assign n20590 = n20589 ^ n14846 ^ n9953 ;
  assign n20591 = ( ~n1728 & n7479 ) | ( ~n1728 & n15318 ) | ( n7479 & n15318 ) ;
  assign n20592 = n5505 ^ n3977 ^ 1'b0 ;
  assign n20593 = ( n4165 & n11184 ) | ( n4165 & ~n20592 ) | ( n11184 & ~n20592 ) ;
  assign n20594 = n7142 ^ n236 ^ 1'b0 ;
  assign n20595 = n2334 & n20594 ;
  assign n20596 = n2020 & ~n8595 ;
  assign n20597 = n8521 & n20596 ;
  assign n20598 = ( n726 & n4460 ) | ( n726 & n20597 ) | ( n4460 & n20597 ) ;
  assign n20599 = n10035 ^ n3977 ^ 1'b0 ;
  assign n20600 = n20598 & n20599 ;
  assign n20601 = n639 ^ n434 ^ 1'b0 ;
  assign n20602 = n20601 ^ n8738 ^ 1'b0 ;
  assign n20603 = n20600 & ~n20602 ;
  assign n20604 = ( n2534 & n9497 ) | ( n2534 & n17086 ) | ( n9497 & n17086 ) ;
  assign n20605 = n20604 ^ n11958 ^ 1'b0 ;
  assign n20606 = n11101 & ~n20605 ;
  assign n20607 = n20606 ^ n5078 ^ 1'b0 ;
  assign n20608 = n20603 & ~n20607 ;
  assign n20612 = n2317 | n7165 ;
  assign n20613 = n20612 ^ n5196 ^ n1665 ;
  assign n20609 = n18912 ^ n10429 ^ 1'b0 ;
  assign n20610 = n6751 & ~n20609 ;
  assign n20611 = n20610 ^ n9963 ^ 1'b0 ;
  assign n20614 = n20613 ^ n20611 ^ n5232 ;
  assign n20615 = ( n2938 & n4604 ) | ( n2938 & n20614 ) | ( n4604 & n20614 ) ;
  assign n20616 = n20615 ^ n12311 ^ n8640 ;
  assign n20617 = ( n5798 & n11068 ) | ( n5798 & ~n16270 ) | ( n11068 & ~n16270 ) ;
  assign n20618 = n15726 & n20617 ;
  assign n20619 = ~n6382 & n6987 ;
  assign n20620 = n20619 ^ n14090 ^ 1'b0 ;
  assign n20621 = n7696 & n7703 ;
  assign n20622 = n1424 & n20621 ;
  assign n20623 = n20622 ^ n5158 ^ 1'b0 ;
  assign n20624 = n20623 ^ n15010 ^ n2170 ;
  assign n20625 = n2946 ^ n866 ^ 1'b0 ;
  assign n20626 = n11368 & ~n20625 ;
  assign n20627 = n20626 ^ n11661 ^ 1'b0 ;
  assign n20628 = n20627 ^ n3626 ^ n2323 ;
  assign n20629 = n20628 ^ n16898 ^ n2565 ;
  assign n20630 = ( n20620 & n20624 ) | ( n20620 & n20629 ) | ( n20624 & n20629 ) ;
  assign n20631 = ( n4293 & n6627 ) | ( n4293 & n19165 ) | ( n6627 & n19165 ) ;
  assign n20632 = n3149 ^ n3101 ^ 1'b0 ;
  assign n20633 = n20632 ^ n3567 ^ 1'b0 ;
  assign n20634 = ~n11980 & n16617 ;
  assign n20635 = n20634 ^ n7235 ^ 1'b0 ;
  assign n20636 = n8478 ^ n7299 ^ 1'b0 ;
  assign n20637 = ~n9798 & n20636 ;
  assign n20638 = ~n631 & n20637 ;
  assign n20639 = n2424 ^ n1749 ^ n556 ;
  assign n20640 = n10896 ^ n6073 ^ 1'b0 ;
  assign n20641 = n8140 & ~n9353 ;
  assign n20642 = n20641 ^ n9272 ^ 1'b0 ;
  assign n20643 = n18143 ^ n17182 ^ n15909 ;
  assign n20644 = ~n853 & n2075 ;
  assign n20645 = ~x101 & n20644 ;
  assign n20646 = n1390 | n7418 ;
  assign n20647 = n15492 & ~n20646 ;
  assign n20648 = ~n1379 & n3726 ;
  assign n20649 = n20648 ^ n3797 ^ 1'b0 ;
  assign n20650 = n14976 & n20649 ;
  assign n20651 = ( x93 & n5416 ) | ( x93 & ~n20650 ) | ( n5416 & ~n20650 ) ;
  assign n20652 = ( ~n12827 & n20647 ) | ( ~n12827 & n20651 ) | ( n20647 & n20651 ) ;
  assign n20653 = ~n20645 & n20652 ;
  assign n20654 = n20653 ^ n10111 ^ 1'b0 ;
  assign n20655 = ~n3514 & n14442 ;
  assign n20656 = n2803 & n20655 ;
  assign n20657 = n5597 ^ n3041 ^ n1280 ;
  assign n20658 = ( ~n4006 & n6691 ) | ( ~n4006 & n9299 ) | ( n6691 & n9299 ) ;
  assign n20659 = ~n11582 & n12661 ;
  assign n20660 = n20659 ^ x77 ^ 1'b0 ;
  assign n20661 = n20660 ^ n1688 ^ n1479 ;
  assign n20662 = n231 & n20661 ;
  assign n20663 = n17432 ^ n12322 ^ n11846 ;
  assign n20664 = n15920 ^ n12357 ^ n6595 ;
  assign n20665 = n7511 | n17984 ;
  assign n20666 = ( ~n20663 & n20664 ) | ( ~n20663 & n20665 ) | ( n20664 & n20665 ) ;
  assign n20667 = n2900 & ~n12582 ;
  assign n20668 = n20667 ^ n184 ^ 1'b0 ;
  assign n20674 = n8156 ^ n5971 ^ n1063 ;
  assign n20669 = ( n1769 & n3599 ) | ( n1769 & ~n9053 ) | ( n3599 & ~n9053 ) ;
  assign n20670 = n20669 ^ n13802 ^ n1600 ;
  assign n20671 = n12203 ^ n4381 ^ n2697 ;
  assign n20672 = n4432 & ~n20671 ;
  assign n20673 = ( n3046 & n20670 ) | ( n3046 & n20672 ) | ( n20670 & n20672 ) ;
  assign n20675 = n20674 ^ n20673 ^ 1'b0 ;
  assign n20676 = ~n3713 & n6354 ;
  assign n20677 = n20676 ^ n5421 ^ 1'b0 ;
  assign n20678 = n2088 | n8028 ;
  assign n20679 = n3537 & ~n20678 ;
  assign n20680 = ~n3819 & n20679 ;
  assign n20681 = n20680 ^ n1455 ^ 1'b0 ;
  assign n20682 = ( n8379 & ~n20677 ) | ( n8379 & n20681 ) | ( ~n20677 & n20681 ) ;
  assign n20683 = ( ~n4835 & n5490 ) | ( ~n4835 & n17651 ) | ( n5490 & n17651 ) ;
  assign n20684 = ( n931 & ~n1608 ) | ( n931 & n13493 ) | ( ~n1608 & n13493 ) ;
  assign n20685 = ~n6815 & n9954 ;
  assign n20688 = n4409 ^ n2843 ^ n580 ;
  assign n20686 = n5427 & ~n7034 ;
  assign n20687 = n13281 | n20686 ;
  assign n20689 = n20688 ^ n20687 ^ 1'b0 ;
  assign n20690 = n2486 | n20689 ;
  assign n20691 = n20685 & ~n20690 ;
  assign n20692 = ( n3362 & n3651 ) | ( n3362 & ~n6256 ) | ( n3651 & ~n6256 ) ;
  assign n20693 = n20692 ^ n1648 ^ 1'b0 ;
  assign n20694 = n13229 | n20693 ;
  assign n20695 = n2835 ^ n1612 ^ n184 ;
  assign n20696 = n20695 ^ n20567 ^ n1683 ;
  assign n20697 = n18316 ^ n17261 ^ 1'b0 ;
  assign n20698 = n19384 ^ n16809 ^ n4736 ;
  assign n20699 = ~n738 & n2051 ;
  assign n20700 = n3556 ^ n3491 ^ n3319 ;
  assign n20701 = ( n648 & n6673 ) | ( n648 & n20700 ) | ( n6673 & n20700 ) ;
  assign n20702 = n1189 | n2712 ;
  assign n20703 = ~n2875 & n20702 ;
  assign n20704 = n20701 & n20703 ;
  assign n20705 = n14168 ^ n1624 ^ 1'b0 ;
  assign n20706 = ( n5144 & ~n16691 ) | ( n5144 & n20705 ) | ( ~n16691 & n20705 ) ;
  assign n20707 = ( n3014 & n11019 ) | ( n3014 & n17267 ) | ( n11019 & n17267 ) ;
  assign n20708 = n20707 ^ n1024 ^ 1'b0 ;
  assign n20709 = n1830 ^ n1779 ^ n302 ;
  assign n20710 = n18644 ^ n14577 ^ n2704 ;
  assign n20711 = n20710 ^ n12533 ^ n11669 ;
  assign n20712 = n4755 & n20711 ;
  assign n20713 = n20712 ^ n9822 ^ 1'b0 ;
  assign n20714 = ( n6482 & ~n20709 ) | ( n6482 & n20713 ) | ( ~n20709 & n20713 ) ;
  assign n20715 = n20714 ^ n5393 ^ n518 ;
  assign n20716 = n5589 ^ n2951 ^ 1'b0 ;
  assign n20717 = n3195 & n20716 ;
  assign n20718 = n8615 & n20717 ;
  assign n20719 = n5083 & n8275 ;
  assign n20720 = n20719 ^ n14643 ^ 1'b0 ;
  assign n20721 = n16362 ^ n15760 ^ 1'b0 ;
  assign n20722 = n19001 & n19030 ;
  assign n20723 = n20722 ^ n4501 ^ 1'b0 ;
  assign n20724 = ( n1091 & n3835 ) | ( n1091 & n6308 ) | ( n3835 & n6308 ) ;
  assign n20725 = n20724 ^ n11276 ^ 1'b0 ;
  assign n20726 = ( ~n12977 & n13295 ) | ( ~n12977 & n20725 ) | ( n13295 & n20725 ) ;
  assign n20729 = n7575 & ~n19937 ;
  assign n20730 = ~n8391 & n20729 ;
  assign n20731 = ( n7496 & n18448 ) | ( n7496 & n20730 ) | ( n18448 & n20730 ) ;
  assign n20727 = n16295 ^ n4106 ^ 1'b0 ;
  assign n20728 = n4611 | n20727 ;
  assign n20732 = n20731 ^ n20728 ^ 1'b0 ;
  assign n20737 = ~n159 & n7444 ;
  assign n20738 = ( x107 & n1940 ) | ( x107 & ~n20737 ) | ( n1940 & ~n20737 ) ;
  assign n20733 = ~n5385 & n11263 ;
  assign n20734 = n20733 ^ n2269 ^ 1'b0 ;
  assign n20735 = ~n7274 & n12694 ;
  assign n20736 = n20734 & n20735 ;
  assign n20739 = n20738 ^ n20736 ^ n16924 ;
  assign n20740 = ( n3242 & ~n3671 ) | ( n3242 & n20739 ) | ( ~n3671 & n20739 ) ;
  assign n20741 = n10920 ^ n1908 ^ n582 ;
  assign n20742 = n317 & n378 ;
  assign n20743 = ( n5763 & n9282 ) | ( n5763 & ~n12298 ) | ( n9282 & ~n12298 ) ;
  assign n20744 = n3759 & n20743 ;
  assign n20745 = ( n847 & n3691 ) | ( n847 & n20744 ) | ( n3691 & n20744 ) ;
  assign n20746 = ( n2524 & ~n20742 ) | ( n2524 & n20745 ) | ( ~n20742 & n20745 ) ;
  assign n20747 = ( n839 & n1016 ) | ( n839 & ~n14055 ) | ( n1016 & ~n14055 ) ;
  assign n20748 = n10434 & n19333 ;
  assign n20750 = x111 & ~n7898 ;
  assign n20751 = ~n1347 & n20750 ;
  assign n20749 = n544 | n4172 ;
  assign n20752 = n20751 ^ n20749 ^ n10758 ;
  assign n20753 = ~n20748 & n20752 ;
  assign n20755 = n6555 ^ n2211 ^ n1214 ;
  assign n20756 = ~n3562 & n20755 ;
  assign n20757 = ~n4018 & n20756 ;
  assign n20758 = n10716 ^ n8914 ^ 1'b0 ;
  assign n20759 = ~n20757 & n20758 ;
  assign n20761 = n3779 & ~n6361 ;
  assign n20760 = n6223 & ~n9352 ;
  assign n20762 = n20761 ^ n20760 ^ 1'b0 ;
  assign n20763 = n20759 & n20762 ;
  assign n20754 = n4471 | n5751 ;
  assign n20764 = n20763 ^ n20754 ^ 1'b0 ;
  assign n20765 = ~n2876 & n20764 ;
  assign n20766 = ~n1019 & n2195 ;
  assign n20767 = n1298 & n20766 ;
  assign n20768 = n4406 & ~n20767 ;
  assign n20769 = n20768 ^ n373 ^ 1'b0 ;
  assign n20770 = n20377 ^ n18283 ^ 1'b0 ;
  assign n20771 = n20770 ^ n16577 ^ 1'b0 ;
  assign n20772 = n20625 ^ n7858 ^ 1'b0 ;
  assign n20773 = ( n15340 & ~n18406 ) | ( n15340 & n19862 ) | ( ~n18406 & n19862 ) ;
  assign n20777 = ( n13533 & n15805 ) | ( n13533 & n20047 ) | ( n15805 & n20047 ) ;
  assign n20774 = n7289 ^ n6941 ^ n2799 ;
  assign n20775 = ( n8206 & ~n12339 ) | ( n8206 & n20774 ) | ( ~n12339 & n20774 ) ;
  assign n20776 = n20775 ^ n11315 ^ n3791 ;
  assign n20778 = n20777 ^ n20776 ^ 1'b0 ;
  assign n20779 = n1349 ^ n1180 ^ 1'b0 ;
  assign n20780 = n3273 & ~n20779 ;
  assign n20783 = ( n7291 & ~n12571 ) | ( n7291 & n19893 ) | ( ~n12571 & n19893 ) ;
  assign n20784 = n10596 & n20783 ;
  assign n20785 = ~n10695 & n20784 ;
  assign n20781 = ~n3273 & n6914 ;
  assign n20782 = n4505 | n20781 ;
  assign n20786 = n20785 ^ n20782 ^ 1'b0 ;
  assign n20787 = n12118 ^ n2982 ^ n250 ;
  assign n20788 = n939 & n6079 ;
  assign n20789 = n20788 ^ n15073 ^ 1'b0 ;
  assign n20790 = n20789 ^ n15408 ^ n5552 ;
  assign n20791 = n20790 ^ n7748 ^ 1'b0 ;
  assign n20792 = n20787 | n20791 ;
  assign n20793 = n8795 & n14211 ;
  assign n20794 = n20161 ^ n786 ^ 1'b0 ;
  assign n20795 = n10291 ^ n7737 ^ n969 ;
  assign n20796 = n20795 ^ n11400 ^ 1'b0 ;
  assign n20797 = ~n7250 & n20796 ;
  assign n20798 = ( n10822 & n20021 ) | ( n10822 & n20797 ) | ( n20021 & n20797 ) ;
  assign n20799 = ( n20793 & ~n20794 ) | ( n20793 & n20798 ) | ( ~n20794 & n20798 ) ;
  assign n20800 = ( ~n637 & n4547 ) | ( ~n637 & n9356 ) | ( n4547 & n9356 ) ;
  assign n20801 = ( ~n1796 & n8738 ) | ( ~n1796 & n20800 ) | ( n8738 & n20800 ) ;
  assign n20802 = n20801 ^ n18948 ^ n4265 ;
  assign n20803 = n11297 & ~n13200 ;
  assign n20804 = ~n20802 & n20803 ;
  assign n20805 = n7932 & n9638 ;
  assign n20807 = n17011 ^ n329 ^ 1'b0 ;
  assign n20806 = ( ~n1225 & n7812 ) | ( ~n1225 & n12503 ) | ( n7812 & n12503 ) ;
  assign n20808 = n20807 ^ n20806 ^ 1'b0 ;
  assign n20809 = n985 & ~n5837 ;
  assign n20810 = n20809 ^ n2882 ^ 1'b0 ;
  assign n20811 = n20810 ^ n19792 ^ n11468 ;
  assign n20812 = n20811 ^ n17049 ^ n4758 ;
  assign n20813 = n10530 & n13914 ;
  assign n20814 = n6214 & n20813 ;
  assign n20815 = n20814 ^ n3206 ^ 1'b0 ;
  assign n20816 = n14384 ^ n13676 ^ 1'b0 ;
  assign n20817 = n16636 | n20816 ;
  assign n20818 = n13457 ^ n10551 ^ 1'b0 ;
  assign n20819 = ~n20817 & n20818 ;
  assign n20820 = ~n740 & n13295 ;
  assign n20821 = n20820 ^ n19907 ^ 1'b0 ;
  assign n20822 = n20418 & n20821 ;
  assign n20823 = n6194 & ~n19969 ;
  assign n20824 = ~x82 & n20823 ;
  assign n20825 = n4216 & n4500 ;
  assign n20826 = n13885 | n20825 ;
  assign n20827 = ( n2259 & n6356 ) | ( n2259 & ~n6693 ) | ( n6356 & ~n6693 ) ;
  assign n20828 = n17739 ^ n10994 ^ 1'b0 ;
  assign n20829 = n1066 & ~n4332 ;
  assign n20830 = n7627 & n20829 ;
  assign n20831 = n1836 | n20830 ;
  assign n20832 = n19068 ^ n11346 ^ 1'b0 ;
  assign n20833 = n9272 ^ n5150 ^ 1'b0 ;
  assign n20834 = ( n8337 & ~n20645 ) | ( n8337 & n20833 ) | ( ~n20645 & n20833 ) ;
  assign n20835 = n20832 & ~n20834 ;
  assign n20836 = n14959 ^ n150 ^ 1'b0 ;
  assign n20837 = n3807 | n20836 ;
  assign n20838 = n381 & n20354 ;
  assign n20843 = n3085 | n9142 ;
  assign n20844 = n20843 ^ n10655 ^ 1'b0 ;
  assign n20841 = n13238 ^ n5805 ^ 1'b0 ;
  assign n20842 = n20841 ^ n18402 ^ 1'b0 ;
  assign n20839 = n14128 ^ n9110 ^ 1'b0 ;
  assign n20840 = n3334 | n20839 ;
  assign n20845 = n20844 ^ n20842 ^ n20840 ;
  assign n20846 = n7965 ^ n3561 ^ n1163 ;
  assign n20847 = n20846 ^ n13152 ^ 1'b0 ;
  assign n20848 = n9167 ^ n5585 ^ n1720 ;
  assign n20849 = n14227 & ~n20848 ;
  assign n20850 = n9082 ^ n4187 ^ x36 ;
  assign n20855 = ( n4141 & n8498 ) | ( n4141 & n14294 ) | ( n8498 & n14294 ) ;
  assign n20851 = ~n4397 & n6310 ;
  assign n20852 = n20851 ^ n4898 ^ 1'b0 ;
  assign n20853 = n20852 ^ n13723 ^ 1'b0 ;
  assign n20854 = n606 | n20853 ;
  assign n20856 = n20855 ^ n20854 ^ n13501 ;
  assign n20857 = n7128 ^ n3369 ^ n1654 ;
  assign n20858 = n9561 & ~n19352 ;
  assign n20859 = n20858 ^ n17558 ^ 1'b0 ;
  assign n20860 = n20859 ^ n3784 ^ n1234 ;
  assign n20863 = n8314 ^ n6059 ^ 1'b0 ;
  assign n20864 = n159 | n20863 ;
  assign n20861 = n6942 ^ n4339 ^ n2087 ;
  assign n20862 = ( n309 & ~n2794 ) | ( n309 & n20861 ) | ( ~n2794 & n20861 ) ;
  assign n20865 = n20864 ^ n20862 ^ n20149 ;
  assign n20866 = n8975 ^ n1923 ^ 1'b0 ;
  assign n20867 = n14387 & ~n20866 ;
  assign n20868 = n20867 ^ n10593 ^ n6170 ;
  assign n20869 = n20868 ^ n9078 ^ n1286 ;
  assign n20871 = n6253 & ~n9016 ;
  assign n20872 = n4522 & ~n20871 ;
  assign n20873 = n20871 & n20872 ;
  assign n20870 = n15569 & ~n19906 ;
  assign n20874 = n20873 ^ n20870 ^ 1'b0 ;
  assign n20875 = ( n17213 & ~n17387 ) | ( n17213 & n20874 ) | ( ~n17387 & n20874 ) ;
  assign n20876 = n10074 ^ n6081 ^ 1'b0 ;
  assign n20877 = n15900 ^ n13112 ^ n2734 ;
  assign n20879 = ( n674 & ~n2973 ) | ( n674 & n2980 ) | ( ~n2973 & n2980 ) ;
  assign n20878 = n7011 ^ n1205 ^ n394 ;
  assign n20880 = n20879 ^ n20878 ^ 1'b0 ;
  assign n20881 = ~n20877 & n20880 ;
  assign n20882 = n20881 ^ n18359 ^ n4622 ;
  assign n20883 = n18782 ^ n13414 ^ n9117 ;
  assign n20884 = ( n8915 & ~n16273 ) | ( n8915 & n20883 ) | ( ~n16273 & n20883 ) ;
  assign n20885 = n1486 ^ n926 ^ 1'b0 ;
  assign n20886 = ( n8545 & n10889 ) | ( n8545 & n14134 ) | ( n10889 & n14134 ) ;
  assign n20887 = x19 | n4578 ;
  assign n20888 = n20887 ^ n12313 ^ 1'b0 ;
  assign n20889 = n20886 & n20888 ;
  assign n20890 = n1715 | n1933 ;
  assign n20891 = n774 & ~n20890 ;
  assign n20892 = ( n9115 & n15815 ) | ( n9115 & ~n20891 ) | ( n15815 & ~n20891 ) ;
  assign n20893 = n20892 ^ n3902 ^ 1'b0 ;
  assign n20894 = n14376 ^ n4191 ^ 1'b0 ;
  assign n20895 = n317 & ~n20894 ;
  assign n20896 = n14893 ^ n13821 ^ 1'b0 ;
  assign n20897 = n15744 & n20896 ;
  assign n20898 = n20897 ^ n17921 ^ 1'b0 ;
  assign n20899 = n7511 & n12598 ;
  assign n20900 = n20899 ^ n9559 ^ 1'b0 ;
  assign n20901 = ( ~n1522 & n5766 ) | ( ~n1522 & n15153 ) | ( n5766 & n15153 ) ;
  assign n20902 = ( ~n8918 & n20900 ) | ( ~n8918 & n20901 ) | ( n20900 & n20901 ) ;
  assign n20903 = n11500 & ~n20902 ;
  assign n20904 = n20903 ^ n3428 ^ 1'b0 ;
  assign n20905 = n4421 ^ n3411 ^ 1'b0 ;
  assign n20906 = n20905 ^ n3728 ^ n405 ;
  assign n20907 = n3325 & ~n20906 ;
  assign n20909 = ( n747 & n2491 ) | ( n747 & n3021 ) | ( n2491 & n3021 ) ;
  assign n20908 = ~n305 & n8511 ;
  assign n20910 = n20909 ^ n20908 ^ 1'b0 ;
  assign n20911 = n12819 | n19716 ;
  assign n20912 = ~n5234 & n20911 ;
  assign n20913 = n15618 ^ n6938 ^ n4443 ;
  assign n20916 = n10067 ^ n5647 ^ 1'b0 ;
  assign n20914 = n3760 & ~n17520 ;
  assign n20915 = n20914 ^ n12656 ^ 1'b0 ;
  assign n20917 = n20916 ^ n20915 ^ n3215 ;
  assign n20918 = n6123 & ~n15120 ;
  assign n20919 = n20918 ^ n15800 ^ n13321 ;
  assign n20920 = ( n4951 & n11315 ) | ( n4951 & ~n20919 ) | ( n11315 & ~n20919 ) ;
  assign n20921 = ( ~n1711 & n7151 ) | ( ~n1711 & n7562 ) | ( n7151 & n7562 ) ;
  assign n20922 = n20921 ^ n11083 ^ n2361 ;
  assign n20924 = ( ~n415 & n957 ) | ( ~n415 & n12905 ) | ( n957 & n12905 ) ;
  assign n20923 = ~n2818 & n18375 ;
  assign n20925 = n20924 ^ n20923 ^ 1'b0 ;
  assign n20926 = n20925 ^ n17084 ^ n6881 ;
  assign n20927 = n12180 & ~n20926 ;
  assign n20928 = ( ~n3159 & n4414 ) | ( ~n3159 & n5772 ) | ( n4414 & n5772 ) ;
  assign n20929 = n20928 ^ n3474 ^ 1'b0 ;
  assign n20930 = ~n7498 & n20929 ;
  assign n20931 = ( ~n7093 & n8817 ) | ( ~n7093 & n18069 ) | ( n8817 & n18069 ) ;
  assign n20932 = ( n3352 & n18365 ) | ( n3352 & ~n20931 ) | ( n18365 & ~n20931 ) ;
  assign n20933 = n5485 | n7347 ;
  assign n20934 = n8369 & ~n20933 ;
  assign n20935 = ( n890 & ~n2078 ) | ( n890 & n20934 ) | ( ~n2078 & n20934 ) ;
  assign n20936 = ( ~n3468 & n4390 ) | ( ~n3468 & n17005 ) | ( n4390 & n17005 ) ;
  assign n20937 = ( n1330 & ~n2254 ) | ( n1330 & n15345 ) | ( ~n2254 & n15345 ) ;
  assign n20938 = ~n8642 & n20937 ;
  assign n20939 = n743 | n7741 ;
  assign n20942 = n4989 & n9168 ;
  assign n20943 = n2924 & ~n20942 ;
  assign n20940 = n1028 & ~n18517 ;
  assign n20941 = n11414 | n20940 ;
  assign n20944 = n20943 ^ n20941 ^ 1'b0 ;
  assign n20947 = n9994 & n12890 ;
  assign n20948 = ~n13310 & n20947 ;
  assign n20945 = n3338 | n8817 ;
  assign n20946 = ~n9318 & n20945 ;
  assign n20949 = n20948 ^ n20946 ^ 1'b0 ;
  assign n20950 = n7848 | n19436 ;
  assign n20951 = n11857 | n20950 ;
  assign n20952 = n4684 & ~n20951 ;
  assign n20953 = ( n8782 & ~n14754 ) | ( n8782 & n20952 ) | ( ~n14754 & n20952 ) ;
  assign n20954 = n18099 ^ n12776 ^ n790 ;
  assign n20955 = n11133 ^ n7236 ^ n3744 ;
  assign n20956 = n18614 | n20955 ;
  assign n20957 = n9290 ^ n1956 ^ 1'b0 ;
  assign n20958 = ~n142 & n4651 ;
  assign n20959 = n3341 & n20958 ;
  assign n20960 = n8754 & ~n11779 ;
  assign n20961 = n20960 ^ n871 ^ 1'b0 ;
  assign n20962 = ~n1289 & n5709 ;
  assign n20963 = ( n5064 & n6430 ) | ( n5064 & n13702 ) | ( n6430 & n13702 ) ;
  assign n20964 = n12129 & ~n14846 ;
  assign n20965 = n20964 ^ n9107 ^ n1387 ;
  assign n20966 = ~x86 & n413 ;
  assign n20967 = ( n10626 & ~n13563 ) | ( n10626 & n20966 ) | ( ~n13563 & n20966 ) ;
  assign n20968 = n20919 & n20967 ;
  assign n20969 = n20968 ^ n2016 ^ 1'b0 ;
  assign n20970 = n4650 ^ n2788 ^ n1831 ;
  assign n20971 = n438 | n3743 ;
  assign n20972 = n20971 ^ n18365 ^ n8071 ;
  assign n20973 = ~n20970 & n20972 ;
  assign n20974 = n20858 & n20973 ;
  assign n20975 = ( n6069 & n7715 ) | ( n6069 & n7911 ) | ( n7715 & n7911 ) ;
  assign n20976 = ( n4022 & n4164 ) | ( n4022 & ~n20975 ) | ( n4164 & ~n20975 ) ;
  assign n20977 = n2520 | n7762 ;
  assign n20978 = n20976 | n20977 ;
  assign n20979 = ( ~n8479 & n8603 ) | ( ~n8479 & n12412 ) | ( n8603 & n12412 ) ;
  assign n20980 = n10756 ^ n4558 ^ 1'b0 ;
  assign n20981 = ~n8076 & n19906 ;
  assign n20982 = ( n1530 & n15888 ) | ( n1530 & ~n19654 ) | ( n15888 & ~n19654 ) ;
  assign n20983 = n20982 ^ n10726 ^ n664 ;
  assign n20984 = ( ~n2314 & n3705 ) | ( ~n2314 & n8870 ) | ( n3705 & n8870 ) ;
  assign n20985 = n20175 ^ n11246 ^ 1'b0 ;
  assign n20986 = n20985 ^ n20854 ^ n16704 ;
  assign n20987 = ( ~n1084 & n1654 ) | ( ~n1084 & n8292 ) | ( n1654 & n8292 ) ;
  assign n20988 = n8766 ^ n3412 ^ 1'b0 ;
  assign n20989 = ( n9461 & n20987 ) | ( n9461 & ~n20988 ) | ( n20987 & ~n20988 ) ;
  assign n20990 = ( n3841 & n10677 ) | ( n3841 & ~n16724 ) | ( n10677 & ~n16724 ) ;
  assign n20991 = n20990 ^ n8472 ^ n6176 ;
  assign n20992 = n20989 & n20991 ;
  assign n20993 = n8240 | n15451 ;
  assign n20994 = ( n11051 & n13813 ) | ( n11051 & n20993 ) | ( n13813 & n20993 ) ;
  assign n20995 = n8398 & n20994 ;
  assign n20996 = n3843 & ~n6874 ;
  assign n20997 = n20996 ^ n9449 ^ 1'b0 ;
  assign n20998 = ~n3666 & n13834 ;
  assign n20999 = n20998 ^ n5181 ^ 1'b0 ;
  assign n21000 = ~n6986 & n10223 ;
  assign n21001 = n21000 ^ n5302 ^ n5144 ;
  assign n21002 = ( n6700 & n20999 ) | ( n6700 & ~n21001 ) | ( n20999 & ~n21001 ) ;
  assign n21003 = n8037 & n21002 ;
  assign n21004 = n17354 | n17548 ;
  assign n21005 = n10344 ^ n771 ^ 1'b0 ;
  assign n21006 = n3539 ^ n3079 ^ 1'b0 ;
  assign n21007 = ~n332 & n21006 ;
  assign n21008 = ~n14709 & n21007 ;
  assign n21009 = n21008 ^ n5374 ^ 1'b0 ;
  assign n21010 = ( n1481 & n1507 ) | ( n1481 & ~n4228 ) | ( n1507 & ~n4228 ) ;
  assign n21011 = n12539 & n18847 ;
  assign n21012 = n21011 ^ n7758 ^ n7064 ;
  assign n21013 = ( n20207 & ~n21010 ) | ( n20207 & n21012 ) | ( ~n21010 & n21012 ) ;
  assign n21014 = n17041 ^ n8273 ^ n6381 ;
  assign n21019 = n2663 & n2962 ;
  assign n21020 = n21019 ^ n7490 ^ n5248 ;
  assign n21021 = n1511 & n21020 ;
  assign n21022 = ~n14011 & n21021 ;
  assign n21023 = n21022 ^ n17213 ^ 1'b0 ;
  assign n21024 = n21023 ^ n15819 ^ n12927 ;
  assign n21015 = n8718 ^ n4580 ^ 1'b0 ;
  assign n21016 = n6041 & ~n21015 ;
  assign n21017 = n21016 ^ n8804 ^ 1'b0 ;
  assign n21018 = n14384 & n21017 ;
  assign n21025 = n21024 ^ n21018 ^ 1'b0 ;
  assign n21026 = ( n3656 & n16790 ) | ( n3656 & ~n17432 ) | ( n16790 & ~n17432 ) ;
  assign n21027 = n20848 ^ n16679 ^ 1'b0 ;
  assign n21028 = ~n21026 & n21027 ;
  assign n21029 = n14962 ^ n5024 ^ 1'b0 ;
  assign n21030 = n12424 & n21029 ;
  assign n21034 = n15133 ^ n6153 ^ 1'b0 ;
  assign n21035 = n9805 & ~n21034 ;
  assign n21031 = ( n8975 & n9587 ) | ( n8975 & n10635 ) | ( n9587 & n10635 ) ;
  assign n21032 = n17506 ^ n13281 ^ 1'b0 ;
  assign n21033 = n21031 & ~n21032 ;
  assign n21036 = n21035 ^ n21033 ^ n14697 ;
  assign n21037 = ( n2889 & n8781 ) | ( n2889 & ~n12865 ) | ( n8781 & ~n12865 ) ;
  assign n21038 = n21037 ^ n5349 ^ 1'b0 ;
  assign n21040 = n11632 ^ n5225 ^ n1475 ;
  assign n21039 = n1917 | n13642 ;
  assign n21041 = n21040 ^ n21039 ^ 1'b0 ;
  assign n21042 = ~n838 & n8209 ;
  assign n21043 = n21042 ^ n4665 ^ 1'b0 ;
  assign n21044 = n595 | n21043 ;
  assign n21045 = n599 & ~n15196 ;
  assign n21046 = ~n18099 & n21045 ;
  assign n21047 = n8172 ^ n6891 ^ n4601 ;
  assign n21048 = n21046 | n21047 ;
  assign n21049 = n3184 | n21048 ;
  assign n21050 = ( n1299 & n4547 ) | ( n1299 & ~n10330 ) | ( n4547 & ~n10330 ) ;
  assign n21051 = ~n9597 & n9716 ;
  assign n21052 = n21051 ^ n4973 ^ 1'b0 ;
  assign n21053 = n9938 & ~n21052 ;
  assign n21054 = ( n10635 & ~n18973 ) | ( n10635 & n21053 ) | ( ~n18973 & n21053 ) ;
  assign n21055 = ( n1977 & n1989 ) | ( n1977 & n17837 ) | ( n1989 & n17837 ) ;
  assign n21056 = ( n8475 & ~n13358 ) | ( n8475 & n19168 ) | ( ~n13358 & n19168 ) ;
  assign n21057 = n15354 ^ n12712 ^ n12408 ;
  assign n21058 = n21057 ^ n9631 ^ 1'b0 ;
  assign n21059 = n5427 & ~n15706 ;
  assign n21060 = n21059 ^ n7953 ^ 1'b0 ;
  assign n21061 = ( ~n15993 & n18249 ) | ( ~n15993 & n21060 ) | ( n18249 & n21060 ) ;
  assign n21062 = ( n11723 & n15338 ) | ( n11723 & ~n21061 ) | ( n15338 & ~n21061 ) ;
  assign n21063 = n21062 ^ n9487 ^ 1'b0 ;
  assign n21064 = ~n3571 & n21063 ;
  assign n21065 = n14805 ^ n3053 ^ n345 ;
  assign n21066 = ( n2411 & n9082 ) | ( n2411 & ~n21065 ) | ( n9082 & ~n21065 ) ;
  assign n21070 = n15661 ^ n10466 ^ 1'b0 ;
  assign n21071 = n5368 & ~n21070 ;
  assign n21067 = n18835 ^ n7544 ^ 1'b0 ;
  assign n21068 = n11557 & ~n21067 ;
  assign n21069 = ~n5786 & n21068 ;
  assign n21072 = n21071 ^ n21069 ^ n11973 ;
  assign n21074 = n15615 ^ n7173 ^ 1'b0 ;
  assign n21075 = n3416 | n21074 ;
  assign n21073 = n5234 & n8656 ;
  assign n21076 = n21075 ^ n21073 ^ n18316 ;
  assign n21078 = ( ~n3253 & n4048 ) | ( ~n3253 & n6746 ) | ( n4048 & n6746 ) ;
  assign n21077 = n5696 ^ n1113 ^ 1'b0 ;
  assign n21079 = n21078 ^ n21077 ^ n19902 ;
  assign n21080 = n13025 | n21079 ;
  assign n21081 = n21080 ^ n4820 ^ 1'b0 ;
  assign n21082 = n13822 ^ n8680 ^ 1'b0 ;
  assign n21083 = ( n4445 & n20989 ) | ( n4445 & ~n21082 ) | ( n20989 & ~n21082 ) ;
  assign n21084 = n13863 ^ n9115 ^ n8763 ;
  assign n21085 = n6989 & ~n7730 ;
  assign n21086 = n21085 ^ n3053 ^ 1'b0 ;
  assign n21087 = ( ~n6601 & n21084 ) | ( ~n6601 & n21086 ) | ( n21084 & n21086 ) ;
  assign n21088 = n7202 | n13224 ;
  assign n21089 = n21088 ^ n16301 ^ n136 ;
  assign n21090 = n7133 | n19722 ;
  assign n21091 = n950 & ~n21090 ;
  assign n21092 = n4090 ^ n2050 ^ 1'b0 ;
  assign n21093 = n12433 & ~n21092 ;
  assign n21094 = n8613 & n16387 ;
  assign n21095 = n6247 | n7674 ;
  assign n21096 = n21094 | n21095 ;
  assign n21097 = n21096 ^ n11468 ^ 1'b0 ;
  assign n21098 = n21097 ^ n10937 ^ 1'b0 ;
  assign n21099 = n21093 & ~n21098 ;
  assign n21100 = n2592 & n4353 ;
  assign n21101 = ~n21099 & n21100 ;
  assign n21102 = n18098 ^ n813 ^ 1'b0 ;
  assign n21103 = n4976 & ~n20810 ;
  assign n21104 = n21102 & ~n21103 ;
  assign n21105 = ( n8535 & ~n10021 ) | ( n8535 & n11395 ) | ( ~n10021 & n11395 ) ;
  assign n21106 = n21105 ^ n8802 ^ 1'b0 ;
  assign n21107 = n11628 ^ n6039 ^ n3288 ;
  assign n21108 = n21106 & n21107 ;
  assign n21109 = n3349 & n21108 ;
  assign n21110 = ~n21104 & n21109 ;
  assign n21111 = ( n14722 & n17495 ) | ( n14722 & ~n19687 ) | ( n17495 & ~n19687 ) ;
  assign n21112 = n20745 ^ n19362 ^ n9719 ;
  assign n21113 = n20982 ^ n7013 ^ 1'b0 ;
  assign n21114 = n12991 | n21113 ;
  assign n21115 = n8013 | n11616 ;
  assign n21116 = n10661 | n21115 ;
  assign n21117 = n3261 & ~n8882 ;
  assign n21118 = n12260 ^ n5644 ^ n4542 ;
  assign n21119 = n7662 | n18775 ;
  assign n21120 = n21119 ^ n4465 ^ 1'b0 ;
  assign n21121 = n21120 ^ n15587 ^ n2171 ;
  assign n21122 = n21121 ^ n17080 ^ n11064 ;
  assign n21123 = n5267 | n9777 ;
  assign n21124 = n21123 ^ n11315 ^ 1'b0 ;
  assign n21125 = ~n19227 & n21124 ;
  assign n21126 = n21125 ^ n245 ^ 1'b0 ;
  assign n21127 = ~n1533 & n13402 ;
  assign n21128 = n21127 ^ n2378 ^ n1628 ;
  assign n21129 = n243 | n21128 ;
  assign n21130 = n21129 ^ n1076 ^ 1'b0 ;
  assign n21131 = n11289 ^ n7366 ^ n1621 ;
  assign n21132 = ( n1970 & ~n13087 ) | ( n1970 & n21131 ) | ( ~n13087 & n21131 ) ;
  assign n21133 = n14897 ^ n6689 ^ 1'b0 ;
  assign n21134 = n6331 & ~n21133 ;
  assign n21135 = ( n6803 & ~n17514 ) | ( n6803 & n21134 ) | ( ~n17514 & n21134 ) ;
  assign n21136 = n20673 ^ n8988 ^ n7232 ;
  assign n21137 = n12184 | n15388 ;
  assign n21138 = ( n1330 & n3942 ) | ( n1330 & ~n8945 ) | ( n3942 & ~n8945 ) ;
  assign n21139 = n14169 ^ n2955 ^ 1'b0 ;
  assign n21140 = n3537 | n21139 ;
  assign n21141 = n185 & ~n21140 ;
  assign n21142 = ~x104 & n17035 ;
  assign n21143 = n21142 ^ n12546 ^ 1'b0 ;
  assign n21144 = n6379 ^ n3843 ^ 1'b0 ;
  assign n21145 = n21144 ^ n19424 ^ 1'b0 ;
  assign n21146 = n21143 & n21145 ;
  assign n21147 = ( n711 & n3483 ) | ( n711 & n7194 ) | ( n3483 & n7194 ) ;
  assign n21148 = n7994 & ~n11801 ;
  assign n21149 = ~n3545 & n21148 ;
  assign n21150 = n21147 & ~n21149 ;
  assign n21151 = n4469 & n21150 ;
  assign n21152 = n1183 | n4744 ;
  assign n21153 = n2634 & ~n21152 ;
  assign n21154 = n5934 ^ n3812 ^ 1'b0 ;
  assign n21156 = n8944 ^ n4274 ^ 1'b0 ;
  assign n21157 = ~n15894 & n21156 ;
  assign n21158 = n21157 ^ n9438 ^ 1'b0 ;
  assign n21155 = ( n3964 & n7097 ) | ( n3964 & n11818 ) | ( n7097 & n11818 ) ;
  assign n21159 = n21158 ^ n21155 ^ n12177 ;
  assign n21160 = n21159 ^ n17917 ^ n988 ;
  assign n21161 = n20021 ^ n5634 ^ n3566 ;
  assign n21162 = n1849 & ~n9881 ;
  assign n21163 = x66 & ~n18114 ;
  assign n21164 = n7473 & n21163 ;
  assign n21165 = n21164 ^ n17089 ^ 1'b0 ;
  assign n21166 = n2510 | n21165 ;
  assign n21167 = n6732 ^ n3311 ^ 1'b0 ;
  assign n21168 = n21167 ^ n13635 ^ 1'b0 ;
  assign n21169 = n1991 & ~n5318 ;
  assign n21170 = n21169 ^ n536 ^ 1'b0 ;
  assign n21171 = ~n8521 & n21170 ;
  assign n21172 = n21171 ^ n18455 ^ n14626 ;
  assign n21173 = ( n8139 & n8486 ) | ( n8139 & n14096 ) | ( n8486 & n14096 ) ;
  assign n21175 = n5496 ^ n4857 ^ 1'b0 ;
  assign n21176 = ~n14504 & n21175 ;
  assign n21174 = ~n2589 & n3603 ;
  assign n21177 = n21176 ^ n21174 ^ 1'b0 ;
  assign n21178 = n8904 & ~n15893 ;
  assign n21179 = n19178 & n21178 ;
  assign n21180 = x42 & n21179 ;
  assign n21181 = n1404 & ~n4177 ;
  assign n21182 = n21181 ^ n18195 ^ 1'b0 ;
  assign n21184 = n1709 ^ n1456 ^ 1'b0 ;
  assign n21183 = ( n5612 & n8157 ) | ( n5612 & ~n13780 ) | ( n8157 & ~n13780 ) ;
  assign n21185 = n21184 ^ n21183 ^ n4934 ;
  assign n21186 = n21185 ^ n12461 ^ n6730 ;
  assign n21187 = n13205 & ~n21186 ;
  assign n21188 = n21187 ^ n8927 ^ 1'b0 ;
  assign n21189 = n12331 ^ n10813 ^ 1'b0 ;
  assign n21190 = n2423 & n5956 ;
  assign n21191 = n21190 ^ n11613 ^ n9538 ;
  assign n21192 = ( ~n1583 & n3063 ) | ( ~n1583 & n14445 ) | ( n3063 & n14445 ) ;
  assign n21193 = n21192 ^ n12903 ^ n2678 ;
  assign n21194 = n2283 & ~n7603 ;
  assign n21195 = n21194 ^ n6627 ^ 1'b0 ;
  assign n21196 = n12350 ^ n2704 ^ n2038 ;
  assign n21197 = ( n3070 & n21195 ) | ( n3070 & ~n21196 ) | ( n21195 & ~n21196 ) ;
  assign n21198 = n529 | n6174 ;
  assign n21199 = ~n1808 & n12538 ;
  assign n21200 = n21198 & n21199 ;
  assign n21201 = n21200 ^ n7882 ^ 1'b0 ;
  assign n21202 = ~n7288 & n15458 ;
  assign n21203 = ~n21201 & n21202 ;
  assign n21204 = n16835 ^ n4224 ^ 1'b0 ;
  assign n21205 = ~n15876 & n21204 ;
  assign n21206 = ~n2847 & n21205 ;
  assign n21207 = n12225 ^ n11468 ^ n7839 ;
  assign n21208 = n21207 ^ n10268 ^ n7130 ;
  assign n21209 = n21208 ^ n14900 ^ n854 ;
  assign n21213 = ( n1318 & n7546 ) | ( n1318 & n12132 ) | ( n7546 & n12132 ) ;
  assign n21210 = n15664 ^ n11995 ^ n802 ;
  assign n21211 = ~n13963 & n21210 ;
  assign n21212 = ~n7812 & n21211 ;
  assign n21214 = n21213 ^ n21212 ^ n11622 ;
  assign n21215 = n2747 ^ n2242 ^ n896 ;
  assign n21216 = n21215 ^ n9877 ^ n2371 ;
  assign n21217 = n5041 & n6083 ;
  assign n21218 = n21217 ^ n14139 ^ 1'b0 ;
  assign n21219 = ( n2319 & n2980 ) | ( n2319 & ~n12043 ) | ( n2980 & ~n12043 ) ;
  assign n21221 = n9943 ^ n7342 ^ 1'b0 ;
  assign n21220 = n2348 & n11337 ;
  assign n21222 = n21221 ^ n21220 ^ n12035 ;
  assign n21223 = ~n21219 & n21222 ;
  assign n21224 = n21223 ^ n11873 ^ 1'b0 ;
  assign n21232 = n4143 ^ n3264 ^ n1862 ;
  assign n21225 = ~n1732 & n12578 ;
  assign n21226 = n21225 ^ n6749 ^ 1'b0 ;
  assign n21227 = n21226 ^ n11636 ^ 1'b0 ;
  assign n21228 = n9016 ^ n5071 ^ n518 ;
  assign n21229 = ~n12845 & n21228 ;
  assign n21230 = n21229 ^ n454 ^ 1'b0 ;
  assign n21231 = ( n11889 & ~n21227 ) | ( n11889 & n21230 ) | ( ~n21227 & n21230 ) ;
  assign n21233 = n21232 ^ n21231 ^ 1'b0 ;
  assign n21234 = ~n21224 & n21233 ;
  assign n21235 = ( ~n1800 & n4679 ) | ( ~n1800 & n8778 ) | ( n4679 & n8778 ) ;
  assign n21236 = n4568 ^ n4265 ^ 1'b0 ;
  assign n21237 = n724 | n11892 ;
  assign n21238 = n10316 & n15327 ;
  assign n21239 = ( n4420 & n9953 ) | ( n4420 & n10606 ) | ( n9953 & n10606 ) ;
  assign n21240 = n21239 ^ n806 ^ 1'b0 ;
  assign n21241 = n9273 & n10608 ;
  assign n21242 = n8322 & n21241 ;
  assign n21243 = n1311 & n1762 ;
  assign n21244 = ~n3891 & n21243 ;
  assign n21247 = n16205 ^ n12042 ^ 1'b0 ;
  assign n21245 = n19566 | n20175 ;
  assign n21246 = n21245 ^ n199 ^ 1'b0 ;
  assign n21248 = n21247 ^ n21246 ^ n967 ;
  assign n21249 = n10581 ^ n6773 ^ n130 ;
  assign n21250 = ( n4722 & n6621 ) | ( n4722 & n12981 ) | ( n6621 & n12981 ) ;
  assign n21251 = ( n16936 & ~n21249 ) | ( n16936 & n21250 ) | ( ~n21249 & n21250 ) ;
  assign n21252 = n18454 ^ n14385 ^ n12075 ;
  assign n21254 = n13141 ^ n9363 ^ 1'b0 ;
  assign n21255 = n13811 & n21254 ;
  assign n21253 = n2252 & ~n9386 ;
  assign n21256 = n21255 ^ n21253 ^ 1'b0 ;
  assign n21257 = ~n3610 & n7056 ;
  assign n21261 = n780 & n7134 ;
  assign n21262 = n21261 ^ n4977 ^ 1'b0 ;
  assign n21258 = n9934 ^ n1134 ^ 1'b0 ;
  assign n21259 = n2075 & ~n11124 ;
  assign n21260 = n21258 & n21259 ;
  assign n21263 = n21262 ^ n21260 ^ n12214 ;
  assign n21264 = n17192 ^ n2488 ^ 1'b0 ;
  assign n21265 = n3648 ^ x59 ^ 1'b0 ;
  assign n21268 = n8219 ^ n8091 ^ n5680 ;
  assign n21269 = n12870 | n21268 ;
  assign n21270 = n21269 ^ x33 ^ 1'b0 ;
  assign n21266 = n9418 & n14559 ;
  assign n21267 = n21266 ^ n7530 ^ 1'b0 ;
  assign n21271 = n21270 ^ n21267 ^ n14720 ;
  assign n21273 = n6267 ^ n3141 ^ 1'b0 ;
  assign n21272 = n10438 ^ n7125 ^ n6984 ;
  assign n21274 = n21273 ^ n21272 ^ n624 ;
  assign n21275 = n21274 ^ n18841 ^ n17326 ;
  assign n21276 = n21275 ^ n4643 ^ 1'b0 ;
  assign n21277 = n17902 & ~n21276 ;
  assign n21278 = n19995 ^ n10361 ^ n10080 ;
  assign n21279 = ~n10979 & n21278 ;
  assign n21280 = n8580 ^ n4642 ^ n3459 ;
  assign n21281 = n11783 ^ n10157 ^ n4434 ;
  assign n21282 = n18402 ^ n16009 ^ n3406 ;
  assign n21283 = n9720 ^ n5766 ^ 1'b0 ;
  assign n21284 = n9497 & ~n21283 ;
  assign n21290 = n8505 ^ n3904 ^ n2906 ;
  assign n21291 = n21290 ^ n17741 ^ n3902 ;
  assign n21288 = n368 & n6325 ;
  assign n21289 = n21288 ^ n7526 ^ 1'b0 ;
  assign n21292 = n21291 ^ n21289 ^ n9276 ;
  assign n21285 = ( n3795 & ~n3914 ) | ( n3795 & n4675 ) | ( ~n3914 & n4675 ) ;
  assign n21286 = n9380 & n21285 ;
  assign n21287 = ~n16434 & n21286 ;
  assign n21293 = n21292 ^ n21287 ^ n4452 ;
  assign n21294 = ( n11840 & n12664 ) | ( n11840 & n13919 ) | ( n12664 & n13919 ) ;
  assign n21295 = n21294 ^ n18481 ^ n4500 ;
  assign n21296 = ~n9876 & n10977 ;
  assign n21297 = n7017 ^ n2389 ^ n2276 ;
  assign n21298 = ~n7793 & n21297 ;
  assign n21299 = ~n4250 & n21298 ;
  assign n21300 = n6382 ^ n4322 ^ n3990 ;
  assign n21301 = ( ~n6307 & n12120 ) | ( ~n6307 & n21300 ) | ( n12120 & n21300 ) ;
  assign n21302 = ( n15057 & n21299 ) | ( n15057 & n21301 ) | ( n21299 & n21301 ) ;
  assign n21303 = n13068 ^ n5135 ^ 1'b0 ;
  assign n21304 = ~n16199 & n21303 ;
  assign n21305 = ( n2077 & ~n14221 ) | ( n2077 & n21304 ) | ( ~n14221 & n21304 ) ;
  assign n21306 = n21305 ^ n6073 ^ 1'b0 ;
  assign n21307 = n21306 ^ n11633 ^ n1477 ;
  assign n21308 = n10822 & ~n14353 ;
  assign n21309 = ~n17731 & n21308 ;
  assign n21310 = n21309 ^ n7715 ^ 1'b0 ;
  assign n21311 = n16181 ^ n8556 ^ n3679 ;
  assign n21312 = ( n332 & n10407 ) | ( n332 & ~n21311 ) | ( n10407 & ~n21311 ) ;
  assign n21313 = ( n7448 & n13645 ) | ( n7448 & n21312 ) | ( n13645 & n21312 ) ;
  assign n21314 = n6142 & ~n9619 ;
  assign n21315 = n21313 & n21314 ;
  assign n21316 = n2259 & n11363 ;
  assign n21317 = n21316 ^ n2103 ^ 1'b0 ;
  assign n21318 = ~n8453 & n20001 ;
  assign n21319 = ( ~n9285 & n13867 ) | ( ~n9285 & n19480 ) | ( n13867 & n19480 ) ;
  assign n21320 = n7993 & ~n16777 ;
  assign n21321 = n17804 ^ n3560 ^ 1'b0 ;
  assign n21322 = ( x19 & ~n19157 ) | ( x19 & n21321 ) | ( ~n19157 & n21321 ) ;
  assign n21323 = ~n1445 & n8973 ;
  assign n21324 = n19788 ^ n14298 ^ n2097 ;
  assign n21325 = n21324 ^ n19971 ^ n2541 ;
  assign n21326 = n10203 ^ n7262 ^ n4524 ;
  assign n21327 = ( ~n10141 & n11523 ) | ( ~n10141 & n19828 ) | ( n11523 & n19828 ) ;
  assign n21331 = n10058 ^ n1965 ^ n1298 ;
  assign n21332 = ( n8616 & ~n20109 ) | ( n8616 & n21331 ) | ( ~n20109 & n21331 ) ;
  assign n21328 = n3067 | n6460 ;
  assign n21329 = n21328 ^ n2284 ^ 1'b0 ;
  assign n21330 = n21329 ^ n10861 ^ n591 ;
  assign n21333 = n21332 ^ n21330 ^ n11660 ;
  assign n21334 = n18674 ^ n12961 ^ n8805 ;
  assign n21335 = n11131 ^ n3927 ^ 1'b0 ;
  assign n21336 = n21334 & n21335 ;
  assign n21337 = ( ~n2325 & n5016 ) | ( ~n2325 & n11468 ) | ( n5016 & n11468 ) ;
  assign n21338 = ( n2046 & n6255 ) | ( n2046 & n21337 ) | ( n6255 & n21337 ) ;
  assign n21339 = ( ~n1997 & n2607 ) | ( ~n1997 & n6102 ) | ( n2607 & n6102 ) ;
  assign n21340 = n5296 & n21339 ;
  assign n21341 = n6116 & n21340 ;
  assign n21342 = n511 | n6210 ;
  assign n21343 = n209 & ~n21342 ;
  assign n21344 = n21343 ^ n8809 ^ 1'b0 ;
  assign n21345 = ( ~n3609 & n21341 ) | ( ~n3609 & n21344 ) | ( n21341 & n21344 ) ;
  assign n21348 = n7793 | n9096 ;
  assign n21349 = n788 & ~n21348 ;
  assign n21346 = ~n2193 & n18977 ;
  assign n21347 = n21346 ^ n9628 ^ 1'b0 ;
  assign n21350 = n21349 ^ n21347 ^ n12856 ;
  assign n21352 = n1147 | n6221 ;
  assign n21351 = ( n1919 & ~n3652 ) | ( n1919 & n6376 ) | ( ~n3652 & n6376 ) ;
  assign n21353 = n21352 ^ n21351 ^ n11053 ;
  assign n21354 = n15890 & ~n21305 ;
  assign n21355 = n17876 & n21354 ;
  assign n21356 = n11091 ^ n2512 ^ n1170 ;
  assign n21357 = n9800 & n21356 ;
  assign n21358 = n4536 & n21357 ;
  assign n21359 = ~n2419 & n6326 ;
  assign n21360 = n5473 & n21359 ;
  assign n21361 = n3466 & n9440 ;
  assign n21362 = n21360 & n21361 ;
  assign n21363 = n6873 | n8465 ;
  assign n21364 = n5979 & ~n21363 ;
  assign n21365 = ( n1761 & ~n8967 ) | ( n1761 & n21364 ) | ( ~n8967 & n21364 ) ;
  assign n21366 = n7004 ^ n2343 ^ 1'b0 ;
  assign n21367 = ~n5923 & n21366 ;
  assign n21368 = ( n16703 & ~n19461 ) | ( n16703 & n21367 ) | ( ~n19461 & n21367 ) ;
  assign n21369 = n21368 ^ n2261 ^ 1'b0 ;
  assign n21370 = ~n21365 & n21369 ;
  assign n21371 = ( ~n5764 & n6924 ) | ( ~n5764 & n14358 ) | ( n6924 & n14358 ) ;
  assign n21372 = n21371 ^ n11248 ^ n7735 ;
  assign n21373 = n17929 ^ n557 ^ 1'b0 ;
  assign n21374 = n21372 | n21373 ;
  assign n21375 = n12892 ^ n5853 ^ 1'b0 ;
  assign n21377 = n13366 ^ n9391 ^ 1'b0 ;
  assign n21378 = n3773 & ~n21377 ;
  assign n21376 = ( ~n7695 & n9630 ) | ( ~n7695 & n10679 ) | ( n9630 & n10679 ) ;
  assign n21379 = n21378 ^ n21376 ^ n1210 ;
  assign n21380 = ~n570 & n21379 ;
  assign n21381 = n18741 ^ n1486 ^ n1273 ;
  assign n21383 = n5369 & ~n20877 ;
  assign n21384 = ~n16316 & n21383 ;
  assign n21385 = n8781 & n21384 ;
  assign n21382 = n7388 ^ n1303 ^ n1055 ;
  assign n21386 = n21385 ^ n21382 ^ n2481 ;
  assign n21388 = ( n3140 & ~n3175 ) | ( n3140 & n10143 ) | ( ~n3175 & n10143 ) ;
  assign n21389 = n12765 | n21388 ;
  assign n21390 = n21389 ^ n11137 ^ 1'b0 ;
  assign n21387 = n12745 | n20759 ;
  assign n21391 = n21390 ^ n21387 ^ n12644 ;
  assign n21392 = n13508 ^ n8537 ^ n1422 ;
  assign n21393 = n14948 ^ n8729 ^ n6677 ;
  assign n21394 = n9612 ^ n9304 ^ n8167 ;
  assign n21395 = ( ~n21392 & n21393 ) | ( ~n21392 & n21394 ) | ( n21393 & n21394 ) ;
  assign n21396 = n21395 ^ n20339 ^ n6863 ;
  assign n21397 = n12960 ^ n6738 ^ 1'b0 ;
  assign n21398 = n1622 | n21397 ;
  assign n21399 = n21398 ^ n10936 ^ 1'b0 ;
  assign n21400 = ( n1361 & n14885 ) | ( n1361 & n21399 ) | ( n14885 & n21399 ) ;
  assign n21401 = n21400 ^ n13061 ^ 1'b0 ;
  assign n21402 = ( n705 & n5597 ) | ( n705 & ~n18725 ) | ( n5597 & ~n18725 ) ;
  assign n21403 = ( n706 & n14796 ) | ( n706 & ~n19242 ) | ( n14796 & ~n19242 ) ;
  assign n21404 = n21403 ^ n8640 ^ 1'b0 ;
  assign n21405 = n1870 & ~n4516 ;
  assign n21406 = n5307 & n21405 ;
  assign n21407 = n1205 | n4974 ;
  assign n21408 = n21406 & ~n21407 ;
  assign n21410 = ( n3294 & n3543 ) | ( n3294 & ~n8247 ) | ( n3543 & ~n8247 ) ;
  assign n21409 = n4913 & ~n19844 ;
  assign n21411 = n21410 ^ n21409 ^ 1'b0 ;
  assign n21412 = n5197 | n21411 ;
  assign n21413 = n21412 ^ n515 ^ 1'b0 ;
  assign n21414 = n20366 ^ n8281 ^ n7490 ;
  assign n21415 = n21414 ^ n7599 ^ 1'b0 ;
  assign n21416 = n6548 & n18369 ;
  assign n21417 = n21416 ^ n16143 ^ 1'b0 ;
  assign n21418 = n8473 ^ n4780 ^ 1'b0 ;
  assign n21419 = n21418 ^ n13986 ^ n3809 ;
  assign n21420 = ( ~n5927 & n21417 ) | ( ~n5927 & n21419 ) | ( n21417 & n21419 ) ;
  assign n21421 = n9404 ^ n4293 ^ 1'b0 ;
  assign n21422 = ~n3567 & n21421 ;
  assign n21423 = ~n11363 & n21422 ;
  assign n21424 = n19950 ^ n13313 ^ 1'b0 ;
  assign n21425 = ( n7661 & n7842 ) | ( n7661 & n21424 ) | ( n7842 & n21424 ) ;
  assign n21426 = ( n7147 & n9779 ) | ( n7147 & n13011 ) | ( n9779 & n13011 ) ;
  assign n21427 = ~n7205 & n13327 ;
  assign n21428 = ~n17202 & n21427 ;
  assign n21429 = n14819 ^ n4581 ^ 1'b0 ;
  assign n21430 = n4568 ^ n3631 ^ 1'b0 ;
  assign n21431 = n21430 ^ n14674 ^ n7630 ;
  assign n21432 = n197 & ~n1437 ;
  assign n21433 = ~n10915 & n18127 ;
  assign n21434 = n15774 ^ n10413 ^ n957 ;
  assign n21435 = ( n7320 & ~n15735 ) | ( n7320 & n21434 ) | ( ~n15735 & n21434 ) ;
  assign n21436 = n7141 ^ n2820 ^ n523 ;
  assign n21437 = n21436 ^ n10057 ^ 1'b0 ;
  assign n21438 = n21435 & n21437 ;
  assign n21439 = ~n8675 & n12523 ;
  assign n21440 = ~n16079 & n21439 ;
  assign n21441 = n13900 ^ n11119 ^ 1'b0 ;
  assign n21442 = n1860 | n8569 ;
  assign n21443 = n21442 ^ n2018 ^ 1'b0 ;
  assign n21444 = n21443 ^ n4106 ^ n1668 ;
  assign n21445 = n6698 & ~n21444 ;
  assign n21446 = ~n1796 & n21445 ;
  assign n21447 = n664 | n21446 ;
  assign n21448 = n21441 & ~n21447 ;
  assign n21449 = n21351 ^ n7302 ^ 1'b0 ;
  assign n21450 = ~n11265 & n15256 ;
  assign n21451 = ( n1600 & n12183 ) | ( n1600 & ~n21450 ) | ( n12183 & ~n21450 ) ;
  assign n21452 = n21451 ^ n7729 ^ 1'b0 ;
  assign n21453 = n406 & n717 ;
  assign n21454 = n21453 ^ n21337 ^ 1'b0 ;
  assign n21455 = n21454 ^ n20520 ^ n472 ;
  assign n21456 = n15003 ^ n1589 ^ 1'b0 ;
  assign n21457 = n2832 ^ n1900 ^ n562 ;
  assign n21458 = n21457 ^ n15897 ^ 1'b0 ;
  assign n21459 = n6042 & n21458 ;
  assign n21465 = n9115 & ~n14290 ;
  assign n21466 = n21465 ^ n8875 ^ n2700 ;
  assign n21462 = n2288 ^ n1600 ^ n203 ;
  assign n21463 = ~n3661 & n21462 ;
  assign n21464 = n11394 & n21463 ;
  assign n21460 = ( n9294 & ~n14419 ) | ( n9294 & n15173 ) | ( ~n14419 & n15173 ) ;
  assign n21461 = n21460 ^ n13936 ^ 1'b0 ;
  assign n21467 = n21466 ^ n21464 ^ n21461 ;
  assign n21468 = n13809 ^ n4591 ^ 1'b0 ;
  assign n21469 = n21468 ^ n9144 ^ 1'b0 ;
  assign n21470 = ( ~n9751 & n17767 ) | ( ~n9751 & n19512 ) | ( n17767 & n19512 ) ;
  assign n21471 = ~n4538 & n9757 ;
  assign n21472 = n14837 & n21471 ;
  assign n21473 = ~n15985 & n21472 ;
  assign n21474 = ( n178 & n12411 ) | ( n178 & n18637 ) | ( n12411 & n18637 ) ;
  assign n21475 = n14185 | n21474 ;
  assign n21476 = n1019 & ~n21475 ;
  assign n21477 = ( ~n2470 & n9219 ) | ( ~n2470 & n12541 ) | ( n9219 & n12541 ) ;
  assign n21478 = ( ~n2116 & n4438 ) | ( ~n2116 & n21477 ) | ( n4438 & n21477 ) ;
  assign n21479 = ( n11337 & ~n15244 ) | ( n11337 & n18756 ) | ( ~n15244 & n18756 ) ;
  assign n21480 = n20931 ^ n13801 ^ n11842 ;
  assign n21481 = n17040 & ~n17758 ;
  assign n21482 = n18222 & ~n21481 ;
  assign n21483 = n1176 & ~n1338 ;
  assign n21484 = n2928 ^ n2661 ^ x115 ;
  assign n21485 = n6983 & ~n16733 ;
  assign n21486 = ( n2493 & n21484 ) | ( n2493 & ~n21485 ) | ( n21484 & ~n21485 ) ;
  assign n21487 = ( ~n2091 & n5535 ) | ( ~n2091 & n9790 ) | ( n5535 & n9790 ) ;
  assign n21488 = n21487 ^ n20551 ^ n8962 ;
  assign n21489 = n18586 ^ n9646 ^ n2187 ;
  assign n21490 = n18228 | n21489 ;
  assign n21491 = n5934 & n16849 ;
  assign n21492 = n10743 ^ n8393 ^ x67 ;
  assign n21493 = n21492 ^ n12718 ^ n8546 ;
  assign n21494 = ( n1006 & ~n12186 ) | ( n1006 & n21493 ) | ( ~n12186 & n21493 ) ;
  assign n21495 = ( ~n6445 & n7528 ) | ( ~n6445 & n10457 ) | ( n7528 & n10457 ) ;
  assign n21496 = n10759 | n15157 ;
  assign n21497 = n12735 | n21496 ;
  assign n21498 = n6272 | n21497 ;
  assign n21499 = ~n520 & n21498 ;
  assign n21500 = n21495 & n21499 ;
  assign n21501 = ( n129 & n5403 ) | ( n129 & ~n21500 ) | ( n5403 & ~n21500 ) ;
  assign n21502 = n1752 & ~n6973 ;
  assign n21503 = ( n887 & n16911 ) | ( n887 & ~n21502 ) | ( n16911 & ~n21502 ) ;
  assign n21504 = ( n1073 & n16193 ) | ( n1073 & ~n21503 ) | ( n16193 & ~n21503 ) ;
  assign n21505 = n21504 ^ n12359 ^ 1'b0 ;
  assign n21506 = ~n2950 & n11491 ;
  assign n21507 = n21506 ^ n18280 ^ n4846 ;
  assign n21508 = n21507 ^ n15130 ^ n1899 ;
  assign n21509 = n11954 | n12351 ;
  assign n21510 = n21509 ^ n14293 ^ 1'b0 ;
  assign n21511 = n11819 | n20642 ;
  assign n21512 = n21510 & ~n21511 ;
  assign n21513 = n5716 & ~n6730 ;
  assign n21514 = n21513 ^ n20106 ^ 1'b0 ;
  assign n21515 = n21514 ^ n3330 ^ 1'b0 ;
  assign n21516 = n6513 | n21515 ;
  assign n21517 = ~n4237 & n6973 ;
  assign n21518 = n1685 & n12358 ;
  assign n21519 = ~n3091 & n21518 ;
  assign n21520 = n21519 ^ n2884 ^ n2335 ;
  assign n21521 = n13366 & ~n19071 ;
  assign n21522 = n21521 ^ n2694 ^ 1'b0 ;
  assign n21523 = n21522 ^ n16938 ^ n1152 ;
  assign n21524 = ~n13873 & n21232 ;
  assign n21525 = n7627 ^ n3243 ^ n2332 ;
  assign n21526 = n21525 ^ n1361 ^ n1283 ;
  assign n21527 = ( n2887 & n7156 ) | ( n2887 & ~n21526 ) | ( n7156 & ~n21526 ) ;
  assign n21528 = n9335 ^ n6968 ^ n6274 ;
  assign n21529 = n17596 ^ n6905 ^ x25 ;
  assign n21530 = n1660 & ~n21529 ;
  assign n21531 = n2733 & ~n17292 ;
  assign n21532 = n21531 ^ n17497 ^ 1'b0 ;
  assign n21533 = n21532 ^ n157 ^ 1'b0 ;
  assign n21534 = ~n17524 & n21533 ;
  assign n21535 = n21534 ^ n20509 ^ n3062 ;
  assign n21536 = n11782 ^ n7119 ^ 1'b0 ;
  assign n21537 = n21536 ^ n5098 ^ 1'b0 ;
  assign n21538 = n18043 | n21537 ;
  assign n21539 = n2043 & ~n16073 ;
  assign n21540 = n9582 & ~n12285 ;
  assign n21541 = n21540 ^ n10015 ^ 1'b0 ;
  assign n21542 = n5612 & ~n10845 ;
  assign n21543 = n15716 & n21542 ;
  assign n21544 = n13657 ^ n8146 ^ 1'b0 ;
  assign n21545 = x29 & ~n21544 ;
  assign n21546 = ( ~n19038 & n21543 ) | ( ~n19038 & n21545 ) | ( n21543 & n21545 ) ;
  assign n21547 = n17791 ^ n2978 ^ n1152 ;
  assign n21548 = ~n10778 & n18518 ;
  assign n21549 = n16169 ^ n13488 ^ n10256 ;
  assign n21550 = n6584 & n21549 ;
  assign n21551 = n21550 ^ n3089 ^ 1'b0 ;
  assign n21552 = ~n2928 & n3577 ;
  assign n21553 = ~n9102 & n21552 ;
  assign n21554 = n9287 ^ n794 ^ 1'b0 ;
  assign n21555 = n7493 ^ n7266 ^ n3585 ;
  assign n21556 = n16122 ^ n16009 ^ n10439 ;
  assign n21561 = ( ~n11033 & n12700 ) | ( ~n11033 & n16115 ) | ( n12700 & n16115 ) ;
  assign n21557 = n2407 ^ x123 ^ 1'b0 ;
  assign n21558 = n21557 ^ n9221 ^ n8670 ;
  assign n21559 = ~n2619 & n21558 ;
  assign n21560 = n21559 ^ n9553 ^ 1'b0 ;
  assign n21562 = n21561 ^ n21560 ^ n3020 ;
  assign n21563 = n14441 ^ n12923 ^ n1891 ;
  assign n21564 = ( n5182 & n8288 ) | ( n5182 & ~n21563 ) | ( n8288 & ~n21563 ) ;
  assign n21565 = n6862 ^ n412 ^ 1'b0 ;
  assign n21566 = n15381 ^ n5079 ^ 1'b0 ;
  assign n21567 = ~n957 & n21566 ;
  assign n21568 = ~n5100 & n21567 ;
  assign n21569 = ( n5550 & ~n21565 ) | ( n5550 & n21568 ) | ( ~n21565 & n21568 ) ;
  assign n21570 = n684 & n17075 ;
  assign n21571 = n21570 ^ n10917 ^ 1'b0 ;
  assign n21572 = n1290 | n2998 ;
  assign n21573 = ~n5671 & n5807 ;
  assign n21574 = ( n1011 & n12529 ) | ( n1011 & n21573 ) | ( n12529 & n21573 ) ;
  assign n21575 = n21574 ^ n14711 ^ n9806 ;
  assign n21576 = ( n15367 & ~n21572 ) | ( n15367 & n21575 ) | ( ~n21572 & n21575 ) ;
  assign n21577 = n2521 & ~n3915 ;
  assign n21578 = n19771 ^ n12126 ^ n3488 ;
  assign n21579 = ( ~n21406 & n21577 ) | ( ~n21406 & n21578 ) | ( n21577 & n21578 ) ;
  assign n21580 = ( ~n2315 & n3447 ) | ( ~n2315 & n21579 ) | ( n3447 & n21579 ) ;
  assign n21581 = ~n7618 & n21580 ;
  assign n21582 = n21581 ^ n1356 ^ 1'b0 ;
  assign n21583 = n3338 & ~n11020 ;
  assign n21584 = ( n5236 & n10959 ) | ( n5236 & ~n12839 ) | ( n10959 & ~n12839 ) ;
  assign n21585 = ( n2178 & n12116 ) | ( n2178 & n21584 ) | ( n12116 & n21584 ) ;
  assign n21586 = n10301 ^ n3078 ^ 1'b0 ;
  assign n21587 = n17599 ^ n13265 ^ 1'b0 ;
  assign n21588 = n4034 & ~n21587 ;
  assign n21589 = n13121 & ~n15819 ;
  assign n21590 = n20759 ^ n20090 ^ n2290 ;
  assign n21591 = n18098 ^ n15667 ^ n3695 ;
  assign n21592 = n21591 ^ n14807 ^ 1'b0 ;
  assign n21593 = n14014 & n21592 ;
  assign n21594 = n21593 ^ n16152 ^ n5283 ;
  assign n21595 = ( n442 & n10339 ) | ( n442 & ~n17411 ) | ( n10339 & ~n17411 ) ;
  assign n21596 = n1989 & n21595 ;
  assign n21597 = n21596 ^ n7654 ^ 1'b0 ;
  assign n21598 = n4405 & ~n21597 ;
  assign n21599 = ~n4489 & n14725 ;
  assign n21600 = n10300 & n21599 ;
  assign n21601 = n9540 & n21600 ;
  assign n21602 = n10747 ^ n2663 ^ 1'b0 ;
  assign n21603 = n7954 & n10501 ;
  assign n21604 = n21603 ^ n21304 ^ 1'b0 ;
  assign n21605 = ~n2577 & n15301 ;
  assign n21606 = n10719 & ~n17163 ;
  assign n21607 = ~n3727 & n21606 ;
  assign n21612 = n3652 ^ n2072 ^ 1'b0 ;
  assign n21609 = n3136 & ~n3201 ;
  assign n21610 = n21609 ^ n14148 ^ 1'b0 ;
  assign n21608 = n10991 | n12828 ;
  assign n21611 = n21610 ^ n21608 ^ 1'b0 ;
  assign n21613 = n21612 ^ n21611 ^ 1'b0 ;
  assign n21614 = n19221 ^ n795 ^ 1'b0 ;
  assign n21615 = n14353 ^ n7299 ^ n4052 ;
  assign n21616 = ( ~n3255 & n10533 ) | ( ~n3255 & n21615 ) | ( n10533 & n21615 ) ;
  assign n21617 = n19876 & ~n21616 ;
  assign n21618 = n12433 ^ n7468 ^ n1125 ;
  assign n21619 = n11829 ^ n8135 ^ n6191 ;
  assign n21620 = n8503 & n10078 ;
  assign n21621 = ( ~n12337 & n13382 ) | ( ~n12337 & n21620 ) | ( n13382 & n21620 ) ;
  assign n21622 = n6965 & ~n21621 ;
  assign n21623 = n7169 & n21622 ;
  assign n21624 = n4089 | n14701 ;
  assign n21625 = n21624 ^ n11523 ^ 1'b0 ;
  assign n21626 = n12669 ^ n6244 ^ 1'b0 ;
  assign n21627 = n21626 ^ n6177 ^ 1'b0 ;
  assign n21628 = ( n1664 & n3573 ) | ( n1664 & n4717 ) | ( n3573 & n4717 ) ;
  assign n21629 = n18289 ^ n9123 ^ n6218 ;
  assign n21630 = ( ~n907 & n1295 ) | ( ~n907 & n11200 ) | ( n1295 & n11200 ) ;
  assign n21631 = ( n1044 & ~n7486 ) | ( n1044 & n21630 ) | ( ~n7486 & n21630 ) ;
  assign n21632 = ( x59 & ~n1128 ) | ( x59 & n10840 ) | ( ~n1128 & n10840 ) ;
  assign n21633 = n768 & ~n21406 ;
  assign n21634 = ~n950 & n21633 ;
  assign n21635 = ( n5907 & n19144 ) | ( n5907 & n21634 ) | ( n19144 & n21634 ) ;
  assign n21636 = ( n4821 & ~n9230 ) | ( n4821 & n9348 ) | ( ~n9230 & n9348 ) ;
  assign n21637 = ( x117 & ~n3944 ) | ( x117 & n10063 ) | ( ~n3944 & n10063 ) ;
  assign n21638 = n21637 ^ n4805 ^ 1'b0 ;
  assign n21639 = ~n21636 & n21638 ;
  assign n21640 = n21639 ^ n19255 ^ 1'b0 ;
  assign n21641 = n8629 & ~n21640 ;
  assign n21642 = n4254 & n14180 ;
  assign n21643 = n21642 ^ n9509 ^ 1'b0 ;
  assign n21644 = n893 & ~n21643 ;
  assign n21645 = n18226 ^ n4842 ^ 1'b0 ;
  assign n21646 = n17307 ^ n11133 ^ 1'b0 ;
  assign n21647 = n1679 & ~n21646 ;
  assign n21648 = ( n3334 & n6671 ) | ( n3334 & n10568 ) | ( n6671 & n10568 ) ;
  assign n21649 = ( ~n12768 & n21647 ) | ( ~n12768 & n21648 ) | ( n21647 & n21648 ) ;
  assign n21650 = n20744 ^ n18639 ^ 1'b0 ;
  assign n21651 = n6104 ^ n4989 ^ n3390 ;
  assign n21652 = n15257 & ~n21651 ;
  assign n21653 = n14965 ^ n13650 ^ 1'b0 ;
  assign n21654 = n15988 | n19288 ;
  assign n21655 = n21653 & ~n21654 ;
  assign n21656 = ( n7643 & ~n14304 ) | ( n7643 & n21085 ) | ( ~n14304 & n21085 ) ;
  assign n21657 = n13601 | n17583 ;
  assign n21658 = n18973 ^ n18361 ^ 1'b0 ;
  assign n21659 = n6177 & ~n21658 ;
  assign n21660 = ( n15895 & n20057 ) | ( n15895 & ~n21418 ) | ( n20057 & ~n21418 ) ;
  assign n21662 = ( ~n2251 & n4553 ) | ( ~n2251 & n12400 ) | ( n4553 & n12400 ) ;
  assign n21661 = n10092 ^ n6442 ^ n4142 ;
  assign n21663 = n21662 ^ n21661 ^ n3901 ;
  assign n21664 = n416 & ~n21663 ;
  assign n21665 = n21660 & n21664 ;
  assign n21666 = ~n2718 & n18335 ;
  assign n21667 = n21666 ^ n20864 ^ 1'b0 ;
  assign n21668 = ~n11289 & n21667 ;
  assign n21669 = n13551 & ~n20296 ;
  assign n21670 = n3758 ^ n3398 ^ 1'b0 ;
  assign n21671 = n11316 ^ n9617 ^ n9553 ;
  assign n21672 = n13468 & ~n21671 ;
  assign n21673 = n19457 ^ n10876 ^ n2622 ;
  assign n21674 = n21673 ^ n8505 ^ n2905 ;
  assign n21675 = ( n5165 & n15522 ) | ( n5165 & ~n16546 ) | ( n15522 & ~n16546 ) ;
  assign n21676 = n19558 ^ n10283 ^ n9369 ;
  assign n21677 = n21676 ^ n20895 ^ n6716 ;
  assign n21678 = ( ~n16570 & n21675 ) | ( ~n16570 & n21677 ) | ( n21675 & n21677 ) ;
  assign n21679 = n18185 ^ n15938 ^ n3209 ;
  assign n21680 = n7064 ^ n3869 ^ n2178 ;
  assign n21681 = ~n7758 & n14370 ;
  assign n21682 = ( ~n3522 & n11846 ) | ( ~n3522 & n18322 ) | ( n11846 & n18322 ) ;
  assign n21683 = n10880 ^ n4786 ^ n3515 ;
  assign n21684 = ~n8362 & n9093 ;
  assign n21685 = n13567 ^ n12000 ^ 1'b0 ;
  assign n21687 = n15639 ^ n8759 ^ n950 ;
  assign n21686 = n8488 ^ n7114 ^ n4452 ;
  assign n21688 = n21687 ^ n21686 ^ n14957 ;
  assign n21689 = ~n21685 & n21688 ;
  assign n21690 = ( n4796 & n21684 ) | ( n4796 & n21689 ) | ( n21684 & n21689 ) ;
  assign n21691 = n9128 & ~n12765 ;
  assign n21692 = n13775 & n21691 ;
  assign n21693 = ( ~n19562 & n20375 ) | ( ~n19562 & n21692 ) | ( n20375 & n21692 ) ;
  assign n21696 = n14736 ^ n4875 ^ n626 ;
  assign n21695 = ( n3995 & ~n4213 ) | ( n3995 & n17576 ) | ( ~n4213 & n17576 ) ;
  assign n21697 = n21696 ^ n21695 ^ 1'b0 ;
  assign n21698 = n1190 & n21697 ;
  assign n21699 = n8667 & ~n18447 ;
  assign n21700 = ~n21698 & n21699 ;
  assign n21694 = ~n20854 & n21007 ;
  assign n21701 = n21700 ^ n21694 ^ 1'b0 ;
  assign n21702 = ( n3950 & n8431 ) | ( n3950 & ~n10655 ) | ( n8431 & ~n10655 ) ;
  assign n21703 = n6272 ^ n3156 ^ 1'b0 ;
  assign n21704 = ( n2838 & n21702 ) | ( n2838 & ~n21703 ) | ( n21702 & ~n21703 ) ;
  assign n21705 = n9191 ^ n6646 ^ 1'b0 ;
  assign n21706 = n18274 ^ n9553 ^ 1'b0 ;
  assign n21707 = ~n21705 & n21706 ;
  assign n21708 = n6828 ^ n2895 ^ 1'b0 ;
  assign n21709 = n21708 ^ n5225 ^ n2428 ;
  assign n21710 = ( n1553 & ~n21707 ) | ( n1553 & n21709 ) | ( ~n21707 & n21709 ) ;
  assign n21711 = n792 & ~n2545 ;
  assign n21712 = n5459 & n21711 ;
  assign n21713 = n21712 ^ n1145 ^ 1'b0 ;
  assign n21714 = ( ~n6578 & n6974 ) | ( ~n6578 & n12443 ) | ( n6974 & n12443 ) ;
  assign n21716 = n9835 ^ n4144 ^ 1'b0 ;
  assign n21717 = n10448 & ~n16840 ;
  assign n21718 = ~n21716 & n21717 ;
  assign n21719 = ( n6397 & n18427 ) | ( n6397 & ~n21718 ) | ( n18427 & ~n21718 ) ;
  assign n21715 = n16848 | n19158 ;
  assign n21720 = n21719 ^ n21715 ^ n5165 ;
  assign n21721 = ~n6026 & n18494 ;
  assign n21722 = n1062 & n21721 ;
  assign n21723 = n4767 | n14495 ;
  assign n21724 = n21722 & ~n21723 ;
  assign n21725 = n21724 ^ n3051 ^ 1'b0 ;
  assign n21726 = n15441 | n21725 ;
  assign n21727 = ( n12656 & n17805 ) | ( n12656 & ~n21726 ) | ( n17805 & ~n21726 ) ;
  assign n21728 = n3488 | n17354 ;
  assign n21729 = n21728 ^ n10814 ^ n326 ;
  assign n21730 = ( ~n4938 & n9100 ) | ( ~n4938 & n11290 ) | ( n9100 & n11290 ) ;
  assign n21731 = ( n17314 & n20627 ) | ( n17314 & ~n21730 ) | ( n20627 & ~n21730 ) ;
  assign n21733 = n17943 ^ n11846 ^ 1'b0 ;
  assign n21734 = n2534 & ~n21733 ;
  assign n21735 = n10941 ^ n9240 ^ 1'b0 ;
  assign n21736 = n12969 | n21735 ;
  assign n21737 = ( ~n18383 & n21734 ) | ( ~n18383 & n21736 ) | ( n21734 & n21736 ) ;
  assign n21732 = x83 & n19773 ;
  assign n21738 = n21737 ^ n21732 ^ 1'b0 ;
  assign n21739 = n308 | n7080 ;
  assign n21740 = n3085 ^ n1129 ^ 1'b0 ;
  assign n21741 = ( n9984 & ~n21393 ) | ( n9984 & n21740 ) | ( ~n21393 & n21740 ) ;
  assign n21743 = n5191 & ~n17729 ;
  assign n21744 = ~n337 & n21743 ;
  assign n21742 = n8936 & ~n16509 ;
  assign n21745 = n21744 ^ n21742 ^ n642 ;
  assign n21746 = n14987 | n21745 ;
  assign n21751 = ( ~n720 & n5907 ) | ( ~n720 & n21170 ) | ( n5907 & n21170 ) ;
  assign n21752 = n21751 ^ n9683 ^ n4962 ;
  assign n21753 = n21752 ^ n20632 ^ n9581 ;
  assign n21748 = n8601 ^ n543 ^ 1'b0 ;
  assign n21749 = ~n7444 & n21748 ;
  assign n21750 = n21749 ^ n6531 ^ n5046 ;
  assign n21747 = ~n6741 & n9779 ;
  assign n21754 = n21753 ^ n21750 ^ n21747 ;
  assign n21755 = ~n6895 & n11358 ;
  assign n21756 = n21755 ^ n9640 ^ 1'b0 ;
  assign n21757 = n21756 ^ n7327 ^ n4143 ;
  assign n21758 = n2256 & n4326 ;
  assign n21759 = n12214 | n15391 ;
  assign n21760 = n21758 & ~n21759 ;
  assign n21761 = n10162 | n12400 ;
  assign n21762 = n20251 | n21761 ;
  assign n21763 = n21762 ^ n15788 ^ 1'b0 ;
  assign n21764 = n10635 | n21221 ;
  assign n21765 = n1938 & ~n21764 ;
  assign n21766 = n8730 ^ n7994 ^ n7002 ;
  assign n21767 = n21766 ^ n15395 ^ n10059 ;
  assign n21768 = ~n1115 & n9079 ;
  assign n21769 = n21768 ^ n710 ^ 1'b0 ;
  assign n21770 = n21769 ^ n20205 ^ n3530 ;
  assign n21771 = n1762 & ~n18092 ;
  assign n21772 = n21771 ^ n9974 ^ 1'b0 ;
  assign n21773 = n2112 & ~n21772 ;
  assign n21774 = n18002 ^ n6860 ^ n4745 ;
  assign n21775 = n21774 ^ n17123 ^ 1'b0 ;
  assign n21776 = n21775 ^ n9563 ^ n5550 ;
  assign n21777 = ( ~n4112 & n8900 ) | ( ~n4112 & n21776 ) | ( n8900 & n21776 ) ;
  assign n21778 = ( n311 & n21773 ) | ( n311 & ~n21777 ) | ( n21773 & ~n21777 ) ;
  assign n21779 = n2040 ^ n1612 ^ 1'b0 ;
  assign n21780 = ( n2835 & n14711 ) | ( n2835 & n21779 ) | ( n14711 & n21779 ) ;
  assign n21781 = n5449 & ~n7446 ;
  assign n21782 = ~n7147 & n21781 ;
  assign n21783 = n14053 & n17323 ;
  assign n21784 = n17093 ^ n14860 ^ n4325 ;
  assign n21787 = ( x45 & ~n10469 ) | ( x45 & n15414 ) | ( ~n10469 & n15414 ) ;
  assign n21785 = n7089 ^ n3162 ^ 1'b0 ;
  assign n21786 = n15420 & n21785 ;
  assign n21788 = n21787 ^ n21786 ^ 1'b0 ;
  assign n21789 = ( n3747 & n3920 ) | ( n3747 & n21207 ) | ( n3920 & n21207 ) ;
  assign n21790 = n17517 ^ n14036 ^ n2493 ;
  assign n21791 = ( ~n2982 & n11031 ) | ( ~n2982 & n17764 ) | ( n11031 & n17764 ) ;
  assign n21792 = n5047 & n21791 ;
  assign n21793 = n18900 ^ n4461 ^ n3921 ;
  assign n21794 = ( ~n397 & n5356 ) | ( ~n397 & n21793 ) | ( n5356 & n21793 ) ;
  assign n21795 = n11391 ^ n3676 ^ n732 ;
  assign n21796 = ( ~n984 & n10415 ) | ( ~n984 & n21795 ) | ( n10415 & n21795 ) ;
  assign n21797 = ( n3028 & n5518 ) | ( n3028 & n21796 ) | ( n5518 & n21796 ) ;
  assign n21798 = n14040 & n21797 ;
  assign n21799 = n21798 ^ n2509 ^ 1'b0 ;
  assign n21800 = ( ~n2685 & n8146 ) | ( ~n2685 & n8290 ) | ( n8146 & n8290 ) ;
  assign n21802 = ~n2667 & n4917 ;
  assign n21803 = n3036 & n21802 ;
  assign n21804 = ( n7215 & ~n7663 ) | ( n7215 & n21803 ) | ( ~n7663 & n21803 ) ;
  assign n21801 = n2292 & n9109 ;
  assign n21805 = n21804 ^ n21801 ^ n20495 ;
  assign n21806 = n21344 ^ n4142 ^ 1'b0 ;
  assign n21807 = n2867 ^ n641 ^ 1'b0 ;
  assign n21808 = n1341 & ~n21807 ;
  assign n21809 = n21808 ^ n12384 ^ n10344 ;
  assign n21810 = n10235 ^ n861 ^ n412 ;
  assign n21811 = n13545 | n21810 ;
  assign n21812 = n16404 & ~n21811 ;
  assign n21813 = n11142 & n17758 ;
  assign n21817 = n13694 ^ n11099 ^ n2838 ;
  assign n21814 = n8125 ^ n4654 ^ n3273 ;
  assign n21815 = ~n7760 & n21814 ;
  assign n21816 = n21815 ^ n13174 ^ 1'b0 ;
  assign n21818 = n21817 ^ n21816 ^ x49 ;
  assign n21819 = ~n3874 & n9581 ;
  assign n21820 = ~n10219 & n21819 ;
  assign n21821 = n2409 & ~n10496 ;
  assign n21822 = n21821 ^ n6968 ^ 1'b0 ;
  assign n21823 = n3775 & n8771 ;
  assign n21824 = ( ~n4814 & n15613 ) | ( ~n4814 & n15971 ) | ( n15613 & n15971 ) ;
  assign n21825 = n21824 ^ n14911 ^ 1'b0 ;
  assign n21826 = ( ~n7288 & n18921 ) | ( ~n7288 & n20196 ) | ( n18921 & n20196 ) ;
  assign n21827 = n21826 ^ n1771 ^ 1'b0 ;
  assign n21828 = n16008 ^ n13457 ^ n8802 ;
  assign n21829 = n7526 ^ n4008 ^ n3225 ;
  assign n21830 = n18183 & ~n21829 ;
  assign n21831 = n10912 ^ n5585 ^ 1'b0 ;
  assign n21837 = n16570 ^ n11289 ^ 1'b0 ;
  assign n21838 = ~n633 & n21837 ;
  assign n21832 = n2424 | n13149 ;
  assign n21833 = n2075 | n21832 ;
  assign n21834 = n21833 ^ n9675 ^ n1186 ;
  assign n21835 = n1716 & ~n21834 ;
  assign n21836 = ( n2056 & ~n11508 ) | ( n2056 & n21835 ) | ( ~n11508 & n21835 ) ;
  assign n21839 = n21838 ^ n21836 ^ n10356 ;
  assign n21840 = n3516 & ~n21839 ;
  assign n21841 = n21840 ^ n3183 ^ 1'b0 ;
  assign n21842 = n13234 & n19231 ;
  assign n21843 = n21842 ^ n11467 ^ 1'b0 ;
  assign n21844 = n9934 ^ n6590 ^ 1'b0 ;
  assign n21845 = n12573 | n15635 ;
  assign n21846 = n11198 ^ n10365 ^ n8244 ;
  assign n21847 = ( n1548 & n14785 ) | ( n1548 & ~n17166 ) | ( n14785 & ~n17166 ) ;
  assign n21848 = n4534 & n14873 ;
  assign n21849 = n21848 ^ n20810 ^ 1'b0 ;
  assign n21850 = n16956 ^ n14065 ^ 1'b0 ;
  assign n21851 = ~n21849 & n21850 ;
  assign n21852 = n4535 & n21851 ;
  assign n21853 = n6975 ^ n5835 ^ n3537 ;
  assign n21854 = n990 & ~n21853 ;
  assign n21855 = n21854 ^ n1066 ^ 1'b0 ;
  assign n21856 = n18671 ^ n17250 ^ 1'b0 ;
  assign n21857 = ( n9404 & ~n16721 ) | ( n9404 & n21856 ) | ( ~n16721 & n21856 ) ;
  assign n21858 = n21857 ^ n15592 ^ n15203 ;
  assign n21859 = n21858 ^ n20611 ^ x74 ;
  assign n21860 = ( n626 & ~n1950 ) | ( n626 & n5073 ) | ( ~n1950 & n5073 ) ;
  assign n21861 = n21860 ^ n2317 ^ 1'b0 ;
  assign n21862 = ( n1126 & ~n12468 ) | ( n1126 & n14412 ) | ( ~n12468 & n14412 ) ;
  assign n21863 = ( ~n1901 & n5975 ) | ( ~n1901 & n10277 ) | ( n5975 & n10277 ) ;
  assign n21864 = ( n6300 & n6548 ) | ( n6300 & n17308 ) | ( n6548 & n17308 ) ;
  assign n21865 = ( n12320 & n21863 ) | ( n12320 & n21864 ) | ( n21863 & n21864 ) ;
  assign n21867 = ( n580 & n5434 ) | ( n580 & ~n8223 ) | ( n5434 & ~n8223 ) ;
  assign n21866 = n6425 | n11494 ;
  assign n21868 = n21867 ^ n21866 ^ n10012 ;
  assign n21869 = n15318 | n17641 ;
  assign n21870 = n15223 | n18989 ;
  assign n21872 = x120 & ~n12245 ;
  assign n21873 = n21872 ^ n1247 ^ 1'b0 ;
  assign n21871 = n20358 ^ n9545 ^ n4805 ;
  assign n21874 = n21873 ^ n21871 ^ 1'b0 ;
  assign n21875 = n21870 | n21874 ;
  assign n21876 = n12038 & ~n12130 ;
  assign n21880 = ~n3240 & n11469 ;
  assign n21881 = n6048 & n21880 ;
  assign n21877 = n11793 & ~n20316 ;
  assign n21878 = n21877 ^ n13445 ^ n3733 ;
  assign n21879 = n7190 & ~n21878 ;
  assign n21882 = n21881 ^ n21879 ^ 1'b0 ;
  assign n21883 = ( n12763 & n13249 ) | ( n12763 & ~n21882 ) | ( n13249 & ~n21882 ) ;
  assign n21884 = n7169 & n9580 ;
  assign n21885 = n21884 ^ x125 ^ 1'b0 ;
  assign n21886 = n10656 ^ n500 ^ 1'b0 ;
  assign n21887 = ~n1293 & n21886 ;
  assign n21888 = n21887 ^ n14958 ^ n14505 ;
  assign n21889 = n17198 & n21675 ;
  assign n21891 = n1486 | n4695 ;
  assign n21890 = n8354 | n8396 ;
  assign n21892 = n21891 ^ n21890 ^ 1'b0 ;
  assign n21893 = n17188 & ~n21892 ;
  assign n21894 = n12861 & n21893 ;
  assign n21895 = n19972 ^ n4234 ^ 1'b0 ;
  assign n21896 = ~n9821 & n21895 ;
  assign n21897 = ~n2681 & n3081 ;
  assign n21898 = n15406 & n21897 ;
  assign n21899 = n10924 | n11667 ;
  assign n21900 = n21899 ^ n2477 ^ 1'b0 ;
  assign n21901 = n3375 & n19505 ;
  assign n21902 = ( n10161 & n21270 ) | ( n10161 & n21901 ) | ( n21270 & n21901 ) ;
  assign n21904 = n3004 & ~n11149 ;
  assign n21903 = ( n1384 & ~n4378 ) | ( n1384 & n5042 ) | ( ~n4378 & n5042 ) ;
  assign n21905 = n21904 ^ n21903 ^ n7322 ;
  assign n21906 = n14347 ^ n6136 ^ n5701 ;
  assign n21907 = n21906 ^ n19271 ^ n14036 ;
  assign n21908 = n21907 ^ n14369 ^ 1'b0 ;
  assign n21909 = ~n4195 & n21908 ;
  assign n21910 = n10840 ^ n3174 ^ n562 ;
  assign n21911 = n20124 ^ n12449 ^ n5081 ;
  assign n21916 = n9144 & n12341 ;
  assign n21914 = n506 & ~n11118 ;
  assign n21915 = ~n17823 & n21914 ;
  assign n21912 = n14233 ^ n6460 ^ 1'b0 ;
  assign n21913 = n21912 ^ n20511 ^ 1'b0 ;
  assign n21917 = n21916 ^ n21915 ^ n21913 ;
  assign n21918 = n12419 | n20450 ;
  assign n21920 = n10639 & n13902 ;
  assign n21921 = n21920 ^ n8943 ^ n5827 ;
  assign n21919 = n9364 ^ n6780 ^ 1'b0 ;
  assign n21922 = n21921 ^ n21919 ^ 1'b0 ;
  assign n21923 = n21736 ^ n6561 ^ 1'b0 ;
  assign n21924 = n7407 | n21923 ;
  assign n21925 = ~n724 & n19703 ;
  assign n21926 = n21925 ^ n1982 ^ 1'b0 ;
  assign n21927 = n7291 ^ n6006 ^ 1'b0 ;
  assign n21928 = n5881 & n21927 ;
  assign n21929 = n16411 ^ n8814 ^ 1'b0 ;
  assign n21930 = n21577 ^ n11842 ^ n9204 ;
  assign n21931 = ( n2222 & n8281 ) | ( n2222 & n21930 ) | ( n8281 & n21930 ) ;
  assign n21932 = ( n3950 & n10308 ) | ( n3950 & ~n13196 ) | ( n10308 & ~n13196 ) ;
  assign n21933 = n13774 ^ n8505 ^ n5100 ;
  assign n21934 = n20622 ^ n14235 ^ n11151 ;
  assign n21935 = n15690 ^ n9912 ^ n8548 ;
  assign n21936 = ( n7525 & n12392 ) | ( n7525 & ~n21935 ) | ( n12392 & ~n21935 ) ;
  assign n21937 = ( n6658 & ~n12045 ) | ( n6658 & n21936 ) | ( ~n12045 & n21936 ) ;
  assign n21938 = n5629 & n21937 ;
  assign n21939 = n19711 ^ n16181 ^ n11955 ;
  assign n21940 = n21514 ^ n13490 ^ 1'b0 ;
  assign n21941 = n21939 & ~n21940 ;
  assign n21942 = n21826 ^ n7734 ^ 1'b0 ;
  assign n21943 = ( n2373 & n13185 ) | ( n2373 & n17396 ) | ( n13185 & n17396 ) ;
  assign n21944 = n21943 ^ n14633 ^ n8508 ;
  assign n21945 = ~n3896 & n6844 ;
  assign n21946 = ~n4010 & n21945 ;
  assign n21947 = n13650 & ~n21946 ;
  assign n21948 = n11305 & n21947 ;
  assign n21949 = ( n11757 & ~n19893 ) | ( n11757 & n21948 ) | ( ~n19893 & n21948 ) ;
  assign n21950 = n9003 ^ n6475 ^ 1'b0 ;
  assign n21951 = n21950 ^ n9675 ^ n9432 ;
  assign n21952 = n1589 & ~n7396 ;
  assign n21953 = n21545 & ~n21952 ;
  assign n21954 = n21953 ^ n9034 ^ 1'b0 ;
  assign n21955 = ~n4020 & n11453 ;
  assign n21956 = n1620 & ~n8504 ;
  assign n21957 = ~n2082 & n21956 ;
  assign n21958 = n21957 ^ n18819 ^ 1'b0 ;
  assign n21959 = n21955 & n21958 ;
  assign n21960 = n11634 ^ n7379 ^ n3597 ;
  assign n21961 = n21960 ^ n16667 ^ n3364 ;
  assign n21962 = n13035 ^ n7124 ^ n2057 ;
  assign n21963 = n13493 & n18634 ;
  assign n21964 = ~n21962 & n21963 ;
  assign n21965 = n21964 ^ n18329 ^ n13992 ;
  assign n21966 = n2969 ^ n562 ^ 1'b0 ;
  assign n21967 = ~n14807 & n21966 ;
  assign n21968 = n13168 & ~n21967 ;
  assign n21969 = n21968 ^ n11011 ^ 1'b0 ;
  assign n21970 = n14301 ^ n2402 ^ n1246 ;
  assign n21971 = n1306 & n2524 ;
  assign n21972 = ~n21970 & n21971 ;
  assign n21973 = n3880 & n8405 ;
  assign n21974 = n21973 ^ n2542 ^ 1'b0 ;
  assign n21975 = ( n16199 & ~n16555 ) | ( n16199 & n21974 ) | ( ~n16555 & n21974 ) ;
  assign n21976 = n15280 ^ n12856 ^ 1'b0 ;
  assign n21977 = ~n21975 & n21976 ;
  assign n21978 = n1648 & n2094 ;
  assign n21979 = n21978 ^ n15495 ^ 1'b0 ;
  assign n21980 = n6475 & n8441 ;
  assign n21981 = ~n4097 & n21980 ;
  assign n21982 = n11411 ^ n2438 ^ n2137 ;
  assign n21983 = ( ~n4418 & n10703 ) | ( ~n4418 & n16590 ) | ( n10703 & n16590 ) ;
  assign n21984 = ( n1301 & ~n21982 ) | ( n1301 & n21983 ) | ( ~n21982 & n21983 ) ;
  assign n21985 = n4649 ^ n2209 ^ 1'b0 ;
  assign n21986 = n18517 ^ n12160 ^ n9632 ;
  assign n21987 = ( n2599 & n21985 ) | ( n2599 & ~n21986 ) | ( n21985 & ~n21986 ) ;
  assign n21988 = n2493 & ~n2903 ;
  assign n21989 = n21988 ^ n16992 ^ 1'b0 ;
  assign n21990 = n3995 | n21989 ;
  assign n21991 = ( n531 & n2785 ) | ( n531 & ~n12675 ) | ( n2785 & ~n12675 ) ;
  assign n21992 = n10565 ^ n4198 ^ 1'b0 ;
  assign n21993 = n11317 & n21992 ;
  assign n21994 = n8473 ^ n8113 ^ 1'b0 ;
  assign n21995 = n21993 & n21994 ;
  assign n21996 = ~n12355 & n19001 ;
  assign n21997 = n10752 | n19564 ;
  assign n21998 = n21997 ^ n10745 ^ 1'b0 ;
  assign n21999 = ( x21 & ~n6723 ) | ( x21 & n21998 ) | ( ~n6723 & n21998 ) ;
  assign n22000 = n1172 & ~n1553 ;
  assign n22001 = n22000 ^ n607 ^ 1'b0 ;
  assign n22002 = n22001 ^ n6350 ^ 1'b0 ;
  assign n22003 = n18726 ^ n2716 ^ 1'b0 ;
  assign n22004 = n7681 & ~n21484 ;
  assign n22005 = n22004 ^ n3640 ^ 1'b0 ;
  assign n22006 = n22005 ^ n10927 ^ n8603 ;
  assign n22007 = n22006 ^ n8411 ^ n5934 ;
  assign n22008 = ( n3401 & n15024 ) | ( n3401 & ~n21916 ) | ( n15024 & ~n21916 ) ;
  assign n22009 = ~n7551 & n7668 ;
  assign n22010 = ~n621 & n22009 ;
  assign n22011 = n6295 & n22010 ;
  assign n22013 = n441 & n2367 ;
  assign n22012 = ~n6586 & n12664 ;
  assign n22014 = n22013 ^ n22012 ^ 1'b0 ;
  assign n22015 = n19564 ^ n7479 ^ 1'b0 ;
  assign n22016 = n11283 & ~n22015 ;
  assign n22017 = x12 & n13311 ;
  assign n22018 = ~n2373 & n22017 ;
  assign n22019 = ( ~n2383 & n2472 ) | ( ~n2383 & n22018 ) | ( n2472 & n22018 ) ;
  assign n22020 = n9646 & ~n18528 ;
  assign n22021 = ~n20137 & n22020 ;
  assign n22023 = n161 & ~n10688 ;
  assign n22024 = n22023 ^ n5177 ^ 1'b0 ;
  assign n22022 = n8674 ^ n3065 ^ 1'b0 ;
  assign n22025 = n22024 ^ n22022 ^ n8361 ;
  assign n22026 = ( n14396 & n20114 ) | ( n14396 & ~n22025 ) | ( n20114 & ~n22025 ) ;
  assign n22027 = ( n10006 & n11291 ) | ( n10006 & ~n16764 ) | ( n11291 & ~n16764 ) ;
  assign n22028 = n18740 ^ n16198 ^ n15664 ;
  assign n22029 = n15127 ^ n12772 ^ 1'b0 ;
  assign n22030 = n2304 | n15340 ;
  assign n22031 = n19781 & ~n22030 ;
  assign n22032 = n22031 ^ n8639 ^ 1'b0 ;
  assign n22033 = ( ~n2526 & n4230 ) | ( ~n2526 & n15225 ) | ( n4230 & n15225 ) ;
  assign n22034 = n22033 ^ n5297 ^ n5164 ;
  assign n22035 = n4452 | n8372 ;
  assign n22036 = n5898 ^ n1904 ^ 1'b0 ;
  assign n22037 = ( n7737 & ~n11556 ) | ( n7737 & n20355 ) | ( ~n11556 & n20355 ) ;
  assign n22038 = ( n5563 & n22036 ) | ( n5563 & ~n22037 ) | ( n22036 & ~n22037 ) ;
  assign n22039 = n8103 ^ n6767 ^ n5786 ;
  assign n22040 = n22039 ^ n11335 ^ n3804 ;
  assign n22041 = n15120 ^ n2086 ^ 1'b0 ;
  assign n22042 = n22041 ^ n13502 ^ 1'b0 ;
  assign n22043 = ~n5861 & n9087 ;
  assign n22044 = n22043 ^ n14432 ^ 1'b0 ;
  assign n22045 = n2509 | n8273 ;
  assign n22046 = n22045 ^ n2967 ^ 1'b0 ;
  assign n22047 = n15938 ^ n8157 ^ n5393 ;
  assign n22048 = n22047 ^ n20810 ^ n13146 ;
  assign n22049 = n11892 ^ n6256 ^ n1802 ;
  assign n22050 = n22049 ^ n14829 ^ x48 ;
  assign n22051 = n12701 ^ n6832 ^ 1'b0 ;
  assign n22052 = n836 & ~n4457 ;
  assign n22053 = ( n3285 & ~n16222 ) | ( n3285 & n17941 ) | ( ~n16222 & n17941 ) ;
  assign n22054 = n14478 ^ n7766 ^ n3583 ;
  assign n22057 = n13926 ^ n5374 ^ 1'b0 ;
  assign n22058 = n3422 | n22057 ;
  assign n22055 = n7856 ^ n1273 ^ 1'b0 ;
  assign n22056 = n3797 & ~n22055 ;
  assign n22059 = n22058 ^ n22056 ^ n10334 ;
  assign n22060 = n22059 ^ n12890 ^ n1059 ;
  assign n22061 = n5708 & ~n22060 ;
  assign n22062 = n22061 ^ n19302 ^ n15392 ;
  assign n22063 = ( n22053 & n22054 ) | ( n22053 & ~n22062 ) | ( n22054 & ~n22062 ) ;
  assign n22064 = n3797 & n11275 ;
  assign n22065 = n22064 ^ n5530 ^ 1'b0 ;
  assign n22066 = ( n1073 & n5891 ) | ( n1073 & ~n22065 ) | ( n5891 & ~n22065 ) ;
  assign n22067 = n19853 ^ n8870 ^ n1853 ;
  assign n22068 = n18756 & n22067 ;
  assign n22069 = n4100 | n7446 ;
  assign n22070 = n22069 ^ n356 ^ 1'b0 ;
  assign n22071 = n22070 ^ n4106 ^ n1740 ;
  assign n22072 = n19166 & ~n20411 ;
  assign n22073 = n937 & n13053 ;
  assign n22077 = n7477 | n11822 ;
  assign n22078 = n22077 ^ n16955 ^ 1'b0 ;
  assign n22079 = n22078 ^ n13893 ^ n9067 ;
  assign n22080 = n22079 ^ n6288 ^ 1'b0 ;
  assign n22081 = n1170 | n22080 ;
  assign n22074 = n21454 ^ n2072 ^ 1'b0 ;
  assign n22075 = n4491 | n22074 ;
  assign n22076 = n22075 ^ n14945 ^ 1'b0 ;
  assign n22082 = n22081 ^ n22076 ^ n17756 ;
  assign n22083 = ( ~n2075 & n2179 ) | ( ~n2075 & n2475 ) | ( n2179 & n2475 ) ;
  assign n22084 = n11173 & n22083 ;
  assign n22085 = n7758 | n22084 ;
  assign n22086 = ( ~n8521 & n10486 ) | ( ~n8521 & n10948 ) | ( n10486 & n10948 ) ;
  assign n22087 = ( n3796 & n10673 ) | ( n3796 & ~n13230 ) | ( n10673 & ~n13230 ) ;
  assign n22088 = n10897 & ~n20967 ;
  assign n22089 = n9140 | n18342 ;
  assign n22090 = n19933 | n22089 ;
  assign n22091 = n22090 ^ n21190 ^ 1'b0 ;
  assign n22092 = n5679 ^ n714 ^ n488 ;
  assign n22093 = ~n1157 & n22092 ;
  assign n22094 = n22091 & n22093 ;
  assign n22095 = n11585 ^ n2773 ^ n1280 ;
  assign n22096 = ~n7306 & n22095 ;
  assign n22097 = n7056 & ~n11159 ;
  assign n22098 = ( n1506 & ~n10555 ) | ( n1506 & n13394 ) | ( ~n10555 & n13394 ) ;
  assign n22099 = n22098 ^ n19038 ^ n5901 ;
  assign n22100 = n22099 ^ n4193 ^ n1272 ;
  assign n22101 = n5784 | n10533 ;
  assign n22102 = n22101 ^ n16147 ^ 1'b0 ;
  assign n22103 = n8156 ^ n7884 ^ n3286 ;
  assign n22104 = ( n6086 & n13292 ) | ( n6086 & n15386 ) | ( n13292 & n15386 ) ;
  assign n22105 = ( ~n696 & n1299 ) | ( ~n696 & n2130 ) | ( n1299 & n2130 ) ;
  assign n22106 = n399 | n22105 ;
  assign n22107 = n22106 ^ n14034 ^ 1'b0 ;
  assign n22108 = n11337 ^ n5928 ^ 1'b0 ;
  assign n22109 = n22107 & ~n22108 ;
  assign n22110 = ~n774 & n17077 ;
  assign n22111 = n684 & ~n22110 ;
  assign n22112 = ~n2178 & n22111 ;
  assign n22113 = n15496 | n18601 ;
  assign n22114 = n6546 ^ n2616 ^ n1816 ;
  assign n22115 = ( n10327 & n14050 ) | ( n10327 & ~n22114 ) | ( n14050 & ~n22114 ) ;
  assign n22116 = n2661 & ~n8096 ;
  assign n22117 = n22116 ^ n3258 ^ 1'b0 ;
  assign n22118 = ( n410 & n5186 ) | ( n410 & ~n22117 ) | ( n5186 & ~n22117 ) ;
  assign n22119 = n22118 ^ n11428 ^ 1'b0 ;
  assign n22120 = n22115 & n22119 ;
  assign n22121 = n22120 ^ n8599 ^ n3900 ;
  assign n22122 = n9119 & n16316 ;
  assign n22123 = n22122 ^ n5457 ^ 1'b0 ;
  assign n22124 = n22123 ^ n1847 ^ x29 ;
  assign n22125 = n22124 ^ n2491 ^ 1'b0 ;
  assign n22126 = ( ~n11443 & n21183 ) | ( ~n11443 & n22125 ) | ( n21183 & n22125 ) ;
  assign n22127 = n19898 & n22126 ;
  assign n22128 = n9898 ^ n8211 ^ n5203 ;
  assign n22129 = n12984 ^ n9128 ^ n6800 ;
  assign n22130 = n22129 ^ n14724 ^ n9451 ;
  assign n22131 = ( n3076 & n20759 ) | ( n3076 & n22130 ) | ( n20759 & n22130 ) ;
  assign n22132 = ( n729 & n4035 ) | ( n729 & n8157 ) | ( n4035 & n8157 ) ;
  assign n22133 = n11023 ^ n9769 ^ 1'b0 ;
  assign n22134 = ~n22132 & n22133 ;
  assign n22135 = ( ~n5198 & n12263 ) | ( ~n5198 & n12939 ) | ( n12263 & n12939 ) ;
  assign n22136 = ~n17875 & n22135 ;
  assign n22137 = ~n22134 & n22136 ;
  assign n22138 = n14437 ^ n4075 ^ 1'b0 ;
  assign n22139 = ~n3420 & n22138 ;
  assign n22140 = n13011 ^ n5941 ^ n3652 ;
  assign n22142 = n1355 & ~n4640 ;
  assign n22143 = n22142 ^ n1155 ^ 1'b0 ;
  assign n22141 = ( n3088 & n6153 ) | ( n3088 & ~n21167 ) | ( n6153 & ~n21167 ) ;
  assign n22144 = n22143 ^ n22141 ^ n2577 ;
  assign n22145 = ~n4399 & n6810 ;
  assign n22146 = n22145 ^ n11125 ^ 1'b0 ;
  assign n22147 = ~n6712 & n22146 ;
  assign n22148 = n22147 ^ n1557 ^ 1'b0 ;
  assign n22149 = ~n15723 & n22148 ;
  assign n22150 = ~n11618 & n18011 ;
  assign n22151 = n17406 & n22150 ;
  assign n22152 = ~n3836 & n11504 ;
  assign n22153 = n5585 & n22152 ;
  assign n22154 = n4084 | n17656 ;
  assign n22155 = n13405 & ~n22154 ;
  assign n22156 = n2334 & n12327 ;
  assign n22157 = ~n12265 & n22156 ;
  assign n22158 = n22157 ^ n13929 ^ 1'b0 ;
  assign n22159 = n923 & ~n22158 ;
  assign n22160 = n22159 ^ n20208 ^ n7550 ;
  assign n22161 = n3204 & n4216 ;
  assign n22162 = n11223 & n22161 ;
  assign n22163 = n6039 | n22162 ;
  assign n22164 = n11807 ^ n681 ^ 1'b0 ;
  assign n22165 = n18601 & n22164 ;
  assign n22166 = n22165 ^ n19337 ^ n9093 ;
  assign n22167 = ( x58 & x121 ) | ( x58 & n5098 ) | ( x121 & n5098 ) ;
  assign n22168 = n9255 ^ n4910 ^ 1'b0 ;
  assign n22169 = n12145 & ~n22168 ;
  assign n22170 = n6972 | n15097 ;
  assign n22171 = ~n18562 & n22170 ;
  assign n22172 = n22171 ^ n12121 ^ 1'b0 ;
  assign n22173 = n5401 | n7250 ;
  assign n22174 = ( ~n2190 & n14679 ) | ( ~n2190 & n22173 ) | ( n14679 & n22173 ) ;
  assign n22175 = n21775 ^ n6327 ^ n6265 ;
  assign n22176 = ( n7193 & n7518 ) | ( n7193 & ~n20738 ) | ( n7518 & ~n20738 ) ;
  assign n22177 = ( ~n3602 & n8639 ) | ( ~n3602 & n22176 ) | ( n8639 & n22176 ) ;
  assign n22178 = n11925 & n21332 ;
  assign n22179 = ~n22177 & n22178 ;
  assign n22180 = ( n289 & n12273 ) | ( n289 & n22179 ) | ( n12273 & n22179 ) ;
  assign n22181 = ~n1960 & n11646 ;
  assign n22182 = n22181 ^ n1137 ^ 1'b0 ;
  assign n22183 = n7414 & ~n22182 ;
  assign n22184 = n17365 & n22183 ;
  assign n22186 = n199 & n7608 ;
  assign n22187 = n9332 & n22186 ;
  assign n22188 = n22187 ^ n11886 ^ n2357 ;
  assign n22185 = n1475 & n5887 ;
  assign n22189 = n22188 ^ n22185 ^ 1'b0 ;
  assign n22190 = n5642 & n22189 ;
  assign n22191 = ~n374 & n22190 ;
  assign n22192 = n22184 & ~n22191 ;
  assign n22194 = n722 & n1916 ;
  assign n22193 = n9230 & n16851 ;
  assign n22195 = n22194 ^ n22193 ^ 1'b0 ;
  assign n22196 = ~n6103 & n7408 ;
  assign n22197 = ( n649 & n21311 ) | ( n649 & n22196 ) | ( n21311 & n22196 ) ;
  assign n22198 = ~n8695 & n9501 ;
  assign n22199 = n22198 ^ n5288 ^ 1'b0 ;
  assign n22200 = n2652 & n13258 ;
  assign n22201 = n3303 & n14505 ;
  assign n22202 = ~n3754 & n22201 ;
  assign n22203 = n9938 ^ n6108 ^ n2021 ;
  assign n22204 = n22203 ^ n1486 ^ 1'b0 ;
  assign n22205 = ( n11440 & n11833 ) | ( n11440 & n18043 ) | ( n11833 & n18043 ) ;
  assign n22208 = n566 ^ n315 ^ 1'b0 ;
  assign n22209 = n466 & ~n22208 ;
  assign n22210 = ( ~n13400 & n15218 ) | ( ~n13400 & n22209 ) | ( n15218 & n22209 ) ;
  assign n22206 = n10964 ^ n6657 ^ 1'b0 ;
  assign n22207 = ~n1849 & n22206 ;
  assign n22211 = n22210 ^ n22207 ^ n6548 ;
  assign n22212 = n21853 | n22211 ;
  assign n22213 = ( n12212 & n13474 ) | ( n12212 & ~n20559 ) | ( n13474 & ~n20559 ) ;
  assign n22214 = n22213 ^ n6013 ^ 1'b0 ;
  assign n22215 = n22214 ^ n5480 ^ 1'b0 ;
  assign n22216 = n2239 ^ n2033 ^ 1'b0 ;
  assign n22218 = ~n10999 & n19036 ;
  assign n22217 = n13079 ^ n2342 ^ 1'b0 ;
  assign n22219 = n22218 ^ n22217 ^ n12771 ;
  assign n22220 = n19532 ^ n5936 ^ n697 ;
  assign n22221 = ~n3445 & n8426 ;
  assign n22222 = n22221 ^ n20849 ^ 1'b0 ;
  assign n22223 = n8269 | n22222 ;
  assign n22224 = n6827 ^ n6485 ^ n3738 ;
  assign n22225 = n3659 & n22224 ;
  assign n22226 = n15170 | n20686 ;
  assign n22227 = n9697 | n22226 ;
  assign n22228 = n17381 ^ n14043 ^ n6580 ;
  assign n22229 = n22076 ^ n15334 ^ n7256 ;
  assign n22230 = n4141 ^ n2834 ^ 1'b0 ;
  assign n22231 = n22230 ^ n17391 ^ n15951 ;
  assign n22232 = n2744 & ~n5386 ;
  assign n22233 = ( n5674 & ~n7681 ) | ( n5674 & n22232 ) | ( ~n7681 & n22232 ) ;
  assign n22234 = n12745 ^ n8311 ^ 1'b0 ;
  assign n22235 = n21841 & ~n22234 ;
  assign n22236 = n22233 & n22235 ;
  assign n22237 = ( n335 & n5125 ) | ( n335 & ~n22236 ) | ( n5125 & ~n22236 ) ;
  assign n22238 = n2150 | n10948 ;
  assign n22239 = n22238 ^ n8044 ^ 1'b0 ;
  assign n22240 = n5881 & ~n22239 ;
  assign n22241 = n22240 ^ n16385 ^ 1'b0 ;
  assign n22242 = n12661 & n13488 ;
  assign n22243 = n22242 ^ n3553 ^ 1'b0 ;
  assign n22246 = n847 & ~n7601 ;
  assign n22247 = ~n5714 & n22246 ;
  assign n22244 = n15970 ^ n6515 ^ 1'b0 ;
  assign n22245 = ( ~n8770 & n12198 ) | ( ~n8770 & n22244 ) | ( n12198 & n22244 ) ;
  assign n22248 = n22247 ^ n22245 ^ 1'b0 ;
  assign n22249 = n5264 & n9175 ;
  assign n22250 = ( n6409 & n11531 ) | ( n6409 & ~n22249 ) | ( n11531 & ~n22249 ) ;
  assign n22251 = n7851 | n22250 ;
  assign n22252 = n22248 | n22251 ;
  assign n22253 = n4406 & n5253 ;
  assign n22254 = n12292 | n22253 ;
  assign n22255 = n8364 ^ n7122 ^ n5659 ;
  assign n22256 = ~n2089 & n7359 ;
  assign n22257 = ( n14594 & n22255 ) | ( n14594 & ~n22256 ) | ( n22255 & ~n22256 ) ;
  assign n22258 = ( n5592 & n6017 ) | ( n5592 & n6481 ) | ( n6017 & n6481 ) ;
  assign n22259 = n22258 ^ n14445 ^ n13800 ;
  assign n22260 = ( n4214 & ~n8551 ) | ( n4214 & n22259 ) | ( ~n8551 & n22259 ) ;
  assign n22261 = n5879 ^ n393 ^ 1'b0 ;
  assign n22262 = n22261 ^ n1911 ^ n853 ;
  assign n22263 = n11080 ^ n6692 ^ 1'b0 ;
  assign n22265 = n2560 & ~n5763 ;
  assign n22266 = n16316 & n22265 ;
  assign n22267 = n5887 & n22266 ;
  assign n22268 = ( ~n4812 & n7379 ) | ( ~n4812 & n22267 ) | ( n7379 & n22267 ) ;
  assign n22264 = n20950 ^ n2076 ^ n1160 ;
  assign n22269 = n22268 ^ n22264 ^ n18026 ;
  assign n22270 = ( ~n3575 & n3761 ) | ( ~n3575 & n6331 ) | ( n3761 & n6331 ) ;
  assign n22271 = ( n2204 & n17024 ) | ( n2204 & ~n22270 ) | ( n17024 & ~n22270 ) ;
  assign n22272 = ( ~n13741 & n19891 ) | ( ~n13741 & n22271 ) | ( n19891 & n22271 ) ;
  assign n22273 = ~n8260 & n14302 ;
  assign n22274 = n22273 ^ x68 ^ 1'b0 ;
  assign n22275 = n5333 & ~n11771 ;
  assign n22276 = n18134 & n22275 ;
  assign n22277 = ( ~n14134 & n16422 ) | ( ~n14134 & n16896 ) | ( n16422 & n16896 ) ;
  assign n22278 = n4501 | n22277 ;
  assign n22279 = n22278 ^ n16760 ^ 1'b0 ;
  assign n22287 = ( n2008 & ~n3575 ) | ( n2008 & n4946 ) | ( ~n3575 & n4946 ) ;
  assign n22283 = n14445 ^ n2589 ^ 1'b0 ;
  assign n22284 = n8873 | n22283 ;
  assign n22285 = n9735 | n22284 ;
  assign n22286 = ( n11062 & n14794 ) | ( n11062 & n22285 ) | ( n14794 & n22285 ) ;
  assign n22281 = n2565 ^ n1475 ^ 1'b0 ;
  assign n22280 = n18813 ^ n17066 ^ n3374 ;
  assign n22282 = n22281 ^ n22280 ^ n2358 ;
  assign n22288 = n22287 ^ n22286 ^ n22282 ;
  assign n22289 = n2095 | n16509 ;
  assign n22290 = n22289 ^ n556 ^ n153 ;
  assign n22291 = n9115 | n20470 ;
  assign n22292 = n13670 ^ n11428 ^ n8023 ;
  assign n22293 = ( n10775 & ~n22291 ) | ( n10775 & n22292 ) | ( ~n22291 & n22292 ) ;
  assign n22294 = ~n3650 & n11453 ;
  assign n22295 = n5019 & n22294 ;
  assign n22296 = ( n12554 & n21387 ) | ( n12554 & n22295 ) | ( n21387 & n22295 ) ;
  assign n22297 = ( n9481 & n13073 ) | ( n9481 & n22296 ) | ( n13073 & n22296 ) ;
  assign n22298 = n4983 ^ n3817 ^ n1028 ;
  assign n22299 = n9827 ^ n6584 ^ 1'b0 ;
  assign n22300 = ~n22298 & n22299 ;
  assign n22301 = ( n10911 & n19845 ) | ( n10911 & ~n22300 ) | ( n19845 & ~n22300 ) ;
  assign n22302 = n22301 ^ n11786 ^ 1'b0 ;
  assign n22303 = ( ~n16988 & n18098 ) | ( ~n16988 & n22302 ) | ( n18098 & n22302 ) ;
  assign n22304 = n15238 ^ n11292 ^ 1'b0 ;
  assign n22305 = n1148 & ~n11888 ;
  assign n22306 = n22305 ^ n2769 ^ 1'b0 ;
  assign n22307 = n9700 | n22306 ;
  assign n22308 = n16220 ^ n14313 ^ n13962 ;
  assign n22309 = n6326 ^ n2504 ^ n2227 ;
  assign n22310 = n22309 ^ n2277 ^ n1497 ;
  assign n22311 = ( n9577 & n16077 ) | ( n9577 & ~n22310 ) | ( n16077 & ~n22310 ) ;
  assign n22312 = ~n1023 & n16205 ;
  assign n22313 = ( ~n5214 & n10779 ) | ( ~n5214 & n22312 ) | ( n10779 & n22312 ) ;
  assign n22314 = ~n7510 & n9124 ;
  assign n22315 = n6445 & ~n21411 ;
  assign n22316 = n22315 ^ n16256 ^ 1'b0 ;
  assign n22317 = n2934 ^ n2746 ^ 1'b0 ;
  assign n22318 = n6416 & ~n22317 ;
  assign n22319 = n22318 ^ n6284 ^ 1'b0 ;
  assign n22320 = n18556 & ~n22319 ;
  assign n22321 = n22320 ^ n9187 ^ 1'b0 ;
  assign n22322 = ( n1422 & n1908 ) | ( n1422 & n7337 ) | ( n1908 & n7337 ) ;
  assign n22324 = ( n1742 & ~n7052 ) | ( n1742 & n7839 ) | ( ~n7052 & n7839 ) ;
  assign n22325 = ( n18104 & ~n21578 ) | ( n18104 & n22324 ) | ( ~n21578 & n22324 ) ;
  assign n22326 = n2543 & ~n22325 ;
  assign n22327 = ( n3900 & n21966 ) | ( n3900 & n22326 ) | ( n21966 & n22326 ) ;
  assign n22323 = n22098 ^ n18153 ^ 1'b0 ;
  assign n22328 = n22327 ^ n22323 ^ n1355 ;
  assign n22329 = n22328 ^ n9490 ^ n9159 ;
  assign n22330 = n509 & n1991 ;
  assign n22331 = n9692 & n22330 ;
  assign n22332 = n22331 ^ n20265 ^ n13788 ;
  assign n22333 = ( n3163 & n16186 ) | ( n3163 & n22332 ) | ( n16186 & n22332 ) ;
  assign n22334 = n1858 & n6115 ;
  assign n22335 = n22334 ^ n3456 ^ 1'b0 ;
  assign n22336 = n22335 ^ n1765 ^ 1'b0 ;
  assign n22337 = ~n21626 & n22336 ;
  assign n22338 = n8591 ^ n4658 ^ 1'b0 ;
  assign n22339 = ~n11237 & n22338 ;
  assign n22343 = n6972 ^ n1443 ^ n376 ;
  assign n22344 = n22343 ^ n5487 ^ n4480 ;
  assign n22342 = n5989 & n8234 ;
  assign n22345 = n22344 ^ n22342 ^ 1'b0 ;
  assign n22340 = n15865 & n20428 ;
  assign n22341 = ( ~n2386 & n16305 ) | ( ~n2386 & n22340 ) | ( n16305 & n22340 ) ;
  assign n22346 = n22345 ^ n22341 ^ n10018 ;
  assign n22347 = n1933 ^ n351 ^ 1'b0 ;
  assign n22348 = n3504 ^ n680 ^ 1'b0 ;
  assign n22349 = n11548 & ~n22348 ;
  assign n22350 = ~n22347 & n22349 ;
  assign n22351 = ( ~n11634 & n15420 ) | ( ~n11634 & n22350 ) | ( n15420 & n22350 ) ;
  assign n22352 = ( ~x45 & n4377 ) | ( ~x45 & n11297 ) | ( n4377 & n11297 ) ;
  assign n22353 = n19211 ^ n9358 ^ 1'b0 ;
  assign n22354 = n7676 & ~n22353 ;
  assign n22355 = n22354 ^ n15694 ^ n926 ;
  assign n22356 = n22352 & ~n22355 ;
  assign n22357 = n21771 ^ n8190 ^ 1'b0 ;
  assign n22358 = n19354 | n22357 ;
  assign n22359 = n20175 ^ n4497 ^ 1'b0 ;
  assign n22360 = ~n6586 & n22359 ;
  assign n22361 = n2819 & ~n8950 ;
  assign n22362 = n22361 ^ n10313 ^ 1'b0 ;
  assign n22368 = n17763 ^ n15107 ^ 1'b0 ;
  assign n22369 = n2265 | n22368 ;
  assign n22365 = n5611 ^ n4105 ^ 1'b0 ;
  assign n22363 = n6315 & ~n11075 ;
  assign n22364 = n22363 ^ x44 ^ 1'b0 ;
  assign n22366 = n22365 ^ n22364 ^ n5458 ;
  assign n22367 = n5220 & ~n22366 ;
  assign n22370 = n22369 ^ n22367 ^ n13311 ;
  assign n22373 = ~n10716 & n18367 ;
  assign n22371 = n11262 ^ n2037 ^ 1'b0 ;
  assign n22372 = ~n2026 & n22371 ;
  assign n22374 = n22373 ^ n22372 ^ 1'b0 ;
  assign n22375 = n3085 | n19602 ;
  assign n22376 = ( ~n3183 & n4666 ) | ( ~n3183 & n6737 ) | ( n4666 & n6737 ) ;
  assign n22377 = n22376 ^ n8105 ^ 1'b0 ;
  assign n22378 = n5332 & ~n22377 ;
  assign n22379 = ( n15593 & ~n22375 ) | ( n15593 & n22378 ) | ( ~n22375 & n22378 ) ;
  assign n22380 = ~n2981 & n18445 ;
  assign n22381 = n22380 ^ n14501 ^ 1'b0 ;
  assign n22382 = n20658 ^ n9304 ^ 1'b0 ;
  assign n22383 = ( n7722 & ~n16837 ) | ( n7722 & n22382 ) | ( ~n16837 & n22382 ) ;
  assign n22384 = ~n10659 & n12663 ;
  assign n22385 = n22383 & n22384 ;
  assign n22387 = ~n3571 & n10989 ;
  assign n22386 = n291 | n503 ;
  assign n22388 = n22387 ^ n22386 ^ 1'b0 ;
  assign n22389 = n12765 ^ n3787 ^ n503 ;
  assign n22390 = n22389 ^ n14877 ^ n5519 ;
  assign n22391 = n9140 ^ n6733 ^ n3180 ;
  assign n22392 = ( n14722 & ~n19536 ) | ( n14722 & n22391 ) | ( ~n19536 & n22391 ) ;
  assign n22393 = n12592 ^ n6840 ^ 1'b0 ;
  assign n22394 = n19580 ^ n10045 ^ 1'b0 ;
  assign n22395 = n1896 & n22394 ;
  assign n22396 = n22395 ^ n2067 ^ 1'b0 ;
  assign n22397 = ~n11846 & n22396 ;
  assign n22398 = ~n4723 & n17923 ;
  assign n22399 = n1341 & ~n11504 ;
  assign n22400 = n757 & n22399 ;
  assign n22401 = n5665 & n10753 ;
  assign n22402 = n22401 ^ n4474 ^ 1'b0 ;
  assign n22403 = n2855 | n22402 ;
  assign n22404 = ~n7671 & n21702 ;
  assign n22405 = n22403 & n22404 ;
  assign n22406 = ( n2653 & n7424 ) | ( n2653 & ~n22405 ) | ( n7424 & ~n22405 ) ;
  assign n22407 = n22221 ^ n18094 ^ n10659 ;
  assign n22408 = n1709 & ~n2023 ;
  assign n22409 = n4392 ^ n844 ^ 1'b0 ;
  assign n22410 = ~n22408 & n22409 ;
  assign n22411 = ~n1419 & n22410 ;
  assign n22412 = ~n2983 & n12274 ;
  assign n22413 = n9662 ^ n5647 ^ 1'b0 ;
  assign n22414 = ~n18895 & n22413 ;
  assign n22415 = n11269 & n12248 ;
  assign n22416 = n22415 ^ n1636 ^ 1'b0 ;
  assign n22417 = n11313 ^ n7792 ^ 1'b0 ;
  assign n22418 = n6254 | n22417 ;
  assign n22419 = n2445 | n7795 ;
  assign n22420 = n22419 ^ n11162 ^ 1'b0 ;
  assign n22421 = ~n14148 & n15608 ;
  assign n22422 = n22421 ^ n6271 ^ 1'b0 ;
  assign n22423 = n622 & ~n10634 ;
  assign n22424 = n22423 ^ n5153 ^ 1'b0 ;
  assign n22425 = ~n19728 & n22424 ;
  assign n22426 = ( n21196 & ~n22422 ) | ( n21196 & n22425 ) | ( ~n22422 & n22425 ) ;
  assign n22427 = n18517 & ~n18913 ;
  assign n22428 = ~n2565 & n22427 ;
  assign n22429 = n22428 ^ n17721 ^ n924 ;
  assign n22430 = ( n8486 & ~n17563 ) | ( n8486 & n22429 ) | ( ~n17563 & n22429 ) ;
  assign n22431 = n10776 ^ n7781 ^ n3284 ;
  assign n22432 = n16173 ^ n11694 ^ n3078 ;
  assign n22433 = n22432 ^ n12400 ^ 1'b0 ;
  assign n22434 = n7504 & n22433 ;
  assign n22435 = n22434 ^ n20528 ^ 1'b0 ;
  assign n22436 = n7003 ^ n3763 ^ 1'b0 ;
  assign n22437 = n3628 | n22436 ;
  assign n22438 = n22437 ^ n20205 ^ 1'b0 ;
  assign n22439 = n4736 & n22438 ;
  assign n22442 = n7472 & ~n8868 ;
  assign n22443 = n22442 ^ n15880 ^ 1'b0 ;
  assign n22440 = n7747 & ~n13012 ;
  assign n22441 = ~n5785 & n22440 ;
  assign n22444 = n22443 ^ n22441 ^ n14421 ;
  assign n22445 = n20249 ^ n5539 ^ 1'b0 ;
  assign n22446 = ~n22444 & n22445 ;
  assign n22448 = n19477 ^ n19220 ^ n10573 ;
  assign n22447 = ( n8413 & n10472 ) | ( n8413 & n12130 ) | ( n10472 & n12130 ) ;
  assign n22449 = n22448 ^ n22447 ^ 1'b0 ;
  assign n22450 = n22449 ^ n18024 ^ n2279 ;
  assign n22451 = n5957 | n7052 ;
  assign n22452 = n22451 ^ n10090 ^ 1'b0 ;
  assign n22453 = n22452 ^ n21441 ^ 1'b0 ;
  assign n22454 = n13498 ^ n13223 ^ n10005 ;
  assign n22455 = n22454 ^ n4982 ^ n1078 ;
  assign n22456 = n16052 ^ n5225 ^ n532 ;
  assign n22458 = n2310 | n2671 ;
  assign n22459 = n22458 ^ n4896 ^ n3797 ;
  assign n22460 = ( n2747 & n6108 ) | ( n2747 & ~n22459 ) | ( n6108 & ~n22459 ) ;
  assign n22457 = ~n13974 & n16670 ;
  assign n22461 = n22460 ^ n22457 ^ 1'b0 ;
  assign n22462 = n5522 & ~n22461 ;
  assign n22463 = n4956 & n14433 ;
  assign n22464 = n4381 & ~n6056 ;
  assign n22465 = n22464 ^ n2629 ^ 1'b0 ;
  assign n22468 = n5425 & n9952 ;
  assign n22469 = ~n3424 & n22468 ;
  assign n22466 = n1875 & ~n5575 ;
  assign n22467 = n22466 ^ x5 ^ 1'b0 ;
  assign n22470 = n22469 ^ n22467 ^ n17587 ;
  assign n22471 = n15314 ^ n8711 ^ n6447 ;
  assign n22475 = ( n3013 & n6832 ) | ( n3013 & n7273 ) | ( n6832 & n7273 ) ;
  assign n22472 = n13621 & n14626 ;
  assign n22473 = n1019 & n22472 ;
  assign n22474 = n22473 ^ n13027 ^ 1'b0 ;
  assign n22476 = n22475 ^ n22474 ^ n18181 ;
  assign n22477 = ~n4536 & n20871 ;
  assign n22478 = n1318 & ~n19507 ;
  assign n22479 = n22478 ^ n4794 ^ 1'b0 ;
  assign n22480 = ( ~n3182 & n22477 ) | ( ~n3182 & n22479 ) | ( n22477 & n22479 ) ;
  assign n22481 = ( n16069 & ~n16909 ) | ( n16069 & n22480 ) | ( ~n16909 & n22480 ) ;
  assign n22482 = ( n6741 & ~n10447 ) | ( n6741 & n12365 ) | ( ~n10447 & n12365 ) ;
  assign n22483 = n16548 | n22482 ;
  assign n22484 = n11289 ^ n5309 ^ 1'b0 ;
  assign n22485 = n2081 & n22484 ;
  assign n22486 = n10878 ^ n8212 ^ 1'b0 ;
  assign n22487 = n22486 ^ n17281 ^ n6770 ;
  assign n22488 = ( n11450 & ~n20906 ) | ( n11450 & n22487 ) | ( ~n20906 & n22487 ) ;
  assign n22489 = n22488 ^ n15852 ^ 1'b0 ;
  assign n22490 = n22485 & ~n22489 ;
  assign n22491 = n3247 ^ n846 ^ 1'b0 ;
  assign n22492 = n3242 & n22491 ;
  assign n22493 = n22492 ^ n3462 ^ 1'b0 ;
  assign n22494 = n17375 ^ n12091 ^ n11726 ;
  assign n22495 = n13026 ^ n8576 ^ 1'b0 ;
  assign n22496 = n22494 & ~n22495 ;
  assign n22497 = n16417 ^ n14073 ^ 1'b0 ;
  assign n22498 = n9471 & ~n20692 ;
  assign n22499 = ( n4354 & n21103 ) | ( n4354 & ~n22498 ) | ( n21103 & ~n22498 ) ;
  assign n22500 = ~n2341 & n9469 ;
  assign n22501 = ~n15256 & n22500 ;
  assign n22502 = ( n2656 & ~n19308 ) | ( n2656 & n22501 ) | ( ~n19308 & n22501 ) ;
  assign n22503 = n19909 & ~n20885 ;
  assign n22504 = n22503 ^ n8721 ^ 1'b0 ;
  assign n22506 = n10824 ^ n2100 ^ 1'b0 ;
  assign n22507 = n566 | n22506 ;
  assign n22505 = n13761 | n14276 ;
  assign n22508 = n22507 ^ n22505 ^ n1307 ;
  assign n22510 = ( n1745 & n10020 ) | ( n1745 & n15718 ) | ( n10020 & n15718 ) ;
  assign n22509 = n1725 | n3474 ;
  assign n22511 = n22510 ^ n22509 ^ 1'b0 ;
  assign n22512 = n5510 & n14036 ;
  assign n22513 = n22512 ^ n16808 ^ 1'b0 ;
  assign n22514 = n19040 ^ n2103 ^ 1'b0 ;
  assign n22515 = ( n6369 & ~n11386 ) | ( n6369 & n22514 ) | ( ~n11386 & n22514 ) ;
  assign n22520 = n7820 ^ n3719 ^ 1'b0 ;
  assign n22516 = ( x2 & ~n172 ) | ( x2 & n4553 ) | ( ~n172 & n4553 ) ;
  assign n22517 = n3011 ^ n1832 ^ n1279 ;
  assign n22518 = ( n2826 & n22516 ) | ( n2826 & ~n22517 ) | ( n22516 & ~n22517 ) ;
  assign n22519 = n5506 | n22518 ;
  assign n22521 = n22520 ^ n22519 ^ x38 ;
  assign n22522 = x47 & ~n1791 ;
  assign n22523 = n22522 ^ n2187 ^ 1'b0 ;
  assign n22524 = n14753 & ~n22523 ;
  assign n22525 = ( n13459 & n13705 ) | ( n13459 & ~n22524 ) | ( n13705 & ~n22524 ) ;
  assign n22526 = n5589 ^ n726 ^ n387 ;
  assign n22527 = n13933 & ~n22526 ;
  assign n22528 = n5312 & ~n9331 ;
  assign n22529 = n22528 ^ n2917 ^ 1'b0 ;
  assign n22530 = ~n11897 & n22529 ;
  assign n22531 = n10383 ^ n7596 ^ n2659 ;
  assign n22533 = n1778 ^ n1669 ^ n219 ;
  assign n22534 = n22533 ^ n4948 ^ 1'b0 ;
  assign n22535 = n9829 | n22534 ;
  assign n22536 = n12961 | n22535 ;
  assign n22532 = n10288 ^ n8261 ^ 1'b0 ;
  assign n22537 = n22536 ^ n22532 ^ n656 ;
  assign n22538 = n13174 ^ n11611 ^ 1'b0 ;
  assign n22539 = n3920 | n22538 ;
  assign n22540 = x63 & ~n1136 ;
  assign n22541 = n22540 ^ n6462 ^ 1'b0 ;
  assign n22542 = ( n1790 & n2819 ) | ( n1790 & n9205 ) | ( n2819 & n9205 ) ;
  assign n22543 = ( n10937 & n22541 ) | ( n10937 & n22542 ) | ( n22541 & n22542 ) ;
  assign n22544 = n15971 ^ n10404 ^ n10256 ;
  assign n22545 = n22544 ^ n7268 ^ n4875 ;
  assign n22546 = n2254 & ~n11693 ;
  assign n22547 = n22546 ^ n1715 ^ n1399 ;
  assign n22548 = ~n3910 & n22547 ;
  assign n22549 = ( x104 & n3690 ) | ( x104 & n14663 ) | ( n3690 & n14663 ) ;
  assign n22556 = ( n432 & n2802 ) | ( n432 & n16517 ) | ( n2802 & n16517 ) ;
  assign n22550 = n3202 & n7484 ;
  assign n22551 = n22550 ^ n5383 ^ 1'b0 ;
  assign n22552 = n4486 | n7911 ;
  assign n22553 = n21262 & n22552 ;
  assign n22554 = n22553 ^ n12311 ^ 1'b0 ;
  assign n22555 = ( ~n15051 & n22551 ) | ( ~n15051 & n22554 ) | ( n22551 & n22554 ) ;
  assign n22557 = n22556 ^ n22555 ^ n11810 ;
  assign n22558 = n2363 & ~n18588 ;
  assign n22559 = n8369 & n22558 ;
  assign n22560 = n20356 & ~n22559 ;
  assign n22561 = n22560 ^ x72 ^ 1'b0 ;
  assign n22562 = n10319 & ~n22561 ;
  assign n22563 = n15809 & n22562 ;
  assign n22564 = n13398 ^ n8603 ^ 1'b0 ;
  assign n22565 = n3273 & ~n22564 ;
  assign n22566 = n10666 ^ n9795 ^ 1'b0 ;
  assign n22567 = n16287 & n20364 ;
  assign n22568 = ( n3653 & n11341 ) | ( n3653 & ~n14040 ) | ( n11341 & ~n14040 ) ;
  assign n22569 = n2496 & ~n11156 ;
  assign n22570 = ~n17377 & n22569 ;
  assign n22571 = n17493 ^ n3057 ^ 1'b0 ;
  assign n22572 = n2914 | n22571 ;
  assign n22573 = n22572 ^ n10656 ^ n8240 ;
  assign n22574 = n22573 ^ n8389 ^ 1'b0 ;
  assign n22575 = n13411 & n22574 ;
  assign n22576 = n9282 & ~n9491 ;
  assign n22577 = n7502 ^ n5201 ^ 1'b0 ;
  assign n22578 = ~n22576 & n22577 ;
  assign n22579 = n5316 & ~n14586 ;
  assign n22580 = ( ~n4188 & n19099 ) | ( ~n4188 & n22579 ) | ( n19099 & n22579 ) ;
  assign n22581 = n22578 | n22580 ;
  assign n22582 = n10472 ^ n2051 ^ 1'b0 ;
  assign n22583 = n17919 & n22582 ;
  assign n22584 = ( ~n2805 & n4980 ) | ( ~n2805 & n14115 ) | ( n4980 & n14115 ) ;
  assign n22585 = n10066 ^ n6283 ^ 1'b0 ;
  assign n22586 = ~n14733 & n22585 ;
  assign n22587 = n22586 ^ n22095 ^ 1'b0 ;
  assign n22588 = n12335 | n22587 ;
  assign n22589 = n1017 & ~n22588 ;
  assign n22590 = n3667 ^ n2350 ^ 1'b0 ;
  assign n22591 = n3834 ^ n483 ^ 1'b0 ;
  assign n22592 = n12785 & ~n22591 ;
  assign n22593 = n3993 & ~n22047 ;
  assign n22594 = ( n489 & ~n11563 ) | ( n489 & n12923 ) | ( ~n11563 & n12923 ) ;
  assign n22595 = ( n12173 & n22593 ) | ( n12173 & ~n22594 ) | ( n22593 & ~n22594 ) ;
  assign n22596 = n2579 | n2850 ;
  assign n22597 = n16065 & ~n22596 ;
  assign n22598 = ( n22592 & n22595 ) | ( n22592 & n22597 ) | ( n22595 & n22597 ) ;
  assign n22599 = n2556 & ~n5565 ;
  assign n22600 = n22599 ^ n1193 ^ 1'b0 ;
  assign n22601 = n10207 & n22600 ;
  assign n22602 = x41 | n6659 ;
  assign n22603 = ( ~n2073 & n9360 ) | ( ~n2073 & n22602 ) | ( n9360 & n22602 ) ;
  assign n22604 = n22603 ^ n11642 ^ 1'b0 ;
  assign n22605 = ~n10859 & n22604 ;
  assign n22606 = n14152 ^ n5545 ^ 1'b0 ;
  assign n22607 = n22605 & n22606 ;
  assign n22608 = n9387 | n13199 ;
  assign n22609 = n22608 ^ n8828 ^ 1'b0 ;
  assign n22610 = ~n9183 & n9186 ;
  assign n22611 = n2218 & n22610 ;
  assign n22612 = n22611 ^ n12927 ^ n11494 ;
  assign n22613 = n13179 & n15617 ;
  assign n22614 = n9177 ^ n996 ^ x80 ;
  assign n22615 = n4037 | n22614 ;
  assign n22616 = ( n13754 & n16864 ) | ( n13754 & n18892 ) | ( n16864 & n18892 ) ;
  assign n22617 = n22616 ^ n21565 ^ 1'b0 ;
  assign n22618 = n22617 ^ n22284 ^ n10437 ;
  assign n22619 = n14963 ^ n11048 ^ n765 ;
  assign n22620 = ( n2474 & ~n18245 ) | ( n2474 & n22619 ) | ( ~n18245 & n22619 ) ;
  assign n22621 = ( n1148 & n5036 ) | ( n1148 & ~n18778 ) | ( n5036 & ~n18778 ) ;
  assign n22622 = n14667 & ~n22621 ;
  assign n22623 = n22622 ^ n22129 ^ n8408 ;
  assign n22624 = n893 & n17902 ;
  assign n22625 = ~n9380 & n22624 ;
  assign n22626 = x93 & ~n19185 ;
  assign n22627 = ~n9808 & n22626 ;
  assign n22628 = ( ~n2163 & n5779 ) | ( ~n2163 & n8139 ) | ( n5779 & n8139 ) ;
  assign n22629 = n10901 ^ n9189 ^ n209 ;
  assign n22630 = ~n22628 & n22629 ;
  assign n22631 = ( n146 & n1129 ) | ( n146 & n1785 ) | ( n1129 & n1785 ) ;
  assign n22632 = n22631 ^ n16686 ^ n5818 ;
  assign n22633 = ~n2784 & n22632 ;
  assign n22634 = n10563 ^ n4651 ^ 1'b0 ;
  assign n22635 = n9591 & ~n22634 ;
  assign n22641 = n10564 ^ n8234 ^ n2687 ;
  assign n22640 = n11703 ^ n9110 ^ n5559 ;
  assign n22636 = n12774 ^ n7793 ^ n1577 ;
  assign n22637 = n6099 | n22636 ;
  assign n22638 = n22637 ^ n13489 ^ 1'b0 ;
  assign n22639 = n12218 | n22638 ;
  assign n22642 = n22641 ^ n22640 ^ n22639 ;
  assign n22650 = n19461 ^ n16076 ^ 1'b0 ;
  assign n22651 = n2771 & ~n22650 ;
  assign n22652 = n2867 | n12730 ;
  assign n22653 = n22651 | n22652 ;
  assign n22643 = ~n11248 & n20794 ;
  assign n22644 = n11441 & n22643 ;
  assign n22645 = n22644 ^ n2550 ^ 1'b0 ;
  assign n22646 = n20260 ^ n11053 ^ 1'b0 ;
  assign n22647 = ~n12897 & n22646 ;
  assign n22648 = n22647 ^ n3459 ^ 1'b0 ;
  assign n22649 = n22645 & ~n22648 ;
  assign n22654 = n22653 ^ n22649 ^ 1'b0 ;
  assign n22655 = n16780 ^ n10320 ^ 1'b0 ;
  assign n22656 = n5356 & ~n22655 ;
  assign n22657 = n16198 ^ n14736 ^ n6062 ;
  assign n22658 = n22657 ^ n3799 ^ 1'b0 ;
  assign n22659 = n1935 | n22658 ;
  assign n22660 = n22659 ^ n19619 ^ n18902 ;
  assign n22661 = n12774 ^ n7932 ^ n3091 ;
  assign n22662 = n22661 ^ n20310 ^ n11088 ;
  assign n22663 = n20964 ^ n18397 ^ n3735 ;
  assign n22664 = ~n10547 & n11565 ;
  assign n22665 = n22664 ^ n9536 ^ n1855 ;
  assign n22666 = n12352 ^ n6845 ^ n2604 ;
  assign n22667 = n22666 ^ n8926 ^ 1'b0 ;
  assign n22668 = n11031 | n22667 ;
  assign n22669 = n22668 ^ n14186 ^ n3107 ;
  assign n22670 = n15517 ^ n3632 ^ 1'b0 ;
  assign n22671 = ~n7836 & n22670 ;
  assign n22672 = n10913 ^ n2449 ^ n2053 ;
  assign n22673 = n3238 & ~n22672 ;
  assign n22674 = ~n20356 & n22673 ;
  assign n22675 = n6637 ^ x95 ^ 1'b0 ;
  assign n22676 = n13015 & ~n22675 ;
  assign n22677 = ~n5642 & n22676 ;
  assign n22678 = n21015 & n21689 ;
  assign n22679 = ( x11 & n5233 ) | ( x11 & n6804 ) | ( n5233 & n6804 ) ;
  assign n22680 = n4559 ^ n3146 ^ 1'b0 ;
  assign n22681 = n22679 & ~n22680 ;
  assign n22682 = n19632 ^ n5282 ^ 1'b0 ;
  assign n22683 = n6324 & n8886 ;
  assign n22684 = n22683 ^ n18161 ^ n345 ;
  assign n22685 = n9591 & n22684 ;
  assign n22686 = x15 & ~n4219 ;
  assign n22687 = n22686 ^ n2424 ^ 1'b0 ;
  assign n22688 = n22687 ^ n11633 ^ 1'b0 ;
  assign n22689 = n22098 ^ n14071 ^ n5300 ;
  assign n22690 = n22689 ^ n12415 ^ n3587 ;
  assign n22691 = n6914 | n22690 ;
  assign n22692 = n22691 ^ n21120 ^ 1'b0 ;
  assign n22693 = n8908 ^ n145 ^ 1'b0 ;
  assign n22694 = ~n20982 & n22693 ;
  assign n22695 = n10278 ^ n4072 ^ 1'b0 ;
  assign n22696 = n11662 ^ n9019 ^ 1'b0 ;
  assign n22697 = n22696 ^ n3073 ^ n677 ;
  assign n22698 = n1349 & ~n5361 ;
  assign n22699 = ~n8388 & n22698 ;
  assign n22700 = n22697 & ~n22699 ;
  assign n22701 = n21662 ^ n12298 ^ n5668 ;
  assign n22702 = n8067 ^ n656 ^ 1'b0 ;
  assign n22703 = n13919 ^ n5691 ^ n2310 ;
  assign n22705 = n9175 ^ n2059 ^ 1'b0 ;
  assign n22706 = ( ~n1448 & n6335 ) | ( ~n1448 & n22705 ) | ( n6335 & n22705 ) ;
  assign n22707 = n22706 ^ n884 ^ n764 ;
  assign n22704 = ( ~n185 & n4767 ) | ( ~n185 & n11618 ) | ( n4767 & n11618 ) ;
  assign n22708 = n22707 ^ n22704 ^ n10759 ;
  assign n22709 = n20163 ^ n9317 ^ n6819 ;
  assign n22710 = n10647 & ~n22709 ;
  assign n22711 = n1353 | n13276 ;
  assign n22712 = n18989 & ~n22711 ;
  assign n22713 = ( n2619 & ~n8703 ) | ( n2619 & n9155 ) | ( ~n8703 & n9155 ) ;
  assign n22714 = ( n5418 & ~n10856 ) | ( n5418 & n22713 ) | ( ~n10856 & n22713 ) ;
  assign n22715 = ~n11256 & n22714 ;
  assign n22716 = n22715 ^ n7634 ^ 1'b0 ;
  assign n22717 = n1346 & n2902 ;
  assign n22718 = n9484 & ~n22717 ;
  assign n22719 = n22718 ^ n15655 ^ 1'b0 ;
  assign n22720 = ( n9731 & ~n11640 ) | ( n9731 & n14403 ) | ( ~n11640 & n14403 ) ;
  assign n22721 = ~n10459 & n19564 ;
  assign n22724 = ~n319 & n3260 ;
  assign n22725 = n22724 ^ n9279 ^ n673 ;
  assign n22722 = n7114 ^ n6965 ^ 1'b0 ;
  assign n22723 = n3916 | n22722 ;
  assign n22726 = n22725 ^ n22723 ^ n992 ;
  assign n22727 = n22726 ^ n18851 ^ n9387 ;
  assign n22728 = n22727 ^ n9759 ^ n4423 ;
  assign n22729 = n11122 ^ n4587 ^ 1'b0 ;
  assign n22730 = n6005 ^ n4357 ^ 1'b0 ;
  assign n22731 = n22730 ^ n5645 ^ n512 ;
  assign n22732 = ( n16387 & ~n22729 ) | ( n16387 & n22731 ) | ( ~n22729 & n22731 ) ;
  assign n22733 = n9320 & ~n16500 ;
  assign n22734 = n22733 ^ n6619 ^ 1'b0 ;
  assign n22735 = n22734 ^ n6153 ^ n4008 ;
  assign n22736 = n19789 ^ n1617 ^ 1'b0 ;
  assign n22737 = n4016 | n22736 ;
  assign n22738 = ~n12254 & n15092 ;
  assign n22739 = n22738 ^ n2435 ^ 1'b0 ;
  assign n22740 = n6746 & n6795 ;
  assign n22741 = n20513 ^ n13250 ^ n10141 ;
  assign n22742 = n22741 ^ n17560 ^ n1737 ;
  assign n22743 = n10219 ^ n9755 ^ n9611 ;
  assign n22744 = ~n5531 & n7219 ;
  assign n22745 = n22744 ^ n13391 ^ 1'b0 ;
  assign n22746 = n22745 ^ n13253 ^ n3702 ;
  assign n22747 = n11405 ^ n3406 ^ 1'b0 ;
  assign n22748 = n235 | n8032 ;
  assign n22749 = n9900 | n22748 ;
  assign n22750 = n22749 ^ x120 ^ 1'b0 ;
  assign n22751 = ( n13451 & n22747 ) | ( n13451 & ~n22750 ) | ( n22747 & ~n22750 ) ;
  assign n22752 = n19823 ^ n7582 ^ 1'b0 ;
  assign n22753 = ( n6352 & n8796 ) | ( n6352 & n12245 ) | ( n8796 & n12245 ) ;
  assign n22754 = n13722 ^ n13313 ^ n7585 ;
  assign n22755 = n2374 & ~n20469 ;
  assign n22756 = n22755 ^ n14614 ^ n8920 ;
  assign n22757 = n8639 ^ n8372 ^ n2961 ;
  assign n22758 = ( ~n2734 & n3909 ) | ( ~n2734 & n22757 ) | ( n3909 & n22757 ) ;
  assign n22759 = n7195 ^ n3966 ^ 1'b0 ;
  assign n22760 = n21213 & ~n22759 ;
  assign n22761 = ( ~n7087 & n7657 ) | ( ~n7087 & n9286 ) | ( n7657 & n9286 ) ;
  assign n22762 = n5479 & ~n22761 ;
  assign n22763 = n22762 ^ x26 ^ 1'b0 ;
  assign n22764 = ~n9565 & n9925 ;
  assign n22765 = n2016 ^ n1263 ^ 1'b0 ;
  assign n22766 = ( ~n3387 & n17157 ) | ( ~n3387 & n22765 ) | ( n17157 & n22765 ) ;
  assign n22767 = ( n3745 & n22764 ) | ( n3745 & n22766 ) | ( n22764 & n22766 ) ;
  assign n22768 = n1465 | n13737 ;
  assign n22775 = n2742 & n18058 ;
  assign n22776 = n22775 ^ n9318 ^ 1'b0 ;
  assign n22771 = ( n5259 & n7183 ) | ( n5259 & ~n14973 ) | ( n7183 & ~n14973 ) ;
  assign n22772 = ~n747 & n22771 ;
  assign n22773 = n22772 ^ n18763 ^ n4088 ;
  assign n22774 = n22773 ^ n22621 ^ n3368 ;
  assign n22769 = n10548 | n14389 ;
  assign n22770 = n22769 ^ n18021 ^ 1'b0 ;
  assign n22777 = n22776 ^ n22774 ^ n22770 ;
  assign n22778 = n14803 ^ n14707 ^ n8936 ;
  assign n22779 = n22778 ^ n18590 ^ n16670 ;
  assign n22783 = n8173 ^ n6586 ^ 1'b0 ;
  assign n22780 = n18726 ^ n13391 ^ n12612 ;
  assign n22781 = n22780 ^ n14500 ^ 1'b0 ;
  assign n22782 = n22781 ^ n3832 ^ n933 ;
  assign n22784 = n22783 ^ n22782 ^ 1'b0 ;
  assign n22785 = n16581 | n22784 ;
  assign n22786 = n22785 ^ n11370 ^ n8827 ;
  assign n22787 = ~n1588 & n18583 ;
  assign n22788 = n21095 & n22787 ;
  assign n22789 = n20356 & ~n22788 ;
  assign n22790 = n13563 & n22789 ;
  assign n22792 = ( n3435 & n7359 ) | ( n3435 & n12087 ) | ( n7359 & n12087 ) ;
  assign n22791 = n4754 ^ n4281 ^ n4093 ;
  assign n22793 = n22792 ^ n22791 ^ n10689 ;
  assign n22794 = n20470 ^ n10252 ^ 1'b0 ;
  assign n22796 = ~n12379 & n20190 ;
  assign n22797 = ~n3150 & n22796 ;
  assign n22795 = ( ~n2413 & n6639 ) | ( ~n2413 & n14097 ) | ( n6639 & n14097 ) ;
  assign n22798 = n22797 ^ n22795 ^ n3504 ;
  assign n22799 = n5095 & ~n9656 ;
  assign n22800 = n555 & n3200 ;
  assign n22801 = n12488 | n22800 ;
  assign n22802 = n5390 & ~n22801 ;
  assign n22803 = ( n3543 & ~n9950 ) | ( n3543 & n12892 ) | ( ~n9950 & n12892 ) ;
  assign n22804 = ( n13055 & n16760 ) | ( n13055 & ~n22803 ) | ( n16760 & ~n22803 ) ;
  assign n22805 = ( n2663 & n9619 ) | ( n2663 & n11168 ) | ( n9619 & n11168 ) ;
  assign n22806 = n22805 ^ n14168 ^ n2423 ;
  assign n22807 = n10451 ^ n3807 ^ 1'b0 ;
  assign n22808 = ~n22806 & n22807 ;
  assign n22809 = ~n22804 & n22808 ;
  assign n22813 = ~n9745 & n18527 ;
  assign n22814 = n4887 & n22813 ;
  assign n22810 = ( n13460 & n15397 ) | ( n13460 & n20663 ) | ( n15397 & n20663 ) ;
  assign n22811 = n1099 | n22810 ;
  assign n22812 = n4453 & ~n22811 ;
  assign n22815 = n22814 ^ n22812 ^ n725 ;
  assign n22816 = n295 | n999 ;
  assign n22817 = ~n170 & n6290 ;
  assign n22818 = n22817 ^ n7588 ^ 1'b0 ;
  assign n22819 = ( n17158 & n22816 ) | ( n17158 & ~n22818 ) | ( n22816 & ~n22818 ) ;
  assign n22820 = ( n9031 & n11063 ) | ( n9031 & n22819 ) | ( n11063 & n22819 ) ;
  assign n22821 = n22820 ^ x53 ^ 1'b0 ;
  assign n22822 = n11916 ^ n7566 ^ n5016 ;
  assign n22823 = ( n16586 & n19115 ) | ( n16586 & n22822 ) | ( n19115 & n22822 ) ;
  assign n22824 = ~n5047 & n14793 ;
  assign n22825 = n22824 ^ n16166 ^ 1'b0 ;
  assign n22826 = n9434 ^ n2411 ^ 1'b0 ;
  assign n22827 = n12367 ^ n1794 ^ 1'b0 ;
  assign n22828 = n22827 ^ n6054 ^ n4551 ;
  assign n22829 = n22828 ^ n7871 ^ 1'b0 ;
  assign n22830 = n22826 | n22829 ;
  assign n22831 = n16230 ^ n2165 ^ 1'b0 ;
  assign n22832 = x67 & n5715 ;
  assign n22833 = n22832 ^ n3676 ^ 1'b0 ;
  assign n22834 = n22833 ^ n6108 ^ 1'b0 ;
  assign n22835 = n17435 ^ n7324 ^ n5397 ;
  assign n22836 = ( n5864 & n6829 ) | ( n5864 & n14781 ) | ( n6829 & n14781 ) ;
  assign n22837 = n21881 ^ n18450 ^ 1'b0 ;
  assign n22838 = n904 & ~n22837 ;
  assign n22839 = ( n14676 & n22836 ) | ( n14676 & ~n22838 ) | ( n22836 & ~n22838 ) ;
  assign n22840 = ~n7223 & n16820 ;
  assign n22841 = ( n10677 & n11806 ) | ( n10677 & ~n19808 ) | ( n11806 & ~n19808 ) ;
  assign n22842 = n14478 & n22841 ;
  assign n22843 = ~n4141 & n22842 ;
  assign n22844 = n22840 & ~n22843 ;
  assign n22845 = n11202 & n22844 ;
  assign n22846 = ( n3969 & n10904 ) | ( n3969 & n22845 ) | ( n10904 & n22845 ) ;
  assign n22847 = n18737 ^ n4169 ^ 1'b0 ;
  assign n22848 = ( n5962 & ~n13298 ) | ( n5962 & n16297 ) | ( ~n13298 & n16297 ) ;
  assign n22849 = n3778 & ~n10523 ;
  assign n22850 = n22849 ^ n8508 ^ 1'b0 ;
  assign n22851 = ( ~n9222 & n11167 ) | ( ~n9222 & n20371 ) | ( n11167 & n20371 ) ;
  assign n22852 = ( ~n9925 & n12239 ) | ( ~n9925 & n19040 ) | ( n12239 & n19040 ) ;
  assign n22853 = ( n5726 & ~n6891 ) | ( n5726 & n16326 ) | ( ~n6891 & n16326 ) ;
  assign n22854 = ~n547 & n1631 ;
  assign n22855 = n332 & n22854 ;
  assign n22856 = n18771 ^ n7943 ^ n3896 ;
  assign n22857 = n17137 ^ n6382 ^ 1'b0 ;
  assign n22858 = n14397 ^ n10685 ^ 1'b0 ;
  assign n22859 = n11829 & ~n22858 ;
  assign n22860 = n21510 ^ n21304 ^ 1'b0 ;
  assign n22861 = n21195 | n22860 ;
  assign n22862 = ( ~n8819 & n22859 ) | ( ~n8819 & n22861 ) | ( n22859 & n22861 ) ;
  assign n22863 = n10372 & n22862 ;
  assign n22864 = n10748 & n22863 ;
  assign n22865 = n22864 ^ n15366 ^ n10949 ;
  assign n22866 = n16794 ^ n8431 ^ 1'b0 ;
  assign n22867 = n9021 ^ n8121 ^ 1'b0 ;
  assign n22868 = ~n9650 & n22867 ;
  assign n22869 = ~n12005 & n16397 ;
  assign n22870 = ( n10125 & ~n17320 ) | ( n10125 & n19564 ) | ( ~n17320 & n19564 ) ;
  assign n22871 = ( n16904 & n22869 ) | ( n16904 & n22870 ) | ( n22869 & n22870 ) ;
  assign n22872 = ( ~n12333 & n22868 ) | ( ~n12333 & n22871 ) | ( n22868 & n22871 ) ;
  assign n22873 = ( ~n1097 & n10052 ) | ( ~n1097 & n22872 ) | ( n10052 & n22872 ) ;
  assign n22874 = n9847 & n13270 ;
  assign n22875 = n8020 | n8560 ;
  assign n22876 = n15828 & ~n22875 ;
  assign n22877 = n22704 ^ n6793 ^ n6168 ;
  assign n22878 = ( ~n14290 & n19500 ) | ( ~n14290 & n22877 ) | ( n19500 & n22877 ) ;
  assign n22879 = ( n4247 & n9041 ) | ( n4247 & n17250 ) | ( n9041 & n17250 ) ;
  assign n22880 = n11268 ^ n2850 ^ 1'b0 ;
  assign n22881 = ~n22879 & n22880 ;
  assign n22882 = n7913 & n22881 ;
  assign n22883 = n9217 ^ n2103 ^ 1'b0 ;
  assign n22884 = n22883 ^ n15126 ^ 1'b0 ;
  assign n22885 = ( n8656 & n19650 ) | ( n8656 & ~n20773 ) | ( n19650 & ~n20773 ) ;
  assign n22886 = ~n3926 & n22885 ;
  assign n22887 = n6046 & n22886 ;
  assign n22888 = n6674 ^ n4486 ^ n4324 ;
  assign n22889 = n22888 ^ n2511 ^ 1'b0 ;
  assign n22891 = n17359 ^ n16238 ^ 1'b0 ;
  assign n22890 = ~n9748 & n14096 ;
  assign n22892 = n22891 ^ n22890 ^ n14806 ;
  assign n22893 = n10942 & n13393 ;
  assign n22894 = ( ~n16793 & n18161 ) | ( ~n16793 & n22893 ) | ( n18161 & n22893 ) ;
  assign n22895 = n7502 ^ n1612 ^ 1'b0 ;
  assign n22898 = n6794 ^ n3521 ^ n589 ;
  assign n22899 = n22898 ^ n8695 ^ 1'b0 ;
  assign n22896 = ~n7169 & n17314 ;
  assign n22897 = ~n2842 & n22896 ;
  assign n22900 = n22899 ^ n22897 ^ n20093 ;
  assign n22904 = n8677 ^ n2535 ^ n639 ;
  assign n22905 = ( n2897 & n16393 ) | ( n2897 & ~n22904 ) | ( n16393 & ~n22904 ) ;
  assign n22902 = ( n298 & ~n7046 ) | ( n298 & n13736 ) | ( ~n7046 & n13736 ) ;
  assign n22901 = n4515 & n16740 ;
  assign n22903 = n22902 ^ n22901 ^ 1'b0 ;
  assign n22906 = n22905 ^ n22903 ^ 1'b0 ;
  assign n22907 = ( ~n2237 & n9695 ) | ( ~n2237 & n15374 ) | ( n9695 & n15374 ) ;
  assign n22908 = n9989 & n22907 ;
  assign n22909 = n17558 & n22908 ;
  assign n22910 = n22909 ^ n19518 ^ n1093 ;
  assign n22911 = ( n2951 & ~n7909 ) | ( n2951 & n9966 ) | ( ~n7909 & n9966 ) ;
  assign n22912 = ( n8494 & n9595 ) | ( n8494 & ~n22911 ) | ( n9595 & ~n22911 ) ;
  assign n22913 = n1899 | n14396 ;
  assign n22914 = n1313 & ~n22913 ;
  assign n22915 = n13023 | n22914 ;
  assign n22916 = n4723 & ~n22915 ;
  assign n22918 = n5024 ^ n1657 ^ 1'b0 ;
  assign n22917 = ~n1871 & n16375 ;
  assign n22919 = n22918 ^ n22917 ^ 1'b0 ;
  assign n22920 = ( n163 & n14950 ) | ( n163 & ~n22919 ) | ( n14950 & ~n22919 ) ;
  assign n22921 = n16025 ^ n11269 ^ 1'b0 ;
  assign n22922 = ( n6546 & n18161 ) | ( n6546 & n22921 ) | ( n18161 & n22921 ) ;
  assign n22923 = n8825 | n9535 ;
  assign n22924 = n14893 & ~n22923 ;
  assign n22925 = n11326 | n22924 ;
  assign n22926 = ( ~n12015 & n17763 ) | ( ~n12015 & n20663 ) | ( n17763 & n20663 ) ;
  assign n22927 = n22926 ^ n19035 ^ n18716 ;
  assign n22928 = n22927 ^ n11025 ^ 1'b0 ;
  assign n22929 = ~n1025 & n3670 ;
  assign n22930 = ~n3410 & n5720 ;
  assign n22931 = n22930 ^ n22192 ^ 1'b0 ;
  assign n22932 = n4383 | n22931 ;
  assign n22933 = n1885 | n16253 ;
  assign n22934 = n22933 ^ n8151 ^ 1'b0 ;
  assign n22935 = ( n16091 & ~n20737 ) | ( n16091 & n22934 ) | ( ~n20737 & n22934 ) ;
  assign n22936 = n18385 & ~n22935 ;
  assign n22937 = n22936 ^ n3473 ^ 1'b0 ;
  assign n22938 = n4540 | n22800 ;
  assign n22939 = n22938 ^ n730 ^ 1'b0 ;
  assign n22940 = ( n4707 & n6235 ) | ( n4707 & n18112 ) | ( n6235 & n18112 ) ;
  assign n22941 = n1457 | n5071 ;
  assign n22942 = n22941 ^ n9978 ^ 1'b0 ;
  assign n22943 = ( n2185 & n22940 ) | ( n2185 & ~n22942 ) | ( n22940 & ~n22942 ) ;
  assign n22944 = ~n7836 & n19728 ;
  assign n22945 = ( n1408 & n6265 ) | ( n1408 & n7427 ) | ( n6265 & n7427 ) ;
  assign n22946 = n12523 & n16360 ;
  assign n22947 = n18778 ^ n7454 ^ 1'b0 ;
  assign n22948 = n22947 ^ n22644 ^ 1'b0 ;
  assign n22949 = n7092 & ~n22948 ;
  assign n22950 = n18647 ^ n15903 ^ 1'b0 ;
  assign n22951 = n20279 ^ n19910 ^ n5374 ;
  assign n22952 = n22951 ^ n5345 ^ n1292 ;
  assign n22953 = ( n4376 & ~n8054 ) | ( n4376 & n12142 ) | ( ~n8054 & n12142 ) ;
  assign n22954 = n13518 ^ n7151 ^ n4706 ;
  assign n22955 = n2259 ^ x92 ^ 1'b0 ;
  assign n22956 = n22954 & n22955 ;
  assign n22957 = ~n4588 & n8869 ;
  assign n22958 = ( n14759 & ~n18190 ) | ( n14759 & n22957 ) | ( ~n18190 & n22957 ) ;
  assign n22959 = n13801 | n22958 ;
  assign n22960 = n22956 | n22959 ;
  assign n22961 = ( ~n22086 & n22953 ) | ( ~n22086 & n22960 ) | ( n22953 & n22960 ) ;
  assign n22962 = n16950 ^ n13708 ^ n3992 ;
  assign n22963 = n22224 ^ n9554 ^ n2490 ;
  assign n22964 = ( n13878 & n22730 ) | ( n13878 & ~n22963 ) | ( n22730 & ~n22963 ) ;
  assign n22965 = n5139 ^ n4853 ^ 1'b0 ;
  assign n22966 = n9562 & n22965 ;
  assign n22967 = n2482 & ~n11778 ;
  assign n22968 = n3591 & n22967 ;
  assign n22969 = n1922 & ~n22968 ;
  assign n22970 = n22969 ^ n4722 ^ 1'b0 ;
  assign n22972 = n8193 ^ n1197 ^ 1'b0 ;
  assign n22973 = n22972 ^ n9245 ^ n4568 ;
  assign n22971 = n12273 ^ n9159 ^ n4120 ;
  assign n22974 = n22973 ^ n22971 ^ n8958 ;
  assign n22975 = ( n6920 & ~n8118 ) | ( n6920 & n14733 ) | ( ~n8118 & n14733 ) ;
  assign n22976 = n17120 ^ n9666 ^ 1'b0 ;
  assign n22977 = n22975 & ~n22976 ;
  assign n22978 = n22977 ^ n3750 ^ n181 ;
  assign n22979 = n22978 ^ n20253 ^ n8024 ;
  assign n22980 = n9682 ^ n1205 ^ 1'b0 ;
  assign n22981 = n1915 & ~n22980 ;
  assign n22982 = n2475 ^ n2179 ^ 1'b0 ;
  assign n22985 = ( n1203 & ~n1984 ) | ( n1203 & n6161 ) | ( ~n1984 & n6161 ) ;
  assign n22983 = n1875 & ~n16733 ;
  assign n22984 = n22983 ^ n11677 ^ 1'b0 ;
  assign n22986 = n22985 ^ n22984 ^ 1'b0 ;
  assign n22987 = n3550 ^ n900 ^ 1'b0 ;
  assign n22988 = ( n4311 & n18252 ) | ( n4311 & n22987 ) | ( n18252 & n22987 ) ;
  assign n22989 = ( n1551 & n2805 ) | ( n1551 & ~n16525 ) | ( n2805 & ~n16525 ) ;
  assign n22990 = n9654 ^ n7071 ^ 1'b0 ;
  assign n22991 = ( n6155 & n10015 ) | ( n6155 & ~n22990 ) | ( n10015 & ~n22990 ) ;
  assign n22994 = n4674 | n4739 ;
  assign n22995 = n22994 ^ n9900 ^ 1'b0 ;
  assign n22992 = n3002 & ~n8554 ;
  assign n22993 = ~n5939 & n22992 ;
  assign n22996 = n22995 ^ n22993 ^ n1587 ;
  assign n22997 = n6392 ^ n4019 ^ n3173 ;
  assign n22998 = ( ~n10079 & n21143 ) | ( ~n10079 & n22997 ) | ( n21143 & n22997 ) ;
  assign n22999 = ( n4594 & ~n8644 ) | ( n4594 & n22998 ) | ( ~n8644 & n22998 ) ;
  assign n23000 = n14706 ^ n8355 ^ 1'b0 ;
  assign n23001 = n15391 & ~n23000 ;
  assign n23002 = n2151 | n15338 ;
  assign n23003 = n23002 ^ n4411 ^ 1'b0 ;
  assign n23004 = n23003 ^ n18706 ^ n16914 ;
  assign n23005 = n13816 & ~n18961 ;
  assign n23006 = n6768 & n23005 ;
  assign n23007 = n3126 & ~n12241 ;
  assign n23008 = n23007 ^ n5896 ^ 1'b0 ;
  assign n23009 = n8961 | n16201 ;
  assign n23010 = ( n12586 & ~n21201 ) | ( n12586 & n21278 ) | ( ~n21201 & n21278 ) ;
  assign n23011 = n5070 | n18736 ;
  assign n23012 = n23011 ^ n14262 ^ 1'b0 ;
  assign n23013 = n22833 ^ n13255 ^ n12762 ;
  assign n23014 = n14206 & ~n23013 ;
  assign n23015 = n23014 ^ n7644 ^ n7141 ;
  assign n23016 = n6768 & ~n23015 ;
  assign n23017 = n1964 & ~n9738 ;
  assign n23018 = n19489 & n23017 ;
  assign n23019 = n6837 | n18696 ;
  assign n23020 = n13704 ^ n469 ^ x107 ;
  assign n23021 = n1718 ^ n338 ^ 1'b0 ;
  assign n23022 = n23021 ^ n12816 ^ n7741 ;
  assign n23023 = n5741 & ~n19992 ;
  assign n23024 = n7968 | n22287 ;
  assign n23026 = n8601 ^ n8235 ^ 1'b0 ;
  assign n23025 = n9607 & n16078 ;
  assign n23027 = n23026 ^ n23025 ^ 1'b0 ;
  assign n23028 = n23027 ^ n2317 ^ 1'b0 ;
  assign n23029 = n10466 & n23028 ;
  assign n23030 = n22124 ^ n5429 ^ 1'b0 ;
  assign n23031 = ( ~n2185 & n18064 ) | ( ~n2185 & n18660 ) | ( n18064 & n18660 ) ;
  assign n23032 = ( n11062 & ~n23030 ) | ( n11062 & n23031 ) | ( ~n23030 & n23031 ) ;
  assign n23033 = n11315 ^ n4461 ^ n2338 ;
  assign n23034 = n23033 ^ n8191 ^ 1'b0 ;
  assign n23035 = ( ~n8918 & n11221 ) | ( ~n8918 & n16904 ) | ( n11221 & n16904 ) ;
  assign n23036 = ( ~n3212 & n7774 ) | ( ~n3212 & n10409 ) | ( n7774 & n10409 ) ;
  assign n23038 = n5048 ^ n2959 ^ 1'b0 ;
  assign n23039 = ~n10274 & n23038 ;
  assign n23040 = n6079 & n23039 ;
  assign n23041 = n19471 ^ n16992 ^ 1'b0 ;
  assign n23042 = n3468 & ~n23041 ;
  assign n23043 = n23040 & ~n23042 ;
  assign n23037 = ( x101 & n13116 ) | ( x101 & ~n18522 ) | ( n13116 & ~n18522 ) ;
  assign n23044 = n23043 ^ n23037 ^ n4694 ;
  assign n23045 = n22692 ^ n9287 ^ 1'b0 ;
  assign n23046 = ( ~n1738 & n11534 ) | ( ~n1738 & n14226 ) | ( n11534 & n14226 ) ;
  assign n23047 = n12225 ^ n5002 ^ 1'b0 ;
  assign n23048 = n11472 & n23047 ;
  assign n23049 = n20999 & n23048 ;
  assign n23050 = n23049 ^ n7542 ^ 1'b0 ;
  assign n23051 = n2747 & ~n5636 ;
  assign n23052 = n7450 & n23051 ;
  assign n23053 = n23052 ^ n5310 ^ n404 ;
  assign n23054 = n1529 & ~n18503 ;
  assign n23055 = ~n23053 & n23054 ;
  assign n23056 = ( ~n18841 & n23050 ) | ( ~n18841 & n23055 ) | ( n23050 & n23055 ) ;
  assign n23057 = n12637 | n17336 ;
  assign n23058 = n18709 ^ n6682 ^ 1'b0 ;
  assign n23059 = n705 & ~n15010 ;
  assign n23060 = n23059 ^ n4003 ^ 1'b0 ;
  assign n23061 = ~n2154 & n4815 ;
  assign n23062 = n23061 ^ n22930 ^ 1'b0 ;
  assign n23063 = n3491 | n15125 ;
  assign n23064 = n23063 ^ n7789 ^ 1'b0 ;
  assign n23065 = n13338 | n22123 ;
  assign n23066 = n23065 ^ n17094 ^ 1'b0 ;
  assign n23067 = n12272 | n12305 ;
  assign n23068 = n5379 | n23067 ;
  assign n23069 = n23068 ^ n16808 ^ 1'b0 ;
  assign n23070 = n23066 | n23069 ;
  assign n23071 = ( ~n8177 & n19620 ) | ( ~n8177 & n23070 ) | ( n19620 & n23070 ) ;
  assign n23072 = n21181 ^ n20536 ^ n11276 ;
  assign n23073 = n23072 ^ n12486 ^ n8129 ;
  assign n23074 = ~n2324 & n21443 ;
  assign n23075 = ( n4393 & n14271 ) | ( n4393 & ~n23074 ) | ( n14271 & ~n23074 ) ;
  assign n23076 = n9323 ^ x108 ^ 1'b0 ;
  assign n23077 = ( ~n8240 & n10640 ) | ( ~n8240 & n23076 ) | ( n10640 & n23076 ) ;
  assign n23078 = ~n312 & n8778 ;
  assign n23079 = n23078 ^ n3712 ^ 1'b0 ;
  assign n23080 = n23077 | n23079 ;
  assign n23081 = n14705 ^ n13414 ^ n12684 ;
  assign n23082 = n22972 ^ n3716 ^ n3344 ;
  assign n23083 = n23082 ^ n7482 ^ 1'b0 ;
  assign n23084 = n17574 & ~n23083 ;
  assign n23085 = n2399 & n18033 ;
  assign n23086 = ( n20119 & ~n20583 ) | ( n20119 & n23085 ) | ( ~n20583 & n23085 ) ;
  assign n23091 = x104 | n3628 ;
  assign n23092 = n23091 ^ n566 ^ 1'b0 ;
  assign n23087 = n6857 ^ x13 ^ 1'b0 ;
  assign n23088 = ( n6780 & n8290 ) | ( n6780 & ~n23087 ) | ( n8290 & ~n23087 ) ;
  assign n23089 = n23088 ^ n5031 ^ 1'b0 ;
  assign n23090 = ~n13738 & n23089 ;
  assign n23093 = n23092 ^ n23090 ^ n13961 ;
  assign n23094 = x5 | n7912 ;
  assign n23095 = n11432 & ~n22083 ;
  assign n23096 = n23095 ^ n764 ^ 1'b0 ;
  assign n23097 = n6607 & n14220 ;
  assign n23098 = n23097 ^ n1968 ^ 1'b0 ;
  assign n23099 = n11787 ^ n2279 ^ x44 ;
  assign n23100 = n23099 ^ n3204 ^ 1'b0 ;
  assign n23101 = n18664 & n23100 ;
  assign n23102 = n14563 ^ n464 ^ 1'b0 ;
  assign n23105 = ( ~n672 & n894 ) | ( ~n672 & n6558 ) | ( n894 & n6558 ) ;
  assign n23106 = n23105 ^ n9371 ^ n1583 ;
  assign n23103 = n3648 & n10942 ;
  assign n23104 = n988 & n23103 ;
  assign n23107 = n23106 ^ n23104 ^ 1'b0 ;
  assign n23108 = n17157 ^ n9003 ^ n1859 ;
  assign n23109 = n23108 ^ n410 ^ 1'b0 ;
  assign n23110 = ~n11475 & n23109 ;
  assign n23111 = ~n5913 & n23110 ;
  assign n23112 = n23111 ^ n22211 ^ n13816 ;
  assign n23113 = ~n3067 & n4859 ;
  assign n23114 = ~n19476 & n23113 ;
  assign n23115 = ~n2494 & n3830 ;
  assign n23116 = n23115 ^ n17187 ^ 1'b0 ;
  assign n23117 = n542 & n23116 ;
  assign n23118 = n23117 ^ n19146 ^ 1'b0 ;
  assign n23119 = n4039 & n10896 ;
  assign n23120 = n13917 ^ n3042 ^ 1'b0 ;
  assign n23121 = n23120 ^ n7343 ^ n1856 ;
  assign n23122 = ( n616 & n6818 ) | ( n616 & n19254 ) | ( n6818 & n19254 ) ;
  assign n23123 = n9925 ^ n8633 ^ n3647 ;
  assign n23124 = n18864 ^ n916 ^ 1'b0 ;
  assign n23125 = n15314 | n23124 ;
  assign n23126 = n6595 ^ n3366 ^ n1068 ;
  assign n23127 = n23126 ^ n4088 ^ 1'b0 ;
  assign n23128 = n23127 ^ n16084 ^ n14050 ;
  assign n23129 = n17375 ^ n5637 ^ 1'b0 ;
  assign n23130 = n23128 & ~n23129 ;
  assign n23131 = n16384 ^ n14411 ^ 1'b0 ;
  assign n23132 = n23130 & ~n23131 ;
  assign n23133 = n10238 & ~n14347 ;
  assign n23134 = ~n15816 & n23133 ;
  assign n23135 = ~n4092 & n14966 ;
  assign n23136 = ( n7381 & n10547 ) | ( n7381 & ~n15850 ) | ( n10547 & ~n15850 ) ;
  assign n23137 = n6427 ^ n3733 ^ 1'b0 ;
  assign n23138 = ~n988 & n1260 ;
  assign n23139 = ( n1771 & n21196 ) | ( n1771 & n23138 ) | ( n21196 & n23138 ) ;
  assign n23140 = ( n17578 & n23137 ) | ( n17578 & ~n23139 ) | ( n23137 & ~n23139 ) ;
  assign n23141 = ( ~n3806 & n17221 ) | ( ~n3806 & n23140 ) | ( n17221 & n23140 ) ;
  assign n23142 = ( n11583 & n14159 ) | ( n11583 & ~n21198 ) | ( n14159 & ~n21198 ) ;
  assign n23143 = ( n1507 & n6471 ) | ( n1507 & n11676 ) | ( n6471 & n11676 ) ;
  assign n23144 = ~n3976 & n23143 ;
  assign n23145 = n23144 ^ n4367 ^ 1'b0 ;
  assign n23146 = n23142 & ~n23145 ;
  assign n23147 = n7879 ^ n3832 ^ 1'b0 ;
  assign n23148 = n6436 | n23147 ;
  assign n23149 = n12486 ^ n1994 ^ 1'b0 ;
  assign n23150 = ~n23148 & n23149 ;
  assign n23151 = n4472 & ~n15028 ;
  assign n23152 = n23151 ^ n5619 ^ 1'b0 ;
  assign n23153 = n18916 & n23152 ;
  assign n23154 = n23153 ^ n9819 ^ 1'b0 ;
  assign n23155 = n16506 ^ n272 ^ 1'b0 ;
  assign n23156 = ( ~n9028 & n15207 ) | ( ~n9028 & n23155 ) | ( n15207 & n23155 ) ;
  assign n23157 = n17477 ^ n14325 ^ n1329 ;
  assign n23158 = n872 & n9580 ;
  assign n23159 = n2824 | n21929 ;
  assign n23160 = n17876 & ~n23159 ;
  assign n23161 = n5700 | n19129 ;
  assign n23162 = n22532 & ~n23161 ;
  assign n23163 = n15352 ^ n8426 ^ n8177 ;
  assign n23164 = n7018 & n7087 ;
  assign n23165 = n19708 ^ n11978 ^ n5644 ;
  assign n23166 = n23165 ^ n20235 ^ n201 ;
  assign n23167 = n2576 & n19010 ;
  assign n23168 = n9834 | n17142 ;
  assign n23169 = n23168 ^ n3840 ^ 1'b0 ;
  assign n23170 = n1987 | n19168 ;
  assign n23171 = n23170 ^ n21636 ^ 1'b0 ;
  assign n23172 = ( n573 & n23169 ) | ( n573 & n23171 ) | ( n23169 & n23171 ) ;
  assign n23173 = n14364 ^ n8101 ^ n1953 ;
  assign n23174 = ( ~n9681 & n11266 ) | ( ~n9681 & n23173 ) | ( n11266 & n23173 ) ;
  assign n23175 = n23174 ^ n19601 ^ n1024 ;
  assign n23176 = n1599 | n3254 ;
  assign n23177 = n14793 | n23176 ;
  assign n23178 = ~n7051 & n23177 ;
  assign n23179 = n4486 & n23178 ;
  assign n23180 = x85 & n11648 ;
  assign n23181 = n6585 & n23180 ;
  assign n23182 = n4067 ^ n2583 ^ 1'b0 ;
  assign n23183 = n23181 | n23182 ;
  assign n23184 = ( n20184 & n23179 ) | ( n20184 & n23183 ) | ( n23179 & n23183 ) ;
  assign n23185 = n12668 ^ n12139 ^ 1'b0 ;
  assign n23186 = n8870 | n23185 ;
  assign n23187 = n23186 ^ n19717 ^ n13164 ;
  assign n23188 = n7244 & ~n14736 ;
  assign n23189 = n23188 ^ n9358 ^ 1'b0 ;
  assign n23190 = n23189 ^ n10780 ^ n4667 ;
  assign n23191 = n16254 ^ n11962 ^ 1'b0 ;
  assign n23192 = ( ~n1548 & n1926 ) | ( ~n1548 & n1982 ) | ( n1926 & n1982 ) ;
  assign n23193 = n13700 ^ n8334 ^ 1'b0 ;
  assign n23194 = n23192 & ~n23193 ;
  assign n23195 = n5554 | n6895 ;
  assign n23196 = n7957 & ~n23195 ;
  assign n23197 = n21496 ^ n7363 ^ 1'b0 ;
  assign n23198 = n10532 ^ n8708 ^ n343 ;
  assign n23199 = ( n4718 & n8234 ) | ( n4718 & n23198 ) | ( n8234 & n23198 ) ;
  assign n23200 = n23199 ^ n20677 ^ n12663 ;
  assign n23201 = ~n18105 & n23200 ;
  assign n23202 = ( n2241 & n3432 ) | ( n2241 & ~n21839 ) | ( n3432 & ~n21839 ) ;
  assign n23203 = ( n3253 & n5941 ) | ( n3253 & ~n20664 ) | ( n5941 & ~n20664 ) ;
  assign n23204 = n9575 ^ n8767 ^ n6763 ;
  assign n23205 = ~n5756 & n23204 ;
  assign n23206 = n17091 & n23205 ;
  assign n23207 = n23206 ^ n20196 ^ n2004 ;
  assign n23208 = n3134 ^ n285 ^ 1'b0 ;
  assign n23209 = n12440 | n23208 ;
  assign n23210 = n19266 ^ n8024 ^ n4305 ;
  assign n23211 = ~n23209 & n23210 ;
  assign n23212 = n5706 ^ x78 ^ 1'b0 ;
  assign n23213 = n8255 & n23212 ;
  assign n23214 = n23213 ^ n5542 ^ 1'b0 ;
  assign n23215 = n18375 & n23214 ;
  assign n23216 = n6994 & n23215 ;
  assign n23217 = n7230 | n23216 ;
  assign n23218 = n23217 ^ n1567 ^ 1'b0 ;
  assign n23219 = ( x0 & ~n23211 ) | ( x0 & n23218 ) | ( ~n23211 & n23218 ) ;
  assign n23220 = n23027 ^ n20364 ^ 1'b0 ;
  assign n23224 = ( n3716 & n4349 ) | ( n3716 & ~n4460 ) | ( n4349 & ~n4460 ) ;
  assign n23221 = n13398 ^ n7888 ^ n4614 ;
  assign n23222 = n23221 ^ n2534 ^ 1'b0 ;
  assign n23223 = n14385 & ~n23222 ;
  assign n23225 = n23224 ^ n23223 ^ 1'b0 ;
  assign n23226 = n6185 & n11044 ;
  assign n23227 = n23226 ^ n11273 ^ 1'b0 ;
  assign n23228 = n23227 ^ n22105 ^ n14805 ;
  assign n23229 = n8370 ^ n7257 ^ 1'b0 ;
  assign n23230 = ~n11133 & n12248 ;
  assign n23231 = n21195 ^ n8592 ^ n8014 ;
  assign n23232 = n23230 | n23231 ;
  assign n23233 = n2648 & n7660 ;
  assign n23234 = n14909 ^ n7431 ^ 1'b0 ;
  assign n23235 = n23234 ^ n7724 ^ 1'b0 ;
  assign n23236 = n13667 & n23235 ;
  assign n23237 = n23233 & n23236 ;
  assign n23238 = n23237 ^ n1823 ^ 1'b0 ;
  assign n23239 = n6919 ^ n3175 ^ n2171 ;
  assign n23241 = n9422 ^ n1448 ^ 1'b0 ;
  assign n23242 = n7820 & n23241 ;
  assign n23243 = n23242 ^ n7234 ^ 1'b0 ;
  assign n23244 = n4904 & ~n23243 ;
  assign n23240 = n17615 ^ n7748 ^ n1084 ;
  assign n23245 = n23244 ^ n23240 ^ n16103 ;
  assign n23246 = n23239 & n23245 ;
  assign n23247 = n6981 ^ n5338 ^ 1'b0 ;
  assign n23248 = ( n483 & ~n7551 ) | ( n483 & n11479 ) | ( ~n7551 & n11479 ) ;
  assign n23249 = n23248 ^ n9840 ^ n7601 ;
  assign n23250 = ( n8173 & ~n9667 ) | ( n8173 & n20937 ) | ( ~n9667 & n20937 ) ;
  assign n23251 = n23249 & n23250 ;
  assign n23252 = ( n1269 & n10081 ) | ( n1269 & ~n22528 ) | ( n10081 & ~n22528 ) ;
  assign n23253 = n23252 ^ n16209 ^ n8470 ;
  assign n23254 = n14743 ^ n5380 ^ 1'b0 ;
  assign n23255 = n1208 & ~n23254 ;
  assign n23256 = ( n420 & n6046 ) | ( n420 & n21311 ) | ( n6046 & n21311 ) ;
  assign n23257 = n17001 ^ n5525 ^ 1'b0 ;
  assign n23258 = ( n3164 & n13093 ) | ( n3164 & n23257 ) | ( n13093 & n23257 ) ;
  assign n23259 = n21982 ^ n15900 ^ n14683 ;
  assign n23260 = n3723 | n8202 ;
  assign n23261 = n23260 ^ n3507 ^ 1'b0 ;
  assign n23262 = n23261 ^ n8386 ^ 1'b0 ;
  assign n23263 = ~n23259 & n23262 ;
  assign n23264 = ( n2053 & n3764 ) | ( n2053 & n5562 ) | ( n3764 & n5562 ) ;
  assign n23265 = n12697 | n23264 ;
  assign n23266 = ~n11471 & n11833 ;
  assign n23267 = ~n23265 & n23266 ;
  assign n23268 = ~n4731 & n17342 ;
  assign n23269 = n305 | n4036 ;
  assign n23270 = n23269 ^ n13420 ^ n12474 ;
  assign n23271 = n10516 ^ n7850 ^ n3198 ;
  assign n23272 = n14764 & ~n23271 ;
  assign n23273 = ~n20477 & n23272 ;
  assign n23274 = ( n9944 & n12387 ) | ( n9944 & ~n23273 ) | ( n12387 & ~n23273 ) ;
  assign n23275 = n2904 & ~n13208 ;
  assign n23276 = n9249 | n23275 ;
  assign n23277 = n16450 & ~n23276 ;
  assign n23278 = n2964 | n23277 ;
  assign n23279 = n21873 ^ n20219 ^ n4169 ;
  assign n23280 = n10408 ^ n3024 ^ 1'b0 ;
  assign n23281 = n23280 ^ n8118 ^ n3955 ;
  assign n23282 = n21017 & ~n23281 ;
  assign n23283 = ~n16552 & n23282 ;
  assign n23284 = n986 | n5388 ;
  assign n23285 = ( n8942 & ~n9204 ) | ( n8942 & n23284 ) | ( ~n9204 & n23284 ) ;
  assign n23286 = n23285 ^ n4438 ^ n3555 ;
  assign n23287 = n18450 ^ n10780 ^ n5669 ;
  assign n23288 = n13053 ^ n3284 ^ 1'b0 ;
  assign n23289 = n3126 & n11200 ;
  assign n23290 = n3726 & ~n23289 ;
  assign n23291 = n23290 ^ n18887 ^ 1'b0 ;
  assign n23292 = ( n964 & n4403 ) | ( n964 & ~n12860 ) | ( n4403 & ~n12860 ) ;
  assign n23293 = n23292 ^ n3287 ^ 1'b0 ;
  assign n23294 = n7789 & ~n23293 ;
  assign n23295 = ~n2216 & n10534 ;
  assign n23296 = ~n10901 & n23295 ;
  assign n23297 = n17965 & n23296 ;
  assign n23298 = n17396 ^ n9540 ^ n2386 ;
  assign n23299 = n17075 ^ n9365 ^ n8072 ;
  assign n23300 = ~n2192 & n23299 ;
  assign n23305 = n23126 ^ n11690 ^ 1'b0 ;
  assign n23301 = ( n2546 & n5006 ) | ( n2546 & ~n19572 ) | ( n5006 & ~n19572 ) ;
  assign n23302 = n20360 ^ n12887 ^ n10892 ;
  assign n23303 = n2427 & ~n23302 ;
  assign n23304 = n23301 & n23303 ;
  assign n23306 = n23305 ^ n23304 ^ n22518 ;
  assign n23307 = ~n725 & n1382 ;
  assign n23308 = n536 & n23307 ;
  assign n23309 = n14144 & n15144 ;
  assign n23310 = n15417 ^ n14206 ^ n3596 ;
  assign n23311 = n18513 & n23310 ;
  assign n23312 = n10965 ^ n1959 ^ 1'b0 ;
  assign n23313 = n2867 | n23312 ;
  assign n23314 = n23313 ^ n16382 ^ n9060 ;
  assign n23315 = n10016 & ~n23314 ;
  assign n23316 = n7085 ^ x127 ^ 1'b0 ;
  assign n23317 = ~n19394 & n23316 ;
  assign n23318 = n1832 & n19601 ;
  assign n23319 = n23318 ^ n9632 ^ 1'b0 ;
  assign n23320 = n19848 ^ n4127 ^ n1212 ;
  assign n23321 = ( n171 & n4272 ) | ( n171 & ~n23320 ) | ( n4272 & ~n23320 ) ;
  assign n23322 = ~n5139 & n8885 ;
  assign n23323 = ~n7739 & n23322 ;
  assign n23324 = n23323 ^ n4940 ^ n894 ;
  assign n23325 = n11062 ^ n7436 ^ 1'b0 ;
  assign n23326 = n13851 ^ n2489 ^ n760 ;
  assign n23327 = ( n2383 & ~n5387 ) | ( n2383 & n23326 ) | ( ~n5387 & n23326 ) ;
  assign n23328 = n17687 ^ n9753 ^ n3582 ;
  assign n23329 = n21935 | n23328 ;
  assign n23330 = ~n11899 & n23329 ;
  assign n23331 = n1046 & ~n14019 ;
  assign n23332 = ~n3565 & n23331 ;
  assign n23333 = n12351 ^ n8281 ^ x48 ;
  assign n23334 = n3529 & ~n7205 ;
  assign n23335 = n23334 ^ n3908 ^ 1'b0 ;
  assign n23336 = n23335 ^ n21222 ^ n12804 ;
  assign n23337 = n19521 ^ n9204 ^ x101 ;
  assign n23338 = ~n2815 & n4706 ;
  assign n23339 = n23338 ^ n351 ^ 1'b0 ;
  assign n23340 = ( ~n6223 & n11880 ) | ( ~n6223 & n23339 ) | ( n11880 & n23339 ) ;
  assign n23341 = n5576 & n16840 ;
  assign n23342 = n21344 & n23341 ;
  assign n23343 = ~n8979 & n11531 ;
  assign n23344 = n23343 ^ n18369 ^ 1'b0 ;
  assign n23345 = n17961 ^ n9202 ^ 1'b0 ;
  assign n23346 = ~n23344 & n23345 ;
  assign n23347 = ~n11810 & n17627 ;
  assign n23348 = ~n2176 & n23347 ;
  assign n23349 = n7614 | n17155 ;
  assign n23350 = n10228 & ~n23349 ;
  assign n23351 = ( n16864 & n17557 ) | ( n16864 & ~n23350 ) | ( n17557 & ~n23350 ) ;
  assign n23352 = ( n10324 & n21170 ) | ( n10324 & ~n21611 ) | ( n21170 & ~n21611 ) ;
  assign n23353 = n7920 ^ n3145 ^ 1'b0 ;
  assign n23354 = n3216 & ~n9572 ;
  assign n23355 = n23354 ^ n1358 ^ 1'b0 ;
  assign n23356 = n17389 & n23355 ;
  assign n23357 = n23356 ^ n11435 ^ 1'b0 ;
  assign n23358 = ( n1332 & n3351 ) | ( n1332 & ~n4233 ) | ( n3351 & ~n4233 ) ;
  assign n23359 = n18756 ^ n4863 ^ 1'b0 ;
  assign n23360 = n23358 & n23359 ;
  assign n23361 = ( n555 & ~n10709 ) | ( n555 & n12654 ) | ( ~n10709 & n12654 ) ;
  assign n23362 = n7119 | n19686 ;
  assign n23363 = ( ~n10564 & n14250 ) | ( ~n10564 & n23362 ) | ( n14250 & n23362 ) ;
  assign n23364 = n8434 & n10778 ;
  assign n23365 = ( n7256 & n10451 ) | ( n7256 & ~n23364 ) | ( n10451 & ~n23364 ) ;
  assign n23366 = n9004 ^ n3758 ^ n2307 ;
  assign n23367 = n17963 & ~n21510 ;
  assign n23368 = ~n23366 & n23367 ;
  assign n23369 = n7340 & n14357 ;
  assign n23370 = n23369 ^ n8094 ^ 1'b0 ;
  assign n23371 = n8642 & ~n22212 ;
  assign n23372 = n23371 ^ n1668 ^ 1'b0 ;
  assign n23373 = n3486 | n7259 ;
  assign n23374 = n5462 | n17354 ;
  assign n23375 = n3482 | n23374 ;
  assign n23376 = n5494 | n23375 ;
  assign n23377 = ( n10664 & n12549 ) | ( n10664 & ~n15031 ) | ( n12549 & ~n15031 ) ;
  assign n23378 = n23377 ^ n19404 ^ n8562 ;
  assign n23379 = n21367 ^ n20287 ^ n10501 ;
  assign n23380 = n23379 ^ n1814 ^ 1'b0 ;
  assign n23381 = n5008 | n13997 ;
  assign n23382 = n10647 & n12368 ;
  assign n23383 = n23382 ^ n10253 ^ 1'b0 ;
  assign n23384 = ~n19290 & n23383 ;
  assign n23386 = n4328 & n10804 ;
  assign n23385 = ~n2324 & n19370 ;
  assign n23387 = n23386 ^ n23385 ^ 1'b0 ;
  assign n23388 = n1318 ^ n541 ^ 1'b0 ;
  assign n23389 = n13119 | n23388 ;
  assign n23390 = ( ~n394 & n8948 ) | ( ~n394 & n17349 ) | ( n8948 & n17349 ) ;
  assign n23391 = n6594 ^ n3473 ^ 1'b0 ;
  assign n23393 = n19521 ^ n13967 ^ n12870 ;
  assign n23392 = ~n3726 & n18417 ;
  assign n23394 = n23393 ^ n23392 ^ 1'b0 ;
  assign n23395 = n21474 ^ n2051 ^ 1'b0 ;
  assign n23396 = n4706 & ~n23395 ;
  assign n23397 = n11383 ^ n10065 ^ n4851 ;
  assign n23398 = n5025 & ~n23397 ;
  assign n23399 = n23398 ^ n5081 ^ 1'b0 ;
  assign n23400 = ~n4093 & n12763 ;
  assign n23401 = n20649 & n23400 ;
  assign n23402 = n16169 & ~n23401 ;
  assign n23403 = n23402 ^ n13539 ^ 1'b0 ;
  assign n23404 = n19166 ^ n12477 ^ n12008 ;
  assign n23406 = n13585 ^ n6228 ^ n4983 ;
  assign n23405 = n17029 | n18400 ;
  assign n23407 = n23406 ^ n23405 ^ n2559 ;
  assign n23408 = ( n12504 & n12630 ) | ( n12504 & ~n22632 ) | ( n12630 & ~n22632 ) ;
  assign n23409 = n16597 ^ n11381 ^ n9493 ;
  assign n23410 = ( n7973 & n18072 ) | ( n7973 & ~n23409 ) | ( n18072 & ~n23409 ) ;
  assign n23411 = ~n3346 & n22513 ;
  assign n23412 = n14442 ^ n9682 ^ n5249 ;
  assign n23413 = n17677 ^ n7633 ^ 1'b0 ;
  assign n23414 = ( n6156 & n15412 ) | ( n6156 & ~n23413 ) | ( n15412 & ~n23413 ) ;
  assign n23415 = n20320 ^ n19876 ^ 1'b0 ;
  assign n23416 = n20737 ^ n17138 ^ n13288 ;
  assign n23417 = n11594 ^ n9823 ^ 1'b0 ;
  assign n23418 = ( ~n4683 & n13118 ) | ( ~n4683 & n17136 ) | ( n13118 & n17136 ) ;
  assign n23419 = ( n5316 & n6699 ) | ( n5316 & ~n22148 ) | ( n6699 & ~n22148 ) ;
  assign n23420 = n23419 ^ n20268 ^ n19828 ;
  assign n23421 = n12354 ^ n7463 ^ n1677 ;
  assign n23422 = ( ~x106 & n1767 ) | ( ~x106 & n15441 ) | ( n1767 & n15441 ) ;
  assign n23423 = n23422 ^ n314 ^ 1'b0 ;
  assign n23424 = n23423 ^ n17537 ^ n1945 ;
  assign n23426 = n11433 ^ n9379 ^ n1049 ;
  assign n23425 = n5046 | n6529 ;
  assign n23427 = n23426 ^ n23425 ^ 1'b0 ;
  assign n23428 = ~n17511 & n23427 ;
  assign n23429 = n792 & n7425 ;
  assign n23430 = n23429 ^ n4674 ^ 1'b0 ;
  assign n23431 = n23430 ^ n21911 ^ 1'b0 ;
  assign n23432 = n8668 & n23431 ;
  assign n23434 = n4467 & ~n7816 ;
  assign n23435 = n23434 ^ n15495 ^ 1'b0 ;
  assign n23433 = n1660 ^ n892 ^ x25 ;
  assign n23436 = n23435 ^ n23433 ^ n3716 ;
  assign n23437 = ( ~n11031 & n18769 ) | ( ~n11031 & n23436 ) | ( n18769 & n23436 ) ;
  assign n23440 = n3830 | n9828 ;
  assign n23441 = n7467 ^ n2807 ^ 1'b0 ;
  assign n23442 = n23440 & ~n23441 ;
  assign n23439 = n3749 ^ n2002 ^ n1233 ;
  assign n23438 = n9121 ^ n5693 ^ 1'b0 ;
  assign n23443 = n23442 ^ n23439 ^ n23438 ;
  assign n23444 = n23079 ^ n22517 ^ n5379 ;
  assign n23445 = n7024 & ~n20681 ;
  assign n23446 = n17376 ^ n6963 ^ n969 ;
  assign n23447 = n23446 ^ n2002 ^ n199 ;
  assign n23448 = n3496 & n6350 ;
  assign n23449 = n23448 ^ n9408 ^ 1'b0 ;
  assign n23450 = n5026 | n14124 ;
  assign n23451 = n7687 | n23450 ;
  assign n23452 = ( n2217 & n6290 ) | ( n2217 & ~n15918 ) | ( n6290 & ~n15918 ) ;
  assign n23453 = n2751 & n23452 ;
  assign n23454 = ( n437 & n8335 ) | ( n437 & ~n23453 ) | ( n8335 & ~n23453 ) ;
  assign n23455 = ( n16926 & ~n23451 ) | ( n16926 & n23454 ) | ( ~n23451 & n23454 ) ;
  assign n23456 = n23455 ^ n12228 ^ 1'b0 ;
  assign n23457 = n1091 | n6024 ;
  assign n23458 = ( ~n4913 & n9141 ) | ( ~n4913 & n15074 ) | ( n9141 & n15074 ) ;
  assign n23459 = n23458 ^ n3390 ^ 1'b0 ;
  assign n23460 = n23457 & n23459 ;
  assign n23461 = ( n2493 & n2515 ) | ( n2493 & ~n6317 ) | ( n2515 & ~n6317 ) ;
  assign n23462 = ( n2026 & n5935 ) | ( n2026 & n11107 ) | ( n5935 & n11107 ) ;
  assign n23463 = n250 | n7096 ;
  assign n23464 = n16284 & ~n23463 ;
  assign n23465 = n4080 ^ n1025 ^ 1'b0 ;
  assign n23466 = ( n4627 & n23464 ) | ( n4627 & ~n23465 ) | ( n23464 & ~n23465 ) ;
  assign n23467 = n11211 ^ n9008 ^ 1'b0 ;
  assign n23468 = n23467 ^ n13712 ^ 1'b0 ;
  assign n23469 = n10401 | n11216 ;
  assign n23470 = n7143 ^ n5492 ^ 1'b0 ;
  assign n23471 = n5330 ^ x12 ^ 1'b0 ;
  assign n23472 = n22376 | n23471 ;
  assign n23473 = n9788 ^ n402 ^ 1'b0 ;
  assign n23474 = n23472 & ~n23473 ;
  assign n23475 = n9822 & ~n15054 ;
  assign n23476 = n23475 ^ n8348 ^ 1'b0 ;
  assign n23477 = ( n7875 & n23474 ) | ( n7875 & n23476 ) | ( n23474 & n23476 ) ;
  assign n23478 = n19211 & n23477 ;
  assign n23479 = n13690 ^ n11619 ^ 1'b0 ;
  assign n23480 = n23479 ^ n19438 ^ 1'b0 ;
  assign n23485 = ( n3201 & n12924 ) | ( n3201 & ~n12966 ) | ( n12924 & ~n12966 ) ;
  assign n23484 = n19836 ^ n4491 ^ 1'b0 ;
  assign n23486 = n23485 ^ n23484 ^ n2291 ;
  assign n23481 = n8265 ^ n7463 ^ n7362 ;
  assign n23482 = n23481 ^ n18671 ^ 1'b0 ;
  assign n23483 = ~n2924 & n23482 ;
  assign n23487 = n23486 ^ n23483 ^ 1'b0 ;
  assign n23488 = n13466 ^ n11335 ^ 1'b0 ;
  assign n23489 = ~n3825 & n23488 ;
  assign n23490 = n23489 ^ n13800 ^ n1912 ;
  assign n23491 = ~n4721 & n11876 ;
  assign n23492 = n1911 & n3759 ;
  assign n23493 = n8243 & n23492 ;
  assign n23494 = ( ~n3448 & n18232 ) | ( ~n3448 & n23493 ) | ( n18232 & n23493 ) ;
  assign n23495 = ( n4105 & ~n23491 ) | ( n4105 & n23494 ) | ( ~n23491 & n23494 ) ;
  assign n23496 = ( n4048 & n10052 ) | ( n4048 & n18792 ) | ( n10052 & n18792 ) ;
  assign n23497 = n23496 ^ n21814 ^ n16766 ;
  assign n23498 = n6681 ^ n2826 ^ n1295 ;
  assign n23499 = n1392 | n6986 ;
  assign n23500 = n1601 | n7105 ;
  assign n23501 = n23500 ^ n3561 ^ 1'b0 ;
  assign n23502 = n5644 ^ n3359 ^ n328 ;
  assign n23503 = n8885 & n23502 ;
  assign n23504 = n23503 ^ n12793 ^ 1'b0 ;
  assign n23505 = ( ~n18422 & n23501 ) | ( ~n18422 & n23504 ) | ( n23501 & n23504 ) ;
  assign n23506 = ( ~n2917 & n7961 ) | ( ~n2917 & n17506 ) | ( n7961 & n17506 ) ;
  assign n23507 = ( n23499 & ~n23505 ) | ( n23499 & n23506 ) | ( ~n23505 & n23506 ) ;
  assign n23508 = n9493 ^ n8690 ^ n5663 ;
  assign n23509 = n23508 ^ n13542 ^ n10397 ;
  assign n23510 = n9554 & n11880 ;
  assign n23511 = ~n23509 & n23510 ;
  assign n23512 = ~n583 & n17567 ;
  assign n23513 = n9474 & n23512 ;
  assign n23514 = n20681 & ~n23513 ;
  assign n23515 = n3805 & n10247 ;
  assign n23516 = ~n22776 & n23515 ;
  assign n23517 = n19069 ^ n10527 ^ 1'b0 ;
  assign n23518 = n21434 & ~n23517 ;
  assign n23519 = ( ~n586 & n4215 ) | ( ~n586 & n14904 ) | ( n4215 & n14904 ) ;
  assign n23520 = ( n20964 & n22331 ) | ( n20964 & n23519 ) | ( n22331 & n23519 ) ;
  assign n23521 = n4259 ^ n3848 ^ n3593 ;
  assign n23522 = n4765 ^ n1447 ^ 1'b0 ;
  assign n23523 = n160 | n250 ;
  assign n23524 = n23523 ^ n5018 ^ 1'b0 ;
  assign n23525 = ( n7542 & n23522 ) | ( n7542 & ~n23524 ) | ( n23522 & ~n23524 ) ;
  assign n23526 = ( n15143 & n23521 ) | ( n15143 & n23525 ) | ( n23521 & n23525 ) ;
  assign n23527 = ( n684 & ~n8931 ) | ( n684 & n19256 ) | ( ~n8931 & n19256 ) ;
  assign n23528 = ( n2709 & ~n10685 ) | ( n2709 & n16840 ) | ( ~n10685 & n16840 ) ;
  assign n23529 = ( n670 & ~n15046 ) | ( n670 & n23528 ) | ( ~n15046 & n23528 ) ;
  assign n23530 = ~n5733 & n22617 ;
  assign n23531 = n23530 ^ n7823 ^ 1'b0 ;
  assign n23533 = n8814 ^ n3841 ^ 1'b0 ;
  assign n23532 = ( n8507 & n11545 ) | ( n8507 & n16992 ) | ( n11545 & n16992 ) ;
  assign n23534 = n23533 ^ n23532 ^ n1439 ;
  assign n23535 = ( n3369 & ~n9729 ) | ( n3369 & n23534 ) | ( ~n9729 & n23534 ) ;
  assign n23536 = n8659 & ~n10113 ;
  assign n23537 = ~x67 & n23536 ;
  assign n23538 = n21730 ^ n664 ^ 1'b0 ;
  assign n23539 = ~n23537 & n23538 ;
  assign n23540 = n4353 & n23539 ;
  assign n23541 = ~n23535 & n23540 ;
  assign n23542 = n506 | n3154 ;
  assign n23543 = n13429 ^ n10551 ^ n7678 ;
  assign n23544 = ( n7890 & ~n23542 ) | ( n7890 & n23543 ) | ( ~n23542 & n23543 ) ;
  assign n23545 = ~n10636 & n17442 ;
  assign n23547 = ( n6185 & ~n10350 ) | ( n6185 & n10927 ) | ( ~n10350 & n10927 ) ;
  assign n23546 = n18634 ^ n5931 ^ n2185 ;
  assign n23548 = n23547 ^ n23546 ^ n4352 ;
  assign n23549 = ( n10359 & n12357 ) | ( n10359 & ~n22877 ) | ( n12357 & ~n22877 ) ;
  assign n23551 = ( x70 & n8232 ) | ( x70 & n14749 ) | ( n8232 & n14749 ) ;
  assign n23550 = n9829 | n14193 ;
  assign n23552 = n23551 ^ n23550 ^ 1'b0 ;
  assign n23554 = ( n6837 & n7225 ) | ( n6837 & n8510 ) | ( n7225 & n8510 ) ;
  assign n23553 = n21124 ^ n8810 ^ n5086 ;
  assign n23555 = n23554 ^ n23553 ^ n14520 ;
  assign n23556 = ~n6908 & n23555 ;
  assign n23557 = ( n12286 & n23552 ) | ( n12286 & ~n23556 ) | ( n23552 & ~n23556 ) ;
  assign n23558 = n4080 | n4108 ;
  assign n23559 = n23558 ^ n4736 ^ 1'b0 ;
  assign n23560 = ( n505 & n15711 ) | ( n505 & ~n23559 ) | ( n15711 & ~n23559 ) ;
  assign n23561 = n4353 ^ n3022 ^ 1'b0 ;
  assign n23562 = n23561 ^ n16216 ^ n6913 ;
  assign n23563 = n23562 ^ n14676 ^ 1'b0 ;
  assign n23564 = n10674 ^ n9444 ^ 1'b0 ;
  assign n23565 = n11884 & ~n23564 ;
  assign n23566 = n10358 & n21201 ;
  assign n23567 = n7260 & n23566 ;
  assign n23568 = n6891 | n7789 ;
  assign n23569 = ( n2543 & n9759 ) | ( n2543 & ~n23568 ) | ( n9759 & ~n23568 ) ;
  assign n23570 = n13950 | n15610 ;
  assign n23571 = n23570 ^ n19817 ^ 1'b0 ;
  assign n23572 = ( n8914 & n9628 ) | ( n8914 & n23571 ) | ( n9628 & n23571 ) ;
  assign n23573 = n10998 ^ n6198 ^ 1'b0 ;
  assign n23574 = ( n6104 & n8952 ) | ( n6104 & n19608 ) | ( n8952 & n19608 ) ;
  assign n23575 = ( n20321 & ~n23573 ) | ( n20321 & n23574 ) | ( ~n23573 & n23574 ) ;
  assign n23577 = n12000 ^ n8413 ^ 1'b0 ;
  assign n23578 = n5661 & ~n23577 ;
  assign n23576 = n2678 ^ n1246 ^ 1'b0 ;
  assign n23579 = n23578 ^ n23576 ^ n8721 ;
  assign n23581 = ( n4305 & n11515 ) | ( n4305 & ~n14053 ) | ( n11515 & ~n14053 ) ;
  assign n23580 = n438 | n1599 ;
  assign n23582 = n23581 ^ n23580 ^ n14584 ;
  assign n23594 = ( n3666 & n8146 ) | ( n3666 & ~n18265 ) | ( n8146 & ~n18265 ) ;
  assign n23583 = n1360 & ~n2974 ;
  assign n23584 = n1153 & ~n15684 ;
  assign n23585 = n23584 ^ n1572 ^ 1'b0 ;
  assign n23586 = ( n20632 & n23583 ) | ( n20632 & n23585 ) | ( n23583 & n23585 ) ;
  assign n23587 = n6033 | n15414 ;
  assign n23588 = n5115 & n23587 ;
  assign n23589 = ~n146 & n23588 ;
  assign n23590 = n8780 & n23589 ;
  assign n23591 = n23590 ^ n15768 ^ 1'b0 ;
  assign n23592 = ~n23586 & n23591 ;
  assign n23593 = n23592 ^ n14676 ^ n2433 ;
  assign n23595 = n23594 ^ n23593 ^ n22084 ;
  assign n23596 = ~n1227 & n2021 ;
  assign n23597 = n9077 & n23596 ;
  assign n23598 = n2546 & ~n9663 ;
  assign n23599 = n23597 & n23598 ;
  assign n23600 = ~n16305 & n22945 ;
  assign n23601 = n23052 & n23600 ;
  assign n23602 = n11432 | n19420 ;
  assign n23603 = n9923 & n16891 ;
  assign n23604 = n23603 ^ n14111 ^ 1'b0 ;
  assign n23605 = n13248 ^ n10035 ^ n4141 ;
  assign n23608 = ( ~n2845 & n9276 ) | ( ~n2845 & n9711 ) | ( n9276 & n9711 ) ;
  assign n23606 = ( n2520 & ~n4539 ) | ( n2520 & n12902 ) | ( ~n4539 & n12902 ) ;
  assign n23607 = ~n5467 & n23606 ;
  assign n23609 = n23608 ^ n23607 ^ 1'b0 ;
  assign n23610 = n3138 & n23609 ;
  assign n23611 = ~n526 & n15558 ;
  assign n23612 = n23611 ^ n19094 ^ n14236 ;
  assign n23613 = n15756 ^ n9986 ^ 1'b0 ;
  assign n23614 = n10996 & n23613 ;
  assign n23615 = ~n12549 & n16556 ;
  assign n23616 = ~n20146 & n23615 ;
  assign n23617 = n18398 & n19888 ;
  assign n23618 = ( n1522 & ~n4564 ) | ( n1522 & n16071 ) | ( ~n4564 & n16071 ) ;
  assign n23619 = n16152 ^ n8734 ^ n5704 ;
  assign n23620 = n23618 | n23619 ;
  assign n23621 = n19483 ^ n18376 ^ n9478 ;
  assign n23622 = n23621 ^ n15117 ^ n9291 ;
  assign n23623 = n11166 ^ n5125 ^ n511 ;
  assign n23625 = n8670 ^ n4372 ^ 1'b0 ;
  assign n23624 = n3256 | n19519 ;
  assign n23626 = n23625 ^ n23624 ^ 1'b0 ;
  assign n23627 = ~n14636 & n23626 ;
  assign n23628 = n10739 & n15930 ;
  assign n23629 = n23628 ^ n1177 ^ 1'b0 ;
  assign n23630 = n15266 ^ n14353 ^ 1'b0 ;
  assign n23631 = ( n1933 & n13732 ) | ( n1933 & ~n23630 ) | ( n13732 & ~n23630 ) ;
  assign n23632 = n16540 ^ n11860 ^ n775 ;
  assign n23633 = n23535 ^ n13585 ^ 1'b0 ;
  assign n23634 = n22985 ^ n22188 ^ n376 ;
  assign n23635 = n7645 ^ x55 ^ 1'b0 ;
  assign n23636 = ~n7884 & n23635 ;
  assign n23637 = ( ~n13769 & n23634 ) | ( ~n13769 & n23636 ) | ( n23634 & n23636 ) ;
  assign n23638 = n23637 ^ n21835 ^ n4139 ;
  assign n23639 = ( n3665 & ~n6564 ) | ( n3665 & n17075 ) | ( ~n6564 & n17075 ) ;
  assign n23640 = n18374 ^ n12732 ^ 1'b0 ;
  assign n23641 = n23639 & n23640 ;
  assign n23650 = n13056 ^ n12903 ^ n11383 ;
  assign n23651 = n23650 ^ n17281 ^ 1'b0 ;
  assign n23644 = ( n4953 & n6326 ) | ( n4953 & ~n22706 ) | ( n6326 & ~n22706 ) ;
  assign n23642 = ( n2373 & n5159 ) | ( n2373 & n19903 ) | ( n5159 & n19903 ) ;
  assign n23643 = ~n1602 & n23642 ;
  assign n23645 = n23644 ^ n23643 ^ n3048 ;
  assign n23646 = n3816 & n18791 ;
  assign n23647 = n11811 & n23646 ;
  assign n23648 = n23647 ^ n10840 ^ 1'b0 ;
  assign n23649 = n23645 & n23648 ;
  assign n23652 = n23651 ^ n23649 ^ 1'b0 ;
  assign n23653 = n15713 ^ n13517 ^ 1'b0 ;
  assign n23654 = ~n6789 & n15350 ;
  assign n23655 = n23654 ^ n9561 ^ n5149 ;
  assign n23656 = n5711 & n11330 ;
  assign n23657 = ~n9407 & n12987 ;
  assign n23658 = n23261 ^ n12715 ^ n3438 ;
  assign n23659 = n1504 | n23658 ;
  assign n23660 = n23659 ^ n8617 ^ 1'b0 ;
  assign n23661 = n18060 ^ n14687 ^ 1'b0 ;
  assign n23662 = n16702 & n23554 ;
  assign n23663 = n23661 & n23662 ;
  assign n23665 = n18764 ^ n8201 ^ n6250 ;
  assign n23664 = n11400 & ~n14526 ;
  assign n23666 = n23665 ^ n23664 ^ 1'b0 ;
  assign n23667 = n7777 ^ n6176 ^ 1'b0 ;
  assign n23668 = ( n11980 & ~n19958 ) | ( n11980 & n23667 ) | ( ~n19958 & n23667 ) ;
  assign n23669 = n23668 ^ n6501 ^ 1'b0 ;
  assign n23670 = ~n18770 & n23669 ;
  assign n23671 = n12222 ^ n10671 ^ 1'b0 ;
  assign n23672 = n16165 & ~n23671 ;
  assign n23673 = ( ~n1111 & n15174 ) | ( ~n1111 & n21891 ) | ( n15174 & n21891 ) ;
  assign n23674 = n8093 ^ n3490 ^ 1'b0 ;
  assign n23675 = ( n3828 & ~n17319 ) | ( n3828 & n23674 ) | ( ~n17319 & n23674 ) ;
  assign n23676 = n2376 & ~n3202 ;
  assign n23677 = ( ~n1996 & n2390 ) | ( ~n1996 & n10342 ) | ( n2390 & n10342 ) ;
  assign n23678 = ( n4608 & n12577 ) | ( n4608 & n23677 ) | ( n12577 & n23677 ) ;
  assign n23679 = ~n6860 & n16203 ;
  assign n23680 = ~n3141 & n23679 ;
  assign n23681 = n915 & ~n23680 ;
  assign n23682 = n23681 ^ n7568 ^ 1'b0 ;
  assign n23683 = n10534 & ~n13767 ;
  assign n23684 = n844 & n7055 ;
  assign n23685 = n16537 ^ n15345 ^ n9886 ;
  assign n23686 = ( n7582 & n23684 ) | ( n7582 & n23685 ) | ( n23684 & n23685 ) ;
  assign n23687 = ~n23683 & n23686 ;
  assign n23688 = n3461 | n14782 ;
  assign n23689 = n23687 | n23688 ;
  assign n23690 = n16880 ^ n6626 ^ n3703 ;
  assign n23691 = ( n9189 & ~n9660 ) | ( n9189 & n23690 ) | ( ~n9660 & n23690 ) ;
  assign n23692 = n18945 ^ n10861 ^ n2324 ;
  assign n23693 = n14522 & ~n23692 ;
  assign n23694 = n8490 ^ n6836 ^ 1'b0 ;
  assign n23695 = ( n2678 & n3115 ) | ( n2678 & ~n7968 ) | ( n3115 & ~n7968 ) ;
  assign n23696 = n23694 & n23695 ;
  assign n23697 = ~n22340 & n23696 ;
  assign n23698 = n5134 & ~n9339 ;
  assign n23699 = n23698 ^ n21573 ^ 1'b0 ;
  assign n23700 = n11698 & ~n14857 ;
  assign n23701 = ~n10890 & n23700 ;
  assign n23702 = n9657 & n10170 ;
  assign n23703 = n23702 ^ n6731 ^ n3932 ;
  assign n23704 = ( n9363 & n16248 ) | ( n9363 & ~n23703 ) | ( n16248 & ~n23703 ) ;
  assign n23705 = n12273 ^ n5051 ^ n2147 ;
  assign n23706 = n23705 ^ n19343 ^ n2312 ;
  assign n23707 = ( n2046 & n6897 ) | ( n2046 & n18376 ) | ( n6897 & n18376 ) ;
  assign n23708 = n23707 ^ n7187 ^ n5490 ;
  assign n23709 = n1490 | n9015 ;
  assign n23710 = n7859 | n23362 ;
  assign n23711 = n20222 ^ n9964 ^ 1'b0 ;
  assign n23712 = n23711 ^ n20142 ^ 1'b0 ;
  assign n23713 = n23710 & ~n23712 ;
  assign n23716 = ~n2144 & n11400 ;
  assign n23717 = n23716 ^ n8017 ^ 1'b0 ;
  assign n23714 = n5518 | n8215 ;
  assign n23715 = n23714 ^ n2361 ^ 1'b0 ;
  assign n23718 = n23717 ^ n23715 ^ n5304 ;
  assign n23719 = ( n16202 & ~n17798 ) | ( n16202 & n23718 ) | ( ~n17798 & n23718 ) ;
  assign n23720 = ( n6070 & n9587 ) | ( n6070 & n16140 ) | ( n9587 & n16140 ) ;
  assign n23721 = ~n23719 & n23720 ;
  assign n23724 = ( n844 & n4092 ) | ( n844 & n7600 ) | ( n4092 & n7600 ) ;
  assign n23722 = n9359 | n14139 ;
  assign n23723 = n23722 ^ n7069 ^ 1'b0 ;
  assign n23725 = n23724 ^ n23723 ^ n11632 ;
  assign n23726 = ( n294 & n23406 ) | ( n294 & ~n23725 ) | ( n23406 & ~n23725 ) ;
  assign n23727 = n12892 ^ n11278 ^ 1'b0 ;
  assign n23728 = ( ~n3242 & n7734 ) | ( ~n3242 & n10909 ) | ( n7734 & n10909 ) ;
  assign n23729 = n23728 ^ n5483 ^ 1'b0 ;
  assign n23731 = ( n890 & n4442 ) | ( n890 & n4554 ) | ( n4442 & n4554 ) ;
  assign n23730 = ( n1122 & n14418 ) | ( n1122 & n15492 ) | ( n14418 & n15492 ) ;
  assign n23732 = n23731 ^ n23730 ^ n1808 ;
  assign n23733 = ( n1839 & n3626 ) | ( n1839 & ~n13036 ) | ( n3626 & ~n13036 ) ;
  assign n23734 = ( n10443 & ~n18763 ) | ( n10443 & n23733 ) | ( ~n18763 & n23733 ) ;
  assign n23735 = n23734 ^ n16485 ^ 1'b0 ;
  assign n23736 = n23732 & n23735 ;
  assign n23737 = ( n7510 & n11434 ) | ( n7510 & n19124 ) | ( n11434 & n19124 ) ;
  assign n23738 = ~n1916 & n12893 ;
  assign n23739 = n23738 ^ n10673 ^ n2862 ;
  assign n23740 = n23739 ^ n10743 ^ 1'b0 ;
  assign n23741 = n23737 | n23740 ;
  assign n23742 = n12130 ^ n6920 ^ 1'b0 ;
  assign n23743 = n17570 ^ n16226 ^ n12674 ;
  assign n23747 = n10993 & ~n19063 ;
  assign n23748 = ~n12465 & n23747 ;
  assign n23744 = n3049 & n17171 ;
  assign n23745 = n23744 ^ n9448 ^ 1'b0 ;
  assign n23746 = n23745 ^ n14052 ^ n1938 ;
  assign n23749 = n23748 ^ n23746 ^ n20416 ;
  assign n23755 = n13173 ^ n2747 ^ n2450 ;
  assign n23756 = n23755 ^ n10533 ^ 1'b0 ;
  assign n23757 = n13473 & n23756 ;
  assign n23758 = n23757 ^ n8507 ^ 1'b0 ;
  assign n23750 = n11515 ^ n8756 ^ n2523 ;
  assign n23751 = n8660 ^ n7069 ^ 1'b0 ;
  assign n23752 = ~n686 & n23751 ;
  assign n23753 = ( ~n4587 & n23750 ) | ( ~n4587 & n23752 ) | ( n23750 & n23752 ) ;
  assign n23754 = n5631 & ~n23753 ;
  assign n23759 = n23758 ^ n23754 ^ n9366 ;
  assign n23764 = n14705 ^ n8571 ^ 1'b0 ;
  assign n23760 = n6047 ^ n5098 ^ 1'b0 ;
  assign n23761 = ( n5925 & n10877 ) | ( n5925 & ~n23760 ) | ( n10877 & ~n23760 ) ;
  assign n23762 = n9019 | n23761 ;
  assign n23763 = n23762 ^ n16570 ^ 1'b0 ;
  assign n23765 = n23764 ^ n23763 ^ n16368 ;
  assign n23766 = n5991 ^ n1843 ^ 1'b0 ;
  assign n23767 = n4484 ^ n1666 ^ 1'b0 ;
  assign n23768 = n2733 & ~n23767 ;
  assign n23769 = n7229 & n23768 ;
  assign n23770 = n6832 & n23769 ;
  assign n23771 = ~n474 & n23138 ;
  assign n23772 = n8283 & n23771 ;
  assign n23773 = n1917 | n6187 ;
  assign n23774 = n23772 & ~n23773 ;
  assign n23775 = n9313 ^ n8856 ^ 1'b0 ;
  assign n23776 = ~n9222 & n23775 ;
  assign n23777 = ( ~n6409 & n17958 ) | ( ~n6409 & n23776 ) | ( n17958 & n23776 ) ;
  assign n23778 = n19046 ^ n12365 ^ n4632 ;
  assign n23779 = ( n9695 & ~n13295 ) | ( n9695 & n18557 ) | ( ~n13295 & n18557 ) ;
  assign n23780 = ( n12680 & ~n14918 ) | ( n12680 & n23779 ) | ( ~n14918 & n23779 ) ;
  assign n23782 = n17267 ^ n7402 ^ n6643 ;
  assign n23781 = n4209 & n16515 ;
  assign n23783 = n23782 ^ n23781 ^ 1'b0 ;
  assign n23784 = n1332 & n4982 ;
  assign n23785 = n23784 ^ n20584 ^ 1'b0 ;
  assign n23786 = n1414 ^ n951 ^ 1'b0 ;
  assign n23787 = n17773 & n23786 ;
  assign n23788 = ( n1999 & n11925 ) | ( n1999 & n23690 ) | ( n11925 & n23690 ) ;
  assign n23789 = n14958 ^ n5921 ^ n4616 ;
  assign n23790 = ( n4452 & n11133 ) | ( n4452 & ~n23789 ) | ( n11133 & ~n23789 ) ;
  assign n23791 = n19353 ^ n2488 ^ n785 ;
  assign n23792 = n23791 ^ n15306 ^ n2329 ;
  assign n23793 = n14343 ^ n2259 ^ n1946 ;
  assign n23794 = ( n10241 & n17939 ) | ( n10241 & n23793 ) | ( n17939 & n23793 ) ;
  assign n23795 = n10695 ^ n7178 ^ n4634 ;
  assign n23796 = n6492 & n11793 ;
  assign n23797 = n23796 ^ n2688 ^ 1'b0 ;
  assign n23798 = n23795 | n23797 ;
  assign n23799 = n23798 ^ n3967 ^ n1186 ;
  assign n23800 = n2472 ^ x101 ^ 1'b0 ;
  assign n23801 = n23800 ^ n6576 ^ 1'b0 ;
  assign n23802 = ~n8380 & n23801 ;
  assign n23803 = n3953 | n10864 ;
  assign n23804 = n11736 ^ x103 ^ 1'b0 ;
  assign n23805 = n23803 & ~n23804 ;
  assign n23806 = n2725 & ~n7929 ;
  assign n23807 = n692 ^ n405 ^ 1'b0 ;
  assign n23808 = n3080 & ~n23807 ;
  assign n23809 = ( n1096 & n1736 ) | ( n1096 & ~n4022 ) | ( n1736 & ~n4022 ) ;
  assign n23810 = ( ~n14799 & n23791 ) | ( ~n14799 & n23809 ) | ( n23791 & n23809 ) ;
  assign n23811 = ( n829 & n1132 ) | ( n829 & ~n7423 ) | ( n1132 & ~n7423 ) ;
  assign n23812 = ~n5773 & n13939 ;
  assign n23813 = n23812 ^ n7116 ^ 1'b0 ;
  assign n23814 = n23813 ^ n4229 ^ n1771 ;
  assign n23815 = ( n20157 & ~n23811 ) | ( n20157 & n23814 ) | ( ~n23811 & n23814 ) ;
  assign n23817 = ~n165 & n4144 ;
  assign n23818 = ~n5111 & n23817 ;
  assign n23816 = n12430 | n18427 ;
  assign n23819 = n23818 ^ n23816 ^ 1'b0 ;
  assign n23820 = ( n12989 & n13523 ) | ( n12989 & n23819 ) | ( n13523 & n23819 ) ;
  assign n23821 = n3159 & n18474 ;
  assign n23822 = n19054 ^ n5605 ^ n2889 ;
  assign n23823 = n471 | n1221 ;
  assign n23824 = n11156 & ~n23823 ;
  assign n23825 = n18185 ^ n11106 ^ 1'b0 ;
  assign n23826 = ( n23822 & ~n23824 ) | ( n23822 & n23825 ) | ( ~n23824 & n23825 ) ;
  assign n23827 = n12892 ^ n8202 ^ n1359 ;
  assign n23828 = n16549 ^ n9034 ^ x35 ;
  assign n23829 = n11156 | n23828 ;
  assign n23830 = n23827 | n23829 ;
  assign n23831 = n9446 ^ n6997 ^ 1'b0 ;
  assign n23832 = ( n854 & n2443 ) | ( n854 & n23831 ) | ( n2443 & n23831 ) ;
  assign n23833 = n23832 ^ n12395 ^ n1635 ;
  assign n23834 = ~n6610 & n10248 ;
  assign n23835 = ~n23833 & n23834 ;
  assign n23836 = ~n3645 & n12598 ;
  assign n23837 = n23836 ^ n1729 ^ 1'b0 ;
  assign n23838 = ( n5985 & ~n8674 ) | ( n5985 & n23837 ) | ( ~n8674 & n23837 ) ;
  assign n23839 = ( n6926 & n11023 ) | ( n6926 & ~n11337 ) | ( n11023 & ~n11337 ) ;
  assign n23840 = ( ~n3860 & n5012 ) | ( ~n3860 & n5512 ) | ( n5012 & n5512 ) ;
  assign n23841 = n3261 ^ n2784 ^ 1'b0 ;
  assign n23842 = n23840 & n23841 ;
  assign n23843 = n17386 ^ n8624 ^ 1'b0 ;
  assign n23844 = ~n18636 & n23843 ;
  assign n23845 = n12778 & n20114 ;
  assign n23846 = n23845 ^ n16749 ^ 1'b0 ;
  assign n23847 = ~n14806 & n15980 ;
  assign n23848 = ( n11932 & n15080 ) | ( n11932 & n23847 ) | ( n15080 & n23847 ) ;
  assign n23849 = n21574 ^ n13955 ^ n2321 ;
  assign n23850 = ( n3964 & ~n6679 ) | ( n3964 & n16369 ) | ( ~n6679 & n16369 ) ;
  assign n23851 = ( ~n986 & n2416 ) | ( ~n986 & n15225 ) | ( n2416 & n15225 ) ;
  assign n23852 = n23851 ^ n18390 ^ n16931 ;
  assign n23853 = n677 | n5714 ;
  assign n23854 = n23212 ^ n19030 ^ n4135 ;
  assign n23855 = ~n3312 & n21684 ;
  assign n23856 = n5980 & n23855 ;
  assign n23857 = n20241 ^ n2948 ^ 1'b0 ;
  assign n23858 = n9719 ^ n4285 ^ n3592 ;
  assign n23859 = ~n21230 & n23858 ;
  assign n23860 = n2587 & n20439 ;
  assign n23861 = n23860 ^ n6761 ^ 1'b0 ;
  assign n23862 = n15604 & n23861 ;
  assign n23863 = n22351 ^ n6598 ^ 1'b0 ;
  assign n23864 = n15993 ^ n10949 ^ n5247 ;
  assign n23865 = n23864 ^ n4968 ^ n725 ;
  assign n23866 = ( n1076 & n12712 ) | ( n1076 & n17133 ) | ( n12712 & n17133 ) ;
  assign n23868 = n5504 & n11855 ;
  assign n23867 = n3704 & n20761 ;
  assign n23869 = n23868 ^ n23867 ^ n8648 ;
  assign n23870 = ( n9740 & n10213 ) | ( n9740 & n18023 ) | ( n10213 & n18023 ) ;
  assign n23871 = n11609 | n23870 ;
  assign n23872 = n20937 ^ n2624 ^ 1'b0 ;
  assign n23873 = ~n7215 & n23872 ;
  assign n23874 = n17521 | n23873 ;
  assign n23875 = n7598 | n8814 ;
  assign n23876 = x96 | n23875 ;
  assign n23877 = n4594 & ~n20104 ;
  assign n23878 = n23877 ^ n11436 ^ 1'b0 ;
  assign n23879 = n6735 & n7764 ;
  assign n23880 = n822 & n23879 ;
  assign n23881 = n23880 ^ n3251 ^ 1'b0 ;
  assign n23882 = n23881 ^ n20372 ^ n7809 ;
  assign n23883 = ( n13041 & n15587 ) | ( n13041 & n17009 ) | ( n15587 & n17009 ) ;
  assign n23884 = n6540 ^ n4639 ^ n3392 ;
  assign n23885 = n9363 ^ n7104 ^ 1'b0 ;
  assign n23886 = ~n7597 & n23885 ;
  assign n23887 = n13648 ^ n6049 ^ 1'b0 ;
  assign n23888 = ( n308 & n23886 ) | ( n308 & n23887 ) | ( n23886 & n23887 ) ;
  assign n23889 = n3298 | n4174 ;
  assign n23890 = n2033 | n23889 ;
  assign n23891 = n22968 | n23890 ;
  assign n23892 = n5353 ^ n3877 ^ 1'b0 ;
  assign n23893 = n19347 & ~n23892 ;
  assign n23894 = n23891 & n23893 ;
  assign n23895 = n7425 & n12723 ;
  assign n23896 = ~n3588 & n23895 ;
  assign n23897 = n5672 & ~n9387 ;
  assign n23898 = n20625 ^ n8919 ^ n3977 ;
  assign n23899 = n23898 ^ n13298 ^ n9756 ;
  assign n23900 = ( n7783 & ~n9119 ) | ( n7783 & n9759 ) | ( ~n9119 & n9759 ) ;
  assign n23901 = n9664 | n23900 ;
  assign n23902 = ~n2049 & n20879 ;
  assign n23903 = n23902 ^ n6093 ^ 1'b0 ;
  assign n23904 = n23903 ^ n13908 ^ n10487 ;
  assign n23905 = n19792 ^ n8504 ^ n2018 ;
  assign n23906 = n23905 ^ n9950 ^ n2445 ;
  assign n23907 = n8985 ^ n2592 ^ 1'b0 ;
  assign n23908 = n23906 & ~n23907 ;
  assign n23909 = n20184 ^ n4691 ^ 1'b0 ;
  assign n23910 = n183 & n23909 ;
  assign n23911 = n5104 | n11687 ;
  assign n23912 = n2876 | n23911 ;
  assign n23913 = n3529 & n14827 ;
  assign n23914 = ~n23912 & n23913 ;
  assign n23915 = n11693 ^ n4987 ^ 1'b0 ;
  assign n23916 = n537 & ~n23915 ;
  assign n23917 = n23916 ^ n23795 ^ n22467 ;
  assign n23918 = n3631 & ~n23917 ;
  assign n23919 = ~n646 & n9160 ;
  assign n23920 = n12271 ^ n11430 ^ n10210 ;
  assign n23921 = ( n2063 & ~n11684 ) | ( n2063 & n20462 ) | ( ~n11684 & n20462 ) ;
  assign n23922 = ( n4219 & n12217 ) | ( n4219 & n13004 ) | ( n12217 & n13004 ) ;
  assign n23923 = n315 | n23922 ;
  assign n23924 = n19221 & n23923 ;
  assign n23925 = n23924 ^ n4906 ^ 1'b0 ;
  assign n23926 = ( ~n12337 & n23921 ) | ( ~n12337 & n23925 ) | ( n23921 & n23925 ) ;
  assign n23928 = ~n4285 & n13737 ;
  assign n23929 = n23928 ^ n21787 ^ 1'b0 ;
  assign n23930 = ( n6489 & ~n22034 ) | ( n6489 & n23929 ) | ( ~n22034 & n23929 ) ;
  assign n23927 = n19518 ^ n11074 ^ 1'b0 ;
  assign n23931 = n23930 ^ n23927 ^ n1896 ;
  assign n23932 = n8503 ^ n835 ^ 1'b0 ;
  assign n23933 = n23931 & ~n23932 ;
  assign n23934 = n5595 & ~n8362 ;
  assign n23935 = n13705 | n22501 ;
  assign n23936 = n23934 | n23935 ;
  assign n23937 = n23933 & ~n23936 ;
  assign n23938 = n3909 & n23937 ;
  assign n23939 = n6762 ^ n5033 ^ 1'b0 ;
  assign n23940 = ~n6091 & n23939 ;
  assign n23941 = n17188 ^ n13781 ^ n4895 ;
  assign n23942 = ~n1020 & n23941 ;
  assign n23943 = n2147 ^ x86 ^ 1'b0 ;
  assign n23944 = ( ~n6094 & n8062 ) | ( ~n6094 & n8870 ) | ( n8062 & n8870 ) ;
  assign n23945 = ( n17704 & n22814 ) | ( n17704 & n23419 ) | ( n22814 & n23419 ) ;
  assign n23946 = n3469 & ~n16995 ;
  assign n23947 = n10907 ^ n2391 ^ 1'b0 ;
  assign n23948 = n3948 & n11258 ;
  assign n23949 = n23948 ^ n9647 ^ 1'b0 ;
  assign n23950 = x84 & n13128 ;
  assign n23951 = n23949 & n23950 ;
  assign n23952 = n9540 & ~n10823 ;
  assign n23953 = ( n9057 & ~n11586 ) | ( n9057 & n17126 ) | ( ~n11586 & n17126 ) ;
  assign n23954 = ( n4065 & n7278 ) | ( n4065 & ~n23953 ) | ( n7278 & ~n23953 ) ;
  assign n23955 = n23954 ^ n4711 ^ 1'b0 ;
  assign n23956 = ~n23952 & n23955 ;
  assign n23957 = n23956 ^ n20849 ^ 1'b0 ;
  assign n23958 = ~n6067 & n23957 ;
  assign n23959 = n23958 ^ n19618 ^ 1'b0 ;
  assign n23960 = ~n2312 & n5995 ;
  assign n23961 = n23960 ^ n1016 ^ 1'b0 ;
  assign n23962 = n21549 ^ n19885 ^ n2291 ;
  assign n23963 = n2562 | n5704 ;
  assign n23964 = n4344 | n23963 ;
  assign n23965 = n12321 & ~n23964 ;
  assign n23966 = n694 | n4339 ;
  assign n23967 = n23966 ^ n10534 ^ 1'b0 ;
  assign n23968 = ~n10782 & n14821 ;
  assign n23969 = n23968 ^ n3794 ^ n3738 ;
  assign n23970 = n9000 ^ n7840 ^ 1'b0 ;
  assign n23971 = n3194 & ~n23970 ;
  assign n23972 = n9232 | n18435 ;
  assign n23973 = n23971 | n23972 ;
  assign n23974 = n1184 | n9818 ;
  assign n23975 = n23974 ^ n5714 ^ 1'b0 ;
  assign n23976 = n8443 | n20721 ;
  assign n23977 = n23975 | n23976 ;
  assign n23978 = n16074 ^ n13571 ^ 1'b0 ;
  assign n23979 = n22052 ^ n17833 ^ 1'b0 ;
  assign n23980 = ( n3992 & n12358 ) | ( n3992 & ~n14312 ) | ( n12358 & ~n14312 ) ;
  assign n23981 = n23980 ^ n23797 ^ n4575 ;
  assign n23982 = n16876 ^ n10181 ^ 1'b0 ;
  assign n23983 = n23982 ^ n15582 ^ n670 ;
  assign n23987 = ( n14809 & ~n15496 ) | ( n14809 & n18480 ) | ( ~n15496 & n18480 ) ;
  assign n23984 = n9946 | n16837 ;
  assign n23985 = ~n11025 & n23984 ;
  assign n23986 = ~n16209 & n23985 ;
  assign n23988 = n23987 ^ n23986 ^ 1'b0 ;
  assign n23989 = n23988 ^ n5471 ^ 1'b0 ;
  assign n23990 = n20555 ^ n6748 ^ n6328 ;
  assign n23991 = n3510 & ~n23990 ;
  assign n23992 = n23991 ^ n2779 ^ n2420 ;
  assign n23993 = n23992 ^ n23250 ^ n659 ;
  assign n23994 = ~n4161 & n18137 ;
  assign n23995 = n3015 & n5595 ;
  assign n23996 = n23995 ^ n10993 ^ 1'b0 ;
  assign n23997 = ~n1917 & n20924 ;
  assign n23998 = n3414 & n23997 ;
  assign n23999 = n4716 & n11474 ;
  assign n24000 = n10617 & n23999 ;
  assign n24001 = n17604 ^ n7229 ^ 1'b0 ;
  assign n24002 = n9587 ^ n6221 ^ n1583 ;
  assign n24003 = n7733 & n24002 ;
  assign n24004 = n2513 & n24003 ;
  assign n24005 = ( n16957 & n23583 ) | ( n16957 & n24004 ) | ( n23583 & n24004 ) ;
  assign n24007 = n2638 | n5521 ;
  assign n24006 = n13441 & n22194 ;
  assign n24008 = n24007 ^ n24006 ^ n16121 ;
  assign n24009 = n15150 ^ n2658 ^ 1'b0 ;
  assign n24010 = n6819 | n18454 ;
  assign n24011 = n24010 ^ n16938 ^ 1'b0 ;
  assign n24012 = n3549 & n6605 ;
  assign n24013 = ~n19207 & n24012 ;
  assign n24014 = n16990 ^ n680 ^ 1'b0 ;
  assign n24015 = n24013 | n24014 ;
  assign n24016 = n16717 ^ n15024 ^ n4956 ;
  assign n24017 = n1817 & n24016 ;
  assign n24018 = n24017 ^ n21139 ^ 1'b0 ;
  assign n24019 = ~n5390 & n20091 ;
  assign n24020 = ~n15036 & n24019 ;
  assign n24021 = n24020 ^ n8303 ^ 1'b0 ;
  assign n24022 = ( n2121 & n6238 ) | ( n2121 & ~n20313 ) | ( n6238 & ~n20313 ) ;
  assign n24023 = n21708 ^ n18008 ^ n16970 ;
  assign n24024 = n6539 | n9076 ;
  assign n24025 = n24024 ^ n1225 ^ 1'b0 ;
  assign n24026 = ( ~n6469 & n18394 ) | ( ~n6469 & n23739 ) | ( n18394 & n23739 ) ;
  assign n24027 = ( ~n4366 & n24025 ) | ( ~n4366 & n24026 ) | ( n24025 & n24026 ) ;
  assign n24028 = ~n875 & n20196 ;
  assign n24030 = n996 & ~n4936 ;
  assign n24031 = n24030 ^ n275 ^ 1'b0 ;
  assign n24032 = ~n2339 & n24031 ;
  assign n24033 = n24032 ^ n7684 ^ n3402 ;
  assign n24029 = ( n7679 & n15437 ) | ( n7679 & n21610 ) | ( n15437 & n21610 ) ;
  assign n24034 = n24033 ^ n24029 ^ n10709 ;
  assign n24035 = n18534 ^ n14863 ^ n13785 ;
  assign n24036 = n18418 | n24035 ;
  assign n24037 = n24036 ^ n20800 ^ 1'b0 ;
  assign n24038 = ~n2331 & n15546 ;
  assign n24039 = ( n1038 & n7134 ) | ( n1038 & n9929 ) | ( n7134 & n9929 ) ;
  assign n24040 = ( ~n2632 & n3016 ) | ( ~n2632 & n24039 ) | ( n3016 & n24039 ) ;
  assign n24041 = ( n726 & n18156 ) | ( n726 & ~n20380 ) | ( n18156 & ~n20380 ) ;
  assign n24042 = ( n5728 & ~n6066 ) | ( n5728 & n14007 ) | ( ~n6066 & n14007 ) ;
  assign n24043 = ( n1628 & ~n6835 ) | ( n1628 & n17198 ) | ( ~n6835 & n17198 ) ;
  assign n24044 = n24043 ^ n13633 ^ 1'b0 ;
  assign n24045 = n21232 ^ n16013 ^ 1'b0 ;
  assign n24046 = n12157 & ~n24045 ;
  assign n24047 = ~n8125 & n10466 ;
  assign n24048 = ( n2220 & ~n11003 ) | ( n2220 & n24047 ) | ( ~n11003 & n24047 ) ;
  assign n24049 = n921 | n24048 ;
  assign n24050 = n24046 | n24049 ;
  assign n24053 = ~n2923 & n6041 ;
  assign n24054 = ( n5154 & ~n8937 ) | ( n5154 & n24053 ) | ( ~n8937 & n24053 ) ;
  assign n24051 = n6828 ^ n4307 ^ 1'b0 ;
  assign n24052 = n19792 & n24051 ;
  assign n24055 = n24054 ^ n24052 ^ n6596 ;
  assign n24056 = n19663 ^ n4997 ^ 1'b0 ;
  assign n24057 = ~n24055 & n24056 ;
  assign n24058 = n11975 & n23606 ;
  assign n24059 = ~n332 & n1316 ;
  assign n24060 = ~x27 & n24059 ;
  assign n24061 = n6316 ^ n4949 ^ x66 ;
  assign n24062 = n24060 & n24061 ;
  assign n24063 = ( n10184 & ~n13323 ) | ( n10184 & n17580 ) | ( ~n13323 & n17580 ) ;
  assign n24064 = ( n13776 & n24025 ) | ( n13776 & ~n24063 ) | ( n24025 & ~n24063 ) ;
  assign n24065 = n1011 & n2873 ;
  assign n24066 = n24065 ^ n13307 ^ 1'b0 ;
  assign n24067 = n24066 ^ n20394 ^ n313 ;
  assign n24068 = n6685 ^ n5695 ^ 1'b0 ;
  assign n24069 = n3776 & ~n24068 ;
  assign n24070 = n24069 ^ n22807 ^ n3376 ;
  assign n24071 = n11201 ^ n5527 ^ 1'b0 ;
  assign n24072 = ~n11943 & n16454 ;
  assign n24073 = n22244 ^ n1936 ^ 1'b0 ;
  assign n24074 = ~n13740 & n24073 ;
  assign n24075 = ( n21388 & ~n24072 ) | ( n21388 & n24074 ) | ( ~n24072 & n24074 ) ;
  assign n24076 = n1597 | n24075 ;
  assign n24077 = n4213 & ~n24076 ;
  assign n24078 = ( ~n5934 & n15314 ) | ( ~n5934 & n23329 ) | ( n15314 & n23329 ) ;
  assign n24079 = ( n3800 & n10897 ) | ( n3800 & n15641 ) | ( n10897 & n15641 ) ;
  assign n24080 = ( n2409 & ~n3656 ) | ( n2409 & n5195 ) | ( ~n3656 & n5195 ) ;
  assign n24081 = ( n1043 & n1886 ) | ( n1043 & n24080 ) | ( n1886 & n24080 ) ;
  assign n24082 = n5564 ^ n2811 ^ n911 ;
  assign n24083 = n21105 ^ n1588 ^ 1'b0 ;
  assign n24084 = n14580 ^ n6466 ^ n1659 ;
  assign n24085 = ( n1893 & n9359 ) | ( n1893 & n14185 ) | ( n9359 & n14185 ) ;
  assign n24086 = ( ~n11905 & n19717 ) | ( ~n11905 & n24085 ) | ( n19717 & n24085 ) ;
  assign n24087 = n24086 ^ n9435 ^ 1'b0 ;
  assign n24088 = x45 & n24087 ;
  assign n24089 = n18604 ^ n2027 ^ 1'b0 ;
  assign n24090 = n21991 ^ n10049 ^ 1'b0 ;
  assign n24091 = ( n8728 & n10268 ) | ( n8728 & ~n10277 ) | ( n10268 & ~n10277 ) ;
  assign n24093 = n20625 ^ n15699 ^ 1'b0 ;
  assign n24092 = n12794 ^ n7383 ^ 1'b0 ;
  assign n24094 = n24093 ^ n24092 ^ n3813 ;
  assign n24095 = n19631 ^ n8689 ^ 1'b0 ;
  assign n24096 = ( n6328 & n12465 ) | ( n6328 & ~n24095 ) | ( n12465 & ~n24095 ) ;
  assign n24097 = n21708 & n24096 ;
  assign n24098 = ( ~n3539 & n8426 ) | ( ~n3539 & n10501 ) | ( n8426 & n10501 ) ;
  assign n24099 = n24098 ^ n10452 ^ n3640 ;
  assign n24100 = ( n839 & n1179 ) | ( n839 & ~n23948 ) | ( n1179 & ~n23948 ) ;
  assign n24101 = n24100 ^ n19090 ^ 1'b0 ;
  assign n24102 = n24099 & n24101 ;
  assign n24103 = ~n3530 & n12777 ;
  assign n24104 = ~n21228 & n24103 ;
  assign n24105 = n12032 ^ n8166 ^ 1'b0 ;
  assign n24106 = n20748 & ~n24105 ;
  assign n24109 = n3157 & n12592 ;
  assign n24110 = ~n7224 & n24109 ;
  assign n24107 = n7875 ^ n203 ^ 1'b0 ;
  assign n24108 = ~n19609 & n24107 ;
  assign n24111 = n24110 ^ n24108 ^ n16301 ;
  assign n24112 = n14423 ^ n3673 ^ 1'b0 ;
  assign n24113 = ~n170 & n24112 ;
  assign n24114 = n24113 ^ n19130 ^ n15752 ;
  assign n24115 = ( n1066 & n7644 ) | ( n1066 & ~n12962 ) | ( n7644 & ~n12962 ) ;
  assign n24116 = n20110 ^ n12333 ^ 1'b0 ;
  assign n24117 = n9341 | n24116 ;
  assign n24118 = n2652 & n8003 ;
  assign n24119 = n24118 ^ n1061 ^ 1'b0 ;
  assign n24120 = ( n2776 & ~n6338 ) | ( n2776 & n13026 ) | ( ~n6338 & n13026 ) ;
  assign n24121 = n24119 & ~n24120 ;
  assign n24122 = ( n876 & n1903 ) | ( n876 & n6603 ) | ( n1903 & n6603 ) ;
  assign n24124 = n7753 ^ n5759 ^ 1'b0 ;
  assign n24123 = n23328 ^ n1896 ^ 1'b0 ;
  assign n24125 = n24124 ^ n24123 ^ n2696 ;
  assign n24126 = n23081 & n23477 ;
  assign n24127 = ~n7490 & n10770 ;
  assign n24128 = ~n5042 & n6505 ;
  assign n24129 = n24128 ^ n1671 ^ 1'b0 ;
  assign n24130 = n24129 ^ n16515 ^ n3278 ;
  assign n24131 = ( ~n18198 & n24127 ) | ( ~n18198 & n24130 ) | ( n24127 & n24130 ) ;
  assign n24132 = ~n1687 & n22056 ;
  assign n24133 = n4250 ^ n2367 ^ 1'b0 ;
  assign n24134 = n10924 | n24133 ;
  assign n24135 = n19711 ^ n1315 ^ 1'b0 ;
  assign n24136 = n17386 ^ n9123 ^ n3028 ;
  assign n24137 = n9255 ^ n6671 ^ n273 ;
  assign n24140 = ( ~n1663 & n6403 ) | ( ~n1663 & n18288 ) | ( n6403 & n18288 ) ;
  assign n24138 = n17078 & n19083 ;
  assign n24139 = n24138 ^ n14249 ^ 1'b0 ;
  assign n24141 = n24140 ^ n24139 ^ 1'b0 ;
  assign n24142 = ( ~n2487 & n24137 ) | ( ~n2487 & n24141 ) | ( n24137 & n24141 ) ;
  assign n24147 = ( n3212 & ~n5105 ) | ( n3212 & n17329 ) | ( ~n5105 & n17329 ) ;
  assign n24145 = n20157 ^ n8276 ^ 1'b0 ;
  assign n24143 = ~n4567 & n15281 ;
  assign n24144 = n23171 & n24143 ;
  assign n24146 = n24145 ^ n24144 ^ 1'b0 ;
  assign n24148 = n24147 ^ n24146 ^ n23562 ;
  assign n24149 = n5164 & ~n17772 ;
  assign n24155 = n6826 & n7193 ;
  assign n24156 = n12895 & n24155 ;
  assign n24157 = n24156 ^ n9151 ^ n5916 ;
  assign n24150 = n8450 ^ n1809 ^ 1'b0 ;
  assign n24151 = n11004 | n24150 ;
  assign n24152 = n24151 ^ n12483 ^ 1'b0 ;
  assign n24153 = ~n11033 & n24152 ;
  assign n24154 = ( n4982 & n12152 ) | ( n4982 & n24153 ) | ( n12152 & n24153 ) ;
  assign n24158 = n24157 ^ n24154 ^ n8035 ;
  assign n24159 = n3847 & ~n19112 ;
  assign n24160 = n5127 & n24159 ;
  assign n24161 = ( n3153 & n13648 ) | ( n3153 & n14045 ) | ( n13648 & n14045 ) ;
  assign n24162 = n10270 | n24161 ;
  assign n24163 = n12239 | n24162 ;
  assign n24164 = ( n10636 & n21414 ) | ( n10636 & ~n24163 ) | ( n21414 & ~n24163 ) ;
  assign n24165 = n23613 | n24164 ;
  assign n24166 = n10769 ^ n6079 ^ n2052 ;
  assign n24167 = ( ~n11159 & n11374 ) | ( ~n11159 & n19266 ) | ( n11374 & n19266 ) ;
  assign n24168 = ( n5457 & n7655 ) | ( n5457 & n24167 ) | ( n7655 & n24167 ) ;
  assign n24169 = ~n4318 & n9094 ;
  assign n24170 = n2871 & ~n24169 ;
  assign n24171 = n7743 | n15501 ;
  assign n24172 = ( ~n6548 & n23422 ) | ( ~n6548 & n24171 ) | ( n23422 & n24171 ) ;
  assign n24173 = n3755 | n24172 ;
  assign n24174 = n24170 | n24173 ;
  assign n24175 = n6636 & ~n22261 ;
  assign n24176 = n16552 ^ n11471 ^ n11381 ;
  assign n24177 = ~n15097 & n24176 ;
  assign n24178 = n12443 ^ n9306 ^ 1'b0 ;
  assign n24179 = n13509 ^ n332 ^ 1'b0 ;
  assign n24180 = ( n21023 & n24178 ) | ( n21023 & ~n24179 ) | ( n24178 & ~n24179 ) ;
  assign n24181 = n12006 ^ n7642 ^ n6142 ;
  assign n24182 = n9165 ^ n7314 ^ n1460 ;
  assign n24183 = n24182 ^ n2370 ^ 1'b0 ;
  assign n24184 = n23233 ^ n13002 ^ n10184 ;
  assign n24185 = n8422 ^ n7871 ^ n3709 ;
  assign n24186 = ( n10534 & n21213 ) | ( n10534 & ~n24185 ) | ( n21213 & ~n24185 ) ;
  assign n24187 = n489 & n14542 ;
  assign n24188 = ~n4236 & n6613 ;
  assign n24189 = n24188 ^ n7507 ^ 1'b0 ;
  assign n24190 = n5782 & ~n24189 ;
  assign n24191 = ~n11505 & n24190 ;
  assign n24192 = n2607 ^ n563 ^ 1'b0 ;
  assign n24193 = n13134 & n24192 ;
  assign n24196 = ( ~n694 & n8687 ) | ( ~n694 & n11898 ) | ( n8687 & n11898 ) ;
  assign n24194 = n17876 ^ n2819 ^ 1'b0 ;
  assign n24195 = n20878 & ~n24194 ;
  assign n24197 = n24196 ^ n24195 ^ n5474 ;
  assign n24198 = n5815 ^ n2857 ^ 1'b0 ;
  assign n24199 = n11020 | n20188 ;
  assign n24200 = n24198 & ~n24199 ;
  assign n24201 = n24200 ^ n14567 ^ 1'b0 ;
  assign n24202 = n6016 ^ n4040 ^ n556 ;
  assign n24203 = n22250 ^ n14674 ^ 1'b0 ;
  assign n24205 = n8718 ^ n615 ^ 1'b0 ;
  assign n24204 = n3883 | n21189 ;
  assign n24206 = n24205 ^ n24204 ^ 1'b0 ;
  assign n24207 = ( n2352 & n9318 ) | ( n2352 & n16386 ) | ( n9318 & n16386 ) ;
  assign n24208 = n24207 ^ n9832 ^ n4543 ;
  assign n24209 = n17075 ^ n7741 ^ n3377 ;
  assign n24210 = ( ~n4496 & n21011 ) | ( ~n4496 & n24209 ) | ( n21011 & n24209 ) ;
  assign n24211 = ( n1940 & n2511 ) | ( n1940 & ~n24210 ) | ( n2511 & ~n24210 ) ;
  assign n24212 = n15722 | n19443 ;
  assign n24213 = n6665 | n8737 ;
  assign n24214 = n11790 | n24213 ;
  assign n24215 = n3776 & n4717 ;
  assign n24218 = n7330 & n14142 ;
  assign n24219 = n9765 & n24218 ;
  assign n24216 = n828 | n10588 ;
  assign n24217 = n21736 & ~n24216 ;
  assign n24220 = n24219 ^ n24217 ^ n7837 ;
  assign n24221 = ( n199 & ~n2093 ) | ( n199 & n2700 ) | ( ~n2093 & n2700 ) ;
  assign n24222 = ( n6496 & ~n11158 ) | ( n6496 & n24221 ) | ( ~n11158 & n24221 ) ;
  assign n24223 = ( n2369 & n5286 ) | ( n2369 & ~n10753 ) | ( n5286 & ~n10753 ) ;
  assign n24224 = n24223 ^ n12043 ^ n7602 ;
  assign n24225 = n3676 ^ n1441 ^ 1'b0 ;
  assign n24226 = n19880 & n24225 ;
  assign n24227 = n9320 ^ n3934 ^ 1'b0 ;
  assign n24228 = ~n10507 & n24227 ;
  assign n24230 = ( n4101 & n7843 ) | ( n4101 & n12543 ) | ( n7843 & n12543 ) ;
  assign n24229 = n2982 | n8426 ;
  assign n24231 = n24230 ^ n24229 ^ 1'b0 ;
  assign n24233 = n23174 ^ n12738 ^ n8054 ;
  assign n24232 = n182 & n15592 ;
  assign n24234 = n24233 ^ n24232 ^ 1'b0 ;
  assign n24235 = ~n13966 & n16603 ;
  assign n24236 = n24235 ^ n1618 ^ 1'b0 ;
  assign n24237 = n20074 & n24236 ;
  assign n24238 = n20940 ^ n8448 ^ n3821 ;
  assign n24239 = ( ~n3453 & n20099 ) | ( ~n3453 & n24238 ) | ( n20099 & n24238 ) ;
  assign n24241 = n11545 & ~n11851 ;
  assign n24240 = n520 ^ n153 ^ 1'b0 ;
  assign n24242 = n24241 ^ n24240 ^ n9098 ;
  assign n24243 = n326 | n1595 ;
  assign n24244 = n16385 ^ n15809 ^ n8570 ;
  assign n24245 = n7382 & ~n24244 ;
  assign n24246 = n2756 ^ n1038 ^ 1'b0 ;
  assign n24247 = n18207 | n24246 ;
  assign n24248 = n24247 ^ n15776 ^ n3405 ;
  assign n24249 = ( ~n15292 & n24245 ) | ( ~n15292 & n24248 ) | ( n24245 & n24248 ) ;
  assign n24250 = n24249 ^ n14279 ^ n897 ;
  assign n24251 = n2435 & n20509 ;
  assign n24252 = ~n13423 & n24251 ;
  assign n24253 = ( n469 & n11112 ) | ( n469 & n12433 ) | ( n11112 & n12433 ) ;
  assign n24254 = n13980 ^ n1555 ^ 1'b0 ;
  assign n24255 = ~n24253 & n24254 ;
  assign n24256 = ( ~n12891 & n16680 ) | ( ~n12891 & n24255 ) | ( n16680 & n24255 ) ;
  assign n24257 = n12530 ^ n1704 ^ 1'b0 ;
  assign n24258 = n24256 & n24257 ;
  assign n24259 = n3292 & n16854 ;
  assign n24260 = ~n3303 & n24259 ;
  assign n24261 = n562 | n24260 ;
  assign n24262 = n24261 ^ n11773 ^ n10078 ;
  assign n24263 = n8453 ^ n971 ^ 1'b0 ;
  assign n24264 = ( n9252 & ~n10096 ) | ( n9252 & n24263 ) | ( ~n10096 & n24263 ) ;
  assign n24265 = n24264 ^ n14749 ^ 1'b0 ;
  assign n24266 = ~n12618 & n24265 ;
  assign n24267 = n6663 & ~n15449 ;
  assign n24268 = ~n9377 & n24267 ;
  assign n24269 = ( ~n13505 & n14387 ) | ( ~n13505 & n24268 ) | ( n14387 & n24268 ) ;
  assign n24270 = n21860 & n24269 ;
  assign n24271 = n6503 ^ n6084 ^ 1'b0 ;
  assign n24272 = n24271 ^ n8203 ^ n183 ;
  assign n24273 = n7311 ^ n2791 ^ 1'b0 ;
  assign n24274 = n13049 | n24273 ;
  assign n24275 = ~n3464 & n24274 ;
  assign n24276 = n13839 & n24275 ;
  assign n24277 = n16325 ^ n6113 ^ n3277 ;
  assign n24278 = ( n7266 & n22187 ) | ( n7266 & n24264 ) | ( n22187 & n24264 ) ;
  assign n24279 = n8537 ^ n6561 ^ n2154 ;
  assign n24280 = n8843 ^ n6776 ^ 1'b0 ;
  assign n24281 = n1554 & ~n24280 ;
  assign n24282 = ~n1711 & n24281 ;
  assign n24283 = ~n24279 & n24282 ;
  assign n24284 = ( n6494 & n14915 ) | ( n6494 & ~n24283 ) | ( n14915 & ~n24283 ) ;
  assign n24285 = n3536 & n4685 ;
  assign n24286 = n6585 & n24285 ;
  assign n24287 = n19460 ^ n15770 ^ 1'b0 ;
  assign n24288 = n19517 & n24287 ;
  assign n24289 = n7456 & ~n14615 ;
  assign n24290 = ( n5969 & n15085 ) | ( n5969 & ~n24289 ) | ( n15085 & ~n24289 ) ;
  assign n24291 = n24290 ^ n14755 ^ 1'b0 ;
  assign n24292 = ~n22091 & n24291 ;
  assign n24293 = n13018 ^ n2445 ^ 1'b0 ;
  assign n24294 = n24292 & ~n24293 ;
  assign n24295 = n1177 | n7647 ;
  assign n24296 = n2090 & ~n6070 ;
  assign n24297 = n24296 ^ n11693 ^ n6632 ;
  assign n24298 = n21642 ^ n12580 ^ n12513 ;
  assign n24299 = ( ~n6877 & n15530 ) | ( ~n6877 & n24298 ) | ( n15530 & n24298 ) ;
  assign n24301 = n4722 & n10501 ;
  assign n24300 = ( n4221 & n6795 ) | ( n4221 & n12005 ) | ( n6795 & n12005 ) ;
  assign n24302 = n24301 ^ n24300 ^ n15352 ;
  assign n24303 = ( n323 & n8232 ) | ( n323 & n14795 ) | ( n8232 & n14795 ) ;
  assign n24304 = n24303 ^ n13719 ^ n7951 ;
  assign n24305 = ( ~n297 & n19519 ) | ( ~n297 & n20945 ) | ( n19519 & n20945 ) ;
  assign n24306 = n24305 ^ n7481 ^ n1455 ;
  assign n24307 = n907 | n5198 ;
  assign n24308 = n24307 ^ n2395 ^ 1'b0 ;
  assign n24309 = n4161 | n18411 ;
  assign n24310 = n24309 ^ n13026 ^ 1'b0 ;
  assign n24311 = n21737 ^ n7000 ^ 1'b0 ;
  assign n24312 = ~n15524 & n24311 ;
  assign n24313 = n1716 | n7083 ;
  assign n24314 = n14684 | n24313 ;
  assign n24318 = ( ~n2496 & n4910 ) | ( ~n2496 & n5158 ) | ( n4910 & n5158 ) ;
  assign n24315 = ~n2146 & n4751 ;
  assign n24316 = n5195 & n24315 ;
  assign n24317 = n17929 & n24316 ;
  assign n24319 = n24318 ^ n24317 ^ n17134 ;
  assign n24320 = n2886 & ~n8348 ;
  assign n24321 = n5388 & n24320 ;
  assign n24322 = ( n11543 & n14316 ) | ( n11543 & n24321 ) | ( n14316 & n24321 ) ;
  assign n24323 = ( n2709 & n3166 ) | ( n2709 & n6636 ) | ( n3166 & n6636 ) ;
  assign n24324 = ( n5156 & ~n24322 ) | ( n5156 & n24323 ) | ( ~n24322 & n24323 ) ;
  assign n24325 = n12986 ^ n7718 ^ 1'b0 ;
  assign n24326 = n7322 | n24325 ;
  assign n24327 = n24326 ^ n20844 ^ n3016 ;
  assign n24328 = n697 & ~n24327 ;
  assign n24329 = n24328 ^ n8094 ^ 1'b0 ;
  assign n24330 = ( ~n9043 & n9835 ) | ( ~n9043 & n13304 ) | ( n9835 & n13304 ) ;
  assign n24331 = n24330 ^ n22934 ^ n12677 ;
  assign n24332 = ( n12418 & ~n13974 ) | ( n12418 & n24331 ) | ( ~n13974 & n24331 ) ;
  assign n24333 = n24332 ^ n23984 ^ 1'b0 ;
  assign n24334 = n14964 & n24333 ;
  assign n24335 = n22232 ^ n19726 ^ 1'b0 ;
  assign n24336 = ( n7525 & ~n9325 ) | ( n7525 & n11290 ) | ( ~n9325 & n11290 ) ;
  assign n24337 = ( n8844 & n21936 ) | ( n8844 & n24336 ) | ( n21936 & n24336 ) ;
  assign n24338 = n11474 ^ n3476 ^ x100 ;
  assign n24339 = ( n9792 & ~n15486 ) | ( n9792 & n18436 ) | ( ~n15486 & n18436 ) ;
  assign n24340 = ( ~n872 & n14101 ) | ( ~n872 & n24339 ) | ( n14101 & n24339 ) ;
  assign n24342 = n9836 ^ n3320 ^ n1002 ;
  assign n24341 = ~n8593 & n21729 ;
  assign n24343 = n24342 ^ n24341 ^ 1'b0 ;
  assign n24344 = n23144 ^ n14585 ^ 1'b0 ;
  assign n24345 = n17494 ^ n7949 ^ n7836 ;
  assign n24346 = n20845 | n24345 ;
  assign n24347 = n9104 & ~n24346 ;
  assign n24348 = n13969 ^ n2491 ^ 1'b0 ;
  assign n24349 = n15706 ^ n10077 ^ n248 ;
  assign n24352 = n3086 ^ n1613 ^ 1'b0 ;
  assign n24353 = ~n345 & n24352 ;
  assign n24350 = n24030 ^ n3978 ^ 1'b0 ;
  assign n24351 = n8624 & n24350 ;
  assign n24354 = n24353 ^ n24351 ^ n6739 ;
  assign n24355 = n24354 ^ n11552 ^ n9358 ;
  assign n24357 = n4974 | n23053 ;
  assign n24356 = n15039 ^ n3762 ^ n2592 ;
  assign n24358 = n24357 ^ n24356 ^ n23174 ;
  assign n24359 = ( ~n3115 & n4403 ) | ( ~n3115 & n4537 ) | ( n4403 & n4537 ) ;
  assign n24360 = n24359 ^ n13678 ^ n9104 ;
  assign n24361 = ( n8156 & ~n21108 ) | ( n8156 & n24360 ) | ( ~n21108 & n24360 ) ;
  assign n24370 = ~n6353 & n13327 ;
  assign n24362 = ~n4016 & n7685 ;
  assign n24363 = n24362 ^ n19511 ^ 1'b0 ;
  assign n24364 = n559 & n15756 ;
  assign n24365 = n24364 ^ n5453 ^ 1'b0 ;
  assign n24366 = ~n9491 & n24365 ;
  assign n24367 = n24366 ^ n12559 ^ 1'b0 ;
  assign n24368 = ( ~n10813 & n24363 ) | ( ~n10813 & n24367 ) | ( n24363 & n24367 ) ;
  assign n24369 = ~n5436 & n24368 ;
  assign n24371 = n24370 ^ n24369 ^ 1'b0 ;
  assign n24372 = ( n2881 & n24361 ) | ( n2881 & ~n24371 ) | ( n24361 & ~n24371 ) ;
  assign n24373 = n1858 & ~n11892 ;
  assign n24374 = n24373 ^ n23216 ^ 1'b0 ;
  assign n24375 = n24374 ^ n12352 ^ 1'b0 ;
  assign n24376 = n7378 ^ n3697 ^ n1828 ;
  assign n24377 = n24376 ^ n6577 ^ 1'b0 ;
  assign n24378 = n21822 & n24377 ;
  assign n24379 = ~n10911 & n24378 ;
  assign n24380 = n11292 ^ n583 ^ 1'b0 ;
  assign n24381 = n14561 ^ n8631 ^ 1'b0 ;
  assign n24382 = n2488 | n24381 ;
  assign n24384 = ( n2286 & ~n5745 ) | ( n2286 & n14788 ) | ( ~n5745 & n14788 ) ;
  assign n24385 = ( n1418 & n6867 ) | ( n1418 & n24384 ) | ( n6867 & n24384 ) ;
  assign n24383 = ~n3118 & n18279 ;
  assign n24386 = n24385 ^ n24383 ^ 1'b0 ;
  assign n24387 = n24386 ^ n10774 ^ 1'b0 ;
  assign n24388 = n10780 & ~n24387 ;
  assign n24389 = n3487 ^ n1320 ^ 1'b0 ;
  assign n24390 = ( n4181 & n9382 ) | ( n4181 & n24389 ) | ( n9382 & n24389 ) ;
  assign n24391 = n24390 ^ n17791 ^ 1'b0 ;
  assign n24392 = n24388 & ~n24391 ;
  assign n24393 = ( n302 & n5918 ) | ( n302 & n14973 ) | ( n5918 & n14973 ) ;
  assign n24394 = ( n3756 & n7265 ) | ( n3756 & n16385 ) | ( n7265 & n16385 ) ;
  assign n24395 = n19511 ^ n13994 ^ 1'b0 ;
  assign n24396 = ~n24394 & n24395 ;
  assign n24397 = n24396 ^ n13493 ^ n2347 ;
  assign n24398 = ~n4621 & n5645 ;
  assign n24399 = n24398 ^ n11646 ^ 1'b0 ;
  assign n24400 = ( n9061 & ~n20159 ) | ( n9061 & n24399 ) | ( ~n20159 & n24399 ) ;
  assign n24401 = n24400 ^ n3441 ^ 1'b0 ;
  assign n24402 = n14334 & ~n19442 ;
  assign n24403 = n12410 | n19223 ;
  assign n24404 = n10594 | n24403 ;
  assign n24405 = n11821 ^ n7722 ^ 1'b0 ;
  assign n24406 = n10319 & n15521 ;
  assign n24407 = ~n24405 & n24406 ;
  assign n24408 = ( ~n5792 & n12626 ) | ( ~n5792 & n24407 ) | ( n12626 & n24407 ) ;
  assign n24409 = n23522 ^ n15350 ^ 1'b0 ;
  assign n24410 = n180 | n21414 ;
  assign n24411 = n24410 ^ n5951 ^ n3696 ;
  assign n24412 = ( n10472 & ~n11790 ) | ( n10472 & n15384 ) | ( ~n11790 & n15384 ) ;
  assign n24415 = ~n13273 & n15244 ;
  assign n24413 = ( n3173 & n6462 ) | ( n3173 & n10031 ) | ( n6462 & n10031 ) ;
  assign n24414 = n24413 ^ n18063 ^ n11945 ;
  assign n24416 = n24415 ^ n24414 ^ 1'b0 ;
  assign n24417 = ( ~n1647 & n6021 ) | ( ~n1647 & n23304 ) | ( n6021 & n23304 ) ;
  assign n24418 = ( n2087 & ~n3077 ) | ( n2087 & n14200 ) | ( ~n3077 & n14200 ) ;
  assign n24419 = n6663 & ~n10924 ;
  assign n24420 = n24418 & n24419 ;
  assign n24421 = n3480 | n11414 ;
  assign n24422 = n24421 ^ n9324 ^ 1'b0 ;
  assign n24423 = n20005 ^ n3592 ^ 1'b0 ;
  assign n24424 = ~n22705 & n24423 ;
  assign n24425 = n24422 & n24424 ;
  assign n24426 = n24425 ^ n14953 ^ 1'b0 ;
  assign n24427 = n3517 | n15533 ;
  assign n24428 = n16832 & ~n24427 ;
  assign n24429 = n3537 & ~n11162 ;
  assign n24430 = n3551 & n12109 ;
  assign n24431 = n22460 ^ n20322 ^ n643 ;
  assign n24433 = n6084 & n12859 ;
  assign n24434 = ( n1025 & n6695 ) | ( n1025 & n17496 ) | ( n6695 & n17496 ) ;
  assign n24435 = n24433 & ~n24434 ;
  assign n24436 = n24435 ^ n10020 ^ 1'b0 ;
  assign n24437 = ( n5974 & n8052 ) | ( n5974 & n24436 ) | ( n8052 & n24436 ) ;
  assign n24438 = n24437 ^ n24061 ^ n22536 ;
  assign n24432 = ( ~n6766 & n8442 ) | ( ~n6766 & n13560 ) | ( n8442 & n13560 ) ;
  assign n24439 = n24438 ^ n24432 ^ n4231 ;
  assign n24440 = ( n863 & ~n6900 ) | ( n863 & n8023 ) | ( ~n6900 & n8023 ) ;
  assign n24441 = ( n4568 & n7687 ) | ( n4568 & ~n24440 ) | ( n7687 & ~n24440 ) ;
  assign n24442 = n15411 ^ n10909 ^ n8148 ;
  assign n24443 = n9451 ^ n2865 ^ 1'b0 ;
  assign n24444 = n24442 | n24443 ;
  assign n24445 = n24441 | n24444 ;
  assign n24446 = n16699 ^ n9249 ^ n5716 ;
  assign n24447 = n24446 ^ n1005 ^ 1'b0 ;
  assign n24448 = n13648 | n24447 ;
  assign n24449 = n17401 ^ n6635 ^ 1'b0 ;
  assign n24450 = n11475 | n24449 ;
  assign n24451 = n14017 | n21432 ;
  assign n24452 = n24450 & ~n24451 ;
  assign n24453 = n4888 ^ n4191 ^ 1'b0 ;
  assign n24454 = ~n2596 & n24453 ;
  assign n24455 = n9587 ^ n6958 ^ n2598 ;
  assign n24456 = ~n24454 & n24455 ;
  assign n24458 = ( n7128 & n13394 ) | ( n7128 & n14953 ) | ( n13394 & n14953 ) ;
  assign n24459 = ( n1494 & ~n2609 ) | ( n1494 & n24458 ) | ( ~n2609 & n24458 ) ;
  assign n24460 = ( n5604 & ~n11505 ) | ( n5604 & n24459 ) | ( ~n11505 & n24459 ) ;
  assign n24457 = n20817 ^ n2137 ^ n1356 ;
  assign n24461 = n24460 ^ n24457 ^ 1'b0 ;
  assign n24466 = n20755 & n24384 ;
  assign n24467 = n24466 ^ n8689 ^ n4365 ;
  assign n24462 = n927 & ~n5198 ;
  assign n24463 = n24462 ^ n3160 ^ 1'b0 ;
  assign n24464 = n289 & n24463 ;
  assign n24465 = ~n3269 & n24464 ;
  assign n24468 = n24467 ^ n24465 ^ n22488 ;
  assign n24469 = ( ~n7195 & n12932 ) | ( ~n7195 & n24468 ) | ( n12932 & n24468 ) ;
  assign n24471 = n24039 ^ n9809 ^ n2593 ;
  assign n24470 = ( n1260 & ~n4416 ) | ( n1260 & n15901 ) | ( ~n4416 & n15901 ) ;
  assign n24472 = n24471 ^ n24470 ^ n15620 ;
  assign n24473 = n22977 ^ n19403 ^ n3209 ;
  assign n24474 = ~n19789 & n24473 ;
  assign n24475 = ~n8988 & n24474 ;
  assign n24476 = ( n1163 & n4002 ) | ( n1163 & ~n24475 ) | ( n4002 & ~n24475 ) ;
  assign n24477 = n3858 & ~n9941 ;
  assign n24478 = n17267 ^ n9593 ^ n4345 ;
  assign n24479 = n15170 & ~n24478 ;
  assign n24480 = ( n24122 & n24477 ) | ( n24122 & ~n24479 ) | ( n24477 & ~n24479 ) ;
  assign n24481 = ( ~n10879 & n12038 ) | ( ~n10879 & n12337 ) | ( n12038 & n12337 ) ;
  assign n24482 = n6790 & n7227 ;
  assign n24483 = n24481 & n24482 ;
  assign n24484 = n2640 | n23216 ;
  assign n24485 = n24484 ^ n849 ^ 1'b0 ;
  assign n24486 = n13890 ^ n7388 ^ n6238 ;
  assign n24487 = ~n24485 & n24486 ;
  assign n24488 = n7583 ^ n4139 ^ n1382 ;
  assign n24489 = ~n7350 & n11432 ;
  assign n24490 = n24488 & n24489 ;
  assign n24491 = n1806 & ~n12308 ;
  assign n24492 = n24491 ^ n7410 ^ 1'b0 ;
  assign n24493 = n2656 & n15127 ;
  assign n24494 = n4639 & n24493 ;
  assign n24495 = n24494 ^ n22870 ^ 1'b0 ;
  assign n24496 = n2023 & ~n2089 ;
  assign n24497 = ~n8643 & n15807 ;
  assign n24498 = ( ~n11586 & n24496 ) | ( ~n11586 & n24497 ) | ( n24496 & n24497 ) ;
  assign n24499 = ( ~n3187 & n5111 ) | ( ~n3187 & n7876 ) | ( n5111 & n7876 ) ;
  assign n24500 = ( n16957 & n20573 ) | ( n16957 & ~n24499 ) | ( n20573 & ~n24499 ) ;
  assign n24502 = n16110 ^ n9479 ^ n4356 ;
  assign n24501 = n14412 ^ n2757 ^ n495 ;
  assign n24503 = n24502 ^ n24501 ^ n12714 ;
  assign n24505 = n10689 | n13139 ;
  assign n24506 = n8822 & ~n24505 ;
  assign n24504 = ( n2934 & ~n3058 ) | ( n2934 & n3199 ) | ( ~n3058 & n3199 ) ;
  assign n24507 = n24506 ^ n24504 ^ n3724 ;
  assign n24508 = ~n3537 & n24507 ;
  assign n24509 = n17219 ^ n14235 ^ 1'b0 ;
  assign n24510 = ~n1295 & n7008 ;
  assign n24511 = n24510 ^ n2880 ^ 1'b0 ;
  assign n24512 = n916 & ~n24511 ;
  assign n24513 = n2948 ^ n1867 ^ 1'b0 ;
  assign n24514 = ~n24512 & n24513 ;
  assign n24515 = n11941 ^ n11500 ^ n1170 ;
  assign n24516 = ~n12300 & n24515 ;
  assign n24517 = n24516 ^ n24353 ^ 1'b0 ;
  assign n24518 = n4835 & ~n24517 ;
  assign n24519 = n24518 ^ n1282 ^ 1'b0 ;
  assign n24520 = n17692 ^ n6819 ^ n4923 ;
  assign n24521 = n7511 & n16415 ;
  assign n24522 = ~n24520 & n24521 ;
  assign n24523 = n12553 ^ n10826 ^ 1'b0 ;
  assign n24524 = n6381 & ~n24523 ;
  assign n24525 = n24524 ^ n12637 ^ n197 ;
  assign n24526 = n24525 ^ n1177 ^ 1'b0 ;
  assign n24527 = n24522 | n24526 ;
  assign n24528 = n24527 ^ n8751 ^ n2103 ;
  assign n24529 = ( n6870 & ~n11024 ) | ( n6870 & n15459 ) | ( ~n11024 & n15459 ) ;
  assign n24535 = n8024 ^ n1919 ^ n1036 ;
  assign n24530 = ~n17365 & n17396 ;
  assign n24531 = n24530 ^ n1486 ^ 1'b0 ;
  assign n24532 = n23590 ^ n11168 ^ 1'b0 ;
  assign n24533 = n24531 & n24532 ;
  assign n24534 = n24533 ^ n1738 ^ 1'b0 ;
  assign n24536 = n24535 ^ n24534 ^ x9 ;
  assign n24537 = n17110 ^ n11160 ^ n3794 ;
  assign n24538 = n19060 | n24537 ;
  assign n24539 = n5805 & ~n24538 ;
  assign n24540 = n24539 ^ n23668 ^ n16695 ;
  assign n24541 = n20282 ^ n5853 ^ n2112 ;
  assign n24542 = n4981 & ~n24541 ;
  assign n24543 = n13095 ^ n10067 ^ 1'b0 ;
  assign n24544 = n12072 ^ n3371 ^ 1'b0 ;
  assign n24545 = n950 | n24544 ;
  assign n24546 = n24545 ^ n8718 ^ n5708 ;
  assign n24548 = n1872 & n7566 ;
  assign n24549 = ~n22510 & n24548 ;
  assign n24550 = n21803 & n24549 ;
  assign n24547 = n8372 & ~n10568 ;
  assign n24551 = n24550 ^ n24547 ^ 1'b0 ;
  assign n24552 = ~n999 & n24551 ;
  assign n24553 = n181 & ~n657 ;
  assign n24554 = n24553 ^ n24060 ^ 1'b0 ;
  assign n24555 = ( n954 & n16653 ) | ( n954 & ~n24554 ) | ( n16653 & ~n24554 ) ;
  assign n24556 = n24555 ^ n12592 ^ n9305 ;
  assign n24557 = ( ~n3879 & n20446 ) | ( ~n3879 & n24556 ) | ( n20446 & n24556 ) ;
  assign n24558 = ( n605 & n8784 ) | ( n605 & ~n20439 ) | ( n8784 & ~n20439 ) ;
  assign n24559 = n9622 ^ n1118 ^ 1'b0 ;
  assign n24560 = n24559 ^ n11759 ^ 1'b0 ;
  assign n24561 = ( n6568 & n7754 ) | ( n6568 & n14654 ) | ( n7754 & n14654 ) ;
  assign n24562 = n12911 | n24561 ;
  assign n24563 = n24560 | n24562 ;
  assign n24564 = n24563 ^ n17251 ^ n4528 ;
  assign n24565 = ~n11019 & n20798 ;
  assign n24566 = n24271 ^ n6546 ^ 1'b0 ;
  assign n24567 = n9124 | n24566 ;
  assign n24568 = n24567 ^ n20561 ^ n7082 ;
  assign n24569 = n24568 ^ n2335 ^ 1'b0 ;
  assign n24570 = n7750 ^ n3218 ^ n1784 ;
  assign n24571 = n24570 ^ n2646 ^ 1'b0 ;
  assign n24572 = n11382 ^ n5062 ^ 1'b0 ;
  assign n24573 = n24571 & n24572 ;
  assign n24574 = n24573 ^ n8685 ^ 1'b0 ;
  assign n24575 = n15446 & ~n24574 ;
  assign n24576 = ~n9579 & n14358 ;
  assign n24577 = n5665 | n8663 ;
  assign n24578 = n24577 ^ n18528 ^ 1'b0 ;
  assign n24579 = n23430 ^ n19021 ^ 1'b0 ;
  assign n24580 = n7114 ^ n5328 ^ n2114 ;
  assign n24581 = n24580 ^ n10368 ^ 1'b0 ;
  assign n24582 = n5860 & ~n24581 ;
  assign n24583 = ~n24151 & n24582 ;
  assign n24584 = n24583 ^ n17667 ^ 1'b0 ;
  assign n24585 = ( n20510 & ~n24579 ) | ( n20510 & n24584 ) | ( ~n24579 & n24584 ) ;
  assign n24590 = n15653 & n17722 ;
  assign n24587 = ( x34 & n3225 ) | ( x34 & n4658 ) | ( n3225 & n4658 ) ;
  assign n24588 = ~n23720 & n24587 ;
  assign n24589 = n24588 ^ n6539 ^ 1'b0 ;
  assign n24586 = n7044 ^ n4691 ^ 1'b0 ;
  assign n24591 = n24590 ^ n24589 ^ n24586 ;
  assign n24592 = n19807 ^ n15076 ^ n6954 ;
  assign n24593 = n11914 & n11961 ;
  assign n24594 = n24593 ^ n18422 ^ 1'b0 ;
  assign n24596 = n9253 & ~n12972 ;
  assign n24597 = n4161 & n24596 ;
  assign n24595 = n6130 & ~n24559 ;
  assign n24598 = n24597 ^ n24595 ^ 1'b0 ;
  assign n24599 = n5524 & n17215 ;
  assign n24600 = n5095 & n24599 ;
  assign n24601 = ( n7254 & n16807 ) | ( n7254 & n24600 ) | ( n16807 & n24600 ) ;
  assign n24602 = n20964 ^ n3912 ^ 1'b0 ;
  assign n24603 = n4643 | n24602 ;
  assign n24604 = ( ~n2052 & n3530 ) | ( ~n2052 & n3534 ) | ( n3530 & n3534 ) ;
  assign n24605 = n24604 ^ n23401 ^ n10505 ;
  assign n24606 = n6338 ^ n2751 ^ 1'b0 ;
  assign n24607 = ( n2555 & ~n9349 ) | ( n2555 & n23739 ) | ( ~n9349 & n23739 ) ;
  assign n24608 = n353 & ~n11888 ;
  assign n24609 = n24608 ^ n10092 ^ 1'b0 ;
  assign n24610 = n10122 & n24609 ;
  assign n24611 = n24610 ^ n18365 ^ 1'b0 ;
  assign n24612 = n18538 ^ n12502 ^ 1'b0 ;
  assign n24613 = ~n3411 & n4851 ;
  assign n24614 = n7743 ^ n1208 ^ 1'b0 ;
  assign n24615 = n24613 | n24614 ;
  assign n24616 = n6488 ^ n4304 ^ 1'b0 ;
  assign n24617 = ~n937 & n5896 ;
  assign n24618 = n18039 & n24617 ;
  assign n24619 = n24618 ^ n22281 ^ n8427 ;
  assign n24620 = ( n244 & ~n4491 ) | ( n244 & n17620 ) | ( ~n4491 & n17620 ) ;
  assign n24621 = n5356 & ~n9208 ;
  assign n24622 = ( n142 & n1327 ) | ( n142 & ~n16102 ) | ( n1327 & ~n16102 ) ;
  assign n24623 = n7677 | n7795 ;
  assign n24624 = n24622 & ~n24623 ;
  assign n24627 = ~n2203 & n3830 ;
  assign n24628 = n24627 ^ n3026 ^ 1'b0 ;
  assign n24625 = n18818 ^ n7046 ^ 1'b0 ;
  assign n24626 = ( n1228 & n6369 ) | ( n1228 & n24625 ) | ( n6369 & n24625 ) ;
  assign n24629 = n24628 ^ n24626 ^ n9169 ;
  assign n24630 = n20198 ^ n3487 ^ n3462 ;
  assign n24631 = n19414 & n20852 ;
  assign n24632 = n24631 ^ n17106 ^ 1'b0 ;
  assign n24633 = ~n20532 & n24632 ;
  assign n24634 = n21464 ^ n15150 ^ 1'b0 ;
  assign n24635 = ~n2392 & n21545 ;
  assign n24636 = n24635 ^ n10019 ^ 1'b0 ;
  assign n24637 = ~n1888 & n3035 ;
  assign n24638 = ( n10504 & n17926 ) | ( n10504 & ~n24637 ) | ( n17926 & ~n24637 ) ;
  assign n24639 = ( n18073 & n24636 ) | ( n18073 & ~n24638 ) | ( n24636 & ~n24638 ) ;
  assign n24640 = n24639 ^ n2665 ^ 1'b0 ;
  assign n24641 = ~n8320 & n24640 ;
  assign n24642 = ( n1048 & ~n12129 ) | ( n1048 & n16830 ) | ( ~n12129 & n16830 ) ;
  assign n24643 = ~n1359 & n24642 ;
  assign n24644 = n24643 ^ n22972 ^ 1'b0 ;
  assign n24645 = n7093 ^ n5566 ^ 1'b0 ;
  assign n24646 = n6353 ^ n2674 ^ 1'b0 ;
  assign n24647 = n24645 & ~n24646 ;
  assign n24648 = ( n1200 & n2582 ) | ( n1200 & n4688 ) | ( n2582 & n4688 ) ;
  assign n24649 = n316 | n5253 ;
  assign n24650 = n21332 | n24649 ;
  assign n24651 = n24650 ^ n21671 ^ n708 ;
  assign n24652 = n3124 & ~n24651 ;
  assign n24653 = n24652 ^ n17883 ^ n903 ;
  assign n24654 = n24653 ^ n471 ^ 1'b0 ;
  assign n24655 = n24648 | n24654 ;
  assign n24656 = n17412 & n20849 ;
  assign n24657 = n24656 ^ n260 ^ 1'b0 ;
  assign n24658 = n3936 ^ n332 ^ 1'b0 ;
  assign n24659 = n10150 & n24658 ;
  assign n24660 = ~n2512 & n24659 ;
  assign n24661 = n24660 ^ n11076 ^ 1'b0 ;
  assign n24662 = ( n2620 & ~n9490 ) | ( n2620 & n24661 ) | ( ~n9490 & n24661 ) ;
  assign n24663 = ( n3253 & ~n9901 ) | ( n3253 & n10984 ) | ( ~n9901 & n10984 ) ;
  assign n24665 = ( n621 & n1600 ) | ( n621 & n5106 ) | ( n1600 & n5106 ) ;
  assign n24666 = n7130 & ~n10367 ;
  assign n24667 = n24665 & n24666 ;
  assign n24664 = n24450 ^ n24351 ^ n20909 ;
  assign n24668 = n24667 ^ n24664 ^ n5501 ;
  assign n24669 = ( n1987 & ~n2365 ) | ( n1987 & n2614 ) | ( ~n2365 & n2614 ) ;
  assign n24670 = n5262 & ~n24669 ;
  assign n24671 = n1486 | n8071 ;
  assign n24672 = x98 & n19887 ;
  assign n24673 = ( n4040 & ~n8156 ) | ( n4040 & n24672 ) | ( ~n8156 & n24672 ) ;
  assign n24674 = ( ~n7092 & n7361 ) | ( ~n7092 & n15517 ) | ( n7361 & n15517 ) ;
  assign n24679 = n3874 | n22187 ;
  assign n24680 = n24679 ^ n2187 ^ 1'b0 ;
  assign n24681 = n24680 ^ n20631 ^ n14656 ;
  assign n24675 = n21489 ^ n15108 ^ n6781 ;
  assign n24676 = n3086 & n9486 ;
  assign n24677 = n24676 ^ n19711 ^ 1'b0 ;
  assign n24678 = n24675 & ~n24677 ;
  assign n24682 = n24681 ^ n24678 ^ 1'b0 ;
  assign n24683 = ( ~n5271 & n20881 ) | ( ~n5271 & n24682 ) | ( n20881 & n24682 ) ;
  assign n24685 = n13441 ^ n6783 ^ n951 ;
  assign n24684 = n1893 & n7166 ;
  assign n24686 = n24685 ^ n24684 ^ 1'b0 ;
  assign n24687 = ( x123 & n2628 ) | ( x123 & n18175 ) | ( n2628 & n18175 ) ;
  assign n24692 = n5595 | n10301 ;
  assign n24693 = ~n10219 & n24692 ;
  assign n24691 = n13935 | n19054 ;
  assign n24694 = n24693 ^ n24691 ^ 1'b0 ;
  assign n24688 = n9135 ^ n412 ^ 1'b0 ;
  assign n24689 = n9311 & n24688 ;
  assign n24690 = n24689 ^ n18907 ^ 1'b0 ;
  assign n24695 = n24694 ^ n24690 ^ n12251 ;
  assign n24696 = n8223 ^ n7166 ^ n6623 ;
  assign n24697 = ( n6274 & n11519 ) | ( n6274 & ~n24696 ) | ( n11519 & ~n24696 ) ;
  assign n24698 = n8505 | n18067 ;
  assign n24699 = n4976 | n24698 ;
  assign n24700 = n1216 & ~n5461 ;
  assign n24701 = n24700 ^ n1071 ^ 1'b0 ;
  assign n24702 = n18029 & n24701 ;
  assign n24703 = n22830 | n24702 ;
  assign n24704 = n21489 | n22296 ;
  assign n24705 = n5695 | n24704 ;
  assign n24706 = ( n8199 & ~n9446 ) | ( n8199 & n9892 ) | ( ~n9446 & n9892 ) ;
  assign n24707 = n24706 ^ n20736 ^ n8375 ;
  assign n24708 = n12486 ^ n9076 ^ n6239 ;
  assign n24709 = n20502 ^ n16036 ^ 1'b0 ;
  assign n24710 = n24709 ^ n23724 ^ n2746 ;
  assign n24711 = n20067 ^ n7548 ^ 1'b0 ;
  assign n24712 = n8179 & ~n11253 ;
  assign n24713 = ~n24711 & n24712 ;
  assign n24714 = n941 & n14639 ;
  assign n24715 = ~n3482 & n24714 ;
  assign n24716 = n7507 ^ n5558 ^ n512 ;
  assign n24717 = ( n158 & ~n2446 ) | ( n158 & n8796 ) | ( ~n2446 & n8796 ) ;
  assign n24718 = n24717 ^ n10690 ^ 1'b0 ;
  assign n24719 = n11256 ^ n10484 ^ 1'b0 ;
  assign n24720 = ( n2452 & ~n20510 ) | ( n2452 & n24719 ) | ( ~n20510 & n24719 ) ;
  assign n24721 = ( n4716 & n8251 ) | ( n4716 & n9580 ) | ( n8251 & n9580 ) ;
  assign n24722 = n18092 ^ n10543 ^ 1'b0 ;
  assign n24723 = n22422 ^ n6820 ^ n179 ;
  assign n24724 = n7745 ^ n5809 ^ n3827 ;
  assign n24725 = n10515 & ~n11055 ;
  assign n24726 = n24724 & n24725 ;
  assign n24727 = n5570 & n24726 ;
  assign n24728 = n24727 ^ n5536 ^ 1'b0 ;
  assign n24729 = ~n24723 & n24728 ;
  assign n24730 = n16298 ^ n12966 ^ 1'b0 ;
  assign n24731 = n16009 ^ n7599 ^ n3258 ;
  assign n24732 = n16192 | n24731 ;
  assign n24733 = n4725 | n24732 ;
  assign n24734 = n24733 ^ n1368 ^ 1'b0 ;
  assign n24735 = n4838 & ~n18531 ;
  assign n24736 = n2549 & n9936 ;
  assign n24737 = n24736 ^ x95 ^ 1'b0 ;
  assign n24738 = n19449 ^ n3564 ^ n2786 ;
  assign n24739 = ( ~n15508 & n24737 ) | ( ~n15508 & n24738 ) | ( n24737 & n24738 ) ;
  assign n24740 = n14818 & n17722 ;
  assign n24741 = n6444 & n10386 ;
  assign n24742 = n24741 ^ x68 ^ 1'b0 ;
  assign n24743 = n20717 | n24742 ;
  assign n24744 = ~n3816 & n9903 ;
  assign n24745 = n5846 ^ n356 ^ 1'b0 ;
  assign n24746 = ~n1802 & n24745 ;
  assign n24747 = n7377 & n24746 ;
  assign n24748 = n24744 & n24747 ;
  assign n24749 = n1106 & ~n24748 ;
  assign n24750 = n24749 ^ n3451 ^ 1'b0 ;
  assign n24751 = ( ~n10963 & n13953 ) | ( ~n10963 & n15437 ) | ( n13953 & n15437 ) ;
  assign n24752 = n24751 ^ n11526 ^ 1'b0 ;
  assign n24753 = ~n4283 & n24752 ;
  assign n24754 = ~n18521 & n24753 ;
  assign n24755 = n24754 ^ n8072 ^ 1'b0 ;
  assign n24757 = n3810 | n9448 ;
  assign n24758 = n18432 ^ n7904 ^ 1'b0 ;
  assign n24759 = n24757 & ~n24758 ;
  assign n24760 = n1353 | n24759 ;
  assign n24756 = n11483 & n19822 ;
  assign n24761 = n24760 ^ n24756 ^ 1'b0 ;
  assign n24762 = ~n5970 & n16952 ;
  assign n24763 = n24762 ^ n18593 ^ n3374 ;
  assign n24764 = n24763 ^ n12554 ^ n2184 ;
  assign n24765 = n2361 | n9407 ;
  assign n24766 = n24765 ^ n18689 ^ 1'b0 ;
  assign n24767 = ~n24477 & n24766 ;
  assign n24768 = n304 & n2261 ;
  assign n24769 = n2048 & n11474 ;
  assign n24770 = n24768 & n24769 ;
  assign n24771 = n6278 & ~n24770 ;
  assign n24777 = ( ~n1396 & n2116 ) | ( ~n1396 & n12395 ) | ( n2116 & n12395 ) ;
  assign n24772 = n6532 | n10108 ;
  assign n24773 = n2864 | n24772 ;
  assign n24774 = n2799 & n4962 ;
  assign n24775 = ~n3841 & n24774 ;
  assign n24776 = ( ~n8609 & n24773 ) | ( ~n8609 & n24775 ) | ( n24773 & n24775 ) ;
  assign n24778 = n24777 ^ n24776 ^ n14005 ;
  assign n24779 = ( n167 & ~n8837 ) | ( n167 & n12070 ) | ( ~n8837 & n12070 ) ;
  assign n24780 = ( n9473 & n10401 ) | ( n9473 & n24779 ) | ( n10401 & n24779 ) ;
  assign n24781 = n8200 & ~n23580 ;
  assign n24782 = n12440 ^ n1019 ^ 1'b0 ;
  assign n24783 = ~n24781 & n24782 ;
  assign n24784 = n20575 & ~n23364 ;
  assign n24785 = n15315 ^ n2972 ^ n1772 ;
  assign n24786 = n24785 ^ n5951 ^ n3026 ;
  assign n24787 = ( n6571 & n21376 ) | ( n6571 & n24786 ) | ( n21376 & n24786 ) ;
  assign n24788 = n19191 ^ n15874 ^ 1'b0 ;
  assign n24789 = ~n12396 & n24788 ;
  assign n24790 = n24789 ^ n20044 ^ n9850 ;
  assign n24791 = n22425 ^ n11249 ^ 1'b0 ;
  assign n24792 = ( n8632 & n9145 ) | ( n8632 & n24791 ) | ( n9145 & n24791 ) ;
  assign n24793 = n16857 ^ n12791 ^ n4864 ;
  assign n24796 = n10126 & n16979 ;
  assign n24797 = ~n5529 & n24796 ;
  assign n24795 = n21290 ^ n9682 ^ 1'b0 ;
  assign n24794 = n24164 ^ n12731 ^ n3812 ;
  assign n24798 = n24797 ^ n24795 ^ n24794 ;
  assign n24799 = n15965 ^ n10302 ^ n3646 ;
  assign n24800 = n24799 ^ n6354 ^ n1597 ;
  assign n24801 = n4639 | n24800 ;
  assign n24802 = n992 & ~n24801 ;
  assign n24803 = n8546 & ~n16089 ;
  assign n24804 = n24803 ^ n271 ^ 1'b0 ;
  assign n24805 = ~n19005 & n24804 ;
  assign n24806 = n17441 & n24805 ;
  assign n24807 = n607 & ~n1890 ;
  assign n24808 = n3398 & ~n13867 ;
  assign n24809 = n24808 ^ n10465 ^ 1'b0 ;
  assign n24810 = n24809 ^ n12757 ^ n11600 ;
  assign n24811 = ~n24807 & n24810 ;
  assign n24812 = ~n15126 & n22124 ;
  assign n24813 = ( n19394 & n20044 ) | ( n19394 & ~n24812 ) | ( n20044 & ~n24812 ) ;
  assign n24814 = n9253 ^ n5695 ^ n2624 ;
  assign n24815 = n15574 ^ n6287 ^ 1'b0 ;
  assign n24816 = n18439 & ~n24815 ;
  assign n24817 = ~n24814 & n24816 ;
  assign n24818 = ~n23636 & n24817 ;
  assign n24819 = ( ~n8151 & n24477 ) | ( ~n8151 & n24818 ) | ( n24477 & n24818 ) ;
  assign n24820 = ~n1728 & n19719 ;
  assign n24821 = ~n884 & n3743 ;
  assign n24822 = n24820 & n24821 ;
  assign n24823 = ~n3495 & n5927 ;
  assign n24824 = n24823 ^ n10002 ^ 1'b0 ;
  assign n24825 = n8082 ^ n5843 ^ 1'b0 ;
  assign n24826 = n13581 & n24825 ;
  assign n24827 = n24535 ^ n15801 ^ 1'b0 ;
  assign n24828 = n9679 ^ n2114 ^ 1'b0 ;
  assign n24829 = n2432 & n13842 ;
  assign n24830 = n21378 ^ n7977 ^ 1'b0 ;
  assign n24831 = n3147 & n12148 ;
  assign n24832 = n4588 | n9967 ;
  assign n24833 = n24831 | n24832 ;
  assign n24834 = ( n6303 & n19722 ) | ( n6303 & ~n24833 ) | ( n19722 & ~n24833 ) ;
  assign n24835 = ( n16411 & n24830 ) | ( n16411 & n24834 ) | ( n24830 & n24834 ) ;
  assign n24836 = ( n18012 & n24829 ) | ( n18012 & ~n24835 ) | ( n24829 & ~n24835 ) ;
  assign n24837 = n17431 ^ n5790 ^ 1'b0 ;
  assign n24838 = ( n3269 & n11251 ) | ( n3269 & n19439 ) | ( n11251 & n19439 ) ;
  assign n24844 = n11773 ^ n1124 ^ 1'b0 ;
  assign n24845 = n5898 | n24844 ;
  assign n24839 = n16026 ^ n11718 ^ 1'b0 ;
  assign n24841 = n1900 | n19798 ;
  assign n24840 = x85 & n11349 ;
  assign n24842 = n24841 ^ n24840 ^ 1'b0 ;
  assign n24843 = ( n15082 & ~n24839 ) | ( n15082 & n24842 ) | ( ~n24839 & n24842 ) ;
  assign n24846 = n24845 ^ n24843 ^ n2051 ;
  assign n24847 = ( n871 & ~n8706 ) | ( n871 & n24846 ) | ( ~n8706 & n24846 ) ;
  assign n24848 = ( n9929 & n14674 ) | ( n9929 & n14994 ) | ( n14674 & n14994 ) ;
  assign n24849 = n16295 ^ n15781 ^ 1'b0 ;
  assign n24850 = n24848 & ~n24849 ;
  assign n24851 = ~n13351 & n17328 ;
  assign n24852 = n19046 & n24851 ;
  assign n24853 = n10317 ^ n8760 ^ 1'b0 ;
  assign n24854 = n8898 | n24853 ;
  assign n24855 = n5905 | n13208 ;
  assign n24856 = ~n16128 & n16499 ;
  assign n24857 = ~n4002 & n6275 ;
  assign n24858 = n5167 & n24857 ;
  assign n24859 = n24858 ^ n4497 ^ n2438 ;
  assign n24860 = ( n2016 & n20472 ) | ( n2016 & n24859 ) | ( n20472 & n24859 ) ;
  assign n24861 = n18888 ^ n11530 ^ n4372 ;
  assign n24862 = n1243 & ~n6578 ;
  assign n24863 = n24862 ^ n12962 ^ n488 ;
  assign n24864 = ( n8176 & n15644 ) | ( n8176 & ~n24863 ) | ( n15644 & ~n24863 ) ;
  assign n24865 = n8023 | n15734 ;
  assign n24866 = ~n7022 & n24865 ;
  assign n24867 = n24866 ^ n3406 ^ 1'b0 ;
  assign n24868 = ~n834 & n14043 ;
  assign n24869 = n24868 ^ n18147 ^ 1'b0 ;
  assign n24870 = n8303 ^ n2870 ^ 1'b0 ;
  assign n24871 = n20477 & ~n24870 ;
  assign n24872 = ( n13069 & n19950 ) | ( n13069 & n20592 ) | ( n19950 & n20592 ) ;
  assign n24873 = n10597 | n23442 ;
  assign n24874 = ( n14824 & n24872 ) | ( n14824 & ~n24873 ) | ( n24872 & ~n24873 ) ;
  assign n24875 = n19893 ^ n8348 ^ 1'b0 ;
  assign n24876 = n3379 | n24875 ;
  assign n24877 = n20331 & n24876 ;
  assign n24878 = n2777 ^ n2010 ^ 1'b0 ;
  assign n24879 = ~n5911 & n24878 ;
  assign n24880 = n24879 ^ n19726 ^ n15711 ;
  assign n24881 = ( n743 & ~n3774 ) | ( n743 & n13265 ) | ( ~n3774 & n13265 ) ;
  assign n24882 = n24881 ^ n11128 ^ 1'b0 ;
  assign n24891 = n12083 ^ n10716 ^ n3561 ;
  assign n24883 = n5473 | n16006 ;
  assign n24884 = n1691 & ~n24883 ;
  assign n24885 = ( ~n1356 & n4147 ) | ( ~n1356 & n13839 ) | ( n4147 & n13839 ) ;
  assign n24886 = ( ~n1543 & n14205 ) | ( ~n1543 & n24885 ) | ( n14205 & n24885 ) ;
  assign n24887 = n2364 | n3650 ;
  assign n24888 = n24886 & ~n24887 ;
  assign n24889 = ( ~n5879 & n23880 ) | ( ~n5879 & n24471 ) | ( n23880 & n24471 ) ;
  assign n24890 = ( ~n24884 & n24888 ) | ( ~n24884 & n24889 ) | ( n24888 & n24889 ) ;
  assign n24892 = n24891 ^ n24890 ^ 1'b0 ;
  assign n24893 = n14901 ^ n5457 ^ n5252 ;
  assign n24894 = n24893 ^ n17414 ^ 1'b0 ;
  assign n24895 = n12633 | n24894 ;
  assign n24896 = n20792 & ~n24895 ;
  assign n24897 = n4352 ^ n1671 ^ 1'b0 ;
  assign n24898 = ( n16708 & n22707 ) | ( n16708 & ~n24897 ) | ( n22707 & ~n24897 ) ;
  assign n24899 = n24898 ^ n10220 ^ 1'b0 ;
  assign n24900 = ( n2864 & n4737 ) | ( n2864 & n17831 ) | ( n4737 & n17831 ) ;
  assign n24901 = n10221 ^ n1206 ^ 1'b0 ;
  assign n24902 = ( n10609 & n11460 ) | ( n10609 & n24901 ) | ( n11460 & n24901 ) ;
  assign n24903 = n22110 ^ n4267 ^ 1'b0 ;
  assign n24904 = n6706 & n11286 ;
  assign n24905 = n24904 ^ n12279 ^ n1169 ;
  assign n24906 = n12526 ^ n1887 ^ 1'b0 ;
  assign n24907 = ~n8101 & n24906 ;
  assign n24908 = n17291 ^ n4302 ^ n2524 ;
  assign n24909 = n3941 ^ n3281 ^ 1'b0 ;
  assign n24910 = n5033 | n24909 ;
  assign n24911 = n3418 | n24910 ;
  assign n24912 = n3921 & ~n24911 ;
  assign n24913 = ~n24908 & n24912 ;
  assign n24914 = n12155 ^ n3895 ^ 1'b0 ;
  assign n24915 = n8845 & ~n24914 ;
  assign n24916 = n700 & ~n18656 ;
  assign n24917 = n22861 & n24916 ;
  assign n24918 = n24917 ^ n10594 ^ 1'b0 ;
  assign n24919 = n24918 ^ n6397 ^ 1'b0 ;
  assign n24920 = n24915 & n24919 ;
  assign n24921 = n18887 ^ n18680 ^ n4181 ;
  assign n24922 = n21814 ^ n19578 ^ n16660 ;
  assign n24923 = n9452 & ~n24922 ;
  assign n24924 = ~n24244 & n24923 ;
  assign n24925 = n3565 | n24924 ;
  assign n24926 = n24925 ^ n1232 ^ 1'b0 ;
  assign n24927 = n24926 ^ n23081 ^ n4594 ;
  assign n24928 = ( n6934 & n11840 ) | ( n6934 & ~n15663 ) | ( n11840 & ~n15663 ) ;
  assign n24929 = n15233 ^ n988 ^ 1'b0 ;
  assign n24930 = n3314 & n24929 ;
  assign n24931 = n24930 ^ n3982 ^ n1275 ;
  assign n24932 = n24931 ^ n2471 ^ 1'b0 ;
  assign n24933 = n12885 ^ n9881 ^ 1'b0 ;
  assign n24934 = n12998 | n24933 ;
  assign n24935 = ~n660 & n15018 ;
  assign n24936 = ~n24934 & n24935 ;
  assign n24937 = ( n7107 & n9485 ) | ( n7107 & ~n11732 ) | ( n9485 & ~n11732 ) ;
  assign n24938 = n24863 & ~n24937 ;
  assign n24948 = n11703 ^ n4821 ^ 1'b0 ;
  assign n24949 = ( n699 & n16547 ) | ( n699 & ~n24948 ) | ( n16547 & ~n24948 ) ;
  assign n24942 = n1802 | n2417 ;
  assign n24939 = n15860 ^ n3286 ^ 1'b0 ;
  assign n24940 = n24939 ^ n6802 ^ n4512 ;
  assign n24941 = n7782 & n24940 ;
  assign n24943 = n24942 ^ n24941 ^ 1'b0 ;
  assign n24944 = n18069 ^ n8259 ^ 1'b0 ;
  assign n24945 = n16195 & ~n24944 ;
  assign n24946 = ( n1986 & n8895 ) | ( n1986 & ~n24945 ) | ( n8895 & ~n24945 ) ;
  assign n24947 = ( n1139 & n24943 ) | ( n1139 & ~n24946 ) | ( n24943 & ~n24946 ) ;
  assign n24950 = n24949 ^ n24947 ^ n9875 ;
  assign n24953 = n24394 ^ n2194 ^ 1'b0 ;
  assign n24954 = n17615 | n24953 ;
  assign n24951 = n4229 | n17383 ;
  assign n24952 = n24951 ^ n16197 ^ 1'b0 ;
  assign n24955 = n24954 ^ n24952 ^ n3604 ;
  assign n24958 = ( n3022 & ~n8648 ) | ( n3022 & n9782 ) | ( ~n8648 & n9782 ) ;
  assign n24957 = n4585 ^ n4317 ^ 1'b0 ;
  assign n24959 = n24958 ^ n24957 ^ n10756 ;
  assign n24956 = n4455 & ~n22761 ;
  assign n24960 = n24959 ^ n24956 ^ n10141 ;
  assign n24961 = n13009 ^ n12223 ^ 1'b0 ;
  assign n24962 = n24960 & ~n24961 ;
  assign n24963 = ~n7744 & n12789 ;
  assign n24964 = n5946 ^ n4593 ^ 1'b0 ;
  assign n24965 = n5917 & n17957 ;
  assign n24966 = n24964 & n24965 ;
  assign n24967 = n6541 & ~n6985 ;
  assign n24968 = ~n1974 & n24967 ;
  assign n24969 = ( n2545 & n5594 ) | ( n2545 & ~n6897 ) | ( n5594 & ~n6897 ) ;
  assign n24970 = ( n5875 & n9272 ) | ( n5875 & ~n24969 ) | ( n9272 & ~n24969 ) ;
  assign n24971 = n11838 ^ n9446 ^ n1620 ;
  assign n24972 = n579 | n21468 ;
  assign n24973 = n24972 ^ n9345 ^ 1'b0 ;
  assign n24974 = n21039 & ~n24973 ;
  assign n24975 = ~n4522 & n14861 ;
  assign n24976 = n12578 & ~n17071 ;
  assign n24977 = n24976 ^ n20825 ^ 1'b0 ;
  assign n24978 = n7111 | n17875 ;
  assign n24979 = n24978 ^ n4177 ^ 1'b0 ;
  assign n24980 = n3697 ^ n2033 ^ n519 ;
  assign n24981 = ( n11597 & n11792 ) | ( n11597 & n16217 ) | ( n11792 & n16217 ) ;
  assign n24982 = n24981 ^ n6482 ^ n3483 ;
  assign n24983 = ( ~n329 & n10232 ) | ( ~n329 & n24982 ) | ( n10232 & n24982 ) ;
  assign n24984 = ( n11776 & n24980 ) | ( n11776 & n24983 ) | ( n24980 & n24983 ) ;
  assign n24985 = n5568 & ~n10088 ;
  assign n24986 = n24985 ^ n22025 ^ 1'b0 ;
  assign n24987 = n8481 ^ n997 ^ 1'b0 ;
  assign n24988 = n14411 | n24987 ;
  assign n24989 = ( n14808 & ~n24986 ) | ( n14808 & n24988 ) | ( ~n24986 & n24988 ) ;
  assign n24999 = ( n469 & n3006 ) | ( n469 & n13058 ) | ( n3006 & n13058 ) ;
  assign n24996 = ~n3860 & n4335 ;
  assign n24997 = n7038 & n24996 ;
  assign n24993 = n4022 & ~n23328 ;
  assign n24994 = ~n18069 & n24993 ;
  assign n24990 = ( n1898 & n1900 ) | ( n1898 & ~n2606 ) | ( n1900 & ~n2606 ) ;
  assign n24991 = n24990 ^ n18006 ^ n5371 ;
  assign n24992 = n2423 & ~n24991 ;
  assign n24995 = n24994 ^ n24992 ^ 1'b0 ;
  assign n24998 = n24997 ^ n24995 ^ n3845 ;
  assign n25000 = n24999 ^ n24998 ^ n18197 ;
  assign n25001 = n21060 ^ n10041 ^ 1'b0 ;
  assign n25002 = n24791 | n25001 ;
  assign n25003 = ( n15694 & ~n22015 ) | ( n15694 & n25002 ) | ( ~n22015 & n25002 ) ;
  assign n25004 = n24458 ^ n18674 ^ n6462 ;
  assign n25005 = n7627 ^ n1052 ^ n856 ;
  assign n25006 = ( n3013 & ~n7882 ) | ( n3013 & n25005 ) | ( ~n7882 & n25005 ) ;
  assign n25007 = n16066 | n25006 ;
  assign n25008 = ~n1163 & n3722 ;
  assign n25009 = n25008 ^ n9448 ^ 1'b0 ;
  assign n25010 = ( n758 & n8479 ) | ( n758 & n17741 ) | ( n8479 & n17741 ) ;
  assign n25011 = n25010 ^ n5576 ^ 1'b0 ;
  assign n25013 = ( n6424 & ~n6712 ) | ( n6424 & n11246 ) | ( ~n6712 & n11246 ) ;
  assign n25012 = n3841 & ~n6169 ;
  assign n25014 = n25013 ^ n25012 ^ 1'b0 ;
  assign n25018 = n11315 ^ n4819 ^ n3077 ;
  assign n25016 = ( ~n244 & n2146 ) | ( ~n244 & n4550 ) | ( n2146 & n4550 ) ;
  assign n25015 = ( n4428 & n13197 ) | ( n4428 & n15292 ) | ( n13197 & n15292 ) ;
  assign n25017 = n25016 ^ n25015 ^ n24886 ;
  assign n25019 = n25018 ^ n25017 ^ n14685 ;
  assign n25020 = ( n13981 & ~n21327 ) | ( n13981 & n25019 ) | ( ~n21327 & n25019 ) ;
  assign n25021 = n12763 ^ n7399 ^ n6810 ;
  assign n25024 = n6537 & ~n12245 ;
  assign n25025 = n10088 & n25024 ;
  assign n25022 = ( n7473 & n10041 ) | ( n7473 & n13147 ) | ( n10041 & n13147 ) ;
  assign n25023 = ( ~n8606 & n18813 ) | ( ~n8606 & n25022 ) | ( n18813 & n25022 ) ;
  assign n25026 = n25025 ^ n25023 ^ n20138 ;
  assign n25027 = ~n4173 & n8461 ;
  assign n25028 = n1585 & n9206 ;
  assign n25029 = n3816 ^ x25 ^ 1'b0 ;
  assign n25030 = n25028 & n25029 ;
  assign n25031 = n10150 ^ n6762 ^ 1'b0 ;
  assign n25032 = n4240 & ~n25031 ;
  assign n25033 = n2881 | n25032 ;
  assign n25037 = n12434 ^ n11483 ^ 1'b0 ;
  assign n25034 = n22210 ^ n15900 ^ n7230 ;
  assign n25035 = ( ~n673 & n11560 ) | ( ~n673 & n25034 ) | ( n11560 & n25034 ) ;
  assign n25036 = n25035 ^ n7482 ^ 1'b0 ;
  assign n25038 = n25037 ^ n25036 ^ n20686 ;
  assign n25042 = ( n11281 & ~n11952 ) | ( n11281 & n16696 ) | ( ~n11952 & n16696 ) ;
  assign n25043 = n13713 ^ n2242 ^ 1'b0 ;
  assign n25044 = n25042 & ~n25043 ;
  assign n25039 = n3267 & ~n19700 ;
  assign n25040 = n25039 ^ n6448 ^ 1'b0 ;
  assign n25041 = n25040 ^ n24731 ^ n6487 ;
  assign n25045 = n25044 ^ n25041 ^ n3225 ;
  assign n25046 = n2081 & n7731 ;
  assign n25047 = n25046 ^ n12671 ^ 1'b0 ;
  assign n25048 = n5230 & n7030 ;
  assign n25049 = n25048 ^ n6501 ^ 1'b0 ;
  assign n25050 = ~n24750 & n25049 ;
  assign n25051 = n19010 ^ n7548 ^ 1'b0 ;
  assign n25057 = ~n7199 & n8154 ;
  assign n25055 = ( ~n3827 & n8395 ) | ( ~n3827 & n15170 ) | ( n8395 & n15170 ) ;
  assign n25052 = ( n1002 & n4645 ) | ( n1002 & ~n10223 ) | ( n4645 & ~n10223 ) ;
  assign n25053 = n11690 | n25052 ;
  assign n25054 = n25053 ^ n4003 ^ 1'b0 ;
  assign n25056 = n25055 ^ n25054 ^ n2383 ;
  assign n25058 = n25057 ^ n25056 ^ n17632 ;
  assign n25059 = n20367 ^ n13314 ^ 1'b0 ;
  assign n25060 = n8686 & ~n25059 ;
  assign n25061 = ( ~n4917 & n5695 ) | ( ~n4917 & n25060 ) | ( n5695 & n25060 ) ;
  assign n25062 = n12855 ^ n7828 ^ 1'b0 ;
  assign n25063 = n2493 & n25062 ;
  assign n25064 = ~n10394 & n13112 ;
  assign n25065 = ~n21921 & n25064 ;
  assign n25066 = n6337 ^ n4482 ^ n2488 ;
  assign n25067 = n8175 & n10678 ;
  assign n25068 = ( n13087 & n18040 ) | ( n13087 & n25067 ) | ( n18040 & n25067 ) ;
  assign n25069 = n13601 & n14073 ;
  assign n25070 = n4821 ^ n3377 ^ 1'b0 ;
  assign n25071 = n25070 ^ n20188 ^ n9905 ;
  assign n25072 = n1180 ^ n698 ^ 1'b0 ;
  assign n25073 = ~n14058 & n25072 ;
  assign n25074 = n25071 & n25073 ;
  assign n25075 = n9286 ^ n8730 ^ n3875 ;
  assign n25076 = n22542 | n25075 ;
  assign n25077 = n3096 | n25076 ;
  assign n25078 = n25077 ^ n15608 ^ 1'b0 ;
  assign n25079 = n18554 ^ n16561 ^ 1'b0 ;
  assign n25080 = n3149 & n18618 ;
  assign n25081 = n6341 & n25080 ;
  assign n25082 = ( n1817 & ~n12480 ) | ( n1817 & n25081 ) | ( ~n12480 & n25081 ) ;
  assign n25083 = n25082 ^ n8604 ^ 1'b0 ;
  assign n25084 = ( n6858 & n9753 ) | ( n6858 & n9860 ) | ( n9753 & n9860 ) ;
  assign n25085 = n25084 ^ n21364 ^ n19420 ;
  assign n25086 = ( n6809 & ~n7409 ) | ( n6809 & n12789 ) | ( ~n7409 & n12789 ) ;
  assign n25087 = n20327 ^ n8800 ^ 1'b0 ;
  assign n25088 = n17774 & ~n25087 ;
  assign n25089 = n11107 ^ n953 ^ 1'b0 ;
  assign n25090 = n4020 | n25089 ;
  assign n25091 = n1684 & n6744 ;
  assign n25092 = ~n2423 & n25091 ;
  assign n25093 = n25092 ^ n4351 ^ 1'b0 ;
  assign n25094 = n25093 ^ n15827 ^ n13210 ;
  assign n25095 = n6991 ^ n5920 ^ n3273 ;
  assign n25099 = ( ~n1090 & n4239 ) | ( ~n1090 & n8850 ) | ( n4239 & n8850 ) ;
  assign n25096 = ( n11859 & ~n15613 ) | ( n11859 & n16518 ) | ( ~n15613 & n16518 ) ;
  assign n25097 = ~n2849 & n13402 ;
  assign n25098 = ~n25096 & n25097 ;
  assign n25100 = n25099 ^ n25098 ^ 1'b0 ;
  assign n25101 = ( x114 & ~n9542 ) | ( x114 & n25100 ) | ( ~n9542 & n25100 ) ;
  assign n25102 = ( n4195 & n10983 ) | ( n4195 & n18045 ) | ( n10983 & n18045 ) ;
  assign n25103 = ( ~n13782 & n25101 ) | ( ~n13782 & n25102 ) | ( n25101 & n25102 ) ;
  assign n25104 = n17587 ^ n13688 ^ 1'b0 ;
  assign n25105 = ( n1716 & n14173 ) | ( n1716 & ~n25104 ) | ( n14173 & ~n25104 ) ;
  assign n25106 = ( n16072 & ~n17296 ) | ( n16072 & n18006 ) | ( ~n17296 & n18006 ) ;
  assign n25107 = n25106 ^ n12099 ^ n7415 ;
  assign n25108 = n25107 ^ n15285 ^ n14153 ;
  assign n25109 = ~n4374 & n11806 ;
  assign n25110 = n25109 ^ n23645 ^ 1'b0 ;
  assign n25111 = n20686 ^ n7388 ^ 1'b0 ;
  assign n25112 = n3996 & n25111 ;
  assign n25113 = n15695 ^ n15246 ^ 1'b0 ;
  assign n25114 = ( n7757 & n9363 ) | ( n7757 & n15100 ) | ( n9363 & n15100 ) ;
  assign n25118 = n19580 ^ n4157 ^ n743 ;
  assign n25115 = ~n3053 & n23654 ;
  assign n25116 = n25115 ^ n904 ^ 1'b0 ;
  assign n25117 = n25116 ^ n17791 ^ n5590 ;
  assign n25119 = n25118 ^ n25117 ^ n14867 ;
  assign n25121 = n5079 | n7329 ;
  assign n25122 = n25121 ^ n2619 ^ 1'b0 ;
  assign n25120 = ( n2514 & ~n2967 ) | ( n2514 & n10770 ) | ( ~n2967 & n10770 ) ;
  assign n25123 = n25122 ^ n25120 ^ n5238 ;
  assign n25124 = n3934 | n25123 ;
  assign n25125 = ( n6958 & n16217 ) | ( n6958 & ~n18888 ) | ( n16217 & ~n18888 ) ;
  assign n25126 = ~n19185 & n25125 ;
  assign n25127 = n20743 ^ n9298 ^ 1'b0 ;
  assign n25128 = n25126 | n25127 ;
  assign n25129 = n17488 ^ n10028 ^ n9360 ;
  assign n25130 = n23567 | n25129 ;
  assign n25133 = n5814 & n8946 ;
  assign n25132 = ( n220 & n7215 ) | ( n220 & ~n13384 ) | ( n7215 & ~n13384 ) ;
  assign n25131 = n8723 ^ x56 ^ 1'b0 ;
  assign n25134 = n25133 ^ n25132 ^ n25131 ;
  assign n25135 = n19595 ^ n12296 ^ n10115 ;
  assign n25136 = n5308 | n15835 ;
  assign n25137 = ( n575 & n2781 ) | ( n575 & n25136 ) | ( n2781 & n25136 ) ;
  assign n25138 = n20994 & n21891 ;
  assign n25139 = n4076 & n6976 ;
  assign n25140 = n19273 ^ n9327 ^ 1'b0 ;
  assign n25141 = n3807 | n25140 ;
  assign n25142 = n25141 ^ n10578 ^ 1'b0 ;
  assign n25143 = n8667 ^ n2761 ^ 1'b0 ;
  assign n25144 = n4503 & n25143 ;
  assign n25145 = n5751 & n25144 ;
  assign n25146 = ( n732 & n3528 ) | ( n732 & n5748 ) | ( n3528 & n5748 ) ;
  assign n25147 = ( n2009 & n4268 ) | ( n2009 & n5150 ) | ( n4268 & n5150 ) ;
  assign n25148 = n16193 & ~n17560 ;
  assign n25149 = ~n24415 & n25148 ;
  assign n25150 = ( n12354 & n25147 ) | ( n12354 & n25149 ) | ( n25147 & n25149 ) ;
  assign n25151 = ( ~x18 & n6382 ) | ( ~x18 & n25016 ) | ( n6382 & n25016 ) ;
  assign n25152 = n25151 ^ n15722 ^ 1'b0 ;
  assign n25153 = n23521 ^ n7942 ^ 1'b0 ;
  assign n25154 = n7477 ^ n313 ^ 1'b0 ;
  assign n25155 = n1940 & n25154 ;
  assign n25156 = n25155 ^ n9758 ^ n8398 ;
  assign n25157 = n2079 & ~n6555 ;
  assign n25158 = ~n3213 & n25157 ;
  assign n25159 = n25156 | n25158 ;
  assign n25160 = n6482 ^ n6152 ^ n3634 ;
  assign n25161 = n367 | n4705 ;
  assign n25162 = n25161 ^ n4621 ^ 1'b0 ;
  assign n25163 = n25160 & ~n25162 ;
  assign n25164 = n16317 ^ n2355 ^ 1'b0 ;
  assign n25165 = n2406 & n25164 ;
  assign n25166 = n25165 ^ n19268 ^ n5399 ;
  assign n25167 = n1125 | n5377 ;
  assign n25168 = n16465 | n25167 ;
  assign n25169 = n25168 ^ n18107 ^ n11428 ;
  assign n25170 = n12891 ^ n11074 ^ n6454 ;
  assign n25171 = ( n4547 & n17662 ) | ( n4547 & n25170 ) | ( n17662 & n25170 ) ;
  assign n25172 = n25171 ^ n5598 ^ n4863 ;
  assign n25173 = n9694 ^ n2567 ^ 1'b0 ;
  assign n25174 = ~n22515 & n25173 ;
  assign n25175 = n20900 ^ n9977 ^ n2537 ;
  assign n25176 = ( n10009 & ~n12571 ) | ( n10009 & n25175 ) | ( ~n12571 & n25175 ) ;
  assign n25177 = n25176 ^ n20324 ^ n19593 ;
  assign n25178 = n15049 ^ n10827 ^ n4403 ;
  assign n25179 = n25178 ^ n1657 ^ 1'b0 ;
  assign n25180 = ( n10662 & n24207 ) | ( n10662 & ~n25179 ) | ( n24207 & ~n25179 ) ;
  assign n25181 = n21752 ^ n4055 ^ n636 ;
  assign n25182 = n25181 ^ n23513 ^ 1'b0 ;
  assign n25183 = n13074 | n15990 ;
  assign n25184 = n7736 & ~n25183 ;
  assign n25185 = n25184 ^ n1848 ^ 1'b0 ;
  assign n25186 = n4337 ^ n1250 ^ 1'b0 ;
  assign n25187 = ( ~n6282 & n11275 ) | ( ~n6282 & n12358 ) | ( n11275 & n12358 ) ;
  assign n25188 = ~n7280 & n25187 ;
  assign n25189 = ~n2394 & n25188 ;
  assign n25190 = n16366 ^ n5887 ^ n3075 ;
  assign n25191 = n20785 ^ n13938 ^ 1'b0 ;
  assign n25194 = n6691 & n21696 ;
  assign n25192 = n8913 | n15752 ;
  assign n25193 = n4461 | n25192 ;
  assign n25195 = n25194 ^ n25193 ^ n4183 ;
  assign n25196 = n25195 ^ n8292 ^ n180 ;
  assign n25198 = n5731 & n10301 ;
  assign n25197 = n2615 & n21007 ;
  assign n25199 = n25198 ^ n25197 ^ 1'b0 ;
  assign n25200 = n13164 ^ n12115 ^ 1'b0 ;
  assign n25201 = ~n17227 & n25200 ;
  assign n25202 = ~n11563 & n25201 ;
  assign n25203 = n25202 ^ n8925 ^ n4425 ;
  assign n25204 = n25203 ^ n10141 ^ 1'b0 ;
  assign n25205 = n25199 & n25204 ;
  assign n25206 = n4920 & ~n5086 ;
  assign n25207 = n14586 & n25206 ;
  assign n25208 = ( ~n2851 & n6987 ) | ( ~n2851 & n25207 ) | ( n6987 & n25207 ) ;
  assign n25209 = n8886 ^ n6198 ^ n6070 ;
  assign n25210 = ~n5376 & n25209 ;
  assign n25211 = ~n24652 & n25210 ;
  assign n25212 = n14265 ^ n7774 ^ 1'b0 ;
  assign n25213 = ~n1649 & n9462 ;
  assign n25214 = n25213 ^ n21002 ^ 1'b0 ;
  assign n25215 = n12573 ^ n2839 ^ 1'b0 ;
  assign n25216 = ~n1553 & n25215 ;
  assign n25217 = n10625 ^ n7942 ^ n7331 ;
  assign n25218 = ( n2488 & ~n8470 ) | ( n2488 & n25217 ) | ( ~n8470 & n25217 ) ;
  assign n25219 = n24248 & ~n25218 ;
  assign n25220 = n11386 ^ n10998 ^ n9022 ;
  assign n25221 = ~n17188 & n22871 ;
  assign n25222 = ( n3050 & n25220 ) | ( n3050 & ~n25221 ) | ( n25220 & ~n25221 ) ;
  assign n25223 = ( n5979 & n7065 ) | ( n5979 & n11130 ) | ( n7065 & n11130 ) ;
  assign n25224 = n14793 ^ n14520 ^ n10145 ;
  assign n25225 = ( n3269 & ~n8663 ) | ( n3269 & n20671 ) | ( ~n8663 & n20671 ) ;
  assign n25226 = ( ~n3035 & n4624 ) | ( ~n3035 & n6783 ) | ( n4624 & n6783 ) ;
  assign n25227 = n25226 ^ n7627 ^ 1'b0 ;
  assign n25228 = n23988 ^ n288 ^ 1'b0 ;
  assign n25229 = n1955 | n4540 ;
  assign n25230 = n25229 ^ n10823 ^ 1'b0 ;
  assign n25231 = n25230 ^ n23900 ^ n11976 ;
  assign n25232 = ( n3944 & n21676 ) | ( n3944 & n25231 ) | ( n21676 & n25231 ) ;
  assign n25233 = n3325 & ~n10627 ;
  assign n25234 = n25233 ^ n20348 ^ 1'b0 ;
  assign n25235 = ( n14485 & n15304 ) | ( n14485 & ~n25234 ) | ( n15304 & ~n25234 ) ;
  assign n25236 = n22459 ^ n19110 ^ 1'b0 ;
  assign n25237 = ( n1023 & n6429 ) | ( n1023 & n22764 ) | ( n6429 & n22764 ) ;
  assign n25238 = n8470 & ~n23847 ;
  assign n25239 = ~n21176 & n25238 ;
  assign n25240 = n25239 ^ n3220 ^ n2507 ;
  assign n25241 = n8094 ^ n4736 ^ n544 ;
  assign n25242 = n25241 ^ n1405 ^ 1'b0 ;
  assign n25243 = ~n13919 & n25242 ;
  assign n25244 = n17520 ^ n6288 ^ 1'b0 ;
  assign n25245 = ~n11289 & n25244 ;
  assign n25246 = ( ~n3749 & n8097 ) | ( ~n3749 & n11449 ) | ( n8097 & n11449 ) ;
  assign n25247 = n22799 ^ n6275 ^ n5920 ;
  assign n25248 = n4805 ^ n2894 ^ 1'b0 ;
  assign n25249 = ~n1451 & n25248 ;
  assign n25250 = ( n4896 & n15063 ) | ( n4896 & ~n18902 ) | ( n15063 & ~n18902 ) ;
  assign n25251 = n25250 ^ n19824 ^ 1'b0 ;
  assign n25252 = ( ~n23800 & n25249 ) | ( ~n23800 & n25251 ) | ( n25249 & n25251 ) ;
  assign n25253 = ( n3728 & n7497 ) | ( n3728 & ~n22081 ) | ( n7497 & ~n22081 ) ;
  assign n25254 = n20151 ^ n3212 ^ n2252 ;
  assign n25255 = n2301 & ~n4734 ;
  assign n25256 = n4273 & n12093 ;
  assign n25257 = n18247 & n25256 ;
  assign n25258 = n25257 ^ n12798 ^ 1'b0 ;
  assign n25259 = n15571 | n16410 ;
  assign n25260 = n25259 ^ n9982 ^ 1'b0 ;
  assign n25261 = n20090 ^ n1832 ^ 1'b0 ;
  assign n25262 = n5142 & n25261 ;
  assign n25263 = ~n17687 & n25262 ;
  assign n25264 = n25263 ^ n13891 ^ 1'b0 ;
  assign n25265 = n5085 & ~n7473 ;
  assign n25266 = n25265 ^ n7362 ^ 1'b0 ;
  assign n25267 = ( n8770 & n24127 ) | ( n8770 & ~n25266 ) | ( n24127 & ~n25266 ) ;
  assign n25268 = n7780 | n10318 ;
  assign n25269 = n25268 ^ n14559 ^ 1'b0 ;
  assign n25270 = n22883 | n25269 ;
  assign n25271 = ~n2695 & n10089 ;
  assign n25272 = ( n11000 & ~n15760 ) | ( n11000 & n25271 ) | ( ~n15760 & n25271 ) ;
  assign n25273 = ( n18375 & ~n24374 ) | ( n18375 & n25272 ) | ( ~n24374 & n25272 ) ;
  assign n25274 = ~n900 & n15911 ;
  assign n25275 = ( ~n1315 & n2638 ) | ( ~n1315 & n10230 ) | ( n2638 & n10230 ) ;
  assign n25276 = n25275 ^ n5222 ^ 1'b0 ;
  assign n25277 = n9920 & n25276 ;
  assign n25278 = n4286 & ~n10355 ;
  assign n25279 = ~n7102 & n10020 ;
  assign n25280 = n11536 & n25279 ;
  assign n25281 = ( n6582 & n7031 ) | ( n6582 & n7197 ) | ( n7031 & n7197 ) ;
  assign n25282 = n13141 & ~n25281 ;
  assign n25283 = n5106 & n12003 ;
  assign n25287 = n15510 ^ n4229 ^ 1'b0 ;
  assign n25284 = n8646 ^ n4858 ^ 1'b0 ;
  assign n25285 = n9756 & ~n25284 ;
  assign n25286 = n21632 & n25285 ;
  assign n25288 = n25287 ^ n25286 ^ 1'b0 ;
  assign n25289 = ( n12247 & n25283 ) | ( n12247 & n25288 ) | ( n25283 & n25288 ) ;
  assign n25290 = n24298 ^ n16779 ^ n8146 ;
  assign n25291 = n6471 & ~n25081 ;
  assign n25292 = ~n3943 & n25291 ;
  assign n25293 = ~n3646 & n25292 ;
  assign n25294 = n25042 ^ n1927 ^ 1'b0 ;
  assign n25295 = n25294 ^ n9240 ^ 1'b0 ;
  assign n25296 = n22898 ^ n10488 ^ n569 ;
  assign n25297 = n25296 ^ n6069 ^ n3906 ;
  assign n25298 = n25297 ^ n2389 ^ n665 ;
  assign n25299 = n11418 ^ n6353 ^ 1'b0 ;
  assign n25300 = n11807 ^ n5256 ^ 1'b0 ;
  assign n25301 = n25299 | n25300 ;
  assign n25302 = n12830 ^ n11417 ^ n3148 ;
  assign n25303 = n6621 ^ n716 ^ 1'b0 ;
  assign n25304 = n25302 | n25303 ;
  assign n25305 = n19290 ^ n15822 ^ 1'b0 ;
  assign n25306 = n4918 | n11597 ;
  assign n25307 = n25306 ^ n17494 ^ 1'b0 ;
  assign n25311 = ~n4899 & n12875 ;
  assign n25312 = n25311 ^ n8275 ^ 1'b0 ;
  assign n25308 = n2809 ^ n2733 ^ 1'b0 ;
  assign n25309 = n207 & n25308 ;
  assign n25310 = ~n20324 & n25309 ;
  assign n25313 = n25312 ^ n25310 ^ n22727 ;
  assign n25314 = n16193 ^ n12339 ^ n11435 ;
  assign n25315 = n18134 | n24384 ;
  assign n25316 = ( n10898 & n25314 ) | ( n10898 & ~n25315 ) | ( n25314 & ~n25315 ) ;
  assign n25317 = n24757 ^ n18264 ^ 1'b0 ;
  assign n25318 = n2466 ^ n892 ^ 1'b0 ;
  assign n25319 = n7256 ^ n409 ^ 1'b0 ;
  assign n25320 = ( n11956 & ~n14963 ) | ( n11956 & n25319 ) | ( ~n14963 & n25319 ) ;
  assign n25321 = ( n2656 & ~n5545 ) | ( n2656 & n10368 ) | ( ~n5545 & n10368 ) ;
  assign n25322 = ~n8473 & n25321 ;
  assign n25323 = ( n11263 & n23590 ) | ( n11263 & ~n25322 ) | ( n23590 & ~n25322 ) ;
  assign n25324 = n969 & ~n5153 ;
  assign n25325 = ( n8062 & n11651 ) | ( n8062 & ~n25324 ) | ( n11651 & ~n25324 ) ;
  assign n25326 = n6454 ^ n575 ^ 1'b0 ;
  assign n25327 = ( n10814 & ~n23847 ) | ( n10814 & n25326 ) | ( ~n23847 & n25326 ) ;
  assign n25328 = n25327 ^ n5696 ^ n171 ;
  assign n25329 = ( n24810 & n25325 ) | ( n24810 & n25328 ) | ( n25325 & n25328 ) ;
  assign n25331 = n7544 & ~n7577 ;
  assign n25330 = n2884 & ~n14414 ;
  assign n25332 = n25331 ^ n25330 ^ 1'b0 ;
  assign n25333 = n691 | n25332 ;
  assign n25334 = n24524 ^ n3012 ^ 1'b0 ;
  assign n25335 = n20270 ^ n7386 ^ 1'b0 ;
  assign n25336 = n10748 | n25335 ;
  assign n25337 = n23227 ^ n788 ^ n765 ;
  assign n25338 = ( n1817 & n14744 ) | ( n1817 & ~n24427 ) | ( n14744 & ~n24427 ) ;
  assign n25343 = n15707 ^ n7839 ^ n3736 ;
  assign n25342 = n7732 ^ n6973 ^ 1'b0 ;
  assign n25339 = n1548 & n15001 ;
  assign n25340 = n9123 & ~n25339 ;
  assign n25341 = n5339 & n25340 ;
  assign n25344 = n25343 ^ n25342 ^ n25341 ;
  assign n25345 = n16107 ^ n5136 ^ n2391 ;
  assign n25346 = n25345 ^ n4812 ^ n3776 ;
  assign n25347 = n23079 ^ n12121 ^ n712 ;
  assign n25348 = n4904 & n9134 ;
  assign n25349 = n25348 ^ n1002 ^ 1'b0 ;
  assign n25350 = ( ~n4005 & n10472 ) | ( ~n4005 & n18836 ) | ( n10472 & n18836 ) ;
  assign n25351 = n9542 | n12320 ;
  assign n25352 = n25350 | n25351 ;
  assign n25353 = n5165 & n25352 ;
  assign n25354 = n16610 ^ n15237 ^ n13131 ;
  assign n25355 = n25354 ^ n10977 ^ n10194 ;
  assign n25356 = n23471 ^ n10486 ^ n8714 ;
  assign n25357 = n25342 | n25356 ;
  assign n25358 = ( n15827 & n16441 ) | ( n15827 & n19629 ) | ( n16441 & n19629 ) ;
  assign n25359 = ( n9915 & ~n12225 ) | ( n9915 & n25018 ) | ( ~n12225 & n25018 ) ;
  assign n25360 = n6324 ^ n5149 ^ 1'b0 ;
  assign n25361 = n14016 ^ n12691 ^ 1'b0 ;
  assign n25362 = n25361 ^ n12087 ^ n1732 ;
  assign n25363 = n13653 & ~n15983 ;
  assign n25364 = n3916 & n25363 ;
  assign n25365 = n23951 ^ n18907 ^ 1'b0 ;
  assign n25366 = n8756 | n25365 ;
  assign n25367 = ( n481 & n2705 ) | ( n481 & ~n13717 ) | ( n2705 & ~n13717 ) ;
  assign n25368 = ( n9096 & n10706 ) | ( n9096 & ~n25367 ) | ( n10706 & ~n25367 ) ;
  assign n25369 = n360 | n1742 ;
  assign n25370 = n25369 ^ n13767 ^ 1'b0 ;
  assign n25371 = ( n1856 & n25368 ) | ( n1856 & n25370 ) | ( n25368 & n25370 ) ;
  assign n25372 = n16769 ^ n7121 ^ 1'b0 ;
  assign n25373 = ~n25371 & n25372 ;
  assign n25374 = ~n10780 & n25373 ;
  assign n25375 = n23015 | n24322 ;
  assign n25377 = n21124 ^ n6456 ^ n5583 ;
  assign n25378 = n9560 | n10060 ;
  assign n25379 = n25377 | n25378 ;
  assign n25376 = n8175 ^ n6371 ^ n5024 ;
  assign n25380 = n25379 ^ n25376 ^ n22725 ;
  assign n25381 = n22457 ^ n13313 ^ 1'b0 ;
  assign n25382 = ( ~n5655 & n14348 ) | ( ~n5655 & n20701 ) | ( n14348 & n20701 ) ;
  assign n25383 = n25382 ^ n25297 ^ n7388 ;
  assign n25385 = n5543 ^ n4574 ^ 1'b0 ;
  assign n25386 = ~n2691 & n25385 ;
  assign n25384 = n529 | n11396 ;
  assign n25387 = n25386 ^ n25384 ^ 1'b0 ;
  assign n25388 = n2616 & ~n2991 ;
  assign n25389 = n25388 ^ n215 ^ 1'b0 ;
  assign n25390 = n25389 ^ n14628 ^ n2955 ;
  assign n25391 = n25390 ^ n3648 ^ 1'b0 ;
  assign n25392 = n10010 ^ n8256 ^ n3461 ;
  assign n25393 = n25392 ^ n20773 ^ 1'b0 ;
  assign n25394 = ~n8970 & n21143 ;
  assign n25395 = n25394 ^ n7277 ^ 1'b0 ;
  assign n25396 = n16536 & n25395 ;
  assign n25397 = n12819 ^ n10497 ^ 1'b0 ;
  assign n25398 = n16083 ^ n3146 ^ 1'b0 ;
  assign n25399 = n4177 | n25398 ;
  assign n25400 = ~n21597 & n25399 ;
  assign n25401 = ( n11260 & n18129 ) | ( n11260 & n25400 ) | ( n18129 & n25400 ) ;
  assign n25402 = ( n1907 & n7940 ) | ( n1907 & n9404 ) | ( n7940 & n9404 ) ;
  assign n25403 = n25402 ^ n1199 ^ 1'b0 ;
  assign n25404 = ( n4970 & n20389 ) | ( n4970 & n25403 ) | ( n20389 & n25403 ) ;
  assign n25405 = n14328 ^ n12624 ^ n1778 ;
  assign n25406 = ~n5923 & n8559 ;
  assign n25407 = n25406 ^ n4429 ^ 1'b0 ;
  assign n25408 = n953 | n25407 ;
  assign n25409 = n3656 | n4544 ;
  assign n25410 = n7023 & ~n25409 ;
  assign n25411 = n10185 | n15596 ;
  assign n25412 = n2236 | n25411 ;
  assign n25413 = n7645 & n19679 ;
  assign n25414 = n25413 ^ n21752 ^ 1'b0 ;
  assign n25415 = n25414 ^ n2374 ^ 1'b0 ;
  assign n25416 = n8400 ^ n7151 ^ 1'b0 ;
  assign n25417 = ( ~n14175 & n24129 ) | ( ~n14175 & n25416 ) | ( n24129 & n25416 ) ;
  assign n25418 = ~n2086 & n7359 ;
  assign n25419 = n25418 ^ n4055 ^ 1'b0 ;
  assign n25420 = ( n2928 & n8087 ) | ( n2928 & n25419 ) | ( n8087 & n25419 ) ;
  assign n25423 = n11807 & ~n22675 ;
  assign n25421 = n3764 & n25377 ;
  assign n25422 = n25421 ^ n17098 ^ 1'b0 ;
  assign n25424 = n25423 ^ n25422 ^ n22773 ;
  assign n25425 = n14413 ^ n5732 ^ n3927 ;
  assign n25426 = n8076 | n20138 ;
  assign n25427 = n25425 | n25426 ;
  assign n25428 = n6880 | n19443 ;
  assign n25429 = n25428 ^ n8298 ^ 1'b0 ;
  assign n25430 = n15360 ^ n13509 ^ n9363 ;
  assign n25431 = n2795 & n25430 ;
  assign n25432 = ( n4218 & n24368 ) | ( n4218 & n25431 ) | ( n24368 & n25431 ) ;
  assign n25433 = n25076 ^ n13102 ^ n9832 ;
  assign n25434 = ( n8519 & ~n18224 ) | ( n8519 & n21714 ) | ( ~n18224 & n21714 ) ;
  assign n25435 = ( n591 & n6699 ) | ( n591 & ~n25434 ) | ( n6699 & ~n25434 ) ;
  assign n25436 = n2803 & n14582 ;
  assign n25437 = n25436 ^ n16083 ^ 1'b0 ;
  assign n25438 = n21399 | n25437 ;
  assign n25439 = n12745 ^ n5461 ^ x91 ;
  assign n25440 = n19122 ^ n16077 ^ n1759 ;
  assign n25441 = n21007 ^ n10191 ^ 1'b0 ;
  assign n25442 = n25440 & n25441 ;
  assign n25443 = ~n5108 & n21131 ;
  assign n25444 = n25443 ^ n15970 ^ 1'b0 ;
  assign n25445 = ( n6175 & n9183 ) | ( n6175 & ~n17213 ) | ( n9183 & ~n17213 ) ;
  assign n25446 = ( n21052 & n25444 ) | ( n21052 & n25445 ) | ( n25444 & n25445 ) ;
  assign n25447 = n11091 ^ n9528 ^ n838 ;
  assign n25448 = n9064 & n16465 ;
  assign n25449 = n25448 ^ n15678 ^ 1'b0 ;
  assign n25450 = n11247 & ~n18416 ;
  assign n25451 = ( n468 & n19241 ) | ( n468 & n25450 ) | ( n19241 & n25450 ) ;
  assign n25454 = n885 & n3748 ;
  assign n25452 = ~n5791 & n6637 ;
  assign n25453 = n11248 | n25452 ;
  assign n25455 = n25454 ^ n25453 ^ 1'b0 ;
  assign n25456 = ~n1483 & n19426 ;
  assign n25457 = ~n10370 & n12327 ;
  assign n25458 = n25457 ^ n22764 ^ 1'b0 ;
  assign n25459 = ( n12547 & n14839 ) | ( n12547 & ~n25458 ) | ( n14839 & ~n25458 ) ;
  assign n25460 = n8277 | n8809 ;
  assign n25461 = n7925 & n11379 ;
  assign n25462 = ~n869 & n25461 ;
  assign n25463 = ~n6366 & n14118 ;
  assign n25464 = n25463 ^ n13382 ^ 1'b0 ;
  assign n25465 = ( n2317 & n4408 ) | ( n2317 & n5800 ) | ( n4408 & n5800 ) ;
  assign n25466 = n16273 ^ n11399 ^ 1'b0 ;
  assign n25467 = n25466 ^ n19509 ^ 1'b0 ;
  assign n25468 = n25465 & n25467 ;
  assign n25469 = ~n1378 & n25468 ;
  assign n25470 = n25469 ^ n12927 ^ 1'b0 ;
  assign n25471 = n22196 ^ n5372 ^ n1259 ;
  assign n25472 = n20369 ^ n2313 ^ 1'b0 ;
  assign n25473 = n4671 & ~n12745 ;
  assign n25474 = ~n17746 & n25473 ;
  assign n25475 = n21289 | n24968 ;
  assign n25476 = n10947 & ~n25475 ;
  assign n25477 = ( ~n10748 & n25474 ) | ( ~n10748 & n25476 ) | ( n25474 & n25476 ) ;
  assign n25478 = n19808 ^ n2286 ^ n137 ;
  assign n25479 = n25474 | n25478 ;
  assign n25480 = n9272 & n17766 ;
  assign n25481 = ~n16686 & n18257 ;
  assign n25482 = n18838 ^ n16636 ^ n12924 ;
  assign n25483 = n7859 & ~n14870 ;
  assign n25484 = n16259 ^ n7452 ^ n1779 ;
  assign n25485 = n25484 ^ n19893 ^ n9036 ;
  assign n25486 = ( n3302 & n4742 ) | ( n3302 & n19316 ) | ( n4742 & n19316 ) ;
  assign n25487 = n25486 ^ n4146 ^ 1'b0 ;
  assign n25488 = n25485 & ~n25487 ;
  assign n25489 = n14159 & ~n22767 ;
  assign n25490 = ~n15198 & n25489 ;
  assign n25491 = ( n5802 & n6673 ) | ( n5802 & ~n9290 ) | ( n6673 & ~n9290 ) ;
  assign n25492 = n20396 ^ n8346 ^ 1'b0 ;
  assign n25493 = ~n25491 & n25492 ;
  assign n25494 = n6994 ^ n5219 ^ 1'b0 ;
  assign n25495 = n2118 & n25494 ;
  assign n25496 = ~n3252 & n25495 ;
  assign n25497 = n25496 ^ n6897 ^ n3591 ;
  assign n25498 = n18610 ^ n13785 ^ n12412 ;
  assign n25501 = ( ~n2532 & n3124 ) | ( ~n2532 & n17245 ) | ( n3124 & n17245 ) ;
  assign n25499 = n1989 & n6448 ;
  assign n25500 = ~n16027 & n25499 ;
  assign n25502 = n25501 ^ n25500 ^ x26 ;
  assign n25503 = n20096 ^ n5236 ^ n2640 ;
  assign n25504 = n2078 | n20310 ;
  assign n25505 = n6305 | n25504 ;
  assign n25509 = n13931 | n21912 ;
  assign n25510 = n25509 ^ n4801 ^ 1'b0 ;
  assign n25507 = ( n6540 & ~n11766 ) | ( n6540 & n21164 ) | ( ~n11766 & n21164 ) ;
  assign n25508 = n25507 ^ n10172 ^ n2376 ;
  assign n25511 = n25510 ^ n25508 ^ n5016 ;
  assign n25506 = ~n3183 & n7340 ;
  assign n25512 = n25511 ^ n25506 ^ 1'b0 ;
  assign n25513 = n23971 ^ n13842 ^ n6623 ;
  assign n25514 = n25513 ^ n20421 ^ n11337 ;
  assign n25515 = n25514 ^ n9141 ^ 1'b0 ;
  assign n25521 = n2661 | n6705 ;
  assign n25518 = n5395 & n7825 ;
  assign n25519 = n25518 ^ n1555 ^ n364 ;
  assign n25520 = n8417 & n25519 ;
  assign n25516 = n7921 | n10704 ;
  assign n25517 = n10863 & ~n25516 ;
  assign n25522 = n25521 ^ n25520 ^ n25517 ;
  assign n25523 = n6214 ^ n888 ^ 1'b0 ;
  assign n25524 = n328 | n25523 ;
  assign n25525 = n25524 ^ n10139 ^ n1635 ;
  assign n25526 = n8105 ^ n605 ^ 1'b0 ;
  assign n25527 = n10041 & ~n25526 ;
  assign n25528 = ( n16407 & n18948 ) | ( n16407 & ~n25527 ) | ( n18948 & ~n25527 ) ;
  assign n25529 = ~n4725 & n21916 ;
  assign n25530 = n20919 ^ n13429 ^ n13129 ;
  assign n25531 = ( ~n10828 & n25529 ) | ( ~n10828 & n25530 ) | ( n25529 & n25530 ) ;
  assign n25532 = n2385 | n4374 ;
  assign n25533 = n14360 & ~n25532 ;
  assign n25534 = n5699 & n9344 ;
  assign n25535 = n25534 ^ n9478 ^ 1'b0 ;
  assign n25536 = n11846 & ~n25535 ;
  assign n25537 = n19730 & ~n24436 ;
  assign n25538 = ( n2358 & n13965 ) | ( n2358 & ~n14170 ) | ( n13965 & ~n14170 ) ;
  assign n25539 = ( n1497 & ~n12662 ) | ( n1497 & n15790 ) | ( ~n12662 & n15790 ) ;
  assign n25540 = ( n8592 & ~n24072 ) | ( n8592 & n25539 ) | ( ~n24072 & n25539 ) ;
  assign n25541 = n18795 ^ n5814 ^ 1'b0 ;
  assign n25542 = ~n6568 & n11552 ;
  assign n25543 = n25542 ^ n2546 ^ 1'b0 ;
  assign n25544 = ( n6810 & ~n11251 ) | ( n6810 & n20547 ) | ( ~n11251 & n20547 ) ;
  assign n25545 = ( n6072 & ~n25543 ) | ( n6072 & n25544 ) | ( ~n25543 & n25544 ) ;
  assign n25546 = ( n22907 & n25541 ) | ( n22907 & n25545 ) | ( n25541 & n25545 ) ;
  assign n25547 = n16366 ^ n1552 ^ 1'b0 ;
  assign n25548 = ~n7015 & n19963 ;
  assign n25549 = n25548 ^ n21039 ^ 1'b0 ;
  assign n25552 = ~n1001 & n7061 ;
  assign n25553 = n1001 & n25552 ;
  assign n25550 = n18026 ^ n413 ^ 1'b0 ;
  assign n25551 = n4172 | n25550 ;
  assign n25554 = n25553 ^ n25551 ^ 1'b0 ;
  assign n25555 = n13628 & n25554 ;
  assign n25556 = n6803 | n18004 ;
  assign n25557 = n14540 | n25556 ;
  assign n25558 = ( ~n783 & n2798 ) | ( ~n783 & n7739 ) | ( n2798 & n7739 ) ;
  assign n25559 = n25558 ^ n8420 ^ 1'b0 ;
  assign n25560 = ( ~n2513 & n9183 ) | ( ~n2513 & n16520 ) | ( n9183 & n16520 ) ;
  assign n25561 = n25560 ^ n2440 ^ 1'b0 ;
  assign n25562 = n8695 & ~n21200 ;
  assign n25563 = n25562 ^ n19699 ^ n8833 ;
  assign n25564 = n13391 ^ n6481 ^ 1'b0 ;
  assign n25565 = ( n22586 & n25563 ) | ( n22586 & n25564 ) | ( n25563 & n25564 ) ;
  assign n25566 = n9187 ^ n9081 ^ n5471 ;
  assign n25567 = n1322 & n1959 ;
  assign n25568 = n4114 & ~n5718 ;
  assign n25569 = n25568 ^ n9806 ^ 1'b0 ;
  assign n25570 = x91 & n25569 ;
  assign n25571 = n25570 ^ n4902 ^ 1'b0 ;
  assign n25572 = n767 | n22297 ;
  assign n25573 = n25572 ^ n15752 ^ 1'b0 ;
  assign n25574 = n9975 & n22713 ;
  assign n25575 = n25574 ^ n19815 ^ 1'b0 ;
  assign n25576 = n24219 ^ n20482 ^ n532 ;
  assign n25579 = n6086 | n24385 ;
  assign n25580 = n10470 & ~n25579 ;
  assign n25577 = n13871 & n15381 ;
  assign n25578 = n2894 & n25577 ;
  assign n25581 = n25580 ^ n25578 ^ 1'b0 ;
  assign n25582 = ( n7867 & ~n21330 ) | ( n7867 & n25581 ) | ( ~n21330 & n25581 ) ;
  assign n25583 = n9129 ^ n6836 ^ n6091 ;
  assign n25584 = n5507 & ~n11411 ;
  assign n25585 = ( n1443 & n15372 ) | ( n1443 & ~n25584 ) | ( n15372 & ~n25584 ) ;
  assign n25586 = n14930 ^ n10964 ^ 1'b0 ;
  assign n25589 = ~n16742 & n24501 ;
  assign n25587 = ( n2950 & ~n3375 ) | ( n2950 & n9898 ) | ( ~n3375 & n9898 ) ;
  assign n25588 = n25587 ^ n7415 ^ 1'b0 ;
  assign n25590 = n25589 ^ n25588 ^ 1'b0 ;
  assign n25591 = n4776 ^ n2492 ^ 1'b0 ;
  assign n25592 = n7104 | n25591 ;
  assign n25593 = ( ~n9170 & n10482 ) | ( ~n9170 & n25592 ) | ( n10482 & n25592 ) ;
  assign n25594 = n4647 & n25593 ;
  assign n25595 = ~n25590 & n25594 ;
  assign n25596 = n8851 & ~n8946 ;
  assign n25597 = n25596 ^ n8952 ^ 1'b0 ;
  assign n25598 = n875 | n10252 ;
  assign n25599 = ~n7705 & n20631 ;
  assign n25600 = n25052 & n25599 ;
  assign n25601 = n25600 ^ n21952 ^ n1498 ;
  assign n25602 = n17134 ^ n3816 ^ 1'b0 ;
  assign n25603 = ~n518 & n25602 ;
  assign n25604 = n5415 & n16350 ;
  assign n25605 = n25604 ^ n23971 ^ 1'b0 ;
  assign n25606 = n25603 | n25605 ;
  assign n25607 = n15655 ^ n1342 ^ 1'b0 ;
  assign n25608 = ( n5672 & n20994 ) | ( n5672 & ~n25607 ) | ( n20994 & ~n25607 ) ;
  assign n25609 = n7519 | n9264 ;
  assign n25610 = n19242 ^ n3914 ^ x29 ;
  assign n25611 = n12247 ^ n6951 ^ n1331 ;
  assign n25612 = ( n6137 & n10119 ) | ( n6137 & n25611 ) | ( n10119 & n25611 ) ;
  assign n25613 = ( n23870 & n25610 ) | ( n23870 & n25612 ) | ( n25610 & n25612 ) ;
  assign n25614 = ( n1426 & n25609 ) | ( n1426 & ~n25613 ) | ( n25609 & ~n25613 ) ;
  assign n25615 = ~n4116 & n17078 ;
  assign n25616 = ~n3300 & n25615 ;
  assign n25617 = n20609 ^ n5745 ^ 1'b0 ;
  assign n25620 = n14499 ^ n7222 ^ 1'b0 ;
  assign n25618 = n2682 | n10006 ;
  assign n25619 = n25618 ^ n5765 ^ 1'b0 ;
  assign n25621 = n25620 ^ n25619 ^ n18450 ;
  assign n25622 = ( n2712 & ~n6697 ) | ( n2712 & n25621 ) | ( ~n6697 & n25621 ) ;
  assign n25623 = n23328 ^ n6496 ^ n1404 ;
  assign n25624 = n5947 | n25623 ;
  assign n25625 = n25624 ^ n7074 ^ 1'b0 ;
  assign n25626 = n7948 ^ n6669 ^ 1'b0 ;
  assign n25627 = n9966 | n25626 ;
  assign n25628 = ( n18892 & ~n23819 ) | ( n18892 & n25627 ) | ( ~n23819 & n25627 ) ;
  assign n25629 = ( n18763 & n21575 ) | ( n18763 & n25041 ) | ( n21575 & n25041 ) ;
  assign n25630 = n9251 | n11393 ;
  assign n25631 = n25630 ^ n21707 ^ 1'b0 ;
  assign n25632 = n12174 ^ n10203 ^ n392 ;
  assign n25633 = n25632 ^ n22296 ^ 1'b0 ;
  assign n25634 = n12502 & ~n25633 ;
  assign n25635 = n1028 & ~n6578 ;
  assign n25636 = n25635 ^ n22284 ^ 1'b0 ;
  assign n25637 = n25636 ^ n5101 ^ 1'b0 ;
  assign n25638 = n16752 & ~n25637 ;
  assign n25639 = n3543 & ~n7025 ;
  assign n25640 = ( n7003 & ~n12337 ) | ( n7003 & n25639 ) | ( ~n12337 & n25639 ) ;
  assign n25641 = n19613 ^ n12010 ^ n3251 ;
  assign n25642 = ( n1566 & n7928 ) | ( n1566 & ~n25641 ) | ( n7928 & ~n25641 ) ;
  assign n25644 = n1263 | n14330 ;
  assign n25645 = ~n6750 & n25644 ;
  assign n25646 = n14568 & n25645 ;
  assign n25643 = ( ~n12009 & n13571 ) | ( ~n12009 & n16291 ) | ( n13571 & n16291 ) ;
  assign n25647 = n25646 ^ n25643 ^ n9475 ;
  assign n25648 = ( n6043 & ~n8482 ) | ( n6043 & n13938 ) | ( ~n8482 & n13938 ) ;
  assign n25649 = n18598 ^ n17386 ^ 1'b0 ;
  assign n25650 = n25649 ^ n9875 ^ x91 ;
  assign n25651 = n25650 ^ n23015 ^ 1'b0 ;
  assign n25652 = n10404 ^ n7176 ^ 1'b0 ;
  assign n25653 = ~n9938 & n25652 ;
  assign n25654 = n5504 | n25653 ;
  assign n25655 = ( n10114 & n11828 ) | ( n10114 & n25654 ) | ( n11828 & n25654 ) ;
  assign n25657 = n6964 ^ n4970 ^ n1088 ;
  assign n25656 = n5592 & n11122 ;
  assign n25658 = n25657 ^ n25656 ^ 1'b0 ;
  assign n25660 = n6957 ^ n6947 ^ n2487 ;
  assign n25659 = n11482 & n12655 ;
  assign n25661 = n25660 ^ n25659 ^ 1'b0 ;
  assign n25662 = n6223 & ~n14932 ;
  assign n25663 = ( n5548 & n13197 ) | ( n5548 & n25662 ) | ( n13197 & n25662 ) ;
  assign n25664 = n12138 ^ n6131 ^ 1'b0 ;
  assign n25665 = n25663 | n25664 ;
  assign n25666 = n11224 ^ n5414 ^ 1'b0 ;
  assign n25668 = n3730 ^ n2728 ^ 1'b0 ;
  assign n25667 = ( n2655 & n9208 ) | ( n2655 & ~n11869 ) | ( n9208 & ~n11869 ) ;
  assign n25669 = n25668 ^ n25667 ^ 1'b0 ;
  assign n25670 = n21826 ^ n5946 ^ 1'b0 ;
  assign n25671 = ( n5350 & n21714 ) | ( n5350 & n25670 ) | ( n21714 & n25670 ) ;
  assign n25672 = ( n4039 & n4578 ) | ( n4039 & ~n15713 ) | ( n4578 & ~n15713 ) ;
  assign n25673 = ( ~n432 & n7102 ) | ( ~n432 & n25672 ) | ( n7102 & n25672 ) ;
  assign n25674 = n7874 ^ n5900 ^ n2923 ;
  assign n25675 = n23323 ^ n19398 ^ 1'b0 ;
  assign n25678 = n23916 ^ n21466 ^ n18149 ;
  assign n25676 = ~n4233 & n19373 ;
  assign n25677 = ~n3141 & n25676 ;
  assign n25679 = n25678 ^ n25677 ^ 1'b0 ;
  assign n25680 = n17620 & n18369 ;
  assign n25681 = ~n7185 & n25680 ;
  assign n25682 = n25681 ^ n10771 ^ 1'b0 ;
  assign n25683 = n24886 ^ n15911 ^ n1182 ;
  assign n25684 = ~n8621 & n24471 ;
  assign n25685 = n25684 ^ n3995 ^ 1'b0 ;
  assign n25686 = n24219 | n25685 ;
  assign n25687 = ( n10936 & n17201 ) | ( n10936 & n25686 ) | ( n17201 & n25686 ) ;
  assign n25689 = n6842 & n9724 ;
  assign n25690 = n25689 ^ n5269 ^ 1'b0 ;
  assign n25688 = ( n2278 & n15425 ) | ( n2278 & ~n18883 ) | ( n15425 & ~n18883 ) ;
  assign n25691 = n25690 ^ n25688 ^ 1'b0 ;
  assign n25692 = n24434 ^ n21519 ^ n13383 ;
  assign n25693 = n1253 | n13908 ;
  assign n25694 = n13132 | n25693 ;
  assign n25695 = n14604 ^ n2968 ^ 1'b0 ;
  assign n25696 = ~x35 & n1344 ;
  assign n25697 = n1759 | n12553 ;
  assign n25698 = n25697 ^ n1922 ^ 1'b0 ;
  assign n25699 = n25698 ^ n7478 ^ n4002 ;
  assign n25700 = ( n2510 & n25696 ) | ( n2510 & n25699 ) | ( n25696 & n25699 ) ;
  assign n25701 = n5864 & n8408 ;
  assign n25702 = ( n11888 & n13504 ) | ( n11888 & ~n25701 ) | ( n13504 & ~n25701 ) ;
  assign n25703 = n14412 ^ n6043 ^ 1'b0 ;
  assign n25704 = n231 | n1134 ;
  assign n25705 = n25704 ^ n317 ^ 1'b0 ;
  assign n25706 = ( n8383 & ~n19716 ) | ( n8383 & n25705 ) | ( ~n19716 & n25705 ) ;
  assign n25707 = n3913 ^ n2850 ^ n667 ;
  assign n25708 = ( x38 & ~n8725 ) | ( x38 & n25707 ) | ( ~n8725 & n25707 ) ;
  assign n25709 = n16265 ^ n12297 ^ 1'b0 ;
  assign n25710 = ~n2579 & n25709 ;
  assign n25711 = n25710 ^ n22735 ^ 1'b0 ;
  assign n25712 = n24731 | n25711 ;
  assign n25713 = ~n10499 & n21443 ;
  assign n25714 = n24994 & n25713 ;
  assign n25715 = ( n869 & n2089 ) | ( n869 & n5923 ) | ( n2089 & n5923 ) ;
  assign n25716 = n20119 ^ n7342 ^ n2583 ;
  assign n25717 = ~n751 & n20295 ;
  assign n25718 = ( ~n25715 & n25716 ) | ( ~n25715 & n25717 ) | ( n25716 & n25717 ) ;
  assign n25719 = ( ~n1296 & n1828 ) | ( ~n1296 & n16807 ) | ( n1828 & n16807 ) ;
  assign n25720 = n24332 | n25719 ;
  assign n25721 = n17408 ^ n15291 ^ n2296 ;
  assign n25722 = n25721 ^ n18348 ^ n13430 ;
  assign n25723 = n10922 ^ n7472 ^ n6905 ;
  assign n25727 = n9087 & n10447 ;
  assign n25724 = ~n1577 & n6783 ;
  assign n25725 = n25724 ^ n179 ^ 1'b0 ;
  assign n25726 = ( ~n313 & n6001 ) | ( ~n313 & n25725 ) | ( n6001 & n25725 ) ;
  assign n25728 = n25727 ^ n25726 ^ 1'b0 ;
  assign n25729 = n14966 | n22426 ;
  assign n25730 = n16238 | n25729 ;
  assign n25731 = n25730 ^ n437 ^ 1'b0 ;
  assign n25732 = n6411 & n25731 ;
  assign n25733 = n5108 | n5453 ;
  assign n25734 = n12308 & ~n25733 ;
  assign n25735 = ( n643 & n13457 ) | ( n643 & n16128 ) | ( n13457 & n16128 ) ;
  assign n25736 = n23508 ^ n2677 ^ 1'b0 ;
  assign n25737 = n25736 ^ n20865 ^ 1'b0 ;
  assign n25738 = n25735 & ~n25737 ;
  assign n25739 = n16436 ^ n12139 ^ n5061 ;
  assign n25740 = n25739 ^ n3292 ^ n1113 ;
  assign n25741 = n25740 ^ n21232 ^ 1'b0 ;
  assign n25742 = n3274 & ~n13032 ;
  assign n25743 = ~n14964 & n25742 ;
  assign n25744 = x87 & n6228 ;
  assign n25745 = n25744 ^ n14060 ^ 1'b0 ;
  assign n25746 = n25745 ^ n17302 ^ n921 ;
  assign n25747 = n337 & ~n25746 ;
  assign n25748 = n25743 & n25747 ;
  assign n25749 = n25748 ^ n25588 ^ 1'b0 ;
  assign n25750 = n24582 ^ n22958 ^ n6754 ;
  assign n25751 = ( ~n14960 & n16499 ) | ( ~n14960 & n17434 ) | ( n16499 & n17434 ) ;
  assign n25752 = ( n12028 & ~n21695 ) | ( n12028 & n25751 ) | ( ~n21695 & n25751 ) ;
  assign n25753 = ( n3742 & ~n15600 ) | ( n3742 & n17526 ) | ( ~n15600 & n17526 ) ;
  assign n25754 = ( ~n19811 & n20695 ) | ( ~n19811 & n25753 ) | ( n20695 & n25753 ) ;
  assign n25755 = n17618 ^ n7823 ^ n7791 ;
  assign n25756 = n25755 ^ n17509 ^ 1'b0 ;
  assign n25757 = n21046 ^ n7317 ^ 1'b0 ;
  assign n25759 = n2014 | n9391 ;
  assign n25758 = ~n3319 & n5405 ;
  assign n25760 = n25759 ^ n25758 ^ 1'b0 ;
  assign n25761 = ( ~n7030 & n10778 ) | ( ~n7030 & n11073 ) | ( n10778 & n11073 ) ;
  assign n25762 = n25761 ^ n18049 ^ 1'b0 ;
  assign n25763 = n3877 & n25762 ;
  assign n25764 = n1493 & n11885 ;
  assign n25765 = n25764 ^ n4932 ^ 1'b0 ;
  assign n25766 = n16619 ^ n13601 ^ n8439 ;
  assign n25767 = n12934 ^ n10767 ^ 1'b0 ;
  assign n25771 = n986 & ~n3629 ;
  assign n25772 = n25771 ^ n4268 ^ 1'b0 ;
  assign n25768 = n9532 & ~n18145 ;
  assign n25769 = n286 & n25768 ;
  assign n25770 = n25769 ^ n12449 ^ 1'b0 ;
  assign n25773 = n25772 ^ n25770 ^ n1785 ;
  assign n25774 = ~n9246 & n22378 ;
  assign n25775 = ~n5822 & n25774 ;
  assign n25776 = ( ~n5900 & n7040 ) | ( ~n5900 & n9242 ) | ( n7040 & n9242 ) ;
  assign n25777 = n9838 ^ n5177 ^ 1'b0 ;
  assign n25778 = n25776 & n25777 ;
  assign n25780 = ( n3977 & n6991 ) | ( n3977 & n8623 ) | ( n6991 & n8623 ) ;
  assign n25779 = n11266 ^ n7920 ^ n7185 ;
  assign n25781 = n25780 ^ n25779 ^ 1'b0 ;
  assign n25782 = ( n9521 & n16750 ) | ( n9521 & n25781 ) | ( n16750 & n25781 ) ;
  assign n25783 = n25778 & n25782 ;
  assign n25784 = ( n3709 & n13169 ) | ( n3709 & n15281 ) | ( n13169 & n15281 ) ;
  assign n25785 = n25784 ^ n4645 ^ 1'b0 ;
  assign n25786 = n15664 | n25785 ;
  assign n25787 = n6124 ^ n4154 ^ 1'b0 ;
  assign n25788 = ~n25786 & n25787 ;
  assign n25789 = n23485 ^ n23379 ^ n18912 ;
  assign n25790 = n25478 ^ n20976 ^ n20886 ;
  assign n25791 = n14318 ^ n4202 ^ 1'b0 ;
  assign n25792 = n25791 ^ n15903 ^ n3706 ;
  assign n25793 = n7496 ^ n4321 ^ 1'b0 ;
  assign n25794 = n13048 | n19513 ;
  assign n25795 = n10316 | n25794 ;
  assign n25796 = ~n7348 & n25795 ;
  assign n25797 = n6139 & n25796 ;
  assign n25798 = n13253 ^ n4657 ^ 1'b0 ;
  assign n25799 = ~n7568 & n25798 ;
  assign n25800 = n16864 ^ n9176 ^ 1'b0 ;
  assign n25801 = n1893 & n25800 ;
  assign n25802 = ( n1791 & ~n2203 ) | ( n1791 & n25801 ) | ( ~n2203 & n25801 ) ;
  assign n25803 = n2733 & n25802 ;
  assign n25804 = ~n25799 & n25803 ;
  assign n25805 = n7732 ^ n1113 ^ 1'b0 ;
  assign n25806 = n1613 & ~n5314 ;
  assign n25807 = n25806 ^ n10374 ^ 1'b0 ;
  assign n25808 = n25807 ^ n14859 ^ n2526 ;
  assign n25809 = n25808 ^ n17189 ^ n5568 ;
  assign n25810 = n16843 ^ n5601 ^ n5207 ;
  assign n25811 = ~n19593 & n25810 ;
  assign n25812 = n19239 ^ n18108 ^ 1'b0 ;
  assign n25813 = ( ~n13214 & n21492 ) | ( ~n13214 & n25049 ) | ( n21492 & n25049 ) ;
  assign n25814 = ( n6301 & n8391 ) | ( n6301 & ~n25813 ) | ( n8391 & ~n25813 ) ;
  assign n25815 = n9061 ^ n3950 ^ 1'b0 ;
  assign n25816 = n12375 ^ n6324 ^ 1'b0 ;
  assign n25817 = n25815 | n25816 ;
  assign n25818 = n25817 ^ n16332 ^ n4993 ;
  assign n25819 = n19734 ^ n6948 ^ 1'b0 ;
  assign n25820 = ~n3280 & n21674 ;
  assign n25822 = n23971 ^ n12802 ^ n11387 ;
  assign n25821 = ( n20320 & ~n20526 ) | ( n20320 & n24818 ) | ( ~n20526 & n24818 ) ;
  assign n25823 = n25822 ^ n25821 ^ n6986 ;
  assign n25824 = ~n3043 & n7055 ;
  assign n25825 = ~n25823 & n25824 ;
  assign n25826 = n18639 ^ n16486 ^ n11429 ;
  assign n25827 = ( n4985 & ~n12027 ) | ( n4985 & n23275 ) | ( ~n12027 & n23275 ) ;
  assign n25828 = n25827 ^ n18568 ^ n12268 ;
  assign n25829 = n24013 ^ n2212 ^ n756 ;
  assign n25830 = ( n7414 & ~n8273 ) | ( n7414 & n14591 ) | ( ~n8273 & n14591 ) ;
  assign n25831 = n25830 ^ n10308 ^ n2076 ;
  assign n25832 = n25831 ^ n25137 ^ 1'b0 ;
  assign n25833 = n7248 ^ n6153 ^ 1'b0 ;
  assign n25834 = n1250 & n1558 ;
  assign n25835 = n25834 ^ n24140 ^ 1'b0 ;
  assign n25836 = n1289 & ~n25835 ;
  assign n25837 = n25836 ^ n9312 ^ 1'b0 ;
  assign n25838 = n4537 | n6954 ;
  assign n25839 = n25838 ^ n1418 ^ 1'b0 ;
  assign n25840 = n8817 ^ n8699 ^ x91 ;
  assign n25841 = n6086 & n25840 ;
  assign n25842 = n25657 ^ n19381 ^ n2736 ;
  assign n25844 = n3376 ^ n1945 ^ n1102 ;
  assign n25843 = n19338 ^ n18414 ^ n310 ;
  assign n25845 = n25844 ^ n25843 ^ n1286 ;
  assign n25846 = n8968 ^ n8171 ^ 1'b0 ;
  assign n25847 = ~n11361 & n25846 ;
  assign n25848 = n24240 ^ n2633 ^ 1'b0 ;
  assign n25849 = ( n2778 & n13478 ) | ( n2778 & n25848 ) | ( n13478 & n25848 ) ;
  assign n25850 = n25849 ^ n9162 ^ n2653 ;
  assign n25851 = ( ~n4421 & n18011 ) | ( ~n4421 & n25850 ) | ( n18011 & n25850 ) ;
  assign n25852 = n4696 | n25138 ;
  assign n25853 = n3312 & ~n25852 ;
  assign n25854 = n1999 | n9454 ;
  assign n25855 = n25854 ^ n12856 ^ 1'b0 ;
  assign n25856 = n3255 | n21635 ;
  assign n25857 = n25856 ^ n10690 ^ 1'b0 ;
  assign n25858 = n2498 | n23248 ;
  assign n25859 = n3678 | n25858 ;
  assign n25860 = n23724 ^ n13900 ^ n5526 ;
  assign n25861 = ~n179 & n13736 ;
  assign n25862 = n25860 & n25861 ;
  assign n25863 = ( n13273 & n14398 ) | ( n13273 & ~n25862 ) | ( n14398 & ~n25862 ) ;
  assign n25864 = n2516 ^ n1310 ^ n1225 ;
  assign n25865 = n25864 ^ n17837 ^ n13949 ;
  assign n25866 = n12066 ^ n896 ^ n805 ;
  assign n25867 = n25866 ^ n24935 ^ n18562 ;
  assign n25868 = n6312 ^ n3220 ^ 1'b0 ;
  assign n25869 = n11429 & ~n25868 ;
  assign n25870 = n22244 ^ n3622 ^ 1'b0 ;
  assign n25871 = n1463 & ~n25870 ;
  assign n25872 = ( n317 & ~n25869 ) | ( n317 & n25871 ) | ( ~n25869 & n25871 ) ;
  assign n25873 = ( n4442 & n6361 ) | ( n4442 & ~n8769 ) | ( n6361 & ~n8769 ) ;
  assign n25874 = n25873 ^ n9788 ^ 1'b0 ;
  assign n25875 = n6535 | n25874 ;
  assign n25876 = ( ~n6968 & n7677 ) | ( ~n6968 & n18639 ) | ( n7677 & n18639 ) ;
  assign n25877 = n19595 ^ n9286 ^ n3484 ;
  assign n25878 = n5332 & ~n11110 ;
  assign n25879 = n25878 ^ n3072 ^ n768 ;
  assign n25880 = ~n22535 & n25879 ;
  assign n25881 = n13160 ^ n4045 ^ x123 ;
  assign n25883 = n6807 & n12009 ;
  assign n25884 = n10401 & n25883 ;
  assign n25882 = ( n186 & ~n1837 ) | ( n186 & n8780 ) | ( ~n1837 & n8780 ) ;
  assign n25885 = n25884 ^ n25882 ^ 1'b0 ;
  assign n25886 = n10475 & ~n13298 ;
  assign n25887 = n24205 & n25886 ;
  assign n25888 = ( ~n20921 & n25885 ) | ( ~n20921 & n25887 ) | ( n25885 & n25887 ) ;
  assign n25889 = n17344 ^ n7884 ^ n2916 ;
  assign n25890 = ~n3103 & n25889 ;
  assign n25891 = ~n13217 & n25890 ;
  assign n25892 = n25891 ^ n24491 ^ 1'b0 ;
  assign n25893 = n9189 ^ n1081 ^ 1'b0 ;
  assign n25894 = n13204 & n25893 ;
  assign n25895 = ~n2477 & n4002 ;
  assign n25897 = ( n12003 & n19112 ) | ( n12003 & n22749 ) | ( n19112 & n22749 ) ;
  assign n25896 = n9764 | n11952 ;
  assign n25898 = n25897 ^ n25896 ^ 1'b0 ;
  assign n25899 = n1623 | n6568 ;
  assign n25900 = n1873 & ~n2424 ;
  assign n25901 = n1025 & ~n22450 ;
  assign n25902 = n25901 ^ n9260 ^ 1'b0 ;
  assign n25903 = n23789 ^ n11142 ^ 1'b0 ;
  assign n25904 = ( ~n1519 & n17836 ) | ( ~n1519 & n25903 ) | ( n17836 & n25903 ) ;
  assign n25905 = ( n2824 & n15525 ) | ( n2824 & n15588 ) | ( n15525 & n15588 ) ;
  assign n25906 = ( n9017 & n13276 ) | ( n9017 & ~n21891 ) | ( n13276 & ~n21891 ) ;
  assign n25909 = n468 & n2381 ;
  assign n25908 = n6246 & n25510 ;
  assign n25907 = n16001 ^ n12321 ^ n11435 ;
  assign n25910 = n25909 ^ n25908 ^ n25907 ;
  assign n25912 = ( ~n539 & n5470 ) | ( ~n539 & n6038 ) | ( n5470 & n6038 ) ;
  assign n25911 = n10061 & n17825 ;
  assign n25913 = n25912 ^ n25911 ^ 1'b0 ;
  assign n25914 = n12231 & ~n25913 ;
  assign n25915 = n16924 ^ n14139 ^ n7125 ;
  assign n25916 = n25915 ^ n11500 ^ n9570 ;
  assign n25917 = n3236 & n25916 ;
  assign n25918 = ( n1836 & n3452 ) | ( n1836 & ~n11579 ) | ( n3452 & ~n11579 ) ;
  assign n25919 = n7599 & ~n25918 ;
  assign n25920 = ~n15546 & n25919 ;
  assign n25921 = n13214 ^ n7113 ^ n3459 ;
  assign n25922 = n25921 ^ n22366 ^ n2456 ;
  assign n25923 = ( n7812 & ~n25920 ) | ( n7812 & n25922 ) | ( ~n25920 & n25922 ) ;
  assign n25924 = n23186 ^ n11165 ^ n5983 ;
  assign n25925 = n11627 & n24692 ;
  assign n25926 = n25925 ^ n25609 ^ 1'b0 ;
  assign n25927 = n25926 ^ n8647 ^ 1'b0 ;
  assign n25935 = n15285 ^ n1839 ^ 1'b0 ;
  assign n25933 = ~n3710 & n13776 ;
  assign n25934 = n794 & ~n25933 ;
  assign n25928 = n1543 & n21285 ;
  assign n25929 = n25928 ^ n10928 ^ 1'b0 ;
  assign n25930 = n4122 & ~n25929 ;
  assign n25931 = ~n5019 & n25930 ;
  assign n25932 = n25931 ^ n11096 ^ 1'b0 ;
  assign n25936 = n25935 ^ n25934 ^ n25932 ;
  assign n25937 = ( n6293 & n10922 ) | ( n6293 & ~n13335 ) | ( n10922 & ~n13335 ) ;
  assign n25938 = n25937 ^ n23576 ^ n1062 ;
  assign n25939 = n5577 & n8721 ;
  assign n25940 = n11171 & n25939 ;
  assign n25941 = n17909 ^ n15408 ^ 1'b0 ;
  assign n25947 = ~n2252 & n2864 ;
  assign n25948 = ( n9159 & n13727 ) | ( n9159 & n25947 ) | ( n13727 & n25947 ) ;
  assign n25942 = n15315 ^ n13873 ^ 1'b0 ;
  assign n25943 = ~n1261 & n25942 ;
  assign n25944 = ~n1243 & n25943 ;
  assign n25945 = n25944 ^ n551 ^ 1'b0 ;
  assign n25946 = n14765 | n25945 ;
  assign n25949 = n25948 ^ n25946 ^ n11224 ;
  assign n25950 = ( ~n9299 & n15429 ) | ( ~n9299 & n25949 ) | ( n15429 & n25949 ) ;
  assign n25951 = n1079 & ~n10355 ;
  assign n25952 = n16773 | n20211 ;
  assign n25953 = n12971 ^ n3665 ^ n981 ;
  assign n25954 = ( n2069 & n20238 ) | ( n2069 & ~n25953 ) | ( n20238 & ~n25953 ) ;
  assign n25955 = n5810 & ~n10024 ;
  assign n25956 = n25955 ^ n5905 ^ n3028 ;
  assign n25957 = n1394 | n8625 ;
  assign n25958 = n4409 & ~n25957 ;
  assign n25959 = n21469 ^ n5635 ^ 1'b0 ;
  assign n25960 = n1796 & ~n2151 ;
  assign n25961 = ~n4951 & n25960 ;
  assign n25962 = n4722 | n25961 ;
  assign n25963 = n14794 | n25962 ;
  assign n25964 = n3225 | n3366 ;
  assign n25965 = n25964 ^ n2299 ^ 1'b0 ;
  assign n25966 = n25965 ^ n11836 ^ 1'b0 ;
  assign n25967 = n11014 | n25966 ;
  assign n25968 = n25967 ^ n17954 ^ 1'b0 ;
  assign n25969 = n25963 & n25968 ;
  assign n25971 = ( n2691 & n14262 ) | ( n2691 & n20137 ) | ( n14262 & n20137 ) ;
  assign n25970 = n3473 | n5887 ;
  assign n25972 = n25971 ^ n25970 ^ 1'b0 ;
  assign n25973 = n2290 & n15616 ;
  assign n25974 = n14231 ^ n9970 ^ n1172 ;
  assign n25975 = ( n3138 & ~n6483 ) | ( n3138 & n24269 ) | ( ~n6483 & n24269 ) ;
  assign n25976 = n9377 & ~n13026 ;
  assign n25977 = ~n13092 & n25976 ;
  assign n25978 = n20137 & ~n25977 ;
  assign n25979 = ( ~n19524 & n25975 ) | ( ~n19524 & n25978 ) | ( n25975 & n25978 ) ;
  assign n25980 = n9927 & ~n14656 ;
  assign n25981 = n25980 ^ n1628 ^ 1'b0 ;
  assign n25982 = ( n3083 & n19636 ) | ( n3083 & ~n25981 ) | ( n19636 & ~n25981 ) ;
  assign n25983 = n8012 | n20104 ;
  assign n25984 = n1843 | n25983 ;
  assign n25985 = n2245 & n25984 ;
  assign n25986 = n7205 | n13449 ;
  assign n25987 = n428 | n25986 ;
  assign n25988 = n5062 & ~n25329 ;
  assign n25989 = n14078 ^ n8592 ^ n2338 ;
  assign n25990 = ( n7687 & n11286 ) | ( n7687 & ~n12897 ) | ( n11286 & ~n12897 ) ;
  assign n25991 = n25990 ^ n5047 ^ n2570 ;
  assign n25992 = ( n15120 & n23948 ) | ( n15120 & ~n25991 ) | ( n23948 & ~n25991 ) ;
  assign n25993 = n7637 | n25992 ;
  assign n25994 = n25993 ^ n12701 ^ n7741 ;
  assign n25995 = n25994 ^ n23397 ^ n14275 ;
  assign n25996 = ~n1370 & n18011 ;
  assign n25997 = ( n3749 & n10273 ) | ( n3749 & n25996 ) | ( n10273 & n25996 ) ;
  assign n25998 = n25997 ^ n24609 ^ n14094 ;
  assign n26001 = ( ~n3735 & n5224 ) | ( ~n3735 & n8038 ) | ( n5224 & n8038 ) ;
  assign n25999 = n20842 ^ n11873 ^ 1'b0 ;
  assign n26000 = n9253 & n25999 ;
  assign n26002 = n26001 ^ n26000 ^ n7022 ;
  assign n26003 = n26002 ^ n24407 ^ 1'b0 ;
  assign n26004 = n20114 ^ n9619 ^ n1203 ;
  assign n26005 = ( n7290 & n8693 ) | ( n7290 & ~n26004 ) | ( n8693 & ~n26004 ) ;
  assign n26006 = n24723 ^ n6984 ^ n3628 ;
  assign n26007 = n26006 ^ n22788 ^ n2011 ;
  assign n26008 = ( n12054 & n26005 ) | ( n12054 & ~n26007 ) | ( n26005 & ~n26007 ) ;
  assign n26009 = n15473 ^ n3848 ^ 1'b0 ;
  assign n26010 = n12126 & ~n26009 ;
  assign n26011 = n3195 & ~n18158 ;
  assign n26012 = n22477 ^ n1088 ^ 1'b0 ;
  assign n26013 = n17279 ^ n14656 ^ n13752 ;
  assign n26014 = n17780 ^ n4575 ^ 1'b0 ;
  assign n26015 = n21808 & n26014 ;
  assign n26017 = ( ~n863 & n6949 ) | ( ~n863 & n21167 ) | ( n6949 & n21167 ) ;
  assign n26016 = n17052 & ~n22362 ;
  assign n26018 = n26017 ^ n26016 ^ 1'b0 ;
  assign n26019 = ( n17992 & n26015 ) | ( n17992 & ~n26018 ) | ( n26015 & ~n26018 ) ;
  assign n26020 = n3117 & ~n8590 ;
  assign n26021 = n9530 & n26020 ;
  assign n26022 = n2192 | n26021 ;
  assign n26023 = n20624 & ~n26022 ;
  assign n26024 = n26023 ^ n6413 ^ 1'b0 ;
  assign n26025 = n5133 & n24458 ;
  assign n26026 = n26025 ^ n13380 ^ n684 ;
  assign n26027 = n8770 & ~n12710 ;
  assign n26028 = ~n21962 & n26027 ;
  assign n26029 = n25878 ^ n11968 ^ 1'b0 ;
  assign n26030 = ~n8431 & n26029 ;
  assign n26031 = n9797 | n24033 ;
  assign n26032 = n13217 | n26031 ;
  assign n26033 = n26032 ^ n21252 ^ 1'b0 ;
  assign n26034 = n7689 & ~n26033 ;
  assign n26035 = n2701 ^ n1871 ^ 1'b0 ;
  assign n26036 = ~n4418 & n26035 ;
  assign n26037 = n26036 ^ n24465 ^ n12170 ;
  assign n26038 = n19909 ^ n11119 ^ n1225 ;
  assign n26039 = n26038 ^ n7046 ^ n6963 ;
  assign n26040 = n26039 ^ n24890 ^ n23927 ;
  assign n26042 = n4401 | n6262 ;
  assign n26043 = n26042 ^ n4610 ^ 1'b0 ;
  assign n26041 = ( n5985 & ~n16774 ) | ( n5985 & n18351 ) | ( ~n16774 & n18351 ) ;
  assign n26044 = n26043 ^ n26041 ^ n24731 ;
  assign n26045 = ( n3702 & n12747 ) | ( n3702 & ~n24119 ) | ( n12747 & ~n24119 ) ;
  assign n26046 = x67 & n7932 ;
  assign n26047 = n21393 ^ n12470 ^ 1'b0 ;
  assign n26048 = n10301 | n26047 ;
  assign n26049 = n15276 ^ n11395 ^ 1'b0 ;
  assign n26050 = n8241 & ~n9632 ;
  assign n26051 = n26050 ^ n15892 ^ 1'b0 ;
  assign n26052 = n19036 & n26051 ;
  assign n26053 = n26052 ^ n6028 ^ 1'b0 ;
  assign n26056 = n8753 & ~n16914 ;
  assign n26054 = n7781 ^ n6317 ^ n3476 ;
  assign n26055 = ~n15090 & n26054 ;
  assign n26057 = n26056 ^ n26055 ^ n22441 ;
  assign n26058 = n2900 | n15809 ;
  assign n26059 = ( n2321 & ~n7379 ) | ( n2321 & n26058 ) | ( ~n7379 & n26058 ) ;
  assign n26060 = n26059 ^ n19454 ^ n8690 ;
  assign n26061 = ~n4279 & n26060 ;
  assign n26062 = n26061 ^ n1234 ^ 1'b0 ;
  assign n26063 = ( n5636 & n17806 ) | ( n5636 & ~n26062 ) | ( n17806 & ~n26062 ) ;
  assign n26064 = n21275 ^ n8064 ^ n4072 ;
  assign n26065 = ( n297 & n2470 ) | ( n297 & ~n6439 ) | ( n2470 & ~n6439 ) ;
  assign n26066 = n598 & ~n9362 ;
  assign n26067 = ~n21156 & n26066 ;
  assign n26068 = ( n1816 & n16715 ) | ( n1816 & n26067 ) | ( n16715 & n26067 ) ;
  assign n26069 = n13018 ^ n7715 ^ 1'b0 ;
  assign n26071 = ( ~n4282 & n6235 ) | ( ~n4282 & n6985 ) | ( n6235 & n6985 ) ;
  assign n26072 = n10442 | n26071 ;
  assign n26073 = n26072 ^ n14779 ^ 1'b0 ;
  assign n26074 = ~n5301 & n26073 ;
  assign n26075 = n26074 ^ n15309 ^ 1'b0 ;
  assign n26070 = ~n14315 & n16418 ;
  assign n26076 = n26075 ^ n26070 ^ 1'b0 ;
  assign n26077 = ~n4700 & n13407 ;
  assign n26078 = n9676 ^ n2279 ^ n1233 ;
  assign n26079 = n8701 ^ n3846 ^ 1'b0 ;
  assign n26080 = n17709 & n26079 ;
  assign n26081 = ( ~n18014 & n18356 ) | ( ~n18014 & n19716 ) | ( n18356 & n19716 ) ;
  assign n26082 = n26081 ^ n23452 ^ 1'b0 ;
  assign n26083 = n2325 & ~n26082 ;
  assign n26084 = ( ~n12875 & n26080 ) | ( ~n12875 & n26083 ) | ( n26080 & n26083 ) ;
  assign n26085 = n1492 & n3707 ;
  assign n26086 = ~n6060 & n15855 ;
  assign n26087 = n26086 ^ n7365 ^ 1'b0 ;
  assign n26088 = n26087 ^ n12219 ^ n6698 ;
  assign n26089 = ( n8028 & n21128 ) | ( n8028 & n26088 ) | ( n21128 & n26088 ) ;
  assign n26090 = n19708 ^ n12025 ^ 1'b0 ;
  assign n26091 = n18563 & ~n25933 ;
  assign n26092 = n1867 & ~n4720 ;
  assign n26093 = n26092 ^ x80 ^ 1'b0 ;
  assign n26094 = ~n6948 & n26015 ;
  assign n26095 = ~n24374 & n26094 ;
  assign n26096 = n13541 ^ n10567 ^ n10232 ;
  assign n26099 = n21671 ^ n19021 ^ n6750 ;
  assign n26100 = ( ~n988 & n10555 ) | ( ~n988 & n26099 ) | ( n10555 & n26099 ) ;
  assign n26101 = ( n1357 & n5860 ) | ( n1357 & ~n6775 ) | ( n5860 & ~n6775 ) ;
  assign n26102 = n26101 ^ n21349 ^ n16651 ;
  assign n26103 = ( ~n12579 & n26100 ) | ( ~n12579 & n26102 ) | ( n26100 & n26102 ) ;
  assign n26097 = n10909 ^ n7205 ^ n4088 ;
  assign n26098 = ( n3452 & n19804 ) | ( n3452 & n26097 ) | ( n19804 & n26097 ) ;
  assign n26104 = n26103 ^ n26098 ^ n13018 ;
  assign n26105 = n16236 & n22597 ;
  assign n26106 = n18945 ^ n12028 ^ n929 ;
  assign n26107 = ( ~n4733 & n14235 ) | ( ~n4733 & n15051 ) | ( n14235 & n15051 ) ;
  assign n26108 = n26106 & ~n26107 ;
  assign n26109 = n12836 ^ n10830 ^ n3374 ;
  assign n26110 = n25259 | n25865 ;
  assign n26111 = n20335 | n26110 ;
  assign n26112 = n13139 ^ n553 ^ 1'b0 ;
  assign n26113 = ( n10377 & ~n10737 ) | ( n10377 & n20135 ) | ( ~n10737 & n20135 ) ;
  assign n26114 = n13083 ^ n3792 ^ 1'b0 ;
  assign n26115 = ( n9454 & ~n13934 ) | ( n9454 & n18289 ) | ( ~n13934 & n18289 ) ;
  assign n26116 = n9819 | n26115 ;
  assign n26117 = n26116 ^ n14227 ^ 1'b0 ;
  assign n26118 = ~n18669 & n26117 ;
  assign n26119 = n21410 ^ n17443 ^ n2200 ;
  assign n26120 = ( ~n26114 & n26118 ) | ( ~n26114 & n26119 ) | ( n26118 & n26119 ) ;
  assign n26121 = n26120 ^ n16585 ^ n6928 ;
  assign n26122 = ( ~n335 & n23746 ) | ( ~n335 & n25367 ) | ( n23746 & n25367 ) ;
  assign n26123 = ( n17478 & ~n18280 ) | ( n17478 & n26122 ) | ( ~n18280 & n26122 ) ;
  assign n26126 = n13370 ^ n11536 ^ n1582 ;
  assign n26127 = n26126 ^ n15441 ^ n10617 ;
  assign n26128 = n25275 & ~n26127 ;
  assign n26124 = n896 & ~n2697 ;
  assign n26125 = ~n3534 & n26124 ;
  assign n26129 = n26128 ^ n26125 ^ n19552 ;
  assign n26130 = n4549 & n14071 ;
  assign n26131 = ( n1706 & n13414 ) | ( n1706 & ~n26130 ) | ( n13414 & ~n26130 ) ;
  assign n26132 = n13941 & n23110 ;
  assign n26133 = n26132 ^ n2590 ^ 1'b0 ;
  assign n26134 = n10727 & n11473 ;
  assign n26135 = n5738 & n26134 ;
  assign n26140 = n3070 ^ n2882 ^ 1'b0 ;
  assign n26137 = n11240 ^ n6558 ^ n4639 ;
  assign n26136 = n16924 ^ n15080 ^ n5904 ;
  assign n26138 = n26137 ^ n26136 ^ n3441 ;
  assign n26139 = ( ~n3579 & n17841 ) | ( ~n3579 & n26138 ) | ( n17841 & n26138 ) ;
  assign n26141 = n26140 ^ n26139 ^ n10671 ;
  assign n26142 = n14895 & ~n25390 ;
  assign n26143 = n24568 ^ n8795 ^ n763 ;
  assign n26144 = n3329 ^ n1582 ^ 1'b0 ;
  assign n26145 = n4180 & n26144 ;
  assign n26146 = n26145 ^ n6767 ^ n4268 ;
  assign n26147 = n2679 & n6672 ;
  assign n26148 = n26147 ^ n12722 ^ 1'b0 ;
  assign n26149 = ( n8385 & ~n13532 ) | ( n8385 & n18614 ) | ( ~n13532 & n18614 ) ;
  assign n26150 = n26149 ^ n23890 ^ n11218 ;
  assign n26151 = ( n26146 & ~n26148 ) | ( n26146 & n26150 ) | ( ~n26148 & n26150 ) ;
  assign n26152 = n21795 ^ n13969 ^ n7885 ;
  assign n26153 = ~n6421 & n21884 ;
  assign n26154 = n16063 ^ n231 ^ 1'b0 ;
  assign n26155 = n497 & ~n26154 ;
  assign n26156 = n8145 & ~n26155 ;
  assign n26157 = n12025 | n26156 ;
  assign n26158 = n26157 ^ n6649 ^ 1'b0 ;
  assign n26160 = n3733 & ~n4230 ;
  assign n26159 = ~n2461 & n7780 ;
  assign n26161 = n26160 ^ n26159 ^ 1'b0 ;
  assign n26162 = ~n16103 & n26161 ;
  assign n26163 = n19514 ^ n10569 ^ n6860 ;
  assign n26164 = n26163 ^ n22259 ^ 1'b0 ;
  assign n26165 = ( n5246 & n19343 ) | ( n5246 & ~n26164 ) | ( n19343 & ~n26164 ) ;
  assign n26168 = n6767 | n18107 ;
  assign n26169 = n836 | n26168 ;
  assign n26167 = ( n168 & n16662 ) | ( n168 & ~n21557 ) | ( n16662 & ~n21557 ) ;
  assign n26166 = ( ~n12586 & n15866 ) | ( ~n12586 & n19068 ) | ( n15866 & n19068 ) ;
  assign n26170 = n26169 ^ n26167 ^ n26166 ;
  assign n26171 = n26170 ^ n23711 ^ 1'b0 ;
  assign n26173 = n4722 | n9226 ;
  assign n26174 = n7308 & ~n26173 ;
  assign n26175 = n16983 | n26174 ;
  assign n26172 = n19394 ^ n8723 ^ n6827 ;
  assign n26176 = n26175 ^ n26172 ^ n5977 ;
  assign n26177 = n3407 ^ n2539 ^ 1'b0 ;
  assign n26178 = ~n8346 & n26177 ;
  assign n26179 = n26178 ^ n12204 ^ n4186 ;
  assign n26180 = n12632 ^ n10434 ^ n3851 ;
  assign n26181 = ~n20385 & n26180 ;
  assign n26182 = n26181 ^ n22664 ^ 1'b0 ;
  assign n26183 = n18260 ^ n6004 ^ n5050 ;
  assign n26184 = n26183 ^ n8762 ^ 1'b0 ;
  assign n26185 = n6667 & n26184 ;
  assign n26186 = n17069 ^ n3386 ^ 1'b0 ;
  assign n26187 = n21287 | n26186 ;
  assign n26188 = n22532 ^ n6749 ^ 1'b0 ;
  assign n26189 = n7403 & ~n26188 ;
  assign n26190 = ~n9360 & n26189 ;
  assign n26191 = n26190 ^ n20321 ^ 1'b0 ;
  assign n26192 = n18148 ^ n15223 ^ n13232 ;
  assign n26193 = n7814 & n16244 ;
  assign n26194 = n26193 ^ n22819 ^ n5788 ;
  assign n26195 = n13816 | n26194 ;
  assign n26196 = ( n9256 & n12339 ) | ( n9256 & ~n17958 ) | ( n12339 & ~n17958 ) ;
  assign n26197 = ( ~n7967 & n12543 ) | ( ~n7967 & n24020 ) | ( n12543 & n24020 ) ;
  assign n26198 = n5041 ^ n3145 ^ 1'b0 ;
  assign n26199 = n21398 & n25726 ;
  assign n26200 = n19512 ^ n10187 ^ n5187 ;
  assign n26201 = n21274 & ~n25541 ;
  assign n26202 = ( n1003 & n22870 ) | ( n1003 & ~n26201 ) | ( n22870 & ~n26201 ) ;
  assign n26203 = n12198 ^ n9379 ^ n6005 ;
  assign n26204 = n25187 ^ n16771 ^ 1'b0 ;
  assign n26205 = ~n26203 & n26204 ;
  assign n26206 = n13597 ^ n13328 ^ 1'b0 ;
  assign n26207 = n15955 & ~n26206 ;
  assign n26208 = n6856 & n24589 ;
  assign n26209 = ~n481 & n15001 ;
  assign n26210 = n13414 ^ n9873 ^ n1744 ;
  assign n26211 = n26209 & ~n26210 ;
  assign n26212 = ~n13568 & n26211 ;
  assign n26213 = ~n7119 & n26212 ;
  assign n26214 = n14046 ^ n7770 ^ n3484 ;
  assign n26215 = ( n4798 & n26213 ) | ( n4798 & ~n26214 ) | ( n26213 & ~n26214 ) ;
  assign n26216 = n25431 ^ n12379 ^ n9545 ;
  assign n26217 = n5003 ^ n294 ^ 1'b0 ;
  assign n26218 = n26217 ^ n6624 ^ n5195 ;
  assign n26219 = ~x110 & n6193 ;
  assign n26220 = n18014 | n26219 ;
  assign n26221 = ( ~n3078 & n3096 ) | ( ~n3078 & n26220 ) | ( n3096 & n26220 ) ;
  assign n26225 = n10005 & n10247 ;
  assign n26226 = n26225 ^ n9409 ^ 1'b0 ;
  assign n26227 = n6566 & n26226 ;
  assign n26224 = ( ~n4500 & n6064 ) | ( ~n4500 & n19593 ) | ( n6064 & n19593 ) ;
  assign n26222 = ( n934 & n8176 ) | ( n934 & n10377 ) | ( n8176 & n10377 ) ;
  assign n26223 = n26222 ^ n24637 ^ n6087 ;
  assign n26228 = n26227 ^ n26224 ^ n26223 ;
  assign n26229 = n11488 | n22806 ;
  assign n26230 = n26229 ^ n23329 ^ 1'b0 ;
  assign n26231 = ~n13242 & n26230 ;
  assign n26232 = n9017 & ~n26231 ;
  assign n26233 = ~n741 & n11941 ;
  assign n26234 = n25414 ^ n24845 ^ n24137 ;
  assign n26235 = n3006 & n15063 ;
  assign n26236 = ( n5196 & n12861 ) | ( n5196 & n26235 ) | ( n12861 & n26235 ) ;
  assign n26237 = n22602 ^ n3041 ^ 1'b0 ;
  assign n26238 = ( n11018 & n11910 ) | ( n11018 & ~n26237 ) | ( n11910 & ~n26237 ) ;
  assign n26239 = n21801 ^ n13240 ^ 1'b0 ;
  assign n26240 = n26239 ^ n24263 ^ n16585 ;
  assign n26241 = n13149 ^ n4034 ^ n2122 ;
  assign n26242 = n26241 ^ n13713 ^ 1'b0 ;
  assign n26243 = ( n2174 & n5722 ) | ( n2174 & n14077 ) | ( n5722 & n14077 ) ;
  assign n26244 = n15310 & ~n23835 ;
  assign n26245 = ~n26243 & n26244 ;
  assign n26246 = n14634 ^ n2418 ^ n831 ;
  assign n26247 = n8037 | n26246 ;
  assign n26248 = ~n4331 & n13530 ;
  assign n26249 = n26248 ^ n8692 ^ 1'b0 ;
  assign n26250 = ~n3104 & n9298 ;
  assign n26251 = n26250 ^ n22956 ^ 1'b0 ;
  assign n26252 = ( ~n2298 & n4913 ) | ( ~n2298 & n12044 ) | ( n4913 & n12044 ) ;
  assign n26253 = n25176 ^ n22382 ^ 1'b0 ;
  assign n26254 = n9808 & n23489 ;
  assign n26255 = n26254 ^ n13533 ^ 1'b0 ;
  assign n26256 = ( ~n3769 & n22091 ) | ( ~n3769 & n26255 ) | ( n22091 & n26255 ) ;
  assign n26257 = n22124 ^ n4173 ^ 1'b0 ;
  assign n26258 = ( x110 & ~n18300 ) | ( x110 & n26257 ) | ( ~n18300 & n26257 ) ;
  assign n26261 = n20555 ^ n3242 ^ n759 ;
  assign n26260 = n8145 & n18008 ;
  assign n26262 = n26261 ^ n26260 ^ 1'b0 ;
  assign n26263 = n26262 ^ n20354 ^ n3969 ;
  assign n26259 = n978 | n20227 ;
  assign n26264 = n26263 ^ n26259 ^ 1'b0 ;
  assign n26265 = n16938 ^ n16004 ^ 1'b0 ;
  assign n26266 = n12174 & ~n26265 ;
  assign n26267 = n8895 & ~n12538 ;
  assign n26268 = n26267 ^ n6310 ^ 1'b0 ;
  assign n26269 = n13777 ^ n1404 ^ 1'b0 ;
  assign n26270 = n22724 | n26269 ;
  assign n26271 = n26270 ^ n5029 ^ 1'b0 ;
  assign n26272 = ~n529 & n23838 ;
  assign n26273 = n19923 ^ n7627 ^ n1839 ;
  assign n26274 = n12898 ^ n4744 ^ n2488 ;
  assign n26275 = n26274 ^ n20217 ^ 1'b0 ;
  assign n26276 = n2670 | n20555 ;
  assign n26277 = n5066 | n26276 ;
  assign n26278 = n14796 & n20040 ;
  assign n26279 = n26278 ^ n6300 ^ 1'b0 ;
  assign n26280 = n14043 | n21341 ;
  assign n26281 = n2640 & ~n26280 ;
  assign n26282 = ( n3841 & n8745 ) | ( n3841 & ~n26281 ) | ( n8745 & ~n26281 ) ;
  assign n26283 = n9986 ^ n1702 ^ 1'b0 ;
  assign n26284 = n26283 ^ n26006 ^ 1'b0 ;
  assign n26285 = n4644 | n22249 ;
  assign n26286 = n3195 & n26285 ;
  assign n26287 = n8087 & n26286 ;
  assign n26288 = n16843 ^ n9544 ^ 1'b0 ;
  assign n26289 = ( n8008 & ~n12915 ) | ( n8008 & n26288 ) | ( ~n12915 & n26288 ) ;
  assign n26290 = ( n3122 & n5142 ) | ( n3122 & ~n26289 ) | ( n5142 & ~n26289 ) ;
  assign n26291 = n12857 ^ n12066 ^ 1'b0 ;
  assign n26292 = ( n3681 & ~n11447 ) | ( n3681 & n16198 ) | ( ~n11447 & n16198 ) ;
  assign n26293 = n26292 ^ n4607 ^ 1'b0 ;
  assign n26294 = n995 & n26293 ;
  assign n26295 = n15415 ^ n14309 ^ 1'b0 ;
  assign n26296 = ( x73 & ~n16743 ) | ( x73 & n23140 ) | ( ~n16743 & n23140 ) ;
  assign n26297 = n23244 ^ n6519 ^ n5191 ;
  assign n26298 = n7065 ^ n4647 ^ n1992 ;
  assign n26299 = n8644 & ~n8925 ;
  assign n26300 = n24885 ^ n3705 ^ 1'b0 ;
  assign n26301 = ~n11189 & n26300 ;
  assign n26302 = ( n5356 & n26299 ) | ( n5356 & ~n26301 ) | ( n26299 & ~n26301 ) ;
  assign n26304 = n5356 | n7038 ;
  assign n26303 = ~n2707 & n8958 ;
  assign n26305 = n26304 ^ n26303 ^ 1'b0 ;
  assign n26306 = ( ~n6598 & n19170 ) | ( ~n6598 & n21435 ) | ( n19170 & n21435 ) ;
  assign n26307 = n13939 & n15307 ;
  assign n26308 = ( ~n12838 & n21929 ) | ( ~n12838 & n26307 ) | ( n21929 & n26307 ) ;
  assign n26309 = n5342 | n7163 ;
  assign n26310 = n3614 & n12390 ;
  assign n26311 = ~n11528 & n26310 ;
  assign n26312 = ( ~n2284 & n26309 ) | ( ~n2284 & n26311 ) | ( n26309 & n26311 ) ;
  assign n26313 = n14251 ^ n7581 ^ n6784 ;
  assign n26314 = ( n2033 & n6179 ) | ( n2033 & ~n14644 ) | ( n6179 & ~n14644 ) ;
  assign n26315 = n26314 ^ n23542 ^ n21101 ;
  assign n26316 = n14101 ^ n13095 ^ 1'b0 ;
  assign n26317 = ( n5721 & ~n14504 ) | ( n5721 & n17009 ) | ( ~n14504 & n17009 ) ;
  assign n26318 = n26317 ^ n6166 ^ 1'b0 ;
  assign n26319 = n5155 & n26318 ;
  assign n26323 = n9792 ^ x123 ^ 1'b0 ;
  assign n26324 = n5064 | n26323 ;
  assign n26320 = n14449 | n15467 ;
  assign n26321 = n9798 & ~n26320 ;
  assign n26322 = n26321 ^ n21838 ^ n10632 ;
  assign n26325 = n26324 ^ n26322 ^ n14783 ;
  assign n26326 = n477 | n2246 ;
  assign n26327 = ( ~n186 & n22037 ) | ( ~n186 & n26326 ) | ( n22037 & n26326 ) ;
  assign n26328 = n25953 ^ n6883 ^ n4747 ;
  assign n26329 = n7484 & n21349 ;
  assign n26330 = ( n10924 & n23108 ) | ( n10924 & ~n26329 ) | ( n23108 & ~n26329 ) ;
  assign n26331 = n12559 & ~n24426 ;
  assign n26332 = n7235 & n26331 ;
  assign n26333 = n14629 ^ n8703 ^ n5150 ;
  assign n26334 = n26333 ^ n18389 ^ n5577 ;
  assign n26335 = ~n19438 & n26334 ;
  assign n26336 = n26335 ^ n2725 ^ 1'b0 ;
  assign n26337 = n15388 ^ n8855 ^ 1'b0 ;
  assign n26338 = n26337 ^ n18621 ^ n1739 ;
  assign n26339 = n10176 ^ n3198 ^ 1'b0 ;
  assign n26340 = n26339 ^ n20669 ^ n15170 ;
  assign n26341 = n6281 & ~n13536 ;
  assign n26342 = n26341 ^ n8096 ^ n4876 ;
  assign n26343 = n5277 | n18768 ;
  assign n26344 = n9361 & ~n26343 ;
  assign n26345 = n21761 ^ n11317 ^ n3903 ;
  assign n26346 = ( n18052 & n26344 ) | ( n18052 & ~n26345 ) | ( n26344 & ~n26345 ) ;
  assign n26351 = n24777 ^ n1794 ^ 1'b0 ;
  assign n26349 = n8010 | n16652 ;
  assign n26350 = n7085 | n26349 ;
  assign n26347 = ~n13757 & n22987 ;
  assign n26348 = n7237 & n26347 ;
  assign n26352 = n26351 ^ n26350 ^ n26348 ;
  assign n26353 = n5101 | n16777 ;
  assign n26354 = n26353 ^ n8093 ^ 1'b0 ;
  assign n26355 = n26354 ^ n22783 ^ n225 ;
  assign n26356 = n26355 ^ n1126 ^ 1'b0 ;
  assign n26357 = n3831 | n26356 ;
  assign n26358 = n6334 & ~n21999 ;
  assign n26366 = n835 & n1150 ;
  assign n26367 = n4948 & n26366 ;
  assign n26368 = ( n5261 & ~n9500 ) | ( n5261 & n26367 ) | ( ~n9500 & n26367 ) ;
  assign n26369 = ( n9756 & n12305 ) | ( n9756 & ~n26368 ) | ( n12305 & ~n26368 ) ;
  assign n26363 = ( n7189 & n8035 ) | ( n7189 & n11370 ) | ( n8035 & n11370 ) ;
  assign n26364 = n25935 ^ n23451 ^ 1'b0 ;
  assign n26365 = n26363 & n26364 ;
  assign n26370 = n26369 ^ n26365 ^ 1'b0 ;
  assign n26360 = n5489 ^ n3068 ^ n1762 ;
  assign n26359 = n1237 & ~n1439 ;
  assign n26361 = n26360 ^ n26359 ^ 1'b0 ;
  assign n26362 = ( n893 & n2260 ) | ( n893 & ~n26361 ) | ( n2260 & ~n26361 ) ;
  assign n26371 = n26370 ^ n26362 ^ 1'b0 ;
  assign n26372 = n14099 ^ n6149 ^ n4418 ;
  assign n26373 = ~n4275 & n5155 ;
  assign n26374 = n7433 & n26373 ;
  assign n26375 = n26374 ^ n19593 ^ n5976 ;
  assign n26376 = n2681 ^ n2222 ^ 1'b0 ;
  assign n26377 = ~n19478 & n26376 ;
  assign n26378 = ~n10890 & n15168 ;
  assign n26379 = n10679 | n19420 ;
  assign n26380 = n26379 ^ n19382 ^ n13486 ;
  assign n26381 = n17495 | n18540 ;
  assign n26382 = ( n865 & n5364 ) | ( n865 & n9342 ) | ( n5364 & n9342 ) ;
  assign n26383 = n26382 ^ n14809 ^ n637 ;
  assign n26384 = n24370 ^ n9481 ^ 1'b0 ;
  assign n26385 = n24561 ^ n11054 ^ 1'b0 ;
  assign n26386 = n6166 & ~n14918 ;
  assign n26387 = x68 & n26386 ;
  assign n26388 = ~n1899 & n7140 ;
  assign n26389 = n26388 ^ n23668 ^ 1'b0 ;
  assign n26390 = ~n26387 & n26389 ;
  assign n26391 = n13257 ^ n5910 ^ n1890 ;
  assign n26392 = n26391 ^ x42 ^ 1'b0 ;
  assign n26393 = n26390 & n26392 ;
  assign n26394 = n5594 & n25263 ;
  assign n26395 = n26394 ^ n9365 ^ 1'b0 ;
  assign n26396 = n26395 ^ n23212 ^ n21464 ;
  assign n26397 = n26396 ^ n5815 ^ 1'b0 ;
  assign n26398 = n12051 ^ n583 ^ 1'b0 ;
  assign n26399 = n26397 & ~n26398 ;
  assign n26400 = n9348 ^ n5098 ^ n1470 ;
  assign n26401 = n1362 & n1479 ;
  assign n26402 = n26400 & n26401 ;
  assign n26406 = n19906 ^ n11596 ^ 1'b0 ;
  assign n26403 = n5144 & ~n19844 ;
  assign n26404 = ~n6679 & n26403 ;
  assign n26405 = n1422 & n26404 ;
  assign n26407 = n26406 ^ n26405 ^ n1796 ;
  assign n26408 = n16066 ^ n15613 ^ 1'b0 ;
  assign n26409 = ~n18531 & n26408 ;
  assign n26410 = n1014 | n2677 ;
  assign n26411 = n26410 ^ n4640 ^ 1'b0 ;
  assign n26412 = n15843 | n26411 ;
  assign n26413 = n10203 | n26412 ;
  assign n26414 = ( n19676 & n19677 ) | ( n19676 & n26413 ) | ( n19677 & n26413 ) ;
  assign n26415 = ~n566 & n8945 ;
  assign n26416 = ~n816 & n26415 ;
  assign n26417 = n6317 & ~n18060 ;
  assign n26418 = n26416 & n26417 ;
  assign n26419 = ( n15688 & ~n21388 ) | ( n15688 & n26418 ) | ( ~n21388 & n26418 ) ;
  assign n26420 = n26419 ^ n14801 ^ n10261 ;
  assign n26421 = n16105 ^ n7591 ^ n3709 ;
  assign n26422 = ( n6077 & n22716 ) | ( n6077 & ~n26421 ) | ( n22716 & ~n26421 ) ;
  assign n26423 = n2537 | n13919 ;
  assign n26424 = n11877 & ~n26423 ;
  assign n26425 = n9060 & ~n21744 ;
  assign n26426 = n22953 | n26425 ;
  assign n26427 = n26426 ^ n1108 ^ 1'b0 ;
  assign n26428 = n16726 ^ n13201 ^ n7875 ;
  assign n26429 = ~n3809 & n26428 ;
  assign n26430 = n1563 & n5961 ;
  assign n26431 = ~n10904 & n26430 ;
  assign n26432 = n20905 ^ n9436 ^ 1'b0 ;
  assign n26433 = ( n5313 & ~n13300 ) | ( n5313 & n14339 ) | ( ~n13300 & n14339 ) ;
  assign n26434 = ( n13370 & n17001 ) | ( n13370 & ~n17035 ) | ( n17001 & ~n17035 ) ;
  assign n26435 = n3979 ^ n3522 ^ 1'b0 ;
  assign n26436 = ~n3709 & n26435 ;
  assign n26437 = ( n555 & ~n15532 ) | ( n555 & n26436 ) | ( ~n15532 & n26436 ) ;
  assign n26438 = n26437 ^ n25416 ^ n22078 ;
  assign n26440 = n8773 ^ n3035 ^ n744 ;
  assign n26439 = ( n329 & ~n2912 ) | ( n329 & n4748 ) | ( ~n2912 & n4748 ) ;
  assign n26441 = n26440 ^ n26439 ^ n1940 ;
  assign n26442 = n14323 | n17293 ;
  assign n26445 = n4290 & n11829 ;
  assign n26443 = n19619 ^ n17804 ^ n16659 ;
  assign n26444 = ~n15869 & n26443 ;
  assign n26446 = n26445 ^ n26444 ^ n10631 ;
  assign n26447 = ( n10904 & n11496 ) | ( n10904 & ~n20701 ) | ( n11496 & ~n20701 ) ;
  assign n26448 = ( n1952 & n5676 ) | ( n1952 & ~n26447 ) | ( n5676 & ~n26447 ) ;
  assign n26449 = n26448 ^ n16305 ^ n13407 ;
  assign n26450 = n10823 | n23323 ;
  assign n26451 = n7935 & ~n26450 ;
  assign n26452 = n6133 & n15661 ;
  assign n26453 = n18052 ^ n17591 ^ 1'b0 ;
  assign n26454 = ~n19124 & n26453 ;
  assign n26455 = ( n11078 & n26452 ) | ( n11078 & ~n26454 ) | ( n26452 & ~n26454 ) ;
  assign n26456 = ( n7658 & n26451 ) | ( n7658 & ~n26455 ) | ( n26451 & ~n26455 ) ;
  assign n26457 = n11641 | n13012 ;
  assign n26458 = n6194 & ~n26457 ;
  assign n26459 = n7498 & n26458 ;
  assign n26460 = n26459 ^ n13980 ^ n13170 ;
  assign n26462 = ( n4911 & n7840 ) | ( n4911 & n10493 ) | ( n7840 & n10493 ) ;
  assign n26461 = n21790 ^ n15137 ^ n3874 ;
  assign n26463 = n26462 ^ n26461 ^ n21179 ;
  assign n26464 = ( n1905 & n15281 ) | ( n1905 & ~n26463 ) | ( n15281 & ~n26463 ) ;
  assign n26465 = n23466 ^ n3028 ^ 1'b0 ;
  assign n26466 = ~n738 & n26465 ;
  assign n26467 = n5941 ^ n4273 ^ 1'b0 ;
  assign n26468 = ( n2670 & ~n15633 ) | ( n2670 & n26467 ) | ( ~n15633 & n26467 ) ;
  assign n26469 = n5200 ^ n3852 ^ 1'b0 ;
  assign n26470 = n26468 | n26469 ;
  assign n26471 = n2987 & ~n5161 ;
  assign n26472 = ( n5436 & n6343 ) | ( n5436 & ~n15434 ) | ( n6343 & ~n15434 ) ;
  assign n26473 = ~n10095 & n21025 ;
  assign n26474 = n26472 & n26473 ;
  assign n26475 = n22129 ^ n18225 ^ n8767 ;
  assign n26476 = n17146 ^ n7703 ^ n7095 ;
  assign n26477 = n6125 ^ n948 ^ 1'b0 ;
  assign n26478 = n816 & ~n26477 ;
  assign n26479 = n26478 ^ n25654 ^ n21936 ;
  assign n26480 = ( n4159 & n13797 ) | ( n4159 & ~n23032 ) | ( n13797 & ~n23032 ) ;
  assign n26481 = ~n849 & n1586 ;
  assign n26482 = n1239 & n26481 ;
  assign n26483 = ( ~n2760 & n3868 ) | ( ~n2760 & n26482 ) | ( n3868 & n26482 ) ;
  assign n26484 = ~n984 & n5348 ;
  assign n26485 = n26484 ^ n4769 ^ 1'b0 ;
  assign n26486 = ~n26483 & n26485 ;
  assign n26487 = ~n1674 & n11024 ;
  assign n26488 = n4583 & ~n15985 ;
  assign n26489 = n26488 ^ n2212 ^ 1'b0 ;
  assign n26490 = ( n7566 & ~n8002 ) | ( n7566 & n22962 ) | ( ~n8002 & n22962 ) ;
  assign n26491 = n24037 & n26490 ;
  assign n26492 = n26489 & n26491 ;
  assign n26493 = ( n2138 & n8849 ) | ( n2138 & n25221 ) | ( n8849 & n25221 ) ;
  assign n26494 = n26493 ^ n21457 ^ 1'b0 ;
  assign n26495 = ( ~n2427 & n12718 ) | ( ~n2427 & n15911 ) | ( n12718 & n15911 ) ;
  assign n26496 = ( n2632 & n4516 ) | ( n2632 & n22541 ) | ( n4516 & n22541 ) ;
  assign n26497 = n19618 ^ n16121 ^ n13261 ;
  assign n26498 = ( n26495 & n26496 ) | ( n26495 & n26497 ) | ( n26496 & n26497 ) ;
  assign n26499 = ( n11493 & n11741 ) | ( n11493 & n22345 ) | ( n11741 & n22345 ) ;
  assign n26500 = n21116 ^ n359 ^ 1'b0 ;
  assign n26501 = n25422 & n26500 ;
  assign n26502 = n5550 & ~n12568 ;
  assign n26503 = n26502 ^ n21436 ^ n1798 ;
  assign n26504 = n26309 ^ n18934 ^ n11488 ;
  assign n26505 = n24327 ^ n18698 ^ 1'b0 ;
  assign n26506 = ( ~n2237 & n4739 ) | ( ~n2237 & n6595 ) | ( n4739 & n6595 ) ;
  assign n26507 = ( n7871 & n20787 ) | ( n7871 & ~n26506 ) | ( n20787 & ~n26506 ) ;
  assign n26508 = ( n2293 & ~n19666 ) | ( n2293 & n26507 ) | ( ~n19666 & n26507 ) ;
  assign n26509 = n22331 ^ n3269 ^ 1'b0 ;
  assign n26510 = n6545 | n15038 ;
  assign n26511 = n16091 ^ n7371 ^ n6368 ;
  assign n26512 = n3386 & ~n26511 ;
  assign n26513 = ~n9072 & n26512 ;
  assign n26514 = n13297 & ~n16995 ;
  assign n26515 = n24090 | n26514 ;
  assign n26516 = n21210 | n26515 ;
  assign n26517 = n26511 ^ n20924 ^ n11403 ;
  assign n26518 = ( ~n275 & n483 ) | ( ~n275 & n20916 ) | ( n483 & n20916 ) ;
  assign n26519 = n10620 & ~n18540 ;
  assign n26520 = n3065 & n15659 ;
  assign n26521 = n26520 ^ n5150 ^ n1285 ;
  assign n26522 = n23858 ^ n10731 ^ n4635 ;
  assign n26523 = n9743 | n26522 ;
  assign n26524 = n24465 & n26523 ;
  assign n26525 = n5368 ^ n910 ^ 1'b0 ;
  assign n26526 = n23205 ^ n14116 ^ n7411 ;
  assign n26527 = n4282 | n20680 ;
  assign n26528 = n12236 ^ n5683 ^ 1'b0 ;
  assign n26529 = ~n8850 & n26528 ;
  assign n26530 = n26529 ^ n26126 ^ n10944 ;
  assign n26531 = n22601 ^ n10776 ^ 1'b0 ;
  assign n26532 = n26530 & n26531 ;
  assign n26533 = ~n22919 & n23931 ;
  assign n26535 = ~n2367 & n6177 ;
  assign n26536 = n26535 ^ n16683 ^ 1'b0 ;
  assign n26534 = n17835 ^ n9399 ^ n8127 ;
  assign n26537 = n26536 ^ n26534 ^ n19495 ;
  assign n26538 = n9404 & n9520 ;
  assign n26539 = ~n26537 & n26538 ;
  assign n26540 = n20500 ^ n15847 ^ 1'b0 ;
  assign n26541 = n6822 ^ n3825 ^ 1'b0 ;
  assign n26542 = n23581 | n26541 ;
  assign n26543 = n26542 ^ n3760 ^ 1'b0 ;
  assign n26544 = n26540 | n26543 ;
  assign n26549 = n11801 ^ n2057 ^ 1'b0 ;
  assign n26545 = ~n1879 & n3018 ;
  assign n26546 = n8219 & ~n26545 ;
  assign n26547 = n26546 ^ n10979 ^ n10513 ;
  assign n26548 = n6444 | n26547 ;
  assign n26550 = n26549 ^ n26548 ^ 1'b0 ;
  assign n26551 = ~n15247 & n26550 ;
  assign n26552 = ( n16076 & n26544 ) | ( n16076 & n26551 ) | ( n26544 & n26551 ) ;
  assign n26553 = n24129 ^ n14722 ^ n8429 ;
  assign n26554 = n18606 ^ n14735 ^ n12390 ;
  assign n26555 = n1504 | n15449 ;
  assign n26556 = n3724 & ~n26555 ;
  assign n26557 = n9315 & ~n26556 ;
  assign n26558 = n13012 & n26557 ;
  assign n26559 = ~n16383 & n26558 ;
  assign n26560 = ( x40 & n25491 ) | ( x40 & n26559 ) | ( n25491 & n26559 ) ;
  assign n26561 = n15227 ^ n14911 ^ 1'b0 ;
  assign n26562 = n22799 ^ n5281 ^ 1'b0 ;
  assign n26563 = n4556 | n26562 ;
  assign n26564 = ( n20458 & ~n21718 ) | ( n20458 & n21774 ) | ( ~n21718 & n21774 ) ;
  assign n26565 = n17050 ^ n9349 ^ 1'b0 ;
  assign n26566 = n26565 ^ n20004 ^ n7154 ;
  assign n26567 = n23379 ^ n15236 ^ n6337 ;
  assign n26568 = n26567 ^ n6914 ^ 1'b0 ;
  assign n26569 = ~n12562 & n26568 ;
  assign n26570 = ( n12353 & n25508 ) | ( n12353 & ~n26569 ) | ( n25508 & ~n26569 ) ;
  assign n26571 = n19029 ^ n6781 ^ n3370 ;
  assign n26572 = ( n19920 & ~n24661 ) | ( n19920 & n26571 ) | ( ~n24661 & n26571 ) ;
  assign n26573 = ~n2339 & n12093 ;
  assign n26574 = n26573 ^ n6368 ^ 1'b0 ;
  assign n26575 = n5027 & ~n9444 ;
  assign n26576 = n26575 ^ n23674 ^ 1'b0 ;
  assign n26577 = n18888 & ~n26576 ;
  assign n26578 = n1566 & ~n14680 ;
  assign n26579 = n26578 ^ n12557 ^ 1'b0 ;
  assign n26580 = n25808 ^ n19566 ^ 1'b0 ;
  assign n26581 = ( n15400 & ~n24667 ) | ( n15400 & n26580 ) | ( ~n24667 & n26580 ) ;
  assign n26582 = ( ~n11140 & n11534 ) | ( ~n11140 & n15228 ) | ( n11534 & n15228 ) ;
  assign n26583 = n6646 & n16717 ;
  assign n26586 = n13628 ^ n6783 ^ 1'b0 ;
  assign n26584 = n4077 & n16552 ;
  assign n26585 = n26584 ^ n12409 ^ 1'b0 ;
  assign n26587 = n26586 ^ n26585 ^ n9253 ;
  assign n26588 = ( n26582 & ~n26583 ) | ( n26582 & n26587 ) | ( ~n26583 & n26587 ) ;
  assign n26589 = ( n2243 & n6991 ) | ( n2243 & n17702 ) | ( n6991 & n17702 ) ;
  assign n26590 = n4868 & n5716 ;
  assign n26591 = ~n12739 & n26590 ;
  assign n26592 = n26591 ^ n23833 ^ n14634 ;
  assign n26593 = n2568 | n20520 ;
  assign n26594 = n17725 ^ n13394 ^ n8037 ;
  assign n26595 = n372 & ~n1972 ;
  assign n26596 = n23033 ^ n12977 ^ n8393 ;
  assign n26597 = n13954 ^ n1411 ^ 1'b0 ;
  assign n26598 = ( n4795 & n11391 ) | ( n4795 & ~n17521 ) | ( n11391 & ~n17521 ) ;
  assign n26599 = n20159 ^ n18684 ^ 1'b0 ;
  assign n26600 = n8201 & n9826 ;
  assign n26601 = ~n9826 & n26600 ;
  assign n26602 = n15299 | n26601 ;
  assign n26603 = n26601 & ~n26602 ;
  assign n26604 = ( n1412 & n2545 ) | ( n1412 & ~n26603 ) | ( n2545 & ~n26603 ) ;
  assign n26605 = ( n11080 & n19765 ) | ( n11080 & ~n21388 ) | ( n19765 & ~n21388 ) ;
  assign n26607 = ~n2724 & n4076 ;
  assign n26608 = n24336 | n26607 ;
  assign n26606 = n3902 & ~n16192 ;
  assign n26609 = n26608 ^ n26606 ^ 1'b0 ;
  assign n26610 = n9876 ^ n7684 ^ n758 ;
  assign n26611 = n12661 & n26610 ;
  assign n26612 = n5037 | n11501 ;
  assign n26613 = n11414 & ~n26612 ;
  assign n26614 = n16350 ^ n3755 ^ 1'b0 ;
  assign n26615 = n7906 ^ n866 ^ 1'b0 ;
  assign n26616 = n26614 & ~n26615 ;
  assign n26617 = n4052 | n23289 ;
  assign n26618 = n26617 ^ n17185 ^ 1'b0 ;
  assign n26619 = ~n1105 & n14294 ;
  assign n26620 = n11597 ^ n11441 ^ n2252 ;
  assign n26621 = n21082 & n26620 ;
  assign n26622 = ( n21983 & n22309 ) | ( n21983 & n26621 ) | ( n22309 & n26621 ) ;
  assign n26623 = ( x109 & n3707 ) | ( x109 & ~n15191 ) | ( n3707 & ~n15191 ) ;
  assign n26624 = n26623 ^ n21260 ^ n1323 ;
  assign n26625 = ( n5590 & ~n10018 ) | ( n5590 & n10645 ) | ( ~n10018 & n10645 ) ;
  assign n26626 = ( n2032 & n26439 ) | ( n2032 & ~n26625 ) | ( n26439 & ~n26625 ) ;
  assign n26627 = n22998 ^ n21906 ^ n9114 ;
  assign n26628 = n20877 ^ n13371 ^ n12157 ;
  assign n26629 = ( n2296 & ~n7882 ) | ( n2296 & n19720 ) | ( ~n7882 & n19720 ) ;
  assign n26630 = n13580 & ~n26629 ;
  assign n26631 = n16280 & n26630 ;
  assign n26632 = n1362 & n4394 ;
  assign n26633 = n26632 ^ n10779 ^ 1'b0 ;
  assign n26634 = n12710 ^ n10518 ^ 1'b0 ;
  assign n26635 = ~n21067 & n26634 ;
  assign n26636 = n5730 & n18716 ;
  assign n26637 = n1800 & n26636 ;
  assign n26638 = n26637 ^ n13306 ^ n13120 ;
  assign n26639 = n16614 ^ n16013 ^ n9236 ;
  assign n26640 = ( n17784 & n19476 ) | ( n17784 & n20374 ) | ( n19476 & n20374 ) ;
  assign n26641 = ( n322 & ~n5661 ) | ( n322 & n26640 ) | ( ~n5661 & n26640 ) ;
  assign n26642 = n24271 & ~n26482 ;
  assign n26644 = n15665 ^ n7427 ^ n4627 ;
  assign n26643 = n6637 | n19283 ;
  assign n26645 = n26644 ^ n26643 ^ 1'b0 ;
  assign n26648 = n13292 & ~n17275 ;
  assign n26646 = n14752 & n25187 ;
  assign n26647 = n12276 | n26646 ;
  assign n26649 = n26648 ^ n26647 ^ 1'b0 ;
  assign n26650 = n4375 ^ n4191 ^ n3096 ;
  assign n26651 = n26650 ^ n18163 ^ n2560 ;
  assign n26652 = ( n8681 & ~n16126 ) | ( n8681 & n26651 ) | ( ~n16126 & n26651 ) ;
  assign n26653 = n11849 | n13577 ;
  assign n26654 = n12426 & ~n16054 ;
  assign n26655 = ( ~n2417 & n3953 ) | ( ~n2417 & n7726 ) | ( n3953 & n7726 ) ;
  assign n26656 = ( ~n986 & n11866 ) | ( ~n986 & n26655 ) | ( n11866 & n26655 ) ;
  assign n26657 = ( n5592 & n6330 ) | ( n5592 & ~n13050 ) | ( n6330 & ~n13050 ) ;
  assign n26658 = ( n17892 & ~n26656 ) | ( n17892 & n26657 ) | ( ~n26656 & n26657 ) ;
  assign n26659 = n12259 ^ n2181 ^ 1'b0 ;
  assign n26660 = n3781 & n26659 ;
  assign n26661 = n26660 ^ n788 ^ 1'b0 ;
  assign n26662 = ~n803 & n26661 ;
  assign n26663 = n896 | n12269 ;
  assign n26664 = n26663 ^ n10493 ^ 1'b0 ;
  assign n26665 = ( ~n2791 & n8619 ) | ( ~n2791 & n15932 ) | ( n8619 & n15932 ) ;
  assign n26666 = ~n10228 & n26665 ;
  assign n26667 = ~n11841 & n26666 ;
  assign n26668 = n10000 & ~n16739 ;
  assign n26669 = n26668 ^ n22177 ^ 1'b0 ;
  assign n26670 = n6361 | n26669 ;
  assign n26671 = n433 | n22044 ;
  assign n26672 = n26671 ^ n2478 ^ 1'b0 ;
  assign n26673 = n23140 ^ x64 ^ 1'b0 ;
  assign n26674 = n17416 & n26673 ;
  assign n26675 = ( n13454 & ~n24305 ) | ( n13454 & n26674 ) | ( ~n24305 & n26674 ) ;
  assign n26676 = ( n3144 & ~n6083 ) | ( n3144 & n9750 ) | ( ~n6083 & n9750 ) ;
  assign n26677 = x108 & n4558 ;
  assign n26678 = ( ~n5206 & n6699 ) | ( ~n5206 & n26677 ) | ( n6699 & n26677 ) ;
  assign n26679 = ( n15439 & n26676 ) | ( n15439 & ~n26678 ) | ( n26676 & ~n26678 ) ;
  assign n26680 = ~n11618 & n14733 ;
  assign n26681 = ~x99 & n1872 ;
  assign n26682 = ~n236 & n10570 ;
  assign n26683 = n26681 & n26682 ;
  assign n26684 = ( ~n21298 & n26549 ) | ( ~n21298 & n26683 ) | ( n26549 & n26683 ) ;
  assign n26685 = ( n2629 & ~n20987 ) | ( n2629 & n26684 ) | ( ~n20987 & n26684 ) ;
  assign n26686 = ( n5423 & n9713 ) | ( n5423 & n12359 ) | ( n9713 & n12359 ) ;
  assign n26687 = n13204 ^ n5340 ^ n2880 ;
  assign n26688 = n26687 ^ n12902 ^ n5479 ;
  assign n26689 = ( n4883 & ~n26686 ) | ( n4883 & n26688 ) | ( ~n26686 & n26688 ) ;
  assign n26690 = n25580 ^ n4717 ^ 1'b0 ;
  assign n26691 = n4855 & ~n26690 ;
  assign n26692 = n12781 & ~n14572 ;
  assign n26693 = n26692 ^ n18975 ^ 1'b0 ;
  assign n26694 = x44 & n19987 ;
  assign n26695 = ( n5191 & n18761 ) | ( n5191 & n26694 ) | ( n18761 & n26694 ) ;
  assign n26696 = n20802 ^ n3653 ^ n719 ;
  assign n26697 = n24336 ^ n17488 ^ n9253 ;
  assign n26698 = n4055 ^ n1397 ^ 1'b0 ;
  assign n26699 = ~n10497 & n26698 ;
  assign n26700 = ( n5921 & n10792 ) | ( n5921 & n26699 ) | ( n10792 & n26699 ) ;
  assign n26701 = ( ~n20841 & n26697 ) | ( ~n20841 & n26700 ) | ( n26697 & n26700 ) ;
  assign n26702 = ( n8300 & n17141 ) | ( n8300 & ~n22792 ) | ( n17141 & ~n22792 ) ;
  assign n26703 = n26702 ^ n21466 ^ n1618 ;
  assign n26704 = n26703 ^ n9256 ^ 1'b0 ;
  assign n26705 = n10223 & ~n11104 ;
  assign n26706 = n18771 ^ n3123 ^ 1'b0 ;
  assign n26707 = ( n19850 & n26705 ) | ( n19850 & ~n26706 ) | ( n26705 & ~n26706 ) ;
  assign n26708 = n21891 ^ n9332 ^ n2410 ;
  assign n26709 = n14746 ^ n5582 ^ n1752 ;
  assign n26710 = n26709 ^ n7733 ^ 1'b0 ;
  assign n26711 = n18815 | n26710 ;
  assign n26712 = n12836 ^ n10104 ^ n2537 ;
  assign n26713 = n6989 ^ n3120 ^ 1'b0 ;
  assign n26714 = n26712 | n26713 ;
  assign n26715 = n7722 & ~n10695 ;
  assign n26716 = ( x50 & ~n4457 ) | ( x50 & n5516 ) | ( ~n4457 & n5516 ) ;
  assign n26719 = n22765 ^ n21975 ^ 1'b0 ;
  assign n26718 = n17157 & ~n26167 ;
  assign n26720 = n26719 ^ n26718 ^ 1'b0 ;
  assign n26721 = n15982 & n26720 ;
  assign n26722 = n26721 ^ n1369 ^ 1'b0 ;
  assign n26717 = ( ~n5076 & n18852 ) | ( ~n5076 & n24244 ) | ( n18852 & n24244 ) ;
  assign n26723 = n26722 ^ n26717 ^ n1660 ;
  assign n26724 = n9172 ^ n2905 ^ 1'b0 ;
  assign n26725 = n12537 ^ n170 ^ 1'b0 ;
  assign n26726 = n13177 ^ n9895 ^ n9383 ;
  assign n26727 = n11394 ^ n9199 ^ 1'b0 ;
  assign n26728 = n10499 | n26727 ;
  assign n26729 = n26728 ^ n4867 ^ 1'b0 ;
  assign n26730 = n26726 | n26729 ;
  assign n26731 = n25137 ^ n7144 ^ 1'b0 ;
  assign n26732 = ~n26730 & n26731 ;
  assign n26733 = ( n1668 & n17440 ) | ( n1668 & ~n19676 ) | ( n17440 & ~n19676 ) ;
  assign n26734 = n18876 ^ n4748 ^ 1'b0 ;
  assign n26735 = n3961 ^ n2882 ^ 1'b0 ;
  assign n26736 = ( ~n2159 & n13797 ) | ( ~n2159 & n26735 ) | ( n13797 & n26735 ) ;
  assign n26738 = n4711 ^ n1323 ^ 1'b0 ;
  assign n26739 = n4583 & n26738 ;
  assign n26737 = ( ~n5273 & n7843 ) | ( ~n5273 & n17617 ) | ( n7843 & n17617 ) ;
  assign n26740 = n26739 ^ n26737 ^ n14050 ;
  assign n26741 = n5054 & n16418 ;
  assign n26742 = ~n26740 & n26741 ;
  assign n26743 = n26736 & ~n26742 ;
  assign n26744 = n2384 ^ n1474 ^ x85 ;
  assign n26745 = n7349 ^ n6728 ^ n1489 ;
  assign n26746 = n2273 & ~n2578 ;
  assign n26747 = n26746 ^ n16179 ^ 1'b0 ;
  assign n26748 = ~n3971 & n26747 ;
  assign n26749 = ~n26745 & n26748 ;
  assign n26750 = ( ~n12260 & n16375 ) | ( ~n12260 & n26749 ) | ( n16375 & n26749 ) ;
  assign n26751 = n3598 & n22657 ;
  assign n26752 = n26751 ^ n26210 ^ 1'b0 ;
  assign n26753 = n6773 ^ n2968 ^ 1'b0 ;
  assign n26754 = n10977 | n26753 ;
  assign n26755 = n22616 & ~n26754 ;
  assign n26763 = n3184 & ~n7635 ;
  assign n26764 = ~n18747 & n26763 ;
  assign n26760 = n25331 ^ n10855 ^ n1097 ;
  assign n26761 = n26760 ^ n12940 ^ 1'b0 ;
  assign n26762 = ~n15579 & n26761 ;
  assign n26765 = n26764 ^ n26762 ^ n2112 ;
  assign n26756 = n18902 & ~n21290 ;
  assign n26757 = n26416 & n26756 ;
  assign n26758 = n3389 ^ n656 ^ 1'b0 ;
  assign n26759 = ~n26757 & n26758 ;
  assign n26766 = n26765 ^ n26759 ^ 1'b0 ;
  assign n26767 = n12739 & n26766 ;
  assign n26768 = ( n2008 & ~n6218 ) | ( n2008 & n12543 ) | ( ~n6218 & n12543 ) ;
  assign n26769 = n14568 ^ n11017 ^ n2682 ;
  assign n26770 = ( n7588 & n8370 ) | ( n7588 & ~n11563 ) | ( n8370 & ~n11563 ) ;
  assign n26771 = ( n11507 & n26769 ) | ( n11507 & ~n26770 ) | ( n26769 & ~n26770 ) ;
  assign n26772 = n9747 & ~n25162 ;
  assign n26773 = n14335 ^ n2136 ^ 1'b0 ;
  assign n26774 = n21078 & ~n26773 ;
  assign n26775 = n26774 ^ n16931 ^ n16652 ;
  assign n26776 = n26775 ^ n10960 ^ 1'b0 ;
  assign n26777 = n20601 ^ n17343 ^ n4406 ;
  assign n26778 = n15379 ^ n7433 ^ 1'b0 ;
  assign n26779 = n4503 & n26778 ;
  assign n26780 = ( ~n4332 & n26777 ) | ( ~n4332 & n26779 ) | ( n26777 & n26779 ) ;
  assign n26781 = n18048 ^ n11090 ^ 1'b0 ;
  assign n26782 = ~n1226 & n16576 ;
  assign n26783 = ~n11332 & n26782 ;
  assign n26784 = n2215 & ~n16643 ;
  assign n26785 = n26784 ^ n8559 ^ 1'b0 ;
  assign n26786 = n7907 ^ n5934 ^ 1'b0 ;
  assign n26787 = ( n141 & ~n7929 ) | ( n141 & n26786 ) | ( ~n7929 & n26786 ) ;
  assign n26788 = n9549 & n14604 ;
  assign n26789 = n14276 & n26788 ;
  assign n26790 = ~n867 & n24675 ;
  assign n26791 = n26789 & n26790 ;
  assign n26792 = n6576 & ~n26791 ;
  assign n26793 = ~n26787 & n26792 ;
  assign n26794 = n18527 ^ n7596 ^ n7331 ;
  assign n26795 = ~n21891 & n26794 ;
  assign n26796 = n14721 & n26795 ;
  assign n26797 = n26796 ^ n21929 ^ 1'b0 ;
  assign n26798 = n489 & n26797 ;
  assign n26799 = n3098 & n3743 ;
  assign n26800 = n26799 ^ n23922 ^ 1'b0 ;
  assign n26801 = n6331 & ~n7688 ;
  assign n26802 = n26801 ^ n9171 ^ 1'b0 ;
  assign n26803 = n2900 ^ n2842 ^ 1'b0 ;
  assign n26804 = ( ~n11493 & n17546 ) | ( ~n11493 & n26803 ) | ( n17546 & n26803 ) ;
  assign n26805 = n26802 & n26804 ;
  assign n26806 = n6004 & n26805 ;
  assign n26807 = ( n1649 & ~n2293 ) | ( n1649 & n26806 ) | ( ~n2293 & n26806 ) ;
  assign n26808 = n6050 & n7032 ;
  assign n26809 = n26808 ^ n16055 ^ n8239 ;
  assign n26810 = n7562 ^ n7268 ^ n1858 ;
  assign n26811 = n5233 & n16387 ;
  assign n26812 = n26811 ^ n14061 ^ 1'b0 ;
  assign n26813 = n8988 & ~n26812 ;
  assign n26814 = n26813 ^ n2592 ^ 1'b0 ;
  assign n26815 = ( n8283 & n26810 ) | ( n8283 & ~n26814 ) | ( n26810 & ~n26814 ) ;
  assign n26816 = n21436 ^ n570 ^ 1'b0 ;
  assign n26817 = n18579 | n26816 ;
  assign n26818 = n26817 ^ n24917 ^ n13575 ;
  assign n26820 = n5704 ^ n3533 ^ 1'b0 ;
  assign n26821 = n26820 ^ n25147 ^ n10432 ;
  assign n26819 = ~n9666 & n16865 ;
  assign n26822 = n26821 ^ n26819 ^ 1'b0 ;
  assign n26823 = n13318 ^ n7327 ^ 1'b0 ;
  assign n26824 = n22117 | n26823 ;
  assign n26825 = n22594 ^ n17078 ^ n9852 ;
  assign n26827 = ( ~n2325 & n4418 ) | ( ~n2325 & n6974 ) | ( n4418 & n6974 ) ;
  assign n26828 = n26827 ^ n18335 ^ 1'b0 ;
  assign n26829 = n18002 | n26828 ;
  assign n26826 = ~n1485 & n5650 ;
  assign n26830 = n26829 ^ n26826 ^ 1'b0 ;
  assign n26831 = ( n3592 & n26317 ) | ( n3592 & ~n26830 ) | ( n26317 & ~n26830 ) ;
  assign n26836 = ~n15723 & n19124 ;
  assign n26837 = n26836 ^ n16115 ^ n6443 ;
  assign n26832 = n4028 ^ n3944 ^ n1150 ;
  assign n26833 = n6478 & n26832 ;
  assign n26834 = n26833 ^ n6175 ^ 1'b0 ;
  assign n26835 = n26834 ^ n9920 ^ 1'b0 ;
  assign n26838 = n26837 ^ n26835 ^ n5246 ;
  assign n26839 = n6861 & ~n20722 ;
  assign n26840 = n13519 ^ n4331 ^ 1'b0 ;
  assign n26841 = n26839 & ~n26840 ;
  assign n26842 = ~n12663 & n15300 ;
  assign n26843 = n9865 | n20523 ;
  assign n26844 = ( n5052 & n24934 ) | ( n5052 & n26843 ) | ( n24934 & n26843 ) ;
  assign n26845 = ( n18909 & ~n19836 ) | ( n18909 & n26075 ) | ( ~n19836 & n26075 ) ;
  assign n26846 = ( ~n6471 & n16241 ) | ( ~n6471 & n16840 ) | ( n16241 & n16840 ) ;
  assign n26847 = ~n7794 & n26846 ;
  assign n26848 = n17593 ^ n11013 ^ n9387 ;
  assign n26849 = n2373 & n16342 ;
  assign n26850 = n4429 & n26849 ;
  assign n26851 = n1001 & n14500 ;
  assign n26852 = ~n9875 & n26851 ;
  assign n26853 = ( ~n20459 & n26850 ) | ( ~n20459 & n26852 ) | ( n26850 & n26852 ) ;
  assign n26854 = n3798 ^ n896 ^ 1'b0 ;
  assign n26855 = n9170 | n26854 ;
  assign n26856 = n10685 & ~n26855 ;
  assign n26857 = n26856 ^ n11662 ^ 1'b0 ;
  assign n26858 = n15562 ^ n12992 ^ 1'b0 ;
  assign n26859 = ~n1992 & n26858 ;
  assign n26860 = ~n19882 & n23048 ;
  assign n26861 = n4844 | n19716 ;
  assign n26862 = n26861 ^ n18940 ^ 1'b0 ;
  assign n26863 = n12149 ^ n11810 ^ 1'b0 ;
  assign n26864 = n26862 | n26863 ;
  assign n26867 = n22249 ^ n4740 ^ 1'b0 ;
  assign n26868 = n8294 & n26867 ;
  assign n26865 = n3996 & ~n25100 ;
  assign n26866 = n17805 & n26865 ;
  assign n26869 = n26868 ^ n26866 ^ n6519 ;
  assign n26870 = ( n15080 & ~n16181 ) | ( n15080 & n25884 ) | ( ~n16181 & n25884 ) ;
  assign n26873 = n9722 ^ n4961 ^ n1127 ;
  assign n26871 = n11702 | n15796 ;
  assign n26872 = n26871 ^ n8463 ^ 1'b0 ;
  assign n26874 = n26873 ^ n26872 ^ n3050 ;
  assign n26875 = n19618 ^ n2691 ^ 1'b0 ;
  assign n26876 = ~n2103 & n26875 ;
  assign n26877 = ( n1208 & ~n3589 ) | ( n1208 & n19995 ) | ( ~n3589 & n19995 ) ;
  assign n26878 = n26877 ^ n5181 ^ 1'b0 ;
  assign n26879 = n26876 & n26878 ;
  assign n26880 = ~n3167 & n26879 ;
  assign n26881 = ~n5155 & n26880 ;
  assign n26882 = n8751 & n26881 ;
  assign n26883 = n7530 & ~n12735 ;
  assign n26884 = ~n26882 & n26883 ;
  assign n26885 = n4217 & n6731 ;
  assign n26886 = n26885 ^ n1657 ^ 1'b0 ;
  assign n26887 = ~n1829 & n26886 ;
  assign n26888 = ~n13011 & n26887 ;
  assign n26889 = n13330 ^ n9948 ^ 1'b0 ;
  assign n26890 = ( n11086 & n14679 ) | ( n11086 & ~n16867 ) | ( n14679 & ~n16867 ) ;
  assign n26891 = n17022 ^ n8189 ^ n4679 ;
  assign n26892 = n26891 ^ n22782 ^ 1'b0 ;
  assign n26893 = ~n1508 & n5068 ;
  assign n26894 = n18180 & n26893 ;
  assign n26895 = n20380 & n26894 ;
  assign n26896 = n11124 ^ n5868 ^ 1'b0 ;
  assign n26897 = n23868 | n26896 ;
  assign n26898 = n13177 & ~n26897 ;
  assign n26899 = ~n14944 & n17050 ;
  assign n26900 = ~n26898 & n26899 ;
  assign n26901 = n13737 & n18551 ;
  assign n26902 = n9935 & n26901 ;
  assign n26903 = n26902 ^ n7448 ^ 1'b0 ;
  assign n26904 = n7771 & ~n16160 ;
  assign n26905 = n2659 | n11714 ;
  assign n26906 = n26904 | n26905 ;
  assign n26907 = n519 & n26906 ;
  assign n26908 = n533 | n19625 ;
  assign n26909 = n26908 ^ n26107 ^ 1'b0 ;
  assign n26910 = n19500 ^ n17729 ^ n16163 ;
  assign n26911 = n26910 ^ n24292 ^ n10782 ;
  assign n26912 = n5471 & ~n26911 ;
  assign n26913 = n8014 ^ n3537 ^ 1'b0 ;
  assign n26914 = n26913 ^ n25848 ^ n20669 ;
  assign n26915 = n3947 | n12986 ;
  assign n26916 = n14601 ^ n3058 ^ 1'b0 ;
  assign n26917 = ~n2928 & n26916 ;
  assign n26918 = n26917 ^ n10012 ^ n7775 ;
  assign n26919 = n26918 ^ n14328 ^ n5431 ;
  assign n26920 = n26919 ^ n11319 ^ n5477 ;
  assign n26921 = n19043 ^ n14316 ^ n7307 ;
  assign n26922 = ( n4800 & ~n12426 ) | ( n4800 & n26921 ) | ( ~n12426 & n26921 ) ;
  assign n26923 = n12367 & n13601 ;
  assign n26924 = n23927 & n26923 ;
  assign n26925 = n2860 & ~n11497 ;
  assign n26926 = ( ~n6334 & n6533 ) | ( ~n6334 & n22354 ) | ( n6533 & n22354 ) ;
  assign n26927 = n26926 ^ n5154 ^ 1'b0 ;
  assign n26928 = ~n26925 & n26927 ;
  assign n26929 = ( n14951 & ~n16614 ) | ( n14951 & n19350 ) | ( ~n16614 & n19350 ) ;
  assign n26930 = n9171 | n17174 ;
  assign n26933 = n16238 ^ n1974 ^ n662 ;
  assign n26934 = ( n8094 & n11857 ) | ( n8094 & ~n26933 ) | ( n11857 & ~n26933 ) ;
  assign n26931 = n23581 ^ n18104 ^ n8912 ;
  assign n26932 = ( n2121 & n7518 ) | ( n2121 & ~n26931 ) | ( n7518 & ~n26931 ) ;
  assign n26935 = n26934 ^ n26932 ^ n11670 ;
  assign n26936 = n3013 ^ n2784 ^ 1'b0 ;
  assign n26937 = n14563 & ~n26936 ;
  assign n26938 = ( ~n8738 & n12897 ) | ( ~n8738 & n26937 ) | ( n12897 & n26937 ) ;
  assign n26939 = n14029 ^ n9342 ^ 1'b0 ;
  assign n26940 = n316 | n26939 ;
  assign n26941 = n24760 & ~n26940 ;
  assign n26942 = ( ~x122 & n10525 ) | ( ~x122 & n13292 ) | ( n10525 & n13292 ) ;
  assign n26944 = ~n1800 & n2564 ;
  assign n26945 = n26944 ^ n26918 ^ n2706 ;
  assign n26943 = n5595 ^ n3851 ^ 1'b0 ;
  assign n26946 = n26945 ^ n26943 ^ n8771 ;
  assign n26947 = n21492 ^ n21116 ^ n129 ;
  assign n26948 = n26947 ^ n24570 ^ n5805 ;
  assign n26949 = ( n6799 & ~n8670 ) | ( n6799 & n11323 ) | ( ~n8670 & n11323 ) ;
  assign n26950 = n9399 & n26949 ;
  assign n26951 = n26950 ^ n20710 ^ n19035 ;
  assign n26957 = ( n3221 & n14221 ) | ( n3221 & ~n22129 ) | ( n14221 & ~n22129 ) ;
  assign n26952 = n26416 ^ n13763 ^ n10122 ;
  assign n26953 = ( ~n4209 & n6659 ) | ( ~n4209 & n9630 ) | ( n6659 & n9630 ) ;
  assign n26954 = n5071 | n26953 ;
  assign n26955 = n26954 ^ n3144 ^ 1'b0 ;
  assign n26956 = ( n8548 & n26952 ) | ( n8548 & ~n26955 ) | ( n26952 & ~n26955 ) ;
  assign n26958 = n26957 ^ n26956 ^ n12202 ;
  assign n26962 = n14650 ^ n6039 ^ n5408 ;
  assign n26959 = ~n3021 & n5847 ;
  assign n26960 = n26959 ^ n1871 ^ 1'b0 ;
  assign n26961 = n26960 ^ n25093 ^ 1'b0 ;
  assign n26963 = n26962 ^ n26961 ^ n12218 ;
  assign n26964 = n26963 ^ n7766 ^ n960 ;
  assign n26965 = n4462 ^ x53 ^ 1'b0 ;
  assign n26966 = ~n577 & n9367 ;
  assign n26967 = n26966 ^ n14667 ^ 1'b0 ;
  assign n26968 = ~n6427 & n8754 ;
  assign n26969 = n26968 ^ n24935 ^ n14846 ;
  assign n26970 = ( ~n4808 & n8723 ) | ( ~n4808 & n26969 ) | ( n8723 & n26969 ) ;
  assign n26971 = n10546 ^ n3182 ^ n867 ;
  assign n26972 = n26971 ^ n11819 ^ n3695 ;
  assign n26973 = ( ~n23606 & n24949 ) | ( ~n23606 & n26490 ) | ( n24949 & n26490 ) ;
  assign n26974 = n5301 ^ n3771 ^ 1'b0 ;
  assign n26975 = n1349 & ~n26974 ;
  assign n26976 = n26975 ^ n14650 ^ n10253 ;
  assign n26977 = ( ~n6347 & n11746 ) | ( ~n6347 & n16330 ) | ( n11746 & n16330 ) ;
  assign n26980 = n12293 ^ n4900 ^ n3785 ;
  assign n26978 = n10403 & ~n13341 ;
  assign n26979 = ~n11116 & n26978 ;
  assign n26981 = n26980 ^ n26979 ^ n20551 ;
  assign n26982 = n21207 & ~n26981 ;
  assign n26983 = ~n26977 & n26982 ;
  assign n26984 = ( n929 & n9819 ) | ( n929 & ~n26983 ) | ( n9819 & ~n26983 ) ;
  assign n26986 = n15901 ^ n3937 ^ n1355 ;
  assign n26985 = n1246 & ~n17100 ;
  assign n26987 = n26986 ^ n26985 ^ 1'b0 ;
  assign n26988 = ( n12563 & n13767 ) | ( n12563 & n14736 ) | ( n13767 & n14736 ) ;
  assign n26989 = ( n717 & ~n26987 ) | ( n717 & n26988 ) | ( ~n26987 & n26988 ) ;
  assign n26990 = n26989 ^ n23362 ^ n1592 ;
  assign n26991 = n19295 ^ n3550 ^ n631 ;
  assign n26992 = n365 & n26991 ;
  assign n26993 = ~n2894 & n26992 ;
  assign n26994 = n25761 ^ n6864 ^ 1'b0 ;
  assign n26995 = ~n26993 & n26994 ;
  assign n26996 = n5195 & ~n5499 ;
  assign n26997 = n26996 ^ n22130 ^ 1'b0 ;
  assign n26998 = n5816 ^ n434 ^ 1'b0 ;
  assign n26999 = ( ~n244 & n3794 ) | ( ~n244 & n26998 ) | ( n3794 & n26998 ) ;
  assign n27000 = n26999 ^ n201 ^ 1'b0 ;
  assign n27001 = n7228 | n27000 ;
  assign n27002 = n5622 & n24761 ;
  assign n27003 = n866 | n19546 ;
  assign n27004 = ~n8329 & n24750 ;
  assign n27005 = ~n13640 & n27004 ;
  assign n27006 = ( ~n13894 & n27003 ) | ( ~n13894 & n27005 ) | ( n27003 & n27005 ) ;
  assign n27007 = n24862 ^ n5809 ^ n3914 ;
  assign n27008 = ( ~n1797 & n7226 ) | ( ~n1797 & n23179 ) | ( n7226 & n23179 ) ;
  assign n27009 = n15933 ^ n8311 ^ 1'b0 ;
  assign n27010 = ( n6255 & n27008 ) | ( n6255 & n27009 ) | ( n27008 & n27009 ) ;
  assign n27011 = n2176 & ~n6138 ;
  assign n27012 = ~n11379 & n27011 ;
  assign n27013 = n365 & n27012 ;
  assign n27014 = n13108 & ~n27013 ;
  assign n27015 = n27014 ^ n4578 ^ n3392 ;
  assign n27016 = n9584 ^ n1984 ^ n660 ;
  assign n27017 = ( n11298 & n13482 ) | ( n11298 & ~n27016 ) | ( n13482 & ~n27016 ) ;
  assign n27018 = n20797 ^ n1821 ^ 1'b0 ;
  assign n27019 = n22975 & n27018 ;
  assign n27020 = ( n1090 & n5536 ) | ( n1090 & ~n27019 ) | ( n5536 & ~n27019 ) ;
  assign n27021 = ( n20811 & n27017 ) | ( n20811 & n27020 ) | ( n27017 & n27020 ) ;
  assign n27022 = ( n4528 & ~n16524 ) | ( n4528 & n20103 ) | ( ~n16524 & n20103 ) ;
  assign n27023 = n27022 ^ n9092 ^ 1'b0 ;
  assign n27024 = ( ~n7994 & n11657 ) | ( ~n7994 & n27023 ) | ( n11657 & n27023 ) ;
  assign n27025 = n27024 ^ n15122 ^ n9086 ;
  assign n27026 = ~n2640 & n4657 ;
  assign n27027 = n27026 ^ n4498 ^ 1'b0 ;
  assign n27028 = n11004 ^ n7680 ^ 1'b0 ;
  assign n27029 = n6153 | n27028 ;
  assign n27030 = ~n19551 & n27029 ;
  assign n27031 = n9625 & n22422 ;
  assign n27032 = n21712 & n27031 ;
  assign n27033 = n27032 ^ n12337 ^ 1'b0 ;
  assign n27034 = n7511 & ~n27033 ;
  assign n27035 = n5998 | n8184 ;
  assign n27036 = n27035 ^ n12722 ^ n7163 ;
  assign n27037 = n27036 ^ n1626 ^ 1'b0 ;
  assign n27038 = n11778 ^ n6271 ^ 1'b0 ;
  assign n27039 = ( n3768 & ~n10020 ) | ( n3768 & n20795 ) | ( ~n10020 & n20795 ) ;
  assign n27040 = n27039 ^ n10252 ^ 1'b0 ;
  assign n27041 = ( n7722 & n21071 ) | ( n7722 & ~n27040 ) | ( n21071 & ~n27040 ) ;
  assign n27042 = ( n2913 & n8748 ) | ( n2913 & n23442 ) | ( n8748 & n23442 ) ;
  assign n27043 = n25379 ^ n14220 ^ n3578 ;
  assign n27044 = ~n9449 & n27043 ;
  assign n27045 = n18995 ^ n16280 ^ n8037 ;
  assign n27046 = n3976 ^ n1427 ^ 1'b0 ;
  assign n27047 = n2472 & ~n27046 ;
  assign n27048 = n27047 ^ n11919 ^ 1'b0 ;
  assign n27049 = n1299 & ~n27048 ;
  assign n27050 = n2725 & ~n2893 ;
  assign n27051 = n27050 ^ n6839 ^ 1'b0 ;
  assign n27052 = n716 | n27051 ;
  assign n27053 = n6482 | n27052 ;
  assign n27054 = n885 & n17372 ;
  assign n27055 = n27054 ^ n20021 ^ 1'b0 ;
  assign n27056 = n13327 ^ n8519 ^ 1'b0 ;
  assign n27057 = n25466 ^ n6550 ^ 1'b0 ;
  assign n27060 = n8714 ^ n5025 ^ n307 ;
  assign n27058 = n3742 & ~n12408 ;
  assign n27059 = ( ~n4578 & n8631 ) | ( ~n4578 & n27058 ) | ( n8631 & n27058 ) ;
  assign n27061 = n27060 ^ n27059 ^ n9986 ;
  assign n27062 = ( n2935 & ~n12778 ) | ( n2935 & n18452 ) | ( ~n12778 & n18452 ) ;
  assign n27063 = n27062 ^ n1688 ^ 1'b0 ;
  assign n27064 = n4455 | n17727 ;
  assign n27065 = ( n6019 & n15867 ) | ( n6019 & n22467 ) | ( n15867 & n22467 ) ;
  assign n27066 = n27065 ^ n912 ^ 1'b0 ;
  assign n27067 = n27064 | n27066 ;
  assign n27070 = n1362 & n3631 ;
  assign n27068 = ( n18404 & n19177 ) | ( n18404 & n20500 ) | ( n19177 & n20500 ) ;
  assign n27069 = n7460 & n27068 ;
  assign n27071 = n27070 ^ n27069 ^ 1'b0 ;
  assign n27072 = n24039 ^ n20268 ^ 1'b0 ;
  assign n27073 = n2478 | n13173 ;
  assign n27074 = n27073 ^ n9828 ^ 1'b0 ;
  assign n27076 = n11569 ^ n8807 ^ n6187 ;
  assign n27075 = ~n9683 & n17439 ;
  assign n27077 = n27076 ^ n27075 ^ 1'b0 ;
  assign n27078 = ~n4793 & n5250 ;
  assign n27079 = n1070 & n27078 ;
  assign n27080 = ~n1023 & n27079 ;
  assign n27081 = ( ~n2994 & n7769 ) | ( ~n2994 & n11086 ) | ( n7769 & n11086 ) ;
  assign n27082 = n10618 & n27081 ;
  assign n27083 = n27080 | n27082 ;
  assign n27084 = ~n17124 & n26100 ;
  assign n27085 = ( n4667 & n10503 ) | ( n4667 & ~n27084 ) | ( n10503 & ~n27084 ) ;
  assign n27086 = n2153 | n17840 ;
  assign n27087 = n27086 ^ n9745 ^ x3 ;
  assign n27088 = n27087 ^ n18902 ^ n14661 ;
  assign n27089 = ( n6028 & n17537 ) | ( n6028 & ~n27088 ) | ( n17537 & ~n27088 ) ;
  assign n27090 = n24769 ^ n19043 ^ n2363 ;
  assign n27091 = ( n5627 & ~n8576 ) | ( n5627 & n12644 ) | ( ~n8576 & n12644 ) ;
  assign n27092 = ( n5154 & n6918 ) | ( n5154 & n27091 ) | ( n6918 & n27091 ) ;
  assign n27093 = n27092 ^ n26686 ^ n22060 ;
  assign n27094 = ~n14244 & n27093 ;
  assign n27095 = n2435 & ~n11353 ;
  assign n27096 = n3749 & n27095 ;
  assign n27097 = n6072 ^ n3448 ^ 1'b0 ;
  assign n27098 = n27096 | n27097 ;
  assign n27100 = n5510 ^ n621 ^ 1'b0 ;
  assign n27101 = n7095 & ~n27100 ;
  assign n27099 = n3375 | n5616 ;
  assign n27102 = n27101 ^ n27099 ^ 1'b0 ;
  assign n27103 = n1001 | n17547 ;
  assign n27104 = n27103 ^ n26262 ^ 1'b0 ;
  assign n27106 = ( n2420 & n2911 ) | ( n2420 & n3055 ) | ( n2911 & n3055 ) ;
  assign n27105 = n18763 ^ n18367 ^ n4084 ;
  assign n27107 = n27106 ^ n27105 ^ n26812 ;
  assign n27108 = n23922 ^ n18927 ^ n8725 ;
  assign n27109 = x34 & n935 ;
  assign n27110 = ~n935 & n27109 ;
  assign n27111 = n27110 ^ n7055 ^ 1'b0 ;
  assign n27112 = n27111 ^ n6026 ^ n4697 ;
  assign n27113 = n27112 ^ n21824 ^ n646 ;
  assign n27114 = n522 & ~n5867 ;
  assign n27115 = n5909 & n27114 ;
  assign n27116 = n13444 | n27115 ;
  assign n27117 = n22592 | n27116 ;
  assign n27118 = n8877 ^ n4902 ^ n3787 ;
  assign n27119 = ( ~n25889 & n27117 ) | ( ~n25889 & n27118 ) | ( n27117 & n27118 ) ;
  assign n27120 = n23148 ^ n11820 ^ 1'b0 ;
  assign n27121 = n7714 ^ n6433 ^ 1'b0 ;
  assign n27122 = n27121 ^ n20597 ^ n17958 ;
  assign n27123 = n27122 ^ n20575 ^ 1'b0 ;
  assign n27124 = n17735 ^ n1496 ^ 1'b0 ;
  assign n27125 = n2614 ^ n1732 ^ 1'b0 ;
  assign n27126 = n27124 | n27125 ;
  assign n27127 = n18162 ^ n14412 ^ 1'b0 ;
  assign n27128 = n2912 & ~n27127 ;
  assign n27129 = n27128 ^ n14866 ^ 1'b0 ;
  assign n27130 = n23920 & n27129 ;
  assign n27131 = n235 & n27130 ;
  assign n27132 = n20384 ^ n10029 ^ 1'b0 ;
  assign n27133 = n4759 | n9980 ;
  assign n27134 = ~n27132 & n27133 ;
  assign n27135 = n27134 ^ n13327 ^ n8959 ;
  assign n27136 = n13462 | n23545 ;
  assign n27137 = n27135 | n27136 ;
  assign n27138 = n27137 ^ n18707 ^ n10876 ;
  assign n27139 = ( n5403 & ~n17472 ) | ( n5403 & n26615 ) | ( ~n17472 & n26615 ) ;
  assign n27140 = n21238 ^ n15307 ^ 1'b0 ;
  assign n27141 = ~n27139 & n27140 ;
  assign n27142 = ( ~n197 & n4196 ) | ( ~n197 & n14640 ) | ( n4196 & n14640 ) ;
  assign n27143 = ( ~n26932 & n27141 ) | ( ~n26932 & n27142 ) | ( n27141 & n27142 ) ;
  assign n27144 = n6970 ^ n6262 ^ 1'b0 ;
  assign n27145 = n3074 & ~n27144 ;
  assign n27146 = n27145 ^ n12964 ^ 1'b0 ;
  assign n27147 = n7553 & n24738 ;
  assign n27148 = ( n1006 & ~n3544 ) | ( n1006 & n3871 ) | ( ~n3544 & n3871 ) ;
  assign n27149 = n27148 ^ n20902 ^ n14879 ;
  assign n27150 = ~n7982 & n27149 ;
  assign n27151 = n5126 & ~n13955 ;
  assign n27152 = n27151 ^ n17947 ^ 1'b0 ;
  assign n27153 = n13516 | n23107 ;
  assign n27154 = n16687 ^ n15762 ^ n15384 ;
  assign n27155 = n27154 ^ n17982 ^ 1'b0 ;
  assign n27156 = n1795 & n27155 ;
  assign n27157 = n4874 & ~n8065 ;
  assign n27158 = ( n9405 & ~n9528 ) | ( n9405 & n16712 ) | ( ~n9528 & n16712 ) ;
  assign n27159 = n3414 | n21305 ;
  assign n27160 = n25934 & ~n27159 ;
  assign n27161 = ( ~n11094 & n24475 ) | ( ~n11094 & n27160 ) | ( n24475 & n27160 ) ;
  assign n27162 = n6773 & ~n16488 ;
  assign n27163 = n27162 ^ n20988 ^ n6485 ;
  assign n27164 = n7898 ^ n2532 ^ 1'b0 ;
  assign n27165 = n5609 | n27164 ;
  assign n27166 = n27165 ^ n8577 ^ n6098 ;
  assign n27167 = ~n311 & n13774 ;
  assign n27168 = n27167 ^ n18771 ^ 1'b0 ;
  assign n27170 = n1152 & ~n17022 ;
  assign n27171 = ( ~n11629 & n21035 ) | ( ~n11629 & n27170 ) | ( n21035 & n27170 ) ;
  assign n27169 = n4981 | n5548 ;
  assign n27172 = n27171 ^ n27169 ^ n13225 ;
  assign n27178 = n7899 | n17431 ;
  assign n27179 = n27178 ^ n713 ^ 1'b0 ;
  assign n27176 = n3292 & ~n9845 ;
  assign n27177 = n27176 ^ n12323 ^ 1'b0 ;
  assign n27174 = ( n2657 & n4608 ) | ( n2657 & n6967 ) | ( n4608 & n6967 ) ;
  assign n27173 = ( n5518 & n12045 ) | ( n5518 & n20358 ) | ( n12045 & n20358 ) ;
  assign n27175 = n27174 ^ n27173 ^ n6424 ;
  assign n27180 = n27179 ^ n27177 ^ n27175 ;
  assign n27181 = n27180 ^ n16145 ^ 1'b0 ;
  assign n27182 = n27172 & ~n27181 ;
  assign n27183 = n1551 & ~n4788 ;
  assign n27184 = ~n22865 & n27183 ;
  assign n27185 = n4372 & n9658 ;
  assign n27186 = n7126 | n27185 ;
  assign n27187 = n14634 | n27186 ;
  assign n27188 = n5300 & ~n9187 ;
  assign n27189 = ( n5712 & n6980 ) | ( n5712 & ~n8171 ) | ( n6980 & ~n8171 ) ;
  assign n27190 = n27189 ^ n7793 ^ 1'b0 ;
  assign n27191 = ~n18398 & n19125 ;
  assign n27192 = n27190 & n27191 ;
  assign n27193 = ( n5164 & ~n7712 ) | ( n5164 & n10487 ) | ( ~n7712 & n10487 ) ;
  assign n27194 = n2313 & ~n12671 ;
  assign n27195 = n27194 ^ n9743 ^ 1'b0 ;
  assign n27196 = ( n16495 & n27193 ) | ( n16495 & n27195 ) | ( n27193 & n27195 ) ;
  assign n27197 = ( ~n14017 & n14407 ) | ( ~n14017 & n20096 ) | ( n14407 & n20096 ) ;
  assign n27198 = n27197 ^ n26961 ^ n6500 ;
  assign n27199 = n11172 & ~n12027 ;
  assign n27200 = n19277 | n27199 ;
  assign n27201 = ( ~n7895 & n8783 ) | ( ~n7895 & n9538 ) | ( n8783 & n9538 ) ;
  assign n27202 = n12763 ^ n937 ^ 1'b0 ;
  assign n27203 = n3996 & ~n4112 ;
  assign n27204 = n27203 ^ n6230 ^ 1'b0 ;
  assign n27205 = n27204 ^ n637 ^ 1'b0 ;
  assign n27206 = n27205 ^ n14639 ^ 1'b0 ;
  assign n27207 = n20335 ^ n9912 ^ 1'b0 ;
  assign n27208 = n27206 & n27207 ;
  assign n27209 = ~n2921 & n11579 ;
  assign n27210 = n2843 & n27209 ;
  assign n27211 = n3769 | n12946 ;
  assign n27212 = n27210 & ~n27211 ;
  assign n27213 = n19161 ^ n4933 ^ n3560 ;
  assign n27214 = n27213 ^ n2360 ^ 1'b0 ;
  assign n27215 = n9187 ^ n1553 ^ 1'b0 ;
  assign n27216 = ( n768 & ~n6862 ) | ( n768 & n11215 ) | ( ~n6862 & n11215 ) ;
  assign n27220 = n9087 ^ n1486 ^ 1'b0 ;
  assign n27221 = n8330 & ~n27220 ;
  assign n27217 = ~n6125 & n10904 ;
  assign n27218 = ~n8111 & n27217 ;
  assign n27219 = n27218 ^ n14225 ^ 1'b0 ;
  assign n27222 = n27221 ^ n27219 ^ n15951 ;
  assign n27223 = ( n12129 & n15326 ) | ( n12129 & ~n17591 ) | ( n15326 & ~n17591 ) ;
  assign n27224 = ~n7296 & n11151 ;
  assign n27225 = ~n2179 & n5924 ;
  assign n27226 = ~n27224 & n27225 ;
  assign n27227 = n8446 ^ n5424 ^ 1'b0 ;
  assign n27228 = n980 | n3173 ;
  assign n27229 = n27227 & ~n27228 ;
  assign n27230 = n22066 ^ n7452 ^ 1'b0 ;
  assign n27231 = n27229 | n27230 ;
  assign n27232 = n3899 & n4774 ;
  assign n27233 = ~n2950 & n27232 ;
  assign n27234 = n2446 & ~n27233 ;
  assign n27235 = ( n5736 & n6524 ) | ( n5736 & ~n16238 ) | ( n6524 & ~n16238 ) ;
  assign n27236 = n3641 ^ n2736 ^ 1'b0 ;
  assign n27237 = ~n27235 & n27236 ;
  assign n27238 = n7021 & ~n8633 ;
  assign n27239 = n5837 & n27238 ;
  assign n27240 = n6505 & ~n27239 ;
  assign n27241 = n27240 ^ n9262 ^ 1'b0 ;
  assign n27242 = ( n7032 & n21434 ) | ( n7032 & ~n27241 ) | ( n21434 & ~n27241 ) ;
  assign n27243 = n1124 & ~n16239 ;
  assign n27244 = n27243 ^ n8126 ^ 1'b0 ;
  assign n27245 = ( n1811 & n2970 ) | ( n1811 & ~n27244 ) | ( n2970 & ~n27244 ) ;
  assign n27246 = ~n6060 & n7687 ;
  assign n27247 = n2103 & n11799 ;
  assign n27248 = n26897 & n27247 ;
  assign n27249 = ( ~n5345 & n27246 ) | ( ~n5345 & n27248 ) | ( n27246 & n27248 ) ;
  assign n27250 = ( n395 & n1411 ) | ( n395 & ~n11523 ) | ( n1411 & ~n11523 ) ;
  assign n27251 = ( n4026 & n14679 ) | ( n4026 & ~n27250 ) | ( n14679 & ~n27250 ) ;
  assign n27252 = ( n9628 & n14414 ) | ( n9628 & n22518 ) | ( n14414 & n22518 ) ;
  assign n27253 = ( n12239 & n16147 ) | ( n12239 & n18039 ) | ( n16147 & n18039 ) ;
  assign n27254 = ( n436 & ~n6029 ) | ( n436 & n10499 ) | ( ~n6029 & n10499 ) ;
  assign n27255 = n11340 ^ n5212 ^ 1'b0 ;
  assign n27256 = n27255 ^ n17836 ^ n16712 ;
  assign n27257 = ~n9050 & n27256 ;
  assign n27258 = n27254 & n27257 ;
  assign n27259 = n20474 ^ n8796 ^ 1'b0 ;
  assign n27260 = n1554 & ~n27259 ;
  assign n27261 = ~n5634 & n20795 ;
  assign n27262 = n27261 ^ n10058 ^ 1'b0 ;
  assign n27263 = n25745 ^ n8580 ^ 1'b0 ;
  assign n27264 = n17391 & n27263 ;
  assign n27265 = n20526 ^ n10624 ^ 1'b0 ;
  assign n27266 = n17075 ^ n342 ^ 1'b0 ;
  assign n27267 = ~n6963 & n27266 ;
  assign n27268 = ( ~n10729 & n15360 ) | ( ~n10729 & n25961 ) | ( n15360 & n25961 ) ;
  assign n27269 = n1171 & ~n4179 ;
  assign n27270 = n8149 & n27269 ;
  assign n27271 = ~n5698 & n27270 ;
  assign n27272 = ( n1528 & n15272 ) | ( n1528 & n27271 ) | ( n15272 & n27271 ) ;
  assign n27273 = n24692 ^ n10577 ^ n7649 ;
  assign n27274 = n15300 ^ n2093 ^ 1'b0 ;
  assign n27275 = n7940 & n27274 ;
  assign n27276 = n2256 & ~n10259 ;
  assign n27277 = n26567 ^ n18912 ^ n6929 ;
  assign n27278 = n12788 ^ n2862 ^ n2834 ;
  assign n27279 = n23757 ^ n7785 ^ 1'b0 ;
  assign n27280 = ( n8633 & n13339 ) | ( n8633 & ~n16220 ) | ( n13339 & ~n16220 ) ;
  assign n27281 = ( n8144 & n27279 ) | ( n8144 & ~n27280 ) | ( n27279 & ~n27280 ) ;
  assign n27282 = n24924 ^ n16924 ^ n676 ;
  assign n27283 = n12326 ^ n4018 ^ n778 ;
  assign n27284 = n13292 & n17138 ;
  assign n27285 = n20900 & n27284 ;
  assign n27286 = ( n14777 & ~n27283 ) | ( n14777 & n27285 ) | ( ~n27283 & n27285 ) ;
  assign n27287 = n5413 & ~n14375 ;
  assign n27288 = n27287 ^ n9273 ^ 1'b0 ;
  assign n27289 = ( n2270 & n3102 ) | ( n2270 & n15477 ) | ( n3102 & n15477 ) ;
  assign n27290 = n27289 ^ n194 ^ 1'b0 ;
  assign n27291 = n13162 | n27290 ;
  assign n27292 = n6984 ^ n5203 ^ n778 ;
  assign n27293 = n11224 ^ n6084 ^ n599 ;
  assign n27294 = n27293 ^ n10715 ^ 1'b0 ;
  assign n27295 = ~n17326 & n18752 ;
  assign n27296 = n12335 | n22641 ;
  assign n27297 = n16808 & ~n27296 ;
  assign n27298 = ( n12626 & n15035 ) | ( n12626 & ~n15039 ) | ( n15035 & ~n15039 ) ;
  assign n27299 = ( ~n2153 & n10489 ) | ( ~n2153 & n27298 ) | ( n10489 & n27298 ) ;
  assign n27300 = n27299 ^ n3390 ^ 1'b0 ;
  assign n27301 = n2257 | n27300 ;
  assign n27302 = n27301 ^ n18089 ^ 1'b0 ;
  assign n27303 = n757 | n2770 ;
  assign n27304 = n27303 ^ n5981 ^ 1'b0 ;
  assign n27305 = n27304 ^ n8144 ^ 1'b0 ;
  assign n27306 = n10303 | n27305 ;
  assign n27307 = n12659 | n27306 ;
  assign n27308 = ~n553 & n20145 ;
  assign n27309 = ~n3918 & n27308 ;
  assign n27310 = n27309 ^ n14735 ^ n9980 ;
  assign n27311 = n16092 ^ n478 ^ 1'b0 ;
  assign n27312 = ( ~n11246 & n16677 ) | ( ~n11246 & n27311 ) | ( n16677 & n27311 ) ;
  assign n27313 = n27312 ^ n19235 ^ n1865 ;
  assign n27314 = n27313 ^ n9797 ^ n5807 ;
  assign n27315 = n3837 ^ n3255 ^ n561 ;
  assign n27316 = n27315 ^ n7582 ^ n1958 ;
  assign n27317 = n1872 & ~n25844 ;
  assign n27318 = ( n12618 & n27316 ) | ( n12618 & n27317 ) | ( n27316 & n27317 ) ;
  assign n27319 = n16999 ^ n13182 ^ n1055 ;
  assign n27320 = ( n4121 & n10961 ) | ( n4121 & n15707 ) | ( n10961 & n15707 ) ;
  assign n27321 = n7100 & ~n15928 ;
  assign n27322 = n20210 & n27321 ;
  assign n27323 = n9050 ^ n4462 ^ n1690 ;
  assign n27324 = ~n27229 & n27323 ;
  assign n27325 = n27322 & ~n27324 ;
  assign n27326 = ( n8615 & ~n27320 ) | ( n8615 & n27325 ) | ( ~n27320 & n27325 ) ;
  assign n27327 = n6334 & n9975 ;
  assign n27328 = ~n24926 & n27327 ;
  assign n27329 = ( n2913 & ~n6897 ) | ( n2913 & n27328 ) | ( ~n6897 & n27328 ) ;
  assign n27330 = ~n24043 & n27329 ;
  assign n27331 = n20982 ^ n3043 ^ 1'b0 ;
  assign n27332 = n10196 & n27331 ;
  assign n27333 = n25430 ^ n20611 ^ n174 ;
  assign n27334 = n1076 | n3337 ;
  assign n27335 = n27334 ^ n14374 ^ 1'b0 ;
  assign n27336 = n27335 ^ n15150 ^ n5045 ;
  assign n27337 = ( n7202 & ~n9830 ) | ( n7202 & n17654 ) | ( ~n9830 & n17654 ) ;
  assign n27338 = n27337 ^ n11177 ^ n10936 ;
  assign n27339 = n20507 ^ n16971 ^ n11916 ;
  assign n27340 = ( x40 & n1179 ) | ( x40 & ~n4810 ) | ( n1179 & ~n4810 ) ;
  assign n27343 = n10742 & n14700 ;
  assign n27344 = n27343 ^ n11949 ^ 1'b0 ;
  assign n27341 = ( n5804 & n10263 ) | ( n5804 & n12299 ) | ( n10263 & n12299 ) ;
  assign n27342 = n18538 & ~n27341 ;
  assign n27345 = n27344 ^ n27342 ^ 1'b0 ;
  assign n27346 = ~n7981 & n23710 ;
  assign n27347 = n27346 ^ n4867 ^ 1'b0 ;
  assign n27351 = ( n4101 & n17570 ) | ( n4101 & ~n24025 ) | ( n17570 & ~n24025 ) ;
  assign n27348 = n3026 ^ n2367 ^ 1'b0 ;
  assign n27349 = ( n5507 & n11101 ) | ( n5507 & ~n27348 ) | ( n11101 & ~n27348 ) ;
  assign n27350 = n2992 & n27349 ;
  assign n27352 = n27351 ^ n27350 ^ 1'b0 ;
  assign n27353 = n12819 & ~n14483 ;
  assign n27354 = ~n3614 & n27353 ;
  assign n27355 = n12679 | n16248 ;
  assign n27356 = ( n21636 & ~n27354 ) | ( n21636 & n27355 ) | ( ~n27354 & n27355 ) ;
  assign n27357 = ( n2622 & n6312 ) | ( n2622 & n6347 ) | ( n6312 & n6347 ) ;
  assign n27358 = ( ~n624 & n4354 ) | ( ~n624 & n15173 ) | ( n4354 & n15173 ) ;
  assign n27359 = ( n6406 & n8791 ) | ( n6406 & ~n9342 ) | ( n8791 & ~n9342 ) ;
  assign n27360 = n27359 ^ n19798 ^ 1'b0 ;
  assign n27361 = n9539 ^ n3850 ^ n796 ;
  assign n27362 = ~n22214 & n27361 ;
  assign n27363 = n7418 | n20848 ;
  assign n27364 = n27363 ^ n4660 ^ 1'b0 ;
  assign n27365 = n15066 ^ n3161 ^ 1'b0 ;
  assign n27366 = n896 & ~n27365 ;
  assign n27367 = ~n13719 & n27366 ;
  assign n27368 = ~n26101 & n27367 ;
  assign n27369 = n25569 ^ n22588 ^ n3807 ;
  assign n27370 = n27369 ^ n14979 ^ n7479 ;
  assign n27371 = n14413 ^ n9346 ^ n4250 ;
  assign n27372 = n2839 | n5854 ;
  assign n27373 = n8540 & ~n27372 ;
  assign n27374 = n19683 & ~n27373 ;
  assign n27375 = n24151 | n27082 ;
  assign n27376 = n10690 ^ n8755 ^ 1'b0 ;
  assign n27378 = ( ~n3291 & n3666 ) | ( ~n3291 & n11504 ) | ( n3666 & n11504 ) ;
  assign n27377 = n26056 ^ n19394 ^ 1'b0 ;
  assign n27379 = n27378 ^ n27377 ^ n15257 ;
  assign n27380 = n2786 & ~n14567 ;
  assign n27381 = n27380 ^ n12738 ^ n6659 ;
  assign n27382 = ( n710 & ~n8713 ) | ( n710 & n15236 ) | ( ~n8713 & n15236 ) ;
  assign n27383 = n5062 ^ n2377 ^ 1'b0 ;
  assign n27384 = n14130 ^ n7935 ^ n447 ;
  assign n27385 = n4812 & n27384 ;
  assign n27387 = ~n7421 & n16971 ;
  assign n27388 = ( n6136 & n23406 ) | ( n6136 & ~n27387 ) | ( n23406 & ~n27387 ) ;
  assign n27386 = ~n16278 & n25759 ;
  assign n27389 = n27388 ^ n27386 ^ 1'b0 ;
  assign n27390 = n11803 ^ n732 ^ 1'b0 ;
  assign n27391 = n253 & ~n11726 ;
  assign n27392 = n2374 ^ n1574 ^ n1452 ;
  assign n27393 = n27392 ^ n6760 ^ 1'b0 ;
  assign n27394 = n13708 | n15859 ;
  assign n27395 = n27394 ^ n4098 ^ 1'b0 ;
  assign n27396 = ~n7444 & n27395 ;
  assign n27397 = ( ~n8232 & n12991 ) | ( ~n8232 & n25600 ) | ( n12991 & n25600 ) ;
  assign n27401 = ( n4991 & n10115 ) | ( n4991 & n14682 ) | ( n10115 & n14682 ) ;
  assign n27398 = ( ~n13919 & n14839 ) | ( ~n13919 & n20296 ) | ( n14839 & n20296 ) ;
  assign n27399 = n27398 ^ n1426 ^ 1'b0 ;
  assign n27400 = n7774 | n27399 ;
  assign n27402 = n27401 ^ n27400 ^ n18621 ;
  assign n27403 = n27402 ^ n9759 ^ n4534 ;
  assign n27404 = n3998 ^ n3301 ^ 1'b0 ;
  assign n27405 = n23040 & ~n27404 ;
  assign n27406 = ( n632 & ~n4580 ) | ( n632 & n13594 ) | ( ~n4580 & n13594 ) ;
  assign n27407 = n2393 | n16718 ;
  assign n27408 = n6354 | n27407 ;
  assign n27409 = ( n15185 & n24561 ) | ( n15185 & n27408 ) | ( n24561 & n27408 ) ;
  assign n27410 = ( n792 & ~n2402 ) | ( n792 & n11073 ) | ( ~n2402 & n11073 ) ;
  assign n27411 = n4647 & ~n8980 ;
  assign n27412 = n5353 & n27411 ;
  assign n27413 = ( ~n26917 & n27410 ) | ( ~n26917 & n27412 ) | ( n27410 & n27412 ) ;
  assign n27414 = n5681 & ~n12464 ;
  assign n27415 = ~n24636 & n27414 ;
  assign n27416 = n27415 ^ n11650 ^ 1'b0 ;
  assign n27417 = ( n8709 & ~n16838 ) | ( n8709 & n19811 ) | ( ~n16838 & n19811 ) ;
  assign n27418 = n23495 ^ n12811 ^ 1'b0 ;
  assign n27419 = ~n14404 & n22337 ;
  assign n27420 = n27419 ^ n14391 ^ 1'b0 ;
  assign n27421 = n8395 ^ n8096 ^ 1'b0 ;
  assign n27422 = n4578 ^ n2264 ^ n692 ;
  assign n27423 = n3048 & n7030 ;
  assign n27424 = n27423 ^ n6566 ^ 1'b0 ;
  assign n27425 = n6435 ^ n2813 ^ 1'b0 ;
  assign n27426 = n8261 & n27425 ;
  assign n27427 = n10649 ^ n3157 ^ n275 ;
  assign n27428 = n27427 ^ n14597 ^ 1'b0 ;
  assign n27429 = n27426 & ~n27428 ;
  assign n27430 = ( ~n27422 & n27424 ) | ( ~n27422 & n27429 ) | ( n27424 & n27429 ) ;
  assign n27434 = n12601 ^ n10403 ^ 1'b0 ;
  assign n27433 = n20153 ^ n5774 ^ 1'b0 ;
  assign n27431 = ( n6844 & n13201 ) | ( n6844 & n20121 ) | ( n13201 & n20121 ) ;
  assign n27432 = n27431 ^ n20506 ^ n377 ;
  assign n27435 = n27434 ^ n27433 ^ n27432 ;
  assign n27437 = n505 | n3885 ;
  assign n27438 = n15690 | n27437 ;
  assign n27436 = n6646 ^ n2113 ^ n471 ;
  assign n27439 = n27438 ^ n27436 ^ n15338 ;
  assign n27440 = n27439 ^ n1577 ^ 1'b0 ;
  assign n27441 = n4614 & ~n27315 ;
  assign n27442 = n27441 ^ n17365 ^ n15986 ;
  assign n27443 = n27442 ^ n8977 ^ n4236 ;
  assign n27444 = ( ~n8243 & n19394 ) | ( ~n8243 & n19659 ) | ( n19394 & n19659 ) ;
  assign n27445 = x17 & n5942 ;
  assign n27446 = n27445 ^ n19375 ^ 1'b0 ;
  assign n27450 = ~n2453 & n25801 ;
  assign n27451 = n27450 ^ n3838 ^ 1'b0 ;
  assign n27452 = ( n2391 & n3593 ) | ( n2391 & ~n8973 ) | ( n3593 & ~n8973 ) ;
  assign n27453 = n27451 & n27452 ;
  assign n27447 = n1353 | n6029 ;
  assign n27448 = n16710 ^ n13460 ^ 1'b0 ;
  assign n27449 = n27447 | n27448 ;
  assign n27454 = n27453 ^ n27449 ^ n25458 ;
  assign n27455 = n4764 & n27454 ;
  assign n27458 = n25454 ^ n1069 ^ n551 ;
  assign n27456 = n1008 | n10296 ;
  assign n27457 = n1905 & ~n27456 ;
  assign n27459 = n27458 ^ n27457 ^ 1'b0 ;
  assign n27460 = n563 & n22354 ;
  assign n27461 = n27460 ^ n14649 ^ 1'b0 ;
  assign n27462 = n4677 & ~n21399 ;
  assign n27465 = n25736 ^ n18252 ^ n8419 ;
  assign n27464 = n16130 ^ n10470 ^ n9545 ;
  assign n27463 = ~n4767 & n17404 ;
  assign n27466 = n27465 ^ n27464 ^ n27463 ;
  assign n27467 = ~n3609 & n20489 ;
  assign n27468 = n27467 ^ n12319 ^ 1'b0 ;
  assign n27469 = n13627 | n17958 ;
  assign n27470 = n27468 & ~n27469 ;
  assign n27471 = n2769 & ~n27470 ;
  assign n27472 = ~n7238 & n27471 ;
  assign n27478 = n3864 | n8134 ;
  assign n27479 = n27478 ^ n12120 ^ 1'b0 ;
  assign n27477 = ~n3163 & n4832 ;
  assign n27480 = n27479 ^ n27477 ^ 1'b0 ;
  assign n27474 = n11531 & ~n12946 ;
  assign n27475 = n21010 & n27474 ;
  assign n27473 = n5556 ^ n3993 ^ 1'b0 ;
  assign n27476 = n27475 ^ n27473 ^ 1'b0 ;
  assign n27481 = n27480 ^ n27476 ^ n5358 ;
  assign n27483 = n1199 & n15360 ;
  assign n27484 = n15449 & n27483 ;
  assign n27482 = n1443 & n21392 ;
  assign n27485 = n27484 ^ n27482 ^ n2734 ;
  assign n27486 = ~n8415 & n25662 ;
  assign n27487 = n7381 & ~n17192 ;
  assign n27488 = ~n11155 & n27487 ;
  assign n27489 = n8235 ^ n5353 ^ 1'b0 ;
  assign n27490 = n10790 & ~n27489 ;
  assign n27491 = n27490 ^ n9491 ^ n6160 ;
  assign n27492 = n27491 ^ n23695 ^ 1'b0 ;
  assign n27493 = n27488 | n27492 ;
  assign n27494 = n23277 ^ n16756 ^ 1'b0 ;
  assign n27495 = n10087 | n27494 ;
  assign n27496 = n7557 & ~n27495 ;
  assign n27497 = ( n7790 & n13072 ) | ( n7790 & n14591 ) | ( n13072 & n14591 ) ;
  assign n27498 = n27497 ^ n14345 ^ n7604 ;
  assign n27499 = n6066 & ~n27498 ;
  assign n27500 = n27499 ^ n10202 ^ 1'b0 ;
  assign n27501 = n1717 | n7909 ;
  assign n27502 = n18034 & ~n27501 ;
  assign n27503 = ( ~n871 & n25450 ) | ( ~n871 & n27502 ) | ( n25450 & n27502 ) ;
  assign n27504 = n3235 | n10608 ;
  assign n27505 = n2491 & ~n27504 ;
  assign n27506 = n27503 & n27505 ;
  assign n27509 = n12321 | n21085 ;
  assign n27510 = n15023 | n27509 ;
  assign n27507 = n2917 & n6389 ;
  assign n27508 = n27507 ^ n19068 ^ 1'b0 ;
  assign n27511 = n27510 ^ n27508 ^ n1832 ;
  assign n27512 = n19655 ^ n13561 ^ n2963 ;
  assign n27513 = ~n3521 & n6220 ;
  assign n27514 = n27513 ^ n7291 ^ 1'b0 ;
  assign n27515 = ( ~n1373 & n15429 ) | ( ~n1373 & n22918 ) | ( n15429 & n22918 ) ;
  assign n27516 = n19730 & n27515 ;
  assign n27517 = ( x124 & n27514 ) | ( x124 & ~n27516 ) | ( n27514 & ~n27516 ) ;
  assign n27518 = ( ~n15001 & n16371 ) | ( ~n15001 & n25331 ) | ( n16371 & n25331 ) ;
  assign n27519 = n5870 ^ n3012 ^ n1029 ;
  assign n27520 = n27519 ^ n8409 ^ n3088 ;
  assign n27521 = ( n25345 & n26243 ) | ( n25345 & ~n27520 ) | ( n26243 & ~n27520 ) ;
  assign n27522 = n20392 ^ n13275 ^ n1368 ;
  assign n27523 = n27522 ^ n18095 ^ 1'b0 ;
  assign n27524 = ~n23061 & n27523 ;
  assign n27525 = n19052 ^ n13378 ^ 1'b0 ;
  assign n27526 = ( n4034 & n19122 ) | ( n4034 & n22403 ) | ( n19122 & n22403 ) ;
  assign n27527 = n22375 ^ n11866 ^ 1'b0 ;
  assign n27528 = n3504 ^ n1612 ^ n211 ;
  assign n27529 = n12259 ^ n2542 ^ 1'b0 ;
  assign n27530 = n18680 ^ n12469 ^ 1'b0 ;
  assign n27531 = n10849 | n27530 ;
  assign n27532 = ~n5297 & n22467 ;
  assign n27533 = ( ~n2924 & n5439 ) | ( ~n2924 & n27532 ) | ( n5439 & n27532 ) ;
  assign n27534 = n27533 ^ n16865 ^ n5353 ;
  assign n27535 = n5199 | n10568 ;
  assign n27536 = n27535 ^ n16116 ^ 1'b0 ;
  assign n27539 = n12207 ^ n1471 ^ 1'b0 ;
  assign n27540 = n5155 & n27539 ;
  assign n27537 = n5745 ^ n3585 ^ 1'b0 ;
  assign n27538 = ~n15913 & n27537 ;
  assign n27541 = n27540 ^ n27538 ^ n2296 ;
  assign n27542 = n18647 | n25006 ;
  assign n27543 = ~n563 & n4129 ;
  assign n27546 = n4402 | n6254 ;
  assign n27544 = n14549 ^ n13484 ^ 1'b0 ;
  assign n27545 = ( n7165 & n15367 ) | ( n7165 & n27544 ) | ( n15367 & n27544 ) ;
  assign n27547 = n27546 ^ n27545 ^ n26993 ;
  assign n27548 = ( n9986 & n22628 ) | ( n9986 & n27547 ) | ( n22628 & n27547 ) ;
  assign n27549 = n27086 ^ n10058 ^ n2889 ;
  assign n27550 = n1617 & n6853 ;
  assign n27551 = n27550 ^ n20324 ^ 1'b0 ;
  assign n27552 = n1493 & ~n27551 ;
  assign n27553 = n27549 & n27552 ;
  assign n27554 = ~n1406 & n9704 ;
  assign n27555 = n27554 ^ n3932 ^ 1'b0 ;
  assign n27557 = n1301 | n21290 ;
  assign n27558 = n27557 ^ n992 ^ 1'b0 ;
  assign n27556 = n21936 & n27490 ;
  assign n27559 = n27558 ^ n27556 ^ 1'b0 ;
  assign n27560 = ~n24740 & n27559 ;
  assign n27561 = n9385 & n27560 ;
  assign n27562 = n16445 ^ n11221 ^ n3277 ;
  assign n27563 = ( n6987 & ~n17628 ) | ( n6987 & n27562 ) | ( ~n17628 & n27562 ) ;
  assign n27574 = n11130 ^ n7034 ^ n2344 ;
  assign n27575 = n27574 ^ n15796 ^ n12461 ;
  assign n27564 = n14897 | n18014 ;
  assign n27565 = ( n4286 & n8227 ) | ( n4286 & n16725 ) | ( n8227 & n16725 ) ;
  assign n27566 = n18094 ^ n16808 ^ n2186 ;
  assign n27567 = n293 & ~n5781 ;
  assign n27568 = ~n27566 & n27567 ;
  assign n27569 = n4775 | n13802 ;
  assign n27570 = ( n20161 & n27568 ) | ( n20161 & n27569 ) | ( n27568 & n27569 ) ;
  assign n27571 = n7143 & n27570 ;
  assign n27572 = n27571 ^ n8937 ^ 1'b0 ;
  assign n27573 = ( n27564 & ~n27565 ) | ( n27564 & n27572 ) | ( ~n27565 & n27572 ) ;
  assign n27576 = n27575 ^ n27573 ^ n23055 ;
  assign n27577 = n6978 & ~n24723 ;
  assign n27578 = n10499 ^ n4852 ^ 1'b0 ;
  assign n27579 = n27578 ^ n16706 ^ 1'b0 ;
  assign n27581 = n9639 & n27434 ;
  assign n27582 = ~n14072 & n27581 ;
  assign n27580 = ( n2916 & n4726 ) | ( n2916 & ~n12628 ) | ( n4726 & ~n12628 ) ;
  assign n27583 = n27582 ^ n27580 ^ n13928 ;
  assign n27584 = n20561 ^ n163 ^ 1'b0 ;
  assign n27585 = n13339 & ~n27584 ;
  assign n27586 = ~n10953 & n21246 ;
  assign n27587 = n3450 & n27586 ;
  assign n27588 = ~n27585 & n27587 ;
  assign n27589 = ( n15824 & n17218 ) | ( n15824 & n20751 ) | ( n17218 & n20751 ) ;
  assign n27590 = n27589 ^ n5053 ^ 1'b0 ;
  assign n27591 = x116 & n27590 ;
  assign n27592 = n19355 ^ n3565 ^ 1'b0 ;
  assign n27593 = ~n3579 & n27592 ;
  assign n27594 = ~n7863 & n12012 ;
  assign n27595 = n27594 ^ n18411 ^ 1'b0 ;
  assign n27596 = ( n2124 & ~n11576 ) | ( n2124 & n16369 ) | ( ~n11576 & n16369 ) ;
  assign n27597 = ( n6214 & ~n19134 ) | ( n6214 & n27596 ) | ( ~n19134 & n27596 ) ;
  assign n27598 = n14916 ^ n12916 ^ n3698 ;
  assign n27599 = ( n5119 & ~n7550 ) | ( n5119 & n8148 ) | ( ~n7550 & n8148 ) ;
  assign n27600 = ( n734 & n7085 ) | ( n734 & n27599 ) | ( n7085 & n27599 ) ;
  assign n27601 = n27600 ^ n7426 ^ 1'b0 ;
  assign n27602 = n7351 | n14424 ;
  assign n27603 = n3312 & ~n18778 ;
  assign n27604 = n6697 ^ n3445 ^ 1'b0 ;
  assign n27605 = n24997 ^ n22180 ^ 1'b0 ;
  assign n27606 = n20586 | n27605 ;
  assign n27607 = n5785 & n7291 ;
  assign n27608 = n27607 ^ n3495 ^ 1'b0 ;
  assign n27609 = n3700 & n27608 ;
  assign n27610 = n27609 ^ n8439 ^ 1'b0 ;
  assign n27611 = n4575 ^ n2882 ^ 1'b0 ;
  assign n27612 = n4011 & n27611 ;
  assign n27613 = n27612 ^ n11736 ^ n2456 ;
  assign n27614 = n22707 ^ n5681 ^ 1'b0 ;
  assign n27615 = n27613 & ~n27614 ;
  assign n27616 = n5674 | n15302 ;
  assign n27617 = n27616 ^ n25256 ^ 1'b0 ;
  assign n27618 = n27617 ^ n3755 ^ x63 ;
  assign n27622 = n8621 & ~n13788 ;
  assign n27623 = n12490 & n27622 ;
  assign n27619 = n16318 & ~n26439 ;
  assign n27620 = n27619 ^ n5536 ^ 1'b0 ;
  assign n27621 = ( n7954 & ~n22968 ) | ( n7954 & n27620 ) | ( ~n22968 & n27620 ) ;
  assign n27624 = n27623 ^ n27621 ^ n12270 ;
  assign n27625 = n1722 & ~n22185 ;
  assign n27626 = ~n11289 & n27625 ;
  assign n27627 = ( n1614 & n11491 ) | ( n1614 & n27626 ) | ( n11491 & n27626 ) ;
  assign n27628 = n5252 ^ n2153 ^ 1'b0 ;
  assign n27629 = n3048 & ~n27628 ;
  assign n27630 = n4503 ^ n2016 ^ n543 ;
  assign n27631 = ( n16402 & n27629 ) | ( n16402 & n27630 ) | ( n27629 & n27630 ) ;
  assign n27632 = ( n2704 & n27627 ) | ( n2704 & ~n27631 ) | ( n27627 & ~n27631 ) ;
  assign n27633 = n1896 & n8461 ;
  assign n27634 = n14199 ^ n5127 ^ 1'b0 ;
  assign n27635 = n12906 & n12961 ;
  assign n27636 = n27634 & n27635 ;
  assign n27637 = n27636 ^ n25184 ^ n15546 ;
  assign n27638 = n16250 ^ n8904 ^ 1'b0 ;
  assign n27639 = n24223 & ~n27638 ;
  assign n27640 = n20879 ^ n17086 ^ 1'b0 ;
  assign n27641 = ( x10 & ~n3973 ) | ( x10 & n6729 ) | ( ~n3973 & n6729 ) ;
  assign n27642 = n11774 & n27641 ;
  assign n27643 = n27642 ^ n3437 ^ 1'b0 ;
  assign n27644 = n1978 & n5454 ;
  assign n27645 = n27644 ^ n3343 ^ 1'b0 ;
  assign n27646 = ( n7436 & ~n15604 ) | ( n7436 & n18621 ) | ( ~n15604 & n18621 ) ;
  assign n27647 = n4490 ^ n3869 ^ n2141 ;
  assign n27648 = ( ~n14396 & n24365 ) | ( ~n14396 & n27647 ) | ( n24365 & n27647 ) ;
  assign n27649 = n26056 ^ n13112 ^ n2393 ;
  assign n27650 = ( n266 & n15665 ) | ( n266 & ~n27649 ) | ( n15665 & ~n27649 ) ;
  assign n27651 = ( n1772 & ~n2720 ) | ( n1772 & n27650 ) | ( ~n2720 & n27650 ) ;
  assign n27652 = n6022 ^ n3068 ^ x11 ;
  assign n27653 = n19534 ^ n14424 ^ n7853 ;
  assign n27654 = n27653 ^ n17925 ^ n4615 ;
  assign n27655 = n26753 ^ n22836 ^ 1'b0 ;
  assign n27656 = ~n6442 & n27655 ;
  assign n27657 = ~n10140 & n27656 ;
  assign n27658 = ~n23486 & n27657 ;
  assign n27659 = n2205 & ~n12885 ;
  assign n27660 = n9072 & n23873 ;
  assign n27661 = ~n14661 & n27660 ;
  assign n27662 = n15862 ^ n10466 ^ 1'b0 ;
  assign n27663 = ( ~n7952 & n8992 ) | ( ~n7952 & n19035 ) | ( n8992 & n19035 ) ;
  assign n27664 = n26551 ^ n12898 ^ 1'b0 ;
  assign n27665 = ~n21128 & n26102 ;
  assign n27666 = n27665 ^ n12384 ^ 1'b0 ;
  assign n27667 = n27666 ^ n19998 ^ n14096 ;
  assign n27668 = n19483 | n21674 ;
  assign n27669 = n27668 ^ n27422 ^ 1'b0 ;
  assign n27670 = n27669 ^ n20088 ^ 1'b0 ;
  assign n27671 = ~n9898 & n22387 ;
  assign n27672 = n25831 & n27671 ;
  assign n27673 = n12569 & n17130 ;
  assign n27674 = n1242 | n18314 ;
  assign n27675 = n26705 & ~n27674 ;
  assign n27676 = n23273 ^ n18679 ^ 1'b0 ;
  assign n27677 = ~n20188 & n27676 ;
  assign n27678 = n20015 ^ n13053 ^ n2867 ;
  assign n27679 = ( n7694 & n20864 ) | ( n7694 & n27678 ) | ( n20864 & n27678 ) ;
  assign n27680 = ( n16901 & n21838 ) | ( n16901 & n27679 ) | ( n21838 & n27679 ) ;
  assign n27681 = n17885 & n23242 ;
  assign n27682 = ( n4293 & ~n9676 ) | ( n4293 & n21630 ) | ( ~n9676 & n21630 ) ;
  assign n27683 = n4295 | n16928 ;
  assign n27684 = n20783 | n27683 ;
  assign n27685 = n27684 ^ n12931 ^ 1'b0 ;
  assign n27686 = n27682 & ~n27685 ;
  assign n27687 = ( ~n4059 & n9847 ) | ( ~n4059 & n22580 ) | ( n9847 & n22580 ) ;
  assign n27688 = n21887 ^ n14766 ^ n6265 ;
  assign n27689 = ( n4534 & n19451 ) | ( n4534 & n27688 ) | ( n19451 & n27688 ) ;
  assign n27690 = ~n4174 & n10344 ;
  assign n27691 = n2744 & n3787 ;
  assign n27692 = ~n27690 & n27691 ;
  assign n27693 = n6837 ^ n1166 ^ 1'b0 ;
  assign n27694 = n13304 & ~n19586 ;
  assign n27695 = n23923 ^ n19285 ^ 1'b0 ;
  assign n27696 = n1393 | n25241 ;
  assign n27697 = ~n540 & n17046 ;
  assign n27698 = n9427 ^ n6174 ^ n2474 ;
  assign n27699 = ~n27697 & n27698 ;
  assign n27700 = n21273 ^ n18778 ^ n15217 ;
  assign n27701 = n27700 ^ n19566 ^ n17920 ;
  assign n27702 = n7790 | n18427 ;
  assign n27703 = n27702 ^ n3745 ^ 1'b0 ;
  assign n27704 = n6533 & n27703 ;
  assign n27705 = n14627 ^ n7899 ^ 1'b0 ;
  assign n27706 = n2677 & ~n17967 ;
  assign n27707 = ( n5242 & ~n8640 ) | ( n5242 & n27244 ) | ( ~n8640 & n27244 ) ;
  assign n27708 = ~n8555 & n18278 ;
  assign n27709 = n25558 ^ n11286 ^ n6403 ;
  assign n27710 = n277 | n15028 ;
  assign n27711 = n9158 | n27710 ;
  assign n27712 = n27711 ^ n2073 ^ 1'b0 ;
  assign n27713 = n27712 ^ n11104 ^ 1'b0 ;
  assign n27714 = n20392 ^ n2928 ^ 1'b0 ;
  assign n27715 = n2978 & ~n27714 ;
  assign n27716 = ~n8093 & n15504 ;
  assign n27717 = ~n9227 & n25877 ;
  assign n27718 = ~n27716 & n27717 ;
  assign n27719 = n6811 ^ n950 ^ 1'b0 ;
  assign n27720 = n10945 & n27719 ;
  assign n27721 = n27720 ^ n7234 ^ 1'b0 ;
  assign n27724 = n23675 ^ n17917 ^ 1'b0 ;
  assign n27725 = n1843 & ~n27724 ;
  assign n27722 = n7701 ^ n6692 ^ 1'b0 ;
  assign n27723 = n14250 & ~n27722 ;
  assign n27726 = n27725 ^ n27723 ^ n18337 ;
  assign n27727 = n6601 | n9437 ;
  assign n27728 = n3676 & ~n27727 ;
  assign n27729 = ( ~n24924 & n26032 ) | ( ~n24924 & n27728 ) | ( n26032 & n27728 ) ;
  assign n27730 = n25947 ^ n7420 ^ 1'b0 ;
  assign n27731 = ( n2343 & ~n11691 ) | ( n2343 & n27730 ) | ( ~n11691 & n27730 ) ;
  assign n27732 = ( n1722 & n10283 ) | ( n1722 & ~n26038 ) | ( n10283 & ~n26038 ) ;
  assign n27737 = n14082 ^ n13451 ^ 1'b0 ;
  assign n27734 = n6123 ^ n3612 ^ n179 ;
  assign n27733 = ~n4440 & n15051 ;
  assign n27735 = n27734 ^ n27733 ^ 1'b0 ;
  assign n27736 = n27735 ^ n10338 ^ n1578 ;
  assign n27738 = n27737 ^ n27736 ^ n2767 ;
  assign n27739 = ~n1928 & n18376 ;
  assign n27740 = n27739 ^ n1228 ^ 1'b0 ;
  assign n27741 = n3556 & ~n23521 ;
  assign n27742 = n23755 & n27741 ;
  assign n27743 = n15893 ^ n5164 ^ n1486 ;
  assign n27744 = n3088 & n27743 ;
  assign n27745 = n17806 | n24013 ;
  assign n27746 = n19462 | n20110 ;
  assign n27747 = ( n3886 & n20738 ) | ( n3886 & ~n24127 ) | ( n20738 & ~n24127 ) ;
  assign n27748 = n21274 ^ n13767 ^ n6640 ;
  assign n27749 = ( n1285 & ~n3035 ) | ( n1285 & n27748 ) | ( ~n3035 & n27748 ) ;
  assign n27750 = ( n13421 & n14977 ) | ( n13421 & n27749 ) | ( n14977 & n27749 ) ;
  assign n27751 = n6794 ^ n824 ^ 1'b0 ;
  assign n27752 = n2804 & ~n27751 ;
  assign n27753 = n10767 | n27752 ;
  assign n27754 = ( n3050 & n21722 ) | ( n3050 & ~n27753 ) | ( n21722 & ~n27753 ) ;
  assign n27755 = n5948 & ~n15479 ;
  assign n27756 = n6039 | n27755 ;
  assign n27757 = n10499 | n27756 ;
  assign n27758 = n4576 | n27757 ;
  assign n27759 = n18827 ^ n3959 ^ 1'b0 ;
  assign n27760 = n12077 | n27759 ;
  assign n27761 = ~n1196 & n2060 ;
  assign n27762 = n27761 ^ n477 ^ 1'b0 ;
  assign n27763 = n1720 | n12217 ;
  assign n27764 = ( n13516 & ~n27762 ) | ( n13516 & n27763 ) | ( ~n27762 & n27763 ) ;
  assign n27765 = n27764 ^ n14312 ^ 1'b0 ;
  assign n27766 = n15892 | n27765 ;
  assign n27767 = n1890 & ~n18937 ;
  assign n27768 = n27767 ^ n14673 ^ 1'b0 ;
  assign n27769 = ~n5672 & n24799 ;
  assign n27774 = n4776 & n10608 ;
  assign n27775 = n27774 ^ n1468 ^ 1'b0 ;
  assign n27770 = ~n1553 & n9155 ;
  assign n27771 = n10015 & n27770 ;
  assign n27772 = ~n13152 & n27771 ;
  assign n27773 = n27772 ^ n12466 ^ n6090 ;
  assign n27776 = n27775 ^ n27773 ^ n24221 ;
  assign n27777 = n27776 ^ n22883 ^ n17328 ;
  assign n27778 = n15213 & n25285 ;
  assign n27779 = n27778 ^ n3991 ^ 1'b0 ;
  assign n27780 = n27779 ^ n13920 ^ n11510 ;
  assign n27785 = ~n9761 & n10475 ;
  assign n27786 = ~n5333 & n27785 ;
  assign n27782 = ( n3254 & n14531 ) | ( n3254 & n15707 ) | ( n14531 & n15707 ) ;
  assign n27781 = ~n924 & n3599 ;
  assign n27783 = n27782 ^ n27781 ^ n13735 ;
  assign n27784 = ( n11162 & ~n12374 ) | ( n11162 & n27783 ) | ( ~n12374 & n27783 ) ;
  assign n27787 = n27786 ^ n27784 ^ n16911 ;
  assign n27788 = n1900 | n20764 ;
  assign n27789 = ( n6353 & n9764 ) | ( n6353 & ~n27788 ) | ( n9764 & ~n27788 ) ;
  assign n27790 = n27789 ^ n20849 ^ 1'b0 ;
  assign n27791 = n6555 | n27790 ;
  assign n27792 = ~n22481 & n24776 ;
  assign n27793 = ~n20820 & n27792 ;
  assign n27794 = n5836 & n8374 ;
  assign n27795 = ( n1371 & n4976 ) | ( n1371 & ~n5165 ) | ( n4976 & ~n5165 ) ;
  assign n27796 = n16296 ^ n15980 ^ n803 ;
  assign n27797 = n27796 ^ n6910 ^ 1'b0 ;
  assign n27798 = n27795 & n27797 ;
  assign n27799 = n11523 ^ n929 ^ 1'b0 ;
  assign n27800 = x52 & ~n27799 ;
  assign n27801 = n27800 ^ n15860 ^ n849 ;
  assign n27802 = ( ~n9667 & n12360 ) | ( ~n9667 & n16765 ) | ( n12360 & n16765 ) ;
  assign n27803 = n16276 ^ n2273 ^ 1'b0 ;
  assign n27804 = ~n18692 & n27803 ;
  assign n27805 = n22458 ^ n2881 ^ 1'b0 ;
  assign n27806 = n16787 & ~n16902 ;
  assign n27807 = n27806 ^ n10516 ^ 1'b0 ;
  assign n27808 = ( n8240 & n17228 ) | ( n8240 & ~n23339 ) | ( n17228 & ~n23339 ) ;
  assign n27809 = n14804 & ~n27808 ;
  assign n27810 = n27809 ^ n11412 ^ 1'b0 ;
  assign n27811 = ~n4994 & n9757 ;
  assign n27812 = n1624 & n27811 ;
  assign n27813 = n16780 ^ n7396 ^ n1601 ;
  assign n27814 = ( ~n5319 & n7160 ) | ( ~n5319 & n18994 ) | ( n7160 & n18994 ) ;
  assign n27815 = n27814 ^ n17488 ^ n11297 ;
  assign n27816 = n20097 & n27815 ;
  assign n27817 = n4601 ^ x23 ^ 1'b0 ;
  assign n27818 = ~n13828 & n27817 ;
  assign n27819 = n18416 | n18684 ;
  assign n27820 = n7152 ^ n6824 ^ n836 ;
  assign n27821 = n4701 & n15965 ;
  assign n27822 = ~n4868 & n27821 ;
  assign n27823 = n16305 ^ n10501 ^ 1'b0 ;
  assign n27824 = n25042 ^ n5689 ^ 1'b0 ;
  assign n27825 = n3193 | n27824 ;
  assign n27826 = n7059 ^ n5403 ^ 1'b0 ;
  assign n27827 = n12222 ^ n7979 ^ n3691 ;
  assign n27828 = ( ~n13250 & n27826 ) | ( ~n13250 & n27827 ) | ( n27826 & n27827 ) ;
  assign n27829 = ( n2428 & n10174 ) | ( n2428 & ~n14824 ) | ( n10174 & ~n14824 ) ;
  assign n27830 = ~n17245 & n27829 ;
  assign n27831 = ( n27825 & n27828 ) | ( n27825 & n27830 ) | ( n27828 & n27830 ) ;
  assign n27832 = n20614 ^ n8711 ^ 1'b0 ;
  assign n27833 = n23568 & ~n27832 ;
  assign n27834 = n12559 & ~n21620 ;
  assign n27835 = n1815 & ~n12763 ;
  assign n27843 = n23289 ^ n10530 ^ n2567 ;
  assign n27838 = n23606 ^ n5478 ^ 1'b0 ;
  assign n27839 = n3973 & ~n27838 ;
  assign n27840 = ~n7423 & n27839 ;
  assign n27841 = n8919 & n27840 ;
  assign n27836 = n9252 | n10348 ;
  assign n27837 = n27836 ^ n15411 ^ 1'b0 ;
  assign n27842 = n27841 ^ n27837 ^ n4324 ;
  assign n27844 = n27843 ^ n27842 ^ n6811 ;
  assign n27845 = x102 & ~n21356 ;
  assign n27846 = n7893 & n25631 ;
  assign n27847 = n4332 | n6529 ;
  assign n27848 = n11886 & ~n27847 ;
  assign n27849 = ( n2390 & n3385 ) | ( n2390 & n23752 ) | ( n3385 & n23752 ) ;
  assign n27850 = ~n6075 & n7415 ;
  assign n27851 = n27850 ^ n252 ^ 1'b0 ;
  assign n27852 = ( n217 & ~n21804 ) | ( n217 & n27851 ) | ( ~n21804 & n27851 ) ;
  assign n27853 = ( ~n8190 & n8331 ) | ( ~n8190 & n27852 ) | ( n8331 & n27852 ) ;
  assign n27854 = ( ~n1850 & n1925 ) | ( ~n1850 & n19239 ) | ( n1925 & n19239 ) ;
  assign n27855 = ( n10452 & ~n22194 ) | ( n10452 & n26002 ) | ( ~n22194 & n26002 ) ;
  assign n27856 = n27855 ^ n8141 ^ n6558 ;
  assign n27857 = n5968 ^ n5358 ^ n1790 ;
  assign n27858 = n27857 ^ n20871 ^ n5009 ;
  assign n27859 = n23984 ^ n17060 ^ 1'b0 ;
  assign n27860 = n17041 ^ n6937 ^ 1'b0 ;
  assign n27861 = n1334 & n27860 ;
  assign n27862 = n4839 ^ n657 ^ 1'b0 ;
  assign n27863 = n27861 & n27862 ;
  assign n27864 = ( n133 & n2948 ) | ( n133 & n26219 ) | ( n2948 & n26219 ) ;
  assign n27865 = n3598 & n27255 ;
  assign n27866 = n27865 ^ n16574 ^ 1'b0 ;
  assign n27867 = ( ~n6072 & n21985 ) | ( ~n6072 & n27866 ) | ( n21985 & n27866 ) ;
  assign n27868 = n11592 ^ n7920 ^ n5308 ;
  assign n27869 = n11950 ^ n5951 ^ n2857 ;
  assign n27870 = n9883 ^ n6861 ^ 1'b0 ;
  assign n27871 = n23667 | n27870 ;
  assign n27872 = n27871 ^ n11799 ^ n8167 ;
  assign n27873 = ( n27868 & ~n27869 ) | ( n27868 & n27872 ) | ( ~n27869 & n27872 ) ;
  assign n27874 = n2168 | n6719 ;
  assign n27875 = n19283 & ~n27874 ;
  assign n27876 = n27875 ^ n18771 ^ n7142 ;
  assign n27877 = ( n20987 & ~n21716 ) | ( n20987 & n27876 ) | ( ~n21716 & n27876 ) ;
  assign n27878 = ( n8348 & n26530 ) | ( n8348 & n27877 ) | ( n26530 & n27877 ) ;
  assign n27879 = n330 & ~n10280 ;
  assign n27880 = ~n1336 & n27879 ;
  assign n27888 = n22365 ^ n22079 ^ n3242 ;
  assign n27886 = n2980 | n10151 ;
  assign n27887 = n27886 ^ n19674 ^ 1'b0 ;
  assign n27881 = ( ~x19 & n10409 ) | ( ~x19 & n15690 ) | ( n10409 & n15690 ) ;
  assign n27882 = n15330 ^ n9078 ^ n5770 ;
  assign n27883 = n5711 & ~n7919 ;
  assign n27884 = n27883 ^ n22927 ^ 1'b0 ;
  assign n27885 = ( n27881 & n27882 ) | ( n27881 & ~n27884 ) | ( n27882 & ~n27884 ) ;
  assign n27889 = n27888 ^ n27887 ^ n27885 ;
  assign n27890 = ( ~n24496 & n27880 ) | ( ~n24496 & n27889 ) | ( n27880 & n27889 ) ;
  assign n27891 = n16780 ^ n7414 ^ 1'b0 ;
  assign n27892 = n11504 | n27891 ;
  assign n27893 = n12586 ^ n9926 ^ n364 ;
  assign n27894 = n16681 | n27893 ;
  assign n27895 = ~n729 & n5741 ;
  assign n27896 = n16030 & ~n27895 ;
  assign n27897 = n8753 ^ n7156 ^ 1'b0 ;
  assign n27898 = ~n14965 & n16488 ;
  assign n27899 = n14561 ^ n4807 ^ x52 ;
  assign n27900 = n27899 ^ n19482 ^ 1'b0 ;
  assign n27902 = n22535 ^ x33 ^ 1'b0 ;
  assign n27901 = n11772 & ~n19719 ;
  assign n27903 = n27902 ^ n27901 ^ n19859 ;
  assign n27904 = n17827 ^ n6385 ^ 1'b0 ;
  assign n27905 = n27904 ^ n10165 ^ n4788 ;
  assign n27906 = n8994 ^ n2377 ^ 1'b0 ;
  assign n27907 = n3617 | n13071 ;
  assign n27908 = n2204 | n27907 ;
  assign n27909 = n12169 & n27908 ;
  assign n27910 = n27909 ^ n3914 ^ 1'b0 ;
  assign n27911 = n7085 & ~n27910 ;
  assign n27912 = ~n11242 & n16171 ;
  assign n27913 = ~n23555 & n27912 ;
  assign n27914 = n1095 & n27913 ;
  assign n27915 = ~n3847 & n4697 ;
  assign n27916 = ( n7322 & ~n9771 ) | ( n7322 & n15893 ) | ( ~n9771 & n15893 ) ;
  assign n27917 = n17861 | n27916 ;
  assign n27918 = n12628 & ~n27917 ;
  assign n27919 = n27918 ^ n14139 ^ 1'b0 ;
  assign n27920 = n25524 ^ n8393 ^ 1'b0 ;
  assign n27921 = ( n402 & n19917 ) | ( n402 & n27920 ) | ( n19917 & n27920 ) ;
  assign n27922 = n3118 & n9562 ;
  assign n27923 = ( n3392 & n14140 ) | ( n3392 & ~n27922 ) | ( n14140 & ~n27922 ) ;
  assign n27924 = n10769 ^ n8094 ^ n4040 ;
  assign n27925 = n27924 ^ n27329 ^ n20283 ;
  assign n27926 = n11925 ^ n9643 ^ n8534 ;
  assign n27927 = n1234 | n27926 ;
  assign n27928 = n26648 ^ n14052 ^ 1'b0 ;
  assign n27929 = n13657 & ~n27928 ;
  assign n27930 = ( n11341 & n11983 ) | ( n11341 & ~n25770 ) | ( n11983 & ~n25770 ) ;
  assign n27931 = n342 & n27930 ;
  assign n27932 = n20868 & n27931 ;
  assign n27933 = n14472 & n16125 ;
  assign n27934 = ~n19118 & n27933 ;
  assign n27935 = n18122 ^ n13116 ^ 1'b0 ;
  assign n27936 = n6740 | n27935 ;
  assign n27937 = n27936 ^ n20631 ^ 1'b0 ;
  assign n27938 = n3195 | n20934 ;
  assign n27939 = ( n5569 & ~n17298 ) | ( n5569 & n27938 ) | ( ~n17298 & n27938 ) ;
  assign n27940 = n9198 ^ n1958 ^ 1'b0 ;
  assign n27941 = n19616 ^ n17876 ^ n17836 ;
  assign n27942 = ~n9037 & n27941 ;
  assign n27943 = n13799 ^ n3806 ^ n967 ;
  assign n27944 = n27943 ^ n11457 ^ n8003 ;
  assign n27945 = n22447 ^ n20131 ^ n8971 ;
  assign n27946 = ( n7880 & ~n27944 ) | ( n7880 & n27945 ) | ( ~n27944 & n27945 ) ;
  assign n27947 = n6903 | n12521 ;
  assign n27948 = n27947 ^ n5775 ^ 1'b0 ;
  assign n27949 = n27948 ^ n26334 ^ 1'b0 ;
  assign n27950 = n3248 & ~n3282 ;
  assign n27951 = ~n14589 & n27950 ;
  assign n27952 = n27951 ^ n7808 ^ 1'b0 ;
  assign n27953 = n10916 ^ n649 ^ 1'b0 ;
  assign n27954 = n988 | n27953 ;
  assign n27955 = n3186 & n13292 ;
  assign n27956 = n27955 ^ n6375 ^ 1'b0 ;
  assign n27957 = n19543 ^ n6079 ^ 1'b0 ;
  assign n27958 = ( n10551 & n21756 ) | ( n10551 & ~n27957 ) | ( n21756 & ~n27957 ) ;
  assign n27959 = n27958 ^ n7774 ^ n966 ;
  assign n27960 = ~n2438 & n7665 ;
  assign n27961 = n27960 ^ n18829 ^ 1'b0 ;
  assign n27962 = ( n12529 & n19045 ) | ( n12529 & n27961 ) | ( n19045 & n27961 ) ;
  assign n27963 = n7187 & n9307 ;
  assign n27964 = ( n7853 & n18762 ) | ( n7853 & ~n27963 ) | ( n18762 & ~n27963 ) ;
  assign n27965 = n17686 ^ n8479 ^ 1'b0 ;
  assign n27966 = n7292 & n27965 ;
  assign n27967 = n10219 ^ n6545 ^ 1'b0 ;
  assign n27968 = n27966 & ~n27967 ;
  assign n27969 = n27968 ^ n26803 ^ n18286 ;
  assign n27970 = n27969 ^ n9022 ^ n5146 ;
  assign n27971 = ( n2210 & n8478 ) | ( n2210 & n14868 ) | ( n8478 & n14868 ) ;
  assign n27972 = n25484 ^ n16670 ^ 1'b0 ;
  assign n27973 = n10721 ^ n3620 ^ 1'b0 ;
  assign n27974 = n22665 ^ n10438 ^ 1'b0 ;
  assign n27975 = n27973 & n27974 ;
  assign n27976 = n481 | n6913 ;
  assign n27977 = n27976 ^ n19077 ^ 1'b0 ;
  assign n27978 = n8599 & ~n13367 ;
  assign n27979 = n27978 ^ n3037 ^ 1'b0 ;
  assign n27980 = n15494 ^ n6945 ^ 1'b0 ;
  assign n27981 = n821 & ~n27980 ;
  assign n27982 = ( ~n3919 & n27979 ) | ( ~n3919 & n27981 ) | ( n27979 & n27981 ) ;
  assign n27983 = n1340 | n5913 ;
  assign n27984 = n27983 ^ n24339 ^ n5276 ;
  assign n27986 = ~n1742 & n9890 ;
  assign n27987 = n2863 & n27986 ;
  assign n27985 = n1854 | n20466 ;
  assign n27988 = n27987 ^ n27985 ^ n211 ;
  assign n27989 = ( n7842 & n14227 ) | ( n7842 & n23339 ) | ( n14227 & n23339 ) ;
  assign n27990 = n21919 ^ n10369 ^ 1'b0 ;
  assign n27991 = ( n6598 & ~n27989 ) | ( n6598 & n27990 ) | ( ~n27989 & n27990 ) ;
  assign n27992 = ( x111 & n2033 ) | ( x111 & ~n18404 ) | ( n2033 & ~n18404 ) ;
  assign n27993 = n27992 ^ n19737 ^ n10742 ;
  assign n27994 = n27993 ^ n7684 ^ 1'b0 ;
  assign n27995 = n9438 | n17166 ;
  assign n27996 = n27995 ^ n19350 ^ 1'b0 ;
  assign n27997 = ~n10568 & n26200 ;
  assign n27998 = n27997 ^ n778 ^ 1'b0 ;
  assign n27999 = n26128 ^ n15928 ^ 1'b0 ;
  assign n28000 = n11443 ^ n10505 ^ 1'b0 ;
  assign n28001 = n10988 ^ n10702 ^ n2962 ;
  assign n28002 = ~n13304 & n28001 ;
  assign n28003 = n28002 ^ n5403 ^ 1'b0 ;
  assign n28004 = x66 & ~n1996 ;
  assign n28005 = ~n8500 & n9455 ;
  assign n28006 = n28005 ^ n19507 ^ 1'b0 ;
  assign n28007 = ( ~n28003 & n28004 ) | ( ~n28003 & n28006 ) | ( n28004 & n28006 ) ;
  assign n28008 = n10377 ^ n7993 ^ n7639 ;
  assign n28009 = n24842 & n26787 ;
  assign n28010 = n13780 ^ n3835 ^ 1'b0 ;
  assign n28011 = ~n11794 & n25202 ;
  assign n28012 = n4157 & ~n20928 ;
  assign n28013 = n28012 ^ n2246 ^ 1'b0 ;
  assign n28014 = ~n3775 & n10893 ;
  assign n28015 = n28013 & n28014 ;
  assign n28016 = ~n249 & n28015 ;
  assign n28017 = ( n5741 & ~n14495 ) | ( n5741 & n28016 ) | ( ~n14495 & n28016 ) ;
  assign n28018 = n7952 ^ n3519 ^ 1'b0 ;
  assign n28019 = n4724 & n10214 ;
  assign n28020 = n28019 ^ n1924 ^ 1'b0 ;
  assign n28021 = ( n6335 & n28018 ) | ( n6335 & n28020 ) | ( n28018 & n28020 ) ;
  assign n28022 = n5613 ^ n3033 ^ n2845 ;
  assign n28023 = n8362 ^ n3638 ^ 1'b0 ;
  assign n28024 = n8388 & n28023 ;
  assign n28025 = n2137 & n28024 ;
  assign n28026 = n24055 & n28025 ;
  assign n28027 = ( n17435 & ~n28022 ) | ( n17435 & n28026 ) | ( ~n28022 & n28026 ) ;
  assign n28028 = n15992 & n26931 ;
  assign n28029 = ~n9176 & n28028 ;
  assign n28030 = n5739 | n8973 ;
  assign n28031 = n10788 | n28030 ;
  assign n28032 = n5991 & ~n28031 ;
  assign n28033 = ( n268 & ~n28029 ) | ( n268 & n28032 ) | ( ~n28029 & n28032 ) ;
  assign n28034 = ( n6924 & n11028 ) | ( n6924 & ~n14934 ) | ( n11028 & ~n14934 ) ;
  assign n28035 = n28034 ^ n13535 ^ n6091 ;
  assign n28036 = ( ~n13777 & n15554 ) | ( ~n13777 & n23210 ) | ( n15554 & n23210 ) ;
  assign n28037 = n910 | n28036 ;
  assign n28038 = n15321 ^ n4307 ^ 1'b0 ;
  assign n28039 = ( n1496 & n6556 ) | ( n1496 & n13411 ) | ( n6556 & n13411 ) ;
  assign n28040 = n28039 ^ n21757 ^ 1'b0 ;
  assign n28041 = n15598 | n28040 ;
  assign n28042 = n28041 ^ n25324 ^ 1'b0 ;
  assign n28043 = n21371 ^ n236 ^ 1'b0 ;
  assign n28046 = ( ~n10193 & n17320 ) | ( ~n10193 & n26467 ) | ( n17320 & n26467 ) ;
  assign n28044 = ( n3287 & n4056 ) | ( n3287 & n13323 ) | ( n4056 & n13323 ) ;
  assign n28045 = ~n1805 & n28044 ;
  assign n28047 = n28046 ^ n28045 ^ 1'b0 ;
  assign n28048 = ( n794 & ~n10406 ) | ( n794 & n23192 ) | ( ~n10406 & n23192 ) ;
  assign n28049 = ( n1129 & n4063 ) | ( n1129 & ~n5516 ) | ( n4063 & ~n5516 ) ;
  assign n28050 = ( n6587 & ~n13295 ) | ( n6587 & n28049 ) | ( ~n13295 & n28049 ) ;
  assign n28052 = n343 & ~n6918 ;
  assign n28051 = ( n7662 & n8707 ) | ( n7662 & n13769 ) | ( n8707 & n13769 ) ;
  assign n28053 = n28052 ^ n28051 ^ n18429 ;
  assign n28054 = n28053 ^ n2840 ^ n1226 ;
  assign n28055 = ( n1294 & n4336 ) | ( n1294 & ~n5522 ) | ( n4336 & ~n5522 ) ;
  assign n28056 = n28055 ^ n17526 ^ 1'b0 ;
  assign n28057 = ~n26808 & n28056 ;
  assign n28058 = n1626 & n15657 ;
  assign n28059 = n28058 ^ n16537 ^ n16300 ;
  assign n28060 = n3644 & n8860 ;
  assign n28061 = n28060 ^ n17651 ^ 1'b0 ;
  assign n28062 = n18134 ^ n15077 ^ 1'b0 ;
  assign n28063 = ( n14777 & ~n28061 ) | ( n14777 & n28062 ) | ( ~n28061 & n28062 ) ;
  assign n28064 = n2659 | n5764 ;
  assign n28065 = n28064 ^ n19632 ^ 1'b0 ;
  assign n28066 = n13068 & n22906 ;
  assign n28067 = n28066 ^ n5853 ^ 1'b0 ;
  assign n28068 = ( n5545 & n11892 ) | ( n5545 & n11976 ) | ( n11892 & n11976 ) ;
  assign n28069 = ~n5792 & n6337 ;
  assign n28070 = ( n453 & ~n14799 ) | ( n453 & n24893 ) | ( ~n14799 & n24893 ) ;
  assign n28071 = n23599 ^ n9335 ^ 1'b0 ;
  assign n28073 = n11346 ^ n5453 ^ 1'b0 ;
  assign n28072 = ( ~n6104 & n10364 ) | ( ~n6104 & n18692 ) | ( n10364 & n18692 ) ;
  assign n28074 = n28073 ^ n28072 ^ n11932 ;
  assign n28076 = n15938 & n18848 ;
  assign n28075 = ~n6949 & n25466 ;
  assign n28077 = n28076 ^ n28075 ^ 1'b0 ;
  assign n28078 = n7912 ^ n2049 ^ x34 ;
  assign n28079 = n28078 ^ n1947 ^ 1'b0 ;
  assign n28080 = n28077 & n28079 ;
  assign n28081 = n24726 ^ n24156 ^ n1257 ;
  assign n28082 = ( ~n2254 & n12094 ) | ( ~n2254 & n28081 ) | ( n12094 & n28081 ) ;
  assign n28083 = n19730 ^ n16256 ^ n12311 ;
  assign n28084 = n20624 & ~n28083 ;
  assign n28085 = ~n28082 & n28084 ;
  assign n28089 = ( n5288 & n10090 ) | ( n5288 & ~n14057 ) | ( n10090 & ~n14057 ) ;
  assign n28086 = n13479 ^ n1021 ^ 1'b0 ;
  assign n28087 = n12774 & ~n28086 ;
  assign n28088 = ( ~n9501 & n17578 ) | ( ~n9501 & n28087 ) | ( n17578 & n28087 ) ;
  assign n28090 = n28089 ^ n28088 ^ n4966 ;
  assign n28091 = ( n2646 & n12283 ) | ( n2646 & ~n13222 ) | ( n12283 & ~n13222 ) ;
  assign n28092 = n13535 ^ n912 ^ n770 ;
  assign n28093 = n28092 ^ n18614 ^ x33 ;
  assign n28094 = ( n5235 & n28091 ) | ( n5235 & ~n28093 ) | ( n28091 & ~n28093 ) ;
  assign n28095 = ( n2632 & n18937 ) | ( n2632 & n28094 ) | ( n18937 & n28094 ) ;
  assign n28096 = n9830 ^ n3182 ^ 1'b0 ;
  assign n28097 = ( n21489 & n27060 ) | ( n21489 & n28096 ) | ( n27060 & n28096 ) ;
  assign n28098 = n12306 & ~n19971 ;
  assign n28099 = ( n3251 & n5324 ) | ( n3251 & n20265 ) | ( n5324 & n20265 ) ;
  assign n28100 = n19706 ^ n5613 ^ n3704 ;
  assign n28101 = ~n5476 & n28100 ;
  assign n28102 = n5064 | n12320 ;
  assign n28103 = n5467 & ~n28102 ;
  assign n28104 = n15184 ^ n14765 ^ 1'b0 ;
  assign n28105 = n11232 ^ n1379 ^ 1'b0 ;
  assign n28113 = n2026 ^ n1295 ^ 1'b0 ;
  assign n28114 = n1608 & n28113 ;
  assign n28112 = n27468 ^ n16364 ^ n293 ;
  assign n28107 = n18363 ^ n17066 ^ 1'b0 ;
  assign n28106 = n25705 ^ n19117 ^ n8630 ;
  assign n28108 = n28107 ^ n28106 ^ n2436 ;
  assign n28109 = n9541 & n28108 ;
  assign n28110 = n28109 ^ n9034 ^ 1'b0 ;
  assign n28111 = ( ~x90 & n22115 ) | ( ~x90 & n28110 ) | ( n22115 & n28110 ) ;
  assign n28115 = n28114 ^ n28112 ^ n28111 ;
  assign n28116 = n20135 ^ n13948 ^ n7051 ;
  assign n28117 = ( ~n3971 & n21406 ) | ( ~n3971 & n28116 ) | ( n21406 & n28116 ) ;
  assign n28118 = n17082 ^ n15898 ^ n836 ;
  assign n28119 = n3576 ^ n2210 ^ n2079 ;
  assign n28120 = n28119 ^ n13893 ^ 1'b0 ;
  assign n28121 = n5856 ^ n1330 ^ 1'b0 ;
  assign n28122 = n28121 ^ n18048 ^ n1127 ;
  assign n28123 = n6467 ^ n2178 ^ 1'b0 ;
  assign n28124 = n22373 | n28123 ;
  assign n28125 = ~n12190 & n14764 ;
  assign n28126 = n28125 ^ n18367 ^ 1'b0 ;
  assign n28127 = n22774 ^ n20429 ^ x120 ;
  assign n28128 = ( ~n2881 & n3183 ) | ( ~n2881 & n15667 ) | ( n3183 & n15667 ) ;
  assign n28129 = ~n27377 & n28128 ;
  assign n28130 = n22479 & n28129 ;
  assign n28131 = n18995 ^ n9385 ^ n996 ;
  assign n28132 = n3076 & ~n13629 ;
  assign n28133 = n28132 ^ n11985 ^ 1'b0 ;
  assign n28134 = ~n8912 & n28133 ;
  assign n28135 = ~n13498 & n28134 ;
  assign n28136 = n18887 ^ n8857 ^ n5240 ;
  assign n28137 = ( n8219 & n25929 ) | ( n8219 & ~n26001 ) | ( n25929 & ~n26001 ) ;
  assign n28139 = n12293 ^ n6941 ^ 1'b0 ;
  assign n28138 = n18251 & ~n24663 ;
  assign n28140 = n28139 ^ n28138 ^ 1'b0 ;
  assign n28141 = n16936 | n20623 ;
  assign n28142 = n18656 & ~n28141 ;
  assign n28143 = n26706 ^ n11782 ^ n7472 ;
  assign n28144 = n11714 ^ n9741 ^ 1'b0 ;
  assign n28145 = n3784 | n28144 ;
  assign n28146 = ( n4546 & n8087 ) | ( n4546 & n28145 ) | ( n8087 & n28145 ) ;
  assign n28147 = n23809 ^ n7227 ^ n2138 ;
  assign n28148 = n8072 ^ n5536 ^ n4919 ;
  assign n28149 = n1693 & n13667 ;
  assign n28150 = ~n6517 & n28149 ;
  assign n28151 = ~n2304 & n28150 ;
  assign n28152 = n8959 | n14809 ;
  assign n28153 = ( n5478 & n16983 ) | ( n5478 & n28152 ) | ( n16983 & n28152 ) ;
  assign n28154 = n28151 & ~n28153 ;
  assign n28155 = n15402 ^ n8007 ^ n1466 ;
  assign n28156 = n3053 & ~n28155 ;
  assign n28157 = n9521 ^ n8978 ^ 1'b0 ;
  assign n28158 = ~n12996 & n28157 ;
  assign n28159 = n1036 & n18518 ;
  assign n28160 = ~n2016 & n28159 ;
  assign n28161 = n16827 | n28160 ;
  assign n28162 = n28161 ^ n11473 ^ 1'b0 ;
  assign n28163 = ~n23120 & n28162 ;
  assign n28164 = n28163 ^ n6070 ^ 1'b0 ;
  assign n28165 = n14236 ^ n12356 ^ 1'b0 ;
  assign n28166 = n15143 & ~n28165 ;
  assign n28167 = ( n1179 & n1621 ) | ( n1179 & n6905 ) | ( n1621 & n6905 ) ;
  assign n28168 = n11892 ^ n8378 ^ n7307 ;
  assign n28169 = n28168 ^ n10915 ^ 1'b0 ;
  assign n28170 = ( n18726 & n28167 ) | ( n18726 & n28169 ) | ( n28167 & n28169 ) ;
  assign n28171 = n702 | n13635 ;
  assign n28172 = n28171 ^ n23039 ^ 1'b0 ;
  assign n28173 = n28172 ^ n25022 ^ 1'b0 ;
  assign n28174 = n26404 ^ n25770 ^ n8251 ;
  assign n28175 = n13425 | n22005 ;
  assign n28176 = n28175 ^ n13004 ^ n11670 ;
  assign n28177 = ( ~n7024 & n11628 ) | ( ~n7024 & n12104 ) | ( n11628 & n12104 ) ;
  assign n28178 = ~n20658 & n27436 ;
  assign n28179 = n28178 ^ n8062 ^ 1'b0 ;
  assign n28180 = n25092 ^ n7713 ^ 1'b0 ;
  assign n28181 = n5693 | n28180 ;
  assign n28182 = n3450 & n8026 ;
  assign n28183 = n21983 ^ n20615 ^ n8352 ;
  assign n28184 = n27909 & n28183 ;
  assign n28185 = ~n4321 & n28184 ;
  assign n28186 = ( n19711 & ~n24795 ) | ( n19711 & n28185 ) | ( ~n24795 & n28185 ) ;
  assign n28187 = n18714 ^ n16437 ^ 1'b0 ;
  assign n28188 = n19566 ^ n18450 ^ n1827 ;
  assign n28191 = ~n764 & n5144 ;
  assign n28192 = n28191 ^ n19900 ^ 1'b0 ;
  assign n28189 = n17147 ^ n1001 ^ 1'b0 ;
  assign n28190 = n253 & n28189 ;
  assign n28193 = n28192 ^ n28190 ^ n13918 ;
  assign n28194 = ~n4393 & n28193 ;
  assign n28195 = n11686 | n12319 ;
  assign n28196 = n5485 | n28195 ;
  assign n28197 = n3389 | n28196 ;
  assign n28198 = n12739 ^ n2073 ^ 1'b0 ;
  assign n28199 = n8667 & ~n28198 ;
  assign n28200 = ( ~n9689 & n16190 ) | ( ~n9689 & n28199 ) | ( n16190 & n28199 ) ;
  assign n28201 = n13936 | n21866 ;
  assign n28202 = n28200 | n28201 ;
  assign n28203 = n20846 ^ n4462 ^ 1'b0 ;
  assign n28204 = n4151 ^ n4114 ^ 1'b0 ;
  assign n28205 = n9479 ^ n8290 ^ n7366 ;
  assign n28206 = n549 & n7732 ;
  assign n28207 = ~n15835 & n28206 ;
  assign n28208 = ( n7783 & n28205 ) | ( n7783 & n28207 ) | ( n28205 & n28207 ) ;
  assign n28210 = x7 & n2809 ;
  assign n28211 = n2653 & n28210 ;
  assign n28212 = ( n1878 & ~n12218 ) | ( n1878 & n28211 ) | ( ~n12218 & n28211 ) ;
  assign n28209 = ~n12915 & n22716 ;
  assign n28213 = n28212 ^ n28209 ^ 1'b0 ;
  assign n28214 = n11646 ^ n1304 ^ 1'b0 ;
  assign n28215 = n14690 & ~n28214 ;
  assign n28216 = ( ~n1523 & n16859 ) | ( ~n1523 & n28215 ) | ( n16859 & n28215 ) ;
  assign n28217 = n27196 & n28216 ;
  assign n28218 = n28217 ^ n988 ^ 1'b0 ;
  assign n28219 = n3438 & ~n18810 ;
  assign n28220 = ~n9207 & n28219 ;
  assign n28221 = n3370 | n27491 ;
  assign n28222 = n2195 | n28221 ;
  assign n28223 = n12417 ^ n7177 ^ 1'b0 ;
  assign n28224 = n19177 & ~n28223 ;
  assign n28225 = n28224 ^ n17805 ^ 1'b0 ;
  assign n28226 = ( ~n5425 & n5815 ) | ( ~n5425 & n17355 ) | ( n5815 & n17355 ) ;
  assign n28227 = n27566 ^ n25860 ^ n2501 ;
  assign n28228 = n8609 | n15961 ;
  assign n28229 = n28228 ^ n26175 ^ n24618 ;
  assign n28230 = n10661 & ~n16250 ;
  assign n28231 = n11574 & n28230 ;
  assign n28232 = ( n1404 & ~n22561 ) | ( n1404 & n28231 ) | ( ~n22561 & n28231 ) ;
  assign n28233 = n18135 ^ n4923 ^ 1'b0 ;
  assign n28234 = n28233 ^ n28205 ^ n26032 ;
  assign n28235 = n3085 | n6149 ;
  assign n28236 = n26490 ^ n23452 ^ 1'b0 ;
  assign n28237 = n10381 | n12516 ;
  assign n28238 = n12387 & ~n28237 ;
  assign n28240 = n9077 ^ n2193 ^ 1'b0 ;
  assign n28241 = ~n1865 & n28240 ;
  assign n28239 = n18891 & ~n23590 ;
  assign n28242 = n28241 ^ n28239 ^ 1'b0 ;
  assign n28243 = n1111 & ~n28242 ;
  assign n28244 = n26820 ^ n19822 ^ n9493 ;
  assign n28245 = n24413 ^ n304 ^ 1'b0 ;
  assign n28246 = n28245 ^ n15531 ^ n7208 ;
  assign n28247 = n23856 ^ n8125 ^ 1'b0 ;
  assign n28248 = n13440 ^ n5131 ^ n985 ;
  assign n28249 = n28248 ^ n9635 ^ n1820 ;
  assign n28250 = n17276 & ~n28249 ;
  assign n28254 = n11014 ^ n2413 ^ 1'b0 ;
  assign n28255 = n8989 | n28254 ;
  assign n28252 = n8699 ^ n913 ^ 1'b0 ;
  assign n28251 = ( n2253 & ~n15411 ) | ( n2253 & n18614 ) | ( ~n15411 & n18614 ) ;
  assign n28253 = n28252 ^ n28251 ^ n2516 ;
  assign n28256 = n28255 ^ n28253 ^ n11632 ;
  assign n28257 = ( x104 & n14513 ) | ( x104 & n16136 ) | ( n14513 & n16136 ) ;
  assign n28258 = n26354 ^ n22884 ^ 1'b0 ;
  assign n28259 = ~n28257 & n28258 ;
  assign n28260 = ~n1265 & n12064 ;
  assign n28261 = n28260 ^ n19972 ^ 1'b0 ;
  assign n28266 = ~n5656 & n14766 ;
  assign n28267 = ( n8975 & n9020 ) | ( n8975 & ~n28266 ) | ( n9020 & ~n28266 ) ;
  assign n28262 = ~n2326 & n3433 ;
  assign n28263 = n8802 ^ n281 ^ 1'b0 ;
  assign n28264 = n9414 | n28263 ;
  assign n28265 = n28262 | n28264 ;
  assign n28268 = n28267 ^ n28265 ^ n16923 ;
  assign n28269 = n1594 & ~n23818 ;
  assign n28270 = n26289 ^ n13939 ^ n392 ;
  assign n28271 = n14602 ^ n11386 ^ n6407 ;
  assign n28273 = n12961 ^ n4916 ^ 1'b0 ;
  assign n28274 = n15647 | n28273 ;
  assign n28272 = ( n984 & n4409 ) | ( n984 & n8411 ) | ( n4409 & n8411 ) ;
  assign n28275 = n28274 ^ n28272 ^ n409 ;
  assign n28276 = ~n21964 & n28275 ;
  assign n28277 = n1063 | n15146 ;
  assign n28282 = n3467 & n13541 ;
  assign n28283 = n28282 ^ n18652 ^ 1'b0 ;
  assign n28278 = n16353 | n21399 ;
  assign n28279 = n21860 | n28278 ;
  assign n28280 = n26549 ^ n17857 ^ n6544 ;
  assign n28281 = ( n13349 & ~n28279 ) | ( n13349 & n28280 ) | ( ~n28279 & n28280 ) ;
  assign n28284 = n28283 ^ n28281 ^ n16274 ;
  assign n28285 = n4415 & ~n28284 ;
  assign n28286 = n28277 & n28285 ;
  assign n28287 = n24343 ^ n18487 ^ 1'b0 ;
  assign n28288 = n4301 | n28287 ;
  assign n28289 = n21143 ^ n17977 ^ n4233 ;
  assign n28290 = n27755 | n28289 ;
  assign n28291 = n23205 ^ n7858 ^ n5877 ;
  assign n28292 = n25545 ^ n23442 ^ n1709 ;
  assign n28293 = ( n3240 & n7981 ) | ( n3240 & ~n17763 ) | ( n7981 & ~n17763 ) ;
  assign n28294 = n28293 ^ n24922 ^ 1'b0 ;
  assign n28295 = n27018 ^ n15991 ^ n2484 ;
  assign n28296 = ~n2890 & n10920 ;
  assign n28297 = n2214 & n25372 ;
  assign n28298 = n3831 & n28297 ;
  assign n28299 = ( n9128 & ~n13083 ) | ( n9128 & n14005 ) | ( ~n13083 & n14005 ) ;
  assign n28300 = n27503 ^ n26926 ^ 1'b0 ;
  assign n28301 = ~n9728 & n11523 ;
  assign n28302 = n28301 ^ n26139 ^ n24669 ;
  assign n28303 = ( n15542 & ~n15889 ) | ( n15542 & n21591 ) | ( ~n15889 & n21591 ) ;
  assign n28304 = n28303 ^ n20672 ^ n10012 ;
  assign n28305 = n14233 ^ n6903 ^ n4342 ;
  assign n28306 = n2526 & ~n23000 ;
  assign n28307 = ~n9706 & n28306 ;
  assign n28308 = n28307 ^ n8450 ^ 1'b0 ;
  assign n28309 = n1828 & ~n12311 ;
  assign n28310 = n6338 | n27784 ;
  assign n28311 = ~n652 & n11262 ;
  assign n28312 = n28311 ^ n15871 ^ 1'b0 ;
  assign n28313 = n12401 ^ n4109 ^ 1'b0 ;
  assign n28314 = ~n4709 & n28313 ;
  assign n28315 = n28314 ^ n3917 ^ 1'b0 ;
  assign n28316 = ~n19393 & n28315 ;
  assign n28317 = n775 & ~n821 ;
  assign n28318 = n17077 ^ n7274 ^ n6984 ;
  assign n28319 = ~n1460 & n28318 ;
  assign n28320 = ( n21503 & ~n28317 ) | ( n21503 & n28319 ) | ( ~n28317 & n28319 ) ;
  assign n28321 = n11177 ^ n9607 ^ x13 ;
  assign n28322 = ( n2138 & ~n3976 ) | ( n2138 & n28321 ) | ( ~n3976 & n28321 ) ;
  assign n28323 = n17477 ^ n8842 ^ n939 ;
  assign n28324 = n8737 & ~n28323 ;
  assign n28325 = ( ~n1503 & n16216 ) | ( ~n1503 & n26918 ) | ( n16216 & n26918 ) ;
  assign n28326 = n8668 & ~n16680 ;
  assign n28327 = n28326 ^ n5530 ^ 1'b0 ;
  assign n28328 = n17610 ^ n5873 ^ 1'b0 ;
  assign n28329 = n28327 | n28328 ;
  assign n28330 = n1518 & ~n2298 ;
  assign n28331 = n16970 ^ n3802 ^ n1668 ;
  assign n28332 = ( n5710 & n17141 ) | ( n5710 & n24332 ) | ( n17141 & n24332 ) ;
  assign n28333 = ( n6182 & n15596 ) | ( n6182 & n23625 ) | ( n15596 & n23625 ) ;
  assign n28334 = n11064 ^ n5956 ^ n4106 ;
  assign n28335 = n14947 ^ n4689 ^ 1'b0 ;
  assign n28336 = n19147 ^ n16712 ^ 1'b0 ;
  assign n28337 = n23248 & n28336 ;
  assign n28338 = ~n6895 & n18927 ;
  assign n28339 = n28338 ^ n10577 ^ 1'b0 ;
  assign n28340 = n28241 ^ n20972 ^ 1'b0 ;
  assign n28341 = n20680 | n28340 ;
  assign n28342 = n28341 ^ n9712 ^ n1757 ;
  assign n28343 = n16704 ^ n8508 ^ n3631 ;
  assign n28344 = n13834 ^ n824 ^ 1'b0 ;
  assign n28345 = ( ~n24661 & n27737 ) | ( ~n24661 & n28344 ) | ( n27737 & n28344 ) ;
  assign n28346 = n14417 ^ n2090 ^ 1'b0 ;
  assign n28347 = n24739 | n28346 ;
  assign n28348 = n542 & n27943 ;
  assign n28349 = n28348 ^ n5658 ^ 1'b0 ;
  assign n28350 = ( ~n9363 & n20544 ) | ( ~n9363 & n28349 ) | ( n20544 & n28349 ) ;
  assign n28351 = n13294 ^ n9910 ^ n203 ;
  assign n28352 = n18437 | n28351 ;
  assign n28353 = n8219 & ~n9014 ;
  assign n28354 = n28353 ^ n6094 ^ 1'b0 ;
  assign n28355 = n27935 & n28354 ;
  assign n28356 = ~n133 & n28355 ;
  assign n28357 = ~n27570 & n28356 ;
  assign n28358 = ~n10279 & n18469 ;
  assign n28359 = n27930 ^ n27378 ^ 1'b0 ;
  assign n28360 = ~n5780 & n16175 ;
  assign n28361 = n16409 ^ n13628 ^ n4776 ;
  assign n28362 = ( n4567 & n22099 ) | ( n4567 & ~n27224 ) | ( n22099 & ~n27224 ) ;
  assign n28363 = ( ~n568 & n3436 ) | ( ~n568 & n10739 ) | ( n3436 & n10739 ) ;
  assign n28364 = ~n9751 & n28363 ;
  assign n28365 = n14484 ^ n4537 ^ 1'b0 ;
  assign n28366 = n10950 & n28365 ;
  assign n28367 = n28366 ^ n22840 ^ n12758 ;
  assign n28368 = n27012 ^ n16049 ^ n13523 ;
  assign n28369 = n24696 ^ n3595 ^ n1887 ;
  assign n28370 = n28369 ^ n4720 ^ 1'b0 ;
  assign n28371 = n1914 & ~n4210 ;
  assign n28372 = ~n15504 & n28371 ;
  assign n28373 = n3548 ^ n1736 ^ n705 ;
  assign n28374 = ( n8849 & n27887 ) | ( n8849 & n28373 ) | ( n27887 & n28373 ) ;
  assign n28375 = n28374 ^ n10261 ^ 1'b0 ;
  assign n28376 = n20500 | n28375 ;
  assign n28377 = n13973 & ~n22935 ;
  assign n28378 = n28377 ^ n21301 ^ 1'b0 ;
  assign n28379 = n16269 ^ n5320 ^ 1'b0 ;
  assign n28380 = n28379 ^ n10241 ^ n8477 ;
  assign n28381 = ( ~n995 & n3779 ) | ( ~n995 & n26697 ) | ( n3779 & n26697 ) ;
  assign n28382 = ( n4549 & n6613 ) | ( n4549 & ~n28381 ) | ( n6613 & ~n28381 ) ;
  assign n28383 = n16952 ^ n4161 ^ n844 ;
  assign n28384 = n10828 & ~n28383 ;
  assign n28385 = ( n2388 & n3846 ) | ( n2388 & ~n6450 ) | ( n3846 & ~n6450 ) ;
  assign n28386 = n11329 | n28385 ;
  assign n28387 = n14555 & ~n28386 ;
  assign n28388 = ( n2470 & n8066 ) | ( n2470 & n18255 ) | ( n8066 & n18255 ) ;
  assign n28389 = ( ~n11065 & n20386 ) | ( ~n11065 & n28388 ) | ( n20386 & n28388 ) ;
  assign n28390 = n4983 ^ n4581 ^ 1'b0 ;
  assign n28391 = n5167 | n26719 ;
  assign n28392 = ( n9138 & ~n20067 ) | ( n9138 & n20681 ) | ( ~n20067 & n20681 ) ;
  assign n28393 = ( ~n16999 & n23694 ) | ( ~n16999 & n28392 ) | ( n23694 & n28392 ) ;
  assign n28394 = n18869 ^ n16679 ^ n2053 ;
  assign n28395 = n28394 ^ n26694 ^ 1'b0 ;
  assign n28396 = ( n14344 & n28015 ) | ( n14344 & ~n28395 ) | ( n28015 & ~n28395 ) ;
  assign n28397 = n27003 ^ n18818 ^ n433 ;
  assign n28398 = n2153 & ~n19702 ;
  assign n28399 = n4585 | n28398 ;
  assign n28400 = n16347 & n23360 ;
  assign n28401 = n8126 & n28400 ;
  assign n28402 = n18900 ^ n13711 ^ n5401 ;
  assign n28403 = n28402 ^ n27858 ^ 1'b0 ;
  assign n28404 = ~n884 & n28403 ;
  assign n28405 = n18461 ^ n6060 ^ n2807 ;
  assign n28406 = n16750 | n25294 ;
  assign n28407 = n3486 ^ n1909 ^ 1'b0 ;
  assign n28408 = ( ~n1257 & n23280 ) | ( ~n1257 & n28407 ) | ( n23280 & n28407 ) ;
  assign n28409 = n24113 ^ n16126 ^ 1'b0 ;
  assign n28412 = n4639 & ~n8140 ;
  assign n28410 = n3254 ^ n250 ^ 1'b0 ;
  assign n28411 = n28410 ^ n10225 ^ n6751 ;
  assign n28413 = n28412 ^ n28411 ^ n20270 ;
  assign n28414 = n28409 & n28413 ;
  assign n28415 = n16406 ^ n5216 ^ 1'b0 ;
  assign n28416 = n28415 ^ n20438 ^ n7277 ;
  assign n28417 = n11613 & n12992 ;
  assign n28418 = ~n3389 & n28417 ;
  assign n28419 = n13108 ^ n2848 ^ 1'b0 ;
  assign n28420 = n8930 & ~n28419 ;
  assign n28421 = n28420 ^ n9657 ^ 1'b0 ;
  assign n28422 = ~n21324 & n23808 ;
  assign n28423 = ( ~n11023 & n19424 ) | ( ~n11023 & n26957 ) | ( n19424 & n26957 ) ;
  assign n28424 = n21510 ^ n13978 ^ n7943 ;
  assign n28425 = n16864 ^ n12822 ^ n1516 ;
  assign n28428 = n6290 & ~n7108 ;
  assign n28429 = n6388 & n28428 ;
  assign n28426 = n17103 | n24522 ;
  assign n28427 = n8687 & ~n28426 ;
  assign n28430 = n28429 ^ n28427 ^ n22271 ;
  assign n28431 = n20482 ^ n17505 ^ n1691 ;
  assign n28432 = ( n11247 & ~n12909 ) | ( n11247 & n28431 ) | ( ~n12909 & n28431 ) ;
  assign n28433 = n7836 & ~n16077 ;
  assign n28434 = ( n13267 & n15648 ) | ( n13267 & n28433 ) | ( n15648 & n28433 ) ;
  assign n28435 = n3131 ^ n2757 ^ 1'b0 ;
  assign n28436 = n20040 & ~n28435 ;
  assign n28438 = n24473 ^ n2377 ^ n273 ;
  assign n28437 = n12339 & ~n16581 ;
  assign n28439 = n28438 ^ n28437 ^ 1'b0 ;
  assign n28440 = n1863 | n3476 ;
  assign n28441 = n21040 ^ n19256 ^ 1'b0 ;
  assign n28442 = n25367 | n28441 ;
  assign n28443 = n16777 ^ n8253 ^ n2812 ;
  assign n28444 = n25491 ^ n20790 ^ n4409 ;
  assign n28445 = n22816 & ~n27433 ;
  assign n28446 = n14425 ^ n2229 ^ n1441 ;
  assign n28447 = n28446 ^ n23369 ^ n22146 ;
  assign n28449 = ( n512 & n3382 ) | ( n512 & n3709 ) | ( n3382 & n3709 ) ;
  assign n28448 = n8664 & ~n13844 ;
  assign n28450 = n28449 ^ n28448 ^ n18747 ;
  assign n28451 = ( n6108 & n10742 ) | ( n6108 & n24140 ) | ( n10742 & n24140 ) ;
  assign n28452 = n4541 & ~n10494 ;
  assign n28453 = ~n27283 & n28452 ;
  assign n28454 = n2524 & ~n11361 ;
  assign n28455 = n28454 ^ n24525 ^ 1'b0 ;
  assign n28460 = ( n345 & ~n1265 ) | ( n345 & n10221 ) | ( ~n1265 & n10221 ) ;
  assign n28456 = ~n4301 & n8771 ;
  assign n28457 = ~n2935 & n28456 ;
  assign n28458 = n15506 & n28457 ;
  assign n28459 = n12569 & ~n28458 ;
  assign n28461 = n28460 ^ n28459 ^ 1'b0 ;
  assign n28462 = n14504 ^ n5138 ^ n4121 ;
  assign n28463 = n16914 | n18252 ;
  assign n28464 = n9722 & ~n28463 ;
  assign n28465 = n28464 ^ n10658 ^ n4195 ;
  assign n28466 = n8882 & n11889 ;
  assign n28467 = ( ~n1129 & n7654 ) | ( ~n1129 & n18021 ) | ( n7654 & n18021 ) ;
  assign n28468 = n17069 ^ n16928 ^ n16006 ;
  assign n28469 = n17941 ^ n15499 ^ n3200 ;
  assign n28470 = n26214 ^ x60 ^ 1'b0 ;
  assign n28471 = n14093 | n28470 ;
  assign n28472 = n14454 ^ n2964 ^ 1'b0 ;
  assign n28473 = ~n13237 & n26209 ;
  assign n28474 = n28472 & n28473 ;
  assign n28475 = n2401 | n9738 ;
  assign n28476 = n10528 | n28475 ;
  assign n28477 = ~n21177 & n28476 ;
  assign n28478 = n28477 ^ n24873 ^ 1'b0 ;
  assign n28479 = ~n24742 & n27307 ;
  assign n28480 = n28479 ^ n6083 ^ 1'b0 ;
  assign n28481 = n5371 | n24648 ;
  assign n28482 = n16628 & ~n28481 ;
  assign n28483 = n11536 & ~n28482 ;
  assign n28484 = ( n825 & n20022 ) | ( n825 & ~n22426 ) | ( n20022 & ~n22426 ) ;
  assign n28485 = n21793 ^ n16802 ^ n11609 ;
  assign n28486 = n22092 ^ n5665 ^ 1'b0 ;
  assign n28487 = n28485 & n28486 ;
  assign n28488 = n15411 ^ n11447 ^ n7523 ;
  assign n28489 = ( n1609 & n2355 ) | ( n1609 & ~n3998 ) | ( n2355 & ~n3998 ) ;
  assign n28490 = n12412 ^ n12109 ^ n760 ;
  assign n28491 = n28490 ^ n10404 ^ 1'b0 ;
  assign n28492 = n28491 ^ n16261 ^ n9650 ;
  assign n28494 = ( n1419 & n2916 ) | ( n1419 & n8130 ) | ( n2916 & n8130 ) ;
  assign n28493 = ~n4404 & n10219 ;
  assign n28495 = n28494 ^ n28493 ^ 1'b0 ;
  assign n28496 = ~n8171 & n18593 ;
  assign n28497 = n28496 ^ n8153 ^ 1'b0 ;
  assign n28498 = n24302 ^ n23734 ^ 1'b0 ;
  assign n28499 = n28497 & n28498 ;
  assign n28500 = n6375 & ~n23165 ;
  assign n28501 = ~n6792 & n28500 ;
  assign n28502 = ~n5809 & n15930 ;
  assign n28504 = n4920 ^ n4638 ^ 1'b0 ;
  assign n28503 = n17835 ^ n5327 ^ 1'b0 ;
  assign n28505 = n28504 ^ n28503 ^ n26537 ;
  assign n28506 = ~n7635 & n11350 ;
  assign n28507 = n28506 ^ n28022 ^ n22907 ;
  assign n28508 = n22803 ^ n15444 ^ 1'b0 ;
  assign n28509 = n28482 ^ n25209 ^ n7523 ;
  assign n28510 = ( n9454 & n9790 ) | ( n9454 & n14794 ) | ( n9790 & n14794 ) ;
  assign n28511 = n14843 & ~n28510 ;
  assign n28512 = n28511 ^ n22247 ^ 1'b0 ;
  assign n28513 = n28512 ^ n13536 ^ n10309 ;
  assign n28514 = ~n13307 & n28082 ;
  assign n28520 = n15483 ^ n6025 ^ 1'b0 ;
  assign n28521 = ~n4793 & n28520 ;
  assign n28518 = n27117 ^ n8781 ^ n2021 ;
  assign n28517 = n27145 ^ n15757 ^ 1'b0 ;
  assign n28515 = ~n10029 & n13697 ;
  assign n28516 = ~n1629 & n28515 ;
  assign n28519 = n28518 ^ n28517 ^ n28516 ;
  assign n28522 = n28521 ^ n28519 ^ 1'b0 ;
  assign n28523 = n7087 & n28522 ;
  assign n28524 = ~n21734 & n28523 ;
  assign n28525 = ~n8298 & n8378 ;
  assign n28526 = n13750 ^ n8970 ^ 1'b0 ;
  assign n28527 = n28525 | n28526 ;
  assign n28528 = n12059 ^ n11389 ^ n6601 ;
  assign n28529 = n28528 ^ n27304 ^ n1059 ;
  assign n28530 = n10723 ^ n9580 ^ n6913 ;
  assign n28531 = ( n479 & n11487 ) | ( n479 & n26674 ) | ( n11487 & n26674 ) ;
  assign n28532 = n11194 ^ n7024 ^ 1'b0 ;
  assign n28533 = n14418 & ~n28532 ;
  assign n28534 = ( n18769 & n26872 ) | ( n18769 & ~n28533 ) | ( n26872 & ~n28533 ) ;
  assign n28535 = n18787 ^ n17943 ^ n825 ;
  assign n28536 = n16534 & ~n28535 ;
  assign n28537 = n6313 ^ n272 ^ n169 ;
  assign n28538 = n3429 & ~n28537 ;
  assign n28539 = n26983 ^ n14406 ^ 1'b0 ;
  assign n28540 = n28539 ^ n1023 ^ 1'b0 ;
  assign n28541 = ( ~n2638 & n3614 ) | ( ~n2638 & n25769 ) | ( n3614 & n25769 ) ;
  assign n28542 = ~n8964 & n22869 ;
  assign n28543 = n137 & n15024 ;
  assign n28544 = n28543 ^ n2431 ^ 1'b0 ;
  assign n28545 = n28544 ^ n5286 ^ 1'b0 ;
  assign n28546 = n17676 ^ n10835 ^ n9034 ;
  assign n28547 = ~n11222 & n19892 ;
  assign n28548 = n28547 ^ n28107 ^ 1'b0 ;
  assign n28549 = n757 | n18432 ;
  assign n28550 = n28549 ^ n3958 ^ 1'b0 ;
  assign n28551 = n28550 ^ n22076 ^ 1'b0 ;
  assign n28552 = n377 | n1971 ;
  assign n28553 = n22616 & ~n28552 ;
  assign n28554 = n28553 ^ n8752 ^ 1'b0 ;
  assign n28555 = n17895 & n28554 ;
  assign n28556 = n12711 ^ n6219 ^ n1444 ;
  assign n28557 = ~n5118 & n28556 ;
  assign n28558 = ~n28555 & n28557 ;
  assign n28559 = ~n6110 & n19444 ;
  assign n28560 = n12582 ^ n9515 ^ 1'b0 ;
  assign n28561 = n11421 ^ n2636 ^ n2632 ;
  assign n28562 = n691 & n28561 ;
  assign n28563 = n28562 ^ n14596 ^ n680 ;
  assign n28564 = n16069 ^ n9469 ^ 1'b0 ;
  assign n28565 = ( ~n12129 & n22210 ) | ( ~n12129 & n25690 ) | ( n22210 & n25690 ) ;
  assign n28566 = ~n842 & n1308 ;
  assign n28567 = ( ~n8258 & n28565 ) | ( ~n8258 & n28566 ) | ( n28565 & n28566 ) ;
  assign n28568 = n28567 ^ n1408 ^ x30 ;
  assign n28569 = n28568 ^ n26681 ^ 1'b0 ;
  assign n28570 = n2096 ^ n1784 ^ 1'b0 ;
  assign n28571 = n15066 & ~n28570 ;
  assign n28572 = n28571 ^ n4587 ^ n1587 ;
  assign n28573 = n9087 ^ n4896 ^ n1804 ;
  assign n28574 = n9028 & n10772 ;
  assign n28575 = ( ~n18219 & n21525 ) | ( ~n18219 & n28574 ) | ( n21525 & n28574 ) ;
  assign n28576 = n28575 ^ n14682 ^ 1'b0 ;
  assign n28577 = ~n4990 & n28136 ;
  assign n28578 = n16221 & n28577 ;
  assign n28579 = n3612 & ~n15576 ;
  assign n28580 = n28579 ^ n18500 ^ 1'b0 ;
  assign n28581 = n28580 ^ n19485 ^ 1'b0 ;
  assign n28582 = n2277 & ~n3107 ;
  assign n28583 = n11419 & n28582 ;
  assign n28584 = n1044 & ~n23127 ;
  assign n28585 = n28584 ^ n5045 ^ 1'b0 ;
  assign n28587 = n16049 ^ n14421 ^ n5346 ;
  assign n28586 = ~n360 & n14170 ;
  assign n28588 = n28587 ^ n28586 ^ 1'b0 ;
  assign n28589 = n24357 ^ n18981 ^ n18302 ;
  assign n28590 = ( n2402 & n13532 ) | ( n2402 & n24376 ) | ( n13532 & n24376 ) ;
  assign n28591 = ( n5648 & n7782 ) | ( n5648 & ~n18565 ) | ( n7782 & ~n18565 ) ;
  assign n28592 = ( n4139 & n9383 ) | ( n4139 & ~n28591 ) | ( n9383 & ~n28591 ) ;
  assign n28593 = ( n10084 & n13622 ) | ( n10084 & n21911 ) | ( n13622 & n21911 ) ;
  assign n28594 = ( ~n7210 & n21744 ) | ( ~n7210 & n28593 ) | ( n21744 & n28593 ) ;
  assign n28595 = n2510 | n21712 ;
  assign n28596 = n20526 | n28595 ;
  assign n28597 = ( n6636 & ~n16148 ) | ( n6636 & n28596 ) | ( ~n16148 & n28596 ) ;
  assign n28598 = ( n3419 & n5081 ) | ( n3419 & ~n26582 ) | ( n5081 & ~n26582 ) ;
  assign n28600 = ( n5145 & n9260 ) | ( n5145 & n18842 ) | ( n9260 & n18842 ) ;
  assign n28599 = n3186 & ~n8970 ;
  assign n28601 = n28600 ^ n28599 ^ 1'b0 ;
  assign n28602 = n1700 & n14455 ;
  assign n28603 = n28602 ^ n7843 ^ 1'b0 ;
  assign n28604 = n24322 ^ n1872 ^ 1'b0 ;
  assign n28605 = n17978 ^ n10684 ^ 1'b0 ;
  assign n28606 = ~n28604 & n28605 ;
  assign n28607 = ~n3511 & n12334 ;
  assign n28608 = ~n6509 & n28607 ;
  assign n28609 = n28608 ^ n20292 ^ n11242 ;
  assign n28610 = n13746 ^ n7848 ^ 1'b0 ;
  assign n28611 = n12359 ^ n441 ^ 1'b0 ;
  assign n28612 = n12970 ^ n8314 ^ 1'b0 ;
  assign n28613 = ( n9317 & n9883 ) | ( n9317 & n28612 ) | ( n9883 & n28612 ) ;
  assign n28614 = n23793 ^ n3575 ^ n794 ;
  assign n28615 = n28614 ^ n23329 ^ n16803 ;
  assign n28616 = n2609 ^ x118 ^ 1'b0 ;
  assign n28617 = n11213 & n28616 ;
  assign n28618 = ~n729 & n28617 ;
  assign n28619 = n28618 ^ n13479 ^ n2227 ;
  assign n28620 = n19044 ^ n11597 ^ 1'b0 ;
  assign n28621 = n25665 ^ n23921 ^ 1'b0 ;
  assign n28622 = n28620 & ~n28621 ;
  assign n28623 = n14966 ^ n3909 ^ 1'b0 ;
  assign n28624 = n7713 & n28623 ;
  assign n28625 = n28624 ^ n4678 ^ 1'b0 ;
  assign n28626 = n23236 ^ n21105 ^ n8728 ;
  assign n28627 = n19702 ^ n18298 ^ n14021 ;
  assign n28628 = n26239 ^ n7082 ^ x120 ;
  assign n28629 = n27770 ^ n11785 ^ n9632 ;
  assign n28630 = n12316 | n28629 ;
  assign n28631 = ~n23296 & n25507 ;
  assign n28632 = n20348 ^ n13013 ^ n4224 ;
  assign n28633 = n9086 & ~n19708 ;
  assign n28634 = n18639 ^ n12315 ^ n4138 ;
  assign n28635 = n7953 & n17929 ;
  assign n28636 = n28634 & n28635 ;
  assign n28637 = n27877 ^ n22037 ^ n20321 ;
  assign n28638 = n12771 ^ n11994 ^ 1'b0 ;
  assign n28639 = n21752 ^ n17094 ^ n8980 ;
  assign n28640 = n10095 ^ n3474 ^ 1'b0 ;
  assign n28641 = ~n14183 & n28640 ;
  assign n28642 = ( n11758 & n20609 ) | ( n11758 & n28641 ) | ( n20609 & n28641 ) ;
  assign n28643 = n16224 ^ n826 ^ 1'b0 ;
  assign n28644 = n3447 | n28643 ;
  assign n28645 = n28644 ^ n16008 ^ 1'b0 ;
  assign n28646 = ( n1084 & n28205 ) | ( n1084 & ~n28645 ) | ( n28205 & ~n28645 ) ;
  assign n28647 = n21864 ^ n13573 ^ n5747 ;
  assign n28648 = ( n12498 & n19242 ) | ( n12498 & ~n22552 ) | ( n19242 & ~n22552 ) ;
  assign n28649 = n8344 | n21399 ;
  assign n28650 = n28648 & ~n28649 ;
  assign n28651 = n3666 & n16440 ;
  assign n28652 = n28651 ^ n27019 ^ 1'b0 ;
  assign n28653 = n12367 ^ n1952 ^ 1'b0 ;
  assign n28654 = ( n2579 & ~n18546 ) | ( n2579 & n28653 ) | ( ~n18546 & n28653 ) ;
  assign n28655 = n11811 ^ n4510 ^ n2128 ;
  assign n28656 = ( n8420 & ~n14249 ) | ( n8420 & n26237 ) | ( ~n14249 & n26237 ) ;
  assign n28657 = n3810 & n15613 ;
  assign n28658 = ( ~n1543 & n21651 ) | ( ~n1543 & n22049 ) | ( n21651 & n22049 ) ;
  assign n28659 = n28658 ^ n15483 ^ n8629 ;
  assign n28660 = n28659 ^ n20316 ^ n18924 ;
  assign n28662 = ( n9144 & n21749 ) | ( n9144 & ~n24587 ) | ( n21749 & ~n24587 ) ;
  assign n28663 = n28662 ^ n10729 ^ n8701 ;
  assign n28661 = n2070 | n3255 ;
  assign n28664 = n28663 ^ n28661 ^ 1'b0 ;
  assign n28665 = n22515 | n28664 ;
  assign n28666 = n4535 & ~n28665 ;
  assign n28667 = n18423 ^ n15561 ^ 1'b0 ;
  assign n28668 = n9594 | n28667 ;
  assign n28669 = ( n7588 & n18064 ) | ( n7588 & ~n23690 ) | ( n18064 & ~n23690 ) ;
  assign n28675 = n5715 ^ n3225 ^ 1'b0 ;
  assign n28674 = n8225 ^ n7939 ^ n3408 ;
  assign n28670 = n13360 ^ n11341 ^ n3837 ;
  assign n28671 = n28670 ^ n19768 ^ n2695 ;
  assign n28672 = ( n11221 & n11932 ) | ( n11221 & n28671 ) | ( n11932 & n28671 ) ;
  assign n28673 = n28672 ^ n13854 ^ n10750 ;
  assign n28676 = n28675 ^ n28674 ^ n28673 ;
  assign n28677 = n8462 & ~n13032 ;
  assign n28678 = n10291 & n28677 ;
  assign n28679 = ( ~n8592 & n18052 ) | ( ~n8592 & n28678 ) | ( n18052 & n28678 ) ;
  assign n28680 = n28679 ^ n6397 ^ n5066 ;
  assign n28681 = n28680 ^ n21474 ^ n18618 ;
  assign n28682 = ~n4906 & n8059 ;
  assign n28683 = n28682 ^ n2459 ^ 1'b0 ;
  assign n28684 = ~n3924 & n21773 ;
  assign n28685 = n28683 & n28684 ;
  assign n28686 = n12931 & n28685 ;
  assign n28687 = n5647 & n5955 ;
  assign n28688 = n1157 | n13334 ;
  assign n28689 = n21094 & ~n28688 ;
  assign n28690 = ( n12256 & n18835 ) | ( n12256 & ~n28689 ) | ( n18835 & ~n28689 ) ;
  assign n28691 = x58 & n23988 ;
  assign n28692 = n9473 ^ n7085 ^ 1'b0 ;
  assign n28693 = n1624 | n28692 ;
  assign n28694 = ~n3076 & n16702 ;
  assign n28695 = n28693 & n28694 ;
  assign n28696 = ~n1439 & n17508 ;
  assign n28697 = ~n12868 & n28696 ;
  assign n28698 = ~n23609 & n28697 ;
  assign n28699 = n9666 ^ n5292 ^ 1'b0 ;
  assign n28700 = n9992 & n15024 ;
  assign n28701 = n28700 ^ n9323 ^ 1'b0 ;
  assign n28702 = n28701 ^ n25808 ^ 1'b0 ;
  assign n28703 = ( n1646 & n7736 ) | ( n1646 & n20952 ) | ( n7736 & n20952 ) ;
  assign n28704 = n28703 ^ n18707 ^ n16231 ;
  assign n28705 = n28704 ^ n21274 ^ n10608 ;
  assign n28706 = n6620 ^ n1018 ^ 1'b0 ;
  assign n28707 = n11239 ^ n2481 ^ 1'b0 ;
  assign n28708 = ~n13723 & n23758 ;
  assign n28709 = ~n18645 & n28708 ;
  assign n28710 = ( n2471 & n28707 ) | ( n2471 & n28709 ) | ( n28707 & n28709 ) ;
  assign n28711 = n24429 ^ n22271 ^ 1'b0 ;
  assign n28712 = n28711 ^ n24151 ^ n21920 ;
  assign n28713 = ( ~n5647 & n12038 ) | ( ~n5647 & n13321 ) | ( n12038 & n13321 ) ;
  assign n28714 = n28713 ^ n15003 ^ n3398 ;
  assign n28715 = n9384 & n11646 ;
  assign n28716 = n471 | n28715 ;
  assign n28717 = n27835 & ~n28716 ;
  assign n28718 = n28714 | n28717 ;
  assign n28719 = n28718 ^ n1601 ^ 1'b0 ;
  assign n28720 = ~n6106 & n14214 ;
  assign n28721 = ~n1634 & n28720 ;
  assign n28722 = n28721 ^ n1507 ^ 1'b0 ;
  assign n28723 = n2205 & ~n25879 ;
  assign n28724 = ~n20354 & n28723 ;
  assign n28725 = n13986 ^ n1340 ^ 1'b0 ;
  assign n28726 = n28724 | n28725 ;
  assign n28727 = n28216 ^ n23229 ^ 1'b0 ;
  assign n28728 = n11275 & n28727 ;
  assign n28730 = n22679 ^ n13404 ^ n9420 ;
  assign n28731 = n2493 & ~n19564 ;
  assign n28732 = n28730 & n28731 ;
  assign n28729 = n1957 | n13125 ;
  assign n28733 = n28732 ^ n28729 ^ 1'b0 ;
  assign n28734 = n28733 ^ n12634 ^ n10230 ;
  assign n28735 = n4129 & ~n4638 ;
  assign n28736 = n28735 ^ n7585 ^ 1'b0 ;
  assign n28737 = n28736 ^ n24475 ^ n19346 ;
  assign n28738 = n8067 ^ n376 ^ 1'b0 ;
  assign n28739 = n7278 ^ n5382 ^ n3540 ;
  assign n28740 = n7874 & ~n9534 ;
  assign n28741 = n20937 ^ n5792 ^ 1'b0 ;
  assign n28742 = n28741 ^ n22576 ^ 1'b0 ;
  assign n28743 = n9658 | n27582 ;
  assign n28744 = ~n9384 & n28743 ;
  assign n28745 = n17365 & n28744 ;
  assign n28746 = n17565 ^ n7121 ^ 1'b0 ;
  assign n28747 = ~n28745 & n28746 ;
  assign n28748 = n9695 | n27930 ;
  assign n28749 = ( n1119 & n6770 ) | ( n1119 & n12407 ) | ( n6770 & n12407 ) ;
  assign n28750 = ( ~x96 & n15546 ) | ( ~x96 & n20810 ) | ( n15546 & n20810 ) ;
  assign n28751 = n2185 & ~n15222 ;
  assign n28752 = n28751 ^ n2770 ^ 1'b0 ;
  assign n28753 = n8154 & n22617 ;
  assign n28754 = n28753 ^ n9682 ^ 1'b0 ;
  assign n28755 = ~n17269 & n17314 ;
  assign n28756 = n15593 & n28755 ;
  assign n28757 = n18950 & ~n23127 ;
  assign n28758 = ~n1348 & n28757 ;
  assign n28759 = n637 | n5554 ;
  assign n28760 = n28759 ^ n10845 ^ 1'b0 ;
  assign n28761 = n7278 ^ n390 ^ 1'b0 ;
  assign n28762 = n12203 | n28761 ;
  assign n28763 = n28762 ^ n22709 ^ 1'b0 ;
  assign n28764 = ( n2298 & n3104 ) | ( n2298 & n3322 ) | ( n3104 & n3322 ) ;
  assign n28765 = n25496 ^ n21718 ^ n16054 ;
  assign n28766 = n21020 ^ n10682 ^ n5824 ;
  assign n28767 = n808 & n6198 ;
  assign n28768 = n19115 ^ n1452 ^ 1'b0 ;
  assign n28769 = ~n28767 & n28768 ;
  assign n28770 = n28769 ^ n4556 ^ 1'b0 ;
  assign n28771 = n21982 ^ n5561 ^ 1'b0 ;
  assign n28772 = n588 & ~n28771 ;
  assign n28773 = n7548 & n28772 ;
  assign n28774 = n4652 & ~n22441 ;
  assign n28775 = n12235 ^ n8776 ^ n3278 ;
  assign n28776 = n28775 ^ n24501 ^ n3679 ;
  assign n28777 = n10629 ^ n9559 ^ 1'b0 ;
  assign n28778 = n27488 | n28777 ;
  assign n28779 = n28778 ^ n24124 ^ n1288 ;
  assign n28780 = n28319 ^ n16298 ^ n2150 ;
  assign n28781 = n16165 ^ n11564 ^ n10759 ;
  assign n28782 = n28781 ^ n22033 ^ n19334 ;
  assign n28783 = n11932 | n12476 ;
  assign n28784 = n28783 ^ n27452 ^ n21399 ;
  assign n28785 = ( n3037 & ~n8658 ) | ( n3037 & n14690 ) | ( ~n8658 & n14690 ) ;
  assign n28786 = n27782 ^ n15420 ^ 1'b0 ;
  assign n28787 = n3976 & n9378 ;
  assign n28788 = ~n9697 & n28787 ;
  assign n28789 = n3014 & ~n14076 ;
  assign n28790 = n133 & n28789 ;
  assign n28791 = n24546 & ~n28790 ;
  assign n28792 = n28788 & n28791 ;
  assign n28793 = n16347 ^ n13597 ^ 1'b0 ;
  assign n28794 = n3739 | n28793 ;
  assign n28795 = n15023 | n28794 ;
  assign n28796 = ( ~n6947 & n20233 ) | ( ~n6947 & n28795 ) | ( n20233 & n28795 ) ;
  assign n28797 = n12067 ^ n5724 ^ 1'b0 ;
  assign n28798 = n28797 ^ n17089 ^ n184 ;
  assign n28799 = n7789 & n16074 ;
  assign n28800 = n28799 ^ n3117 ^ 1'b0 ;
  assign n28801 = n2633 & n12586 ;
  assign n28802 = n28800 & n28801 ;
  assign n28803 = n28802 ^ n28680 ^ n3835 ;
  assign n28804 = n15022 ^ n1831 ^ 1'b0 ;
  assign n28805 = ( n536 & n8630 ) | ( n536 & ~n28804 ) | ( n8630 & ~n28804 ) ;
  assign n28806 = n28805 ^ n12339 ^ n9338 ;
  assign n28807 = ( ~n13744 & n22806 ) | ( ~n13744 & n28806 ) | ( n22806 & n28806 ) ;
  assign n28808 = ~n550 & n24956 ;
  assign n28809 = ( n1248 & n3755 ) | ( n1248 & n20283 ) | ( n3755 & n20283 ) ;
  assign n28811 = ( n3975 & ~n5629 ) | ( n3975 & n11930 ) | ( ~n5629 & n11930 ) ;
  assign n28810 = n3967 & n12885 ;
  assign n28812 = n28811 ^ n28810 ^ 1'b0 ;
  assign n28813 = n875 | n7758 ;
  assign n28814 = n6104 | n28813 ;
  assign n28816 = ( n2524 & n8788 ) | ( n2524 & n9092 ) | ( n8788 & n9092 ) ;
  assign n28817 = n28816 ^ n21410 ^ 1'b0 ;
  assign n28815 = n2770 | n8756 ;
  assign n28818 = n28817 ^ n28815 ^ 1'b0 ;
  assign n28822 = n2950 & n17384 ;
  assign n28819 = ( n10227 & n16740 ) | ( n10227 & ~n28340 ) | ( n16740 & ~n28340 ) ;
  assign n28820 = n28819 ^ n8448 ^ n1431 ;
  assign n28821 = n2255 & ~n28820 ;
  assign n28823 = n28822 ^ n28821 ^ 1'b0 ;
  assign n28824 = ( n1501 & n6038 ) | ( n1501 & n7232 ) | ( n6038 & n7232 ) ;
  assign n28825 = ~n6864 & n24198 ;
  assign n28826 = n421 & ~n8064 ;
  assign n28827 = ~n16344 & n28826 ;
  assign n28828 = ( n28824 & n28825 ) | ( n28824 & n28827 ) | ( n28825 & n28827 ) ;
  assign n28829 = ( n13598 & ~n22009 ) | ( n13598 & n24982 ) | ( ~n22009 & n24982 ) ;
  assign n28830 = n19836 ^ n7049 ^ 1'b0 ;
  assign n28831 = ( ~n1727 & n19334 ) | ( ~n1727 & n28830 ) | ( n19334 & n28830 ) ;
  assign n28832 = n28831 ^ n26344 ^ n15952 ;
  assign n28833 = ~n7655 & n28832 ;
  assign n28834 = ~n5859 & n22412 ;
  assign n28835 = ( n23486 & n28767 ) | ( n23486 & ~n28834 ) | ( n28767 & ~n28834 ) ;
  assign n28836 = n12626 ^ n9500 ^ 1'b0 ;
  assign n28837 = n5216 & ~n28836 ;
  assign n28838 = n28837 ^ n19791 ^ n9490 ;
  assign n28839 = ~n5152 & n17266 ;
  assign n28840 = ~n6833 & n28839 ;
  assign n28841 = ( ~n4456 & n12502 ) | ( ~n4456 & n28840 ) | ( n12502 & n28840 ) ;
  assign n28842 = n11493 | n28841 ;
  assign n28843 = ( n662 & ~n11821 ) | ( n662 & n20496 ) | ( ~n11821 & n20496 ) ;
  assign n28844 = n3840 & n28843 ;
  assign n28846 = ( n3082 & n10709 ) | ( n3082 & ~n28083 ) | ( n10709 & ~n28083 ) ;
  assign n28845 = n5268 | n23661 ;
  assign n28847 = n28846 ^ n28845 ^ 1'b0 ;
  assign n28848 = n13741 ^ n8783 ^ n8004 ;
  assign n28849 = n28848 ^ n27020 ^ 1'b0 ;
  assign n28850 = ~n22192 & n28849 ;
  assign n28851 = n28850 ^ n9370 ^ 1'b0 ;
  assign n28852 = n2950 | n18610 ;
  assign n28853 = n28852 ^ n18561 ^ 1'b0 ;
  assign n28854 = n136 & n12145 ;
  assign n28855 = ~n9001 & n11604 ;
  assign n28856 = n11818 ^ n11659 ^ n10253 ;
  assign n28857 = n28856 ^ n13718 ^ n11035 ;
  assign n28858 = n28857 ^ n4919 ^ 1'b0 ;
  assign n28859 = n28858 ^ n17308 ^ 1'b0 ;
  assign n28860 = ( n5969 & n6290 ) | ( n5969 & ~n20408 ) | ( n6290 & ~n20408 ) ;
  assign n28861 = n19346 ^ n4102 ^ 1'b0 ;
  assign n28862 = n26890 ^ n21728 ^ 1'b0 ;
  assign n28863 = n292 & ~n28862 ;
  assign n28864 = ~n3699 & n13009 ;
  assign n28865 = n28864 ^ n20061 ^ 1'b0 ;
  assign n28866 = n2056 & n27304 ;
  assign n28867 = n28866 ^ n1049 ^ 1'b0 ;
  assign n28868 = n13657 ^ n4632 ^ 1'b0 ;
  assign n28869 = ~n28867 & n28868 ;
  assign n28870 = n19124 | n28869 ;
  assign n28871 = ( n323 & n6603 ) | ( n323 & ~n22126 ) | ( n6603 & ~n22126 ) ;
  assign n28872 = n20942 ^ n13412 ^ n965 ;
  assign n28873 = n28872 ^ n11930 ^ n1260 ;
  assign n28874 = n25271 ^ n22401 ^ n19920 ;
  assign n28875 = ( n1471 & ~n3560 ) | ( n1471 & n13314 ) | ( ~n3560 & n13314 ) ;
  assign n28876 = n20400 ^ n9435 ^ 1'b0 ;
  assign n28877 = n8690 ^ n8388 ^ 1'b0 ;
  assign n28878 = ~n4484 & n16285 ;
  assign n28879 = n21496 & n28878 ;
  assign n28880 = n21558 ^ n11044 ^ 1'b0 ;
  assign n28881 = ~n11300 & n28880 ;
  assign n28882 = n16661 ^ n8817 ^ 1'b0 ;
  assign n28883 = ~n25761 & n28882 ;
  assign n28884 = ~n3736 & n28883 ;
  assign n28885 = n28884 ^ n21422 ^ 1'b0 ;
  assign n28886 = ( n1817 & ~n7743 ) | ( n1817 & n20883 ) | ( ~n7743 & n20883 ) ;
  assign n28887 = n28886 ^ n25299 ^ 1'b0 ;
  assign n28888 = n28887 ^ n10896 ^ x70 ;
  assign n28889 = ( n293 & n13366 ) | ( n293 & n15578 ) | ( n13366 & n15578 ) ;
  assign n28890 = n24719 ^ n23413 ^ n7793 ;
  assign n28891 = ( n18989 & n28889 ) | ( n18989 & n28890 ) | ( n28889 & n28890 ) ;
  assign n28892 = n17314 | n22065 ;
  assign n28893 = n28892 ^ n26161 ^ n4508 ;
  assign n28894 = n8752 ^ n4521 ^ 1'b0 ;
  assign n28895 = n14895 ^ n8035 ^ n7661 ;
  assign n28896 = ( ~n13747 & n15043 ) | ( ~n13747 & n15504 ) | ( n15043 & n15504 ) ;
  assign n28897 = ( n11864 & ~n28895 ) | ( n11864 & n28896 ) | ( ~n28895 & n28896 ) ;
  assign n28898 = ( n6954 & n8292 ) | ( n6954 & n20115 ) | ( n8292 & n20115 ) ;
  assign n28899 = n12878 & n26214 ;
  assign n28900 = n313 | n3207 ;
  assign n28901 = n28900 ^ n2338 ^ 1'b0 ;
  assign n28902 = n28901 ^ n17920 ^ 1'b0 ;
  assign n28903 = n7896 & ~n28902 ;
  assign n28904 = n7739 & ~n20424 ;
  assign n28905 = ( n15052 & n16524 ) | ( n15052 & ~n28265 ) | ( n16524 & ~n28265 ) ;
  assign n28906 = n28905 ^ n19052 ^ n17697 ;
  assign n28907 = ( ~n1597 & n2109 ) | ( ~n1597 & n13249 ) | ( n2109 & n13249 ) ;
  assign n28908 = ~n26855 & n28907 ;
  assign n28909 = n18149 ^ n9858 ^ 1'b0 ;
  assign n28910 = n12441 & n22807 ;
  assign n28911 = n4744 & n28910 ;
  assign n28912 = ( ~n4918 & n28596 ) | ( ~n4918 & n28911 ) | ( n28596 & n28911 ) ;
  assign n28913 = n19619 ^ n16054 ^ 1'b0 ;
  assign n28915 = n2195 & ~n8701 ;
  assign n28914 = ~n3022 & n27535 ;
  assign n28916 = n28915 ^ n28914 ^ n26786 ;
  assign n28917 = ( n3552 & n6688 ) | ( n3552 & n16645 ) | ( n6688 & n16645 ) ;
  assign n28918 = n28917 ^ n14861 ^ 1'b0 ;
  assign n28919 = n27074 ^ n7641 ^ 1'b0 ;
  assign n28920 = n10228 | n28919 ;
  assign n28921 = n9689 & n25701 ;
  assign n28922 = n9137 | n21040 ;
  assign n28923 = n8977 ^ n4576 ^ 1'b0 ;
  assign n28924 = n20672 ^ n7962 ^ n7697 ;
  assign n28925 = ( n21671 & n22523 ) | ( n21671 & ~n27433 ) | ( n22523 & ~n27433 ) ;
  assign n28926 = n17185 ^ n10040 ^ 1'b0 ;
  assign n28927 = n3780 ^ n814 ^ 1'b0 ;
  assign n28928 = n2894 & n28927 ;
  assign n28929 = n8335 & n27377 ;
  assign n28930 = n14694 & ~n28929 ;
  assign n28931 = ( ~n12138 & n17941 ) | ( ~n12138 & n28634 ) | ( n17941 & n28634 ) ;
  assign n28932 = n28931 ^ n15510 ^ n4149 ;
  assign n28933 = n12099 | n28932 ;
  assign n28934 = n28933 ^ n17954 ^ 1'b0 ;
  assign n28935 = ~n11091 & n17414 ;
  assign n28937 = n1873 & n11804 ;
  assign n28936 = n24386 ^ n2219 ^ 1'b0 ;
  assign n28938 = n28937 ^ n28936 ^ n11128 ;
  assign n28939 = n28935 | n28938 ;
  assign n28940 = n28939 ^ n28715 ^ 1'b0 ;
  assign n28941 = ( x58 & n4189 ) | ( x58 & ~n11597 ) | ( n4189 & ~n11597 ) ;
  assign n28942 = ( n2655 & n4259 ) | ( n2655 & ~n10369 ) | ( n4259 & ~n10369 ) ;
  assign n28943 = n21838 ^ n8711 ^ n7750 ;
  assign n28944 = n5974 ^ n3111 ^ n164 ;
  assign n28945 = n12207 ^ n10076 ^ n7463 ;
  assign n28946 = ( n2834 & n28944 ) | ( n2834 & ~n28945 ) | ( n28944 & ~n28945 ) ;
  assign n28947 = n11411 ^ n7998 ^ 1'b0 ;
  assign n28948 = n28824 ^ n2189 ^ 1'b0 ;
  assign n28949 = n12054 ^ n10731 ^ 1'b0 ;
  assign n28950 = n9551 | n28949 ;
  assign n28951 = n28950 ^ n17071 ^ 1'b0 ;
  assign n28952 = n4815 | n9735 ;
  assign n28953 = n28952 ^ n24064 ^ 1'b0 ;
  assign n28954 = ~n23764 & n28953 ;
  assign n28955 = n25517 ^ n21434 ^ n6656 ;
  assign n28956 = n18086 ^ n11435 ^ 1'b0 ;
  assign n28957 = n28955 | n28956 ;
  assign n28958 = n4401 ^ n888 ^ n581 ;
  assign n28959 = ( n4403 & n7681 ) | ( n4403 & n28958 ) | ( n7681 & n28958 ) ;
  assign n28960 = n22668 ^ n11956 ^ 1'b0 ;
  assign n28962 = n23181 ^ n6485 ^ n2450 ;
  assign n28961 = n20339 ^ n3826 ^ n2424 ;
  assign n28963 = n28962 ^ n28961 ^ n20092 ;
  assign n28964 = n20276 ^ n12136 ^ 1'b0 ;
  assign n28965 = n24053 & ~n28255 ;
  assign n28966 = n24546 & n28965 ;
  assign n28967 = n28966 ^ n26872 ^ 1'b0 ;
  assign n28968 = ( n10441 & n28964 ) | ( n10441 & ~n28967 ) | ( n28964 & ~n28967 ) ;
  assign n28969 = n10201 & ~n12691 ;
  assign n28970 = n3664 & n10480 ;
  assign n28971 = ~n13072 & n28970 ;
  assign n28972 = ( n826 & n9359 ) | ( n826 & ~n28971 ) | ( n9359 & ~n28971 ) ;
  assign n28973 = n858 & n20450 ;
  assign n28974 = n28972 & n28973 ;
  assign n28975 = n21567 ^ n13349 ^ n12554 ;
  assign n28976 = n8782 & ~n28975 ;
  assign n28977 = n28976 ^ n19040 ^ 1'b0 ;
  assign n28978 = n13860 ^ n9479 ^ n1205 ;
  assign n28979 = n13657 ^ n9058 ^ 1'b0 ;
  assign n28980 = n15807 & ~n28979 ;
  assign n28981 = n28978 & n28980 ;
  assign n28982 = n28981 ^ n26363 ^ n4414 ;
  assign n28983 = ( ~n6151 & n15532 ) | ( ~n6151 & n28982 ) | ( n15532 & n28982 ) ;
  assign n28984 = n7838 & ~n19707 ;
  assign n28985 = n18003 ^ n16721 ^ 1'b0 ;
  assign n28986 = n8482 ^ n4541 ^ x71 ;
  assign n28987 = n8346 | n28986 ;
  assign n28988 = n20356 | n28987 ;
  assign n28989 = n28988 ^ n20569 ^ 1'b0 ;
  assign n28990 = n11694 & n17083 ;
  assign n28991 = n28990 ^ n780 ^ 1'b0 ;
  assign n28992 = ~n18014 & n28991 ;
  assign n28993 = ( n14762 & ~n27763 ) | ( n14762 & n28992 ) | ( ~n27763 & n28992 ) ;
  assign n28994 = n13071 ^ n11867 ^ n2055 ;
  assign n28995 = n4960 ^ n4220 ^ 1'b0 ;
  assign n28996 = ~n12072 & n28995 ;
  assign n28997 = n1590 & n2190 ;
  assign n28998 = n28997 ^ n20887 ^ 1'b0 ;
  assign n28999 = n8207 ^ n4667 ^ 1'b0 ;
  assign n29000 = n24918 & ~n28999 ;
  assign n29001 = ( n511 & n11950 ) | ( n511 & ~n15866 ) | ( n11950 & ~n15866 ) ;
  assign n29002 = n29001 ^ n20110 ^ 1'b0 ;
  assign n29003 = n6646 & ~n29002 ;
  assign n29004 = n19071 ^ n16035 ^ n5868 ;
  assign n29005 = n29004 ^ n10982 ^ n3980 ;
  assign n29006 = n24960 ^ n14011 ^ n3220 ;
  assign n29007 = n7836 & ~n18104 ;
  assign n29008 = n11583 ^ n8942 ^ n3662 ;
  assign n29009 = ( n17898 & ~n19844 ) | ( n17898 & n29008 ) | ( ~n19844 & n29008 ) ;
  assign n29010 = n4161 ^ n1083 ^ 1'b0 ;
  assign n29011 = ~n9137 & n29010 ;
  assign n29012 = ( n2661 & ~n3892 ) | ( n2661 & n29011 ) | ( ~n3892 & n29011 ) ;
  assign n29013 = ( n9471 & n26583 ) | ( n9471 & n29012 ) | ( n26583 & n29012 ) ;
  assign n29014 = n12955 ^ n3452 ^ n281 ;
  assign n29018 = ~n4100 & n10046 ;
  assign n29019 = n29018 ^ n22365 ^ 1'b0 ;
  assign n29016 = n4204 & ~n4271 ;
  assign n29017 = n29016 ^ n10295 ^ 1'b0 ;
  assign n29020 = n29019 ^ n29017 ^ n3632 ;
  assign n29015 = n6533 & ~n24434 ;
  assign n29021 = n29020 ^ n29015 ^ 1'b0 ;
  assign n29022 = n16835 & ~n29021 ;
  assign n29023 = n28266 ^ n27072 ^ n25271 ;
  assign n29024 = n4660 | n29023 ;
  assign n29025 = n18207 & ~n29024 ;
  assign n29026 = n24433 ^ n11549 ^ n9539 ;
  assign n29027 = ~n14721 & n29026 ;
  assign n29028 = n29027 ^ n3159 ^ 1'b0 ;
  assign n29029 = n18891 ^ n5538 ^ n4196 ;
  assign n29030 = ~n19872 & n24269 ;
  assign n29031 = ~n23975 & n29030 ;
  assign n29032 = n9367 & ~n29031 ;
  assign n29033 = n20658 & n29032 ;
  assign n29034 = ( n9865 & ~n11065 ) | ( n9865 & n29033 ) | ( ~n11065 & n29033 ) ;
  assign n29035 = n17227 ^ n13836 ^ n1834 ;
  assign n29036 = ( n3475 & ~n8084 ) | ( n3475 & n11881 ) | ( ~n8084 & n11881 ) ;
  assign n29037 = ( n3809 & n19900 ) | ( n3809 & n29036 ) | ( n19900 & n29036 ) ;
  assign n29038 = n9695 ^ n6287 ^ 1'b0 ;
  assign n29039 = ~n3238 & n5865 ;
  assign n29040 = ( n10099 & n12056 ) | ( n10099 & ~n29039 ) | ( n12056 & ~n29039 ) ;
  assign n29041 = ( x22 & n8119 ) | ( x22 & ~n29040 ) | ( n8119 & ~n29040 ) ;
  assign n29042 = n11911 & ~n23299 ;
  assign n29043 = n3451 | n29042 ;
  assign n29044 = n29041 | n29043 ;
  assign n29045 = n16076 ^ n3138 ^ 1'b0 ;
  assign n29046 = n15273 & ~n29045 ;
  assign n29047 = ~n12347 & n29046 ;
  assign n29048 = n29047 ^ n15181 ^ 1'b0 ;
  assign n29049 = n8769 & n28245 ;
  assign n29050 = n17049 | n28633 ;
  assign n29051 = n29050 ^ n20544 ^ 1'b0 ;
  assign n29052 = ( n4796 & n5296 ) | ( n4796 & n21332 ) | ( n5296 & n21332 ) ;
  assign n29053 = ( n4918 & n26155 ) | ( n4918 & ~n29052 ) | ( n26155 & ~n29052 ) ;
  assign n29054 = ( n5634 & ~n15949 ) | ( n5634 & n20567 ) | ( ~n15949 & n20567 ) ;
  assign n29055 = n29054 ^ n3150 ^ n1811 ;
  assign n29056 = ( n1533 & ~n22963 ) | ( n1533 & n26960 ) | ( ~n22963 & n26960 ) ;
  assign n29057 = n17089 ^ n9000 ^ 1'b0 ;
  assign n29058 = n4287 | n18912 ;
  assign n29059 = n16976 | n22141 ;
  assign n29060 = n29059 ^ n15805 ^ 1'b0 ;
  assign n29061 = n3453 & ~n8084 ;
  assign n29062 = ~n6699 & n29061 ;
  assign n29063 = n21026 ^ n1693 ^ 1'b0 ;
  assign n29064 = n13030 & ~n16547 ;
  assign n29065 = ~n14457 & n29064 ;
  assign n29070 = ( ~n1899 & n3937 ) | ( ~n1899 & n8462 ) | ( n3937 & n8462 ) ;
  assign n29069 = ( n4863 & ~n13341 ) | ( n4863 & n16807 ) | ( ~n13341 & n16807 ) ;
  assign n29067 = n2455 & n11515 ;
  assign n29066 = ~n9291 & n23130 ;
  assign n29068 = n29067 ^ n29066 ^ 1'b0 ;
  assign n29071 = n29070 ^ n29069 ^ n29068 ;
  assign n29072 = n23574 ^ n4110 ^ 1'b0 ;
  assign n29073 = n291 & n29072 ;
  assign n29074 = n1996 ^ n345 ^ 1'b0 ;
  assign n29075 = n26919 ^ n9360 ^ 1'b0 ;
  assign n29076 = n5527 & n29075 ;
  assign n29077 = n29076 ^ n2637 ^ 1'b0 ;
  assign n29078 = n4150 ^ n2573 ^ n2144 ;
  assign n29079 = ~n27229 & n29078 ;
  assign n29080 = n29079 ^ n8465 ^ 1'b0 ;
  assign n29081 = ( n9915 & ~n11686 ) | ( n9915 & n29080 ) | ( ~n11686 & n29080 ) ;
  assign n29082 = n6773 ^ n531 ^ 1'b0 ;
  assign n29083 = n26416 | n29082 ;
  assign n29084 = ( n6043 & n10428 ) | ( n6043 & ~n21384 ) | ( n10428 & ~n21384 ) ;
  assign n29085 = n16914 ^ n13360 ^ n2304 ;
  assign n29086 = n16518 | n29085 ;
  assign n29087 = n4877 | n29086 ;
  assign n29088 = n29084 | n29087 ;
  assign n29089 = ( ~n9096 & n29083 ) | ( ~n9096 & n29088 ) | ( n29083 & n29088 ) ;
  assign n29090 = n10780 ^ n10059 ^ 1'b0 ;
  assign n29091 = n2426 & ~n29090 ;
  assign n29092 = ~n7299 & n14661 ;
  assign n29093 = n17250 ^ n12559 ^ 1'b0 ;
  assign n29094 = ~n29092 & n29093 ;
  assign n29095 = n19241 ^ n8667 ^ n3877 ;
  assign n29096 = n7033 ^ n4931 ^ n1284 ;
  assign n29097 = n29096 ^ n16107 ^ n14460 ;
  assign n29098 = ( n7409 & n11548 ) | ( n7409 & n15240 ) | ( n11548 & n15240 ) ;
  assign n29099 = n29098 ^ n24862 ^ n14578 ;
  assign n29100 = n2705 & n23675 ;
  assign n29101 = ( n7180 & n29099 ) | ( n7180 & ~n29100 ) | ( n29099 & ~n29100 ) ;
  assign n29102 = ~n2170 & n10901 ;
  assign n29103 = n29102 ^ n28832 ^ n4601 ;
  assign n29104 = ( ~n4968 & n12774 ) | ( ~n4968 & n26379 ) | ( n12774 & n26379 ) ;
  assign n29105 = ~n3956 & n22988 ;
  assign n29106 = ~n2016 & n29105 ;
  assign n29107 = ~n17106 & n18962 ;
  assign n29108 = n1476 & n29107 ;
  assign n29109 = n29108 ^ n15096 ^ 1'b0 ;
  assign n29110 = n16498 ^ n1742 ^ 1'b0 ;
  assign n29111 = n19302 & n29110 ;
  assign n29112 = n16167 ^ n2935 ^ 1'b0 ;
  assign n29113 = n20764 & n29112 ;
  assign n29114 = n3744 & n29113 ;
  assign n29115 = n11428 & n13378 ;
  assign n29116 = ~n12503 & n29115 ;
  assign n29117 = ( n1994 & n3763 ) | ( n1994 & n29116 ) | ( n3763 & n29116 ) ;
  assign n29118 = n9637 | n29117 ;
  assign n29119 = n1276 & ~n6798 ;
  assign n29120 = n29119 ^ n1651 ^ 1'b0 ;
  assign n29121 = n29120 ^ n15501 ^ n14293 ;
  assign n29122 = n29121 ^ n14472 ^ n11411 ;
  assign n29123 = n24332 ^ n22619 ^ n4022 ;
  assign n29124 = ~n1763 & n4884 ;
  assign n29125 = n10156 & n29124 ;
  assign n29126 = ( n3628 & n26855 ) | ( n3628 & ~n29125 ) | ( n26855 & ~n29125 ) ;
  assign n29127 = n29126 ^ n20972 ^ n2094 ;
  assign n29128 = n1669 & ~n1885 ;
  assign n29129 = n29128 ^ n5026 ^ 1'b0 ;
  assign n29130 = ( n904 & n7546 ) | ( n904 & ~n10304 ) | ( n7546 & ~n10304 ) ;
  assign n29131 = n27490 ^ n18536 ^ 1'b0 ;
  assign n29132 = n29130 & n29131 ;
  assign n29133 = n20088 ^ x19 ^ 1'b0 ;
  assign n29134 = n3794 | n29133 ;
  assign n29135 = n11075 ^ n1442 ^ 1'b0 ;
  assign n29136 = n9847 & ~n29135 ;
  assign n29137 = n28512 ^ n6807 ^ n4020 ;
  assign n29138 = ( n9128 & ~n9675 ) | ( n9128 & n11075 ) | ( ~n9675 & n11075 ) ;
  assign n29139 = n29138 ^ n15438 ^ n4542 ;
  assign n29141 = n12091 ^ n5561 ^ 1'b0 ;
  assign n29140 = n5967 & n27132 ;
  assign n29142 = n29141 ^ n29140 ^ 1'b0 ;
  assign n29143 = n13925 ^ n5681 ^ n4663 ;
  assign n29145 = ( n6499 & n10057 ) | ( n6499 & ~n20400 ) | ( n10057 & ~n20400 ) ;
  assign n29144 = n4434 & n24260 ;
  assign n29146 = n29145 ^ n29144 ^ n6617 ;
  assign n29147 = ( ~n29142 & n29143 ) | ( ~n29142 & n29146 ) | ( n29143 & n29146 ) ;
  assign n29148 = n9236 | n17472 ;
  assign n29149 = n19064 | n29148 ;
  assign n29150 = n9347 | n18812 ;
  assign n29151 = n6934 | n28286 ;
  assign n29152 = n29150 & ~n29151 ;
  assign n29153 = n9296 & n16724 ;
  assign n29154 = n29153 ^ n2584 ^ 1'b0 ;
  assign n29155 = n3253 ^ n287 ^ 1'b0 ;
  assign n29156 = ~n3512 & n29155 ;
  assign n29157 = ~n13278 & n29156 ;
  assign n29158 = ~n13092 & n29157 ;
  assign n29159 = n967 & n12787 ;
  assign n29160 = n29158 & n29159 ;
  assign n29161 = ~n10701 & n29160 ;
  assign n29162 = n413 & ~n16230 ;
  assign n29163 = ( ~n3828 & n23204 ) | ( ~n3828 & n28073 ) | ( n23204 & n28073 ) ;
  assign n29164 = n5669 & ~n21858 ;
  assign n29165 = n14981 & n21916 ;
  assign n29166 = n16363 ^ n3828 ^ 1'b0 ;
  assign n29167 = n28006 ^ n25529 ^ n16199 ;
  assign n29168 = x16 & ~n20166 ;
  assign n29169 = n4230 & n29168 ;
  assign n29170 = n5708 ^ n1942 ^ n1268 ;
  assign n29171 = n29170 ^ n6047 ^ 1'b0 ;
  assign n29172 = ~n16410 & n29171 ;
  assign n29173 = n14897 | n14977 ;
  assign n29174 = n29173 ^ n2964 ^ 1'b0 ;
  assign n29175 = n22613 ^ n14472 ^ 1'b0 ;
  assign n29176 = ~n3836 & n29175 ;
  assign n29177 = n15333 & n19517 ;
  assign n29178 = n29177 ^ n11244 ^ 1'b0 ;
  assign n29179 = n29178 ^ n25195 ^ n7909 ;
  assign n29182 = ( n5711 & n11272 ) | ( n5711 & n14276 ) | ( n11272 & n14276 ) ;
  assign n29180 = n3285 | n10113 ;
  assign n29181 = n7549 & ~n29180 ;
  assign n29183 = n29182 ^ n29181 ^ n11544 ;
  assign n29184 = ( n14567 & ~n17982 ) | ( n14567 & n22731 ) | ( ~n17982 & n22731 ) ;
  assign n29185 = ~n1029 & n14661 ;
  assign n29186 = ~n18009 & n29185 ;
  assign n29187 = n17274 ^ n6048 ^ 1'b0 ;
  assign n29188 = n10749 | n29187 ;
  assign n29189 = n2215 & n5932 ;
  assign n29190 = n29189 ^ n28612 ^ n6955 ;
  assign n29191 = ~n6667 & n20331 ;
  assign n29192 = n29191 ^ n20408 ^ 1'b0 ;
  assign n29193 = n29192 ^ n18905 ^ 1'b0 ;
  assign n29194 = ~n29190 & n29193 ;
  assign n29195 = n1083 & ~n19953 ;
  assign n29196 = n734 & n5482 ;
  assign n29197 = n29196 ^ n2663 ^ 1'b0 ;
  assign n29198 = n29197 ^ n28030 ^ n6864 ;
  assign n29199 = n20102 ^ n11940 ^ 1'b0 ;
  assign n29200 = n29199 ^ n26128 ^ n20711 ;
  assign n29201 = n2192 & n5516 ;
  assign n29202 = n29201 ^ n6319 ^ 1'b0 ;
  assign n29203 = ~n24675 & n29202 ;
  assign n29204 = n4713 | n17166 ;
  assign n29205 = ( ~n1376 & n5181 ) | ( ~n1376 & n14612 ) | ( n5181 & n14612 ) ;
  assign n29206 = ( n3598 & n18279 ) | ( n3598 & n29205 ) | ( n18279 & n29205 ) ;
  assign n29207 = n11873 ^ n3854 ^ 1'b0 ;
  assign n29208 = ~n15313 & n24485 ;
  assign n29209 = n18114 ^ n11387 ^ n1068 ;
  assign n29211 = ( n866 & n2253 ) | ( n866 & ~n20262 ) | ( n2253 & ~n20262 ) ;
  assign n29210 = n18195 ^ n7929 ^ n6236 ;
  assign n29212 = n29211 ^ n29210 ^ n5393 ;
  assign n29213 = n10581 ^ n9991 ^ 1'b0 ;
  assign n29214 = n15137 ^ n6166 ^ n4392 ;
  assign n29215 = ( ~n8920 & n9910 ) | ( ~n8920 & n29214 ) | ( n9910 & n29214 ) ;
  assign n29216 = n28395 | n29215 ;
  assign n29217 = ( ~n4649 & n29213 ) | ( ~n4649 & n29216 ) | ( n29213 & n29216 ) ;
  assign n29218 = ( n1388 & ~n8985 ) | ( n1388 & n9380 ) | ( ~n8985 & n9380 ) ;
  assign n29219 = ( n288 & n786 ) | ( n288 & ~n29218 ) | ( n786 & ~n29218 ) ;
  assign n29220 = ( n14299 & n16622 ) | ( n14299 & n29219 ) | ( n16622 & n29219 ) ;
  assign n29221 = ( n3159 & n23779 ) | ( n3159 & n29220 ) | ( n23779 & n29220 ) ;
  assign n29222 = n4055 ^ n2270 ^ 1'b0 ;
  assign n29223 = n1814 & n7594 ;
  assign n29224 = n29223 ^ n11665 ^ 1'b0 ;
  assign n29225 = ~n17062 & n22387 ;
  assign n29226 = n29225 ^ n20509 ^ 1'b0 ;
  assign n29227 = ( n2636 & ~n4234 ) | ( n2636 & n8691 ) | ( ~n4234 & n8691 ) ;
  assign n29228 = n3662 & ~n24298 ;
  assign n29229 = n29228 ^ n23496 ^ n7308 ;
  assign n29230 = n16393 ^ n14950 ^ 1'b0 ;
  assign n29231 = n5793 | n11454 ;
  assign n29232 = n29231 ^ n2850 ^ 1'b0 ;
  assign n29233 = ( ~n7441 & n18196 ) | ( ~n7441 & n29232 ) | ( n18196 & n29232 ) ;
  assign n29234 = n8847 ^ n6841 ^ 1'b0 ;
  assign n29235 = ~n6025 & n29234 ;
  assign n29236 = ( n14531 & n22721 ) | ( n14531 & ~n29235 ) | ( n22721 & ~n29235 ) ;
  assign n29237 = n15084 ^ n12024 ^ 1'b0 ;
  assign n29238 = n20104 | n29237 ;
  assign n29239 = n413 | n29238 ;
  assign n29240 = n19077 & ~n25052 ;
  assign n29241 = ~n14082 & n29240 ;
  assign n29242 = ~n8655 & n9819 ;
  assign n29243 = n29242 ^ n4568 ^ 1'b0 ;
  assign n29244 = ~n4864 & n7973 ;
  assign n29245 = n29244 ^ n22488 ^ 1'b0 ;
  assign n29246 = n14307 ^ n9135 ^ n4537 ;
  assign n29247 = n18791 ^ n18033 ^ 1'b0 ;
  assign n29248 = n29247 ^ n12926 ^ n4077 ;
  assign n29249 = ~n19179 & n29248 ;
  assign n29250 = n29249 ^ n14255 ^ n11482 ;
  assign n29251 = n15854 ^ n3766 ^ 1'b0 ;
  assign n29252 = n29251 ^ n11053 ^ n5694 ;
  assign n29253 = n9411 & n9642 ;
  assign n29254 = ~n7225 & n29253 ;
  assign n29255 = n10480 | n21615 ;
  assign n29256 = n29254 & n29255 ;
  assign n29257 = n29256 ^ n11547 ^ n4144 ;
  assign n29258 = n1366 & n29257 ;
  assign n29259 = n8103 & n10449 ;
  assign n29260 = n4252 | n26715 ;
  assign n29261 = n29260 ^ n25813 ^ 1'b0 ;
  assign n29262 = n6850 & n22351 ;
  assign n29263 = n29262 ^ n25271 ^ 1'b0 ;
  assign n29264 = n19356 ^ n10918 ^ 1'b0 ;
  assign n29265 = n8760 & n29264 ;
  assign n29266 = n2045 | n9855 ;
  assign n29267 = n29265 | n29266 ;
  assign n29268 = ( n6695 & n15770 ) | ( n6695 & n28116 ) | ( n15770 & n28116 ) ;
  assign n29269 = n9208 & ~n29268 ;
  assign n29270 = n25010 ^ n17701 ^ 1'b0 ;
  assign n29271 = ( n652 & n4654 ) | ( n652 & n19524 ) | ( n4654 & n19524 ) ;
  assign n29272 = ( n12409 & n16691 ) | ( n12409 & n25326 ) | ( n16691 & n25326 ) ;
  assign n29273 = n9260 ^ n6792 ^ n3684 ;
  assign n29274 = ( n3378 & n18631 ) | ( n3378 & ~n28717 ) | ( n18631 & ~n28717 ) ;
  assign n29275 = n13267 ^ n577 ^ n305 ;
  assign n29276 = n18338 & n29275 ;
  assign n29277 = n29276 ^ n3234 ^ 1'b0 ;
  assign n29278 = ~n133 & n3070 ;
  assign n29279 = ~n3070 & n29278 ;
  assign n29280 = ( n4514 & n7586 ) | ( n4514 & n29279 ) | ( n7586 & n29279 ) ;
  assign n29281 = n29280 ^ n17094 ^ 1'b0 ;
  assign n29282 = n20452 & n26667 ;
  assign n29283 = n29282 ^ n4331 ^ 1'b0 ;
  assign n29284 = n14424 ^ n4396 ^ n1739 ;
  assign n29285 = ~n5781 & n13648 ;
  assign n29286 = n15687 ^ n6072 ^ n2801 ;
  assign n29287 = n29286 ^ n24127 ^ n4190 ;
  assign n29288 = ( ~n20672 & n29285 ) | ( ~n20672 & n29287 ) | ( n29285 & n29287 ) ;
  assign n29289 = n5912 & ~n8724 ;
  assign n29290 = ( n9992 & ~n28741 ) | ( n9992 & n29289 ) | ( ~n28741 & n29289 ) ;
  assign n29291 = n29290 ^ n28937 ^ n12563 ;
  assign n29292 = n157 | n2736 ;
  assign n29293 = n10601 ^ n7024 ^ 1'b0 ;
  assign n29294 = ( n16148 & n29292 ) | ( n16148 & ~n29293 ) | ( n29292 & ~n29293 ) ;
  assign n29295 = n16074 & n24054 ;
  assign n29296 = ~n18598 & n29295 ;
  assign n29297 = ~n5587 & n29296 ;
  assign n29298 = n770 & n5483 ;
  assign n29299 = ~n6786 & n29298 ;
  assign n29300 = ( ~n8435 & n11242 ) | ( ~n8435 & n29299 ) | ( n11242 & n29299 ) ;
  assign n29301 = n29300 ^ n28714 ^ n13444 ;
  assign n29304 = n6749 & ~n6884 ;
  assign n29305 = n29304 ^ n19500 ^ 1'b0 ;
  assign n29302 = n17836 ^ n8766 ^ 1'b0 ;
  assign n29303 = n24506 | n29302 ;
  assign n29306 = n29305 ^ n29303 ^ n3903 ;
  assign n29307 = ( n15374 & ~n19432 ) | ( n15374 & n29306 ) | ( ~n19432 & n29306 ) ;
  assign n29308 = n19507 ^ n10313 ^ 1'b0 ;
  assign n29309 = ~n21164 & n22533 ;
  assign n29310 = ~n12968 & n29309 ;
  assign n29311 = n29310 ^ n19091 ^ n3678 ;
  assign n29312 = ~n29308 & n29311 ;
  assign n29313 = n29312 ^ n7726 ^ 1'b0 ;
  assign n29315 = n9124 & ~n9845 ;
  assign n29316 = n29315 ^ n17185 ^ n12986 ;
  assign n29317 = ( n4512 & n16535 ) | ( n4512 & n29316 ) | ( n16535 & n29316 ) ;
  assign n29314 = n7154 ^ n4421 ^ n3666 ;
  assign n29318 = n29317 ^ n29314 ^ 1'b0 ;
  assign n29319 = n10456 ^ n2661 ^ n472 ;
  assign n29322 = n14411 ^ n2466 ^ 1'b0 ;
  assign n29320 = ~n3926 & n17343 ;
  assign n29321 = n29320 ^ n25769 ^ n18410 ;
  assign n29323 = n29322 ^ n29321 ^ 1'b0 ;
  assign n29324 = n3711 & n29323 ;
  assign n29325 = n26817 ^ n7062 ^ n2934 ;
  assign n29326 = n29325 ^ n9385 ^ 1'b0 ;
  assign n29327 = ( ~n24457 & n29324 ) | ( ~n24457 & n29326 ) | ( n29324 & n29326 ) ;
  assign n29328 = ( n6899 & n12286 ) | ( n6899 & n22828 ) | ( n12286 & n22828 ) ;
  assign n29329 = n29328 ^ n17719 ^ n15913 ;
  assign n29330 = ( n9207 & n23683 ) | ( n9207 & ~n29329 ) | ( n23683 & ~n29329 ) ;
  assign n29331 = n5384 ^ n4050 ^ 1'b0 ;
  assign n29332 = n23284 ^ n17599 ^ n3522 ;
  assign n29333 = n24455 & n28630 ;
  assign n29334 = ~n23409 & n29333 ;
  assign n29335 = n8286 | n9221 ;
  assign n29336 = n26901 | n29335 ;
  assign n29337 = ( n1942 & n14271 ) | ( n1942 & ~n22022 ) | ( n14271 & ~n22022 ) ;
  assign n29338 = n19837 ^ n17265 ^ n5245 ;
  assign n29339 = ~n25712 & n29338 ;
  assign n29340 = n29337 & n29339 ;
  assign n29341 = n6436 | n21230 ;
  assign n29342 = n29341 ^ n27322 ^ 1'b0 ;
  assign n29343 = n4312 ^ n2236 ^ 1'b0 ;
  assign n29350 = n6182 & n24706 ;
  assign n29347 = ~n1157 & n14247 ;
  assign n29348 = n29347 ^ n5329 ^ 1'b0 ;
  assign n29345 = ( n9539 & n11044 ) | ( n9539 & ~n15713 ) | ( n11044 & ~n15713 ) ;
  assign n29344 = n2204 & n18437 ;
  assign n29346 = n29345 ^ n29344 ^ 1'b0 ;
  assign n29349 = n29348 ^ n29346 ^ n6568 ;
  assign n29351 = n29350 ^ n29349 ^ n25466 ;
  assign n29352 = n2108 | n13105 ;
  assign n29353 = n11754 & ~n23052 ;
  assign n29354 = ( ~n12701 & n13974 ) | ( ~n12701 & n14586 ) | ( n13974 & n14586 ) ;
  assign n29355 = ( n7770 & n29353 ) | ( n7770 & ~n29354 ) | ( n29353 & ~n29354 ) ;
  assign n29356 = ( ~n775 & n29352 ) | ( ~n775 & n29355 ) | ( n29352 & n29355 ) ;
  assign n29357 = ( ~n10268 & n19684 ) | ( ~n10268 & n20902 ) | ( n19684 & n20902 ) ;
  assign n29358 = ( ~n2346 & n6085 ) | ( ~n2346 & n9391 ) | ( n6085 & n9391 ) ;
  assign n29359 = n29358 ^ n9407 ^ n7747 ;
  assign n29360 = n3836 ^ n828 ^ 1'b0 ;
  assign n29361 = n1509 & n29360 ;
  assign n29362 = ( ~n12196 & n12269 ) | ( ~n12196 & n29361 ) | ( n12269 & n29361 ) ;
  assign n29363 = n13008 & ~n16953 ;
  assign n29364 = ~n16291 & n29363 ;
  assign n29365 = n16381 ^ n15898 ^ n12403 ;
  assign n29366 = ~n12562 & n29365 ;
  assign n29367 = ~n9382 & n29366 ;
  assign n29368 = n7361 & ~n11773 ;
  assign n29369 = ~n8812 & n29368 ;
  assign n29370 = n18793 & ~n29369 ;
  assign n29371 = n29370 ^ n5865 ^ 1'b0 ;
  assign n29372 = n27058 ^ n9737 ^ n3995 ;
  assign n29373 = ~n937 & n13393 ;
  assign n29374 = n29373 ^ n5184 ^ 1'b0 ;
  assign n29375 = n1452 | n29374 ;
  assign n29376 = ( n1501 & n12242 ) | ( n1501 & n15329 ) | ( n12242 & n15329 ) ;
  assign n29377 = ~n9061 & n17086 ;
  assign n29378 = n6614 & n6799 ;
  assign n29379 = n29378 ^ n427 ^ 1'b0 ;
  assign n29380 = ( n2499 & n3678 ) | ( n2499 & ~n29379 ) | ( n3678 & ~n29379 ) ;
  assign n29382 = n9258 ^ n4750 ^ 1'b0 ;
  assign n29383 = ~n15805 & n29382 ;
  assign n29384 = ~n13447 & n29383 ;
  assign n29381 = n1690 & ~n11803 ;
  assign n29385 = n29384 ^ n29381 ^ 1'b0 ;
  assign n29386 = n5907 ^ n4158 ^ 1'b0 ;
  assign n29387 = x92 & n29386 ;
  assign n29388 = n13735 ^ n3619 ^ 1'b0 ;
  assign n29389 = n29387 & ~n29388 ;
  assign n29390 = n22187 ^ n14948 ^ 1'b0 ;
  assign n29391 = ( ~n5456 & n17910 ) | ( ~n5456 & n29390 ) | ( n17910 & n29390 ) ;
  assign n29392 = n1308 & n20886 ;
  assign n29393 = n29392 ^ n2857 ^ 1'b0 ;
  assign n29394 = n10565 ^ n3202 ^ 1'b0 ;
  assign n29395 = ( n7848 & ~n27987 ) | ( n7848 & n29394 ) | ( ~n27987 & n29394 ) ;
  assign n29396 = n23693 & ~n29395 ;
  assign n29397 = n29396 ^ n2866 ^ 1'b0 ;
  assign n29398 = n13296 ^ n8601 ^ 1'b0 ;
  assign n29399 = ~n738 & n29398 ;
  assign n29400 = ( n2029 & n9077 ) | ( n2029 & ~n12961 ) | ( n9077 & ~n12961 ) ;
  assign n29401 = n9272 & ~n11609 ;
  assign n29402 = n22304 & n29401 ;
  assign n29403 = ~n6937 & n29402 ;
  assign n29405 = n456 | n7898 ;
  assign n29406 = n27255 | n29405 ;
  assign n29404 = n3512 | n22721 ;
  assign n29407 = n29406 ^ n29404 ^ 1'b0 ;
  assign n29408 = n1624 | n10540 ;
  assign n29409 = n29408 ^ x124 ^ 1'b0 ;
  assign n29410 = n26322 ^ n5910 ^ 1'b0 ;
  assign n29411 = x1 & ~n29410 ;
  assign n29412 = n25822 ^ n20794 ^ n10128 ;
  assign n29413 = n27051 ^ n18467 ^ n14696 ;
  assign n29414 = n18116 ^ n8390 ^ n8078 ;
  assign n29415 = ( n1176 & n6379 ) | ( n1176 & ~n26220 ) | ( n6379 & ~n26220 ) ;
  assign n29416 = n8764 | n21052 ;
  assign n29417 = n29416 ^ n28762 ^ 1'b0 ;
  assign n29418 = n3334 | n29417 ;
  assign n29419 = n25352 ^ n11511 ^ 1'b0 ;
  assign n29420 = n1251 & n14928 ;
  assign n29422 = ( n6108 & ~n12129 ) | ( n6108 & n14788 ) | ( ~n12129 & n14788 ) ;
  assign n29421 = n25974 & ~n28272 ;
  assign n29423 = n29422 ^ n29421 ^ 1'b0 ;
  assign n29424 = ( n4304 & n19822 ) | ( n4304 & ~n22578 ) | ( n19822 & ~n22578 ) ;
  assign n29425 = n13998 & ~n29424 ;
  assign n29426 = ( n5342 & n9950 ) | ( n5342 & ~n29373 ) | ( n9950 & ~n29373 ) ;
  assign n29427 = n27235 ^ n17296 ^ n15569 ;
  assign n29428 = n12302 & n26537 ;
  assign n29429 = ~n676 & n11109 ;
  assign n29430 = ~n29428 & n29429 ;
  assign n29431 = ~n7867 & n29430 ;
  assign n29432 = n1867 & ~n25198 ;
  assign n29433 = n29432 ^ n11313 ^ 1'b0 ;
  assign n29434 = n10307 & ~n29433 ;
  assign n29435 = n29434 ^ n22396 ^ 1'b0 ;
  assign n29436 = n29435 ^ n20013 ^ n4824 ;
  assign n29437 = ( ~n20093 & n20655 ) | ( ~n20093 & n21673 ) | ( n20655 & n21673 ) ;
  assign n29439 = n3416 | n9336 ;
  assign n29440 = n29439 ^ n28675 ^ 1'b0 ;
  assign n29441 = ~n11179 & n25272 ;
  assign n29442 = ~n19880 & n29441 ;
  assign n29443 = ( ~n15329 & n29440 ) | ( ~n15329 & n29442 ) | ( n29440 & n29442 ) ;
  assign n29438 = n5704 | n5854 ;
  assign n29444 = n29443 ^ n29438 ^ 1'b0 ;
  assign n29445 = ~n4350 & n19740 ;
  assign n29446 = n29445 ^ n9471 ^ 1'b0 ;
  assign n29448 = n2684 ^ x118 ^ 1'b0 ;
  assign n29449 = n7042 & ~n29448 ;
  assign n29450 = ( n7689 & ~n14915 ) | ( n7689 & n29449 ) | ( ~n14915 & n29449 ) ;
  assign n29447 = ~n3420 & n5066 ;
  assign n29451 = n29450 ^ n29447 ^ 1'b0 ;
  assign n29452 = n881 | n1068 ;
  assign n29453 = n18916 ^ n18240 ^ 1'b0 ;
  assign n29454 = n12207 | n29453 ;
  assign n29455 = n4725 & n24613 ;
  assign n29456 = ~n6430 & n29455 ;
  assign n29457 = ( n3410 & n16298 ) | ( n3410 & ~n19181 ) | ( n16298 & ~n19181 ) ;
  assign n29458 = n26615 ^ n25266 ^ n9954 ;
  assign n29459 = ( ~n1171 & n6383 ) | ( ~n1171 & n12204 ) | ( n6383 & n12204 ) ;
  assign n29460 = n25745 ^ n23986 ^ n162 ;
  assign n29461 = n1725 & n13533 ;
  assign n29462 = n11688 & ~n19760 ;
  assign n29463 = n29462 ^ n18637 ^ 1'b0 ;
  assign n29464 = ( n8118 & n9261 ) | ( n8118 & n16147 ) | ( n9261 & n16147 ) ;
  assign n29465 = n15088 | n29464 ;
  assign n29466 = n29463 & ~n29465 ;
  assign n29467 = n871 & n7352 ;
  assign n29468 = ~n3560 & n29467 ;
  assign n29469 = n9296 ^ n2071 ^ 1'b0 ;
  assign n29470 = n18891 & ~n29469 ;
  assign n29471 = n29470 ^ n2312 ^ 1'b0 ;
  assign n29472 = n10174 & ~n29471 ;
  assign n29473 = n7257 | n12070 ;
  assign n29474 = ( n11531 & n23426 ) | ( n11531 & ~n29473 ) | ( n23426 & ~n29473 ) ;
  assign n29475 = ( ~n1664 & n14706 ) | ( ~n1664 & n21349 ) | ( n14706 & n21349 ) ;
  assign n29476 = n256 | n1714 ;
  assign n29477 = ( ~n6826 & n9687 ) | ( ~n6826 & n29476 ) | ( n9687 & n29476 ) ;
  assign n29478 = ~n4245 & n29088 ;
  assign n29479 = n11500 ^ n4793 ^ 1'b0 ;
  assign n29480 = n22672 ^ n147 ^ 1'b0 ;
  assign n29481 = ~n1729 & n22592 ;
  assign n29482 = n29481 ^ n409 ^ 1'b0 ;
  assign n29483 = ~n1665 & n7983 ;
  assign n29484 = ~n29482 & n29483 ;
  assign n29485 = n1865 ^ n1671 ^ 1'b0 ;
  assign n29486 = n2870 & ~n29485 ;
  assign n29487 = ~n11503 & n29486 ;
  assign n29488 = n29487 ^ n20036 ^ 1'b0 ;
  assign n29489 = n352 | n16251 ;
  assign n29490 = ~n6624 & n12038 ;
  assign n29491 = n29490 ^ n18835 ^ 1'b0 ;
  assign n29492 = n19507 ^ n17015 ^ 1'b0 ;
  assign n29493 = ( n2272 & n21804 ) | ( n2272 & n29492 ) | ( n21804 & n29492 ) ;
  assign n29494 = ( n23581 & n29491 ) | ( n23581 & ~n29493 ) | ( n29491 & ~n29493 ) ;
  assign n29495 = n1976 | n11442 ;
  assign n29496 = n10444 & ~n29495 ;
  assign n29497 = n29496 ^ n21313 ^ n11053 ;
  assign n29498 = n29497 ^ n13776 ^ 1'b0 ;
  assign n29499 = n12375 | n14654 ;
  assign n29500 = ( n4386 & ~n23795 ) | ( n4386 & n25239 ) | ( ~n23795 & n25239 ) ;
  assign n29503 = n14446 ^ n5396 ^ 1'b0 ;
  assign n29504 = n11143 & n29503 ;
  assign n29505 = n11487 ^ n6778 ^ n4860 ;
  assign n29506 = n29505 ^ n14495 ^ 1'b0 ;
  assign n29507 = n29504 | n29506 ;
  assign n29501 = ~n7637 & n9248 ;
  assign n29502 = n29501 ^ n10448 ^ 1'b0 ;
  assign n29508 = n29507 ^ n29502 ^ 1'b0 ;
  assign n29510 = n23618 ^ n10593 ^ n9666 ;
  assign n29511 = n22690 ^ n9840 ^ 1'b0 ;
  assign n29512 = ~n29510 & n29511 ;
  assign n29509 = n581 & ~n3605 ;
  assign n29513 = n29512 ^ n29509 ^ 1'b0 ;
  assign n29514 = n6172 & n13088 ;
  assign n29515 = n21015 & n23733 ;
  assign n29516 = n895 ^ n872 ^ 1'b0 ;
  assign n29517 = n18224 ^ n12139 ^ 1'b0 ;
  assign n29518 = ( n957 & n13189 ) | ( n957 & ~n29517 ) | ( n13189 & ~n29517 ) ;
  assign n29519 = n29353 ^ n20576 ^ n11021 ;
  assign n29520 = n24791 ^ n6927 ^ 1'b0 ;
  assign n29521 = ~n4333 & n29520 ;
  assign n29522 = ( ~n25795 & n26706 ) | ( ~n25795 & n29521 ) | ( n26706 & n29521 ) ;
  assign n29523 = n25341 ^ n21312 ^ n6849 ;
  assign n29524 = n6200 & ~n19489 ;
  assign n29525 = n575 & ~n6134 ;
  assign n29526 = n6736 & n29525 ;
  assign n29527 = n12600 ^ n7694 ^ 1'b0 ;
  assign n29528 = ~n949 & n12787 ;
  assign n29529 = ~n20802 & n29528 ;
  assign n29530 = n19826 ^ n16136 ^ n10897 ;
  assign n29531 = n7472 ^ n7288 ^ 1'b0 ;
  assign n29532 = ( ~n1636 & n4773 ) | ( ~n1636 & n9662 ) | ( n4773 & n9662 ) ;
  assign n29533 = ( n1685 & ~n9144 ) | ( n1685 & n29532 ) | ( ~n9144 & n29532 ) ;
  assign n29537 = n3509 & ~n28321 ;
  assign n29538 = n29537 ^ n14584 ^ 1'b0 ;
  assign n29534 = n4555 | n8718 ;
  assign n29535 = n415 & ~n29534 ;
  assign n29536 = ( ~n14243 & n24444 ) | ( ~n14243 & n29535 ) | ( n24444 & n29535 ) ;
  assign n29539 = n29538 ^ n29536 ^ 1'b0 ;
  assign n29540 = n10924 ^ n10784 ^ n6672 ;
  assign n29541 = n22483 ^ n2141 ^ 1'b0 ;
  assign n29542 = ~n17371 & n29541 ;
  assign n29543 = n28539 ^ n16837 ^ 1'b0 ;
  assign n29544 = n26558 | n29543 ;
  assign n29545 = n19427 ^ n3335 ^ 1'b0 ;
  assign n29546 = ~n29544 & n29545 ;
  assign n29547 = n189 & n24066 ;
  assign n29548 = x91 & ~n29547 ;
  assign n29549 = n5227 & n15535 ;
  assign n29550 = n29549 ^ n24886 ^ 1'b0 ;
  assign n29551 = ( n22372 & n22424 ) | ( n22372 & n29550 ) | ( n22424 & n29550 ) ;
  assign n29552 = ( ~n22090 & n29548 ) | ( ~n22090 & n29551 ) | ( n29548 & n29551 ) ;
  assign n29553 = n18062 ^ n12425 ^ n7620 ;
  assign n29554 = ( n541 & ~n2151 ) | ( n541 & n13764 ) | ( ~n2151 & n13764 ) ;
  assign n29555 = n12573 & n21356 ;
  assign n29556 = n6965 & n7090 ;
  assign n29557 = ~n3231 & n4974 ;
  assign n29558 = n29557 ^ n8270 ^ 1'b0 ;
  assign n29559 = n29558 ^ n7375 ^ 1'b0 ;
  assign n29560 = n7252 & ~n29559 ;
  assign n29561 = n29560 ^ n21541 ^ 1'b0 ;
  assign n29562 = n440 | n29561 ;
  assign n29563 = n8507 & ~n17823 ;
  assign n29564 = n7087 & ~n20153 ;
  assign n29565 = n22620 ^ n263 ^ 1'b0 ;
  assign n29566 = n9087 & ~n21298 ;
  assign n29567 = n23772 & n29566 ;
  assign n29568 = n29567 ^ n25545 ^ n2880 ;
  assign n29569 = ( n1606 & n6016 ) | ( n1606 & n19509 ) | ( n6016 & n19509 ) ;
  assign n29570 = n17755 ^ n16944 ^ n2118 ;
  assign n29571 = ( ~n10816 & n23427 ) | ( ~n10816 & n29570 ) | ( n23427 & n29570 ) ;
  assign n29572 = ~n3992 & n28373 ;
  assign n29573 = n29572 ^ n12926 ^ 1'b0 ;
  assign n29574 = ( n1097 & n4678 ) | ( n1097 & ~n29573 ) | ( n4678 & ~n29573 ) ;
  assign n29575 = n7570 & n15589 ;
  assign n29576 = n13891 & ~n29575 ;
  assign n29577 = ( n440 & n13391 ) | ( n440 & ~n24680 ) | ( n13391 & ~n24680 ) ;
  assign n29578 = ( n1255 & n23718 ) | ( n1255 & n29577 ) | ( n23718 & n29577 ) ;
  assign n29579 = n17040 | n29578 ;
  assign n29580 = n29579 ^ n4434 ^ 1'b0 ;
  assign n29581 = n13018 & n20235 ;
  assign n29582 = n29581 ^ n2301 ^ 1'b0 ;
  assign n29583 = n15057 | n29582 ;
  assign n29584 = ~n3207 & n17326 ;
  assign n29585 = n29584 ^ n5307 ^ 1'b0 ;
  assign n29586 = ( n7783 & n16762 ) | ( n7783 & ~n20867 ) | ( n16762 & ~n20867 ) ;
  assign n29587 = ~n13120 & n20517 ;
  assign n29588 = n23933 ^ n8475 ^ n1112 ;
  assign n29589 = n3136 & ~n4112 ;
  assign n29590 = ~n23797 & n29589 ;
  assign n29591 = n29590 ^ n20781 ^ 1'b0 ;
  assign n29592 = ( ~n10384 & n24013 ) | ( ~n10384 & n29591 ) | ( n24013 & n29591 ) ;
  assign n29593 = n18049 ^ n11794 ^ n2722 ;
  assign n29594 = n29593 ^ n18990 ^ 1'b0 ;
  assign n29595 = n23451 ^ n21291 ^ 1'b0 ;
  assign n29596 = n25653 & ~n29595 ;
  assign n29598 = n16909 ^ n13994 ^ n2456 ;
  assign n29599 = n8881 ^ n6635 ^ 1'b0 ;
  assign n29600 = n29598 | n29599 ;
  assign n29597 = n19775 & ~n21538 ;
  assign n29601 = n29600 ^ n29597 ^ 1'b0 ;
  assign n29604 = n7431 ^ n3186 ^ 1'b0 ;
  assign n29605 = n445 & n29604 ;
  assign n29602 = n16800 | n17091 ;
  assign n29603 = ~n27104 & n29602 ;
  assign n29606 = n29605 ^ n29603 ^ 1'b0 ;
  assign n29608 = n18008 ^ n3408 ^ 1'b0 ;
  assign n29609 = n8176 ^ n615 ^ 1'b0 ;
  assign n29610 = n29608 & n29609 ;
  assign n29607 = n16960 & n26286 ;
  assign n29611 = n29610 ^ n29607 ^ n15992 ;
  assign n29612 = n24357 ^ n13653 ^ n7051 ;
  assign n29613 = n10868 ^ n9474 ^ n461 ;
  assign n29614 = n29613 ^ n24467 ^ n909 ;
  assign n29615 = n29614 ^ n24580 ^ n5387 ;
  assign n29616 = ( ~n16389 & n20523 ) | ( ~n16389 & n23809 ) | ( n20523 & n23809 ) ;
  assign n29617 = n10301 ^ n3035 ^ n1118 ;
  assign n29618 = ( n27763 & n29616 ) | ( n27763 & n29617 ) | ( n29616 & n29617 ) ;
  assign n29619 = ~n878 & n3177 ;
  assign n29620 = ~n7911 & n29619 ;
  assign n29622 = n2466 & ~n12098 ;
  assign n29621 = n2897 | n9655 ;
  assign n29623 = n29622 ^ n29621 ^ 1'b0 ;
  assign n29624 = n16830 | n18639 ;
  assign n29625 = n29624 ^ n15163 ^ 1'b0 ;
  assign n29626 = n24326 ^ n14058 ^ n9655 ;
  assign n29627 = n18020 ^ n5056 ^ n3364 ;
  assign n29628 = ( n8664 & ~n11264 ) | ( n8664 & n29627 ) | ( ~n11264 & n29627 ) ;
  assign n29629 = n28051 ^ n5031 ^ n4610 ;
  assign n29630 = ( n1331 & n7727 ) | ( n1331 & ~n11642 ) | ( n7727 & ~n11642 ) ;
  assign n29631 = n29630 ^ n3517 ^ 1'b0 ;
  assign n29632 = ( n2160 & n26391 ) | ( n2160 & ~n29631 ) | ( n26391 & ~n29631 ) ;
  assign n29633 = n16796 ^ n10316 ^ n9208 ;
  assign n29634 = ( n1922 & n29538 ) | ( n1922 & ~n29633 ) | ( n29538 & ~n29633 ) ;
  assign n29635 = n10708 ^ n4351 ^ 1'b0 ;
  assign n29636 = n6847 | n29635 ;
  assign n29637 = n21446 ^ n14437 ^ x70 ;
  assign n29638 = ( n29634 & n29636 ) | ( n29634 & ~n29637 ) | ( n29636 & ~n29637 ) ;
  assign n29639 = ( x78 & n7083 ) | ( x78 & n12885 ) | ( n7083 & n12885 ) ;
  assign n29640 = ~n13964 & n28215 ;
  assign n29641 = n29640 ^ n11494 ^ 1'b0 ;
  assign n29642 = n8551 ^ n1228 ^ 1'b0 ;
  assign n29643 = n11195 ^ n3206 ^ 1'b0 ;
  assign n29644 = n9363 | n29643 ;
  assign n29645 = n29644 ^ n13577 ^ 1'b0 ;
  assign n29646 = ~n20537 & n29645 ;
  assign n29647 = n16433 & n29646 ;
  assign n29648 = n29647 ^ n29401 ^ 1'b0 ;
  assign n29649 = n11811 ^ n2496 ^ 1'b0 ;
  assign n29650 = n26224 ^ n12927 ^ n12677 ;
  assign n29651 = ( n9270 & n19071 ) | ( n9270 & n21272 ) | ( n19071 & n21272 ) ;
  assign n29652 = n8951 & n29651 ;
  assign n29653 = n26160 ^ n16136 ^ n2489 ;
  assign n29654 = n8548 ^ n5716 ^ n2161 ;
  assign n29655 = n29654 ^ n22885 ^ n3891 ;
  assign n29656 = n7987 ^ n7249 ^ 1'b0 ;
  assign n29657 = ( n4900 & ~n12973 ) | ( n4900 & n29656 ) | ( ~n12973 & n29656 ) ;
  assign n29658 = n27852 ^ n11003 ^ n6380 ;
  assign n29659 = n11055 ^ n7673 ^ 1'b0 ;
  assign n29660 = ~n26367 & n29659 ;
  assign n29661 = n18036 ^ n925 ^ 1'b0 ;
  assign n29662 = ~n20166 & n29661 ;
  assign n29663 = n19944 ^ n8119 ^ 1'b0 ;
  assign n29664 = n11526 & ~n29663 ;
  assign n29665 = n6903 | n11976 ;
  assign n29666 = n27875 & ~n29665 ;
  assign n29667 = n23430 ^ n11003 ^ 1'b0 ;
  assign n29668 = n20526 ^ n11091 ^ n351 ;
  assign n29669 = n29668 ^ n17372 ^ n1566 ;
  assign n29670 = ( n5073 & n10365 ) | ( n5073 & n21801 ) | ( n10365 & n21801 ) ;
  assign n29671 = ( ~n5847 & n9261 ) | ( ~n5847 & n19815 ) | ( n9261 & n19815 ) ;
  assign n29672 = n9102 & n17900 ;
  assign n29673 = n13920 & n29672 ;
  assign n29674 = ( n22062 & n25070 ) | ( n22062 & n29673 ) | ( n25070 & n29673 ) ;
  assign n29675 = ( n18723 & n20852 ) | ( n18723 & n27918 ) | ( n20852 & n27918 ) ;
  assign n29677 = n16768 ^ n2183 ^ n343 ;
  assign n29678 = n29677 ^ n6215 ^ 1'b0 ;
  assign n29676 = n731 & ~n2606 ;
  assign n29679 = n29678 ^ n29676 ^ 1'b0 ;
  assign n29681 = n1475 & ~n7194 ;
  assign n29680 = n7782 & n17392 ;
  assign n29682 = n29681 ^ n29680 ^ 1'b0 ;
  assign n29683 = n17776 ^ n9324 ^ 1'b0 ;
  assign n29684 = n9212 & n29683 ;
  assign n29685 = n27808 ^ n3955 ^ 1'b0 ;
  assign n29686 = ~n15069 & n29685 ;
  assign n29687 = n29686 ^ n6985 ^ n3587 ;
  assign n29688 = n3872 & n8395 ;
  assign n29689 = ~n14711 & n29688 ;
  assign n29690 = ( x115 & ~n2749 ) | ( x115 & n9630 ) | ( ~n2749 & n9630 ) ;
  assign n29691 = ( ~n5551 & n13599 ) | ( ~n5551 & n29690 ) | ( n13599 & n29690 ) ;
  assign n29692 = n8232 ^ n5398 ^ n5033 ;
  assign n29693 = ( n1509 & ~n20745 ) | ( n1509 & n29692 ) | ( ~n20745 & n29692 ) ;
  assign n29694 = n7728 & ~n9125 ;
  assign n29695 = n29694 ^ n9261 ^ n372 ;
  assign n29696 = ( ~n2914 & n11693 ) | ( ~n2914 & n21891 ) | ( n11693 & n21891 ) ;
  assign n29697 = n9158 ^ n3078 ^ 1'b0 ;
  assign n29698 = n2906 & ~n29697 ;
  assign n29699 = n21485 ^ n17936 ^ n15815 ;
  assign n29700 = n15875 & ~n29699 ;
  assign n29701 = ~n29698 & n29700 ;
  assign n29702 = n698 | n13182 ;
  assign n29706 = n26482 ^ n5836 ^ 1'b0 ;
  assign n29703 = n4585 | n9531 ;
  assign n29704 = n10165 | n29703 ;
  assign n29705 = ~n783 & n29704 ;
  assign n29707 = n29706 ^ n29705 ^ 1'b0 ;
  assign n29708 = n16979 ^ n5939 ^ n4189 ;
  assign n29709 = n18671 & ~n25871 ;
  assign n29710 = ( n6359 & ~n9646 ) | ( n6359 & n15045 ) | ( ~n9646 & n15045 ) ;
  assign n29711 = n15859 ^ n4275 ^ n1312 ;
  assign n29712 = n8505 ^ n850 ^ n376 ;
  assign n29713 = n5349 & ~n29712 ;
  assign n29714 = n29713 ^ n8910 ^ n4147 ;
  assign n29715 = n4221 & n29714 ;
  assign n29716 = n29715 ^ n26127 ^ 1'b0 ;
  assign n29717 = ~n1448 & n7906 ;
  assign n29718 = n29717 ^ n11610 ^ n7419 ;
  assign n29719 = n11110 & ~n29718 ;
  assign n29720 = n5008 ^ n3887 ^ 1'b0 ;
  assign n29721 = n29719 & ~n29720 ;
  assign n29722 = n17526 & ~n26241 ;
  assign n29723 = ( n468 & n748 ) | ( n468 & n1583 ) | ( n748 & n1583 ) ;
  assign n29724 = ( n777 & n9751 ) | ( n777 & n29723 ) | ( n9751 & n29723 ) ;
  assign n29725 = ( n9310 & ~n16687 ) | ( n9310 & n29724 ) | ( ~n16687 & n29724 ) ;
  assign n29726 = n3382 & ~n23464 ;
  assign n29727 = ( n5499 & ~n15522 ) | ( n5499 & n20673 ) | ( ~n15522 & n20673 ) ;
  assign n29728 = n29727 ^ n17111 ^ 1'b0 ;
  assign n29729 = n18614 ^ n15361 ^ n1260 ;
  assign n29730 = n4522 ^ n2521 ^ n1371 ;
  assign n29731 = ( n5140 & ~n14525 ) | ( n5140 & n29730 ) | ( ~n14525 & n29730 ) ;
  assign n29732 = ( n14227 & n23204 ) | ( n14227 & ~n29731 ) | ( n23204 & ~n29731 ) ;
  assign n29733 = n4629 | n10932 ;
  assign n29734 = n29733 ^ n12543 ^ 1'b0 ;
  assign n29735 = n18494 ^ n10993 ^ n3595 ;
  assign n29736 = n3141 | n29735 ;
  assign n29737 = n13315 ^ n8979 ^ n5909 ;
  assign n29738 = n21866 | n29737 ;
  assign n29739 = n29738 ^ x50 ^ 1'b0 ;
  assign n29740 = n2622 & ~n18316 ;
  assign n29741 = n1100 & n20583 ;
  assign n29742 = n7420 | n23127 ;
  assign n29743 = n3683 & n8182 ;
  assign n29744 = n7635 ^ n3904 ^ 1'b0 ;
  assign n29745 = ~n3044 & n10989 ;
  assign n29746 = n29745 ^ n5081 ^ 1'b0 ;
  assign n29747 = n29746 ^ n17113 ^ n5610 ;
  assign n29748 = ( ~n9656 & n29744 ) | ( ~n9656 & n29747 ) | ( n29744 & n29747 ) ;
  assign n29749 = ( n3406 & ~n7895 ) | ( n3406 & n29748 ) | ( ~n7895 & n29748 ) ;
  assign n29750 = ( n6918 & ~n9495 ) | ( n6918 & n17488 ) | ( ~n9495 & n17488 ) ;
  assign n29751 = ( n6384 & n20743 ) | ( n6384 & ~n29750 ) | ( n20743 & ~n29750 ) ;
  assign n29752 = n18892 ^ n4654 ^ 1'b0 ;
  assign n29753 = ~n27981 & n29752 ;
  assign n29755 = n16390 ^ n11611 ^ n4180 ;
  assign n29754 = ( n4239 & n5909 ) | ( n4239 & n7687 ) | ( n5909 & n7687 ) ;
  assign n29756 = n29755 ^ n29754 ^ 1'b0 ;
  assign n29757 = ~n6091 & n29756 ;
  assign n29758 = ~n4164 & n11613 ;
  assign n29759 = ~n14350 & n29758 ;
  assign n29760 = n29493 ^ n11080 ^ 1'b0 ;
  assign n29761 = ~n4002 & n29760 ;
  assign n29762 = n13896 ^ n10447 ^ n2767 ;
  assign n29763 = ~n8254 & n8837 ;
  assign n29764 = ~n29762 & n29763 ;
  assign n29765 = n15248 | n16004 ;
  assign n29766 = n29765 ^ n15375 ^ 1'b0 ;
  assign n29770 = ( n4643 & n5637 ) | ( n4643 & n6918 ) | ( n5637 & n6918 ) ;
  assign n29771 = ( ~n16743 & n24151 ) | ( ~n16743 & n29770 ) | ( n24151 & n29770 ) ;
  assign n29767 = ( ~n265 & n1901 ) | ( ~n265 & n2059 ) | ( n1901 & n2059 ) ;
  assign n29768 = n29767 ^ n6152 ^ n3113 ;
  assign n29769 = n29768 ^ n12402 ^ n11151 ;
  assign n29772 = n29771 ^ n29769 ^ n989 ;
  assign n29773 = ( n1660 & n7548 ) | ( n1660 & ~n10968 ) | ( n7548 & ~n10968 ) ;
  assign n29774 = n29773 ^ n15669 ^ n4895 ;
  assign n29775 = ( n18257 & n26006 ) | ( n18257 & ~n29774 ) | ( n26006 & ~n29774 ) ;
  assign n29776 = n29775 ^ n17683 ^ n2785 ;
  assign n29777 = ( n595 & n2622 ) | ( n595 & n4173 ) | ( n2622 & n4173 ) ;
  assign n29778 = n29777 ^ n28485 ^ n21498 ;
  assign n29779 = n8066 ^ n7140 ^ n6336 ;
  assign n29780 = n29779 ^ n19685 ^ 1'b0 ;
  assign n29781 = n18247 ^ n17535 ^ n2861 ;
  assign n29782 = n2163 ^ n1599 ^ 1'b0 ;
  assign n29783 = n7485 & n29782 ;
  assign n29784 = n10959 ^ n266 ^ 1'b0 ;
  assign n29785 = n29783 & ~n29784 ;
  assign n29786 = n10930 & ~n11216 ;
  assign n29787 = n1608 ^ n370 ^ 1'b0 ;
  assign n29789 = n5762 | n5780 ;
  assign n29788 = ~n17836 & n29737 ;
  assign n29790 = n29789 ^ n29788 ^ n5892 ;
  assign n29791 = n4748 & n23603 ;
  assign n29792 = n29791 ^ n5769 ^ n5456 ;
  assign n29793 = n17066 | n27427 ;
  assign n29794 = n28262 ^ n9172 ^ 1'b0 ;
  assign n29795 = n12707 ^ n2138 ^ 1'b0 ;
  assign n29796 = n9500 ^ n7225 ^ 1'b0 ;
  assign n29797 = n2489 | n29796 ;
  assign n29798 = n29797 ^ n14829 ^ 1'b0 ;
  assign n29799 = ( n4541 & ~n13367 ) | ( n4541 & n17539 ) | ( ~n13367 & n17539 ) ;
  assign n29800 = n29799 ^ n519 ^ 1'b0 ;
  assign n29801 = n15605 & n29800 ;
  assign n29802 = ( n8593 & n9622 ) | ( n8593 & ~n15233 ) | ( n9622 & ~n15233 ) ;
  assign n29803 = n16158 ^ n1266 ^ 1'b0 ;
  assign n29804 = n29802 & ~n29803 ;
  assign n29805 = n2374 | n10953 ;
  assign n29806 = n9148 | n29805 ;
  assign n29807 = n1284 & ~n9779 ;
  assign n29808 = n29807 ^ n6083 ^ 1'b0 ;
  assign n29809 = n16397 ^ n6156 ^ n2446 ;
  assign n29810 = n16938 ^ n15361 ^ n3349 ;
  assign n29811 = n29810 ^ n29349 ^ n20282 ;
  assign n29812 = n5395 ^ n1316 ^ 1'b0 ;
  assign n29813 = n21332 ^ n194 ^ 1'b0 ;
  assign n29814 = n9800 & n29813 ;
  assign n29815 = n29814 ^ n10970 ^ n2804 ;
  assign n29816 = n29815 ^ n23214 ^ n12344 ;
  assign n29817 = n369 & ~n4396 ;
  assign n29818 = ~n15052 & n29817 ;
  assign n29819 = ( n29812 & n29816 ) | ( n29812 & ~n29818 ) | ( n29816 & ~n29818 ) ;
  assign n29820 = n13379 ^ n10893 ^ n5824 ;
  assign n29821 = ~n637 & n29820 ;
  assign n29822 = ( n6024 & n19738 ) | ( n6024 & ~n29821 ) | ( n19738 & ~n29821 ) ;
  assign n29823 = ~n8350 & n22556 ;
  assign n29824 = ~n13267 & n29823 ;
  assign n29825 = n29824 ^ n29668 ^ n21787 ;
  assign n29826 = n29825 ^ n24198 ^ n3683 ;
  assign n29827 = n5716 & n15818 ;
  assign n29828 = ~n17173 & n29827 ;
  assign n29829 = n1774 & ~n12094 ;
  assign n29830 = n24952 ^ n4450 ^ 1'b0 ;
  assign n29832 = n15125 ^ n3108 ^ 1'b0 ;
  assign n29833 = n1956 | n29832 ;
  assign n29834 = n11913 & ~n29833 ;
  assign n29835 = ~n3636 & n29834 ;
  assign n29831 = ~n4957 & n20992 ;
  assign n29836 = n29835 ^ n29831 ^ 1'b0 ;
  assign n29837 = n8925 ^ n2205 ^ 1'b0 ;
  assign n29838 = n5306 & ~n20466 ;
  assign n29839 = n29837 & n29838 ;
  assign n29840 = n10000 & ~n29839 ;
  assign n29841 = ~n8164 & n29840 ;
  assign n29844 = n5215 ^ n5009 ^ 1'b0 ;
  assign n29845 = n7671 | n29844 ;
  assign n29843 = ~n5648 & n8466 ;
  assign n29846 = n29845 ^ n29843 ^ 1'b0 ;
  assign n29842 = n18055 ^ n18015 ^ n15397 ;
  assign n29847 = n29846 ^ n29842 ^ n326 ;
  assign n29848 = ( n229 & n1196 ) | ( n229 & ~n10415 ) | ( n1196 & ~n10415 ) ;
  assign n29849 = ( ~n10291 & n18219 ) | ( ~n10291 & n29848 ) | ( n18219 & n29848 ) ;
  assign n29850 = n6437 & ~n29849 ;
  assign n29851 = n29850 ^ n9115 ^ 1'b0 ;
  assign n29852 = n29851 ^ n22963 ^ n17528 ;
  assign n29853 = n29852 ^ n9305 ^ 1'b0 ;
  assign n29854 = n16341 ^ n13004 ^ 1'b0 ;
  assign n29855 = n24835 ^ n12255 ^ 1'b0 ;
  assign n29856 = n25535 ^ n6038 ^ n4110 ;
  assign n29857 = ( ~n4011 & n10174 ) | ( ~n4011 & n29856 ) | ( n10174 & n29856 ) ;
  assign n29858 = n21210 ^ n3395 ^ n1788 ;
  assign n29859 = n639 | n25807 ;
  assign n29860 = n29859 ^ n15758 ^ 1'b0 ;
  assign n29861 = n25549 ^ n21695 ^ 1'b0 ;
  assign n29862 = n21020 & n29861 ;
  assign n29863 = n3014 & ~n4546 ;
  assign n29864 = n2252 & n29863 ;
  assign n29865 = n25696 ^ n9701 ^ 1'b0 ;
  assign n29866 = ~n14749 & n29865 ;
  assign n29867 = n26075 & n29802 ;
  assign n29868 = n21147 ^ n8413 ^ 1'b0 ;
  assign n29869 = ( ~n21937 & n24770 ) | ( ~n21937 & n29868 ) | ( n24770 & n29868 ) ;
  assign n29874 = ( ~n1618 & n9519 ) | ( ~n1618 & n12793 ) | ( n9519 & n12793 ) ;
  assign n29875 = ( n9651 & n10902 ) | ( n9651 & n29874 ) | ( n10902 & n29874 ) ;
  assign n29870 = n2014 & n2551 ;
  assign n29871 = n29870 ^ n6673 ^ 1'b0 ;
  assign n29872 = ( n2303 & n6638 ) | ( n2303 & ~n29505 ) | ( n6638 & ~n29505 ) ;
  assign n29873 = ( n19304 & ~n29871 ) | ( n19304 & n29872 ) | ( ~n29871 & n29872 ) ;
  assign n29876 = n29875 ^ n29873 ^ n8184 ;
  assign n29877 = ( ~n2016 & n17319 ) | ( ~n2016 & n26829 ) | ( n17319 & n26829 ) ;
  assign n29878 = n29877 ^ n197 ^ 1'b0 ;
  assign n29879 = ( ~n14402 & n15068 ) | ( ~n14402 & n17591 ) | ( n15068 & n17591 ) ;
  assign n29880 = n10748 ^ n3927 ^ 1'b0 ;
  assign n29881 = n22956 & ~n29880 ;
  assign n29882 = n29774 ^ n7298 ^ 1'b0 ;
  assign n29883 = n16421 & n29882 ;
  assign n29884 = n15807 ^ n2871 ^ 1'b0 ;
  assign n29885 = n6311 & n6783 ;
  assign n29886 = n29885 ^ n2277 ^ 1'b0 ;
  assign n29887 = n29886 ^ n4508 ^ 1'b0 ;
  assign n29888 = ~n2388 & n25272 ;
  assign n29889 = n26821 & ~n29888 ;
  assign n29890 = n5034 & ~n7884 ;
  assign n29891 = ( ~n2724 & n4148 ) | ( ~n2724 & n29890 ) | ( n4148 & n29890 ) ;
  assign n29892 = n9577 & ~n29891 ;
  assign n29893 = ( n8870 & n9371 ) | ( n8870 & ~n16239 ) | ( n9371 & ~n16239 ) ;
  assign n29894 = n29893 ^ n26625 ^ n8058 ;
  assign n29895 = n18709 ^ n4306 ^ 1'b0 ;
  assign n29896 = n25386 ^ n13994 ^ n13402 ;
  assign n29897 = ( n13811 & n29895 ) | ( n13811 & n29896 ) | ( n29895 & n29896 ) ;
  assign n29898 = n13827 ^ n7601 ^ n468 ;
  assign n29899 = n29898 ^ n12861 ^ n8921 ;
  assign n29900 = n29899 ^ n3589 ^ 1'b0 ;
  assign n29901 = ( n2428 & n7418 ) | ( n2428 & ~n14690 ) | ( n7418 & ~n14690 ) ;
  assign n29902 = n24928 & n29901 ;
  assign n29903 = n11586 & ~n14140 ;
  assign n29904 = n25736 & n29903 ;
  assign n29905 = n3197 & ~n4996 ;
  assign n29906 = n29905 ^ n3773 ^ 1'b0 ;
  assign n29907 = n3267 & ~n16835 ;
  assign n29908 = n24488 & n29907 ;
  assign n29909 = ( n23192 & ~n29906 ) | ( n23192 & n29908 ) | ( ~n29906 & n29908 ) ;
  assign n29910 = ( n11540 & n23588 ) | ( n11540 & ~n29909 ) | ( n23588 & ~n29909 ) ;
  assign n29911 = ~n8613 & n19711 ;
  assign n29912 = n29910 & n29911 ;
  assign n29913 = ( n3729 & n10441 ) | ( n3729 & ~n16477 ) | ( n10441 & ~n16477 ) ;
  assign n29914 = n29913 ^ n29254 ^ n17929 ;
  assign n29915 = n1600 & n6083 ;
  assign n29916 = ~n27315 & n29915 ;
  assign n29917 = n29442 | n29916 ;
  assign n29918 = ( n11260 & n13571 ) | ( n11260 & ~n15029 ) | ( n13571 & ~n15029 ) ;
  assign n29919 = ( ~n6845 & n11992 ) | ( ~n6845 & n24099 ) | ( n11992 & n24099 ) ;
  assign n29920 = n27129 ^ n8034 ^ n7785 ;
  assign n29923 = ~n895 & n16084 ;
  assign n29921 = n11185 & n16756 ;
  assign n29922 = n29921 ^ n10093 ^ n4002 ;
  assign n29924 = n29923 ^ n29922 ^ n21577 ;
  assign n29925 = n29924 ^ n23752 ^ n16002 ;
  assign n29926 = n28817 ^ n24954 ^ n1310 ;
  assign n29927 = n1724 & ~n29926 ;
  assign n29928 = n7276 & n29927 ;
  assign n29929 = ( n3231 & n7272 ) | ( n3231 & ~n14293 ) | ( n7272 & ~n14293 ) ;
  assign n29930 = n2718 | n9195 ;
  assign n29931 = n7806 | n29930 ;
  assign n29932 = n29929 | n29931 ;
  assign n29933 = n5979 ^ n2906 ^ 1'b0 ;
  assign n29934 = ~n1240 & n6924 ;
  assign n29935 = n29934 ^ n13886 ^ 1'b0 ;
  assign n29938 = n17876 ^ n12408 ^ 1'b0 ;
  assign n29936 = ~n17420 & n25791 ;
  assign n29937 = n29936 ^ n11281 ^ 1'b0 ;
  assign n29939 = n29938 ^ n29937 ^ n16146 ;
  assign n29941 = n134 | n3517 ;
  assign n29942 = n9881 & ~n29941 ;
  assign n29940 = n2342 | n16281 ;
  assign n29943 = n29942 ^ n29940 ^ 1'b0 ;
  assign n29944 = ( ~n14045 & n24091 ) | ( ~n14045 & n29943 ) | ( n24091 & n29943 ) ;
  assign n29945 = ~n12881 & n14478 ;
  assign n29946 = n29945 ^ n15792 ^ 1'b0 ;
  assign n29947 = ( n13493 & n19765 ) | ( n13493 & n29946 ) | ( n19765 & n29946 ) ;
  assign n29952 = n625 | n15767 ;
  assign n29953 = n25879 & ~n29952 ;
  assign n29948 = ( n649 & n692 ) | ( n649 & n3311 ) | ( n692 & n3311 ) ;
  assign n29949 = n17534 ^ n14821 ^ n11722 ;
  assign n29950 = n29949 ^ n16779 ^ 1'b0 ;
  assign n29951 = n29948 | n29950 ;
  assign n29954 = n29953 ^ n29951 ^ n19685 ;
  assign n29955 = n16835 ^ n10735 ^ n829 ;
  assign n29956 = ( n17381 & n23183 ) | ( n17381 & n25780 ) | ( n23183 & n25780 ) ;
  assign n29957 = n2433 & n21161 ;
  assign n29958 = n3605 | n21746 ;
  assign n29959 = n11673 & ~n29958 ;
  assign n29960 = n20001 & ~n29959 ;
  assign n29961 = n14269 ^ n4374 ^ 1'b0 ;
  assign n29962 = ~n11630 & n29961 ;
  assign n29963 = n11759 ^ n6990 ^ 1'b0 ;
  assign n29964 = n6297 ^ n4717 ^ 1'b0 ;
  assign n29969 = n5302 ^ n4460 ^ 1'b0 ;
  assign n29970 = n5162 & ~n29969 ;
  assign n29971 = n29970 ^ n5806 ^ n3821 ;
  assign n29972 = n1619 & ~n21972 ;
  assign n29973 = n29972 ^ n5628 ^ 1'b0 ;
  assign n29974 = ( n16660 & n29971 ) | ( n16660 & ~n29973 ) | ( n29971 & ~n29973 ) ;
  assign n29965 = ( n10301 & ~n15406 ) | ( n10301 & n23668 ) | ( ~n15406 & n23668 ) ;
  assign n29966 = n29965 ^ n12459 ^ 1'b0 ;
  assign n29967 = n22737 ^ n11500 ^ 1'b0 ;
  assign n29968 = n29966 & ~n29967 ;
  assign n29975 = n29974 ^ n29968 ^ n25356 ;
  assign n29976 = ( ~n6223 & n11237 ) | ( ~n6223 & n19468 ) | ( n11237 & n19468 ) ;
  assign n29977 = n19853 | n23941 ;
  assign n29978 = n29977 ^ n1186 ^ 1'b0 ;
  assign n29979 = n29978 ^ n10871 ^ n2940 ;
  assign n29981 = ~n5653 & n11066 ;
  assign n29982 = n29981 ^ n7104 ^ 1'b0 ;
  assign n29980 = n26292 ^ n3721 ^ 1'b0 ;
  assign n29983 = n29982 ^ n29980 ^ n23732 ;
  assign n29984 = n659 & ~n12861 ;
  assign n29985 = n13969 & ~n16192 ;
  assign n29986 = n4056 & ~n9852 ;
  assign n29987 = ~n29985 & n29986 ;
  assign n29988 = ~n1192 & n1332 ;
  assign n29989 = n6226 & n29988 ;
  assign n29990 = ( n5969 & n12539 ) | ( n5969 & n18088 ) | ( n12539 & n18088 ) ;
  assign n29991 = n18252 | n29990 ;
  assign n29992 = ~n12991 & n25194 ;
  assign n29993 = n29991 & n29992 ;
  assign n29994 = n2417 & n8555 ;
  assign n29995 = n13201 ^ n13069 ^ n5833 ;
  assign n29996 = n9403 ^ n229 ^ 1'b0 ;
  assign n29997 = ~n5098 & n29996 ;
  assign n29998 = ( n2978 & n12935 ) | ( n2978 & n29997 ) | ( n12935 & n29997 ) ;
  assign n29999 = ( ~n13881 & n26071 ) | ( ~n13881 & n29373 ) | ( n26071 & n29373 ) ;
  assign n30000 = n12474 ^ n5981 ^ n2803 ;
  assign n30001 = n26425 ^ n16557 ^ n10835 ;
  assign n30002 = n30001 ^ n11716 ^ n3729 ;
  assign n30003 = n11096 ^ n6352 ^ 1'b0 ;
  assign n30004 = n3254 | n30003 ;
  assign n30005 = n13174 & ~n30004 ;
  assign n30006 = n6774 ^ n3836 ^ 1'b0 ;
  assign n30007 = n10555 | n30006 ;
  assign n30008 = n18008 ^ n1473 ^ 1'b0 ;
  assign n30009 = n8934 & n30008 ;
  assign n30010 = n30009 ^ n10948 ^ n5371 ;
  assign n30011 = n15526 | n30010 ;
  assign n30012 = n8056 & ~n30011 ;
  assign n30013 = ( ~x15 & n11512 ) | ( ~x15 & n18586 ) | ( n11512 & n18586 ) ;
  assign n30014 = n2696 & ~n30013 ;
  assign n30015 = n30014 ^ n2112 ^ 1'b0 ;
  assign n30016 = n2884 & ~n5751 ;
  assign n30017 = n30016 ^ n8013 ^ 1'b0 ;
  assign n30018 = ( ~n14483 & n21181 ) | ( ~n14483 & n30017 ) | ( n21181 & n30017 ) ;
  assign n30019 = ( n7884 & ~n17965 ) | ( n7884 & n30018 ) | ( ~n17965 & n30018 ) ;
  assign n30020 = ( n1583 & n3687 ) | ( n1583 & ~n18551 ) | ( n3687 & ~n18551 ) ;
  assign n30021 = n10884 ^ n6073 ^ 1'b0 ;
  assign n30022 = ~n11496 & n30021 ;
  assign n30023 = n30022 ^ n4527 ^ 1'b0 ;
  assign n30024 = n14811 & n30023 ;
  assign n30025 = n7670 & ~n11359 ;
  assign n30026 = n18026 ^ n12731 ^ 1'b0 ;
  assign n30027 = ( n30024 & n30025 ) | ( n30024 & n30026 ) | ( n30025 & n30026 ) ;
  assign n30028 = n27627 ^ n16577 ^ n3602 ;
  assign n30029 = n10750 ^ n9087 ^ 1'b0 ;
  assign n30030 = ( n863 & ~n18940 ) | ( n863 & n30029 ) | ( ~n18940 & n30029 ) ;
  assign n30031 = ~n16712 & n29227 ;
  assign n30032 = n7263 | n12188 ;
  assign n30033 = n30032 ^ n11867 ^ 1'b0 ;
  assign n30034 = n30033 ^ n8491 ^ 1'b0 ;
  assign n30035 = n10195 ^ n7575 ^ 1'b0 ;
  assign n30036 = ~n30034 & n30035 ;
  assign n30037 = n24265 ^ n3877 ^ n145 ;
  assign n30038 = ( ~n537 & n15854 ) | ( ~n537 & n26493 ) | ( n15854 & n26493 ) ;
  assign n30042 = n2668 | n4396 ;
  assign n30043 = n4268 | n30042 ;
  assign n30039 = n16940 & n24195 ;
  assign n30040 = n30039 ^ n6827 ^ 1'b0 ;
  assign n30041 = ~n3995 & n30040 ;
  assign n30044 = n30043 ^ n30041 ^ n13747 ;
  assign n30045 = ( ~n7893 & n14591 ) | ( ~n7893 & n23199 ) | ( n14591 & n23199 ) ;
  assign n30046 = ( n7065 & n22487 ) | ( n7065 & ~n30045 ) | ( n22487 & ~n30045 ) ;
  assign n30047 = n21975 ^ n4415 ^ n529 ;
  assign n30048 = ( n4454 & ~n24799 ) | ( n4454 & n30047 ) | ( ~n24799 & n30047 ) ;
  assign n30049 = n29922 | n30048 ;
  assign n30050 = n4404 ^ n305 ^ 1'b0 ;
  assign n30051 = n1862 & n30050 ;
  assign n30052 = n30051 ^ n11583 ^ 1'b0 ;
  assign n30053 = n11582 | n13869 ;
  assign n30054 = n30053 ^ n6477 ^ 1'b0 ;
  assign n30055 = n4484 | n30054 ;
  assign n30056 = n18076 | n30055 ;
  assign n30057 = n11331 | n22996 ;
  assign n30058 = n17067 | n30057 ;
  assign n30059 = n14870 ^ n7083 ^ 1'b0 ;
  assign n30060 = n5168 | n30059 ;
  assign n30061 = n21558 ^ n5412 ^ 1'b0 ;
  assign n30062 = n20755 ^ n2900 ^ 1'b0 ;
  assign n30063 = ~n5009 & n8437 ;
  assign n30068 = n10359 ^ n696 ^ 1'b0 ;
  assign n30069 = n11096 & n30068 ;
  assign n30065 = n23186 ^ n5849 ^ n1066 ;
  assign n30064 = n9854 | n13312 ;
  assign n30066 = n30065 ^ n30064 ^ 1'b0 ;
  assign n30067 = ( ~n407 & n5522 ) | ( ~n407 & n30066 ) | ( n5522 & n30066 ) ;
  assign n30070 = n30069 ^ n30067 ^ n3068 ;
  assign n30071 = ( n4949 & ~n9367 ) | ( n4949 & n23127 ) | ( ~n9367 & n23127 ) ;
  assign n30072 = ~n2421 & n2716 ;
  assign n30073 = n30072 ^ n5716 ^ 1'b0 ;
  assign n30074 = n16830 | n17558 ;
  assign n30075 = n20114 | n30074 ;
  assign n30076 = ( n23451 & n30073 ) | ( n23451 & n30075 ) | ( n30073 & n30075 ) ;
  assign n30077 = n20649 | n30076 ;
  assign n30078 = n4475 | n7059 ;
  assign n30079 = n30078 ^ n14111 ^ 1'b0 ;
  assign n30080 = n17295 ^ n13836 ^ 1'b0 ;
  assign n30081 = n17035 & n30080 ;
  assign n30082 = ( ~n1656 & n5720 ) | ( ~n1656 & n21653 ) | ( n5720 & n21653 ) ;
  assign n30084 = n11013 | n17080 ;
  assign n30085 = n30084 ^ n15141 ^ 1'b0 ;
  assign n30086 = n30085 ^ n14034 ^ n6867 ;
  assign n30083 = n17213 ^ n13079 ^ n1011 ;
  assign n30087 = n30086 ^ n30083 ^ 1'b0 ;
  assign n30090 = n16846 | n25275 ;
  assign n30088 = n3385 | n16081 ;
  assign n30089 = n605 | n30088 ;
  assign n30091 = n30090 ^ n30089 ^ n23355 ;
  assign n30092 = ( n2200 & n13616 ) | ( n2200 & n17025 ) | ( n13616 & n17025 ) ;
  assign n30093 = ( n4840 & n25569 ) | ( n4840 & n30092 ) | ( n25569 & n30092 ) ;
  assign n30094 = n4542 | n15888 ;
  assign n30095 = n11594 & ~n30094 ;
  assign n30096 = n20203 & n28859 ;
  assign n30097 = n30095 & n30096 ;
  assign n30098 = n8754 ^ n7907 ^ n5843 ;
  assign n30099 = n25609 & ~n30098 ;
  assign n30100 = n30099 ^ n15318 ^ 1'b0 ;
  assign n30101 = n30100 ^ n4405 ^ 1'b0 ;
  assign n30102 = n11401 ^ n2710 ^ 1'b0 ;
  assign n30103 = n22726 & ~n30102 ;
  assign n30104 = n2294 & n11266 ;
  assign n30105 = ~n3362 & n30104 ;
  assign n30106 = ~x115 & n30105 ;
  assign n30107 = n8377 ^ n6871 ^ n4139 ;
  assign n30108 = n26629 ^ n15051 ^ n10630 ;
  assign n30109 = n14178 ^ n4723 ^ n2744 ;
  assign n30110 = ~n2369 & n5313 ;
  assign n30111 = n24814 ^ n10124 ^ n5539 ;
  assign n30112 = ( n5546 & ~n6015 ) | ( n5546 & n9923 ) | ( ~n6015 & n9923 ) ;
  assign n30113 = n30112 ^ n28518 ^ n17164 ;
  assign n30114 = ( n25784 & n30111 ) | ( n25784 & n30113 ) | ( n30111 & n30113 ) ;
  assign n30115 = ( ~n500 & n3603 ) | ( ~n500 & n30114 ) | ( n3603 & n30114 ) ;
  assign n30116 = ( ~n10191 & n14722 ) | ( ~n10191 & n29322 ) | ( n14722 & n29322 ) ;
  assign n30117 = n12804 & n30116 ;
  assign n30118 = n22376 ^ n11108 ^ 1'b0 ;
  assign n30119 = ~n28040 & n30118 ;
  assign n30120 = ( n1498 & ~n6183 ) | ( n1498 & n29948 ) | ( ~n6183 & n29948 ) ;
  assign n30121 = ~n14991 & n24515 ;
  assign n30122 = n30120 & n30121 ;
  assign n30123 = ~n22408 & n24798 ;
  assign n30124 = n30122 & n30123 ;
  assign n30125 = n24386 ^ n22491 ^ n10223 ;
  assign n30126 = n4224 & n30125 ;
  assign n30127 = ( n5225 & n18637 ) | ( n5225 & n24033 ) | ( n18637 & n24033 ) ;
  assign n30129 = n19674 ^ n15140 ^ 1'b0 ;
  assign n30130 = ~n6593 & n30129 ;
  assign n30128 = n9713 ^ n5466 ^ 1'b0 ;
  assign n30131 = n30130 ^ n30128 ^ n25965 ;
  assign n30132 = n15854 ^ n6174 ^ 1'b0 ;
  assign n30133 = x87 & n30132 ;
  assign n30134 = n4906 | n10386 ;
  assign n30135 = n30133 | n30134 ;
  assign n30136 = n30135 ^ n17111 ^ n12598 ;
  assign n30137 = ( n5491 & n19063 ) | ( n5491 & n26223 ) | ( n19063 & n26223 ) ;
  assign n30138 = n29189 ^ n11068 ^ n2753 ;
  assign n30139 = n30138 ^ n11548 ^ n2282 ;
  assign n30140 = n13143 ^ n10367 ^ n3821 ;
  assign n30141 = n16358 ^ n7502 ^ 1'b0 ;
  assign n30142 = n30140 & ~n30141 ;
  assign n30143 = ~n7730 & n21823 ;
  assign n30144 = ~n6975 & n30143 ;
  assign n30145 = n13650 ^ n7202 ^ n2185 ;
  assign n30146 = n25549 & n25935 ;
  assign n30147 = n30146 ^ n16773 ^ 1'b0 ;
  assign n30148 = ( n23594 & n30145 ) | ( n23594 & n30147 ) | ( n30145 & n30147 ) ;
  assign n30149 = ( n2741 & ~n4234 ) | ( n2741 & n5587 ) | ( ~n4234 & n5587 ) ;
  assign n30150 = n28732 ^ n17177 ^ n15051 ;
  assign n30151 = n30150 ^ n11718 ^ n8985 ;
  assign n30152 = n2493 & ~n9465 ;
  assign n30154 = n6677 ^ n4776 ^ 1'b0 ;
  assign n30153 = n5083 & ~n6690 ;
  assign n30155 = n30154 ^ n30153 ^ n24153 ;
  assign n30156 = n15360 ^ n10656 ^ 1'b0 ;
  assign n30157 = ( n5619 & ~n26873 ) | ( n5619 & n30156 ) | ( ~n26873 & n30156 ) ;
  assign n30158 = n5299 & n30157 ;
  assign n30159 = n25891 ^ n14679 ^ n10698 ;
  assign n30160 = n7436 & ~n20377 ;
  assign n30161 = n30159 & n30160 ;
  assign n30162 = n20426 ^ n18016 ^ 1'b0 ;
  assign n30163 = n17119 ^ n1750 ^ 1'b0 ;
  assign n30164 = n26283 ^ n12447 ^ n7891 ;
  assign n30165 = ( n7843 & ~n23986 ) | ( n7843 & n30164 ) | ( ~n23986 & n30164 ) ;
  assign n30166 = ~n4946 & n8398 ;
  assign n30167 = ~n3140 & n30166 ;
  assign n30168 = n24515 ^ n9687 ^ 1'b0 ;
  assign n30169 = n16128 ^ n9079 ^ 1'b0 ;
  assign n30170 = ( n2417 & n7054 ) | ( n2417 & n27817 ) | ( n7054 & n27817 ) ;
  assign n30171 = n2227 & n13928 ;
  assign n30172 = ( n644 & n7071 ) | ( n644 & n30171 ) | ( n7071 & n30171 ) ;
  assign n30173 = n14529 ^ n9233 ^ 1'b0 ;
  assign n30174 = n30172 | n30173 ;
  assign n30175 = n14808 & n30174 ;
  assign n30176 = n23281 ^ n16446 ^ 1'b0 ;
  assign n30177 = n9676 | n10234 ;
  assign n30178 = n25813 | n30177 ;
  assign n30179 = n22271 ^ n12852 ^ 1'b0 ;
  assign n30180 = n16417 & ~n30179 ;
  assign n30181 = n30180 ^ n7624 ^ 1'b0 ;
  assign n30182 = ~n22479 & n30181 ;
  assign n30183 = n10201 | n18571 ;
  assign n30184 = n3836 | n17038 ;
  assign n30185 = n30184 ^ n8369 ^ 1'b0 ;
  assign n30186 = x93 | n4700 ;
  assign n30187 = ~n3785 & n9134 ;
  assign n30188 = n30187 ^ n3566 ^ 1'b0 ;
  assign n30189 = n30188 ^ n11594 ^ n3757 ;
  assign n30191 = n15562 ^ n15205 ^ 1'b0 ;
  assign n30190 = n9225 & n19073 ;
  assign n30192 = n30191 ^ n30190 ^ 1'b0 ;
  assign n30193 = n19853 ^ n17848 ^ n4688 ;
  assign n30194 = ~n30192 & n30193 ;
  assign n30195 = ( n21787 & ~n30189 ) | ( n21787 & n30194 ) | ( ~n30189 & n30194 ) ;
  assign n30196 = n10293 ^ n9847 ^ n3988 ;
  assign n30197 = n5231 ^ n3768 ^ 1'b0 ;
  assign n30198 = n545 & ~n2374 ;
  assign n30199 = ~n30197 & n30198 ;
  assign n30200 = ( ~n22890 & n30196 ) | ( ~n22890 & n30199 ) | ( n30196 & n30199 ) ;
  assign n30201 = ( n2603 & n26363 ) | ( n2603 & n29737 ) | ( n26363 & n29737 ) ;
  assign n30202 = n11193 ^ n1343 ^ 1'b0 ;
  assign n30203 = n6248 | n30202 ;
  assign n30204 = ( n7082 & n11332 ) | ( n7082 & n15203 ) | ( n11332 & n15203 ) ;
  assign n30205 = n30204 ^ n23669 ^ n11335 ;
  assign n30206 = n12444 & ~n30205 ;
  assign n30207 = n30206 ^ n14901 ^ 1'b0 ;
  assign n30208 = ( n9071 & n30203 ) | ( n9071 & ~n30207 ) | ( n30203 & ~n30207 ) ;
  assign n30209 = ( n4006 & n7236 ) | ( n4006 & n18534 ) | ( n7236 & n18534 ) ;
  assign n30210 = n30060 & n30209 ;
  assign n30211 = n1899 | n25082 ;
  assign n30212 = ( ~n1700 & n4260 ) | ( ~n1700 & n5868 ) | ( n4260 & n5868 ) ;
  assign n30213 = n21948 & ~n30212 ;
  assign n30214 = ~n16892 & n17462 ;
  assign n30215 = n15034 & n30214 ;
  assign n30216 = n26787 ^ n12416 ^ 1'b0 ;
  assign n30217 = n21450 | n30216 ;
  assign n30218 = n23746 ^ n18104 ^ 1'b0 ;
  assign n30219 = ( n913 & n8450 ) | ( n913 & ~n27589 ) | ( n8450 & ~n27589 ) ;
  assign n30220 = ( n2190 & n4016 ) | ( n2190 & n5780 ) | ( n4016 & n5780 ) ;
  assign n30221 = ( n2429 & n21857 ) | ( n2429 & n30220 ) | ( n21857 & n30220 ) ;
  assign n30222 = n25044 ^ n13881 ^ n3599 ;
  assign n30223 = n6379 ^ n5762 ^ n3760 ;
  assign n30224 = n30223 ^ n10948 ^ n5186 ;
  assign n30225 = n7624 & ~n25746 ;
  assign n30226 = n20615 & n30225 ;
  assign n30230 = n4184 & n7541 ;
  assign n30231 = n30230 ^ n14574 ^ 1'b0 ;
  assign n30232 = n30231 ^ n28116 ^ 1'b0 ;
  assign n30233 = n2190 & n30232 ;
  assign n30234 = ( n850 & n15273 ) | ( n850 & n30233 ) | ( n15273 & n30233 ) ;
  assign n30227 = ~n1465 & n5025 ;
  assign n30228 = n14290 & n30227 ;
  assign n30229 = n6111 | n30228 ;
  assign n30235 = n30234 ^ n30229 ^ 1'b0 ;
  assign n30236 = n27432 ^ n3829 ^ 1'b0 ;
  assign n30237 = n11440 ^ n8052 ^ n4778 ;
  assign n30238 = ( n12465 & n20470 ) | ( n12465 & n30237 ) | ( n20470 & n30237 ) ;
  assign n30239 = ( n16697 & n27490 ) | ( n16697 & ~n30238 ) | ( n27490 & ~n30238 ) ;
  assign n30240 = n13649 & ~n25402 ;
  assign n30241 = ~x95 & n30240 ;
  assign n30242 = n30241 ^ n13524 ^ 1'b0 ;
  assign n30243 = n30242 ^ n19659 ^ 1'b0 ;
  assign n30245 = n4545 & ~n5569 ;
  assign n30246 = n30245 ^ n6464 ^ 1'b0 ;
  assign n30244 = ( n1835 & n5051 ) | ( n1835 & n9259 ) | ( n5051 & n9259 ) ;
  assign n30247 = n30246 ^ n30244 ^ n15494 ;
  assign n30248 = n21522 ^ n17528 ^ 1'b0 ;
  assign n30249 = n8473 | n9065 ;
  assign n30250 = ~n5985 & n30249 ;
  assign n30251 = n30250 ^ n16001 ^ 1'b0 ;
  assign n30252 = ( n23509 & n26404 ) | ( n23509 & n27305 ) | ( n26404 & n27305 ) ;
  assign n30253 = n30252 ^ n28292 ^ 1'b0 ;
  assign n30254 = n3257 & n5277 ;
  assign n30255 = n30254 ^ n12196 ^ 1'b0 ;
  assign n30256 = n1078 & ~n9255 ;
  assign n30257 = n30256 ^ n1687 ^ 1'b0 ;
  assign n30258 = n4621 | n11247 ;
  assign n30259 = n30257 | n30258 ;
  assign n30261 = n16813 ^ n8992 ^ n8505 ;
  assign n30260 = n6154 | n19521 ;
  assign n30262 = n30261 ^ n30260 ^ 1'b0 ;
  assign n30263 = n30262 ^ n19385 ^ 1'b0 ;
  assign n30264 = n30259 & ~n30263 ;
  assign n30265 = n4765 ^ n2433 ^ n2361 ;
  assign n30266 = n13541 & n30265 ;
  assign n30267 = n30266 ^ n4298 ^ 1'b0 ;
  assign n30268 = n10448 & ~n30267 ;
  assign n30269 = n5165 ^ n409 ^ 1'b0 ;
  assign n30270 = n30268 & n30269 ;
  assign n30271 = n6418 | n13345 ;
  assign n30272 = n22766 ^ n10597 ^ n5177 ;
  assign n30273 = n30272 ^ n14224 ^ 1'b0 ;
  assign n30274 = ~n20976 & n30051 ;
  assign n30275 = n30274 ^ n19475 ^ n2706 ;
  assign n30276 = ( n2062 & n17054 ) | ( n2062 & ~n23240 ) | ( n17054 & ~n23240 ) ;
  assign n30277 = n16712 | n30276 ;
  assign n30278 = n4498 | n30277 ;
  assign n30279 = n5700 & n30278 ;
  assign n30282 = ( n248 & n3352 ) | ( n248 & ~n10832 ) | ( n3352 & ~n10832 ) ;
  assign n30280 = n27193 ^ n7937 ^ 1'b0 ;
  assign n30281 = n7187 & n30280 ;
  assign n30283 = n30282 ^ n30281 ^ n13212 ;
  assign n30284 = n18836 ^ n11246 ^ n4429 ;
  assign n30285 = n30284 ^ n21853 ^ n10902 ;
  assign n30286 = ~n5655 & n17149 ;
  assign n30287 = n30286 ^ n1226 ^ 1'b0 ;
  assign n30290 = n10145 ^ n2323 ^ 1'b0 ;
  assign n30289 = ~n17351 & n29752 ;
  assign n30291 = n30290 ^ n30289 ^ 1'b0 ;
  assign n30292 = n30291 ^ n16662 ^ n397 ;
  assign n30288 = ~n3167 & n27869 ;
  assign n30293 = n30292 ^ n30288 ^ 1'b0 ;
  assign n30294 = n24977 | n30293 ;
  assign n30295 = n30294 ^ n3035 ^ 1'b0 ;
  assign n30296 = n9231 & n14118 ;
  assign n30297 = n30296 ^ n7585 ^ 1'b0 ;
  assign n30298 = ( n1901 & n13071 ) | ( n1901 & n19379 ) | ( n13071 & n19379 ) ;
  assign n30299 = n30298 ^ n12268 ^ 1'b0 ;
  assign n30300 = n21630 ^ n19885 ^ n19804 ;
  assign n30301 = n6496 & n9744 ;
  assign n30302 = ~n25621 & n30301 ;
  assign n30303 = ( n7676 & n16840 ) | ( n7676 & ~n22488 ) | ( n16840 & ~n22488 ) ;
  assign n30304 = n3768 & ~n9871 ;
  assign n30305 = n6887 ^ n3569 ^ 1'b0 ;
  assign n30306 = ( n24434 & ~n30304 ) | ( n24434 & n30305 ) | ( ~n30304 & n30305 ) ;
  assign n30307 = n30306 ^ n8211 ^ n5259 ;
  assign n30309 = n4488 & ~n15233 ;
  assign n30308 = ~n4028 & n16494 ;
  assign n30310 = n30309 ^ n30308 ^ 1'b0 ;
  assign n30311 = n6752 & ~n17547 ;
  assign n30312 = n30311 ^ n13856 ^ 1'b0 ;
  assign n30313 = ~n3956 & n21790 ;
  assign n30314 = n30313 ^ n16988 ^ 1'b0 ;
  assign n30315 = n29966 ^ n18265 ^ 1'b0 ;
  assign n30316 = n7695 ^ n3805 ^ n266 ;
  assign n30317 = n15216 | n30316 ;
  assign n30318 = n30317 ^ n28211 ^ 1'b0 ;
  assign n30319 = n30318 ^ n15913 ^ n1225 ;
  assign n30320 = x108 & ~n2040 ;
  assign n30321 = ~n4522 & n30320 ;
  assign n30322 = n30321 ^ n15815 ^ 1'b0 ;
  assign n30323 = ~n24669 & n27427 ;
  assign n30324 = n19523 ^ n13164 ^ n9332 ;
  assign n30325 = n19142 ^ n2011 ^ 1'b0 ;
  assign n30326 = n3349 & ~n6867 ;
  assign n30327 = ~n733 & n30326 ;
  assign n30328 = n30327 ^ n19653 ^ 1'b0 ;
  assign n30329 = n30325 & n30328 ;
  assign n30330 = ~n25218 & n25292 ;
  assign n30331 = x72 & n11273 ;
  assign n30332 = n17491 ^ n12865 ^ 1'b0 ;
  assign n30335 = n1857 & n13851 ;
  assign n30336 = ~n9162 & n30335 ;
  assign n30333 = n11616 ^ n2112 ^ n250 ;
  assign n30334 = ( x126 & ~n1465 ) | ( x126 & n30333 ) | ( ~n1465 & n30333 ) ;
  assign n30337 = n30336 ^ n30334 ^ n2863 ;
  assign n30338 = n23992 ^ n6462 ^ 1'b0 ;
  assign n30339 = n20879 ^ n18838 ^ 1'b0 ;
  assign n30341 = n20551 ^ n15580 ^ 1'b0 ;
  assign n30340 = n5558 | n26163 ;
  assign n30342 = n30341 ^ n30340 ^ n12931 ;
  assign n30344 = n7152 | n11679 ;
  assign n30345 = n12674 & ~n30344 ;
  assign n30343 = n6489 & ~n24726 ;
  assign n30346 = n30345 ^ n30343 ^ n1194 ;
  assign n30347 = ( n3992 & ~n9226 ) | ( n3992 & n10114 ) | ( ~n9226 & n10114 ) ;
  assign n30348 = n30347 ^ n19950 ^ n11832 ;
  assign n30350 = n22296 ^ n13518 ^ n1422 ;
  assign n30349 = ~n2499 & n21156 ;
  assign n30351 = n30350 ^ n30349 ^ 1'b0 ;
  assign n30352 = ~n9368 & n29997 ;
  assign n30353 = ~n28645 & n30352 ;
  assign n30354 = ( n4151 & n6504 ) | ( n4151 & ~n13353 ) | ( n6504 & ~n13353 ) ;
  assign n30355 = n30354 ^ n5001 ^ 1'b0 ;
  assign n30356 = ~n19308 & n30355 ;
  assign n30357 = n11995 & ~n15473 ;
  assign n30358 = n30357 ^ n23329 ^ 1'b0 ;
  assign n30359 = ( n10439 & n18145 ) | ( n10439 & n30358 ) | ( n18145 & n30358 ) ;
  assign n30360 = n8390 & n20442 ;
  assign n30361 = ~n26436 & n30360 ;
  assign n30362 = ~n14863 & n25717 ;
  assign n30363 = n30361 & n30362 ;
  assign n30364 = n30363 ^ n26803 ^ n19036 ;
  assign n30365 = n26610 ^ n20776 ^ n15332 ;
  assign n30366 = ( n13621 & ~n28193 ) | ( n13621 & n28629 ) | ( ~n28193 & n28629 ) ;
  assign n30367 = n24201 & n29491 ;
  assign n30368 = n14504 & n30367 ;
  assign n30369 = n9588 | n30368 ;
  assign n30370 = n29491 ^ n22194 ^ n3286 ;
  assign n30371 = ( ~n4161 & n13994 ) | ( ~n4161 & n23725 ) | ( n13994 & n23725 ) ;
  assign n30372 = n23732 ^ n10207 ^ n1220 ;
  assign n30373 = n11956 & n24631 ;
  assign n30374 = ( n7511 & ~n29088 ) | ( n7511 & n30373 ) | ( ~n29088 & n30373 ) ;
  assign n30375 = n10575 | n11754 ;
  assign n30376 = n30375 ^ n20251 ^ 1'b0 ;
  assign n30377 = n4357 & ~n12421 ;
  assign n30378 = n30376 & ~n30377 ;
  assign n30379 = ( n847 & ~n8851 ) | ( n847 & n15332 ) | ( ~n8851 & n15332 ) ;
  assign n30380 = n3015 & ~n6226 ;
  assign n30381 = n30379 & n30380 ;
  assign n30382 = n14464 | n20446 ;
  assign n30383 = n30382 ^ n14046 ^ 1'b0 ;
  assign n30384 = ~n1100 & n4859 ;
  assign n30385 = n18568 ^ n15447 ^ n4238 ;
  assign n30386 = ( n15855 & n19045 ) | ( n15855 & n19685 ) | ( n19045 & n19685 ) ;
  assign n30387 = ~n3756 & n5780 ;
  assign n30388 = ( n13212 & ~n30119 ) | ( n13212 & n30387 ) | ( ~n30119 & n30387 ) ;
  assign n30389 = n22881 ^ n10873 ^ 1'b0 ;
  assign n30390 = n129 & ~n29692 ;
  assign n30391 = n30390 ^ n4386 ^ 1'b0 ;
  assign n30392 = ~n4765 & n30391 ;
  assign n30393 = ~n17044 & n29365 ;
  assign n30394 = n13362 ^ n3456 ^ 1'b0 ;
  assign n30395 = n2793 | n6382 ;
  assign n30396 = n10854 & ~n30395 ;
  assign n30397 = n10982 ^ n2103 ^ 1'b0 ;
  assign n30398 = n405 & n30397 ;
  assign n30399 = ( ~n2593 & n6545 ) | ( ~n2593 & n9779 ) | ( n6545 & n9779 ) ;
  assign n30400 = n30399 ^ n14472 ^ n10890 ;
  assign n30401 = n2544 & ~n17115 ;
  assign n30402 = ( n2694 & n28341 ) | ( n2694 & ~n30401 ) | ( n28341 & ~n30401 ) ;
  assign n30403 = n30402 ^ n25437 ^ n8859 ;
  assign n30404 = ( ~n12403 & n14826 ) | ( ~n12403 & n30403 ) | ( n14826 & n30403 ) ;
  assign n30405 = n10903 ^ n9177 ^ 1'b0 ;
  assign n30406 = n17641 ^ n14903 ^ n2431 ;
  assign n30407 = n13321 & n27361 ;
  assign n30408 = n7750 | n19556 ;
  assign n30409 = n30408 ^ n2108 ^ 1'b0 ;
  assign n30410 = n6262 ^ n3965 ^ 1'b0 ;
  assign n30411 = n5786 & ~n10706 ;
  assign n30412 = n30411 ^ n18490 ^ 1'b0 ;
  assign n30413 = n30412 ^ n22172 ^ 1'b0 ;
  assign n30414 = n30410 & ~n30413 ;
  assign n30415 = n27299 ^ n21858 ^ n3838 ;
  assign n30416 = n27979 ^ n16645 ^ n5722 ;
  assign n30417 = ( n21435 & ~n21998 ) | ( n21435 & n30416 ) | ( ~n21998 & n30416 ) ;
  assign n30418 = n18015 | n30417 ;
  assign n30419 = ( n20354 & n23221 ) | ( n20354 & n28215 ) | ( n23221 & n28215 ) ;
  assign n30420 = n15210 & ~n18577 ;
  assign n30421 = ( ~n3956 & n22510 ) | ( ~n3956 & n30420 ) | ( n22510 & n30420 ) ;
  assign n30422 = n30333 ^ n26548 ^ n5438 ;
  assign n30423 = ( n8521 & n10625 ) | ( n8521 & ~n11164 ) | ( n10625 & ~n11164 ) ;
  assign n30424 = ~n4985 & n8764 ;
  assign n30425 = n16326 & ~n30424 ;
  assign n30426 = n9800 & n11938 ;
  assign n30427 = ( n2197 & n2545 ) | ( n2197 & n3734 ) | ( n2545 & n3734 ) ;
  assign n30428 = n30427 ^ n6289 ^ n3982 ;
  assign n30429 = n1362 & ~n7754 ;
  assign n30430 = n30428 & n30429 ;
  assign n30431 = ( n10040 & n23495 ) | ( n10040 & ~n30430 ) | ( n23495 & ~n30430 ) ;
  assign n30432 = n17042 & n30431 ;
  assign n30433 = n30432 ^ n15852 ^ 1'b0 ;
  assign n30434 = n526 & ~n9935 ;
  assign n30435 = n30434 ^ n6089 ^ 1'b0 ;
  assign n30436 = n4130 & n30435 ;
  assign n30437 = ~n1522 & n30436 ;
  assign n30438 = n24053 | n30437 ;
  assign n30439 = n22182 ^ n12208 ^ 1'b0 ;
  assign n30440 = ~n30438 & n30439 ;
  assign n30441 = ( n10505 & ~n25508 ) | ( n10505 & n27023 ) | ( ~n25508 & n27023 ) ;
  assign n30442 = ( x19 & n1504 ) | ( x19 & n15433 ) | ( n1504 & n15433 ) ;
  assign n30443 = n2331 & ~n2862 ;
  assign n30444 = n8528 ^ n6699 ^ n5341 ;
  assign n30445 = n20304 ^ n9712 ^ 1'b0 ;
  assign n30446 = n28556 & n30445 ;
  assign n30447 = n16261 & n30446 ;
  assign n30450 = ( n1669 & ~n5039 ) | ( n1669 & n6456 ) | ( ~n5039 & n6456 ) ;
  assign n30448 = ( n3113 & ~n5782 ) | ( n3113 & n6793 ) | ( ~n5782 & n6793 ) ;
  assign n30449 = n7363 & n30448 ;
  assign n30451 = n30450 ^ n30449 ^ 1'b0 ;
  assign n30452 = n19636 ^ n18312 ^ n17024 ;
  assign n30453 = n7874 & ~n23711 ;
  assign n30454 = ~n30452 & n30453 ;
  assign n30457 = n15647 ^ n5015 ^ n1511 ;
  assign n30458 = n30457 ^ n17131 ^ n13146 ;
  assign n30455 = ~n5139 & n8391 ;
  assign n30456 = n30455 ^ n28907 ^ 1'b0 ;
  assign n30459 = n30458 ^ n30456 ^ n8604 ;
  assign n30460 = n23491 ^ n9347 ^ n1894 ;
  assign n30461 = ( ~n1818 & n5146 ) | ( ~n1818 & n23477 ) | ( n5146 & n23477 ) ;
  assign n30462 = n30461 ^ n26709 ^ n18908 ;
  assign n30463 = ( n5096 & n9046 ) | ( n5096 & n19167 ) | ( n9046 & n19167 ) ;
  assign n30464 = ( n16319 & ~n16687 ) | ( n16319 & n30463 ) | ( ~n16687 & n30463 ) ;
  assign n30465 = n30464 ^ n10577 ^ n3063 ;
  assign n30466 = n5230 & ~n22510 ;
  assign n30467 = n1882 & n30466 ;
  assign n30468 = ( n254 & ~n1677 ) | ( n254 & n11772 ) | ( ~n1677 & n11772 ) ;
  assign n30469 = n30119 & n30468 ;
  assign n30470 = n30469 ^ n28215 ^ 1'b0 ;
  assign n30471 = n3203 & ~n24735 ;
  assign n30472 = n30471 ^ n2701 ^ 1'b0 ;
  assign n30473 = n13203 | n24733 ;
  assign n30474 = ~n20447 & n30473 ;
  assign n30475 = ~n22448 & n23491 ;
  assign n30476 = n30475 ^ n3029 ^ 1'b0 ;
  assign n30477 = n9504 & n12109 ;
  assign n30478 = ( ~n5454 & n18397 ) | ( ~n5454 & n30477 ) | ( n18397 & n30477 ) ;
  assign n30482 = x95 & ~n3979 ;
  assign n30483 = n30482 ^ n948 ^ 1'b0 ;
  assign n30484 = ~n7859 & n30483 ;
  assign n30485 = n17444 ^ n10072 ^ 1'b0 ;
  assign n30486 = n30484 | n30485 ;
  assign n30479 = n8491 ^ n5583 ^ 1'b0 ;
  assign n30480 = n3934 & n30479 ;
  assign n30481 = n30480 ^ n767 ^ 1'b0 ;
  assign n30487 = n30486 ^ n30481 ^ n17883 ;
  assign n30488 = n1619 & n22360 ;
  assign n30489 = n30488 ^ n4960 ^ 1'b0 ;
  assign n30490 = n30489 ^ n21399 ^ n8814 ;
  assign n30491 = n29190 ^ n26830 ^ n26073 ;
  assign n30492 = n13737 ^ n3739 ^ 1'b0 ;
  assign n30493 = ( n18099 & ~n18867 ) | ( n18099 & n30492 ) | ( ~n18867 & n30492 ) ;
  assign n30494 = n19564 ^ n8360 ^ 1'b0 ;
  assign n30495 = ~n12480 & n30494 ;
  assign n30496 = n30495 ^ n24096 ^ n19817 ;
  assign n30497 = n10944 & ~n30496 ;
  assign n30498 = ~n3194 & n10225 ;
  assign n30499 = n5419 | n19859 ;
  assign n30500 = ~n30498 & n30499 ;
  assign n30501 = n24454 ^ n15453 ^ 1'b0 ;
  assign n30502 = n26032 ^ n24957 ^ n297 ;
  assign n30503 = n12715 & n26571 ;
  assign n30504 = n11703 ^ n11540 ^ n975 ;
  assign n30505 = ( ~n15982 & n20710 ) | ( ~n15982 & n23189 ) | ( n20710 & n23189 ) ;
  assign n30506 = n30505 ^ n26987 ^ n1384 ;
  assign n30507 = ( n6053 & n6138 ) | ( n6053 & n10690 ) | ( n6138 & n10690 ) ;
  assign n30508 = n2546 & n30507 ;
  assign n30509 = n2674 & n30508 ;
  assign n30510 = n30509 ^ n20989 ^ 1'b0 ;
  assign n30511 = n1829 | n13920 ;
  assign n30512 = n12441 | n30511 ;
  assign n30513 = ( ~n16045 & n25162 ) | ( ~n16045 & n30477 ) | ( n25162 & n30477 ) ;
  assign n30514 = n9355 ^ n1129 ^ 1'b0 ;
  assign n30515 = n8450 & ~n30514 ;
  assign n30516 = n30515 ^ n18624 ^ n16597 ;
  assign n30517 = n1664 ^ n1113 ^ 1'b0 ;
  assign n30518 = n30517 ^ n18555 ^ 1'b0 ;
  assign n30519 = n30518 ^ n25230 ^ n20031 ;
  assign n30520 = n8557 ^ n5295 ^ 1'b0 ;
  assign n30521 = ( n369 & n19124 ) | ( n369 & n30520 ) | ( n19124 & n30520 ) ;
  assign n30522 = ( n1996 & n3593 ) | ( n1996 & n8223 ) | ( n3593 & n8223 ) ;
  assign n30523 = n12603 ^ n5278 ^ 1'b0 ;
  assign n30524 = n30522 & ~n30523 ;
  assign n30525 = ( n9490 & n21078 ) | ( n9490 & n30524 ) | ( n21078 & n30524 ) ;
  assign n30526 = n17735 | n28001 ;
  assign n30527 = n5456 & ~n17174 ;
  assign n30528 = ~n16772 & n30527 ;
  assign n30529 = n17091 ^ n16667 ^ 1'b0 ;
  assign n30530 = n9260 & ~n30529 ;
  assign n30531 = n21226 ^ n14105 ^ 1'b0 ;
  assign n30532 = x5 & ~n30531 ;
  assign n30533 = n17578 ^ n3686 ^ 1'b0 ;
  assign n30534 = n16723 & n19460 ;
  assign n30535 = n30533 & n30534 ;
  assign n30536 = ( n6320 & n19229 ) | ( n6320 & n22805 ) | ( n19229 & n22805 ) ;
  assign n30537 = n27842 ^ n24442 ^ n19604 ;
  assign n30538 = n13478 ^ n7403 ^ 1'b0 ;
  assign n30539 = n30538 ^ n13801 ^ n12297 ;
  assign n30540 = ( n14344 & ~n21543 ) | ( n14344 & n30539 ) | ( ~n21543 & n30539 ) ;
  assign n30541 = ( n3835 & ~n10273 ) | ( n3835 & n11084 ) | ( ~n10273 & n11084 ) ;
  assign n30542 = ~n15025 & n23289 ;
  assign n30543 = n13616 ^ n11547 ^ 1'b0 ;
  assign n30544 = n6095 | n30543 ;
  assign n30545 = n13345 | n28535 ;
  assign n30546 = n22114 | n30545 ;
  assign n30547 = n27348 ^ n24694 ^ n20222 ;
  assign n30548 = n20157 ^ n10662 ^ 1'b0 ;
  assign n30549 = n5725 | n30548 ;
  assign n30550 = ( n30546 & n30547 ) | ( n30546 & n30549 ) | ( n30547 & n30549 ) ;
  assign n30551 = n30550 ^ n2485 ^ 1'b0 ;
  assign n30552 = n5818 | n7142 ;
  assign n30553 = n7642 ^ n4976 ^ n3937 ;
  assign n30554 = n30553 ^ n18518 ^ n18077 ;
  assign n30555 = n30554 ^ n426 ^ 1'b0 ;
  assign n30556 = n30552 | n30555 ;
  assign n30557 = ~n12944 & n15437 ;
  assign n30558 = ( ~n1510 & n9348 ) | ( ~n1510 & n16397 ) | ( n9348 & n16397 ) ;
  assign n30559 = n20557 ^ n20349 ^ n13297 ;
  assign n30560 = n3338 ^ n1971 ^ 1'b0 ;
  assign n30561 = ( n6855 & n15665 ) | ( n6855 & ~n30560 ) | ( n15665 & ~n30560 ) ;
  assign n30562 = n28456 ^ n11653 ^ x120 ;
  assign n30563 = n8715 & n20044 ;
  assign n30564 = n11265 ^ n5989 ^ 1'b0 ;
  assign n30565 = n3934 & ~n30564 ;
  assign n30566 = n30565 ^ n1600 ^ 1'b0 ;
  assign n30567 = n24571 & n30566 ;
  assign n30568 = n14879 ^ n13539 ^ 1'b0 ;
  assign n30569 = n1865 & n30568 ;
  assign n30571 = n6822 ^ n4273 ^ 1'b0 ;
  assign n30570 = ~n3019 & n9629 ;
  assign n30572 = n30571 ^ n30570 ^ 1'b0 ;
  assign n30573 = n3381 & ~n19655 ;
  assign n30574 = ( ~n3204 & n9941 ) | ( ~n3204 & n18961 ) | ( n9941 & n18961 ) ;
  assign n30575 = n3768 & ~n30574 ;
  assign n30576 = n30477 ^ n8584 ^ 1'b0 ;
  assign n30577 = n30575 & n30576 ;
  assign n30578 = n22129 ^ n11315 ^ 1'b0 ;
  assign n30579 = ( n916 & n8946 ) | ( n916 & n30578 ) | ( n8946 & n30578 ) ;
  assign n30580 = n30029 ^ n11691 ^ 1'b0 ;
  assign n30581 = n8442 & n30580 ;
  assign n30582 = n17766 & n30581 ;
  assign n30583 = n30579 & n30582 ;
  assign n30584 = n30577 & n30583 ;
  assign n30585 = ( n7130 & n11684 ) | ( n7130 & n13848 ) | ( n11684 & n13848 ) ;
  assign n30586 = ( n8822 & n22774 ) | ( n8822 & n30585 ) | ( n22774 & n30585 ) ;
  assign n30587 = n20592 ^ n14061 ^ n4973 ;
  assign n30588 = n30587 ^ n7482 ^ 1'b0 ;
  assign n30589 = ( n14334 & ~n21196 ) | ( n14334 & n30588 ) | ( ~n21196 & n30588 ) ;
  assign n30591 = n17947 & ~n26174 ;
  assign n30590 = n14893 | n19939 ;
  assign n30592 = n30591 ^ n30590 ^ 1'b0 ;
  assign n30593 = n6243 & n9467 ;
  assign n30594 = n30593 ^ n3424 ^ 1'b0 ;
  assign n30595 = n593 | n12766 ;
  assign n30596 = n24568 & ~n30595 ;
  assign n30597 = ( n11633 & n12666 ) | ( n11633 & ~n18278 ) | ( n12666 & ~n18278 ) ;
  assign n30598 = n30597 ^ n13366 ^ n7512 ;
  assign n30599 = n22904 ^ n13894 ^ 1'b0 ;
  assign n30600 = n30599 ^ n14838 ^ n11983 ;
  assign n30601 = n30600 ^ n8699 ^ 1'b0 ;
  assign n30602 = n29464 ^ n22403 ^ n11003 ;
  assign n30603 = n25823 ^ n189 ^ 1'b0 ;
  assign n30604 = n12009 ^ n5232 ^ 1'b0 ;
  assign n30606 = ( ~x66 & n6204 ) | ( ~x66 & n11158 ) | ( n6204 & n11158 ) ;
  assign n30605 = ( ~n4036 & n7979 ) | ( ~n4036 & n23586 ) | ( n7979 & n23586 ) ;
  assign n30607 = n30606 ^ n30605 ^ n4407 ;
  assign n30608 = n3514 | n4876 ;
  assign n30609 = n30608 ^ n24486 ^ 1'b0 ;
  assign n30613 = n903 & n4753 ;
  assign n30610 = n13965 ^ n11146 ^ 1'b0 ;
  assign n30611 = n11643 | n30610 ;
  assign n30612 = n1796 & ~n30611 ;
  assign n30614 = n30613 ^ n30612 ^ 1'b0 ;
  assign n30615 = n4932 | n18163 ;
  assign n30616 = n30615 ^ n21758 ^ 1'b0 ;
  assign n30617 = n12969 ^ n9114 ^ n6571 ;
  assign n30618 = n30617 ^ n30376 ^ 1'b0 ;
  assign n30619 = x80 & n30618 ;
  assign n30620 = n4939 ^ n1927 ^ n203 ;
  assign n30621 = ( ~n297 & n6492 ) | ( ~n297 & n30620 ) | ( n6492 & n30620 ) ;
  assign n30622 = n30621 ^ n3853 ^ 1'b0 ;
  assign n30623 = n2229 & n30622 ;
  assign n30624 = n30623 ^ n20163 ^ n15487 ;
  assign n30625 = n30624 ^ n22947 ^ n17134 ;
  assign n30626 = ( ~n6435 & n6687 ) | ( ~n6435 & n12018 ) | ( n6687 & n12018 ) ;
  assign n30627 = n30626 ^ n11013 ^ 1'b0 ;
  assign n30628 = ( n2612 & ~n3352 ) | ( n2612 & n8258 ) | ( ~n3352 & n8258 ) ;
  assign n30629 = ( n8835 & ~n18262 ) | ( n8835 & n30628 ) | ( ~n18262 & n30628 ) ;
  assign n30630 = n20700 ^ n9287 ^ n3110 ;
  assign n30631 = n3410 & ~n23261 ;
  assign n30632 = ~n29345 & n30631 ;
  assign n30633 = ( ~n1452 & n27503 ) | ( ~n1452 & n30632 ) | ( n27503 & n30632 ) ;
  assign n30634 = n961 & ~n10125 ;
  assign n30635 = n30634 ^ n27985 ^ 1'b0 ;
  assign n30636 = ( n12181 & n13327 ) | ( n12181 & ~n28945 ) | ( n13327 & ~n28945 ) ;
  assign n30638 = n8335 | n13663 ;
  assign n30639 = n20709 | n30638 ;
  assign n30637 = n24884 ^ n9782 ^ n2898 ;
  assign n30640 = n30639 ^ n30637 ^ n18547 ;
  assign n30641 = ( n394 & ~n18680 ) | ( n394 & n25458 ) | ( ~n18680 & n25458 ) ;
  assign n30642 = ( ~n7231 & n10994 ) | ( ~n7231 & n19236 ) | ( n10994 & n19236 ) ;
  assign n30643 = ( n14119 & ~n15690 ) | ( n14119 & n16509 ) | ( ~n15690 & n16509 ) ;
  assign n30644 = n16960 ^ n3507 ^ n953 ;
  assign n30645 = n18526 & ~n30644 ;
  assign n30646 = n3985 & n30645 ;
  assign n30647 = n12512 ^ n8035 ^ n4443 ;
  assign n30648 = ~n28541 & n30647 ;
  assign n30649 = n30648 ^ n6413 ^ 1'b0 ;
  assign n30650 = ~n16508 & n30086 ;
  assign n30651 = n3836 & n30650 ;
  assign n30652 = n18367 ^ n18044 ^ n17809 ;
  assign n30653 = ~n1388 & n2904 ;
  assign n30654 = n24940 ^ n6328 ^ 1'b0 ;
  assign n30655 = n30620 ^ n21881 ^ n16803 ;
  assign n30656 = n30655 ^ n6855 ^ n5527 ;
  assign n30657 = n30076 & n30656 ;
  assign n30658 = ( n8012 & n12747 ) | ( n8012 & ~n14525 ) | ( n12747 & ~n14525 ) ;
  assign n30659 = n3349 ^ n3288 ^ n197 ;
  assign n30660 = ~n9867 & n11086 ;
  assign n30661 = ~n16915 & n30660 ;
  assign n30662 = n9501 & ~n15088 ;
  assign n30663 = ~n28006 & n30662 ;
  assign n30664 = n20484 ^ n10040 ^ 1'b0 ;
  assign n30665 = ~n11801 & n30664 ;
  assign n30666 = ~n9296 & n30665 ;
  assign n30667 = n2653 | n5724 ;
  assign n30668 = n30667 ^ n17878 ^ 1'b0 ;
  assign n30669 = ( x66 & ~n1603 ) | ( x66 & n15016 ) | ( ~n1603 & n15016 ) ;
  assign n30670 = ( n1890 & ~n21791 ) | ( n1890 & n26571 ) | ( ~n21791 & n26571 ) ;
  assign n30671 = ( n8710 & ~n14928 ) | ( n8710 & n30670 ) | ( ~n14928 & n30670 ) ;
  assign n30674 = ( n2163 & n5240 ) | ( n2163 & n9403 ) | ( n5240 & n9403 ) ;
  assign n30675 = n23952 & n30674 ;
  assign n30676 = n30675 ^ n11892 ^ 1'b0 ;
  assign n30677 = ~n6363 & n30676 ;
  assign n30672 = n3843 & n6742 ;
  assign n30673 = n30672 ^ n15778 ^ 1'b0 ;
  assign n30678 = n30677 ^ n30673 ^ n15386 ;
  assign n30679 = n7588 ^ n2948 ^ 1'b0 ;
  assign n30680 = n16259 & n30679 ;
  assign n30681 = ( ~n759 & n20249 ) | ( ~n759 & n30680 ) | ( n20249 & n30680 ) ;
  assign n30682 = ( n10769 & n11836 ) | ( n10769 & n16287 ) | ( n11836 & n16287 ) ;
  assign n30683 = n13676 | n30682 ;
  assign n30684 = ~n1916 & n15784 ;
  assign n30685 = ~n11688 & n30684 ;
  assign n30686 = n14080 ^ n12817 ^ 1'b0 ;
  assign n30687 = n14652 & ~n30686 ;
  assign n30688 = n7838 ^ n7331 ^ n2421 ;
  assign n30691 = ~n12419 & n26160 ;
  assign n30692 = n30691 ^ n21275 ^ 1'b0 ;
  assign n30689 = n7863 | n11144 ;
  assign n30690 = n5482 & ~n30689 ;
  assign n30693 = n30692 ^ n30690 ^ 1'b0 ;
  assign n30694 = n2169 & ~n21662 ;
  assign n30695 = n30694 ^ n8201 ^ 1'b0 ;
  assign n30696 = ~n576 & n11387 ;
  assign n30697 = n30696 ^ n29143 ^ 1'b0 ;
  assign n30698 = ( n3977 & n4700 ) | ( n3977 & n30697 ) | ( n4700 & n30697 ) ;
  assign n30699 = ( n2008 & n2112 ) | ( n2008 & n26337 ) | ( n2112 & n26337 ) ;
  assign n30700 = ( n17123 & n19429 ) | ( n17123 & n30699 ) | ( n19429 & n30699 ) ;
  assign n30701 = n15703 & ~n30700 ;
  assign n30702 = n17721 ^ n7073 ^ 1'b0 ;
  assign n30703 = n25049 & ~n30702 ;
  assign n30704 = n8527 & n30703 ;
  assign n30705 = ~n7343 & n14774 ;
  assign n30706 = n30705 ^ n17094 ^ 1'b0 ;
  assign n30707 = ( ~n5622 & n16837 ) | ( ~n5622 & n30706 ) | ( n16837 & n30706 ) ;
  assign n30708 = ( n3817 & n9543 ) | ( n3817 & n10704 ) | ( n9543 & n10704 ) ;
  assign n30709 = ( ~n3231 & n7113 ) | ( ~n3231 & n30708 ) | ( n7113 & n30708 ) ;
  assign n30710 = ( n8277 & n18264 ) | ( n8277 & ~n21384 ) | ( n18264 & ~n21384 ) ;
  assign n30711 = x72 & n3644 ;
  assign n30712 = n30711 ^ n2475 ^ 1'b0 ;
  assign n30713 = n20320 ^ n4949 ^ 1'b0 ;
  assign n30714 = n23578 & n30713 ;
  assign n30715 = n28612 ^ n14318 ^ 1'b0 ;
  assign n30716 = ~n17560 & n30715 ;
  assign n30717 = ( n3551 & n7337 ) | ( n3551 & n15241 ) | ( n7337 & n15241 ) ;
  assign n30718 = n30717 ^ n4401 ^ n3912 ;
  assign n30719 = ( n16614 & ~n17988 ) | ( n16614 & n30718 ) | ( ~n17988 & n30718 ) ;
  assign n30720 = n15740 ^ n12225 ^ 1'b0 ;
  assign n30721 = n8459 ^ n6093 ^ 1'b0 ;
  assign n30722 = n17146 ^ n2273 ^ 1'b0 ;
  assign n30723 = n4429 | n30722 ;
  assign n30724 = ( ~n24841 & n30721 ) | ( ~n24841 & n30723 ) | ( n30721 & n30723 ) ;
  assign n30725 = n30724 ^ n14352 ^ n7347 ;
  assign n30726 = n30725 ^ n26448 ^ n24244 ;
  assign n30727 = ( ~n7288 & n18652 ) | ( ~n7288 & n26036 ) | ( n18652 & n26036 ) ;
  assign n30728 = ( n464 & n7108 ) | ( n464 & n29503 ) | ( n7108 & n29503 ) ;
  assign n30729 = n30728 ^ n19543 ^ n17856 ;
  assign n30730 = n12707 ^ n4509 ^ n4231 ;
  assign n30731 = ( n2276 & n8422 ) | ( n2276 & ~n12712 ) | ( n8422 & ~n12712 ) ;
  assign n30732 = n30731 ^ n19328 ^ 1'b0 ;
  assign n30733 = n30730 & n30732 ;
  assign n30734 = ( n1422 & n7236 ) | ( n1422 & ~n8674 ) | ( n7236 & ~n8674 ) ;
  assign n30735 = n14665 & n30734 ;
  assign n30736 = n10016 | n30735 ;
  assign n30737 = n11271 & n18260 ;
  assign n30738 = n30737 ^ n6881 ^ 1'b0 ;
  assign n30739 = n3820 & n8878 ;
  assign n30740 = n16875 ^ n10291 ^ 1'b0 ;
  assign n30741 = n30739 & n30740 ;
  assign n30742 = n10857 & n14196 ;
  assign n30743 = n30742 ^ n21239 ^ 1'b0 ;
  assign n30744 = n1227 | n3762 ;
  assign n30745 = n30744 ^ n9910 ^ 1'b0 ;
  assign n30746 = n4282 & n10344 ;
  assign n30747 = ~n10344 & n30746 ;
  assign n30748 = ( ~n383 & n9901 ) | ( ~n383 & n30747 ) | ( n9901 & n30747 ) ;
  assign n30749 = ( n3311 & ~n25907 ) | ( n3311 & n30748 ) | ( ~n25907 & n30748 ) ;
  assign n30750 = ( n28134 & ~n30745 ) | ( n28134 & n30749 ) | ( ~n30745 & n30749 ) ;
  assign n30751 = n17158 ^ n826 ^ 1'b0 ;
  assign n30752 = n19631 ^ n15726 ^ 1'b0 ;
  assign n30753 = n12322 ^ n7890 ^ n5134 ;
  assign n30754 = n30753 ^ n15547 ^ 1'b0 ;
  assign n30755 = n1408 & n30754 ;
  assign n30756 = n30755 ^ x26 ^ 1'b0 ;
  assign n30757 = n8919 | n19998 ;
  assign n30760 = n1790 & n20567 ;
  assign n30761 = ~n9683 & n30760 ;
  assign n30762 = n30761 ^ n9958 ^ 1'b0 ;
  assign n30758 = n13900 ^ n4796 ^ 1'b0 ;
  assign n30759 = n18709 & ~n30758 ;
  assign n30763 = n30762 ^ n30759 ^ n3369 ;
  assign n30764 = n7640 ^ n2434 ^ 1'b0 ;
  assign n30765 = n17311 ^ n14683 ^ 1'b0 ;
  assign n30766 = n3727 & n30765 ;
  assign n30767 = n9036 & n11372 ;
  assign n30768 = ~n6272 & n30767 ;
  assign n30769 = n27107 ^ n3838 ^ 1'b0 ;
  assign n30770 = n30768 | n30769 ;
  assign n30771 = n6696 | n20781 ;
  assign n30772 = n10117 & ~n30771 ;
  assign n30773 = n9291 ^ n7708 ^ 1'b0 ;
  assign n30774 = ~n15684 & n30773 ;
  assign n30775 = n30774 ^ n27913 ^ n5167 ;
  assign n30776 = ( x92 & ~n16504 ) | ( x92 & n18981 ) | ( ~n16504 & n18981 ) ;
  assign n30778 = ~n4306 & n9259 ;
  assign n30777 = n2844 | n7463 ;
  assign n30779 = n30778 ^ n30777 ^ 1'b0 ;
  assign n30780 = n30779 ^ n5353 ^ n4932 ;
  assign n30781 = n30776 & ~n30780 ;
  assign n30782 = n20369 ^ n17039 ^ 1'b0 ;
  assign n30783 = n17027 ^ n3644 ^ 1'b0 ;
  assign n30784 = ( n177 & n11630 ) | ( n177 & ~n30783 ) | ( n11630 & ~n30783 ) ;
  assign n30785 = n7884 ^ n2696 ^ 1'b0 ;
  assign n30786 = n26259 ^ n8177 ^ n7100 ;
  assign n30787 = n509 & ~n7614 ;
  assign n30788 = n30787 ^ n23739 ^ 1'b0 ;
  assign n30789 = ~n1650 & n22422 ;
  assign n30790 = ~n12857 & n30789 ;
  assign n30791 = n11738 & ~n30790 ;
  assign n30792 = n29227 | n30791 ;
  assign n30793 = n30792 ^ n11224 ^ 1'b0 ;
  assign n30794 = n4868 ^ x11 ^ 1'b0 ;
  assign n30795 = ~n1902 & n29202 ;
  assign n30798 = ~n17727 & n29602 ;
  assign n30799 = n12196 & n30798 ;
  assign n30796 = ~n2377 & n3011 ;
  assign n30797 = n30796 ^ n6620 ^ 1'b0 ;
  assign n30800 = n30799 ^ n30797 ^ n27169 ;
  assign n30801 = ~n2595 & n23733 ;
  assign n30802 = n30801 ^ n10813 ^ 1'b0 ;
  assign n30803 = n30800 | n30802 ;
  assign n30804 = ( n1830 & ~n4911 ) | ( n1830 & n12418 ) | ( ~n4911 & n12418 ) ;
  assign n30805 = ( n7606 & n12416 ) | ( n7606 & n14879 ) | ( n12416 & n14879 ) ;
  assign n30806 = n30805 ^ n18240 ^ n7205 ;
  assign n30807 = n30806 ^ n26759 ^ 1'b0 ;
  assign n30808 = ~n5139 & n5942 ;
  assign n30809 = n30808 ^ n1602 ^ 1'b0 ;
  assign n30810 = n14044 | n16845 ;
  assign n30811 = ( n21667 & n22467 ) | ( n21667 & n22826 ) | ( n22467 & n22826 ) ;
  assign n30812 = n30811 ^ n16486 ^ n1371 ;
  assign n30813 = ( n30809 & ~n30810 ) | ( n30809 & n30812 ) | ( ~n30810 & n30812 ) ;
  assign n30814 = n21673 ^ n6692 ^ 1'b0 ;
  assign n30815 = n6280 & ~n7502 ;
  assign n30816 = n30815 ^ n20047 ^ 1'b0 ;
  assign n30817 = n30816 ^ n20247 ^ n9974 ;
  assign n30818 = n24353 ^ n11480 ^ n5917 ;
  assign n30819 = n30818 ^ n29791 ^ n28685 ;
  assign n30821 = n6036 | n17936 ;
  assign n30820 = n2050 & ~n6578 ;
  assign n30822 = n30821 ^ n30820 ^ 1'b0 ;
  assign n30824 = n1880 & ~n4856 ;
  assign n30825 = n30824 ^ n7071 ^ n834 ;
  assign n30823 = ~n3029 & n12070 ;
  assign n30826 = n30825 ^ n30823 ^ 1'b0 ;
  assign n30827 = n3987 | n11457 ;
  assign n30828 = n6373 | n30827 ;
  assign n30829 = n3727 & ~n26810 ;
  assign n30830 = n30829 ^ n3530 ^ 1'b0 ;
  assign n30831 = n8607 ^ n2723 ^ n532 ;
  assign n30833 = n3910 & n4039 ;
  assign n30834 = n2072 & ~n30833 ;
  assign n30832 = n3289 & ~n15000 ;
  assign n30835 = n30834 ^ n30832 ^ n4627 ;
  assign n30836 = ( n4883 & n8216 ) | ( n4883 & n15626 ) | ( n8216 & n15626 ) ;
  assign n30837 = n28696 ^ n20564 ^ n7832 ;
  assign n30838 = n9975 ^ n4660 ^ n2685 ;
  assign n30839 = n720 & n30838 ;
  assign n30840 = n30839 ^ n9832 ^ 1'b0 ;
  assign n30841 = n30840 ^ n13780 ^ n12207 ;
  assign n30842 = n24814 ^ n22141 ^ n6158 ;
  assign n30843 = ~n2865 & n26977 ;
  assign n30844 = ~n26135 & n27924 ;
  assign n30845 = n30844 ^ n5137 ^ 1'b0 ;
  assign n30846 = n22953 ^ n10108 ^ x16 ;
  assign n30847 = n6004 ^ n2153 ^ 1'b0 ;
  assign n30848 = ~n10076 & n30847 ;
  assign n30849 = ( ~n10876 & n20793 ) | ( ~n10876 & n30848 ) | ( n20793 & n30848 ) ;
  assign n30850 = ( n1265 & n22152 ) | ( n1265 & n30849 ) | ( n22152 & n30849 ) ;
  assign n30851 = ( n2214 & n8918 ) | ( n2214 & n12987 ) | ( n8918 & n12987 ) ;
  assign n30852 = n26194 ^ n1606 ^ 1'b0 ;
  assign n30853 = ( n20742 & n27495 ) | ( n20742 & ~n30852 ) | ( n27495 & ~n30852 ) ;
  assign n30854 = ( ~n23482 & n25392 ) | ( ~n23482 & n30853 ) | ( n25392 & n30853 ) ;
  assign n30855 = ( ~n4107 & n15663 ) | ( ~n4107 & n21989 ) | ( n15663 & n21989 ) ;
  assign n30856 = ( n6403 & n15758 ) | ( n6403 & n22396 ) | ( n15758 & n22396 ) ;
  assign n30857 = ( n11738 & n15106 ) | ( n11738 & ~n15479 ) | ( n15106 & ~n15479 ) ;
  assign n30858 = n30857 ^ n15813 ^ n8604 ;
  assign n30859 = ( n26898 & n30856 ) | ( n26898 & n30858 ) | ( n30856 & n30858 ) ;
  assign n30860 = ( n14358 & ~n18699 ) | ( n14358 & n30859 ) | ( ~n18699 & n30859 ) ;
  assign n30861 = n1157 & n4076 ;
  assign n30862 = n3369 ^ n883 ^ 1'b0 ;
  assign n30863 = n9387 & n30862 ;
  assign n30864 = n17260 | n28759 ;
  assign n30865 = n16037 ^ n15580 ^ 1'b0 ;
  assign n30866 = ~n771 & n1852 ;
  assign n30867 = n10777 ^ n7090 ^ n4751 ;
  assign n30868 = n9173 & ~n30867 ;
  assign n30869 = ( n22822 & ~n25636 ) | ( n22822 & n30868 ) | ( ~n25636 & n30868 ) ;
  assign n30870 = ( n6425 & ~n25198 ) | ( n6425 & n30301 ) | ( ~n25198 & n30301 ) ;
  assign n30871 = ( n5277 & n13189 ) | ( n5277 & ~n30870 ) | ( n13189 & ~n30870 ) ;
  assign n30872 = n203 & ~n17493 ;
  assign n30873 = n27510 ^ n6778 ^ 1'b0 ;
  assign n30874 = n6539 | n24934 ;
  assign n30875 = n30874 ^ n13953 ^ 1'b0 ;
  assign n30876 = ( n3828 & n29192 ) | ( n3828 & n30875 ) | ( n29192 & n30875 ) ;
  assign n30877 = n6719 | n9778 ;
  assign n30878 = n5975 | n30877 ;
  assign n30879 = n5733 | n30878 ;
  assign n30880 = ( ~n2805 & n3405 ) | ( ~n2805 & n6671 ) | ( n3405 & n6671 ) ;
  assign n30881 = n6414 ^ n2711 ^ 1'b0 ;
  assign n30883 = n9414 | n12887 ;
  assign n30884 = ( ~n13908 & n25165 ) | ( ~n13908 & n30883 ) | ( n25165 & n30883 ) ;
  assign n30882 = n12365 & n25332 ;
  assign n30885 = n30884 ^ n30882 ^ 1'b0 ;
  assign n30886 = ~n1200 & n3057 ;
  assign n30887 = n30886 ^ n2817 ^ 1'b0 ;
  assign n30888 = n30887 ^ n17314 ^ n2773 ;
  assign n30889 = n30888 ^ n15481 ^ n8925 ;
  assign n30890 = n15338 ^ n10998 ^ n7055 ;
  assign n30891 = ( n8583 & n20067 ) | ( n8583 & ~n30890 ) | ( n20067 & ~n30890 ) ;
  assign n30892 = ( n11249 & n29714 ) | ( n11249 & ~n30891 ) | ( n29714 & ~n30891 ) ;
  assign n30893 = n5098 ^ n4724 ^ 1'b0 ;
  assign n30894 = n2440 | n30893 ;
  assign n30895 = n8162 & n30894 ;
  assign n30896 = ( n3898 & ~n27355 ) | ( n3898 & n30895 ) | ( ~n27355 & n30895 ) ;
  assign n30897 = ( ~n610 & n3118 ) | ( ~n610 & n14562 ) | ( n3118 & n14562 ) ;
  assign n30898 = n30897 ^ n28091 ^ 1'b0 ;
  assign n30899 = n13918 & n30898 ;
  assign n30900 = n30899 ^ n16517 ^ 1'b0 ;
  assign n30901 = n30900 ^ n29824 ^ n25474 ;
  assign n30902 = ( n6539 & n12966 ) | ( n6539 & ~n22891 ) | ( n12966 & ~n22891 ) ;
  assign n30903 = n11803 ^ n5979 ^ 1'b0 ;
  assign n30904 = n23838 & n30903 ;
  assign n30905 = n20536 & n30904 ;
  assign n30906 = n4707 ^ n3910 ^ 1'b0 ;
  assign n30907 = n17442 & ~n30906 ;
  assign n30908 = n1566 & n30907 ;
  assign n30909 = n12663 & n30908 ;
  assign n30910 = n21695 ^ n14261 ^ 1'b0 ;
  assign n30911 = n5472 & n30910 ;
  assign n30912 = n24230 ^ n4209 ^ 1'b0 ;
  assign n30913 = n2472 & n30912 ;
  assign n30914 = ~n30911 & n30913 ;
  assign n30915 = n21687 ^ n18750 ^ 1'b0 ;
  assign n30919 = n7624 & ~n10816 ;
  assign n30916 = n5434 ^ n2676 ^ 1'b0 ;
  assign n30917 = ~n435 & n30916 ;
  assign n30918 = n30917 ^ n1483 ^ 1'b0 ;
  assign n30920 = n30919 ^ n30918 ^ n8442 ;
  assign n30921 = n4736 & n27438 ;
  assign n30922 = ~n3456 & n30921 ;
  assign n30923 = ( n7753 & n9296 ) | ( n7753 & ~n30922 ) | ( n9296 & ~n30922 ) ;
  assign n30924 = ( ~n8311 & n14432 ) | ( ~n8311 & n14869 ) | ( n14432 & n14869 ) ;
  assign n30925 = n4448 ^ n702 ^ 1'b0 ;
  assign n30926 = n4057 ^ n1053 ^ n752 ;
  assign n30927 = n1189 | n1239 ;
  assign n30928 = n30926 | n30927 ;
  assign n30929 = ( ~n30924 & n30925 ) | ( ~n30924 & n30928 ) | ( n30925 & n30928 ) ;
  assign n30930 = n17559 & n18844 ;
  assign n30931 = n13752 ^ n3082 ^ 1'b0 ;
  assign n30932 = n27881 & n30931 ;
  assign n30933 = n30932 ^ n12663 ^ 1'b0 ;
  assign n30934 = ( x35 & n30930 ) | ( x35 & n30933 ) | ( n30930 & n30933 ) ;
  assign n30935 = ( n6903 & ~n10090 ) | ( n6903 & n14656 ) | ( ~n10090 & n14656 ) ;
  assign n30936 = n19995 ^ n3385 ^ n3305 ;
  assign n30937 = n5356 & ~n7497 ;
  assign n30938 = n30937 ^ n1048 ^ 1'b0 ;
  assign n30939 = n195 & ~n29121 ;
  assign n30940 = n18796 & n30939 ;
  assign n30941 = n21171 ^ n138 ^ 1'b0 ;
  assign n30942 = n21804 | n30941 ;
  assign n30943 = n19694 ^ n3097 ^ 1'b0 ;
  assign n30944 = n15733 & n30943 ;
  assign n30945 = ( n11160 & ~n21464 ) | ( n11160 & n28076 ) | ( ~n21464 & n28076 ) ;
  assign n30946 = n19273 ^ n5566 ^ n2637 ;
  assign n30947 = n7795 & n14604 ;
  assign n30948 = n30947 ^ n16457 ^ 1'b0 ;
  assign n30949 = n21403 ^ n1291 ^ 1'b0 ;
  assign n30950 = ( n6991 & ~n16751 ) | ( n6991 & n20561 ) | ( ~n16751 & n20561 ) ;
  assign n30951 = n30950 ^ n15171 ^ 1'b0 ;
  assign n30952 = n4230 ^ n217 ^ 1'b0 ;
  assign n30953 = n2402 | n30952 ;
  assign n30954 = n30953 ^ n12066 ^ 1'b0 ;
  assign n30955 = n9297 ^ n5601 ^ x48 ;
  assign n30956 = ~n18300 & n30955 ;
  assign n30957 = n30956 ^ n4786 ^ 1'b0 ;
  assign n30958 = n3020 & ~n18464 ;
  assign n30959 = n1681 & n30958 ;
  assign n30960 = n30959 ^ n8734 ^ 1'b0 ;
  assign n30961 = n16891 ^ n8850 ^ n5357 ;
  assign n30962 = n28741 ^ n9344 ^ n6509 ;
  assign n30963 = ( ~n4910 & n30961 ) | ( ~n4910 & n30962 ) | ( n30961 & n30962 ) ;
  assign n30964 = n21742 ^ n20918 ^ 1'b0 ;
  assign n30965 = n30964 ^ n27141 ^ n21465 ;
  assign n30966 = n10729 | n17110 ;
  assign n30967 = n30966 ^ n1704 ^ 1'b0 ;
  assign n30968 = n30967 ^ n25653 ^ n13451 ;
  assign n30969 = n24692 ^ n703 ^ n673 ;
  assign n30970 = n30969 ^ n16486 ^ n7807 ;
  assign n30971 = n3677 | n8788 ;
  assign n30972 = n6442 ^ n480 ^ 1'b0 ;
  assign n30973 = n30971 | n30972 ;
  assign n30974 = n30973 ^ n10972 ^ n10526 ;
  assign n30975 = n7144 & n22768 ;
  assign n30976 = n6633 & n19356 ;
  assign n30977 = ( n5278 & ~n8002 ) | ( n5278 & n19808 ) | ( ~n8002 & n19808 ) ;
  assign n30978 = n2835 & ~n3478 ;
  assign n30979 = ~n12189 & n30978 ;
  assign n30980 = n30979 ^ n11708 ^ 1'b0 ;
  assign n30981 = n24365 ^ n16106 ^ n10765 ;
  assign n30982 = n30981 ^ n8405 ^ n6659 ;
  assign n30983 = n2206 ^ n265 ^ 1'b0 ;
  assign n30984 = n18538 & ~n22327 ;
  assign n30986 = n5785 & n17109 ;
  assign n30987 = ~n5345 & n30986 ;
  assign n30988 = n24075 | n30987 ;
  assign n30989 = n30988 ^ n924 ^ 1'b0 ;
  assign n30985 = n4239 & ~n10571 ;
  assign n30990 = n30989 ^ n30985 ^ n22143 ;
  assign n30991 = x43 & ~n30575 ;
  assign n30992 = n15381 | n18398 ;
  assign n30993 = n30992 ^ n26866 ^ n2980 ;
  assign n30994 = n23809 ^ n16275 ^ 1'b0 ;
  assign n30995 = n30993 | n30994 ;
  assign n30996 = n23979 ^ n3354 ^ 1'b0 ;
  assign n30997 = n7207 & ~n30996 ;
  assign n30998 = ~n5134 & n9162 ;
  assign n30999 = n13851 ^ n9639 ^ n2445 ;
  assign n31000 = n30999 ^ n11441 ^ 1'b0 ;
  assign n31001 = n27578 ^ n16944 ^ 1'b0 ;
  assign n31002 = ~n24613 & n27427 ;
  assign n31003 = n21703 ^ n10045 ^ n2270 ;
  assign n31004 = ( n13567 & n22714 ) | ( n13567 & n31003 ) | ( n22714 & n31003 ) ;
  assign n31005 = n890 | n13636 ;
  assign n31006 = n31005 ^ n27436 ^ n6571 ;
  assign n31007 = ( n11319 & n12486 ) | ( n11319 & n31006 ) | ( n12486 & n31006 ) ;
  assign n31008 = n21139 ^ n3950 ^ 1'b0 ;
  assign n31009 = n4366 & ~n31008 ;
  assign n31010 = n15768 ^ n6182 ^ 1'b0 ;
  assign n31011 = n2900 & ~n31010 ;
  assign n31012 = n26390 ^ n17278 ^ n11553 ;
  assign n31013 = n25784 ^ n4812 ^ n1946 ;
  assign n31014 = n31012 & n31013 ;
  assign n31015 = n30880 ^ n4033 ^ n3044 ;
  assign n31016 = n20645 ^ n9312 ^ 1'b0 ;
  assign n31017 = n4583 & n31016 ;
  assign n31018 = n31017 ^ n24818 ^ x47 ;
  assign n31019 = n30108 & n31018 ;
  assign n31020 = ( ~n8761 & n30677 ) | ( ~n8761 & n31019 ) | ( n30677 & n31019 ) ;
  assign n31021 = n6294 ^ n2838 ^ 1'b0 ;
  assign n31022 = n31021 ^ n30857 ^ n7919 ;
  assign n31023 = n31022 ^ n1976 ^ 1'b0 ;
  assign n31025 = n9014 ^ n8895 ^ n7671 ;
  assign n31024 = ~n4033 & n15731 ;
  assign n31026 = n31025 ^ n31024 ^ n22668 ;
  assign n31027 = n1115 | n6637 ;
  assign n31028 = n6411 | n31027 ;
  assign n31029 = n31028 ^ n22126 ^ 1'b0 ;
  assign n31030 = n31029 ^ n22881 ^ n373 ;
  assign n31032 = ( n2370 & ~n5521 ) | ( n2370 & n15760 ) | ( ~n5521 & n15760 ) ;
  assign n31031 = n26058 ^ n21285 ^ n14291 ;
  assign n31033 = n31032 ^ n31031 ^ n23988 ;
  assign n31034 = n6987 & ~n21444 ;
  assign n31035 = n31034 ^ x105 ^ 1'b0 ;
  assign n31036 = n9251 | n15451 ;
  assign n31037 = n2363 & n8495 ;
  assign n31038 = n31037 ^ n22898 ^ 1'b0 ;
  assign n31039 = n4571 & ~n31038 ;
  assign n31040 = n31039 ^ n13922 ^ 1'b0 ;
  assign n31041 = ~n10855 & n14466 ;
  assign n31042 = n31040 & n31041 ;
  assign n31043 = ~n23107 & n31042 ;
  assign n31044 = n20645 ^ n19843 ^ 1'b0 ;
  assign n31045 = n12225 & ~n31044 ;
  assign n31046 = ( n3418 & n5814 ) | ( n3418 & n17540 ) | ( n5814 & n17540 ) ;
  assign n31047 = n7603 ^ n1525 ^ n225 ;
  assign n31048 = n2119 | n17241 ;
  assign n31049 = n31048 ^ n10293 ^ 1'b0 ;
  assign n31050 = ( ~n2551 & n29433 ) | ( ~n2551 & n31049 ) | ( n29433 & n31049 ) ;
  assign n31051 = n21696 ^ n1248 ^ 1'b0 ;
  assign n31052 = ~n5129 & n31051 ;
  assign n31053 = n25122 ^ n1926 ^ 1'b0 ;
  assign n31054 = n31052 & n31053 ;
  assign n31055 = n31054 ^ n7116 ^ n3728 ;
  assign n31056 = n13104 | n26459 ;
  assign n31057 = x85 & ~n3457 ;
  assign n31058 = ( n8252 & ~n19517 ) | ( n8252 & n26145 ) | ( ~n19517 & n26145 ) ;
  assign n31059 = n16555 & n31058 ;
  assign n31060 = n31059 ^ n3728 ^ 1'b0 ;
  assign n31061 = n31060 ^ n8440 ^ n2681 ;
  assign n31062 = n31061 ^ n10125 ^ x86 ;
  assign n31063 = ( n1609 & n31057 ) | ( n1609 & ~n31062 ) | ( n31057 & ~n31062 ) ;
  assign n31064 = ( n1460 & n6879 ) | ( n1460 & ~n17354 ) | ( n6879 & ~n17354 ) ;
  assign n31065 = ( ~n1470 & n4039 ) | ( ~n1470 & n31064 ) | ( n4039 & n31064 ) ;
  assign n31066 = n31065 ^ n19290 ^ n8283 ;
  assign n31067 = n17426 | n18957 ;
  assign n31068 = n31066 | n31067 ;
  assign n31069 = n4408 & n13100 ;
  assign n31070 = n26051 ^ n25339 ^ 1'b0 ;
  assign n31071 = n981 | n31070 ;
  assign n31072 = n13468 ^ n10005 ^ n7382 ;
  assign n31073 = n10630 ^ n9685 ^ 1'b0 ;
  assign n31074 = ~n31072 & n31073 ;
  assign n31075 = n12283 ^ n6705 ^ n580 ;
  assign n31076 = n18823 ^ n11640 ^ 1'b0 ;
  assign n31077 = n31075 | n31076 ;
  assign n31078 = n22867 ^ n14441 ^ n11596 ;
  assign n31079 = n31078 ^ n7022 ^ n2935 ;
  assign n31081 = ( n5764 & n6149 ) | ( n5764 & n11741 ) | ( n6149 & n11741 ) ;
  assign n31080 = n29504 ^ n15380 ^ n7166 ;
  assign n31082 = n31081 ^ n31080 ^ n10968 ;
  assign n31083 = ( n5948 & n8754 ) | ( n5948 & ~n15046 ) | ( n8754 & ~n15046 ) ;
  assign n31084 = n25339 ^ n12138 ^ 1'b0 ;
  assign n31085 = n19878 ^ n7309 ^ 1'b0 ;
  assign n31086 = n31085 ^ n7231 ^ n1509 ;
  assign n31087 = n16969 ^ x97 ^ 1'b0 ;
  assign n31088 = ~n17496 & n31087 ;
  assign n31089 = n25517 & n31088 ;
  assign n31090 = n11110 & n30999 ;
  assign n31091 = n31090 ^ n26804 ^ 1'b0 ;
  assign n31092 = n3947 & ~n31091 ;
  assign n31093 = ~n7748 & n31092 ;
  assign n31094 = n4445 & ~n18049 ;
  assign n31095 = n4527 ^ n4106 ^ 1'b0 ;
  assign n31096 = n4358 & ~n31095 ;
  assign n31097 = ~n31094 & n31096 ;
  assign n31098 = n23412 & n31097 ;
  assign n31099 = n22968 & n31098 ;
  assign n31100 = n27641 ^ n4720 ^ 1'b0 ;
  assign n31101 = n1544 & ~n8064 ;
  assign n31102 = n29369 & n31101 ;
  assign n31103 = ~n5070 & n16017 ;
  assign n31104 = n31103 ^ n29096 ^ 1'b0 ;
  assign n31105 = n8078 ^ n971 ^ 1'b0 ;
  assign n31106 = n31105 ^ n26591 ^ n5089 ;
  assign n31107 = ( ~n7747 & n9953 ) | ( ~n7747 & n16712 ) | ( n9953 & n16712 ) ;
  assign n31109 = ~n2144 & n4739 ;
  assign n31108 = ( n2106 & n11022 ) | ( n2106 & ~n15310 ) | ( n11022 & ~n15310 ) ;
  assign n31110 = n31109 ^ n31108 ^ n29874 ;
  assign n31111 = n16996 ^ n16504 ^ n10299 ;
  assign n31112 = ( n1357 & n6427 ) | ( n1357 & ~n31111 ) | ( n6427 & ~n31111 ) ;
  assign n31113 = n302 | n3704 ;
  assign n31114 = n31113 ^ n26421 ^ 1'b0 ;
  assign n31115 = n2462 & n24422 ;
  assign n31116 = n31115 ^ n5773 ^ 1'b0 ;
  assign n31117 = n31116 ^ n11714 ^ 1'b0 ;
  assign n31118 = n3216 & n31117 ;
  assign n31119 = n31118 ^ n505 ^ 1'b0 ;
  assign n31124 = n8151 ^ n3073 ^ n2687 ;
  assign n31120 = n18945 ^ n11524 ^ n9121 ;
  assign n31121 = n30708 ^ n4531 ^ n836 ;
  assign n31122 = n18116 ^ n15734 ^ n15404 ;
  assign n31123 = ( ~n31120 & n31121 ) | ( ~n31120 & n31122 ) | ( n31121 & n31122 ) ;
  assign n31125 = n31124 ^ n31123 ^ n19005 ;
  assign n31126 = n16464 ^ n8570 ^ n7703 ;
  assign n31127 = n13944 ^ n9794 ^ 1'b0 ;
  assign n31128 = n17256 ^ n11830 ^ n8184 ;
  assign n31129 = ( n7161 & n14158 ) | ( n7161 & n16181 ) | ( n14158 & n16181 ) ;
  assign n31130 = ( n10919 & n16379 ) | ( n10919 & ~n18736 ) | ( n16379 & ~n18736 ) ;
  assign n31131 = ( ~n31128 & n31129 ) | ( ~n31128 & n31130 ) | ( n31129 & n31130 ) ;
  assign n31132 = n10653 & ~n27922 ;
  assign n31133 = n31132 ^ n2441 ^ 1'b0 ;
  assign n31134 = n31133 ^ n18664 ^ n16338 ;
  assign n31135 = n17384 ^ n1375 ^ 1'b0 ;
  assign n31136 = n31135 ^ n2593 ^ n2556 ;
  assign n31137 = n24890 ^ n19534 ^ n2711 ;
  assign n31138 = x60 & n9287 ;
  assign n31139 = n31138 ^ n18993 ^ 1'b0 ;
  assign n31140 = n31137 & ~n31139 ;
  assign n31141 = ( n4890 & n10265 ) | ( n4890 & n26100 ) | ( n10265 & n26100 ) ;
  assign n31142 = ~n1268 & n14953 ;
  assign n31143 = n27294 & n31142 ;
  assign n31144 = n31141 & n31143 ;
  assign n31145 = n18309 ^ n10642 ^ n5070 ;
  assign n31146 = n3969 | n31145 ;
  assign n31147 = n31146 ^ n8842 ^ 1'b0 ;
  assign n31148 = n2900 & ~n23499 ;
  assign n31149 = n31147 & n31148 ;
  assign n31153 = n5295 & ~n8052 ;
  assign n31154 = n31153 ^ n12365 ^ n7660 ;
  assign n31155 = n31154 ^ n15535 ^ n11428 ;
  assign n31150 = n3462 & n27966 ;
  assign n31151 = n31150 ^ n25519 ^ 1'b0 ;
  assign n31152 = n1382 & ~n31151 ;
  assign n31156 = n31155 ^ n31152 ^ 1'b0 ;
  assign n31157 = n19620 ^ n11013 ^ n10184 ;
  assign n31158 = n6064 & n12949 ;
  assign n31159 = n31158 ^ n23750 ^ 1'b0 ;
  assign n31160 = n31159 ^ n21795 ^ n4724 ;
  assign n31161 = ( n343 & n10689 ) | ( n343 & ~n17369 ) | ( n10689 & ~n17369 ) ;
  assign n31162 = ( ~n10827 & n22750 ) | ( ~n10827 & n30373 ) | ( n22750 & n30373 ) ;
  assign n31163 = ( n6546 & n31161 ) | ( n6546 & n31162 ) | ( n31161 & n31162 ) ;
  assign n31164 = n7743 & n14886 ;
  assign n31165 = n156 & ~n5747 ;
  assign n31166 = n31165 ^ n7401 ^ 1'b0 ;
  assign n31167 = ( n28252 & n31164 ) | ( n28252 & n31166 ) | ( n31164 & n31166 ) ;
  assign n31168 = n29394 & n31167 ;
  assign n31169 = ( n16422 & n31163 ) | ( n16422 & n31168 ) | ( n31163 & n31168 ) ;
  assign n31170 = n25869 ^ n21334 ^ 1'b0 ;
  assign n31171 = n29737 ^ n15791 ^ n9902 ;
  assign n31172 = n15893 | n31171 ;
  assign n31173 = ( n10609 & n18435 ) | ( n10609 & n31172 ) | ( n18435 & n31172 ) ;
  assign n31175 = n6948 & ~n9466 ;
  assign n31174 = n10852 & ~n15105 ;
  assign n31176 = n31175 ^ n31174 ^ 1'b0 ;
  assign n31177 = n31176 ^ n29699 ^ n15273 ;
  assign n31178 = ~n146 & n17930 ;
  assign n31179 = n9352 & n31178 ;
  assign n31180 = n18474 ^ n12356 ^ 1'b0 ;
  assign n31181 = n31180 ^ n17028 ^ n7765 ;
  assign n31182 = n21703 ^ n13038 ^ 1'b0 ;
  assign n31183 = n4434 & ~n31182 ;
  assign n31184 = n31183 ^ n9315 ^ 1'b0 ;
  assign n31185 = ~n31181 & n31184 ;
  assign n31186 = n18722 ^ n8540 ^ n7272 ;
  assign n31187 = n6226 & n23653 ;
  assign n31188 = ~n962 & n31187 ;
  assign n31189 = n6424 & ~n18787 ;
  assign n31190 = n4381 & n6019 ;
  assign n31191 = n6692 & n31190 ;
  assign n31192 = ( ~n2653 & n26850 ) | ( ~n2653 & n31191 ) | ( n26850 & n31191 ) ;
  assign n31193 = n31192 ^ n31080 ^ n25491 ;
  assign n31194 = ( ~n332 & n3169 ) | ( ~n332 & n5978 ) | ( n3169 & n5978 ) ;
  assign n31195 = n26739 ^ n24196 ^ n5411 ;
  assign n31196 = n31195 ^ n30089 ^ 1'b0 ;
  assign n31197 = ( n2325 & ~n5824 ) | ( n2325 & n7589 ) | ( ~n5824 & n7589 ) ;
  assign n31198 = ( n21826 & n23467 ) | ( n21826 & ~n31197 ) | ( n23467 & ~n31197 ) ;
  assign n31199 = n25271 ^ n18932 ^ 1'b0 ;
  assign n31200 = n29202 ^ n9005 ^ n5312 ;
  assign n31201 = ~n17997 & n31200 ;
  assign n31202 = n2904 & n26825 ;
  assign n31203 = n31202 ^ n9250 ^ 1'b0 ;
  assign n31204 = n1190 & ~n1898 ;
  assign n31205 = n31204 ^ n24537 ^ 1'b0 ;
  assign n31206 = n10830 ^ n10078 ^ 1'b0 ;
  assign n31207 = ~n3392 & n6837 ;
  assign n31208 = n22173 ^ n3823 ^ n1614 ;
  assign n31209 = n12462 & n29727 ;
  assign n31210 = ~n1738 & n15023 ;
  assign n31211 = n31210 ^ n25668 ^ n2708 ;
  assign n31212 = n17514 ^ n13902 ^ 1'b0 ;
  assign n31213 = n3182 & ~n31212 ;
  assign n31214 = ( n3897 & n3926 ) | ( n3897 & n4035 ) | ( n3926 & n4035 ) ;
  assign n31215 = n31214 ^ n6588 ^ 1'b0 ;
  assign n31216 = n4057 & n29076 ;
  assign n31217 = n31216 ^ n8922 ^ 1'b0 ;
  assign n31218 = n31217 ^ n2928 ^ x54 ;
  assign n31219 = n15894 | n19710 ;
  assign n31220 = ~n3474 & n5122 ;
  assign n31221 = n31220 ^ n3047 ^ 1'b0 ;
  assign n31222 = n31221 ^ n3723 ^ 1'b0 ;
  assign n31223 = n19987 ^ n16500 ^ n7554 ;
  assign n31224 = ~n5875 & n31223 ;
  assign n31225 = ~n31222 & n31224 ;
  assign n31226 = ~n15494 & n18756 ;
  assign n31227 = n31226 ^ n14865 ^ 1'b0 ;
  assign n31228 = n4513 | n30003 ;
  assign n31229 = n16495 & ~n31228 ;
  assign n31230 = n11411 | n19043 ;
  assign n31231 = n25807 | n26203 ;
  assign n31232 = ( n13882 & n17681 ) | ( n13882 & ~n22066 ) | ( n17681 & ~n22066 ) ;
  assign n31233 = ( n9183 & n14300 ) | ( n9183 & n31232 ) | ( n14300 & n31232 ) ;
  assign n31234 = n24371 ^ n1853 ^ 1'b0 ;
  assign n31236 = n23537 ^ n1500 ^ 1'b0 ;
  assign n31237 = n31236 ^ n21274 ^ n12503 ;
  assign n31235 = n15030 ^ n9455 ^ n8812 ;
  assign n31238 = n31237 ^ n31235 ^ n2111 ;
  assign n31239 = n5649 & ~n13307 ;
  assign n31240 = n27902 ^ n3992 ^ 1'b0 ;
  assign n31241 = n31239 & n31240 ;
  assign n31242 = ( n1147 & n29150 ) | ( n1147 & n31241 ) | ( n29150 & n31241 ) ;
  assign n31243 = n8304 ^ n1718 ^ 1'b0 ;
  assign n31244 = ~n12748 & n31243 ;
  assign n31245 = n9227 ^ n8888 ^ 1'b0 ;
  assign n31246 = n18262 | n31245 ;
  assign n31247 = n29644 ^ n9918 ^ 1'b0 ;
  assign n31248 = ~n21983 & n31247 ;
  assign n31249 = n7583 & n29104 ;
  assign n31250 = n29117 & n31249 ;
  assign n31251 = n19761 ^ n19356 ^ n4985 ;
  assign n31252 = n2744 | n11118 ;
  assign n31253 = ( ~n3085 & n12710 ) | ( ~n3085 & n28972 ) | ( n12710 & n28972 ) ;
  assign n31254 = n604 & n22520 ;
  assign n31255 = n19791 & n31254 ;
  assign n31256 = ( n9970 & n25107 ) | ( n9970 & ~n31255 ) | ( n25107 & ~n31255 ) ;
  assign n31257 = ( n8432 & n22971 ) | ( n8432 & n28550 ) | ( n22971 & n28550 ) ;
  assign n31258 = ( n519 & ~n13291 ) | ( n519 & n22845 ) | ( ~n13291 & n22845 ) ;
  assign n31259 = ( n5103 & ~n11806 ) | ( n5103 & n31258 ) | ( ~n11806 & n31258 ) ;
  assign n31260 = ( n4524 & n14158 ) | ( n4524 & ~n16190 ) | ( n14158 & ~n16190 ) ;
  assign n31261 = n3126 | n31260 ;
  assign n31262 = n1617 | n31261 ;
  assign n31263 = n13054 & n31262 ;
  assign n31264 = n31263 ^ n24525 ^ n2026 ;
  assign n31265 = ( n3102 & ~n12001 ) | ( n3102 & n17535 ) | ( ~n12001 & n17535 ) ;
  assign n31266 = n10407 & n19963 ;
  assign n31267 = n31266 ^ n15511 ^ 1'b0 ;
  assign n31268 = n31265 & n31267 ;
  assign n31269 = n9402 & ~n14574 ;
  assign n31270 = ~n13164 & n24399 ;
  assign n31271 = n4241 | n31270 ;
  assign n31272 = n16037 & ~n31271 ;
  assign n31273 = n25623 ^ n16181 ^ 1'b0 ;
  assign n31274 = ( n30282 & n31272 ) | ( n30282 & ~n31273 ) | ( n31272 & ~n31273 ) ;
  assign n31275 = ( ~n4336 & n10057 ) | ( ~n4336 & n16338 ) | ( n10057 & n16338 ) ;
  assign n31276 = ( n6744 & ~n16049 ) | ( n6744 & n31275 ) | ( ~n16049 & n31275 ) ;
  assign n31277 = n13058 ^ n1032 ^ 1'b0 ;
  assign n31278 = ( n10403 & n10472 ) | ( n10403 & ~n31277 ) | ( n10472 & ~n31277 ) ;
  assign n31279 = ( n4815 & n20751 ) | ( n4815 & n22803 ) | ( n20751 & n22803 ) ;
  assign n31280 = n8389 ^ n3804 ^ 1'b0 ;
  assign n31281 = n29600 | n31280 ;
  assign n31282 = n148 & n21536 ;
  assign n31283 = ( n20043 & ~n31281 ) | ( n20043 & n31282 ) | ( ~n31281 & n31282 ) ;
  assign n31284 = ( ~n2020 & n9217 ) | ( ~n2020 & n12207 ) | ( n9217 & n12207 ) ;
  assign n31285 = n15284 | n31284 ;
  assign n31286 = n5198 | n23705 ;
  assign n31287 = ( ~n3435 & n5419 ) | ( ~n3435 & n24219 ) | ( n5419 & n24219 ) ;
  assign n31288 = n15052 & n31287 ;
  assign n31289 = n31288 ^ n8372 ^ 1'b0 ;
  assign n31290 = n2716 & n30565 ;
  assign n31291 = n31290 ^ n10587 ^ 1'b0 ;
  assign n31293 = n17384 ^ n11794 ^ 1'b0 ;
  assign n31294 = n4889 & ~n31293 ;
  assign n31292 = n16504 | n22121 ;
  assign n31295 = n31294 ^ n31292 ^ 1'b0 ;
  assign n31296 = ~n5242 & n5566 ;
  assign n31297 = ~n10979 & n31296 ;
  assign n31298 = ( n5769 & ~n12260 ) | ( n5769 & n21742 ) | ( ~n12260 & n21742 ) ;
  assign n31299 = n17389 ^ n9516 ^ n7639 ;
  assign n31300 = ( n1896 & ~n5137 ) | ( n1896 & n16742 ) | ( ~n5137 & n16742 ) ;
  assign n31301 = ~n359 & n31300 ;
  assign n31302 = n18247 & ~n19006 ;
  assign n31303 = ~n15495 & n31302 ;
  assign n31304 = n31303 ^ n7990 ^ 1'b0 ;
  assign n31305 = ( n8379 & n18348 ) | ( n8379 & n23222 ) | ( n18348 & n23222 ) ;
  assign n31306 = n6290 | n14941 ;
  assign n31307 = ( n807 & n23573 ) | ( n807 & n31306 ) | ( n23573 & n31306 ) ;
  assign n31308 = n13460 & ~n31138 ;
  assign n31309 = ( n10731 & n28720 ) | ( n10731 & n31308 ) | ( n28720 & n31308 ) ;
  assign n31310 = ~n19288 & n31309 ;
  assign n31311 = n31310 ^ n10989 ^ 1'b0 ;
  assign n31312 = n8529 ^ n1593 ^ 1'b0 ;
  assign n31313 = n10973 & ~n31312 ;
  assign n31314 = ( n15481 & n19850 ) | ( n15481 & n23022 ) | ( n19850 & n23022 ) ;
  assign n31315 = ( n13345 & n23013 ) | ( n13345 & n31314 ) | ( n23013 & n31314 ) ;
  assign n31316 = n8358 ^ n785 ^ 1'b0 ;
  assign n31317 = ~n31315 & n31316 ;
  assign n31318 = ~n5339 & n18058 ;
  assign n31319 = n19285 ^ n10004 ^ 1'b0 ;
  assign n31320 = ( n19937 & n26659 ) | ( n19937 & ~n31319 ) | ( n26659 & ~n31319 ) ;
  assign n31321 = n25041 ^ n11677 ^ n7330 ;
  assign n31322 = n6516 | n28510 ;
  assign n31323 = n2492 & ~n31322 ;
  assign n31324 = ( n8348 & n23214 ) | ( n8348 & n31323 ) | ( n23214 & n31323 ) ;
  assign n31325 = n3802 ^ n3445 ^ 1'b0 ;
  assign n31326 = n9021 & ~n31325 ;
  assign n31327 = n26715 | n31326 ;
  assign n31328 = n10313 ^ n375 ^ 1'b0 ;
  assign n31329 = n21061 ^ n19581 ^ n8790 ;
  assign n31330 = ( n18250 & n31328 ) | ( n18250 & ~n31329 ) | ( n31328 & ~n31329 ) ;
  assign n31331 = n8689 | n25084 ;
  assign n31333 = n15207 ^ n9322 ^ n3057 ;
  assign n31332 = ~n313 & n15541 ;
  assign n31334 = n31333 ^ n31332 ^ 1'b0 ;
  assign n31335 = n31334 ^ n23599 ^ 1'b0 ;
  assign n31336 = n31331 | n31335 ;
  assign n31337 = n4312 ^ n3918 ^ 1'b0 ;
  assign n31338 = n9070 | n31337 ;
  assign n31339 = ( ~n896 & n4105 ) | ( ~n896 & n19532 ) | ( n4105 & n19532 ) ;
  assign n31340 = n31339 ^ n29547 ^ x30 ;
  assign n31341 = n26252 ^ n268 ^ 1'b0 ;
  assign n31342 = n31340 | n31341 ;
  assign n31343 = n8209 & ~n8767 ;
  assign n31344 = n2682 & n31343 ;
  assign n31345 = n4787 & ~n31344 ;
  assign n31346 = ~n15343 & n31345 ;
  assign n31347 = n8794 ^ n3074 ^ 1'b0 ;
  assign n31348 = n31346 | n31347 ;
  assign n31349 = n11684 ^ n11677 ^ n2395 ;
  assign n31350 = ( n18998 & ~n25331 ) | ( n18998 & n25878 ) | ( ~n25331 & n25878 ) ;
  assign n31351 = n8094 & n11332 ;
  assign n31352 = ~n5368 & n31351 ;
  assign n31353 = n31352 ^ n3469 ^ 1'b0 ;
  assign n31354 = ( ~n11080 & n31350 ) | ( ~n11080 & n31353 ) | ( n31350 & n31353 ) ;
  assign n31355 = ( n1784 & n7967 ) | ( n1784 & ~n31354 ) | ( n7967 & ~n31354 ) ;
  assign n31356 = ~n511 & n9966 ;
  assign n31357 = ( n1407 & n1980 ) | ( n1407 & ~n4425 ) | ( n1980 & ~n4425 ) ;
  assign n31358 = ( ~n23935 & n31356 ) | ( ~n23935 & n31357 ) | ( n31356 & n31357 ) ;
  assign n31359 = n22092 ^ n3481 ^ n1653 ;
  assign n31360 = ( ~n786 & n31358 ) | ( ~n786 & n31359 ) | ( n31358 & n31359 ) ;
  assign n31361 = n131 | n4175 ;
  assign n31362 = n31361 ^ n8958 ^ 1'b0 ;
  assign n31363 = n31362 ^ n13222 ^ n5162 ;
  assign n31364 = n25905 ^ n2109 ^ 1'b0 ;
  assign n31365 = n12844 & n31364 ;
  assign n31366 = ( n10077 & n31363 ) | ( n10077 & n31365 ) | ( n31363 & n31365 ) ;
  assign n31367 = n10260 ^ n8409 ^ n3995 ;
  assign n31368 = ( x41 & n1765 ) | ( x41 & n7097 ) | ( n1765 & n7097 ) ;
  assign n31369 = ~n6855 & n10911 ;
  assign n31370 = ~n31368 & n31369 ;
  assign n31371 = ( n648 & ~n31367 ) | ( n648 & n31370 ) | ( ~n31367 & n31370 ) ;
  assign n31372 = ( n2108 & n20846 ) | ( n2108 & ~n31371 ) | ( n20846 & ~n31371 ) ;
  assign n31375 = n11534 ^ n9966 ^ n6102 ;
  assign n31376 = ~n4684 & n10589 ;
  assign n31377 = n31375 & n31376 ;
  assign n31373 = n17569 ^ n8128 ^ 1'b0 ;
  assign n31374 = n607 & n31373 ;
  assign n31378 = n31377 ^ n31374 ^ n26906 ;
  assign n31379 = n1908 & n18526 ;
  assign n31382 = n10051 ^ n7939 ^ n5262 ;
  assign n31381 = n14259 & ~n15598 ;
  assign n31383 = n31382 ^ n31381 ^ 1'b0 ;
  assign n31380 = n10289 | n18839 ;
  assign n31384 = n31383 ^ n31380 ^ 1'b0 ;
  assign n31385 = ~n13011 & n14496 ;
  assign n31386 = n20400 & n31385 ;
  assign n31387 = n13427 & ~n19562 ;
  assign n31388 = n31386 & n31387 ;
  assign n31389 = n9168 | n13351 ;
  assign n31390 = n22791 & n23407 ;
  assign n31391 = ~n31389 & n31390 ;
  assign n31392 = n14977 | n31391 ;
  assign n31393 = n31392 ^ n30446 ^ 1'b0 ;
  assign n31394 = n23192 ^ n9353 ^ 1'b0 ;
  assign n31395 = n11076 & ~n31394 ;
  assign n31396 = ( n24786 & n31192 ) | ( n24786 & n31395 ) | ( n31192 & n31395 ) ;
  assign n31397 = ( n6276 & ~n14554 ) | ( n6276 & n31396 ) | ( ~n14554 & n31396 ) ;
  assign n31398 = ~n3077 & n10185 ;
  assign n31399 = ( ~n12212 & n24060 ) | ( ~n12212 & n30550 ) | ( n24060 & n30550 ) ;
  assign n31400 = n26411 ^ n9395 ^ n2193 ;
  assign n31401 = n19489 ^ n5154 ^ 1'b0 ;
  assign n31402 = n16147 ^ n7691 ^ n3947 ;
  assign n31403 = ~n19566 & n31402 ;
  assign n31404 = ~n26655 & n31403 ;
  assign n31405 = ( n3473 & ~n31401 ) | ( n3473 & n31404 ) | ( ~n31401 & n31404 ) ;
  assign n31406 = n4844 ^ n3160 ^ n1633 ;
  assign n31407 = n27014 ^ n892 ^ 1'b0 ;
  assign n31408 = n31406 | n31407 ;
  assign n31409 = n10601 & ~n23127 ;
  assign n31410 = n16016 & n31409 ;
  assign n31411 = n1404 & n31410 ;
  assign n31412 = n10365 & n29017 ;
  assign n31413 = n30333 & n31412 ;
  assign n31414 = n31413 ^ n681 ^ 1'b0 ;
  assign n31415 = n30553 & ~n31414 ;
  assign n31416 = ( n2487 & ~n14251 ) | ( n2487 & n19783 ) | ( ~n14251 & n19783 ) ;
  assign n31417 = n31416 ^ n8148 ^ 1'b0 ;
  assign n31418 = n2786 & n31417 ;
  assign n31419 = ( n7059 & ~n17434 ) | ( n7059 & n31418 ) | ( ~n17434 & n31418 ) ;
  assign n31421 = n8107 | n11256 ;
  assign n31420 = n22865 & ~n25138 ;
  assign n31422 = n31421 ^ n31420 ^ 1'b0 ;
  assign n31423 = n12962 & ~n31422 ;
  assign n31424 = n10925 | n18813 ;
  assign n31425 = ( ~n6525 & n11528 ) | ( ~n6525 & n19709 ) | ( n11528 & n19709 ) ;
  assign n31426 = ~n11771 & n31425 ;
  assign n31427 = ~n2697 & n31426 ;
  assign n31428 = n9177 | n26115 ;
  assign n31429 = n12882 & n18504 ;
  assign n31430 = n30947 ^ n2226 ^ 1'b0 ;
  assign n31431 = n6792 & ~n31430 ;
  assign n31432 = ~n4724 & n31431 ;
  assign n31433 = n25098 ^ n12024 ^ n4629 ;
  assign n31434 = n8107 ^ n5221 ^ 1'b0 ;
  assign n31435 = n31433 | n31434 ;
  assign n31438 = n6731 ^ n3256 ^ n3113 ;
  assign n31436 = n12274 ^ n4224 ^ n235 ;
  assign n31437 = n31436 ^ n14053 ^ n4390 ;
  assign n31439 = n31438 ^ n31437 ^ n6632 ;
  assign n31440 = n27488 ^ n7207 ^ n3900 ;
  assign n31441 = ( ~n1472 & n31396 ) | ( ~n1472 & n31440 ) | ( n31396 & n31440 ) ;
  assign n31442 = ( ~n10266 & n13893 ) | ( ~n10266 & n14292 ) | ( n13893 & n14292 ) ;
  assign n31443 = ( n15874 & n16525 ) | ( n15874 & ~n19853 ) | ( n16525 & ~n19853 ) ;
  assign n31444 = ~n23992 & n30045 ;
  assign n31445 = ( n10081 & ~n31443 ) | ( n10081 & n31444 ) | ( ~n31443 & n31444 ) ;
  assign n31446 = n28212 ^ n14087 ^ n9431 ;
  assign n31447 = n31446 ^ n11500 ^ n243 ;
  assign n31448 = ~n8098 & n14934 ;
  assign n31449 = n31448 ^ n13871 ^ 1'b0 ;
  assign n31450 = n11014 ^ n10320 ^ 1'b0 ;
  assign n31451 = n10671 & ~n31450 ;
  assign n31452 = ~n20642 & n31451 ;
  assign n31453 = ( ~n8408 & n31449 ) | ( ~n8408 & n31452 ) | ( n31449 & n31452 ) ;
  assign n31454 = n29692 ^ n1709 ^ 1'b0 ;
  assign n31455 = ~n5474 & n31454 ;
  assign n31456 = n31455 ^ n30437 ^ n10868 ;
  assign n31457 = ~n524 & n31456 ;
  assign n31458 = n31457 ^ n6415 ^ 1'b0 ;
  assign n31459 = ( n4657 & n11913 ) | ( n4657 & ~n16754 ) | ( n11913 & ~n16754 ) ;
  assign n31460 = n10733 & ~n17647 ;
  assign n31461 = ~n7828 & n31460 ;
  assign n31462 = ~n31459 & n31461 ;
  assign n31463 = n2315 | n31462 ;
  assign n31464 = n31463 ^ n18376 ^ 1'b0 ;
  assign n31466 = n11149 & n13741 ;
  assign n31467 = n5826 & n31466 ;
  assign n31465 = ~n28204 & n28340 ;
  assign n31468 = n31467 ^ n31465 ^ 1'b0 ;
  assign n31469 = n4187 & ~n13312 ;
  assign n31470 = n21327 & n31469 ;
  assign n31471 = n31470 ^ n25486 ^ 1'b0 ;
  assign n31472 = n21110 | n28678 ;
  assign n31473 = n31472 ^ n22247 ^ 1'b0 ;
  assign y0 = x12 ;
  assign y1 = x20 ;
  assign y2 = x23 ;
  assign y3 = x25 ;
  assign y4 = x42 ;
  assign y5 = x53 ;
  assign y6 = x57 ;
  assign y7 = x64 ;
  assign y8 = x71 ;
  assign y9 = x72 ;
  assign y10 = x75 ;
  assign y11 = x91 ;
  assign y12 = x94 ;
  assign y13 = x102 ;
  assign y14 = x103 ;
  assign y15 = x106 ;
  assign y16 = x127 ;
  assign y17 = n129 ;
  assign y18 = ~n130 ;
  assign y19 = ~n131 ;
  assign y20 = ~n133 ;
  assign y21 = ~n134 ;
  assign y22 = n137 ;
  assign y23 = ~n138 ;
  assign y24 = n143 ;
  assign y25 = ~1'b0 ;
  assign y26 = ~n146 ;
  assign y27 = ~1'b0 ;
  assign y28 = ~n150 ;
  assign y29 = n151 ;
  assign y30 = ~n157 ;
  assign y31 = ~n160 ;
  assign y32 = n164 ;
  assign y33 = ~n169 ;
  assign y34 = ~n170 ;
  assign y35 = n176 ;
  assign y36 = n178 ;
  assign y37 = ~n179 ;
  assign y38 = n181 ;
  assign y39 = ~n190 ;
  assign y40 = n194 ;
  assign y41 = n195 ;
  assign y42 = n199 ;
  assign y43 = ~1'b0 ;
  assign y44 = n201 ;
  assign y45 = n207 ;
  assign y46 = n215 ;
  assign y47 = ~n218 ;
  assign y48 = ~n219 ;
  assign y49 = ~1'b0 ;
  assign y50 = ~x66 ;
  assign y51 = n222 ;
  assign y52 = ~n227 ;
  assign y53 = ~n230 ;
  assign y54 = ~n244 ;
  assign y55 = n247 ;
  assign y56 = ~n248 ;
  assign y57 = ~n249 ;
  assign y58 = n259 ;
  assign y59 = n260 ;
  assign y60 = ~1'b0 ;
  assign y61 = n266 ;
  assign y62 = ~n267 ;
  assign y63 = ~n277 ;
  assign y64 = n285 ;
  assign y65 = ~n286 ;
  assign y66 = n287 ;
  assign y67 = ~n305 ;
  assign y68 = ~n312 ;
  assign y69 = n314 ;
  assign y70 = ~n325 ;
  assign y71 = n330 ;
  assign y72 = ~1'b0 ;
  assign y73 = ~n334 ;
  assign y74 = n337 ;
  assign y75 = n342 ;
  assign y76 = n346 ;
  assign y77 = ~n364 ;
  assign y78 = n365 ;
  assign y79 = ~n367 ;
  assign y80 = n370 ;
  assign y81 = ~n390 ;
  assign y82 = n393 ;
  assign y83 = ~n399 ;
  assign y84 = n406 ;
  assign y85 = ~n408 ;
  assign y86 = n416 ;
  assign y87 = ~n418 ;
  assign y88 = n421 ;
  assign y89 = ~n426 ;
  assign y90 = ~n435 ;
  assign y91 = ~1'b0 ;
  assign y92 = ~1'b0 ;
  assign y93 = n437 ;
  assign y94 = n438 ;
  assign y95 = ~n447 ;
  assign y96 = ~n450 ;
  assign y97 = ~n456 ;
  assign y98 = ~n465 ;
  assign y99 = ~1'b0 ;
  assign y100 = ~n471 ;
  assign y101 = ~n476 ;
  assign y102 = ~n478 ;
  assign y103 = n480 ;
  assign y104 = n484 ;
  assign y105 = ~n486 ;
  assign y106 = n489 ;
  assign y107 = n495 ;
  assign y108 = ~n499 ;
  assign y109 = n501 ;
  assign y110 = ~n503 ;
  assign y111 = n509 ;
  assign y112 = n512 ;
  assign y113 = ~1'b0 ;
  assign y114 = n515 ;
  assign y115 = n519 ;
  assign y116 = ~n524 ;
  assign y117 = n526 ;
  assign y118 = ~n527 ;
  assign y119 = ~n533 ;
  assign y120 = n542 ;
  assign y121 = ~n557 ;
  assign y122 = n563 ;
  assign y123 = n570 ;
  assign y124 = ~1'b0 ;
  assign y125 = ~n576 ;
  assign y126 = ~n577 ;
  assign y127 = ~n579 ;
  assign y128 = n581 ;
  assign y129 = ~n583 ;
  assign y130 = n588 ;
  assign y131 = ~n589 ;
  assign y132 = n598 ;
  assign y133 = ~n600 ;
  assign y134 = n601 ;
  assign y135 = n602 ;
  assign y136 = ~1'b0 ;
  assign y137 = ~n606 ;
  assign y138 = ~n610 ;
  assign y139 = ~n619 ;
  assign y140 = ~n621 ;
  assign y141 = n626 ;
  assign y142 = n628 ;
  assign y143 = n631 ;
  assign y144 = ~n639 ;
  assign y145 = ~n650 ;
  assign y146 = ~n657 ;
  assign y147 = ~n659 ;
  assign y148 = n688 ;
  assign y149 = ~n692 ;
  assign y150 = n696 ;
  assign y151 = n697 ;
  assign y152 = n700 ;
  assign y153 = ~1'b0 ;
  assign y154 = n720 ;
  assign y155 = n722 ;
  assign y156 = ~n724 ;
  assign y157 = ~n728 ;
  assign y158 = n729 ;
  assign y159 = ~1'b0 ;
  assign y160 = n731 ;
  assign y161 = n732 ;
  assign y162 = ~1'b0 ;
  assign y163 = ~n740 ;
  assign y164 = n741 ;
  assign y165 = ~n746 ;
  assign y166 = ~n752 ;
  assign y167 = ~n753 ;
  assign y168 = ~n757 ;
  assign y169 = ~n764 ;
  assign y170 = ~n777 ;
  assign y171 = n780 ;
  assign y172 = ~n782 ;
  assign y173 = ~n783 ;
  assign y174 = ~n785 ;
  assign y175 = ~n788 ;
  assign y176 = n792 ;
  assign y177 = n796 ;
  assign y178 = ~1'b0 ;
  assign y179 = n800 ;
  assign y180 = n806 ;
  assign y181 = n808 ;
  assign y182 = ~n811 ;
  assign y183 = n814 ;
  assign y184 = n816 ;
  assign y185 = ~1'b0 ;
  assign y186 = ~n817 ;
  assign y187 = ~1'b0 ;
  assign y188 = ~1'b0 ;
  assign y189 = ~n826 ;
  assign y190 = n830 ;
  assign y191 = n832 ;
  assign y192 = ~1'b0 ;
  assign y193 = n835 ;
  assign y194 = ~n840 ;
  assign y195 = n847 ;
  assign y196 = n858 ;
  assign y197 = ~n859 ;
  assign y198 = ~n867 ;
  assign y199 = n871 ;
  assign y200 = ~n878 ;
  assign y201 = n886 ;
  assign y202 = n892 ;
  assign y203 = n894 ;
  assign y204 = n896 ;
  assign y205 = ~1'b0 ;
  assign y206 = n760 ;
  assign y207 = n900 ;
  assign y208 = n905 ;
  assign y209 = ~n907 ;
  assign y210 = ~n910 ;
  assign y211 = n912 ;
  assign y212 = n915 ;
  assign y213 = ~n916 ;
  assign y214 = ~n921 ;
  assign y215 = n927 ;
  assign y216 = n941 ;
  assign y217 = ~n948 ;
  assign y218 = n955 ;
  assign y219 = n956 ;
  assign y220 = n961 ;
  assign y221 = n965 ;
  assign y222 = n967 ;
  assign y223 = ~n971 ;
  assign y224 = n974 ;
  assign y225 = n976 ;
  assign y226 = ~n980 ;
  assign y227 = n986 ;
  assign y228 = n990 ;
  assign y229 = n997 ;
  assign y230 = ~n998 ;
  assign y231 = ~n1001 ;
  assign y232 = ~n1004 ;
  assign y233 = ~1'b0 ;
  assign y234 = n1005 ;
  assign y235 = ~1'b0 ;
  assign y236 = n1015 ;
  assign y237 = n1021 ;
  assign y238 = n1030 ;
  assign y239 = ~n1032 ;
  assign y240 = ~n1040 ;
  assign y241 = n1044 ;
  assign y242 = n1049 ;
  assign y243 = ~n1057 ;
  assign y244 = ~1'b0 ;
  assign y245 = n1063 ;
  assign y246 = n1071 ;
  assign y247 = n1095 ;
  assign y248 = ~n1099 ;
  assign y249 = n1100 ;
  assign y250 = n1104 ;
  assign y251 = n1106 ;
  assign y252 = ~n1111 ;
  assign y253 = ~n1114 ;
  assign y254 = ~n1115 ;
  assign y255 = ~n1120 ;
  assign y256 = n1126 ;
  assign y257 = ~n1127 ;
  assign y258 = ~n1130 ;
  assign y259 = ~n1139 ;
  assign y260 = ~n1142 ;
  assign y261 = n1148 ;
  assign y262 = ~1'b0 ;
  assign y263 = n1150 ;
  assign y264 = n1153 ;
  assign y265 = ~n1157 ;
  assign y266 = n1168 ;
  assign y267 = ~n1174 ;
  assign y268 = ~1'b0 ;
  assign y269 = ~n1177 ;
  assign y270 = ~n1183 ;
  assign y271 = ~x84 ;
  assign y272 = n1191 ;
  assign y273 = ~n1193 ;
  assign y274 = ~n1205 ;
  assign y275 = n1206 ;
  assign y276 = ~1'b0 ;
  assign y277 = n1214 ;
  assign y278 = ~n1221 ;
  assign y279 = ~n1227 ;
  assign y280 = ~1'b0 ;
  assign y281 = n1233 ;
  assign y282 = ~1'b0 ;
  assign y283 = n1235 ;
  assign y284 = n1237 ;
  assign y285 = ~n1239 ;
  assign y286 = ~n1242 ;
  assign y287 = ~n1243 ;
  assign y288 = ~n1253 ;
  assign y289 = ~n1262 ;
  assign y290 = n1264 ;
  assign y291 = ~n1266 ;
  assign y292 = n1276 ;
  assign y293 = ~n1283 ;
  assign y294 = n1284 ;
  assign y295 = ~n1288 ;
  assign y296 = n1289 ;
  assign y297 = ~n896 ;
  assign y298 = ~n1296 ;
  assign y299 = n1306 ;
  assign y300 = ~n1313 ;
  assign y301 = n1314 ;
  assign y302 = ~1'b0 ;
  assign y303 = n1318 ;
  assign y304 = n1324 ;
  assign y305 = ~1'b0 ;
  assign y306 = ~n1326 ;
  assign y307 = n1340 ;
  assign y308 = n1341 ;
  assign y309 = ~n1346 ;
  assign y310 = ~1'b0 ;
  assign y311 = ~1'b0 ;
  assign y312 = n1349 ;
  assign y313 = ~1'b0 ;
  assign y314 = ~n1353 ;
  assign y315 = ~n1354 ;
  assign y316 = ~n1359 ;
  assign y317 = n1369 ;
  assign y318 = n1373 ;
  assign y319 = ~n1378 ;
  assign y320 = ~n1380 ;
  assign y321 = n1382 ;
  assign y322 = ~n1390 ;
  assign y323 = ~n1394 ;
  assign y324 = ~n1395 ;
  assign y325 = ~n1396 ;
  assign y326 = ~n1397 ;
  assign y327 = ~n1401 ;
  assign y328 = n1405 ;
  assign y329 = ~n1406 ;
  assign y330 = ~n1414 ;
  assign y331 = ~n1418 ;
  assign y332 = ~n1425 ;
  assign y333 = ~n1426 ;
  assign y334 = ~n1430 ;
  assign y335 = ~n1433 ;
  assign y336 = ~1'b0 ;
  assign y337 = ~n1441 ;
  assign y338 = ~n1442 ;
  assign y339 = n1447 ;
  assign y340 = ~n1450 ;
  assign y341 = n1454 ;
  assign y342 = ~n1457 ;
  assign y343 = n1459 ;
  assign y344 = n1466 ;
  assign y345 = ~n1468 ;
  assign y346 = ~1'b0 ;
  assign y347 = n1476 ;
  assign y348 = n1479 ;
  assign y349 = ~n1485 ;
  assign y350 = n1493 ;
  assign y351 = n1500 ;
  assign y352 = ~n1508 ;
  assign y353 = ~1'b0 ;
  assign y354 = ~n1515 ;
  assign y355 = ~n1518 ;
  assign y356 = ~n1522 ;
  assign y357 = n1524 ;
  assign y358 = ~1'b0 ;
  assign y359 = n1529 ;
  assign y360 = ~n1534 ;
  assign y361 = ~n1205 ;
  assign y362 = n1544 ;
  assign y363 = n1551 ;
  assign y364 = ~n1555 ;
  assign y365 = n1559 ;
  assign y366 = ~1'b0 ;
  assign y367 = n1563 ;
  assign y368 = n1566 ;
  assign y369 = n1567 ;
  assign y370 = n1570 ;
  assign y371 = ~n1571 ;
  assign y372 = ~1'b0 ;
  assign y373 = ~n1582 ;
  assign y374 = ~1'b0 ;
  assign y375 = n1586 ;
  assign y376 = ~n1589 ;
  assign y377 = n1590 ;
  assign y378 = ~1'b0 ;
  assign y379 = ~1'b0 ;
  assign y380 = n1593 ;
  assign y381 = ~n1597 ;
  assign y382 = n1600 ;
  assign y383 = n1613 ;
  assign y384 = ~n1616 ;
  assign y385 = ~1'b0 ;
  assign y386 = n1617 ;
  assign y387 = n1618 ;
  assign y388 = n1631 ;
  assign y389 = ~n1634 ;
  assign y390 = ~n1636 ;
  assign y391 = ~1'b0 ;
  assign y392 = n1641 ;
  assign y393 = ~1'b0 ;
  assign y394 = n1648 ;
  assign y395 = ~n1657 ;
  assign y396 = ~1'b0 ;
  assign y397 = n1663 ;
  assign y398 = ~n1665 ;
  assign y399 = n1666 ;
  assign y400 = n1681 ;
  assign y401 = ~n1687 ;
  assign y402 = ~n1697 ;
  assign y403 = n1699 ;
  assign y404 = n1700 ;
  assign y405 = n1703 ;
  assign y406 = ~n1704 ;
  assign y407 = n1708 ;
  assign y408 = ~n1711 ;
  assign y409 = ~1'b0 ;
  assign y410 = n1714 ;
  assign y411 = ~n1715 ;
  assign y412 = n1718 ;
  assign y413 = ~n1720 ;
  assign y414 = n1724 ;
  assign y415 = ~n1729 ;
  assign y416 = ~n1732 ;
  assign y417 = ~n1734 ;
  assign y418 = ~n1738 ;
  assign y419 = ~n1739 ;
  assign y420 = ~1'b0 ;
  assign y421 = ~n1742 ;
  assign y422 = ~n1747 ;
  assign y423 = n1748 ;
  assign y424 = ~n1750 ;
  assign y425 = ~n1754 ;
  assign y426 = ~1'b0 ;
  assign y427 = n1762 ;
  assign y428 = ~n1763 ;
  assign y429 = ~n1764 ;
  assign y430 = ~n1765 ;
  assign y431 = ~n1780 ;
  assign y432 = ~1'b0 ;
  assign y433 = ~n1790 ;
  assign y434 = n1796 ;
  assign y435 = ~n1805 ;
  assign y436 = ~n1809 ;
  assign y437 = ~n1821 ;
  assign y438 = ~n1826 ;
  assign y439 = ~n1829 ;
  assign y440 = ~n1831 ;
  assign y441 = n1833 ;
  assign y442 = n1844 ;
  assign y443 = ~1'b0 ;
  assign y444 = ~n1849 ;
  assign y445 = ~1'b0 ;
  assign y446 = n1854 ;
  assign y447 = n1857 ;
  assign y448 = ~1'b0 ;
  assign y449 = n1858 ;
  assign y450 = ~n1863 ;
  assign y451 = ~1'b0 ;
  assign y452 = n1867 ;
  assign y453 = n1873 ;
  assign y454 = ~1'b0 ;
  assign y455 = n1875 ;
  assign y456 = ~n1885 ;
  assign y457 = ~n1887 ;
  assign y458 = n1888 ;
  assign y459 = n1893 ;
  assign y460 = ~n1895 ;
  assign y461 = ~n1898 ;
  assign y462 = ~n1899 ;
  assign y463 = ~n1900 ;
  assign y464 = n1902 ;
  assign y465 = n1905 ;
  assign y466 = ~n1909 ;
  assign y467 = n1914 ;
  assign y468 = ~n1917 ;
  assign y469 = ~1'b0 ;
  assign y470 = n1918 ;
  assign y471 = n1920 ;
  assign y472 = n1923 ;
  assign y473 = ~n1926 ;
  assign y474 = ~n1928 ;
  assign y475 = n1931 ;
  assign y476 = ~n1935 ;
  assign y477 = n1936 ;
  assign y478 = ~n1943 ;
  assign y479 = ~n1947 ;
  assign y480 = n1953 ;
  assign y481 = ~1'b0 ;
  assign y482 = n1962 ;
  assign y483 = ~1'b0 ;
  assign y484 = 1'b0 ;
  assign y485 = ~n1967 ;
  assign y486 = ~n1969 ;
  assign y487 = n1988 ;
  assign y488 = n1989 ;
  assign y489 = n1997 ;
  assign y490 = n2000 ;
  assign y491 = n2014 ;
  assign y492 = ~n2023 ;
  assign y493 = ~n2025 ;
  assign y494 = ~1'b0 ;
  assign y495 = ~n2035 ;
  assign y496 = ~1'b0 ;
  assign y497 = n2037 ;
  assign y498 = ~n2040 ;
  assign y499 = ~1'b0 ;
  assign y500 = ~n2045 ;
  assign y501 = ~n2051 ;
  assign y502 = n2060 ;
  assign y503 = n2061 ;
  assign y504 = ~n2071 ;
  assign y505 = n2072 ;
  assign y506 = n2075 ;
  assign y507 = n2079 ;
  assign y508 = n2085 ;
  assign y509 = ~n2086 ;
  assign y510 = n2093 ;
  assign y511 = ~n2095 ;
  assign y512 = ~n2096 ;
  assign y513 = ~1'b0 ;
  assign y514 = n2098 ;
  assign y515 = ~n2100 ;
  assign y516 = n2102 ;
  assign y517 = n2117 ;
  assign y518 = n2118 ;
  assign y519 = ~n2119 ;
  assign y520 = n2126 ;
  assign y521 = n2134 ;
  assign y522 = ~n2136 ;
  assign y523 = ~1'b0 ;
  assign y524 = n2137 ;
  assign y525 = ~1'b0 ;
  assign y526 = ~n2140 ;
  assign y527 = ~n2146 ;
  assign y528 = ~n2152 ;
  assign y529 = n2154 ;
  assign y530 = ~n2163 ;
  assign y531 = ~n2168 ;
  assign y532 = n2169 ;
  assign y533 = n2181 ;
  assign y534 = n2187 ;
  assign y535 = n2194 ;
  assign y536 = n2195 ;
  assign y537 = ~n2196 ;
  assign y538 = ~n2198 ;
  assign y539 = x19 ;
  assign y540 = ~n2199 ;
  assign y541 = n2201 ;
  assign y542 = n2209 ;
  assign y543 = n2211 ;
  assign y544 = ~1'b0 ;
  assign y545 = n2213 ;
  assign y546 = n2215 ;
  assign y547 = ~n2216 ;
  assign y548 = n2223 ;
  assign y549 = n2224 ;
  assign y550 = n2232 ;
  assign y551 = ~1'b0 ;
  assign y552 = ~n2242 ;
  assign y553 = ~n2247 ;
  assign y554 = n2252 ;
  assign y555 = n2254 ;
  assign y556 = n2255 ;
  assign y557 = ~n2257 ;
  assign y558 = n2259 ;
  assign y559 = n2261 ;
  assign y560 = n2274 ;
  assign y561 = ~1'b0 ;
  assign y562 = ~1'b0 ;
  assign y563 = ~n2276 ;
  assign y564 = n2277 ;
  assign y565 = ~1'b0 ;
  assign y566 = ~n2281 ;
  assign y567 = n2289 ;
  assign y568 = n2295 ;
  assign y569 = n2304 ;
  assign y570 = ~n2312 ;
  assign y571 = ~n2315 ;
  assign y572 = ~n2317 ;
  assign y573 = ~n2326 ;
  assign y574 = ~n2337 ;
  assign y575 = ~n2339 ;
  assign y576 = ~n2341 ;
  assign y577 = ~n2342 ;
  assign y578 = ~1'b0 ;
  assign y579 = ~n2353 ;
  assign y580 = ~n2364 ;
  assign y581 = ~n2374 ;
  assign y582 = n2376 ;
  assign y583 = ~n2377 ;
  assign y584 = n2378 ;
  assign y585 = ~n2385 ;
  assign y586 = ~n2392 ;
  assign y587 = n2398 ;
  assign y588 = ~n2401 ;
  assign y589 = ~1'b0 ;
  assign y590 = n2409 ;
  assign y591 = n2414 ;
  assign y592 = ~n2421 ;
  assign y593 = n2423 ;
  assign y594 = n2427 ;
  assign y595 = n2433 ;
  assign y596 = n2435 ;
  assign y597 = ~n2438 ;
  assign y598 = ~n2449 ;
  assign y599 = n2451 ;
  assign y600 = ~1'b0 ;
  assign y601 = n2455 ;
  assign y602 = n1456 ;
  assign y603 = ~n2461 ;
  assign y604 = ~1'b0 ;
  assign y605 = n2462 ;
  assign y606 = ~n2463 ;
  assign y607 = n2464 ;
  assign y608 = ~1'b0 ;
  assign y609 = ~n2466 ;
  assign y610 = n2468 ;
  assign y611 = n2472 ;
  assign y612 = ~n2477 ;
  assign y613 = ~n2478 ;
  assign y614 = n2479 ;
  assign y615 = ~n2486 ;
  assign y616 = n2491 ;
  assign y617 = n2493 ;
  assign y618 = ~n2499 ;
  assign y619 = ~n2504 ;
  assign y620 = ~n2512 ;
  assign y621 = n2534 ;
  assign y622 = ~n2537 ;
  assign y623 = ~n2547 ;
  assign y624 = n2549 ;
  assign y625 = ~n2554 ;
  assign y626 = ~n2557 ;
  assign y627 = ~n2562 ;
  assign y628 = ~n2567 ;
  assign y629 = n2575 ;
  assign y630 = ~n2582 ;
  assign y631 = n2602 ;
  assign y632 = n2607 ;
  assign y633 = n2615 ;
  assign y634 = ~1'b0 ;
  assign y635 = n2616 ;
  assign y636 = n2618 ;
  assign y637 = ~n2619 ;
  assign y638 = n2622 ;
  assign y639 = ~n2625 ;
  assign y640 = ~n2626 ;
  assign y641 = n2635 ;
  assign y642 = ~n2640 ;
  assign y643 = n2641 ;
  assign y644 = ~1'b0 ;
  assign y645 = ~1'b0 ;
  assign y646 = n2644 ;
  assign y647 = ~n2649 ;
  assign y648 = ~n2659 ;
  assign y649 = ~n2660 ;
  assign y650 = n2665 ;
  assign y651 = ~1'b0 ;
  assign y652 = ~n2667 ;
  assign y653 = ~n2668 ;
  assign y654 = ~n2670 ;
  assign y655 = ~n2673 ;
  assign y656 = n2674 ;
  assign y657 = ~1'b0 ;
  assign y658 = n2679 ;
  assign y659 = ~n2682 ;
  assign y660 = n2683 ;
  assign y661 = ~n2684 ;
  assign y662 = ~n2703 ;
  assign y663 = ~n2707 ;
  assign y664 = n2710 ;
  assign y665 = ~1'b0 ;
  assign y666 = n2711 ;
  assign y667 = ~n2714 ;
  assign y668 = n2716 ;
  assign y669 = n2726 ;
  assign y670 = ~n2728 ;
  assign y671 = ~n2731 ;
  assign y672 = n2733 ;
  assign y673 = n2739 ;
  assign y674 = ~n2740 ;
  assign y675 = n2741 ;
  assign y676 = n2742 ;
  assign y677 = ~n2754 ;
  assign y678 = n2757 ;
  assign y679 = n2759 ;
  assign y680 = n2773 ;
  assign y681 = ~n2778 ;
  assign y682 = ~n2783 ;
  assign y683 = ~n2791 ;
  assign y684 = ~n2793 ;
  assign y685 = ~1'b0 ;
  assign y686 = n2796 ;
  assign y687 = ~n298 ;
  assign y688 = n2799 ;
  assign y689 = n2804 ;
  assign y690 = ~1'b0 ;
  assign y691 = ~1'b0 ;
  assign y692 = n2807 ;
  assign y693 = ~n2815 ;
  assign y694 = ~n2817 ;
  assign y695 = ~n2818 ;
  assign y696 = ~n2820 ;
  assign y697 = n2823 ;
  assign y698 = ~n2824 ;
  assign y699 = ~n2839 ;
  assign y700 = ~n2843 ;
  assign y701 = ~n2853 ;
  assign y702 = ~n2854 ;
  assign y703 = ~n2859 ;
  assign y704 = ~1'b0 ;
  assign y705 = ~n2860 ;
  assign y706 = ~n2867 ;
  assign y707 = ~n2869 ;
  assign y708 = n2873 ;
  assign y709 = ~n2875 ;
  assign y710 = ~n2878 ;
  assign y711 = ~n2883 ;
  assign y712 = n2892 ;
  assign y713 = ~n2893 ;
  assign y714 = n2895 ;
  assign y715 = ~n2897 ;
  assign y716 = n2900 ;
  assign y717 = ~n2903 ;
  assign y718 = ~1'b0 ;
  assign y719 = ~n2908 ;
  assign y720 = n2912 ;
  assign y721 = ~n2913 ;
  assign y722 = n2915 ;
  assign y723 = ~n2916 ;
  assign y724 = ~n2918 ;
  assign y725 = ~n2919 ;
  assign y726 = n2923 ;
  assign y727 = ~n2924 ;
  assign y728 = n2930 ;
  assign y729 = ~n2935 ;
  assign y730 = n2937 ;
  assign y731 = ~n2949 ;
  assign y732 = ~n2954 ;
  assign y733 = ~n2959 ;
  assign y734 = n2965 ;
  assign y735 = ~1'b0 ;
  assign y736 = ~n2981 ;
  assign y737 = ~1'b0 ;
  assign y738 = ~n2989 ;
  assign y739 = n2992 ;
  assign y740 = ~n2996 ;
  assign y741 = ~n3001 ;
  assign y742 = ~n3008 ;
  assign y743 = ~1'b0 ;
  assign y744 = n3011 ;
  assign y745 = n3013 ;
  assign y746 = n3015 ;
  assign y747 = ~n3019 ;
  assign y748 = ~n3022 ;
  assign y749 = ~n3029 ;
  assign y750 = n3039 ;
  assign y751 = ~n3043 ;
  assign y752 = ~n3045 ;
  assign y753 = n3047 ;
  assign y754 = ~1'b0 ;
  assign y755 = ~1'b0 ;
  assign y756 = n3057 ;
  assign y757 = ~1'b0 ;
  assign y758 = n3059 ;
  assign y759 = n3064 ;
  assign y760 = ~n3072 ;
  assign y761 = n3074 ;
  assign y762 = ~1'b0 ;
  assign y763 = ~n3079 ;
  assign y764 = ~n3084 ;
  assign y765 = ~n3087 ;
  assign y766 = n3088 ;
  assign y767 = n3091 ;
  assign y768 = ~n3092 ;
  assign y769 = ~n3094 ;
  assign y770 = n3099 ;
  assign y771 = ~n3103 ;
  assign y772 = n3108 ;
  assign y773 = ~n3118 ;
  assign y774 = ~n3119 ;
  assign y775 = n3120 ;
  assign y776 = ~n3121 ;
  assign y777 = n3126 ;
  assign y778 = n3129 ;
  assign y779 = n3133 ;
  assign y780 = ~n3137 ;
  assign y781 = n3142 ;
  assign y782 = ~n3154 ;
  assign y783 = n3157 ;
  assign y784 = ~n3161 ;
  assign y785 = ~1'b0 ;
  assign y786 = ~n3162 ;
  assign y787 = n3163 ;
  assign y788 = ~n3165 ;
  assign y789 = ~1'b0 ;
  assign y790 = ~n3167 ;
  assign y791 = ~n3183 ;
  assign y792 = n3186 ;
  assign y793 = n3190 ;
  assign y794 = n3202 ;
  assign y795 = n3204 ;
  assign y796 = ~1'b0 ;
  assign y797 = n3205 ;
  assign y798 = ~n3206 ;
  assign y799 = ~n3207 ;
  assign y800 = n3210 ;
  assign y801 = n3216 ;
  assign y802 = ~n3222 ;
  assign y803 = n3238 ;
  assign y804 = ~n3241 ;
  assign y805 = n3242 ;
  assign y806 = ~1'b0 ;
  assign y807 = ~1'b0 ;
  assign y808 = ~n3245 ;
  assign y809 = ~n3254 ;
  assign y810 = ~n3256 ;
  assign y811 = n3257 ;
  assign y812 = ~1'b0 ;
  assign y813 = n3258 ;
  assign y814 = ~1'b0 ;
  assign y815 = ~n3261 ;
  assign y816 = n376 ;
  assign y817 = n3262 ;
  assign y818 = n3263 ;
  assign y819 = n3264 ;
  assign y820 = n3267 ;
  assign y821 = n3270 ;
  assign y822 = ~n3285 ;
  assign y823 = ~1'b0 ;
  assign y824 = n3287 ;
  assign y825 = n3292 ;
  assign y826 = ~n3298 ;
  assign y827 = ~n3299 ;
  assign y828 = ~1'b0 ;
  assign y829 = n3301 ;
  assign y830 = n3303 ;
  assign y831 = ~n3307 ;
  assign y832 = n3314 ;
  assign y833 = n3320 ;
  assign y834 = ~n243 ;
  assign y835 = ~1'b0 ;
  assign y836 = ~n3323 ;
  assign y837 = n3328 ;
  assign y838 = ~n3330 ;
  assign y839 = n3331 ;
  assign y840 = n3335 ;
  assign y841 = n3337 ;
  assign y842 = ~n3351 ;
  assign y843 = n3352 ;
  assign y844 = ~n3356 ;
  assign y845 = n3357 ;
  assign y846 = ~n3362 ;
  assign y847 = ~n3370 ;
  assign y848 = n3371 ;
  assign y849 = ~n3375 ;
  assign y850 = n3386 ;
  assign y851 = n3390 ;
  assign y852 = ~n3391 ;
  assign y853 = ~n3393 ;
  assign y854 = n3407 ;
  assign y855 = n3415 ;
  assign y856 = ~n3416 ;
  assign y857 = n3426 ;
  assign y858 = n3438 ;
  assign y859 = ~n3445 ;
  assign y860 = n3448 ;
  assign y861 = ~1'b0 ;
  assign y862 = ~n3451 ;
  assign y863 = n3453 ;
  assign y864 = n3456 ;
  assign y865 = ~1'b0 ;
  assign y866 = ~n3458 ;
  assign y867 = n3462 ;
  assign y868 = ~1'b0 ;
  assign y869 = ~n3464 ;
  assign y870 = n3466 ;
  assign y871 = n3467 ;
  assign y872 = n3470 ;
  assign y873 = ~n3474 ;
  assign y874 = ~n3478 ;
  assign y875 = ~n3480 ;
  assign y876 = ~n3488 ;
  assign y877 = ~n3491 ;
  assign y878 = n3509 ;
  assign y879 = n3513 ;
  assign y880 = ~n3514 ;
  assign y881 = ~n3517 ;
  assign y882 = ~n3521 ;
  assign y883 = n3526 ;
  assign y884 = ~n2399 ;
  assign y885 = n3529 ;
  assign y886 = ~1'b0 ;
  assign y887 = n3531 ;
  assign y888 = ~n3541 ;
  assign y889 = n3552 ;
  assign y890 = 1'b0 ;
  assign y891 = ~n3553 ;
  assign y892 = ~1'b0 ;
  assign y893 = ~1'b0 ;
  assign y894 = ~1'b0 ;
  assign y895 = n3556 ;
  assign y896 = n3561 ;
  assign y897 = ~n3565 ;
  assign y898 = ~n3576 ;
  assign y899 = n3577 ;
  assign y900 = ~n3582 ;
  assign y901 = ~n3585 ;
  assign y902 = n3600 ;
  assign y903 = ~n3607 ;
  assign y904 = n3612 ;
  assign y905 = ~1'b0 ;
  assign y906 = ~n3617 ;
  assign y907 = ~n3619 ;
  assign y908 = ~1'b0 ;
  assign y909 = ~1'b0 ;
  assign y910 = ~n3622 ;
  assign y911 = ~n3625 ;
  assign y912 = ~n3631 ;
  assign y913 = ~n3632 ;
  assign y914 = ~n3634 ;
  assign y915 = n3635 ;
  assign y916 = n3644 ;
  assign y917 = ~n3650 ;
  assign y918 = n3659 ;
  assign y919 = n3662 ;
  assign y920 = n3664 ;
  assign y921 = n3666 ;
  assign y922 = n3670 ;
  assign y923 = n3673 ;
  assign y924 = n3693 ;
  assign y925 = ~n3699 ;
  assign y926 = n3700 ;
  assign y927 = ~1'b0 ;
  assign y928 = ~n3704 ;
  assign y929 = ~n3715 ;
  assign y930 = n3722 ;
  assign y931 = n3726 ;
  assign y932 = n3727 ;
  assign y933 = n3733 ;
  assign y934 = n3734 ;
  assign y935 = ~n3736 ;
  assign y936 = ~n3739 ;
  assign y937 = ~1'b0 ;
  assign y938 = n3742 ;
  assign y939 = n3743 ;
  assign y940 = n3745 ;
  assign y941 = n3752 ;
  assign y942 = ~1'b0 ;
  assign y943 = ~n3757 ;
  assign y944 = n3760 ;
  assign y945 = n3764 ;
  assign y946 = ~n3768 ;
  assign y947 = ~n3769 ;
  assign y948 = n3771 ;
  assign y949 = n3773 ;
  assign y950 = n969 ;
  assign y951 = ~n3775 ;
  assign y952 = n3783 ;
  assign y953 = n3787 ;
  assign y954 = ~n3789 ;
  assign y955 = ~n3795 ;
  assign y956 = n3796 ;
  assign y957 = n3804 ;
  assign y958 = n3805 ;
  assign y959 = n3811 ;
  assign y960 = ~n3815 ;
  assign y961 = ~1'b0 ;
  assign y962 = ~1'b0 ;
  assign y963 = n3816 ;
  assign y964 = n3830 ;
  assign y965 = n3832 ;
  assign y966 = ~1'b0 ;
  assign y967 = n3834 ;
  assign y968 = n3840 ;
  assign y969 = ~1'b0 ;
  assign y970 = n3843 ;
  assign y971 = n3847 ;
  assign y972 = n3848 ;
  assign y973 = ~n1873 ;
  assign y974 = n3852 ;
  assign y975 = n3853 ;
  assign y976 = n3858 ;
  assign y977 = ~1'b0 ;
  assign y978 = ~n3864 ;
  assign y979 = ~n3872 ;
  assign y980 = n3880 ;
  assign y981 = n3887 ;
  assign y982 = n3888 ;
  assign y983 = n3895 ;
  assign y984 = ~n3896 ;
  assign y985 = n3899 ;
  assign y986 = n3902 ;
  assign y987 = ~n3914 ;
  assign y988 = ~1'b0 ;
  assign y989 = n3917 ;
  assign y990 = n3921 ;
  assign y991 = ~1'b0 ;
  assign y992 = ~1'b0 ;
  assign y993 = ~n3926 ;
  assign y994 = n3927 ;
  assign y995 = ~n3930 ;
  assign y996 = n3947 ;
  assign y997 = n3950 ;
  assign y998 = n3959 ;
  assign y999 = n3965 ;
  assign y1000 = n3966 ;
  assign y1001 = ~n3975 ;
  assign y1002 = ~n3979 ;
  assign y1003 = n3981 ;
  assign y1004 = n3984 ;
  assign y1005 = ~n3988 ;
  assign y1006 = n3989 ;
  assign y1007 = ~n3992 ;
  assign y1008 = ~n3995 ;
  assign y1009 = n3996 ;
  assign y1010 = n4004 ;
  assign y1011 = ~1'b0 ;
  assign y1012 = n4011 ;
  assign y1013 = ~n4012 ;
  assign y1014 = ~n4014 ;
  assign y1015 = n4015 ;
  assign y1016 = ~n4028 ;
  assign y1017 = n4029 ;
  assign y1018 = ~1'b0 ;
  assign y1019 = ~1'b0 ;
  assign y1020 = ~n4031 ;
  assign y1021 = ~n4035 ;
  assign y1022 = ~n2950 ;
  assign y1023 = n4047 ;
  assign y1024 = ~1'b0 ;
  assign y1025 = ~n4051 ;
  assign y1026 = ~n4052 ;
  assign y1027 = n4056 ;
  assign y1028 = ~1'b0 ;
  assign y1029 = n4057 ;
  assign y1030 = n4063 ;
  assign y1031 = ~n4066 ;
  assign y1032 = n4067 ;
  assign y1033 = n4068 ;
  assign y1034 = n4069 ;
  assign y1035 = ~1'b0 ;
  assign y1036 = ~1'b0 ;
  assign y1037 = n4077 ;
  assign y1038 = n4079 ;
  assign y1039 = ~n4083 ;
  assign y1040 = ~n4084 ;
  assign y1041 = ~n4089 ;
  assign y1042 = ~n4090 ;
  assign y1043 = ~1'b0 ;
  assign y1044 = n4094 ;
  assign y1045 = ~1'b0 ;
  assign y1046 = ~n4100 ;
  assign y1047 = ~n4108 ;
  assign y1048 = ~n4116 ;
  assign y1049 = ~n4118 ;
  assign y1050 = n4122 ;
  assign y1051 = n4125 ;
  assign y1052 = n4130 ;
  assign y1053 = n4134 ;
  assign y1054 = n4138 ;
  assign y1055 = ~n4145 ;
  assign y1056 = n4146 ;
  assign y1057 = ~n4155 ;
  assign y1058 = ~n4164 ;
  assign y1059 = ~n4166 ;
  assign y1060 = n4170 ;
  assign y1061 = ~1'b0 ;
  assign y1062 = ~n4174 ;
  assign y1063 = ~n4175 ;
  assign y1064 = ~n4182 ;
  assign y1065 = n4184 ;
  assign y1066 = ~n4200 ;
  assign y1067 = ~n4203 ;
  assign y1068 = n4209 ;
  assign y1069 = n4217 ;
  assign y1070 = ~n4219 ;
  assign y1071 = n4220 ;
  assign y1072 = n4221 ;
  assign y1073 = n4224 ;
  assign y1074 = n3253 ;
  assign y1075 = ~n4226 ;
  assign y1076 = ~n4229 ;
  assign y1077 = n4230 ;
  assign y1078 = ~n4237 ;
  assign y1079 = ~n4241 ;
  assign y1080 = ~n4243 ;
  assign y1081 = ~n4252 ;
  assign y1082 = ~n4254 ;
  assign y1083 = ~1'b0 ;
  assign y1084 = ~n4279 ;
  assign y1085 = ~n4283 ;
  assign y1086 = n4286 ;
  assign y1087 = ~n4292 ;
  assign y1088 = ~n4295 ;
  assign y1089 = n4299 ;
  assign y1090 = ~n4301 ;
  assign y1091 = n4303 ;
  assign y1092 = ~n4306 ;
  assign y1093 = ~n4307 ;
  assign y1094 = ~n4312 ;
  assign y1095 = n4314 ;
  assign y1096 = ~n4332 ;
  assign y1097 = ~n4334 ;
  assign y1098 = ~1'b0 ;
  assign y1099 = ~n4339 ;
  assign y1100 = n4345 ;
  assign y1101 = ~n4351 ;
  assign y1102 = ~1'b0 ;
  assign y1103 = ~1'b0 ;
  assign y1104 = n4353 ;
  assign y1105 = n4361 ;
  assign y1106 = ~n4367 ;
  assign y1107 = ~n4369 ;
  assign y1108 = ~1'b0 ;
  assign y1109 = n4373 ;
  assign y1110 = n4380 ;
  assign y1111 = n4382 ;
  assign y1112 = ~n4385 ;
  assign y1113 = n4392 ;
  assign y1114 = n4394 ;
  assign y1115 = ~n4396 ;
  assign y1116 = ~1'b0 ;
  assign y1117 = ~n4397 ;
  assign y1118 = ~n4404 ;
  assign y1119 = ~n4405 ;
  assign y1120 = n4406 ;
  assign y1121 = ~n4411 ;
  assign y1122 = n4415 ;
  assign y1123 = ~1'b0 ;
  assign y1124 = ~n4417 ;
  assign y1125 = n4428 ;
  assign y1126 = ~n4429 ;
  assign y1127 = ~n4431 ;
  assign y1128 = ~1'b0 ;
  assign y1129 = ~n4450 ;
  assign y1130 = ~1'b0 ;
  assign y1131 = ~n4452 ;
  assign y1132 = ~n4455 ;
  assign y1133 = ~1'b0 ;
  assign y1134 = ~n4463 ;
  assign y1135 = n4464 ;
  assign y1136 = n4465 ;
  assign y1137 = n4472 ;
  assign y1138 = ~n1180 ;
  assign y1139 = n4474 ;
  assign y1140 = ~n4475 ;
  assign y1141 = n4478 ;
  assign y1142 = ~n4479 ;
  assign y1143 = ~n4484 ;
  assign y1144 = n4489 ;
  assign y1145 = n4493 ;
  assign y1146 = n4494 ;
  assign y1147 = ~n4497 ;
  assign y1148 = ~n4513 ;
  assign y1149 = n4518 ;
  assign y1150 = n4522 ;
  assign y1151 = ~n4524 ;
  assign y1152 = n4527 ;
  assign y1153 = n4531 ;
  assign y1154 = ~1'b0 ;
  assign y1155 = ~n4532 ;
  assign y1156 = ~n4540 ;
  assign y1157 = n4541 ;
  assign y1158 = ~n4544 ;
  assign y1159 = n4545 ;
  assign y1160 = n4550 ;
  assign y1161 = ~n4554 ;
  assign y1162 = ~n4556 ;
  assign y1163 = n4570 ;
  assign y1164 = n4571 ;
  assign y1165 = n4583 ;
  assign y1166 = ~n4588 ;
  assign y1167 = n4602 ;
  assign y1168 = ~1'b0 ;
  assign y1169 = ~n4611 ;
  assign y1170 = ~n4612 ;
  assign y1171 = ~n4621 ;
  assign y1172 = n4623 ;
  assign y1173 = n4626 ;
  assign y1174 = n4636 ;
  assign y1175 = ~n4638 ;
  assign y1176 = ~1'b0 ;
  assign y1177 = ~n4639 ;
  assign y1178 = ~n4645 ;
  assign y1179 = ~1'b0 ;
  assign y1180 = n4649 ;
  assign y1181 = n4651 ;
  assign y1182 = ~n4065 ;
  assign y1183 = ~n4652 ;
  assign y1184 = ~n4655 ;
  assign y1185 = n4658 ;
  assign y1186 = ~n4660 ;
  assign y1187 = ~n4665 ;
  assign y1188 = n4671 ;
  assign y1189 = n4685 ;
  assign y1190 = ~n4698 ;
  assign y1191 = ~n4703 ;
  assign y1192 = ~n4344 ;
  assign y1193 = n4710 ;
  assign y1194 = n4711 ;
  assign y1195 = ~n4712 ;
  assign y1196 = n4714 ;
  assign y1197 = ~n4720 ;
  assign y1198 = ~n4730 ;
  assign y1199 = n4732 ;
  assign y1200 = ~n4734 ;
  assign y1201 = ~n4738 ;
  assign y1202 = n4751 ;
  assign y1203 = n4757 ;
  assign y1204 = ~n4762 ;
  assign y1205 = ~n4764 ;
  assign y1206 = n4769 ;
  assign y1207 = n4773 ;
  assign y1208 = n4774 ;
  assign y1209 = n4776 ;
  assign y1210 = n4778 ;
  assign y1211 = ~n4782 ;
  assign y1212 = ~n4784 ;
  assign y1213 = n4787 ;
  assign y1214 = ~1'b0 ;
  assign y1215 = n4790 ;
  assign y1216 = n4792 ;
  assign y1217 = n4794 ;
  assign y1218 = ~n4803 ;
  assign y1219 = n4805 ;
  assign y1220 = n4807 ;
  assign y1221 = n4812 ;
  assign y1222 = ~n4816 ;
  assign y1223 = n4822 ;
  assign y1224 = n4827 ;
  assign y1225 = n4831 ;
  assign y1226 = n4832 ;
  assign y1227 = n4835 ;
  assign y1228 = ~n4837 ;
  assign y1229 = n4848 ;
  assign y1230 = ~1'b0 ;
  assign y1231 = ~n4853 ;
  assign y1232 = ~n4854 ;
  assign y1233 = ~n4856 ;
  assign y1234 = n4865 ;
  assign y1235 = n4868 ;
  assign y1236 = n4870 ;
  assign y1237 = ~n4877 ;
  assign y1238 = ~1'b0 ;
  assign y1239 = n4885 ;
  assign y1240 = ~n4891 ;
  assign y1241 = n4893 ;
  assign y1242 = ~n4898 ;
  assign y1243 = ~1'b0 ;
  assign y1244 = ~n4899 ;
  assign y1245 = ~n4903 ;
  assign y1246 = n4904 ;
  assign y1247 = ~n4908 ;
  assign y1248 = ~1'b0 ;
  assign y1249 = n4910 ;
  assign y1250 = ~n4916 ;
  assign y1251 = n4920 ;
  assign y1252 = ~n4922 ;
  assign y1253 = n4929 ;
  assign y1254 = ~n4932 ;
  assign y1255 = ~n4943 ;
  assign y1256 = ~n4944 ;
  assign y1257 = ~n4947 ;
  assign y1258 = n4949 ;
  assign y1259 = ~n4950 ;
  assign y1260 = n4956 ;
  assign y1261 = ~n4964 ;
  assign y1262 = ~n4971 ;
  assign y1263 = ~1'b0 ;
  assign y1264 = n4973 ;
  assign y1265 = n4975 ;
  assign y1266 = n4984 ;
  assign y1267 = n4987 ;
  assign y1268 = ~n4992 ;
  assign y1269 = ~n4996 ;
  assign y1270 = ~n4997 ;
  assign y1271 = ~1'b0 ;
  assign y1272 = ~n4999 ;
  assign y1273 = ~n5001 ;
  assign y1274 = n5002 ;
  assign y1275 = n5003 ;
  assign y1276 = n5010 ;
  assign y1277 = n5012 ;
  assign y1278 = ~1'b0 ;
  assign y1279 = n5014 ;
  assign y1280 = ~n5019 ;
  assign y1281 = ~n5020 ;
  assign y1282 = n5023 ;
  assign y1283 = ~n5024 ;
  assign y1284 = n5025 ;
  assign y1285 = ~n5029 ;
  assign y1286 = ~1'b0 ;
  assign y1287 = ~n5030 ;
  assign y1288 = ~n5033 ;
  assign y1289 = ~n5037 ;
  assign y1290 = ~n5043 ;
  assign y1291 = ~n5046 ;
  assign y1292 = ~n5047 ;
  assign y1293 = n5053 ;
  assign y1294 = n5054 ;
  assign y1295 = ~n5056 ;
  assign y1296 = ~1'b0 ;
  assign y1297 = n5057 ;
  assign y1298 = n5059 ;
  assign y1299 = ~1'b0 ;
  assign y1300 = n5060 ;
  assign y1301 = ~n5064 ;
  assign y1302 = n5066 ;
  assign y1303 = ~n5074 ;
  assign y1304 = ~n5078 ;
  assign y1305 = ~1'b0 ;
  assign y1306 = ~n5079 ;
  assign y1307 = n5080 ;
  assign y1308 = n5085 ;
  assign y1309 = ~n5091 ;
  assign y1310 = n5092 ;
  assign y1311 = ~n5101 ;
  assign y1312 = n5102 ;
  assign y1313 = ~1'b0 ;
  assign y1314 = ~n5104 ;
  assign y1315 = ~n5106 ;
  assign y1316 = n5115 ;
  assign y1317 = ~n5118 ;
  assign y1318 = n5123 ;
  assign y1319 = ~n5128 ;
  assign y1320 = ~n5129 ;
  assign y1321 = ~n5132 ;
  assign y1322 = ~1'b0 ;
  assign y1323 = ~n5139 ;
  assign y1324 = 1'b0 ;
  assign y1325 = n5141 ;
  assign y1326 = ~n5147 ;
  assign y1327 = n5154 ;
  assign y1328 = ~n5161 ;
  assign y1329 = ~n5165 ;
  assign y1330 = n5169 ;
  assign y1331 = ~n5171 ;
  assign y1332 = n5172 ;
  assign y1333 = n5174 ;
  assign y1334 = ~1'b0 ;
  assign y1335 = ~n5176 ;
  assign y1336 = ~n5180 ;
  assign y1337 = ~1'b0 ;
  assign y1338 = ~1'b0 ;
  assign y1339 = ~n5181 ;
  assign y1340 = n5184 ;
  assign y1341 = ~n5197 ;
  assign y1342 = ~n5201 ;
  assign y1343 = n5215 ;
  assign y1344 = ~n5221 ;
  assign y1345 = n5222 ;
  assign y1346 = ~n5229 ;
  assign y1347 = ~n5239 ;
  assign y1348 = n5243 ;
  assign y1349 = n5244 ;
  assign y1350 = ~n5247 ;
  assign y1351 = ~n5253 ;
  assign y1352 = ~n5254 ;
  assign y1353 = n5255 ;
  assign y1354 = n3953 ;
  assign y1355 = n5256 ;
  assign y1356 = n5260 ;
  assign y1357 = ~1'b0 ;
  assign y1358 = ~1'b0 ;
  assign y1359 = ~1'b0 ;
  assign y1360 = ~n5268 ;
  assign y1361 = ~1'b0 ;
  assign y1362 = n5273 ;
  assign y1363 = n5279 ;
  assign y1364 = ~n5283 ;
  assign y1365 = ~n5285 ;
  assign y1366 = ~n293 ;
  assign y1367 = ~1'b0 ;
  assign y1368 = n5299 ;
  assign y1369 = ~n5301 ;
  assign y1370 = n5305 ;
  assign y1371 = n5306 ;
  assign y1372 = n5309 ;
  assign y1373 = ~n5321 ;
  assign y1374 = ~1'b0 ;
  assign y1375 = ~n5337 ;
  assign y1376 = ~n5340 ;
  assign y1377 = n5348 ;
  assign y1378 = ~n5349 ;
  assign y1379 = n5352 ;
  assign y1380 = ~1'b0 ;
  assign y1381 = n5360 ;
  assign y1382 = ~1'b0 ;
  assign y1383 = ~n5361 ;
  assign y1384 = n5369 ;
  assign y1385 = ~n5376 ;
  assign y1386 = ~n5377 ;
  assign y1387 = n5380 ;
  assign y1388 = n5383 ;
  assign y1389 = ~n5385 ;
  assign y1390 = n5386 ;
  assign y1391 = ~n5390 ;
  assign y1392 = n5398 ;
  assign y1393 = ~n5401 ;
  assign y1394 = n5405 ;
  assign y1395 = n5413 ;
  assign y1396 = n5415 ;
  assign y1397 = ~n5429 ;
  assign y1398 = ~n5436 ;
  assign y1399 = n5440 ;
  assign y1400 = ~n5448 ;
  assign y1401 = n5449 ;
  assign y1402 = ~n5453 ;
  assign y1403 = n5456 ;
  assign y1404 = ~n5462 ;
  assign y1405 = ~n5469 ;
  assign y1406 = ~1'b0 ;
  assign y1407 = n5474 ;
  assign y1408 = n5475 ;
  assign y1409 = ~1'b0 ;
  assign y1410 = n5479 ;
  assign y1411 = n5482 ;
  assign y1412 = ~n3079 ;
  assign y1413 = ~1'b0 ;
  assign y1414 = ~n5485 ;
  assign y1415 = ~n5486 ;
  assign y1416 = ~1'b0 ;
  assign y1417 = n5502 ;
  assign y1418 = n5510 ;
  assign y1419 = ~n5515 ;
  assign y1420 = n5524 ;
  assign y1421 = n5527 ;
  assign y1422 = n5532 ;
  assign y1423 = n5539 ;
  assign y1424 = n5540 ;
  assign y1425 = n1332 ;
  assign y1426 = n5543 ;
  assign y1427 = ~n5546 ;
  assign y1428 = ~n5560 ;
  assign y1429 = 1'b0 ;
  assign y1430 = ~1'b0 ;
  assign y1431 = ~n5561 ;
  assign y1432 = n5566 ;
  assign y1433 = n5573 ;
  assign y1434 = n5576 ;
  assign y1435 = n5577 ;
  assign y1436 = n5581 ;
  assign y1437 = ~n5582 ;
  assign y1438 = n5590 ;
  assign y1439 = n5594 ;
  assign y1440 = n5595 ;
  assign y1441 = ~n5600 ;
  assign y1442 = ~1'b0 ;
  assign y1443 = ~n5609 ;
  assign y1444 = n5612 ;
  assign y1445 = ~1'b0 ;
  assign y1446 = n5620 ;
  assign y1447 = n5624 ;
  assign y1448 = ~n5625 ;
  assign y1449 = ~n5633 ;
  assign y1450 = ~n5634 ;
  assign y1451 = n5639 ;
  assign y1452 = ~n5643 ;
  assign y1453 = ~n5654 ;
  assign y1454 = ~n5655 ;
  assign y1455 = ~n5656 ;
  assign y1456 = n5660 ;
  assign y1457 = n5663 ;
  assign y1458 = ~n5665 ;
  assign y1459 = n5667 ;
  assign y1460 = ~1'b0 ;
  assign y1461 = ~n4767 ;
  assign y1462 = ~1'b0 ;
  assign y1463 = n5671 ;
  assign y1464 = n5681 ;
  assign y1465 = ~n5683 ;
  assign y1466 = ~n5684 ;
  assign y1467 = n5687 ;
  assign y1468 = ~n5689 ;
  assign y1469 = ~n5702 ;
  assign y1470 = ~n5703 ;
  assign y1471 = ~n5704 ;
  assign y1472 = ~n5705 ;
  assign y1473 = ~1'b0 ;
  assign y1474 = n5709 ;
  assign y1475 = n5711 ;
  assign y1476 = n5715 ;
  assign y1477 = n5716 ;
  assign y1478 = ~n5718 ;
  assign y1479 = ~n5724 ;
  assign y1480 = ~n5733 ;
  assign y1481 = n5737 ;
  assign y1482 = ~1'b0 ;
  assign y1483 = ~n5743 ;
  assign y1484 = ~n5744 ;
  assign y1485 = ~n5745 ;
  assign y1486 = ~1'b0 ;
  assign y1487 = n5750 ;
  assign y1488 = ~n5752 ;
  assign y1489 = ~n1887 ;
  assign y1490 = n5760 ;
  assign y1491 = n5761 ;
  assign y1492 = ~n5763 ;
  assign y1493 = ~n5766 ;
  assign y1494 = ~n5767 ;
  assign y1495 = ~n5770 ;
  assign y1496 = n5782 ;
  assign y1497 = 1'b0 ;
  assign y1498 = n5785 ;
  assign y1499 = n5786 ;
  assign y1500 = ~n5787 ;
  assign y1501 = n5788 ;
  assign y1502 = ~n5794 ;
  assign y1503 = ~n5798 ;
  assign y1504 = ~n5804 ;
  assign y1505 = n5809 ;
  assign y1506 = n5810 ;
  assign y1507 = ~n5813 ;
  assign y1508 = n5821 ;
  assign y1509 = n5828 ;
  assign y1510 = n5829 ;
  assign y1511 = n5831 ;
  assign y1512 = n5834 ;
  assign y1513 = ~n5836 ;
  assign y1514 = ~n5838 ;
  assign y1515 = ~n5839 ;
  assign y1516 = ~n5841 ;
  assign y1517 = n5860 ;
  assign y1518 = ~n5861 ;
  assign y1519 = n5873 ;
  assign y1520 = ~1'b0 ;
  assign y1521 = ~n5875 ;
  assign y1522 = ~n5877 ;
  assign y1523 = n5881 ;
  assign y1524 = ~n5887 ;
  assign y1525 = ~1'b0 ;
  assign y1526 = ~n5889 ;
  assign y1527 = n5890 ;
  assign y1528 = ~n2179 ;
  assign y1529 = n5902 ;
  assign y1530 = ~n5910 ;
  assign y1531 = ~1'b0 ;
  assign y1532 = ~n5913 ;
  assign y1533 = n5917 ;
  assign y1534 = ~n5923 ;
  assign y1535 = n5927 ;
  assign y1536 = n5928 ;
  assign y1537 = ~1'b0 ;
  assign y1538 = n5937 ;
  assign y1539 = n5942 ;
  assign y1540 = ~n5944 ;
  assign y1541 = ~n5952 ;
  assign y1542 = ~n5957 ;
  assign y1543 = n5963 ;
  assign y1544 = n5967 ;
  assign y1545 = ~n5973 ;
  assign y1546 = ~n5979 ;
  assign y1547 = ~n5987 ;
  assign y1548 = n5989 ;
  assign y1549 = ~n5991 ;
  assign y1550 = n5995 ;
  assign y1551 = ~n5996 ;
  assign y1552 = ~n6003 ;
  assign y1553 = n6007 ;
  assign y1554 = ~1'b0 ;
  assign y1555 = ~n6010 ;
  assign y1556 = ~n6011 ;
  assign y1557 = ~n6026 ;
  assign y1558 = ~1'b0 ;
  assign y1559 = ~1'b0 ;
  assign y1560 = ~n6030 ;
  assign y1561 = n6031 ;
  assign y1562 = ~1'b0 ;
  assign y1563 = n6032 ;
  assign y1564 = ~n6035 ;
  assign y1565 = ~n6044 ;
  assign y1566 = ~n6047 ;
  assign y1567 = ~1'b0 ;
  assign y1568 = n6049 ;
  assign y1569 = n6051 ;
  assign y1570 = n6052 ;
  assign y1571 = ~n6056 ;
  assign y1572 = ~n6058 ;
  assign y1573 = n6064 ;
  assign y1574 = n6066 ;
  assign y1575 = n6068 ;
  assign y1576 = ~n6075 ;
  assign y1577 = ~n6080 ;
  assign y1578 = ~n6081 ;
  assign y1579 = ~n6086 ;
  assign y1580 = ~1'b0 ;
  assign y1581 = n6090 ;
  assign y1582 = ~n6097 ;
  assign y1583 = ~n6099 ;
  assign y1584 = ~n6111 ;
  assign y1585 = ~n6116 ;
  assign y1586 = ~n6119 ;
  assign y1587 = ~1'b0 ;
  assign y1588 = n6121 ;
  assign y1589 = ~n6122 ;
  assign y1590 = n6124 ;
  assign y1591 = ~n6126 ;
  assign y1592 = n6130 ;
  assign y1593 = ~n6131 ;
  assign y1594 = ~n6134 ;
  assign y1595 = ~n6138 ;
  assign y1596 = ~n6150 ;
  assign y1597 = ~n6154 ;
  assign y1598 = ~n6158 ;
  assign y1599 = n6162 ;
  assign y1600 = n6166 ;
  assign y1601 = ~1'b0 ;
  assign y1602 = ~n6169 ;
  assign y1603 = n6171 ;
  assign y1604 = ~n6172 ;
  assign y1605 = ~n6179 ;
  assign y1606 = n6182 ;
  assign y1607 = n6185 ;
  assign y1608 = ~1'b0 ;
  assign y1609 = n6194 ;
  assign y1610 = ~n6203 ;
  assign y1611 = n6206 ;
  assign y1612 = ~n6216 ;
  assign y1613 = n6224 ;
  assign y1614 = ~x104 ;
  assign y1615 = n6228 ;
  assign y1616 = n6243 ;
  assign y1617 = n6252 ;
  assign y1618 = n6256 ;
  assign y1619 = ~n6259 ;
  assign y1620 = ~n6264 ;
  assign y1621 = ~n6274 ;
  assign y1622 = n6275 ;
  assign y1623 = ~n6280 ;
  assign y1624 = ~1'b0 ;
  assign y1625 = ~n6287 ;
  assign y1626 = ~n6288 ;
  assign y1627 = ~1'b0 ;
  assign y1628 = ~n6289 ;
  assign y1629 = ~n6304 ;
  assign y1630 = n6311 ;
  assign y1631 = n6315 ;
  assign y1632 = ~n6322 ;
  assign y1633 = ~n6323 ;
  assign y1634 = ~1'b0 ;
  assign y1635 = n6334 ;
  assign y1636 = ~n6337 ;
  assign y1637 = ~n6338 ;
  assign y1638 = n6339 ;
  assign y1639 = ~1'b0 ;
  assign y1640 = n6350 ;
  assign y1641 = ~n6360 ;
  assign y1642 = ~n6361 ;
  assign y1643 = n6364 ;
  assign y1644 = ~n6366 ;
  assign y1645 = ~n6370 ;
  assign y1646 = n6375 ;
  assign y1647 = n6386 ;
  assign y1648 = n6389 ;
  assign y1649 = ~n6390 ;
  assign y1650 = ~n6391 ;
  assign y1651 = n6394 ;
  assign y1652 = n6395 ;
  assign y1653 = n6396 ;
  assign y1654 = ~1'b0 ;
  assign y1655 = n6416 ;
  assign y1656 = n6417 ;
  assign y1657 = n6420 ;
  assign y1658 = n6431 ;
  assign y1659 = ~1'b0 ;
  assign y1660 = ~n6436 ;
  assign y1661 = n6445 ;
  assign y1662 = ~n2911 ;
  assign y1663 = n6448 ;
  assign y1664 = n6453 ;
  assign y1665 = n6458 ;
  assign y1666 = ~n6467 ;
  assign y1667 = n6475 ;
  assign y1668 = n6478 ;
  assign y1669 = ~n6488 ;
  assign y1670 = n6489 ;
  assign y1671 = n6493 ;
  assign y1672 = n6505 ;
  assign y1673 = ~n6512 ;
  assign y1674 = ~n6515 ;
  assign y1675 = ~1'b0 ;
  assign y1676 = ~n6517 ;
  assign y1677 = ~n6520 ;
  assign y1678 = n6527 ;
  assign y1679 = ~1'b0 ;
  assign y1680 = ~n6528 ;
  assign y1681 = ~n6531 ;
  assign y1682 = n6534 ;
  assign y1683 = ~n6545 ;
  assign y1684 = n6548 ;
  assign y1685 = ~n6553 ;
  assign y1686 = n6560 ;
  assign y1687 = n6561 ;
  assign y1688 = n6573 ;
  assign y1689 = ~n6574 ;
  assign y1690 = n6576 ;
  assign y1691 = ~1'b0 ;
  assign y1692 = ~n6578 ;
  assign y1693 = n6581 ;
  assign y1694 = n6584 ;
  assign y1695 = ~n6599 ;
  assign y1696 = n6600 ;
  assign y1697 = n6601 ;
  assign y1698 = n6605 ;
  assign y1699 = n6607 ;
  assign y1700 = ~n6610 ;
  assign y1701 = ~n6611 ;
  assign y1702 = n6614 ;
  assign y1703 = n6621 ;
  assign y1704 = ~n6624 ;
  assign y1705 = ~n6630 ;
  assign y1706 = n6633 ;
  assign y1707 = ~n6637 ;
  assign y1708 = n6642 ;
  assign y1709 = ~n6652 ;
  assign y1710 = ~1'b0 ;
  assign y1711 = n6653 ;
  assign y1712 = n6655 ;
  assign y1713 = ~1'b0 ;
  assign y1714 = ~n6657 ;
  assign y1715 = n6662 ;
  assign y1716 = n6663 ;
  assign y1717 = n6668 ;
  assign y1718 = n6677 ;
  assign y1719 = n6683 ;
  assign y1720 = ~n6684 ;
  assign y1721 = ~n6685 ;
  assign y1722 = ~1'b0 ;
  assign y1723 = n6686 ;
  assign y1724 = n6687 ;
  assign y1725 = n6689 ;
  assign y1726 = ~n6696 ;
  assign y1727 = ~1'b0 ;
  assign y1728 = n6698 ;
  assign y1729 = ~n6705 ;
  assign y1730 = n6706 ;
  assign y1731 = ~n6709 ;
  assign y1732 = ~n6711 ;
  assign y1733 = n6718 ;
  assign y1734 = n6721 ;
  assign y1735 = ~n6722 ;
  assign y1736 = n6727 ;
  assign y1737 = ~n6733 ;
  assign y1738 = ~n6738 ;
  assign y1739 = ~n6740 ;
  assign y1740 = ~1'b0 ;
  assign y1741 = ~n6743 ;
  assign y1742 = ~n2982 ;
  assign y1743 = ~n6748 ;
  assign y1744 = n6749 ;
  assign y1745 = ~1'b0 ;
  assign y1746 = n6752 ;
  assign y1747 = ~n6757 ;
  assign y1748 = ~n6758 ;
  assign y1749 = n6761 ;
  assign y1750 = ~n6768 ;
  assign y1751 = n6771 ;
  assign y1752 = n6774 ;
  assign y1753 = ~n6787 ;
  assign y1754 = n6792 ;
  assign y1755 = ~n6797 ;
  assign y1756 = ~n6798 ;
  assign y1757 = n6799 ;
  assign y1758 = n6806 ;
  assign y1759 = ~1'b0 ;
  assign y1760 = ~1'b0 ;
  assign y1761 = n6808 ;
  assign y1762 = ~n6816 ;
  assign y1763 = ~n6819 ;
  assign y1764 = ~n6823 ;
  assign y1765 = ~n6825 ;
  assign y1766 = n6833 ;
  assign y1767 = ~n6834 ;
  assign y1768 = n6837 ;
  assign y1769 = n6839 ;
  assign y1770 = ~1'b0 ;
  assign y1771 = n6841 ;
  assign y1772 = n6844 ;
  assign y1773 = n6851 ;
  assign y1774 = ~n6855 ;
  assign y1775 = n6856 ;
  assign y1776 = ~n6859 ;
  assign y1777 = ~n6867 ;
  assign y1778 = ~n6872 ;
  assign y1779 = ~n6873 ;
  assign y1780 = n6875 ;
  assign y1781 = n6878 ;
  assign y1782 = ~n6880 ;
  assign y1783 = n6889 ;
  assign y1784 = ~n6898 ;
  assign y1785 = ~n6907 ;
  assign y1786 = ~n6910 ;
  assign y1787 = ~n6911 ;
  assign y1788 = ~n6919 ;
  assign y1789 = ~1'b0 ;
  assign y1790 = n6920 ;
  assign y1791 = ~1'b0 ;
  assign y1792 = ~n6921 ;
  assign y1793 = ~n6922 ;
  assign y1794 = n6924 ;
  assign y1795 = ~n6927 ;
  assign y1796 = n6936 ;
  assign y1797 = n6940 ;
  assign y1798 = ~n6948 ;
  assign y1799 = ~n6960 ;
  assign y1800 = n6961 ;
  assign y1801 = ~n6967 ;
  assign y1802 = n6982 ;
  assign y1803 = n6987 ;
  assign y1804 = ~1'b0 ;
  assign y1805 = n6996 ;
  assign y1806 = ~n7000 ;
  assign y1807 = n7004 ;
  assign y1808 = ~n7014 ;
  assign y1809 = ~n7015 ;
  assign y1810 = 1'b0 ;
  assign y1811 = ~n7017 ;
  assign y1812 = n7021 ;
  assign y1813 = ~n7022 ;
  assign y1814 = ~n7027 ;
  assign y1815 = n7035 ;
  assign y1816 = n7039 ;
  assign y1817 = ~n7043 ;
  assign y1818 = ~n7045 ;
  assign y1819 = ~n7050 ;
  assign y1820 = ~n7052 ;
  assign y1821 = n7058 ;
  assign y1822 = ~n7069 ;
  assign y1823 = ~n7076 ;
  assign y1824 = ~n7081 ;
  assign y1825 = ~n7083 ;
  assign y1826 = n7087 ;
  assign y1827 = n7091 ;
  assign y1828 = n7094 ;
  assign y1829 = ~n7111 ;
  assign y1830 = n7112 ;
  assign y1831 = ~n7120 ;
  assign y1832 = ~n7126 ;
  assign y1833 = n7132 ;
  assign y1834 = ~n7137 ;
  assign y1835 = ~n7138 ;
  assign y1836 = n7149 ;
  assign y1837 = ~n7157 ;
  assign y1838 = ~n7160 ;
  assign y1839 = ~n7175 ;
  assign y1840 = ~n7176 ;
  assign y1841 = ~n7178 ;
  assign y1842 = n7182 ;
  assign y1843 = ~n7185 ;
  assign y1844 = n7190 ;
  assign y1845 = n7194 ;
  assign y1846 = ~n7201 ;
  assign y1847 = ~1'b0 ;
  assign y1848 = n7203 ;
  assign y1849 = ~n7216 ;
  assign y1850 = n7222 ;
  assign y1851 = ~n7230 ;
  assign y1852 = n7233 ;
  assign y1853 = ~n7234 ;
  assign y1854 = ~1'b0 ;
  assign y1855 = ~1'b0 ;
  assign y1856 = n7238 ;
  assign y1857 = n7243 ;
  assign y1858 = ~n7249 ;
  assign y1859 = ~n7271 ;
  assign y1860 = ~n7281 ;
  assign y1861 = ~n7285 ;
  assign y1862 = n7286 ;
  assign y1863 = n7291 ;
  assign y1864 = ~n7293 ;
  assign y1865 = n7294 ;
  assign y1866 = ~1'b0 ;
  assign y1867 = ~n7296 ;
  assign y1868 = ~1'b0 ;
  assign y1869 = n7298 ;
  assign y1870 = ~n7300 ;
  assign y1871 = ~n7306 ;
  assign y1872 = n7309 ;
  assign y1873 = ~1'b0 ;
  assign y1874 = n7326 ;
  assign y1875 = n7327 ;
  assign y1876 = ~n7332 ;
  assign y1877 = n7333 ;
  assign y1878 = ~n7334 ;
  assign y1879 = n7336 ;
  assign y1880 = ~1'b0 ;
  assign y1881 = ~n7339 ;
  assign y1882 = ~1'b0 ;
  assign y1883 = n7345 ;
  assign y1884 = ~n7350 ;
  assign y1885 = ~n7362 ;
  assign y1886 = n7363 ;
  assign y1887 = n7368 ;
  assign y1888 = n7370 ;
  assign y1889 = n7374 ;
  assign y1890 = n7375 ;
  assign y1891 = ~1'b0 ;
  assign y1892 = ~n7378 ;
  assign y1893 = n7380 ;
  assign y1894 = n7385 ;
  assign y1895 = ~n7386 ;
  assign y1896 = ~1'b0 ;
  assign y1897 = ~n7391 ;
  assign y1898 = ~1'b0 ;
  assign y1899 = n7392 ;
  assign y1900 = n7404 ;
  assign y1901 = ~n7412 ;
  assign y1902 = ~n7416 ;
  assign y1903 = ~n7417 ;
  assign y1904 = ~n7418 ;
  assign y1905 = ~n7419 ;
  assign y1906 = ~n7423 ;
  assign y1907 = ~n7428 ;
  assign y1908 = n7431 ;
  assign y1909 = ~1'b0 ;
  assign y1910 = n7436 ;
  assign y1911 = n7447 ;
  assign y1912 = n7459 ;
  assign y1913 = ~1'b0 ;
  assign y1914 = n7460 ;
  assign y1915 = n7470 ;
  assign y1916 = n7475 ;
  assign y1917 = ~n3173 ;
  assign y1918 = ~1'b0 ;
  assign y1919 = n7492 ;
  assign y1920 = ~n7495 ;
  assign y1921 = n7496 ;
  assign y1922 = ~1'b0 ;
  assign y1923 = ~1'b0 ;
  assign y1924 = ~n7497 ;
  assign y1925 = ~n7502 ;
  assign y1926 = ~1'b0 ;
  assign y1927 = ~n7503 ;
  assign y1928 = n7504 ;
  assign y1929 = n7506 ;
  assign y1930 = ~n7510 ;
  assign y1931 = ~n7513 ;
  assign y1932 = ~n7515 ;
  assign y1933 = ~n7522 ;
  assign y1934 = n7524 ;
  assign y1935 = ~n7525 ;
  assign y1936 = n7527 ;
  assign y1937 = n7531 ;
  assign y1938 = ~n7533 ;
  assign y1939 = ~n7538 ;
  assign y1940 = n7545 ;
  assign y1941 = n7552 ;
  assign y1942 = n7558 ;
  assign y1943 = n7560 ;
  assign y1944 = n7570 ;
  assign y1945 = ~1'b0 ;
  assign y1946 = ~n7587 ;
  assign y1947 = n7590 ;
  assign y1948 = n7592 ;
  assign y1949 = n7594 ;
  assign y1950 = n7599 ;
  assign y1951 = n7605 ;
  assign y1952 = n7607 ;
  assign y1953 = n7609 ;
  assign y1954 = ~n7618 ;
  assign y1955 = ~1'b0 ;
  assign y1956 = n7624 ;
  assign y1957 = n7638 ;
  assign y1958 = ~1'b0 ;
  assign y1959 = ~1'b0 ;
  assign y1960 = n7645 ;
  assign y1961 = ~n7647 ;
  assign y1962 = ~1'b0 ;
  assign y1963 = n7653 ;
  assign y1964 = ~n7657 ;
  assign y1965 = n7664 ;
  assign y1966 = n7665 ;
  assign y1967 = ~n7668 ;
  assign y1968 = ~1'b0 ;
  assign y1969 = ~n7669 ;
  assign y1970 = n1441 ;
  assign y1971 = n7670 ;
  assign y1972 = ~n7673 ;
  assign y1973 = ~n7682 ;
  assign y1974 = ~n7687 ;
  assign y1975 = ~n7688 ;
  assign y1976 = ~n7690 ;
  assign y1977 = ~n7699 ;
  assign y1978 = ~1'b0 ;
  assign y1979 = ~n7705 ;
  assign y1980 = ~n7708 ;
  assign y1981 = n7713 ;
  assign y1982 = n7719 ;
  assign y1983 = ~1'b0 ;
  assign y1984 = n7720 ;
  assign y1985 = n7731 ;
  assign y1986 = n7732 ;
  assign y1987 = ~n7740 ;
  assign y1988 = ~1'b0 ;
  assign y1989 = ~n7743 ;
  assign y1990 = n7744 ;
  assign y1991 = ~n7750 ;
  assign y1992 = ~n7758 ;
  assign y1993 = ~n7760 ;
  assign y1994 = ~n7762 ;
  assign y1995 = n7763 ;
  assign y1996 = ~n7768 ;
  assign y1997 = n3620 ;
  assign y1998 = ~n7775 ;
  assign y1999 = n7778 ;
  assign y2000 = ~n7795 ;
  assign y2001 = n7797 ;
  assign y2002 = n7802 ;
  assign y2003 = ~1'b0 ;
  assign y2004 = ~n7806 ;
  assign y2005 = ~n7813 ;
  assign y2006 = n7826 ;
  assign y2007 = ~n7829 ;
  assign y2008 = n7834 ;
  assign y2009 = n7840 ;
  assign y2010 = n7846 ;
  assign y2011 = ~n7851 ;
  assign y2012 = n7852 ;
  assign y2013 = ~n7853 ;
  assign y2014 = ~n7854 ;
  assign y2015 = n7857 ;
  assign y2016 = n7864 ;
  assign y2017 = ~n7866 ;
  assign y2018 = n2619 ;
  assign y2019 = n7869 ;
  assign y2020 = n7871 ;
  assign y2021 = n7874 ;
  assign y2022 = ~n7875 ;
  assign y2023 = ~n7878 ;
  assign y2024 = ~n7883 ;
  assign y2025 = n7885 ;
  assign y2026 = n7886 ;
  assign y2027 = n7889 ;
  assign y2028 = ~n7900 ;
  assign y2029 = ~1'b0 ;
  assign y2030 = ~1'b0 ;
  assign y2031 = ~n7902 ;
  assign y2032 = n7910 ;
  assign y2033 = ~n7914 ;
  assign y2034 = ~n7921 ;
  assign y2035 = ~n7923 ;
  assign y2036 = n7925 ;
  assign y2037 = n7937 ;
  assign y2038 = ~n7946 ;
  assign y2039 = ~1'b0 ;
  assign y2040 = ~n7948 ;
  assign y2041 = ~n7959 ;
  assign y2042 = ~n7968 ;
  assign y2043 = n7973 ;
  assign y2044 = ~n7975 ;
  assign y2045 = ~n7977 ;
  assign y2046 = n7980 ;
  assign y2047 = ~n7981 ;
  assign y2048 = ~n7986 ;
  assign y2049 = ~n7995 ;
  assign y2050 = ~n7996 ;
  assign y2051 = n8006 ;
  assign y2052 = n8016 ;
  assign y2053 = ~n8019 ;
  assign y2054 = ~n8022 ;
  assign y2055 = ~n8030 ;
  assign y2056 = n8033 ;
  assign y2057 = ~1'b0 ;
  assign y2058 = ~1'b0 ;
  assign y2059 = 1'b0 ;
  assign y2060 = n8034 ;
  assign y2061 = ~n8051 ;
  assign y2062 = ~1'b0 ;
  assign y2063 = ~n8069 ;
  assign y2064 = ~n8079 ;
  assign y2065 = ~1'b0 ;
  assign y2066 = ~n8081 ;
  assign y2067 = ~n8082 ;
  assign y2068 = ~n8083 ;
  assign y2069 = ~n8089 ;
  assign y2070 = ~n8092 ;
  assign y2071 = ~1'b0 ;
  assign y2072 = ~n8104 ;
  assign y2073 = ~n8105 ;
  assign y2074 = ~n8110 ;
  assign y2075 = ~n8113 ;
  assign y2076 = ~n8114 ;
  assign y2077 = n8123 ;
  assign y2078 = n8131 ;
  assign y2079 = n8142 ;
  assign y2080 = ~n8144 ;
  assign y2081 = ~1'b0 ;
  assign y2082 = n8147 ;
  assign y2083 = ~n8148 ;
  assign y2084 = n8149 ;
  assign y2085 = n8154 ;
  assign y2086 = n8157 ;
  assign y2087 = ~1'b0 ;
  assign y2088 = n8158 ;
  assign y2089 = ~n8159 ;
  assign y2090 = ~1'b0 ;
  assign y2091 = n8163 ;
  assign y2092 = ~1'b0 ;
  assign y2093 = n8165 ;
  assign y2094 = ~n8166 ;
  assign y2095 = ~n8169 ;
  assign y2096 = ~1'b0 ;
  assign y2097 = ~n8171 ;
  assign y2098 = n8176 ;
  assign y2099 = ~n8178 ;
  assign y2100 = ~n8180 ;
  assign y2101 = ~n8181 ;
  assign y2102 = n8187 ;
  assign y2103 = ~n8197 ;
  assign y2104 = n8200 ;
  assign y2105 = n8207 ;
  assign y2106 = ~n8210 ;
  assign y2107 = ~1'b0 ;
  assign y2108 = ~n8211 ;
  assign y2109 = ~n8214 ;
  assign y2110 = ~n8217 ;
  assign y2111 = ~n8222 ;
  assign y2112 = ~1'b0 ;
  assign y2113 = n8225 ;
  assign y2114 = ~n8233 ;
  assign y2115 = n8237 ;
  assign y2116 = n8241 ;
  assign y2117 = ~1'b0 ;
  assign y2118 = n8246 ;
  assign y2119 = n8257 ;
  assign y2120 = ~n8260 ;
  assign y2121 = ~n8273 ;
  assign y2122 = n8275 ;
  assign y2123 = n8283 ;
  assign y2124 = n8285 ;
  assign y2125 = ~1'b0 ;
  assign y2126 = ~1'b0 ;
  assign y2127 = ~n8286 ;
  assign y2128 = n8296 ;
  assign y2129 = ~n8308 ;
  assign y2130 = n8310 ;
  assign y2131 = ~1'b0 ;
  assign y2132 = ~n8312 ;
  assign y2133 = n8316 ;
  assign y2134 = n8319 ;
  assign y2135 = ~n8321 ;
  assign y2136 = n8324 ;
  assign y2137 = ~1'b0 ;
  assign y2138 = n8327 ;
  assign y2139 = ~n8339 ;
  assign y2140 = ~n8346 ;
  assign y2141 = ~n8350 ;
  assign y2142 = n8351 ;
  assign y2143 = ~1'b0 ;
  assign y2144 = ~n8360 ;
  assign y2145 = n8362 ;
  assign y2146 = n8364 ;
  assign y2147 = n8371 ;
  assign y2148 = ~1'b0 ;
  assign y2149 = n8378 ;
  assign y2150 = n8382 ;
  assign y2151 = ~n8386 ;
  assign y2152 = n2377 ;
  assign y2153 = ~n8387 ;
  assign y2154 = n8388 ;
  assign y2155 = ~n8389 ;
  assign y2156 = ~n8399 ;
  assign y2157 = ~n8404 ;
  assign y2158 = n8417 ;
  assign y2159 = ~n8436 ;
  assign y2160 = n8441 ;
  assign y2161 = n8444 ;
  assign y2162 = ~1'b0 ;
  assign y2163 = n8447 ;
  assign y2164 = ~n8449 ;
  assign y2165 = n8450 ;
  assign y2166 = ~n5062 ;
  assign y2167 = ~n8451 ;
  assign y2168 = ~n8457 ;
  assign y2169 = n8460 ;
  assign y2170 = ~n8471 ;
  assign y2171 = ~n8473 ;
  assign y2172 = n8474 ;
  assign y2173 = ~1'b0 ;
  assign y2174 = n8478 ;
  assign y2175 = ~1'b0 ;
  assign y2176 = ~1'b0 ;
  assign y2177 = ~n8481 ;
  assign y2178 = 1'b0 ;
  assign y2179 = n8483 ;
  assign y2180 = ~1'b0 ;
  assign y2181 = ~1'b0 ;
  assign y2182 = ~n8485 ;
  assign y2183 = n8489 ;
  assign y2184 = ~1'b0 ;
  assign y2185 = n8502 ;
  assign y2186 = ~1'b0 ;
  assign y2187 = ~1'b0 ;
  assign y2188 = n8511 ;
  assign y2189 = n8513 ;
  assign y2190 = ~1'b0 ;
  assign y2191 = ~n8514 ;
  assign y2192 = n8518 ;
  assign y2193 = n8520 ;
  assign y2194 = ~n8523 ;
  assign y2195 = ~n8530 ;
  assign y2196 = n8532 ;
  assign y2197 = ~1'b0 ;
  assign y2198 = n8535 ;
  assign y2199 = ~n8547 ;
  assign y2200 = ~n8554 ;
  assign y2201 = ~n8560 ;
  assign y2202 = ~1'b0 ;
  assign y2203 = n8567 ;
  assign y2204 = ~n8573 ;
  assign y2205 = n8575 ;
  assign y2206 = n8576 ;
  assign y2207 = ~n8580 ;
  assign y2208 = ~1'b0 ;
  assign y2209 = n8586 ;
  assign y2210 = ~n8589 ;
  assign y2211 = ~n8590 ;
  assign y2212 = n8591 ;
  assign y2213 = ~n8595 ;
  assign y2214 = ~1'b0 ;
  assign y2215 = ~1'b0 ;
  assign y2216 = ~n8596 ;
  assign y2217 = n8600 ;
  assign y2218 = ~n8603 ;
  assign y2219 = ~n8609 ;
  assign y2220 = ~n8613 ;
  assign y2221 = n8621 ;
  assign y2222 = n8624 ;
  assign y2223 = ~1'b0 ;
  assign y2224 = ~1'b0 ;
  assign y2225 = n8627 ;
  assign y2226 = n8628 ;
  assign y2227 = ~n8631 ;
  assign y2228 = ~1'b0 ;
  assign y2229 = ~n8637 ;
  assign y2230 = n8638 ;
  assign y2231 = ~n8639 ;
  assign y2232 = ~n8643 ;
  assign y2233 = n8646 ;
  assign y2234 = ~1'b0 ;
  assign y2235 = ~n8649 ;
  assign y2236 = ~n8650 ;
  assign y2237 = ~n8655 ;
  assign y2238 = n8657 ;
  assign y2239 = n8665 ;
  assign y2240 = ~n8666 ;
  assign y2241 = n8668 ;
  assign y2242 = ~1'b0 ;
  assign y2243 = ~n8672 ;
  assign y2244 = ~n8675 ;
  assign y2245 = n8683 ;
  assign y2246 = ~n8685 ;
  assign y2247 = ~1'b0 ;
  assign y2248 = n8689 ;
  assign y2249 = ~n8695 ;
  assign y2250 = n8698 ;
  assign y2251 = n8700 ;
  assign y2252 = ~n8705 ;
  assign y2253 = n8708 ;
  assign y2254 = ~1'b0 ;
  assign y2255 = ~1'b0 ;
  assign y2256 = n8716 ;
  assign y2257 = n8722 ;
  assign y2258 = ~n8724 ;
  assign y2259 = n8728 ;
  assign y2260 = ~n8733 ;
  assign y2261 = ~n8735 ;
  assign y2262 = ~n8744 ;
  assign y2263 = ~n8746 ;
  assign y2264 = ~n8750 ;
  assign y2265 = ~1'b0 ;
  assign y2266 = ~n8752 ;
  assign y2267 = ~n8755 ;
  assign y2268 = ~n8756 ;
  assign y2269 = n8760 ;
  assign y2270 = n8762 ;
  assign y2271 = ~n8764 ;
  assign y2272 = n8769 ;
  assign y2273 = n8770 ;
  assign y2274 = n8774 ;
  assign y2275 = n8777 ;
  assign y2276 = n8782 ;
  assign y2277 = ~n8796 ;
  assign y2278 = n8798 ;
  assign y2279 = ~n8799 ;
  assign y2280 = ~n8800 ;
  assign y2281 = n8801 ;
  assign y2282 = ~1'b0 ;
  assign y2283 = ~n8804 ;
  assign y2284 = n8808 ;
  assign y2285 = n8810 ;
  assign y2286 = ~n8813 ;
  assign y2287 = n8818 ;
  assign y2288 = ~n8819 ;
  assign y2289 = ~n8823 ;
  assign y2290 = n8830 ;
  assign y2291 = n8837 ;
  assign y2292 = ~n8838 ;
  assign y2293 = n8839 ;
  assign y2294 = ~1'b0 ;
  assign y2295 = ~n8841 ;
  assign y2296 = ~n8846 ;
  assign y2297 = ~1'b0 ;
  assign y2298 = n8851 ;
  assign y2299 = ~n8856 ;
  assign y2300 = ~1'b0 ;
  assign y2301 = ~1'b0 ;
  assign y2302 = n8860 ;
  assign y2303 = ~n8862 ;
  assign y2304 = ~n8863 ;
  assign y2305 = ~n4663 ;
  assign y2306 = ~n8865 ;
  assign y2307 = n8866 ;
  assign y2308 = n8867 ;
  assign y2309 = n8872 ;
  assign y2310 = ~n8873 ;
  assign y2311 = n8880 ;
  assign y2312 = ~n8881 ;
  assign y2313 = ~n8884 ;
  assign y2314 = n8885 ;
  assign y2315 = ~n8891 ;
  assign y2316 = n8892 ;
  assign y2317 = ~1'b0 ;
  assign y2318 = n8904 ;
  assign y2319 = ~1'b0 ;
  assign y2320 = ~n8905 ;
  assign y2321 = ~n8906 ;
  assign y2322 = ~1'b0 ;
  assign y2323 = ~n8913 ;
  assign y2324 = n8917 ;
  assign y2325 = ~n8928 ;
  assign y2326 = ~n8929 ;
  assign y2327 = n8930 ;
  assign y2328 = ~n8938 ;
  assign y2329 = ~n8942 ;
  assign y2330 = n8962 ;
  assign y2331 = ~n8963 ;
  assign y2332 = ~n8966 ;
  assign y2333 = ~n8968 ;
  assign y2334 = ~n8974 ;
  assign y2335 = ~n8979 ;
  assign y2336 = ~n8987 ;
  assign y2337 = ~1'b0 ;
  assign y2338 = n8988 ;
  assign y2339 = n8993 ;
  assign y2340 = n8995 ;
  assign y2341 = n8999 ;
  assign y2342 = ~1'b0 ;
  assign y2343 = ~1'b0 ;
  assign y2344 = ~n9002 ;
  assign y2345 = n9009 ;
  assign y2346 = n9012 ;
  assign y2347 = ~n9014 ;
  assign y2348 = ~n9019 ;
  assign y2349 = ~n9025 ;
  assign y2350 = n9026 ;
  assign y2351 = ~n9027 ;
  assign y2352 = n9029 ;
  assign y2353 = ~1'b0 ;
  assign y2354 = ~n9041 ;
  assign y2355 = ~n9048 ;
  assign y2356 = ~n9050 ;
  assign y2357 = n9051 ;
  assign y2358 = ~n9052 ;
  assign y2359 = ~n9053 ;
  assign y2360 = ~n9055 ;
  assign y2361 = ~n9068 ;
  assign y2362 = ~1'b0 ;
  assign y2363 = n9072 ;
  assign y2364 = 1'b0 ;
  assign y2365 = n9084 ;
  assign y2366 = n9090 ;
  assign y2367 = n9103 ;
  assign y2368 = ~n9112 ;
  assign y2369 = n9130 ;
  assign y2370 = ~n4585 ;
  assign y2371 = ~n9133 ;
  assign y2372 = ~n9137 ;
  assign y2373 = ~n9142 ;
  assign y2374 = n9154 ;
  assign y2375 = ~n9164 ;
  assign y2376 = ~n9179 ;
  assign y2377 = ~1'b0 ;
  assign y2378 = ~n9184 ;
  assign y2379 = n9190 ;
  assign y2380 = ~1'b0 ;
  assign y2381 = n9199 ;
  assign y2382 = ~1'b0 ;
  assign y2383 = n9202 ;
  assign y2384 = ~n9209 ;
  assign y2385 = ~n9213 ;
  assign y2386 = n9214 ;
  assign y2387 = ~1'b0 ;
  assign y2388 = ~n9216 ;
  assign y2389 = n9225 ;
  assign y2390 = ~n9227 ;
  assign y2391 = n9230 ;
  assign y2392 = n9231 ;
  assign y2393 = ~n9232 ;
  assign y2394 = ~n9233 ;
  assign y2395 = n9238 ;
  assign y2396 = n9239 ;
  assign y2397 = n9241 ;
  assign y2398 = ~n9243 ;
  assign y2399 = n9244 ;
  assign y2400 = ~1'b0 ;
  assign y2401 = ~n9246 ;
  assign y2402 = n2026 ;
  assign y2403 = ~n9249 ;
  assign y2404 = ~1'b0 ;
  assign y2405 = ~n9251 ;
  assign y2406 = ~n9252 ;
  assign y2407 = n9263 ;
  assign y2408 = n9265 ;
  assign y2409 = n9271 ;
  assign y2410 = n9274 ;
  assign y2411 = n9275 ;
  assign y2412 = n9280 ;
  assign y2413 = n9288 ;
  assign y2414 = ~n9291 ;
  assign y2415 = n9292 ;
  assign y2416 = n9296 ;
  assign y2417 = n9298 ;
  assign y2418 = n9299 ;
  assign y2419 = n9301 ;
  assign y2420 = n9302 ;
  assign y2421 = ~n9304 ;
  assign y2422 = n9307 ;
  assign y2423 = ~n9309 ;
  assign y2424 = n9311 ;
  assign y2425 = n9315 ;
  assign y2426 = ~n9318 ;
  assign y2427 = n9320 ;
  assign y2428 = n9328 ;
  assign y2429 = n9330 ;
  assign y2430 = ~n9334 ;
  assign y2431 = ~1'b0 ;
  assign y2432 = ~n9343 ;
  assign y2433 = ~n9348 ;
  assign y2434 = n9351 ;
  assign y2435 = ~n9355 ;
  assign y2436 = ~n9360 ;
  assign y2437 = ~n9365 ;
  assign y2438 = ~1'b0 ;
  assign y2439 = ~1'b0 ;
  assign y2440 = ~n9368 ;
  assign y2441 = ~n9373 ;
  assign y2442 = n9374 ;
  assign y2443 = ~n9375 ;
  assign y2444 = n9381 ;
  assign y2445 = n9383 ;
  assign y2446 = ~n9384 ;
  assign y2447 = ~1'b0 ;
  assign y2448 = ~n9386 ;
  assign y2449 = n9389 ;
  assign y2450 = ~n9390 ;
  assign y2451 = n9392 ;
  assign y2452 = n9396 ;
  assign y2453 = ~n9400 ;
  assign y2454 = n9402 ;
  assign y2455 = n9415 ;
  assign y2456 = n9418 ;
  assign y2457 = n9420 ;
  assign y2458 = ~n9424 ;
  assign y2459 = n9425 ;
  assign y2460 = n9428 ;
  assign y2461 = ~n9430 ;
  assign y2462 = ~n9433 ;
  assign y2463 = ~n9438 ;
  assign y2464 = ~1'b0 ;
  assign y2465 = n9441 ;
  assign y2466 = ~1'b0 ;
  assign y2467 = n9442 ;
  assign y2468 = ~n9454 ;
  assign y2469 = n9455 ;
  assign y2470 = ~n9456 ;
  assign y2471 = n9460 ;
  assign y2472 = ~n9464 ;
  assign y2473 = ~n9468 ;
  assign y2474 = ~n9475 ;
  assign y2475 = n9480 ;
  assign y2476 = ~n9483 ;
  assign y2477 = ~1'b0 ;
  assign y2478 = n9484 ;
  assign y2479 = n9486 ;
  assign y2480 = ~1'b0 ;
  assign y2481 = ~n9487 ;
  assign y2482 = ~n9488 ;
  assign y2483 = n9492 ;
  assign y2484 = ~n9496 ;
  assign y2485 = ~1'b0 ;
  assign y2486 = ~n9499 ;
  assign y2487 = ~n9500 ;
  assign y2488 = n9501 ;
  assign y2489 = n9508 ;
  assign y2490 = ~1'b0 ;
  assign y2491 = ~n9509 ;
  assign y2492 = ~n9514 ;
  assign y2493 = n9520 ;
  assign y2494 = n9521 ;
  assign y2495 = n9523 ;
  assign y2496 = ~n9524 ;
  assign y2497 = ~n9531 ;
  assign y2498 = ~n9535 ;
  assign y2499 = n9537 ;
  assign y2500 = n9541 ;
  assign y2501 = ~n9542 ;
  assign y2502 = ~n9544 ;
  assign y2503 = ~n9551 ;
  assign y2504 = ~n9556 ;
  assign y2505 = n9569 ;
  assign y2506 = ~n9572 ;
  assign y2507 = n9578 ;
  assign y2508 = n6540 ;
  assign y2509 = n9582 ;
  assign y2510 = ~n9583 ;
  assign y2511 = 1'b0 ;
  assign y2512 = ~n9598 ;
  assign y2513 = ~n9599 ;
  assign y2514 = ~n9604 ;
  assign y2515 = ~n9606 ;
  assign y2516 = n9615 ;
  assign y2517 = ~n9619 ;
  assign y2518 = n9624 ;
  assign y2519 = ~1'b0 ;
  assign y2520 = ~n5612 ;
  assign y2521 = n9635 ;
  assign y2522 = n9636 ;
  assign y2523 = n9643 ;
  assign y2524 = n9653 ;
  assign y2525 = n9658 ;
  assign y2526 = ~n9663 ;
  assign y2527 = ~1'b0 ;
  assign y2528 = ~n9666 ;
  assign y2529 = ~n9676 ;
  assign y2530 = ~1'b0 ;
  assign y2531 = n9688 ;
  assign y2532 = ~n9701 ;
  assign y2533 = n9703 ;
  assign y2534 = n9709 ;
  assign y2535 = ~n9714 ;
  assign y2536 = n3738 ;
  assign y2537 = n9715 ;
  assign y2538 = n9716 ;
  assign y2539 = n9718 ;
  assign y2540 = n9725 ;
  assign y2541 = n9727 ;
  assign y2542 = ~1'b0 ;
  assign y2543 = ~1'b0 ;
  assign y2544 = n9733 ;
  assign y2545 = ~n9738 ;
  assign y2546 = ~1'b0 ;
  assign y2547 = n9741 ;
  assign y2548 = n9744 ;
  assign y2549 = ~n9745 ;
  assign y2550 = n6697 ;
  assign y2551 = ~n9754 ;
  assign y2552 = n9757 ;
  assign y2553 = n9760 ;
  assign y2554 = ~n9762 ;
  assign y2555 = ~n9764 ;
  assign y2556 = ~n9773 ;
  assign y2557 = ~n9775 ;
  assign y2558 = ~n9778 ;
  assign y2559 = n9784 ;
  assign y2560 = ~n9786 ;
  assign y2561 = n9788 ;
  assign y2562 = n9808 ;
  assign y2563 = ~1'b0 ;
  assign y2564 = ~n9809 ;
  assign y2565 = ~n9816 ;
  assign y2566 = n9825 ;
  assign y2567 = n9826 ;
  assign y2568 = n9827 ;
  assign y2569 = ~1'b0 ;
  assign y2570 = ~n9838 ;
  assign y2571 = n9839 ;
  assign y2572 = ~1'b0 ;
  assign y2573 = n9843 ;
  assign y2574 = n9853 ;
  assign y2575 = ~n9854 ;
  assign y2576 = ~n9861 ;
  assign y2577 = ~n9863 ;
  assign y2578 = ~1'b0 ;
  assign y2579 = ~n9867 ;
  assign y2580 = ~1'b0 ;
  assign y2581 = n9869 ;
  assign y2582 = ~n9871 ;
  assign y2583 = n9877 ;
  assign y2584 = ~n9878 ;
  assign y2585 = n9882 ;
  assign y2586 = n9885 ;
  assign y2587 = ~n9888 ;
  assign y2588 = n9893 ;
  assign y2589 = ~n9899 ;
  assign y2590 = ~n9902 ;
  assign y2591 = n9903 ;
  assign y2592 = ~1'b0 ;
  assign y2593 = ~n9906 ;
  assign y2594 = n9907 ;
  assign y2595 = n9912 ;
  assign y2596 = n9913 ;
  assign y2597 = n9914 ;
  assign y2598 = ~n9918 ;
  assign y2599 = n9927 ;
  assign y2600 = ~n9929 ;
  assign y2601 = n9930 ;
  assign y2602 = ~n9940 ;
  assign y2603 = ~n9943 ;
  assign y2604 = ~n9951 ;
  assign y2605 = n9955 ;
  assign y2606 = ~n9956 ;
  assign y2607 = n9960 ;
  assign y2608 = n9973 ;
  assign y2609 = ~1'b0 ;
  assign y2610 = n9975 ;
  assign y2611 = ~n9976 ;
  assign y2612 = ~n9983 ;
  assign y2613 = ~n9984 ;
  assign y2614 = n9987 ;
  assign y2615 = n9989 ;
  assign y2616 = ~1'b0 ;
  assign y2617 = n9994 ;
  assign y2618 = n10000 ;
  assign y2619 = ~n10004 ;
  assign y2620 = ~1'b0 ;
  assign y2621 = ~n10006 ;
  assign y2622 = ~n10008 ;
  assign y2623 = ~n10011 ;
  assign y2624 = ~n10016 ;
  assign y2625 = ~n10026 ;
  assign y2626 = ~n3392 ;
  assign y2627 = ~n10029 ;
  assign y2628 = n10033 ;
  assign y2629 = n10036 ;
  assign y2630 = ~n10037 ;
  assign y2631 = ~n10045 ;
  assign y2632 = ~n10051 ;
  assign y2633 = n10053 ;
  assign y2634 = n10061 ;
  assign y2635 = n10063 ;
  assign y2636 = n10067 ;
  assign y2637 = n10075 ;
  assign y2638 = ~1'b0 ;
  assign y2639 = n10078 ;
  assign y2640 = ~n10082 ;
  assign y2641 = n10083 ;
  assign y2642 = ~n10094 ;
  assign y2643 = ~1'b0 ;
  assign y2644 = ~n10098 ;
  assign y2645 = n10099 ;
  assign y2646 = n10102 ;
  assign y2647 = n10103 ;
  assign y2648 = n10112 ;
  assign y2649 = ~1'b0 ;
  assign y2650 = ~n10118 ;
  assign y2651 = ~n10120 ;
  assign y2652 = ~n10127 ;
  assign y2653 = ~1'b0 ;
  assign y2654 = ~n10131 ;
  assign y2655 = ~1'b0 ;
  assign y2656 = ~n10140 ;
  assign y2657 = ~n10143 ;
  assign y2658 = ~n10147 ;
  assign y2659 = n10149 ;
  assign y2660 = n10150 ;
  assign y2661 = ~n10151 ;
  assign y2662 = ~1'b0 ;
  assign y2663 = ~n10152 ;
  assign y2664 = n2027 ;
  assign y2665 = ~n10157 ;
  assign y2666 = ~1'b0 ;
  assign y2667 = n10159 ;
  assign y2668 = ~n10164 ;
  assign y2669 = n10168 ;
  assign y2670 = n10172 ;
  assign y2671 = ~1'b0 ;
  assign y2672 = ~n10178 ;
  assign y2673 = n10179 ;
  assign y2674 = n10180 ;
  assign y2675 = ~n10181 ;
  assign y2676 = n10189 ;
  assign y2677 = n10195 ;
  assign y2678 = ~n10200 ;
  assign y2679 = n10205 ;
  assign y2680 = ~n10208 ;
  assign y2681 = n10214 ;
  assign y2682 = ~n10218 ;
  assign y2683 = ~1'b0 ;
  assign y2684 = ~1'b0 ;
  assign y2685 = ~n10220 ;
  assign y2686 = n10226 ;
  assign y2687 = ~n10235 ;
  assign y2688 = n10238 ;
  assign y2689 = n4331 ;
  assign y2690 = ~n10239 ;
  assign y2691 = n10242 ;
  assign y2692 = n10243 ;
  assign y2693 = ~n10244 ;
  assign y2694 = ~n10250 ;
  assign y2695 = ~n10255 ;
  assign y2696 = ~n10261 ;
  assign y2697 = ~n10264 ;
  assign y2698 = n10267 ;
  assign y2699 = n10272 ;
  assign y2700 = ~n10276 ;
  assign y2701 = ~n10284 ;
  assign y2702 = ~n10287 ;
  assign y2703 = ~1'b0 ;
  assign y2704 = ~n10289 ;
  assign y2705 = n10297 ;
  assign y2706 = n10300 ;
  assign y2707 = ~n10303 ;
  assign y2708 = n10307 ;
  assign y2709 = ~n10314 ;
  assign y2710 = ~n10315 ;
  assign y2711 = ~n10318 ;
  assign y2712 = n10319 ;
  assign y2713 = n10320 ;
  assign y2714 = ~n10331 ;
  assign y2715 = n10333 ;
  assign y2716 = ~n10343 ;
  assign y2717 = n10345 ;
  assign y2718 = ~n10349 ;
  assign y2719 = n10353 ;
  assign y2720 = ~n10354 ;
  assign y2721 = ~1'b0 ;
  assign y2722 = n10356 ;
  assign y2723 = n10358 ;
  assign y2724 = ~n10363 ;
  assign y2725 = n10369 ;
  assign y2726 = n10371 ;
  assign y2727 = n10372 ;
  assign y2728 = ~n10378 ;
  assign y2729 = ~n10380 ;
  assign y2730 = ~n10381 ;
  assign y2731 = ~1'b0 ;
  assign y2732 = ~n10385 ;
  assign y2733 = ~1'b0 ;
  assign y2734 = ~n10388 ;
  assign y2735 = ~n10389 ;
  assign y2736 = ~n10392 ;
  assign y2737 = ~1'b0 ;
  assign y2738 = ~1'b0 ;
  assign y2739 = ~n10393 ;
  assign y2740 = ~n10394 ;
  assign y2741 = ~n10395 ;
  assign y2742 = n10398 ;
  assign y2743 = n10399 ;
  assign y2744 = ~n10405 ;
  assign y2745 = n10419 ;
  assign y2746 = ~1'b0 ;
  assign y2747 = n10420 ;
  assign y2748 = ~1'b0 ;
  assign y2749 = ~1'b0 ;
  assign y2750 = n10421 ;
  assign y2751 = n10425 ;
  assign y2752 = n10427 ;
  assign y2753 = ~n10442 ;
  assign y2754 = n10443 ;
  assign y2755 = n10446 ;
  assign y2756 = n10452 ;
  assign y2757 = n10453 ;
  assign y2758 = n10454 ;
  assign y2759 = ~n10461 ;
  assign y2760 = ~n10462 ;
  assign y2761 = n10463 ;
  assign y2762 = ~n10468 ;
  assign y2763 = n10478 ;
  assign y2764 = n10480 ;
  assign y2765 = ~n10485 ;
  assign y2766 = n10491 ;
  assign y2767 = ~n10498 ;
  assign y2768 = ~n10499 ;
  assign y2769 = n10500 ;
  assign y2770 = n10508 ;
  assign y2771 = ~n10521 ;
  assign y2772 = ~n10523 ;
  assign y2773 = n10527 ;
  assign y2774 = n10532 ;
  assign y2775 = ~n10539 ;
  assign y2776 = ~n10540 ;
  assign y2777 = ~n10548 ;
  assign y2778 = n10550 ;
  assign y2779 = n10553 ;
  assign y2780 = ~n10557 ;
  assign y2781 = ~n10560 ;
  assign y2782 = ~1'b0 ;
  assign y2783 = ~n10574 ;
  assign y2784 = n10580 ;
  assign y2785 = n10583 ;
  assign y2786 = ~n10586 ;
  assign y2787 = ~n10588 ;
  assign y2788 = n10590 ;
  assign y2789 = ~1'b0 ;
  assign y2790 = n10591 ;
  assign y2791 = n10596 ;
  assign y2792 = ~n10600 ;
  assign y2793 = n10602 ;
  assign y2794 = n10604 ;
  assign y2795 = ~n10606 ;
  assign y2796 = n10611 ;
  assign y2797 = ~n10613 ;
  assign y2798 = ~n10614 ;
  assign y2799 = ~n10615 ;
  assign y2800 = n10617 ;
  assign y2801 = n10619 ;
  assign y2802 = ~n10622 ;
  assign y2803 = ~n10629 ;
  assign y2804 = ~n10630 ;
  assign y2805 = ~n10639 ;
  assign y2806 = n10648 ;
  assign y2807 = ~n10651 ;
  assign y2808 = n10653 ;
  assign y2809 = ~n1870 ;
  assign y2810 = ~n10660 ;
  assign y2811 = n10663 ;
  assign y2812 = n2628 ;
  assign y2813 = ~n10664 ;
  assign y2814 = ~1'b0 ;
  assign y2815 = n10669 ;
  assign y2816 = n10670 ;
  assign y2817 = n10672 ;
  assign y2818 = n10674 ;
  assign y2819 = ~n10681 ;
  assign y2820 = ~n10682 ;
  assign y2821 = n10683 ;
  assign y2822 = n10685 ;
  assign y2823 = ~1'b0 ;
  assign y2824 = n10692 ;
  assign y2825 = ~n10694 ;
  assign y2826 = n10699 ;
  assign y2827 = ~n10701 ;
  assign y2828 = n10712 ;
  assign y2829 = n10719 ;
  assign y2830 = ~n10732 ;
  assign y2831 = n10733 ;
  assign y2832 = ~n10736 ;
  assign y2833 = n10738 ;
  assign y2834 = n10761 ;
  assign y2835 = ~1'b0 ;
  assign y2836 = n10764 ;
  assign y2837 = ~n10770 ;
  assign y2838 = ~n10777 ;
  assign y2839 = n10778 ;
  assign y2840 = n10780 ;
  assign y2841 = ~1'b0 ;
  assign y2842 = ~1'b0 ;
  assign y2843 = ~1'b0 ;
  assign y2844 = n10786 ;
  assign y2845 = ~n10788 ;
  assign y2846 = ~n10789 ;
  assign y2847 = n10791 ;
  assign y2848 = ~n10794 ;
  assign y2849 = n10795 ;
  assign y2850 = n10797 ;
  assign y2851 = n10799 ;
  assign y2852 = ~n10801 ;
  assign y2853 = n10803 ;
  assign y2854 = ~n10813 ;
  assign y2855 = ~n10823 ;
  assign y2856 = n10833 ;
  assign y2857 = n10834 ;
  assign y2858 = ~n10836 ;
  assign y2859 = n10838 ;
  assign y2860 = n10841 ;
  assign y2861 = ~n10843 ;
  assign y2862 = n10850 ;
  assign y2863 = ~n10855 ;
  assign y2864 = ~n10867 ;
  assign y2865 = ~1'b0 ;
  assign y2866 = ~1'b0 ;
  assign y2867 = n10869 ;
  assign y2868 = ~n10875 ;
  assign y2869 = n10882 ;
  assign y2870 = n10885 ;
  assign y2871 = ~n10886 ;
  assign y2872 = n10888 ;
  assign y2873 = n10893 ;
  assign y2874 = ~n10900 ;
  assign y2875 = ~n10916 ;
  assign y2876 = n10918 ;
  assign y2877 = ~n10932 ;
  assign y2878 = n10936 ;
  assign y2879 = ~n10941 ;
  assign y2880 = ~1'b0 ;
  assign y2881 = ~n10944 ;
  assign y2882 = ~n10946 ;
  assign y2883 = ~n10962 ;
  assign y2884 = ~1'b0 ;
  assign y2885 = n10966 ;
  assign y2886 = ~n10969 ;
  assign y2887 = n10976 ;
  assign y2888 = ~n10977 ;
  assign y2889 = n10980 ;
  assign y2890 = ~1'b0 ;
  assign y2891 = ~n10982 ;
  assign y2892 = ~n10987 ;
  assign y2893 = n10996 ;
  assign y2894 = ~n10999 ;
  assign y2895 = ~n11002 ;
  assign y2896 = ~n11005 ;
  assign y2897 = n11006 ;
  assign y2898 = ~1'b0 ;
  assign y2899 = n11010 ;
  assign y2900 = ~n11011 ;
  assign y2901 = ~1'b0 ;
  assign y2902 = n11013 ;
  assign y2903 = ~n11015 ;
  assign y2904 = ~n11019 ;
  assign y2905 = ~n11020 ;
  assign y2906 = n11024 ;
  assign y2907 = n11036 ;
  assign y2908 = ~1'b0 ;
  assign y2909 = ~n11041 ;
  assign y2910 = n11043 ;
  assign y2911 = n11057 ;
  assign y2912 = ~n11058 ;
  assign y2913 = n11066 ;
  assign y2914 = ~n11069 ;
  assign y2915 = n11071 ;
  assign y2916 = ~1'b0 ;
  assign y2917 = ~n11077 ;
  assign y2918 = ~n11079 ;
  assign y2919 = ~n11080 ;
  assign y2920 = n6954 ;
  assign y2921 = n11081 ;
  assign y2922 = ~n11087 ;
  assign y2923 = ~n11092 ;
  assign y2924 = ~1'b0 ;
  assign y2925 = ~n11095 ;
  assign y2926 = n11102 ;
  assign y2927 = ~n11106 ;
  assign y2928 = n11107 ;
  assign y2929 = n11108 ;
  assign y2930 = n11109 ;
  assign y2931 = n11110 ;
  assign y2932 = ~n11114 ;
  assign y2933 = n11115 ;
  assign y2934 = n11120 ;
  assign y2935 = ~n11124 ;
  assign y2936 = ~n11127 ;
  assign y2937 = ~1'b0 ;
  assign y2938 = ~n11129 ;
  assign y2939 = n11131 ;
  assign y2940 = ~n11134 ;
  assign y2941 = n11136 ;
  assign y2942 = ~n11138 ;
  assign y2943 = n11139 ;
  assign y2944 = n11142 ;
  assign y2945 = n11146 ;
  assign y2946 = n11148 ;
  assign y2947 = n11150 ;
  assign y2948 = ~n11152 ;
  assign y2949 = ~n11154 ;
  assign y2950 = ~n11162 ;
  assign y2951 = ~n11168 ;
  assign y2952 = ~n11170 ;
  assign y2953 = n11173 ;
  assign y2954 = n11175 ;
  assign y2955 = ~1'b0 ;
  assign y2956 = n11176 ;
  assign y2957 = ~n11180 ;
  assign y2958 = n11181 ;
  assign y2959 = n11187 ;
  assign y2960 = n11191 ;
  assign y2961 = n11194 ;
  assign y2962 = ~n11196 ;
  assign y2963 = n11197 ;
  assign y2964 = ~n11199 ;
  assign y2965 = ~n11206 ;
  assign y2966 = n11208 ;
  assign y2967 = n11209 ;
  assign y2968 = ~n11216 ;
  assign y2969 = n11219 ;
  assign y2970 = n11229 ;
  assign y2971 = n11232 ;
  assign y2972 = ~n11236 ;
  assign y2973 = ~n11248 ;
  assign y2974 = ~n11253 ;
  assign y2975 = n11255 ;
  assign y2976 = ~n11261 ;
  assign y2977 = n11262 ;
  assign y2978 = ~n11267 ;
  assign y2979 = n11271 ;
  assign y2980 = ~n11274 ;
  assign y2981 = ~n11280 ;
  assign y2982 = ~1'b0 ;
  assign y2983 = ~n11283 ;
  assign y2984 = n11292 ;
  assign y2985 = n11293 ;
  assign y2986 = n11297 ;
  assign y2987 = ~n11299 ;
  assign y2988 = ~n11302 ;
  assign y2989 = n11306 ;
  assign y2990 = ~n11307 ;
  assign y2991 = n11308 ;
  assign y2992 = ~1'b0 ;
  assign y2993 = n11313 ;
  assign y2994 = ~n11318 ;
  assign y2995 = ~n11328 ;
  assign y2996 = ~1'b0 ;
  assign y2997 = ~n11333 ;
  assign y2998 = ~n11336 ;
  assign y2999 = n11339 ;
  assign y3000 = n11342 ;
  assign y3001 = ~n11347 ;
  assign y3002 = ~1'b0 ;
  assign y3003 = n11349 ;
  assign y3004 = ~n11353 ;
  assign y3005 = n11356 ;
  assign y3006 = ~n11361 ;
  assign y3007 = ~n11364 ;
  assign y3008 = n11367 ;
  assign y3009 = n11368 ;
  assign y3010 = n11376 ;
  assign y3011 = ~n11377 ;
  assign y3012 = ~1'b0 ;
  assign y3013 = ~n11385 ;
  assign y3014 = n11392 ;
  assign y3015 = ~n11397 ;
  assign y3016 = ~1'b0 ;
  assign y3017 = ~n11399 ;
  assign y3018 = n11410 ;
  assign y3019 = ~n11413 ;
  assign y3020 = ~n11416 ;
  assign y3021 = ~1'b0 ;
  assign y3022 = ~1'b0 ;
  assign y3023 = ~n11424 ;
  assign y3024 = n11425 ;
  assign y3025 = n11427 ;
  assign y3026 = n11434 ;
  assign y3027 = n11438 ;
  assign y3028 = n3565 ;
  assign y3029 = n11439 ;
  assign y3030 = n11444 ;
  assign y3031 = ~1'b0 ;
  assign y3032 = n11446 ;
  assign y3033 = ~1'b0 ;
  assign y3034 = ~n11455 ;
  assign y3035 = ~n11457 ;
  assign y3036 = ~n11458 ;
  assign y3037 = ~n11463 ;
  assign y3038 = n11466 ;
  assign y3039 = n11473 ;
  assign y3040 = n11474 ;
  assign y3041 = ~n11477 ;
  assign y3042 = n11483 ;
  assign y3043 = ~n11485 ;
  assign y3044 = ~n11486 ;
  assign y3045 = ~n11489 ;
  assign y3046 = ~n11493 ;
  assign y3047 = ~1'b0 ;
  assign y3048 = n11498 ;
  assign y3049 = ~n11503 ;
  assign y3050 = n11505 ;
  assign y3051 = n11513 ;
  assign y3052 = n11514 ;
  assign y3053 = ~n11533 ;
  assign y3054 = ~1'b0 ;
  assign y3055 = n11537 ;
  assign y3056 = ~n11550 ;
  assign y3057 = ~n11556 ;
  assign y3058 = ~1'b0 ;
  assign y3059 = ~n11558 ;
  assign y3060 = n11568 ;
  assign y3061 = ~n11572 ;
  assign y3062 = ~n11583 ;
  assign y3063 = ~n11590 ;
  assign y3064 = n11593 ;
  assign y3065 = n11605 ;
  assign y3066 = n11615 ;
  assign y3067 = ~n11619 ;
  assign y3068 = ~1'b0 ;
  assign y3069 = ~n11624 ;
  assign y3070 = n11627 ;
  assign y3071 = ~n11635 ;
  assign y3072 = ~n11638 ;
  assign y3073 = n11642 ;
  assign y3074 = ~n11644 ;
  assign y3075 = n11645 ;
  assign y3076 = ~1'b0 ;
  assign y3077 = ~1'b0 ;
  assign y3078 = n11652 ;
  assign y3079 = n11655 ;
  assign y3080 = ~n11663 ;
  assign y3081 = n11664 ;
  assign y3082 = ~n11666 ;
  assign y3083 = ~n11669 ;
  assign y3084 = ~1'b0 ;
  assign y3085 = ~n11672 ;
  assign y3086 = ~n11674 ;
  assign y3087 = n11698 ;
  assign y3088 = ~1'b0 ;
  assign y3089 = ~1'b0 ;
  assign y3090 = n11700 ;
  assign y3091 = ~n11701 ;
  assign y3092 = ~n11702 ;
  assign y3093 = ~n11705 ;
  assign y3094 = ~1'b0 ;
  assign y3095 = n11706 ;
  assign y3096 = n11710 ;
  assign y3097 = ~1'b0 ;
  assign y3098 = n11715 ;
  assign y3099 = ~1'b0 ;
  assign y3100 = ~1'b0 ;
  assign y3101 = n11721 ;
  assign y3102 = ~n11723 ;
  assign y3103 = ~1'b0 ;
  assign y3104 = ~n11726 ;
  assign y3105 = ~1'b0 ;
  assign y3106 = n11729 ;
  assign y3107 = ~n11730 ;
  assign y3108 = n11734 ;
  assign y3109 = ~1'b0 ;
  assign y3110 = ~n11744 ;
  assign y3111 = ~1'b0 ;
  assign y3112 = ~1'b0 ;
  assign y3113 = ~1'b0 ;
  assign y3114 = ~1'b0 ;
  assign y3115 = n11745 ;
  assign y3116 = ~n11752 ;
  assign y3117 = ~n11755 ;
  assign y3118 = ~1'b0 ;
  assign y3119 = ~n11759 ;
  assign y3120 = n11761 ;
  assign y3121 = ~n11762 ;
  assign y3122 = n11768 ;
  assign y3123 = ~1'b0 ;
  assign y3124 = n11770 ;
  assign y3125 = ~n11771 ;
  assign y3126 = n11774 ;
  assign y3127 = ~n4157 ;
  assign y3128 = n11775 ;
  assign y3129 = ~1'b0 ;
  assign y3130 = ~1'b0 ;
  assign y3131 = ~n11779 ;
  assign y3132 = n11786 ;
  assign y3133 = ~n11788 ;
  assign y3134 = n11790 ;
  assign y3135 = ~n11794 ;
  assign y3136 = ~1'b0 ;
  assign y3137 = ~n11797 ;
  assign y3138 = ~n11808 ;
  assign y3139 = ~n11810 ;
  assign y3140 = ~1'b0 ;
  assign y3141 = n11813 ;
  assign y3142 = ~n11817 ;
  assign y3143 = n11823 ;
  assign y3144 = n11824 ;
  assign y3145 = n11826 ;
  assign y3146 = n11833 ;
  assign y3147 = n11836 ;
  assign y3148 = ~1'b0 ;
  assign y3149 = n11841 ;
  assign y3150 = ~n11843 ;
  assign y3151 = n11844 ;
  assign y3152 = ~n11853 ;
  assign y3153 = ~n11854 ;
  assign y3154 = n11862 ;
  assign y3155 = ~n11871 ;
  assign y3156 = n11875 ;
  assign y3157 = n11879 ;
  assign y3158 = n11880 ;
  assign y3159 = n11882 ;
  assign y3160 = ~1'b0 ;
  assign y3161 = ~1'b0 ;
  assign y3162 = n11885 ;
  assign y3163 = ~n11893 ;
  assign y3164 = n11896 ;
  assign y3165 = ~1'b0 ;
  assign y3166 = ~n11903 ;
  assign y3167 = ~n11905 ;
  assign y3168 = n11911 ;
  assign y3169 = n11913 ;
  assign y3170 = ~n11919 ;
  assign y3171 = ~n11921 ;
  assign y3172 = n11926 ;
  assign y3173 = n11933 ;
  assign y3174 = ~n11938 ;
  assign y3175 = n11939 ;
  assign y3176 = ~n3695 ;
  assign y3177 = ~n11943 ;
  assign y3178 = ~1'b0 ;
  assign y3179 = n11951 ;
  assign y3180 = n11953 ;
  assign y3181 = ~n11954 ;
  assign y3182 = n11958 ;
  assign y3183 = ~n11960 ;
  assign y3184 = ~n11962 ;
  assign y3185 = ~1'b0 ;
  assign y3186 = n11964 ;
  assign y3187 = ~n11966 ;
  assign y3188 = ~n11968 ;
  assign y3189 = ~n11969 ;
  assign y3190 = ~1'b0 ;
  assign y3191 = n11970 ;
  assign y3192 = ~1'b0 ;
  assign y3193 = ~n11976 ;
  assign y3194 = ~n8510 ;
  assign y3195 = ~n11977 ;
  assign y3196 = ~n11979 ;
  assign y3197 = n11982 ;
  assign y3198 = n11985 ;
  assign y3199 = ~n11990 ;
  assign y3200 = ~1'b0 ;
  assign y3201 = ~n11993 ;
  assign y3202 = ~n11998 ;
  assign y3203 = ~n12002 ;
  assign y3204 = n12004 ;
  assign y3205 = ~1'b0 ;
  assign y3206 = n12012 ;
  assign y3207 = n12014 ;
  assign y3208 = n12017 ;
  assign y3209 = n12019 ;
  assign y3210 = n12023 ;
  assign y3211 = ~n12025 ;
  assign y3212 = n12034 ;
  assign y3213 = ~1'b0 ;
  assign y3214 = n12037 ;
  assign y3215 = ~1'b0 ;
  assign y3216 = n12039 ;
  assign y3217 = n12046 ;
  assign y3218 = ~n12048 ;
  assign y3219 = ~n12052 ;
  assign y3220 = ~1'b0 ;
  assign y3221 = n12055 ;
  assign y3222 = ~n12057 ;
  assign y3223 = ~n12059 ;
  assign y3224 = n12060 ;
  assign y3225 = ~n12062 ;
  assign y3226 = ~1'b0 ;
  assign y3227 = ~1'b0 ;
  assign y3228 = n12064 ;
  assign y3229 = n12069 ;
  assign y3230 = ~n12079 ;
  assign y3231 = n12080 ;
  assign y3232 = ~n12081 ;
  assign y3233 = ~1'b0 ;
  assign y3234 = ~n12085 ;
  assign y3235 = ~1'b0 ;
  assign y3236 = ~1'b0 ;
  assign y3237 = ~1'b0 ;
  assign y3238 = ~1'b0 ;
  assign y3239 = ~n12097 ;
  assign y3240 = ~n12099 ;
  assign y3241 = n12100 ;
  assign y3242 = n12101 ;
  assign y3243 = ~n12106 ;
  assign y3244 = ~n12107 ;
  assign y3245 = ~n12110 ;
  assign y3246 = ~n12117 ;
  assign y3247 = n12119 ;
  assign y3248 = n12125 ;
  assign y3249 = n12131 ;
  assign y3250 = ~n12132 ;
  assign y3251 = ~n12141 ;
  assign y3252 = ~n12147 ;
  assign y3253 = n12151 ;
  assign y3254 = n12156 ;
  assign y3255 = ~1'b0 ;
  assign y3256 = n12163 ;
  assign y3257 = n12165 ;
  assign y3258 = n12167 ;
  assign y3259 = ~n12172 ;
  assign y3260 = n12176 ;
  assign y3261 = ~n12188 ;
  assign y3262 = ~n12190 ;
  assign y3263 = n12192 ;
  assign y3264 = ~n12194 ;
  assign y3265 = ~1'b0 ;
  assign y3266 = ~1'b0 ;
  assign y3267 = n12200 ;
  assign y3268 = n12205 ;
  assign y3269 = ~1'b0 ;
  assign y3270 = ~1'b0 ;
  assign y3271 = ~n12208 ;
  assign y3272 = ~1'b0 ;
  assign y3273 = n12210 ;
  assign y3274 = ~n12223 ;
  assign y3275 = ~n2361 ;
  assign y3276 = n12226 ;
  assign y3277 = ~n12228 ;
  assign y3278 = n12234 ;
  assign y3279 = ~n12237 ;
  assign y3280 = n12243 ;
  assign y3281 = n12248 ;
  assign y3282 = ~n12249 ;
  assign y3283 = n12253 ;
  assign y3284 = ~n12254 ;
  assign y3285 = ~1'b0 ;
  assign y3286 = ~n12267 ;
  assign y3287 = ~n12272 ;
  assign y3288 = ~n12276 ;
  assign y3289 = n12281 ;
  assign y3290 = n12282 ;
  assign y3291 = ~n12284 ;
  assign y3292 = n12288 ;
  assign y3293 = n12289 ;
  assign y3294 = n12290 ;
  assign y3295 = n12292 ;
  assign y3296 = ~n12294 ;
  assign y3297 = ~n12300 ;
  assign y3298 = ~n12301 ;
  assign y3299 = ~n12302 ;
  assign y3300 = ~n12304 ;
  assign y3301 = ~n12310 ;
  assign y3302 = ~1'b0 ;
  assign y3303 = n12313 ;
  assign y3304 = ~n11839 ;
  assign y3305 = ~n12317 ;
  assign y3306 = ~n12324 ;
  assign y3307 = ~n12333 ;
  assign y3308 = ~1'b0 ;
  assign y3309 = ~1'b0 ;
  assign y3310 = ~1'b0 ;
  assign y3311 = n12334 ;
  assign y3312 = ~n12335 ;
  assign y3313 = n12336 ;
  assign y3314 = n12337 ;
  assign y3315 = n12342 ;
  assign y3316 = ~n12343 ;
  assign y3317 = ~n12347 ;
  assign y3318 = ~n12355 ;
  assign y3319 = ~n12360 ;
  assign y3320 = n12362 ;
  assign y3321 = ~1'b0 ;
  assign y3322 = n12363 ;
  assign y3323 = n12365 ;
  assign y3324 = ~n12369 ;
  assign y3325 = ~n12370 ;
  assign y3326 = ~n12371 ;
  assign y3327 = n12376 ;
  assign y3328 = n12380 ;
  assign y3329 = ~n12381 ;
  assign y3330 = n12385 ;
  assign y3331 = n12390 ;
  assign y3332 = ~n12391 ;
  assign y3333 = ~n12393 ;
  assign y3334 = ~1'b0 ;
  assign y3335 = ~1'b0 ;
  assign y3336 = n12399 ;
  assign y3337 = n12404 ;
  assign y3338 = ~n12405 ;
  assign y3339 = n12406 ;
  assign y3340 = ~n12413 ;
  assign y3341 = ~1'b0 ;
  assign y3342 = ~n12417 ;
  assign y3343 = ~n12419 ;
  assign y3344 = ~n12423 ;
  assign y3345 = ~1'b0 ;
  assign y3346 = n12427 ;
  assign y3347 = n12429 ;
  assign y3348 = n12431 ;
  assign y3349 = ~1'b0 ;
  assign y3350 = n12432 ;
  assign y3351 = n12434 ;
  assign y3352 = n12438 ;
  assign y3353 = ~n12440 ;
  assign y3354 = ~1'b0 ;
  assign y3355 = ~1'b0 ;
  assign y3356 = ~1'b0 ;
  assign y3357 = ~n12442 ;
  assign y3358 = n12444 ;
  assign y3359 = ~n12455 ;
  assign y3360 = n12456 ;
  assign y3361 = ~1'b0 ;
  assign y3362 = n12458 ;
  assign y3363 = ~n12460 ;
  assign y3364 = ~n12469 ;
  assign y3365 = n12470 ;
  assign y3366 = ~1'b0 ;
  assign y3367 = ~n12479 ;
  assign y3368 = ~n12481 ;
  assign y3369 = n12489 ;
  assign y3370 = ~n12492 ;
  assign y3371 = ~n12496 ;
  assign y3372 = n12500 ;
  assign y3373 = n12506 ;
  assign y3374 = ~1'b0 ;
  assign y3375 = n12508 ;
  assign y3376 = ~n12511 ;
  assign y3377 = n12514 ;
  assign y3378 = ~n12515 ;
  assign y3379 = ~1'b0 ;
  assign y3380 = ~n12519 ;
  assign y3381 = ~n12522 ;
  assign y3382 = n12523 ;
  assign y3383 = n12524 ;
  assign y3384 = n12531 ;
  assign y3385 = n12535 ;
  assign y3386 = n12542 ;
  assign y3387 = 1'b0 ;
  assign y3388 = n12545 ;
  assign y3389 = n1617 ;
  assign y3390 = ~n12548 ;
  assign y3391 = n12551 ;
  assign y3392 = ~1'b0 ;
  assign y3393 = n12559 ;
  assign y3394 = ~n12562 ;
  assign y3395 = n12566 ;
  assign y3396 = ~n12567 ;
  assign y3397 = n12569 ;
  assign y3398 = n12575 ;
  assign y3399 = ~n12581 ;
  assign y3400 = ~1'b0 ;
  assign y3401 = ~n12582 ;
  assign y3402 = ~n12583 ;
  assign y3403 = n12588 ;
  assign y3404 = ~n12596 ;
  assign y3405 = n12597 ;
  assign y3406 = 1'b0 ;
  assign y3407 = n12600 ;
  assign y3408 = ~n12603 ;
  assign y3409 = n12606 ;
  assign y3410 = ~1'b0 ;
  assign y3411 = ~n12614 ;
  assign y3412 = n12620 ;
  assign y3413 = ~n12621 ;
  assign y3414 = ~n12622 ;
  assign y3415 = ~n12625 ;
  assign y3416 = ~n12631 ;
  assign y3417 = n12639 ;
  assign y3418 = n12641 ;
  assign y3419 = ~n12642 ;
  assign y3420 = n12647 ;
  assign y3421 = n12650 ;
  assign y3422 = n12655 ;
  assign y3423 = ~n12662 ;
  assign y3424 = ~n12665 ;
  assign y3425 = ~n12682 ;
  assign y3426 = n12683 ;
  assign y3427 = ~n12688 ;
  assign y3428 = n12691 ;
  assign y3429 = n12694 ;
  assign y3430 = ~n12695 ;
  assign y3431 = n12698 ;
  assign y3432 = n12702 ;
  assign y3433 = n12708 ;
  assign y3434 = ~n12716 ;
  assign y3435 = ~n12717 ;
  assign y3436 = n12720 ;
  assign y3437 = n725 ;
  assign y3438 = n12721 ;
  assign y3439 = ~n12727 ;
  assign y3440 = n12734 ;
  assign y3441 = ~n12735 ;
  assign y3442 = n12737 ;
  assign y3443 = n12741 ;
  assign y3444 = n12742 ;
  assign y3445 = n12744 ;
  assign y3446 = n12749 ;
  assign y3447 = ~n12752 ;
  assign y3448 = n12754 ;
  assign y3449 = n12756 ;
  assign y3450 = n12759 ;
  assign y3451 = ~n12766 ;
  assign y3452 = n12767 ;
  assign y3453 = ~1'b0 ;
  assign y3454 = n12769 ;
  assign y3455 = ~n12770 ;
  assign y3456 = n11346 ;
  assign y3457 = n12777 ;
  assign y3458 = ~n12779 ;
  assign y3459 = n12780 ;
  assign y3460 = ~1'b0 ;
  assign y3461 = n12787 ;
  assign y3462 = n12790 ;
  assign y3463 = n12797 ;
  assign y3464 = ~n12799 ;
  assign y3465 = ~n12801 ;
  assign y3466 = n12806 ;
  assign y3467 = n2051 ;
  assign y3468 = ~n12807 ;
  assign y3469 = n12808 ;
  assign y3470 = ~n12810 ;
  assign y3471 = n12813 ;
  assign y3472 = ~n12815 ;
  assign y3473 = n12817 ;
  assign y3474 = n12821 ;
  assign y3475 = n12824 ;
  assign y3476 = ~n12825 ;
  assign y3477 = ~n12828 ;
  assign y3478 = ~n12830 ;
  assign y3479 = ~1'b0 ;
  assign y3480 = ~n12831 ;
  assign y3481 = n12832 ;
  assign y3482 = ~n12833 ;
  assign y3483 = ~n12834 ;
  assign y3484 = n12840 ;
  assign y3485 = ~1'b0 ;
  assign y3486 = ~1'b0 ;
  assign y3487 = ~n12841 ;
  assign y3488 = n12846 ;
  assign y3489 = ~1'b0 ;
  assign y3490 = ~1'b0 ;
  assign y3491 = ~n12851 ;
  assign y3492 = n12852 ;
  assign y3493 = ~n12855 ;
  assign y3494 = ~n12862 ;
  assign y3495 = ~n12863 ;
  assign y3496 = ~1'b0 ;
  assign y3497 = ~n12868 ;
  assign y3498 = ~n12876 ;
  assign y3499 = n12878 ;
  assign y3500 = ~n12881 ;
  assign y3501 = ~1'b0 ;
  assign y3502 = ~n12882 ;
  assign y3503 = n12885 ;
  assign y3504 = n12886 ;
  assign y3505 = ~1'b0 ;
  assign y3506 = n12900 ;
  assign y3507 = n12901 ;
  assign y3508 = n12906 ;
  assign y3509 = ~n12913 ;
  assign y3510 = n12918 ;
  assign y3511 = ~1'b0 ;
  assign y3512 = ~n12921 ;
  assign y3513 = ~n12922 ;
  assign y3514 = n12923 ;
  assign y3515 = n12930 ;
  assign y3516 = ~n12937 ;
  assign y3517 = ~n12945 ;
  assign y3518 = n12949 ;
  assign y3519 = n12950 ;
  assign y3520 = ~n12956 ;
  assign y3521 = n12957 ;
  assign y3522 = ~n12959 ;
  assign y3523 = n12968 ;
  assign y3524 = ~n12983 ;
  assign y3525 = ~n12991 ;
  assign y3526 = ~n12993 ;
  assign y3527 = ~1'b0 ;
  assign y3528 = ~n12995 ;
  assign y3529 = n12997 ;
  assign y3530 = ~1'b0 ;
  assign y3531 = n13000 ;
  assign y3532 = ~1'b0 ;
  assign y3533 = n13007 ;
  assign y3534 = n13009 ;
  assign y3535 = ~n13011 ;
  assign y3536 = n13015 ;
  assign y3537 = ~n13023 ;
  assign y3538 = n13024 ;
  assign y3539 = ~n13025 ;
  assign y3540 = ~n13029 ;
  assign y3541 = ~1'b0 ;
  assign y3542 = n13030 ;
  assign y3543 = n13031 ;
  assign y3544 = ~n13032 ;
  assign y3545 = ~n13039 ;
  assign y3546 = n13042 ;
  assign y3547 = n13043 ;
  assign y3548 = ~n13045 ;
  assign y3549 = ~1'b0 ;
  assign y3550 = n13052 ;
  assign y3551 = n13054 ;
  assign y3552 = ~n13059 ;
  assign y3553 = ~n13060 ;
  assign y3554 = ~n13065 ;
  assign y3555 = n13076 ;
  assign y3556 = ~n13077 ;
  assign y3557 = n13089 ;
  assign y3558 = ~n13096 ;
  assign y3559 = n13098 ;
  assign y3560 = ~1'b0 ;
  assign y3561 = ~n13101 ;
  assign y3562 = n13103 ;
  assign y3563 = ~n13111 ;
  assign y3564 = n13114 ;
  assign y3565 = ~1'b0 ;
  assign y3566 = ~1'b0 ;
  assign y3567 = ~1'b0 ;
  assign y3568 = n13122 ;
  assign y3569 = n13123 ;
  assign y3570 = ~n13125 ;
  assign y3571 = ~n13131 ;
  assign y3572 = ~n13136 ;
  assign y3573 = ~n13145 ;
  assign y3574 = ~n13148 ;
  assign y3575 = ~n13151 ;
  assign y3576 = ~1'b0 ;
  assign y3577 = ~n13156 ;
  assign y3578 = n13159 ;
  assign y3579 = ~1'b0 ;
  assign y3580 = ~n13165 ;
  assign y3581 = n13166 ;
  assign y3582 = ~n13176 ;
  assign y3583 = ~1'b0 ;
  assign y3584 = n11483 ;
  assign y3585 = ~n13178 ;
  assign y3586 = ~1'b0 ;
  assign y3587 = n13180 ;
  assign y3588 = n13181 ;
  assign y3589 = ~n13184 ;
  assign y3590 = n13187 ;
  assign y3591 = n13190 ;
  assign y3592 = ~n13191 ;
  assign y3593 = n13195 ;
  assign y3594 = ~n13199 ;
  assign y3595 = ~1'b0 ;
  assign y3596 = ~n13200 ;
  assign y3597 = n13205 ;
  assign y3598 = n13228 ;
  assign y3599 = n13235 ;
  assign y3600 = n13236 ;
  assign y3601 = ~n13237 ;
  assign y3602 = 1'b0 ;
  assign y3603 = ~n13246 ;
  assign y3604 = n13248 ;
  assign y3605 = ~n13252 ;
  assign y3606 = n13254 ;
  assign y3607 = ~1'b0 ;
  assign y3608 = ~n13262 ;
  assign y3609 = ~1'b0 ;
  assign y3610 = ~n13271 ;
  assign y3611 = ~n13278 ;
  assign y3612 = ~n13280 ;
  assign y3613 = ~n13284 ;
  assign y3614 = ~n13287 ;
  assign y3615 = n13292 ;
  assign y3616 = ~n13302 ;
  assign y3617 = ~n13320 ;
  assign y3618 = ~n13322 ;
  assign y3619 = ~n13324 ;
  assign y3620 = ~n13325 ;
  assign y3621 = n4604 ;
  assign y3622 = n13328 ;
  assign y3623 = ~n13331 ;
  assign y3624 = ~1'b0 ;
  assign y3625 = ~1'b0 ;
  assign y3626 = n13332 ;
  assign y3627 = ~1'b0 ;
  assign y3628 = ~n13338 ;
  assign y3629 = n13342 ;
  assign y3630 = n13348 ;
  assign y3631 = ~n13354 ;
  assign y3632 = n13356 ;
  assign y3633 = ~n13358 ;
  assign y3634 = n13363 ;
  assign y3635 = ~1'b0 ;
  assign y3636 = ~n13365 ;
  assign y3637 = n13368 ;
  assign y3638 = n13372 ;
  assign y3639 = ~n13381 ;
  assign y3640 = ~n13385 ;
  assign y3641 = n13388 ;
  assign y3642 = ~n13390 ;
  assign y3643 = n13393 ;
  assign y3644 = ~n13401 ;
  assign y3645 = n13410 ;
  assign y3646 = n13415 ;
  assign y3647 = n13418 ;
  assign y3648 = ~n13426 ;
  assign y3649 = ~n13431 ;
  assign y3650 = n13433 ;
  assign y3651 = ~1'b0 ;
  assign y3652 = n13434 ;
  assign y3653 = n13437 ;
  assign y3654 = n13440 ;
  assign y3655 = ~n13443 ;
  assign y3656 = ~n13445 ;
  assign y3657 = ~n13450 ;
  assign y3658 = ~n13455 ;
  assign y3659 = ~n13466 ;
  assign y3660 = ~1'b0 ;
  assign y3661 = ~1'b0 ;
  assign y3662 = n13467 ;
  assign y3663 = ~n13470 ;
  assign y3664 = n13471 ;
  assign y3665 = ~n13475 ;
  assign y3666 = n13480 ;
  assign y3667 = n13488 ;
  assign y3668 = ~n13489 ;
  assign y3669 = ~n13490 ;
  assign y3670 = n13491 ;
  assign y3671 = ~n13492 ;
  assign y3672 = n13495 ;
  assign y3673 = n13496 ;
  assign y3674 = ~1'b0 ;
  assign y3675 = ~n13502 ;
  assign y3676 = n13506 ;
  assign y3677 = n13507 ;
  assign y3678 = ~n13515 ;
  assign y3679 = n13521 ;
  assign y3680 = n13525 ;
  assign y3681 = ~1'b0 ;
  assign y3682 = n13527 ;
  assign y3683 = ~n13528 ;
  assign y3684 = ~n9189 ;
  assign y3685 = ~n13531 ;
  assign y3686 = n13533 ;
  assign y3687 = n13539 ;
  assign y3688 = ~1'b0 ;
  assign y3689 = ~1'b0 ;
  assign y3690 = n13540 ;
  assign y3691 = ~n13545 ;
  assign y3692 = n13546 ;
  assign y3693 = n4056 ;
  assign y3694 = ~1'b0 ;
  assign y3695 = ~n13548 ;
  assign y3696 = ~n13550 ;
  assign y3697 = n13553 ;
  assign y3698 = ~1'b0 ;
  assign y3699 = n13555 ;
  assign y3700 = ~n13556 ;
  assign y3701 = n13559 ;
  assign y3702 = ~n13562 ;
  assign y3703 = n13565 ;
  assign y3704 = ~n13566 ;
  assign y3705 = ~n13576 ;
  assign y3706 = n13579 ;
  assign y3707 = n13580 ;
  assign y3708 = n13582 ;
  assign y3709 = n13586 ;
  assign y3710 = ~n13588 ;
  assign y3711 = ~n9208 ;
  assign y3712 = n13590 ;
  assign y3713 = n13592 ;
  assign y3714 = n13601 ;
  assign y3715 = n13602 ;
  assign y3716 = ~n13605 ;
  assign y3717 = ~1'b0 ;
  assign y3718 = n13606 ;
  assign y3719 = n13607 ;
  assign y3720 = ~n13610 ;
  assign y3721 = n13612 ;
  assign y3722 = n13614 ;
  assign y3723 = ~n13616 ;
  assign y3724 = n13619 ;
  assign y3725 = n13623 ;
  assign y3726 = n13625 ;
  assign y3727 = ~1'b0 ;
  assign y3728 = n13631 ;
  assign y3729 = n13639 ;
  assign y3730 = ~n13647 ;
  assign y3731 = ~1'b0 ;
  assign y3732 = ~n13651 ;
  assign y3733 = ~n13654 ;
  assign y3734 = ~n13656 ;
  assign y3735 = n13660 ;
  assign y3736 = ~n13665 ;
  assign y3737 = n13671 ;
  assign y3738 = ~n13673 ;
  assign y3739 = ~n13674 ;
  assign y3740 = ~1'b0 ;
  assign y3741 = n13677 ;
  assign y3742 = ~n6187 ;
  assign y3743 = n13681 ;
  assign y3744 = ~n13683 ;
  assign y3745 = ~n13684 ;
  assign y3746 = ~1'b0 ;
  assign y3747 = ~n13689 ;
  assign y3748 = n13698 ;
  assign y3749 = ~n13699 ;
  assign y3750 = n13703 ;
  assign y3751 = ~n13715 ;
  assign y3752 = ~n13719 ;
  assign y3753 = n13720 ;
  assign y3754 = ~n13724 ;
  assign y3755 = ~n13726 ;
  assign y3756 = ~n13728 ;
  assign y3757 = n13729 ;
  assign y3758 = n13730 ;
  assign y3759 = ~n13734 ;
  assign y3760 = n13742 ;
  assign y3761 = ~n13745 ;
  assign y3762 = n13746 ;
  assign y3763 = ~1'b0 ;
  assign y3764 = n13749 ;
  assign y3765 = ~n13756 ;
  assign y3766 = ~n13757 ;
  assign y3767 = ~n13759 ;
  assign y3768 = ~1'b0 ;
  assign y3769 = ~n13762 ;
  assign y3770 = ~n13766 ;
  assign y3771 = n13768 ;
  assign y3772 = n13771 ;
  assign y3773 = ~n13773 ;
  assign y3774 = n13774 ;
  assign y3775 = ~1'b0 ;
  assign y3776 = n13777 ;
  assign y3777 = n13783 ;
  assign y3778 = ~n13784 ;
  assign y3779 = n13786 ;
  assign y3780 = n13790 ;
  assign y3781 = ~n13793 ;
  assign y3782 = ~n13794 ;
  assign y3783 = ~n13795 ;
  assign y3784 = n13796 ;
  assign y3785 = ~n13806 ;
  assign y3786 = n13810 ;
  assign y3787 = ~n3053 ;
  assign y3788 = n13818 ;
  assign y3789 = ~1'b0 ;
  assign y3790 = n1690 ;
  assign y3791 = n13819 ;
  assign y3792 = ~n13821 ;
  assign y3793 = ~n13823 ;
  assign y3794 = ~n13825 ;
  assign y3795 = ~n13831 ;
  assign y3796 = n13836 ;
  assign y3797 = ~1'b0 ;
  assign y3798 = ~n13843 ;
  assign y3799 = n13847 ;
  assign y3800 = n13849 ;
  assign y3801 = ~1'b0 ;
  assign y3802 = ~n13852 ;
  assign y3803 = n13855 ;
  assign y3804 = ~n13857 ;
  assign y3805 = ~n13858 ;
  assign y3806 = n13864 ;
  assign y3807 = ~n13865 ;
  assign y3808 = ~n13869 ;
  assign y3809 = ~1'b0 ;
  assign y3810 = ~n13872 ;
  assign y3811 = ~n13876 ;
  assign y3812 = ~n13880 ;
  assign y3813 = 1'b0 ;
  assign y3814 = ~n13884 ;
  assign y3815 = ~1'b0 ;
  assign y3816 = ~n13887 ;
  assign y3817 = ~n13889 ;
  assign y3818 = ~1'b0 ;
  assign y3819 = n13891 ;
  assign y3820 = ~n13892 ;
  assign y3821 = ~n13899 ;
  assign y3822 = n13903 ;
  assign y3823 = ~n13905 ;
  assign y3824 = ~n13907 ;
  assign y3825 = ~1'b0 ;
  assign y3826 = ~1'b0 ;
  assign y3827 = n13909 ;
  assign y3828 = n13913 ;
  assign y3829 = ~n3126 ;
  assign y3830 = ~1'b0 ;
  assign y3831 = n13918 ;
  assign y3832 = n13923 ;
  assign y3833 = ~1'b0 ;
  assign y3834 = ~1'b0 ;
  assign y3835 = ~n13924 ;
  assign y3836 = n13929 ;
  assign y3837 = ~1'b0 ;
  assign y3838 = n13930 ;
  assign y3839 = ~n13935 ;
  assign y3840 = ~n13936 ;
  assign y3841 = ~n13941 ;
  assign y3842 = n13943 ;
  assign y3843 = n13945 ;
  assign y3844 = ~n13949 ;
  assign y3845 = n13951 ;
  assign y3846 = ~n13955 ;
  assign y3847 = ~n13957 ;
  assign y3848 = n13958 ;
  assign y3849 = ~n13971 ;
  assign y3850 = n13973 ;
  assign y3851 = ~n13977 ;
  assign y3852 = ~n13978 ;
  assign y3853 = ~n13982 ;
  assign y3854 = n11202 ;
  assign y3855 = ~n13991 ;
  assign y3856 = ~n13996 ;
  assign y3857 = ~n13998 ;
  assign y3858 = ~1'b0 ;
  assign y3859 = ~n13999 ;
  assign y3860 = ~1'b0 ;
  assign y3861 = ~n14000 ;
  assign y3862 = ~1'b0 ;
  assign y3863 = n9819 ;
  assign y3864 = n14001 ;
  assign y3865 = ~n14009 ;
  assign y3866 = ~n14012 ;
  assign y3867 = n14014 ;
  assign y3868 = ~n14019 ;
  assign y3869 = n14023 ;
  assign y3870 = ~n14027 ;
  assign y3871 = ~n14031 ;
  assign y3872 = ~n14037 ;
  assign y3873 = ~n14042 ;
  assign y3874 = ~n14047 ;
  assign y3875 = ~n14052 ;
  assign y3876 = ~n14054 ;
  assign y3877 = n14059 ;
  assign y3878 = ~n14063 ;
  assign y3879 = ~1'b0 ;
  assign y3880 = ~n14075 ;
  assign y3881 = ~n14076 ;
  assign y3882 = ~n14084 ;
  assign y3883 = n14085 ;
  assign y3884 = ~n14086 ;
  assign y3885 = ~n14100 ;
  assign y3886 = ~n14103 ;
  assign y3887 = n14105 ;
  assign y3888 = ~n14120 ;
  assign y3889 = ~n14122 ;
  assign y3890 = ~1'b0 ;
  assign y3891 = ~n12279 ;
  assign y3892 = ~n14125 ;
  assign y3893 = ~n14127 ;
  assign y3894 = ~n14128 ;
  assign y3895 = ~1'b0 ;
  assign y3896 = n7071 ;
  assign y3897 = ~n14133 ;
  assign y3898 = n2478 ;
  assign y3899 = n14137 ;
  assign y3900 = ~n14140 ;
  assign y3901 = n14141 ;
  assign y3902 = ~n14143 ;
  assign y3903 = n14144 ;
  assign y3904 = ~n14145 ;
  assign y3905 = ~n14150 ;
  assign y3906 = n14151 ;
  assign y3907 = ~1'b0 ;
  assign y3908 = ~1'b0 ;
  assign y3909 = ~n14155 ;
  assign y3910 = n14161 ;
  assign y3911 = n14163 ;
  assign y3912 = ~n14164 ;
  assign y3913 = n14165 ;
  assign y3914 = n14166 ;
  assign y3915 = ~1'b0 ;
  assign y3916 = ~n14167 ;
  assign y3917 = n14170 ;
  assign y3918 = ~n14174 ;
  assign y3919 = ~n14176 ;
  assign y3920 = ~1'b0 ;
  assign y3921 = n14177 ;
  assign y3922 = ~n14181 ;
  assign y3923 = ~n14184 ;
  assign y3924 = ~1'b0 ;
  assign y3925 = ~n14189 ;
  assign y3926 = n14196 ;
  assign y3927 = ~n14202 ;
  assign y3928 = ~1'b0 ;
  assign y3929 = ~n14203 ;
  assign y3930 = ~n14204 ;
  assign y3931 = ~n14212 ;
  assign y3932 = ~n14215 ;
  assign y3933 = ~n14217 ;
  assign y3934 = ~n14218 ;
  assign y3935 = ~n14219 ;
  assign y3936 = n14220 ;
  assign y3937 = ~1'b0 ;
  assign y3938 = ~n14229 ;
  assign y3939 = ~1'b0 ;
  assign y3940 = n14236 ;
  assign y3941 = n14237 ;
  assign y3942 = ~1'b0 ;
  assign y3943 = n14239 ;
  assign y3944 = ~n14242 ;
  assign y3945 = n14246 ;
  assign y3946 = ~n14253 ;
  assign y3947 = ~n14254 ;
  assign y3948 = ~n14257 ;
  assign y3949 = n14259 ;
  assign y3950 = n14260 ;
  assign y3951 = n14263 ;
  assign y3952 = ~1'b0 ;
  assign y3953 = ~n14269 ;
  assign y3954 = ~n14272 ;
  assign y3955 = ~1'b0 ;
  assign y3956 = ~n14274 ;
  assign y3957 = ~n14277 ;
  assign y3958 = ~n14280 ;
  assign y3959 = ~n14281 ;
  assign y3960 = ~n14286 ;
  assign y3961 = ~n14288 ;
  assign y3962 = n14296 ;
  assign y3963 = ~1'b0 ;
  assign y3964 = ~1'b0 ;
  assign y3965 = ~n14297 ;
  assign y3966 = n14310 ;
  assign y3967 = ~n14312 ;
  assign y3968 = ~n14315 ;
  assign y3969 = ~n14318 ;
  assign y3970 = n14319 ;
  assign y3971 = n14321 ;
  assign y3972 = n14331 ;
  assign y3973 = n14332 ;
  assign y3974 = ~n14336 ;
  assign y3975 = ~1'b0 ;
  assign y3976 = n14337 ;
  assign y3977 = ~n14340 ;
  assign y3978 = ~n14346 ;
  assign y3979 = n14359 ;
  assign y3980 = n14362 ;
  assign y3981 = ~1'b0 ;
  assign y3982 = ~n14367 ;
  assign y3983 = ~n14368 ;
  assign y3984 = ~n14369 ;
  assign y3985 = n14372 ;
  assign y3986 = ~n14379 ;
  assign y3987 = n14382 ;
  assign y3988 = n14384 ;
  assign y3989 = n14393 ;
  assign y3990 = ~n970 ;
  assign y3991 = ~1'b0 ;
  assign y3992 = n14394 ;
  assign y3993 = ~n14399 ;
  assign y3994 = n14401 ;
  assign y3995 = n14406 ;
  assign y3996 = ~n14409 ;
  assign y3997 = n14417 ;
  assign y3998 = n14422 ;
  assign y3999 = ~n14429 ;
  assign y4000 = ~n14430 ;
  assign y4001 = ~1'b0 ;
  assign y4002 = n14432 ;
  assign y4003 = ~n14434 ;
  assign y4004 = ~n14435 ;
  assign y4005 = ~n14438 ;
  assign y4006 = ~n14439 ;
  assign y4007 = ~n14443 ;
  assign y4008 = ~n14444 ;
  assign y4009 = n14448 ;
  assign y4010 = ~1'b0 ;
  assign y4011 = n14456 ;
  assign y4012 = ~n14458 ;
  assign y4013 = ~n14464 ;
  assign y4014 = ~n14467 ;
  assign y4015 = n14470 ;
  assign y4016 = n14474 ;
  assign y4017 = ~n14480 ;
  assign y4018 = ~n14487 ;
  assign y4019 = ~n14489 ;
  assign y4020 = ~n14494 ;
  assign y4021 = n14496 ;
  assign y4022 = ~n14497 ;
  assign y4023 = ~1'b0 ;
  assign y4024 = n14500 ;
  assign y4025 = n14506 ;
  assign y4026 = ~n14509 ;
  assign y4027 = n14516 ;
  assign y4028 = ~1'b0 ;
  assign y4029 = ~n14517 ;
  assign y4030 = n14518 ;
  assign y4031 = n14523 ;
  assign y4032 = ~n14524 ;
  assign y4033 = ~n14526 ;
  assign y4034 = n246 ;
  assign y4035 = ~n14527 ;
  assign y4036 = n14528 ;
  assign y4037 = n14532 ;
  assign y4038 = ~n14535 ;
  assign y4039 = ~1'b0 ;
  assign y4040 = ~n14538 ;
  assign y4041 = n14541 ;
  assign y4042 = n14547 ;
  assign y4043 = ~n14550 ;
  assign y4044 = n14553 ;
  assign y4045 = n14556 ;
  assign y4046 = ~n14566 ;
  assign y4047 = ~n14571 ;
  assign y4048 = ~n14572 ;
  assign y4049 = ~n14575 ;
  assign y4050 = ~n14576 ;
  assign y4051 = ~1'b0 ;
  assign y4052 = ~1'b0 ;
  assign y4053 = n14579 ;
  assign y4054 = n14585 ;
  assign y4055 = ~n14589 ;
  assign y4056 = n14595 ;
  assign y4057 = n14597 ;
  assign y4058 = ~n14599 ;
  assign y4059 = ~n14600 ;
  assign y4060 = n14603 ;
  assign y4061 = ~1'b0 ;
  assign y4062 = ~1'b0 ;
  assign y4063 = ~n14606 ;
  assign y4064 = n14608 ;
  assign y4065 = ~1'b0 ;
  assign y4066 = ~n14610 ;
  assign y4067 = n14611 ;
  assign y4068 = ~n14617 ;
  assign y4069 = n14619 ;
  assign y4070 = n14620 ;
  assign y4071 = ~n14623 ;
  assign y4072 = ~n14624 ;
  assign y4073 = ~n14625 ;
  assign y4074 = ~n14630 ;
  assign y4075 = n14637 ;
  assign y4076 = n14645 ;
  assign y4077 = ~1'b0 ;
  assign y4078 = ~n14646 ;
  assign y4079 = ~n14647 ;
  assign y4080 = n14653 ;
  assign y4081 = ~n14660 ;
  assign y4082 = n14661 ;
  assign y4083 = ~n14664 ;
  assign y4084 = ~n14666 ;
  assign y4085 = ~n14670 ;
  assign y4086 = n14675 ;
  assign y4087 = ~n14677 ;
  assign y4088 = n14681 ;
  assign y4089 = n14688 ;
  assign y4090 = n14691 ;
  assign y4091 = n14694 ;
  assign y4092 = ~n14695 ;
  assign y4093 = n14702 ;
  assign y4094 = ~n14704 ;
  assign y4095 = ~1'b0 ;
  assign y4096 = ~1'b0 ;
  assign y4097 = ~1'b0 ;
  assign y4098 = ~n14708 ;
  assign y4099 = ~n14709 ;
  assign y4100 = ~n14717 ;
  assign y4101 = ~n14719 ;
  assign y4102 = ~n14721 ;
  assign y4103 = ~n14726 ;
  assign y4104 = n14728 ;
  assign y4105 = n14730 ;
  assign y4106 = n14731 ;
  assign y4107 = n14732 ;
  assign y4108 = n14755 ;
  assign y4109 = n14756 ;
  assign y4110 = ~1'b0 ;
  assign y4111 = n14761 ;
  assign y4112 = ~n14765 ;
  assign y4113 = ~n14772 ;
  assign y4114 = n14774 ;
  assign y4115 = ~n14776 ;
  assign y4116 = n14780 ;
  assign y4117 = ~n14782 ;
  assign y4118 = ~1'b0 ;
  assign y4119 = n14784 ;
  assign y4120 = n14786 ;
  assign y4121 = ~1'b0 ;
  assign y4122 = ~n14791 ;
  assign y4123 = n14796 ;
  assign y4124 = n14804 ;
  assign y4125 = ~n14810 ;
  assign y4126 = n14813 ;
  assign y4127 = ~n4707 ;
  assign y4128 = n14636 ;
  assign y4129 = n14814 ;
  assign y4130 = n14815 ;
  assign y4131 = n14825 ;
  assign y4132 = ~n14828 ;
  assign y4133 = ~1'b0 ;
  assign y4134 = n14836 ;
  assign y4135 = n14843 ;
  assign y4136 = n14848 ;
  assign y4137 = ~n14849 ;
  assign y4138 = ~n14851 ;
  assign y4139 = n14853 ;
  assign y4140 = ~n14855 ;
  assign y4141 = ~1'b0 ;
  assign y4142 = ~n14857 ;
  assign y4143 = ~n14863 ;
  assign y4144 = ~1'b0 ;
  assign y4145 = ~1'b0 ;
  assign y4146 = ~n14872 ;
  assign y4147 = ~n14875 ;
  assign y4148 = ~n14887 ;
  assign y4149 = ~n14896 ;
  assign y4150 = ~n14902 ;
  assign y4151 = ~n14906 ;
  assign y4152 = n14908 ;
  assign y4153 = n14910 ;
  assign y4154 = ~n14912 ;
  assign y4155 = ~n14913 ;
  assign y4156 = n14922 ;
  assign y4157 = n14924 ;
  assign y4158 = ~1'b0 ;
  assign y4159 = n14936 ;
  assign y4160 = ~n14940 ;
  assign y4161 = ~1'b0 ;
  assign y4162 = ~n14945 ;
  assign y4163 = n14946 ;
  assign y4164 = n14036 ;
  assign y4165 = n14957 ;
  assign y4166 = ~n14961 ;
  assign y4167 = n14967 ;
  assign y4168 = ~n14969 ;
  assign y4169 = n14975 ;
  assign y4170 = ~n14977 ;
  assign y4171 = ~n14978 ;
  assign y4172 = n14980 ;
  assign y4173 = ~n14982 ;
  assign y4174 = n2352 ;
  assign y4175 = ~n14986 ;
  assign y4176 = n14989 ;
  assign y4177 = ~n14991 ;
  assign y4178 = n14997 ;
  assign y4179 = n14998 ;
  assign y4180 = ~1'b0 ;
  assign y4181 = ~n15000 ;
  assign y4182 = n15002 ;
  assign y4183 = n15003 ;
  assign y4184 = n15007 ;
  assign y4185 = ~n15009 ;
  assign y4186 = ~n15010 ;
  assign y4187 = ~n15021 ;
  assign y4188 = n15026 ;
  assign y4189 = ~1'b0 ;
  assign y4190 = ~1'b0 ;
  assign y4191 = ~n15033 ;
  assign y4192 = n15047 ;
  assign y4193 = n15048 ;
  assign y4194 = n15052 ;
  assign y4195 = n15057 ;
  assign y4196 = ~1'b0 ;
  assign y4197 = ~n15058 ;
  assign y4198 = n15059 ;
  assign y4199 = n15063 ;
  assign y4200 = n15078 ;
  assign y4201 = ~n15079 ;
  assign y4202 = ~n15084 ;
  assign y4203 = n15089 ;
  assign y4204 = ~n15090 ;
  assign y4205 = n15099 ;
  assign y4206 = ~1'b0 ;
  assign y4207 = ~n15101 ;
  assign y4208 = ~1'b0 ;
  assign y4209 = ~n15105 ;
  assign y4210 = n15109 ;
  assign y4211 = n15112 ;
  assign y4212 = ~n15114 ;
  assign y4213 = ~n15119 ;
  assign y4214 = 1'b0 ;
  assign y4215 = ~n15121 ;
  assign y4216 = n15124 ;
  assign y4217 = ~n15135 ;
  assign y4218 = ~1'b0 ;
  assign y4219 = ~n15138 ;
  assign y4220 = ~n15144 ;
  assign y4221 = ~n15151 ;
  assign y4222 = ~1'b0 ;
  assign y4223 = ~n15152 ;
  assign y4224 = n15155 ;
  assign y4225 = ~n15164 ;
  assign y4226 = ~n15167 ;
  assign y4227 = n15175 ;
  assign y4228 = ~n15176 ;
  assign y4229 = ~n15177 ;
  assign y4230 = ~1'b0 ;
  assign y4231 = n15179 ;
  assign y4232 = ~1'b0 ;
  assign y4233 = n15184 ;
  assign y4234 = ~n15189 ;
  assign y4235 = ~1'b0 ;
  assign y4236 = ~1'b0 ;
  assign y4237 = n15200 ;
  assign y4238 = ~n15202 ;
  assign y4239 = ~n15208 ;
  assign y4240 = n3610 ;
  assign y4241 = ~n15211 ;
  assign y4242 = n15213 ;
  assign y4243 = ~n15222 ;
  assign y4244 = n15224 ;
  assign y4245 = n15227 ;
  assign y4246 = n15229 ;
  assign y4247 = n15231 ;
  assign y4248 = n15235 ;
  assign y4249 = n15242 ;
  assign y4250 = ~n15250 ;
  assign y4251 = n15252 ;
  assign y4252 = ~1'b0 ;
  assign y4253 = ~n15262 ;
  assign y4254 = ~n15264 ;
  assign y4255 = n15265 ;
  assign y4256 = ~n15267 ;
  assign y4257 = ~1'b0 ;
  assign y4258 = ~n15269 ;
  assign y4259 = n15270 ;
  assign y4260 = ~n15271 ;
  assign y4261 = ~n15275 ;
  assign y4262 = n15280 ;
  assign y4263 = n15282 ;
  assign y4264 = ~1'b0 ;
  assign y4265 = n15286 ;
  assign y4266 = ~n15288 ;
  assign y4267 = n15289 ;
  assign y4268 = ~n15295 ;
  assign y4269 = n15312 ;
  assign y4270 = ~n15320 ;
  assign y4271 = ~n15322 ;
  assign y4272 = ~n15325 ;
  assign y4273 = ~n15327 ;
  assign y4274 = ~n15328 ;
  assign y4275 = ~1'b0 ;
  assign y4276 = ~n15335 ;
  assign y4277 = ~n15341 ;
  assign y4278 = ~1'b0 ;
  assign y4279 = ~n15349 ;
  assign y4280 = ~n15355 ;
  assign y4281 = n15356 ;
  assign y4282 = ~n15362 ;
  assign y4283 = ~1'b0 ;
  assign y4284 = ~1'b0 ;
  assign y4285 = ~n15364 ;
  assign y4286 = ~1'b0 ;
  assign y4287 = ~1'b0 ;
  assign y4288 = ~1'b0 ;
  assign y4289 = ~n15368 ;
  assign y4290 = ~n15373 ;
  assign y4291 = ~n15379 ;
  assign y4292 = ~n15387 ;
  assign y4293 = ~n15390 ;
  assign y4294 = n15401 ;
  assign y4295 = n15402 ;
  assign y4296 = ~n15405 ;
  assign y4297 = ~n15407 ;
  assign y4298 = n15412 ;
  assign y4299 = n15420 ;
  assign y4300 = n15421 ;
  assign y4301 = n15426 ;
  assign y4302 = n15427 ;
  assign y4303 = ~n15436 ;
  assign y4304 = ~1'b0 ;
  assign y4305 = n15445 ;
  assign y4306 = ~n15448 ;
  assign y4307 = n15458 ;
  assign y4308 = ~n15461 ;
  assign y4309 = n15464 ;
  assign y4310 = n15465 ;
  assign y4311 = n15466 ;
  assign y4312 = n15474 ;
  assign y4313 = ~n15475 ;
  assign y4314 = n15484 ;
  assign y4315 = n15488 ;
  assign y4316 = ~n15494 ;
  assign y4317 = ~n15500 ;
  assign y4318 = ~n15503 ;
  assign y4319 = n15509 ;
  assign y4320 = n15513 ;
  assign y4321 = n15516 ;
  assign y4322 = n15518 ;
  assign y4323 = ~1'b0 ;
  assign y4324 = ~n15526 ;
  assign y4325 = n15528 ;
  assign y4326 = n15533 ;
  assign y4327 = ~n11819 ;
  assign y4328 = n15541 ;
  assign y4329 = ~n15544 ;
  assign y4330 = ~1'b0 ;
  assign y4331 = n15547 ;
  assign y4332 = ~n15551 ;
  assign y4333 = ~1'b0 ;
  assign y4334 = ~n15553 ;
  assign y4335 = n15560 ;
  assign y4336 = ~1'b0 ;
  assign y4337 = ~n15561 ;
  assign y4338 = ~n15563 ;
  assign y4339 = ~n15564 ;
  assign y4340 = n15572 ;
  assign y4341 = ~n15577 ;
  assign y4342 = n15583 ;
  assign y4343 = ~1'b0 ;
  assign y4344 = ~1'b0 ;
  assign y4345 = ~n15584 ;
  assign y4346 = ~n15591 ;
  assign y4347 = n15592 ;
  assign y4348 = ~n15594 ;
  assign y4349 = ~n15595 ;
  assign y4350 = n15603 ;
  assign y4351 = ~n15606 ;
  assign y4352 = ~n15609 ;
  assign y4353 = ~n15611 ;
  assign y4354 = n15612 ;
  assign y4355 = n15615 ;
  assign y4356 = n15623 ;
  assign y4357 = ~n15625 ;
  assign y4358 = n15630 ;
  assign y4359 = n15634 ;
  assign y4360 = ~n15637 ;
  assign y4361 = n15638 ;
  assign y4362 = ~n15643 ;
  assign y4363 = n15645 ;
  assign y4364 = ~n15649 ;
  assign y4365 = n15650 ;
  assign y4366 = ~n15651 ;
  assign y4367 = ~n15654 ;
  assign y4368 = ~n15664 ;
  assign y4369 = n15666 ;
  assign y4370 = ~n15672 ;
  assign y4371 = n15680 ;
  assign y4372 = ~1'b0 ;
  assign y4373 = n15686 ;
  assign y4374 = n15687 ;
  assign y4375 = ~n15689 ;
  assign y4376 = ~1'b0 ;
  assign y4377 = ~n15692 ;
  assign y4378 = ~n15695 ;
  assign y4379 = ~n15696 ;
  assign y4380 = ~n15698 ;
  assign y4381 = ~n15699 ;
  assign y4382 = n15701 ;
  assign y4383 = n15704 ;
  assign y4384 = n15711 ;
  assign y4385 = ~n15715 ;
  assign y4386 = n15717 ;
  assign y4387 = ~n15720 ;
  assign y4388 = n15722 ;
  assign y4389 = ~n15723 ;
  assign y4390 = n15728 ;
  assign y4391 = ~n15729 ;
  assign y4392 = n15732 ;
  assign y4393 = ~n15737 ;
  assign y4394 = n15738 ;
  assign y4395 = n15745 ;
  assign y4396 = ~n15747 ;
  assign y4397 = n15748 ;
  assign y4398 = n15750 ;
  assign y4399 = n15753 ;
  assign y4400 = ~n15764 ;
  assign y4401 = ~n15767 ;
  assign y4402 = ~1'b0 ;
  assign y4403 = n15771 ;
  assign y4404 = ~n15773 ;
  assign y4405 = n15775 ;
  assign y4406 = ~1'b0 ;
  assign y4407 = ~n15777 ;
  assign y4408 = n15780 ;
  assign y4409 = ~n15781 ;
  assign y4410 = n15782 ;
  assign y4411 = n15784 ;
  assign y4412 = ~n13987 ;
  assign y4413 = ~1'b0 ;
  assign y4414 = n15785 ;
  assign y4415 = ~n15786 ;
  assign y4416 = ~1'b0 ;
  assign y4417 = n15794 ;
  assign y4418 = ~n15797 ;
  assign y4419 = n12861 ;
  assign y4420 = n15799 ;
  assign y4421 = ~n15802 ;
  assign y4422 = n15803 ;
  assign y4423 = ~1'b0 ;
  assign y4424 = n15806 ;
  assign y4425 = ~1'b0 ;
  assign y4426 = n15808 ;
  assign y4427 = n15811 ;
  assign y4428 = ~1'b0 ;
  assign y4429 = ~1'b0 ;
  assign y4430 = ~n15817 ;
  assign y4431 = n15822 ;
  assign y4432 = ~n15826 ;
  assign y4433 = ~n15829 ;
  assign y4434 = ~1'b0 ;
  assign y4435 = n15830 ;
  assign y4436 = n15831 ;
  assign y4437 = n15833 ;
  assign y4438 = ~n15834 ;
  assign y4439 = ~n15837 ;
  assign y4440 = n15842 ;
  assign y4441 = ~n15843 ;
  assign y4442 = ~1'b0 ;
  assign y4443 = ~n15846 ;
  assign y4444 = n15857 ;
  assign y4445 = ~n15859 ;
  assign y4446 = ~n15864 ;
  assign y4447 = n15870 ;
  assign y4448 = n15877 ;
  assign y4449 = ~n15879 ;
  assign y4450 = ~1'b0 ;
  assign y4451 = n15881 ;
  assign y4452 = n15882 ;
  assign y4453 = ~n15883 ;
  assign y4454 = ~1'b0 ;
  assign y4455 = ~1'b0 ;
  assign y4456 = ~n15885 ;
  assign y4457 = n15886 ;
  assign y4458 = n15890 ;
  assign y4459 = ~n15899 ;
  assign y4460 = ~n15904 ;
  assign y4461 = ~n15906 ;
  assign y4462 = n15915 ;
  assign y4463 = n15927 ;
  assign y4464 = ~n15931 ;
  assign y4465 = ~n15934 ;
  assign y4466 = n15935 ;
  assign y4467 = ~1'b0 ;
  assign y4468 = n15936 ;
  assign y4469 = n15939 ;
  assign y4470 = ~1'b0 ;
  assign y4471 = n15940 ;
  assign y4472 = ~n15941 ;
  assign y4473 = ~1'b0 ;
  assign y4474 = ~1'b0 ;
  assign y4475 = ~n12860 ;
  assign y4476 = n15956 ;
  assign y4477 = ~1'b0 ;
  assign y4478 = ~n15958 ;
  assign y4479 = n15960 ;
  assign y4480 = n15962 ;
  assign y4481 = n15965 ;
  assign y4482 = ~1'b0 ;
  assign y4483 = n15967 ;
  assign y4484 = n15968 ;
  assign y4485 = n15969 ;
  assign y4486 = ~n15973 ;
  assign y4487 = ~n10355 ;
  assign y4488 = ~n15974 ;
  assign y4489 = ~n13261 ;
  assign y4490 = ~n15976 ;
  assign y4491 = ~n15978 ;
  assign y4492 = ~n15987 ;
  assign y4493 = ~n15988 ;
  assign y4494 = ~n15990 ;
  assign y4495 = ~n15992 ;
  assign y4496 = n14043 ;
  assign y4497 = ~n15994 ;
  assign y4498 = ~n15997 ;
  assign y4499 = ~n15999 ;
  assign y4500 = n16000 ;
  assign y4501 = ~1'b0 ;
  assign y4502 = ~1'b0 ;
  assign y4503 = n16003 ;
  assign y4504 = ~n16004 ;
  assign y4505 = ~n16007 ;
  assign y4506 = n16016 ;
  assign y4507 = n16017 ;
  assign y4508 = n16020 ;
  assign y4509 = ~n16024 ;
  assign y4510 = n16033 ;
  assign y4511 = ~n16038 ;
  assign y4512 = n16043 ;
  assign y4513 = ~n16046 ;
  assign y4514 = ~n16050 ;
  assign y4515 = ~n16057 ;
  assign y4516 = ~n16058 ;
  assign y4517 = ~n16059 ;
  assign y4518 = n16061 ;
  assign y4519 = ~n16063 ;
  assign y4520 = n16070 ;
  assign y4521 = n16073 ;
  assign y4522 = n16074 ;
  assign y4523 = n16078 ;
  assign y4524 = ~n16081 ;
  assign y4525 = ~n16084 ;
  assign y4526 = ~n16086 ;
  assign y4527 = n16088 ;
  assign y4528 = ~n16093 ;
  assign y4529 = n16095 ;
  assign y4530 = ~1'b0 ;
  assign y4531 = n16096 ;
  assign y4532 = ~n16098 ;
  assign y4533 = n16099 ;
  assign y4534 = ~1'b0 ;
  assign y4535 = n16101 ;
  assign y4536 = n16108 ;
  assign y4537 = ~n16109 ;
  assign y4538 = ~n16111 ;
  assign y4539 = ~n16120 ;
  assign y4540 = ~n16123 ;
  assign y4541 = ~1'b0 ;
  assign y4542 = ~1'b0 ;
  assign y4543 = ~n16127 ;
  assign y4544 = ~n16132 ;
  assign y4545 = n16135 ;
  assign y4546 = n16137 ;
  assign y4547 = ~1'b0 ;
  assign y4548 = n16145 ;
  assign y4549 = ~n16151 ;
  assign y4550 = n16153 ;
  assign y4551 = n16154 ;
  assign y4552 = n16155 ;
  assign y4553 = n16156 ;
  assign y4554 = ~1'b0 ;
  assign y4555 = n16167 ;
  assign y4556 = ~n16168 ;
  assign y4557 = ~n16170 ;
  assign y4558 = n16174 ;
  assign y4559 = n16175 ;
  assign y4560 = n16176 ;
  assign y4561 = ~n16178 ;
  assign y4562 = n16182 ;
  assign y4563 = ~n16183 ;
  assign y4564 = n16188 ;
  assign y4565 = n16189 ;
  assign y4566 = n16203 ;
  assign y4567 = n16206 ;
  assign y4568 = n16207 ;
  assign y4569 = n6906 ;
  assign y4570 = n16212 ;
  assign y4571 = ~1'b0 ;
  assign y4572 = n16228 ;
  assign y4573 = n16235 ;
  assign y4574 = n16237 ;
  assign y4575 = ~1'b0 ;
  assign y4576 = n16243 ;
  assign y4577 = ~n16246 ;
  assign y4578 = ~n16251 ;
  assign y4579 = ~n16257 ;
  assign y4580 = ~1'b0 ;
  assign y4581 = n16260 ;
  assign y4582 = ~n16262 ;
  assign y4583 = n16267 ;
  assign y4584 = n16275 ;
  assign y4585 = ~n16278 ;
  assign y4586 = ~n16283 ;
  assign y4587 = ~n16290 ;
  assign y4588 = ~n16299 ;
  assign y4589 = ~n16302 ;
  assign y4590 = ~n16303 ;
  assign y4591 = ~1'b0 ;
  assign y4592 = ~n16306 ;
  assign y4593 = ~n16307 ;
  assign y4594 = n16309 ;
  assign y4595 = n16311 ;
  assign y4596 = ~1'b0 ;
  assign y4597 = n16315 ;
  assign y4598 = n16318 ;
  assign y4599 = ~n16322 ;
  assign y4600 = ~n16323 ;
  assign y4601 = n16326 ;
  assign y4602 = n16334 ;
  assign y4603 = n16337 ;
  assign y4604 = n16339 ;
  assign y4605 = ~n16343 ;
  assign y4606 = ~n16345 ;
  assign y4607 = n16348 ;
  assign y4608 = n16352 ;
  assign y4609 = ~1'b0 ;
  assign y4610 = ~n16353 ;
  assign y4611 = n16356 ;
  assign y4612 = n16357 ;
  assign y4613 = ~n16361 ;
  assign y4614 = ~n16367 ;
  assign y4615 = ~n16373 ;
  assign y4616 = ~1'b0 ;
  assign y4617 = n16374 ;
  assign y4618 = n16377 ;
  assign y4619 = ~1'b0 ;
  assign y4620 = n16380 ;
  assign y4621 = ~n16383 ;
  assign y4622 = n16384 ;
  assign y4623 = n16391 ;
  assign y4624 = n16395 ;
  assign y4625 = n16399 ;
  assign y4626 = ~1'b0 ;
  assign y4627 = ~n16401 ;
  assign y4628 = n16405 ;
  assign y4629 = ~1'b0 ;
  assign y4630 = n16414 ;
  assign y4631 = ~n16420 ;
  assign y4632 = ~n16423 ;
  assign y4633 = ~n16424 ;
  assign y4634 = n16425 ;
  assign y4635 = n16426 ;
  assign y4636 = n16427 ;
  assign y4637 = ~1'b0 ;
  assign y4638 = n16429 ;
  assign y4639 = ~n16431 ;
  assign y4640 = n16433 ;
  assign y4641 = ~n16446 ;
  assign y4642 = n16453 ;
  assign y4643 = n16455 ;
  assign y4644 = ~1'b0 ;
  assign y4645 = ~n16456 ;
  assign y4646 = ~n16461 ;
  assign y4647 = ~n16466 ;
  assign y4648 = ~n16468 ;
  assign y4649 = ~1'b0 ;
  assign y4650 = n16469 ;
  assign y4651 = ~n8082 ;
  assign y4652 = n16472 ;
  assign y4653 = ~n16473 ;
  assign y4654 = n16474 ;
  assign y4655 = ~n16475 ;
  assign y4656 = n3471 ;
  assign y4657 = ~n16476 ;
  assign y4658 = ~n16480 ;
  assign y4659 = ~n16484 ;
  assign y4660 = n16485 ;
  assign y4661 = ~n16489 ;
  assign y4662 = ~n16491 ;
  assign y4663 = n16499 ;
  assign y4664 = n16503 ;
  assign y4665 = ~n16508 ;
  assign y4666 = n16510 ;
  assign y4667 = n16512 ;
  assign y4668 = ~1'b0 ;
  assign y4669 = ~1'b0 ;
  assign y4670 = n16522 ;
  assign y4671 = ~n16531 ;
  assign y4672 = ~n16532 ;
  assign y4673 = n16539 ;
  assign y4674 = n16542 ;
  assign y4675 = ~n16543 ;
  assign y4676 = ~n16549 ;
  assign y4677 = n16553 ;
  assign y4678 = n16556 ;
  assign y4679 = n16558 ;
  assign y4680 = n16562 ;
  assign y4681 = n16564 ;
  assign y4682 = ~n16567 ;
  assign y4683 = n16568 ;
  assign y4684 = n16569 ;
  assign y4685 = n16572 ;
  assign y4686 = n16573 ;
  assign y4687 = ~1'b0 ;
  assign y4688 = n16575 ;
  assign y4689 = n16578 ;
  assign y4690 = ~n16582 ;
  assign y4691 = n16583 ;
  assign y4692 = ~n16588 ;
  assign y4693 = n16592 ;
  assign y4694 = ~1'b0 ;
  assign y4695 = n16593 ;
  assign y4696 = ~n16596 ;
  assign y4697 = n16599 ;
  assign y4698 = ~n16600 ;
  assign y4699 = ~n16604 ;
  assign y4700 = ~n16609 ;
  assign y4701 = ~n16611 ;
  assign y4702 = ~1'b0 ;
  assign y4703 = n16615 ;
  assign y4704 = n16616 ;
  assign y4705 = n16617 ;
  assign y4706 = ~1'b0 ;
  assign y4707 = n16620 ;
  assign y4708 = n16621 ;
  assign y4709 = n16629 ;
  assign y4710 = n16630 ;
  assign y4711 = ~n16632 ;
  assign y4712 = ~1'b0 ;
  assign y4713 = n16634 ;
  assign y4714 = n16639 ;
  assign y4715 = ~n16640 ;
  assign y4716 = n16641 ;
  assign y4717 = n16647 ;
  assign y4718 = ~n16654 ;
  assign y4719 = ~n16657 ;
  assign y4720 = ~n16661 ;
  assign y4721 = ~n16663 ;
  assign y4722 = ~n16664 ;
  assign y4723 = n16666 ;
  assign y4724 = ~n16670 ;
  assign y4725 = ~n16673 ;
  assign y4726 = n16688 ;
  assign y4727 = n16692 ;
  assign y4728 = n16693 ;
  assign y4729 = n16701 ;
  assign y4730 = n16702 ;
  assign y4731 = n16710 ;
  assign y4732 = n16711 ;
  assign y4733 = n16719 ;
  assign y4734 = ~n16726 ;
  assign y4735 = ~n16727 ;
  assign y4736 = n16730 ;
  assign y4737 = ~n16735 ;
  assign y4738 = ~1'b0 ;
  assign y4739 = ~n16737 ;
  assign y4740 = ~n16739 ;
  assign y4741 = n16741 ;
  assign y4742 = n16745 ;
  assign y4743 = n16747 ;
  assign y4744 = ~n16749 ;
  assign y4745 = n16753 ;
  assign y4746 = ~n16761 ;
  assign y4747 = n16771 ;
  assign y4748 = ~n16775 ;
  assign y4749 = n16778 ;
  assign y4750 = ~n16780 ;
  assign y4751 = ~n16782 ;
  assign y4752 = ~1'b0 ;
  assign y4753 = ~n16784 ;
  assign y4754 = ~1'b0 ;
  assign y4755 = n16785 ;
  assign y4756 = n16789 ;
  assign y4757 = ~n16800 ;
  assign y4758 = ~1'b0 ;
  assign y4759 = ~n16806 ;
  assign y4760 = ~n16810 ;
  assign y4761 = n16812 ;
  assign y4762 = n16814 ;
  assign y4763 = ~n16816 ;
  assign y4764 = ~n16818 ;
  assign y4765 = ~n16823 ;
  assign y4766 = ~n16827 ;
  assign y4767 = ~1'b0 ;
  assign y4768 = ~n16829 ;
  assign y4769 = ~n16830 ;
  assign y4770 = ~n16833 ;
  assign y4771 = ~n16834 ;
  assign y4772 = ~n16836 ;
  assign y4773 = ~n16839 ;
  assign y4774 = n16840 ;
  assign y4775 = ~n16842 ;
  assign y4776 = n16844 ;
  assign y4777 = ~1'b0 ;
  assign y4778 = ~1'b0 ;
  assign y4779 = ~1'b0 ;
  assign y4780 = ~n16845 ;
  assign y4781 = n16849 ;
  assign y4782 = ~1'b0 ;
  assign y4783 = ~1'b0 ;
  assign y4784 = n16852 ;
  assign y4785 = n16858 ;
  assign y4786 = ~n16860 ;
  assign y4787 = ~n16861 ;
  assign y4788 = ~n16866 ;
  assign y4789 = n16869 ;
  assign y4790 = n16870 ;
  assign y4791 = ~n16871 ;
  assign y4792 = ~1'b0 ;
  assign y4793 = ~1'b0 ;
  assign y4794 = ~n16875 ;
  assign y4795 = ~n16884 ;
  assign y4796 = n16886 ;
  assign y4797 = ~n16888 ;
  assign y4798 = ~n16895 ;
  assign y4799 = ~n16899 ;
  assign y4800 = ~n16902 ;
  assign y4801 = ~n16906 ;
  assign y4802 = n16907 ;
  assign y4803 = ~n16910 ;
  assign y4804 = ~n16917 ;
  assign y4805 = ~1'b0 ;
  assign y4806 = n16918 ;
  assign y4807 = ~n16920 ;
  assign y4808 = n16921 ;
  assign y4809 = ~n16925 ;
  assign y4810 = n16934 ;
  assign y4811 = ~n16936 ;
  assign y4812 = ~1'b0 ;
  assign y4813 = ~1'b0 ;
  assign y4814 = n16945 ;
  assign y4815 = n16948 ;
  assign y4816 = ~n16953 ;
  assign y4817 = ~n16963 ;
  assign y4818 = ~1'b0 ;
  assign y4819 = n16964 ;
  assign y4820 = ~n16965 ;
  assign y4821 = n16967 ;
  assign y4822 = ~1'b0 ;
  assign y4823 = n16969 ;
  assign y4824 = ~n16972 ;
  assign y4825 = ~n16975 ;
  assign y4826 = n16981 ;
  assign y4827 = ~n16986 ;
  assign y4828 = ~n16989 ;
  assign y4829 = n16991 ;
  assign y4830 = n17003 ;
  assign y4831 = ~n17008 ;
  assign y4832 = ~1'b0 ;
  assign y4833 = ~n17013 ;
  assign y4834 = n17017 ;
  assign y4835 = n17020 ;
  assign y4836 = n17021 ;
  assign y4837 = ~n17026 ;
  assign y4838 = n17029 ;
  assign y4839 = n17031 ;
  assign y4840 = n17033 ;
  assign y4841 = ~1'b0 ;
  assign y4842 = n17034 ;
  assign y4843 = n17036 ;
  assign y4844 = ~n17038 ;
  assign y4845 = ~1'b0 ;
  assign y4846 = ~1'b0 ;
  assign y4847 = ~1'b0 ;
  assign y4848 = ~1'b0 ;
  assign y4849 = ~n17040 ;
  assign y4850 = n17042 ;
  assign y4851 = n12152 ;
  assign y4852 = n17043 ;
  assign y4853 = ~n17044 ;
  assign y4854 = ~n17047 ;
  assign y4855 = n17050 ;
  assign y4856 = n17055 ;
  assign y4857 = ~n17056 ;
  assign y4858 = n17058 ;
  assign y4859 = ~n17062 ;
  assign y4860 = ~n17072 ;
  assign y4861 = ~n17073 ;
  assign y4862 = ~1'b0 ;
  assign y4863 = n17088 ;
  assign y4864 = ~1'b0 ;
  assign y4865 = ~1'b0 ;
  assign y4866 = n17091 ;
  assign y4867 = ~1'b0 ;
  assign y4868 = ~n17096 ;
  assign y4869 = ~n17100 ;
  assign y4870 = n17101 ;
  assign y4871 = n17105 ;
  assign y4872 = n17109 ;
  assign y4873 = ~n17114 ;
  assign y4874 = ~n17116 ;
  assign y4875 = ~n17119 ;
  assign y4876 = n17122 ;
  assign y4877 = ~1'b0 ;
  assign y4878 = ~n17125 ;
  assign y4879 = ~n17127 ;
  assign y4880 = ~n17132 ;
  assign y4881 = n17139 ;
  assign y4882 = ~n17140 ;
  assign y4883 = ~n17143 ;
  assign y4884 = ~n17148 ;
  assign y4885 = ~n17151 ;
  assign y4886 = n5195 ;
  assign y4887 = ~1'b0 ;
  assign y4888 = ~n17167 ;
  assign y4889 = n17169 ;
  assign y4890 = ~n17170 ;
  assign y4891 = n17172 ;
  assign y4892 = n17175 ;
  assign y4893 = ~n17176 ;
  assign y4894 = ~n17178 ;
  assign y4895 = ~1'b0 ;
  assign y4896 = n17180 ;
  assign y4897 = n17181 ;
  assign y4898 = n17186 ;
  assign y4899 = ~n17191 ;
  assign y4900 = n17193 ;
  assign y4901 = n17196 ;
  assign y4902 = ~1'b0 ;
  assign y4903 = ~1'b0 ;
  assign y4904 = n17200 ;
  assign y4905 = n17205 ;
  assign y4906 = ~n17207 ;
  assign y4907 = n17208 ;
  assign y4908 = n17210 ;
  assign y4909 = ~1'b0 ;
  assign y4910 = ~n17211 ;
  assign y4911 = ~n17215 ;
  assign y4912 = ~n17216 ;
  assign y4913 = n17219 ;
  assign y4914 = ~n17223 ;
  assign y4915 = ~n17226 ;
  assign y4916 = ~n17229 ;
  assign y4917 = ~n17231 ;
  assign y4918 = n17234 ;
  assign y4919 = ~n17236 ;
  assign y4920 = ~1'b0 ;
  assign y4921 = ~n3811 ;
  assign y4922 = n17239 ;
  assign y4923 = n17240 ;
  assign y4924 = ~1'b0 ;
  assign y4925 = ~n17241 ;
  assign y4926 = ~1'b0 ;
  assign y4927 = n17243 ;
  assign y4928 = n17244 ;
  assign y4929 = n17246 ;
  assign y4930 = n17248 ;
  assign y4931 = ~n17249 ;
  assign y4932 = n17253 ;
  assign y4933 = ~n17254 ;
  assign y4934 = 1'b0 ;
  assign y4935 = ~n17255 ;
  assign y4936 = ~n17257 ;
  assign y4937 = n17258 ;
  assign y4938 = ~1'b0 ;
  assign y4939 = ~1'b0 ;
  assign y4940 = ~n17262 ;
  assign y4941 = ~n17263 ;
  assign y4942 = ~n17269 ;
  assign y4943 = n17272 ;
  assign y4944 = n17274 ;
  assign y4945 = ~n17275 ;
  assign y4946 = n17277 ;
  assign y4947 = ~n17283 ;
  assign y4948 = 1'b0 ;
  assign y4949 = ~n17285 ;
  assign y4950 = n17287 ;
  assign y4951 = ~n17289 ;
  assign y4952 = ~n17294 ;
  assign y4953 = ~n17299 ;
  assign y4954 = n17305 ;
  assign y4955 = ~n17310 ;
  assign y4956 = n17311 ;
  assign y4957 = n17312 ;
  assign y4958 = n17315 ;
  assign y4959 = ~n17316 ;
  assign y4960 = ~n17330 ;
  assign y4961 = ~n17332 ;
  assign y4962 = ~n17339 ;
  assign y4963 = ~n17348 ;
  assign y4964 = ~n17352 ;
  assign y4965 = ~n17356 ;
  assign y4966 = ~n17358 ;
  assign y4967 = n17360 ;
  assign y4968 = ~n17361 ;
  assign y4969 = ~n17364 ;
  assign y4970 = ~n17366 ;
  assign y4971 = ~n17371 ;
  assign y4972 = ~n17372 ;
  assign y4973 = ~n17380 ;
  assign y4974 = n4376 ;
  assign y4975 = n17392 ;
  assign y4976 = ~n17395 ;
  assign y4977 = n17398 ;
  assign y4978 = ~n17400 ;
  assign y4979 = ~1'b0 ;
  assign y4980 = n17403 ;
  assign y4981 = n17409 ;
  assign y4982 = n17412 ;
  assign y4983 = n17413 ;
  assign y4984 = n17414 ;
  assign y4985 = ~n17417 ;
  assign y4986 = ~n17419 ;
  assign y4987 = ~n17420 ;
  assign y4988 = n17422 ;
  assign y4989 = n17425 ;
  assign y4990 = ~n17427 ;
  assign y4991 = ~1'b0 ;
  assign y4992 = ~n17428 ;
  assign y4993 = n17429 ;
  assign y4994 = ~n17437 ;
  assign y4995 = n17439 ;
  assign y4996 = ~n17444 ;
  assign y4997 = n17446 ;
  assign y4998 = ~1'b0 ;
  assign y4999 = ~n17451 ;
  assign y5000 = ~n17452 ;
  assign y5001 = n17454 ;
  assign y5002 = ~n17456 ;
  assign y5003 = ~n17457 ;
  assign y5004 = ~n17460 ;
  assign y5005 = n17462 ;
  assign y5006 = n17464 ;
  assign y5007 = n17466 ;
  assign y5008 = ~n17467 ;
  assign y5009 = ~n17468 ;
  assign y5010 = ~n1034 ;
  assign y5011 = n17469 ;
  assign y5012 = ~n17472 ;
  assign y5013 = ~n17474 ;
  assign y5014 = ~n17480 ;
  assign y5015 = n17485 ;
  assign y5016 = ~n14890 ;
  assign y5017 = n17499 ;
  assign y5018 = n17500 ;
  assign y5019 = ~n4374 ;
  assign y5020 = n17501 ;
  assign y5021 = ~n17502 ;
  assign y5022 = ~n17507 ;
  assign y5023 = ~n17510 ;
  assign y5024 = ~n14709 ;
  assign y5025 = n17514 ;
  assign y5026 = n7060 ;
  assign y5027 = ~n17516 ;
  assign y5028 = ~n17519 ;
  assign y5029 = ~n17525 ;
  assign y5030 = n17526 ;
  assign y5031 = ~n17527 ;
  assign y5032 = n17529 ;
  assign y5033 = ~1'b0 ;
  assign y5034 = n17530 ;
  assign y5035 = n17532 ;
  assign y5036 = ~n17533 ;
  assign y5037 = ~n17536 ;
  assign y5038 = ~n17538 ;
  assign y5039 = ~n17542 ;
  assign y5040 = ~1'b0 ;
  assign y5041 = n17544 ;
  assign y5042 = ~n17545 ;
  assign y5043 = ~n17549 ;
  assign y5044 = n17552 ;
  assign y5045 = ~n17554 ;
  assign y5046 = n17555 ;
  assign y5047 = n17561 ;
  assign y5048 = ~1'b0 ;
  assign y5049 = n17562 ;
  assign y5050 = ~n17564 ;
  assign y5051 = n17565 ;
  assign y5052 = n17567 ;
  assign y5053 = ~n17568 ;
  assign y5054 = ~1'b0 ;
  assign y5055 = n17570 ;
  assign y5056 = ~n17575 ;
  assign y5057 = n17581 ;
  assign y5058 = ~1'b0 ;
  assign y5059 = ~1'b0 ;
  assign y5060 = n2870 ;
  assign y5061 = ~n8740 ;
  assign y5062 = n17585 ;
  assign y5063 = n17586 ;
  assign y5064 = ~1'b0 ;
  assign y5065 = n17588 ;
  assign y5066 = ~n17595 ;
  assign y5067 = n17601 ;
  assign y5068 = n17606 ;
  assign y5069 = ~n17608 ;
  assign y5070 = ~1'b0 ;
  assign y5071 = n17614 ;
  assign y5072 = ~n17616 ;
  assign y5073 = ~n17622 ;
  assign y5074 = ~n17623 ;
  assign y5075 = ~n17624 ;
  assign y5076 = n17625 ;
  assign y5077 = n17630 ;
  assign y5078 = ~n17633 ;
  assign y5079 = n17637 ;
  assign y5080 = ~1'b0 ;
  assign y5081 = ~n17642 ;
  assign y5082 = ~n17646 ;
  assign y5083 = ~n17649 ;
  assign y5084 = ~n17652 ;
  assign y5085 = n17660 ;
  assign y5086 = ~n17663 ;
  assign y5087 = ~n17668 ;
  assign y5088 = n17674 ;
  assign y5089 = ~1'b0 ;
  assign y5090 = ~n17679 ;
  assign y5091 = n17682 ;
  assign y5092 = n17683 ;
  assign y5093 = n17684 ;
  assign y5094 = ~n17689 ;
  assign y5095 = ~n17690 ;
  assign y5096 = ~n17691 ;
  assign y5097 = ~n17694 ;
  assign y5098 = ~n17698 ;
  assign y5099 = ~n17706 ;
  assign y5100 = n17710 ;
  assign y5101 = ~n17712 ;
  assign y5102 = ~n17713 ;
  assign y5103 = ~n17714 ;
  assign y5104 = ~1'b0 ;
  assign y5105 = ~1'b0 ;
  assign y5106 = ~1'b0 ;
  assign y5107 = n17720 ;
  assign y5108 = n17724 ;
  assign y5109 = n17726 ;
  assign y5110 = ~n17728 ;
  assign y5111 = ~n17730 ;
  assign y5112 = ~n17731 ;
  assign y5113 = n17732 ;
  assign y5114 = n17734 ;
  assign y5115 = n17736 ;
  assign y5116 = n17743 ;
  assign y5117 = n3269 ;
  assign y5118 = ~1'b0 ;
  assign y5119 = n17744 ;
  assign y5120 = ~n17745 ;
  assign y5121 = n17747 ;
  assign y5122 = n17748 ;
  assign y5123 = n17750 ;
  assign y5124 = ~n17753 ;
  assign y5125 = ~n17754 ;
  assign y5126 = n17761 ;
  assign y5127 = ~n17765 ;
  assign y5128 = ~n17770 ;
  assign y5129 = n17775 ;
  assign y5130 = n17776 ;
  assign y5131 = n17781 ;
  assign y5132 = ~n17787 ;
  assign y5133 = ~n17788 ;
  assign y5134 = ~1'b0 ;
  assign y5135 = ~n17790 ;
  assign y5136 = n17791 ;
  assign y5137 = n17792 ;
  assign y5138 = n17794 ;
  assign y5139 = ~1'b0 ;
  assign y5140 = ~n17795 ;
  assign y5141 = n17796 ;
  assign y5142 = n17799 ;
  assign y5143 = ~n17808 ;
  assign y5144 = n17814 ;
  assign y5145 = n17817 ;
  assign y5146 = ~n17820 ;
  assign y5147 = ~n17821 ;
  assign y5148 = ~n17838 ;
  assign y5149 = ~n17839 ;
  assign y5150 = n11528 ;
  assign y5151 = n17842 ;
  assign y5152 = n17843 ;
  assign y5153 = ~n17845 ;
  assign y5154 = n17846 ;
  assign y5155 = n17847 ;
  assign y5156 = ~n17851 ;
  assign y5157 = ~1'b0 ;
  assign y5158 = n17859 ;
  assign y5159 = ~n17860 ;
  assign y5160 = n17862 ;
  assign y5161 = ~n17865 ;
  assign y5162 = ~n17866 ;
  assign y5163 = n17868 ;
  assign y5164 = n17871 ;
  assign y5165 = n17873 ;
  assign y5166 = n17874 ;
  assign y5167 = n17879 ;
  assign y5168 = ~n17880 ;
  assign y5169 = n17884 ;
  assign y5170 = ~n17886 ;
  assign y5171 = ~n17888 ;
  assign y5172 = ~n17890 ;
  assign y5173 = ~n17891 ;
  assign y5174 = ~n17896 ;
  assign y5175 = ~n17899 ;
  assign y5176 = n17900 ;
  assign y5177 = ~n17901 ;
  assign y5178 = ~1'b0 ;
  assign y5179 = ~n17905 ;
  assign y5180 = ~1'b0 ;
  assign y5181 = n17906 ;
  assign y5182 = ~n17907 ;
  assign y5183 = ~1'b0 ;
  assign y5184 = ~n17912 ;
  assign y5185 = n17913 ;
  assign y5186 = n17916 ;
  assign y5187 = ~n17917 ;
  assign y5188 = n17920 ;
  assign y5189 = ~1'b0 ;
  assign y5190 = ~n17921 ;
  assign y5191 = n17922 ;
  assign y5192 = n17923 ;
  assign y5193 = n17924 ;
  assign y5194 = n17926 ;
  assign y5195 = ~n17928 ;
  assign y5196 = n17931 ;
  assign y5197 = n17932 ;
  assign y5198 = n17934 ;
  assign y5199 = n17935 ;
  assign y5200 = ~n17936 ;
  assign y5201 = n17937 ;
  assign y5202 = n17938 ;
  assign y5203 = ~1'b0 ;
  assign y5204 = ~n17942 ;
  assign y5205 = n17945 ;
  assign y5206 = n17949 ;
  assign y5207 = ~n17951 ;
  assign y5208 = ~1'b0 ;
  assign y5209 = ~n17953 ;
  assign y5210 = ~n17960 ;
  assign y5211 = n17961 ;
  assign y5212 = ~n17971 ;
  assign y5213 = ~n17973 ;
  assign y5214 = n17975 ;
  assign y5215 = ~n17978 ;
  assign y5216 = n17985 ;
  assign y5217 = ~n17987 ;
  assign y5218 = ~n17991 ;
  assign y5219 = n17994 ;
  assign y5220 = ~n17999 ;
  assign y5221 = ~1'b0 ;
  assign y5222 = n18001 ;
  assign y5223 = ~n18004 ;
  assign y5224 = n18007 ;
  assign y5225 = ~n18010 ;
  assign y5226 = ~n18018 ;
  assign y5227 = n18019 ;
  assign y5228 = ~n18029 ;
  assign y5229 = n18032 ;
  assign y5230 = ~n18036 ;
  assign y5231 = ~n18037 ;
  assign y5232 = n18047 ;
  assign y5233 = n18051 ;
  assign y5234 = n18056 ;
  assign y5235 = ~n18061 ;
  assign y5236 = ~n18065 ;
  assign y5237 = ~n18067 ;
  assign y5238 = ~n18068 ;
  assign y5239 = n18071 ;
  assign y5240 = ~n18080 ;
  assign y5241 = ~n18085 ;
  assign y5242 = ~n18086 ;
  assign y5243 = ~n18095 ;
  assign y5244 = ~n18100 ;
  assign y5245 = ~n18102 ;
  assign y5246 = ~n18103 ;
  assign y5247 = ~1'b0 ;
  assign y5248 = ~n18110 ;
  assign y5249 = n18111 ;
  assign y5250 = n18113 ;
  assign y5251 = n18117 ;
  assign y5252 = n18118 ;
  assign y5253 = n18120 ;
  assign y5254 = ~n18123 ;
  assign y5255 = n18124 ;
  assign y5256 = ~n18125 ;
  assign y5257 = n18130 ;
  assign y5258 = ~1'b0 ;
  assign y5259 = ~1'b0 ;
  assign y5260 = n18132 ;
  assign y5261 = n18136 ;
  assign y5262 = n18137 ;
  assign y5263 = ~n18141 ;
  assign y5264 = ~n18142 ;
  assign y5265 = ~1'b0 ;
  assign y5266 = ~n18155 ;
  assign y5267 = n18157 ;
  assign y5268 = n18159 ;
  assign y5269 = ~n18164 ;
  assign y5270 = ~n18166 ;
  assign y5271 = ~n18173 ;
  assign y5272 = ~n18174 ;
  assign y5273 = ~n18178 ;
  assign y5274 = ~1'b0 ;
  assign y5275 = ~n18179 ;
  assign y5276 = n18183 ;
  assign y5277 = n18188 ;
  assign y5278 = ~n18189 ;
  assign y5279 = n18192 ;
  assign y5280 = n18193 ;
  assign y5281 = ~n18195 ;
  assign y5282 = n18200 ;
  assign y5283 = ~n18201 ;
  assign y5284 = ~n18203 ;
  assign y5285 = ~n18206 ;
  assign y5286 = ~1'b0 ;
  assign y5287 = n18208 ;
  assign y5288 = n18209 ;
  assign y5289 = ~n18211 ;
  assign y5290 = ~n18213 ;
  assign y5291 = ~n18215 ;
  assign y5292 = n18218 ;
  assign y5293 = ~n18227 ;
  assign y5294 = n18228 ;
  assign y5295 = ~n18230 ;
  assign y5296 = ~n18234 ;
  assign y5297 = ~1'b0 ;
  assign y5298 = ~1'b0 ;
  assign y5299 = n18235 ;
  assign y5300 = ~n18237 ;
  assign y5301 = n18239 ;
  assign y5302 = ~n18242 ;
  assign y5303 = ~n18243 ;
  assign y5304 = n18248 ;
  assign y5305 = ~n18258 ;
  assign y5306 = ~n18261 ;
  assign y5307 = ~n18267 ;
  assign y5308 = ~1'b0 ;
  assign y5309 = ~1'b0 ;
  assign y5310 = ~n18272 ;
  assign y5311 = ~n18273 ;
  assign y5312 = n18276 ;
  assign y5313 = ~n18283 ;
  assign y5314 = ~n18285 ;
  assign y5315 = n18291 ;
  assign y5316 = ~n18293 ;
  assign y5317 = n18295 ;
  assign y5318 = ~n18296 ;
  assign y5319 = n18299 ;
  assign y5320 = ~n18300 ;
  assign y5321 = n18303 ;
  assign y5322 = ~n18304 ;
  assign y5323 = ~n18306 ;
  assign y5324 = n18311 ;
  assign y5325 = ~1'b0 ;
  assign y5326 = ~n18315 ;
  assign y5327 = n18318 ;
  assign y5328 = n18320 ;
  assign y5329 = ~n18321 ;
  assign y5330 = n18326 ;
  assign y5331 = ~1'b0 ;
  assign y5332 = ~n18327 ;
  assign y5333 = n18332 ;
  assign y5334 = n18333 ;
  assign y5335 = ~1'b0 ;
  assign y5336 = ~n18336 ;
  assign y5337 = n18337 ;
  assign y5338 = ~1'b0 ;
  assign y5339 = n18338 ;
  assign y5340 = n18339 ;
  assign y5341 = n994 ;
  assign y5342 = ~1'b0 ;
  assign y5343 = ~n18341 ;
  assign y5344 = n18343 ;
  assign y5345 = ~n18345 ;
  assign y5346 = ~1'b0 ;
  assign y5347 = n18347 ;
  assign y5348 = ~n18350 ;
  assign y5349 = ~n6246 ;
  assign y5350 = n18352 ;
  assign y5351 = n18353 ;
  assign y5352 = ~n18354 ;
  assign y5353 = n18357 ;
  assign y5354 = ~1'b0 ;
  assign y5355 = ~1'b0 ;
  assign y5356 = ~n18359 ;
  assign y5357 = ~n18364 ;
  assign y5358 = ~n18372 ;
  assign y5359 = ~n18373 ;
  assign y5360 = n18374 ;
  assign y5361 = n18379 ;
  assign y5362 = ~n18381 ;
  assign y5363 = n18385 ;
  assign y5364 = n18388 ;
  assign y5365 = n18398 ;
  assign y5366 = ~1'b0 ;
  assign y5367 = ~1'b0 ;
  assign y5368 = n18399 ;
  assign y5369 = n18405 ;
  assign y5370 = ~n18408 ;
  assign y5371 = n18409 ;
  assign y5372 = ~n18411 ;
  assign y5373 = ~n18418 ;
  assign y5374 = n18419 ;
  assign y5375 = ~n18421 ;
  assign y5376 = ~n18425 ;
  assign y5377 = n18430 ;
  assign y5378 = n18431 ;
  assign y5379 = n18445 ;
  assign y5380 = ~n18447 ;
  assign y5381 = ~n18458 ;
  assign y5382 = ~1'b0 ;
  assign y5383 = ~n18460 ;
  assign y5384 = ~n18463 ;
  assign y5385 = n18470 ;
  assign y5386 = ~n18471 ;
  assign y5387 = n18475 ;
  assign y5388 = n18476 ;
  assign y5389 = ~n18477 ;
  assign y5390 = n18478 ;
  assign y5391 = ~n18483 ;
  assign y5392 = n18488 ;
  assign y5393 = ~n18493 ;
  assign y5394 = n18499 ;
  assign y5395 = ~n18502 ;
  assign y5396 = n18507 ;
  assign y5397 = ~n18508 ;
  assign y5398 = ~n18509 ;
  assign y5399 = n18512 ;
  assign y5400 = ~n18515 ;
  assign y5401 = ~n18516 ;
  assign y5402 = ~1'b0 ;
  assign y5403 = n18519 ;
  assign y5404 = n18520 ;
  assign y5405 = n18523 ;
  assign y5406 = ~n18524 ;
  assign y5407 = n18526 ;
  assign y5408 = ~1'b0 ;
  assign y5409 = n18530 ;
  assign y5410 = ~1'b0 ;
  assign y5411 = n18533 ;
  assign y5412 = n18535 ;
  assign y5413 = ~n18539 ;
  assign y5414 = n18542 ;
  assign y5415 = ~n18544 ;
  assign y5416 = n18549 ;
  assign y5417 = n18555 ;
  assign y5418 = n18556 ;
  assign y5419 = ~n18558 ;
  assign y5420 = n18559 ;
  assign y5421 = ~n18562 ;
  assign y5422 = ~n18567 ;
  assign y5423 = ~n18572 ;
  assign y5424 = ~n18573 ;
  assign y5425 = ~n18575 ;
  assign y5426 = ~n18582 ;
  assign y5427 = ~1'b0 ;
  assign y5428 = ~n18584 ;
  assign y5429 = n18592 ;
  assign y5430 = n18593 ;
  assign y5431 = ~1'b0 ;
  assign y5432 = 1'b0 ;
  assign y5433 = n18594 ;
  assign y5434 = n18596 ;
  assign y5435 = n18597 ;
  assign y5436 = ~n18600 ;
  assign y5437 = n18605 ;
  assign y5438 = n8067 ;
  assign y5439 = n18607 ;
  assign y5440 = n18608 ;
  assign y5441 = ~n18610 ;
  assign y5442 = ~1'b0 ;
  assign y5443 = ~1'b0 ;
  assign y5444 = ~1'b0 ;
  assign y5445 = n18611 ;
  assign y5446 = n18613 ;
  assign y5447 = n18617 ;
  assign y5448 = ~n18622 ;
  assign y5449 = n18628 ;
  assign y5450 = ~n18630 ;
  assign y5451 = n18633 ;
  assign y5452 = n18634 ;
  assign y5453 = ~n18638 ;
  assign y5454 = n18640 ;
  assign y5455 = ~n18642 ;
  assign y5456 = ~n18643 ;
  assign y5457 = n18648 ;
  assign y5458 = n18653 ;
  assign y5459 = ~n18654 ;
  assign y5460 = n18657 ;
  assign y5461 = ~n18662 ;
  assign y5462 = ~n18666 ;
  assign y5463 = ~n18668 ;
  assign y5464 = ~n18669 ;
  assign y5465 = ~n18670 ;
  assign y5466 = ~n18673 ;
  assign y5467 = ~1'b0 ;
  assign y5468 = n18675 ;
  assign y5469 = ~n18677 ;
  assign y5470 = ~1'b0 ;
  assign y5471 = ~n18679 ;
  assign y5472 = ~1'b0 ;
  assign y5473 = ~n18682 ;
  assign y5474 = ~n18686 ;
  assign y5475 = ~1'b0 ;
  assign y5476 = n18687 ;
  assign y5477 = ~n18693 ;
  assign y5478 = ~n18695 ;
  assign y5479 = ~n18700 ;
  assign y5480 = n18702 ;
  assign y5481 = n18703 ;
  assign y5482 = n18708 ;
  assign y5483 = ~n18710 ;
  assign y5484 = n18715 ;
  assign y5485 = ~n18718 ;
  assign y5486 = n18721 ;
  assign y5487 = ~n18722 ;
  assign y5488 = ~n18728 ;
  assign y5489 = n18730 ;
  assign y5490 = ~1'b0 ;
  assign y5491 = ~n18735 ;
  assign y5492 = ~n18742 ;
  assign y5493 = ~n18743 ;
  assign y5494 = ~n18744 ;
  assign y5495 = n18746 ;
  assign y5496 = 1'b0 ;
  assign y5497 = n18748 ;
  assign y5498 = n18750 ;
  assign y5499 = n18757 ;
  assign y5500 = ~n18765 ;
  assign y5501 = n18766 ;
  assign y5502 = n18770 ;
  assign y5503 = ~1'b0 ;
  assign y5504 = ~1'b0 ;
  assign y5505 = ~n18779 ;
  assign y5506 = n15027 ;
  assign y5507 = ~n18780 ;
  assign y5508 = ~n18781 ;
  assign y5509 = n18783 ;
  assign y5510 = ~n18785 ;
  assign y5511 = ~n18786 ;
  assign y5512 = ~n18788 ;
  assign y5513 = ~n18789 ;
  assign y5514 = n18793 ;
  assign y5515 = n18794 ;
  assign y5516 = n18797 ;
  assign y5517 = n18799 ;
  assign y5518 = ~n18801 ;
  assign y5519 = n18803 ;
  assign y5520 = ~1'b0 ;
  assign y5521 = ~n18804 ;
  assign y5522 = ~n18809 ;
  assign y5523 = ~n18816 ;
  assign y5524 = ~n18819 ;
  assign y5525 = n18822 ;
  assign y5526 = n18825 ;
  assign y5527 = ~n18831 ;
  assign y5528 = ~n18832 ;
  assign y5529 = n18840 ;
  assign y5530 = ~n18845 ;
  assign y5531 = n18849 ;
  assign y5532 = ~1'b0 ;
  assign y5533 = ~1'b0 ;
  assign y5534 = ~n18854 ;
  assign y5535 = n18855 ;
  assign y5536 = ~n18859 ;
  assign y5537 = ~n18860 ;
  assign y5538 = ~1'b0 ;
  assign y5539 = ~n18863 ;
  assign y5540 = n18871 ;
  assign y5541 = n18873 ;
  assign y5542 = ~n18877 ;
  assign y5543 = ~n18879 ;
  assign y5544 = ~1'b0 ;
  assign y5545 = n18881 ;
  assign y5546 = n18884 ;
  assign y5547 = n18885 ;
  assign y5548 = ~n18894 ;
  assign y5549 = ~n18896 ;
  assign y5550 = ~n18899 ;
  assign y5551 = ~1'b0 ;
  assign y5552 = n18906 ;
  assign y5553 = n18910 ;
  assign y5554 = n18914 ;
  assign y5555 = n18916 ;
  assign y5556 = ~n18922 ;
  assign y5557 = n18925 ;
  assign y5558 = ~n18926 ;
  assign y5559 = n18927 ;
  assign y5560 = n18929 ;
  assign y5561 = ~n18931 ;
  assign y5562 = n18941 ;
  assign y5563 = ~n18942 ;
  assign y5564 = ~n18947 ;
  assign y5565 = n18950 ;
  assign y5566 = n18951 ;
  assign y5567 = ~n18954 ;
  assign y5568 = ~n18957 ;
  assign y5569 = n18959 ;
  assign y5570 = n18963 ;
  assign y5571 = ~n18968 ;
  assign y5572 = ~n18969 ;
  assign y5573 = n18972 ;
  assign y5574 = ~n18973 ;
  assign y5575 = n18974 ;
  assign y5576 = n18976 ;
  assign y5577 = ~1'b0 ;
  assign y5578 = n18977 ;
  assign y5579 = 1'b0 ;
  assign y5580 = ~n18979 ;
  assign y5581 = ~1'b0 ;
  assign y5582 = n18980 ;
  assign y5583 = n18982 ;
  assign y5584 = ~n18985 ;
  assign y5585 = ~1'b0 ;
  assign y5586 = ~n18987 ;
  assign y5587 = ~n18990 ;
  assign y5588 = n18993 ;
  assign y5589 = ~1'b0 ;
  assign y5590 = ~n8934 ;
  assign y5591 = n18996 ;
  assign y5592 = ~n19000 ;
  assign y5593 = ~n19004 ;
  assign y5594 = n19007 ;
  assign y5595 = ~1'b0 ;
  assign y5596 = ~1'b0 ;
  assign y5597 = ~n19008 ;
  assign y5598 = n19009 ;
  assign y5599 = ~n19011 ;
  assign y5600 = ~n19014 ;
  assign y5601 = n19015 ;
  assign y5602 = ~n19018 ;
  assign y5603 = n19028 ;
  assign y5604 = n19033 ;
  assign y5605 = ~n19034 ;
  assign y5606 = n19047 ;
  assign y5607 = n19049 ;
  assign y5608 = n19053 ;
  assign y5609 = n19056 ;
  assign y5610 = ~n19058 ;
  assign y5611 = ~n19062 ;
  assign y5612 = ~1'b0 ;
  assign y5613 = n1450 ;
  assign y5614 = ~n19067 ;
  assign y5615 = ~n19070 ;
  assign y5616 = ~n19074 ;
  assign y5617 = ~n19076 ;
  assign y5618 = ~1'b0 ;
  assign y5619 = n19077 ;
  assign y5620 = ~1'b0 ;
  assign y5621 = ~n19080 ;
  assign y5622 = n19082 ;
  assign y5623 = n19083 ;
  assign y5624 = ~n19084 ;
  assign y5625 = ~1'b0 ;
  assign y5626 = ~n19085 ;
  assign y5627 = n19086 ;
  assign y5628 = n19088 ;
  assign y5629 = n19093 ;
  assign y5630 = ~n19097 ;
  assign y5631 = n19100 ;
  assign y5632 = n19101 ;
  assign y5633 = n19102 ;
  assign y5634 = n19105 ;
  assign y5635 = n19106 ;
  assign y5636 = n19108 ;
  assign y5637 = ~n19109 ;
  assign y5638 = ~n19114 ;
  assign y5639 = n19116 ;
  assign y5640 = ~1'b0 ;
  assign y5641 = ~n19120 ;
  assign y5642 = n19121 ;
  assign y5643 = ~n19123 ;
  assign y5644 = n19126 ;
  assign y5645 = n19128 ;
  assign y5646 = ~n19129 ;
  assign y5647 = ~1'b0 ;
  assign y5648 = ~n19132 ;
  assign y5649 = ~n19133 ;
  assign y5650 = ~n19137 ;
  assign y5651 = n19139 ;
  assign y5652 = ~1'b0 ;
  assign y5653 = n19141 ;
  assign y5654 = ~n19143 ;
  assign y5655 = ~n19147 ;
  assign y5656 = n19149 ;
  assign y5657 = n19151 ;
  assign y5658 = ~n19152 ;
  assign y5659 = ~n19154 ;
  assign y5660 = ~n19156 ;
  assign y5661 = n19159 ;
  assign y5662 = n19160 ;
  assign y5663 = n19163 ;
  assign y5664 = n19171 ;
  assign y5665 = n19173 ;
  assign y5666 = n19174 ;
  assign y5667 = ~n19183 ;
  assign y5668 = ~n19185 ;
  assign y5669 = n19187 ;
  assign y5670 = ~n19188 ;
  assign y5671 = n19189 ;
  assign y5672 = ~n19191 ;
  assign y5673 = ~n19193 ;
  assign y5674 = ~n19195 ;
  assign y5675 = ~n19199 ;
  assign y5676 = n19201 ;
  assign y5677 = ~n19202 ;
  assign y5678 = n19206 ;
  assign y5679 = ~1'b0 ;
  assign y5680 = ~1'b0 ;
  assign y5681 = ~n19209 ;
  assign y5682 = ~n19210 ;
  assign y5683 = n19214 ;
  assign y5684 = ~1'b0 ;
  assign y5685 = ~1'b0 ;
  assign y5686 = ~n19216 ;
  assign y5687 = ~n19222 ;
  assign y5688 = ~n19223 ;
  assign y5689 = ~n19225 ;
  assign y5690 = ~n19227 ;
  assign y5691 = ~1'b0 ;
  assign y5692 = n19231 ;
  assign y5693 = ~n19234 ;
  assign y5694 = ~n19237 ;
  assign y5695 = n19244 ;
  assign y5696 = ~n19247 ;
  assign y5697 = n19249 ;
  assign y5698 = n19250 ;
  assign y5699 = ~n19255 ;
  assign y5700 = n19257 ;
  assign y5701 = n19258 ;
  assign y5702 = n19259 ;
  assign y5703 = ~1'b0 ;
  assign y5704 = n19263 ;
  assign y5705 = ~n19270 ;
  assign y5706 = ~n19275 ;
  assign y5707 = n19282 ;
  assign y5708 = ~n19288 ;
  assign y5709 = n19289 ;
  assign y5710 = ~1'b0 ;
  assign y5711 = ~1'b0 ;
  assign y5712 = n19291 ;
  assign y5713 = n19293 ;
  assign y5714 = ~n19300 ;
  assign y5715 = n19301 ;
  assign y5716 = ~n19309 ;
  assign y5717 = n19310 ;
  assign y5718 = ~n19311 ;
  assign y5719 = n19321 ;
  assign y5720 = ~n19322 ;
  assign y5721 = ~n19323 ;
  assign y5722 = ~n19324 ;
  assign y5723 = ~n19326 ;
  assign y5724 = n19328 ;
  assign y5725 = n19329 ;
  assign y5726 = n19331 ;
  assign y5727 = n19332 ;
  assign y5728 = ~n19335 ;
  assign y5729 = ~n19339 ;
  assign y5730 = n19340 ;
  assign y5731 = n19341 ;
  assign y5732 = ~n19342 ;
  assign y5733 = ~n19344 ;
  assign y5734 = n19345 ;
  assign y5735 = ~n19358 ;
  assign y5736 = ~n19360 ;
  assign y5737 = ~1'b0 ;
  assign y5738 = ~n19361 ;
  assign y5739 = n19363 ;
  assign y5740 = ~n19364 ;
  assign y5741 = n19365 ;
  assign y5742 = n19366 ;
  assign y5743 = ~n19368 ;
  assign y5744 = n19370 ;
  assign y5745 = ~1'b0 ;
  assign y5746 = ~n19376 ;
  assign y5747 = 1'b0 ;
  assign y5748 = n19385 ;
  assign y5749 = n19388 ;
  assign y5750 = n19390 ;
  assign y5751 = ~1'b0 ;
  assign y5752 = ~n19391 ;
  assign y5753 = ~n19396 ;
  assign y5754 = ~n19397 ;
  assign y5755 = n19399 ;
  assign y5756 = ~n19407 ;
  assign y5757 = ~n19408 ;
  assign y5758 = n19412 ;
  assign y5759 = 1'b0 ;
  assign y5760 = n19422 ;
  assign y5761 = ~n19428 ;
  assign y5762 = ~n19430 ;
  assign y5763 = ~n19435 ;
  assign y5764 = ~n19438 ;
  assign y5765 = n19440 ;
  assign y5766 = n19444 ;
  assign y5767 = ~1'b0 ;
  assign y5768 = ~n19445 ;
  assign y5769 = ~1'b0 ;
  assign y5770 = ~n19447 ;
  assign y5771 = n19453 ;
  assign y5772 = ~1'b0 ;
  assign y5773 = n19460 ;
  assign y5774 = ~n19464 ;
  assign y5775 = n19465 ;
  assign y5776 = ~1'b0 ;
  assign y5777 = ~n19467 ;
  assign y5778 = n19469 ;
  assign y5779 = ~n19472 ;
  assign y5780 = n19473 ;
  assign y5781 = ~n19485 ;
  assign y5782 = n19493 ;
  assign y5783 = ~n19497 ;
  assign y5784 = ~n19503 ;
  assign y5785 = n19504 ;
  assign y5786 = n19506 ;
  assign y5787 = n19520 ;
  assign y5788 = n19522 ;
  assign y5789 = ~n19527 ;
  assign y5790 = ~1'b0 ;
  assign y5791 = n19530 ;
  assign y5792 = n19531 ;
  assign y5793 = n19535 ;
  assign y5794 = n19538 ;
  assign y5795 = ~n19540 ;
  assign y5796 = n19542 ;
  assign y5797 = n19549 ;
  assign y5798 = ~n19551 ;
  assign y5799 = n19554 ;
  assign y5800 = ~n19555 ;
  assign y5801 = ~n19559 ;
  assign y5802 = n19560 ;
  assign y5803 = ~n19562 ;
  assign y5804 = ~n19567 ;
  assign y5805 = n19571 ;
  assign y5806 = ~n19573 ;
  assign y5807 = n19574 ;
  assign y5808 = n19582 ;
  assign y5809 = ~n19589 ;
  assign y5810 = ~n19591 ;
  assign y5811 = ~n19594 ;
  assign y5812 = n19600 ;
  assign y5813 = n19601 ;
  assign y5814 = ~n19603 ;
  assign y5815 = n19605 ;
  assign y5816 = ~1'b0 ;
  assign y5817 = n19607 ;
  assign y5818 = n19610 ;
  assign y5819 = n19611 ;
  assign y5820 = ~n19617 ;
  assign y5821 = n19624 ;
  assign y5822 = n19627 ;
  assign y5823 = ~1'b0 ;
  assign y5824 = ~1'b0 ;
  assign y5825 = ~n17749 ;
  assign y5826 = ~n19638 ;
  assign y5827 = ~n19639 ;
  assign y5828 = ~n19640 ;
  assign y5829 = n19641 ;
  assign y5830 = ~n19647 ;
  assign y5831 = n19651 ;
  assign y5832 = ~n19653 ;
  assign y5833 = n19656 ;
  assign y5834 = ~n19657 ;
  assign y5835 = ~n19660 ;
  assign y5836 = ~n19667 ;
  assign y5837 = ~n19669 ;
  assign y5838 = ~1'b0 ;
  assign y5839 = ~n19673 ;
  assign y5840 = n19675 ;
  assign y5841 = n19680 ;
  assign y5842 = ~n19681 ;
  assign y5843 = ~n19682 ;
  assign y5844 = ~n19687 ;
  assign y5845 = n19688 ;
  assign y5846 = n19689 ;
  assign y5847 = ~1'b0 ;
  assign y5848 = n19694 ;
  assign y5849 = ~n19695 ;
  assign y5850 = ~n19701 ;
  assign y5851 = ~n19704 ;
  assign y5852 = n19705 ;
  assign y5853 = ~n19708 ;
  assign y5854 = n19712 ;
  assign y5855 = ~n19713 ;
  assign y5856 = n19715 ;
  assign y5857 = n19718 ;
  assign y5858 = ~n19723 ;
  assign y5859 = n19724 ;
  assign y5860 = n19727 ;
  assign y5861 = n19732 ;
  assign y5862 = ~n19735 ;
  assign y5863 = n19740 ;
  assign y5864 = ~n19742 ;
  assign y5865 = ~n19744 ;
  assign y5866 = n19745 ;
  assign y5867 = n19746 ;
  assign y5868 = ~n19749 ;
  assign y5869 = ~1'b0 ;
  assign y5870 = ~n19751 ;
  assign y5871 = ~n19754 ;
  assign y5872 = ~1'b0 ;
  assign y5873 = ~n19756 ;
  assign y5874 = n19758 ;
  assign y5875 = n19759 ;
  assign y5876 = ~n19764 ;
  assign y5877 = ~n19767 ;
  assign y5878 = ~n19770 ;
  assign y5879 = n19772 ;
  assign y5880 = ~1'b0 ;
  assign y5881 = n19773 ;
  assign y5882 = ~n19777 ;
  assign y5883 = n19778 ;
  assign y5884 = ~n19779 ;
  assign y5885 = n19781 ;
  assign y5886 = n19785 ;
  assign y5887 = n19786 ;
  assign y5888 = ~n19789 ;
  assign y5889 = n19790 ;
  assign y5890 = ~n19797 ;
  assign y5891 = ~n19799 ;
  assign y5892 = n19802 ;
  assign y5893 = n19806 ;
  assign y5894 = ~n19809 ;
  assign y5895 = ~n19812 ;
  assign y5896 = n19818 ;
  assign y5897 = n19820 ;
  assign y5898 = ~n19825 ;
  assign y5899 = ~n19830 ;
  assign y5900 = ~1'b0 ;
  assign y5901 = ~1'b0 ;
  assign y5902 = ~n19832 ;
  assign y5903 = n19834 ;
  assign y5904 = ~n19841 ;
  assign y5905 = ~n19842 ;
  assign y5906 = n19843 ;
  assign y5907 = ~1'b0 ;
  assign y5908 = ~n19849 ;
  assign y5909 = n19852 ;
  assign y5910 = ~n19855 ;
  assign y5911 = n19856 ;
  assign y5912 = n19857 ;
  assign y5913 = ~n19864 ;
  assign y5914 = ~n19866 ;
  assign y5915 = ~n19872 ;
  assign y5916 = ~n19874 ;
  assign y5917 = n19877 ;
  assign y5918 = ~n19879 ;
  assign y5919 = n19881 ;
  assign y5920 = ~n19882 ;
  assign y5921 = ~n19884 ;
  assign y5922 = ~1'b0 ;
  assign y5923 = n19892 ;
  assign y5924 = ~n19899 ;
  assign y5925 = ~1'b0 ;
  assign y5926 = ~n19904 ;
  assign y5927 = n19908 ;
  assign y5928 = n19912 ;
  assign y5929 = ~n19916 ;
  assign y5930 = ~n19918 ;
  assign y5931 = n15210 ;
  assign y5932 = n19922 ;
  assign y5933 = ~n19925 ;
  assign y5934 = ~n19927 ;
  assign y5935 = n19929 ;
  assign y5936 = ~1'b0 ;
  assign y5937 = ~1'b0 ;
  assign y5938 = ~n19930 ;
  assign y5939 = ~n8331 ;
  assign y5940 = ~1'b0 ;
  assign y5941 = n19934 ;
  assign y5942 = n19936 ;
  assign y5943 = ~1'b0 ;
  assign y5944 = ~n19938 ;
  assign y5945 = ~n19939 ;
  assign y5946 = ~n19940 ;
  assign y5947 = n19942 ;
  assign y5948 = ~n19944 ;
  assign y5949 = ~n19948 ;
  assign y5950 = ~n19953 ;
  assign y5951 = n19956 ;
  assign y5952 = ~n19961 ;
  assign y5953 = n19962 ;
  assign y5954 = ~n19965 ;
  assign y5955 = ~n19969 ;
  assign y5956 = n19973 ;
  assign y5957 = ~n19975 ;
  assign y5958 = n5730 ;
  assign y5959 = n19976 ;
  assign y5960 = ~n19977 ;
  assign y5961 = ~1'b0 ;
  assign y5962 = n19979 ;
  assign y5963 = ~n19984 ;
  assign y5964 = ~n19988 ;
  assign y5965 = ~n19989 ;
  assign y5966 = n19991 ;
  assign y5967 = n19993 ;
  assign y5968 = n20000 ;
  assign y5969 = ~n20003 ;
  assign y5970 = ~n20010 ;
  assign y5971 = ~1'b0 ;
  assign y5972 = n20011 ;
  assign y5973 = ~n20016 ;
  assign y5974 = n11961 ;
  assign y5975 = ~n20017 ;
  assign y5976 = ~1'b0 ;
  assign y5977 = 1'b0 ;
  assign y5978 = n20018 ;
  assign y5979 = ~n20019 ;
  assign y5980 = ~n20024 ;
  assign y5981 = ~1'b0 ;
  assign y5982 = ~n20025 ;
  assign y5983 = n20029 ;
  assign y5984 = n20030 ;
  assign y5985 = n20034 ;
  assign y5986 = n20038 ;
  assign y5987 = ~n20042 ;
  assign y5988 = n20053 ;
  assign y5989 = ~n20054 ;
  assign y5990 = ~n20055 ;
  assign y5991 = n20060 ;
  assign y5992 = ~n20065 ;
  assign y5993 = n20068 ;
  assign y5994 = ~n20072 ;
  assign y5995 = n20074 ;
  assign y5996 = n20076 ;
  assign y5997 = n20078 ;
  assign y5998 = n20080 ;
  assign y5999 = n20081 ;
  assign y6000 = n20086 ;
  assign y6001 = ~n20094 ;
  assign y6002 = n20098 ;
  assign y6003 = ~n20105 ;
  assign y6004 = ~n20107 ;
  assign y6005 = n20110 ;
  assign y6006 = ~1'b0 ;
  assign y6007 = ~1'b0 ;
  assign y6008 = ~n20117 ;
  assign y6009 = ~n20118 ;
  assign y6010 = ~n20125 ;
  assign y6011 = n20133 ;
  assign y6012 = ~n20138 ;
  assign y6013 = n20145 ;
  assign y6014 = ~n20146 ;
  assign y6015 = ~n20152 ;
  assign y6016 = ~n20154 ;
  assign y6017 = ~n20158 ;
  assign y6018 = ~n20171 ;
  assign y6019 = n20172 ;
  assign y6020 = ~n20176 ;
  assign y6021 = n20177 ;
  assign y6022 = ~n20178 ;
  assign y6023 = ~1'b0 ;
  assign y6024 = n20179 ;
  assign y6025 = n20184 ;
  assign y6026 = n20187 ;
  assign y6027 = ~n20193 ;
  assign y6028 = ~1'b0 ;
  assign y6029 = ~n20194 ;
  assign y6030 = n20195 ;
  assign y6031 = n20199 ;
  assign y6032 = ~1'b0 ;
  assign y6033 = ~1'b0 ;
  assign y6034 = n20201 ;
  assign y6035 = ~n20205 ;
  assign y6036 = n20216 ;
  assign y6037 = n20220 ;
  assign y6038 = ~n20222 ;
  assign y6039 = n20224 ;
  assign y6040 = ~n20228 ;
  assign y6041 = ~n20234 ;
  assign y6042 = n20236 ;
  assign y6043 = n20242 ;
  assign y6044 = ~1'b0 ;
  assign y6045 = ~1'b0 ;
  assign y6046 = ~1'b0 ;
  assign y6047 = ~n20244 ;
  assign y6048 = ~n20246 ;
  assign y6049 = n20256 ;
  assign y6050 = ~n20257 ;
  assign y6051 = n20259 ;
  assign y6052 = ~n20264 ;
  assign y6053 = n20267 ;
  assign y6054 = n20271 ;
  assign y6055 = n20272 ;
  assign y6056 = n20275 ;
  assign y6057 = ~n20278 ;
  assign y6058 = ~1'b0 ;
  assign y6059 = n20280 ;
  assign y6060 = ~n20285 ;
  assign y6061 = ~n20289 ;
  assign y6062 = ~n20290 ;
  assign y6063 = ~n20294 ;
  assign y6064 = n20299 ;
  assign y6065 = ~1'b0 ;
  assign y6066 = ~n20300 ;
  assign y6067 = n20301 ;
  assign y6068 = ~n20303 ;
  assign y6069 = ~n20306 ;
  assign y6070 = ~n20310 ;
  assign y6071 = n20312 ;
  assign y6072 = n20315 ;
  assign y6073 = ~n20318 ;
  assign y6074 = n20323 ;
  assign y6075 = ~n20328 ;
  assign y6076 = ~n20329 ;
  assign y6077 = ~n20330 ;
  assign y6078 = ~n20331 ;
  assign y6079 = ~n20334 ;
  assign y6080 = n20336 ;
  assign y6081 = n20337 ;
  assign y6082 = ~n20340 ;
  assign y6083 = n20341 ;
  assign y6084 = ~n20343 ;
  assign y6085 = n20347 ;
  assign y6086 = ~1'b0 ;
  assign y6087 = n20350 ;
  assign y6088 = n20351 ;
  assign y6089 = n20352 ;
  assign y6090 = 1'b0 ;
  assign y6091 = ~1'b0 ;
  assign y6092 = ~1'b0 ;
  assign y6093 = ~n20362 ;
  assign y6094 = n20363 ;
  assign y6095 = n20364 ;
  assign y6096 = 1'b0 ;
  assign y6097 = n20373 ;
  assign y6098 = ~n20379 ;
  assign y6099 = n20383 ;
  assign y6100 = ~n20385 ;
  assign y6101 = ~n20390 ;
  assign y6102 = n20391 ;
  assign y6103 = ~1'b0 ;
  assign y6104 = ~1'b0 ;
  assign y6105 = ~n20396 ;
  assign y6106 = n20398 ;
  assign y6107 = ~n7356 ;
  assign y6108 = ~1'b0 ;
  assign y6109 = n20399 ;
  assign y6110 = ~n20403 ;
  assign y6111 = ~n20404 ;
  assign y6112 = ~n20405 ;
  assign y6113 = ~n20409 ;
  assign y6114 = n20410 ;
  assign y6115 = ~n20413 ;
  assign y6116 = ~n20417 ;
  assign y6117 = n20420 ;
  assign y6118 = n20426 ;
  assign y6119 = ~n20430 ;
  assign y6120 = n20431 ;
  assign y6121 = ~n20437 ;
  assign y6122 = ~n20439 ;
  assign y6123 = n20441 ;
  assign y6124 = n20444 ;
  assign y6125 = n20450 ;
  assign y6126 = ~n20453 ;
  assign y6127 = ~n20455 ;
  assign y6128 = ~n20463 ;
  assign y6129 = ~n20467 ;
  assign y6130 = n20468 ;
  assign y6131 = ~n20473 ;
  assign y6132 = ~n20476 ;
  assign y6133 = ~n20479 ;
  assign y6134 = ~1'b0 ;
  assign y6135 = n20481 ;
  assign y6136 = ~n20487 ;
  assign y6137 = n20492 ;
  assign y6138 = ~n20493 ;
  assign y6139 = n20498 ;
  assign y6140 = ~1'b0 ;
  assign y6141 = ~1'b0 ;
  assign y6142 = n20504 ;
  assign y6143 = ~n20514 ;
  assign y6144 = ~n20521 ;
  assign y6145 = ~n20522 ;
  assign y6146 = ~n20524 ;
  assign y6147 = ~1'b0 ;
  assign y6148 = n20527 ;
  assign y6149 = n20529 ;
  assign y6150 = ~n20530 ;
  assign y6151 = n20533 ;
  assign y6152 = ~n20541 ;
  assign y6153 = n20545 ;
  assign y6154 = ~1'b0 ;
  assign y6155 = ~n20550 ;
  assign y6156 = ~1'b0 ;
  assign y6157 = ~n20553 ;
  assign y6158 = ~1'b0 ;
  assign y6159 = n20563 ;
  assign y6160 = ~n20565 ;
  assign y6161 = n20566 ;
  assign y6162 = n20569 ;
  assign y6163 = ~1'b0 ;
  assign y6164 = ~n20571 ;
  assign y6165 = ~n20578 ;
  assign y6166 = ~n20579 ;
  assign y6167 = ~n20580 ;
  assign y6168 = ~n20587 ;
  assign y6169 = ~n20590 ;
  assign y6170 = n20591 ;
  assign y6171 = ~n20593 ;
  assign y6172 = n20595 ;
  assign y6173 = n20608 ;
  assign y6174 = ~1'b0 ;
  assign y6175 = n20616 ;
  assign y6176 = ~n20618 ;
  assign y6177 = n20630 ;
  assign y6178 = n20631 ;
  assign y6179 = n20633 ;
  assign y6180 = 1'b0 ;
  assign y6181 = n20635 ;
  assign y6182 = ~1'b0 ;
  assign y6183 = ~1'b0 ;
  assign y6184 = ~n20638 ;
  assign y6185 = n20639 ;
  assign y6186 = ~n20640 ;
  assign y6187 = ~n20642 ;
  assign y6188 = ~n20643 ;
  assign y6189 = ~n20654 ;
  assign y6190 = ~1'b0 ;
  assign y6191 = n20656 ;
  assign y6192 = n20657 ;
  assign y6193 = ~n20658 ;
  assign y6194 = n13551 ;
  assign y6195 = n20662 ;
  assign y6196 = ~n20666 ;
  assign y6197 = ~1'b0 ;
  assign y6198 = ~n20668 ;
  assign y6199 = ~n20675 ;
  assign y6200 = n20682 ;
  assign y6201 = ~n20683 ;
  assign y6202 = ~n20684 ;
  assign y6203 = ~n20691 ;
  assign y6204 = ~n20694 ;
  assign y6205 = ~n20696 ;
  assign y6206 = ~n20697 ;
  assign y6207 = n20698 ;
  assign y6208 = n20699 ;
  assign y6209 = ~1'b0 ;
  assign y6210 = ~n20704 ;
  assign y6211 = n20706 ;
  assign y6212 = n8282 ;
  assign y6213 = n20708 ;
  assign y6214 = ~n20715 ;
  assign y6215 = ~n20718 ;
  assign y6216 = ~n20720 ;
  assign y6217 = ~1'b0 ;
  assign y6218 = ~1'b0 ;
  assign y6219 = ~n20721 ;
  assign y6220 = n20723 ;
  assign y6221 = n20726 ;
  assign y6222 = ~n20732 ;
  assign y6223 = ~n20740 ;
  assign y6224 = ~n20741 ;
  assign y6225 = ~n20746 ;
  assign y6226 = ~n20747 ;
  assign y6227 = n20753 ;
  assign y6228 = n20765 ;
  assign y6229 = ~n20769 ;
  assign y6230 = ~n20771 ;
  assign y6231 = ~n20772 ;
  assign y6232 = ~n20773 ;
  assign y6233 = n20778 ;
  assign y6234 = ~1'b0 ;
  assign y6235 = n20780 ;
  assign y6236 = ~n20786 ;
  assign y6237 = ~n20792 ;
  assign y6238 = n20799 ;
  assign y6239 = ~1'b0 ;
  assign y6240 = ~n20804 ;
  assign y6241 = n20805 ;
  assign y6242 = ~1'b0 ;
  assign y6243 = n20808 ;
  assign y6244 = n20812 ;
  assign y6245 = n20815 ;
  assign y6246 = n20819 ;
  assign y6247 = n20822 ;
  assign y6248 = ~n20824 ;
  assign y6249 = ~n20826 ;
  assign y6250 = n20827 ;
  assign y6251 = ~n20828 ;
  assign y6252 = ~n20831 ;
  assign y6253 = n20835 ;
  assign y6254 = ~n20837 ;
  assign y6255 = ~1'b0 ;
  assign y6256 = ~1'b0 ;
  assign y6257 = n20838 ;
  assign y6258 = ~n20845 ;
  assign y6259 = ~n20847 ;
  assign y6260 = n20849 ;
  assign y6261 = n20850 ;
  assign y6262 = ~n20856 ;
  assign y6263 = ~n8873 ;
  assign y6264 = ~n8503 ;
  assign y6265 = n20857 ;
  assign y6266 = n20860 ;
  assign y6267 = n20865 ;
  assign y6268 = ~n20869 ;
  assign y6269 = ~n20875 ;
  assign y6270 = ~1'b0 ;
  assign y6271 = ~n20876 ;
  assign y6272 = ~n20882 ;
  assign y6273 = ~n20884 ;
  assign y6274 = ~n20885 ;
  assign y6275 = ~1'b0 ;
  assign y6276 = n20889 ;
  assign y6277 = ~n20893 ;
  assign y6278 = ~1'b0 ;
  assign y6279 = ~1'b0 ;
  assign y6280 = ~n20895 ;
  assign y6281 = ~n20898 ;
  assign y6282 = ~1'b0 ;
  assign y6283 = n20904 ;
  assign y6284 = ~n20907 ;
  assign y6285 = n20910 ;
  assign y6286 = ~n20912 ;
  assign y6287 = ~n20913 ;
  assign y6288 = ~n20917 ;
  assign y6289 = n20920 ;
  assign y6290 = ~n20922 ;
  assign y6291 = ~n20927 ;
  assign y6292 = n20930 ;
  assign y6293 = n20932 ;
  assign y6294 = ~n20935 ;
  assign y6295 = n20936 ;
  assign y6296 = ~n20938 ;
  assign y6297 = n20939 ;
  assign y6298 = ~n20944 ;
  assign y6299 = n20949 ;
  assign y6300 = ~n20953 ;
  assign y6301 = ~n20954 ;
  assign y6302 = ~n20956 ;
  assign y6303 = ~n20957 ;
  assign y6304 = ~n20959 ;
  assign y6305 = ~n20961 ;
  assign y6306 = n6160 ;
  assign y6307 = ~n20962 ;
  assign y6308 = n20963 ;
  assign y6309 = ~n20965 ;
  assign y6310 = ~1'b0 ;
  assign y6311 = ~n20969 ;
  assign y6312 = ~n20974 ;
  assign y6313 = n20978 ;
  assign y6314 = ~n20979 ;
  assign y6315 = n20980 ;
  assign y6316 = ~n20981 ;
  assign y6317 = ~1'b0 ;
  assign y6318 = n20983 ;
  assign y6319 = n20984 ;
  assign y6320 = n20986 ;
  assign y6321 = n20992 ;
  assign y6322 = ~1'b0 ;
  assign y6323 = n20995 ;
  assign y6324 = ~1'b0 ;
  assign y6325 = n20997 ;
  assign y6326 = n21003 ;
  assign y6327 = ~n21004 ;
  assign y6328 = n21005 ;
  assign y6329 = n21009 ;
  assign y6330 = n21013 ;
  assign y6331 = n21014 ;
  assign y6332 = n21025 ;
  assign y6333 = ~1'b0 ;
  assign y6334 = n21028 ;
  assign y6335 = n21030 ;
  assign y6336 = n21036 ;
  assign y6337 = n21038 ;
  assign y6338 = ~n3312 ;
  assign y6339 = n21041 ;
  assign y6340 = ~n21044 ;
  assign y6341 = ~1'b0 ;
  assign y6342 = n21049 ;
  assign y6343 = n21050 ;
  assign y6344 = n21054 ;
  assign y6345 = n21055 ;
  assign y6346 = n21056 ;
  assign y6347 = n21058 ;
  assign y6348 = ~1'b0 ;
  assign y6349 = ~1'b0 ;
  assign y6350 = ~1'b0 ;
  assign y6351 = n21064 ;
  assign y6352 = ~n15480 ;
  assign y6353 = ~n21066 ;
  assign y6354 = ~n21072 ;
  assign y6355 = n21076 ;
  assign y6356 = ~n21081 ;
  assign y6357 = n11004 ;
  assign y6358 = n21083 ;
  assign y6359 = ~n21087 ;
  assign y6360 = n21089 ;
  assign y6361 = ~n21091 ;
  assign y6362 = ~n21101 ;
  assign y6363 = ~n21110 ;
  assign y6364 = n21111 ;
  assign y6365 = ~n21112 ;
  assign y6366 = ~n21114 ;
  assign y6367 = n21116 ;
  assign y6368 = ~n21117 ;
  assign y6369 = n21118 ;
  assign y6370 = n21122 ;
  assign y6371 = n21126 ;
  assign y6372 = ~n21130 ;
  assign y6373 = ~1'b0 ;
  assign y6374 = n21132 ;
  assign y6375 = ~n21135 ;
  assign y6376 = n21136 ;
  assign y6377 = n21137 ;
  assign y6378 = n21138 ;
  assign y6379 = ~n21141 ;
  assign y6380 = n21146 ;
  assign y6381 = ~n21151 ;
  assign y6382 = ~n21153 ;
  assign y6383 = ~n21154 ;
  assign y6384 = n21160 ;
  assign y6385 = n21161 ;
  assign y6386 = ~1'b0 ;
  assign y6387 = n21162 ;
  assign y6388 = ~n21166 ;
  assign y6389 = n21168 ;
  assign y6390 = ~1'b0 ;
  assign y6391 = ~n21172 ;
  assign y6392 = ~n21173 ;
  assign y6393 = ~n21177 ;
  assign y6394 = ~n21180 ;
  assign y6395 = n21182 ;
  assign y6396 = n21188 ;
  assign y6397 = ~n21189 ;
  assign y6398 = ~n21191 ;
  assign y6399 = n21193 ;
  assign y6400 = n21197 ;
  assign y6401 = ~n21203 ;
  assign y6402 = ~n21206 ;
  assign y6403 = ~1'b0 ;
  assign y6404 = n21209 ;
  assign y6405 = n21214 ;
  assign y6406 = ~n21216 ;
  assign y6407 = ~n21218 ;
  assign y6408 = n21234 ;
  assign y6409 = n21235 ;
  assign y6410 = ~n21236 ;
  assign y6411 = ~n21237 ;
  assign y6412 = ~n21238 ;
  assign y6413 = n21240 ;
  assign y6414 = ~n21242 ;
  assign y6415 = ~1'b0 ;
  assign y6416 = ~n21244 ;
  assign y6417 = n21248 ;
  assign y6418 = ~n21251 ;
  assign y6419 = ~n21252 ;
  assign y6420 = ~n21256 ;
  assign y6421 = n21257 ;
  assign y6422 = ~1'b0 ;
  assign y6423 = n21263 ;
  assign y6424 = n21264 ;
  assign y6425 = n21265 ;
  assign y6426 = ~n21271 ;
  assign y6427 = ~1'b0 ;
  assign y6428 = n21277 ;
  assign y6429 = ~n21279 ;
  assign y6430 = n21280 ;
  assign y6431 = n21281 ;
  assign y6432 = n21282 ;
  assign y6433 = n21284 ;
  assign y6434 = ~1'b0 ;
  assign y6435 = n21293 ;
  assign y6436 = n21295 ;
  assign y6437 = ~n21296 ;
  assign y6438 = ~n21302 ;
  assign y6439 = n21307 ;
  assign y6440 = ~1'b0 ;
  assign y6441 = ~1'b0 ;
  assign y6442 = n21310 ;
  assign y6443 = ~n21315 ;
  assign y6444 = ~n21317 ;
  assign y6445 = ~n21318 ;
  assign y6446 = n21319 ;
  assign y6447 = n21320 ;
  assign y6448 = ~n21322 ;
  assign y6449 = ~n21323 ;
  assign y6450 = ~1'b0 ;
  assign y6451 = n21325 ;
  assign y6452 = ~n21326 ;
  assign y6453 = n21327 ;
  assign y6454 = ~n21333 ;
  assign y6455 = ~1'b0 ;
  assign y6456 = n21336 ;
  assign y6457 = ~n21338 ;
  assign y6458 = ~n21345 ;
  assign y6459 = ~n21350 ;
  assign y6460 = n21353 ;
  assign y6461 = ~n21355 ;
  assign y6462 = ~n21358 ;
  assign y6463 = ~n21362 ;
  assign y6464 = n21370 ;
  assign y6465 = ~n21374 ;
  assign y6466 = ~n21375 ;
  assign y6467 = ~n21380 ;
  assign y6468 = ~n21381 ;
  assign y6469 = n21386 ;
  assign y6470 = ~n21391 ;
  assign y6471 = ~1'b0 ;
  assign y6472 = ~n21396 ;
  assign y6473 = n21401 ;
  assign y6474 = ~n21402 ;
  assign y6475 = ~n21404 ;
  assign y6476 = ~1'b0 ;
  assign y6477 = ~n21408 ;
  assign y6478 = ~n21413 ;
  assign y6479 = n21415 ;
  assign y6480 = ~1'b0 ;
  assign y6481 = ~n21420 ;
  assign y6482 = ~n21423 ;
  assign y6483 = ~n21425 ;
  assign y6484 = ~n21426 ;
  assign y6485 = ~1'b0 ;
  assign y6486 = ~n21428 ;
  assign y6487 = n21429 ;
  assign y6488 = ~n21431 ;
  assign y6489 = ~n21432 ;
  assign y6490 = n21433 ;
  assign y6491 = n21438 ;
  assign y6492 = ~n21440 ;
  assign y6493 = ~n21448 ;
  assign y6494 = n21449 ;
  assign y6495 = ~n21452 ;
  assign y6496 = n21455 ;
  assign y6497 = n21456 ;
  assign y6498 = ~n21459 ;
  assign y6499 = ~n21467 ;
  assign y6500 = ~n21469 ;
  assign y6501 = ~n21470 ;
  assign y6502 = ~n21473 ;
  assign y6503 = ~n15379 ;
  assign y6504 = ~n21476 ;
  assign y6505 = n21478 ;
  assign y6506 = ~n21479 ;
  assign y6507 = n21480 ;
  assign y6508 = ~n21482 ;
  assign y6509 = n21483 ;
  assign y6510 = n21486 ;
  assign y6511 = n21488 ;
  assign y6512 = ~n21490 ;
  assign y6513 = ~n21491 ;
  assign y6514 = ~1'b0 ;
  assign y6515 = ~1'b0 ;
  assign y6516 = n21494 ;
  assign y6517 = n21501 ;
  assign y6518 = n21505 ;
  assign y6519 = ~n21508 ;
  assign y6520 = ~n21512 ;
  assign y6521 = ~n21516 ;
  assign y6522 = ~n21517 ;
  assign y6523 = ~n21520 ;
  assign y6524 = n21523 ;
  assign y6525 = ~1'b0 ;
  assign y6526 = ~n21524 ;
  assign y6527 = n21527 ;
  assign y6528 = ~n21528 ;
  assign y6529 = ~n21530 ;
  assign y6530 = n21535 ;
  assign y6531 = ~n21538 ;
  assign y6532 = n21539 ;
  assign y6533 = ~n21541 ;
  assign y6534 = n21546 ;
  assign y6535 = ~n21547 ;
  assign y6536 = n21548 ;
  assign y6537 = ~1'b0 ;
  assign y6538 = n21551 ;
  assign y6539 = ~1'b0 ;
  assign y6540 = ~n21553 ;
  assign y6541 = n21554 ;
  assign y6542 = ~n21555 ;
  assign y6543 = ~n21556 ;
  assign y6544 = ~n21562 ;
  assign y6545 = ~1'b0 ;
  assign y6546 = ~1'b0 ;
  assign y6547 = ~n16679 ;
  assign y6548 = ~n21564 ;
  assign y6549 = n21569 ;
  assign y6550 = ~n21571 ;
  assign y6551 = ~n21576 ;
  assign y6552 = ~1'b0 ;
  assign y6553 = n21582 ;
  assign y6554 = ~1'b0 ;
  assign y6555 = n21583 ;
  assign y6556 = ~n21585 ;
  assign y6557 = n21586 ;
  assign y6558 = ~1'b0 ;
  assign y6559 = n21588 ;
  assign y6560 = n21589 ;
  assign y6561 = n21590 ;
  assign y6562 = ~n21594 ;
  assign y6563 = ~n21598 ;
  assign y6564 = x84 ;
  assign y6565 = ~n21601 ;
  assign y6566 = ~1'b0 ;
  assign y6567 = n21602 ;
  assign y6568 = n21604 ;
  assign y6569 = ~n21605 ;
  assign y6570 = ~n21607 ;
  assign y6571 = ~1'b0 ;
  assign y6572 = ~1'b0 ;
  assign y6573 = ~n21613 ;
  assign y6574 = ~n21614 ;
  assign y6575 = ~n21617 ;
  assign y6576 = ~n21618 ;
  assign y6577 = ~n21619 ;
  assign y6578 = ~n21623 ;
  assign y6579 = ~1'b0 ;
  assign y6580 = n21625 ;
  assign y6581 = n21627 ;
  assign y6582 = ~n21628 ;
  assign y6583 = n21629 ;
  assign y6584 = n21631 ;
  assign y6585 = n21632 ;
  assign y6586 = ~n21635 ;
  assign y6587 = ~1'b0 ;
  assign y6588 = n21641 ;
  assign y6589 = n21644 ;
  assign y6590 = ~1'b0 ;
  assign y6591 = ~n21645 ;
  assign y6592 = n21649 ;
  assign y6593 = n21650 ;
  assign y6594 = ~n21652 ;
  assign y6595 = ~1'b0 ;
  assign y6596 = ~n21655 ;
  assign y6597 = ~1'b0 ;
  assign y6598 = ~n21656 ;
  assign y6599 = ~n21657 ;
  assign y6600 = n21659 ;
  assign y6601 = ~n21665 ;
  assign y6602 = n21668 ;
  assign y6603 = ~1'b0 ;
  assign y6604 = n21669 ;
  assign y6605 = n21670 ;
  assign y6606 = ~1'b0 ;
  assign y6607 = n21672 ;
  assign y6608 = ~1'b0 ;
  assign y6609 = ~1'b0 ;
  assign y6610 = ~n21674 ;
  assign y6611 = ~n21678 ;
  assign y6612 = n21679 ;
  assign y6613 = n21680 ;
  assign y6614 = ~n21681 ;
  assign y6615 = ~1'b0 ;
  assign y6616 = n21682 ;
  assign y6617 = ~n21683 ;
  assign y6618 = n21690 ;
  assign y6619 = ~n21693 ;
  assign y6620 = n21701 ;
  assign y6621 = ~n21704 ;
  assign y6622 = ~n21710 ;
  assign y6623 = ~n21713 ;
  assign y6624 = n21714 ;
  assign y6625 = n21720 ;
  assign y6626 = n21727 ;
  assign y6627 = n21729 ;
  assign y6628 = n21731 ;
  assign y6629 = n7154 ;
  assign y6630 = n21738 ;
  assign y6631 = ~1'b0 ;
  assign y6632 = ~n21739 ;
  assign y6633 = ~n21741 ;
  assign y6634 = ~n21746 ;
  assign y6635 = n21754 ;
  assign y6636 = n21757 ;
  assign y6637 = ~n21760 ;
  assign y6638 = n21763 ;
  assign y6639 = ~n21765 ;
  assign y6640 = ~n21767 ;
  assign y6641 = n21770 ;
  assign y6642 = ~n21778 ;
  assign y6643 = ~n21780 ;
  assign y6644 = ~n21782 ;
  assign y6645 = n21783 ;
  assign y6646 = ~n4576 ;
  assign y6647 = ~1'b0 ;
  assign y6648 = n21784 ;
  assign y6649 = ~n21788 ;
  assign y6650 = n21789 ;
  assign y6651 = n21790 ;
  assign y6652 = ~1'b0 ;
  assign y6653 = ~n21792 ;
  assign y6654 = n21794 ;
  assign y6655 = ~n21799 ;
  assign y6656 = ~1'b0 ;
  assign y6657 = ~1'b0 ;
  assign y6658 = ~1'b0 ;
  assign y6659 = ~n21800 ;
  assign y6660 = n21805 ;
  assign y6661 = n21806 ;
  assign y6662 = n21809 ;
  assign y6663 = ~1'b0 ;
  assign y6664 = ~1'b0 ;
  assign y6665 = ~n21812 ;
  assign y6666 = ~1'b0 ;
  assign y6667 = ~n21813 ;
  assign y6668 = ~n21818 ;
  assign y6669 = ~n21820 ;
  assign y6670 = n21822 ;
  assign y6671 = n21823 ;
  assign y6672 = n21825 ;
  assign y6673 = ~n21827 ;
  assign y6674 = n21828 ;
  assign y6675 = ~n21830 ;
  assign y6676 = ~n21831 ;
  assign y6677 = n21841 ;
  assign y6678 = ~n21843 ;
  assign y6679 = n21844 ;
  assign y6680 = ~n21845 ;
  assign y6681 = ~n21846 ;
  assign y6682 = ~n21847 ;
  assign y6683 = ~n21852 ;
  assign y6684 = ~n21855 ;
  assign y6685 = n21859 ;
  assign y6686 = ~n21861 ;
  assign y6687 = ~n21862 ;
  assign y6688 = ~n21865 ;
  assign y6689 = n21868 ;
  assign y6690 = ~n21869 ;
  assign y6691 = ~n21875 ;
  assign y6692 = ~1'b0 ;
  assign y6693 = n21876 ;
  assign y6694 = ~n21883 ;
  assign y6695 = ~n21885 ;
  assign y6696 = ~n21888 ;
  assign y6697 = ~n21889 ;
  assign y6698 = n21894 ;
  assign y6699 = n21896 ;
  assign y6700 = ~n21898 ;
  assign y6701 = ~n21900 ;
  assign y6702 = n21902 ;
  assign y6703 = ~n21905 ;
  assign y6704 = n21909 ;
  assign y6705 = ~1'b0 ;
  assign y6706 = ~n21910 ;
  assign y6707 = n21911 ;
  assign y6708 = ~n21917 ;
  assign y6709 = n21918 ;
  assign y6710 = ~n21922 ;
  assign y6711 = ~1'b0 ;
  assign y6712 = ~n21924 ;
  assign y6713 = ~n21926 ;
  assign y6714 = n21928 ;
  assign y6715 = ~n21929 ;
  assign y6716 = ~n21931 ;
  assign y6717 = ~n21932 ;
  assign y6718 = n21933 ;
  assign y6719 = ~n21934 ;
  assign y6720 = ~n21938 ;
  assign y6721 = ~1'b0 ;
  assign y6722 = n21941 ;
  assign y6723 = n21942 ;
  assign y6724 = n21944 ;
  assign y6725 = ~n21949 ;
  assign y6726 = n21951 ;
  assign y6727 = ~1'b0 ;
  assign y6728 = ~1'b0 ;
  assign y6729 = ~n21954 ;
  assign y6730 = n21959 ;
  assign y6731 = ~n21961 ;
  assign y6732 = n21965 ;
  assign y6733 = n21969 ;
  assign y6734 = ~n21972 ;
  assign y6735 = n21977 ;
  assign y6736 = ~n21979 ;
  assign y6737 = ~n21981 ;
  assign y6738 = ~n21984 ;
  assign y6739 = ~n21987 ;
  assign y6740 = ~n21990 ;
  assign y6741 = ~n21991 ;
  assign y6742 = n21995 ;
  assign y6743 = ~1'b0 ;
  assign y6744 = ~n21996 ;
  assign y6745 = ~1'b0 ;
  assign y6746 = n21999 ;
  assign y6747 = ~n22002 ;
  assign y6748 = n22003 ;
  assign y6749 = ~n22007 ;
  assign y6750 = n22008 ;
  assign y6751 = ~1'b0 ;
  assign y6752 = ~n22011 ;
  assign y6753 = n22014 ;
  assign y6754 = n22016 ;
  assign y6755 = ~n22019 ;
  assign y6756 = ~1'b0 ;
  assign y6757 = ~n22021 ;
  assign y6758 = ~n22026 ;
  assign y6759 = ~n22027 ;
  assign y6760 = n22028 ;
  assign y6761 = ~n22029 ;
  assign y6762 = n22032 ;
  assign y6763 = ~1'b0 ;
  assign y6764 = n22034 ;
  assign y6765 = n22035 ;
  assign y6766 = ~n22038 ;
  assign y6767 = n22040 ;
  assign y6768 = n22042 ;
  assign y6769 = ~n22044 ;
  assign y6770 = ~n22046 ;
  assign y6771 = n22048 ;
  assign y6772 = n22050 ;
  assign y6773 = ~n22051 ;
  assign y6774 = ~1'b0 ;
  assign y6775 = ~n22052 ;
  assign y6776 = ~n22063 ;
  assign y6777 = n22066 ;
  assign y6778 = ~n22068 ;
  assign y6779 = n22071 ;
  assign y6780 = n22072 ;
  assign y6781 = ~n22073 ;
  assign y6782 = ~1'b0 ;
  assign y6783 = ~n22082 ;
  assign y6784 = ~n22085 ;
  assign y6785 = n22086 ;
  assign y6786 = n22087 ;
  assign y6787 = ~n22088 ;
  assign y6788 = ~n22094 ;
  assign y6789 = ~1'b0 ;
  assign y6790 = ~n22096 ;
  assign y6791 = ~n22097 ;
  assign y6792 = ~n22100 ;
  assign y6793 = n22102 ;
  assign y6794 = n22103 ;
  assign y6795 = n22104 ;
  assign y6796 = n22109 ;
  assign y6797 = ~n22112 ;
  assign y6798 = n22113 ;
  assign y6799 = ~n22121 ;
  assign y6800 = n22127 ;
  assign y6801 = n22128 ;
  assign y6802 = ~n22131 ;
  assign y6803 = ~n22137 ;
  assign y6804 = ~1'b0 ;
  assign y6805 = n22139 ;
  assign y6806 = ~1'b0 ;
  assign y6807 = ~n12927 ;
  assign y6808 = ~n22140 ;
  assign y6809 = ~n22144 ;
  assign y6810 = ~n22149 ;
  assign y6811 = ~n22151 ;
  assign y6812 = ~n22153 ;
  assign y6813 = ~n22155 ;
  assign y6814 = ~n22160 ;
  assign y6815 = ~n22163 ;
  assign y6816 = ~n22166 ;
  assign y6817 = n22167 ;
  assign y6818 = n22169 ;
  assign y6819 = n22172 ;
  assign y6820 = ~n22174 ;
  assign y6821 = n9908 ;
  assign y6822 = ~n568 ;
  assign y6823 = n22175 ;
  assign y6824 = ~1'b0 ;
  assign y6825 = n22180 ;
  assign y6826 = ~n22192 ;
  assign y6827 = ~n22195 ;
  assign y6828 = n22197 ;
  assign y6829 = ~n22199 ;
  assign y6830 = ~n22200 ;
  assign y6831 = ~n22202 ;
  assign y6832 = n22204 ;
  assign y6833 = ~1'b0 ;
  assign y6834 = ~n22205 ;
  assign y6835 = ~n22212 ;
  assign y6836 = n22215 ;
  assign y6837 = n22216 ;
  assign y6838 = ~n22219 ;
  assign y6839 = ~n22220 ;
  assign y6840 = ~n22223 ;
  assign y6841 = n22225 ;
  assign y6842 = n22227 ;
  assign y6843 = ~n22228 ;
  assign y6844 = n22229 ;
  assign y6845 = ~n22231 ;
  assign y6846 = n22237 ;
  assign y6847 = n22241 ;
  assign y6848 = ~1'b0 ;
  assign y6849 = ~n22243 ;
  assign y6850 = n22252 ;
  assign y6851 = ~n22254 ;
  assign y6852 = n22257 ;
  assign y6853 = n22260 ;
  assign y6854 = n22262 ;
  assign y6855 = n22263 ;
  assign y6856 = n22269 ;
  assign y6857 = ~n22272 ;
  assign y6858 = n22274 ;
  assign y6859 = ~n22276 ;
  assign y6860 = n22279 ;
  assign y6861 = ~n22288 ;
  assign y6862 = ~n22290 ;
  assign y6863 = n22293 ;
  assign y6864 = ~n22297 ;
  assign y6865 = ~n22303 ;
  assign y6866 = ~1'b0 ;
  assign y6867 = n22304 ;
  assign y6868 = ~1'b0 ;
  assign y6869 = n22307 ;
  assign y6870 = n22308 ;
  assign y6871 = ~n22311 ;
  assign y6872 = ~n22313 ;
  assign y6873 = ~n22314 ;
  assign y6874 = n222 ;
  assign y6875 = n22316 ;
  assign y6876 = ~n22321 ;
  assign y6877 = ~n22322 ;
  assign y6878 = ~n22329 ;
  assign y6879 = ~n22333 ;
  assign y6880 = ~1'b0 ;
  assign y6881 = n22337 ;
  assign y6882 = n22339 ;
  assign y6883 = ~n22346 ;
  assign y6884 = n22351 ;
  assign y6885 = ~n22356 ;
  assign y6886 = ~n22358 ;
  assign y6887 = n22360 ;
  assign y6888 = ~1'b0 ;
  assign y6889 = ~n22362 ;
  assign y6890 = ~n22370 ;
  assign y6891 = ~n22374 ;
  assign y6892 = ~n22379 ;
  assign y6893 = ~1'b0 ;
  assign y6894 = n22381 ;
  assign y6895 = ~n22385 ;
  assign y6896 = n22388 ;
  assign y6897 = ~n22390 ;
  assign y6898 = ~n22392 ;
  assign y6899 = ~n22393 ;
  assign y6900 = ~n22397 ;
  assign y6901 = ~1'b0 ;
  assign y6902 = n22398 ;
  assign y6903 = ~1'b0 ;
  assign y6904 = ~n22400 ;
  assign y6905 = ~n22406 ;
  assign y6906 = ~n22407 ;
  assign y6907 = n22411 ;
  assign y6908 = n22412 ;
  assign y6909 = ~n22414 ;
  assign y6910 = n22416 ;
  assign y6911 = ~n22418 ;
  assign y6912 = ~n22420 ;
  assign y6913 = ~n22426 ;
  assign y6914 = n22430 ;
  assign y6915 = ~n22431 ;
  assign y6916 = n22435 ;
  assign y6917 = n22439 ;
  assign y6918 = n22446 ;
  assign y6919 = ~n22450 ;
  assign y6920 = n22453 ;
  assign y6921 = ~n22455 ;
  assign y6922 = ~n22456 ;
  assign y6923 = n22462 ;
  assign y6924 = ~n22463 ;
  assign y6925 = ~n22465 ;
  assign y6926 = ~1'b0 ;
  assign y6927 = ~n22470 ;
  assign y6928 = n22471 ;
  assign y6929 = ~n22476 ;
  assign y6930 = ~n22481 ;
  assign y6931 = ~n22483 ;
  assign y6932 = n22490 ;
  assign y6933 = ~1'b0 ;
  assign y6934 = ~n22493 ;
  assign y6935 = n22496 ;
  assign y6936 = ~1'b0 ;
  assign y6937 = ~n22497 ;
  assign y6938 = ~n22499 ;
  assign y6939 = n22502 ;
  assign y6940 = n22504 ;
  assign y6941 = ~1'b0 ;
  assign y6942 = n18723 ;
  assign y6943 = ~n22508 ;
  assign y6944 = ~n22511 ;
  assign y6945 = 1'b0 ;
  assign y6946 = ~1'b0 ;
  assign y6947 = ~1'b0 ;
  assign y6948 = n22513 ;
  assign y6949 = ~n22515 ;
  assign y6950 = ~n22521 ;
  assign y6951 = n22525 ;
  assign y6952 = n22527 ;
  assign y6953 = n22530 ;
  assign y6954 = n22531 ;
  assign y6955 = n22537 ;
  assign y6956 = ~1'b0 ;
  assign y6957 = ~n22539 ;
  assign y6958 = ~1'b0 ;
  assign y6959 = n22543 ;
  assign y6960 = n22545 ;
  assign y6961 = ~n22548 ;
  assign y6962 = n22549 ;
  assign y6963 = ~n22557 ;
  assign y6964 = ~n22563 ;
  assign y6965 = n22565 ;
  assign y6966 = ~n22566 ;
  assign y6967 = ~n22567 ;
  assign y6968 = n21321 ;
  assign y6969 = ~n22568 ;
  assign y6970 = ~n22570 ;
  assign y6971 = n22575 ;
  assign y6972 = n22581 ;
  assign y6973 = n22583 ;
  assign y6974 = n22584 ;
  assign y6975 = n22589 ;
  assign y6976 = ~n22590 ;
  assign y6977 = n22598 ;
  assign y6978 = ~1'b0 ;
  assign y6979 = n22601 ;
  assign y6980 = n22607 ;
  assign y6981 = ~n22609 ;
  assign y6982 = ~n22612 ;
  assign y6983 = n22613 ;
  assign y6984 = n22615 ;
  assign y6985 = n22618 ;
  assign y6986 = ~n22620 ;
  assign y6987 = ~n22623 ;
  assign y6988 = ~n22625 ;
  assign y6989 = ~n22627 ;
  assign y6990 = ~n22630 ;
  assign y6991 = ~n22633 ;
  assign y6992 = ~n22635 ;
  assign y6993 = ~n22642 ;
  assign y6994 = n22654 ;
  assign y6995 = ~1'b0 ;
  assign y6996 = n22656 ;
  assign y6997 = ~n22660 ;
  assign y6998 = n22662 ;
  assign y6999 = ~n22663 ;
  assign y7000 = ~n22665 ;
  assign y7001 = ~n22669 ;
  assign y7002 = n22671 ;
  assign y7003 = ~n22674 ;
  assign y7004 = ~n22677 ;
  assign y7005 = ~1'b0 ;
  assign y7006 = ~n22678 ;
  assign y7007 = ~n22681 ;
  assign y7008 = ~n22682 ;
  assign y7009 = ~n22685 ;
  assign y7010 = ~n22688 ;
  assign y7011 = n22692 ;
  assign y7012 = n22694 ;
  assign y7013 = n22695 ;
  assign y7014 = ~n22700 ;
  assign y7015 = n22701 ;
  assign y7016 = ~n22702 ;
  assign y7017 = n22703 ;
  assign y7018 = n22708 ;
  assign y7019 = n22710 ;
  assign y7020 = ~n22712 ;
  assign y7021 = n22716 ;
  assign y7022 = ~n22719 ;
  assign y7023 = n22720 ;
  assign y7024 = ~n22721 ;
  assign y7025 = n22728 ;
  assign y7026 = n22732 ;
  assign y7027 = ~n22735 ;
  assign y7028 = ~n22737 ;
  assign y7029 = ~n22739 ;
  assign y7030 = ~n22740 ;
  assign y7031 = ~1'b0 ;
  assign y7032 = ~n22742 ;
  assign y7033 = n22743 ;
  assign y7034 = ~n22746 ;
  assign y7035 = ~n22751 ;
  assign y7036 = ~1'b0 ;
  assign y7037 = ~n22752 ;
  assign y7038 = ~n22753 ;
  assign y7039 = n22754 ;
  assign y7040 = n8762 ;
  assign y7041 = ~n22756 ;
  assign y7042 = n22758 ;
  assign y7043 = n22760 ;
  assign y7044 = ~1'b0 ;
  assign y7045 = ~n22763 ;
  assign y7046 = ~1'b0 ;
  assign y7047 = ~n22767 ;
  assign y7048 = ~n22768 ;
  assign y7049 = n22777 ;
  assign y7050 = ~n22779 ;
  assign y7051 = n22786 ;
  assign y7052 = ~n22790 ;
  assign y7053 = n22793 ;
  assign y7054 = n22794 ;
  assign y7055 = n22798 ;
  assign y7056 = ~1'b0 ;
  assign y7057 = n22799 ;
  assign y7058 = ~n10777 ;
  assign y7059 = ~n22802 ;
  assign y7060 = ~n22809 ;
  assign y7061 = n22815 ;
  assign y7062 = ~n22821 ;
  assign y7063 = n22823 ;
  assign y7064 = ~n22825 ;
  assign y7065 = ~n22830 ;
  assign y7066 = ~n22831 ;
  assign y7067 = n22834 ;
  assign y7068 = n22835 ;
  assign y7069 = n22839 ;
  assign y7070 = ~n22846 ;
  assign y7071 = ~n22847 ;
  assign y7072 = ~n22848 ;
  assign y7073 = ~n22850 ;
  assign y7074 = ~1'b0 ;
  assign y7075 = n22851 ;
  assign y7076 = n6477 ;
  assign y7077 = n22852 ;
  assign y7078 = n22853 ;
  assign y7079 = ~n22855 ;
  assign y7080 = ~1'b0 ;
  assign y7081 = ~1'b0 ;
  assign y7082 = n22856 ;
  assign y7083 = n22857 ;
  assign y7084 = n22865 ;
  assign y7085 = n22866 ;
  assign y7086 = n22873 ;
  assign y7087 = ~n22874 ;
  assign y7088 = ~n22876 ;
  assign y7089 = n22878 ;
  assign y7090 = n22882 ;
  assign y7091 = ~n22884 ;
  assign y7092 = ~n22887 ;
  assign y7093 = ~n22889 ;
  assign y7094 = n22892 ;
  assign y7095 = n22894 ;
  assign y7096 = ~1'b0 ;
  assign y7097 = ~1'b0 ;
  assign y7098 = n22895 ;
  assign y7099 = n22900 ;
  assign y7100 = n22906 ;
  assign y7101 = ~n22910 ;
  assign y7102 = n22912 ;
  assign y7103 = ~1'b0 ;
  assign y7104 = ~n22916 ;
  assign y7105 = ~n22920 ;
  assign y7106 = ~n22922 ;
  assign y7107 = ~n22925 ;
  assign y7108 = n22928 ;
  assign y7109 = ~n22929 ;
  assign y7110 = ~1'b0 ;
  assign y7111 = ~n22932 ;
  assign y7112 = n22937 ;
  assign y7113 = ~n22939 ;
  assign y7114 = ~n22943 ;
  assign y7115 = n22944 ;
  assign y7116 = n22945 ;
  assign y7117 = n22946 ;
  assign y7118 = n22949 ;
  assign y7119 = ~n22950 ;
  assign y7120 = ~1'b0 ;
  assign y7121 = n22952 ;
  assign y7122 = n22961 ;
  assign y7123 = ~n22962 ;
  assign y7124 = n22964 ;
  assign y7125 = ~1'b0 ;
  assign y7126 = n22966 ;
  assign y7127 = ~1'b0 ;
  assign y7128 = n22970 ;
  assign y7129 = ~n22974 ;
  assign y7130 = ~n13493 ;
  assign y7131 = n22979 ;
  assign y7132 = n22981 ;
  assign y7133 = ~n22982 ;
  assign y7134 = ~1'b0 ;
  assign y7135 = ~1'b0 ;
  assign y7136 = ~n22986 ;
  assign y7137 = n22988 ;
  assign y7138 = ~n22989 ;
  assign y7139 = ~1'b0 ;
  assign y7140 = ~1'b0 ;
  assign y7141 = n22991 ;
  assign y7142 = ~n22996 ;
  assign y7143 = n22999 ;
  assign y7144 = ~n23001 ;
  assign y7145 = n23004 ;
  assign y7146 = ~n23006 ;
  assign y7147 = ~1'b0 ;
  assign y7148 = ~1'b0 ;
  assign y7149 = ~n23008 ;
  assign y7150 = ~n23009 ;
  assign y7151 = n23010 ;
  assign y7152 = n23012 ;
  assign y7153 = n13918 ;
  assign y7154 = n23016 ;
  assign y7155 = ~n23018 ;
  assign y7156 = n23019 ;
  assign y7157 = ~n23020 ;
  assign y7158 = n23022 ;
  assign y7159 = ~n23023 ;
  assign y7160 = ~1'b0 ;
  assign y7161 = n23024 ;
  assign y7162 = n23029 ;
  assign y7163 = n23032 ;
  assign y7164 = ~n23034 ;
  assign y7165 = n23035 ;
  assign y7166 = n23036 ;
  assign y7167 = n23044 ;
  assign y7168 = ~1'b0 ;
  assign y7169 = ~1'b0 ;
  assign y7170 = ~1'b0 ;
  assign y7171 = ~1'b0 ;
  assign y7172 = ~n23045 ;
  assign y7173 = ~n23046 ;
  assign y7174 = n23056 ;
  assign y7175 = ~n23057 ;
  assign y7176 = n23058 ;
  assign y7177 = n23060 ;
  assign y7178 = n23062 ;
  assign y7179 = n23064 ;
  assign y7180 = ~n23071 ;
  assign y7181 = n23073 ;
  assign y7182 = n702 ;
  assign y7183 = ~n23075 ;
  assign y7184 = ~n23080 ;
  assign y7185 = ~n23081 ;
  assign y7186 = n23084 ;
  assign y7187 = ~n23086 ;
  assign y7188 = ~n23093 ;
  assign y7189 = n23094 ;
  assign y7190 = n23096 ;
  assign y7191 = n23098 ;
  assign y7192 = n23101 ;
  assign y7193 = ~1'b0 ;
  assign y7194 = ~n23102 ;
  assign y7195 = ~n23107 ;
  assign y7196 = ~n23112 ;
  assign y7197 = ~n23114 ;
  assign y7198 = n23118 ;
  assign y7199 = ~n23119 ;
  assign y7200 = n23121 ;
  assign y7201 = n23122 ;
  assign y7202 = n23123 ;
  assign y7203 = ~n23125 ;
  assign y7204 = ~1'b0 ;
  assign y7205 = n23132 ;
  assign y7206 = ~n23134 ;
  assign y7207 = ~1'b0 ;
  assign y7208 = ~n23135 ;
  assign y7209 = n23136 ;
  assign y7210 = n23141 ;
  assign y7211 = n23146 ;
  assign y7212 = n23150 ;
  assign y7213 = ~1'b0 ;
  assign y7214 = n23154 ;
  assign y7215 = ~n23156 ;
  assign y7216 = ~n23157 ;
  assign y7217 = n23158 ;
  assign y7218 = ~1'b0 ;
  assign y7219 = ~n23160 ;
  assign y7220 = ~n23162 ;
  assign y7221 = ~n23163 ;
  assign y7222 = n23164 ;
  assign y7223 = n23166 ;
  assign y7224 = n23167 ;
  assign y7225 = ~1'b0 ;
  assign y7226 = ~n23172 ;
  assign y7227 = ~n23175 ;
  assign y7228 = ~n1968 ;
  assign y7229 = ~n23184 ;
  assign y7230 = n23187 ;
  assign y7231 = n23190 ;
  assign y7232 = ~n23191 ;
  assign y7233 = n23194 ;
  assign y7234 = ~n23196 ;
  assign y7235 = n23197 ;
  assign y7236 = n23201 ;
  assign y7237 = n23202 ;
  assign y7238 = n23203 ;
  assign y7239 = ~n23207 ;
  assign y7240 = n23219 ;
  assign y7241 = ~1'b0 ;
  assign y7242 = ~1'b0 ;
  assign y7243 = n23220 ;
  assign y7244 = ~1'b0 ;
  assign y7245 = n23225 ;
  assign y7246 = ~n23228 ;
  assign y7247 = n23229 ;
  assign y7248 = n23232 ;
  assign y7249 = n23238 ;
  assign y7250 = ~1'b0 ;
  assign y7251 = n23246 ;
  assign y7252 = ~n23247 ;
  assign y7253 = ~n23251 ;
  assign y7254 = ~n23253 ;
  assign y7255 = ~1'b0 ;
  assign y7256 = ~1'b0 ;
  assign y7257 = n23255 ;
  assign y7258 = ~n23256 ;
  assign y7259 = ~n23258 ;
  assign y7260 = ~1'b0 ;
  assign y7261 = ~1'b0 ;
  assign y7262 = n23263 ;
  assign y7263 = ~1'b0 ;
  assign y7264 = ~n23267 ;
  assign y7265 = ~n23268 ;
  assign y7266 = n23270 ;
  assign y7267 = n23274 ;
  assign y7268 = ~n23278 ;
  assign y7269 = ~n23279 ;
  assign y7270 = ~n23283 ;
  assign y7271 = ~1'b0 ;
  assign y7272 = n23286 ;
  assign y7273 = ~n23287 ;
  assign y7274 = n23288 ;
  assign y7275 = 1'b0 ;
  assign y7276 = n23291 ;
  assign y7277 = n23294 ;
  assign y7278 = ~1'b0 ;
  assign y7279 = ~n23297 ;
  assign y7280 = ~n23298 ;
  assign y7281 = ~n23300 ;
  assign y7282 = n23306 ;
  assign y7283 = ~1'b0 ;
  assign y7284 = ~n23308 ;
  assign y7285 = ~1'b0 ;
  assign y7286 = ~n23309 ;
  assign y7287 = ~n23311 ;
  assign y7288 = ~1'b0 ;
  assign y7289 = ~n23315 ;
  assign y7290 = n23317 ;
  assign y7291 = n23319 ;
  assign y7292 = ~n23321 ;
  assign y7293 = n23324 ;
  assign y7294 = n23325 ;
  assign y7295 = n23327 ;
  assign y7296 = ~1'b0 ;
  assign y7297 = ~n23330 ;
  assign y7298 = ~n23332 ;
  assign y7299 = n23333 ;
  assign y7300 = n23336 ;
  assign y7301 = n23337 ;
  assign y7302 = n23340 ;
  assign y7303 = ~n23342 ;
  assign y7304 = n23346 ;
  assign y7305 = ~n23348 ;
  assign y7306 = n23351 ;
  assign y7307 = ~n23352 ;
  assign y7308 = ~n23353 ;
  assign y7309 = ~1'b0 ;
  assign y7310 = ~n23357 ;
  assign y7311 = n23360 ;
  assign y7312 = ~1'b0 ;
  assign y7313 = n23361 ;
  assign y7314 = n23363 ;
  assign y7315 = ~n23365 ;
  assign y7316 = ~n23368 ;
  assign y7317 = ~n23370 ;
  assign y7318 = n23372 ;
  assign y7319 = n23373 ;
  assign y7320 = n23376 ;
  assign y7321 = n23378 ;
  assign y7322 = n23380 ;
  assign y7323 = n23381 ;
  assign y7324 = n23384 ;
  assign y7325 = n23387 ;
  assign y7326 = ~n23389 ;
  assign y7327 = ~1'b0 ;
  assign y7328 = ~n23390 ;
  assign y7329 = ~n23391 ;
  assign y7330 = ~n23394 ;
  assign y7331 = n23396 ;
  assign y7332 = ~n23399 ;
  assign y7333 = ~1'b0 ;
  assign y7334 = ~n23403 ;
  assign y7335 = ~n23404 ;
  assign y7336 = n23407 ;
  assign y7337 = ~n23408 ;
  assign y7338 = ~n23410 ;
  assign y7339 = ~1'b0 ;
  assign y7340 = n23411 ;
  assign y7341 = n23412 ;
  assign y7342 = n23414 ;
  assign y7343 = ~n23415 ;
  assign y7344 = ~n23416 ;
  assign y7345 = ~n23417 ;
  assign y7346 = ~1'b0 ;
  assign y7347 = ~n23418 ;
  assign y7348 = n23420 ;
  assign y7349 = ~n23421 ;
  assign y7350 = n23424 ;
  assign y7351 = n2934 ;
  assign y7352 = n23428 ;
  assign y7353 = n23432 ;
  assign y7354 = ~n23437 ;
  assign y7355 = ~n23443 ;
  assign y7356 = ~n23444 ;
  assign y7357 = ~n23445 ;
  assign y7358 = ~n23447 ;
  assign y7359 = n23449 ;
  assign y7360 = ~1'b0 ;
  assign y7361 = n23456 ;
  assign y7362 = n23460 ;
  assign y7363 = ~n23461 ;
  assign y7364 = n23462 ;
  assign y7365 = n23466 ;
  assign y7366 = ~n23468 ;
  assign y7367 = ~n23469 ;
  assign y7368 = n23470 ;
  assign y7369 = n23478 ;
  assign y7370 = n23480 ;
  assign y7371 = ~n23487 ;
  assign y7372 = ~n23490 ;
  assign y7373 = n23495 ;
  assign y7374 = n23497 ;
  assign y7375 = n23498 ;
  assign y7376 = ~n23507 ;
  assign y7377 = ~n23511 ;
  assign y7378 = ~n23514 ;
  assign y7379 = ~n23516 ;
  assign y7380 = n23518 ;
  assign y7381 = ~n23520 ;
  assign y7382 = ~n23526 ;
  assign y7383 = n23527 ;
  assign y7384 = ~n23529 ;
  assign y7385 = ~n23531 ;
  assign y7386 = ~n23541 ;
  assign y7387 = ~n23544 ;
  assign y7388 = ~n23545 ;
  assign y7389 = ~n23548 ;
  assign y7390 = ~n23549 ;
  assign y7391 = n23557 ;
  assign y7392 = ~n23560 ;
  assign y7393 = ~1'b0 ;
  assign y7394 = ~n23563 ;
  assign y7395 = n23565 ;
  assign y7396 = ~n23567 ;
  assign y7397 = ~n23569 ;
  assign y7398 = n23572 ;
  assign y7399 = ~n23575 ;
  assign y7400 = ~n23579 ;
  assign y7401 = n23582 ;
  assign y7402 = n23595 ;
  assign y7403 = ~n23599 ;
  assign y7404 = ~n23601 ;
  assign y7405 = ~n23602 ;
  assign y7406 = ~n23604 ;
  assign y7407 = ~n23605 ;
  assign y7408 = ~n23610 ;
  assign y7409 = n23612 ;
  assign y7410 = n23614 ;
  assign y7411 = ~n23616 ;
  assign y7412 = ~n23617 ;
  assign y7413 = n23620 ;
  assign y7414 = n23622 ;
  assign y7415 = n23623 ;
  assign y7416 = n23627 ;
  assign y7417 = ~1'b0 ;
  assign y7418 = n23629 ;
  assign y7419 = ~1'b0 ;
  assign y7420 = ~n23631 ;
  assign y7421 = ~n23632 ;
  assign y7422 = ~n23633 ;
  assign y7423 = ~n23638 ;
  assign y7424 = n23641 ;
  assign y7425 = ~1'b0 ;
  assign y7426 = n23652 ;
  assign y7427 = n23653 ;
  assign y7428 = ~n23655 ;
  assign y7429 = n23656 ;
  assign y7430 = n8344 ;
  assign y7431 = n23657 ;
  assign y7432 = n23660 ;
  assign y7433 = ~n23663 ;
  assign y7434 = ~n23666 ;
  assign y7435 = n23670 ;
  assign y7436 = ~1'b0 ;
  assign y7437 = ~n23672 ;
  assign y7438 = ~n23673 ;
  assign y7439 = n23675 ;
  assign y7440 = ~n23676 ;
  assign y7441 = n23678 ;
  assign y7442 = n23682 ;
  assign y7443 = n23689 ;
  assign y7444 = ~1'b0 ;
  assign y7445 = ~n23691 ;
  assign y7446 = ~n23693 ;
  assign y7447 = ~n23697 ;
  assign y7448 = n23699 ;
  assign y7449 = ~n23701 ;
  assign y7450 = ~1'b0 ;
  assign y7451 = ~n23704 ;
  assign y7452 = n23706 ;
  assign y7453 = ~n23708 ;
  assign y7454 = n23709 ;
  assign y7455 = n23713 ;
  assign y7456 = n23721 ;
  assign y7457 = ~n23726 ;
  assign y7458 = ~n23727 ;
  assign y7459 = n23729 ;
  assign y7460 = ~1'b0 ;
  assign y7461 = n23736 ;
  assign y7462 = ~n23741 ;
  assign y7463 = ~n23742 ;
  assign y7464 = n23743 ;
  assign y7465 = ~n23749 ;
  assign y7466 = ~n23759 ;
  assign y7467 = n23765 ;
  assign y7468 = n23766 ;
  assign y7469 = ~n23770 ;
  assign y7470 = ~n23774 ;
  assign y7471 = n23777 ;
  assign y7472 = n23778 ;
  assign y7473 = n23780 ;
  assign y7474 = ~n23783 ;
  assign y7475 = n23785 ;
  assign y7476 = n23787 ;
  assign y7477 = n23788 ;
  assign y7478 = ~n23790 ;
  assign y7479 = n23792 ;
  assign y7480 = ~n23794 ;
  assign y7481 = ~n23799 ;
  assign y7482 = n23802 ;
  assign y7483 = n23805 ;
  assign y7484 = ~n23806 ;
  assign y7485 = n23808 ;
  assign y7486 = ~n23810 ;
  assign y7487 = n23815 ;
  assign y7488 = ~n23820 ;
  assign y7489 = ~n23821 ;
  assign y7490 = ~n23826 ;
  assign y7491 = n23830 ;
  assign y7492 = ~n23835 ;
  assign y7493 = ~1'b0 ;
  assign y7494 = n23838 ;
  assign y7495 = n23839 ;
  assign y7496 = n23842 ;
  assign y7497 = n3121 ;
  assign y7498 = n23844 ;
  assign y7499 = n23846 ;
  assign y7500 = ~n23848 ;
  assign y7501 = n23849 ;
  assign y7502 = ~n23850 ;
  assign y7503 = ~n23852 ;
  assign y7504 = n23853 ;
  assign y7505 = n23854 ;
  assign y7506 = ~n23856 ;
  assign y7507 = ~n23857 ;
  assign y7508 = n23859 ;
  assign y7509 = n23862 ;
  assign y7510 = n23863 ;
  assign y7511 = n23865 ;
  assign y7512 = ~n23866 ;
  assign y7513 = n23869 ;
  assign y7514 = n23871 ;
  assign y7515 = n23874 ;
  assign y7516 = n9571 ;
  assign y7517 = n23876 ;
  assign y7518 = n23878 ;
  assign y7519 = ~n23882 ;
  assign y7520 = ~n23883 ;
  assign y7521 = ~n23884 ;
  assign y7522 = ~n23888 ;
  assign y7523 = n23894 ;
  assign y7524 = ~1'b0 ;
  assign y7525 = ~n23896 ;
  assign y7526 = n23897 ;
  assign y7527 = ~n23899 ;
  assign y7528 = n23901 ;
  assign y7529 = n23904 ;
  assign y7530 = n23908 ;
  assign y7531 = n23910 ;
  assign y7532 = ~n23914 ;
  assign y7533 = ~n23918 ;
  assign y7534 = n23919 ;
  assign y7535 = n23920 ;
  assign y7536 = n23926 ;
  assign y7537 = ~n23938 ;
  assign y7538 = ~1'b0 ;
  assign y7539 = n23940 ;
  assign y7540 = n23942 ;
  assign y7541 = ~n23943 ;
  assign y7542 = ~n23944 ;
  assign y7543 = n23945 ;
  assign y7544 = ~1'b0 ;
  assign y7545 = ~n23946 ;
  assign y7546 = ~n23947 ;
  assign y7547 = ~n23951 ;
  assign y7548 = n23959 ;
  assign y7549 = n23961 ;
  assign y7550 = n23962 ;
  assign y7551 = ~n23965 ;
  assign y7552 = ~n23967 ;
  assign y7553 = ~n23969 ;
  assign y7554 = n23973 ;
  assign y7555 = n23977 ;
  assign y7556 = ~n23978 ;
  assign y7557 = n23979 ;
  assign y7558 = n23981 ;
  assign y7559 = ~n23983 ;
  assign y7560 = ~n13937 ;
  assign y7561 = ~n23989 ;
  assign y7562 = ~n23993 ;
  assign y7563 = n23994 ;
  assign y7564 = ~n23996 ;
  assign y7565 = ~n23998 ;
  assign y7566 = ~n24000 ;
  assign y7567 = ~n24001 ;
  assign y7568 = ~n24005 ;
  assign y7569 = ~n24008 ;
  assign y7570 = n24009 ;
  assign y7571 = ~n24011 ;
  assign y7572 = ~n24015 ;
  assign y7573 = n24018 ;
  assign y7574 = ~1'b0 ;
  assign y7575 = ~n24021 ;
  assign y7576 = n24022 ;
  assign y7577 = n24023 ;
  assign y7578 = n24027 ;
  assign y7579 = n24028 ;
  assign y7580 = ~n24034 ;
  assign y7581 = n24037 ;
  assign y7582 = ~1'b0 ;
  assign y7583 = n24038 ;
  assign y7584 = ~n24040 ;
  assign y7585 = n24041 ;
  assign y7586 = ~n24042 ;
  assign y7587 = n24044 ;
  assign y7588 = n24050 ;
  assign y7589 = ~1'b0 ;
  assign y7590 = n24057 ;
  assign y7591 = n24058 ;
  assign y7592 = ~n24062 ;
  assign y7593 = n24064 ;
  assign y7594 = n24067 ;
  assign y7595 = ~n24070 ;
  assign y7596 = ~1'b0 ;
  assign y7597 = ~n24071 ;
  assign y7598 = ~n24077 ;
  assign y7599 = ~n24078 ;
  assign y7600 = n24079 ;
  assign y7601 = ~n24081 ;
  assign y7602 = ~n24082 ;
  assign y7603 = ~n24083 ;
  assign y7604 = ~n24084 ;
  assign y7605 = n24088 ;
  assign y7606 = n24089 ;
  assign y7607 = ~n24090 ;
  assign y7608 = n24091 ;
  assign y7609 = n24094 ;
  assign y7610 = ~n24097 ;
  assign y7611 = ~1'b0 ;
  assign y7612 = n24102 ;
  assign y7613 = ~n24104 ;
  assign y7614 = n24106 ;
  assign y7615 = n24111 ;
  assign y7616 = ~n24114 ;
  assign y7617 = n24115 ;
  assign y7618 = ~n24117 ;
  assign y7619 = ~1'b0 ;
  assign y7620 = ~1'b0 ;
  assign y7621 = ~n24121 ;
  assign y7622 = n24122 ;
  assign y7623 = ~n24125 ;
  assign y7624 = ~n24126 ;
  assign y7625 = ~n24131 ;
  assign y7626 = ~1'b0 ;
  assign y7627 = ~1'b0 ;
  assign y7628 = n24132 ;
  assign y7629 = n24134 ;
  assign y7630 = ~n24135 ;
  assign y7631 = n24136 ;
  assign y7632 = ~n24142 ;
  assign y7633 = ~n24148 ;
  assign y7634 = n24149 ;
  assign y7635 = ~n24158 ;
  assign y7636 = ~n24160 ;
  assign y7637 = ~1'b0 ;
  assign y7638 = ~1'b0 ;
  assign y7639 = n24165 ;
  assign y7640 = ~n24166 ;
  assign y7641 = n24168 ;
  assign y7642 = n24174 ;
  assign y7643 = n24175 ;
  assign y7644 = ~1'b0 ;
  assign y7645 = ~n24177 ;
  assign y7646 = n24180 ;
  assign y7647 = ~n24181 ;
  assign y7648 = ~n24183 ;
  assign y7649 = n24184 ;
  assign y7650 = n24186 ;
  assign y7651 = ~1'b0 ;
  assign y7652 = n24187 ;
  assign y7653 = ~n24191 ;
  assign y7654 = n24193 ;
  assign y7655 = ~1'b0 ;
  assign y7656 = ~n24197 ;
  assign y7657 = n24201 ;
  assign y7658 = ~n24202 ;
  assign y7659 = ~n24203 ;
  assign y7660 = ~n24206 ;
  assign y7661 = ~1'b0 ;
  assign y7662 = ~1'b0 ;
  assign y7663 = ~n19382 ;
  assign y7664 = ~n24208 ;
  assign y7665 = n24211 ;
  assign y7666 = n24212 ;
  assign y7667 = n24214 ;
  assign y7668 = ~1'b0 ;
  assign y7669 = n24215 ;
  assign y7670 = n24220 ;
  assign y7671 = ~n24222 ;
  assign y7672 = ~n24224 ;
  assign y7673 = n24226 ;
  assign y7674 = n24228 ;
  assign y7675 = n24231 ;
  assign y7676 = n24234 ;
  assign y7677 = n24237 ;
  assign y7678 = ~n24239 ;
  assign y7679 = n24242 ;
  assign y7680 = ~n24243 ;
  assign y7681 = ~n24250 ;
  assign y7682 = n10444 ;
  assign y7683 = ~n24252 ;
  assign y7684 = ~1'b0 ;
  assign y7685 = n24258 ;
  assign y7686 = ~n24262 ;
  assign y7687 = n24266 ;
  assign y7688 = n24270 ;
  assign y7689 = n24272 ;
  assign y7690 = ~1'b0 ;
  assign y7691 = ~1'b0 ;
  assign y7692 = ~1'b0 ;
  assign y7693 = ~1'b0 ;
  assign y7694 = ~n24276 ;
  assign y7695 = n24277 ;
  assign y7696 = ~n24278 ;
  assign y7697 = n24284 ;
  assign y7698 = ~n24286 ;
  assign y7699 = ~1'b0 ;
  assign y7700 = n24288 ;
  assign y7701 = n24294 ;
  assign y7702 = ~n24295 ;
  assign y7703 = n24297 ;
  assign y7704 = n24299 ;
  assign y7705 = n24302 ;
  assign y7706 = n24304 ;
  assign y7707 = n24306 ;
  assign y7708 = ~n24308 ;
  assign y7709 = ~n24310 ;
  assign y7710 = n24312 ;
  assign y7711 = n24314 ;
  assign y7712 = ~1'b0 ;
  assign y7713 = n24319 ;
  assign y7714 = ~n24324 ;
  assign y7715 = ~1'b0 ;
  assign y7716 = ~n24329 ;
  assign y7717 = n24334 ;
  assign y7718 = ~n24335 ;
  assign y7719 = ~1'b0 ;
  assign y7720 = n24337 ;
  assign y7721 = ~n24338 ;
  assign y7722 = ~n24340 ;
  assign y7723 = n24343 ;
  assign y7724 = ~n24344 ;
  assign y7725 = ~n24347 ;
  assign y7726 = n24348 ;
  assign y7727 = n24349 ;
  assign y7728 = n24355 ;
  assign y7729 = ~n24358 ;
  assign y7730 = ~n24372 ;
  assign y7731 = n24375 ;
  assign y7732 = ~n24379 ;
  assign y7733 = ~n24380 ;
  assign y7734 = ~n24382 ;
  assign y7735 = n24392 ;
  assign y7736 = ~n24393 ;
  assign y7737 = ~n24397 ;
  assign y7738 = n24401 ;
  assign y7739 = ~n24402 ;
  assign y7740 = n24404 ;
  assign y7741 = 1'b0 ;
  assign y7742 = n24408 ;
  assign y7743 = n24409 ;
  assign y7744 = ~n24411 ;
  assign y7745 = ~n24412 ;
  assign y7746 = ~n24416 ;
  assign y7747 = ~n24417 ;
  assign y7748 = ~1'b0 ;
  assign y7749 = ~n24420 ;
  assign y7750 = ~1'b0 ;
  assign y7751 = ~n24426 ;
  assign y7752 = ~n24428 ;
  assign y7753 = n8195 ;
  assign y7754 = ~1'b0 ;
  assign y7755 = ~n24429 ;
  assign y7756 = ~1'b0 ;
  assign y7757 = ~n7536 ;
  assign y7758 = ~n24430 ;
  assign y7759 = ~n24431 ;
  assign y7760 = n24439 ;
  assign y7761 = n24445 ;
  assign y7762 = ~1'b0 ;
  assign y7763 = ~1'b0 ;
  assign y7764 = ~n24448 ;
  assign y7765 = ~n24452 ;
  assign y7766 = ~1'b0 ;
  assign y7767 = ~n24456 ;
  assign y7768 = n24461 ;
  assign y7769 = n24469 ;
  assign y7770 = ~n24472 ;
  assign y7771 = ~n24476 ;
  assign y7772 = n24480 ;
  assign y7773 = ~n24483 ;
  assign y7774 = n24487 ;
  assign y7775 = ~n24490 ;
  assign y7776 = n24492 ;
  assign y7777 = ~n24495 ;
  assign y7778 = ~n24498 ;
  assign y7779 = n24500 ;
  assign y7780 = ~n24503 ;
  assign y7781 = n24508 ;
  assign y7782 = n24509 ;
  assign y7783 = ~1'b0 ;
  assign y7784 = n24514 ;
  assign y7785 = ~n24519 ;
  assign y7786 = ~n24528 ;
  assign y7787 = ~n24529 ;
  assign y7788 = n24536 ;
  assign y7789 = n24540 ;
  assign y7790 = n24542 ;
  assign y7791 = 1'b0 ;
  assign y7792 = n24543 ;
  assign y7793 = n24546 ;
  assign y7794 = n24552 ;
  assign y7795 = ~n24557 ;
  assign y7796 = ~n24558 ;
  assign y7797 = n24564 ;
  assign y7798 = n24565 ;
  assign y7799 = ~1'b0 ;
  assign y7800 = ~n24569 ;
  assign y7801 = n24575 ;
  assign y7802 = ~n24576 ;
  assign y7803 = n24578 ;
  assign y7804 = n24585 ;
  assign y7805 = ~n24591 ;
  assign y7806 = ~n24592 ;
  assign y7807 = n24594 ;
  assign y7808 = n24598 ;
  assign y7809 = ~1'b0 ;
  assign y7810 = ~1'b0 ;
  assign y7811 = ~n24601 ;
  assign y7812 = n24603 ;
  assign y7813 = ~n24605 ;
  assign y7814 = ~n24606 ;
  assign y7815 = ~n24607 ;
  assign y7816 = n24611 ;
  assign y7817 = n24612 ;
  assign y7818 = ~n24615 ;
  assign y7819 = n24616 ;
  assign y7820 = n24619 ;
  assign y7821 = n24620 ;
  assign y7822 = n24621 ;
  assign y7823 = ~n12538 ;
  assign y7824 = ~1'b0 ;
  assign y7825 = ~n24624 ;
  assign y7826 = ~n24629 ;
  assign y7827 = ~n24630 ;
  assign y7828 = ~n24633 ;
  assign y7829 = ~n24634 ;
  assign y7830 = n24641 ;
  assign y7831 = n24644 ;
  assign y7832 = n24647 ;
  assign y7833 = ~n24655 ;
  assign y7834 = ~n24657 ;
  assign y7835 = ~n9205 ;
  assign y7836 = n24662 ;
  assign y7837 = ~n24663 ;
  assign y7838 = n24668 ;
  assign y7839 = ~n24670 ;
  assign y7840 = ~1'b0 ;
  assign y7841 = ~1'b0 ;
  assign y7842 = n24671 ;
  assign y7843 = n4607 ;
  assign y7844 = ~n24673 ;
  assign y7845 = n24674 ;
  assign y7846 = n24683 ;
  assign y7847 = ~n24686 ;
  assign y7848 = ~1'b0 ;
  assign y7849 = ~n24687 ;
  assign y7850 = n24695 ;
  assign y7851 = ~n24697 ;
  assign y7852 = n24699 ;
  assign y7853 = n24703 ;
  assign y7854 = ~1'b0 ;
  assign y7855 = n24705 ;
  assign y7856 = ~n24707 ;
  assign y7857 = ~n24708 ;
  assign y7858 = ~n24710 ;
  assign y7859 = ~n24713 ;
  assign y7860 = ~n24715 ;
  assign y7861 = ~1'b0 ;
  assign y7862 = ~n24716 ;
  assign y7863 = ~n24718 ;
  assign y7864 = n24720 ;
  assign y7865 = n24721 ;
  assign y7866 = ~n24722 ;
  assign y7867 = 1'b0 ;
  assign y7868 = n24729 ;
  assign y7869 = ~1'b0 ;
  assign y7870 = ~1'b0 ;
  assign y7871 = n23471 ;
  assign y7872 = n24730 ;
  assign y7873 = n24734 ;
  assign y7874 = ~n24735 ;
  assign y7875 = n24739 ;
  assign y7876 = ~n24740 ;
  assign y7877 = n24743 ;
  assign y7878 = n24750 ;
  assign y7879 = n24755 ;
  assign y7880 = ~n24761 ;
  assign y7881 = n24764 ;
  assign y7882 = n24767 ;
  assign y7883 = n24771 ;
  assign y7884 = n24778 ;
  assign y7885 = ~n24780 ;
  assign y7886 = n24783 ;
  assign y7887 = n24784 ;
  assign y7888 = ~1'b0 ;
  assign y7889 = n24787 ;
  assign y7890 = n24790 ;
  assign y7891 = ~n24792 ;
  assign y7892 = ~n24793 ;
  assign y7893 = n24798 ;
  assign y7894 = ~1'b0 ;
  assign y7895 = ~n24802 ;
  assign y7896 = ~n24806 ;
  assign y7897 = ~1'b0 ;
  assign y7898 = ~n24811 ;
  assign y7899 = n24813 ;
  assign y7900 = ~1'b0 ;
  assign y7901 = ~n24819 ;
  assign y7902 = ~n24822 ;
  assign y7903 = ~n24824 ;
  assign y7904 = n24826 ;
  assign y7905 = ~n24827 ;
  assign y7906 = ~n24828 ;
  assign y7907 = ~n24836 ;
  assign y7908 = ~n24837 ;
  assign y7909 = n24838 ;
  assign y7910 = n24847 ;
  assign y7911 = n24850 ;
  assign y7912 = ~n24852 ;
  assign y7913 = ~n24854 ;
  assign y7914 = n24855 ;
  assign y7915 = ~n24856 ;
  assign y7916 = ~n24860 ;
  assign y7917 = n24861 ;
  assign y7918 = n24864 ;
  assign y7919 = ~n24867 ;
  assign y7920 = ~1'b0 ;
  assign y7921 = n24869 ;
  assign y7922 = ~1'b0 ;
  assign y7923 = n24871 ;
  assign y7924 = n24874 ;
  assign y7925 = ~n24877 ;
  assign y7926 = ~n24880 ;
  assign y7927 = n24882 ;
  assign y7928 = n24892 ;
  assign y7929 = n24896 ;
  assign y7930 = ~1'b0 ;
  assign y7931 = n24899 ;
  assign y7932 = ~n24900 ;
  assign y7933 = n24902 ;
  assign y7934 = n24903 ;
  assign y7935 = ~n24905 ;
  assign y7936 = ~n19307 ;
  assign y7937 = n24907 ;
  assign y7938 = ~n24913 ;
  assign y7939 = n24920 ;
  assign y7940 = ~n24921 ;
  assign y7941 = n24927 ;
  assign y7942 = ~n24928 ;
  assign y7943 = ~1'b0 ;
  assign y7944 = n24932 ;
  assign y7945 = ~1'b0 ;
  assign y7946 = ~n24936 ;
  assign y7947 = ~n24938 ;
  assign y7948 = ~n24950 ;
  assign y7949 = ~n24955 ;
  assign y7950 = ~1'b0 ;
  assign y7951 = n24962 ;
  assign y7952 = n24963 ;
  assign y7953 = ~1'b0 ;
  assign y7954 = ~n24966 ;
  assign y7955 = n24968 ;
  assign y7956 = ~n24970 ;
  assign y7957 = n24971 ;
  assign y7958 = ~n24974 ;
  assign y7959 = n24975 ;
  assign y7960 = ~n24977 ;
  assign y7961 = ~n24979 ;
  assign y7962 = n24984 ;
  assign y7963 = n24989 ;
  assign y7964 = ~n25000 ;
  assign y7965 = ~n25003 ;
  assign y7966 = ~n25004 ;
  assign y7967 = ~n25007 ;
  assign y7968 = n25009 ;
  assign y7969 = ~1'b0 ;
  assign y7970 = ~n25011 ;
  assign y7971 = n25014 ;
  assign y7972 = ~n25020 ;
  assign y7973 = ~n25021 ;
  assign y7974 = ~n25026 ;
  assign y7975 = ~n25027 ;
  assign y7976 = ~1'b0 ;
  assign y7977 = ~1'b0 ;
  assign y7978 = ~1'b0 ;
  assign y7979 = n25030 ;
  assign y7980 = ~1'b0 ;
  assign y7981 = ~n25033 ;
  assign y7982 = ~1'b0 ;
  assign y7983 = n25038 ;
  assign y7984 = ~n25045 ;
  assign y7985 = n25047 ;
  assign y7986 = ~1'b0 ;
  assign y7987 = ~1'b0 ;
  assign y7988 = ~n25050 ;
  assign y7989 = n25051 ;
  assign y7990 = ~n25058 ;
  assign y7991 = ~n7031 ;
  assign y7992 = n25061 ;
  assign y7993 = n25063 ;
  assign y7994 = ~1'b0 ;
  assign y7995 = ~1'b0 ;
  assign y7996 = ~n25065 ;
  assign y7997 = ~1'b0 ;
  assign y7998 = n25066 ;
  assign y7999 = n25068 ;
  assign y8000 = ~1'b0 ;
  assign y8001 = ~n25069 ;
  assign y8002 = ~n25074 ;
  assign y8003 = ~1'b0 ;
  assign y8004 = n25078 ;
  assign y8005 = n25079 ;
  assign y8006 = ~n25083 ;
  assign y8007 = n25085 ;
  assign y8008 = ~1'b0 ;
  assign y8009 = n25086 ;
  assign y8010 = n25088 ;
  assign y8011 = ~n25090 ;
  assign y8012 = ~1'b0 ;
  assign y8013 = ~n25094 ;
  assign y8014 = ~n25095 ;
  assign y8015 = ~n25103 ;
  assign y8016 = n25105 ;
  assign y8017 = ~n25108 ;
  assign y8018 = ~n25110 ;
  assign y8019 = ~n25112 ;
  assign y8020 = ~1'b0 ;
  assign y8021 = n25113 ;
  assign y8022 = ~1'b0 ;
  assign y8023 = n25114 ;
  assign y8024 = n25119 ;
  assign y8025 = n16148 ;
  assign y8026 = n25124 ;
  assign y8027 = ~1'b0 ;
  assign y8028 = ~n25128 ;
  assign y8029 = n25130 ;
  assign y8030 = ~n25134 ;
  assign y8031 = n25135 ;
  assign y8032 = n25137 ;
  assign y8033 = ~n25138 ;
  assign y8034 = ~1'b0 ;
  assign y8035 = ~1'b0 ;
  assign y8036 = ~1'b0 ;
  assign y8037 = ~n25139 ;
  assign y8038 = ~n25142 ;
  assign y8039 = ~n25145 ;
  assign y8040 = n25146 ;
  assign y8041 = ~n25150 ;
  assign y8042 = n25152 ;
  assign y8043 = ~1'b0 ;
  assign y8044 = ~n25153 ;
  assign y8045 = n25159 ;
  assign y8046 = ~1'b0 ;
  assign y8047 = n25163 ;
  assign y8048 = ~n16627 ;
  assign y8049 = n25166 ;
  assign y8050 = n25169 ;
  assign y8051 = ~n25172 ;
  assign y8052 = n25174 ;
  assign y8053 = ~n25177 ;
  assign y8054 = ~n25180 ;
  assign y8055 = ~n25182 ;
  assign y8056 = n25185 ;
  assign y8057 = ~n25186 ;
  assign y8058 = ~1'b0 ;
  assign y8059 = ~1'b0 ;
  assign y8060 = ~n25189 ;
  assign y8061 = ~1'b0 ;
  assign y8062 = ~n25190 ;
  assign y8063 = ~n25191 ;
  assign y8064 = n13012 ;
  assign y8065 = ~n25196 ;
  assign y8066 = n25205 ;
  assign y8067 = n25208 ;
  assign y8068 = ~n25211 ;
  assign y8069 = ~n25212 ;
  assign y8070 = ~n25214 ;
  assign y8071 = n25216 ;
  assign y8072 = n25219 ;
  assign y8073 = ~n25222 ;
  assign y8074 = n25223 ;
  assign y8075 = n25224 ;
  assign y8076 = ~n25225 ;
  assign y8077 = ~1'b0 ;
  assign y8078 = n25227 ;
  assign y8079 = ~1'b0 ;
  assign y8080 = n25228 ;
  assign y8081 = n25232 ;
  assign y8082 = n25235 ;
  assign y8083 = n25236 ;
  assign y8084 = ~n25237 ;
  assign y8085 = ~n25240 ;
  assign y8086 = ~1'b0 ;
  assign y8087 = n25243 ;
  assign y8088 = n25245 ;
  assign y8089 = ~n25246 ;
  assign y8090 = n25247 ;
  assign y8091 = ~n25252 ;
  assign y8092 = n25253 ;
  assign y8093 = n25254 ;
  assign y8094 = n25255 ;
  assign y8095 = ~1'b0 ;
  assign y8096 = ~n25258 ;
  assign y8097 = n25260 ;
  assign y8098 = n25264 ;
  assign y8099 = n25267 ;
  assign y8100 = n25270 ;
  assign y8101 = n25273 ;
  assign y8102 = n25274 ;
  assign y8103 = ~1'b0 ;
  assign y8104 = n25277 ;
  assign y8105 = ~n25278 ;
  assign y8106 = n25280 ;
  assign y8107 = ~n25282 ;
  assign y8108 = ~n25289 ;
  assign y8109 = n25290 ;
  assign y8110 = ~n25293 ;
  assign y8111 = ~n25295 ;
  assign y8112 = ~n25298 ;
  assign y8113 = ~n25301 ;
  assign y8114 = ~n25304 ;
  assign y8115 = n25305 ;
  assign y8116 = ~n25307 ;
  assign y8117 = ~n25313 ;
  assign y8118 = ~n25316 ;
  assign y8119 = ~1'b0 ;
  assign y8120 = ~1'b0 ;
  assign y8121 = ~n25317 ;
  assign y8122 = ~n25318 ;
  assign y8123 = ~1'b0 ;
  assign y8124 = n25320 ;
  assign y8125 = ~n25323 ;
  assign y8126 = ~n25329 ;
  assign y8127 = n25333 ;
  assign y8128 = ~n25334 ;
  assign y8129 = ~1'b0 ;
  assign y8130 = ~1'b0 ;
  assign y8131 = ~n25336 ;
  assign y8132 = ~n25337 ;
  assign y8133 = n25338 ;
  assign y8134 = n25344 ;
  assign y8135 = n25346 ;
  assign y8136 = ~n25347 ;
  assign y8137 = ~1'b0 ;
  assign y8138 = n25349 ;
  assign y8139 = ~1'b0 ;
  assign y8140 = ~n25353 ;
  assign y8141 = ~n25355 ;
  assign y8142 = ~n25357 ;
  assign y8143 = ~n25358 ;
  assign y8144 = ~n25359 ;
  assign y8145 = n25360 ;
  assign y8146 = n25362 ;
  assign y8147 = ~n25364 ;
  assign y8148 = ~n25366 ;
  assign y8149 = ~1'b0 ;
  assign y8150 = ~n25374 ;
  assign y8151 = ~n25375 ;
  assign y8152 = n25380 ;
  assign y8153 = n25381 ;
  assign y8154 = ~n25383 ;
  assign y8155 = 1'b0 ;
  assign y8156 = ~n3174 ;
  assign y8157 = n25387 ;
  assign y8158 = n25391 ;
  assign y8159 = n25393 ;
  assign y8160 = n25396 ;
  assign y8161 = ~n25397 ;
  assign y8162 = ~n25401 ;
  assign y8163 = n25404 ;
  assign y8164 = ~n25405 ;
  assign y8165 = ~n25408 ;
  assign y8166 = ~n25410 ;
  assign y8167 = n25412 ;
  assign y8168 = ~1'b0 ;
  assign y8169 = ~1'b0 ;
  assign y8170 = ~n25415 ;
  assign y8171 = n25417 ;
  assign y8172 = ~n25420 ;
  assign y8173 = ~n25424 ;
  assign y8174 = ~1'b0 ;
  assign y8175 = n25427 ;
  assign y8176 = n25429 ;
  assign y8177 = ~n25432 ;
  assign y8178 = ~n25433 ;
  assign y8179 = ~n25435 ;
  assign y8180 = n25438 ;
  assign y8181 = ~n25439 ;
  assign y8182 = n25442 ;
  assign y8183 = ~1'b0 ;
  assign y8184 = ~n25446 ;
  assign y8185 = n25447 ;
  assign y8186 = ~n25449 ;
  assign y8187 = n25451 ;
  assign y8188 = ~1'b0 ;
  assign y8189 = n25455 ;
  assign y8190 = n25456 ;
  assign y8191 = ~n25459 ;
  assign y8192 = ~n25460 ;
  assign y8193 = n10735 ;
  assign y8194 = ~n25462 ;
  assign y8195 = ~1'b0 ;
  assign y8196 = ~n25464 ;
  assign y8197 = n25470 ;
  assign y8198 = ~n25471 ;
  assign y8199 = n142 ;
  assign y8200 = ~n25472 ;
  assign y8201 = ~n25477 ;
  assign y8202 = n25479 ;
  assign y8203 = ~1'b0 ;
  assign y8204 = n25480 ;
  assign y8205 = ~n25481 ;
  assign y8206 = n25482 ;
  assign y8207 = ~n25483 ;
  assign y8208 = ~1'b0 ;
  assign y8209 = ~1'b0 ;
  assign y8210 = n25488 ;
  assign y8211 = ~n25490 ;
  assign y8212 = n25493 ;
  assign y8213 = n25497 ;
  assign y8214 = ~n25498 ;
  assign y8215 = n25502 ;
  assign y8216 = n25503 ;
  assign y8217 = ~1'b0 ;
  assign y8218 = n25505 ;
  assign y8219 = ~n25512 ;
  assign y8220 = ~n25515 ;
  assign y8221 = n25522 ;
  assign y8222 = ~n25525 ;
  assign y8223 = ~n25528 ;
  assign y8224 = ~n25531 ;
  assign y8225 = n6274 ;
  assign y8226 = ~n25533 ;
  assign y8227 = n25536 ;
  assign y8228 = ~1'b0 ;
  assign y8229 = n25537 ;
  assign y8230 = ~n25538 ;
  assign y8231 = ~n25540 ;
  assign y8232 = n25546 ;
  assign y8233 = n25547 ;
  assign y8234 = n25549 ;
  assign y8235 = ~1'b0 ;
  assign y8236 = n25555 ;
  assign y8237 = n25557 ;
  assign y8238 = n25559 ;
  assign y8239 = ~n25561 ;
  assign y8240 = n25565 ;
  assign y8241 = n25566 ;
  assign y8242 = ~n25567 ;
  assign y8243 = ~1'b0 ;
  assign y8244 = n25571 ;
  assign y8245 = ~n25573 ;
  assign y8246 = ~n25575 ;
  assign y8247 = ~n25576 ;
  assign y8248 = n25582 ;
  assign y8249 = n25583 ;
  assign y8250 = n25585 ;
  assign y8251 = n12306 ;
  assign y8252 = ~n25586 ;
  assign y8253 = ~n25595 ;
  assign y8254 = n25597 ;
  assign y8255 = ~n25598 ;
  assign y8256 = n25601 ;
  assign y8257 = n25606 ;
  assign y8258 = n25608 ;
  assign y8259 = n25614 ;
  assign y8260 = ~1'b0 ;
  assign y8261 = ~1'b0 ;
  assign y8262 = ~1'b0 ;
  assign y8263 = ~n25616 ;
  assign y8264 = n25617 ;
  assign y8265 = ~n25622 ;
  assign y8266 = n25625 ;
  assign y8267 = ~n25628 ;
  assign y8268 = ~n25629 ;
  assign y8269 = n25631 ;
  assign y8270 = n25634 ;
  assign y8271 = ~1'b0 ;
  assign y8272 = n25638 ;
  assign y8273 = n25640 ;
  assign y8274 = ~n25642 ;
  assign y8275 = ~n25647 ;
  assign y8276 = n25648 ;
  assign y8277 = n25651 ;
  assign y8278 = n25655 ;
  assign y8279 = ~n25658 ;
  assign y8280 = ~n25661 ;
  assign y8281 = ~n25665 ;
  assign y8282 = n25666 ;
  assign y8283 = n25669 ;
  assign y8284 = n25671 ;
  assign y8285 = ~n25673 ;
  assign y8286 = n25674 ;
  assign y8287 = n25675 ;
  assign y8288 = ~1'b0 ;
  assign y8289 = n25679 ;
  assign y8290 = ~1'b0 ;
  assign y8291 = ~n25682 ;
  assign y8292 = n25683 ;
  assign y8293 = ~n25687 ;
  assign y8294 = n25691 ;
  assign y8295 = ~n25692 ;
  assign y8296 = n5745 ;
  assign y8297 = n25694 ;
  assign y8298 = ~1'b0 ;
  assign y8299 = ~1'b0 ;
  assign y8300 = n25695 ;
  assign y8301 = ~n25700 ;
  assign y8302 = ~n25702 ;
  assign y8303 = n25703 ;
  assign y8304 = ~n25706 ;
  assign y8305 = n25708 ;
  assign y8306 = ~1'b0 ;
  assign y8307 = ~n25712 ;
  assign y8308 = ~n25714 ;
  assign y8309 = ~1'b0 ;
  assign y8310 = ~n25718 ;
  assign y8311 = n25720 ;
  assign y8312 = ~n25722 ;
  assign y8313 = ~n25723 ;
  assign y8314 = ~n25728 ;
  assign y8315 = n25732 ;
  assign y8316 = ~n25734 ;
  assign y8317 = n25738 ;
  assign y8318 = ~n25741 ;
  assign y8319 = n25749 ;
  assign y8320 = n25750 ;
  assign y8321 = n25752 ;
  assign y8322 = ~n25754 ;
  assign y8323 = n25756 ;
  assign y8324 = ~n25757 ;
  assign y8325 = ~n25760 ;
  assign y8326 = n25763 ;
  assign y8327 = n25765 ;
  assign y8328 = ~n25766 ;
  assign y8329 = ~n25767 ;
  assign y8330 = ~n25773 ;
  assign y8331 = ~n25775 ;
  assign y8332 = n25783 ;
  assign y8333 = n25788 ;
  assign y8334 = ~n25789 ;
  assign y8335 = ~n25790 ;
  assign y8336 = n25792 ;
  assign y8337 = n25793 ;
  assign y8338 = ~n25797 ;
  assign y8339 = ~n25804 ;
  assign y8340 = n25805 ;
  assign y8341 = ~1'b0 ;
  assign y8342 = ~n25809 ;
  assign y8343 = n25811 ;
  assign y8344 = ~n25812 ;
  assign y8345 = n25814 ;
  assign y8346 = n25818 ;
  assign y8347 = n25819 ;
  assign y8348 = n25820 ;
  assign y8349 = ~1'b0 ;
  assign y8350 = ~n25825 ;
  assign y8351 = n23004 ;
  assign y8352 = ~n25826 ;
  assign y8353 = n25828 ;
  assign y8354 = n25829 ;
  assign y8355 = n25832 ;
  assign y8356 = ~n25833 ;
  assign y8357 = n25837 ;
  assign y8358 = ~n25839 ;
  assign y8359 = ~1'b0 ;
  assign y8360 = n25841 ;
  assign y8361 = n25842 ;
  assign y8362 = ~n25845 ;
  assign y8363 = ~n25847 ;
  assign y8364 = ~n25851 ;
  assign y8365 = ~n25853 ;
  assign y8366 = ~n25855 ;
  assign y8367 = n25857 ;
  assign y8368 = n25859 ;
  assign y8369 = n25863 ;
  assign y8370 = ~n25865 ;
  assign y8371 = n25867 ;
  assign y8372 = n8354 ;
  assign y8373 = n25872 ;
  assign y8374 = ~1'b0 ;
  assign y8375 = ~n25875 ;
  assign y8376 = ~1'b0 ;
  assign y8377 = ~n25876 ;
  assign y8378 = n25877 ;
  assign y8379 = ~n25880 ;
  assign y8380 = n25881 ;
  assign y8381 = n25888 ;
  assign y8382 = n25892 ;
  assign y8383 = n25894 ;
  assign y8384 = ~n25895 ;
  assign y8385 = n25898 ;
  assign y8386 = n25899 ;
  assign y8387 = ~n25900 ;
  assign y8388 = n25902 ;
  assign y8389 = ~n25904 ;
  assign y8390 = ~n25905 ;
  assign y8391 = n25906 ;
  assign y8392 = ~n25910 ;
  assign y8393 = ~1'b0 ;
  assign y8394 = ~n25914 ;
  assign y8395 = n25917 ;
  assign y8396 = ~1'b0 ;
  assign y8397 = n25923 ;
  assign y8398 = ~n25924 ;
  assign y8399 = n25927 ;
  assign y8400 = ~n25936 ;
  assign y8401 = n25938 ;
  assign y8402 = ~1'b0 ;
  assign y8403 = ~1'b0 ;
  assign y8404 = ~n25940 ;
  assign y8405 = ~n25941 ;
  assign y8406 = n25950 ;
  assign y8407 = ~n25951 ;
  assign y8408 = n25952 ;
  assign y8409 = n25954 ;
  assign y8410 = n25956 ;
  assign y8411 = ~n25958 ;
  assign y8412 = n25959 ;
  assign y8413 = n25969 ;
  assign y8414 = n25972 ;
  assign y8415 = ~n25973 ;
  assign y8416 = n25974 ;
  assign y8417 = n25979 ;
  assign y8418 = n25982 ;
  assign y8419 = ~n25985 ;
  assign y8420 = n25987 ;
  assign y8421 = ~1'b0 ;
  assign y8422 = ~n25988 ;
  assign y8423 = ~1'b0 ;
  assign y8424 = ~1'b0 ;
  assign y8425 = n25989 ;
  assign y8426 = ~n25995 ;
  assign y8427 = ~n25998 ;
  assign y8428 = n26003 ;
  assign y8429 = ~n26008 ;
  assign y8430 = n26010 ;
  assign y8431 = ~1'b0 ;
  assign y8432 = ~n26011 ;
  assign y8433 = ~1'b0 ;
  assign y8434 = ~n26012 ;
  assign y8435 = ~n26013 ;
  assign y8436 = ~n26019 ;
  assign y8437 = n26024 ;
  assign y8438 = ~n26026 ;
  assign y8439 = ~n26028 ;
  assign y8440 = n26030 ;
  assign y8441 = n26034 ;
  assign y8442 = n26037 ;
  assign y8443 = ~n13984 ;
  assign y8444 = n26040 ;
  assign y8445 = ~n26044 ;
  assign y8446 = ~n26045 ;
  assign y8447 = n26046 ;
  assign y8448 = ~n26048 ;
  assign y8449 = ~n26049 ;
  assign y8450 = ~n26053 ;
  assign y8451 = n26057 ;
  assign y8452 = ~n26063 ;
  assign y8453 = ~n26064 ;
  assign y8454 = ~n26065 ;
  assign y8455 = ~n26068 ;
  assign y8456 = ~n26069 ;
  assign y8457 = ~1'b0 ;
  assign y8458 = n26076 ;
  assign y8459 = n26077 ;
  assign y8460 = ~n26078 ;
  assign y8461 = n26084 ;
  assign y8462 = ~n26085 ;
  assign y8463 = ~n26089 ;
  assign y8464 = n26090 ;
  assign y8465 = ~n26091 ;
  assign y8466 = ~n26093 ;
  assign y8467 = ~1'b0 ;
  assign y8468 = ~n26095 ;
  assign y8469 = ~1'b0 ;
  assign y8470 = ~n26096 ;
  assign y8471 = ~n26104 ;
  assign y8472 = ~n26105 ;
  assign y8473 = ~n26108 ;
  assign y8474 = n26109 ;
  assign y8475 = ~1'b0 ;
  assign y8476 = ~1'b0 ;
  assign y8477 = n26111 ;
  assign y8478 = n26112 ;
  assign y8479 = ~n26113 ;
  assign y8480 = n26121 ;
  assign y8481 = ~n26123 ;
  assign y8482 = ~n26129 ;
  assign y8483 = ~n26131 ;
  assign y8484 = ~n26133 ;
  assign y8485 = ~n26135 ;
  assign y8486 = ~1'b0 ;
  assign y8487 = ~n26141 ;
  assign y8488 = n26142 ;
  assign y8489 = n26143 ;
  assign y8490 = ~n24891 ;
  assign y8491 = n26151 ;
  assign y8492 = n26152 ;
  assign y8493 = ~n26153 ;
  assign y8494 = n26158 ;
  assign y8495 = ~n26162 ;
  assign y8496 = n26165 ;
  assign y8497 = n26171 ;
  assign y8498 = ~n26176 ;
  assign y8499 = ~n26179 ;
  assign y8500 = ~n26182 ;
  assign y8501 = n26185 ;
  assign y8502 = ~n26187 ;
  assign y8503 = ~n26191 ;
  assign y8504 = ~n26192 ;
  assign y8505 = n26195 ;
  assign y8506 = n26196 ;
  assign y8507 = ~1'b0 ;
  assign y8508 = ~1'b0 ;
  assign y8509 = n26197 ;
  assign y8510 = n26198 ;
  assign y8511 = ~n26199 ;
  assign y8512 = n26200 ;
  assign y8513 = n26202 ;
  assign y8514 = n26205 ;
  assign y8515 = n26207 ;
  assign y8516 = ~1'b0 ;
  assign y8517 = ~1'b0 ;
  assign y8518 = n26208 ;
  assign y8519 = ~n26215 ;
  assign y8520 = n26216 ;
  assign y8521 = ~n26218 ;
  assign y8522 = ~n26221 ;
  assign y8523 = n26228 ;
  assign y8524 = n26232 ;
  assign y8525 = ~1'b0 ;
  assign y8526 = ~1'b0 ;
  assign y8527 = ~1'b0 ;
  assign y8528 = n26233 ;
  assign y8529 = ~n26234 ;
  assign y8530 = n26236 ;
  assign y8531 = ~n26238 ;
  assign y8532 = n26240 ;
  assign y8533 = n26242 ;
  assign y8534 = ~n26245 ;
  assign y8535 = n26247 ;
  assign y8536 = n26249 ;
  assign y8537 = ~n26251 ;
  assign y8538 = n26252 ;
  assign y8539 = n26253 ;
  assign y8540 = ~n26256 ;
  assign y8541 = n26258 ;
  assign y8542 = n26264 ;
  assign y8543 = n26266 ;
  assign y8544 = ~n26268 ;
  assign y8545 = n26271 ;
  assign y8546 = n26272 ;
  assign y8547 = n26273 ;
  assign y8548 = ~n26275 ;
  assign y8549 = ~1'b0 ;
  assign y8550 = n26277 ;
  assign y8551 = ~1'b0 ;
  assign y8552 = ~n26279 ;
  assign y8553 = n26282 ;
  assign y8554 = n26284 ;
  assign y8555 = n26287 ;
  assign y8556 = ~n26290 ;
  assign y8557 = n26291 ;
  assign y8558 = n26294 ;
  assign y8559 = ~1'b0 ;
  assign y8560 = n26295 ;
  assign y8561 = n26296 ;
  assign y8562 = ~n26297 ;
  assign y8563 = n26298 ;
  assign y8564 = ~n26302 ;
  assign y8565 = ~1'b0 ;
  assign y8566 = ~n26305 ;
  assign y8567 = ~n26306 ;
  assign y8568 = ~n26308 ;
  assign y8569 = ~n26312 ;
  assign y8570 = n26313 ;
  assign y8571 = ~n26315 ;
  assign y8572 = n26316 ;
  assign y8573 = ~1'b0 ;
  assign y8574 = ~1'b0 ;
  assign y8575 = 1'b0 ;
  assign y8576 = n26319 ;
  assign y8577 = ~1'b0 ;
  assign y8578 = n26325 ;
  assign y8579 = n26327 ;
  assign y8580 = n26328 ;
  assign y8581 = ~n26330 ;
  assign y8582 = ~1'b0 ;
  assign y8583 = ~n26332 ;
  assign y8584 = ~n26336 ;
  assign y8585 = n26338 ;
  assign y8586 = ~n26340 ;
  assign y8587 = n26342 ;
  assign y8588 = ~n26346 ;
  assign y8589 = n26352 ;
  assign y8590 = ~n26357 ;
  assign y8591 = n26358 ;
  assign y8592 = n23326 ;
  assign y8593 = ~n26371 ;
  assign y8594 = ~n26372 ;
  assign y8595 = n26375 ;
  assign y8596 = ~1'b0 ;
  assign y8597 = ~1'b0 ;
  assign y8598 = n26377 ;
  assign y8599 = n26378 ;
  assign y8600 = n26380 ;
  assign y8601 = n26381 ;
  assign y8602 = ~n26383 ;
  assign y8603 = ~n26384 ;
  assign y8604 = n26385 ;
  assign y8605 = ~1'b0 ;
  assign y8606 = n26393 ;
  assign y8607 = n26399 ;
  assign y8608 = ~n26402 ;
  assign y8609 = ~n26407 ;
  assign y8610 = ~n26409 ;
  assign y8611 = ~n26414 ;
  assign y8612 = n26420 ;
  assign y8613 = ~n26422 ;
  assign y8614 = ~n26424 ;
  assign y8615 = ~n26427 ;
  assign y8616 = ~1'b0 ;
  assign y8617 = n26429 ;
  assign y8618 = ~n26431 ;
  assign y8619 = n26432 ;
  assign y8620 = n26433 ;
  assign y8621 = ~n26434 ;
  assign y8622 = ~n26438 ;
  assign y8623 = n26441 ;
  assign y8624 = ~n26442 ;
  assign y8625 = ~1'b0 ;
  assign y8626 = ~1'b0 ;
  assign y8627 = ~n26446 ;
  assign y8628 = ~n26449 ;
  assign y8629 = n26456 ;
  assign y8630 = n26460 ;
  assign y8631 = n26464 ;
  assign y8632 = n26466 ;
  assign y8633 = ~n26470 ;
  assign y8634 = ~n26471 ;
  assign y8635 = ~n26474 ;
  assign y8636 = ~1'b0 ;
  assign y8637 = n26475 ;
  assign y8638 = ~n26476 ;
  assign y8639 = ~n26479 ;
  assign y8640 = ~n26480 ;
  assign y8641 = n26486 ;
  assign y8642 = ~1'b0 ;
  assign y8643 = ~n26487 ;
  assign y8644 = ~n26492 ;
  assign y8645 = n26494 ;
  assign y8646 = ~n26498 ;
  assign y8647 = ~n26499 ;
  assign y8648 = ~n23552 ;
  assign y8649 = n26501 ;
  assign y8650 = ~1'b0 ;
  assign y8651 = ~1'b0 ;
  assign y8652 = ~1'b0 ;
  assign y8653 = ~1'b0 ;
  assign y8654 = ~n26503 ;
  assign y8655 = n26504 ;
  assign y8656 = ~n26505 ;
  assign y8657 = ~n26508 ;
  assign y8658 = n26509 ;
  assign y8659 = ~n26510 ;
  assign y8660 = ~n26513 ;
  assign y8661 = n26516 ;
  assign y8662 = ~1'b0 ;
  assign y8663 = ~n26517 ;
  assign y8664 = ~n26518 ;
  assign y8665 = ~n26519 ;
  assign y8666 = ~n26521 ;
  assign y8667 = ~n26524 ;
  assign y8668 = ~1'b0 ;
  assign y8669 = ~1'b0 ;
  assign y8670 = ~n26525 ;
  assign y8671 = n26526 ;
  assign y8672 = ~n18196 ;
  assign y8673 = ~n26527 ;
  assign y8674 = n26532 ;
  assign y8675 = n26533 ;
  assign y8676 = ~n26539 ;
  assign y8677 = ~n2754 ;
  assign y8678 = n26552 ;
  assign y8679 = ~n26553 ;
  assign y8680 = n10884 ;
  assign y8681 = n26554 ;
  assign y8682 = ~n26560 ;
  assign y8683 = ~1'b0 ;
  assign y8684 = n26561 ;
  assign y8685 = ~n26563 ;
  assign y8686 = ~1'b0 ;
  assign y8687 = ~1'b0 ;
  assign y8688 = n26564 ;
  assign y8689 = ~n26566 ;
  assign y8690 = ~1'b0 ;
  assign y8691 = ~n26570 ;
  assign y8692 = n26572 ;
  assign y8693 = n26574 ;
  assign y8694 = n26577 ;
  assign y8695 = n26579 ;
  assign y8696 = n26581 ;
  assign y8697 = ~n26588 ;
  assign y8698 = n26589 ;
  assign y8699 = n26592 ;
  assign y8700 = ~n26593 ;
  assign y8701 = ~n26594 ;
  assign y8702 = ~1'b0 ;
  assign y8703 = ~1'b0 ;
  assign y8704 = ~n26595 ;
  assign y8705 = ~1'b0 ;
  assign y8706 = n26596 ;
  assign y8707 = ~n26597 ;
  assign y8708 = ~n26598 ;
  assign y8709 = n26599 ;
  assign y8710 = n26604 ;
  assign y8711 = ~n26605 ;
  assign y8712 = ~1'b0 ;
  assign y8713 = ~1'b0 ;
  assign y8714 = ~n26609 ;
  assign y8715 = n26611 ;
  assign y8716 = ~n26613 ;
  assign y8717 = ~n20987 ;
  assign y8718 = n26616 ;
  assign y8719 = n26618 ;
  assign y8720 = ~1'b0 ;
  assign y8721 = ~1'b0 ;
  assign y8722 = ~n26619 ;
  assign y8723 = n26622 ;
  assign y8724 = ~n26624 ;
  assign y8725 = ~n26626 ;
  assign y8726 = n26627 ;
  assign y8727 = ~n26628 ;
  assign y8728 = ~n26631 ;
  assign y8729 = ~1'b0 ;
  assign y8730 = n26633 ;
  assign y8731 = n26635 ;
  assign y8732 = ~1'b0 ;
  assign y8733 = n26638 ;
  assign y8734 = n26639 ;
  assign y8735 = ~n26641 ;
  assign y8736 = ~1'b0 ;
  assign y8737 = n26642 ;
  assign y8738 = n26645 ;
  assign y8739 = n26649 ;
  assign y8740 = ~n26652 ;
  assign y8741 = n26653 ;
  assign y8742 = ~n26654 ;
  assign y8743 = n26658 ;
  assign y8744 = n26662 ;
  assign y8745 = ~n26664 ;
  assign y8746 = n26667 ;
  assign y8747 = n26670 ;
  assign y8748 = ~n26672 ;
  assign y8749 = ~n26675 ;
  assign y8750 = ~n26679 ;
  assign y8751 = ~n26680 ;
  assign y8752 = n26685 ;
  assign y8753 = ~n26689 ;
  assign y8754 = ~1'b0 ;
  assign y8755 = n26691 ;
  assign y8756 = ~1'b0 ;
  assign y8757 = n26693 ;
  assign y8758 = n26695 ;
  assign y8759 = ~n26696 ;
  assign y8760 = n26701 ;
  assign y8761 = n26704 ;
  assign y8762 = ~n26707 ;
  assign y8763 = ~n26708 ;
  assign y8764 = ~n26711 ;
  assign y8765 = ~n26714 ;
  assign y8766 = ~1'b0 ;
  assign y8767 = ~n26715 ;
  assign y8768 = n26716 ;
  assign y8769 = n26723 ;
  assign y8770 = ~n26724 ;
  assign y8771 = ~1'b0 ;
  assign y8772 = ~n26725 ;
  assign y8773 = n26732 ;
  assign y8774 = n26733 ;
  assign y8775 = ~n26734 ;
  assign y8776 = ~n26743 ;
  assign y8777 = ~n26744 ;
  assign y8778 = ~n26750 ;
  assign y8779 = n26752 ;
  assign y8780 = ~n26755 ;
  assign y8781 = ~1'b0 ;
  assign y8782 = n26767 ;
  assign y8783 = n26768 ;
  assign y8784 = n26771 ;
  assign y8785 = n26772 ;
  assign y8786 = n26776 ;
  assign y8787 = n26780 ;
  assign y8788 = n26781 ;
  assign y8789 = ~n26783 ;
  assign y8790 = ~n26785 ;
  assign y8791 = ~n26793 ;
  assign y8792 = n26798 ;
  assign y8793 = n26800 ;
  assign y8794 = ~n26807 ;
  assign y8795 = n26809 ;
  assign y8796 = ~n26815 ;
  assign y8797 = ~n26818 ;
  assign y8798 = ~n26822 ;
  assign y8799 = ~1'b0 ;
  assign y8800 = ~n26824 ;
  assign y8801 = ~1'b0 ;
  assign y8802 = ~1'b0 ;
  assign y8803 = ~1'b0 ;
  assign y8804 = n26825 ;
  assign y8805 = ~n26831 ;
  assign y8806 = n26838 ;
  assign y8807 = ~1'b0 ;
  assign y8808 = ~1'b0 ;
  assign y8809 = n26841 ;
  assign y8810 = n26842 ;
  assign y8811 = ~1'b0 ;
  assign y8812 = ~n26844 ;
  assign y8813 = ~n26845 ;
  assign y8814 = ~n26847 ;
  assign y8815 = ~n26848 ;
  assign y8816 = ~n26853 ;
  assign y8817 = ~n26857 ;
  assign y8818 = n26859 ;
  assign y8819 = n26860 ;
  assign y8820 = ~n26864 ;
  assign y8821 = n26869 ;
  assign y8822 = ~n26870 ;
  assign y8823 = ~n26874 ;
  assign y8824 = ~n26884 ;
  assign y8825 = n26888 ;
  assign y8826 = ~n26889 ;
  assign y8827 = n26890 ;
  assign y8828 = ~n26892 ;
  assign y8829 = ~n26895 ;
  assign y8830 = ~n26900 ;
  assign y8831 = ~n26903 ;
  assign y8832 = n26907 ;
  assign y8833 = ~1'b0 ;
  assign y8834 = n26909 ;
  assign y8835 = ~n26912 ;
  assign y8836 = n26914 ;
  assign y8837 = n13830 ;
  assign y8838 = n26915 ;
  assign y8839 = ~n26920 ;
  assign y8840 = n26922 ;
  assign y8841 = ~1'b0 ;
  assign y8842 = ~1'b0 ;
  assign y8843 = ~n26924 ;
  assign y8844 = ~1'b0 ;
  assign y8845 = n26928 ;
  assign y8846 = n26929 ;
  assign y8847 = ~n26930 ;
  assign y8848 = ~n26935 ;
  assign y8849 = ~n26938 ;
  assign y8850 = n26941 ;
  assign y8851 = n26942 ;
  assign y8852 = ~1'b0 ;
  assign y8853 = n9236 ;
  assign y8854 = ~1'b0 ;
  assign y8855 = ~n26946 ;
  assign y8856 = ~n26948 ;
  assign y8857 = n26951 ;
  assign y8858 = ~n26958 ;
  assign y8859 = ~n26964 ;
  assign y8860 = ~n26965 ;
  assign y8861 = ~n26967 ;
  assign y8862 = ~1'b0 ;
  assign y8863 = ~1'b0 ;
  assign y8864 = ~n26970 ;
  assign y8865 = ~n26972 ;
  assign y8866 = ~n26973 ;
  assign y8867 = n26976 ;
  assign y8868 = n26984 ;
  assign y8869 = n26990 ;
  assign y8870 = ~1'b0 ;
  assign y8871 = n26995 ;
  assign y8872 = n26997 ;
  assign y8873 = ~n27001 ;
  assign y8874 = n27002 ;
  assign y8875 = ~n27006 ;
  assign y8876 = ~n27007 ;
  assign y8877 = ~n27010 ;
  assign y8878 = ~n27015 ;
  assign y8879 = n27021 ;
  assign y8880 = n27025 ;
  assign y8881 = n27027 ;
  assign y8882 = ~n27030 ;
  assign y8883 = n27034 ;
  assign y8884 = n27037 ;
  assign y8885 = n27038 ;
  assign y8886 = n27041 ;
  assign y8887 = n27042 ;
  assign y8888 = ~n27044 ;
  assign y8889 = n27045 ;
  assign y8890 = ~1'b0 ;
  assign y8891 = n27049 ;
  assign y8892 = ~1'b0 ;
  assign y8893 = n27053 ;
  assign y8894 = n27055 ;
  assign y8895 = ~n27056 ;
  assign y8896 = n27057 ;
  assign y8897 = ~n27061 ;
  assign y8898 = ~n16760 ;
  assign y8899 = ~n27063 ;
  assign y8900 = ~n27067 ;
  assign y8901 = ~n27071 ;
  assign y8902 = n27072 ;
  assign y8903 = ~n27074 ;
  assign y8904 = ~n27077 ;
  assign y8905 = n27083 ;
  assign y8906 = ~n27085 ;
  assign y8907 = n27089 ;
  assign y8908 = ~n27090 ;
  assign y8909 = n27094 ;
  assign y8910 = ~n27098 ;
  assign y8911 = n27102 ;
  assign y8912 = ~n27104 ;
  assign y8913 = ~1'b0 ;
  assign y8914 = ~1'b0 ;
  assign y8915 = n27107 ;
  assign y8916 = ~n27108 ;
  assign y8917 = ~n27113 ;
  assign y8918 = ~n27119 ;
  assign y8919 = n27120 ;
  assign y8920 = n27123 ;
  assign y8921 = ~n27126 ;
  assign y8922 = ~n27131 ;
  assign y8923 = ~1'b0 ;
  assign y8924 = ~1'b0 ;
  assign y8925 = n27138 ;
  assign y8926 = n27143 ;
  assign y8927 = n12426 ;
  assign y8928 = ~n27146 ;
  assign y8929 = n27147 ;
  assign y8930 = ~n27150 ;
  assign y8931 = ~n27152 ;
  assign y8932 = ~n27153 ;
  assign y8933 = ~1'b0 ;
  assign y8934 = n27156 ;
  assign y8935 = ~n27157 ;
  assign y8936 = n27158 ;
  assign y8937 = ~n27161 ;
  assign y8938 = ~n27163 ;
  assign y8939 = n27166 ;
  assign y8940 = ~n27168 ;
  assign y8941 = n27182 ;
  assign y8942 = ~n27184 ;
  assign y8943 = ~1'b0 ;
  assign y8944 = n27187 ;
  assign y8945 = ~n27188 ;
  assign y8946 = ~n27192 ;
  assign y8947 = n27196 ;
  assign y8948 = n27198 ;
  assign y8949 = n27200 ;
  assign y8950 = ~n27201 ;
  assign y8951 = n27202 ;
  assign y8952 = n27208 ;
  assign y8953 = ~1'b0 ;
  assign y8954 = ~n27212 ;
  assign y8955 = ~n27214 ;
  assign y8956 = ~n27215 ;
  assign y8957 = n27216 ;
  assign y8958 = n27222 ;
  assign y8959 = ~n27223 ;
  assign y8960 = ~n27226 ;
  assign y8961 = ~n27231 ;
  assign y8962 = n27234 ;
  assign y8963 = ~1'b0 ;
  assign y8964 = n27237 ;
  assign y8965 = ~n27242 ;
  assign y8966 = ~n27245 ;
  assign y8967 = ~n27249 ;
  assign y8968 = n27251 ;
  assign y8969 = ~n27252 ;
  assign y8970 = n27253 ;
  assign y8971 = ~n27258 ;
  assign y8972 = n27260 ;
  assign y8973 = ~n27262 ;
  assign y8974 = n27264 ;
  assign y8975 = n27265 ;
  assign y8976 = n27267 ;
  assign y8977 = n27268 ;
  assign y8978 = ~n27272 ;
  assign y8979 = ~n27273 ;
  assign y8980 = ~1'b0 ;
  assign y8981 = n27275 ;
  assign y8982 = ~1'b0 ;
  assign y8983 = ~1'b0 ;
  assign y8984 = ~n27276 ;
  assign y8985 = n27277 ;
  assign y8986 = ~n27278 ;
  assign y8987 = n27281 ;
  assign y8988 = n27282 ;
  assign y8989 = ~n27286 ;
  assign y8990 = ~n27288 ;
  assign y8991 = ~n27291 ;
  assign y8992 = ~1'b0 ;
  assign y8993 = ~1'b0 ;
  assign y8994 = ~1'b0 ;
  assign y8995 = ~n27292 ;
  assign y8996 = ~1'b0 ;
  assign y8997 = n27294 ;
  assign y8998 = ~n27295 ;
  assign y8999 = ~n3941 ;
  assign y9000 = ~1'b0 ;
  assign y9001 = ~1'b0 ;
  assign y9002 = ~n27297 ;
  assign y9003 = n27302 ;
  assign y9004 = n27307 ;
  assign y9005 = n27310 ;
  assign y9006 = ~n27314 ;
  assign y9007 = ~n27318 ;
  assign y9008 = n27319 ;
  assign y9009 = ~n27326 ;
  assign y9010 = ~n27330 ;
  assign y9011 = ~1'b0 ;
  assign y9012 = ~1'b0 ;
  assign y9013 = n27332 ;
  assign y9014 = ~n27333 ;
  assign y9015 = n27336 ;
  assign y9016 = ~n27338 ;
  assign y9017 = n27339 ;
  assign y9018 = n27340 ;
  assign y9019 = ~n27345 ;
  assign y9020 = ~1'b0 ;
  assign y9021 = ~n27347 ;
  assign y9022 = n27352 ;
  assign y9023 = 1'b0 ;
  assign y9024 = ~n27356 ;
  assign y9025 = n27357 ;
  assign y9026 = ~n27358 ;
  assign y9027 = n27360 ;
  assign y9028 = n27362 ;
  assign y9029 = ~n27364 ;
  assign y9030 = ~1'b0 ;
  assign y9031 = ~n27368 ;
  assign y9032 = n27370 ;
  assign y9033 = ~n27371 ;
  assign y9034 = ~n27374 ;
  assign y9035 = n27375 ;
  assign y9036 = ~1'b0 ;
  assign y9037 = ~1'b0 ;
  assign y9038 = n27376 ;
  assign y9039 = ~1'b0 ;
  assign y9040 = n27379 ;
  assign y9041 = n27381 ;
  assign y9042 = ~n27382 ;
  assign y9043 = ~n16880 ;
  assign y9044 = n27383 ;
  assign y9045 = n27385 ;
  assign y9046 = ~n27389 ;
  assign y9047 = ~n27390 ;
  assign y9048 = ~n27391 ;
  assign y9049 = n23818 ;
  assign y9050 = ~n27393 ;
  assign y9051 = ~n27396 ;
  assign y9052 = ~n27397 ;
  assign y9053 = ~n27403 ;
  assign y9054 = ~1'b0 ;
  assign y9055 = ~1'b0 ;
  assign y9056 = ~1'b0 ;
  assign y9057 = n27405 ;
  assign y9058 = ~n27406 ;
  assign y9059 = n27409 ;
  assign y9060 = ~n27413 ;
  assign y9061 = ~n27416 ;
  assign y9062 = n27417 ;
  assign y9063 = ~n27418 ;
  assign y9064 = ~1'b0 ;
  assign y9065 = n27420 ;
  assign y9066 = 1'b0 ;
  assign y9067 = ~n27421 ;
  assign y9068 = ~n27430 ;
  assign y9069 = ~n27435 ;
  assign y9070 = ~n27440 ;
  assign y9071 = ~n27443 ;
  assign y9072 = n27444 ;
  assign y9073 = ~n27446 ;
  assign y9074 = n27455 ;
  assign y9075 = n27459 ;
  assign y9076 = ~n27461 ;
  assign y9077 = ~n27462 ;
  assign y9078 = ~n27466 ;
  assign y9079 = n27472 ;
  assign y9080 = ~n27481 ;
  assign y9081 = n27485 ;
  assign y9082 = n27486 ;
  assign y9083 = ~n27493 ;
  assign y9084 = n27496 ;
  assign y9085 = ~n27500 ;
  assign y9086 = ~n27506 ;
  assign y9087 = ~n27511 ;
  assign y9088 = ~n27512 ;
  assign y9089 = n27517 ;
  assign y9090 = ~n27518 ;
  assign y9091 = n27521 ;
  assign y9092 = n27524 ;
  assign y9093 = ~1'b0 ;
  assign y9094 = n27525 ;
  assign y9095 = ~1'b0 ;
  assign y9096 = ~n27526 ;
  assign y9097 = n27527 ;
  assign y9098 = n27528 ;
  assign y9099 = n27529 ;
  assign y9100 = ~1'b0 ;
  assign y9101 = ~1'b0 ;
  assign y9102 = ~n27531 ;
  assign y9103 = ~1'b0 ;
  assign y9104 = n27534 ;
  assign y9105 = n27536 ;
  assign y9106 = n27541 ;
  assign y9107 = n27542 ;
  assign y9108 = n27543 ;
  assign y9109 = ~n27548 ;
  assign y9110 = ~n27553 ;
  assign y9111 = ~n27555 ;
  assign y9112 = n16259 ;
  assign y9113 = ~n27561 ;
  assign y9114 = n27563 ;
  assign y9115 = ~n27576 ;
  assign y9116 = ~n27577 ;
  assign y9117 = ~n27579 ;
  assign y9118 = n17766 ;
  assign y9119 = ~n27583 ;
  assign y9120 = ~n27588 ;
  assign y9121 = n27591 ;
  assign y9122 = n27593 ;
  assign y9123 = ~n14573 ;
  assign y9124 = n27595 ;
  assign y9125 = ~n27597 ;
  assign y9126 = n27598 ;
  assign y9127 = ~n27601 ;
  assign y9128 = ~n27602 ;
  assign y9129 = ~n27603 ;
  assign y9130 = ~n27604 ;
  assign y9131 = ~n27606 ;
  assign y9132 = ~n27610 ;
  assign y9133 = n4452 ;
  assign y9134 = ~1'b0 ;
  assign y9135 = n27615 ;
  assign y9136 = ~n27618 ;
  assign y9137 = ~n27624 ;
  assign y9138 = ~n27632 ;
  assign y9139 = n27633 ;
  assign y9140 = ~n27637 ;
  assign y9141 = ~1'b0 ;
  assign y9142 = ~n27639 ;
  assign y9143 = ~n27640 ;
  assign y9144 = n27643 ;
  assign y9145 = n27645 ;
  assign y9146 = ~n27646 ;
  assign y9147 = n27648 ;
  assign y9148 = ~n27651 ;
  assign y9149 = ~n27652 ;
  assign y9150 = ~n27654 ;
  assign y9151 = ~n27658 ;
  assign y9152 = ~1'b0 ;
  assign y9153 = n27659 ;
  assign y9154 = ~n27661 ;
  assign y9155 = ~n27662 ;
  assign y9156 = ~n27663 ;
  assign y9157 = ~n27664 ;
  assign y9158 = n27667 ;
  assign y9159 = ~n27670 ;
  assign y9160 = n27672 ;
  assign y9161 = ~n27673 ;
  assign y9162 = ~1'b0 ;
  assign y9163 = ~n27675 ;
  assign y9164 = n27677 ;
  assign y9165 = ~1'b0 ;
  assign y9166 = ~n27680 ;
  assign y9167 = ~n27681 ;
  assign y9168 = ~n27686 ;
  assign y9169 = n27687 ;
  assign y9170 = n27689 ;
  assign y9171 = ~n27692 ;
  assign y9172 = ~1'b0 ;
  assign y9173 = n27693 ;
  assign y9174 = ~n27694 ;
  assign y9175 = ~n27695 ;
  assign y9176 = n27696 ;
  assign y9177 = ~n27699 ;
  assign y9178 = n3360 ;
  assign y9179 = ~n27701 ;
  assign y9180 = ~1'b0 ;
  assign y9181 = ~1'b0 ;
  assign y9182 = n27704 ;
  assign y9183 = n27705 ;
  assign y9184 = ~n27706 ;
  assign y9185 = n27707 ;
  assign y9186 = ~n27708 ;
  assign y9187 = n27709 ;
  assign y9188 = ~n27713 ;
  assign y9189 = n27715 ;
  assign y9190 = ~n27718 ;
  assign y9191 = ~1'b0 ;
  assign y9192 = n27721 ;
  assign y9193 = n27726 ;
  assign y9194 = n27729 ;
  assign y9195 = n27731 ;
  assign y9196 = ~n27732 ;
  assign y9197 = ~n4070 ;
  assign y9198 = ~n27738 ;
  assign y9199 = n27740 ;
  assign y9200 = ~n27742 ;
  assign y9201 = ~n27744 ;
  assign y9202 = n27745 ;
  assign y9203 = n27746 ;
  assign y9204 = n27747 ;
  assign y9205 = ~n27750 ;
  assign y9206 = ~n27754 ;
  assign y9207 = n27758 ;
  assign y9208 = ~n27760 ;
  assign y9209 = ~1'b0 ;
  assign y9210 = ~n27766 ;
  assign y9211 = ~n27768 ;
  assign y9212 = ~n27769 ;
  assign y9213 = n9058 ;
  assign y9214 = n6800 ;
  assign y9215 = n27777 ;
  assign y9216 = ~n27780 ;
  assign y9217 = ~n27787 ;
  assign y9218 = ~n27791 ;
  assign y9219 = ~n27793 ;
  assign y9220 = n27794 ;
  assign y9221 = ~1'b0 ;
  assign y9222 = n27798 ;
  assign y9223 = n27801 ;
  assign y9224 = ~n27802 ;
  assign y9225 = ~n27804 ;
  assign y9226 = ~n27805 ;
  assign y9227 = ~n26161 ;
  assign y9228 = ~n27807 ;
  assign y9229 = ~n27810 ;
  assign y9230 = ~n27812 ;
  assign y9231 = ~n27813 ;
  assign y9232 = ~n27816 ;
  assign y9233 = ~n27818 ;
  assign y9234 = n25915 ;
  assign y9235 = ~n27819 ;
  assign y9236 = n27820 ;
  assign y9237 = ~n27822 ;
  assign y9238 = ~1'b0 ;
  assign y9239 = ~1'b0 ;
  assign y9240 = ~1'b0 ;
  assign y9241 = ~n27823 ;
  assign y9242 = ~n27831 ;
  assign y9243 = n27833 ;
  assign y9244 = n27834 ;
  assign y9245 = n27835 ;
  assign y9246 = n27844 ;
  assign y9247 = ~1'b0 ;
  assign y9248 = ~1'b0 ;
  assign y9249 = ~n27845 ;
  assign y9250 = ~n27846 ;
  assign y9251 = ~n27848 ;
  assign y9252 = n27849 ;
  assign y9253 = n27853 ;
  assign y9254 = ~n27854 ;
  assign y9255 = n27856 ;
  assign y9256 = ~n27858 ;
  assign y9257 = n27859 ;
  assign y9258 = n27863 ;
  assign y9259 = ~n27864 ;
  assign y9260 = n27867 ;
  assign y9261 = ~n27873 ;
  assign y9262 = ~n27878 ;
  assign y9263 = ~n27890 ;
  assign y9264 = ~n27892 ;
  assign y9265 = ~n18427 ;
  assign y9266 = ~n27894 ;
  assign y9267 = n27896 ;
  assign y9268 = n27897 ;
  assign y9269 = ~n27898 ;
  assign y9270 = n27900 ;
  assign y9271 = ~n27903 ;
  assign y9272 = ~n27905 ;
  assign y9273 = n27906 ;
  assign y9274 = n27911 ;
  assign y9275 = ~n27914 ;
  assign y9276 = n27915 ;
  assign y9277 = ~n27919 ;
  assign y9278 = ~n27921 ;
  assign y9279 = n27923 ;
  assign y9280 = ~n27925 ;
  assign y9281 = ~n27927 ;
  assign y9282 = n27929 ;
  assign y9283 = ~n27932 ;
  assign y9284 = ~n27934 ;
  assign y9285 = ~n27937 ;
  assign y9286 = n27939 ;
  assign y9287 = ~n10515 ;
  assign y9288 = ~n27940 ;
  assign y9289 = ~n27942 ;
  assign y9290 = ~n27946 ;
  assign y9291 = n27949 ;
  assign y9292 = ~n27952 ;
  assign y9293 = ~n27954 ;
  assign y9294 = ~n27956 ;
  assign y9295 = ~1'b0 ;
  assign y9296 = n27959 ;
  assign y9297 = ~n27962 ;
  assign y9298 = n27964 ;
  assign y9299 = ~n27970 ;
  assign y9300 = n27971 ;
  assign y9301 = ~n27972 ;
  assign y9302 = ~1'b0 ;
  assign y9303 = ~1'b0 ;
  assign y9304 = n27975 ;
  assign y9305 = n27977 ;
  assign y9306 = n8144 ;
  assign y9307 = n27982 ;
  assign y9308 = ~n27984 ;
  assign y9309 = ~n27988 ;
  assign y9310 = n27991 ;
  assign y9311 = ~n27994 ;
  assign y9312 = ~n27996 ;
  assign y9313 = n27998 ;
  assign y9314 = ~1'b0 ;
  assign y9315 = ~n27999 ;
  assign y9316 = n28000 ;
  assign y9317 = n28007 ;
  assign y9318 = n28008 ;
  assign y9319 = ~n28009 ;
  assign y9320 = 1'b0 ;
  assign y9321 = ~n9877 ;
  assign y9322 = ~n28010 ;
  assign y9323 = ~n28011 ;
  assign y9324 = ~1'b0 ;
  assign y9325 = n28017 ;
  assign y9326 = n28021 ;
  assign y9327 = ~n28027 ;
  assign y9328 = ~n28033 ;
  assign y9329 = n28035 ;
  assign y9330 = n28037 ;
  assign y9331 = ~n28038 ;
  assign y9332 = ~n28042 ;
  assign y9333 = n28043 ;
  assign y9334 = n28047 ;
  assign y9335 = n28048 ;
  assign y9336 = n28050 ;
  assign y9337 = n28054 ;
  assign y9338 = n28057 ;
  assign y9339 = ~n28059 ;
  assign y9340 = n28063 ;
  assign y9341 = ~1'b0 ;
  assign y9342 = ~n28065 ;
  assign y9343 = ~n28067 ;
  assign y9344 = ~1'b0 ;
  assign y9345 = ~n28068 ;
  assign y9346 = ~n28069 ;
  assign y9347 = ~n28070 ;
  assign y9348 = ~n28071 ;
  assign y9349 = n28074 ;
  assign y9350 = n28080 ;
  assign y9351 = ~n28085 ;
  assign y9352 = n28090 ;
  assign y9353 = n28095 ;
  assign y9354 = n28097 ;
  assign y9355 = ~n28098 ;
  assign y9356 = n28099 ;
  assign y9357 = ~n28101 ;
  assign y9358 = ~n28103 ;
  assign y9359 = ~1'b0 ;
  assign y9360 = ~n28104 ;
  assign y9361 = ~1'b0 ;
  assign y9362 = ~n28105 ;
  assign y9363 = n28115 ;
  assign y9364 = ~n28117 ;
  assign y9365 = n28118 ;
  assign y9366 = n28120 ;
  assign y9367 = n28122 ;
  assign y9368 = ~1'b0 ;
  assign y9369 = ~n28124 ;
  assign y9370 = n28126 ;
  assign y9371 = ~n28127 ;
  assign y9372 = ~n28130 ;
  assign y9373 = n28131 ;
  assign y9374 = ~n28135 ;
  assign y9375 = n28136 ;
  assign y9376 = n28137 ;
  assign y9377 = ~1'b0 ;
  assign y9378 = n28140 ;
  assign y9379 = ~1'b0 ;
  assign y9380 = ~n28142 ;
  assign y9381 = ~n28143 ;
  assign y9382 = n28146 ;
  assign y9383 = n28147 ;
  assign y9384 = n28148 ;
  assign y9385 = ~n28154 ;
  assign y9386 = n28156 ;
  assign y9387 = n28158 ;
  assign y9388 = n28164 ;
  assign y9389 = n28166 ;
  assign y9390 = ~n28170 ;
  assign y9391 = n28173 ;
  assign y9392 = ~n28174 ;
  assign y9393 = ~n28176 ;
  assign y9394 = n28177 ;
  assign y9395 = n28179 ;
  assign y9396 = ~1'b0 ;
  assign y9397 = ~n28181 ;
  assign y9398 = ~1'b0 ;
  assign y9399 = ~n28182 ;
  assign y9400 = ~1'b0 ;
  assign y9401 = n28186 ;
  assign y9402 = ~n28187 ;
  assign y9403 = ~n28188 ;
  assign y9404 = n28194 ;
  assign y9405 = n28197 ;
  assign y9406 = n28202 ;
  assign y9407 = n28203 ;
  assign y9408 = ~n28204 ;
  assign y9409 = ~n28208 ;
  assign y9410 = ~n28213 ;
  assign y9411 = ~1'b0 ;
  assign y9412 = n28218 ;
  assign y9413 = ~n28220 ;
  assign y9414 = n28222 ;
  assign y9415 = ~n28225 ;
  assign y9416 = ~n28226 ;
  assign y9417 = n28227 ;
  assign y9418 = ~n28229 ;
  assign y9419 = ~n28232 ;
  assign y9420 = n28234 ;
  assign y9421 = n28235 ;
  assign y9422 = n28236 ;
  assign y9423 = ~n28238 ;
  assign y9424 = n28243 ;
  assign y9425 = ~n28244 ;
  assign y9426 = ~n28246 ;
  assign y9427 = n28247 ;
  assign y9428 = n28250 ;
  assign y9429 = ~n28256 ;
  assign y9430 = n28259 ;
  assign y9431 = ~1'b0 ;
  assign y9432 = ~1'b0 ;
  assign y9433 = ~n28261 ;
  assign y9434 = n28268 ;
  assign y9435 = ~n28269 ;
  assign y9436 = n28270 ;
  assign y9437 = ~n28271 ;
  assign y9438 = ~n28276 ;
  assign y9439 = ~n28286 ;
  assign y9440 = ~1'b0 ;
  assign y9441 = ~n28288 ;
  assign y9442 = ~1'b0 ;
  assign y9443 = n28290 ;
  assign y9444 = n28291 ;
  assign y9445 = ~n28292 ;
  assign y9446 = n28294 ;
  assign y9447 = ~n28295 ;
  assign y9448 = ~n28296 ;
  assign y9449 = ~1'b0 ;
  assign y9450 = ~n28298 ;
  assign y9451 = n28299 ;
  assign y9452 = ~n28300 ;
  assign y9453 = n28302 ;
  assign y9454 = ~n28304 ;
  assign y9455 = n28305 ;
  assign y9456 = n28308 ;
  assign y9457 = n28309 ;
  assign y9458 = ~n28310 ;
  assign y9459 = n28312 ;
  assign y9460 = n28316 ;
  assign y9461 = ~1'b0 ;
  assign y9462 = n28320 ;
  assign y9463 = ~n28322 ;
  assign y9464 = ~n28324 ;
  assign y9465 = ~n28325 ;
  assign y9466 = ~1'b0 ;
  assign y9467 = ~n28329 ;
  assign y9468 = n28330 ;
  assign y9469 = n28331 ;
  assign y9470 = n28332 ;
  assign y9471 = ~n28333 ;
  assign y9472 = n25939 ;
  assign y9473 = ~n28334 ;
  assign y9474 = ~n28335 ;
  assign y9475 = ~1'b0 ;
  assign y9476 = ~1'b0 ;
  assign y9477 = n28337 ;
  assign y9478 = ~n28339 ;
  assign y9479 = ~n28342 ;
  assign y9480 = n28343 ;
  assign y9481 = n28345 ;
  assign y9482 = n28347 ;
  assign y9483 = ~n28350 ;
  assign y9484 = n28352 ;
  assign y9485 = ~n28357 ;
  assign y9486 = ~n28358 ;
  assign y9487 = ~n28359 ;
  assign y9488 = ~n28360 ;
  assign y9489 = ~1'b0 ;
  assign y9490 = n28361 ;
  assign y9491 = ~n28362 ;
  assign y9492 = ~n28364 ;
  assign y9493 = n28367 ;
  assign y9494 = ~n28368 ;
  assign y9495 = n28370 ;
  assign y9496 = ~n28372 ;
  assign y9497 = ~n28376 ;
  assign y9498 = n28378 ;
  assign y9499 = n28380 ;
  assign y9500 = n28382 ;
  assign y9501 = ~n28384 ;
  assign y9502 = n28387 ;
  assign y9503 = ~n28389 ;
  assign y9504 = ~1'b0 ;
  assign y9505 = ~1'b0 ;
  assign y9506 = ~n28390 ;
  assign y9507 = ~n28391 ;
  assign y9508 = ~n28393 ;
  assign y9509 = n28396 ;
  assign y9510 = ~n22195 ;
  assign y9511 = n28397 ;
  assign y9512 = ~n28399 ;
  assign y9513 = ~1'b0 ;
  assign y9514 = ~n28401 ;
  assign y9515 = n28404 ;
  assign y9516 = ~1'b0 ;
  assign y9517 = ~n28405 ;
  assign y9518 = ~n28406 ;
  assign y9519 = ~n28408 ;
  assign y9520 = ~n28414 ;
  assign y9521 = n28416 ;
  assign y9522 = ~n28418 ;
  assign y9523 = ~1'b0 ;
  assign y9524 = ~n28421 ;
  assign y9525 = ~n28422 ;
  assign y9526 = ~n28423 ;
  assign y9527 = ~n28424 ;
  assign y9528 = n28425 ;
  assign y9529 = n28430 ;
  assign y9530 = ~n28432 ;
  assign y9531 = n28434 ;
  assign y9532 = n28436 ;
  assign y9533 = ~1'b0 ;
  assign y9534 = ~n28439 ;
  assign y9535 = ~n28440 ;
  assign y9536 = ~n28442 ;
  assign y9537 = ~n28443 ;
  assign y9538 = n28444 ;
  assign y9539 = n28445 ;
  assign y9540 = ~n28447 ;
  assign y9541 = ~n28450 ;
  assign y9542 = n28451 ;
  assign y9543 = ~1'b0 ;
  assign y9544 = ~n28453 ;
  assign y9545 = ~1'b0 ;
  assign y9546 = ~n28455 ;
  assign y9547 = ~n28461 ;
  assign y9548 = ~n28462 ;
  assign y9549 = n28465 ;
  assign y9550 = ~n28466 ;
  assign y9551 = ~n28467 ;
  assign y9552 = n28468 ;
  assign y9553 = ~n28469 ;
  assign y9554 = ~n28471 ;
  assign y9555 = ~n28474 ;
  assign y9556 = ~n28478 ;
  assign y9557 = ~1'b0 ;
  assign y9558 = ~n28480 ;
  assign y9559 = n28483 ;
  assign y9560 = n28484 ;
  assign y9561 = ~n28487 ;
  assign y9562 = n28488 ;
  assign y9563 = n28489 ;
  assign y9564 = n28492 ;
  assign y9565 = n28495 ;
  assign y9566 = n28499 ;
  assign y9567 = ~n28501 ;
  assign y9568 = n28502 ;
  assign y9569 = ~n28505 ;
  assign y9570 = n28507 ;
  assign y9571 = n28508 ;
  assign y9572 = ~n28509 ;
  assign y9573 = ~n28513 ;
  assign y9574 = n28514 ;
  assign y9575 = n11011 ;
  assign y9576 = ~1'b0 ;
  assign y9577 = ~n28524 ;
  assign y9578 = ~n28527 ;
  assign y9579 = ~n28529 ;
  assign y9580 = ~n28530 ;
  assign y9581 = ~n28531 ;
  assign y9582 = ~n28534 ;
  assign y9583 = ~n28536 ;
  assign y9584 = ~n10884 ;
  assign y9585 = ~1'b0 ;
  assign y9586 = ~n28538 ;
  assign y9587 = ~n28540 ;
  assign y9588 = ~n28541 ;
  assign y9589 = n28542 ;
  assign y9590 = ~n28545 ;
  assign y9591 = ~n28546 ;
  assign y9592 = ~n28548 ;
  assign y9593 = n28551 ;
  assign y9594 = ~n28558 ;
  assign y9595 = ~n28559 ;
  assign y9596 = n28560 ;
  assign y9597 = n28563 ;
  assign y9598 = ~n28564 ;
  assign y9599 = n28569 ;
  assign y9600 = ~n28572 ;
  assign y9601 = ~n28573 ;
  assign y9602 = n28576 ;
  assign y9603 = ~n28578 ;
  assign y9604 = n28581 ;
  assign y9605 = ~n28583 ;
  assign y9606 = n28585 ;
  assign y9607 = n28588 ;
  assign y9608 = n28589 ;
  assign y9609 = ~n28590 ;
  assign y9610 = n28592 ;
  assign y9611 = ~n28594 ;
  assign y9612 = ~n28597 ;
  assign y9613 = n28598 ;
  assign y9614 = ~1'b0 ;
  assign y9615 = ~1'b0 ;
  assign y9616 = ~n28601 ;
  assign y9617 = ~n28603 ;
  assign y9618 = n28606 ;
  assign y9619 = ~n28609 ;
  assign y9620 = n28610 ;
  assign y9621 = ~n28611 ;
  assign y9622 = ~n28613 ;
  assign y9623 = n28615 ;
  assign y9624 = ~n28619 ;
  assign y9625 = ~1'b0 ;
  assign y9626 = ~1'b0 ;
  assign y9627 = n28622 ;
  assign y9628 = n28625 ;
  assign y9629 = n28626 ;
  assign y9630 = n28627 ;
  assign y9631 = ~n28628 ;
  assign y9632 = n28630 ;
  assign y9633 = ~n28631 ;
  assign y9634 = n28632 ;
  assign y9635 = ~n28633 ;
  assign y9636 = ~1'b0 ;
  assign y9637 = ~1'b0 ;
  assign y9638 = ~1'b0 ;
  assign y9639 = ~n28636 ;
  assign y9640 = ~n28637 ;
  assign y9641 = ~n28638 ;
  assign y9642 = n28639 ;
  assign y9643 = ~n28642 ;
  assign y9644 = ~n28646 ;
  assign y9645 = n28647 ;
  assign y9646 = ~1'b0 ;
  assign y9647 = n28650 ;
  assign y9648 = 1'b0 ;
  assign y9649 = ~1'b0 ;
  assign y9650 = n28652 ;
  assign y9651 = n28654 ;
  assign y9652 = n28655 ;
  assign y9653 = ~n28656 ;
  assign y9654 = ~n28657 ;
  assign y9655 = n28660 ;
  assign y9656 = ~1'b0 ;
  assign y9657 = ~1'b0 ;
  assign y9658 = ~n28666 ;
  assign y9659 = ~n28668 ;
  assign y9660 = ~1'b0 ;
  assign y9661 = ~n28669 ;
  assign y9662 = n28676 ;
  assign y9663 = ~n28681 ;
  assign y9664 = ~n28686 ;
  assign y9665 = n28687 ;
  assign y9666 = ~n28690 ;
  assign y9667 = ~n28691 ;
  assign y9668 = ~n28695 ;
  assign y9669 = ~1'b0 ;
  assign y9670 = ~n28698 ;
  assign y9671 = ~n28699 ;
  assign y9672 = n28702 ;
  assign y9673 = n28705 ;
  assign y9674 = ~n28706 ;
  assign y9675 = ~n28710 ;
  assign y9676 = ~n28712 ;
  assign y9677 = ~n28719 ;
  assign y9678 = n28722 ;
  assign y9679 = ~n28726 ;
  assign y9680 = n28728 ;
  assign y9681 = n28734 ;
  assign y9682 = n28737 ;
  assign y9683 = n28738 ;
  assign y9684 = ~n28739 ;
  assign y9685 = n28740 ;
  assign y9686 = ~n28742 ;
  assign y9687 = ~1'b0 ;
  assign y9688 = n28747 ;
  assign y9689 = ~1'b0 ;
  assign y9690 = ~1'b0 ;
  assign y9691 = n28748 ;
  assign y9692 = ~n28749 ;
  assign y9693 = n28750 ;
  assign y9694 = n28752 ;
  assign y9695 = n25151 ;
  assign y9696 = ~n28754 ;
  assign y9697 = ~1'b0 ;
  assign y9698 = ~n28756 ;
  assign y9699 = ~n28758 ;
  assign y9700 = ~1'b0 ;
  assign y9701 = n28760 ;
  assign y9702 = ~n28763 ;
  assign y9703 = ~n28764 ;
  assign y9704 = n28765 ;
  assign y9705 = n28766 ;
  assign y9706 = ~n760 ;
  assign y9707 = ~1'b0 ;
  assign y9708 = n28770 ;
  assign y9709 = ~n28773 ;
  assign y9710 = n28774 ;
  assign y9711 = ~1'b0 ;
  assign y9712 = ~n28776 ;
  assign y9713 = n28779 ;
  assign y9714 = n28780 ;
  assign y9715 = ~n28782 ;
  assign y9716 = n28784 ;
  assign y9717 = n28785 ;
  assign y9718 = ~1'b0 ;
  assign y9719 = ~1'b0 ;
  assign y9720 = ~n28786 ;
  assign y9721 = ~n28792 ;
  assign y9722 = n28796 ;
  assign y9723 = n28798 ;
  assign y9724 = n28803 ;
  assign y9725 = n28807 ;
  assign y9726 = ~n28808 ;
  assign y9727 = n28809 ;
  assign y9728 = n28812 ;
  assign y9729 = n28814 ;
  assign y9730 = ~1'b0 ;
  assign y9731 = n28818 ;
  assign y9732 = ~n28823 ;
  assign y9733 = ~n28828 ;
  assign y9734 = n28829 ;
  assign y9735 = ~1'b0 ;
  assign y9736 = ~n28833 ;
  assign y9737 = ~n28835 ;
  assign y9738 = n28838 ;
  assign y9739 = ~1'b0 ;
  assign y9740 = n28842 ;
  assign y9741 = n28844 ;
  assign y9742 = n28847 ;
  assign y9743 = n28851 ;
  assign y9744 = ~n28853 ;
  assign y9745 = ~n28854 ;
  assign y9746 = ~n28855 ;
  assign y9747 = n28859 ;
  assign y9748 = n28860 ;
  assign y9749 = n28861 ;
  assign y9750 = n28863 ;
  assign y9751 = n28865 ;
  assign y9752 = ~1'b0 ;
  assign y9753 = n28870 ;
  assign y9754 = ~n28871 ;
  assign y9755 = n28873 ;
  assign y9756 = n28874 ;
  assign y9757 = ~n28875 ;
  assign y9758 = n28876 ;
  assign y9759 = n28877 ;
  assign y9760 = ~n28879 ;
  assign y9761 = n28881 ;
  assign y9762 = ~n28885 ;
  assign y9763 = ~1'b0 ;
  assign y9764 = n28888 ;
  assign y9765 = ~n28891 ;
  assign y9766 = n28893 ;
  assign y9767 = ~n28894 ;
  assign y9768 = ~n28897 ;
  assign y9769 = ~n28898 ;
  assign y9770 = ~1'b0 ;
  assign y9771 = ~n28899 ;
  assign y9772 = n28903 ;
  assign y9773 = n28904 ;
  assign y9774 = ~1'b0 ;
  assign y9775 = ~n28906 ;
  assign y9776 = n28908 ;
  assign y9777 = n28909 ;
  assign y9778 = n28912 ;
  assign y9779 = n28913 ;
  assign y9780 = n28916 ;
  assign y9781 = n28918 ;
  assign y9782 = ~n28920 ;
  assign y9783 = n28921 ;
  assign y9784 = ~n28922 ;
  assign y9785 = n28923 ;
  assign y9786 = n28924 ;
  assign y9787 = ~n28925 ;
  assign y9788 = n28926 ;
  assign y9789 = n28928 ;
  assign y9790 = n28930 ;
  assign y9791 = ~1'b0 ;
  assign y9792 = ~n28934 ;
  assign y9793 = ~n28940 ;
  assign y9794 = n28941 ;
  assign y9795 = n28942 ;
  assign y9796 = ~n28943 ;
  assign y9797 = ~n28946 ;
  assign y9798 = ~n28947 ;
  assign y9799 = ~n28948 ;
  assign y9800 = ~n28951 ;
  assign y9801 = n28954 ;
  assign y9802 = ~n28957 ;
  assign y9803 = ~1'b0 ;
  assign y9804 = n28959 ;
  assign y9805 = ~n28960 ;
  assign y9806 = n28963 ;
  assign y9807 = n28968 ;
  assign y9808 = ~1'b0 ;
  assign y9809 = n28969 ;
  assign y9810 = ~n28974 ;
  assign y9811 = n28977 ;
  assign y9812 = ~1'b0 ;
  assign y9813 = n28983 ;
  assign y9814 = ~n28984 ;
  assign y9815 = ~n28985 ;
  assign y9816 = n28989 ;
  assign y9817 = ~n28993 ;
  assign y9818 = n28994 ;
  assign y9819 = n28996 ;
  assign y9820 = ~1'b0 ;
  assign y9821 = ~n28998 ;
  assign y9822 = n29000 ;
  assign y9823 = n29003 ;
  assign y9824 = ~n29005 ;
  assign y9825 = n29006 ;
  assign y9826 = ~n29007 ;
  assign y9827 = ~n29009 ;
  assign y9828 = ~n29013 ;
  assign y9829 = ~n29014 ;
  assign y9830 = 1'b0 ;
  assign y9831 = n29022 ;
  assign y9832 = ~n29025 ;
  assign y9833 = n19734 ;
  assign y9834 = n29028 ;
  assign y9835 = n29029 ;
  assign y9836 = ~n29034 ;
  assign y9837 = ~n29035 ;
  assign y9838 = ~n29037 ;
  assign y9839 = ~n29038 ;
  assign y9840 = n29044 ;
  assign y9841 = n29048 ;
  assign y9842 = ~n29049 ;
  assign y9843 = ~n29051 ;
  assign y9844 = ~n29053 ;
  assign y9845 = ~n29055 ;
  assign y9846 = ~n29056 ;
  assign y9847 = ~n29057 ;
  assign y9848 = n29058 ;
  assign y9849 = n29060 ;
  assign y9850 = ~n29062 ;
  assign y9851 = ~1'b0 ;
  assign y9852 = ~n29063 ;
  assign y9853 = ~1'b0 ;
  assign y9854 = ~n29065 ;
  assign y9855 = ~n29071 ;
  assign y9856 = ~n29073 ;
  assign y9857 = ~n29074 ;
  assign y9858 = n29077 ;
  assign y9859 = n29081 ;
  assign y9860 = n29089 ;
  assign y9861 = n29091 ;
  assign y9862 = ~1'b0 ;
  assign y9863 = ~1'b0 ;
  assign y9864 = n29094 ;
  assign y9865 = ~n29095 ;
  assign y9866 = ~n29097 ;
  assign y9867 = ~n29101 ;
  assign y9868 = ~n29103 ;
  assign y9869 = n29104 ;
  assign y9870 = ~1'b0 ;
  assign y9871 = ~n29106 ;
  assign y9872 = ~1'b0 ;
  assign y9873 = ~n29109 ;
  assign y9874 = n29111 ;
  assign y9875 = n29114 ;
  assign y9876 = ~n29118 ;
  assign y9877 = ~n29122 ;
  assign y9878 = ~n29123 ;
  assign y9879 = n29127 ;
  assign y9880 = ~1'b0 ;
  assign y9881 = n29129 ;
  assign y9882 = n29132 ;
  assign y9883 = ~n29134 ;
  assign y9884 = ~n29136 ;
  assign y9885 = n29137 ;
  assign y9886 = n29139 ;
  assign y9887 = ~n29147 ;
  assign y9888 = n29149 ;
  assign y9889 = ~n29152 ;
  assign y9890 = n29154 ;
  assign y9891 = ~n29161 ;
  assign y9892 = 1'b0 ;
  assign y9893 = n29162 ;
  assign y9894 = n29163 ;
  assign y9895 = ~n29164 ;
  assign y9896 = n29165 ;
  assign y9897 = ~n29166 ;
  assign y9898 = n29167 ;
  assign y9899 = ~n29169 ;
  assign y9900 = ~1'b0 ;
  assign y9901 = n29172 ;
  assign y9902 = ~n29174 ;
  assign y9903 = n29176 ;
  assign y9904 = n21561 ;
  assign y9905 = ~n29179 ;
  assign y9906 = n29183 ;
  assign y9907 = ~n29184 ;
  assign y9908 = ~n29186 ;
  assign y9909 = ~1'b0 ;
  assign y9910 = ~n29188 ;
  assign y9911 = n29194 ;
  assign y9912 = ~n29195 ;
  assign y9913 = n29198 ;
  assign y9914 = ~n29200 ;
  assign y9915 = ~n29203 ;
  assign y9916 = n29204 ;
  assign y9917 = n29206 ;
  assign y9918 = ~n29207 ;
  assign y9919 = ~n29208 ;
  assign y9920 = ~1'b0 ;
  assign y9921 = ~n9109 ;
  assign y9922 = ~1'b0 ;
  assign y9923 = ~1'b0 ;
  assign y9924 = ~n29209 ;
  assign y9925 = n29212 ;
  assign y9926 = ~n29217 ;
  assign y9927 = ~n29221 ;
  assign y9928 = n29222 ;
  assign y9929 = ~1'b0 ;
  assign y9930 = ~n29224 ;
  assign y9931 = ~1'b0 ;
  assign y9932 = ~n29226 ;
  assign y9933 = ~n29227 ;
  assign y9934 = ~n29229 ;
  assign y9935 = n29230 ;
  assign y9936 = ~n29233 ;
  assign y9937 = ~n29236 ;
  assign y9938 = ~n29239 ;
  assign y9939 = ~n29241 ;
  assign y9940 = n29243 ;
  assign y9941 = n29245 ;
  assign y9942 = ~n29246 ;
  assign y9943 = ~n29250 ;
  assign y9944 = n29252 ;
  assign y9945 = ~n29258 ;
  assign y9946 = n29259 ;
  assign y9947 = n29261 ;
  assign y9948 = n29263 ;
  assign y9949 = n29267 ;
  assign y9950 = n29269 ;
  assign y9951 = ~1'b0 ;
  assign y9952 = n29270 ;
  assign y9953 = ~n29271 ;
  assign y9954 = ~n29272 ;
  assign y9955 = n29273 ;
  assign y9956 = n13868 ;
  assign y9957 = n29274 ;
  assign y9958 = ~n29277 ;
  assign y9959 = ~1'b0 ;
  assign y9960 = ~n29281 ;
  assign y9961 = n29283 ;
  assign y9962 = ~n29284 ;
  assign y9963 = ~n29288 ;
  assign y9964 = n29291 ;
  assign y9965 = n29294 ;
  assign y9966 = ~n29297 ;
  assign y9967 = n29301 ;
  assign y9968 = ~n29307 ;
  assign y9969 = ~1'b0 ;
  assign y9970 = n29313 ;
  assign y9971 = ~1'b0 ;
  assign y9972 = ~1'b0 ;
  assign y9973 = ~n29318 ;
  assign y9974 = ~n29319 ;
  assign y9975 = n29327 ;
  assign y9976 = ~n29330 ;
  assign y9977 = n29331 ;
  assign y9978 = ~n29332 ;
  assign y9979 = ~n29334 ;
  assign y9980 = n29336 ;
  assign y9981 = ~n29340 ;
  assign y9982 = ~1'b0 ;
  assign y9983 = ~n29342 ;
  assign y9984 = ~n29343 ;
  assign y9985 = n29351 ;
  assign y9986 = n29356 ;
  assign y9987 = ~n29357 ;
  assign y9988 = ~n29359 ;
  assign y9989 = n29362 ;
  assign y9990 = ~n29364 ;
  assign y9991 = ~n29367 ;
  assign y9992 = ~1'b0 ;
  assign y9993 = ~1'b0 ;
  assign y9994 = n29371 ;
  assign y9995 = n19346 ;
  assign y9996 = n29372 ;
  assign y9997 = n29375 ;
  assign y9998 = n29376 ;
  assign y9999 = ~n29377 ;
  assign y10000 = ~n29380 ;
  assign y10001 = n29385 ;
  assign y10002 = ~1'b0 ;
  assign y10003 = ~1'b0 ;
  assign y10004 = ~n29013 ;
  assign y10005 = n29389 ;
  assign y10006 = n29391 ;
  assign y10007 = n29393 ;
  assign y10008 = ~n29397 ;
  assign y10009 = ~n29399 ;
  assign y10010 = ~n29400 ;
  assign y10011 = ~n29403 ;
  assign y10012 = n29407 ;
  assign y10013 = n29409 ;
  assign y10014 = n29411 ;
  assign y10015 = ~1'b0 ;
  assign y10016 = ~n29412 ;
  assign y10017 = n29413 ;
  assign y10018 = ~n29414 ;
  assign y10019 = n29415 ;
  assign y10020 = ~n29418 ;
  assign y10021 = ~n29419 ;
  assign y10022 = ~1'b0 ;
  assign y10023 = n29420 ;
  assign y10024 = n29423 ;
  assign y10025 = n29425 ;
  assign y10026 = n29426 ;
  assign y10027 = n29427 ;
  assign y10028 = ~n29431 ;
  assign y10029 = ~n29436 ;
  assign y10030 = n29437 ;
  assign y10031 = ~n29444 ;
  assign y10032 = n29446 ;
  assign y10033 = ~n29451 ;
  assign y10034 = ~n29452 ;
  assign y10035 = ~n29454 ;
  assign y10036 = ~n29456 ;
  assign y10037 = ~1'b0 ;
  assign y10038 = n29457 ;
  assign y10039 = n29458 ;
  assign y10040 = ~n29459 ;
  assign y10041 = ~n29460 ;
  assign y10042 = ~n29461 ;
  assign y10043 = ~n29466 ;
  assign y10044 = ~n29468 ;
  assign y10045 = n9562 ;
  assign y10046 = n29472 ;
  assign y10047 = n29474 ;
  assign y10048 = ~n29475 ;
  assign y10049 = n29477 ;
  assign y10050 = ~n29478 ;
  assign y10051 = n29479 ;
  assign y10052 = ~n29480 ;
  assign y10053 = ~n29484 ;
  assign y10054 = ~n29488 ;
  assign y10055 = ~1'b0 ;
  assign y10056 = n29489 ;
  assign y10057 = n20840 ;
  assign y10058 = n29494 ;
  assign y10059 = ~n29498 ;
  assign y10060 = n29499 ;
  assign y10061 = n29500 ;
  assign y10062 = 1'b0 ;
  assign y10063 = ~n29508 ;
  assign y10064 = ~n29513 ;
  assign y10065 = n29514 ;
  assign y10066 = ~n29515 ;
  assign y10067 = n29516 ;
  assign y10068 = n29518 ;
  assign y10069 = n29519 ;
  assign y10070 = ~n29522 ;
  assign y10071 = n29523 ;
  assign y10072 = ~n29524 ;
  assign y10073 = ~n29526 ;
  assign y10074 = ~n29527 ;
  assign y10075 = ~n29529 ;
  assign y10076 = ~1'b0 ;
  assign y10077 = n29530 ;
  assign y10078 = ~n29531 ;
  assign y10079 = n29533 ;
  assign y10080 = n29539 ;
  assign y10081 = ~n29540 ;
  assign y10082 = n29542 ;
  assign y10083 = n29546 ;
  assign y10084 = ~1'b0 ;
  assign y10085 = ~1'b0 ;
  assign y10086 = n29552 ;
  assign y10087 = n29553 ;
  assign y10088 = n29554 ;
  assign y10089 = ~n29555 ;
  assign y10090 = n15025 ;
  assign y10091 = n29556 ;
  assign y10092 = ~n29562 ;
  assign y10093 = ~1'b0 ;
  assign y10094 = n29563 ;
  assign y10095 = ~1'b0 ;
  assign y10096 = n29564 ;
  assign y10097 = ~n29565 ;
  assign y10098 = ~n29568 ;
  assign y10099 = n29569 ;
  assign y10100 = n29571 ;
  assign y10101 = n29574 ;
  assign y10102 = ~1'b0 ;
  assign y10103 = n29576 ;
  assign y10104 = n29580 ;
  assign y10105 = ~n29583 ;
  assign y10106 = ~n2455 ;
  assign y10107 = ~n29585 ;
  assign y10108 = n29586 ;
  assign y10109 = n29587 ;
  assign y10110 = n29588 ;
  assign y10111 = ~1'b0 ;
  assign y10112 = n29592 ;
  assign y10113 = ~1'b0 ;
  assign y10114 = ~n29594 ;
  assign y10115 = n29596 ;
  assign y10116 = n29601 ;
  assign y10117 = ~n29606 ;
  assign y10118 = n29611 ;
  assign y10119 = n29612 ;
  assign y10120 = ~1'b0 ;
  assign y10121 = n29615 ;
  assign y10122 = ~n29618 ;
  assign y10123 = ~n29620 ;
  assign y10124 = ~1'b0 ;
  assign y10125 = n4865 ;
  assign y10126 = ~n29623 ;
  assign y10127 = ~n29625 ;
  assign y10128 = n29626 ;
  assign y10129 = ~n29628 ;
  assign y10130 = n29629 ;
  assign y10131 = n29632 ;
  assign y10132 = ~n29638 ;
  assign y10133 = n29639 ;
  assign y10134 = n29641 ;
  assign y10135 = ~n29642 ;
  assign y10136 = ~n29648 ;
  assign y10137 = n29649 ;
  assign y10138 = ~n29650 ;
  assign y10139 = ~n29652 ;
  assign y10140 = ~n29653 ;
  assign y10141 = n29655 ;
  assign y10142 = ~n29657 ;
  assign y10143 = n29658 ;
  assign y10144 = n29660 ;
  assign y10145 = n29662 ;
  assign y10146 = ~1'b0 ;
  assign y10147 = n29664 ;
  assign y10148 = ~n29666 ;
  assign y10149 = n29667 ;
  assign y10150 = n29669 ;
  assign y10151 = n29670 ;
  assign y10152 = ~n29671 ;
  assign y10153 = n29674 ;
  assign y10154 = n29675 ;
  assign y10155 = ~1'b0 ;
  assign y10156 = ~1'b0 ;
  assign y10157 = ~n29679 ;
  assign y10158 = n29682 ;
  assign y10159 = n29684 ;
  assign y10160 = n29687 ;
  assign y10161 = ~n29689 ;
  assign y10162 = n29691 ;
  assign y10163 = n29693 ;
  assign y10164 = ~n29695 ;
  assign y10165 = ~n29696 ;
  assign y10166 = ~1'b0 ;
  assign y10167 = ~n29701 ;
  assign y10168 = ~1'b0 ;
  assign y10169 = ~n29702 ;
  assign y10170 = ~n29707 ;
  assign y10171 = ~n29708 ;
  assign y10172 = ~1'b0 ;
  assign y10173 = ~n29709 ;
  assign y10174 = ~n29710 ;
  assign y10175 = n29711 ;
  assign y10176 = ~1'b0 ;
  assign y10177 = n29716 ;
  assign y10178 = n29721 ;
  assign y10179 = ~1'b0 ;
  assign y10180 = n29722 ;
  assign y10181 = ~n29725 ;
  assign y10182 = ~n29726 ;
  assign y10183 = ~n29728 ;
  assign y10184 = ~n29729 ;
  assign y10185 = n29732 ;
  assign y10186 = n29734 ;
  assign y10187 = n29736 ;
  assign y10188 = n29739 ;
  assign y10189 = ~n29740 ;
  assign y10190 = n29741 ;
  assign y10191 = n29742 ;
  assign y10192 = ~n29743 ;
  assign y10193 = n29749 ;
  assign y10194 = ~n29751 ;
  assign y10195 = ~n29753 ;
  assign y10196 = n29757 ;
  assign y10197 = 1'b0 ;
  assign y10198 = ~n29759 ;
  assign y10199 = n29761 ;
  assign y10200 = ~n29764 ;
  assign y10201 = ~n29766 ;
  assign y10202 = n29772 ;
  assign y10203 = n29776 ;
  assign y10204 = ~1'b0 ;
  assign y10205 = ~n29778 ;
  assign y10206 = ~n29780 ;
  assign y10207 = n29781 ;
  assign y10208 = ~1'b0 ;
  assign y10209 = n29785 ;
  assign y10210 = ~n29786 ;
  assign y10211 = ~n29787 ;
  assign y10212 = n29790 ;
  assign y10213 = ~n29792 ;
  assign y10214 = ~n29793 ;
  assign y10215 = n29794 ;
  assign y10216 = n29795 ;
  assign y10217 = ~n29798 ;
  assign y10218 = n29801 ;
  assign y10219 = n29804 ;
  assign y10220 = n29806 ;
  assign y10221 = ~1'b0 ;
  assign y10222 = ~n29808 ;
  assign y10223 = n29809 ;
  assign y10224 = n29811 ;
  assign y10225 = ~n29819 ;
  assign y10226 = n29822 ;
  assign y10227 = ~n29826 ;
  assign y10228 = ~n29828 ;
  assign y10229 = n29829 ;
  assign y10230 = n29830 ;
  assign y10231 = n29836 ;
  assign y10232 = ~n29841 ;
  assign y10233 = n29847 ;
  assign y10234 = n29853 ;
  assign y10235 = n29854 ;
  assign y10236 = n29855 ;
  assign y10237 = ~n29857 ;
  assign y10238 = ~n29858 ;
  assign y10239 = n29860 ;
  assign y10240 = n29862 ;
  assign y10241 = ~n29864 ;
  assign y10242 = n29866 ;
  assign y10243 = ~1'b0 ;
  assign y10244 = ~n29867 ;
  assign y10245 = ~n29869 ;
  assign y10246 = ~n29876 ;
  assign y10247 = n29878 ;
  assign y10248 = n29879 ;
  assign y10249 = n29881 ;
  assign y10250 = n29883 ;
  assign y10251 = ~1'b0 ;
  assign y10252 = ~n29884 ;
  assign y10253 = ~n29887 ;
  assign y10254 = ~n29889 ;
  assign y10255 = ~n29892 ;
  assign y10256 = n29894 ;
  assign y10257 = n29897 ;
  assign y10258 = ~n29900 ;
  assign y10259 = n29902 ;
  assign y10260 = ~1'b0 ;
  assign y10261 = ~n29904 ;
  assign y10262 = ~n29912 ;
  assign y10263 = n29914 ;
  assign y10264 = ~n29917 ;
  assign y10265 = n29918 ;
  assign y10266 = n29919 ;
  assign y10267 = ~n29920 ;
  assign y10268 = n29925 ;
  assign y10269 = ~n29928 ;
  assign y10270 = n29932 ;
  assign y10271 = n29933 ;
  assign y10272 = ~n29935 ;
  assign y10273 = n29939 ;
  assign y10274 = n29944 ;
  assign y10275 = ~n29947 ;
  assign y10276 = n29954 ;
  assign y10277 = n29955 ;
  assign y10278 = ~n29956 ;
  assign y10279 = ~1'b0 ;
  assign y10280 = ~n29957 ;
  assign y10281 = n29960 ;
  assign y10282 = n29962 ;
  assign y10283 = n29963 ;
  assign y10284 = ~n29964 ;
  assign y10285 = ~n29975 ;
  assign y10286 = ~n29976 ;
  assign y10287 = ~n29979 ;
  assign y10288 = ~n29983 ;
  assign y10289 = n29984 ;
  assign y10290 = ~n29987 ;
  assign y10291 = ~n29989 ;
  assign y10292 = ~n29993 ;
  assign y10293 = ~1'b0 ;
  assign y10294 = ~n29994 ;
  assign y10295 = ~n29995 ;
  assign y10296 = n29998 ;
  assign y10297 = ~n29999 ;
  assign y10298 = n30000 ;
  assign y10299 = ~n30002 ;
  assign y10300 = ~n30005 ;
  assign y10301 = ~n30007 ;
  assign y10302 = ~1'b0 ;
  assign y10303 = ~n30012 ;
  assign y10304 = ~n30015 ;
  assign y10305 = ~n30019 ;
  assign y10306 = n30020 ;
  assign y10307 = n30027 ;
  assign y10308 = n30028 ;
  assign y10309 = ~n30030 ;
  assign y10310 = ~n30031 ;
  assign y10311 = n30036 ;
  assign y10312 = ~1'b0 ;
  assign y10313 = ~1'b0 ;
  assign y10314 = ~1'b0 ;
  assign y10315 = ~n30037 ;
  assign y10316 = ~n30038 ;
  assign y10317 = ~n30044 ;
  assign y10318 = ~n30046 ;
  assign y10319 = ~n28938 ;
  assign y10320 = n30049 ;
  assign y10321 = ~n30052 ;
  assign y10322 = n30056 ;
  assign y10323 = n30058 ;
  assign y10324 = ~n30060 ;
  assign y10325 = ~1'b0 ;
  assign y10326 = n30061 ;
  assign y10327 = n30062 ;
  assign y10328 = n30063 ;
  assign y10329 = n30070 ;
  assign y10330 = ~n30071 ;
  assign y10331 = n30077 ;
  assign y10332 = ~1'b0 ;
  assign y10333 = ~n30079 ;
  assign y10334 = n30081 ;
  assign y10335 = ~1'b0 ;
  assign y10336 = ~1'b0 ;
  assign y10337 = n30082 ;
  assign y10338 = n30087 ;
  assign y10339 = ~n30091 ;
  assign y10340 = n30093 ;
  assign y10341 = ~n30097 ;
  assign y10342 = n30101 ;
  assign y10343 = ~1'b0 ;
  assign y10344 = n30103 ;
  assign y10345 = ~n30106 ;
  assign y10346 = n30107 ;
  assign y10347 = ~n30108 ;
  assign y10348 = n30109 ;
  assign y10349 = n30110 ;
  assign y10350 = n30115 ;
  assign y10351 = ~n30117 ;
  assign y10352 = ~1'b0 ;
  assign y10353 = n30119 ;
  assign y10354 = ~n30124 ;
  assign y10355 = n30126 ;
  assign y10356 = ~n30127 ;
  assign y10357 = n30131 ;
  assign y10358 = ~n30136 ;
  assign y10359 = n30137 ;
  assign y10360 = n30139 ;
  assign y10361 = n30142 ;
  assign y10362 = ~1'b0 ;
  assign y10363 = ~n30144 ;
  assign y10364 = ~1'b0 ;
  assign y10365 = ~1'b0 ;
  assign y10366 = ~n30148 ;
  assign y10367 = ~n30149 ;
  assign y10368 = n30151 ;
  assign y10369 = n30152 ;
  assign y10370 = n30155 ;
  assign y10371 = n7076 ;
  assign y10372 = n30158 ;
  assign y10373 = ~n30161 ;
  assign y10374 = n30162 ;
  assign y10375 = ~n30163 ;
  assign y10376 = n30165 ;
  assign y10377 = ~n30167 ;
  assign y10378 = n30168 ;
  assign y10379 = n30169 ;
  assign y10380 = n30170 ;
  assign y10381 = ~n30175 ;
  assign y10382 = n30176 ;
  assign y10383 = n30178 ;
  assign y10384 = n30182 ;
  assign y10385 = n30183 ;
  assign y10386 = ~n30185 ;
  assign y10387 = n30186 ;
  assign y10388 = n30195 ;
  assign y10389 = ~n30200 ;
  assign y10390 = n30201 ;
  assign y10391 = ~n30208 ;
  assign y10392 = n30210 ;
  assign y10393 = ~1'b0 ;
  assign y10394 = n30211 ;
  assign y10395 = ~n30213 ;
  assign y10396 = ~n30215 ;
  assign y10397 = ~n30217 ;
  assign y10398 = ~n30218 ;
  assign y10399 = n30219 ;
  assign y10400 = n30221 ;
  assign y10401 = n30222 ;
  assign y10402 = ~n30224 ;
  assign y10403 = ~n30226 ;
  assign y10404 = ~1'b0 ;
  assign y10405 = n30235 ;
  assign y10406 = ~1'b0 ;
  assign y10407 = n30236 ;
  assign y10408 = n30239 ;
  assign y10409 = ~n30243 ;
  assign y10410 = n30247 ;
  assign y10411 = ~n30248 ;
  assign y10412 = n30251 ;
  assign y10413 = n30253 ;
  assign y10414 = n30255 ;
  assign y10415 = ~1'b0 ;
  assign y10416 = n30264 ;
  assign y10417 = n30270 ;
  assign y10418 = n30271 ;
  assign y10419 = ~n30273 ;
  assign y10420 = ~n30275 ;
  assign y10421 = ~n30279 ;
  assign y10422 = n30283 ;
  assign y10423 = n30285 ;
  assign y10424 = ~1'b0 ;
  assign y10425 = ~1'b0 ;
  assign y10426 = n30287 ;
  assign y10427 = n30295 ;
  assign y10428 = ~n30297 ;
  assign y10429 = ~n30299 ;
  assign y10430 = n6447 ;
  assign y10431 = n30300 ;
  assign y10432 = n30302 ;
  assign y10433 = n30303 ;
  assign y10434 = ~n30307 ;
  assign y10435 = n30310 ;
  assign y10436 = ~n30312 ;
  assign y10437 = ~1'b0 ;
  assign y10438 = n30314 ;
  assign y10439 = ~n30315 ;
  assign y10440 = n15521 ;
  assign y10441 = ~n30319 ;
  assign y10442 = ~n30322 ;
  assign y10443 = ~n30323 ;
  assign y10444 = n30324 ;
  assign y10445 = ~1'b0 ;
  assign y10446 = n30329 ;
  assign y10447 = ~n30330 ;
  assign y10448 = ~n30331 ;
  assign y10449 = n30332 ;
  assign y10450 = ~n30337 ;
  assign y10451 = n30338 ;
  assign y10452 = ~n30339 ;
  assign y10453 = ~n30342 ;
  assign y10454 = n30346 ;
  assign y10455 = n30348 ;
  assign y10456 = ~1'b0 ;
  assign y10457 = ~n30351 ;
  assign y10458 = ~n30353 ;
  assign y10459 = n30356 ;
  assign y10460 = ~n27162 ;
  assign y10461 = n30359 ;
  assign y10462 = n30364 ;
  assign y10463 = ~n30365 ;
  assign y10464 = n30366 ;
  assign y10465 = ~1'b0 ;
  assign y10466 = ~1'b0 ;
  assign y10467 = ~1'b0 ;
  assign y10468 = ~1'b0 ;
  assign y10469 = ~1'b0 ;
  assign y10470 = ~n30369 ;
  assign y10471 = n30370 ;
  assign y10472 = n30371 ;
  assign y10473 = ~n30372 ;
  assign y10474 = ~n30374 ;
  assign y10475 = ~n30378 ;
  assign y10476 = ~n12241 ;
  assign y10477 = ~n30381 ;
  assign y10478 = n30383 ;
  assign y10479 = ~1'b0 ;
  assign y10480 = n30384 ;
  assign y10481 = n30385 ;
  assign y10482 = ~1'b0 ;
  assign y10483 = n30386 ;
  assign y10484 = ~n30388 ;
  assign y10485 = ~n30389 ;
  assign y10486 = ~n30392 ;
  assign y10487 = ~1'b0 ;
  assign y10488 = n30393 ;
  assign y10489 = ~n30394 ;
  assign y10490 = ~n30396 ;
  assign y10491 = n30398 ;
  assign y10492 = ~n14736 ;
  assign y10493 = n30400 ;
  assign y10494 = ~n30404 ;
  assign y10495 = ~n30405 ;
  assign y10496 = ~n30406 ;
  assign y10497 = n30407 ;
  assign y10498 = n30409 ;
  assign y10499 = ~1'b0 ;
  assign y10500 = ~1'b0 ;
  assign y10501 = n30414 ;
  assign y10502 = ~n30415 ;
  assign y10503 = n30418 ;
  assign y10504 = n30419 ;
  assign y10505 = ~n30421 ;
  assign y10506 = n30422 ;
  assign y10507 = ~n30423 ;
  assign y10508 = n30425 ;
  assign y10509 = ~1'b0 ;
  assign y10510 = n30426 ;
  assign y10511 = ~n30433 ;
  assign y10512 = n30440 ;
  assign y10513 = n30441 ;
  assign y10514 = n30442 ;
  assign y10515 = ~n30443 ;
  assign y10516 = n30444 ;
  assign y10517 = ~n30447 ;
  assign y10518 = ~1'b0 ;
  assign y10519 = ~1'b0 ;
  assign y10520 = n30451 ;
  assign y10521 = ~n30454 ;
  assign y10522 = ~1'b0 ;
  assign y10523 = n30459 ;
  assign y10524 = n30460 ;
  assign y10525 = ~n30462 ;
  assign y10526 = ~n30465 ;
  assign y10527 = ~n30467 ;
  assign y10528 = ~n30470 ;
  assign y10529 = ~1'b0 ;
  assign y10530 = n30472 ;
  assign y10531 = ~1'b0 ;
  assign y10532 = n30474 ;
  assign y10533 = n30476 ;
  assign y10534 = ~n30478 ;
  assign y10535 = ~n30487 ;
  assign y10536 = n30490 ;
  assign y10537 = n30491 ;
  assign y10538 = ~n30493 ;
  assign y10539 = ~1'b0 ;
  assign y10540 = ~1'b0 ;
  assign y10541 = ~1'b0 ;
  assign y10542 = n30497 ;
  assign y10543 = ~1'b0 ;
  assign y10544 = n30500 ;
  assign y10545 = n30501 ;
  assign y10546 = n30502 ;
  assign y10547 = ~n30503 ;
  assign y10548 = n30504 ;
  assign y10549 = n30506 ;
  assign y10550 = ~1'b0 ;
  assign y10551 = ~n30510 ;
  assign y10552 = n30512 ;
  assign y10553 = ~1'b0 ;
  assign y10554 = n30513 ;
  assign y10555 = ~n30516 ;
  assign y10556 = n30519 ;
  assign y10557 = ~n30521 ;
  assign y10558 = ~n30525 ;
  assign y10559 = n30526 ;
  assign y10560 = ~n30528 ;
  assign y10561 = n30530 ;
  assign y10562 = ~1'b0 ;
  assign y10563 = n30532 ;
  assign y10564 = ~1'b0 ;
  assign y10565 = n30535 ;
  assign y10566 = ~n30536 ;
  assign y10567 = n30537 ;
  assign y10568 = n30540 ;
  assign y10569 = ~n30541 ;
  assign y10570 = ~n30542 ;
  assign y10571 = ~n30544 ;
  assign y10572 = ~1'b0 ;
  assign y10573 = ~n30551 ;
  assign y10574 = ~n30556 ;
  assign y10575 = ~1'b0 ;
  assign y10576 = ~n30557 ;
  assign y10577 = ~n30558 ;
  assign y10578 = n30559 ;
  assign y10579 = n30561 ;
  assign y10580 = ~n30562 ;
  assign y10581 = ~n30563 ;
  assign y10582 = ~1'b0 ;
  assign y10583 = n30567 ;
  assign y10584 = ~1'b0 ;
  assign y10585 = n30569 ;
  assign y10586 = n30572 ;
  assign y10587 = ~n30573 ;
  assign y10588 = ~n30584 ;
  assign y10589 = ~n30586 ;
  assign y10590 = ~n30589 ;
  assign y10591 = n30592 ;
  assign y10592 = ~1'b0 ;
  assign y10593 = ~1'b0 ;
  assign y10594 = ~n30594 ;
  assign y10595 = ~n30596 ;
  assign y10596 = n30598 ;
  assign y10597 = n30601 ;
  assign y10598 = ~n30602 ;
  assign y10599 = ~n30603 ;
  assign y10600 = ~n30604 ;
  assign y10601 = n30607 ;
  assign y10602 = ~n30609 ;
  assign y10603 = n30614 ;
  assign y10604 = ~n30616 ;
  assign y10605 = ~1'b0 ;
  assign y10606 = ~n30619 ;
  assign y10607 = n30625 ;
  assign y10608 = n30627 ;
  assign y10609 = ~n30629 ;
  assign y10610 = ~n30630 ;
  assign y10611 = ~n30633 ;
  assign y10612 = ~1'b0 ;
  assign y10613 = n30635 ;
  assign y10614 = ~1'b0 ;
  assign y10615 = ~n16536 ;
  assign y10616 = n30636 ;
  assign y10617 = n30640 ;
  assign y10618 = n30641 ;
  assign y10619 = ~n30642 ;
  assign y10620 = n30643 ;
  assign y10621 = ~1'b0 ;
  assign y10622 = ~n30646 ;
  assign y10623 = n30649 ;
  assign y10624 = ~n30651 ;
  assign y10625 = ~1'b0 ;
  assign y10626 = ~n30652 ;
  assign y10627 = n30653 ;
  assign y10628 = n30654 ;
  assign y10629 = n30657 ;
  assign y10630 = ~n30658 ;
  assign y10631 = n30659 ;
  assign y10632 = ~n30661 ;
  assign y10633 = ~n30663 ;
  assign y10634 = n30666 ;
  assign y10635 = n30668 ;
  assign y10636 = ~1'b0 ;
  assign y10637 = ~n30669 ;
  assign y10638 = n30671 ;
  assign y10639 = ~n30678 ;
  assign y10640 = n30681 ;
  assign y10641 = ~n30683 ;
  assign y10642 = ~n30685 ;
  assign y10643 = n30687 ;
  assign y10644 = ~n30688 ;
  assign y10645 = ~n30693 ;
  assign y10646 = ~n30695 ;
  assign y10647 = ~n30698 ;
  assign y10648 = n30701 ;
  assign y10649 = n30704 ;
  assign y10650 = n30707 ;
  assign y10651 = n30709 ;
  assign y10652 = n30710 ;
  assign y10653 = ~n30712 ;
  assign y10654 = ~1'b0 ;
  assign y10655 = n30714 ;
  assign y10656 = n30716 ;
  assign y10657 = ~1'b0 ;
  assign y10658 = ~n30719 ;
  assign y10659 = n30720 ;
  assign y10660 = n30726 ;
  assign y10661 = n30727 ;
  assign y10662 = n30729 ;
  assign y10663 = n30733 ;
  assign y10664 = n30736 ;
  assign y10665 = n30738 ;
  assign y10666 = n30741 ;
  assign y10667 = ~n30743 ;
  assign y10668 = n30750 ;
  assign y10669 = n30751 ;
  assign y10670 = n30752 ;
  assign y10671 = n30756 ;
  assign y10672 = ~n30757 ;
  assign y10673 = n30763 ;
  assign y10674 = n30764 ;
  assign y10675 = n30766 ;
  assign y10676 = ~n30770 ;
  assign y10677 = ~1'b0 ;
  assign y10678 = ~n30772 ;
  assign y10679 = ~n30775 ;
  assign y10680 = n30781 ;
  assign y10681 = ~n30782 ;
  assign y10682 = ~n30784 ;
  assign y10683 = ~n30785 ;
  assign y10684 = n30786 ;
  assign y10685 = ~n30788 ;
  assign y10686 = n30793 ;
  assign y10687 = n30794 ;
  assign y10688 = n30795 ;
  assign y10689 = ~n30803 ;
  assign y10690 = n30804 ;
  assign y10691 = ~n30807 ;
  assign y10692 = n30813 ;
  assign y10693 = ~n30814 ;
  assign y10694 = ~n30817 ;
  assign y10695 = n30819 ;
  assign y10696 = n30822 ;
  assign y10697 = n30826 ;
  assign y10698 = ~1'b0 ;
  assign y10699 = n30828 ;
  assign y10700 = n30830 ;
  assign y10701 = n30831 ;
  assign y10702 = ~n30835 ;
  assign y10703 = ~n30836 ;
  assign y10704 = ~n30837 ;
  assign y10705 = n30841 ;
  assign y10706 = ~n30842 ;
  assign y10707 = n30843 ;
  assign y10708 = n30845 ;
  assign y10709 = ~1'b0 ;
  assign y10710 = ~1'b0 ;
  assign y10711 = 1'b0 ;
  assign y10712 = ~n30846 ;
  assign y10713 = n30850 ;
  assign y10714 = n30851 ;
  assign y10715 = ~n30854 ;
  assign y10716 = n30855 ;
  assign y10717 = ~n30860 ;
  assign y10718 = n30861 ;
  assign y10719 = ~1'b0 ;
  assign y10720 = ~n30863 ;
  assign y10721 = n30864 ;
  assign y10722 = ~n30865 ;
  assign y10723 = ~n30866 ;
  assign y10724 = n30869 ;
  assign y10725 = ~n30871 ;
  assign y10726 = ~n30872 ;
  assign y10727 = n30873 ;
  assign y10728 = n30876 ;
  assign y10729 = ~1'b0 ;
  assign y10730 = n30879 ;
  assign y10731 = ~n30880 ;
  assign y10732 = n30881 ;
  assign y10733 = ~n30885 ;
  assign y10734 = ~n28939 ;
  assign y10735 = n30889 ;
  assign y10736 = n30892 ;
  assign y10737 = n30896 ;
  assign y10738 = n30901 ;
  assign y10739 = ~n30902 ;
  assign y10740 = ~n30905 ;
  assign y10741 = ~n30909 ;
  assign y10742 = ~n30914 ;
  assign y10743 = ~n30915 ;
  assign y10744 = ~1'b0 ;
  assign y10745 = ~n30920 ;
  assign y10746 = n30923 ;
  assign y10747 = ~n30929 ;
  assign y10748 = ~n30934 ;
  assign y10749 = ~n30935 ;
  assign y10750 = ~n30936 ;
  assign y10751 = ~1'b0 ;
  assign y10752 = ~n30938 ;
  assign y10753 = ~n30940 ;
  assign y10754 = ~n30942 ;
  assign y10755 = n30944 ;
  assign y10756 = n30945 ;
  assign y10757 = ~n30946 ;
  assign y10758 = ~n30948 ;
  assign y10759 = ~n30949 ;
  assign y10760 = ~n30951 ;
  assign y10761 = n30954 ;
  assign y10762 = n30957 ;
  assign y10763 = ~1'b0 ;
  assign y10764 = ~1'b0 ;
  assign y10765 = n30960 ;
  assign y10766 = ~1'b0 ;
  assign y10767 = ~n30963 ;
  assign y10768 = n30965 ;
  assign y10769 = ~1'b0 ;
  assign y10770 = ~n30968 ;
  assign y10771 = ~n30970 ;
  assign y10772 = ~n30974 ;
  assign y10773 = ~1'b0 ;
  assign y10774 = ~1'b0 ;
  assign y10775 = n30975 ;
  assign y10776 = n30976 ;
  assign y10777 = n30977 ;
  assign y10778 = n30980 ;
  assign y10779 = ~n30982 ;
  assign y10780 = ~n30983 ;
  assign y10781 = ~n30984 ;
  assign y10782 = n30990 ;
  assign y10783 = n30991 ;
  assign y10784 = ~1'b0 ;
  assign y10785 = ~n30995 ;
  assign y10786 = n30997 ;
  assign y10787 = ~1'b0 ;
  assign y10788 = ~n30998 ;
  assign y10789 = ~n31000 ;
  assign y10790 = n31001 ;
  assign y10791 = ~n31002 ;
  assign y10792 = ~n31004 ;
  assign y10793 = n31007 ;
  assign y10794 = ~1'b0 ;
  assign y10795 = n31009 ;
  assign y10796 = n31011 ;
  assign y10797 = n31014 ;
  assign y10798 = ~1'b0 ;
  assign y10799 = ~n31015 ;
  assign y10800 = n31020 ;
  assign y10801 = n31023 ;
  assign y10802 = n31026 ;
  assign y10803 = ~n31030 ;
  assign y10804 = ~n31033 ;
  assign y10805 = ~1'b0 ;
  assign y10806 = ~n31035 ;
  assign y10807 = ~n31036 ;
  assign y10808 = ~n31043 ;
  assign y10809 = n31045 ;
  assign y10810 = n31046 ;
  assign y10811 = ~n31047 ;
  assign y10812 = ~n31050 ;
  assign y10813 = n31055 ;
  assign y10814 = ~n31056 ;
  assign y10815 = n31063 ;
  assign y10816 = n31068 ;
  assign y10817 = n31069 ;
  assign y10818 = ~n31071 ;
  assign y10819 = n31074 ;
  assign y10820 = n31077 ;
  assign y10821 = ~n31079 ;
  assign y10822 = n31082 ;
  assign y10823 = ~n31083 ;
  assign y10824 = ~n31084 ;
  assign y10825 = n31086 ;
  assign y10826 = ~n31089 ;
  assign y10827 = ~n31093 ;
  assign y10828 = ~n31099 ;
  assign y10829 = ~n31100 ;
  assign y10830 = ~n31102 ;
  assign y10831 = n31104 ;
  assign y10832 = n31106 ;
  assign y10833 = n31107 ;
  assign y10834 = ~n31110 ;
  assign y10835 = ~n31112 ;
  assign y10836 = n31114 ;
  assign y10837 = n31119 ;
  assign y10838 = ~1'b0 ;
  assign y10839 = n2541 ;
  assign y10840 = ~n31125 ;
  assign y10841 = ~n31126 ;
  assign y10842 = ~n31127 ;
  assign y10843 = n31131 ;
  assign y10844 = ~n31134 ;
  assign y10845 = ~n31136 ;
  assign y10846 = n31140 ;
  assign y10847 = ~1'b0 ;
  assign y10848 = ~n31144 ;
  assign y10849 = ~n31149 ;
  assign y10850 = ~n31156 ;
  assign y10851 = n31157 ;
  assign y10852 = ~n31160 ;
  assign y10853 = n31169 ;
  assign y10854 = ~n31170 ;
  assign y10855 = ~n31173 ;
  assign y10856 = n31177 ;
  assign y10857 = ~n31179 ;
  assign y10858 = n31185 ;
  assign y10859 = ~n31186 ;
  assign y10860 = ~1'b0 ;
  assign y10861 = ~n31188 ;
  assign y10862 = ~n31189 ;
  assign y10863 = n31193 ;
  assign y10864 = ~n31194 ;
  assign y10865 = n31196 ;
  assign y10866 = ~n31198 ;
  assign y10867 = ~n31199 ;
  assign y10868 = ~n31201 ;
  assign y10869 = n31203 ;
  assign y10870 = n31205 ;
  assign y10871 = n31206 ;
  assign y10872 = ~n31207 ;
  assign y10873 = n31208 ;
  assign y10874 = ~n31209 ;
  assign y10875 = ~n31211 ;
  assign y10876 = ~n31213 ;
  assign y10877 = n31215 ;
  assign y10878 = n31218 ;
  assign y10879 = ~n31219 ;
  assign y10880 = ~n31225 ;
  assign y10881 = ~n31227 ;
  assign y10882 = ~n31229 ;
  assign y10883 = n31230 ;
  assign y10884 = ~n31231 ;
  assign y10885 = ~n31233 ;
  assign y10886 = ~n31234 ;
  assign y10887 = n31238 ;
  assign y10888 = ~n31242 ;
  assign y10889 = ~n6934 ;
  assign y10890 = n31244 ;
  assign y10891 = ~n31246 ;
  assign y10892 = n31248 ;
  assign y10893 = ~1'b0 ;
  assign y10894 = ~n31250 ;
  assign y10895 = ~n31251 ;
  assign y10896 = n31252 ;
  assign y10897 = ~n31253 ;
  assign y10898 = n31256 ;
  assign y10899 = ~n31257 ;
  assign y10900 = n31259 ;
  assign y10901 = ~1'b0 ;
  assign y10902 = ~n31264 ;
  assign y10903 = ~1'b0 ;
  assign y10904 = ~n31268 ;
  assign y10905 = ~n31269 ;
  assign y10906 = ~n31274 ;
  assign y10907 = n31276 ;
  assign y10908 = ~n31278 ;
  assign y10909 = ~n31279 ;
  assign y10910 = ~n31283 ;
  assign y10911 = ~n31285 ;
  assign y10912 = ~n31286 ;
  assign y10913 = ~n31289 ;
  assign y10914 = n31291 ;
  assign y10915 = n31295 ;
  assign y10916 = ~n31297 ;
  assign y10917 = ~n31298 ;
  assign y10918 = n31299 ;
  assign y10919 = ~n31301 ;
  assign y10920 = n31304 ;
  assign y10921 = ~n31305 ;
  assign y10922 = n31307 ;
  assign y10923 = ~n31311 ;
  assign y10924 = ~1'b0 ;
  assign y10925 = n31313 ;
  assign y10926 = n31317 ;
  assign y10927 = n31318 ;
  assign y10928 = ~n31320 ;
  assign y10929 = ~n31321 ;
  assign y10930 = ~n31324 ;
  assign y10931 = n31327 ;
  assign y10932 = n31330 ;
  assign y10933 = ~n31336 ;
  assign y10934 = ~1'b0 ;
  assign y10935 = ~n31338 ;
  assign y10936 = ~n31342 ;
  assign y10937 = ~n31348 ;
  assign y10938 = n31349 ;
  assign y10939 = ~n31355 ;
  assign y10940 = n31360 ;
  assign y10941 = n31366 ;
  assign y10942 = n31372 ;
  assign y10943 = n31378 ;
  assign y10944 = ~n31379 ;
  assign y10945 = ~n31384 ;
  assign y10946 = ~n31388 ;
  assign y10947 = ~1'b0 ;
  assign y10948 = n31393 ;
  assign y10949 = ~n147 ;
  assign y10950 = n31397 ;
  assign y10951 = ~n31398 ;
  assign y10952 = ~n31399 ;
  assign y10953 = n31400 ;
  assign y10954 = ~n31405 ;
  assign y10955 = ~1'b0 ;
  assign y10956 = ~n31408 ;
  assign y10957 = ~n31411 ;
  assign y10958 = ~1'b0 ;
  assign y10959 = ~n31415 ;
  assign y10960 = ~n31419 ;
  assign y10961 = ~n31423 ;
  assign y10962 = n31424 ;
  assign y10963 = n31427 ;
  assign y10964 = ~n31428 ;
  assign y10965 = ~1'b0 ;
  assign y10966 = n31429 ;
  assign y10967 = ~n31432 ;
  assign y10968 = ~1'b0 ;
  assign y10969 = ~n31435 ;
  assign y10970 = n31439 ;
  assign y10971 = n31441 ;
  assign y10972 = ~n31442 ;
  assign y10973 = n31445 ;
  assign y10974 = n31447 ;
  assign y10975 = n31453 ;
  assign y10976 = n31458 ;
  assign y10977 = n31464 ;
  assign y10978 = n31468 ;
  assign y10979 = n31471 ;
  assign y10980 = ~n31473 ;
endmodule
