module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 ;
  wire n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10951 , n10952 , n10953 ;
  assign n25 = x21 & x22 ;
  assign n26 = ~x1 & ~x2 ;
  assign n27 = ~x0 & n26 ;
  assign n28 = ~x3 & n27 ;
  assign n29 = ~x4 & n28 ;
  assign n30 = ~x5 & n29 ;
  assign n31 = ~x6 & n30 ;
  assign n32 = ~x7 & n31 ;
  assign n33 = ~x8 & n32 ;
  assign n34 = ~x9 & n33 ;
  assign n35 = ~x10 & n34 ;
  assign n36 = ~x11 & n35 ;
  assign n37 = ~x12 & n36 ;
  assign n38 = ~x13 & n37 ;
  assign n39 = ~x14 & n38 ;
  assign n40 = ~x15 & n39 ;
  assign n41 = ~x16 & n40 ;
  assign n42 = ~x17 & n41 ;
  assign n43 = ~x18 & n42 ;
  assign n44 = ~x19 & n43 ;
  assign n45 = ~x20 & n44 ;
  assign n46 = ~x21 & n45 ;
  assign n47 = x21 & ~n45 ;
  assign n48 = ~n46 & ~n47 ;
  assign n49 = ~x22 & n48 ;
  assign n50 = ~n25 & ~n49 ;
  assign n51 = x20 & x22 ;
  assign n52 = x20 & ~n44 ;
  assign n53 = ~n45 & ~n52 ;
  assign n54 = ~x22 & n53 ;
  assign n55 = ~n51 & ~n54 ;
  assign n56 = n50 & n55 ;
  assign n57 = x15 & x22 ;
  assign n58 = ~x22 & ~n40 ;
  assign n59 = x15 & ~n39 ;
  assign n60 = n58 & ~n59 ;
  assign n61 = ~n57 & ~n60 ;
  assign n62 = n56 & n61 ;
  assign n63 = ~x22 & ~n43 ;
  assign n64 = x19 & ~n63 ;
  assign n65 = ~x19 & n63 ;
  assign n66 = ~n64 & ~n65 ;
  assign n67 = x18 & x22 ;
  assign n68 = x18 & ~n42 ;
  assign n69 = n63 & ~n68 ;
  assign n70 = ~n67 & ~n69 ;
  assign n71 = ~n66 & ~n70 ;
  assign n72 = ~x22 & ~n41 ;
  assign n73 = x17 & ~n72 ;
  assign n74 = ~x17 & n72 ;
  assign n75 = ~n73 & ~n74 ;
  assign n76 = x16 & ~n58 ;
  assign n77 = ~x16 & n58 ;
  assign n78 = ~n76 & ~n77 ;
  assign n79 = ~n75 & n78 ;
  assign n80 = n71 & n79 ;
  assign n81 = n62 & n80 ;
  assign n82 = n75 & n78 ;
  assign n83 = n71 & n82 ;
  assign n84 = n50 & ~n55 ;
  assign n85 = n61 & n84 ;
  assign n86 = n83 & n85 ;
  assign n87 = ~n66 & n70 ;
  assign n88 = n82 & n87 ;
  assign n89 = n85 & n88 ;
  assign n90 = ~n61 & n84 ;
  assign n91 = n66 & ~n70 ;
  assign n92 = n82 & n91 ;
  assign n93 = n90 & n92 ;
  assign n94 = ~n50 & n55 ;
  assign n95 = ~n61 & n94 ;
  assign n96 = n75 & ~n78 ;
  assign n97 = n87 & n96 ;
  assign n98 = n95 & n97 ;
  assign n99 = ~n50 & ~n55 ;
  assign n100 = ~n61 & n99 ;
  assign n101 = n79 & n87 ;
  assign n102 = n100 & n101 ;
  assign n103 = n61 & n99 ;
  assign n104 = n80 & n103 ;
  assign n105 = n56 & ~n61 ;
  assign n106 = n79 & n91 ;
  assign n107 = n105 & n106 ;
  assign n108 = n80 & n95 ;
  assign n109 = n97 & n100 ;
  assign n110 = ~n75 & ~n78 ;
  assign n111 = n91 & n110 ;
  assign n112 = n100 & n111 ;
  assign n113 = n103 & n111 ;
  assign n114 = n97 & n103 ;
  assign n115 = n103 & n106 ;
  assign n116 = ~n114 & ~n115 ;
  assign n117 = n80 & n85 ;
  assign n118 = n71 & n96 ;
  assign n119 = n103 & n118 ;
  assign n120 = ~n117 & ~n119 ;
  assign n121 = n80 & n90 ;
  assign n122 = n91 & n96 ;
  assign n123 = n85 & n122 ;
  assign n124 = ~n121 & ~n123 ;
  assign n125 = n101 & n103 ;
  assign n126 = n87 & n110 ;
  assign n127 = n103 & n126 ;
  assign n128 = ~n125 & ~n127 ;
  assign n129 = n105 & n111 ;
  assign n130 = n80 & n100 ;
  assign n131 = ~n129 & ~n130 ;
  assign n132 = n128 & n131 ;
  assign n133 = n124 & n132 ;
  assign n134 = n120 & n133 ;
  assign n135 = n116 & n134 ;
  assign n136 = ~n113 & n135 ;
  assign n137 = ~n112 & n136 ;
  assign n138 = ~n109 & n137 ;
  assign n139 = ~n108 & n138 ;
  assign n140 = ~n107 & n139 ;
  assign n141 = n85 & n118 ;
  assign n142 = n95 & n126 ;
  assign n143 = n62 & n126 ;
  assign n144 = n90 & n97 ;
  assign n145 = n66 & n70 ;
  assign n146 = n82 & n145 ;
  assign n147 = n90 & n146 ;
  assign n148 = n61 & n94 ;
  assign n149 = n126 & n148 ;
  assign n150 = n83 & n100 ;
  assign n151 = n100 & n118 ;
  assign n152 = n92 & n148 ;
  assign n153 = n83 & n103 ;
  assign n154 = ~n152 & ~n153 ;
  assign n155 = ~n151 & n154 ;
  assign n156 = ~n150 & n155 ;
  assign n157 = ~n149 & n156 ;
  assign n158 = ~n147 & n157 ;
  assign n159 = ~n144 & n158 ;
  assign n160 = ~n143 & n159 ;
  assign n161 = n83 & n95 ;
  assign n162 = n110 & n145 ;
  assign n163 = n103 & n162 ;
  assign n164 = ~n161 & ~n163 ;
  assign n165 = n85 & n126 ;
  assign n166 = n92 & n95 ;
  assign n167 = n95 & n101 ;
  assign n168 = n96 & n145 ;
  assign n169 = n100 & n168 ;
  assign n170 = n71 & n110 ;
  assign n171 = n103 & n170 ;
  assign n172 = ~n169 & ~n171 ;
  assign n173 = ~n167 & n172 ;
  assign n174 = ~n166 & n173 ;
  assign n175 = ~n165 & n174 ;
  assign n176 = n164 & n175 ;
  assign n177 = n160 & n176 ;
  assign n178 = ~n142 & n177 ;
  assign n179 = ~n141 & n178 ;
  assign n180 = n79 & n145 ;
  assign n181 = n90 & n180 ;
  assign n182 = n95 & n106 ;
  assign n183 = n103 & n122 ;
  assign n184 = ~n182 & ~n183 ;
  assign n185 = ~n181 & n184 ;
  assign n186 = n105 & n122 ;
  assign n187 = n90 & n170 ;
  assign n188 = n146 & n148 ;
  assign n189 = n100 & n146 ;
  assign n190 = n92 & n105 ;
  assign n191 = n85 & n101 ;
  assign n192 = n95 & n122 ;
  assign n193 = n83 & n148 ;
  assign n194 = n100 & n162 ;
  assign n195 = n100 & n106 ;
  assign n196 = n100 & n122 ;
  assign n197 = n103 & n168 ;
  assign n198 = n97 & n105 ;
  assign n199 = n90 & n101 ;
  assign n200 = n95 & n118 ;
  assign n201 = n80 & n148 ;
  assign n202 = n100 & n126 ;
  assign n203 = n88 & n100 ;
  assign n204 = ~n202 & ~n203 ;
  assign n205 = ~n201 & n204 ;
  assign n206 = ~n200 & n205 ;
  assign n207 = ~n199 & n206 ;
  assign n208 = ~n198 & n207 ;
  assign n209 = n90 & n162 ;
  assign n210 = n80 & n105 ;
  assign n211 = ~n209 & ~n210 ;
  assign n212 = n105 & n162 ;
  assign n213 = n105 & n180 ;
  assign n214 = ~n212 & ~n213 ;
  assign n215 = n211 & n214 ;
  assign n216 = n208 & n215 ;
  assign n217 = ~n197 & n216 ;
  assign n218 = ~n196 & n217 ;
  assign n219 = ~n195 & n218 ;
  assign n220 = ~n194 & n219 ;
  assign n221 = ~n193 & n220 ;
  assign n222 = ~n192 & n221 ;
  assign n223 = ~n191 & n222 ;
  assign n224 = ~n190 & n223 ;
  assign n225 = ~n189 & n224 ;
  assign n226 = ~n188 & n225 ;
  assign n227 = ~n187 & n226 ;
  assign n228 = ~n186 & n227 ;
  assign n229 = n148 & n168 ;
  assign n230 = n95 & n170 ;
  assign n231 = ~n229 & ~n230 ;
  assign n232 = n88 & n148 ;
  assign n233 = n62 & n168 ;
  assign n234 = ~n232 & ~n233 ;
  assign n235 = n231 & n234 ;
  assign n236 = n228 & n235 ;
  assign n237 = n185 & n236 ;
  assign n238 = n179 & n237 ;
  assign n239 = n140 & n238 ;
  assign n240 = ~n104 & n239 ;
  assign n241 = ~n102 & n240 ;
  assign n242 = ~n98 & n241 ;
  assign n243 = ~n93 & n242 ;
  assign n244 = ~n89 & n243 ;
  assign n245 = ~n86 & n244 ;
  assign n246 = ~n81 & n245 ;
  assign n247 = ~x22 & ~n29 ;
  assign n248 = x5 & ~n247 ;
  assign n249 = ~x5 & n247 ;
  assign n250 = ~n248 & ~n249 ;
  assign n251 = x4 & x22 ;
  assign n252 = x4 & ~n28 ;
  assign n253 = n247 & ~n252 ;
  assign n254 = ~n251 & ~n253 ;
  assign n255 = n250 & ~n254 ;
  assign n256 = ~n250 & n254 ;
  assign n257 = ~n255 & ~n256 ;
  assign n258 = ~x22 & ~n27 ;
  assign n259 = x3 & ~n258 ;
  assign n260 = ~x3 & n258 ;
  assign n261 = ~n259 & ~n260 ;
  assign n262 = x2 & x22 ;
  assign n263 = ~x0 & ~x1 ;
  assign n264 = x2 & ~n263 ;
  assign n265 = n258 & ~n264 ;
  assign n266 = ~n262 & ~n265 ;
  assign n267 = n261 & ~n266 ;
  assign n268 = ~n261 & n266 ;
  assign n269 = ~n267 & ~n268 ;
  assign n270 = n257 & ~n269 ;
  assign n271 = n105 & n126 ;
  assign n272 = n83 & n90 ;
  assign n273 = n88 & n90 ;
  assign n274 = n97 & n148 ;
  assign n275 = n95 & n180 ;
  assign n276 = ~n186 & ~n275 ;
  assign n277 = n90 & n106 ;
  assign n278 = ~n86 & ~n277 ;
  assign n279 = n154 & n278 ;
  assign n280 = n276 & n279 ;
  assign n281 = ~n112 & n280 ;
  assign n282 = ~n274 & n281 ;
  assign n283 = ~n166 & n282 ;
  assign n284 = ~n273 & n283 ;
  assign n285 = ~n272 & n284 ;
  assign n286 = ~n271 & n285 ;
  assign n287 = n148 & n170 ;
  assign n288 = n95 & n111 ;
  assign n289 = ~n196 & ~n288 ;
  assign n290 = n85 & n162 ;
  assign n291 = ~n89 & ~n290 ;
  assign n292 = n100 & n180 ;
  assign n293 = ~n104 & ~n292 ;
  assign n294 = ~n182 & n293 ;
  assign n295 = n291 & n294 ;
  assign n296 = n289 & n295 ;
  assign n297 = ~n287 & n296 ;
  assign n298 = ~n187 & n297 ;
  assign n299 = n62 & n146 ;
  assign n300 = ~n98 & ~n299 ;
  assign n301 = n62 & n122 ;
  assign n302 = n111 & n148 ;
  assign n303 = n103 & n180 ;
  assign n304 = n122 & n148 ;
  assign n305 = ~n303 & ~n304 ;
  assign n306 = ~n230 & n305 ;
  assign n307 = ~n302 & n306 ;
  assign n308 = ~n143 & n307 ;
  assign n309 = ~n301 & n308 ;
  assign n310 = n85 & n168 ;
  assign n311 = n88 & n95 ;
  assign n312 = n88 & n103 ;
  assign n313 = ~n163 & ~n312 ;
  assign n314 = ~n150 & n313 ;
  assign n315 = ~n311 & n314 ;
  assign n316 = ~n310 & n315 ;
  assign n317 = n83 & n105 ;
  assign n318 = n148 & n162 ;
  assign n319 = ~n317 & ~n318 ;
  assign n320 = n105 & n146 ;
  assign n321 = ~n125 & ~n320 ;
  assign n322 = n85 & n170 ;
  assign n323 = n106 & n148 ;
  assign n324 = ~n322 & ~n323 ;
  assign n325 = n101 & n148 ;
  assign n326 = n62 & n88 ;
  assign n327 = ~n167 & ~n201 ;
  assign n328 = ~n326 & n327 ;
  assign n329 = ~n192 & n328 ;
  assign n330 = ~n191 & n329 ;
  assign n331 = n85 & n146 ;
  assign n332 = n85 & n111 ;
  assign n333 = n85 & n180 ;
  assign n334 = n85 & n92 ;
  assign n335 = n95 & n162 ;
  assign n336 = n90 & n122 ;
  assign n337 = ~n335 & ~n336 ;
  assign n338 = ~n334 & n337 ;
  assign n339 = ~n333 & n338 ;
  assign n340 = ~n332 & n339 ;
  assign n341 = ~n331 & n340 ;
  assign n342 = n62 & n170 ;
  assign n343 = n62 & n101 ;
  assign n344 = ~n102 & ~n343 ;
  assign n345 = n148 & n180 ;
  assign n346 = n344 & ~n345 ;
  assign n347 = ~n342 & n346 ;
  assign n348 = ~n81 & ~n190 ;
  assign n349 = n347 & n348 ;
  assign n350 = n341 & n349 ;
  assign n351 = n330 & n350 ;
  assign n352 = ~n149 & n351 ;
  assign n353 = ~n108 & n352 ;
  assign n354 = ~n121 & n353 ;
  assign n355 = ~n198 & n354 ;
  assign n356 = n131 & n355 ;
  assign n357 = ~n325 & n356 ;
  assign n358 = n324 & n357 ;
  assign n359 = n321 & n358 ;
  assign n360 = n234 & n359 ;
  assign n361 = n319 & n360 ;
  assign n362 = n316 & n361 ;
  assign n363 = n309 & n362 ;
  assign n364 = n300 & n363 ;
  assign n365 = n298 & n364 ;
  assign n366 = n286 & n365 ;
  assign n367 = ~n183 & n366 ;
  assign n368 = ~n109 & n367 ;
  assign n369 = n100 & n170 ;
  assign n370 = ~n167 & ~n325 ;
  assign n371 = ~n149 & ~n312 ;
  assign n372 = ~n182 & ~n302 ;
  assign n373 = n371 & n372 ;
  assign n374 = n289 & n373 ;
  assign n375 = n116 & n374 ;
  assign n376 = ~n183 & n375 ;
  assign n377 = ~n203 & n376 ;
  assign n378 = n370 & n377 ;
  assign n379 = ~n142 & n378 ;
  assign n380 = n92 & n100 ;
  assign n381 = ~n112 & ~n232 ;
  assign n382 = ~n311 & n381 ;
  assign n383 = n92 & n103 ;
  assign n384 = ~n113 & ~n383 ;
  assign n385 = ~n195 & n384 ;
  assign n386 = ~n274 & n385 ;
  assign n387 = n382 & n386 ;
  assign n388 = ~n380 & n387 ;
  assign n389 = ~n98 & n388 ;
  assign n390 = n103 & n146 ;
  assign n391 = ~n230 & ~n390 ;
  assign n392 = n118 & n148 ;
  assign n393 = n128 & n164 ;
  assign n394 = ~n102 & n393 ;
  assign n395 = ~n194 & n394 ;
  assign n396 = ~n200 & n395 ;
  assign n397 = ~n392 & n396 ;
  assign n398 = ~n193 & n397 ;
  assign n399 = n391 & n398 ;
  assign n400 = n389 & n399 ;
  assign n401 = ~n197 & n400 ;
  assign n402 = ~n119 & n401 ;
  assign n403 = ~n104 & n402 ;
  assign n404 = ~n151 & n403 ;
  assign n405 = ~n189 & n404 ;
  assign n406 = ~n109 & n405 ;
  assign n407 = ~n130 & ~n169 ;
  assign n408 = ~n153 & ~n202 ;
  assign n409 = ~n150 & n408 ;
  assign n410 = ~n287 & n409 ;
  assign n411 = ~n201 & n410 ;
  assign n412 = ~n108 & n411 ;
  assign n413 = n407 & n412 ;
  assign n414 = n406 & n413 ;
  assign n415 = n379 & n414 ;
  assign n416 = ~n303 & n415 ;
  assign n417 = ~n171 & n416 ;
  assign n418 = ~n292 & n417 ;
  assign n419 = ~n369 & n418 ;
  assign n420 = n62 & n97 ;
  assign n421 = n95 & n146 ;
  assign n422 = n90 & n126 ;
  assign n423 = ~n165 & ~n422 ;
  assign n424 = n90 & n118 ;
  assign n425 = ~n272 & ~n424 ;
  assign n426 = ~n141 & n425 ;
  assign n427 = n423 & n426 ;
  assign n428 = ~n121 & n427 ;
  assign n429 = ~n229 & ~n318 ;
  assign n430 = ~n199 & n429 ;
  assign n431 = ~n187 & n430 ;
  assign n432 = ~n117 & n431 ;
  assign n433 = n95 & n168 ;
  assign n434 = ~n275 & ~n433 ;
  assign n435 = ~n335 & ~n345 ;
  assign n436 = n324 & n435 ;
  assign n437 = n434 & n436 ;
  assign n438 = n432 & n437 ;
  assign n439 = n428 & n438 ;
  assign n440 = ~n188 & n439 ;
  assign n441 = ~n421 & n440 ;
  assign n442 = ~n86 & n441 ;
  assign n443 = n88 & n105 ;
  assign n444 = n101 & n105 ;
  assign n445 = n62 & n83 ;
  assign n446 = n105 & n170 ;
  assign n447 = n62 & n118 ;
  assign n448 = ~n152 & ~n304 ;
  assign n449 = ~n210 & ~n331 ;
  assign n450 = ~n166 & ~n192 ;
  assign n451 = ~n147 & n450 ;
  assign n452 = n105 & n118 ;
  assign n453 = ~n317 & ~n452 ;
  assign n454 = n451 & n453 ;
  assign n455 = n449 & n454 ;
  assign n456 = n448 & n455 ;
  assign n457 = ~n81 & n456 ;
  assign n458 = ~n342 & n457 ;
  assign n459 = ~n447 & n458 ;
  assign n460 = ~n446 & n459 ;
  assign n461 = ~n445 & n460 ;
  assign n462 = ~n143 & n461 ;
  assign n463 = ~n271 & n462 ;
  assign n464 = ~n444 & n463 ;
  assign n465 = ~n443 & n464 ;
  assign n466 = n442 & n465 ;
  assign n467 = ~n343 & n466 ;
  assign n468 = ~n420 & n467 ;
  assign n469 = ~n198 & n468 ;
  assign n470 = n90 & n168 ;
  assign n471 = ~n93 & ~n310 ;
  assign n472 = ~n470 & n471 ;
  assign n473 = ~n333 & n472 ;
  assign n474 = ~n290 & n473 ;
  assign n475 = ~n209 & n474 ;
  assign n476 = ~n181 & n475 ;
  assign n477 = ~n334 & n476 ;
  assign n478 = n85 & n97 ;
  assign n479 = n90 & n111 ;
  assign n480 = ~n191 & ~n479 ;
  assign n481 = n85 & n106 ;
  assign n482 = ~n332 & ~n336 ;
  assign n483 = ~n481 & n482 ;
  assign n484 = n480 & n483 ;
  assign n485 = ~n277 & n484 ;
  assign n486 = ~n273 & n485 ;
  assign n487 = ~n144 & n486 ;
  assign n488 = ~n89 & n487 ;
  assign n489 = ~n478 & n488 ;
  assign n490 = n442 & n489 ;
  assign n491 = n450 & n490 ;
  assign n492 = n448 & n491 ;
  assign n493 = n477 & n492 ;
  assign n494 = ~n123 & n493 ;
  assign n495 = ~n469 & ~n494 ;
  assign n496 = x14 & x22 ;
  assign n497 = x14 & ~n38 ;
  assign n498 = ~n39 & ~n497 ;
  assign n499 = ~x22 & n498 ;
  assign n500 = ~n496 & ~n499 ;
  assign n501 = ~x22 & ~n37 ;
  assign n502 = x13 & ~n501 ;
  assign n503 = ~x13 & n501 ;
  assign n504 = ~n502 & ~n503 ;
  assign n505 = ~n500 & n504 ;
  assign n506 = n500 & ~n504 ;
  assign n507 = ~n505 & ~n506 ;
  assign n508 = n495 & n507 ;
  assign n509 = ~n495 & ~n507 ;
  assign n510 = ~n508 & ~n509 ;
  assign n511 = ~n419 & n510 ;
  assign n512 = n469 & ~n494 ;
  assign n513 = ~n469 & n494 ;
  assign n514 = ~n512 & ~n513 ;
  assign n515 = n469 & n494 ;
  assign n516 = n419 & ~n515 ;
  assign n517 = n514 & ~n516 ;
  assign n518 = ~n500 & n517 ;
  assign n519 = ~n419 & ~n495 ;
  assign n520 = ~n514 & ~n519 ;
  assign n521 = n500 & ~n519 ;
  assign n522 = ~n520 & ~n521 ;
  assign n523 = ~n518 & n522 ;
  assign n524 = ~n419 & ~n504 ;
  assign n525 = n523 & ~n524 ;
  assign n526 = ~n523 & n524 ;
  assign n527 = n62 & n111 ;
  assign n528 = n62 & n180 ;
  assign n529 = n62 & n106 ;
  assign n530 = ~n213 & ~n529 ;
  assign n531 = ~n183 & n530 ;
  assign n532 = ~n196 & n531 ;
  assign n533 = ~n342 & n532 ;
  assign n534 = ~n200 & ~n392 ;
  assign n535 = ~n271 & n534 ;
  assign n536 = ~n209 & ~n446 ;
  assign n537 = ~n212 & n536 ;
  assign n538 = ~n202 & ~n369 ;
  assign n539 = ~n102 & n538 ;
  assign n540 = n537 & n539 ;
  assign n541 = n535 & n540 ;
  assign n542 = n533 & n541 ;
  assign n543 = n160 & n542 ;
  assign n544 = ~n104 & n543 ;
  assign n545 = ~n323 & n544 ;
  assign n546 = ~n528 & n545 ;
  assign n547 = ~n142 & ~n195 ;
  assign n548 = ~n166 & n547 ;
  assign n549 = ~n312 & n548 ;
  assign n550 = ~n335 & n549 ;
  assign n551 = ~n187 & n550 ;
  assign n552 = ~n445 & n551 ;
  assign n553 = ~n93 & ~n171 ;
  assign n554 = ~n89 & n553 ;
  assign n555 = ~n478 & n554 ;
  assign n556 = ~n444 & n555 ;
  assign n557 = ~n193 & ~n318 ;
  assign n558 = ~n304 & n557 ;
  assign n559 = ~n424 & n558 ;
  assign n560 = ~n273 & ~n322 ;
  assign n561 = ~n331 & n560 ;
  assign n562 = n140 & ~n203 ;
  assign n563 = ~n334 & n562 ;
  assign n564 = n62 & n162 ;
  assign n565 = ~n161 & ~n564 ;
  assign n566 = n563 & n565 ;
  assign n567 = n561 & n566 ;
  assign n568 = n559 & n567 ;
  assign n569 = n556 & n568 ;
  assign n570 = n552 & n569 ;
  assign n571 = n546 & n570 ;
  assign n572 = n330 & n571 ;
  assign n573 = ~n527 & n572 ;
  assign n574 = n62 & n92 ;
  assign n575 = n116 & n348 ;
  assign n576 = ~n195 & n575 ;
  assign n577 = ~n109 & n576 ;
  assign n578 = ~n147 & n577 ;
  assign n579 = ~n273 & n578 ;
  assign n580 = ~n481 & n579 ;
  assign n581 = ~n529 & n580 ;
  assign n582 = ~n197 & ~n312 ;
  assign n583 = ~n89 & n582 ;
  assign n584 = ~n292 & ~n380 ;
  assign n585 = n449 & n584 ;
  assign n586 = ~n202 & n585 ;
  assign n587 = ~n323 & n586 ;
  assign n588 = ~n304 & n587 ;
  assign n589 = ~n129 & n588 ;
  assign n590 = n128 & n407 ;
  assign n591 = n480 & n590 ;
  assign n592 = n589 & n591 ;
  assign n593 = ~n383 & n592 ;
  assign n594 = ~n163 & n593 ;
  assign n595 = ~n104 & n594 ;
  assign n596 = ~n192 & n595 ;
  assign n597 = ~n332 & n596 ;
  assign n598 = ~n301 & n597 ;
  assign n599 = ~n369 & n598 ;
  assign n600 = ~n326 & n599 ;
  assign n601 = ~n183 & ~n189 ;
  assign n602 = ~n112 & n601 ;
  assign n603 = ~n144 & n602 ;
  assign n604 = n600 & n603 ;
  assign n605 = n319 & n604 ;
  assign n606 = n583 & n605 ;
  assign n607 = n581 & n606 ;
  assign n608 = ~n166 & n607 ;
  assign n609 = ~n421 & n608 ;
  assign n610 = ~n574 & n609 ;
  assign n611 = ~n186 & n610 ;
  assign n612 = ~n287 & ~n390 ;
  assign n613 = ~n151 & ~n478 ;
  assign n614 = n612 & n613 ;
  assign n615 = ~n171 & n614 ;
  assign n616 = ~n150 & n615 ;
  assign n617 = ~n275 & n616 ;
  assign n618 = ~n277 & n617 ;
  assign n619 = ~n188 & ~n447 ;
  assign n620 = ~n113 & ~n203 ;
  assign n621 = ~n452 & n620 ;
  assign n622 = ~n102 & ~n303 ;
  assign n623 = ~n345 & n622 ;
  assign n624 = n231 & n623 ;
  assign n625 = ~n119 & n624 ;
  assign n626 = ~n196 & n625 ;
  assign n627 = ~n446 & n626 ;
  assign n628 = ~n107 & n627 ;
  assign n629 = ~n194 & n628 ;
  assign n630 = ~n433 & n629 ;
  assign n631 = n154 & n630 ;
  assign n632 = n621 & n631 ;
  assign n633 = n619 & n632 ;
  assign n634 = n618 & n633 ;
  assign n635 = n611 & n634 ;
  assign n636 = n337 & n635 ;
  assign n637 = ~n527 & n636 ;
  assign n638 = ~n342 & n637 ;
  assign n639 = ~n573 & ~n638 ;
  assign n640 = ~n469 & ~n639 ;
  assign n641 = ~x22 & ~n35 ;
  assign n642 = x11 & ~n641 ;
  assign n643 = ~x11 & n641 ;
  assign n644 = ~n642 & ~n643 ;
  assign n645 = ~n419 & ~n644 ;
  assign n646 = ~n640 & n645 ;
  assign n647 = n640 & ~n645 ;
  assign n648 = ~n646 & ~n647 ;
  assign n649 = x12 & x22 ;
  assign n650 = x12 & ~n36 ;
  assign n651 = n501 & ~n650 ;
  assign n652 = ~n649 & ~n651 ;
  assign n653 = ~n419 & ~n652 ;
  assign n654 = n648 & n653 ;
  assign n655 = ~n646 & ~n654 ;
  assign n656 = ~n525 & ~n655 ;
  assign n657 = ~n526 & n656 ;
  assign n658 = ~n525 & ~n657 ;
  assign n659 = ~n514 & ~n516 ;
  assign n660 = ~n500 & n659 ;
  assign n661 = n500 & n520 ;
  assign n662 = n514 & ~n519 ;
  assign n663 = n504 & n662 ;
  assign n664 = ~n504 & n517 ;
  assign n665 = ~n663 & ~n664 ;
  assign n666 = ~n661 & n665 ;
  assign n667 = ~n660 & n666 ;
  assign n668 = n573 & ~n638 ;
  assign n669 = ~n573 & n638 ;
  assign n670 = ~n668 & ~n669 ;
  assign n671 = n573 & n638 ;
  assign n672 = n469 & ~n671 ;
  assign n673 = n670 & ~n672 ;
  assign n674 = ~n500 & n673 ;
  assign n675 = ~n640 & ~n670 ;
  assign n676 = n500 & ~n640 ;
  assign n677 = ~n675 & ~n676 ;
  assign n678 = ~n674 & n677 ;
  assign n679 = ~n645 & n678 ;
  assign n680 = ~n504 & n659 ;
  assign n681 = n504 & n520 ;
  assign n682 = n652 & n662 ;
  assign n683 = n517 & ~n652 ;
  assign n684 = ~n682 & ~n683 ;
  assign n685 = ~n681 & n684 ;
  assign n686 = ~n680 & n685 ;
  assign n687 = n645 & ~n678 ;
  assign n688 = ~n679 & ~n687 ;
  assign n689 = n686 & n688 ;
  assign n690 = ~n679 & ~n689 ;
  assign n691 = n667 & ~n690 ;
  assign n692 = ~n667 & n690 ;
  assign n693 = ~n691 & ~n692 ;
  assign n694 = ~n648 & ~n653 ;
  assign n695 = ~n654 & ~n694 ;
  assign n696 = n693 & n695 ;
  assign n697 = ~n691 & ~n696 ;
  assign n698 = ~n655 & ~n657 ;
  assign n699 = ~n526 & n658 ;
  assign n700 = ~n698 & ~n699 ;
  assign n701 = ~n697 & n700 ;
  assign n702 = n697 & ~n700 ;
  assign n703 = ~n701 & ~n702 ;
  assign n704 = ~n197 & ~n390 ;
  assign n705 = ~n194 & n704 ;
  assign n706 = ~n334 & n705 ;
  assign n707 = ~n141 & n706 ;
  assign n708 = ~n445 & n707 ;
  assign n709 = ~n343 & n708 ;
  assign n710 = ~n320 & n709 ;
  assign n711 = n105 & n168 ;
  assign n712 = ~n98 & ~n142 ;
  assign n713 = ~n191 & n712 ;
  assign n714 = ~n711 & n713 ;
  assign n715 = ~n312 & ~n470 ;
  assign n716 = ~n478 & n715 ;
  assign n717 = ~n481 & n716 ;
  assign n718 = ~n326 & n717 ;
  assign n719 = ~n210 & n718 ;
  assign n720 = n451 & n719 ;
  assign n721 = n714 & n720 ;
  assign n722 = ~n114 & n721 ;
  assign n723 = ~n479 & n722 ;
  assign n724 = ~n272 & n723 ;
  assign n725 = ~n181 & n724 ;
  assign n726 = ~n81 & n725 ;
  assign n727 = ~n213 & n726 ;
  assign n728 = ~n107 & ~n273 ;
  assign n729 = ~n323 & n620 ;
  assign n730 = ~n325 & n729 ;
  assign n731 = ~n193 & n730 ;
  assign n732 = ~n123 & n731 ;
  assign n733 = ~n152 & ~n186 ;
  assign n734 = ~n190 & n733 ;
  assign n735 = ~n187 & ~n447 ;
  assign n736 = n734 & n735 ;
  assign n737 = n732 & n736 ;
  assign n738 = n728 & n737 ;
  assign n739 = ~n163 & n738 ;
  assign n740 = ~n232 & n739 ;
  assign n741 = ~n117 & n740 ;
  assign n742 = ~n527 & n741 ;
  assign n743 = ~n420 & n742 ;
  assign n744 = ~n112 & ~n288 ;
  assign n745 = ~n422 & n744 ;
  assign n746 = ~n290 & n745 ;
  assign n747 = ~n143 & n746 ;
  assign n748 = ~n446 & n747 ;
  assign n749 = ~n189 & ~n380 ;
  assign n750 = ~n277 & n749 ;
  assign n751 = ~n229 & ~n275 ;
  assign n752 = ~n200 & n751 ;
  assign n753 = n750 & n752 ;
  assign n754 = n748 & n753 ;
  assign n755 = n743 & n754 ;
  assign n756 = n727 & n755 ;
  assign n757 = n710 & n756 ;
  assign n758 = ~n383 & n757 ;
  assign n759 = ~n201 & n758 ;
  assign n760 = ~n108 & n759 ;
  assign n761 = ~n212 & n760 ;
  assign n762 = ~n141 & ~n201 ;
  assign n763 = ~n212 & n762 ;
  assign n764 = ~n452 & n763 ;
  assign n765 = ~n144 & ~n161 ;
  assign n766 = ~n322 & n765 ;
  assign n767 = ~n198 & n766 ;
  assign n768 = ~n86 & ~n151 ;
  assign n769 = ~n445 & n768 ;
  assign n770 = ~n109 & ~n153 ;
  assign n771 = ~n187 & n770 ;
  assign n772 = n769 & n771 ;
  assign n773 = n623 & n772 ;
  assign n774 = n767 & n773 ;
  assign n775 = ~n194 & n774 ;
  assign n776 = ~n325 & n775 ;
  assign n777 = ~n392 & n776 ;
  assign n778 = ~n108 & n777 ;
  assign n779 = ~n290 & n778 ;
  assign n780 = ~n81 & n779 ;
  assign n781 = ~n200 & ~n274 ;
  assign n782 = ~n98 & ~n150 ;
  assign n783 = ~n119 & ~n311 ;
  assign n784 = ~n433 & ~n564 ;
  assign n785 = n276 & n784 ;
  assign n786 = n124 & n785 ;
  assign n787 = ~n233 & n786 ;
  assign n788 = ~n343 & n787 ;
  assign n789 = ~n272 & n788 ;
  assign n790 = ~n181 & n789 ;
  assign n791 = n600 & n790 ;
  assign n792 = n783 & n791 ;
  assign n793 = n782 & n792 ;
  assign n794 = n781 & n793 ;
  assign n795 = n780 & n794 ;
  assign n796 = n764 & n795 ;
  assign n797 = ~n147 & n796 ;
  assign n798 = n553 & n797 ;
  assign n799 = ~n333 & n798 ;
  assign n800 = ~n711 & n799 ;
  assign n801 = ~n271 & n800 ;
  assign n802 = ~n761 & ~n801 ;
  assign n803 = ~n573 & ~n802 ;
  assign n804 = ~x22 & ~n33 ;
  assign n805 = x9 & ~n804 ;
  assign n806 = ~x9 & n804 ;
  assign n807 = ~n805 & ~n806 ;
  assign n808 = ~n419 & ~n807 ;
  assign n809 = ~n803 & n808 ;
  assign n810 = n803 & ~n808 ;
  assign n811 = ~n809 & ~n810 ;
  assign n812 = x10 & x22 ;
  assign n813 = x10 & ~n34 ;
  assign n814 = n641 & ~n813 ;
  assign n815 = ~n812 & ~n814 ;
  assign n816 = ~n419 & ~n815 ;
  assign n817 = n811 & n816 ;
  assign n818 = ~n809 & ~n817 ;
  assign n819 = ~n670 & ~n672 ;
  assign n820 = ~n500 & n819 ;
  assign n821 = n500 & n675 ;
  assign n822 = ~n640 & n670 ;
  assign n823 = n504 & n822 ;
  assign n824 = ~n504 & n673 ;
  assign n825 = ~n823 & ~n824 ;
  assign n826 = ~n821 & n825 ;
  assign n827 = ~n820 & n826 ;
  assign n828 = ~n652 & n659 ;
  assign n829 = n520 & n652 ;
  assign n830 = n644 & n662 ;
  assign n831 = n517 & ~n644 ;
  assign n832 = ~n830 & ~n831 ;
  assign n833 = ~n829 & n832 ;
  assign n834 = ~n828 & n833 ;
  assign n835 = n827 & n834 ;
  assign n836 = n761 & ~n801 ;
  assign n837 = ~n761 & n801 ;
  assign n838 = ~n836 & ~n837 ;
  assign n839 = n761 & n801 ;
  assign n840 = n573 & ~n839 ;
  assign n841 = n838 & ~n840 ;
  assign n842 = ~n500 & n841 ;
  assign n843 = ~n803 & ~n838 ;
  assign n844 = n500 & ~n803 ;
  assign n845 = ~n843 & ~n844 ;
  assign n846 = ~n842 & n845 ;
  assign n847 = ~n808 & n846 ;
  assign n848 = ~n504 & n819 ;
  assign n849 = n504 & n675 ;
  assign n850 = n652 & n822 ;
  assign n851 = ~n652 & n673 ;
  assign n852 = ~n850 & ~n851 ;
  assign n853 = ~n849 & n852 ;
  assign n854 = ~n848 & n853 ;
  assign n855 = n808 & ~n846 ;
  assign n856 = ~n847 & ~n855 ;
  assign n857 = n854 & n856 ;
  assign n858 = ~n847 & ~n857 ;
  assign n859 = ~n827 & ~n834 ;
  assign n860 = ~n835 & ~n859 ;
  assign n861 = ~n858 & n860 ;
  assign n862 = ~n835 & ~n861 ;
  assign n863 = ~n818 & ~n862 ;
  assign n864 = ~n818 & ~n863 ;
  assign n865 = ~n862 & ~n863 ;
  assign n866 = ~n864 & ~n865 ;
  assign n867 = ~n686 & ~n688 ;
  assign n868 = ~n689 & ~n867 ;
  assign n869 = ~n866 & n868 ;
  assign n870 = ~n863 & ~n869 ;
  assign n871 = ~n693 & ~n695 ;
  assign n872 = ~n696 & ~n871 ;
  assign n873 = ~n870 & n872 ;
  assign n874 = ~n644 & n659 ;
  assign n875 = n520 & n644 ;
  assign n876 = n662 & n815 ;
  assign n877 = n517 & ~n815 ;
  assign n878 = ~n876 & ~n877 ;
  assign n879 = ~n875 & n878 ;
  assign n880 = ~n874 & n879 ;
  assign n881 = ~n141 & ~n421 ;
  assign n882 = n120 & n881 ;
  assign n883 = ~n527 & n882 ;
  assign n884 = ~n213 & n883 ;
  assign n885 = ~n271 & n884 ;
  assign n886 = ~n149 & ~n445 ;
  assign n887 = ~n197 & n886 ;
  assign n888 = ~n325 & n887 ;
  assign n889 = ~n320 & n888 ;
  assign n890 = n278 & n889 ;
  assign n891 = n298 & n890 ;
  assign n892 = n885 & n891 ;
  assign n893 = ~n127 & n892 ;
  assign n894 = ~n171 & n893 ;
  assign n895 = ~n161 & n894 ;
  assign n896 = ~n479 & n895 ;
  assign n897 = ~n470 & n896 ;
  assign n898 = ~n129 & n897 ;
  assign n899 = ~n345 & ~n443 ;
  assign n900 = ~n322 & n899 ;
  assign n901 = ~n420 & n900 ;
  assign n902 = ~n102 & n382 ;
  assign n903 = ~n191 & n902 ;
  assign n904 = ~n564 & n903 ;
  assign n905 = ~n342 & n904 ;
  assign n906 = ~n114 & ~n302 ;
  assign n907 = n537 & n613 ;
  assign n908 = n906 & n907 ;
  assign n909 = n905 & n908 ;
  assign n910 = n901 & n909 ;
  assign n911 = ~n194 & n910 ;
  assign n912 = ~n274 & n911 ;
  assign n913 = ~n123 & n912 ;
  assign n914 = ~n152 & ~n189 ;
  assign n915 = ~n193 & n914 ;
  assign n916 = ~n167 & n915 ;
  assign n917 = ~n108 & n916 ;
  assign n918 = ~n711 & n917 ;
  assign n919 = ~n317 & n918 ;
  assign n920 = ~n165 & ~n369 ;
  assign n921 = ~n210 & n920 ;
  assign n922 = ~n130 & ~n380 ;
  assign n923 = ~n326 & n922 ;
  assign n924 = n471 & n548 ;
  assign n925 = n923 & n924 ;
  assign n926 = n921 & n925 ;
  assign n927 = n300 & n926 ;
  assign n928 = n919 & n927 ;
  assign n929 = n913 & n928 ;
  assign n930 = n898 & n929 ;
  assign n931 = ~n275 & n930 ;
  assign n932 = ~n230 & n931 ;
  assign n933 = ~n233 & n932 ;
  assign n934 = ~n528 & n933 ;
  assign n935 = ~n144 & ~n335 ;
  assign n936 = ~n422 & n935 ;
  assign n937 = ~n130 & n936 ;
  assign n938 = ~n325 & n937 ;
  assign n939 = ~n193 & n938 ;
  assign n940 = ~n209 & n939 ;
  assign n941 = ~n334 & n940 ;
  assign n942 = ~n332 & n941 ;
  assign n943 = ~n108 & ~n232 ;
  assign n944 = ~n343 & n943 ;
  assign n945 = ~n444 & ~n446 ;
  assign n946 = n944 & n945 ;
  assign n947 = ~n119 & n946 ;
  assign n948 = ~n302 & n947 ;
  assign n949 = ~n421 & n948 ;
  assign n950 = ~n290 & n949 ;
  assign n951 = ~n165 & ~n277 ;
  assign n952 = ~n149 & n951 ;
  assign n953 = ~n166 & n952 ;
  assign n954 = ~n143 & n953 ;
  assign n955 = ~n197 & ~n383 ;
  assign n956 = ~n369 & n955 ;
  assign n957 = ~n203 & n956 ;
  assign n958 = ~n392 & n957 ;
  assign n959 = ~n104 & ~n153 ;
  assign n960 = ~n171 & n959 ;
  assign n961 = ~n424 & n960 ;
  assign n962 = n231 & n961 ;
  assign n963 = n958 & n962 ;
  assign n964 = n901 & n963 ;
  assign n965 = ~n303 & n964 ;
  assign n966 = ~n151 & n965 ;
  assign n967 = ~n195 & n966 ;
  assign n968 = ~n147 & n967 ;
  assign n969 = n762 & n968 ;
  assign n970 = ~n198 & n969 ;
  assign n971 = ~n312 & n970 ;
  assign n972 = ~n150 & n971 ;
  assign n973 = ~n527 & n972 ;
  assign n974 = ~n326 & n973 ;
  assign n975 = n954 & n974 ;
  assign n976 = n116 & n975 ;
  assign n977 = n950 & n976 ;
  assign n978 = n942 & n977 ;
  assign n979 = n589 & n978 ;
  assign n980 = ~n274 & n979 ;
  assign n981 = ~n478 & n980 ;
  assign n982 = ~n342 & n981 ;
  assign n983 = ~n934 & ~n982 ;
  assign n984 = ~n761 & ~n983 ;
  assign n985 = ~x22 & ~n31 ;
  assign n986 = x7 & ~n985 ;
  assign n987 = ~x7 & n985 ;
  assign n988 = ~n986 & ~n987 ;
  assign n989 = ~n419 & ~n988 ;
  assign n990 = ~n984 & n989 ;
  assign n991 = n984 & ~n989 ;
  assign n992 = ~n990 & ~n991 ;
  assign n993 = x8 & x22 ;
  assign n994 = x8 & ~n32 ;
  assign n995 = n804 & ~n994 ;
  assign n996 = ~n993 & ~n995 ;
  assign n997 = n992 & ~n996 ;
  assign n998 = ~n419 & n997 ;
  assign n999 = ~n990 & ~n998 ;
  assign n1000 = n880 & ~n999 ;
  assign n1001 = n659 & ~n815 ;
  assign n1002 = n520 & n815 ;
  assign n1003 = n662 & n807 ;
  assign n1004 = n517 & ~n807 ;
  assign n1005 = ~n1003 & ~n1004 ;
  assign n1006 = ~n1002 & n1005 ;
  assign n1007 = ~n1001 & n1006 ;
  assign n1008 = ~n838 & ~n840 ;
  assign n1009 = ~n500 & n1008 ;
  assign n1010 = n500 & n843 ;
  assign n1011 = ~n803 & n838 ;
  assign n1012 = n504 & n1011 ;
  assign n1013 = ~n504 & n841 ;
  assign n1014 = ~n1012 & ~n1013 ;
  assign n1015 = ~n1010 & n1014 ;
  assign n1016 = ~n1009 & n1015 ;
  assign n1017 = ~n652 & n819 ;
  assign n1018 = n652 & n675 ;
  assign n1019 = n644 & n822 ;
  assign n1020 = ~n644 & n673 ;
  assign n1021 = ~n1019 & ~n1020 ;
  assign n1022 = ~n1018 & n1021 ;
  assign n1023 = ~n1017 & n1022 ;
  assign n1024 = n1016 & ~n1023 ;
  assign n1025 = ~n1016 & n1023 ;
  assign n1026 = ~n1024 & ~n1025 ;
  assign n1027 = n1007 & ~n1026 ;
  assign n1028 = n1016 & n1023 ;
  assign n1029 = ~n1027 & ~n1028 ;
  assign n1030 = n880 & ~n1000 ;
  assign n1031 = ~n999 & ~n1000 ;
  assign n1032 = ~n1030 & ~n1031 ;
  assign n1033 = ~n1029 & ~n1032 ;
  assign n1034 = ~n1000 & ~n1033 ;
  assign n1035 = ~n811 & ~n816 ;
  assign n1036 = ~n817 & ~n1035 ;
  assign n1037 = ~n1034 & n1036 ;
  assign n1038 = n1034 & ~n1036 ;
  assign n1039 = ~n1037 & ~n1038 ;
  assign n1040 = n858 & ~n860 ;
  assign n1041 = ~n861 & ~n1040 ;
  assign n1042 = n1039 & n1041 ;
  assign n1043 = ~n1037 & ~n1042 ;
  assign n1044 = ~n866 & ~n869 ;
  assign n1045 = n868 & ~n869 ;
  assign n1046 = ~n1044 & ~n1045 ;
  assign n1047 = ~n1043 & n1046 ;
  assign n1048 = n1043 & ~n1046 ;
  assign n1049 = ~n1047 & ~n1048 ;
  assign n1050 = ~n644 & n819 ;
  assign n1051 = n644 & n675 ;
  assign n1052 = n815 & n822 ;
  assign n1053 = n673 & ~n815 ;
  assign n1054 = ~n1052 & ~n1053 ;
  assign n1055 = ~n1051 & n1054 ;
  assign n1056 = ~n1050 & n1055 ;
  assign n1057 = n659 & ~n807 ;
  assign n1058 = n520 & n807 ;
  assign n1059 = n662 & n996 ;
  assign n1060 = n517 & ~n996 ;
  assign n1061 = ~n1059 & ~n1060 ;
  assign n1062 = ~n1058 & n1061 ;
  assign n1063 = ~n1057 & n1062 ;
  assign n1064 = n1056 & n1063 ;
  assign n1065 = ~n323 & ~n470 ;
  assign n1066 = ~n310 & n1065 ;
  assign n1067 = ~n201 & ~n421 ;
  assign n1068 = ~n528 & n1067 ;
  assign n1069 = ~n150 & ~n318 ;
  assign n1070 = ~n478 & n1069 ;
  assign n1071 = ~n447 & n1070 ;
  assign n1072 = n1068 & n1071 ;
  assign n1073 = n1066 & n1072 ;
  assign n1074 = n958 & n1073 ;
  assign n1075 = n124 & n1074 ;
  assign n1076 = ~n171 & n1075 ;
  assign n1077 = ~n302 & n1076 ;
  assign n1078 = ~n187 & n1077 ;
  assign n1079 = ~n444 & n1078 ;
  assign n1080 = ~n93 & n370 ;
  assign n1081 = ~n210 & n1080 ;
  assign n1082 = n423 & n1081 ;
  assign n1083 = ~n199 & n1082 ;
  assign n1084 = n435 & ~n443 ;
  assign n1085 = ~n151 & n1084 ;
  assign n1086 = ~n189 & n1085 ;
  assign n1087 = ~n193 & n1086 ;
  assign n1088 = ~n479 & n1087 ;
  assign n1089 = ~n333 & n1088 ;
  assign n1090 = ~n320 & n1089 ;
  assign n1091 = ~n198 & ~n574 ;
  assign n1092 = ~n115 & ~n311 ;
  assign n1093 = n1091 & n1092 ;
  assign n1094 = n584 & n1093 ;
  assign n1095 = n533 & n1094 ;
  assign n1096 = n300 & n1095 ;
  assign n1097 = n1090 & n1096 ;
  assign n1098 = n1083 & n1097 ;
  assign n1099 = n286 & n1098 ;
  assign n1100 = n1079 & n1099 ;
  assign n1101 = ~n163 & n1100 ;
  assign n1102 = ~n108 & n1101 ;
  assign n1103 = ~n181 & n1102 ;
  assign n1104 = ~n141 & n1103 ;
  assign n1105 = ~n527 & n1104 ;
  assign n1106 = n434 & n1091 ;
  assign n1107 = n782 & n1106 ;
  assign n1108 = ~n195 & n1107 ;
  assign n1109 = ~n369 & n1108 ;
  assign n1110 = n621 & n923 ;
  assign n1111 = n289 & n1110 ;
  assign n1112 = n1083 & n1111 ;
  assign n1113 = n1109 & n1112 ;
  assign n1114 = ~n104 & n1113 ;
  assign n1115 = ~n171 & n1114 ;
  assign n1116 = ~n125 & n1115 ;
  assign n1117 = ~n188 & n1116 ;
  assign n1118 = ~n144 & n1117 ;
  assign n1119 = ~n290 & n1118 ;
  assign n1120 = ~n301 & n1119 ;
  assign n1121 = n612 & n886 ;
  assign n1122 = ~n169 & n1121 ;
  assign n1123 = ~n189 & n1122 ;
  assign n1124 = ~n323 & n1123 ;
  assign n1125 = ~n274 & n1124 ;
  assign n1126 = ~n527 & n1125 ;
  assign n1127 = ~n711 & n1126 ;
  assign n1128 = n535 & n944 ;
  assign n1129 = ~n299 & n1128 ;
  assign n1130 = n1127 & n1129 ;
  assign n1131 = n450 & n1130 ;
  assign n1132 = ~n142 & n1131 ;
  assign n1133 = ~n311 & n1132 ;
  assign n1134 = ~n233 & n1133 ;
  assign n1135 = ~n320 & n1134 ;
  assign n1136 = ~n129 & n1135 ;
  assign n1137 = ~n190 & n1136 ;
  assign n1138 = ~n183 & ~n383 ;
  assign n1139 = ~n117 & n1138 ;
  assign n1140 = ~n86 & n1139 ;
  assign n1141 = n735 & n1140 ;
  assign n1142 = n426 & n1141 ;
  assign n1143 = n480 & n1142 ;
  assign n1144 = n341 & n1143 ;
  assign n1145 = n116 & n1144 ;
  assign n1146 = n1137 & n1145 ;
  assign n1147 = n1120 & n1146 ;
  assign n1148 = ~n127 & n1147 ;
  assign n1149 = ~n194 & n1148 ;
  assign n1150 = ~n310 & n1149 ;
  assign n1151 = ~n1105 & ~n1150 ;
  assign n1152 = ~n934 & ~n1151 ;
  assign n1153 = n1105 & ~n1152 ;
  assign n1154 = ~n1105 & n1152 ;
  assign n1155 = x6 & x22 ;
  assign n1156 = x6 & ~n30 ;
  assign n1157 = n985 & ~n1156 ;
  assign n1158 = ~n1155 & ~n1157 ;
  assign n1159 = ~n419 & ~n1158 ;
  assign n1160 = ~n1153 & n1159 ;
  assign n1161 = ~n1154 & n1160 ;
  assign n1162 = ~n1153 & ~n1161 ;
  assign n1163 = ~n1056 & ~n1063 ;
  assign n1164 = ~n1064 & ~n1163 ;
  assign n1165 = ~n1162 & n1164 ;
  assign n1166 = ~n1064 & ~n1165 ;
  assign n1167 = n934 & ~n982 ;
  assign n1168 = ~n934 & n982 ;
  assign n1169 = ~n1167 & ~n1168 ;
  assign n1170 = n934 & n982 ;
  assign n1171 = n761 & ~n1170 ;
  assign n1172 = n1169 & ~n1171 ;
  assign n1173 = ~n500 & n1172 ;
  assign n1174 = ~n984 & ~n1169 ;
  assign n1175 = n500 & ~n984 ;
  assign n1176 = ~n1174 & ~n1175 ;
  assign n1177 = ~n1173 & n1176 ;
  assign n1178 = ~n989 & n1177 ;
  assign n1179 = ~n504 & n1008 ;
  assign n1180 = n504 & n843 ;
  assign n1181 = n652 & n1011 ;
  assign n1182 = ~n652 & n841 ;
  assign n1183 = ~n1181 & ~n1182 ;
  assign n1184 = ~n1180 & n1183 ;
  assign n1185 = ~n1179 & n1184 ;
  assign n1186 = n989 & ~n1177 ;
  assign n1187 = ~n1178 & ~n1186 ;
  assign n1188 = n1185 & n1187 ;
  assign n1189 = ~n1178 & ~n1188 ;
  assign n1190 = ~n1166 & ~n1189 ;
  assign n1191 = ~n1166 & ~n1190 ;
  assign n1192 = ~n1189 & ~n1190 ;
  assign n1193 = ~n1191 & ~n1192 ;
  assign n1194 = ~n419 & ~n998 ;
  assign n1195 = ~n996 & n1194 ;
  assign n1196 = n992 & ~n998 ;
  assign n1197 = ~n1195 & ~n1196 ;
  assign n1198 = ~n1193 & ~n1197 ;
  assign n1199 = ~n1190 & ~n1198 ;
  assign n1200 = ~n854 & ~n856 ;
  assign n1201 = ~n857 & ~n1200 ;
  assign n1202 = ~n1199 & n1201 ;
  assign n1203 = ~n1029 & ~n1033 ;
  assign n1204 = ~n1032 & ~n1033 ;
  assign n1205 = ~n1203 & ~n1204 ;
  assign n1206 = n1199 & ~n1201 ;
  assign n1207 = ~n1202 & ~n1206 ;
  assign n1208 = ~n1205 & n1207 ;
  assign n1209 = ~n1202 & ~n1208 ;
  assign n1210 = ~n1039 & ~n1041 ;
  assign n1211 = ~n1042 & ~n1210 ;
  assign n1212 = ~n1209 & n1211 ;
  assign n1213 = n1207 & ~n1208 ;
  assign n1214 = ~n1205 & ~n1208 ;
  assign n1215 = ~n1213 & ~n1214 ;
  assign n1216 = ~n1169 & ~n1171 ;
  assign n1217 = ~n500 & n1216 ;
  assign n1218 = n500 & n1174 ;
  assign n1219 = ~n984 & n1169 ;
  assign n1220 = n504 & n1219 ;
  assign n1221 = ~n504 & n1172 ;
  assign n1222 = ~n1220 & ~n1221 ;
  assign n1223 = ~n1218 & n1222 ;
  assign n1224 = ~n1217 & n1223 ;
  assign n1225 = ~n815 & n819 ;
  assign n1226 = n675 & n815 ;
  assign n1227 = n807 & n822 ;
  assign n1228 = n673 & ~n807 ;
  assign n1229 = ~n1227 & ~n1228 ;
  assign n1230 = ~n1226 & n1229 ;
  assign n1231 = ~n1225 & n1230 ;
  assign n1232 = n659 & ~n996 ;
  assign n1233 = n520 & n996 ;
  assign n1234 = n662 & n988 ;
  assign n1235 = n517 & ~n988 ;
  assign n1236 = ~n1234 & ~n1235 ;
  assign n1237 = ~n1233 & n1236 ;
  assign n1238 = ~n1232 & n1237 ;
  assign n1239 = n1231 & ~n1238 ;
  assign n1240 = ~n1231 & n1238 ;
  assign n1241 = ~n1239 & ~n1240 ;
  assign n1242 = n1224 & ~n1241 ;
  assign n1243 = n1231 & n1238 ;
  assign n1244 = ~n1242 & ~n1243 ;
  assign n1245 = ~n1185 & ~n1187 ;
  assign n1246 = ~n1188 & ~n1245 ;
  assign n1247 = ~n1244 & n1246 ;
  assign n1248 = ~n1244 & ~n1247 ;
  assign n1249 = n1246 & ~n1247 ;
  assign n1250 = ~n1248 & ~n1249 ;
  assign n1251 = n1162 & ~n1164 ;
  assign n1252 = ~n1165 & ~n1251 ;
  assign n1253 = ~n1250 & n1252 ;
  assign n1254 = ~n1247 & ~n1253 ;
  assign n1255 = n1007 & ~n1027 ;
  assign n1256 = ~n1026 & ~n1027 ;
  assign n1257 = ~n1255 & ~n1256 ;
  assign n1258 = ~n1254 & ~n1257 ;
  assign n1259 = ~n1254 & ~n1258 ;
  assign n1260 = ~n1257 & ~n1258 ;
  assign n1261 = ~n1259 & ~n1260 ;
  assign n1262 = ~n1193 & ~n1198 ;
  assign n1263 = ~n1197 & ~n1198 ;
  assign n1264 = ~n1262 & ~n1263 ;
  assign n1265 = ~n1261 & ~n1264 ;
  assign n1266 = ~n1258 & ~n1265 ;
  assign n1267 = ~n1215 & ~n1266 ;
  assign n1268 = ~n1215 & ~n1267 ;
  assign n1269 = ~n1266 & ~n1267 ;
  assign n1270 = ~n1268 & ~n1269 ;
  assign n1271 = ~n652 & n1008 ;
  assign n1272 = n652 & n843 ;
  assign n1273 = n644 & n1011 ;
  assign n1274 = ~n644 & n841 ;
  assign n1275 = ~n1273 & ~n1274 ;
  assign n1276 = ~n1272 & n1275 ;
  assign n1277 = ~n1271 & n1276 ;
  assign n1278 = ~n1154 & n1162 ;
  assign n1279 = n1159 & ~n1161 ;
  assign n1280 = ~n1278 & ~n1279 ;
  assign n1281 = n1277 & ~n1280 ;
  assign n1282 = ~n250 & ~n419 ;
  assign n1283 = ~n1105 & n1282 ;
  assign n1284 = n1105 & ~n1282 ;
  assign n1285 = n1105 & ~n1150 ;
  assign n1286 = ~n1105 & n1150 ;
  assign n1287 = ~n1285 & ~n1286 ;
  assign n1288 = n1105 & n1150 ;
  assign n1289 = n934 & ~n1288 ;
  assign n1290 = n1287 & ~n1289 ;
  assign n1291 = ~n500 & n1290 ;
  assign n1292 = ~n1152 & ~n1287 ;
  assign n1293 = n500 & ~n1152 ;
  assign n1294 = ~n1292 & ~n1293 ;
  assign n1295 = ~n1291 & n1294 ;
  assign n1296 = ~n1283 & n1295 ;
  assign n1297 = ~n1284 & n1296 ;
  assign n1298 = ~n1283 & ~n1297 ;
  assign n1299 = ~n1277 & n1280 ;
  assign n1300 = ~n1281 & ~n1299 ;
  assign n1301 = ~n1298 & n1300 ;
  assign n1302 = ~n1281 & ~n1301 ;
  assign n1303 = ~n504 & n1216 ;
  assign n1304 = n504 & n1174 ;
  assign n1305 = n652 & n1219 ;
  assign n1306 = ~n652 & n1172 ;
  assign n1307 = ~n1305 & ~n1306 ;
  assign n1308 = ~n1304 & n1307 ;
  assign n1309 = ~n1303 & n1308 ;
  assign n1310 = ~n644 & n1008 ;
  assign n1311 = n644 & n843 ;
  assign n1312 = n815 & n1011 ;
  assign n1313 = ~n815 & n841 ;
  assign n1314 = ~n1312 & ~n1313 ;
  assign n1315 = ~n1311 & n1314 ;
  assign n1316 = ~n1310 & n1315 ;
  assign n1317 = n1309 & n1316 ;
  assign n1318 = ~n807 & n819 ;
  assign n1319 = n675 & n807 ;
  assign n1320 = n822 & n996 ;
  assign n1321 = n673 & ~n996 ;
  assign n1322 = ~n1320 & ~n1321 ;
  assign n1323 = ~n1319 & n1322 ;
  assign n1324 = ~n1318 & n1323 ;
  assign n1325 = n1309 & ~n1316 ;
  assign n1326 = ~n1309 & n1316 ;
  assign n1327 = ~n1325 & ~n1326 ;
  assign n1328 = n1324 & ~n1327 ;
  assign n1329 = ~n1317 & ~n1328 ;
  assign n1330 = ~n1224 & n1241 ;
  assign n1331 = ~n1242 & ~n1330 ;
  assign n1332 = ~n1329 & n1331 ;
  assign n1333 = n659 & ~n988 ;
  assign n1334 = n520 & n988 ;
  assign n1335 = n662 & n1158 ;
  assign n1336 = n517 & ~n1158 ;
  assign n1337 = ~n1335 & ~n1336 ;
  assign n1338 = ~n1334 & n1337 ;
  assign n1339 = ~n1333 & n1338 ;
  assign n1340 = ~n254 & ~n419 ;
  assign n1341 = ~n1105 & n1340 ;
  assign n1342 = n1105 & ~n1340 ;
  assign n1343 = ~n1287 & ~n1289 ;
  assign n1344 = ~n500 & n1343 ;
  assign n1345 = n500 & n1292 ;
  assign n1346 = ~n1152 & n1287 ;
  assign n1347 = n504 & n1346 ;
  assign n1348 = ~n504 & n1290 ;
  assign n1349 = ~n1347 & ~n1348 ;
  assign n1350 = ~n1345 & n1349 ;
  assign n1351 = ~n1344 & n1350 ;
  assign n1352 = ~n1341 & n1351 ;
  assign n1353 = ~n1342 & n1352 ;
  assign n1354 = ~n1341 & ~n1353 ;
  assign n1355 = n1339 & ~n1354 ;
  assign n1356 = ~n1339 & n1354 ;
  assign n1357 = ~n1355 & ~n1356 ;
  assign n1358 = ~n815 & n1008 ;
  assign n1359 = n815 & n843 ;
  assign n1360 = n807 & n1011 ;
  assign n1361 = ~n807 & n841 ;
  assign n1362 = ~n1360 & ~n1361 ;
  assign n1363 = ~n1359 & n1362 ;
  assign n1364 = ~n1358 & n1363 ;
  assign n1365 = ~n652 & n1216 ;
  assign n1366 = n652 & n1174 ;
  assign n1367 = n644 & n1219 ;
  assign n1368 = ~n644 & n1172 ;
  assign n1369 = ~n1367 & ~n1368 ;
  assign n1370 = ~n1366 & n1369 ;
  assign n1371 = ~n1365 & n1370 ;
  assign n1372 = n1364 & n1371 ;
  assign n1373 = n819 & ~n996 ;
  assign n1374 = n675 & n996 ;
  assign n1375 = n822 & n988 ;
  assign n1376 = n673 & ~n988 ;
  assign n1377 = ~n1375 & ~n1376 ;
  assign n1378 = ~n1374 & n1377 ;
  assign n1379 = ~n1373 & n1378 ;
  assign n1380 = ~n1364 & n1371 ;
  assign n1381 = n1364 & ~n1371 ;
  assign n1382 = ~n1380 & ~n1381 ;
  assign n1383 = n1379 & ~n1382 ;
  assign n1384 = ~n1372 & ~n1383 ;
  assign n1385 = n1357 & ~n1384 ;
  assign n1386 = ~n1355 & ~n1385 ;
  assign n1387 = n1329 & ~n1331 ;
  assign n1388 = ~n1332 & ~n1387 ;
  assign n1389 = ~n1386 & n1388 ;
  assign n1390 = ~n1332 & ~n1389 ;
  assign n1391 = ~n1302 & ~n1390 ;
  assign n1392 = ~n1302 & ~n1391 ;
  assign n1393 = ~n1390 & ~n1391 ;
  assign n1394 = ~n1392 & ~n1393 ;
  assign n1395 = n1252 & ~n1253 ;
  assign n1396 = ~n1250 & ~n1253 ;
  assign n1397 = ~n1395 & ~n1396 ;
  assign n1398 = ~n1394 & ~n1397 ;
  assign n1399 = ~n1391 & ~n1398 ;
  assign n1400 = ~n1261 & n1264 ;
  assign n1401 = n1261 & ~n1264 ;
  assign n1402 = ~n1400 & ~n1401 ;
  assign n1403 = ~n1399 & ~n1402 ;
  assign n1404 = ~n1394 & ~n1398 ;
  assign n1405 = ~n1397 & ~n1398 ;
  assign n1406 = ~n1404 & ~n1405 ;
  assign n1407 = ~n1284 & n1298 ;
  assign n1408 = n1295 & ~n1297 ;
  assign n1409 = ~n1407 & ~n1408 ;
  assign n1410 = n1324 & ~n1328 ;
  assign n1411 = ~n1327 & ~n1328 ;
  assign n1412 = ~n1410 & ~n1411 ;
  assign n1413 = ~n1409 & ~n1412 ;
  assign n1414 = ~n1409 & ~n1413 ;
  assign n1415 = ~n1412 & ~n1413 ;
  assign n1416 = ~n1414 & ~n1415 ;
  assign n1417 = n659 & ~n1158 ;
  assign n1418 = n520 & n1158 ;
  assign n1419 = n250 & n662 ;
  assign n1420 = ~n250 & n517 ;
  assign n1421 = ~n1419 & ~n1420 ;
  assign n1422 = ~n1418 & n1421 ;
  assign n1423 = ~n1417 & n1422 ;
  assign n1424 = ~n261 & ~n419 ;
  assign n1425 = ~n196 & n784 ;
  assign n1426 = ~n149 & n1425 ;
  assign n1427 = ~n275 & n1426 ;
  assign n1428 = ~n98 & n1427 ;
  assign n1429 = ~n187 & n1428 ;
  assign n1430 = ~n322 & n1429 ;
  assign n1431 = ~n527 & n1430 ;
  assign n1432 = ~n528 & n1431 ;
  assign n1433 = ~n195 & ~n325 ;
  assign n1434 = ~n290 & n1433 ;
  assign n1435 = n407 & n559 ;
  assign n1436 = n1434 & n1435 ;
  assign n1437 = n943 & n1436 ;
  assign n1438 = n619 & n1437 ;
  assign n1439 = ~n312 & n1438 ;
  assign n1440 = ~n189 & n1439 ;
  assign n1441 = ~n392 & n1440 ;
  assign n1442 = ~n209 & n1441 ;
  assign n1443 = ~n342 & n1442 ;
  assign n1444 = ~n299 & ~n335 ;
  assign n1445 = ~n421 & n1444 ;
  assign n1446 = ~n147 & n1445 ;
  assign n1447 = ~n478 & n1446 ;
  assign n1448 = ~n331 & n1447 ;
  assign n1449 = ~n191 & n1448 ;
  assign n1450 = ~n317 & n1449 ;
  assign n1451 = ~n129 & n1450 ;
  assign n1452 = n348 & n1451 ;
  assign n1453 = n1443 & n1452 ;
  assign n1454 = n396 & n1453 ;
  assign n1455 = n1432 & n1454 ;
  assign n1456 = ~n153 & n1455 ;
  assign n1457 = ~n183 & n1456 ;
  assign n1458 = ~n93 & n1457 ;
  assign n1459 = ~n336 & n1458 ;
  assign n1460 = ~n233 & n1459 ;
  assign n1461 = ~n574 & n1460 ;
  assign n1462 = ~n186 & n1461 ;
  assign n1463 = ~n500 & n1462 ;
  assign n1464 = ~n1105 & ~n1463 ;
  assign n1465 = n1424 & n1464 ;
  assign n1466 = ~n504 & n1343 ;
  assign n1467 = n504 & n1292 ;
  assign n1468 = n652 & n1346 ;
  assign n1469 = ~n652 & n1290 ;
  assign n1470 = ~n1468 & ~n1469 ;
  assign n1471 = ~n1467 & n1470 ;
  assign n1472 = ~n1466 & n1471 ;
  assign n1473 = ~n1424 & ~n1464 ;
  assign n1474 = ~n1465 & ~n1473 ;
  assign n1475 = n1472 & n1474 ;
  assign n1476 = ~n1465 & ~n1475 ;
  assign n1477 = n1423 & ~n1476 ;
  assign n1478 = ~n1423 & n1476 ;
  assign n1479 = ~n1477 & ~n1478 ;
  assign n1480 = ~n807 & n1008 ;
  assign n1481 = n807 & n843 ;
  assign n1482 = n996 & n1011 ;
  assign n1483 = n841 & ~n996 ;
  assign n1484 = ~n1482 & ~n1483 ;
  assign n1485 = ~n1481 & n1484 ;
  assign n1486 = ~n1480 & n1485 ;
  assign n1487 = ~n644 & n1216 ;
  assign n1488 = n644 & n1174 ;
  assign n1489 = n815 & n1219 ;
  assign n1490 = ~n815 & n1172 ;
  assign n1491 = ~n1489 & ~n1490 ;
  assign n1492 = ~n1488 & n1491 ;
  assign n1493 = ~n1487 & n1492 ;
  assign n1494 = n1486 & n1493 ;
  assign n1495 = n819 & ~n988 ;
  assign n1496 = n675 & n988 ;
  assign n1497 = n822 & n1158 ;
  assign n1498 = n673 & ~n1158 ;
  assign n1499 = ~n1497 & ~n1498 ;
  assign n1500 = ~n1496 & n1499 ;
  assign n1501 = ~n1495 & n1500 ;
  assign n1502 = ~n1486 & n1493 ;
  assign n1503 = n1486 & ~n1493 ;
  assign n1504 = ~n1502 & ~n1503 ;
  assign n1505 = n1501 & ~n1504 ;
  assign n1506 = ~n1494 & ~n1505 ;
  assign n1507 = n1479 & ~n1506 ;
  assign n1508 = ~n1477 & ~n1507 ;
  assign n1509 = ~n1416 & ~n1508 ;
  assign n1510 = ~n1413 & ~n1509 ;
  assign n1511 = n1298 & ~n1300 ;
  assign n1512 = ~n1301 & ~n1511 ;
  assign n1513 = ~n1510 & n1512 ;
  assign n1514 = n1510 & ~n1512 ;
  assign n1515 = ~n1513 & ~n1514 ;
  assign n1516 = n1386 & ~n1388 ;
  assign n1517 = ~n1389 & ~n1516 ;
  assign n1518 = n1515 & n1517 ;
  assign n1519 = ~n1513 & ~n1518 ;
  assign n1520 = ~n1406 & ~n1519 ;
  assign n1521 = n1406 & ~n1519 ;
  assign n1522 = ~n1406 & n1519 ;
  assign n1523 = ~n1521 & ~n1522 ;
  assign n1524 = n1105 & ~n1462 ;
  assign n1525 = ~n1462 & ~n1524 ;
  assign n1526 = ~n500 & n1525 ;
  assign n1527 = n500 & n1524 ;
  assign n1528 = n504 & ~n1105 ;
  assign n1529 = n1462 & ~n1528 ;
  assign n1530 = ~n1527 & ~n1529 ;
  assign n1531 = ~n1526 & n1530 ;
  assign n1532 = ~n261 & n659 ;
  assign n1533 = n261 & ~n519 ;
  assign n1534 = ~n662 & ~n1533 ;
  assign n1535 = ~n1532 & n1534 ;
  assign n1536 = n519 & n1535 ;
  assign n1537 = n1531 & n1536 ;
  assign n1538 = ~n250 & n659 ;
  assign n1539 = n250 & n520 ;
  assign n1540 = n254 & n662 ;
  assign n1541 = ~n254 & n517 ;
  assign n1542 = ~n1540 & ~n1541 ;
  assign n1543 = ~n1539 & n1542 ;
  assign n1544 = ~n1538 & n1543 ;
  assign n1545 = n1537 & n1544 ;
  assign n1546 = ~n815 & n1216 ;
  assign n1547 = n815 & n1174 ;
  assign n1548 = n807 & n1219 ;
  assign n1549 = ~n807 & n1172 ;
  assign n1550 = ~n1548 & ~n1549 ;
  assign n1551 = ~n1547 & n1550 ;
  assign n1552 = ~n1546 & n1551 ;
  assign n1553 = ~n996 & n1008 ;
  assign n1554 = n843 & n996 ;
  assign n1555 = n988 & n1011 ;
  assign n1556 = n841 & ~n988 ;
  assign n1557 = ~n1555 & ~n1556 ;
  assign n1558 = ~n1554 & n1557 ;
  assign n1559 = ~n1553 & n1558 ;
  assign n1560 = n819 & ~n1158 ;
  assign n1561 = n675 & n1158 ;
  assign n1562 = n250 & n822 ;
  assign n1563 = ~n250 & n673 ;
  assign n1564 = ~n1562 & ~n1563 ;
  assign n1565 = ~n1561 & n1564 ;
  assign n1566 = ~n1560 & n1565 ;
  assign n1567 = n1559 & ~n1566 ;
  assign n1568 = ~n1559 & n1566 ;
  assign n1569 = ~n1567 & ~n1568 ;
  assign n1570 = n1552 & ~n1569 ;
  assign n1571 = n1559 & n1566 ;
  assign n1572 = ~n1570 & ~n1571 ;
  assign n1573 = ~n1537 & ~n1544 ;
  assign n1574 = ~n1545 & ~n1573 ;
  assign n1575 = ~n1572 & n1574 ;
  assign n1576 = ~n1545 & ~n1575 ;
  assign n1577 = ~n1342 & n1354 ;
  assign n1578 = n1351 & ~n1353 ;
  assign n1579 = ~n1577 & ~n1578 ;
  assign n1580 = n1576 & ~n1579 ;
  assign n1581 = ~n1576 & n1579 ;
  assign n1582 = ~n1580 & ~n1581 ;
  assign n1583 = n1379 & ~n1383 ;
  assign n1584 = ~n1382 & ~n1383 ;
  assign n1585 = ~n1583 & ~n1584 ;
  assign n1586 = ~n1582 & ~n1585 ;
  assign n1587 = ~n1576 & ~n1579 ;
  assign n1588 = ~n1586 & ~n1587 ;
  assign n1589 = ~n1357 & n1384 ;
  assign n1590 = ~n1385 & ~n1589 ;
  assign n1591 = ~n1588 & n1590 ;
  assign n1592 = n1416 & ~n1508 ;
  assign n1593 = ~n1416 & n1508 ;
  assign n1594 = ~n1592 & ~n1593 ;
  assign n1595 = n1588 & ~n1590 ;
  assign n1596 = ~n1591 & ~n1595 ;
  assign n1597 = ~n1594 & n1596 ;
  assign n1598 = ~n1591 & ~n1597 ;
  assign n1599 = ~n1515 & ~n1517 ;
  assign n1600 = ~n1518 & ~n1599 ;
  assign n1601 = ~n1598 & n1600 ;
  assign n1602 = ~n652 & n1343 ;
  assign n1603 = n652 & n1292 ;
  assign n1604 = n644 & n1346 ;
  assign n1605 = ~n644 & n1290 ;
  assign n1606 = ~n1604 & ~n1605 ;
  assign n1607 = ~n1603 & n1606 ;
  assign n1608 = ~n1602 & n1607 ;
  assign n1609 = ~n254 & n659 ;
  assign n1610 = n254 & n520 ;
  assign n1611 = n261 & n662 ;
  assign n1612 = ~n261 & n517 ;
  assign n1613 = ~n1611 & ~n1612 ;
  assign n1614 = ~n1610 & n1613 ;
  assign n1615 = ~n1609 & n1614 ;
  assign n1616 = n1608 & n1615 ;
  assign n1617 = ~n1531 & ~n1536 ;
  assign n1618 = ~n1537 & ~n1617 ;
  assign n1619 = ~n1608 & ~n1615 ;
  assign n1620 = ~n1616 & ~n1619 ;
  assign n1621 = n1618 & n1620 ;
  assign n1622 = ~n1616 & ~n1621 ;
  assign n1623 = ~n1472 & ~n1474 ;
  assign n1624 = ~n1475 & ~n1623 ;
  assign n1625 = ~n1622 & n1624 ;
  assign n1626 = n1622 & ~n1624 ;
  assign n1627 = ~n1625 & ~n1626 ;
  assign n1628 = n1501 & ~n1505 ;
  assign n1629 = ~n1504 & ~n1505 ;
  assign n1630 = ~n1628 & ~n1629 ;
  assign n1631 = n1627 & ~n1630 ;
  assign n1632 = ~n1625 & ~n1631 ;
  assign n1633 = ~n1479 & n1506 ;
  assign n1634 = ~n1507 & ~n1633 ;
  assign n1635 = ~n1632 & n1634 ;
  assign n1636 = n1632 & ~n1634 ;
  assign n1637 = ~n1635 & ~n1636 ;
  assign n1638 = n1582 & n1585 ;
  assign n1639 = ~n1586 & ~n1638 ;
  assign n1640 = n1637 & n1639 ;
  assign n1641 = ~n1635 & ~n1640 ;
  assign n1642 = n1594 & ~n1596 ;
  assign n1643 = ~n1597 & ~n1642 ;
  assign n1644 = ~n1641 & n1643 ;
  assign n1645 = ~n652 & n1525 ;
  assign n1646 = n652 & n1524 ;
  assign n1647 = n644 & ~n1105 ;
  assign n1648 = n1462 & ~n1647 ;
  assign n1649 = ~n1646 & ~n1648 ;
  assign n1650 = ~n1645 & n1649 ;
  assign n1651 = ~n261 & n819 ;
  assign n1652 = n261 & ~n640 ;
  assign n1653 = ~n822 & ~n1652 ;
  assign n1654 = ~n1651 & n1653 ;
  assign n1655 = n640 & n1654 ;
  assign n1656 = n1650 & n1655 ;
  assign n1657 = ~n807 & n1216 ;
  assign n1658 = n807 & n1174 ;
  assign n1659 = n996 & n1219 ;
  assign n1660 = ~n996 & n1172 ;
  assign n1661 = ~n1659 & ~n1660 ;
  assign n1662 = ~n1658 & n1661 ;
  assign n1663 = ~n1657 & n1662 ;
  assign n1664 = ~n988 & n1008 ;
  assign n1665 = n843 & n988 ;
  assign n1666 = n1011 & n1158 ;
  assign n1667 = n841 & ~n1158 ;
  assign n1668 = ~n1666 & ~n1667 ;
  assign n1669 = ~n1665 & n1668 ;
  assign n1670 = ~n1664 & n1669 ;
  assign n1671 = n1663 & ~n1670 ;
  assign n1672 = ~n1663 & n1670 ;
  assign n1673 = ~n1671 & ~n1672 ;
  assign n1674 = n1656 & ~n1673 ;
  assign n1675 = n1663 & n1670 ;
  assign n1676 = ~n1674 & ~n1675 ;
  assign n1677 = ~n250 & n819 ;
  assign n1678 = n250 & n675 ;
  assign n1679 = n254 & n822 ;
  assign n1680 = ~n254 & n673 ;
  assign n1681 = ~n1679 & ~n1680 ;
  assign n1682 = ~n1678 & n1681 ;
  assign n1683 = ~n1677 & n1682 ;
  assign n1684 = ~n504 & n1525 ;
  assign n1685 = n504 & n1524 ;
  assign n1686 = n652 & ~n1105 ;
  assign n1687 = n1462 & ~n1686 ;
  assign n1688 = ~n1685 & ~n1687 ;
  assign n1689 = ~n1684 & n1688 ;
  assign n1690 = ~n644 & n1343 ;
  assign n1691 = n644 & n1292 ;
  assign n1692 = n815 & n1346 ;
  assign n1693 = ~n815 & n1290 ;
  assign n1694 = ~n1692 & ~n1693 ;
  assign n1695 = ~n1691 & n1694 ;
  assign n1696 = ~n1690 & n1695 ;
  assign n1697 = n1689 & ~n1696 ;
  assign n1698 = ~n1689 & n1696 ;
  assign n1699 = ~n1697 & ~n1698 ;
  assign n1700 = n1683 & ~n1699 ;
  assign n1701 = n1689 & n1696 ;
  assign n1702 = ~n1700 & ~n1701 ;
  assign n1703 = ~n1676 & ~n1702 ;
  assign n1704 = ~n1676 & ~n1703 ;
  assign n1705 = ~n1702 & ~n1703 ;
  assign n1706 = ~n1704 & ~n1705 ;
  assign n1707 = n1552 & ~n1570 ;
  assign n1708 = ~n1569 & ~n1570 ;
  assign n1709 = ~n1707 & ~n1708 ;
  assign n1710 = ~n1706 & ~n1709 ;
  assign n1711 = ~n1703 & ~n1710 ;
  assign n1712 = n1572 & ~n1574 ;
  assign n1713 = ~n1575 & ~n1712 ;
  assign n1714 = ~n1711 & n1713 ;
  assign n1715 = n1627 & ~n1631 ;
  assign n1716 = ~n1630 & ~n1631 ;
  assign n1717 = ~n1715 & ~n1716 ;
  assign n1718 = n1711 & ~n1713 ;
  assign n1719 = ~n1714 & ~n1718 ;
  assign n1720 = ~n1717 & n1719 ;
  assign n1721 = ~n1714 & ~n1720 ;
  assign n1722 = ~n1637 & ~n1639 ;
  assign n1723 = ~n1640 & ~n1722 ;
  assign n1724 = ~n1721 & n1723 ;
  assign n1725 = ~n519 & ~n1535 ;
  assign n1726 = ~n996 & n1216 ;
  assign n1727 = n996 & n1174 ;
  assign n1728 = n988 & n1219 ;
  assign n1729 = ~n988 & n1172 ;
  assign n1730 = ~n1728 & ~n1729 ;
  assign n1731 = ~n1727 & n1730 ;
  assign n1732 = ~n1726 & n1731 ;
  assign n1733 = ~n815 & n1343 ;
  assign n1734 = n815 & n1292 ;
  assign n1735 = n807 & n1346 ;
  assign n1736 = ~n807 & n1290 ;
  assign n1737 = ~n1735 & ~n1736 ;
  assign n1738 = ~n1734 & n1737 ;
  assign n1739 = ~n1733 & n1738 ;
  assign n1740 = n1008 & ~n1158 ;
  assign n1741 = n843 & n1158 ;
  assign n1742 = n250 & n1011 ;
  assign n1743 = ~n250 & n841 ;
  assign n1744 = ~n1742 & ~n1743 ;
  assign n1745 = ~n1741 & n1744 ;
  assign n1746 = ~n1740 & n1745 ;
  assign n1747 = n1739 & ~n1746 ;
  assign n1748 = ~n1739 & n1746 ;
  assign n1749 = ~n1747 & ~n1748 ;
  assign n1750 = n1732 & ~n1749 ;
  assign n1751 = n1739 & n1746 ;
  assign n1752 = ~n1750 & ~n1751 ;
  assign n1753 = ~n1536 & ~n1752 ;
  assign n1754 = ~n1725 & n1753 ;
  assign n1755 = ~n1536 & ~n1754 ;
  assign n1756 = ~n1725 & n1755 ;
  assign n1757 = ~n1752 & ~n1754 ;
  assign n1758 = ~n1756 & ~n1757 ;
  assign n1759 = ~n1656 & n1673 ;
  assign n1760 = ~n1674 & ~n1759 ;
  assign n1761 = ~n1758 & n1760 ;
  assign n1762 = ~n1754 & ~n1761 ;
  assign n1763 = n1618 & ~n1621 ;
  assign n1764 = ~n1619 & n1622 ;
  assign n1765 = ~n1763 & ~n1764 ;
  assign n1766 = ~n1762 & n1765 ;
  assign n1767 = n1762 & ~n1765 ;
  assign n1768 = ~n1766 & ~n1767 ;
  assign n1769 = ~n1706 & ~n1710 ;
  assign n1770 = ~n1709 & ~n1710 ;
  assign n1771 = ~n1769 & ~n1770 ;
  assign n1772 = ~n1768 & ~n1771 ;
  assign n1773 = ~n1762 & ~n1765 ;
  assign n1774 = ~n1772 & ~n1773 ;
  assign n1775 = n1717 & ~n1719 ;
  assign n1776 = ~n1720 & ~n1775 ;
  assign n1777 = ~n1774 & n1776 ;
  assign n1778 = ~n644 & n1525 ;
  assign n1779 = n644 & n1524 ;
  assign n1780 = n815 & ~n1105 ;
  assign n1781 = n1462 & ~n1780 ;
  assign n1782 = ~n1779 & ~n1781 ;
  assign n1783 = ~n1778 & n1782 ;
  assign n1784 = ~n807 & n1343 ;
  assign n1785 = n807 & n1292 ;
  assign n1786 = n996 & n1346 ;
  assign n1787 = ~n996 & n1290 ;
  assign n1788 = ~n1786 & ~n1787 ;
  assign n1789 = ~n1785 & n1788 ;
  assign n1790 = ~n1784 & n1789 ;
  assign n1791 = n1783 & n1790 ;
  assign n1792 = ~n988 & n1216 ;
  assign n1793 = n988 & n1174 ;
  assign n1794 = n1158 & n1219 ;
  assign n1795 = ~n1158 & n1172 ;
  assign n1796 = ~n1794 & ~n1795 ;
  assign n1797 = ~n1793 & n1796 ;
  assign n1798 = ~n1792 & n1797 ;
  assign n1799 = n1783 & ~n1790 ;
  assign n1800 = ~n1783 & n1790 ;
  assign n1801 = ~n1799 & ~n1800 ;
  assign n1802 = n1798 & ~n1801 ;
  assign n1803 = ~n1791 & ~n1802 ;
  assign n1804 = ~n254 & n819 ;
  assign n1805 = n254 & n675 ;
  assign n1806 = n261 & n822 ;
  assign n1807 = ~n261 & n673 ;
  assign n1808 = ~n1806 & ~n1807 ;
  assign n1809 = ~n1805 & n1808 ;
  assign n1810 = ~n1804 & n1809 ;
  assign n1811 = ~n1650 & ~n1655 ;
  assign n1812 = ~n1656 & ~n1811 ;
  assign n1813 = n1810 & ~n1812 ;
  assign n1814 = ~n1810 & n1812 ;
  assign n1815 = ~n1813 & ~n1814 ;
  assign n1816 = ~n1803 & ~n1815 ;
  assign n1817 = n1810 & n1812 ;
  assign n1818 = ~n1816 & ~n1817 ;
  assign n1819 = n1683 & ~n1700 ;
  assign n1820 = ~n1699 & ~n1700 ;
  assign n1821 = ~n1819 & ~n1820 ;
  assign n1822 = ~n1818 & ~n1821 ;
  assign n1823 = ~n1758 & ~n1761 ;
  assign n1824 = n1760 & ~n1761 ;
  assign n1825 = ~n1823 & ~n1824 ;
  assign n1826 = ~n1818 & ~n1822 ;
  assign n1827 = ~n1821 & ~n1822 ;
  assign n1828 = ~n1826 & ~n1827 ;
  assign n1829 = ~n1825 & ~n1828 ;
  assign n1830 = ~n1822 & ~n1829 ;
  assign n1831 = ~n250 & n1008 ;
  assign n1832 = n250 & n843 ;
  assign n1833 = n254 & n1011 ;
  assign n1834 = ~n254 & n841 ;
  assign n1835 = ~n1833 & ~n1834 ;
  assign n1836 = ~n1832 & n1835 ;
  assign n1837 = ~n1831 & n1836 ;
  assign n1838 = ~n815 & n1525 ;
  assign n1839 = n815 & n1524 ;
  assign n1840 = n807 & ~n1105 ;
  assign n1841 = n1462 & ~n1840 ;
  assign n1842 = ~n1839 & ~n1841 ;
  assign n1843 = ~n1838 & n1842 ;
  assign n1844 = ~n261 & n1008 ;
  assign n1845 = n261 & ~n803 ;
  assign n1846 = ~n1011 & ~n1845 ;
  assign n1847 = ~n1844 & n1846 ;
  assign n1848 = n803 & n1847 ;
  assign n1849 = n1843 & n1848 ;
  assign n1850 = n1837 & n1849 ;
  assign n1851 = ~n1837 & n1849 ;
  assign n1852 = n1837 & ~n1849 ;
  assign n1853 = ~n1851 & ~n1852 ;
  assign n1854 = ~n261 & ~n670 ;
  assign n1855 = ~n1853 & n1854 ;
  assign n1856 = ~n1850 & ~n1855 ;
  assign n1857 = ~n1732 & n1749 ;
  assign n1858 = ~n1750 & ~n1857 ;
  assign n1859 = ~n1856 & n1858 ;
  assign n1860 = n1856 & ~n1858 ;
  assign n1861 = ~n1859 & ~n1860 ;
  assign n1862 = n1803 & n1815 ;
  assign n1863 = ~n1816 & ~n1862 ;
  assign n1864 = ~n1861 & ~n1863 ;
  assign n1865 = n1861 & n1863 ;
  assign n1866 = ~n254 & n1008 ;
  assign n1867 = n254 & n843 ;
  assign n1868 = n261 & n1011 ;
  assign n1869 = ~n261 & n841 ;
  assign n1870 = ~n1868 & ~n1869 ;
  assign n1871 = ~n1867 & n1870 ;
  assign n1872 = ~n1866 & n1871 ;
  assign n1873 = ~n996 & n1343 ;
  assign n1874 = n996 & n1292 ;
  assign n1875 = n988 & n1346 ;
  assign n1876 = ~n988 & n1290 ;
  assign n1877 = ~n1875 & ~n1876 ;
  assign n1878 = ~n1874 & n1877 ;
  assign n1879 = ~n1873 & n1878 ;
  assign n1880 = ~n1158 & n1216 ;
  assign n1881 = n1158 & n1174 ;
  assign n1882 = n250 & n1219 ;
  assign n1883 = ~n250 & n1172 ;
  assign n1884 = ~n1882 & ~n1883 ;
  assign n1885 = ~n1881 & n1884 ;
  assign n1886 = ~n1880 & n1885 ;
  assign n1887 = n1879 & ~n1886 ;
  assign n1888 = ~n1879 & n1886 ;
  assign n1889 = ~n1887 & ~n1888 ;
  assign n1890 = n1872 & ~n1889 ;
  assign n1891 = n1879 & n1886 ;
  assign n1892 = ~n1890 & ~n1891 ;
  assign n1893 = ~n1798 & n1801 ;
  assign n1894 = ~n1802 & ~n1893 ;
  assign n1895 = ~n1892 & n1894 ;
  assign n1896 = n1853 & ~n1854 ;
  assign n1897 = ~n1855 & ~n1896 ;
  assign n1898 = ~n1892 & ~n1895 ;
  assign n1899 = n1894 & ~n1895 ;
  assign n1900 = ~n1898 & ~n1899 ;
  assign n1901 = n1897 & ~n1900 ;
  assign n1902 = ~n1895 & ~n1901 ;
  assign n1903 = ~n803 & ~n1847 ;
  assign n1904 = ~n996 & n1525 ;
  assign n1905 = n996 & n1524 ;
  assign n1906 = n988 & ~n1105 ;
  assign n1907 = n1462 & ~n1906 ;
  assign n1908 = ~n1905 & ~n1907 ;
  assign n1909 = ~n1904 & n1908 ;
  assign n1910 = ~n261 & n1216 ;
  assign n1911 = n261 & ~n984 ;
  assign n1912 = ~n1219 & ~n1911 ;
  assign n1913 = ~n1910 & n1912 ;
  assign n1914 = n984 & n1913 ;
  assign n1915 = n1909 & n1914 ;
  assign n1916 = ~n1848 & n1915 ;
  assign n1917 = ~n1903 & n1916 ;
  assign n1918 = ~n1158 & n1343 ;
  assign n1919 = n1158 & n1292 ;
  assign n1920 = n250 & n1346 ;
  assign n1921 = ~n250 & n1290 ;
  assign n1922 = ~n1920 & ~n1921 ;
  assign n1923 = ~n1919 & n1922 ;
  assign n1924 = ~n1918 & n1923 ;
  assign n1925 = ~n254 & n1216 ;
  assign n1926 = n254 & n1174 ;
  assign n1927 = n261 & n1219 ;
  assign n1928 = ~n261 & n1172 ;
  assign n1929 = ~n1927 & ~n1928 ;
  assign n1930 = ~n1926 & n1929 ;
  assign n1931 = ~n1925 & n1930 ;
  assign n1932 = n1924 & n1931 ;
  assign n1933 = ~n1909 & ~n1914 ;
  assign n1934 = ~n1915 & ~n1933 ;
  assign n1935 = ~n1924 & ~n1931 ;
  assign n1936 = ~n1932 & ~n1935 ;
  assign n1937 = n1934 & n1936 ;
  assign n1938 = ~n1932 & ~n1937 ;
  assign n1939 = n1915 & ~n1917 ;
  assign n1940 = ~n1848 & ~n1917 ;
  assign n1941 = ~n1903 & n1940 ;
  assign n1942 = ~n1939 & ~n1941 ;
  assign n1943 = ~n1938 & ~n1942 ;
  assign n1944 = ~n1917 & ~n1943 ;
  assign n1945 = ~n250 & n1216 ;
  assign n1946 = n250 & n1174 ;
  assign n1947 = n254 & n1219 ;
  assign n1948 = ~n254 & n1172 ;
  assign n1949 = ~n1947 & ~n1948 ;
  assign n1950 = ~n1946 & n1949 ;
  assign n1951 = ~n1945 & n1950 ;
  assign n1952 = ~n988 & n1343 ;
  assign n1953 = n988 & n1292 ;
  assign n1954 = n1158 & n1346 ;
  assign n1955 = ~n1158 & n1290 ;
  assign n1956 = ~n1954 & ~n1955 ;
  assign n1957 = ~n1953 & n1956 ;
  assign n1958 = ~n1952 & n1957 ;
  assign n1959 = ~n807 & n1525 ;
  assign n1960 = n807 & n1524 ;
  assign n1961 = n996 & ~n1105 ;
  assign n1962 = n1462 & ~n1961 ;
  assign n1963 = ~n1960 & ~n1962 ;
  assign n1964 = ~n1959 & n1963 ;
  assign n1965 = ~n1958 & n1964 ;
  assign n1966 = n1958 & ~n1964 ;
  assign n1967 = ~n1965 & ~n1966 ;
  assign n1968 = ~n1951 & n1967 ;
  assign n1969 = n1951 & ~n1967 ;
  assign n1970 = ~n988 & n1525 ;
  assign n1971 = n988 & n1524 ;
  assign n1972 = ~n1105 & n1158 ;
  assign n1973 = n1462 & ~n1972 ;
  assign n1974 = ~n1971 & ~n1973 ;
  assign n1975 = ~n1970 & n1974 ;
  assign n1976 = ~n250 & n1343 ;
  assign n1977 = n250 & n1292 ;
  assign n1978 = n254 & n1346 ;
  assign n1979 = ~n254 & n1290 ;
  assign n1980 = ~n1978 & ~n1979 ;
  assign n1981 = ~n1977 & n1980 ;
  assign n1982 = ~n1976 & n1981 ;
  assign n1983 = n1975 & ~n1982 ;
  assign n1984 = ~n1975 & n1982 ;
  assign n1985 = ~n1983 & ~n1984 ;
  assign n1986 = ~n1158 & n1525 ;
  assign n1987 = n1158 & n1524 ;
  assign n1988 = n250 & ~n1105 ;
  assign n1989 = n1462 & ~n1988 ;
  assign n1990 = ~n1987 & ~n1989 ;
  assign n1991 = ~n1986 & n1990 ;
  assign n1992 = ~n261 & n1343 ;
  assign n1993 = n261 & ~n1152 ;
  assign n1994 = ~n1346 & ~n1993 ;
  assign n1995 = ~n1992 & n1994 ;
  assign n1996 = n1152 & n1995 ;
  assign n1997 = n1991 & n1996 ;
  assign n1998 = n1985 & ~n1997 ;
  assign n1999 = ~n1985 & n1997 ;
  assign n2000 = ~n254 & n1343 ;
  assign n2001 = n254 & n1292 ;
  assign n2002 = ~n261 & n1290 ;
  assign n2003 = ~n1152 & ~n1995 ;
  assign n2004 = ~n250 & n1525 ;
  assign n2005 = n250 & n1524 ;
  assign n2006 = ~n254 & ~n1462 ;
  assign n2007 = n1105 & n1462 ;
  assign n2008 = n254 & ~n2007 ;
  assign n2009 = ~n2006 & ~n2008 ;
  assign n2010 = ~n2005 & ~n2009 ;
  assign n2011 = ~n2004 & n2010 ;
  assign n2012 = n261 & ~n1105 ;
  assign n2013 = ~n2006 & n2012 ;
  assign n2014 = ~n2011 & ~n2013 ;
  assign n2015 = ~n1996 & ~n2014 ;
  assign n2016 = ~n2003 & n2015 ;
  assign n2017 = n2011 & n2013 ;
  assign n2018 = ~n2016 & ~n2017 ;
  assign n2019 = ~n1991 & ~n1996 ;
  assign n2020 = ~n1997 & ~n2019 ;
  assign n2021 = n2018 & ~n2020 ;
  assign n2022 = n261 & n1346 ;
  assign n2023 = ~n2021 & ~n2022 ;
  assign n2024 = ~n2002 & n2023 ;
  assign n2025 = ~n2001 & n2024 ;
  assign n2026 = ~n2000 & n2025 ;
  assign n2027 = ~n2018 & n2020 ;
  assign n2028 = ~n2026 & ~n2027 ;
  assign n2029 = ~n261 & ~n1169 ;
  assign n2030 = n2028 & ~n2029 ;
  assign n2031 = ~n1999 & ~n2030 ;
  assign n2032 = ~n1998 & n2031 ;
  assign n2033 = ~n2028 & n2029 ;
  assign n2034 = ~n2032 & ~n2033 ;
  assign n2035 = n1934 & ~n1937 ;
  assign n2036 = ~n1935 & n1938 ;
  assign n2037 = ~n2035 & ~n2036 ;
  assign n2038 = n2034 & n2037 ;
  assign n2039 = n1975 & n1982 ;
  assign n2040 = ~n1999 & ~n2039 ;
  assign n2041 = ~n2038 & ~n2040 ;
  assign n2042 = ~n2034 & ~n2037 ;
  assign n2043 = ~n2041 & ~n2042 ;
  assign n2044 = ~n1938 & ~n1943 ;
  assign n2045 = ~n1942 & ~n1943 ;
  assign n2046 = ~n2044 & ~n2045 ;
  assign n2047 = n2043 & n2046 ;
  assign n2048 = ~n1969 & ~n2047 ;
  assign n2049 = ~n1968 & n2048 ;
  assign n2050 = ~n2043 & ~n2046 ;
  assign n2051 = ~n2049 & ~n2050 ;
  assign n2052 = ~n1944 & ~n2051 ;
  assign n2053 = n1944 & n2051 ;
  assign n2054 = n1872 & ~n1890 ;
  assign n2055 = ~n1889 & ~n1890 ;
  assign n2056 = ~n2054 & ~n2055 ;
  assign n2057 = ~n1843 & ~n1848 ;
  assign n2058 = ~n1849 & ~n2057 ;
  assign n2059 = n1958 & n1964 ;
  assign n2060 = ~n1969 & ~n2059 ;
  assign n2061 = n2058 & ~n2060 ;
  assign n2062 = ~n2058 & n2060 ;
  assign n2063 = ~n2061 & ~n2062 ;
  assign n2064 = ~n2056 & n2063 ;
  assign n2065 = n2056 & ~n2063 ;
  assign n2066 = ~n2064 & ~n2065 ;
  assign n2067 = ~n2053 & n2066 ;
  assign n2068 = ~n2052 & ~n2067 ;
  assign n2069 = ~n2061 & ~n2064 ;
  assign n2070 = ~n2068 & ~n2069 ;
  assign n2071 = n2068 & n2069 ;
  assign n2072 = ~n1897 & n1900 ;
  assign n2073 = ~n1901 & ~n2072 ;
  assign n2074 = ~n2071 & n2073 ;
  assign n2075 = ~n2070 & ~n2074 ;
  assign n2076 = n1902 & n2075 ;
  assign n2077 = ~n1865 & ~n2076 ;
  assign n2078 = ~n1864 & n2077 ;
  assign n2079 = ~n1902 & ~n2075 ;
  assign n2080 = ~n2078 & ~n2079 ;
  assign n2081 = ~n1859 & ~n1865 ;
  assign n2082 = ~n2080 & ~n2081 ;
  assign n2083 = n2080 & n2081 ;
  assign n2084 = n1825 & n1828 ;
  assign n2085 = ~n1829 & ~n2084 ;
  assign n2086 = ~n2083 & n2085 ;
  assign n2087 = ~n2082 & ~n2086 ;
  assign n2088 = n1830 & n2087 ;
  assign n2089 = n1768 & n1771 ;
  assign n2090 = ~n2088 & ~n2089 ;
  assign n2091 = ~n1772 & n2090 ;
  assign n2092 = ~n1830 & ~n2087 ;
  assign n2093 = ~n2091 & ~n2092 ;
  assign n2094 = n1774 & ~n1776 ;
  assign n2095 = ~n1777 & ~n2094 ;
  assign n2096 = ~n2093 & n2095 ;
  assign n2097 = ~n1777 & ~n2096 ;
  assign n2098 = n1721 & ~n1723 ;
  assign n2099 = ~n1724 & ~n2098 ;
  assign n2100 = ~n2097 & n2099 ;
  assign n2101 = ~n1724 & ~n2100 ;
  assign n2102 = n1641 & ~n1643 ;
  assign n2103 = ~n1644 & ~n2102 ;
  assign n2104 = ~n2101 & n2103 ;
  assign n2105 = ~n1644 & ~n2104 ;
  assign n2106 = n1598 & ~n1600 ;
  assign n2107 = ~n1601 & ~n2106 ;
  assign n2108 = ~n2105 & n2107 ;
  assign n2109 = ~n1601 & ~n2108 ;
  assign n2110 = ~n1523 & ~n2109 ;
  assign n2111 = ~n1520 & ~n2110 ;
  assign n2112 = n1399 & n1402 ;
  assign n2113 = ~n1403 & ~n2112 ;
  assign n2114 = ~n2111 & n2113 ;
  assign n2115 = ~n1403 & ~n2114 ;
  assign n2116 = ~n1270 & ~n2115 ;
  assign n2117 = ~n1267 & ~n2116 ;
  assign n2118 = n1209 & ~n1211 ;
  assign n2119 = ~n1212 & ~n2118 ;
  assign n2120 = ~n2117 & n2119 ;
  assign n2121 = ~n1212 & ~n2120 ;
  assign n2122 = ~n1049 & ~n2121 ;
  assign n2123 = ~n1043 & ~n1046 ;
  assign n2124 = ~n2122 & ~n2123 ;
  assign n2125 = n870 & ~n872 ;
  assign n2126 = ~n873 & ~n2125 ;
  assign n2127 = ~n2124 & n2126 ;
  assign n2128 = ~n873 & ~n2127 ;
  assign n2129 = ~n703 & ~n2128 ;
  assign n2130 = ~n697 & ~n700 ;
  assign n2131 = ~n2129 & ~n2130 ;
  assign n2132 = n658 & ~n2131 ;
  assign n2133 = ~n658 & n2131 ;
  assign n2134 = ~n2132 & ~n2133 ;
  assign n2135 = n511 & n2134 ;
  assign n2136 = ~n511 & ~n2134 ;
  assign n2137 = ~n2135 & ~n2136 ;
  assign n2138 = ~n368 & ~n2137 ;
  assign n2139 = n368 & n2137 ;
  assign n2140 = ~n109 & ~n443 ;
  assign n2141 = ~n194 & n2140 ;
  assign n2142 = ~n229 & ~n304 ;
  assign n2143 = ~n333 & n2142 ;
  assign n2144 = ~n301 & n2143 ;
  assign n2145 = ~n317 & n2144 ;
  assign n2146 = n735 & n2145 ;
  assign n2147 = ~n201 & n2146 ;
  assign n2148 = ~n193 & n2147 ;
  assign n2149 = ~n142 & n2148 ;
  assign n2150 = ~n181 & n2149 ;
  assign n2151 = ~n165 & n2150 ;
  assign n2152 = ~n564 & n2151 ;
  assign n2153 = ~n711 & n2152 ;
  assign n2154 = ~n390 & n601 ;
  assign n2155 = ~n272 & n2154 ;
  assign n2156 = ~n331 & n2155 ;
  assign n2157 = ~n336 & n943 ;
  assign n2158 = ~n117 & n2157 ;
  assign n2159 = n530 & n2158 ;
  assign n2160 = n451 & n2159 ;
  assign n2161 = n1066 & n2160 ;
  assign n2162 = n2156 & n2161 ;
  assign n2163 = n961 & n2162 ;
  assign n2164 = n728 & n2163 ;
  assign n2165 = ~n129 & n2164 ;
  assign n2166 = ~n115 & n767 ;
  assign n2167 = ~n274 & n2166 ;
  assign n2168 = ~n433 & n2167 ;
  assign n2169 = ~n332 & n2168 ;
  assign n2170 = ~n123 & n2169 ;
  assign n2171 = ~n528 & n2170 ;
  assign n2172 = n128 & n783 ;
  assign n2173 = n372 & n2172 ;
  assign n2174 = n748 & n2173 ;
  assign n2175 = n2171 & n2174 ;
  assign n2176 = n2165 & n2175 ;
  assign n2177 = n2153 & n2176 ;
  assign n2178 = n2141 & n2177 ;
  assign n2179 = ~n303 & n2178 ;
  assign n2180 = ~n203 & n2179 ;
  assign n2181 = ~n152 & n2180 ;
  assign n2182 = ~n479 & n2181 ;
  assign n2183 = ~n342 & n2182 ;
  assign n2184 = ~n190 & n2183 ;
  assign n2185 = n703 & n2128 ;
  assign n2186 = ~n2129 & ~n2185 ;
  assign n2187 = ~n2184 & ~n2186 ;
  assign n2188 = n120 & n769 ;
  assign n2189 = n294 & n2188 ;
  assign n2190 = n449 & n2189 ;
  assign n2191 = n612 & n2190 ;
  assign n2192 = n714 & n2191 ;
  assign n2193 = n942 & n2192 ;
  assign n2194 = n581 & n2193 ;
  assign n2195 = n1079 & n2194 ;
  assign n2196 = ~n433 & n2195 ;
  assign n2197 = ~n272 & n2196 ;
  assign n2198 = ~n333 & n2197 ;
  assign n2199 = ~n143 & n2198 ;
  assign n2200 = ~n212 & n2199 ;
  assign n2201 = n2124 & ~n2126 ;
  assign n2202 = ~n2127 & ~n2201 ;
  assign n2203 = ~n2200 & ~n2202 ;
  assign n2204 = n2200 & n2202 ;
  assign n2205 = n306 & n2158 ;
  assign n2206 = n211 & n2205 ;
  assign n2207 = n276 & n2206 ;
  assign n2208 = n612 & n2207 ;
  assign n2209 = n2141 & n2208 ;
  assign n2210 = n330 & n2209 ;
  assign n2211 = ~n196 & n2210 ;
  assign n2212 = ~n369 & n2211 ;
  assign n2213 = ~n200 & n2212 ;
  assign n2214 = ~n181 & n2213 ;
  assign n2215 = ~n229 & n881 ;
  assign n2216 = ~n422 & n2215 ;
  assign n2217 = ~n123 & n2216 ;
  assign n2218 = ~n86 & n2217 ;
  assign n2219 = ~n213 & n2218 ;
  assign n2220 = n556 & n603 ;
  assign n2221 = n2219 & n2220 ;
  assign n2222 = ~n202 & n2221 ;
  assign n2223 = ~n392 & n2222 ;
  assign n2224 = ~n98 & n2223 ;
  assign n2225 = ~n711 & n2224 ;
  assign n2226 = ~n153 & ~n481 ;
  assign n2227 = ~n446 & n2226 ;
  assign n2228 = ~n277 & ~n288 ;
  assign n2229 = ~n420 & n2228 ;
  assign n2230 = n453 & n2229 ;
  assign n2231 = n2227 & n2230 ;
  assign n2232 = n131 & n2231 ;
  assign n2233 = n552 & n2232 ;
  assign n2234 = n619 & n2233 ;
  assign n2235 = n2225 & n2234 ;
  assign n2236 = n2214 & n2235 ;
  assign n2237 = ~n292 & n2236 ;
  assign n2238 = ~n311 & n2237 ;
  assign n2239 = ~n529 & n2238 ;
  assign n2240 = n1049 & n2121 ;
  assign n2241 = ~n2122 & ~n2240 ;
  assign n2242 = ~n2239 & ~n2241 ;
  assign n2243 = n371 & n2227 ;
  assign n2244 = n426 & n2243 ;
  assign n2245 = ~n114 & n2244 ;
  assign n2246 = ~n163 & n2245 ;
  assign n2247 = ~n104 & n2246 ;
  assign n2248 = ~n334 & n2247 ;
  assign n2249 = ~n310 & n2248 ;
  assign n2250 = ~n342 & n2249 ;
  assign n2251 = ~n574 & n2250 ;
  assign n2252 = ~n422 & ~n527 ;
  assign n2253 = ~n212 & n2252 ;
  assign n2254 = ~n127 & n2214 ;
  assign n2255 = ~n271 & n2254 ;
  assign n2256 = ~n190 & n2255 ;
  assign n2257 = n1434 & n2256 ;
  assign n2258 = n2253 & n2257 ;
  assign n2259 = n300 & n2258 ;
  assign n2260 = n2171 & n2259 ;
  assign n2261 = n2251 & n2260 ;
  assign n2262 = n955 & n2261 ;
  assign n2263 = ~n151 & n2262 ;
  assign n2264 = ~n318 & n2263 ;
  assign n2265 = ~n142 & n2264 ;
  assign n2266 = ~n335 & n2265 ;
  assign n2267 = ~n288 & n2266 ;
  assign n2268 = n2117 & ~n2119 ;
  assign n2269 = ~n2120 & ~n2268 ;
  assign n2270 = ~n2267 & ~n2269 ;
  assign n2271 = n2267 & n2269 ;
  assign n2272 = ~n113 & ~n202 ;
  assign n2273 = ~n98 & n2272 ;
  assign n2274 = ~n147 & n2273 ;
  assign n2275 = ~n209 & n2274 ;
  assign n2276 = ~n332 & n2275 ;
  assign n2277 = ~n191 & n2276 ;
  assign n2278 = ~n143 & n2277 ;
  assign n2279 = n116 & n1091 ;
  assign n2280 = n919 & n2279 ;
  assign n2281 = n619 & n2280 ;
  assign n2282 = n344 & n2281 ;
  assign n2283 = ~n312 & n2282 ;
  assign n2284 = ~n433 & n2283 ;
  assign n2285 = ~n422 & n2284 ;
  assign n2286 = ~n322 & n2285 ;
  assign n2287 = ~n81 & n898 ;
  assign n2288 = ~n301 & n2287 ;
  assign n2289 = ~n192 & ~n203 ;
  assign n2290 = ~n121 & n2289 ;
  assign n2291 = ~n186 & n2290 ;
  assign n2292 = ~n444 & n2291 ;
  assign n2293 = n2288 & n2292 ;
  assign n2294 = n2286 & n2293 ;
  assign n2295 = n2278 & n2294 ;
  assign n2296 = ~n303 & n2295 ;
  assign n2297 = ~n383 & n2296 ;
  assign n2298 = ~n169 & n2297 ;
  assign n2299 = ~n194 & n2298 ;
  assign n2300 = ~n273 & n2299 ;
  assign n2301 = n425 & n2300 ;
  assign n2302 = ~n420 & n2301 ;
  assign n2303 = n1270 & n2115 ;
  assign n2304 = ~n2116 & ~n2303 ;
  assign n2305 = ~n2302 & ~n2304 ;
  assign n2306 = ~n188 & n483 ;
  assign n2307 = ~n711 & n2306 ;
  assign n2308 = ~n320 & n2307 ;
  assign n2309 = n278 & n734 ;
  assign n2310 = n906 & n2309 ;
  assign n2311 = ~n144 & n2310 ;
  assign n2312 = ~n89 & n2311 ;
  assign n2313 = ~n301 & n2312 ;
  assign n2314 = ~n444 & n2313 ;
  assign n2315 = ~n113 & ~n121 ;
  assign n2316 = ~n81 & ~n323 ;
  assign n2317 = ~n213 & n2316 ;
  assign n2318 = n407 & n2317 ;
  assign n2319 = n2315 & n2318 ;
  assign n2320 = n1081 & n2319 ;
  assign n2321 = n319 & n2320 ;
  assign n2322 = n289 & n2321 ;
  assign n2323 = n2314 & n2322 ;
  assign n2324 = n970 & n2323 ;
  assign n2325 = n905 & n2324 ;
  assign n2326 = n2308 & n2325 ;
  assign n2327 = ~n127 & n2326 ;
  assign n2328 = ~n192 & n2327 ;
  assign n2329 = ~n470 & n2328 ;
  assign n2330 = n2111 & ~n2113 ;
  assign n2331 = ~n2114 & ~n2330 ;
  assign n2332 = ~n2329 & ~n2331 ;
  assign n2333 = n2329 & n2331 ;
  assign n2334 = n116 & ~n287 ;
  assign n2335 = ~n392 & n2334 ;
  assign n2336 = ~n288 & n2335 ;
  assign n2337 = ~n199 & n2336 ;
  assign n2338 = ~n528 & n2337 ;
  assign n2339 = ~n210 & n2338 ;
  assign n2340 = ~n230 & ~n424 ;
  assign n2341 = ~n529 & n2340 ;
  assign n2342 = ~n169 & ~n212 ;
  assign n2343 = n2341 & n2342 ;
  assign n2344 = n885 & n2343 ;
  assign n2345 = ~n163 & n2344 ;
  assign n2346 = ~n302 & n2345 ;
  assign n2347 = ~n323 & n2346 ;
  assign n2348 = ~n304 & n2347 ;
  assign n2349 = ~n166 & n2348 ;
  assign n2350 = ~n478 & n2349 ;
  assign n2351 = n357 & n423 ;
  assign n2352 = n2350 & n2351 ;
  assign n2353 = n728 & n2352 ;
  assign n2354 = n2339 & n2353 ;
  assign n2355 = ~n171 & n2354 ;
  assign n2356 = ~n196 & n2355 ;
  assign n2357 = ~n369 & n2356 ;
  assign n2358 = ~n142 & n2357 ;
  assign n2359 = ~n322 & n2358 ;
  assign n2360 = ~n447 & n2359 ;
  assign n2361 = n1523 & n2109 ;
  assign n2362 = ~n2110 & ~n2361 ;
  assign n2363 = ~n2360 & ~n2362 ;
  assign n2364 = n539 & n2229 ;
  assign n2365 = n881 & n2364 ;
  assign n2366 = n386 & n2365 ;
  assign n2367 = ~n335 & n2366 ;
  assign n2368 = ~n89 & n2367 ;
  assign n2369 = ~n301 & n2368 ;
  assign n2370 = ~n198 & n2369 ;
  assign n2371 = n391 & n448 ;
  assign n2372 = ~n273 & n2371 ;
  assign n2373 = ~n93 & n2372 ;
  assign n2374 = ~n199 & n2373 ;
  assign n2375 = ~n342 & n2374 ;
  assign n2376 = n565 & n2375 ;
  assign n2377 = n2370 & n2376 ;
  assign n2378 = n727 & n2377 ;
  assign n2379 = n961 & n2378 ;
  assign n2380 = n124 & n2379 ;
  assign n2381 = ~n203 & n2380 ;
  assign n2382 = ~n194 & n2381 ;
  assign n2383 = ~n201 & n2382 ;
  assign n2384 = ~n311 & n2383 ;
  assign n2385 = ~n209 & n2384 ;
  assign n2386 = ~n233 & n2385 ;
  assign n2387 = ~n529 & n2386 ;
  assign n2388 = ~n317 & n2387 ;
  assign n2389 = ~n271 & n2388 ;
  assign n2390 = n2105 & ~n2107 ;
  assign n2391 = ~n2108 & ~n2390 ;
  assign n2392 = ~n2389 & ~n2391 ;
  assign n2393 = ~n528 & ~n574 ;
  assign n2394 = ~n310 & n2393 ;
  assign n2395 = ~n86 & n2394 ;
  assign n2396 = ~n452 & n2395 ;
  assign n2397 = ~n271 & ~n424 ;
  assign n2398 = n945 & n2397 ;
  assign n2399 = n2396 & n2398 ;
  assign n2400 = n2253 & n2399 ;
  assign n2401 = n348 & n2400 ;
  assign n2402 = n2308 & n2401 ;
  assign n2403 = n901 & n2402 ;
  assign n2404 = ~n334 & n2403 ;
  assign n2405 = ~n333 & n2404 ;
  assign n2406 = ~n447 & n2405 ;
  assign n2407 = ~n198 & n2406 ;
  assign n2408 = ~n326 & ~n479 ;
  assign n2409 = n371 & n781 ;
  assign n2410 = n2408 & n2409 ;
  assign n2411 = n2375 & n2410 ;
  assign n2412 = n300 & n2411 ;
  assign n2413 = n298 & n2412 ;
  assign n2414 = n958 & n2413 ;
  assign n2415 = n2407 & n2414 ;
  assign n2416 = n140 & n2415 ;
  assign n2417 = ~n303 & n2416 ;
  assign n2418 = ~n189 & n2417 ;
  assign n2419 = ~n232 & n2418 ;
  assign n2420 = ~n335 & n2419 ;
  assign n2421 = ~n213 & n2420 ;
  assign n2422 = n2101 & ~n2103 ;
  assign n2423 = ~n2104 & ~n2422 ;
  assign n2424 = ~n2421 & ~n2423 ;
  assign n2425 = n2421 & n2423 ;
  assign n2426 = ~n127 & n1092 ;
  assign n2427 = ~n202 & n2426 ;
  assign n2428 = ~n322 & n2427 ;
  assign n2429 = ~n529 & n2428 ;
  assign n2430 = ~n151 & ~n287 ;
  assign n2431 = ~n345 & n2430 ;
  assign n2432 = ~n336 & n2431 ;
  assign n2433 = ~n107 & n2432 ;
  assign n2434 = n2429 & n2433 ;
  assign n2435 = ~n318 & n2434 ;
  assign n2436 = ~n433 & n2435 ;
  assign n2437 = ~n334 & n2436 ;
  assign n2438 = ~n527 & n2437 ;
  assign n2439 = ~n129 & n2438 ;
  assign n2440 = n231 & n2397 ;
  assign n2441 = n449 & n2440 ;
  assign n2442 = n2314 & n2441 ;
  assign n2443 = n2439 & n2442 ;
  assign n2444 = n764 & n2443 ;
  assign n2445 = ~n312 & n2444 ;
  assign n2446 = ~n183 & n2445 ;
  assign n2447 = ~n109 & n2446 ;
  assign n2448 = ~n167 & n2447 ;
  assign n2449 = ~n98 & n2448 ;
  assign n2450 = ~n199 & n2449 ;
  assign n2451 = ~n332 & n2450 ;
  assign n2452 = ~n420 & n2451 ;
  assign n2453 = n2097 & ~n2099 ;
  assign n2454 = ~n2100 & ~n2453 ;
  assign n2455 = ~n2452 & ~n2454 ;
  assign n2456 = n2452 & n2454 ;
  assign n2457 = ~n2093 & ~n2096 ;
  assign n2458 = n2095 & ~n2096 ;
  assign n2459 = ~n2457 & ~n2458 ;
  assign n2460 = n752 & n1071 ;
  assign n2461 = n889 & n2460 ;
  assign n2462 = n348 & n2461 ;
  assign n2463 = n2370 & n2462 ;
  assign n2464 = n714 & n2463 ;
  assign n2465 = n2165 & n2464 ;
  assign n2466 = ~n392 & n2465 ;
  assign n2467 = ~n167 & n2466 ;
  assign n2468 = ~n333 & n2467 ;
  assign n2469 = ~n165 & n2468 ;
  assign n2470 = ~n574 & n2469 ;
  assign n2471 = ~n2459 & n2470 ;
  assign n2472 = ~n2455 & ~n2471 ;
  assign n2473 = ~n2456 & n2472 ;
  assign n2474 = ~n2455 & ~n2473 ;
  assign n2475 = ~n2424 & ~n2474 ;
  assign n2476 = ~n2425 & n2475 ;
  assign n2477 = ~n2424 & ~n2476 ;
  assign n2478 = n2389 & n2391 ;
  assign n2479 = ~n2392 & ~n2478 ;
  assign n2480 = ~n2477 & n2479 ;
  assign n2481 = ~n2392 & ~n2480 ;
  assign n2482 = n2360 & n2362 ;
  assign n2483 = ~n2363 & ~n2482 ;
  assign n2484 = ~n2481 & n2483 ;
  assign n2485 = ~n2363 & ~n2484 ;
  assign n2486 = ~n2332 & ~n2485 ;
  assign n2487 = ~n2333 & n2486 ;
  assign n2488 = ~n2332 & ~n2487 ;
  assign n2489 = ~n2302 & ~n2305 ;
  assign n2490 = ~n2304 & ~n2305 ;
  assign n2491 = ~n2489 & ~n2490 ;
  assign n2492 = ~n2488 & ~n2491 ;
  assign n2493 = ~n2305 & ~n2492 ;
  assign n2494 = ~n2270 & ~n2493 ;
  assign n2495 = ~n2271 & n2494 ;
  assign n2496 = ~n2270 & ~n2495 ;
  assign n2497 = n2239 & n2241 ;
  assign n2498 = ~n2242 & ~n2497 ;
  assign n2499 = ~n2496 & n2498 ;
  assign n2500 = ~n2242 & ~n2499 ;
  assign n2501 = ~n2203 & ~n2500 ;
  assign n2502 = ~n2204 & n2501 ;
  assign n2503 = ~n2203 & ~n2502 ;
  assign n2504 = n2184 & n2186 ;
  assign n2505 = ~n2187 & ~n2504 ;
  assign n2506 = ~n2503 & n2505 ;
  assign n2507 = ~n2187 & ~n2506 ;
  assign n2508 = ~n2138 & ~n2507 ;
  assign n2509 = ~n2139 & n2508 ;
  assign n2510 = ~n2138 & ~n2509 ;
  assign n2511 = ~n383 & n771 ;
  assign n2512 = ~n163 & n2511 ;
  assign n2513 = ~n202 & n2512 ;
  assign n2514 = ~n149 & n2513 ;
  assign n2515 = ~n343 & n2514 ;
  assign n2516 = n453 & n1066 ;
  assign n2517 = n2314 & n2516 ;
  assign n2518 = n1443 & n2517 ;
  assign n2519 = n2515 & n2518 ;
  assign n2520 = n628 & n2519 ;
  assign n2521 = n124 & n2520 ;
  assign n2522 = ~n274 & n2521 ;
  assign n2523 = n920 & n2522 ;
  assign n2524 = ~n527 & n2523 ;
  assign n2525 = ~n529 & n2524 ;
  assign n2526 = ~n198 & n2525 ;
  assign n2527 = n2510 & n2526 ;
  assign n2528 = ~n2510 & ~n2526 ;
  assign n2529 = ~n2527 & ~n2528 ;
  assign n2530 = n270 & ~n2529 ;
  assign n2531 = ~n254 & n261 ;
  assign n2532 = n254 & ~n261 ;
  assign n2533 = ~n2531 & ~n2532 ;
  assign n2534 = ~n257 & n269 ;
  assign n2535 = n2533 & n2534 ;
  assign n2536 = n2503 & ~n2505 ;
  assign n2537 = ~n2506 & ~n2536 ;
  assign n2538 = n2535 & n2537 ;
  assign n2539 = ~n2507 & ~n2509 ;
  assign n2540 = ~n2139 & n2510 ;
  assign n2541 = ~n2539 & ~n2540 ;
  assign n2542 = n269 & ~n2533 ;
  assign n2543 = ~n2541 & n2542 ;
  assign n2544 = ~n2538 & ~n2543 ;
  assign n2545 = ~n2530 & n2544 ;
  assign n2546 = ~n257 & ~n269 ;
  assign n2547 = n2537 & ~n2541 ;
  assign n2548 = ~n2500 & ~n2502 ;
  assign n2549 = ~n2204 & n2503 ;
  assign n2550 = ~n2548 & ~n2549 ;
  assign n2551 = n2537 & ~n2550 ;
  assign n2552 = n2496 & ~n2498 ;
  assign n2553 = ~n2499 & ~n2552 ;
  assign n2554 = ~n2550 & n2553 ;
  assign n2555 = ~n2493 & ~n2495 ;
  assign n2556 = ~n2271 & n2496 ;
  assign n2557 = ~n2555 & ~n2556 ;
  assign n2558 = n2553 & ~n2557 ;
  assign n2559 = ~n2488 & ~n2492 ;
  assign n2560 = ~n2491 & ~n2492 ;
  assign n2561 = ~n2559 & ~n2560 ;
  assign n2562 = ~n2557 & ~n2561 ;
  assign n2563 = ~n2485 & ~n2487 ;
  assign n2564 = ~n2333 & n2488 ;
  assign n2565 = ~n2563 & ~n2564 ;
  assign n2566 = ~n2561 & ~n2565 ;
  assign n2567 = n2481 & ~n2483 ;
  assign n2568 = ~n2484 & ~n2567 ;
  assign n2569 = ~n2565 & n2568 ;
  assign n2570 = n2477 & ~n2479 ;
  assign n2571 = ~n2480 & ~n2570 ;
  assign n2572 = n2568 & n2571 ;
  assign n2573 = ~n2474 & ~n2476 ;
  assign n2574 = ~n2425 & n2477 ;
  assign n2575 = ~n2573 & ~n2574 ;
  assign n2576 = n2571 & ~n2575 ;
  assign n2577 = ~n2471 & ~n2473 ;
  assign n2578 = ~n2456 & n2474 ;
  assign n2579 = ~n2577 & ~n2578 ;
  assign n2580 = ~n2575 & ~n2579 ;
  assign n2581 = n2459 & ~n2470 ;
  assign n2582 = ~n2471 & ~n2581 ;
  assign n2583 = ~n2579 & ~n2582 ;
  assign n2584 = n2575 & n2583 ;
  assign n2585 = ~n2580 & ~n2584 ;
  assign n2586 = ~n2571 & n2575 ;
  assign n2587 = ~n2585 & ~n2586 ;
  assign n2588 = ~n2576 & n2587 ;
  assign n2589 = ~n2576 & ~n2588 ;
  assign n2590 = ~n2568 & ~n2571 ;
  assign n2591 = ~n2589 & ~n2590 ;
  assign n2592 = ~n2572 & n2591 ;
  assign n2593 = ~n2572 & ~n2592 ;
  assign n2594 = n2565 & ~n2568 ;
  assign n2595 = ~n2569 & ~n2594 ;
  assign n2596 = ~n2593 & n2595 ;
  assign n2597 = ~n2569 & ~n2596 ;
  assign n2598 = n2561 & n2565 ;
  assign n2599 = ~n2566 & ~n2598 ;
  assign n2600 = ~n2597 & n2599 ;
  assign n2601 = ~n2566 & ~n2600 ;
  assign n2602 = n2557 & n2561 ;
  assign n2603 = ~n2562 & ~n2602 ;
  assign n2604 = ~n2601 & n2603 ;
  assign n2605 = ~n2562 & ~n2604 ;
  assign n2606 = ~n2553 & n2557 ;
  assign n2607 = ~n2558 & ~n2606 ;
  assign n2608 = ~n2605 & n2607 ;
  assign n2609 = ~n2558 & ~n2608 ;
  assign n2610 = n2550 & ~n2553 ;
  assign n2611 = ~n2554 & ~n2610 ;
  assign n2612 = ~n2609 & n2611 ;
  assign n2613 = ~n2554 & ~n2612 ;
  assign n2614 = ~n2537 & n2550 ;
  assign n2615 = ~n2551 & ~n2614 ;
  assign n2616 = ~n2613 & n2615 ;
  assign n2617 = ~n2551 & ~n2616 ;
  assign n2618 = ~n2537 & n2541 ;
  assign n2619 = ~n2547 & ~n2618 ;
  assign n2620 = ~n2617 & n2619 ;
  assign n2621 = ~n2547 & ~n2620 ;
  assign n2622 = ~n2529 & ~n2541 ;
  assign n2623 = n2529 & n2541 ;
  assign n2624 = ~n2622 & ~n2623 ;
  assign n2625 = ~n2621 & n2624 ;
  assign n2626 = n2621 & ~n2624 ;
  assign n2627 = ~n2625 & ~n2626 ;
  assign n2628 = n2546 & n2627 ;
  assign n2629 = n2545 & ~n2628 ;
  assign n2630 = ~n250 & ~n2629 ;
  assign n2631 = n250 & n2629 ;
  assign n2632 = ~n2630 & ~n2631 ;
  assign n2633 = n644 & ~n652 ;
  assign n2634 = ~n644 & n652 ;
  assign n2635 = ~n2633 & ~n2634 ;
  assign n2636 = ~n2582 & ~n2635 ;
  assign n2637 = ~n500 & ~n2636 ;
  assign n2638 = n504 & ~n652 ;
  assign n2639 = ~n504 & n652 ;
  assign n2640 = ~n2638 & ~n2639 ;
  assign n2641 = n2635 & ~n2640 ;
  assign n2642 = ~n2582 & n2641 ;
  assign n2643 = n507 & ~n2635 ;
  assign n2644 = ~n2579 & n2643 ;
  assign n2645 = ~n2642 & ~n2644 ;
  assign n2646 = n2579 & ~n2582 ;
  assign n2647 = ~n2579 & n2582 ;
  assign n2648 = ~n2646 & ~n2647 ;
  assign n2649 = ~n507 & ~n2635 ;
  assign n2650 = ~n2648 & n2649 ;
  assign n2651 = n2645 & ~n2650 ;
  assign n2652 = ~n500 & ~n2651 ;
  assign n2653 = ~n500 & ~n2652 ;
  assign n2654 = ~n2651 & ~n2652 ;
  assign n2655 = ~n2653 & ~n2654 ;
  assign n2656 = n2637 & ~n2655 ;
  assign n2657 = ~n2637 & n2655 ;
  assign n2658 = ~n2656 & ~n2657 ;
  assign n2659 = n807 & ~n996 ;
  assign n2660 = ~n807 & n996 ;
  assign n2661 = ~n2659 & ~n2660 ;
  assign n2662 = n644 & ~n815 ;
  assign n2663 = ~n644 & n815 ;
  assign n2664 = ~n2662 & ~n2663 ;
  assign n2665 = ~n2661 & ~n2664 ;
  assign n2666 = n807 & ~n815 ;
  assign n2667 = ~n807 & n815 ;
  assign n2668 = ~n2666 & ~n2667 ;
  assign n2669 = n2661 & ~n2664 ;
  assign n2670 = n2668 & n2669 ;
  assign n2671 = ~n2575 & n2670 ;
  assign n2672 = n2661 & ~n2668 ;
  assign n2673 = n2571 & n2672 ;
  assign n2674 = ~n2661 & n2664 ;
  assign n2675 = n2568 & n2674 ;
  assign n2676 = ~n2673 & ~n2675 ;
  assign n2677 = ~n2671 & n2676 ;
  assign n2678 = ~n2665 & n2677 ;
  assign n2679 = ~n2589 & ~n2592 ;
  assign n2680 = ~n2590 & n2593 ;
  assign n2681 = ~n2679 & ~n2680 ;
  assign n2682 = n2677 & n2681 ;
  assign n2683 = ~n2678 & ~n2682 ;
  assign n2684 = n644 & ~n2683 ;
  assign n2685 = ~n644 & n2683 ;
  assign n2686 = ~n2684 & ~n2685 ;
  assign n2687 = n2658 & n2686 ;
  assign n2688 = ~n2582 & ~n2661 ;
  assign n2689 = ~n644 & ~n2688 ;
  assign n2690 = ~n2582 & n2672 ;
  assign n2691 = ~n2579 & n2674 ;
  assign n2692 = ~n2690 & ~n2691 ;
  assign n2693 = ~n2648 & n2665 ;
  assign n2694 = n2692 & ~n2693 ;
  assign n2695 = ~n644 & ~n2694 ;
  assign n2696 = n644 & n2694 ;
  assign n2697 = ~n2695 & ~n2696 ;
  assign n2698 = n2689 & n2697 ;
  assign n2699 = ~n2575 & n2674 ;
  assign n2700 = ~n2582 & n2670 ;
  assign n2701 = ~n2579 & n2672 ;
  assign n2702 = ~n2700 & ~n2701 ;
  assign n2703 = ~n2699 & n2702 ;
  assign n2704 = ~n2665 & n2703 ;
  assign n2705 = n2575 & ~n2647 ;
  assign n2706 = ~n2575 & n2647 ;
  assign n2707 = ~n2705 & ~n2706 ;
  assign n2708 = n2703 & ~n2707 ;
  assign n2709 = ~n2704 & ~n2708 ;
  assign n2710 = n644 & ~n2709 ;
  assign n2711 = ~n644 & n2709 ;
  assign n2712 = ~n2710 & ~n2711 ;
  assign n2713 = n2698 & n2712 ;
  assign n2714 = n2636 & n2713 ;
  assign n2715 = n2713 & ~n2714 ;
  assign n2716 = n2636 & ~n2714 ;
  assign n2717 = ~n2715 & ~n2716 ;
  assign n2718 = ~n2575 & n2672 ;
  assign n2719 = n2571 & n2674 ;
  assign n2720 = ~n2579 & n2670 ;
  assign n2721 = ~n2719 & ~n2720 ;
  assign n2722 = ~n2718 & n2721 ;
  assign n2723 = ~n2585 & ~n2588 ;
  assign n2724 = ~n2586 & n2589 ;
  assign n2725 = ~n2723 & ~n2724 ;
  assign n2726 = n2665 & ~n2725 ;
  assign n2727 = n2722 & ~n2726 ;
  assign n2728 = ~n644 & ~n2727 ;
  assign n2729 = n644 & n2727 ;
  assign n2730 = ~n2728 & ~n2729 ;
  assign n2731 = ~n2717 & n2730 ;
  assign n2732 = ~n2714 & ~n2731 ;
  assign n2733 = ~n2658 & ~n2686 ;
  assign n2734 = ~n2687 & ~n2733 ;
  assign n2735 = ~n2732 & n2734 ;
  assign n2736 = ~n2687 & ~n2735 ;
  assign n2737 = ~n2565 & n2674 ;
  assign n2738 = n2571 & n2670 ;
  assign n2739 = n2568 & n2672 ;
  assign n2740 = ~n2738 & ~n2739 ;
  assign n2741 = ~n2737 & n2740 ;
  assign n2742 = n2593 & ~n2595 ;
  assign n2743 = ~n2596 & ~n2742 ;
  assign n2744 = n2665 & n2743 ;
  assign n2745 = n2741 & ~n2744 ;
  assign n2746 = ~n644 & ~n2745 ;
  assign n2747 = n644 & n2745 ;
  assign n2748 = ~n2746 & ~n2747 ;
  assign n2749 = ~n2575 & n2643 ;
  assign n2750 = ~n507 & n2635 ;
  assign n2751 = n2640 & n2750 ;
  assign n2752 = ~n2582 & n2751 ;
  assign n2753 = ~n2579 & n2641 ;
  assign n2754 = ~n2752 & ~n2753 ;
  assign n2755 = ~n2749 & n2754 ;
  assign n2756 = ~n2649 & n2755 ;
  assign n2757 = ~n2707 & n2755 ;
  assign n2758 = ~n2756 & ~n2757 ;
  assign n2759 = n500 & ~n2758 ;
  assign n2760 = ~n500 & n2758 ;
  assign n2761 = ~n2759 & ~n2760 ;
  assign n2762 = n2656 & n2761 ;
  assign n2763 = ~n2656 & ~n2761 ;
  assign n2764 = ~n2762 & ~n2763 ;
  assign n2765 = n2748 & n2764 ;
  assign n2766 = ~n2748 & ~n2764 ;
  assign n2767 = ~n2765 & ~n2766 ;
  assign n2768 = n2736 & ~n2767 ;
  assign n2769 = ~n2736 & n2767 ;
  assign n2770 = ~n2768 & ~n2769 ;
  assign n2771 = n988 & ~n996 ;
  assign n2772 = ~n988 & n996 ;
  assign n2773 = ~n2771 & ~n2772 ;
  assign n2774 = n250 & ~n1158 ;
  assign n2775 = ~n250 & n1158 ;
  assign n2776 = ~n2774 & ~n2775 ;
  assign n2777 = n2773 & ~n2776 ;
  assign n2778 = n2553 & n2777 ;
  assign n2779 = n988 & ~n1158 ;
  assign n2780 = ~n988 & n1158 ;
  assign n2781 = ~n2779 & ~n2780 ;
  assign n2782 = ~n2773 & n2776 ;
  assign n2783 = n2781 & n2782 ;
  assign n2784 = ~n2561 & n2783 ;
  assign n2785 = n2776 & ~n2781 ;
  assign n2786 = ~n2557 & n2785 ;
  assign n2787 = ~n2784 & ~n2786 ;
  assign n2788 = ~n2778 & n2787 ;
  assign n2789 = n2605 & ~n2607 ;
  assign n2790 = ~n2608 & ~n2789 ;
  assign n2791 = n2788 & ~n2790 ;
  assign n2792 = ~n2773 & ~n2776 ;
  assign n2793 = n2788 & ~n2792 ;
  assign n2794 = ~n2791 & ~n2793 ;
  assign n2795 = n996 & ~n2794 ;
  assign n2796 = ~n996 & n2794 ;
  assign n2797 = ~n2795 & ~n2796 ;
  assign n2798 = n2770 & n2797 ;
  assign n2799 = ~n2557 & n2777 ;
  assign n2800 = ~n2565 & n2783 ;
  assign n2801 = ~n2561 & n2785 ;
  assign n2802 = ~n2800 & ~n2801 ;
  assign n2803 = ~n2799 & n2802 ;
  assign n2804 = n2601 & ~n2603 ;
  assign n2805 = ~n2604 & ~n2804 ;
  assign n2806 = n2792 & n2805 ;
  assign n2807 = n2803 & ~n2806 ;
  assign n2808 = ~n996 & ~n2807 ;
  assign n2809 = ~n2807 & ~n2808 ;
  assign n2810 = ~n996 & ~n2808 ;
  assign n2811 = ~n2809 & ~n2810 ;
  assign n2812 = n2732 & ~n2734 ;
  assign n2813 = ~n2735 & ~n2812 ;
  assign n2814 = ~n2811 & n2813 ;
  assign n2815 = ~n2717 & ~n2731 ;
  assign n2816 = n2730 & ~n2731 ;
  assign n2817 = ~n2815 & ~n2816 ;
  assign n2818 = ~n2561 & n2777 ;
  assign n2819 = n2568 & n2783 ;
  assign n2820 = ~n2565 & n2785 ;
  assign n2821 = ~n2819 & ~n2820 ;
  assign n2822 = ~n2818 & n2821 ;
  assign n2823 = n2597 & ~n2599 ;
  assign n2824 = ~n2600 & ~n2823 ;
  assign n2825 = n2822 & ~n2824 ;
  assign n2826 = ~n2792 & n2822 ;
  assign n2827 = ~n2825 & ~n2826 ;
  assign n2828 = n996 & ~n2827 ;
  assign n2829 = ~n996 & n2827 ;
  assign n2830 = ~n2828 & ~n2829 ;
  assign n2831 = ~n2817 & n2830 ;
  assign n2832 = ~n2565 & n2777 ;
  assign n2833 = n2571 & n2783 ;
  assign n2834 = n2568 & n2785 ;
  assign n2835 = ~n2833 & ~n2834 ;
  assign n2836 = ~n2832 & n2835 ;
  assign n2837 = n2743 & n2792 ;
  assign n2838 = n2836 & ~n2837 ;
  assign n2839 = ~n996 & ~n2838 ;
  assign n2840 = ~n2838 & ~n2839 ;
  assign n2841 = ~n996 & ~n2839 ;
  assign n2842 = ~n2840 & ~n2841 ;
  assign n2843 = ~n2698 & ~n2712 ;
  assign n2844 = ~n2713 & ~n2843 ;
  assign n2845 = ~n2842 & n2844 ;
  assign n2846 = ~n2689 & ~n2697 ;
  assign n2847 = ~n2698 & ~n2846 ;
  assign n2848 = ~n2575 & n2783 ;
  assign n2849 = n2571 & n2785 ;
  assign n2850 = n2568 & n2777 ;
  assign n2851 = ~n2849 & ~n2850 ;
  assign n2852 = ~n2848 & n2851 ;
  assign n2853 = ~n2792 & n2852 ;
  assign n2854 = n2681 & n2852 ;
  assign n2855 = ~n2853 & ~n2854 ;
  assign n2856 = n996 & ~n2855 ;
  assign n2857 = ~n996 & n2855 ;
  assign n2858 = ~n2856 & ~n2857 ;
  assign n2859 = n2847 & n2858 ;
  assign n2860 = ~n2582 & n2785 ;
  assign n2861 = ~n2579 & n2777 ;
  assign n2862 = ~n2860 & ~n2861 ;
  assign n2863 = ~n2648 & n2792 ;
  assign n2864 = n2862 & ~n2863 ;
  assign n2865 = ~n996 & ~n2864 ;
  assign n2866 = ~n996 & ~n2865 ;
  assign n2867 = ~n2864 & ~n2865 ;
  assign n2868 = ~n2866 & ~n2867 ;
  assign n2869 = ~n2582 & ~n2776 ;
  assign n2870 = ~n996 & ~n2869 ;
  assign n2871 = ~n2868 & n2870 ;
  assign n2872 = ~n2575 & n2777 ;
  assign n2873 = ~n2582 & n2783 ;
  assign n2874 = ~n2579 & n2785 ;
  assign n2875 = ~n2873 & ~n2874 ;
  assign n2876 = ~n2872 & n2875 ;
  assign n2877 = ~n2707 & n2876 ;
  assign n2878 = ~n2792 & n2876 ;
  assign n2879 = ~n2877 & ~n2878 ;
  assign n2880 = n996 & ~n2879 ;
  assign n2881 = ~n996 & n2879 ;
  assign n2882 = ~n2880 & ~n2881 ;
  assign n2883 = n2871 & n2882 ;
  assign n2884 = n2688 & n2883 ;
  assign n2885 = n2883 & ~n2884 ;
  assign n2886 = n2688 & ~n2884 ;
  assign n2887 = ~n2885 & ~n2886 ;
  assign n2888 = ~n2575 & n2785 ;
  assign n2889 = n2571 & n2777 ;
  assign n2890 = ~n2579 & n2783 ;
  assign n2891 = ~n2889 & ~n2890 ;
  assign n2892 = ~n2888 & n2891 ;
  assign n2893 = ~n2725 & n2792 ;
  assign n2894 = n2892 & ~n2893 ;
  assign n2895 = ~n996 & ~n2894 ;
  assign n2896 = ~n996 & ~n2895 ;
  assign n2897 = ~n2894 & ~n2895 ;
  assign n2898 = ~n2896 & ~n2897 ;
  assign n2899 = ~n2887 & ~n2898 ;
  assign n2900 = ~n2884 & ~n2899 ;
  assign n2901 = ~n2847 & ~n2858 ;
  assign n2902 = ~n2859 & ~n2901 ;
  assign n2903 = ~n2900 & n2902 ;
  assign n2904 = ~n2859 & ~n2903 ;
  assign n2905 = ~n2842 & ~n2845 ;
  assign n2906 = n2844 & ~n2845 ;
  assign n2907 = ~n2905 & ~n2906 ;
  assign n2908 = ~n2904 & ~n2907 ;
  assign n2909 = ~n2845 & ~n2908 ;
  assign n2910 = ~n2817 & ~n2831 ;
  assign n2911 = n2830 & ~n2831 ;
  assign n2912 = ~n2910 & ~n2911 ;
  assign n2913 = ~n2909 & ~n2912 ;
  assign n2914 = ~n2831 & ~n2913 ;
  assign n2915 = ~n2811 & ~n2814 ;
  assign n2916 = n2813 & ~n2814 ;
  assign n2917 = ~n2915 & ~n2916 ;
  assign n2918 = ~n2914 & ~n2917 ;
  assign n2919 = ~n2814 & ~n2918 ;
  assign n2920 = n2770 & ~n2798 ;
  assign n2921 = n2797 & ~n2798 ;
  assign n2922 = ~n2920 & ~n2921 ;
  assign n2923 = ~n2919 & ~n2922 ;
  assign n2924 = ~n2798 & ~n2923 ;
  assign n2925 = ~n2561 & n2674 ;
  assign n2926 = n2568 & n2670 ;
  assign n2927 = ~n2565 & n2672 ;
  assign n2928 = ~n2926 & ~n2927 ;
  assign n2929 = ~n2925 & n2928 ;
  assign n2930 = n2665 & n2824 ;
  assign n2931 = n2929 & ~n2930 ;
  assign n2932 = ~n644 & ~n2931 ;
  assign n2933 = n644 & n2931 ;
  assign n2934 = ~n2932 & ~n2933 ;
  assign n2935 = ~n2575 & n2641 ;
  assign n2936 = n2571 & n2643 ;
  assign n2937 = ~n2579 & n2751 ;
  assign n2938 = ~n2936 & ~n2937 ;
  assign n2939 = ~n2935 & n2938 ;
  assign n2940 = n2649 & ~n2725 ;
  assign n2941 = n2939 & ~n2940 ;
  assign n2942 = ~n500 & ~n2941 ;
  assign n2943 = ~n2941 & ~n2942 ;
  assign n2944 = ~n500 & ~n2942 ;
  assign n2945 = ~n2943 & ~n2944 ;
  assign n2946 = ~n500 & ~n2582 ;
  assign n2947 = ~n2762 & ~n2946 ;
  assign n2948 = n2762 & n2946 ;
  assign n2949 = ~n2945 & ~n2948 ;
  assign n2950 = ~n2947 & n2949 ;
  assign n2951 = ~n2945 & ~n2950 ;
  assign n2952 = ~n2948 & ~n2950 ;
  assign n2953 = ~n2947 & n2952 ;
  assign n2954 = ~n2951 & ~n2953 ;
  assign n2955 = n2934 & ~n2954 ;
  assign n2956 = n2934 & ~n2955 ;
  assign n2957 = ~n2954 & ~n2955 ;
  assign n2958 = ~n2956 & ~n2957 ;
  assign n2959 = ~n2765 & ~n2769 ;
  assign n2960 = n2958 & n2959 ;
  assign n2961 = ~n2958 & ~n2959 ;
  assign n2962 = ~n2960 & ~n2961 ;
  assign n2963 = n2609 & ~n2611 ;
  assign n2964 = ~n2612 & ~n2963 ;
  assign n2965 = ~n2550 & n2777 ;
  assign n2966 = ~n2557 & n2783 ;
  assign n2967 = n2553 & n2785 ;
  assign n2968 = ~n2966 & ~n2967 ;
  assign n2969 = ~n2965 & n2968 ;
  assign n2970 = ~n2964 & n2969 ;
  assign n2971 = ~n2792 & n2969 ;
  assign n2972 = ~n2970 & ~n2971 ;
  assign n2973 = n996 & ~n2972 ;
  assign n2974 = ~n996 & n2972 ;
  assign n2975 = ~n2973 & ~n2974 ;
  assign n2976 = n2962 & n2975 ;
  assign n2977 = n2962 & ~n2976 ;
  assign n2978 = n2975 & ~n2976 ;
  assign n2979 = ~n2977 & ~n2978 ;
  assign n2980 = ~n2924 & ~n2979 ;
  assign n2981 = ~n2924 & ~n2980 ;
  assign n2982 = ~n2979 & ~n2980 ;
  assign n2983 = ~n2981 & ~n2982 ;
  assign n2984 = n2632 & ~n2983 ;
  assign n2985 = n2632 & ~n2984 ;
  assign n2986 = ~n2983 & ~n2984 ;
  assign n2987 = ~n2985 & ~n2986 ;
  assign n2988 = ~n2919 & ~n2923 ;
  assign n2989 = ~n2922 & ~n2923 ;
  assign n2990 = ~n2988 & ~n2989 ;
  assign n2991 = n270 & ~n2541 ;
  assign n2992 = n2535 & ~n2550 ;
  assign n2993 = n2537 & n2542 ;
  assign n2994 = ~n2992 & ~n2993 ;
  assign n2995 = ~n2991 & n2994 ;
  assign n2996 = n2617 & ~n2619 ;
  assign n2997 = ~n2620 & ~n2996 ;
  assign n2998 = n2546 & n2997 ;
  assign n2999 = n2995 & ~n2998 ;
  assign n3000 = ~n250 & ~n2999 ;
  assign n3001 = n250 & n2999 ;
  assign n3002 = ~n3000 & ~n3001 ;
  assign n3003 = ~n2990 & n3002 ;
  assign n3004 = n3002 & ~n3003 ;
  assign n3005 = ~n2990 & ~n3003 ;
  assign n3006 = ~n3004 & ~n3005 ;
  assign n3007 = ~n2914 & n2917 ;
  assign n3008 = n2914 & ~n2917 ;
  assign n3009 = ~n3007 & ~n3008 ;
  assign n3010 = n270 & n2537 ;
  assign n3011 = n2535 & n2553 ;
  assign n3012 = n2542 & ~n2550 ;
  assign n3013 = ~n3011 & ~n3012 ;
  assign n3014 = ~n3010 & n3013 ;
  assign n3015 = ~n2546 & n3014 ;
  assign n3016 = n2613 & ~n2615 ;
  assign n3017 = ~n2616 & ~n3016 ;
  assign n3018 = n3014 & ~n3017 ;
  assign n3019 = ~n3015 & ~n3018 ;
  assign n3020 = n250 & ~n3019 ;
  assign n3021 = ~n250 & n3019 ;
  assign n3022 = ~n3020 & ~n3021 ;
  assign n3023 = ~n3009 & n3022 ;
  assign n3024 = ~n2909 & ~n2913 ;
  assign n3025 = ~n2912 & ~n2913 ;
  assign n3026 = ~n3024 & ~n3025 ;
  assign n3027 = n270 & ~n2550 ;
  assign n3028 = n2535 & ~n2557 ;
  assign n3029 = n2542 & n2553 ;
  assign n3030 = ~n3028 & ~n3029 ;
  assign n3031 = ~n3027 & n3030 ;
  assign n3032 = ~n2546 & n3031 ;
  assign n3033 = ~n2964 & n3031 ;
  assign n3034 = ~n3032 & ~n3033 ;
  assign n3035 = n250 & ~n3034 ;
  assign n3036 = ~n250 & n3034 ;
  assign n3037 = ~n3035 & ~n3036 ;
  assign n3038 = ~n3026 & n3037 ;
  assign n3039 = ~n2904 & n2907 ;
  assign n3040 = n2904 & ~n2907 ;
  assign n3041 = ~n3039 & ~n3040 ;
  assign n3042 = n270 & n2553 ;
  assign n3043 = n2535 & ~n2561 ;
  assign n3044 = n2542 & ~n2557 ;
  assign n3045 = ~n3043 & ~n3044 ;
  assign n3046 = ~n3042 & n3045 ;
  assign n3047 = ~n2546 & n3046 ;
  assign n3048 = ~n2790 & n3046 ;
  assign n3049 = ~n3047 & ~n3048 ;
  assign n3050 = n250 & ~n3049 ;
  assign n3051 = ~n250 & n3049 ;
  assign n3052 = ~n3050 & ~n3051 ;
  assign n3053 = ~n3041 & n3052 ;
  assign n3054 = n270 & ~n2557 ;
  assign n3055 = n2535 & ~n2565 ;
  assign n3056 = n2542 & ~n2561 ;
  assign n3057 = ~n3055 & ~n3056 ;
  assign n3058 = ~n3054 & n3057 ;
  assign n3059 = n2546 & n2805 ;
  assign n3060 = n3058 & ~n3059 ;
  assign n3061 = ~n250 & ~n3060 ;
  assign n3062 = n250 & n3060 ;
  assign n3063 = ~n3061 & ~n3062 ;
  assign n3064 = n2900 & ~n2902 ;
  assign n3065 = ~n2903 & ~n3064 ;
  assign n3066 = n3063 & n3065 ;
  assign n3067 = ~n2887 & ~n2899 ;
  assign n3068 = ~n2898 & ~n2899 ;
  assign n3069 = ~n3067 & ~n3068 ;
  assign n3070 = n270 & ~n2561 ;
  assign n3071 = n2535 & n2568 ;
  assign n3072 = n2542 & ~n2565 ;
  assign n3073 = ~n3071 & ~n3072 ;
  assign n3074 = ~n3070 & n3073 ;
  assign n3075 = ~n2546 & n3074 ;
  assign n3076 = ~n2824 & n3074 ;
  assign n3077 = ~n3075 & ~n3076 ;
  assign n3078 = n250 & ~n3077 ;
  assign n3079 = ~n250 & n3077 ;
  assign n3080 = ~n3078 & ~n3079 ;
  assign n3081 = ~n3069 & n3080 ;
  assign n3082 = n270 & ~n2565 ;
  assign n3083 = n2535 & n2571 ;
  assign n3084 = n2542 & n2568 ;
  assign n3085 = ~n3083 & ~n3084 ;
  assign n3086 = ~n3082 & n3085 ;
  assign n3087 = n2546 & n2743 ;
  assign n3088 = n3086 & ~n3087 ;
  assign n3089 = ~n250 & ~n3088 ;
  assign n3090 = n250 & n3088 ;
  assign n3091 = ~n3089 & ~n3090 ;
  assign n3092 = ~n2871 & ~n2882 ;
  assign n3093 = ~n2883 & ~n3092 ;
  assign n3094 = n3091 & n3093 ;
  assign n3095 = n2868 & ~n2870 ;
  assign n3096 = ~n2871 & ~n3095 ;
  assign n3097 = n2535 & ~n2575 ;
  assign n3098 = n2542 & n2571 ;
  assign n3099 = n270 & n2568 ;
  assign n3100 = ~n3098 & ~n3099 ;
  assign n3101 = ~n3097 & n3100 ;
  assign n3102 = ~n2546 & n3101 ;
  assign n3103 = n2681 & n3101 ;
  assign n3104 = ~n3102 & ~n3103 ;
  assign n3105 = n250 & ~n3104 ;
  assign n3106 = ~n250 & n3104 ;
  assign n3107 = ~n3105 & ~n3106 ;
  assign n3108 = n3096 & n3107 ;
  assign n3109 = ~n269 & ~n2582 ;
  assign n3110 = ~n250 & ~n3109 ;
  assign n3111 = n2542 & ~n2582 ;
  assign n3112 = n270 & ~n2579 ;
  assign n3113 = ~n3111 & ~n3112 ;
  assign n3114 = n2546 & ~n2648 ;
  assign n3115 = n3113 & ~n3114 ;
  assign n3116 = ~n250 & ~n3115 ;
  assign n3117 = n250 & n3115 ;
  assign n3118 = ~n3116 & ~n3117 ;
  assign n3119 = n3110 & n3118 ;
  assign n3120 = n270 & ~n2575 ;
  assign n3121 = n2535 & ~n2582 ;
  assign n3122 = n2542 & ~n2579 ;
  assign n3123 = ~n3121 & ~n3122 ;
  assign n3124 = ~n3120 & n3123 ;
  assign n3125 = ~n2546 & n3124 ;
  assign n3126 = ~n2707 & n3124 ;
  assign n3127 = ~n3125 & ~n3126 ;
  assign n3128 = n250 & ~n3127 ;
  assign n3129 = ~n250 & n3127 ;
  assign n3130 = ~n3128 & ~n3129 ;
  assign n3131 = n3119 & n3130 ;
  assign n3132 = n2869 & n3131 ;
  assign n3133 = n3131 & ~n3132 ;
  assign n3134 = n2869 & ~n3132 ;
  assign n3135 = ~n3133 & ~n3134 ;
  assign n3136 = n2542 & ~n2575 ;
  assign n3137 = n270 & n2571 ;
  assign n3138 = n2535 & ~n2579 ;
  assign n3139 = ~n3137 & ~n3138 ;
  assign n3140 = ~n3136 & n3139 ;
  assign n3141 = n2546 & ~n2725 ;
  assign n3142 = n3140 & ~n3141 ;
  assign n3143 = ~n250 & ~n3142 ;
  assign n3144 = n250 & n3142 ;
  assign n3145 = ~n3143 & ~n3144 ;
  assign n3146 = ~n3135 & n3145 ;
  assign n3147 = ~n3132 & ~n3146 ;
  assign n3148 = ~n3096 & ~n3107 ;
  assign n3149 = ~n3108 & ~n3148 ;
  assign n3150 = ~n3147 & n3149 ;
  assign n3151 = ~n3108 & ~n3150 ;
  assign n3152 = ~n3091 & ~n3093 ;
  assign n3153 = ~n3094 & ~n3152 ;
  assign n3154 = ~n3151 & n3153 ;
  assign n3155 = ~n3094 & ~n3154 ;
  assign n3156 = ~n3069 & ~n3081 ;
  assign n3157 = n3080 & ~n3081 ;
  assign n3158 = ~n3156 & ~n3157 ;
  assign n3159 = ~n3155 & ~n3158 ;
  assign n3160 = ~n3081 & ~n3159 ;
  assign n3161 = ~n3063 & ~n3065 ;
  assign n3162 = ~n3066 & ~n3161 ;
  assign n3163 = ~n3160 & n3162 ;
  assign n3164 = ~n3066 & ~n3163 ;
  assign n3165 = ~n3041 & ~n3053 ;
  assign n3166 = n3052 & ~n3053 ;
  assign n3167 = ~n3165 & ~n3166 ;
  assign n3168 = ~n3164 & ~n3167 ;
  assign n3169 = ~n3053 & ~n3168 ;
  assign n3170 = ~n3026 & ~n3038 ;
  assign n3171 = n3037 & ~n3038 ;
  assign n3172 = ~n3170 & ~n3171 ;
  assign n3173 = ~n3169 & ~n3172 ;
  assign n3174 = ~n3038 & ~n3173 ;
  assign n3175 = n3009 & ~n3022 ;
  assign n3176 = ~n3023 & ~n3175 ;
  assign n3177 = ~n3174 & n3176 ;
  assign n3178 = ~n3023 & ~n3177 ;
  assign n3179 = ~n3006 & ~n3178 ;
  assign n3180 = ~n3003 & ~n3179 ;
  assign n3181 = n2987 & n3180 ;
  assign n3182 = ~n2987 & ~n3180 ;
  assign n3183 = ~n3181 & ~n3182 ;
  assign n3184 = x0 & ~x22 ;
  assign n3185 = x1 & ~n3184 ;
  assign n3186 = ~x1 & n3184 ;
  assign n3187 = ~n3185 & ~n3186 ;
  assign n3188 = ~n266 & n3187 ;
  assign n3189 = n266 & ~n3187 ;
  assign n3190 = ~n3188 & ~n3189 ;
  assign n3191 = x0 & ~n3190 ;
  assign n3192 = x0 & n3190 ;
  assign n3193 = ~n299 & n784 ;
  assign n3194 = n460 & n3193 ;
  assign n3195 = n406 & n3194 ;
  assign n3196 = n2219 & n3195 ;
  assign n3197 = n2308 & n3196 ;
  assign n3198 = n2393 & n3197 ;
  assign n3199 = n951 & n3198 ;
  assign n3200 = ~n479 & n3199 ;
  assign n3201 = ~n272 & n3200 ;
  assign n3202 = ~n187 & n3201 ;
  assign n3203 = ~n233 & n3202 ;
  assign n3204 = ~n212 & n3203 ;
  assign n3205 = ~n275 & n783 ;
  assign n3206 = ~n301 & n3205 ;
  assign n3207 = n175 & n3206 ;
  assign n3208 = n2141 & n3207 ;
  assign n3209 = ~n390 & n3208 ;
  assign n3210 = ~n201 & n3209 ;
  assign n3211 = ~n188 & n3210 ;
  assign n3212 = ~n345 & n3211 ;
  assign n3213 = ~n422 & n3212 ;
  assign n3214 = ~n310 & n3213 ;
  assign n3215 = ~n89 & n3214 ;
  assign n3216 = ~n333 & n3215 ;
  assign n3217 = ~n81 & n3216 ;
  assign n3218 = ~n317 & n3217 ;
  assign n3219 = n719 & n2341 ;
  assign n3220 = n131 & n3219 ;
  assign n3221 = n743 & n3220 ;
  assign n3222 = n3218 & n3221 ;
  assign n3223 = n185 & n3222 ;
  assign n3224 = ~n125 & n3223 ;
  assign n3225 = ~n151 & n3224 ;
  assign n3226 = ~n195 & n3225 ;
  assign n3227 = ~n202 & n3226 ;
  assign n3228 = ~n161 & n3227 ;
  assign n3229 = ~n421 & n3228 ;
  assign n3230 = ~n336 & n3229 ;
  assign n3231 = ~n452 & n3230 ;
  assign n3232 = n2527 & n3231 ;
  assign n3233 = n3204 & n3232 ;
  assign n3234 = ~n109 & ~n380 ;
  assign n3235 = n324 & n398 ;
  assign n3236 = n1140 & n3235 ;
  assign n3237 = n372 & n3236 ;
  assign n3238 = n412 & n3237 ;
  assign n3239 = n289 & n3238 ;
  assign n3240 = n460 & n3239 ;
  assign n3241 = n477 & n3240 ;
  assign n3242 = n428 & n3241 ;
  assign n3243 = n3234 & n3242 ;
  assign n3244 = ~n115 & n3243 ;
  assign n3245 = ~n3233 & n3244 ;
  assign n3246 = n3233 & ~n3244 ;
  assign n3247 = ~n3245 & ~n3246 ;
  assign n3248 = n3192 & n3247 ;
  assign n3249 = n263 & ~n3190 ;
  assign n3250 = ~n2527 & n3231 ;
  assign n3251 = n2527 & ~n3231 ;
  assign n3252 = ~n3250 & ~n3251 ;
  assign n3253 = n3249 & n3252 ;
  assign n3254 = ~n3204 & ~n3232 ;
  assign n3255 = ~n3233 & ~n3254 ;
  assign n3256 = ~x0 & ~n3187 ;
  assign n3257 = ~n3255 & n3256 ;
  assign n3258 = ~n3253 & ~n3257 ;
  assign n3259 = ~n3248 & n3258 ;
  assign n3260 = ~n3191 & n3259 ;
  assign n3261 = n3252 & ~n3255 ;
  assign n3262 = ~n2529 & n3252 ;
  assign n3263 = ~n2622 & ~n2625 ;
  assign n3264 = n2529 & ~n3252 ;
  assign n3265 = ~n3262 & ~n3264 ;
  assign n3266 = ~n3263 & n3265 ;
  assign n3267 = ~n3262 & ~n3266 ;
  assign n3268 = ~n3252 & n3255 ;
  assign n3269 = ~n3261 & ~n3268 ;
  assign n3270 = ~n3267 & n3269 ;
  assign n3271 = ~n3261 & ~n3270 ;
  assign n3272 = ~n3247 & n3255 ;
  assign n3273 = n3247 & ~n3255 ;
  assign n3274 = ~n3272 & ~n3273 ;
  assign n3275 = ~n3271 & n3274 ;
  assign n3276 = n3271 & ~n3274 ;
  assign n3277 = ~n3275 & ~n3276 ;
  assign n3278 = n3259 & ~n3277 ;
  assign n3279 = ~n3260 & ~n3278 ;
  assign n3280 = n266 & ~n3279 ;
  assign n3281 = ~n266 & n3279 ;
  assign n3282 = ~n3280 & ~n3281 ;
  assign n3283 = n3183 & n3282 ;
  assign n3284 = n3006 & n3178 ;
  assign n3285 = ~n3179 & ~n3284 ;
  assign n3286 = n3192 & ~n3255 ;
  assign n3287 = ~n2529 & n3249 ;
  assign n3288 = n3252 & n3256 ;
  assign n3289 = ~n3287 & ~n3288 ;
  assign n3290 = ~n3286 & n3289 ;
  assign n3291 = ~n3191 & n3290 ;
  assign n3292 = n3267 & ~n3269 ;
  assign n3293 = ~n3270 & ~n3292 ;
  assign n3294 = n3290 & ~n3293 ;
  assign n3295 = ~n3291 & ~n3294 ;
  assign n3296 = n266 & ~n3295 ;
  assign n3297 = ~n266 & n3295 ;
  assign n3298 = ~n3296 & ~n3297 ;
  assign n3299 = n3285 & n3298 ;
  assign n3300 = n3174 & ~n3176 ;
  assign n3301 = n3192 & n3252 ;
  assign n3302 = ~n2541 & n3249 ;
  assign n3303 = ~n2529 & n3256 ;
  assign n3304 = ~n3302 & ~n3303 ;
  assign n3305 = ~n3301 & n3304 ;
  assign n3306 = n3263 & ~n3265 ;
  assign n3307 = ~n3266 & ~n3306 ;
  assign n3308 = n3191 & n3307 ;
  assign n3309 = n3305 & ~n3308 ;
  assign n3310 = ~n266 & ~n3309 ;
  assign n3311 = ~n3309 & ~n3310 ;
  assign n3312 = ~n266 & ~n3310 ;
  assign n3313 = ~n3311 & ~n3312 ;
  assign n3314 = n2537 & n3192 ;
  assign n3315 = n2553 & n3249 ;
  assign n3316 = ~n2550 & n3256 ;
  assign n3317 = ~n3315 & ~n3316 ;
  assign n3318 = ~n3314 & n3317 ;
  assign n3319 = ~n266 & ~n3318 ;
  assign n3320 = n3017 & n3191 ;
  assign n3321 = n3318 & ~n3320 ;
  assign n3322 = n266 & n3321 ;
  assign n3323 = ~n266 & n3191 ;
  assign n3324 = n3017 & n3323 ;
  assign n3325 = ~n2550 & n3192 ;
  assign n3326 = ~n2557 & n3249 ;
  assign n3327 = n2553 & n3256 ;
  assign n3328 = ~n3326 & ~n3327 ;
  assign n3329 = ~n3325 & n3328 ;
  assign n3330 = ~n266 & ~n3329 ;
  assign n3331 = n2964 & n3191 ;
  assign n3332 = n3329 & ~n3331 ;
  assign n3333 = n266 & n3332 ;
  assign n3334 = n2964 & n3323 ;
  assign n3335 = n2553 & n3192 ;
  assign n3336 = ~n2561 & n3249 ;
  assign n3337 = ~n2557 & n3256 ;
  assign n3338 = ~n3336 & ~n3337 ;
  assign n3339 = ~n3335 & n3338 ;
  assign n3340 = ~n266 & ~n3339 ;
  assign n3341 = n2790 & n3191 ;
  assign n3342 = n3339 & ~n3341 ;
  assign n3343 = n266 & n3342 ;
  assign n3344 = n2790 & n3323 ;
  assign n3345 = n3147 & ~n3149 ;
  assign n3346 = ~n2561 & n3192 ;
  assign n3347 = n2568 & n3249 ;
  assign n3348 = ~n2565 & n3256 ;
  assign n3349 = ~n3347 & ~n3348 ;
  assign n3350 = ~n3346 & n3349 ;
  assign n3351 = ~n266 & ~n3350 ;
  assign n3352 = n2824 & n3191 ;
  assign n3353 = n3350 & ~n3352 ;
  assign n3354 = n266 & n3353 ;
  assign n3355 = n2824 & n3323 ;
  assign n3356 = ~n3119 & ~n3130 ;
  assign n3357 = ~n2575 & n3249 ;
  assign n3358 = n2571 & n3256 ;
  assign n3359 = n2568 & n3192 ;
  assign n3360 = ~n3358 & ~n3359 ;
  assign n3361 = ~n3357 & n3360 ;
  assign n3362 = ~n266 & ~n3361 ;
  assign n3363 = ~n2681 & n3191 ;
  assign n3364 = n3361 & ~n3363 ;
  assign n3365 = n266 & n3364 ;
  assign n3366 = ~n2681 & n3323 ;
  assign n3367 = x0 & ~n2582 ;
  assign n3368 = n2707 & n3323 ;
  assign n3369 = ~n2575 & n3192 ;
  assign n3370 = ~n2582 & n3249 ;
  assign n3371 = ~n2579 & n3256 ;
  assign n3372 = ~n3370 & ~n3371 ;
  assign n3373 = ~n3369 & n3372 ;
  assign n3374 = ~n266 & ~n3373 ;
  assign n3375 = ~n2648 & n3323 ;
  assign n3376 = ~n2579 & n3192 ;
  assign n3377 = ~n2582 & n3256 ;
  assign n3378 = ~n266 & ~n3377 ;
  assign n3379 = ~n3376 & n3378 ;
  assign n3380 = ~n3375 & n3379 ;
  assign n3381 = ~n3374 & n3380 ;
  assign n3382 = ~n3368 & n3381 ;
  assign n3383 = ~n3367 & n3382 ;
  assign n3384 = ~n3109 & ~n3383 ;
  assign n3385 = ~n2575 & n3256 ;
  assign n3386 = n2571 & n3192 ;
  assign n3387 = ~n2579 & n3249 ;
  assign n3388 = ~n3386 & ~n3387 ;
  assign n3389 = ~n3385 & n3388 ;
  assign n3390 = ~n2725 & n3191 ;
  assign n3391 = n3389 & ~n3390 ;
  assign n3392 = ~n266 & ~n3391 ;
  assign n3393 = n266 & n3391 ;
  assign n3394 = ~n3392 & ~n3393 ;
  assign n3395 = ~n3384 & n3394 ;
  assign n3396 = n3109 & n3383 ;
  assign n3397 = ~n3395 & ~n3396 ;
  assign n3398 = ~n3110 & ~n3118 ;
  assign n3399 = ~n3119 & ~n3398 ;
  assign n3400 = n3397 & ~n3399 ;
  assign n3401 = ~n3366 & ~n3400 ;
  assign n3402 = ~n3365 & n3401 ;
  assign n3403 = ~n3362 & n3402 ;
  assign n3404 = ~n3397 & n3399 ;
  assign n3405 = ~n3403 & ~n3404 ;
  assign n3406 = ~n2565 & n3192 ;
  assign n3407 = n2571 & n3249 ;
  assign n3408 = n2568 & n3256 ;
  assign n3409 = ~n3407 & ~n3408 ;
  assign n3410 = ~n3406 & n3409 ;
  assign n3411 = n2743 & n3191 ;
  assign n3412 = n3410 & ~n3411 ;
  assign n3413 = ~n266 & ~n3412 ;
  assign n3414 = ~n3412 & ~n3413 ;
  assign n3415 = ~n266 & ~n3413 ;
  assign n3416 = ~n3414 & ~n3415 ;
  assign n3417 = n3405 & n3416 ;
  assign n3418 = ~n3131 & ~n3417 ;
  assign n3419 = ~n3356 & n3418 ;
  assign n3420 = ~n3405 & ~n3416 ;
  assign n3421 = ~n3419 & ~n3420 ;
  assign n3422 = ~n3135 & ~n3146 ;
  assign n3423 = n3145 & ~n3146 ;
  assign n3424 = ~n3422 & ~n3423 ;
  assign n3425 = n3421 & n3424 ;
  assign n3426 = ~n3355 & ~n3425 ;
  assign n3427 = ~n3354 & n3426 ;
  assign n3428 = ~n3351 & n3427 ;
  assign n3429 = ~n3421 & ~n3424 ;
  assign n3430 = ~n3428 & ~n3429 ;
  assign n3431 = ~n2557 & n3192 ;
  assign n3432 = ~n2565 & n3249 ;
  assign n3433 = ~n2561 & n3256 ;
  assign n3434 = ~n3432 & ~n3433 ;
  assign n3435 = ~n3431 & n3434 ;
  assign n3436 = n2805 & n3191 ;
  assign n3437 = n3435 & ~n3436 ;
  assign n3438 = ~n266 & ~n3437 ;
  assign n3439 = ~n3437 & ~n3438 ;
  assign n3440 = ~n266 & ~n3438 ;
  assign n3441 = ~n3439 & ~n3440 ;
  assign n3442 = n3430 & n3441 ;
  assign n3443 = ~n3150 & ~n3442 ;
  assign n3444 = ~n3345 & n3443 ;
  assign n3445 = ~n3430 & ~n3441 ;
  assign n3446 = ~n3444 & ~n3445 ;
  assign n3447 = n3151 & ~n3153 ;
  assign n3448 = ~n3154 & ~n3447 ;
  assign n3449 = n3446 & ~n3448 ;
  assign n3450 = ~n3344 & ~n3449 ;
  assign n3451 = ~n3343 & n3450 ;
  assign n3452 = ~n3340 & n3451 ;
  assign n3453 = ~n3446 & n3448 ;
  assign n3454 = ~n3452 & ~n3453 ;
  assign n3455 = ~n3155 & ~n3159 ;
  assign n3456 = ~n3158 & ~n3159 ;
  assign n3457 = ~n3455 & ~n3456 ;
  assign n3458 = n3454 & n3457 ;
  assign n3459 = ~n3334 & ~n3458 ;
  assign n3460 = ~n3333 & n3459 ;
  assign n3461 = ~n3330 & n3460 ;
  assign n3462 = ~n3454 & ~n3457 ;
  assign n3463 = ~n3461 & ~n3462 ;
  assign n3464 = n3160 & ~n3162 ;
  assign n3465 = ~n3163 & ~n3464 ;
  assign n3466 = n3463 & ~n3465 ;
  assign n3467 = ~n3324 & ~n3466 ;
  assign n3468 = ~n3322 & n3467 ;
  assign n3469 = ~n3319 & n3468 ;
  assign n3470 = ~n3463 & n3465 ;
  assign n3471 = ~n3469 & ~n3470 ;
  assign n3472 = n3164 & n3167 ;
  assign n3473 = ~n3168 & ~n3472 ;
  assign n3474 = ~n3471 & n3473 ;
  assign n3475 = ~n2541 & n3192 ;
  assign n3476 = ~n2550 & n3249 ;
  assign n3477 = n2537 & n3256 ;
  assign n3478 = ~n3476 & ~n3477 ;
  assign n3479 = ~n3475 & n3478 ;
  assign n3480 = n2997 & n3191 ;
  assign n3481 = n3479 & ~n3480 ;
  assign n3482 = n266 & ~n3481 ;
  assign n3483 = ~n266 & n3481 ;
  assign n3484 = ~n3482 & ~n3483 ;
  assign n3485 = ~n3474 & n3484 ;
  assign n3486 = n3471 & ~n3473 ;
  assign n3487 = ~n3485 & ~n3486 ;
  assign n3488 = n3169 & n3172 ;
  assign n3489 = ~n3173 & ~n3488 ;
  assign n3490 = ~n3487 & ~n3489 ;
  assign n3491 = ~n2529 & n3192 ;
  assign n3492 = n2537 & n3249 ;
  assign n3493 = ~n2541 & n3256 ;
  assign n3494 = ~n3492 & ~n3493 ;
  assign n3495 = ~n3491 & n3494 ;
  assign n3496 = n2627 & n3191 ;
  assign n3497 = n3495 & ~n3496 ;
  assign n3498 = ~n266 & ~n3497 ;
  assign n3499 = n266 & n3497 ;
  assign n3500 = ~n3498 & ~n3499 ;
  assign n3501 = ~n3490 & n3500 ;
  assign n3502 = n3487 & n3489 ;
  assign n3503 = ~n3501 & ~n3502 ;
  assign n3504 = n3313 & n3503 ;
  assign n3505 = ~n3177 & ~n3504 ;
  assign n3506 = ~n3300 & n3505 ;
  assign n3507 = ~n3313 & ~n3503 ;
  assign n3508 = ~n3506 & ~n3507 ;
  assign n3509 = n3285 & ~n3299 ;
  assign n3510 = n3298 & ~n3299 ;
  assign n3511 = ~n3509 & ~n3510 ;
  assign n3512 = ~n3508 & ~n3511 ;
  assign n3513 = ~n3299 & ~n3512 ;
  assign n3514 = n3183 & ~n3283 ;
  assign n3515 = n3282 & ~n3283 ;
  assign n3516 = ~n3514 & ~n3515 ;
  assign n3517 = ~n3513 & ~n3516 ;
  assign n3518 = ~n3283 & ~n3517 ;
  assign n3519 = ~n2984 & ~n3182 ;
  assign n3520 = n270 & n3252 ;
  assign n3521 = n2535 & ~n2541 ;
  assign n3522 = ~n2529 & n2542 ;
  assign n3523 = ~n3521 & ~n3522 ;
  assign n3524 = ~n3520 & n3523 ;
  assign n3525 = n2546 & n3307 ;
  assign n3526 = n3524 & ~n3525 ;
  assign n3527 = ~n250 & ~n3526 ;
  assign n3528 = n250 & n3526 ;
  assign n3529 = ~n3527 & ~n3528 ;
  assign n3530 = ~n2976 & ~n2980 ;
  assign n3531 = ~n2955 & ~n2961 ;
  assign n3532 = ~n2557 & n2674 ;
  assign n3533 = ~n2565 & n2670 ;
  assign n3534 = ~n2561 & n2672 ;
  assign n3535 = ~n3533 & ~n3534 ;
  assign n3536 = ~n3532 & n3535 ;
  assign n3537 = n2665 & n2805 ;
  assign n3538 = n3536 & ~n3537 ;
  assign n3539 = ~n644 & ~n3538 ;
  assign n3540 = n644 & n3538 ;
  assign n3541 = ~n3539 & ~n3540 ;
  assign n3542 = ~n500 & ~n2579 ;
  assign n3543 = ~n2575 & n2751 ;
  assign n3544 = n2571 & n2641 ;
  assign n3545 = n2568 & n2643 ;
  assign n3546 = ~n3544 & ~n3545 ;
  assign n3547 = ~n3543 & n3546 ;
  assign n3548 = n2649 & ~n2681 ;
  assign n3549 = n3547 & ~n3548 ;
  assign n3550 = ~n500 & ~n3549 ;
  assign n3551 = n3542 & ~n3550 ;
  assign n3552 = n3542 & ~n3551 ;
  assign n3553 = n500 & n3549 ;
  assign n3554 = ~n3550 & ~n3553 ;
  assign n3555 = ~n3551 & n3554 ;
  assign n3556 = ~n3552 & ~n3555 ;
  assign n3557 = ~n2952 & ~n3556 ;
  assign n3558 = ~n2952 & ~n3557 ;
  assign n3559 = ~n3556 & ~n3557 ;
  assign n3560 = ~n3558 & ~n3559 ;
  assign n3561 = n3541 & ~n3560 ;
  assign n3562 = n3541 & ~n3561 ;
  assign n3563 = ~n3560 & ~n3561 ;
  assign n3564 = ~n3562 & ~n3563 ;
  assign n3565 = ~n3531 & n3564 ;
  assign n3566 = n3531 & ~n3564 ;
  assign n3567 = ~n3565 & ~n3566 ;
  assign n3568 = n2537 & n2777 ;
  assign n3569 = n2553 & n2783 ;
  assign n3570 = ~n2550 & n2785 ;
  assign n3571 = ~n3569 & ~n3570 ;
  assign n3572 = ~n3568 & n3571 ;
  assign n3573 = ~n3017 & n3572 ;
  assign n3574 = ~n2792 & n3572 ;
  assign n3575 = ~n3573 & ~n3574 ;
  assign n3576 = n996 & ~n3575 ;
  assign n3577 = ~n996 & n3575 ;
  assign n3578 = ~n3576 & ~n3577 ;
  assign n3579 = ~n3567 & n3578 ;
  assign n3580 = n3567 & ~n3578 ;
  assign n3581 = ~n3579 & ~n3580 ;
  assign n3582 = ~n3530 & n3581 ;
  assign n3583 = n3530 & ~n3581 ;
  assign n3584 = ~n3582 & ~n3583 ;
  assign n3585 = n3529 & n3584 ;
  assign n3586 = ~n3529 & ~n3584 ;
  assign n3587 = ~n3585 & ~n3586 ;
  assign n3588 = ~n3519 & n3587 ;
  assign n3589 = n3519 & ~n3587 ;
  assign n3590 = ~n3588 & ~n3589 ;
  assign n3591 = ~n323 & n477 ;
  assign n3592 = ~n123 & n3591 ;
  assign n3593 = n489 & n3592 ;
  assign n3594 = n460 & n3593 ;
  assign n3595 = n389 & n3594 ;
  assign n3596 = n379 & n3595 ;
  assign n3597 = ~n163 & n3596 ;
  assign n3598 = ~n194 & n3597 ;
  assign n3599 = ~n199 & n3598 ;
  assign n3600 = n3233 & n3244 ;
  assign n3601 = ~n3599 & ~n3600 ;
  assign n3602 = n3599 & n3600 ;
  assign n3603 = ~n3601 & ~n3602 ;
  assign n3604 = n3192 & ~n3603 ;
  assign n3605 = n3249 & ~n3255 ;
  assign n3606 = n3247 & n3256 ;
  assign n3607 = ~n3605 & ~n3606 ;
  assign n3608 = ~n3604 & n3607 ;
  assign n3609 = ~n3191 & n3608 ;
  assign n3610 = ~n3273 & ~n3275 ;
  assign n3611 = ~n3247 & n3603 ;
  assign n3612 = n3247 & ~n3603 ;
  assign n3613 = ~n3611 & ~n3612 ;
  assign n3614 = ~n3610 & n3613 ;
  assign n3615 = n3610 & ~n3613 ;
  assign n3616 = ~n3614 & ~n3615 ;
  assign n3617 = n3608 & ~n3616 ;
  assign n3618 = ~n3609 & ~n3617 ;
  assign n3619 = n266 & ~n3618 ;
  assign n3620 = ~n266 & n3618 ;
  assign n3621 = ~n3619 & ~n3620 ;
  assign n3622 = n3590 & n3621 ;
  assign n3623 = ~n3590 & ~n3621 ;
  assign n3624 = ~n3622 & ~n3623 ;
  assign n3625 = ~n3518 & n3624 ;
  assign n3626 = n3518 & ~n3624 ;
  assign n3627 = ~n3625 & ~n3626 ;
  assign n3628 = ~n246 & n3627 ;
  assign n3629 = ~n89 & ~n481 ;
  assign n3630 = ~n711 & n3629 ;
  assign n3631 = ~n271 & n3630 ;
  assign n3632 = ~n129 & n3631 ;
  assign n3633 = n781 & n3632 ;
  assign n3634 = ~n114 & n3633 ;
  assign n3635 = ~n125 & n3634 ;
  assign n3636 = ~n161 & n3635 ;
  assign n3637 = ~n288 & n3636 ;
  assign n3638 = ~n108 & n3637 ;
  assign n3639 = ~n334 & n3638 ;
  assign n3640 = ~n117 & n3639 ;
  assign n3641 = ~n81 & n3640 ;
  assign n3642 = n347 & n480 ;
  assign n3643 = n1109 & n3642 ;
  assign n3644 = ~n192 & n3643 ;
  assign n3645 = ~n230 & n3644 ;
  assign n3646 = ~n470 & n3645 ;
  assign n3647 = ~n528 & n3646 ;
  assign n3648 = ~n420 & n3647 ;
  assign n3649 = ~n446 & n3648 ;
  assign n3650 = ~n190 & n3649 ;
  assign n3651 = n764 & n3650 ;
  assign n3652 = ~n392 & n3651 ;
  assign n3653 = ~n273 & n3652 ;
  assign n3654 = n2429 & n3653 ;
  assign n3655 = n3641 & n3654 ;
  assign n3656 = n955 & n3655 ;
  assign n3657 = ~n112 & n3656 ;
  assign n3658 = ~n229 & n3657 ;
  assign n3659 = ~n302 & n3658 ;
  assign n3660 = ~n421 & n3659 ;
  assign n3661 = ~n121 & n3660 ;
  assign n3662 = ~n272 & n3661 ;
  assign n3663 = ~n310 & n3662 ;
  assign n3664 = ~n445 & n3663 ;
  assign n3665 = ~n317 & n3664 ;
  assign n3666 = n3513 & ~n3515 ;
  assign n3667 = ~n3514 & n3666 ;
  assign n3668 = ~n3517 & ~n3667 ;
  assign n3669 = n372 & n2253 ;
  assign n3670 = n2278 & n3669 ;
  assign n3671 = ~n119 & n3670 ;
  assign n3672 = ~n478 & n3671 ;
  assign n3673 = ~n331 & n3672 ;
  assign n3674 = ~n452 & n3673 ;
  assign n3675 = n316 & n788 ;
  assign n3676 = ~n112 & n3675 ;
  assign n3677 = ~n130 & n3676 ;
  assign n3678 = n435 & n2397 ;
  assign n3679 = n2408 & n3678 ;
  assign n3680 = n319 & n3679 ;
  assign n3681 = n3677 & n3680 ;
  assign n3682 = n3674 & n3681 ;
  assign n3683 = n2339 & n3682 ;
  assign n3684 = ~n390 & n3683 ;
  assign n3685 = ~n125 & n3684 ;
  assign n3686 = ~n292 & n3685 ;
  assign n3687 = ~n194 & n3686 ;
  assign n3688 = ~n149 & n3687 ;
  assign n3689 = ~n193 & n3688 ;
  assign n3690 = ~n277 & n3689 ;
  assign n3691 = n3508 & n3511 ;
  assign n3692 = ~n3512 & ~n3691 ;
  assign n3693 = ~n3690 & n3692 ;
  assign n3694 = ~n3668 & ~n3693 ;
  assign n3695 = ~n3665 & ~n3694 ;
  assign n3696 = n3668 & n3693 ;
  assign n3697 = ~n3695 & ~n3696 ;
  assign n3698 = ~n246 & ~n3628 ;
  assign n3699 = n3627 & ~n3628 ;
  assign n3700 = ~n3698 & ~n3699 ;
  assign n3701 = ~n3697 & ~n3700 ;
  assign n3702 = ~n3628 & ~n3701 ;
  assign n3703 = n214 & n565 ;
  assign n3704 = ~n325 & n3703 ;
  assign n3705 = ~n98 & n3704 ;
  assign n3706 = ~n288 & n3705 ;
  assign n3707 = ~n182 & n3706 ;
  assign n3708 = ~n420 & n3707 ;
  assign n3709 = ~n444 & n3708 ;
  assign n3710 = n328 & ~n443 ;
  assign n3711 = n309 & n3710 ;
  assign n3712 = n1137 & n3711 ;
  assign n3713 = n3709 & n3712 ;
  assign n3714 = n2393 & n3713 ;
  assign n3715 = ~n197 & n3714 ;
  assign n3716 = ~n292 & n3715 ;
  assign n3717 = ~n152 & n3716 ;
  assign n3718 = ~n193 & n3717 ;
  assign n3719 = ~n529 & n3718 ;
  assign n3720 = ~n186 & n3719 ;
  assign n3721 = ~n107 & n3720 ;
  assign n3722 = ~n198 & n3721 ;
  assign n3723 = ~n3602 & n3722 ;
  assign n3724 = n3602 & ~n3722 ;
  assign n3725 = ~n3723 & ~n3724 ;
  assign n3726 = n3192 & n3725 ;
  assign n3727 = n3247 & n3249 ;
  assign n3728 = n3256 & ~n3603 ;
  assign n3729 = ~n3727 & ~n3728 ;
  assign n3730 = ~n3726 & n3729 ;
  assign n3731 = ~n3612 & ~n3614 ;
  assign n3732 = n3603 & ~n3725 ;
  assign n3733 = ~n3603 & n3725 ;
  assign n3734 = ~n3732 & ~n3733 ;
  assign n3735 = ~n3731 & n3734 ;
  assign n3736 = n3731 & ~n3734 ;
  assign n3737 = ~n3735 & ~n3736 ;
  assign n3738 = n3191 & n3737 ;
  assign n3739 = n3730 & ~n3738 ;
  assign n3740 = ~n266 & ~n3739 ;
  assign n3741 = ~n3739 & ~n3740 ;
  assign n3742 = ~n266 & ~n3740 ;
  assign n3743 = ~n3741 & ~n3742 ;
  assign n3744 = ~n3585 & ~n3588 ;
  assign n3745 = ~n2541 & n2777 ;
  assign n3746 = ~n2550 & n2783 ;
  assign n3747 = n2537 & n2785 ;
  assign n3748 = ~n3746 & ~n3747 ;
  assign n3749 = ~n3745 & n3748 ;
  assign n3750 = n2792 & n2997 ;
  assign n3751 = n3749 & ~n3750 ;
  assign n3752 = ~n996 & ~n3751 ;
  assign n3753 = ~n3751 & ~n3752 ;
  assign n3754 = ~n996 & ~n3752 ;
  assign n3755 = ~n3753 & ~n3754 ;
  assign n3756 = ~n3531 & ~n3564 ;
  assign n3757 = ~n3561 & ~n3756 ;
  assign n3758 = ~n3551 & ~n3557 ;
  assign n3759 = ~n2565 & n2643 ;
  assign n3760 = n2571 & n2751 ;
  assign n3761 = n2568 & n2641 ;
  assign n3762 = ~n3760 & ~n3761 ;
  assign n3763 = ~n3759 & n3762 ;
  assign n3764 = n2649 & n2743 ;
  assign n3765 = n3763 & ~n3764 ;
  assign n3766 = ~n500 & n2575 ;
  assign n3767 = ~n3765 & n3766 ;
  assign n3768 = n3765 & ~n3766 ;
  assign n3769 = ~n3767 & ~n3768 ;
  assign n3770 = ~n3758 & n3769 ;
  assign n3771 = n3758 & ~n3769 ;
  assign n3772 = ~n3770 & ~n3771 ;
  assign n3773 = n2553 & n2674 ;
  assign n3774 = ~n2561 & n2670 ;
  assign n3775 = ~n2557 & n2672 ;
  assign n3776 = ~n3774 & ~n3775 ;
  assign n3777 = ~n3773 & n3776 ;
  assign n3778 = ~n2665 & n3777 ;
  assign n3779 = ~n2790 & n3777 ;
  assign n3780 = ~n3778 & ~n3779 ;
  assign n3781 = n644 & ~n3780 ;
  assign n3782 = ~n644 & n3780 ;
  assign n3783 = ~n3781 & ~n3782 ;
  assign n3784 = n3772 & n3783 ;
  assign n3785 = n3772 & ~n3784 ;
  assign n3786 = n3783 & ~n3784 ;
  assign n3787 = ~n3785 & ~n3786 ;
  assign n3788 = ~n3757 & ~n3787 ;
  assign n3789 = ~n3757 & ~n3788 ;
  assign n3790 = ~n3787 & ~n3788 ;
  assign n3791 = ~n3789 & ~n3790 ;
  assign n3792 = ~n3755 & ~n3791 ;
  assign n3793 = ~n3755 & ~n3792 ;
  assign n3794 = ~n3791 & ~n3792 ;
  assign n3795 = ~n3793 & ~n3794 ;
  assign n3796 = ~n3579 & ~n3582 ;
  assign n3797 = n3795 & n3796 ;
  assign n3798 = ~n3795 & ~n3796 ;
  assign n3799 = ~n3797 & ~n3798 ;
  assign n3800 = n270 & ~n3255 ;
  assign n3801 = ~n2529 & n2535 ;
  assign n3802 = n2542 & n3252 ;
  assign n3803 = ~n3801 & ~n3802 ;
  assign n3804 = ~n3800 & n3803 ;
  assign n3805 = ~n2546 & n3804 ;
  assign n3806 = ~n3293 & n3804 ;
  assign n3807 = ~n3805 & ~n3806 ;
  assign n3808 = n250 & ~n3807 ;
  assign n3809 = ~n250 & n3807 ;
  assign n3810 = ~n3808 & ~n3809 ;
  assign n3811 = n3799 & n3810 ;
  assign n3812 = n3799 & ~n3811 ;
  assign n3813 = n3810 & ~n3811 ;
  assign n3814 = ~n3812 & ~n3813 ;
  assign n3815 = ~n3744 & ~n3814 ;
  assign n3816 = ~n3744 & ~n3815 ;
  assign n3817 = ~n3814 & ~n3815 ;
  assign n3818 = ~n3816 & ~n3817 ;
  assign n3819 = ~n3743 & ~n3818 ;
  assign n3820 = ~n3743 & ~n3819 ;
  assign n3821 = ~n3818 & ~n3819 ;
  assign n3822 = ~n3820 & ~n3821 ;
  assign n3823 = ~n3622 & ~n3625 ;
  assign n3824 = n3822 & n3823 ;
  assign n3825 = ~n3822 & ~n3823 ;
  assign n3826 = ~n3824 & ~n3825 ;
  assign n3827 = n214 & n1068 ;
  assign n3828 = n781 & n3827 ;
  assign n3829 = n1434 & n3828 ;
  assign n3830 = n2286 & n3829 ;
  assign n3831 = n618 & n3830 ;
  assign n3832 = n598 & n3831 ;
  assign n3833 = n185 & n3832 ;
  assign n3834 = ~n230 & n3833 ;
  assign n3835 = ~n123 & n3834 ;
  assign n3836 = ~n320 & n3835 ;
  assign n3837 = ~n3826 & n3836 ;
  assign n3838 = n3826 & ~n3836 ;
  assign n3839 = ~n3837 & ~n3838 ;
  assign n3840 = ~n3702 & n3839 ;
  assign n3841 = n3702 & ~n3839 ;
  assign n3842 = ~n3840 & ~n3841 ;
  assign n3843 = ~n3697 & ~n3701 ;
  assign n3844 = ~n3700 & ~n3701 ;
  assign n3845 = ~n3843 & ~n3844 ;
  assign n3846 = n3842 & ~n3845 ;
  assign n3847 = n3842 & ~n3846 ;
  assign n3848 = ~n3845 & ~n3846 ;
  assign n3849 = ~n3847 & ~n3848 ;
  assign n7676 = ~n3849 & x24 ;
  assign n3850 = ~x21 & ~x22 ;
  assign n3851 = x1 & x2 ;
  assign n3852 = x0 & n3851 ;
  assign n3853 = x3 & n3852 ;
  assign n3854 = x4 & n3853 ;
  assign n3855 = x5 & n3854 ;
  assign n3856 = x6 & n3855 ;
  assign n3857 = x7 & n3856 ;
  assign n3858 = x8 & n3857 ;
  assign n3859 = x9 & n3858 ;
  assign n3860 = x10 & n3859 ;
  assign n3861 = x11 & n3860 ;
  assign n3862 = x12 & n3861 ;
  assign n3863 = x13 & n3862 ;
  assign n3864 = x14 & n3863 ;
  assign n3865 = x15 & n3864 ;
  assign n3866 = x16 & n3865 ;
  assign n3867 = x17 & n3866 ;
  assign n3868 = x18 & n3867 ;
  assign n3869 = x19 & n3868 ;
  assign n3870 = x20 & n3869 ;
  assign n3871 = x21 & n3870 ;
  assign n3872 = ~x21 & ~n3870 ;
  assign n3873 = ~n3871 & ~n3872 ;
  assign n3874 = x22 & n3873 ;
  assign n3875 = ~n3850 & ~n3874 ;
  assign n3876 = ~x20 & ~x22 ;
  assign n3877 = ~x20 & ~n3869 ;
  assign n3878 = ~n3870 & ~n3877 ;
  assign n3879 = x22 & n3878 ;
  assign n3880 = ~n3876 & ~n3879 ;
  assign n3881 = n3875 & n3880 ;
  assign n3882 = ~x15 & ~x22 ;
  assign n3883 = x22 & ~n3865 ;
  assign n3884 = ~x15 & ~n3864 ;
  assign n3885 = n3883 & ~n3884 ;
  assign n3886 = ~n3882 & ~n3885 ;
  assign n3887 = n3881 & n3886 ;
  assign n3888 = x22 & ~n3868 ;
  assign n3889 = ~x19 & ~n3888 ;
  assign n3890 = x19 & n3888 ;
  assign n3891 = ~n3889 & ~n3890 ;
  assign n3892 = ~x18 & ~x22 ;
  assign n3893 = ~x18 & ~n3867 ;
  assign n3894 = n3888 & ~n3893 ;
  assign n3895 = ~n3892 & ~n3894 ;
  assign n3896 = ~n3891 & ~n3895 ;
  assign n3897 = x22 & ~n3866 ;
  assign n3898 = ~x17 & ~n3897 ;
  assign n3899 = x17 & n3897 ;
  assign n3900 = ~n3898 & ~n3899 ;
  assign n3901 = ~x16 & ~n3883 ;
  assign n3902 = x16 & n3883 ;
  assign n3903 = ~n3901 & ~n3902 ;
  assign n3904 = ~n3900 & n3903 ;
  assign n3905 = n3896 & n3904 ;
  assign n3906 = n3887 & n3905 ;
  assign n3907 = n3900 & n3903 ;
  assign n3908 = n3896 & n3907 ;
  assign n3909 = n3875 & ~n3880 ;
  assign n3910 = n3886 & n3909 ;
  assign n3911 = n3908 & n3910 ;
  assign n3912 = ~n3891 & n3895 ;
  assign n3913 = n3907 & n3912 ;
  assign n3914 = n3910 & n3913 ;
  assign n3915 = ~n3886 & n3909 ;
  assign n3916 = n3891 & ~n3895 ;
  assign n3917 = n3907 & n3916 ;
  assign n3918 = n3915 & n3917 ;
  assign n3919 = ~n3875 & n3880 ;
  assign n3920 = ~n3886 & n3919 ;
  assign n3921 = n3900 & ~n3903 ;
  assign n3922 = n3912 & n3921 ;
  assign n3923 = n3920 & n3922 ;
  assign n3924 = ~n3875 & ~n3880 ;
  assign n3925 = ~n3886 & n3924 ;
  assign n3926 = n3904 & n3912 ;
  assign n3927 = n3925 & n3926 ;
  assign n3928 = n3886 & n3924 ;
  assign n3929 = n3905 & n3928 ;
  assign n3930 = n3881 & ~n3886 ;
  assign n3931 = n3904 & n3916 ;
  assign n3932 = n3930 & n3931 ;
  assign n3933 = n3905 & n3920 ;
  assign n3934 = n3922 & n3925 ;
  assign n3935 = ~n3900 & ~n3903 ;
  assign n3936 = n3916 & n3935 ;
  assign n3937 = n3925 & n3936 ;
  assign n3938 = n3928 & n3936 ;
  assign n3939 = n3922 & n3928 ;
  assign n3940 = n3928 & n3931 ;
  assign n3941 = ~n3939 & ~n3940 ;
  assign n3942 = n3905 & n3910 ;
  assign n3943 = n3896 & n3921 ;
  assign n3944 = n3928 & n3943 ;
  assign n3945 = ~n3942 & ~n3944 ;
  assign n3946 = n3905 & n3915 ;
  assign n3947 = n3916 & n3921 ;
  assign n3948 = n3910 & n3947 ;
  assign n3949 = ~n3946 & ~n3948 ;
  assign n3950 = n3926 & n3928 ;
  assign n3951 = n3912 & n3935 ;
  assign n3952 = n3928 & n3951 ;
  assign n3953 = ~n3950 & ~n3952 ;
  assign n3954 = n3930 & n3936 ;
  assign n3955 = n3905 & n3925 ;
  assign n3956 = ~n3954 & ~n3955 ;
  assign n3957 = n3953 & n3956 ;
  assign n3958 = n3949 & n3957 ;
  assign n3959 = n3945 & n3958 ;
  assign n3960 = n3941 & n3959 ;
  assign n3961 = ~n3938 & n3960 ;
  assign n3962 = ~n3937 & n3961 ;
  assign n3963 = ~n3934 & n3962 ;
  assign n3964 = ~n3933 & n3963 ;
  assign n3965 = ~n3932 & n3964 ;
  assign n3966 = n3910 & n3943 ;
  assign n3967 = n3920 & n3951 ;
  assign n3968 = n3887 & n3951 ;
  assign n3969 = n3915 & n3922 ;
  assign n3970 = n3891 & n3895 ;
  assign n3971 = n3907 & n3970 ;
  assign n3972 = n3915 & n3971 ;
  assign n3973 = n3886 & n3919 ;
  assign n3974 = n3951 & n3973 ;
  assign n3975 = n3908 & n3925 ;
  assign n3976 = n3925 & n3943 ;
  assign n3977 = n3917 & n3973 ;
  assign n3978 = n3908 & n3928 ;
  assign n3979 = ~n3977 & ~n3978 ;
  assign n3980 = ~n3976 & n3979 ;
  assign n3981 = ~n3975 & n3980 ;
  assign n3982 = ~n3974 & n3981 ;
  assign n3983 = ~n3972 & n3982 ;
  assign n3984 = ~n3969 & n3983 ;
  assign n3985 = ~n3968 & n3984 ;
  assign n3986 = n3908 & n3920 ;
  assign n3987 = n3935 & n3970 ;
  assign n3988 = n3928 & n3987 ;
  assign n3989 = ~n3986 & ~n3988 ;
  assign n3990 = n3910 & n3951 ;
  assign n3991 = n3917 & n3920 ;
  assign n3992 = n3920 & n3926 ;
  assign n3993 = n3921 & n3970 ;
  assign n3994 = n3925 & n3993 ;
  assign n3995 = n3896 & n3935 ;
  assign n3996 = n3928 & n3995 ;
  assign n3997 = ~n3994 & ~n3996 ;
  assign n3998 = ~n3992 & n3997 ;
  assign n3999 = ~n3991 & n3998 ;
  assign n4000 = ~n3990 & n3999 ;
  assign n4001 = n3989 & n4000 ;
  assign n4002 = n3985 & n4001 ;
  assign n4003 = ~n3967 & n4002 ;
  assign n4004 = ~n3966 & n4003 ;
  assign n4005 = n3904 & n3970 ;
  assign n4006 = n3915 & n4005 ;
  assign n4007 = n3920 & n3931 ;
  assign n4008 = n3928 & n3947 ;
  assign n4009 = ~n4007 & ~n4008 ;
  assign n4010 = ~n4006 & n4009 ;
  assign n4011 = n3930 & n3947 ;
  assign n4012 = n3915 & n3995 ;
  assign n4013 = n3971 & n3973 ;
  assign n4014 = n3925 & n3971 ;
  assign n4015 = n3917 & n3930 ;
  assign n4016 = n3910 & n3926 ;
  assign n4017 = n3920 & n3947 ;
  assign n4018 = n3908 & n3973 ;
  assign n4019 = n3925 & n3987 ;
  assign n4020 = n3925 & n3931 ;
  assign n4021 = n3925 & n3947 ;
  assign n4022 = n3928 & n3993 ;
  assign n4023 = n3922 & n3930 ;
  assign n4024 = n3915 & n3926 ;
  assign n4025 = n3920 & n3943 ;
  assign n4026 = n3905 & n3973 ;
  assign n4027 = n3925 & n3951 ;
  assign n4028 = n3913 & n3925 ;
  assign n4029 = ~n4027 & ~n4028 ;
  assign n4030 = ~n4026 & n4029 ;
  assign n4031 = ~n4025 & n4030 ;
  assign n4032 = ~n4024 & n4031 ;
  assign n4033 = ~n4023 & n4032 ;
  assign n4034 = n3915 & n3987 ;
  assign n4035 = n3905 & n3930 ;
  assign n4036 = ~n4034 & ~n4035 ;
  assign n4037 = n3930 & n3987 ;
  assign n4038 = n3930 & n4005 ;
  assign n4039 = ~n4037 & ~n4038 ;
  assign n4040 = n4036 & n4039 ;
  assign n4041 = n4033 & n4040 ;
  assign n4042 = ~n4022 & n4041 ;
  assign n4043 = ~n4021 & n4042 ;
  assign n4044 = ~n4020 & n4043 ;
  assign n4045 = ~n4019 & n4044 ;
  assign n4046 = ~n4018 & n4045 ;
  assign n4047 = ~n4017 & n4046 ;
  assign n4048 = ~n4016 & n4047 ;
  assign n4049 = ~n4015 & n4048 ;
  assign n4050 = ~n4014 & n4049 ;
  assign n4051 = ~n4013 & n4050 ;
  assign n4052 = ~n4012 & n4051 ;
  assign n4053 = ~n4011 & n4052 ;
  assign n4054 = n3973 & n3993 ;
  assign n4055 = n3920 & n3995 ;
  assign n4056 = ~n4054 & ~n4055 ;
  assign n4057 = n3913 & n3973 ;
  assign n4058 = n3887 & n3993 ;
  assign n4059 = ~n4057 & ~n4058 ;
  assign n4060 = n4056 & n4059 ;
  assign n4061 = n4053 & n4060 ;
  assign n4062 = n4010 & n4061 ;
  assign n4063 = n4004 & n4062 ;
  assign n4064 = n3965 & n4063 ;
  assign n4065 = ~n3929 & n4064 ;
  assign n4066 = ~n3927 & n4065 ;
  assign n4067 = ~n3923 & n4066 ;
  assign n4068 = ~n3918 & n4067 ;
  assign n4069 = ~n3914 & n4068 ;
  assign n4070 = ~n3911 & n4069 ;
  assign n4071 = ~n3906 & n4070 ;
  assign n4072 = x22 & ~n3854 ;
  assign n4073 = ~x5 & ~n4072 ;
  assign n4074 = x5 & n4072 ;
  assign n4075 = ~n4073 & ~n4074 ;
  assign n4076 = ~x4 & ~x22 ;
  assign n4077 = ~x4 & ~n3853 ;
  assign n4078 = n4072 & ~n4077 ;
  assign n4079 = ~n4076 & ~n4078 ;
  assign n4080 = n4075 & ~n4079 ;
  assign n4081 = ~n4075 & n4079 ;
  assign n4082 = ~n4080 & ~n4081 ;
  assign n4083 = x22 & ~n3852 ;
  assign n4084 = ~x3 & ~n4083 ;
  assign n4085 = x3 & n4083 ;
  assign n4086 = ~n4084 & ~n4085 ;
  assign n4087 = ~x2 & ~x22 ;
  assign n4088 = x0 & x1 ;
  assign n4089 = ~x2 & ~n4088 ;
  assign n4090 = n4083 & ~n4089 ;
  assign n4091 = ~n4087 & ~n4090 ;
  assign n4092 = n4086 & ~n4091 ;
  assign n4093 = ~n4086 & n4091 ;
  assign n4094 = ~n4092 & ~n4093 ;
  assign n4095 = n4082 & ~n4094 ;
  assign n4096 = n3930 & n3951 ;
  assign n4097 = n3908 & n3915 ;
  assign n4098 = n3913 & n3915 ;
  assign n4099 = n3922 & n3973 ;
  assign n4100 = n3920 & n4005 ;
  assign n4101 = ~n4011 & ~n4100 ;
  assign n4102 = n3915 & n3931 ;
  assign n4103 = ~n3911 & ~n4102 ;
  assign n4104 = n3979 & n4103 ;
  assign n4105 = n4101 & n4104 ;
  assign n4106 = ~n3937 & n4105 ;
  assign n4107 = ~n4099 & n4106 ;
  assign n4108 = ~n3991 & n4107 ;
  assign n4109 = ~n4098 & n4108 ;
  assign n4110 = ~n4097 & n4109 ;
  assign n4111 = ~n4096 & n4110 ;
  assign n4112 = n3973 & n3995 ;
  assign n4113 = n3920 & n3936 ;
  assign n4114 = ~n4021 & ~n4113 ;
  assign n4115 = n3910 & n3987 ;
  assign n4116 = ~n3914 & ~n4115 ;
  assign n4117 = n3925 & n4005 ;
  assign n4118 = ~n3929 & ~n4117 ;
  assign n4119 = ~n4007 & n4118 ;
  assign n4120 = n4116 & n4119 ;
  assign n4121 = n4114 & n4120 ;
  assign n4122 = ~n4112 & n4121 ;
  assign n4123 = ~n4012 & n4122 ;
  assign n4124 = n3887 & n3971 ;
  assign n4125 = ~n3923 & ~n4124 ;
  assign n4126 = n3887 & n3947 ;
  assign n4127 = n3936 & n3973 ;
  assign n4128 = n3928 & n4005 ;
  assign n4129 = n3947 & n3973 ;
  assign n4130 = ~n4128 & ~n4129 ;
  assign n4131 = ~n4055 & n4130 ;
  assign n4132 = ~n4127 & n4131 ;
  assign n4133 = ~n3968 & n4132 ;
  assign n4134 = ~n4126 & n4133 ;
  assign n4135 = n3910 & n3993 ;
  assign n4136 = n3913 & n3920 ;
  assign n4137 = n3913 & n3928 ;
  assign n4138 = ~n3988 & ~n4137 ;
  assign n4139 = ~n3975 & n4138 ;
  assign n4140 = ~n4136 & n4139 ;
  assign n4141 = ~n4135 & n4140 ;
  assign n4142 = n3908 & n3930 ;
  assign n4143 = n3973 & n3987 ;
  assign n4144 = ~n4142 & ~n4143 ;
  assign n4145 = n3930 & n3971 ;
  assign n4146 = ~n3950 & ~n4145 ;
  assign n4147 = n3910 & n3995 ;
  assign n4148 = n3931 & n3973 ;
  assign n4149 = ~n4147 & ~n4148 ;
  assign n4150 = n3926 & n3973 ;
  assign n4151 = n3887 & n3913 ;
  assign n4152 = ~n3992 & ~n4026 ;
  assign n4153 = ~n4151 & n4152 ;
  assign n4154 = ~n4017 & n4153 ;
  assign n4155 = ~n4016 & n4154 ;
  assign n4156 = n3910 & n3971 ;
  assign n4157 = n3910 & n3936 ;
  assign n4158 = n3910 & n4005 ;
  assign n4159 = n3910 & n3917 ;
  assign n4160 = n3920 & n3987 ;
  assign n4161 = n3915 & n3947 ;
  assign n4162 = ~n4160 & ~n4161 ;
  assign n4163 = ~n4159 & n4162 ;
  assign n4164 = ~n4158 & n4163 ;
  assign n4165 = ~n4157 & n4164 ;
  assign n4166 = ~n4156 & n4165 ;
  assign n4167 = n3887 & n3995 ;
  assign n4168 = n3887 & n3926 ;
  assign n4169 = ~n3927 & ~n4168 ;
  assign n4170 = n3973 & n4005 ;
  assign n4171 = n4169 & ~n4170 ;
  assign n4172 = ~n4167 & n4171 ;
  assign n4173 = ~n3906 & ~n4015 ;
  assign n4174 = n4172 & n4173 ;
  assign n4175 = n4166 & n4174 ;
  assign n4176 = n4155 & n4175 ;
  assign n4177 = ~n3974 & n4176 ;
  assign n4178 = ~n3933 & n4177 ;
  assign n4179 = ~n3946 & n4178 ;
  assign n4180 = ~n4023 & n4179 ;
  assign n4181 = n3956 & n4180 ;
  assign n4182 = ~n4150 & n4181 ;
  assign n4183 = n4149 & n4182 ;
  assign n4184 = n4146 & n4183 ;
  assign n4185 = n4059 & n4184 ;
  assign n4186 = n4144 & n4185 ;
  assign n4187 = n4141 & n4186 ;
  assign n4188 = n4134 & n4187 ;
  assign n4189 = n4125 & n4188 ;
  assign n4190 = n4123 & n4189 ;
  assign n4191 = n4111 & n4190 ;
  assign n4192 = ~n4008 & n4191 ;
  assign n4193 = ~n3934 & n4192 ;
  assign n4194 = n3925 & n3995 ;
  assign n4195 = ~n3992 & ~n4150 ;
  assign n4196 = ~n3974 & ~n4137 ;
  assign n4197 = ~n4007 & ~n4127 ;
  assign n4198 = n4196 & n4197 ;
  assign n4199 = n4114 & n4198 ;
  assign n4200 = n3941 & n4199 ;
  assign n4201 = ~n4008 & n4200 ;
  assign n4202 = ~n4028 & n4201 ;
  assign n4203 = n4195 & n4202 ;
  assign n4204 = ~n3967 & n4203 ;
  assign n4205 = n3917 & n3925 ;
  assign n4206 = ~n3937 & ~n4057 ;
  assign n4207 = ~n4136 & n4206 ;
  assign n4208 = n3917 & n3928 ;
  assign n4209 = ~n3938 & ~n4208 ;
  assign n4210 = ~n4020 & n4209 ;
  assign n4211 = ~n4099 & n4210 ;
  assign n4212 = n4207 & n4211 ;
  assign n4213 = ~n4205 & n4212 ;
  assign n4214 = ~n3923 & n4213 ;
  assign n4215 = n3928 & n3971 ;
  assign n4216 = ~n4055 & ~n4215 ;
  assign n4217 = n3943 & n3973 ;
  assign n4218 = n3953 & n3989 ;
  assign n4219 = ~n3927 & n4218 ;
  assign n4220 = ~n4019 & n4219 ;
  assign n4221 = ~n4025 & n4220 ;
  assign n4222 = ~n4217 & n4221 ;
  assign n4223 = ~n4018 & n4222 ;
  assign n4224 = n4216 & n4223 ;
  assign n4225 = n4214 & n4224 ;
  assign n4226 = ~n4022 & n4225 ;
  assign n4227 = ~n3944 & n4226 ;
  assign n4228 = ~n3929 & n4227 ;
  assign n4229 = ~n3976 & n4228 ;
  assign n4230 = ~n4014 & n4229 ;
  assign n4231 = ~n3934 & n4230 ;
  assign n4232 = ~n3955 & ~n3994 ;
  assign n4233 = ~n3978 & ~n4027 ;
  assign n4234 = ~n3975 & n4233 ;
  assign n4235 = ~n4112 & n4234 ;
  assign n4236 = ~n4026 & n4235 ;
  assign n4237 = ~n3933 & n4236 ;
  assign n4238 = n4232 & n4237 ;
  assign n4239 = n4231 & n4238 ;
  assign n4240 = n4204 & n4239 ;
  assign n4241 = ~n4128 & n4240 ;
  assign n4242 = ~n3996 & n4241 ;
  assign n4243 = ~n4117 & n4242 ;
  assign n4244 = ~n4194 & n4243 ;
  assign n4245 = n3887 & n3922 ;
  assign n4246 = n3920 & n3971 ;
  assign n4247 = n3915 & n3951 ;
  assign n4248 = ~n3990 & ~n4247 ;
  assign n4249 = n3915 & n3943 ;
  assign n4250 = ~n4097 & ~n4249 ;
  assign n4251 = ~n3966 & n4250 ;
  assign n4252 = n4248 & n4251 ;
  assign n4253 = ~n3946 & n4252 ;
  assign n4254 = ~n4054 & ~n4143 ;
  assign n4255 = ~n4024 & n4254 ;
  assign n4256 = ~n4012 & n4255 ;
  assign n4257 = ~n3942 & n4256 ;
  assign n4258 = n3920 & n3993 ;
  assign n4259 = ~n4100 & ~n4258 ;
  assign n4260 = ~n4160 & ~n4170 ;
  assign n4261 = n4149 & n4260 ;
  assign n4262 = n4259 & n4261 ;
  assign n4263 = n4257 & n4262 ;
  assign n4264 = n4253 & n4263 ;
  assign n4265 = ~n4013 & n4264 ;
  assign n4266 = ~n4246 & n4265 ;
  assign n4267 = ~n3911 & n4266 ;
  assign n4268 = n3913 & n3930 ;
  assign n4269 = n3926 & n3930 ;
  assign n4270 = n3887 & n3908 ;
  assign n4271 = n3930 & n3995 ;
  assign n4272 = n3887 & n3943 ;
  assign n4273 = ~n3977 & ~n4129 ;
  assign n4274 = ~n4035 & ~n4156 ;
  assign n4275 = ~n3991 & ~n4017 ;
  assign n4276 = ~n3972 & n4275 ;
  assign n4277 = n3930 & n3943 ;
  assign n4278 = ~n4142 & ~n4277 ;
  assign n4279 = n4276 & n4278 ;
  assign n4280 = n4274 & n4279 ;
  assign n4281 = n4273 & n4280 ;
  assign n4282 = ~n3906 & n4281 ;
  assign n4283 = ~n4167 & n4282 ;
  assign n4284 = ~n4272 & n4283 ;
  assign n4285 = ~n4271 & n4284 ;
  assign n4286 = ~n4270 & n4285 ;
  assign n4287 = ~n3968 & n4286 ;
  assign n4288 = ~n4096 & n4287 ;
  assign n4289 = ~n4269 & n4288 ;
  assign n4290 = ~n4268 & n4289 ;
  assign n4291 = n4267 & n4290 ;
  assign n4292 = ~n4168 & n4291 ;
  assign n4293 = ~n4245 & n4292 ;
  assign n4294 = ~n4023 & n4293 ;
  assign n4295 = n3915 & n3993 ;
  assign n4296 = ~n3918 & ~n4135 ;
  assign n4297 = ~n4295 & n4296 ;
  assign n4298 = ~n4158 & n4297 ;
  assign n4299 = ~n4115 & n4298 ;
  assign n4300 = ~n4034 & n4299 ;
  assign n4301 = ~n4006 & n4300 ;
  assign n4302 = ~n4159 & n4301 ;
  assign n4303 = n3910 & n3922 ;
  assign n4304 = n3915 & n3936 ;
  assign n4305 = ~n4016 & ~n4304 ;
  assign n4306 = n3910 & n3931 ;
  assign n4307 = ~n4157 & ~n4161 ;
  assign n4308 = ~n4306 & n4307 ;
  assign n4309 = n4305 & n4308 ;
  assign n4310 = ~n4102 & n4309 ;
  assign n4311 = ~n4098 & n4310 ;
  assign n4312 = ~n3969 & n4311 ;
  assign n4313 = ~n3914 & n4312 ;
  assign n4314 = ~n4303 & n4313 ;
  assign n4315 = n4267 & n4314 ;
  assign n4316 = n4275 & n4315 ;
  assign n4317 = n4273 & n4316 ;
  assign n4318 = n4302 & n4317 ;
  assign n4319 = ~n3948 & n4318 ;
  assign n4320 = ~n4294 & ~n4319 ;
  assign n4321 = ~x14 & ~x22 ;
  assign n4322 = ~x14 & ~n3863 ;
  assign n4323 = ~n3864 & ~n4322 ;
  assign n4324 = x22 & n4323 ;
  assign n4325 = ~n4321 & ~n4324 ;
  assign n4326 = x22 & ~n3862 ;
  assign n4327 = ~x13 & ~n4326 ;
  assign n4328 = x13 & n4326 ;
  assign n4329 = ~n4327 & ~n4328 ;
  assign n4330 = ~n4325 & n4329 ;
  assign n4331 = n4325 & ~n4329 ;
  assign n4332 = ~n4330 & ~n4331 ;
  assign n4333 = n4320 & n4332 ;
  assign n4334 = ~n4320 & ~n4332 ;
  assign n4335 = ~n4333 & ~n4334 ;
  assign n4336 = ~n4244 & n4335 ;
  assign n4337 = n4294 & ~n4319 ;
  assign n4338 = ~n4294 & n4319 ;
  assign n4339 = ~n4337 & ~n4338 ;
  assign n4340 = n4294 & n4319 ;
  assign n4341 = n4244 & ~n4340 ;
  assign n4342 = n4339 & ~n4341 ;
  assign n4343 = ~n4325 & n4342 ;
  assign n4344 = ~n4244 & ~n4320 ;
  assign n4345 = ~n4339 & ~n4344 ;
  assign n4346 = n4325 & ~n4344 ;
  assign n4347 = ~n4345 & ~n4346 ;
  assign n4348 = ~n4343 & n4347 ;
  assign n4349 = ~n4244 & ~n4329 ;
  assign n4350 = n4348 & ~n4349 ;
  assign n4351 = ~n4348 & n4349 ;
  assign n4352 = n3887 & n3936 ;
  assign n4353 = n3887 & n4005 ;
  assign n4354 = n3887 & n3931 ;
  assign n4355 = ~n4038 & ~n4354 ;
  assign n4356 = ~n4008 & n4355 ;
  assign n4357 = ~n4021 & n4356 ;
  assign n4358 = ~n4167 & n4357 ;
  assign n4359 = ~n4025 & ~n4217 ;
  assign n4360 = ~n4096 & n4359 ;
  assign n4361 = ~n4034 & ~n4271 ;
  assign n4362 = ~n4037 & n4361 ;
  assign n4363 = ~n4027 & ~n4194 ;
  assign n4364 = ~n3927 & n4363 ;
  assign n4365 = n4362 & n4364 ;
  assign n4366 = n4360 & n4365 ;
  assign n4367 = n4358 & n4366 ;
  assign n4368 = n3985 & n4367 ;
  assign n4369 = ~n3929 & n4368 ;
  assign n4370 = ~n4148 & n4369 ;
  assign n4371 = ~n4353 & n4370 ;
  assign n4372 = ~n3967 & ~n4020 ;
  assign n4373 = ~n3991 & n4372 ;
  assign n4374 = ~n4137 & n4373 ;
  assign n4375 = ~n4160 & n4374 ;
  assign n4376 = ~n4012 & n4375 ;
  assign n4377 = ~n4270 & n4376 ;
  assign n4378 = ~n3918 & ~n3996 ;
  assign n4379 = ~n3914 & n4378 ;
  assign n4380 = ~n4303 & n4379 ;
  assign n4381 = ~n4269 & n4380 ;
  assign n4382 = ~n4018 & ~n4143 ;
  assign n4383 = ~n4129 & n4382 ;
  assign n4384 = ~n4249 & n4383 ;
  assign n4385 = ~n4098 & ~n4147 ;
  assign n4386 = ~n4156 & n4385 ;
  assign n4387 = n3965 & ~n4028 ;
  assign n4388 = ~n4159 & n4387 ;
  assign n4389 = n3887 & n3987 ;
  assign n4390 = ~n3986 & ~n4389 ;
  assign n4391 = n4388 & n4390 ;
  assign n4392 = n4386 & n4391 ;
  assign n4393 = n4384 & n4392 ;
  assign n4394 = n4381 & n4393 ;
  assign n4395 = n4377 & n4394 ;
  assign n4396 = n4371 & n4395 ;
  assign n4397 = n4155 & n4396 ;
  assign n4398 = ~n4352 & n4397 ;
  assign n4399 = n3887 & n3917 ;
  assign n4400 = n3941 & n4173 ;
  assign n4401 = ~n4020 & n4400 ;
  assign n4402 = ~n3934 & n4401 ;
  assign n4403 = ~n3972 & n4402 ;
  assign n4404 = ~n4098 & n4403 ;
  assign n4405 = ~n4306 & n4404 ;
  assign n4406 = ~n4354 & n4405 ;
  assign n4407 = ~n4022 & ~n4137 ;
  assign n4408 = ~n3914 & n4407 ;
  assign n4409 = ~n4117 & ~n4205 ;
  assign n4410 = n4274 & n4409 ;
  assign n4411 = ~n4027 & n4410 ;
  assign n4412 = ~n4148 & n4411 ;
  assign n4413 = ~n4129 & n4412 ;
  assign n4414 = ~n3954 & n4413 ;
  assign n4415 = n3953 & n4232 ;
  assign n4416 = n4305 & n4415 ;
  assign n4417 = n4414 & n4416 ;
  assign n4418 = ~n4208 & n4417 ;
  assign n4419 = ~n3988 & n4418 ;
  assign n4420 = ~n3929 & n4419 ;
  assign n4421 = ~n4017 & n4420 ;
  assign n4422 = ~n4157 & n4421 ;
  assign n4423 = ~n4126 & n4422 ;
  assign n4424 = ~n4194 & n4423 ;
  assign n4425 = ~n4151 & n4424 ;
  assign n4426 = ~n4008 & ~n4014 ;
  assign n4427 = ~n3937 & n4426 ;
  assign n4428 = ~n3969 & n4427 ;
  assign n4429 = n4425 & n4428 ;
  assign n4430 = n4144 & n4429 ;
  assign n4431 = n4408 & n4430 ;
  assign n4432 = n4406 & n4431 ;
  assign n4433 = ~n3991 & n4432 ;
  assign n4434 = ~n4246 & n4433 ;
  assign n4435 = ~n4399 & n4434 ;
  assign n4436 = ~n4011 & n4435 ;
  assign n4437 = ~n4112 & ~n4215 ;
  assign n4438 = ~n3976 & ~n4303 ;
  assign n4439 = n4437 & n4438 ;
  assign n4440 = ~n3996 & n4439 ;
  assign n4441 = ~n3975 & n4440 ;
  assign n4442 = ~n4100 & n4441 ;
  assign n4443 = ~n4102 & n4442 ;
  assign n4444 = ~n4013 & ~n4272 ;
  assign n4445 = ~n3938 & ~n4028 ;
  assign n4446 = ~n4277 & n4445 ;
  assign n4447 = ~n3927 & ~n4128 ;
  assign n4448 = ~n4170 & n4447 ;
  assign n4449 = n4056 & n4448 ;
  assign n4450 = ~n3944 & n4449 ;
  assign n4451 = ~n4021 & n4450 ;
  assign n4452 = ~n4271 & n4451 ;
  assign n4453 = ~n3932 & n4452 ;
  assign n4454 = ~n4019 & n4453 ;
  assign n4455 = ~n4258 & n4454 ;
  assign n4456 = n3979 & n4455 ;
  assign n4457 = n4446 & n4456 ;
  assign n4458 = n4444 & n4457 ;
  assign n4459 = n4443 & n4458 ;
  assign n4460 = n4436 & n4459 ;
  assign n4461 = n4162 & n4460 ;
  assign n4462 = ~n4352 & n4461 ;
  assign n4463 = ~n4167 & n4462 ;
  assign n4464 = ~n4398 & ~n4463 ;
  assign n4465 = ~n4294 & ~n4464 ;
  assign n4466 = x22 & ~n3860 ;
  assign n4467 = ~x11 & ~n4466 ;
  assign n4468 = x11 & n4466 ;
  assign n4469 = ~n4467 & ~n4468 ;
  assign n4470 = ~n4244 & ~n4469 ;
  assign n4471 = ~n4465 & n4470 ;
  assign n4472 = n4465 & ~n4470 ;
  assign n4473 = ~n4471 & ~n4472 ;
  assign n4474 = ~x12 & ~x22 ;
  assign n4475 = ~x12 & ~n3861 ;
  assign n4476 = n4326 & ~n4475 ;
  assign n4477 = ~n4474 & ~n4476 ;
  assign n4478 = ~n4244 & ~n4477 ;
  assign n4479 = n4473 & n4478 ;
  assign n4480 = ~n4471 & ~n4479 ;
  assign n4481 = ~n4350 & ~n4480 ;
  assign n4482 = ~n4351 & n4481 ;
  assign n4483 = ~n4350 & ~n4482 ;
  assign n4484 = ~n4339 & ~n4341 ;
  assign n4485 = ~n4325 & n4484 ;
  assign n4486 = n4325 & n4345 ;
  assign n4487 = n4339 & ~n4344 ;
  assign n4488 = n4329 & n4487 ;
  assign n4489 = ~n4329 & n4342 ;
  assign n4490 = ~n4488 & ~n4489 ;
  assign n4491 = ~n4486 & n4490 ;
  assign n4492 = ~n4485 & n4491 ;
  assign n4493 = n4398 & ~n4463 ;
  assign n4494 = ~n4398 & n4463 ;
  assign n4495 = ~n4493 & ~n4494 ;
  assign n4496 = n4398 & n4463 ;
  assign n4497 = n4294 & ~n4496 ;
  assign n4498 = n4495 & ~n4497 ;
  assign n4499 = ~n4325 & n4498 ;
  assign n4500 = ~n4465 & ~n4495 ;
  assign n4501 = n4325 & ~n4465 ;
  assign n4502 = ~n4500 & ~n4501 ;
  assign n4503 = ~n4499 & n4502 ;
  assign n4504 = ~n4470 & n4503 ;
  assign n4505 = ~n4329 & n4484 ;
  assign n4506 = n4329 & n4345 ;
  assign n4507 = n4477 & n4487 ;
  assign n4508 = n4342 & ~n4477 ;
  assign n4509 = ~n4507 & ~n4508 ;
  assign n4510 = ~n4506 & n4509 ;
  assign n4511 = ~n4505 & n4510 ;
  assign n4512 = n4470 & ~n4503 ;
  assign n4513 = ~n4504 & ~n4512 ;
  assign n4514 = n4511 & n4513 ;
  assign n4515 = ~n4504 & ~n4514 ;
  assign n4516 = n4492 & ~n4515 ;
  assign n4517 = ~n4492 & n4515 ;
  assign n4518 = ~n4516 & ~n4517 ;
  assign n4519 = ~n4473 & ~n4478 ;
  assign n4520 = ~n4479 & ~n4519 ;
  assign n4521 = n4518 & n4520 ;
  assign n4522 = ~n4516 & ~n4521 ;
  assign n4523 = ~n4480 & ~n4482 ;
  assign n4524 = ~n4351 & n4483 ;
  assign n4525 = ~n4523 & ~n4524 ;
  assign n4526 = ~n4522 & n4525 ;
  assign n4527 = n4522 & ~n4525 ;
  assign n4528 = ~n4526 & ~n4527 ;
  assign n4529 = ~n4022 & ~n4215 ;
  assign n4530 = ~n4019 & n4529 ;
  assign n4531 = ~n4159 & n4530 ;
  assign n4532 = ~n3966 & n4531 ;
  assign n4533 = ~n4270 & n4532 ;
  assign n4534 = ~n4168 & n4533 ;
  assign n4535 = ~n4145 & n4534 ;
  assign n4536 = n3930 & n3993 ;
  assign n4537 = ~n3923 & ~n3967 ;
  assign n4538 = ~n4016 & n4537 ;
  assign n4539 = ~n4536 & n4538 ;
  assign n4540 = ~n4137 & ~n4295 ;
  assign n4541 = ~n4303 & n4540 ;
  assign n4542 = ~n4306 & n4541 ;
  assign n4543 = ~n4151 & n4542 ;
  assign n4544 = ~n4035 & n4543 ;
  assign n4545 = n4276 & n4544 ;
  assign n4546 = n4539 & n4545 ;
  assign n4547 = ~n3939 & n4546 ;
  assign n4548 = ~n4304 & n4547 ;
  assign n4549 = ~n4097 & n4548 ;
  assign n4550 = ~n4006 & n4549 ;
  assign n4551 = ~n3906 & n4550 ;
  assign n4552 = ~n4038 & n4551 ;
  assign n4553 = ~n3932 & ~n4098 ;
  assign n4554 = ~n4148 & n4445 ;
  assign n4555 = ~n4150 & n4554 ;
  assign n4556 = ~n4018 & n4555 ;
  assign n4557 = ~n3948 & n4556 ;
  assign n4558 = ~n3977 & ~n4011 ;
  assign n4559 = ~n4015 & n4558 ;
  assign n4560 = ~n4012 & ~n4272 ;
  assign n4561 = n4559 & n4560 ;
  assign n4562 = n4557 & n4561 ;
  assign n4563 = n4553 & n4562 ;
  assign n4564 = ~n3988 & n4563 ;
  assign n4565 = ~n4057 & n4564 ;
  assign n4566 = ~n3942 & n4565 ;
  assign n4567 = ~n4352 & n4566 ;
  assign n4568 = ~n4245 & n4567 ;
  assign n4569 = ~n3937 & ~n4113 ;
  assign n4570 = ~n4247 & n4569 ;
  assign n4571 = ~n4115 & n4570 ;
  assign n4572 = ~n3968 & n4571 ;
  assign n4573 = ~n4271 & n4572 ;
  assign n4574 = ~n4014 & ~n4205 ;
  assign n4575 = ~n4102 & n4574 ;
  assign n4576 = ~n4054 & ~n4100 ;
  assign n4577 = ~n4025 & n4576 ;
  assign n4578 = n4575 & n4577 ;
  assign n4579 = n4573 & n4578 ;
  assign n4580 = n4568 & n4579 ;
  assign n4581 = n4552 & n4580 ;
  assign n4582 = n4535 & n4581 ;
  assign n4583 = ~n4208 & n4582 ;
  assign n4584 = ~n4026 & n4583 ;
  assign n4585 = ~n3933 & n4584 ;
  assign n4586 = ~n4037 & n4585 ;
  assign n4587 = ~n3966 & ~n4026 ;
  assign n4588 = ~n4037 & n4587 ;
  assign n4589 = ~n4277 & n4588 ;
  assign n4590 = ~n3969 & ~n3986 ;
  assign n4591 = ~n4147 & n4590 ;
  assign n4592 = ~n4023 & n4591 ;
  assign n4593 = ~n3911 & ~n3976 ;
  assign n4594 = ~n4270 & n4593 ;
  assign n4595 = ~n3934 & ~n3978 ;
  assign n4596 = ~n4012 & n4595 ;
  assign n4597 = n4594 & n4596 ;
  assign n4598 = n4448 & n4597 ;
  assign n4599 = n4592 & n4598 ;
  assign n4600 = ~n4019 & n4599 ;
  assign n4601 = ~n4150 & n4600 ;
  assign n4602 = ~n4217 & n4601 ;
  assign n4603 = ~n3933 & n4602 ;
  assign n4604 = ~n4115 & n4603 ;
  assign n4605 = ~n3906 & n4604 ;
  assign n4606 = ~n4025 & ~n4099 ;
  assign n4607 = ~n3923 & ~n3975 ;
  assign n4608 = ~n3944 & ~n4136 ;
  assign n4609 = ~n4258 & ~n4389 ;
  assign n4610 = n4101 & n4609 ;
  assign n4611 = n3949 & n4610 ;
  assign n4612 = ~n4058 & n4611 ;
  assign n4613 = ~n4168 & n4612 ;
  assign n4614 = ~n4097 & n4613 ;
  assign n4615 = ~n4006 & n4614 ;
  assign n4616 = n4425 & n4615 ;
  assign n4617 = n4608 & n4616 ;
  assign n4618 = n4607 & n4617 ;
  assign n4619 = n4606 & n4618 ;
  assign n4620 = n4605 & n4619 ;
  assign n4621 = n4589 & n4620 ;
  assign n4622 = ~n3972 & n4621 ;
  assign n4623 = n4378 & n4622 ;
  assign n4624 = ~n4158 & n4623 ;
  assign n4625 = ~n4536 & n4624 ;
  assign n4626 = ~n4096 & n4625 ;
  assign n4627 = ~n4586 & ~n4626 ;
  assign n4628 = ~n4398 & ~n4627 ;
  assign n4629 = x22 & ~n3858 ;
  assign n4630 = ~x9 & ~n4629 ;
  assign n4631 = x9 & n4629 ;
  assign n4632 = ~n4630 & ~n4631 ;
  assign n4633 = ~n4244 & ~n4632 ;
  assign n4634 = ~n4628 & n4633 ;
  assign n4635 = n4628 & ~n4633 ;
  assign n4636 = ~n4634 & ~n4635 ;
  assign n4637 = ~x10 & ~x22 ;
  assign n4638 = ~x10 & ~n3859 ;
  assign n4639 = n4466 & ~n4638 ;
  assign n4640 = ~n4637 & ~n4639 ;
  assign n4641 = ~n4244 & ~n4640 ;
  assign n4642 = n4636 & n4641 ;
  assign n4643 = ~n4634 & ~n4642 ;
  assign n4644 = ~n4495 & ~n4497 ;
  assign n4645 = ~n4325 & n4644 ;
  assign n4646 = n4325 & n4500 ;
  assign n4647 = ~n4465 & n4495 ;
  assign n4648 = n4329 & n4647 ;
  assign n4649 = ~n4329 & n4498 ;
  assign n4650 = ~n4648 & ~n4649 ;
  assign n4651 = ~n4646 & n4650 ;
  assign n4652 = ~n4645 & n4651 ;
  assign n4653 = ~n4477 & n4484 ;
  assign n4654 = n4345 & n4477 ;
  assign n4655 = n4469 & n4487 ;
  assign n4656 = n4342 & ~n4469 ;
  assign n4657 = ~n4655 & ~n4656 ;
  assign n4658 = ~n4654 & n4657 ;
  assign n4659 = ~n4653 & n4658 ;
  assign n4660 = n4652 & n4659 ;
  assign n4661 = n4586 & ~n4626 ;
  assign n4662 = ~n4586 & n4626 ;
  assign n4663 = ~n4661 & ~n4662 ;
  assign n4664 = n4586 & n4626 ;
  assign n4665 = n4398 & ~n4664 ;
  assign n4666 = n4663 & ~n4665 ;
  assign n4667 = ~n4325 & n4666 ;
  assign n4668 = ~n4628 & ~n4663 ;
  assign n4669 = n4325 & ~n4628 ;
  assign n4670 = ~n4668 & ~n4669 ;
  assign n4671 = ~n4667 & n4670 ;
  assign n4672 = ~n4633 & n4671 ;
  assign n4673 = ~n4329 & n4644 ;
  assign n4674 = n4329 & n4500 ;
  assign n4675 = n4477 & n4647 ;
  assign n4676 = ~n4477 & n4498 ;
  assign n4677 = ~n4675 & ~n4676 ;
  assign n4678 = ~n4674 & n4677 ;
  assign n4679 = ~n4673 & n4678 ;
  assign n4680 = n4633 & ~n4671 ;
  assign n4681 = ~n4672 & ~n4680 ;
  assign n4682 = n4679 & n4681 ;
  assign n4683 = ~n4672 & ~n4682 ;
  assign n4684 = ~n4652 & ~n4659 ;
  assign n4685 = ~n4660 & ~n4684 ;
  assign n4686 = ~n4683 & n4685 ;
  assign n4687 = ~n4660 & ~n4686 ;
  assign n4688 = ~n4643 & ~n4687 ;
  assign n4689 = ~n4643 & ~n4688 ;
  assign n4690 = ~n4687 & ~n4688 ;
  assign n4691 = ~n4689 & ~n4690 ;
  assign n4692 = ~n4511 & ~n4513 ;
  assign n4693 = ~n4514 & ~n4692 ;
  assign n4694 = ~n4691 & n4693 ;
  assign n4695 = ~n4688 & ~n4694 ;
  assign n4696 = ~n4518 & ~n4520 ;
  assign n4697 = ~n4521 & ~n4696 ;
  assign n4698 = ~n4695 & n4697 ;
  assign n4699 = ~n4469 & n4484 ;
  assign n4700 = n4345 & n4469 ;
  assign n4701 = n4487 & n4640 ;
  assign n4702 = n4342 & ~n4640 ;
  assign n4703 = ~n4701 & ~n4702 ;
  assign n4704 = ~n4700 & n4703 ;
  assign n4705 = ~n4699 & n4704 ;
  assign n4706 = ~n3966 & ~n4246 ;
  assign n4707 = n3945 & n4706 ;
  assign n4708 = ~n4352 & n4707 ;
  assign n4709 = ~n4038 & n4708 ;
  assign n4710 = ~n4096 & n4709 ;
  assign n4711 = ~n3974 & ~n4270 ;
  assign n4712 = ~n4022 & n4711 ;
  assign n4713 = ~n4150 & n4712 ;
  assign n4714 = ~n4145 & n4713 ;
  assign n4715 = n4103 & n4714 ;
  assign n4716 = n4123 & n4715 ;
  assign n4717 = n4710 & n4716 ;
  assign n4718 = ~n3952 & n4717 ;
  assign n4719 = ~n3996 & n4718 ;
  assign n4720 = ~n3986 & n4719 ;
  assign n4721 = ~n4304 & n4720 ;
  assign n4722 = ~n4295 & n4721 ;
  assign n4723 = ~n3954 & n4722 ;
  assign n4724 = ~n4170 & ~n4268 ;
  assign n4725 = ~n4147 & n4724 ;
  assign n4726 = ~n4245 & n4725 ;
  assign n4727 = ~n3927 & n4207 ;
  assign n4728 = ~n4016 & n4727 ;
  assign n4729 = ~n4389 & n4728 ;
  assign n4730 = ~n4167 & n4729 ;
  assign n4731 = ~n3939 & ~n4127 ;
  assign n4732 = n4362 & n4438 ;
  assign n4733 = n4731 & n4732 ;
  assign n4734 = n4730 & n4733 ;
  assign n4735 = n4726 & n4734 ;
  assign n4736 = ~n4019 & n4735 ;
  assign n4737 = ~n4099 & n4736 ;
  assign n4738 = ~n3948 & n4737 ;
  assign n4739 = ~n3977 & ~n4014 ;
  assign n4740 = ~n4018 & n4739 ;
  assign n4741 = ~n3992 & n4740 ;
  assign n4742 = ~n3933 & n4741 ;
  assign n4743 = ~n4536 & n4742 ;
  assign n4744 = ~n4142 & n4743 ;
  assign n4745 = ~n3990 & ~n4194 ;
  assign n4746 = ~n4035 & n4745 ;
  assign n4747 = ~n3955 & ~n4205 ;
  assign n4748 = ~n4151 & n4747 ;
  assign n4749 = n4296 & n4373 ;
  assign n4750 = n4748 & n4749 ;
  assign n4751 = n4746 & n4750 ;
  assign n4752 = n4125 & n4751 ;
  assign n4753 = n4744 & n4752 ;
  assign n4754 = n4738 & n4753 ;
  assign n4755 = n4723 & n4754 ;
  assign n4756 = ~n4100 & n4755 ;
  assign n4757 = ~n4055 & n4756 ;
  assign n4758 = ~n4058 & n4757 ;
  assign n4759 = ~n4353 & n4758 ;
  assign n4760 = ~n3969 & ~n4160 ;
  assign n4761 = ~n4247 & n4760 ;
  assign n4762 = ~n3955 & n4761 ;
  assign n4763 = ~n4150 & n4762 ;
  assign n4764 = ~n4018 & n4763 ;
  assign n4765 = ~n4034 & n4764 ;
  assign n4766 = ~n4159 & n4765 ;
  assign n4767 = ~n4157 & n4766 ;
  assign n4768 = ~n3933 & ~n4057 ;
  assign n4769 = ~n4168 & n4768 ;
  assign n4770 = ~n4269 & ~n4271 ;
  assign n4771 = n4769 & n4770 ;
  assign n4772 = ~n3944 & n4771 ;
  assign n4773 = ~n4127 & n4772 ;
  assign n4774 = ~n4246 & n4773 ;
  assign n4775 = ~n4115 & n4774 ;
  assign n4776 = ~n3990 & ~n4102 ;
  assign n4777 = ~n3974 & n4776 ;
  assign n4778 = ~n3991 & n4777 ;
  assign n4779 = ~n3968 & n4778 ;
  assign n4780 = ~n4022 & ~n4208 ;
  assign n4781 = ~n4194 & n4780 ;
  assign n4782 = ~n4028 & n4781 ;
  assign n4783 = ~n4217 & n4782 ;
  assign n4784 = ~n3929 & ~n3978 ;
  assign n4785 = ~n3996 & n4784 ;
  assign n4786 = ~n4249 & n4785 ;
  assign n4787 = n4056 & n4786 ;
  assign n4788 = n4783 & n4787 ;
  assign n4789 = n4726 & n4788 ;
  assign n4790 = ~n4128 & n4789 ;
  assign n4791 = ~n3976 & n4790 ;
  assign n4792 = ~n4020 & n4791 ;
  assign n4793 = ~n3972 & n4792 ;
  assign n4794 = n4587 & n4793 ;
  assign n4795 = ~n4023 & n4794 ;
  assign n4796 = ~n4137 & n4795 ;
  assign n4797 = ~n3975 & n4796 ;
  assign n4798 = ~n4352 & n4797 ;
  assign n4799 = ~n4151 & n4798 ;
  assign n4800 = n4779 & n4799 ;
  assign n4801 = n3941 & n4800 ;
  assign n4802 = n4775 & n4801 ;
  assign n4803 = n4767 & n4802 ;
  assign n4804 = n4414 & n4803 ;
  assign n4805 = ~n4099 & n4804 ;
  assign n4806 = ~n4303 & n4805 ;
  assign n4807 = ~n4167 & n4806 ;
  assign n4808 = ~n4759 & ~n4807 ;
  assign n4809 = ~n4586 & ~n4808 ;
  assign n4810 = x22 & ~n3856 ;
  assign n4811 = ~x7 & ~n4810 ;
  assign n4812 = x7 & n4810 ;
  assign n4813 = ~n4811 & ~n4812 ;
  assign n4814 = ~n4244 & ~n4813 ;
  assign n4815 = ~n4809 & n4814 ;
  assign n4816 = n4809 & ~n4814 ;
  assign n4817 = ~n4815 & ~n4816 ;
  assign n4818 = ~x8 & ~x22 ;
  assign n4819 = ~x8 & ~n3857 ;
  assign n4820 = n4629 & ~n4819 ;
  assign n4821 = ~n4818 & ~n4820 ;
  assign n4822 = n4817 & ~n4821 ;
  assign n4823 = ~n4244 & n4822 ;
  assign n4824 = ~n4815 & ~n4823 ;
  assign n4825 = n4705 & ~n4824 ;
  assign n4826 = n4484 & ~n4640 ;
  assign n4827 = n4345 & n4640 ;
  assign n4828 = n4487 & n4632 ;
  assign n4829 = n4342 & ~n4632 ;
  assign n4830 = ~n4828 & ~n4829 ;
  assign n4831 = ~n4827 & n4830 ;
  assign n4832 = ~n4826 & n4831 ;
  assign n4833 = ~n4663 & ~n4665 ;
  assign n4834 = ~n4325 & n4833 ;
  assign n4835 = n4325 & n4668 ;
  assign n4836 = ~n4628 & n4663 ;
  assign n4837 = n4329 & n4836 ;
  assign n4838 = ~n4329 & n4666 ;
  assign n4839 = ~n4837 & ~n4838 ;
  assign n4840 = ~n4835 & n4839 ;
  assign n4841 = ~n4834 & n4840 ;
  assign n4842 = ~n4477 & n4644 ;
  assign n4843 = n4477 & n4500 ;
  assign n4844 = n4469 & n4647 ;
  assign n4845 = ~n4469 & n4498 ;
  assign n4846 = ~n4844 & ~n4845 ;
  assign n4847 = ~n4843 & n4846 ;
  assign n4848 = ~n4842 & n4847 ;
  assign n4849 = n4841 & ~n4848 ;
  assign n4850 = ~n4841 & n4848 ;
  assign n4851 = ~n4849 & ~n4850 ;
  assign n4852 = n4832 & ~n4851 ;
  assign n4853 = n4841 & n4848 ;
  assign n4854 = ~n4852 & ~n4853 ;
  assign n4855 = n4705 & ~n4825 ;
  assign n4856 = ~n4824 & ~n4825 ;
  assign n4857 = ~n4855 & ~n4856 ;
  assign n4858 = ~n4854 & ~n4857 ;
  assign n4859 = ~n4825 & ~n4858 ;
  assign n4860 = ~n4636 & ~n4641 ;
  assign n4861 = ~n4642 & ~n4860 ;
  assign n4862 = ~n4859 & n4861 ;
  assign n4863 = n4859 & ~n4861 ;
  assign n4864 = ~n4862 & ~n4863 ;
  assign n4865 = n4683 & ~n4685 ;
  assign n4866 = ~n4686 & ~n4865 ;
  assign n4867 = n4864 & n4866 ;
  assign n4868 = ~n4862 & ~n4867 ;
  assign n4869 = ~n4691 & ~n4694 ;
  assign n4870 = n4693 & ~n4694 ;
  assign n4871 = ~n4869 & ~n4870 ;
  assign n4872 = ~n4868 & n4871 ;
  assign n4873 = n4868 & ~n4871 ;
  assign n4874 = ~n4872 & ~n4873 ;
  assign n4875 = ~n4469 & n4644 ;
  assign n4876 = n4469 & n4500 ;
  assign n4877 = n4640 & n4647 ;
  assign n4878 = n4498 & ~n4640 ;
  assign n4879 = ~n4877 & ~n4878 ;
  assign n4880 = ~n4876 & n4879 ;
  assign n4881 = ~n4875 & n4880 ;
  assign n4882 = n4484 & ~n4632 ;
  assign n4883 = n4345 & n4632 ;
  assign n4884 = n4487 & n4821 ;
  assign n4885 = n4342 & ~n4821 ;
  assign n4886 = ~n4884 & ~n4885 ;
  assign n4887 = ~n4883 & n4886 ;
  assign n4888 = ~n4882 & n4887 ;
  assign n4889 = n4881 & n4888 ;
  assign n4890 = ~n4148 & ~n4295 ;
  assign n4891 = ~n4135 & n4890 ;
  assign n4892 = ~n4026 & ~n4246 ;
  assign n4893 = ~n4353 & n4892 ;
  assign n4894 = ~n3975 & ~n4143 ;
  assign n4895 = ~n4303 & n4894 ;
  assign n4896 = ~n4272 & n4895 ;
  assign n4897 = n4893 & n4896 ;
  assign n4898 = n4891 & n4897 ;
  assign n4899 = n4783 & n4898 ;
  assign n4900 = n3949 & n4899 ;
  assign n4901 = ~n3996 & n4900 ;
  assign n4902 = ~n4127 & n4901 ;
  assign n4903 = ~n4012 & n4902 ;
  assign n4904 = ~n4269 & n4903 ;
  assign n4905 = ~n3918 & n4195 ;
  assign n4906 = ~n4035 & n4905 ;
  assign n4907 = n4248 & n4906 ;
  assign n4908 = ~n4024 & n4907 ;
  assign n4909 = n4260 & ~n4268 ;
  assign n4910 = ~n3976 & n4909 ;
  assign n4911 = ~n4014 & n4910 ;
  assign n4912 = ~n4018 & n4911 ;
  assign n4913 = ~n4304 & n4912 ;
  assign n4914 = ~n4158 & n4913 ;
  assign n4915 = ~n4145 & n4914 ;
  assign n4916 = ~n4023 & ~n4399 ;
  assign n4917 = ~n3940 & ~n4136 ;
  assign n4918 = n4916 & n4917 ;
  assign n4919 = n4409 & n4918 ;
  assign n4920 = n4358 & n4919 ;
  assign n4921 = n4125 & n4920 ;
  assign n4922 = n4915 & n4921 ;
  assign n4923 = n4908 & n4922 ;
  assign n4924 = n4111 & n4923 ;
  assign n4925 = n4904 & n4924 ;
  assign n4926 = ~n3988 & n4925 ;
  assign n4927 = ~n3933 & n4926 ;
  assign n4928 = ~n4006 & n4927 ;
  assign n4929 = ~n3966 & n4928 ;
  assign n4930 = ~n4352 & n4929 ;
  assign n4931 = n4259 & n4916 ;
  assign n4932 = n4607 & n4931 ;
  assign n4933 = ~n4020 & n4932 ;
  assign n4934 = ~n4194 & n4933 ;
  assign n4935 = n4446 & n4748 ;
  assign n4936 = n4114 & n4935 ;
  assign n4937 = n4908 & n4936 ;
  assign n4938 = n4934 & n4937 ;
  assign n4939 = ~n3929 & n4938 ;
  assign n4940 = ~n3996 & n4939 ;
  assign n4941 = ~n3950 & n4940 ;
  assign n4942 = ~n4013 & n4941 ;
  assign n4943 = ~n3969 & n4942 ;
  assign n4944 = ~n4115 & n4943 ;
  assign n4945 = ~n4126 & n4944 ;
  assign n4946 = n4437 & n4711 ;
  assign n4947 = ~n3994 & n4946 ;
  assign n4948 = ~n4014 & n4947 ;
  assign n4949 = ~n4148 & n4948 ;
  assign n4950 = ~n4099 & n4949 ;
  assign n4951 = ~n4352 & n4950 ;
  assign n4952 = ~n4536 & n4951 ;
  assign n4953 = n4360 & n4769 ;
  assign n4954 = ~n4124 & n4953 ;
  assign n4955 = n4952 & n4954 ;
  assign n4956 = n4275 & n4955 ;
  assign n4957 = ~n3967 & n4956 ;
  assign n4958 = ~n4136 & n4957 ;
  assign n4959 = ~n4058 & n4958 ;
  assign n4960 = ~n4145 & n4959 ;
  assign n4961 = ~n3954 & n4960 ;
  assign n4962 = ~n4015 & n4961 ;
  assign n4963 = ~n4008 & ~n4208 ;
  assign n4964 = ~n3942 & n4963 ;
  assign n4965 = ~n3911 & n4964 ;
  assign n4966 = n4560 & n4965 ;
  assign n4967 = n4251 & n4966 ;
  assign n4968 = n4305 & n4967 ;
  assign n4969 = n4166 & n4968 ;
  assign n4970 = n3941 & n4969 ;
  assign n4971 = n4962 & n4970 ;
  assign n4972 = n4945 & n4971 ;
  assign n4973 = ~n3952 & n4972 ;
  assign n4974 = ~n4019 & n4973 ;
  assign n4975 = ~n4135 & n4974 ;
  assign n4976 = ~n4930 & ~n4975 ;
  assign n4977 = ~n4759 & ~n4976 ;
  assign n4978 = n4930 & ~n4977 ;
  assign n4979 = ~n4930 & n4977 ;
  assign n4980 = ~x6 & ~x22 ;
  assign n4981 = ~x6 & ~n3855 ;
  assign n4982 = n4810 & ~n4981 ;
  assign n4983 = ~n4980 & ~n4982 ;
  assign n4984 = ~n4244 & ~n4983 ;
  assign n4985 = ~n4978 & n4984 ;
  assign n4986 = ~n4979 & n4985 ;
  assign n4987 = ~n4978 & ~n4986 ;
  assign n4988 = ~n4881 & ~n4888 ;
  assign n4989 = ~n4889 & ~n4988 ;
  assign n4990 = ~n4987 & n4989 ;
  assign n4991 = ~n4889 & ~n4990 ;
  assign n4992 = n4759 & ~n4807 ;
  assign n4993 = ~n4759 & n4807 ;
  assign n4994 = ~n4992 & ~n4993 ;
  assign n4995 = n4759 & n4807 ;
  assign n4996 = n4586 & ~n4995 ;
  assign n4997 = n4994 & ~n4996 ;
  assign n4998 = ~n4325 & n4997 ;
  assign n4999 = ~n4809 & ~n4994 ;
  assign n5000 = n4325 & ~n4809 ;
  assign n5001 = ~n4999 & ~n5000 ;
  assign n5002 = ~n4998 & n5001 ;
  assign n5003 = ~n4814 & n5002 ;
  assign n5004 = ~n4329 & n4833 ;
  assign n5005 = n4329 & n4668 ;
  assign n5006 = n4477 & n4836 ;
  assign n5007 = ~n4477 & n4666 ;
  assign n5008 = ~n5006 & ~n5007 ;
  assign n5009 = ~n5005 & n5008 ;
  assign n5010 = ~n5004 & n5009 ;
  assign n5011 = n4814 & ~n5002 ;
  assign n5012 = ~n5003 & ~n5011 ;
  assign n5013 = n5010 & n5012 ;
  assign n5014 = ~n5003 & ~n5013 ;
  assign n5015 = ~n4991 & ~n5014 ;
  assign n5016 = ~n4991 & ~n5015 ;
  assign n5017 = ~n5014 & ~n5015 ;
  assign n5018 = ~n5016 & ~n5017 ;
  assign n5019 = ~n4244 & ~n4823 ;
  assign n5020 = ~n4821 & n5019 ;
  assign n5021 = n4817 & ~n4823 ;
  assign n5022 = ~n5020 & ~n5021 ;
  assign n5023 = ~n5018 & ~n5022 ;
  assign n5024 = ~n5015 & ~n5023 ;
  assign n5025 = ~n4679 & ~n4681 ;
  assign n5026 = ~n4682 & ~n5025 ;
  assign n5027 = ~n5024 & n5026 ;
  assign n5028 = ~n4854 & ~n4858 ;
  assign n5029 = ~n4857 & ~n4858 ;
  assign n5030 = ~n5028 & ~n5029 ;
  assign n5031 = n5024 & ~n5026 ;
  assign n5032 = ~n5027 & ~n5031 ;
  assign n5033 = ~n5030 & n5032 ;
  assign n5034 = ~n5027 & ~n5033 ;
  assign n5035 = ~n4864 & ~n4866 ;
  assign n5036 = ~n4867 & ~n5035 ;
  assign n5037 = ~n5034 & n5036 ;
  assign n5038 = n5032 & ~n5033 ;
  assign n5039 = ~n5030 & ~n5033 ;
  assign n5040 = ~n5038 & ~n5039 ;
  assign n5041 = ~n4994 & ~n4996 ;
  assign n5042 = ~n4325 & n5041 ;
  assign n5043 = n4325 & n4999 ;
  assign n5044 = ~n4809 & n4994 ;
  assign n5045 = n4329 & n5044 ;
  assign n5046 = ~n4329 & n4997 ;
  assign n5047 = ~n5045 & ~n5046 ;
  assign n5048 = ~n5043 & n5047 ;
  assign n5049 = ~n5042 & n5048 ;
  assign n5050 = ~n4640 & n4644 ;
  assign n5051 = n4500 & n4640 ;
  assign n5052 = n4632 & n4647 ;
  assign n5053 = n4498 & ~n4632 ;
  assign n5054 = ~n5052 & ~n5053 ;
  assign n5055 = ~n5051 & n5054 ;
  assign n5056 = ~n5050 & n5055 ;
  assign n5057 = n4484 & ~n4821 ;
  assign n5058 = n4345 & n4821 ;
  assign n5059 = n4487 & n4813 ;
  assign n5060 = n4342 & ~n4813 ;
  assign n5061 = ~n5059 & ~n5060 ;
  assign n5062 = ~n5058 & n5061 ;
  assign n5063 = ~n5057 & n5062 ;
  assign n5064 = n5056 & ~n5063 ;
  assign n5065 = ~n5056 & n5063 ;
  assign n5066 = ~n5064 & ~n5065 ;
  assign n5067 = n5049 & ~n5066 ;
  assign n5068 = n5056 & n5063 ;
  assign n5069 = ~n5067 & ~n5068 ;
  assign n5070 = ~n5010 & ~n5012 ;
  assign n5071 = ~n5013 & ~n5070 ;
  assign n5072 = ~n5069 & n5071 ;
  assign n5073 = ~n5069 & ~n5072 ;
  assign n5074 = n5071 & ~n5072 ;
  assign n5075 = ~n5073 & ~n5074 ;
  assign n5076 = n4987 & ~n4989 ;
  assign n5077 = ~n4990 & ~n5076 ;
  assign n5078 = ~n5075 & n5077 ;
  assign n5079 = ~n5072 & ~n5078 ;
  assign n5080 = n4832 & ~n4852 ;
  assign n5081 = ~n4851 & ~n4852 ;
  assign n5082 = ~n5080 & ~n5081 ;
  assign n5083 = ~n5079 & ~n5082 ;
  assign n5084 = ~n5079 & ~n5083 ;
  assign n5085 = ~n5082 & ~n5083 ;
  assign n5086 = ~n5084 & ~n5085 ;
  assign n5087 = ~n5018 & ~n5023 ;
  assign n5088 = ~n5022 & ~n5023 ;
  assign n5089 = ~n5087 & ~n5088 ;
  assign n5090 = ~n5086 & ~n5089 ;
  assign n5091 = ~n5083 & ~n5090 ;
  assign n5092 = ~n5040 & ~n5091 ;
  assign n5093 = ~n5040 & ~n5092 ;
  assign n5094 = ~n5091 & ~n5092 ;
  assign n5095 = ~n5093 & ~n5094 ;
  assign n5096 = ~n4477 & n4833 ;
  assign n5097 = n4477 & n4668 ;
  assign n5098 = n4469 & n4836 ;
  assign n5099 = ~n4469 & n4666 ;
  assign n5100 = ~n5098 & ~n5099 ;
  assign n5101 = ~n5097 & n5100 ;
  assign n5102 = ~n5096 & n5101 ;
  assign n5103 = ~n4979 & n4987 ;
  assign n5104 = n4984 & ~n4986 ;
  assign n5105 = ~n5103 & ~n5104 ;
  assign n5106 = n5102 & ~n5105 ;
  assign n5107 = ~n4075 & ~n4244 ;
  assign n5108 = ~n4930 & n5107 ;
  assign n5109 = n4930 & ~n5107 ;
  assign n5110 = n4930 & ~n4975 ;
  assign n5111 = ~n4930 & n4975 ;
  assign n5112 = ~n5110 & ~n5111 ;
  assign n5113 = n4930 & n4975 ;
  assign n5114 = n4759 & ~n5113 ;
  assign n5115 = n5112 & ~n5114 ;
  assign n5116 = ~n4325 & n5115 ;
  assign n5117 = ~n4977 & ~n5112 ;
  assign n5118 = n4325 & ~n4977 ;
  assign n5119 = ~n5117 & ~n5118 ;
  assign n5120 = ~n5116 & n5119 ;
  assign n5121 = ~n5108 & n5120 ;
  assign n5122 = ~n5109 & n5121 ;
  assign n5123 = ~n5108 & ~n5122 ;
  assign n5124 = ~n5102 & n5105 ;
  assign n5125 = ~n5106 & ~n5124 ;
  assign n5126 = ~n5123 & n5125 ;
  assign n5127 = ~n5106 & ~n5126 ;
  assign n5128 = ~n4329 & n5041 ;
  assign n5129 = n4329 & n4999 ;
  assign n5130 = n4477 & n5044 ;
  assign n5131 = ~n4477 & n4997 ;
  assign n5132 = ~n5130 & ~n5131 ;
  assign n5133 = ~n5129 & n5132 ;
  assign n5134 = ~n5128 & n5133 ;
  assign n5135 = ~n4469 & n4833 ;
  assign n5136 = n4469 & n4668 ;
  assign n5137 = n4640 & n4836 ;
  assign n5138 = ~n4640 & n4666 ;
  assign n5139 = ~n5137 & ~n5138 ;
  assign n5140 = ~n5136 & n5139 ;
  assign n5141 = ~n5135 & n5140 ;
  assign n5142 = n5134 & n5141 ;
  assign n5143 = ~n4632 & n4644 ;
  assign n5144 = n4500 & n4632 ;
  assign n5145 = n4647 & n4821 ;
  assign n5146 = n4498 & ~n4821 ;
  assign n5147 = ~n5145 & ~n5146 ;
  assign n5148 = ~n5144 & n5147 ;
  assign n5149 = ~n5143 & n5148 ;
  assign n5150 = n5134 & ~n5141 ;
  assign n5151 = ~n5134 & n5141 ;
  assign n5152 = ~n5150 & ~n5151 ;
  assign n5153 = n5149 & ~n5152 ;
  assign n5154 = ~n5142 & ~n5153 ;
  assign n5155 = ~n5049 & n5066 ;
  assign n5156 = ~n5067 & ~n5155 ;
  assign n5157 = ~n5154 & n5156 ;
  assign n5158 = n4484 & ~n4813 ;
  assign n5159 = n4345 & n4813 ;
  assign n5160 = n4487 & n4983 ;
  assign n5161 = n4342 & ~n4983 ;
  assign n5162 = ~n5160 & ~n5161 ;
  assign n5163 = ~n5159 & n5162 ;
  assign n5164 = ~n5158 & n5163 ;
  assign n5165 = ~n4079 & ~n4244 ;
  assign n5166 = ~n4930 & n5165 ;
  assign n5167 = n4930 & ~n5165 ;
  assign n5168 = ~n5112 & ~n5114 ;
  assign n5169 = ~n4325 & n5168 ;
  assign n5170 = n4325 & n5117 ;
  assign n5171 = ~n4977 & n5112 ;
  assign n5172 = n4329 & n5171 ;
  assign n5173 = ~n4329 & n5115 ;
  assign n5174 = ~n5172 & ~n5173 ;
  assign n5175 = ~n5170 & n5174 ;
  assign n5176 = ~n5169 & n5175 ;
  assign n5177 = ~n5166 & n5176 ;
  assign n5178 = ~n5167 & n5177 ;
  assign n5179 = ~n5166 & ~n5178 ;
  assign n5180 = n5164 & ~n5179 ;
  assign n5181 = ~n5164 & n5179 ;
  assign n5182 = ~n5180 & ~n5181 ;
  assign n5183 = ~n4640 & n4833 ;
  assign n5184 = n4640 & n4668 ;
  assign n5185 = n4632 & n4836 ;
  assign n5186 = ~n4632 & n4666 ;
  assign n5187 = ~n5185 & ~n5186 ;
  assign n5188 = ~n5184 & n5187 ;
  assign n5189 = ~n5183 & n5188 ;
  assign n5190 = ~n4477 & n5041 ;
  assign n5191 = n4477 & n4999 ;
  assign n5192 = n4469 & n5044 ;
  assign n5193 = ~n4469 & n4997 ;
  assign n5194 = ~n5192 & ~n5193 ;
  assign n5195 = ~n5191 & n5194 ;
  assign n5196 = ~n5190 & n5195 ;
  assign n5197 = n5189 & n5196 ;
  assign n5198 = n4644 & ~n4821 ;
  assign n5199 = n4500 & n4821 ;
  assign n5200 = n4647 & n4813 ;
  assign n5201 = n4498 & ~n4813 ;
  assign n5202 = ~n5200 & ~n5201 ;
  assign n5203 = ~n5199 & n5202 ;
  assign n5204 = ~n5198 & n5203 ;
  assign n5205 = ~n5189 & n5196 ;
  assign n5206 = n5189 & ~n5196 ;
  assign n5207 = ~n5205 & ~n5206 ;
  assign n5208 = n5204 & ~n5207 ;
  assign n5209 = ~n5197 & ~n5208 ;
  assign n5210 = n5182 & ~n5209 ;
  assign n5211 = ~n5180 & ~n5210 ;
  assign n5212 = n5154 & ~n5156 ;
  assign n5213 = ~n5157 & ~n5212 ;
  assign n5214 = ~n5211 & n5213 ;
  assign n5215 = ~n5157 & ~n5214 ;
  assign n5216 = ~n5127 & ~n5215 ;
  assign n5217 = ~n5127 & ~n5216 ;
  assign n5218 = ~n5215 & ~n5216 ;
  assign n5219 = ~n5217 & ~n5218 ;
  assign n5220 = n5077 & ~n5078 ;
  assign n5221 = ~n5075 & ~n5078 ;
  assign n5222 = ~n5220 & ~n5221 ;
  assign n5223 = ~n5219 & ~n5222 ;
  assign n5224 = ~n5216 & ~n5223 ;
  assign n5225 = ~n5086 & n5089 ;
  assign n5226 = n5086 & ~n5089 ;
  assign n5227 = ~n5225 & ~n5226 ;
  assign n5228 = ~n5224 & ~n5227 ;
  assign n5229 = ~n5219 & ~n5223 ;
  assign n5230 = ~n5222 & ~n5223 ;
  assign n5231 = ~n5229 & ~n5230 ;
  assign n5232 = ~n5109 & n5123 ;
  assign n5233 = n5120 & ~n5122 ;
  assign n5234 = ~n5232 & ~n5233 ;
  assign n5235 = n5149 & ~n5153 ;
  assign n5236 = ~n5152 & ~n5153 ;
  assign n5237 = ~n5235 & ~n5236 ;
  assign n5238 = ~n5234 & ~n5237 ;
  assign n5239 = ~n5234 & ~n5238 ;
  assign n5240 = ~n5237 & ~n5238 ;
  assign n5241 = ~n5239 & ~n5240 ;
  assign n5242 = n4484 & ~n4983 ;
  assign n5243 = n4345 & n4983 ;
  assign n5244 = n4075 & n4487 ;
  assign n5245 = ~n4075 & n4342 ;
  assign n5246 = ~n5244 & ~n5245 ;
  assign n5247 = ~n5243 & n5246 ;
  assign n5248 = ~n5242 & n5247 ;
  assign n5249 = ~n4086 & ~n4244 ;
  assign n5250 = ~n4021 & n4609 ;
  assign n5251 = ~n3974 & n5250 ;
  assign n5252 = ~n4100 & n5251 ;
  assign n5253 = ~n3923 & n5252 ;
  assign n5254 = ~n4012 & n5253 ;
  assign n5255 = ~n4147 & n5254 ;
  assign n5256 = ~n4352 & n5255 ;
  assign n5257 = ~n4353 & n5256 ;
  assign n5258 = ~n4020 & ~n4150 ;
  assign n5259 = ~n4115 & n5258 ;
  assign n5260 = n4232 & n4384 ;
  assign n5261 = n5259 & n5260 ;
  assign n5262 = n4768 & n5261 ;
  assign n5263 = n4444 & n5262 ;
  assign n5264 = ~n4137 & n5263 ;
  assign n5265 = ~n4014 & n5264 ;
  assign n5266 = ~n4217 & n5265 ;
  assign n5267 = ~n4034 & n5266 ;
  assign n5268 = ~n4167 & n5267 ;
  assign n5269 = ~n4124 & ~n4160 ;
  assign n5270 = ~n4246 & n5269 ;
  assign n5271 = ~n3972 & n5270 ;
  assign n5272 = ~n4303 & n5271 ;
  assign n5273 = ~n4156 & n5272 ;
  assign n5274 = ~n4016 & n5273 ;
  assign n5275 = ~n4142 & n5274 ;
  assign n5276 = ~n3954 & n5275 ;
  assign n5277 = n4173 & n5276 ;
  assign n5278 = n5268 & n5277 ;
  assign n5279 = n4221 & n5278 ;
  assign n5280 = n5257 & n5279 ;
  assign n5281 = ~n3978 & n5280 ;
  assign n5282 = ~n4008 & n5281 ;
  assign n5283 = ~n3918 & n5282 ;
  assign n5284 = ~n4161 & n5283 ;
  assign n5285 = ~n4058 & n5284 ;
  assign n5286 = ~n4399 & n5285 ;
  assign n5287 = ~n4011 & n5286 ;
  assign n5288 = ~n4325 & n5287 ;
  assign n5289 = ~n4930 & ~n5288 ;
  assign n5290 = n5249 & n5289 ;
  assign n5291 = ~n4329 & n5168 ;
  assign n5292 = n4329 & n5117 ;
  assign n5293 = n4477 & n5171 ;
  assign n5294 = ~n4477 & n5115 ;
  assign n5295 = ~n5293 & ~n5294 ;
  assign n5296 = ~n5292 & n5295 ;
  assign n5297 = ~n5291 & n5296 ;
  assign n5298 = ~n5249 & ~n5289 ;
  assign n5299 = ~n5290 & ~n5298 ;
  assign n5300 = n5297 & n5299 ;
  assign n5301 = ~n5290 & ~n5300 ;
  assign n5302 = n5248 & ~n5301 ;
  assign n5303 = ~n5248 & n5301 ;
  assign n5304 = ~n5302 & ~n5303 ;
  assign n5305 = ~n4632 & n4833 ;
  assign n5306 = n4632 & n4668 ;
  assign n5307 = n4821 & n4836 ;
  assign n5308 = n4666 & ~n4821 ;
  assign n5309 = ~n5307 & ~n5308 ;
  assign n5310 = ~n5306 & n5309 ;
  assign n5311 = ~n5305 & n5310 ;
  assign n5312 = ~n4469 & n5041 ;
  assign n5313 = n4469 & n4999 ;
  assign n5314 = n4640 & n5044 ;
  assign n5315 = ~n4640 & n4997 ;
  assign n5316 = ~n5314 & ~n5315 ;
  assign n5317 = ~n5313 & n5316 ;
  assign n5318 = ~n5312 & n5317 ;
  assign n5319 = n5311 & n5318 ;
  assign n5320 = n4644 & ~n4813 ;
  assign n5321 = n4500 & n4813 ;
  assign n5322 = n4647 & n4983 ;
  assign n5323 = n4498 & ~n4983 ;
  assign n5324 = ~n5322 & ~n5323 ;
  assign n5325 = ~n5321 & n5324 ;
  assign n5326 = ~n5320 & n5325 ;
  assign n5327 = ~n5311 & n5318 ;
  assign n5328 = n5311 & ~n5318 ;
  assign n5329 = ~n5327 & ~n5328 ;
  assign n5330 = n5326 & ~n5329 ;
  assign n5331 = ~n5319 & ~n5330 ;
  assign n5332 = n5304 & ~n5331 ;
  assign n5333 = ~n5302 & ~n5332 ;
  assign n5334 = ~n5241 & ~n5333 ;
  assign n5335 = ~n5238 & ~n5334 ;
  assign n5336 = n5123 & ~n5125 ;
  assign n5337 = ~n5126 & ~n5336 ;
  assign n5338 = ~n5335 & n5337 ;
  assign n5339 = n5335 & ~n5337 ;
  assign n5340 = ~n5338 & ~n5339 ;
  assign n5341 = n5211 & ~n5213 ;
  assign n5342 = ~n5214 & ~n5341 ;
  assign n5343 = n5340 & n5342 ;
  assign n5344 = ~n5338 & ~n5343 ;
  assign n5345 = ~n5231 & ~n5344 ;
  assign n5346 = n5231 & ~n5344 ;
  assign n5347 = ~n5231 & n5344 ;
  assign n5348 = ~n5346 & ~n5347 ;
  assign n5349 = n4930 & ~n5287 ;
  assign n5350 = ~n5287 & ~n5349 ;
  assign n5351 = ~n4325 & n5350 ;
  assign n5352 = n4325 & n5349 ;
  assign n5353 = n4329 & ~n4930 ;
  assign n5354 = n5287 & ~n5353 ;
  assign n5355 = ~n5352 & ~n5354 ;
  assign n5356 = ~n5351 & n5355 ;
  assign n5357 = ~n4086 & n4484 ;
  assign n5358 = n4086 & ~n4344 ;
  assign n5359 = ~n4487 & ~n5358 ;
  assign n5360 = ~n5357 & n5359 ;
  assign n5361 = n4344 & n5360 ;
  assign n5362 = n5356 & n5361 ;
  assign n5363 = ~n4075 & n4484 ;
  assign n5364 = n4075 & n4345 ;
  assign n5365 = n4079 & n4487 ;
  assign n5366 = ~n4079 & n4342 ;
  assign n5367 = ~n5365 & ~n5366 ;
  assign n5368 = ~n5364 & n5367 ;
  assign n5369 = ~n5363 & n5368 ;
  assign n5370 = n5362 & n5369 ;
  assign n5371 = ~n4640 & n5041 ;
  assign n5372 = n4640 & n4999 ;
  assign n5373 = n4632 & n5044 ;
  assign n5374 = ~n4632 & n4997 ;
  assign n5375 = ~n5373 & ~n5374 ;
  assign n5376 = ~n5372 & n5375 ;
  assign n5377 = ~n5371 & n5376 ;
  assign n5378 = ~n4821 & n4833 ;
  assign n5379 = n4668 & n4821 ;
  assign n5380 = n4813 & n4836 ;
  assign n5381 = n4666 & ~n4813 ;
  assign n5382 = ~n5380 & ~n5381 ;
  assign n5383 = ~n5379 & n5382 ;
  assign n5384 = ~n5378 & n5383 ;
  assign n5385 = n4644 & ~n4983 ;
  assign n5386 = n4500 & n4983 ;
  assign n5387 = n4075 & n4647 ;
  assign n5388 = ~n4075 & n4498 ;
  assign n5389 = ~n5387 & ~n5388 ;
  assign n5390 = ~n5386 & n5389 ;
  assign n5391 = ~n5385 & n5390 ;
  assign n5392 = n5384 & ~n5391 ;
  assign n5393 = ~n5384 & n5391 ;
  assign n5394 = ~n5392 & ~n5393 ;
  assign n5395 = n5377 & ~n5394 ;
  assign n5396 = n5384 & n5391 ;
  assign n5397 = ~n5395 & ~n5396 ;
  assign n5398 = ~n5362 & ~n5369 ;
  assign n5399 = ~n5370 & ~n5398 ;
  assign n5400 = ~n5397 & n5399 ;
  assign n5401 = ~n5370 & ~n5400 ;
  assign n5402 = ~n5167 & n5179 ;
  assign n5403 = n5176 & ~n5178 ;
  assign n5404 = ~n5402 & ~n5403 ;
  assign n5405 = n5401 & ~n5404 ;
  assign n5406 = ~n5401 & n5404 ;
  assign n5407 = ~n5405 & ~n5406 ;
  assign n5408 = n5204 & ~n5208 ;
  assign n5409 = ~n5207 & ~n5208 ;
  assign n5410 = ~n5408 & ~n5409 ;
  assign n5411 = ~n5407 & ~n5410 ;
  assign n5412 = ~n5401 & ~n5404 ;
  assign n5413 = ~n5411 & ~n5412 ;
  assign n5414 = ~n5182 & n5209 ;
  assign n5415 = ~n5210 & ~n5414 ;
  assign n5416 = ~n5413 & n5415 ;
  assign n5417 = n5241 & ~n5333 ;
  assign n5418 = ~n5241 & n5333 ;
  assign n5419 = ~n5417 & ~n5418 ;
  assign n5420 = n5413 & ~n5415 ;
  assign n5421 = ~n5416 & ~n5420 ;
  assign n5422 = ~n5419 & n5421 ;
  assign n5423 = ~n5416 & ~n5422 ;
  assign n5424 = ~n5340 & ~n5342 ;
  assign n5425 = ~n5343 & ~n5424 ;
  assign n5426 = ~n5423 & n5425 ;
  assign n5427 = ~n4477 & n5168 ;
  assign n5428 = n4477 & n5117 ;
  assign n5429 = n4469 & n5171 ;
  assign n5430 = ~n4469 & n5115 ;
  assign n5431 = ~n5429 & ~n5430 ;
  assign n5432 = ~n5428 & n5431 ;
  assign n5433 = ~n5427 & n5432 ;
  assign n5434 = ~n4079 & n4484 ;
  assign n5435 = n4079 & n4345 ;
  assign n5436 = n4086 & n4487 ;
  assign n5437 = ~n4086 & n4342 ;
  assign n5438 = ~n5436 & ~n5437 ;
  assign n5439 = ~n5435 & n5438 ;
  assign n5440 = ~n5434 & n5439 ;
  assign n5441 = n5433 & n5440 ;
  assign n5442 = ~n5356 & ~n5361 ;
  assign n5443 = ~n5362 & ~n5442 ;
  assign n5444 = ~n5433 & ~n5440 ;
  assign n5445 = ~n5441 & ~n5444 ;
  assign n5446 = n5443 & n5445 ;
  assign n5447 = ~n5441 & ~n5446 ;
  assign n5448 = ~n5297 & ~n5299 ;
  assign n5449 = ~n5300 & ~n5448 ;
  assign n5450 = ~n5447 & n5449 ;
  assign n5451 = n5447 & ~n5449 ;
  assign n5452 = ~n5450 & ~n5451 ;
  assign n5453 = n5326 & ~n5330 ;
  assign n5454 = ~n5329 & ~n5330 ;
  assign n5455 = ~n5453 & ~n5454 ;
  assign n5456 = n5452 & ~n5455 ;
  assign n5457 = ~n5450 & ~n5456 ;
  assign n5458 = ~n5304 & n5331 ;
  assign n5459 = ~n5332 & ~n5458 ;
  assign n5460 = ~n5457 & n5459 ;
  assign n5461 = n5457 & ~n5459 ;
  assign n5462 = ~n5460 & ~n5461 ;
  assign n5463 = n5407 & n5410 ;
  assign n5464 = ~n5411 & ~n5463 ;
  assign n5465 = n5462 & n5464 ;
  assign n5466 = ~n5460 & ~n5465 ;
  assign n5467 = n5419 & ~n5421 ;
  assign n5468 = ~n5422 & ~n5467 ;
  assign n5469 = ~n5466 & n5468 ;
  assign n5470 = ~n4477 & n5350 ;
  assign n5471 = n4477 & n5349 ;
  assign n5472 = n4469 & ~n4930 ;
  assign n5473 = n5287 & ~n5472 ;
  assign n5474 = ~n5471 & ~n5473 ;
  assign n5475 = ~n5470 & n5474 ;
  assign n5476 = ~n4086 & n4644 ;
  assign n5477 = n4086 & ~n4465 ;
  assign n5478 = ~n4647 & ~n5477 ;
  assign n5479 = ~n5476 & n5478 ;
  assign n5480 = n4465 & n5479 ;
  assign n5481 = n5475 & n5480 ;
  assign n5482 = ~n4632 & n5041 ;
  assign n5483 = n4632 & n4999 ;
  assign n5484 = n4821 & n5044 ;
  assign n5485 = ~n4821 & n4997 ;
  assign n5486 = ~n5484 & ~n5485 ;
  assign n5487 = ~n5483 & n5486 ;
  assign n5488 = ~n5482 & n5487 ;
  assign n5489 = ~n4813 & n4833 ;
  assign n5490 = n4668 & n4813 ;
  assign n5491 = n4836 & n4983 ;
  assign n5492 = n4666 & ~n4983 ;
  assign n5493 = ~n5491 & ~n5492 ;
  assign n5494 = ~n5490 & n5493 ;
  assign n5495 = ~n5489 & n5494 ;
  assign n5496 = n5488 & ~n5495 ;
  assign n5497 = ~n5488 & n5495 ;
  assign n5498 = ~n5496 & ~n5497 ;
  assign n5499 = n5481 & ~n5498 ;
  assign n5500 = n5488 & n5495 ;
  assign n5501 = ~n5499 & ~n5500 ;
  assign n5502 = ~n4075 & n4644 ;
  assign n5503 = n4075 & n4500 ;
  assign n5504 = n4079 & n4647 ;
  assign n5505 = ~n4079 & n4498 ;
  assign n5506 = ~n5504 & ~n5505 ;
  assign n5507 = ~n5503 & n5506 ;
  assign n5508 = ~n5502 & n5507 ;
  assign n5509 = ~n4329 & n5350 ;
  assign n5510 = n4329 & n5349 ;
  assign n5511 = n4477 & ~n4930 ;
  assign n5512 = n5287 & ~n5511 ;
  assign n5513 = ~n5510 & ~n5512 ;
  assign n5514 = ~n5509 & n5513 ;
  assign n5515 = ~n4469 & n5168 ;
  assign n5516 = n4469 & n5117 ;
  assign n5517 = n4640 & n5171 ;
  assign n5518 = ~n4640 & n5115 ;
  assign n5519 = ~n5517 & ~n5518 ;
  assign n5520 = ~n5516 & n5519 ;
  assign n5521 = ~n5515 & n5520 ;
  assign n5522 = n5514 & ~n5521 ;
  assign n5523 = ~n5514 & n5521 ;
  assign n5524 = ~n5522 & ~n5523 ;
  assign n5525 = n5508 & ~n5524 ;
  assign n5526 = n5514 & n5521 ;
  assign n5527 = ~n5525 & ~n5526 ;
  assign n5528 = ~n5501 & ~n5527 ;
  assign n5529 = ~n5501 & ~n5528 ;
  assign n5530 = ~n5527 & ~n5528 ;
  assign n5531 = ~n5529 & ~n5530 ;
  assign n5532 = n5377 & ~n5395 ;
  assign n5533 = ~n5394 & ~n5395 ;
  assign n5534 = ~n5532 & ~n5533 ;
  assign n5535 = ~n5531 & ~n5534 ;
  assign n5536 = ~n5528 & ~n5535 ;
  assign n5537 = n5397 & ~n5399 ;
  assign n5538 = ~n5400 & ~n5537 ;
  assign n5539 = ~n5536 & n5538 ;
  assign n5540 = n5452 & ~n5456 ;
  assign n5541 = ~n5455 & ~n5456 ;
  assign n5542 = ~n5540 & ~n5541 ;
  assign n5543 = n5536 & ~n5538 ;
  assign n5544 = ~n5539 & ~n5543 ;
  assign n5545 = ~n5542 & n5544 ;
  assign n5546 = ~n5539 & ~n5545 ;
  assign n5547 = ~n5462 & ~n5464 ;
  assign n5548 = ~n5465 & ~n5547 ;
  assign n5549 = ~n5546 & n5548 ;
  assign n5550 = ~n4344 & ~n5360 ;
  assign n5551 = ~n4821 & n5041 ;
  assign n5552 = n4821 & n4999 ;
  assign n5553 = n4813 & n5044 ;
  assign n5554 = ~n4813 & n4997 ;
  assign n5555 = ~n5553 & ~n5554 ;
  assign n5556 = ~n5552 & n5555 ;
  assign n5557 = ~n5551 & n5556 ;
  assign n5558 = ~n4640 & n5168 ;
  assign n5559 = n4640 & n5117 ;
  assign n5560 = n4632 & n5171 ;
  assign n5561 = ~n4632 & n5115 ;
  assign n5562 = ~n5560 & ~n5561 ;
  assign n5563 = ~n5559 & n5562 ;
  assign n5564 = ~n5558 & n5563 ;
  assign n5565 = n4833 & ~n4983 ;
  assign n5566 = n4668 & n4983 ;
  assign n5567 = n4075 & n4836 ;
  assign n5568 = ~n4075 & n4666 ;
  assign n5569 = ~n5567 & ~n5568 ;
  assign n5570 = ~n5566 & n5569 ;
  assign n5571 = ~n5565 & n5570 ;
  assign n5572 = n5564 & ~n5571 ;
  assign n5573 = ~n5564 & n5571 ;
  assign n5574 = ~n5572 & ~n5573 ;
  assign n5575 = n5557 & ~n5574 ;
  assign n5576 = n5564 & n5571 ;
  assign n5577 = ~n5575 & ~n5576 ;
  assign n5578 = ~n5361 & ~n5577 ;
  assign n5579 = ~n5550 & n5578 ;
  assign n5580 = ~n5361 & ~n5579 ;
  assign n5581 = ~n5550 & n5580 ;
  assign n5582 = ~n5577 & ~n5579 ;
  assign n5583 = ~n5581 & ~n5582 ;
  assign n5584 = ~n5481 & n5498 ;
  assign n5585 = ~n5499 & ~n5584 ;
  assign n5586 = ~n5583 & n5585 ;
  assign n5587 = ~n5579 & ~n5586 ;
  assign n5588 = n5443 & ~n5446 ;
  assign n5589 = ~n5444 & n5447 ;
  assign n5590 = ~n5588 & ~n5589 ;
  assign n5591 = ~n5587 & n5590 ;
  assign n5592 = n5587 & ~n5590 ;
  assign n5593 = ~n5591 & ~n5592 ;
  assign n5594 = ~n5531 & ~n5535 ;
  assign n5595 = ~n5534 & ~n5535 ;
  assign n5596 = ~n5594 & ~n5595 ;
  assign n5597 = ~n5593 & ~n5596 ;
  assign n5598 = ~n5587 & ~n5590 ;
  assign n5599 = ~n5597 & ~n5598 ;
  assign n5600 = n5542 & ~n5544 ;
  assign n5601 = ~n5545 & ~n5600 ;
  assign n5602 = ~n5599 & n5601 ;
  assign n5603 = ~n4469 & n5350 ;
  assign n5604 = n4469 & n5349 ;
  assign n5605 = n4640 & ~n4930 ;
  assign n5606 = n5287 & ~n5605 ;
  assign n5607 = ~n5604 & ~n5606 ;
  assign n5608 = ~n5603 & n5607 ;
  assign n5609 = ~n4632 & n5168 ;
  assign n5610 = n4632 & n5117 ;
  assign n5611 = n4821 & n5171 ;
  assign n5612 = ~n4821 & n5115 ;
  assign n5613 = ~n5611 & ~n5612 ;
  assign n5614 = ~n5610 & n5613 ;
  assign n5615 = ~n5609 & n5614 ;
  assign n5616 = n5608 & n5615 ;
  assign n5617 = ~n4813 & n5041 ;
  assign n5618 = n4813 & n4999 ;
  assign n5619 = n4983 & n5044 ;
  assign n5620 = ~n4983 & n4997 ;
  assign n5621 = ~n5619 & ~n5620 ;
  assign n5622 = ~n5618 & n5621 ;
  assign n5623 = ~n5617 & n5622 ;
  assign n5624 = n5608 & ~n5615 ;
  assign n5625 = ~n5608 & n5615 ;
  assign n5626 = ~n5624 & ~n5625 ;
  assign n5627 = n5623 & ~n5626 ;
  assign n5628 = ~n5616 & ~n5627 ;
  assign n5629 = ~n4079 & n4644 ;
  assign n5630 = n4079 & n4500 ;
  assign n5631 = n4086 & n4647 ;
  assign n5632 = ~n4086 & n4498 ;
  assign n5633 = ~n5631 & ~n5632 ;
  assign n5634 = ~n5630 & n5633 ;
  assign n5635 = ~n5629 & n5634 ;
  assign n5636 = ~n5475 & ~n5480 ;
  assign n5637 = ~n5481 & ~n5636 ;
  assign n5638 = n5635 & ~n5637 ;
  assign n5639 = ~n5635 & n5637 ;
  assign n5640 = ~n5638 & ~n5639 ;
  assign n5641 = ~n5628 & ~n5640 ;
  assign n5642 = n5635 & n5637 ;
  assign n5643 = ~n5641 & ~n5642 ;
  assign n5644 = n5508 & ~n5525 ;
  assign n5645 = ~n5524 & ~n5525 ;
  assign n5646 = ~n5644 & ~n5645 ;
  assign n5647 = ~n5643 & ~n5646 ;
  assign n5648 = ~n5583 & ~n5586 ;
  assign n5649 = n5585 & ~n5586 ;
  assign n5650 = ~n5648 & ~n5649 ;
  assign n5651 = ~n5643 & ~n5647 ;
  assign n5652 = ~n5646 & ~n5647 ;
  assign n5653 = ~n5651 & ~n5652 ;
  assign n5654 = ~n5650 & ~n5653 ;
  assign n5655 = ~n5647 & ~n5654 ;
  assign n5656 = ~n4075 & n4833 ;
  assign n5657 = n4075 & n4668 ;
  assign n5658 = n4079 & n4836 ;
  assign n5659 = ~n4079 & n4666 ;
  assign n5660 = ~n5658 & ~n5659 ;
  assign n5661 = ~n5657 & n5660 ;
  assign n5662 = ~n5656 & n5661 ;
  assign n5663 = ~n4640 & n5350 ;
  assign n5664 = n4640 & n5349 ;
  assign n5665 = n4632 & ~n4930 ;
  assign n5666 = n5287 & ~n5665 ;
  assign n5667 = ~n5664 & ~n5666 ;
  assign n5668 = ~n5663 & n5667 ;
  assign n5669 = ~n4086 & n4833 ;
  assign n5670 = n4086 & ~n4628 ;
  assign n5671 = ~n4836 & ~n5670 ;
  assign n5672 = ~n5669 & n5671 ;
  assign n5673 = n4628 & n5672 ;
  assign n5674 = n5668 & n5673 ;
  assign n5675 = n5662 & n5674 ;
  assign n5676 = ~n5662 & n5674 ;
  assign n5677 = n5662 & ~n5674 ;
  assign n5678 = ~n5676 & ~n5677 ;
  assign n5679 = ~n4086 & ~n4495 ;
  assign n5680 = ~n5678 & n5679 ;
  assign n5681 = ~n5675 & ~n5680 ;
  assign n5682 = ~n5557 & n5574 ;
  assign n5683 = ~n5575 & ~n5682 ;
  assign n5684 = ~n5681 & n5683 ;
  assign n5685 = n5681 & ~n5683 ;
  assign n5686 = ~n5684 & ~n5685 ;
  assign n5687 = n5628 & n5640 ;
  assign n5688 = ~n5641 & ~n5687 ;
  assign n5689 = ~n5686 & ~n5688 ;
  assign n5690 = n5686 & n5688 ;
  assign n5691 = ~n4079 & n4833 ;
  assign n5692 = n4079 & n4668 ;
  assign n5693 = n4086 & n4836 ;
  assign n5694 = ~n4086 & n4666 ;
  assign n5695 = ~n5693 & ~n5694 ;
  assign n5696 = ~n5692 & n5695 ;
  assign n5697 = ~n5691 & n5696 ;
  assign n5698 = ~n4821 & n5168 ;
  assign n5699 = n4821 & n5117 ;
  assign n5700 = n4813 & n5171 ;
  assign n5701 = ~n4813 & n5115 ;
  assign n5702 = ~n5700 & ~n5701 ;
  assign n5703 = ~n5699 & n5702 ;
  assign n5704 = ~n5698 & n5703 ;
  assign n5705 = ~n4983 & n5041 ;
  assign n5706 = n4983 & n4999 ;
  assign n5707 = n4075 & n5044 ;
  assign n5708 = ~n4075 & n4997 ;
  assign n5709 = ~n5707 & ~n5708 ;
  assign n5710 = ~n5706 & n5709 ;
  assign n5711 = ~n5705 & n5710 ;
  assign n5712 = n5704 & ~n5711 ;
  assign n5713 = ~n5704 & n5711 ;
  assign n5714 = ~n5712 & ~n5713 ;
  assign n5715 = n5697 & ~n5714 ;
  assign n5716 = n5704 & n5711 ;
  assign n5717 = ~n5715 & ~n5716 ;
  assign n5718 = ~n5623 & n5626 ;
  assign n5719 = ~n5627 & ~n5718 ;
  assign n5720 = ~n5717 & n5719 ;
  assign n5721 = n5678 & ~n5679 ;
  assign n5722 = ~n5680 & ~n5721 ;
  assign n5723 = ~n5717 & ~n5720 ;
  assign n5724 = n5719 & ~n5720 ;
  assign n5725 = ~n5723 & ~n5724 ;
  assign n5726 = n5722 & ~n5725 ;
  assign n5727 = ~n5720 & ~n5726 ;
  assign n5728 = ~n4628 & ~n5672 ;
  assign n5729 = ~n4821 & n5350 ;
  assign n5730 = n4821 & n5349 ;
  assign n5731 = n4813 & ~n4930 ;
  assign n5732 = n5287 & ~n5731 ;
  assign n5733 = ~n5730 & ~n5732 ;
  assign n5734 = ~n5729 & n5733 ;
  assign n5735 = ~n4086 & n5041 ;
  assign n5736 = n4086 & ~n4809 ;
  assign n5737 = ~n5044 & ~n5736 ;
  assign n5738 = ~n5735 & n5737 ;
  assign n5739 = n4809 & n5738 ;
  assign n5740 = n5734 & n5739 ;
  assign n5741 = ~n5673 & n5740 ;
  assign n5742 = ~n5728 & n5741 ;
  assign n5743 = ~n4983 & n5168 ;
  assign n5744 = n4983 & n5117 ;
  assign n5745 = n4075 & n5171 ;
  assign n5746 = ~n4075 & n5115 ;
  assign n5747 = ~n5745 & ~n5746 ;
  assign n5748 = ~n5744 & n5747 ;
  assign n5749 = ~n5743 & n5748 ;
  assign n5750 = ~n4079 & n5041 ;
  assign n5751 = n4079 & n4999 ;
  assign n5752 = n4086 & n5044 ;
  assign n5753 = ~n4086 & n4997 ;
  assign n5754 = ~n5752 & ~n5753 ;
  assign n5755 = ~n5751 & n5754 ;
  assign n5756 = ~n5750 & n5755 ;
  assign n5757 = n5749 & n5756 ;
  assign n5758 = ~n5734 & ~n5739 ;
  assign n5759 = ~n5740 & ~n5758 ;
  assign n5760 = ~n5749 & ~n5756 ;
  assign n5761 = ~n5757 & ~n5760 ;
  assign n5762 = n5759 & n5761 ;
  assign n5763 = ~n5757 & ~n5762 ;
  assign n5764 = n5740 & ~n5742 ;
  assign n5765 = ~n5673 & ~n5742 ;
  assign n5766 = ~n5728 & n5765 ;
  assign n5767 = ~n5764 & ~n5766 ;
  assign n5768 = ~n5763 & ~n5767 ;
  assign n5769 = ~n5742 & ~n5768 ;
  assign n5770 = ~n4075 & n5041 ;
  assign n5771 = n4075 & n4999 ;
  assign n5772 = n4079 & n5044 ;
  assign n5773 = ~n4079 & n4997 ;
  assign n5774 = ~n5772 & ~n5773 ;
  assign n5775 = ~n5771 & n5774 ;
  assign n5776 = ~n5770 & n5775 ;
  assign n5777 = ~n4813 & n5168 ;
  assign n5778 = n4813 & n5117 ;
  assign n5779 = n4983 & n5171 ;
  assign n5780 = ~n4983 & n5115 ;
  assign n5781 = ~n5779 & ~n5780 ;
  assign n5782 = ~n5778 & n5781 ;
  assign n5783 = ~n5777 & n5782 ;
  assign n5784 = ~n4632 & n5350 ;
  assign n5785 = n4632 & n5349 ;
  assign n5786 = n4821 & ~n4930 ;
  assign n5787 = n5287 & ~n5786 ;
  assign n5788 = ~n5785 & ~n5787 ;
  assign n5789 = ~n5784 & n5788 ;
  assign n5790 = ~n5783 & n5789 ;
  assign n5791 = n5783 & ~n5789 ;
  assign n5792 = ~n5790 & ~n5791 ;
  assign n5793 = ~n5776 & n5792 ;
  assign n5794 = n5776 & ~n5792 ;
  assign n5795 = ~n4813 & n5350 ;
  assign n5796 = n4813 & n5349 ;
  assign n5797 = ~n4930 & n4983 ;
  assign n5798 = n5287 & ~n5797 ;
  assign n5799 = ~n5796 & ~n5798 ;
  assign n5800 = ~n5795 & n5799 ;
  assign n5801 = ~n4075 & n5168 ;
  assign n5802 = n4075 & n5117 ;
  assign n5803 = n4079 & n5171 ;
  assign n5804 = ~n4079 & n5115 ;
  assign n5805 = ~n5803 & ~n5804 ;
  assign n5806 = ~n5802 & n5805 ;
  assign n5807 = ~n5801 & n5806 ;
  assign n5808 = n5800 & ~n5807 ;
  assign n5809 = ~n5800 & n5807 ;
  assign n5810 = ~n5808 & ~n5809 ;
  assign n5811 = ~n4983 & n5350 ;
  assign n5812 = n4983 & n5349 ;
  assign n5813 = n4075 & ~n4930 ;
  assign n5814 = n5287 & ~n5813 ;
  assign n5815 = ~n5812 & ~n5814 ;
  assign n5816 = ~n5811 & n5815 ;
  assign n5817 = ~n4086 & n5168 ;
  assign n5818 = n4086 & ~n4977 ;
  assign n5819 = ~n5171 & ~n5818 ;
  assign n5820 = ~n5817 & n5819 ;
  assign n5821 = n4977 & n5820 ;
  assign n5822 = n5816 & n5821 ;
  assign n5823 = n5810 & ~n5822 ;
  assign n5824 = ~n5810 & n5822 ;
  assign n5825 = ~n4079 & n5168 ;
  assign n5826 = n4079 & n5117 ;
  assign n5827 = ~n4086 & n5115 ;
  assign n5828 = ~n4977 & ~n5820 ;
  assign n5829 = ~n4075 & n5350 ;
  assign n5830 = n4075 & n5349 ;
  assign n5831 = ~n4079 & ~n5287 ;
  assign n5832 = n4930 & n5287 ;
  assign n5833 = n4079 & ~n5832 ;
  assign n5834 = ~n5831 & ~n5833 ;
  assign n5835 = ~n5830 & ~n5834 ;
  assign n5836 = ~n5829 & n5835 ;
  assign n5837 = n4086 & ~n4930 ;
  assign n5838 = ~n5831 & n5837 ;
  assign n5839 = ~n5836 & ~n5838 ;
  assign n5840 = ~n5821 & ~n5839 ;
  assign n5841 = ~n5828 & n5840 ;
  assign n5842 = n5836 & n5838 ;
  assign n5843 = ~n5841 & ~n5842 ;
  assign n5844 = ~n5816 & ~n5821 ;
  assign n5845 = ~n5822 & ~n5844 ;
  assign n5846 = n5843 & ~n5845 ;
  assign n5847 = n4086 & n5171 ;
  assign n5848 = ~n5846 & ~n5847 ;
  assign n5849 = ~n5827 & n5848 ;
  assign n5850 = ~n5826 & n5849 ;
  assign n5851 = ~n5825 & n5850 ;
  assign n5852 = ~n5843 & n5845 ;
  assign n5853 = ~n5851 & ~n5852 ;
  assign n5854 = ~n4086 & ~n4994 ;
  assign n5855 = n5853 & ~n5854 ;
  assign n5856 = ~n5824 & ~n5855 ;
  assign n5857 = ~n5823 & n5856 ;
  assign n5858 = ~n5853 & n5854 ;
  assign n5859 = ~n5857 & ~n5858 ;
  assign n5860 = n5759 & ~n5762 ;
  assign n5861 = ~n5760 & n5763 ;
  assign n5862 = ~n5860 & ~n5861 ;
  assign n5863 = n5859 & n5862 ;
  assign n5864 = n5800 & n5807 ;
  assign n5865 = ~n5824 & ~n5864 ;
  assign n5866 = ~n5863 & ~n5865 ;
  assign n5867 = ~n5859 & ~n5862 ;
  assign n5868 = ~n5866 & ~n5867 ;
  assign n5869 = ~n5763 & ~n5768 ;
  assign n5870 = ~n5767 & ~n5768 ;
  assign n5871 = ~n5869 & ~n5870 ;
  assign n5872 = n5868 & n5871 ;
  assign n5873 = ~n5794 & ~n5872 ;
  assign n5874 = ~n5793 & n5873 ;
  assign n5875 = ~n5868 & ~n5871 ;
  assign n5876 = ~n5874 & ~n5875 ;
  assign n5877 = ~n5769 & ~n5876 ;
  assign n5878 = n5769 & n5876 ;
  assign n5879 = n5697 & ~n5715 ;
  assign n5880 = ~n5714 & ~n5715 ;
  assign n5881 = ~n5879 & ~n5880 ;
  assign n5882 = ~n5668 & ~n5673 ;
  assign n5883 = ~n5674 & ~n5882 ;
  assign n5884 = n5783 & n5789 ;
  assign n5885 = ~n5794 & ~n5884 ;
  assign n5886 = n5883 & ~n5885 ;
  assign n5887 = ~n5883 & n5885 ;
  assign n5888 = ~n5886 & ~n5887 ;
  assign n5889 = ~n5881 & n5888 ;
  assign n5890 = n5881 & ~n5888 ;
  assign n5891 = ~n5889 & ~n5890 ;
  assign n5892 = ~n5878 & n5891 ;
  assign n5893 = ~n5877 & ~n5892 ;
  assign n5894 = ~n5886 & ~n5889 ;
  assign n5895 = ~n5893 & ~n5894 ;
  assign n5896 = n5893 & n5894 ;
  assign n5897 = ~n5722 & n5725 ;
  assign n5898 = ~n5726 & ~n5897 ;
  assign n5899 = ~n5896 & n5898 ;
  assign n5900 = ~n5895 & ~n5899 ;
  assign n5901 = n5727 & n5900 ;
  assign n5902 = ~n5690 & ~n5901 ;
  assign n5903 = ~n5689 & n5902 ;
  assign n5904 = ~n5727 & ~n5900 ;
  assign n5905 = ~n5903 & ~n5904 ;
  assign n5906 = ~n5684 & ~n5690 ;
  assign n5907 = ~n5905 & ~n5906 ;
  assign n5908 = n5905 & n5906 ;
  assign n5909 = n5650 & n5653 ;
  assign n5910 = ~n5654 & ~n5909 ;
  assign n5911 = ~n5908 & n5910 ;
  assign n5912 = ~n5907 & ~n5911 ;
  assign n5913 = n5655 & n5912 ;
  assign n5914 = n5593 & n5596 ;
  assign n5915 = ~n5913 & ~n5914 ;
  assign n5916 = ~n5597 & n5915 ;
  assign n5917 = ~n5655 & ~n5912 ;
  assign n5918 = ~n5916 & ~n5917 ;
  assign n5919 = n5599 & ~n5601 ;
  assign n5920 = ~n5602 & ~n5919 ;
  assign n5921 = ~n5918 & n5920 ;
  assign n5922 = ~n5602 & ~n5921 ;
  assign n5923 = n5546 & ~n5548 ;
  assign n5924 = ~n5549 & ~n5923 ;
  assign n5925 = ~n5922 & n5924 ;
  assign n5926 = ~n5549 & ~n5925 ;
  assign n5927 = n5466 & ~n5468 ;
  assign n5928 = ~n5469 & ~n5927 ;
  assign n5929 = ~n5926 & n5928 ;
  assign n5930 = ~n5469 & ~n5929 ;
  assign n5931 = n5423 & ~n5425 ;
  assign n5932 = ~n5426 & ~n5931 ;
  assign n5933 = ~n5930 & n5932 ;
  assign n5934 = ~n5426 & ~n5933 ;
  assign n5935 = ~n5348 & ~n5934 ;
  assign n5936 = ~n5345 & ~n5935 ;
  assign n5937 = n5224 & n5227 ;
  assign n5938 = ~n5228 & ~n5937 ;
  assign n5939 = ~n5936 & n5938 ;
  assign n5940 = ~n5228 & ~n5939 ;
  assign n5941 = ~n5095 & ~n5940 ;
  assign n5942 = ~n5092 & ~n5941 ;
  assign n5943 = n5034 & ~n5036 ;
  assign n5944 = ~n5037 & ~n5943 ;
  assign n5945 = ~n5942 & n5944 ;
  assign n5946 = ~n5037 & ~n5945 ;
  assign n5947 = ~n4874 & ~n5946 ;
  assign n5948 = ~n4868 & ~n4871 ;
  assign n5949 = ~n5947 & ~n5948 ;
  assign n5950 = n4695 & ~n4697 ;
  assign n5951 = ~n4698 & ~n5950 ;
  assign n5952 = ~n5949 & n5951 ;
  assign n5953 = ~n4698 & ~n5952 ;
  assign n5954 = ~n4528 & ~n5953 ;
  assign n5955 = ~n4522 & ~n4525 ;
  assign n5956 = ~n5954 & ~n5955 ;
  assign n5957 = n4483 & ~n5956 ;
  assign n5958 = ~n4483 & n5956 ;
  assign n5959 = ~n5957 & ~n5958 ;
  assign n5960 = n4336 & n5959 ;
  assign n5961 = ~n4336 & ~n5959 ;
  assign n5962 = ~n5960 & ~n5961 ;
  assign n5963 = ~n4193 & ~n5962 ;
  assign n5964 = n4193 & n5962 ;
  assign n5965 = ~n3934 & ~n4268 ;
  assign n5966 = ~n4019 & n5965 ;
  assign n5967 = ~n4054 & ~n4129 ;
  assign n5968 = ~n4158 & n5967 ;
  assign n5969 = ~n4126 & n5968 ;
  assign n5970 = ~n4142 & n5969 ;
  assign n5971 = n4560 & n5970 ;
  assign n5972 = ~n4026 & n5971 ;
  assign n5973 = ~n4018 & n5972 ;
  assign n5974 = ~n3967 & n5973 ;
  assign n5975 = ~n4006 & n5974 ;
  assign n5976 = ~n3990 & n5975 ;
  assign n5977 = ~n4389 & n5976 ;
  assign n5978 = ~n4536 & n5977 ;
  assign n5979 = ~n4215 & n4426 ;
  assign n5980 = ~n4097 & n5979 ;
  assign n5981 = ~n4156 & n5980 ;
  assign n5982 = ~n4161 & n4768 ;
  assign n5983 = ~n3942 & n5982 ;
  assign n5984 = n4355 & n5983 ;
  assign n5985 = n4276 & n5984 ;
  assign n5986 = n4891 & n5985 ;
  assign n5987 = n5981 & n5986 ;
  assign n5988 = n4786 & n5987 ;
  assign n5989 = n4553 & n5988 ;
  assign n5990 = ~n3954 & n5989 ;
  assign n5991 = ~n3940 & n4592 ;
  assign n5992 = ~n4099 & n5991 ;
  assign n5993 = ~n4258 & n5992 ;
  assign n5994 = ~n4157 & n5993 ;
  assign n5995 = ~n3948 & n5994 ;
  assign n5996 = ~n4353 & n5995 ;
  assign n5997 = n3953 & n4608 ;
  assign n5998 = n4197 & n5997 ;
  assign n5999 = n4573 & n5998 ;
  assign n6000 = n5996 & n5999 ;
  assign n6001 = n5990 & n6000 ;
  assign n6002 = n5978 & n6001 ;
  assign n6003 = n5966 & n6002 ;
  assign n6004 = ~n4128 & n6003 ;
  assign n6005 = ~n4028 & n6004 ;
  assign n6006 = ~n3977 & n6005 ;
  assign n6007 = ~n4304 & n6006 ;
  assign n6008 = ~n4167 & n6007 ;
  assign n6009 = ~n4015 & n6008 ;
  assign n6010 = n4528 & n5953 ;
  assign n6011 = ~n5954 & ~n6010 ;
  assign n6012 = ~n6009 & ~n6011 ;
  assign n6013 = n3945 & n4594 ;
  assign n6014 = n4119 & n6013 ;
  assign n6015 = n4274 & n6014 ;
  assign n6016 = n4437 & n6015 ;
  assign n6017 = n4539 & n6016 ;
  assign n6018 = n4767 & n6017 ;
  assign n6019 = n4406 & n6018 ;
  assign n6020 = n4904 & n6019 ;
  assign n6021 = ~n4258 & n6020 ;
  assign n6022 = ~n4097 & n6021 ;
  assign n6023 = ~n4158 & n6022 ;
  assign n6024 = ~n3968 & n6023 ;
  assign n6025 = ~n4037 & n6024 ;
  assign n6026 = n5949 & ~n5951 ;
  assign n6027 = ~n5952 & ~n6026 ;
  assign n6028 = ~n6025 & ~n6027 ;
  assign n6029 = n6025 & n6027 ;
  assign n6030 = n4131 & n5983 ;
  assign n6031 = n4036 & n6030 ;
  assign n6032 = n4101 & n6031 ;
  assign n6033 = n4437 & n6032 ;
  assign n6034 = n5966 & n6033 ;
  assign n6035 = n4155 & n6034 ;
  assign n6036 = ~n4021 & n6035 ;
  assign n6037 = ~n4194 & n6036 ;
  assign n6038 = ~n4025 & n6037 ;
  assign n6039 = ~n4006 & n6038 ;
  assign n6040 = ~n4054 & n4706 ;
  assign n6041 = ~n4247 & n6040 ;
  assign n6042 = ~n3948 & n6041 ;
  assign n6043 = ~n3911 & n6042 ;
  assign n6044 = ~n4038 & n6043 ;
  assign n6045 = n4381 & n4428 ;
  assign n6046 = n6044 & n6045 ;
  assign n6047 = ~n4027 & n6046 ;
  assign n6048 = ~n4217 & n6047 ;
  assign n6049 = ~n3923 & n6048 ;
  assign n6050 = ~n4536 & n6049 ;
  assign n6051 = ~n3978 & ~n4306 ;
  assign n6052 = ~n4271 & n6051 ;
  assign n6053 = ~n4102 & ~n4113 ;
  assign n6054 = ~n4245 & n6053 ;
  assign n6055 = n4278 & n6054 ;
  assign n6056 = n6052 & n6055 ;
  assign n6057 = n3956 & n6056 ;
  assign n6058 = n4377 & n6057 ;
  assign n6059 = n4444 & n6058 ;
  assign n6060 = n6050 & n6059 ;
  assign n6061 = n6039 & n6060 ;
  assign n6062 = ~n4117 & n6061 ;
  assign n6063 = ~n4136 & n6062 ;
  assign n6064 = ~n4354 & n6063 ;
  assign n6065 = n4874 & n5946 ;
  assign n6066 = ~n5947 & ~n6065 ;
  assign n6067 = ~n6064 & ~n6066 ;
  assign n6068 = n4196 & n6052 ;
  assign n6069 = n4251 & n6068 ;
  assign n6070 = ~n3939 & n6069 ;
  assign n6071 = ~n3988 & n6070 ;
  assign n6072 = ~n3929 & n6071 ;
  assign n6073 = ~n4159 & n6072 ;
  assign n6074 = ~n4135 & n6073 ;
  assign n6075 = ~n4167 & n6074 ;
  assign n6076 = ~n4399 & n6075 ;
  assign n6077 = ~n4247 & ~n4352 ;
  assign n6078 = ~n4037 & n6077 ;
  assign n6079 = ~n3952 & n6039 ;
  assign n6080 = ~n4096 & n6079 ;
  assign n6081 = ~n4015 & n6080 ;
  assign n6082 = n5259 & n6081 ;
  assign n6083 = n6078 & n6082 ;
  assign n6084 = n4125 & n6083 ;
  assign n6085 = n5996 & n6084 ;
  assign n6086 = n6076 & n6085 ;
  assign n6087 = n4780 & n6086 ;
  assign n6088 = ~n3976 & n6087 ;
  assign n6089 = ~n4143 & n6088 ;
  assign n6090 = ~n3967 & n6089 ;
  assign n6091 = ~n4160 & n6090 ;
  assign n6092 = ~n4113 & n6091 ;
  assign n6093 = n5942 & ~n5944 ;
  assign n6094 = ~n5945 & ~n6093 ;
  assign n6095 = ~n6092 & ~n6094 ;
  assign n6096 = n6092 & n6094 ;
  assign n6097 = ~n3938 & ~n4027 ;
  assign n6098 = ~n3923 & n6097 ;
  assign n6099 = ~n3972 & n6098 ;
  assign n6100 = ~n4034 & n6099 ;
  assign n6101 = ~n4157 & n6100 ;
  assign n6102 = ~n4016 & n6101 ;
  assign n6103 = ~n3968 & n6102 ;
  assign n6104 = n3941 & n4916 ;
  assign n6105 = n4744 & n6104 ;
  assign n6106 = n4444 & n6105 ;
  assign n6107 = n4169 & n6106 ;
  assign n6108 = ~n4137 & n6107 ;
  assign n6109 = ~n4258 & n6108 ;
  assign n6110 = ~n4247 & n6109 ;
  assign n6111 = ~n4147 & n6110 ;
  assign n6112 = ~n3906 & n4723 ;
  assign n6113 = ~n4126 & n6112 ;
  assign n6114 = ~n4017 & ~n4028 ;
  assign n6115 = ~n3946 & n6114 ;
  assign n6116 = ~n4011 & n6115 ;
  assign n6117 = ~n4269 & n6116 ;
  assign n6118 = n6113 & n6117 ;
  assign n6119 = n6111 & n6118 ;
  assign n6120 = n6103 & n6119 ;
  assign n6121 = ~n4128 & n6120 ;
  assign n6122 = ~n4208 & n6121 ;
  assign n6123 = ~n3994 & n6122 ;
  assign n6124 = ~n4019 & n6123 ;
  assign n6125 = ~n4098 & n6124 ;
  assign n6126 = n4250 & n6125 ;
  assign n6127 = ~n4245 & n6126 ;
  assign n6128 = n5095 & n5940 ;
  assign n6129 = ~n5941 & ~n6128 ;
  assign n6130 = ~n6127 & ~n6129 ;
  assign n6131 = ~n4013 & n4308 ;
  assign n6132 = ~n4536 & n6131 ;
  assign n6133 = ~n4145 & n6132 ;
  assign n6134 = n4103 & n4559 ;
  assign n6135 = n4731 & n6134 ;
  assign n6136 = ~n3969 & n6135 ;
  assign n6137 = ~n3914 & n6136 ;
  assign n6138 = ~n4126 & n6137 ;
  assign n6139 = ~n4269 & n6138 ;
  assign n6140 = ~n3938 & ~n3946 ;
  assign n6141 = ~n3906 & ~n4148 ;
  assign n6142 = ~n4038 & n6141 ;
  assign n6143 = n4232 & n6142 ;
  assign n6144 = n6140 & n6143 ;
  assign n6145 = n4906 & n6144 ;
  assign n6146 = n4144 & n6145 ;
  assign n6147 = n4114 & n6146 ;
  assign n6148 = n6139 & n6147 ;
  assign n6149 = n4795 & n6148 ;
  assign n6150 = n4730 & n6149 ;
  assign n6151 = n6133 & n6150 ;
  assign n6152 = ~n3952 & n6151 ;
  assign n6153 = ~n4017 & n6152 ;
  assign n6154 = ~n4295 & n6153 ;
  assign n6155 = n5936 & ~n5938 ;
  assign n6156 = ~n5939 & ~n6155 ;
  assign n6157 = ~n6154 & ~n6156 ;
  assign n6158 = n6154 & n6156 ;
  assign n6159 = n3941 & ~n4112 ;
  assign n6160 = ~n4217 & n6159 ;
  assign n6161 = ~n4113 & n6160 ;
  assign n6162 = ~n4024 & n6161 ;
  assign n6163 = ~n4353 & n6162 ;
  assign n6164 = ~n4035 & n6163 ;
  assign n6165 = ~n4055 & ~n4249 ;
  assign n6166 = ~n4354 & n6165 ;
  assign n6167 = ~n3994 & ~n4037 ;
  assign n6168 = n6166 & n6167 ;
  assign n6169 = n4710 & n6168 ;
  assign n6170 = ~n3988 & n6169 ;
  assign n6171 = ~n4127 & n6170 ;
  assign n6172 = ~n4148 & n6171 ;
  assign n6173 = ~n4129 & n6172 ;
  assign n6174 = ~n3991 & n6173 ;
  assign n6175 = ~n4303 & n6174 ;
  assign n6176 = n4182 & n4248 ;
  assign n6177 = n6175 & n6176 ;
  assign n6178 = n4553 & n6177 ;
  assign n6179 = n6164 & n6178 ;
  assign n6180 = ~n3996 & n6179 ;
  assign n6181 = ~n4021 & n6180 ;
  assign n6182 = ~n4194 & n6181 ;
  assign n6183 = ~n3967 & n6182 ;
  assign n6184 = ~n4147 & n6183 ;
  assign n6185 = ~n4272 & n6184 ;
  assign n6186 = n5348 & n5934 ;
  assign n6187 = ~n5935 & ~n6186 ;
  assign n6188 = ~n6185 & ~n6187 ;
  assign n6189 = n4364 & n6054 ;
  assign n6190 = n4706 & n6189 ;
  assign n6191 = n4211 & n6190 ;
  assign n6192 = ~n4160 & n6191 ;
  assign n6193 = ~n3914 & n6192 ;
  assign n6194 = ~n4126 & n6193 ;
  assign n6195 = ~n4023 & n6194 ;
  assign n6196 = n4216 & n4273 ;
  assign n6197 = ~n4098 & n6196 ;
  assign n6198 = ~n3918 & n6197 ;
  assign n6199 = ~n4024 & n6198 ;
  assign n6200 = ~n4167 & n6199 ;
  assign n6201 = n4390 & n6200 ;
  assign n6202 = n6195 & n6201 ;
  assign n6203 = n4552 & n6202 ;
  assign n6204 = n4786 & n6203 ;
  assign n6205 = n3949 & n6204 ;
  assign n6206 = ~n4028 & n6205 ;
  assign n6207 = ~n4019 & n6206 ;
  assign n6208 = ~n4026 & n6207 ;
  assign n6209 = ~n4136 & n6208 ;
  assign n6210 = ~n4034 & n6209 ;
  assign n6211 = ~n4058 & n6210 ;
  assign n6212 = ~n4354 & n6211 ;
  assign n6213 = ~n4142 & n6212 ;
  assign n6214 = ~n4096 & n6213 ;
  assign n6215 = n5930 & ~n5932 ;
  assign n6216 = ~n5933 & ~n6215 ;
  assign n6217 = ~n6214 & ~n6216 ;
  assign n6218 = ~n4353 & ~n4399 ;
  assign n6219 = ~n4135 & n6218 ;
  assign n6220 = ~n3911 & n6219 ;
  assign n6221 = ~n4277 & n6220 ;
  assign n6222 = ~n4096 & ~n4249 ;
  assign n6223 = n4770 & n6222 ;
  assign n6224 = n6221 & n6223 ;
  assign n6225 = n6078 & n6224 ;
  assign n6226 = n4173 & n6225 ;
  assign n6227 = n6133 & n6226 ;
  assign n6228 = n4726 & n6227 ;
  assign n6229 = ~n4159 & n6228 ;
  assign n6230 = ~n4158 & n6229 ;
  assign n6231 = ~n4272 & n6230 ;
  assign n6232 = ~n4023 & n6231 ;
  assign n6233 = ~n4151 & ~n4304 ;
  assign n6234 = n4196 & n4606 ;
  assign n6235 = n6233 & n6234 ;
  assign n6236 = n6200 & n6235 ;
  assign n6237 = n4125 & n6236 ;
  assign n6238 = n4123 & n6237 ;
  assign n6239 = n4783 & n6238 ;
  assign n6240 = n6232 & n6239 ;
  assign n6241 = n3965 & n6240 ;
  assign n6242 = ~n4128 & n6241 ;
  assign n6243 = ~n4014 & n6242 ;
  assign n6244 = ~n4057 & n6243 ;
  assign n6245 = ~n4160 & n6244 ;
  assign n6246 = ~n4038 & n6245 ;
  assign n6247 = n5926 & ~n5928 ;
  assign n6248 = ~n5929 & ~n6247 ;
  assign n6249 = ~n6246 & ~n6248 ;
  assign n6250 = n6246 & n6248 ;
  assign n6251 = ~n3952 & n4917 ;
  assign n6252 = ~n4027 & n6251 ;
  assign n6253 = ~n4147 & n6252 ;
  assign n6254 = ~n4354 & n6253 ;
  assign n6255 = ~n3976 & ~n4112 ;
  assign n6256 = ~n4170 & n6255 ;
  assign n6257 = ~n4161 & n6256 ;
  assign n6258 = ~n3932 & n6257 ;
  assign n6259 = n6254 & n6258 ;
  assign n6260 = ~n4143 & n6259 ;
  assign n6261 = ~n4258 & n6260 ;
  assign n6262 = ~n4159 & n6261 ;
  assign n6263 = ~n4352 & n6262 ;
  assign n6264 = ~n3954 & n6263 ;
  assign n6265 = n4056 & n6222 ;
  assign n6266 = n4274 & n6265 ;
  assign n6267 = n6139 & n6266 ;
  assign n6268 = n6264 & n6267 ;
  assign n6269 = n4589 & n6268 ;
  assign n6270 = ~n4137 & n6269 ;
  assign n6271 = ~n4008 & n6270 ;
  assign n6272 = ~n3934 & n6271 ;
  assign n6273 = ~n3992 & n6272 ;
  assign n6274 = ~n3923 & n6273 ;
  assign n6275 = ~n4024 & n6274 ;
  assign n6276 = ~n4157 & n6275 ;
  assign n6277 = ~n4245 & n6276 ;
  assign n6278 = n5922 & ~n5924 ;
  assign n6279 = ~n5925 & ~n6278 ;
  assign n6280 = ~n6277 & ~n6279 ;
  assign n6281 = n6277 & n6279 ;
  assign n6282 = ~n5918 & ~n5921 ;
  assign n6283 = n5920 & ~n5921 ;
  assign n6284 = ~n6282 & ~n6283 ;
  assign n6285 = n4577 & n4896 ;
  assign n6286 = n4714 & n6285 ;
  assign n6287 = n4173 & n6286 ;
  assign n6288 = n6195 & n6287 ;
  assign n6289 = n4539 & n6288 ;
  assign n6290 = n5990 & n6289 ;
  assign n6291 = ~n4217 & n6290 ;
  assign n6292 = ~n3992 & n6291 ;
  assign n6293 = ~n4158 & n6292 ;
  assign n6294 = ~n3990 & n6293 ;
  assign n6295 = ~n4399 & n6294 ;
  assign n6296 = ~n6284 & n6295 ;
  assign n6297 = ~n6280 & ~n6296 ;
  assign n6298 = ~n6281 & n6297 ;
  assign n6299 = ~n6280 & ~n6298 ;
  assign n6300 = ~n6249 & ~n6299 ;
  assign n6301 = ~n6250 & n6300 ;
  assign n6302 = ~n6249 & ~n6301 ;
  assign n6303 = n6214 & n6216 ;
  assign n6304 = ~n6217 & ~n6303 ;
  assign n6305 = ~n6302 & n6304 ;
  assign n6306 = ~n6217 & ~n6305 ;
  assign n6307 = n6185 & n6187 ;
  assign n6308 = ~n6188 & ~n6307 ;
  assign n6309 = ~n6306 & n6308 ;
  assign n6310 = ~n6188 & ~n6309 ;
  assign n6311 = ~n6157 & ~n6310 ;
  assign n6312 = ~n6158 & n6311 ;
  assign n6313 = ~n6157 & ~n6312 ;
  assign n6314 = ~n6127 & ~n6130 ;
  assign n6315 = ~n6129 & ~n6130 ;
  assign n6316 = ~n6314 & ~n6315 ;
  assign n6317 = ~n6313 & ~n6316 ;
  assign n6318 = ~n6130 & ~n6317 ;
  assign n6319 = ~n6095 & ~n6318 ;
  assign n6320 = ~n6096 & n6319 ;
  assign n6321 = ~n6095 & ~n6320 ;
  assign n6322 = n6064 & n6066 ;
  assign n6323 = ~n6067 & ~n6322 ;
  assign n6324 = ~n6321 & n6323 ;
  assign n6325 = ~n6067 & ~n6324 ;
  assign n6326 = ~n6028 & ~n6325 ;
  assign n6327 = ~n6029 & n6326 ;
  assign n6328 = ~n6028 & ~n6327 ;
  assign n6329 = n6009 & n6011 ;
  assign n6330 = ~n6012 & ~n6329 ;
  assign n6331 = ~n6328 & n6330 ;
  assign n6332 = ~n6012 & ~n6331 ;
  assign n6333 = ~n5963 & ~n6332 ;
  assign n6334 = ~n5964 & n6333 ;
  assign n6335 = ~n5963 & ~n6334 ;
  assign n6336 = ~n4208 & n4596 ;
  assign n6337 = ~n3988 & n6336 ;
  assign n6338 = ~n4027 & n6337 ;
  assign n6339 = ~n3974 & n6338 ;
  assign n6340 = ~n4168 & n6339 ;
  assign n6341 = n4278 & n4891 ;
  assign n6342 = n6139 & n6341 ;
  assign n6343 = n5268 & n6342 ;
  assign n6344 = n6340 & n6343 ;
  assign n6345 = n4453 & n6344 ;
  assign n6346 = n3949 & n6345 ;
  assign n6347 = ~n4099 & n6346 ;
  assign n6348 = n4745 & n6347 ;
  assign n6349 = ~n4352 & n6348 ;
  assign n6350 = ~n4354 & n6349 ;
  assign n6351 = ~n4023 & n6350 ;
  assign n6352 = n6335 & n6351 ;
  assign n6353 = ~n6335 & ~n6351 ;
  assign n6354 = ~n6352 & ~n6353 ;
  assign n6355 = n4095 & ~n6354 ;
  assign n6356 = ~n4079 & n4086 ;
  assign n6357 = n4079 & ~n4086 ;
  assign n6358 = ~n6356 & ~n6357 ;
  assign n6359 = ~n4082 & n4094 ;
  assign n6360 = n6358 & n6359 ;
  assign n6361 = n6328 & ~n6330 ;
  assign n6362 = ~n6331 & ~n6361 ;
  assign n6363 = n6360 & n6362 ;
  assign n6364 = ~n6332 & ~n6334 ;
  assign n6365 = ~n5964 & n6335 ;
  assign n6366 = ~n6364 & ~n6365 ;
  assign n6367 = n4094 & ~n6358 ;
  assign n6368 = ~n6366 & n6367 ;
  assign n6369 = ~n6363 & ~n6368 ;
  assign n6370 = ~n6355 & n6369 ;
  assign n6371 = ~n4082 & ~n4094 ;
  assign n6372 = n6362 & ~n6366 ;
  assign n6373 = ~n6325 & ~n6327 ;
  assign n6374 = ~n6029 & n6328 ;
  assign n6375 = ~n6373 & ~n6374 ;
  assign n6376 = n6362 & ~n6375 ;
  assign n6377 = n6321 & ~n6323 ;
  assign n6378 = ~n6324 & ~n6377 ;
  assign n6379 = ~n6375 & n6378 ;
  assign n6380 = ~n6318 & ~n6320 ;
  assign n6381 = ~n6096 & n6321 ;
  assign n6382 = ~n6380 & ~n6381 ;
  assign n6383 = n6378 & ~n6382 ;
  assign n6384 = ~n6313 & ~n6317 ;
  assign n6385 = ~n6316 & ~n6317 ;
  assign n6386 = ~n6384 & ~n6385 ;
  assign n6387 = ~n6382 & ~n6386 ;
  assign n6388 = ~n6310 & ~n6312 ;
  assign n6389 = ~n6158 & n6313 ;
  assign n6390 = ~n6388 & ~n6389 ;
  assign n6391 = ~n6386 & ~n6390 ;
  assign n6392 = n6306 & ~n6308 ;
  assign n6393 = ~n6309 & ~n6392 ;
  assign n6394 = ~n6390 & n6393 ;
  assign n6395 = n6302 & ~n6304 ;
  assign n6396 = ~n6305 & ~n6395 ;
  assign n6397 = n6393 & n6396 ;
  assign n6398 = ~n6299 & ~n6301 ;
  assign n6399 = ~n6250 & n6302 ;
  assign n6400 = ~n6398 & ~n6399 ;
  assign n6401 = n6396 & ~n6400 ;
  assign n6402 = ~n6296 & ~n6298 ;
  assign n6403 = ~n6281 & n6299 ;
  assign n6404 = ~n6402 & ~n6403 ;
  assign n6405 = ~n6400 & ~n6404 ;
  assign n6406 = n6284 & ~n6295 ;
  assign n6407 = ~n6296 & ~n6406 ;
  assign n6408 = ~n6404 & ~n6407 ;
  assign n6409 = n6400 & n6408 ;
  assign n6410 = ~n6405 & ~n6409 ;
  assign n6411 = ~n6396 & n6400 ;
  assign n6412 = ~n6410 & ~n6411 ;
  assign n6413 = ~n6401 & n6412 ;
  assign n6414 = ~n6401 & ~n6413 ;
  assign n6415 = ~n6393 & ~n6396 ;
  assign n6416 = ~n6414 & ~n6415 ;
  assign n6417 = ~n6397 & n6416 ;
  assign n6418 = ~n6397 & ~n6417 ;
  assign n6419 = n6390 & ~n6393 ;
  assign n6420 = ~n6394 & ~n6419 ;
  assign n6421 = ~n6418 & n6420 ;
  assign n6422 = ~n6394 & ~n6421 ;
  assign n6423 = n6386 & n6390 ;
  assign n6424 = ~n6391 & ~n6423 ;
  assign n6425 = ~n6422 & n6424 ;
  assign n6426 = ~n6391 & ~n6425 ;
  assign n6427 = n6382 & n6386 ;
  assign n6428 = ~n6387 & ~n6427 ;
  assign n6429 = ~n6426 & n6428 ;
  assign n6430 = ~n6387 & ~n6429 ;
  assign n6431 = ~n6378 & n6382 ;
  assign n6432 = ~n6383 & ~n6431 ;
  assign n6433 = ~n6430 & n6432 ;
  assign n6434 = ~n6383 & ~n6433 ;
  assign n6435 = n6375 & ~n6378 ;
  assign n6436 = ~n6379 & ~n6435 ;
  assign n6437 = ~n6434 & n6436 ;
  assign n6438 = ~n6379 & ~n6437 ;
  assign n6439 = ~n6362 & n6375 ;
  assign n6440 = ~n6376 & ~n6439 ;
  assign n6441 = ~n6438 & n6440 ;
  assign n6442 = ~n6376 & ~n6441 ;
  assign n6443 = ~n6362 & n6366 ;
  assign n6444 = ~n6372 & ~n6443 ;
  assign n6445 = ~n6442 & n6444 ;
  assign n6446 = ~n6372 & ~n6445 ;
  assign n6447 = ~n6354 & ~n6366 ;
  assign n6448 = n6354 & n6366 ;
  assign n6449 = ~n6447 & ~n6448 ;
  assign n6450 = ~n6446 & n6449 ;
  assign n6451 = n6446 & ~n6449 ;
  assign n6452 = ~n6450 & ~n6451 ;
  assign n6453 = n6371 & n6452 ;
  assign n6454 = n6370 & ~n6453 ;
  assign n6455 = ~n4075 & ~n6454 ;
  assign n6456 = n4075 & n6454 ;
  assign n6457 = ~n6455 & ~n6456 ;
  assign n6458 = n4469 & ~n4477 ;
  assign n6459 = ~n4469 & n4477 ;
  assign n6460 = ~n6458 & ~n6459 ;
  assign n6461 = ~n6407 & ~n6460 ;
  assign n6462 = ~n4325 & ~n6461 ;
  assign n6463 = n4329 & ~n4477 ;
  assign n6464 = ~n4329 & n4477 ;
  assign n6465 = ~n6463 & ~n6464 ;
  assign n6466 = n6460 & ~n6465 ;
  assign n6467 = ~n6407 & n6466 ;
  assign n6468 = n4332 & ~n6460 ;
  assign n6469 = ~n6404 & n6468 ;
  assign n6470 = ~n6467 & ~n6469 ;
  assign n6471 = n6404 & ~n6407 ;
  assign n6472 = ~n6404 & n6407 ;
  assign n6473 = ~n6471 & ~n6472 ;
  assign n6474 = ~n4332 & ~n6460 ;
  assign n6475 = ~n6473 & n6474 ;
  assign n6476 = n6470 & ~n6475 ;
  assign n6477 = ~n4325 & ~n6476 ;
  assign n6478 = ~n4325 & ~n6477 ;
  assign n6479 = ~n6476 & ~n6477 ;
  assign n6480 = ~n6478 & ~n6479 ;
  assign n6481 = n6462 & ~n6480 ;
  assign n6482 = ~n6462 & n6480 ;
  assign n6483 = ~n6481 & ~n6482 ;
  assign n6484 = n4632 & ~n4821 ;
  assign n6485 = ~n4632 & n4821 ;
  assign n6486 = ~n6484 & ~n6485 ;
  assign n6487 = n4469 & ~n4640 ;
  assign n6488 = ~n4469 & n4640 ;
  assign n6489 = ~n6487 & ~n6488 ;
  assign n6490 = ~n6486 & ~n6489 ;
  assign n6491 = n4632 & ~n4640 ;
  assign n6492 = ~n4632 & n4640 ;
  assign n6493 = ~n6491 & ~n6492 ;
  assign n6494 = n6486 & ~n6489 ;
  assign n6495 = n6493 & n6494 ;
  assign n6496 = ~n6400 & n6495 ;
  assign n6497 = n6486 & ~n6493 ;
  assign n6498 = n6396 & n6497 ;
  assign n6499 = ~n6486 & n6489 ;
  assign n6500 = n6393 & n6499 ;
  assign n6501 = ~n6498 & ~n6500 ;
  assign n6502 = ~n6496 & n6501 ;
  assign n6503 = ~n6490 & n6502 ;
  assign n6504 = ~n6414 & ~n6417 ;
  assign n6505 = ~n6415 & n6418 ;
  assign n6506 = ~n6504 & ~n6505 ;
  assign n6507 = n6502 & n6506 ;
  assign n6508 = ~n6503 & ~n6507 ;
  assign n6509 = n4469 & ~n6508 ;
  assign n6510 = ~n4469 & n6508 ;
  assign n6511 = ~n6509 & ~n6510 ;
  assign n6512 = n6483 & n6511 ;
  assign n6513 = ~n6407 & ~n6486 ;
  assign n6514 = ~n4469 & ~n6513 ;
  assign n6515 = ~n6407 & n6497 ;
  assign n6516 = ~n6404 & n6499 ;
  assign n6517 = ~n6515 & ~n6516 ;
  assign n6518 = ~n6473 & n6490 ;
  assign n6519 = n6517 & ~n6518 ;
  assign n6520 = ~n4469 & ~n6519 ;
  assign n6521 = n4469 & n6519 ;
  assign n6522 = ~n6520 & ~n6521 ;
  assign n6523 = n6514 & n6522 ;
  assign n6524 = ~n6400 & n6499 ;
  assign n6525 = ~n6407 & n6495 ;
  assign n6526 = ~n6404 & n6497 ;
  assign n6527 = ~n6525 & ~n6526 ;
  assign n6528 = ~n6524 & n6527 ;
  assign n6529 = ~n6490 & n6528 ;
  assign n6530 = n6400 & ~n6472 ;
  assign n6531 = ~n6400 & n6472 ;
  assign n6532 = ~n6530 & ~n6531 ;
  assign n6533 = n6528 & ~n6532 ;
  assign n6534 = ~n6529 & ~n6533 ;
  assign n6535 = n4469 & ~n6534 ;
  assign n6536 = ~n4469 & n6534 ;
  assign n6537 = ~n6535 & ~n6536 ;
  assign n6538 = n6523 & n6537 ;
  assign n6539 = n6461 & n6538 ;
  assign n6540 = n6538 & ~n6539 ;
  assign n6541 = n6461 & ~n6539 ;
  assign n6542 = ~n6540 & ~n6541 ;
  assign n6543 = ~n6400 & n6497 ;
  assign n6544 = n6396 & n6499 ;
  assign n6545 = ~n6404 & n6495 ;
  assign n6546 = ~n6544 & ~n6545 ;
  assign n6547 = ~n6543 & n6546 ;
  assign n6548 = ~n6410 & ~n6413 ;
  assign n6549 = ~n6411 & n6414 ;
  assign n6550 = ~n6548 & ~n6549 ;
  assign n6551 = n6490 & ~n6550 ;
  assign n6552 = n6547 & ~n6551 ;
  assign n6553 = ~n4469 & ~n6552 ;
  assign n6554 = n4469 & n6552 ;
  assign n6555 = ~n6553 & ~n6554 ;
  assign n6556 = ~n6542 & n6555 ;
  assign n6557 = ~n6539 & ~n6556 ;
  assign n6558 = ~n6483 & ~n6511 ;
  assign n6559 = ~n6512 & ~n6558 ;
  assign n6560 = ~n6557 & n6559 ;
  assign n6561 = ~n6512 & ~n6560 ;
  assign n6562 = ~n6390 & n6499 ;
  assign n6563 = n6396 & n6495 ;
  assign n6564 = n6393 & n6497 ;
  assign n6565 = ~n6563 & ~n6564 ;
  assign n6566 = ~n6562 & n6565 ;
  assign n6567 = n6418 & ~n6420 ;
  assign n6568 = ~n6421 & ~n6567 ;
  assign n6569 = n6490 & n6568 ;
  assign n6570 = n6566 & ~n6569 ;
  assign n6571 = ~n4469 & ~n6570 ;
  assign n6572 = n4469 & n6570 ;
  assign n6573 = ~n6571 & ~n6572 ;
  assign n6574 = ~n6400 & n6468 ;
  assign n6575 = ~n4332 & n6460 ;
  assign n6576 = n6465 & n6575 ;
  assign n6577 = ~n6407 & n6576 ;
  assign n6578 = ~n6404 & n6466 ;
  assign n6579 = ~n6577 & ~n6578 ;
  assign n6580 = ~n6574 & n6579 ;
  assign n6581 = ~n6474 & n6580 ;
  assign n6582 = ~n6532 & n6580 ;
  assign n6583 = ~n6581 & ~n6582 ;
  assign n6584 = n4325 & ~n6583 ;
  assign n6585 = ~n4325 & n6583 ;
  assign n6586 = ~n6584 & ~n6585 ;
  assign n6587 = n6481 & n6586 ;
  assign n6588 = ~n6481 & ~n6586 ;
  assign n6589 = ~n6587 & ~n6588 ;
  assign n6590 = n6573 & n6589 ;
  assign n6591 = ~n6573 & ~n6589 ;
  assign n6592 = ~n6590 & ~n6591 ;
  assign n6593 = n6561 & ~n6592 ;
  assign n6594 = ~n6561 & n6592 ;
  assign n6595 = ~n6593 & ~n6594 ;
  assign n6596 = n4813 & ~n4821 ;
  assign n6597 = ~n4813 & n4821 ;
  assign n6598 = ~n6596 & ~n6597 ;
  assign n6599 = n4075 & ~n4983 ;
  assign n6600 = ~n4075 & n4983 ;
  assign n6601 = ~n6599 & ~n6600 ;
  assign n6602 = n6598 & ~n6601 ;
  assign n6603 = n6378 & n6602 ;
  assign n6604 = n4813 & ~n4983 ;
  assign n6605 = ~n4813 & n4983 ;
  assign n6606 = ~n6604 & ~n6605 ;
  assign n6607 = ~n6598 & n6601 ;
  assign n6608 = n6606 & n6607 ;
  assign n6609 = ~n6386 & n6608 ;
  assign n6610 = n6601 & ~n6606 ;
  assign n6611 = ~n6382 & n6610 ;
  assign n6612 = ~n6609 & ~n6611 ;
  assign n6613 = ~n6603 & n6612 ;
  assign n6614 = n6430 & ~n6432 ;
  assign n6615 = ~n6433 & ~n6614 ;
  assign n6616 = n6613 & ~n6615 ;
  assign n6617 = ~n6598 & ~n6601 ;
  assign n6618 = n6613 & ~n6617 ;
  assign n6619 = ~n6616 & ~n6618 ;
  assign n6620 = n4821 & ~n6619 ;
  assign n6621 = ~n4821 & n6619 ;
  assign n6622 = ~n6620 & ~n6621 ;
  assign n6623 = n6595 & n6622 ;
  assign n6624 = ~n6382 & n6602 ;
  assign n6625 = ~n6390 & n6608 ;
  assign n6626 = ~n6386 & n6610 ;
  assign n6627 = ~n6625 & ~n6626 ;
  assign n6628 = ~n6624 & n6627 ;
  assign n6629 = n6426 & ~n6428 ;
  assign n6630 = ~n6429 & ~n6629 ;
  assign n6631 = n6617 & n6630 ;
  assign n6632 = n6628 & ~n6631 ;
  assign n6633 = ~n4821 & ~n6632 ;
  assign n6634 = ~n6632 & ~n6633 ;
  assign n6635 = ~n4821 & ~n6633 ;
  assign n6636 = ~n6634 & ~n6635 ;
  assign n6637 = n6557 & ~n6559 ;
  assign n6638 = ~n6560 & ~n6637 ;
  assign n6639 = ~n6636 & n6638 ;
  assign n6640 = ~n6542 & ~n6556 ;
  assign n6641 = n6555 & ~n6556 ;
  assign n6642 = ~n6640 & ~n6641 ;
  assign n6643 = ~n6386 & n6602 ;
  assign n6644 = n6393 & n6608 ;
  assign n6645 = ~n6390 & n6610 ;
  assign n6646 = ~n6644 & ~n6645 ;
  assign n6647 = ~n6643 & n6646 ;
  assign n6648 = n6422 & ~n6424 ;
  assign n6649 = ~n6425 & ~n6648 ;
  assign n6650 = n6647 & ~n6649 ;
  assign n6651 = ~n6617 & n6647 ;
  assign n6652 = ~n6650 & ~n6651 ;
  assign n6653 = n4821 & ~n6652 ;
  assign n6654 = ~n4821 & n6652 ;
  assign n6655 = ~n6653 & ~n6654 ;
  assign n6656 = ~n6642 & n6655 ;
  assign n6657 = ~n6390 & n6602 ;
  assign n6658 = n6396 & n6608 ;
  assign n6659 = n6393 & n6610 ;
  assign n6660 = ~n6658 & ~n6659 ;
  assign n6661 = ~n6657 & n6660 ;
  assign n6662 = n6568 & n6617 ;
  assign n6663 = n6661 & ~n6662 ;
  assign n6664 = ~n4821 & ~n6663 ;
  assign n6665 = ~n6663 & ~n6664 ;
  assign n6666 = ~n4821 & ~n6664 ;
  assign n6667 = ~n6665 & ~n6666 ;
  assign n6668 = ~n6523 & ~n6537 ;
  assign n6669 = ~n6538 & ~n6668 ;
  assign n6670 = ~n6667 & n6669 ;
  assign n6671 = ~n6514 & ~n6522 ;
  assign n6672 = ~n6523 & ~n6671 ;
  assign n6673 = ~n6400 & n6608 ;
  assign n6674 = n6396 & n6610 ;
  assign n6675 = n6393 & n6602 ;
  assign n6676 = ~n6674 & ~n6675 ;
  assign n6677 = ~n6673 & n6676 ;
  assign n6678 = ~n6617 & n6677 ;
  assign n6679 = n6506 & n6677 ;
  assign n6680 = ~n6678 & ~n6679 ;
  assign n6681 = n4821 & ~n6680 ;
  assign n6682 = ~n4821 & n6680 ;
  assign n6683 = ~n6681 & ~n6682 ;
  assign n6684 = n6672 & n6683 ;
  assign n6685 = ~n6407 & n6610 ;
  assign n6686 = ~n6404 & n6602 ;
  assign n6687 = ~n6685 & ~n6686 ;
  assign n6688 = ~n6473 & n6617 ;
  assign n6689 = n6687 & ~n6688 ;
  assign n6690 = ~n4821 & ~n6689 ;
  assign n6691 = ~n4821 & ~n6690 ;
  assign n6692 = ~n6689 & ~n6690 ;
  assign n6693 = ~n6691 & ~n6692 ;
  assign n6694 = ~n6407 & ~n6601 ;
  assign n6695 = ~n4821 & ~n6694 ;
  assign n6696 = ~n6693 & n6695 ;
  assign n6697 = ~n6400 & n6602 ;
  assign n6698 = ~n6407 & n6608 ;
  assign n6699 = ~n6404 & n6610 ;
  assign n6700 = ~n6698 & ~n6699 ;
  assign n6701 = ~n6697 & n6700 ;
  assign n6702 = ~n6532 & n6701 ;
  assign n6703 = ~n6617 & n6701 ;
  assign n6704 = ~n6702 & ~n6703 ;
  assign n6705 = n4821 & ~n6704 ;
  assign n6706 = ~n4821 & n6704 ;
  assign n6707 = ~n6705 & ~n6706 ;
  assign n6708 = n6696 & n6707 ;
  assign n6709 = n6513 & n6708 ;
  assign n6710 = n6708 & ~n6709 ;
  assign n6711 = n6513 & ~n6709 ;
  assign n6712 = ~n6710 & ~n6711 ;
  assign n6713 = ~n6400 & n6610 ;
  assign n6714 = n6396 & n6602 ;
  assign n6715 = ~n6404 & n6608 ;
  assign n6716 = ~n6714 & ~n6715 ;
  assign n6717 = ~n6713 & n6716 ;
  assign n6718 = ~n6550 & n6617 ;
  assign n6719 = n6717 & ~n6718 ;
  assign n6720 = ~n4821 & ~n6719 ;
  assign n6721 = ~n4821 & ~n6720 ;
  assign n6722 = ~n6719 & ~n6720 ;
  assign n6723 = ~n6721 & ~n6722 ;
  assign n6724 = ~n6712 & ~n6723 ;
  assign n6725 = ~n6709 & ~n6724 ;
  assign n6726 = ~n6672 & ~n6683 ;
  assign n6727 = ~n6684 & ~n6726 ;
  assign n6728 = ~n6725 & n6727 ;
  assign n6729 = ~n6684 & ~n6728 ;
  assign n6730 = ~n6667 & ~n6670 ;
  assign n6731 = n6669 & ~n6670 ;
  assign n6732 = ~n6730 & ~n6731 ;
  assign n6733 = ~n6729 & ~n6732 ;
  assign n6734 = ~n6670 & ~n6733 ;
  assign n6735 = ~n6642 & ~n6656 ;
  assign n6736 = n6655 & ~n6656 ;
  assign n6737 = ~n6735 & ~n6736 ;
  assign n6738 = ~n6734 & ~n6737 ;
  assign n6739 = ~n6656 & ~n6738 ;
  assign n6740 = ~n6636 & ~n6639 ;
  assign n6741 = n6638 & ~n6639 ;
  assign n6742 = ~n6740 & ~n6741 ;
  assign n6743 = ~n6739 & ~n6742 ;
  assign n6744 = ~n6639 & ~n6743 ;
  assign n6745 = n6595 & ~n6623 ;
  assign n6746 = n6622 & ~n6623 ;
  assign n6747 = ~n6745 & ~n6746 ;
  assign n6748 = ~n6744 & ~n6747 ;
  assign n6749 = ~n6623 & ~n6748 ;
  assign n6750 = ~n6386 & n6499 ;
  assign n6751 = n6393 & n6495 ;
  assign n6752 = ~n6390 & n6497 ;
  assign n6753 = ~n6751 & ~n6752 ;
  assign n6754 = ~n6750 & n6753 ;
  assign n6755 = n6490 & n6649 ;
  assign n6756 = n6754 & ~n6755 ;
  assign n6757 = ~n4469 & ~n6756 ;
  assign n6758 = n4469 & n6756 ;
  assign n6759 = ~n6757 & ~n6758 ;
  assign n6760 = ~n6400 & n6466 ;
  assign n6761 = n6396 & n6468 ;
  assign n6762 = ~n6404 & n6576 ;
  assign n6763 = ~n6761 & ~n6762 ;
  assign n6764 = ~n6760 & n6763 ;
  assign n6765 = n6474 & ~n6550 ;
  assign n6766 = n6764 & ~n6765 ;
  assign n6767 = ~n4325 & ~n6766 ;
  assign n6768 = ~n6766 & ~n6767 ;
  assign n6769 = ~n4325 & ~n6767 ;
  assign n6770 = ~n6768 & ~n6769 ;
  assign n6771 = ~n4325 & ~n6407 ;
  assign n6772 = ~n6587 & ~n6771 ;
  assign n6773 = n6587 & n6771 ;
  assign n6774 = ~n6770 & ~n6773 ;
  assign n6775 = ~n6772 & n6774 ;
  assign n6776 = ~n6770 & ~n6775 ;
  assign n6777 = ~n6773 & ~n6775 ;
  assign n6778 = ~n6772 & n6777 ;
  assign n6779 = ~n6776 & ~n6778 ;
  assign n6780 = n6759 & ~n6779 ;
  assign n6781 = n6759 & ~n6780 ;
  assign n6782 = ~n6779 & ~n6780 ;
  assign n6783 = ~n6781 & ~n6782 ;
  assign n6784 = ~n6590 & ~n6594 ;
  assign n6785 = n6783 & n6784 ;
  assign n6786 = ~n6783 & ~n6784 ;
  assign n6787 = ~n6785 & ~n6786 ;
  assign n6788 = n6434 & ~n6436 ;
  assign n6789 = ~n6437 & ~n6788 ;
  assign n6790 = ~n6375 & n6602 ;
  assign n6791 = ~n6382 & n6608 ;
  assign n6792 = n6378 & n6610 ;
  assign n6793 = ~n6791 & ~n6792 ;
  assign n6794 = ~n6790 & n6793 ;
  assign n6795 = ~n6789 & n6794 ;
  assign n6796 = ~n6617 & n6794 ;
  assign n6797 = ~n6795 & ~n6796 ;
  assign n6798 = n4821 & ~n6797 ;
  assign n6799 = ~n4821 & n6797 ;
  assign n6800 = ~n6798 & ~n6799 ;
  assign n6801 = n6787 & n6800 ;
  assign n6802 = n6787 & ~n6801 ;
  assign n6803 = n6800 & ~n6801 ;
  assign n6804 = ~n6802 & ~n6803 ;
  assign n6805 = ~n6749 & ~n6804 ;
  assign n6806 = ~n6749 & ~n6805 ;
  assign n6807 = ~n6804 & ~n6805 ;
  assign n6808 = ~n6806 & ~n6807 ;
  assign n6809 = n6457 & ~n6808 ;
  assign n6810 = n6457 & ~n6809 ;
  assign n6811 = ~n6808 & ~n6809 ;
  assign n6812 = ~n6810 & ~n6811 ;
  assign n6813 = ~n6744 & ~n6748 ;
  assign n6814 = ~n6747 & ~n6748 ;
  assign n6815 = ~n6813 & ~n6814 ;
  assign n6816 = n4095 & ~n6366 ;
  assign n6817 = n6360 & ~n6375 ;
  assign n6818 = n6362 & n6367 ;
  assign n6819 = ~n6817 & ~n6818 ;
  assign n6820 = ~n6816 & n6819 ;
  assign n6821 = n6442 & ~n6444 ;
  assign n6822 = ~n6445 & ~n6821 ;
  assign n6823 = n6371 & n6822 ;
  assign n6824 = n6820 & ~n6823 ;
  assign n6825 = ~n4075 & ~n6824 ;
  assign n6826 = n4075 & n6824 ;
  assign n6827 = ~n6825 & ~n6826 ;
  assign n6828 = ~n6815 & n6827 ;
  assign n6829 = n6827 & ~n6828 ;
  assign n6830 = ~n6815 & ~n6828 ;
  assign n6831 = ~n6829 & ~n6830 ;
  assign n6832 = ~n6739 & n6742 ;
  assign n6833 = n6739 & ~n6742 ;
  assign n6834 = ~n6832 & ~n6833 ;
  assign n6835 = n4095 & n6362 ;
  assign n6836 = n6360 & n6378 ;
  assign n6837 = n6367 & ~n6375 ;
  assign n6838 = ~n6836 & ~n6837 ;
  assign n6839 = ~n6835 & n6838 ;
  assign n6840 = ~n6371 & n6839 ;
  assign n6841 = n6438 & ~n6440 ;
  assign n6842 = ~n6441 & ~n6841 ;
  assign n6843 = n6839 & ~n6842 ;
  assign n6844 = ~n6840 & ~n6843 ;
  assign n6845 = n4075 & ~n6844 ;
  assign n6846 = ~n4075 & n6844 ;
  assign n6847 = ~n6845 & ~n6846 ;
  assign n6848 = ~n6834 & n6847 ;
  assign n6849 = ~n6734 & ~n6738 ;
  assign n6850 = ~n6737 & ~n6738 ;
  assign n6851 = ~n6849 & ~n6850 ;
  assign n6852 = n4095 & ~n6375 ;
  assign n6853 = n6360 & ~n6382 ;
  assign n6854 = n6367 & n6378 ;
  assign n6855 = ~n6853 & ~n6854 ;
  assign n6856 = ~n6852 & n6855 ;
  assign n6857 = ~n6371 & n6856 ;
  assign n6858 = ~n6789 & n6856 ;
  assign n6859 = ~n6857 & ~n6858 ;
  assign n6860 = n4075 & ~n6859 ;
  assign n6861 = ~n4075 & n6859 ;
  assign n6862 = ~n6860 & ~n6861 ;
  assign n6863 = ~n6851 & n6862 ;
  assign n6864 = ~n6729 & n6732 ;
  assign n6865 = n6729 & ~n6732 ;
  assign n6866 = ~n6864 & ~n6865 ;
  assign n6867 = n4095 & n6378 ;
  assign n6868 = n6360 & ~n6386 ;
  assign n6869 = n6367 & ~n6382 ;
  assign n6870 = ~n6868 & ~n6869 ;
  assign n6871 = ~n6867 & n6870 ;
  assign n6872 = ~n6371 & n6871 ;
  assign n6873 = ~n6615 & n6871 ;
  assign n6874 = ~n6872 & ~n6873 ;
  assign n6875 = n4075 & ~n6874 ;
  assign n6876 = ~n4075 & n6874 ;
  assign n6877 = ~n6875 & ~n6876 ;
  assign n6878 = ~n6866 & n6877 ;
  assign n6879 = n4095 & ~n6382 ;
  assign n6880 = n6360 & ~n6390 ;
  assign n6881 = n6367 & ~n6386 ;
  assign n6882 = ~n6880 & ~n6881 ;
  assign n6883 = ~n6879 & n6882 ;
  assign n6884 = n6371 & n6630 ;
  assign n6885 = n6883 & ~n6884 ;
  assign n6886 = ~n4075 & ~n6885 ;
  assign n6887 = n4075 & n6885 ;
  assign n6888 = ~n6886 & ~n6887 ;
  assign n6889 = n6725 & ~n6727 ;
  assign n6890 = ~n6728 & ~n6889 ;
  assign n6891 = n6888 & n6890 ;
  assign n6892 = ~n6712 & ~n6724 ;
  assign n6893 = ~n6723 & ~n6724 ;
  assign n6894 = ~n6892 & ~n6893 ;
  assign n6895 = n4095 & ~n6386 ;
  assign n6896 = n6360 & n6393 ;
  assign n6897 = n6367 & ~n6390 ;
  assign n6898 = ~n6896 & ~n6897 ;
  assign n6899 = ~n6895 & n6898 ;
  assign n6900 = ~n6371 & n6899 ;
  assign n6901 = ~n6649 & n6899 ;
  assign n6902 = ~n6900 & ~n6901 ;
  assign n6903 = n4075 & ~n6902 ;
  assign n6904 = ~n4075 & n6902 ;
  assign n6905 = ~n6903 & ~n6904 ;
  assign n6906 = ~n6894 & n6905 ;
  assign n6907 = n4095 & ~n6390 ;
  assign n6908 = n6360 & n6396 ;
  assign n6909 = n6367 & n6393 ;
  assign n6910 = ~n6908 & ~n6909 ;
  assign n6911 = ~n6907 & n6910 ;
  assign n6912 = n6371 & n6568 ;
  assign n6913 = n6911 & ~n6912 ;
  assign n6914 = ~n4075 & ~n6913 ;
  assign n6915 = n4075 & n6913 ;
  assign n6916 = ~n6914 & ~n6915 ;
  assign n6917 = ~n6696 & ~n6707 ;
  assign n6918 = ~n6708 & ~n6917 ;
  assign n6919 = n6916 & n6918 ;
  assign n6920 = n6693 & ~n6695 ;
  assign n6921 = ~n6696 & ~n6920 ;
  assign n6922 = n6360 & ~n6400 ;
  assign n6923 = n6367 & n6396 ;
  assign n6924 = n4095 & n6393 ;
  assign n6925 = ~n6923 & ~n6924 ;
  assign n6926 = ~n6922 & n6925 ;
  assign n6927 = ~n6371 & n6926 ;
  assign n6928 = n6506 & n6926 ;
  assign n6929 = ~n6927 & ~n6928 ;
  assign n6930 = n4075 & ~n6929 ;
  assign n6931 = ~n4075 & n6929 ;
  assign n6932 = ~n6930 & ~n6931 ;
  assign n6933 = n6921 & n6932 ;
  assign n6934 = ~n4094 & ~n6407 ;
  assign n6935 = ~n4075 & ~n6934 ;
  assign n6936 = n6367 & ~n6407 ;
  assign n6937 = n4095 & ~n6404 ;
  assign n6938 = ~n6936 & ~n6937 ;
  assign n6939 = n6371 & ~n6473 ;
  assign n6940 = n6938 & ~n6939 ;
  assign n6941 = ~n4075 & ~n6940 ;
  assign n6942 = n4075 & n6940 ;
  assign n6943 = ~n6941 & ~n6942 ;
  assign n6944 = n6935 & n6943 ;
  assign n6945 = n4095 & ~n6400 ;
  assign n6946 = n6360 & ~n6407 ;
  assign n6947 = n6367 & ~n6404 ;
  assign n6948 = ~n6946 & ~n6947 ;
  assign n6949 = ~n6945 & n6948 ;
  assign n6950 = ~n6371 & n6949 ;
  assign n6951 = ~n6532 & n6949 ;
  assign n6952 = ~n6950 & ~n6951 ;
  assign n6953 = n4075 & ~n6952 ;
  assign n6954 = ~n4075 & n6952 ;
  assign n6955 = ~n6953 & ~n6954 ;
  assign n6956 = n6944 & n6955 ;
  assign n6957 = n6694 & n6956 ;
  assign n6958 = n6956 & ~n6957 ;
  assign n6959 = n6694 & ~n6957 ;
  assign n6960 = ~n6958 & ~n6959 ;
  assign n6961 = n6367 & ~n6400 ;
  assign n6962 = n4095 & n6396 ;
  assign n6963 = n6360 & ~n6404 ;
  assign n6964 = ~n6962 & ~n6963 ;
  assign n6965 = ~n6961 & n6964 ;
  assign n6966 = n6371 & ~n6550 ;
  assign n6967 = n6965 & ~n6966 ;
  assign n6968 = ~n4075 & ~n6967 ;
  assign n6969 = n4075 & n6967 ;
  assign n6970 = ~n6968 & ~n6969 ;
  assign n6971 = ~n6960 & n6970 ;
  assign n6972 = ~n6957 & ~n6971 ;
  assign n6973 = ~n6921 & ~n6932 ;
  assign n6974 = ~n6933 & ~n6973 ;
  assign n6975 = ~n6972 & n6974 ;
  assign n6976 = ~n6933 & ~n6975 ;
  assign n6977 = ~n6916 & ~n6918 ;
  assign n6978 = ~n6919 & ~n6977 ;
  assign n6979 = ~n6976 & n6978 ;
  assign n6980 = ~n6919 & ~n6979 ;
  assign n6981 = ~n6894 & ~n6906 ;
  assign n6982 = n6905 & ~n6906 ;
  assign n6983 = ~n6981 & ~n6982 ;
  assign n6984 = ~n6980 & ~n6983 ;
  assign n6985 = ~n6906 & ~n6984 ;
  assign n6986 = ~n6888 & ~n6890 ;
  assign n6987 = ~n6891 & ~n6986 ;
  assign n6988 = ~n6985 & n6987 ;
  assign n6989 = ~n6891 & ~n6988 ;
  assign n6990 = ~n6866 & ~n6878 ;
  assign n6991 = n6877 & ~n6878 ;
  assign n6992 = ~n6990 & ~n6991 ;
  assign n6993 = ~n6989 & ~n6992 ;
  assign n6994 = ~n6878 & ~n6993 ;
  assign n6995 = ~n6851 & ~n6863 ;
  assign n6996 = n6862 & ~n6863 ;
  assign n6997 = ~n6995 & ~n6996 ;
  assign n6998 = ~n6994 & ~n6997 ;
  assign n6999 = ~n6863 & ~n6998 ;
  assign n7000 = n6834 & ~n6847 ;
  assign n7001 = ~n6848 & ~n7000 ;
  assign n7002 = ~n6999 & n7001 ;
  assign n7003 = ~n6848 & ~n7002 ;
  assign n7004 = ~n6831 & ~n7003 ;
  assign n7005 = ~n6828 & ~n7004 ;
  assign n7006 = n6812 & n7005 ;
  assign n7007 = ~n6812 & ~n7005 ;
  assign n7008 = ~n7006 & ~n7007 ;
  assign n7009 = ~x0 & x22 ;
  assign n7010 = ~x1 & ~n7009 ;
  assign n7011 = x1 & n7009 ;
  assign n7012 = ~n7010 & ~n7011 ;
  assign n7013 = ~n4091 & n7012 ;
  assign n7014 = n4091 & ~n7012 ;
  assign n7015 = ~n7013 & ~n7014 ;
  assign n7016 = ~x0 & ~n7015 ;
  assign n7017 = ~x0 & n7015 ;
  assign n7018 = ~n4124 & n4609 ;
  assign n7019 = n4285 & n7018 ;
  assign n7020 = n4231 & n7019 ;
  assign n7021 = n6044 & n7020 ;
  assign n7022 = n6133 & n7021 ;
  assign n7023 = n6218 & n7022 ;
  assign n7024 = n4776 & n7023 ;
  assign n7025 = ~n4304 & n7024 ;
  assign n7026 = ~n4097 & n7025 ;
  assign n7027 = ~n4012 & n7026 ;
  assign n7028 = ~n4058 & n7027 ;
  assign n7029 = ~n4037 & n7028 ;
  assign n7030 = ~n4100 & n4608 ;
  assign n7031 = ~n4126 & n7030 ;
  assign n7032 = n4000 & n7031 ;
  assign n7033 = n5966 & n7032 ;
  assign n7034 = ~n4215 & n7033 ;
  assign n7035 = ~n4026 & n7034 ;
  assign n7036 = ~n4013 & n7035 ;
  assign n7037 = ~n4170 & n7036 ;
  assign n7038 = ~n4247 & n7037 ;
  assign n7039 = ~n4135 & n7038 ;
  assign n7040 = ~n3914 & n7039 ;
  assign n7041 = ~n4158 & n7040 ;
  assign n7042 = ~n3906 & n7041 ;
  assign n7043 = ~n4142 & n7042 ;
  assign n7044 = n4544 & n6166 ;
  assign n7045 = n3956 & n7044 ;
  assign n7046 = n4568 & n7045 ;
  assign n7047 = n7043 & n7046 ;
  assign n7048 = n4010 & n7047 ;
  assign n7049 = ~n3950 & n7048 ;
  assign n7050 = ~n3976 & n7049 ;
  assign n7051 = ~n4020 & n7050 ;
  assign n7052 = ~n4027 & n7051 ;
  assign n7053 = ~n3986 & n7052 ;
  assign n7054 = ~n4246 & n7053 ;
  assign n7055 = ~n4161 & n7054 ;
  assign n7056 = ~n4277 & n7055 ;
  assign n7057 = n6352 & n7056 ;
  assign n7058 = n7029 & n7057 ;
  assign n7059 = ~n3934 & ~n4205 ;
  assign n7060 = n4149 & n4223 ;
  assign n7061 = n4965 & n7060 ;
  assign n7062 = n4197 & n7061 ;
  assign n7063 = n4237 & n7062 ;
  assign n7064 = n4114 & n7063 ;
  assign n7065 = n4285 & n7064 ;
  assign n7066 = n4302 & n7065 ;
  assign n7067 = n4253 & n7066 ;
  assign n7068 = n7059 & n7067 ;
  assign n7069 = ~n3940 & n7068 ;
  assign n7070 = ~n7058 & n7069 ;
  assign n7071 = n7058 & ~n7069 ;
  assign n7072 = ~n7070 & ~n7071 ;
  assign n7073 = n7017 & n7072 ;
  assign n7074 = n4088 & ~n7015 ;
  assign n7075 = ~n6352 & n7056 ;
  assign n7076 = n6352 & ~n7056 ;
  assign n7077 = ~n7075 & ~n7076 ;
  assign n7078 = n7074 & n7077 ;
  assign n7079 = ~n7029 & ~n7057 ;
  assign n7080 = ~n7058 & ~n7079 ;
  assign n7081 = x0 & ~n7012 ;
  assign n7082 = ~n7080 & n7081 ;
  assign n7083 = ~n7078 & ~n7082 ;
  assign n7084 = ~n7073 & n7083 ;
  assign n7085 = ~n7016 & n7084 ;
  assign n7086 = n7077 & ~n7080 ;
  assign n7087 = ~n6354 & n7077 ;
  assign n7088 = ~n6447 & ~n6450 ;
  assign n7089 = n6354 & ~n7077 ;
  assign n7090 = ~n7087 & ~n7089 ;
  assign n7091 = ~n7088 & n7090 ;
  assign n7092 = ~n7087 & ~n7091 ;
  assign n7093 = ~n7077 & n7080 ;
  assign n7094 = ~n7086 & ~n7093 ;
  assign n7095 = ~n7092 & n7094 ;
  assign n7096 = ~n7086 & ~n7095 ;
  assign n7097 = ~n7072 & n7080 ;
  assign n7098 = n7072 & ~n7080 ;
  assign n7099 = ~n7097 & ~n7098 ;
  assign n7100 = ~n7096 & n7099 ;
  assign n7101 = n7096 & ~n7099 ;
  assign n7102 = ~n7100 & ~n7101 ;
  assign n7103 = n7084 & ~n7102 ;
  assign n7104 = ~n7085 & ~n7103 ;
  assign n7105 = n4091 & ~n7104 ;
  assign n7106 = ~n4091 & n7104 ;
  assign n7107 = ~n7105 & ~n7106 ;
  assign n7108 = n7008 & n7107 ;
  assign n7109 = n6831 & n7003 ;
  assign n7110 = ~n7004 & ~n7109 ;
  assign n7111 = n7017 & ~n7080 ;
  assign n7112 = ~n6354 & n7074 ;
  assign n7113 = n7077 & n7081 ;
  assign n7114 = ~n7112 & ~n7113 ;
  assign n7115 = ~n7111 & n7114 ;
  assign n7116 = ~n7016 & n7115 ;
  assign n7117 = n7092 & ~n7094 ;
  assign n7118 = ~n7095 & ~n7117 ;
  assign n7119 = n7115 & ~n7118 ;
  assign n7120 = ~n7116 & ~n7119 ;
  assign n7121 = n4091 & ~n7120 ;
  assign n7122 = ~n4091 & n7120 ;
  assign n7123 = ~n7121 & ~n7122 ;
  assign n7124 = n7110 & n7123 ;
  assign n7125 = n6999 & ~n7001 ;
  assign n7126 = n7017 & n7077 ;
  assign n7127 = ~n6366 & n7074 ;
  assign n7128 = ~n6354 & n7081 ;
  assign n7129 = ~n7127 & ~n7128 ;
  assign n7130 = ~n7126 & n7129 ;
  assign n7131 = n7088 & ~n7090 ;
  assign n7132 = ~n7091 & ~n7131 ;
  assign n7133 = n7016 & n7132 ;
  assign n7134 = n7130 & ~n7133 ;
  assign n7135 = ~n4091 & ~n7134 ;
  assign n7136 = ~n7134 & ~n7135 ;
  assign n7137 = ~n4091 & ~n7135 ;
  assign n7138 = ~n7136 & ~n7137 ;
  assign n7139 = n6362 & n7017 ;
  assign n7140 = n6378 & n7074 ;
  assign n7141 = ~n6375 & n7081 ;
  assign n7142 = ~n7140 & ~n7141 ;
  assign n7143 = ~n7139 & n7142 ;
  assign n7144 = ~n4091 & ~n7143 ;
  assign n7145 = n6842 & n7016 ;
  assign n7146 = n7143 & ~n7145 ;
  assign n7147 = n4091 & n7146 ;
  assign n7148 = ~n4091 & n7016 ;
  assign n7149 = n6842 & n7148 ;
  assign n7150 = ~n6375 & n7017 ;
  assign n7151 = ~n6382 & n7074 ;
  assign n7152 = n6378 & n7081 ;
  assign n7153 = ~n7151 & ~n7152 ;
  assign n7154 = ~n7150 & n7153 ;
  assign n7155 = ~n4091 & ~n7154 ;
  assign n7156 = n6789 & n7016 ;
  assign n7157 = n7154 & ~n7156 ;
  assign n7158 = n4091 & n7157 ;
  assign n7159 = n6789 & n7148 ;
  assign n7160 = n6378 & n7017 ;
  assign n7161 = ~n6386 & n7074 ;
  assign n7162 = ~n6382 & n7081 ;
  assign n7163 = ~n7161 & ~n7162 ;
  assign n7164 = ~n7160 & n7163 ;
  assign n7165 = ~n4091 & ~n7164 ;
  assign n7166 = n6615 & n7016 ;
  assign n7167 = n7164 & ~n7166 ;
  assign n7168 = n4091 & n7167 ;
  assign n7169 = n6615 & n7148 ;
  assign n7170 = n6972 & ~n6974 ;
  assign n7171 = ~n6386 & n7017 ;
  assign n7172 = n6393 & n7074 ;
  assign n7173 = ~n6390 & n7081 ;
  assign n7174 = ~n7172 & ~n7173 ;
  assign n7175 = ~n7171 & n7174 ;
  assign n7176 = ~n4091 & ~n7175 ;
  assign n7177 = n6649 & n7016 ;
  assign n7178 = n7175 & ~n7177 ;
  assign n7179 = n4091 & n7178 ;
  assign n7180 = n6649 & n7148 ;
  assign n7181 = ~n6944 & ~n6955 ;
  assign n7182 = ~n6400 & n7074 ;
  assign n7183 = n6396 & n7081 ;
  assign n7184 = n6393 & n7017 ;
  assign n7185 = ~n7183 & ~n7184 ;
  assign n7186 = ~n7182 & n7185 ;
  assign n7187 = ~n4091 & ~n7186 ;
  assign n7188 = ~n6506 & n7016 ;
  assign n7189 = n7186 & ~n7188 ;
  assign n7190 = n4091 & n7189 ;
  assign n7191 = ~n6506 & n7148 ;
  assign n7192 = ~x0 & ~n6407 ;
  assign n7193 = n6532 & n7148 ;
  assign n7194 = ~n6400 & n7017 ;
  assign n7195 = ~n6407 & n7074 ;
  assign n7196 = ~n6404 & n7081 ;
  assign n7197 = ~n7195 & ~n7196 ;
  assign n7198 = ~n7194 & n7197 ;
  assign n7199 = ~n4091 & ~n7198 ;
  assign n7200 = ~n6473 & n7148 ;
  assign n7201 = ~n6404 & n7017 ;
  assign n7202 = ~n6407 & n7081 ;
  assign n7203 = ~n4091 & ~n7202 ;
  assign n7204 = ~n7201 & n7203 ;
  assign n7205 = ~n7200 & n7204 ;
  assign n7206 = ~n7199 & n7205 ;
  assign n7207 = ~n7193 & n7206 ;
  assign n7208 = ~n7192 & n7207 ;
  assign n7209 = ~n6934 & ~n7208 ;
  assign n7210 = ~n6400 & n7081 ;
  assign n7211 = n6396 & n7017 ;
  assign n7212 = ~n6404 & n7074 ;
  assign n7213 = ~n7211 & ~n7212 ;
  assign n7214 = ~n7210 & n7213 ;
  assign n7215 = ~n6550 & n7016 ;
  assign n7216 = n7214 & ~n7215 ;
  assign n7217 = ~n4091 & ~n7216 ;
  assign n7218 = n4091 & n7216 ;
  assign n7219 = ~n7217 & ~n7218 ;
  assign n7220 = ~n7209 & n7219 ;
  assign n7221 = n6934 & n7208 ;
  assign n7222 = ~n7220 & ~n7221 ;
  assign n7223 = ~n6935 & ~n6943 ;
  assign n7224 = ~n6944 & ~n7223 ;
  assign n7225 = n7222 & ~n7224 ;
  assign n7226 = ~n7191 & ~n7225 ;
  assign n7227 = ~n7190 & n7226 ;
  assign n7228 = ~n7187 & n7227 ;
  assign n7229 = ~n7222 & n7224 ;
  assign n7230 = ~n7228 & ~n7229 ;
  assign n7231 = ~n6390 & n7017 ;
  assign n7232 = n6396 & n7074 ;
  assign n7233 = n6393 & n7081 ;
  assign n7234 = ~n7232 & ~n7233 ;
  assign n7235 = ~n7231 & n7234 ;
  assign n7236 = n6568 & n7016 ;
  assign n7237 = n7235 & ~n7236 ;
  assign n7238 = ~n4091 & ~n7237 ;
  assign n7239 = ~n7237 & ~n7238 ;
  assign n7240 = ~n4091 & ~n7238 ;
  assign n7241 = ~n7239 & ~n7240 ;
  assign n7242 = n7230 & n7241 ;
  assign n7243 = ~n6956 & ~n7242 ;
  assign n7244 = ~n7181 & n7243 ;
  assign n7245 = ~n7230 & ~n7241 ;
  assign n7246 = ~n7244 & ~n7245 ;
  assign n7247 = ~n6960 & ~n6971 ;
  assign n7248 = n6970 & ~n6971 ;
  assign n7249 = ~n7247 & ~n7248 ;
  assign n7250 = n7246 & n7249 ;
  assign n7251 = ~n7180 & ~n7250 ;
  assign n7252 = ~n7179 & n7251 ;
  assign n7253 = ~n7176 & n7252 ;
  assign n7254 = ~n7246 & ~n7249 ;
  assign n7255 = ~n7253 & ~n7254 ;
  assign n7256 = ~n6382 & n7017 ;
  assign n7257 = ~n6390 & n7074 ;
  assign n7258 = ~n6386 & n7081 ;
  assign n7259 = ~n7257 & ~n7258 ;
  assign n7260 = ~n7256 & n7259 ;
  assign n7261 = n6630 & n7016 ;
  assign n7262 = n7260 & ~n7261 ;
  assign n7263 = ~n4091 & ~n7262 ;
  assign n7264 = ~n7262 & ~n7263 ;
  assign n7265 = ~n4091 & ~n7263 ;
  assign n7266 = ~n7264 & ~n7265 ;
  assign n7267 = n7255 & n7266 ;
  assign n7268 = ~n6975 & ~n7267 ;
  assign n7269 = ~n7170 & n7268 ;
  assign n7270 = ~n7255 & ~n7266 ;
  assign n7271 = ~n7269 & ~n7270 ;
  assign n7272 = n6976 & ~n6978 ;
  assign n7273 = ~n6979 & ~n7272 ;
  assign n7274 = n7271 & ~n7273 ;
  assign n7275 = ~n7169 & ~n7274 ;
  assign n7276 = ~n7168 & n7275 ;
  assign n7277 = ~n7165 & n7276 ;
  assign n7278 = ~n7271 & n7273 ;
  assign n7279 = ~n7277 & ~n7278 ;
  assign n7280 = ~n6980 & ~n6984 ;
  assign n7281 = ~n6983 & ~n6984 ;
  assign n7282 = ~n7280 & ~n7281 ;
  assign n7283 = n7279 & n7282 ;
  assign n7284 = ~n7159 & ~n7283 ;
  assign n7285 = ~n7158 & n7284 ;
  assign n7286 = ~n7155 & n7285 ;
  assign n7287 = ~n7279 & ~n7282 ;
  assign n7288 = ~n7286 & ~n7287 ;
  assign n7289 = n6985 & ~n6987 ;
  assign n7290 = ~n6988 & ~n7289 ;
  assign n7291 = n7288 & ~n7290 ;
  assign n7292 = ~n7149 & ~n7291 ;
  assign n7293 = ~n7147 & n7292 ;
  assign n7294 = ~n7144 & n7293 ;
  assign n7295 = ~n7288 & n7290 ;
  assign n7296 = ~n7294 & ~n7295 ;
  assign n7297 = n6989 & n6992 ;
  assign n7298 = ~n6993 & ~n7297 ;
  assign n7299 = ~n7296 & n7298 ;
  assign n7300 = ~n6366 & n7017 ;
  assign n7301 = ~n6375 & n7074 ;
  assign n7302 = n6362 & n7081 ;
  assign n7303 = ~n7301 & ~n7302 ;
  assign n7304 = ~n7300 & n7303 ;
  assign n7305 = n6822 & n7016 ;
  assign n7306 = n7304 & ~n7305 ;
  assign n7307 = n4091 & ~n7306 ;
  assign n7308 = ~n4091 & n7306 ;
  assign n7309 = ~n7307 & ~n7308 ;
  assign n7310 = ~n7299 & n7309 ;
  assign n7311 = n7296 & ~n7298 ;
  assign n7312 = ~n7310 & ~n7311 ;
  assign n7313 = n6994 & n6997 ;
  assign n7314 = ~n6998 & ~n7313 ;
  assign n7315 = ~n7312 & ~n7314 ;
  assign n7316 = ~n6354 & n7017 ;
  assign n7317 = n6362 & n7074 ;
  assign n7318 = ~n6366 & n7081 ;
  assign n7319 = ~n7317 & ~n7318 ;
  assign n7320 = ~n7316 & n7319 ;
  assign n7321 = n6452 & n7016 ;
  assign n7322 = n7320 & ~n7321 ;
  assign n7323 = ~n4091 & ~n7322 ;
  assign n7324 = n4091 & n7322 ;
  assign n7325 = ~n7323 & ~n7324 ;
  assign n7326 = ~n7315 & n7325 ;
  assign n7327 = n7312 & n7314 ;
  assign n7328 = ~n7326 & ~n7327 ;
  assign n7329 = n7138 & n7328 ;
  assign n7330 = ~n7002 & ~n7329 ;
  assign n7331 = ~n7125 & n7330 ;
  assign n7332 = ~n7138 & ~n7328 ;
  assign n7333 = ~n7331 & ~n7332 ;
  assign n7334 = n7110 & ~n7124 ;
  assign n7335 = n7123 & ~n7124 ;
  assign n7336 = ~n7334 & ~n7335 ;
  assign n7337 = ~n7333 & ~n7336 ;
  assign n7338 = ~n7124 & ~n7337 ;
  assign n7339 = n7008 & ~n7108 ;
  assign n7340 = n7107 & ~n7108 ;
  assign n7341 = ~n7339 & ~n7340 ;
  assign n7342 = ~n7338 & ~n7341 ;
  assign n7343 = ~n7108 & ~n7342 ;
  assign n7344 = ~n6809 & ~n7007 ;
  assign n7345 = n4095 & n7077 ;
  assign n7346 = n6360 & ~n6366 ;
  assign n7347 = ~n6354 & n6367 ;
  assign n7348 = ~n7346 & ~n7347 ;
  assign n7349 = ~n7345 & n7348 ;
  assign n7350 = n6371 & n7132 ;
  assign n7351 = n7349 & ~n7350 ;
  assign n7352 = ~n4075 & ~n7351 ;
  assign n7353 = n4075 & n7351 ;
  assign n7354 = ~n7352 & ~n7353 ;
  assign n7355 = ~n6801 & ~n6805 ;
  assign n7356 = ~n6780 & ~n6786 ;
  assign n7357 = ~n6382 & n6499 ;
  assign n7358 = ~n6390 & n6495 ;
  assign n7359 = ~n6386 & n6497 ;
  assign n7360 = ~n7358 & ~n7359 ;
  assign n7361 = ~n7357 & n7360 ;
  assign n7362 = n6490 & n6630 ;
  assign n7363 = n7361 & ~n7362 ;
  assign n7364 = ~n4469 & ~n7363 ;
  assign n7365 = n4469 & n7363 ;
  assign n7366 = ~n7364 & ~n7365 ;
  assign n7367 = ~n4325 & ~n6404 ;
  assign n7368 = ~n6400 & n6576 ;
  assign n7369 = n6396 & n6466 ;
  assign n7370 = n6393 & n6468 ;
  assign n7371 = ~n7369 & ~n7370 ;
  assign n7372 = ~n7368 & n7371 ;
  assign n7373 = n6474 & ~n6506 ;
  assign n7374 = n7372 & ~n7373 ;
  assign n7375 = ~n4325 & ~n7374 ;
  assign n7376 = n7367 & ~n7375 ;
  assign n7377 = n7367 & ~n7376 ;
  assign n7378 = n4325 & n7374 ;
  assign n7379 = ~n7375 & ~n7378 ;
  assign n7380 = ~n7376 & n7379 ;
  assign n7381 = ~n7377 & ~n7380 ;
  assign n7382 = ~n6777 & ~n7381 ;
  assign n7383 = ~n6777 & ~n7382 ;
  assign n7384 = ~n7381 & ~n7382 ;
  assign n7385 = ~n7383 & ~n7384 ;
  assign n7386 = n7366 & ~n7385 ;
  assign n7387 = n7366 & ~n7386 ;
  assign n7388 = ~n7385 & ~n7386 ;
  assign n7389 = ~n7387 & ~n7388 ;
  assign n7390 = ~n7356 & n7389 ;
  assign n7391 = n7356 & ~n7389 ;
  assign n7392 = ~n7390 & ~n7391 ;
  assign n7393 = n6362 & n6602 ;
  assign n7394 = n6378 & n6608 ;
  assign n7395 = ~n6375 & n6610 ;
  assign n7396 = ~n7394 & ~n7395 ;
  assign n7397 = ~n7393 & n7396 ;
  assign n7398 = ~n6842 & n7397 ;
  assign n7399 = ~n6617 & n7397 ;
  assign n7400 = ~n7398 & ~n7399 ;
  assign n7401 = n4821 & ~n7400 ;
  assign n7402 = ~n4821 & n7400 ;
  assign n7403 = ~n7401 & ~n7402 ;
  assign n7404 = ~n7392 & n7403 ;
  assign n7405 = n7392 & ~n7403 ;
  assign n7406 = ~n7404 & ~n7405 ;
  assign n7407 = ~n7355 & n7406 ;
  assign n7408 = n7355 & ~n7406 ;
  assign n7409 = ~n7407 & ~n7408 ;
  assign n7410 = n7354 & n7409 ;
  assign n7411 = ~n7354 & ~n7409 ;
  assign n7412 = ~n7410 & ~n7411 ;
  assign n7413 = ~n7344 & n7412 ;
  assign n7414 = n7344 & ~n7412 ;
  assign n7415 = ~n7413 & ~n7414 ;
  assign n7416 = ~n4148 & n4302 ;
  assign n7417 = ~n3948 & n7416 ;
  assign n7418 = n4314 & n7417 ;
  assign n7419 = n4285 & n7418 ;
  assign n7420 = n4214 & n7419 ;
  assign n7421 = n4204 & n7420 ;
  assign n7422 = ~n3988 & n7421 ;
  assign n7423 = ~n4019 & n7422 ;
  assign n7424 = ~n4024 & n7423 ;
  assign n7425 = n7058 & n7069 ;
  assign n7426 = ~n7424 & ~n7425 ;
  assign n7427 = n7424 & n7425 ;
  assign n7428 = ~n7426 & ~n7427 ;
  assign n7429 = n7017 & ~n7428 ;
  assign n7430 = n7074 & ~n7080 ;
  assign n7431 = n7072 & n7081 ;
  assign n7432 = ~n7430 & ~n7431 ;
  assign n7433 = ~n7429 & n7432 ;
  assign n7434 = ~n7016 & n7433 ;
  assign n7435 = ~n7098 & ~n7100 ;
  assign n7436 = ~n7072 & n7428 ;
  assign n7437 = n7072 & ~n7428 ;
  assign n7438 = ~n7436 & ~n7437 ;
  assign n7439 = ~n7435 & n7438 ;
  assign n7440 = n7435 & ~n7438 ;
  assign n7441 = ~n7439 & ~n7440 ;
  assign n7442 = n7433 & ~n7441 ;
  assign n7443 = ~n7434 & ~n7442 ;
  assign n7444 = n4091 & ~n7443 ;
  assign n7445 = ~n4091 & n7443 ;
  assign n7446 = ~n7444 & ~n7445 ;
  assign n7447 = n7415 & n7446 ;
  assign n7448 = ~n7415 & ~n7446 ;
  assign n7449 = ~n7447 & ~n7448 ;
  assign n7450 = ~n7343 & n7449 ;
  assign n7451 = n7343 & ~n7449 ;
  assign n7452 = ~n7450 & ~n7451 ;
  assign n7453 = ~n4071 & n7452 ;
  assign n7454 = ~n3914 & ~n4306 ;
  assign n7455 = ~n4536 & n7454 ;
  assign n7456 = ~n4096 & n7455 ;
  assign n7457 = ~n3954 & n7456 ;
  assign n7458 = n4606 & n7457 ;
  assign n7459 = ~n3939 & n7458 ;
  assign n7460 = ~n3950 & n7459 ;
  assign n7461 = ~n3986 & n7460 ;
  assign n7462 = ~n4113 & n7461 ;
  assign n7463 = ~n3933 & n7462 ;
  assign n7464 = ~n4159 & n7463 ;
  assign n7465 = ~n3942 & n7464 ;
  assign n7466 = ~n3906 & n7465 ;
  assign n7467 = n4172 & n4305 ;
  assign n7468 = n4934 & n7467 ;
  assign n7469 = ~n4017 & n7468 ;
  assign n7470 = ~n4055 & n7469 ;
  assign n7471 = ~n4295 & n7470 ;
  assign n7472 = ~n4353 & n7471 ;
  assign n7473 = ~n4245 & n7472 ;
  assign n7474 = ~n4271 & n7473 ;
  assign n7475 = ~n4015 & n7474 ;
  assign n7476 = n4589 & n7475 ;
  assign n7477 = ~n4217 & n7476 ;
  assign n7478 = ~n4098 & n7477 ;
  assign n7479 = n6254 & n7478 ;
  assign n7480 = n7466 & n7479 ;
  assign n7481 = n4780 & n7480 ;
  assign n7482 = ~n3937 & n7481 ;
  assign n7483 = ~n4054 & n7482 ;
  assign n7484 = ~n4127 & n7483 ;
  assign n7485 = ~n4246 & n7484 ;
  assign n7486 = ~n3946 & n7485 ;
  assign n7487 = ~n4097 & n7486 ;
  assign n7488 = ~n4135 & n7487 ;
  assign n7489 = ~n4270 & n7488 ;
  assign n7490 = ~n4142 & n7489 ;
  assign n7491 = n7338 & ~n7340 ;
  assign n7492 = ~n7339 & n7491 ;
  assign n7493 = ~n7342 & ~n7492 ;
  assign n7494 = n4197 & n6078 ;
  assign n7495 = n6103 & n7494 ;
  assign n7496 = ~n3944 & n7495 ;
  assign n7497 = ~n4303 & n7496 ;
  assign n7498 = ~n4156 & n7497 ;
  assign n7499 = ~n4277 & n7498 ;
  assign n7500 = n4141 & n4613 ;
  assign n7501 = ~n3937 & n7500 ;
  assign n7502 = ~n3955 & n7501 ;
  assign n7503 = n4260 & n6222 ;
  assign n7504 = n6233 & n7503 ;
  assign n7505 = n4144 & n7504 ;
  assign n7506 = n7502 & n7505 ;
  assign n7507 = n7499 & n7506 ;
  assign n7508 = n6164 & n7507 ;
  assign n7509 = ~n4215 & n7508 ;
  assign n7510 = ~n3950 & n7509 ;
  assign n7511 = ~n4117 & n7510 ;
  assign n7512 = ~n4019 & n7511 ;
  assign n7513 = ~n3974 & n7512 ;
  assign n7514 = ~n4018 & n7513 ;
  assign n7515 = ~n4102 & n7514 ;
  assign n7516 = n7333 & n7336 ;
  assign n7517 = ~n7337 & ~n7516 ;
  assign n7518 = ~n7515 & n7517 ;
  assign n7519 = ~n7493 & ~n7518 ;
  assign n7520 = ~n7490 & ~n7519 ;
  assign n7521 = n7493 & n7518 ;
  assign n7522 = ~n7520 & ~n7521 ;
  assign n7523 = ~n4071 & ~n7453 ;
  assign n7524 = n7452 & ~n7453 ;
  assign n7525 = ~n7523 & ~n7524 ;
  assign n7526 = ~n7522 & ~n7525 ;
  assign n7527 = ~n7453 & ~n7526 ;
  assign n7528 = n4039 & n4390 ;
  assign n7529 = ~n4150 & n7528 ;
  assign n7530 = ~n3923 & n7529 ;
  assign n7531 = ~n4113 & n7530 ;
  assign n7532 = ~n4007 & n7531 ;
  assign n7533 = ~n4245 & n7532 ;
  assign n7534 = ~n4269 & n7533 ;
  assign n7535 = n4153 & ~n4268 ;
  assign n7536 = n4134 & n7535 ;
  assign n7537 = n4962 & n7536 ;
  assign n7538 = n7534 & n7537 ;
  assign n7539 = n6218 & n7538 ;
  assign n7540 = ~n4022 & n7539 ;
  assign n7541 = ~n4117 & n7540 ;
  assign n7542 = ~n3977 & n7541 ;
  assign n7543 = ~n4018 & n7542 ;
  assign n7544 = ~n4354 & n7543 ;
  assign n7545 = ~n4011 & n7544 ;
  assign n7546 = ~n3932 & n7545 ;
  assign n7547 = ~n4023 & n7546 ;
  assign n7548 = ~n7427 & n7547 ;
  assign n7549 = n7427 & ~n7547 ;
  assign n7550 = ~n7548 & ~n7549 ;
  assign n7551 = n7017 & n7550 ;
  assign n7552 = n7072 & n7074 ;
  assign n7553 = n7081 & ~n7428 ;
  assign n7554 = ~n7552 & ~n7553 ;
  assign n7555 = ~n7551 & n7554 ;
  assign n7556 = ~n7437 & ~n7439 ;
  assign n7557 = n7428 & ~n7550 ;
  assign n7558 = ~n7428 & n7550 ;
  assign n7559 = ~n7557 & ~n7558 ;
  assign n7560 = ~n7556 & n7559 ;
  assign n7561 = n7556 & ~n7559 ;
  assign n7562 = ~n7560 & ~n7561 ;
  assign n7563 = n7016 & n7562 ;
  assign n7564 = n7555 & ~n7563 ;
  assign n7565 = ~n4091 & ~n7564 ;
  assign n7566 = ~n7564 & ~n7565 ;
  assign n7567 = ~n4091 & ~n7565 ;
  assign n7568 = ~n7566 & ~n7567 ;
  assign n7569 = ~n7410 & ~n7413 ;
  assign n7570 = ~n6366 & n6602 ;
  assign n7571 = ~n6375 & n6608 ;
  assign n7572 = n6362 & n6610 ;
  assign n7573 = ~n7571 & ~n7572 ;
  assign n7574 = ~n7570 & n7573 ;
  assign n7575 = n6617 & n6822 ;
  assign n7576 = n7574 & ~n7575 ;
  assign n7577 = ~n4821 & ~n7576 ;
  assign n7578 = ~n7576 & ~n7577 ;
  assign n7579 = ~n4821 & ~n7577 ;
  assign n7580 = ~n7578 & ~n7579 ;
  assign n7581 = ~n7356 & ~n7389 ;
  assign n7582 = ~n7386 & ~n7581 ;
  assign n7583 = ~n7376 & ~n7382 ;
  assign n7584 = ~n6390 & n6468 ;
  assign n7585 = n6396 & n6576 ;
  assign n7586 = n6393 & n6466 ;
  assign n7587 = ~n7585 & ~n7586 ;
  assign n7588 = ~n7584 & n7587 ;
  assign n7589 = n6474 & n6568 ;
  assign n7590 = n7588 & ~n7589 ;
  assign n7591 = ~n4325 & n6400 ;
  assign n7592 = ~n7590 & n7591 ;
  assign n7593 = n7590 & ~n7591 ;
  assign n7594 = ~n7592 & ~n7593 ;
  assign n7595 = ~n7583 & n7594 ;
  assign n7596 = n7583 & ~n7594 ;
  assign n7597 = ~n7595 & ~n7596 ;
  assign n7598 = n6378 & n6499 ;
  assign n7599 = ~n6386 & n6495 ;
  assign n7600 = ~n6382 & n6497 ;
  assign n7601 = ~n7599 & ~n7600 ;
  assign n7602 = ~n7598 & n7601 ;
  assign n7603 = ~n6490 & n7602 ;
  assign n7604 = ~n6615 & n7602 ;
  assign n7605 = ~n7603 & ~n7604 ;
  assign n7606 = n4469 & ~n7605 ;
  assign n7607 = ~n4469 & n7605 ;
  assign n7608 = ~n7606 & ~n7607 ;
  assign n7609 = n7597 & n7608 ;
  assign n7610 = n7597 & ~n7609 ;
  assign n7611 = n7608 & ~n7609 ;
  assign n7612 = ~n7610 & ~n7611 ;
  assign n7613 = ~n7582 & ~n7612 ;
  assign n7614 = ~n7582 & ~n7613 ;
  assign n7615 = ~n7612 & ~n7613 ;
  assign n7616 = ~n7614 & ~n7615 ;
  assign n7617 = ~n7580 & ~n7616 ;
  assign n7618 = ~n7580 & ~n7617 ;
  assign n7619 = ~n7616 & ~n7617 ;
  assign n7620 = ~n7618 & ~n7619 ;
  assign n7621 = ~n7404 & ~n7407 ;
  assign n7622 = n7620 & n7621 ;
  assign n7623 = ~n7620 & ~n7621 ;
  assign n7624 = ~n7622 & ~n7623 ;
  assign n7625 = n4095 & ~n7080 ;
  assign n7626 = ~n6354 & n6360 ;
  assign n7627 = n6367 & n7077 ;
  assign n7628 = ~n7626 & ~n7627 ;
  assign n7629 = ~n7625 & n7628 ;
  assign n7630 = ~n6371 & n7629 ;
  assign n7631 = ~n7118 & n7629 ;
  assign n7632 = ~n7630 & ~n7631 ;
  assign n7633 = n4075 & ~n7632 ;
  assign n7634 = ~n4075 & n7632 ;
  assign n7635 = ~n7633 & ~n7634 ;
  assign n7636 = n7624 & n7635 ;
  assign n7637 = n7624 & ~n7636 ;
  assign n7638 = n7635 & ~n7636 ;
  assign n7639 = ~n7637 & ~n7638 ;
  assign n7640 = ~n7569 & ~n7639 ;
  assign n7641 = ~n7569 & ~n7640 ;
  assign n7642 = ~n7639 & ~n7640 ;
  assign n7643 = ~n7641 & ~n7642 ;
  assign n7644 = ~n7568 & ~n7643 ;
  assign n7645 = ~n7568 & ~n7644 ;
  assign n7646 = ~n7643 & ~n7644 ;
  assign n7647 = ~n7645 & ~n7646 ;
  assign n7648 = ~n7447 & ~n7450 ;
  assign n7649 = n7647 & n7648 ;
  assign n7650 = ~n7647 & ~n7648 ;
  assign n7651 = ~n7649 & ~n7650 ;
  assign n7652 = n4039 & n4893 ;
  assign n7653 = n4606 & n7652 ;
  assign n7654 = n5259 & n7653 ;
  assign n7655 = n6111 & n7654 ;
  assign n7656 = n4443 & n7655 ;
  assign n7657 = n4423 & n7656 ;
  assign n7658 = n4010 & n7657 ;
  assign n7659 = ~n4055 & n7658 ;
  assign n7660 = ~n3948 & n7659 ;
  assign n7661 = ~n4145 & n7660 ;
  assign n7662 = ~n7651 & n7661 ;
  assign n7663 = n7651 & ~n7661 ;
  assign n7664 = ~n7662 & ~n7663 ;
  assign n7665 = ~n7527 & n7664 ;
  assign n7666 = n7527 & ~n7664 ;
  assign n7667 = ~n7665 & ~n7666 ;
  assign n7668 = ~n7522 & ~n7526 ;
  assign n7669 = ~n7525 & ~n7526 ;
  assign n7670 = ~n7668 & ~n7669 ;
  assign n7671 = n7667 & ~n7670 ;
  assign n7672 = n7667 & ~n7671 ;
  assign n7673 = ~n7670 & ~n7671 ;
  assign n7674 = ~n7672 & ~n7673 ;
  assign n7677 = n7674 & ~x24 ;
  assign n7678 = ~n7676 & ~n7677 ;
  assign n7679 = ~n3838 & ~n3840 ;
  assign n7680 = n3602 & n3722 ;
  assign n7681 = n211 & n2408 ;
  assign n7682 = n432 & n7681 ;
  assign n7683 = n728 & n7682 ;
  assign n7684 = ~n144 & n7683 ;
  assign n7685 = ~n93 & n7684 ;
  assign n7686 = ~n141 & n7685 ;
  assign n7687 = ~n143 & n7686 ;
  assign n7688 = n291 & n530 ;
  assign n7689 = n790 & n7688 ;
  assign n7690 = n1451 & n7689 ;
  assign n7691 = n7687 & n7690 ;
  assign n7692 = n2407 & n7691 ;
  assign n7693 = n951 & n7692 ;
  assign n7694 = ~n470 & n7693 ;
  assign n7695 = ~n445 & n7694 ;
  assign n7696 = ~n342 & n7695 ;
  assign n7697 = ~n301 & n7696 ;
  assign n7698 = ~n7680 & n7697 ;
  assign n7699 = n7680 & ~n7697 ;
  assign n7700 = ~n7698 & ~n7699 ;
  assign n7701 = n3192 & n7700 ;
  assign n7702 = n3249 & ~n3603 ;
  assign n7703 = n3256 & n3725 ;
  assign n7704 = ~n7702 & ~n7703 ;
  assign n7705 = ~n7701 & n7704 ;
  assign n7706 = ~n3733 & ~n3735 ;
  assign n7707 = ~n3725 & ~n7700 ;
  assign n7708 = n3725 & n7700 ;
  assign n7709 = ~n7707 & ~n7708 ;
  assign n7710 = ~n7706 & n7709 ;
  assign n7711 = n7706 & ~n7709 ;
  assign n7712 = ~n7710 & ~n7711 ;
  assign n7713 = n3191 & n7712 ;
  assign n7714 = n7705 & ~n7713 ;
  assign n7715 = ~n266 & ~n7714 ;
  assign n7716 = ~n7714 & ~n7715 ;
  assign n7717 = ~n266 & ~n7715 ;
  assign n7718 = ~n7716 & ~n7717 ;
  assign n7719 = ~n3811 & ~n3815 ;
  assign n7720 = ~n2529 & n2777 ;
  assign n7721 = n2537 & n2783 ;
  assign n7722 = ~n2541 & n2785 ;
  assign n7723 = ~n7721 & ~n7722 ;
  assign n7724 = ~n7720 & n7723 ;
  assign n7725 = n2627 & n2792 ;
  assign n7726 = n7724 & ~n7725 ;
  assign n7727 = ~n996 & ~n7726 ;
  assign n7728 = ~n7726 & ~n7727 ;
  assign n7729 = ~n996 & ~n7727 ;
  assign n7730 = ~n7728 & ~n7729 ;
  assign n7731 = ~n3784 & ~n3788 ;
  assign n7732 = ~n500 & ~n2575 ;
  assign n7733 = n3765 & n7732 ;
  assign n7734 = ~n3770 & ~n7733 ;
  assign n7735 = ~n2561 & n2643 ;
  assign n7736 = n2568 & n2751 ;
  assign n7737 = ~n2565 & n2641 ;
  assign n7738 = ~n7736 & ~n7737 ;
  assign n7739 = ~n7735 & n7738 ;
  assign n7740 = n2649 & n2824 ;
  assign n7741 = n7739 & ~n7740 ;
  assign n7742 = ~n500 & ~n2571 ;
  assign n7743 = ~n7741 & n7742 ;
  assign n7744 = n7741 & ~n7742 ;
  assign n7745 = ~n7743 & ~n7744 ;
  assign n7746 = ~n7734 & n7745 ;
  assign n7747 = ~n7734 & ~n7746 ;
  assign n7748 = n7745 & ~n7746 ;
  assign n7749 = ~n7747 & ~n7748 ;
  assign n7750 = ~n2550 & n2674 ;
  assign n7751 = ~n2557 & n2670 ;
  assign n7752 = n2553 & n2672 ;
  assign n7753 = ~n7751 & ~n7752 ;
  assign n7754 = ~n7750 & n7753 ;
  assign n7755 = ~n2665 & n7754 ;
  assign n7756 = ~n2964 & n7754 ;
  assign n7757 = ~n7755 & ~n7756 ;
  assign n7758 = n644 & ~n7757 ;
  assign n7759 = ~n644 & n7757 ;
  assign n7760 = ~n7758 & ~n7759 ;
  assign n7761 = ~n7749 & n7760 ;
  assign n7762 = ~n7749 & ~n7761 ;
  assign n7763 = n7760 & ~n7761 ;
  assign n7764 = ~n7762 & ~n7763 ;
  assign n7765 = ~n7731 & ~n7764 ;
  assign n7766 = ~n7731 & ~n7765 ;
  assign n7767 = ~n7764 & ~n7765 ;
  assign n7768 = ~n7766 & ~n7767 ;
  assign n7769 = ~n7730 & ~n7768 ;
  assign n7770 = ~n7730 & ~n7769 ;
  assign n7771 = ~n7768 & ~n7769 ;
  assign n7772 = ~n7770 & ~n7771 ;
  assign n7773 = ~n3792 & ~n3798 ;
  assign n7774 = n7772 & n7773 ;
  assign n7775 = ~n7772 & ~n7773 ;
  assign n7776 = ~n7774 & ~n7775 ;
  assign n7777 = n270 & n3247 ;
  assign n7778 = n2535 & n3252 ;
  assign n7779 = n2542 & ~n3255 ;
  assign n7780 = ~n7778 & ~n7779 ;
  assign n7781 = ~n7777 & n7780 ;
  assign n7782 = ~n2546 & n7781 ;
  assign n7783 = ~n3277 & n7781 ;
  assign n7784 = ~n7782 & ~n7783 ;
  assign n7785 = n250 & ~n7784 ;
  assign n7786 = ~n250 & n7784 ;
  assign n7787 = ~n7785 & ~n7786 ;
  assign n7788 = n7776 & n7787 ;
  assign n7789 = n7776 & ~n7788 ;
  assign n7790 = n7787 & ~n7788 ;
  assign n7791 = ~n7789 & ~n7790 ;
  assign n7792 = ~n7719 & ~n7791 ;
  assign n7793 = ~n7719 & ~n7792 ;
  assign n7794 = ~n7791 & ~n7792 ;
  assign n7795 = ~n7793 & ~n7794 ;
  assign n7796 = ~n7718 & ~n7795 ;
  assign n7797 = ~n7718 & ~n7796 ;
  assign n7798 = ~n7795 & ~n7796 ;
  assign n7799 = ~n7797 & ~n7798 ;
  assign n7800 = ~n3819 & ~n3825 ;
  assign n7801 = n7799 & n7800 ;
  assign n7802 = ~n7799 & ~n7800 ;
  assign n7803 = ~n7801 & ~n7802 ;
  assign n7804 = ~n115 & ~n380 ;
  assign n7805 = ~n336 & n7804 ;
  assign n7806 = ~n233 & n7805 ;
  assign n7807 = n612 & n2315 ;
  assign n7808 = n2251 & n7807 ;
  assign n7809 = n224 & n7808 ;
  assign n7810 = n728 & n7809 ;
  assign n7811 = n7806 & n7810 ;
  assign n7812 = n185 & n7811 ;
  assign n7813 = n3206 & n7812 ;
  assign n7814 = ~n150 & n7813 ;
  assign n7815 = ~n130 & n7814 ;
  assign n7816 = ~n302 & n7815 ;
  assign n7817 = ~n166 & n7816 ;
  assign n7818 = ~n93 & n7817 ;
  assign n7819 = ~n420 & n7818 ;
  assign n7820 = ~n7803 & n7819 ;
  assign n7821 = n7803 & ~n7819 ;
  assign n7822 = ~n7820 & ~n7821 ;
  assign n7823 = ~n7679 & n7822 ;
  assign n7824 = n7679 & ~n7822 ;
  assign n7825 = ~n7823 & ~n7824 ;
  assign n7826 = n3846 & n7825 ;
  assign n7827 = ~n3846 & ~n7825 ;
  assign n7828 = ~n7826 & ~n7827 ;
  assign n7829 = x22 & ~x23 ;
  assign n7830 = ~x22 & x23 ;
  assign n7831 = ~n7829 & ~n7830 ;
  assign n7832 = ~n3849 & ~n7831 ;
  assign n7833 = ~n7828 & n7832 ;
  assign n7834 = n7828 & ~n7832 ;
  assign n7835 = ~n7833 & ~n7834 ;
  assign n7991 = ~n7835 & x25 ;
  assign n7836 = ~n7663 & ~n7665 ;
  assign n7837 = n7427 & n7547 ;
  assign n7838 = n4036 & n6233 ;
  assign n7839 = n4257 & n7838 ;
  assign n7840 = n4553 & n7839 ;
  assign n7841 = ~n3969 & n7840 ;
  assign n7842 = ~n3918 & n7841 ;
  assign n7843 = ~n3966 & n7842 ;
  assign n7844 = ~n3968 & n7843 ;
  assign n7845 = n4116 & n4355 ;
  assign n7846 = n4615 & n7845 ;
  assign n7847 = n5276 & n7846 ;
  assign n7848 = n7844 & n7847 ;
  assign n7849 = n6232 & n7848 ;
  assign n7850 = n4776 & n7849 ;
  assign n7851 = ~n4295 & n7850 ;
  assign n7852 = ~n4270 & n7851 ;
  assign n7853 = ~n4167 & n7852 ;
  assign n7854 = ~n4126 & n7853 ;
  assign n7855 = ~n7837 & n7854 ;
  assign n7856 = n7837 & ~n7854 ;
  assign n7857 = ~n7855 & ~n7856 ;
  assign n7858 = n7017 & n7857 ;
  assign n7859 = n7074 & ~n7428 ;
  assign n7860 = n7081 & n7550 ;
  assign n7861 = ~n7859 & ~n7860 ;
  assign n7862 = ~n7858 & n7861 ;
  assign n7863 = ~n7558 & ~n7560 ;
  assign n7864 = ~n7550 & ~n7857 ;
  assign n7865 = n7550 & n7857 ;
  assign n7866 = ~n7864 & ~n7865 ;
  assign n7867 = ~n7863 & n7866 ;
  assign n7868 = n7863 & ~n7866 ;
  assign n7869 = ~n7867 & ~n7868 ;
  assign n7870 = n7016 & n7869 ;
  assign n7871 = n7862 & ~n7870 ;
  assign n7872 = ~n4091 & ~n7871 ;
  assign n7873 = ~n7871 & ~n7872 ;
  assign n7874 = ~n4091 & ~n7872 ;
  assign n7875 = ~n7873 & ~n7874 ;
  assign n7876 = ~n7636 & ~n7640 ;
  assign n7877 = ~n6354 & n6602 ;
  assign n7878 = n6362 & n6608 ;
  assign n7879 = ~n6366 & n6610 ;
  assign n7880 = ~n7878 & ~n7879 ;
  assign n7881 = ~n7877 & n7880 ;
  assign n7882 = n6452 & n6617 ;
  assign n7883 = n7881 & ~n7882 ;
  assign n7884 = ~n4821 & ~n7883 ;
  assign n7885 = ~n7883 & ~n7884 ;
  assign n7886 = ~n4821 & ~n7884 ;
  assign n7887 = ~n7885 & ~n7886 ;
  assign n7888 = ~n7609 & ~n7613 ;
  assign n7889 = ~n4325 & ~n6400 ;
  assign n7890 = n7590 & n7889 ;
  assign n7891 = ~n7595 & ~n7890 ;
  assign n7892 = ~n6386 & n6468 ;
  assign n7893 = n6393 & n6576 ;
  assign n7894 = ~n6390 & n6466 ;
  assign n7895 = ~n7893 & ~n7894 ;
  assign n7896 = ~n7892 & n7895 ;
  assign n7897 = n6474 & n6649 ;
  assign n7898 = n7896 & ~n7897 ;
  assign n7899 = ~n4325 & ~n6396 ;
  assign n7900 = ~n7898 & n7899 ;
  assign n7901 = n7898 & ~n7899 ;
  assign n7902 = ~n7900 & ~n7901 ;
  assign n7903 = ~n7891 & n7902 ;
  assign n7904 = ~n7891 & ~n7903 ;
  assign n7905 = n7902 & ~n7903 ;
  assign n7906 = ~n7904 & ~n7905 ;
  assign n7907 = ~n6375 & n6499 ;
  assign n7908 = ~n6382 & n6495 ;
  assign n7909 = n6378 & n6497 ;
  assign n7910 = ~n7908 & ~n7909 ;
  assign n7911 = ~n7907 & n7910 ;
  assign n7912 = ~n6490 & n7911 ;
  assign n7913 = ~n6789 & n7911 ;
  assign n7914 = ~n7912 & ~n7913 ;
  assign n7915 = n4469 & ~n7914 ;
  assign n7916 = ~n4469 & n7914 ;
  assign n7917 = ~n7915 & ~n7916 ;
  assign n7918 = ~n7906 & n7917 ;
  assign n7919 = ~n7906 & ~n7918 ;
  assign n7920 = n7917 & ~n7918 ;
  assign n7921 = ~n7919 & ~n7920 ;
  assign n7922 = ~n7888 & ~n7921 ;
  assign n7923 = ~n7888 & ~n7922 ;
  assign n7924 = ~n7921 & ~n7922 ;
  assign n7925 = ~n7923 & ~n7924 ;
  assign n7926 = ~n7887 & ~n7925 ;
  assign n7927 = ~n7887 & ~n7926 ;
  assign n7928 = ~n7925 & ~n7926 ;
  assign n7929 = ~n7927 & ~n7928 ;
  assign n7930 = ~n7617 & ~n7623 ;
  assign n7931 = n7929 & n7930 ;
  assign n7932 = ~n7929 & ~n7930 ;
  assign n7933 = ~n7931 & ~n7932 ;
  assign n7934 = n4095 & n7072 ;
  assign n7935 = n6360 & n7077 ;
  assign n7936 = n6367 & ~n7080 ;
  assign n7937 = ~n7935 & ~n7936 ;
  assign n7938 = ~n7934 & n7937 ;
  assign n7939 = ~n6371 & n7938 ;
  assign n7940 = ~n7102 & n7938 ;
  assign n7941 = ~n7939 & ~n7940 ;
  assign n7942 = n4075 & ~n7941 ;
  assign n7943 = ~n4075 & n7941 ;
  assign n7944 = ~n7942 & ~n7943 ;
  assign n7945 = n7933 & n7944 ;
  assign n7946 = n7933 & ~n7945 ;
  assign n7947 = n7944 & ~n7945 ;
  assign n7948 = ~n7946 & ~n7947 ;
  assign n7949 = ~n7876 & ~n7948 ;
  assign n7950 = ~n7876 & ~n7949 ;
  assign n7951 = ~n7948 & ~n7949 ;
  assign n7952 = ~n7950 & ~n7951 ;
  assign n7953 = ~n7875 & ~n7952 ;
  assign n7954 = ~n7875 & ~n7953 ;
  assign n7955 = ~n7952 & ~n7953 ;
  assign n7956 = ~n7954 & ~n7955 ;
  assign n7957 = ~n7644 & ~n7650 ;
  assign n7958 = n7956 & n7957 ;
  assign n7959 = ~n7956 & ~n7957 ;
  assign n7960 = ~n7958 & ~n7959 ;
  assign n7961 = ~n3940 & ~n4205 ;
  assign n7962 = ~n4161 & n7961 ;
  assign n7963 = ~n4058 & n7962 ;
  assign n7964 = n4437 & n6140 ;
  assign n7965 = n6076 & n7964 ;
  assign n7966 = n4049 & n7965 ;
  assign n7967 = n4553 & n7966 ;
  assign n7968 = n7963 & n7967 ;
  assign n7969 = n4010 & n7968 ;
  assign n7970 = n7031 & n7969 ;
  assign n7971 = ~n3975 & n7970 ;
  assign n7972 = ~n3955 & n7971 ;
  assign n7973 = ~n4127 & n7972 ;
  assign n7974 = ~n3991 & n7973 ;
  assign n7975 = ~n3918 & n7974 ;
  assign n7976 = ~n4245 & n7975 ;
  assign n7977 = ~n7960 & n7976 ;
  assign n7978 = n7960 & ~n7976 ;
  assign n7979 = ~n7977 & ~n7978 ;
  assign n7980 = ~n7836 & n7979 ;
  assign n7981 = n7836 & ~n7979 ;
  assign n7982 = ~n7980 & ~n7981 ;
  assign n7983 = n7671 & n7982 ;
  assign n7984 = ~n7671 & ~n7982 ;
  assign n7985 = ~n7983 & ~n7984 ;
  assign n7986 = ~n7674 & ~n7831 ;
  assign n7987 = ~n7985 & n7986 ;
  assign n7988 = n7985 & ~n7986 ;
  assign n7989 = ~n7987 & ~n7988 ;
  assign n7992 = n7989 & ~x25 ;
  assign n7993 = ~n7991 & ~n7992 ;
  assign n7994 = ~n7821 & ~n7823 ;
  assign n7995 = n321 & ~n383 ;
  assign n7996 = ~n104 & n7995 ;
  assign n7997 = ~n203 & n7996 ;
  assign n7998 = ~n117 & n7997 ;
  assign n7999 = ~n107 & n7998 ;
  assign n8000 = n391 & n583 ;
  assign n8001 = n780 & n8000 ;
  assign n8002 = n7999 & n8001 ;
  assign n8003 = n3674 & n8002 ;
  assign n8004 = ~n288 & n8003 ;
  assign n8005 = ~n433 & n8004 ;
  assign n8006 = ~n479 & n8005 ;
  assign n8007 = ~n273 & n8006 ;
  assign n8008 = ~n121 & n8007 ;
  assign n8009 = ~n481 & n8008 ;
  assign n8010 = ~n301 & n8009 ;
  assign n8011 = ~n7796 & ~n7802 ;
  assign n8012 = n3249 & n3725 ;
  assign n8013 = n3256 & n7700 ;
  assign n8014 = ~n8012 & ~n8013 ;
  assign n8015 = ~n3725 & ~n7710 ;
  assign n8016 = n7700 & ~n8015 ;
  assign n8017 = ~n7700 & ~n7710 ;
  assign n8018 = ~n8016 & ~n8017 ;
  assign n8019 = n3191 & n8018 ;
  assign n8020 = n8014 & ~n8019 ;
  assign n8021 = ~n266 & ~n8020 ;
  assign n8022 = ~n8020 & ~n8021 ;
  assign n8023 = ~n266 & ~n8021 ;
  assign n8024 = ~n8022 & ~n8023 ;
  assign n8025 = ~n7788 & ~n7792 ;
  assign n8026 = n2777 & n3252 ;
  assign n8027 = ~n2541 & n2783 ;
  assign n8028 = ~n2529 & n2785 ;
  assign n8029 = ~n8027 & ~n8028 ;
  assign n8030 = ~n8026 & n8029 ;
  assign n8031 = n2792 & n3307 ;
  assign n8032 = n8030 & ~n8031 ;
  assign n8033 = ~n996 & ~n8032 ;
  assign n8034 = ~n8032 & ~n8033 ;
  assign n8035 = ~n996 & ~n8033 ;
  assign n8036 = ~n8034 & ~n8035 ;
  assign n8037 = ~n7761 & ~n7765 ;
  assign n8038 = ~n500 & n7741 ;
  assign n8039 = n2571 & n8038 ;
  assign n8040 = ~n7746 & ~n8039 ;
  assign n8041 = ~n2557 & n2643 ;
  assign n8042 = ~n2565 & n2751 ;
  assign n8043 = ~n2561 & n2641 ;
  assign n8044 = ~n8042 & ~n8043 ;
  assign n8045 = ~n8041 & n8044 ;
  assign n8046 = n2649 & n2805 ;
  assign n8047 = n8045 & ~n8046 ;
  assign n8048 = ~n500 & ~n2568 ;
  assign n8049 = ~n8047 & n8048 ;
  assign n8050 = n8047 & ~n8048 ;
  assign n8051 = ~n8049 & ~n8050 ;
  assign n8052 = ~n8040 & n8051 ;
  assign n8053 = ~n8040 & ~n8052 ;
  assign n8054 = n8051 & ~n8052 ;
  assign n8055 = ~n8053 & ~n8054 ;
  assign n8056 = n2537 & n2674 ;
  assign n8057 = n2553 & n2670 ;
  assign n8058 = ~n2550 & n2672 ;
  assign n8059 = ~n8057 & ~n8058 ;
  assign n8060 = ~n8056 & n8059 ;
  assign n8061 = ~n2665 & n8060 ;
  assign n8062 = ~n3017 & n8060 ;
  assign n8063 = ~n8061 & ~n8062 ;
  assign n8064 = n644 & ~n8063 ;
  assign n8065 = ~n644 & n8063 ;
  assign n8066 = ~n8064 & ~n8065 ;
  assign n8067 = ~n8055 & n8066 ;
  assign n8068 = ~n8055 & ~n8067 ;
  assign n8069 = n8066 & ~n8067 ;
  assign n8070 = ~n8068 & ~n8069 ;
  assign n8071 = ~n8037 & ~n8070 ;
  assign n8072 = ~n8037 & ~n8071 ;
  assign n8073 = ~n8070 & ~n8071 ;
  assign n8074 = ~n8072 & ~n8073 ;
  assign n8075 = ~n8036 & ~n8074 ;
  assign n8076 = ~n8036 & ~n8075 ;
  assign n8077 = ~n8074 & ~n8075 ;
  assign n8078 = ~n8076 & ~n8077 ;
  assign n8079 = ~n7769 & ~n7775 ;
  assign n8080 = n8078 & n8079 ;
  assign n8081 = ~n8078 & ~n8079 ;
  assign n8082 = ~n8080 & ~n8081 ;
  assign n8083 = n270 & ~n3603 ;
  assign n8084 = n2535 & ~n3255 ;
  assign n8085 = n2542 & n3247 ;
  assign n8086 = ~n8084 & ~n8085 ;
  assign n8087 = ~n8083 & n8086 ;
  assign n8088 = ~n2546 & n8087 ;
  assign n8089 = ~n3616 & n8087 ;
  assign n8090 = ~n8088 & ~n8089 ;
  assign n8091 = n250 & ~n8090 ;
  assign n8092 = ~n250 & n8090 ;
  assign n8093 = ~n8091 & ~n8092 ;
  assign n8094 = n8082 & n8093 ;
  assign n8095 = n8082 & ~n8094 ;
  assign n8096 = n8093 & ~n8094 ;
  assign n8097 = ~n8095 & ~n8096 ;
  assign n8098 = ~n8025 & ~n8097 ;
  assign n8099 = ~n8025 & ~n8098 ;
  assign n8100 = ~n8097 & ~n8098 ;
  assign n8101 = ~n8099 & ~n8100 ;
  assign n8102 = ~n8024 & ~n8101 ;
  assign n8103 = ~n8024 & ~n8102 ;
  assign n8104 = ~n8101 & ~n8102 ;
  assign n8105 = ~n8103 & ~n8104 ;
  assign n8106 = ~n8011 & n8105 ;
  assign n8107 = n8011 & ~n8105 ;
  assign n8108 = ~n8106 & ~n8107 ;
  assign n8109 = ~n8010 & ~n8108 ;
  assign n8110 = n8010 & n8108 ;
  assign n8111 = ~n7994 & ~n8110 ;
  assign n8112 = ~n8109 & n8111 ;
  assign n8113 = ~n7994 & ~n8112 ;
  assign n8114 = ~n8109 & ~n8112 ;
  assign n8115 = ~n8110 & n8114 ;
  assign n8116 = ~n8113 & ~n8115 ;
  assign n8117 = ~n7826 & n8116 ;
  assign n8118 = n7826 & ~n8116 ;
  assign n8119 = ~n8117 & ~n8118 ;
  assign n8120 = n3849 & ~n7828 ;
  assign n8121 = ~n7831 & ~n8120 ;
  assign n8122 = ~n8119 & n8121 ;
  assign n8123 = n8119 & ~n8121 ;
  assign n8124 = ~n8122 & ~n8123 ;
  assign n8257 = ~n8124 & x26 ;
  assign n8125 = ~n7978 & ~n7980 ;
  assign n8126 = n4146 & ~n4208 ;
  assign n8127 = ~n3929 & n8126 ;
  assign n8128 = ~n4028 & n8127 ;
  assign n8129 = ~n3942 & n8128 ;
  assign n8130 = ~n3932 & n8129 ;
  assign n8131 = n4216 & n4408 ;
  assign n8132 = n4605 & n8131 ;
  assign n8133 = n8130 & n8132 ;
  assign n8134 = n7499 & n8133 ;
  assign n8135 = ~n4113 & n8134 ;
  assign n8136 = ~n4258 & n8135 ;
  assign n8137 = ~n4304 & n8136 ;
  assign n8138 = ~n4098 & n8137 ;
  assign n8139 = ~n3946 & n8138 ;
  assign n8140 = ~n4306 & n8139 ;
  assign n8141 = ~n4126 & n8140 ;
  assign n8142 = ~n7953 & ~n7959 ;
  assign n8143 = n7074 & n7550 ;
  assign n8144 = n7081 & n7857 ;
  assign n8145 = ~n8143 & ~n8144 ;
  assign n8146 = ~n7550 & ~n7867 ;
  assign n8147 = n7857 & ~n8146 ;
  assign n8148 = ~n7857 & ~n7867 ;
  assign n8149 = ~n8147 & ~n8148 ;
  assign n8150 = n7016 & n8149 ;
  assign n8151 = n8145 & ~n8150 ;
  assign n8152 = ~n4091 & ~n8151 ;
  assign n8153 = ~n8151 & ~n8152 ;
  assign n8154 = ~n4091 & ~n8152 ;
  assign n8155 = ~n8153 & ~n8154 ;
  assign n8156 = ~n7945 & ~n7949 ;
  assign n8157 = n6602 & n7077 ;
  assign n8158 = ~n6366 & n6608 ;
  assign n8159 = ~n6354 & n6610 ;
  assign n8160 = ~n8158 & ~n8159 ;
  assign n8161 = ~n8157 & n8160 ;
  assign n8162 = n6617 & n7132 ;
  assign n8163 = n8161 & ~n8162 ;
  assign n8164 = ~n4821 & ~n8163 ;
  assign n8165 = ~n8163 & ~n8164 ;
  assign n8166 = ~n4821 & ~n8164 ;
  assign n8167 = ~n8165 & ~n8166 ;
  assign n8168 = ~n7918 & ~n7922 ;
  assign n8169 = ~n4325 & n7898 ;
  assign n8170 = n6396 & n8169 ;
  assign n8171 = ~n7903 & ~n8170 ;
  assign n8172 = ~n6382 & n6468 ;
  assign n8173 = ~n6390 & n6576 ;
  assign n8174 = ~n6386 & n6466 ;
  assign n8175 = ~n8173 & ~n8174 ;
  assign n8176 = ~n8172 & n8175 ;
  assign n8177 = n6474 & n6630 ;
  assign n8178 = n8176 & ~n8177 ;
  assign n8179 = ~n4325 & ~n6393 ;
  assign n8180 = ~n8178 & n8179 ;
  assign n8181 = n8178 & ~n8179 ;
  assign n8182 = ~n8180 & ~n8181 ;
  assign n8183 = ~n8171 & n8182 ;
  assign n8184 = ~n8171 & ~n8183 ;
  assign n8185 = n8182 & ~n8183 ;
  assign n8186 = ~n8184 & ~n8185 ;
  assign n8187 = n6362 & n6499 ;
  assign n8188 = n6378 & n6495 ;
  assign n8189 = ~n6375 & n6497 ;
  assign n8190 = ~n8188 & ~n8189 ;
  assign n8191 = ~n8187 & n8190 ;
  assign n8192 = ~n6490 & n8191 ;
  assign n8193 = ~n6842 & n8191 ;
  assign n8194 = ~n8192 & ~n8193 ;
  assign n8195 = n4469 & ~n8194 ;
  assign n8196 = ~n4469 & n8194 ;
  assign n8197 = ~n8195 & ~n8196 ;
  assign n8198 = ~n8186 & n8197 ;
  assign n8199 = ~n8186 & ~n8198 ;
  assign n8200 = n8197 & ~n8198 ;
  assign n8201 = ~n8199 & ~n8200 ;
  assign n8202 = ~n8168 & ~n8201 ;
  assign n8203 = ~n8168 & ~n8202 ;
  assign n8204 = ~n8201 & ~n8202 ;
  assign n8205 = ~n8203 & ~n8204 ;
  assign n8206 = ~n8167 & ~n8205 ;
  assign n8207 = ~n8167 & ~n8206 ;
  assign n8208 = ~n8205 & ~n8206 ;
  assign n8209 = ~n8207 & ~n8208 ;
  assign n8210 = ~n7926 & ~n7932 ;
  assign n8211 = n8209 & n8210 ;
  assign n8212 = ~n8209 & ~n8210 ;
  assign n8213 = ~n8211 & ~n8212 ;
  assign n8214 = n4095 & ~n7428 ;
  assign n8215 = n6360 & ~n7080 ;
  assign n8216 = n6367 & n7072 ;
  assign n8217 = ~n8215 & ~n8216 ;
  assign n8218 = ~n8214 & n8217 ;
  assign n8219 = ~n6371 & n8218 ;
  assign n8220 = ~n7441 & n8218 ;
  assign n8221 = ~n8219 & ~n8220 ;
  assign n8222 = n4075 & ~n8221 ;
  assign n8223 = ~n4075 & n8221 ;
  assign n8224 = ~n8222 & ~n8223 ;
  assign n8225 = n8213 & n8224 ;
  assign n8226 = n8213 & ~n8225 ;
  assign n8227 = n8224 & ~n8225 ;
  assign n8228 = ~n8226 & ~n8227 ;
  assign n8229 = ~n8156 & ~n8228 ;
  assign n8230 = ~n8156 & ~n8229 ;
  assign n8231 = ~n8228 & ~n8229 ;
  assign n8232 = ~n8230 & ~n8231 ;
  assign n8233 = ~n8155 & ~n8232 ;
  assign n8234 = ~n8155 & ~n8233 ;
  assign n8235 = ~n8232 & ~n8233 ;
  assign n8236 = ~n8234 & ~n8235 ;
  assign n8237 = ~n8142 & n8236 ;
  assign n8238 = n8142 & ~n8236 ;
  assign n8239 = ~n8237 & ~n8238 ;
  assign n8240 = ~n8141 & ~n8239 ;
  assign n8241 = n8141 & n8239 ;
  assign n8242 = ~n8125 & ~n8241 ;
  assign n8243 = ~n8240 & n8242 ;
  assign n8244 = ~n8125 & ~n8243 ;
  assign n8245 = ~n8240 & ~n8243 ;
  assign n8246 = ~n8241 & n8245 ;
  assign n8247 = ~n8244 & ~n8246 ;
  assign n8248 = ~n7983 & n8247 ;
  assign n8249 = n7983 & ~n8247 ;
  assign n8250 = ~n8248 & ~n8249 ;
  assign n8251 = n7674 & ~n7985 ;
  assign n8252 = ~n7831 & ~n8251 ;
  assign n8253 = ~n8250 & n8252 ;
  assign n8254 = n8250 & ~n8252 ;
  assign n8255 = ~n8253 & ~n8254 ;
  assign n8258 = n8255 & ~x26 ;
  assign n8259 = ~n8257 & ~n8258 ;
  assign n8260 = n2315 & n3632 ;
  assign n8261 = n372 & n8260 ;
  assign n8262 = n921 & n8261 ;
  assign n8263 = n2171 & n8262 ;
  assign n8264 = n1443 & n8263 ;
  assign n8265 = n710 & n8264 ;
  assign n8266 = n330 & n8265 ;
  assign n8267 = ~n292 & n8266 ;
  assign n8268 = ~n150 & n8267 ;
  assign n8269 = ~n345 & n8268 ;
  assign n8270 = ~n86 & n8269 ;
  assign n8271 = ~n233 & n8270 ;
  assign n8272 = ~n213 & n8271 ;
  assign n8273 = ~n8011 & ~n8105 ;
  assign n8274 = ~n8102 & ~n8273 ;
  assign n8275 = ~n8094 & ~n8098 ;
  assign n8276 = n3249 & n7700 ;
  assign n8277 = n3191 & n8016 ;
  assign n8278 = ~n8276 & ~n8277 ;
  assign n8279 = ~n266 & ~n8278 ;
  assign n8280 = ~n8278 & ~n8279 ;
  assign n8281 = ~n266 & ~n8279 ;
  assign n8282 = ~n8280 & ~n8281 ;
  assign n8283 = n2777 & ~n3255 ;
  assign n8284 = ~n2529 & n2783 ;
  assign n8285 = n2785 & n3252 ;
  assign n8286 = ~n8284 & ~n8285 ;
  assign n8287 = ~n8283 & n8286 ;
  assign n8288 = n2792 & n3293 ;
  assign n8289 = n8287 & ~n8288 ;
  assign n8290 = ~n996 & ~n8289 ;
  assign n8291 = ~n8289 & ~n8290 ;
  assign n8292 = ~n996 & ~n8290 ;
  assign n8293 = ~n8291 & ~n8292 ;
  assign n8294 = ~n8067 & ~n8071 ;
  assign n8295 = ~n500 & n8047 ;
  assign n8296 = n2568 & n8295 ;
  assign n8297 = ~n8052 & ~n8296 ;
  assign n8298 = n2553 & n2643 ;
  assign n8299 = ~n2561 & n2751 ;
  assign n8300 = ~n2557 & n2641 ;
  assign n8301 = ~n8299 & ~n8300 ;
  assign n8302 = ~n8298 & n8301 ;
  assign n8303 = n2649 & n2790 ;
  assign n8304 = n8302 & ~n8303 ;
  assign n8305 = ~n500 & n2565 ;
  assign n8306 = ~n8304 & n8305 ;
  assign n8307 = n8304 & ~n8305 ;
  assign n8308 = ~n8306 & ~n8307 ;
  assign n8309 = ~n8297 & n8308 ;
  assign n8310 = ~n8297 & ~n8309 ;
  assign n8311 = n8308 & ~n8309 ;
  assign n8312 = ~n8310 & ~n8311 ;
  assign n8313 = ~n2541 & n2674 ;
  assign n8314 = ~n2550 & n2670 ;
  assign n8315 = n2537 & n2672 ;
  assign n8316 = ~n8314 & ~n8315 ;
  assign n8317 = ~n8313 & n8316 ;
  assign n8318 = ~n2665 & n8317 ;
  assign n8319 = ~n2997 & n8317 ;
  assign n8320 = ~n8318 & ~n8319 ;
  assign n8321 = n644 & ~n8320 ;
  assign n8322 = ~n644 & n8320 ;
  assign n8323 = ~n8321 & ~n8322 ;
  assign n8324 = ~n8312 & n8323 ;
  assign n8325 = n8312 & ~n8323 ;
  assign n8326 = ~n8324 & ~n8325 ;
  assign n8327 = ~n8294 & n8326 ;
  assign n8328 = n8294 & ~n8326 ;
  assign n8329 = ~n8327 & ~n8328 ;
  assign n8330 = ~n8293 & n8329 ;
  assign n8331 = ~n8293 & ~n8330 ;
  assign n8332 = n8329 & ~n8330 ;
  assign n8333 = ~n8331 & ~n8332 ;
  assign n8334 = ~n8075 & ~n8081 ;
  assign n8335 = n8333 & n8334 ;
  assign n8336 = ~n8333 & ~n8334 ;
  assign n8337 = ~n8335 & ~n8336 ;
  assign n8338 = n270 & n3725 ;
  assign n8339 = n2535 & n3247 ;
  assign n8340 = n2542 & ~n3603 ;
  assign n8341 = ~n8339 & ~n8340 ;
  assign n8342 = ~n8338 & n8341 ;
  assign n8343 = ~n2546 & n8342 ;
  assign n8344 = ~n3737 & n8342 ;
  assign n8345 = ~n8343 & ~n8344 ;
  assign n8346 = n250 & ~n8345 ;
  assign n8347 = ~n250 & n8345 ;
  assign n8348 = ~n8346 & ~n8347 ;
  assign n8349 = n8337 & n8348 ;
  assign n8350 = ~n8337 & ~n8348 ;
  assign n8351 = ~n8349 & ~n8350 ;
  assign n8352 = ~n8282 & n8351 ;
  assign n8353 = n8282 & ~n8351 ;
  assign n8354 = ~n8352 & ~n8353 ;
  assign n8355 = ~n8275 & n8354 ;
  assign n8356 = n8275 & ~n8354 ;
  assign n8357 = ~n8355 & ~n8356 ;
  assign n8358 = ~n8274 & n8357 ;
  assign n8359 = n8274 & ~n8357 ;
  assign n8360 = ~n8358 & ~n8359 ;
  assign n8361 = ~n8272 & n8360 ;
  assign n8362 = ~n8272 & ~n8361 ;
  assign n8363 = n8360 & ~n8361 ;
  assign n8364 = ~n8362 & ~n8363 ;
  assign n8365 = ~n8114 & ~n8364 ;
  assign n8366 = n8114 & ~n8363 ;
  assign n8367 = ~n8362 & n8366 ;
  assign n8368 = ~n8365 & ~n8367 ;
  assign n8369 = n8118 & n8368 ;
  assign n8370 = n8368 & ~n8369 ;
  assign n8371 = n8118 & ~n8369 ;
  assign n8372 = ~n8370 & ~n8371 ;
  assign n8373 = ~n8119 & n8120 ;
  assign n8374 = ~n7831 & ~n8373 ;
  assign n8375 = ~n8372 & n8374 ;
  assign n8376 = n8372 & ~n8374 ;
  assign n8377 = ~n8375 & ~n8376 ;
  assign n8497 = n8377 & x27 ;
  assign n8378 = n6140 & n7457 ;
  assign n8379 = n4197 & n8378 ;
  assign n8380 = n4746 & n8379 ;
  assign n8381 = n5996 & n8380 ;
  assign n8382 = n5268 & n8381 ;
  assign n8383 = n4535 & n8382 ;
  assign n8384 = n4155 & n8383 ;
  assign n8385 = ~n4117 & n8384 ;
  assign n8386 = ~n3975 & n8385 ;
  assign n8387 = ~n4170 & n8386 ;
  assign n8388 = ~n3911 & n8387 ;
  assign n8389 = ~n4058 & n8388 ;
  assign n8390 = ~n4038 & n8389 ;
  assign n8391 = ~n8142 & ~n8236 ;
  assign n8392 = ~n8233 & ~n8391 ;
  assign n8393 = ~n8225 & ~n8229 ;
  assign n8394 = n7074 & n7857 ;
  assign n8395 = n7016 & n8147 ;
  assign n8396 = ~n8394 & ~n8395 ;
  assign n8397 = ~n4091 & ~n8396 ;
  assign n8398 = ~n8396 & ~n8397 ;
  assign n8399 = ~n4091 & ~n8397 ;
  assign n8400 = ~n8398 & ~n8399 ;
  assign n8401 = n6602 & ~n7080 ;
  assign n8402 = ~n6354 & n6608 ;
  assign n8403 = n6610 & n7077 ;
  assign n8404 = ~n8402 & ~n8403 ;
  assign n8405 = ~n8401 & n8404 ;
  assign n8406 = n6617 & n7118 ;
  assign n8407 = n8405 & ~n8406 ;
  assign n8408 = ~n4821 & ~n8407 ;
  assign n8409 = ~n8407 & ~n8408 ;
  assign n8410 = ~n4821 & ~n8408 ;
  assign n8411 = ~n8409 & ~n8410 ;
  assign n8412 = ~n8198 & ~n8202 ;
  assign n8413 = ~n4325 & n8178 ;
  assign n8414 = n6393 & n8413 ;
  assign n8415 = ~n8183 & ~n8414 ;
  assign n8416 = n6378 & n6468 ;
  assign n8417 = ~n6386 & n6576 ;
  assign n8418 = ~n6382 & n6466 ;
  assign n8419 = ~n8417 & ~n8418 ;
  assign n8420 = ~n8416 & n8419 ;
  assign n8421 = n6474 & n6615 ;
  assign n8422 = n8420 & ~n8421 ;
  assign n8423 = ~n4325 & n6390 ;
  assign n8424 = ~n8422 & n8423 ;
  assign n8425 = n8422 & ~n8423 ;
  assign n8426 = ~n8424 & ~n8425 ;
  assign n8427 = ~n8415 & n8426 ;
  assign n8428 = ~n8415 & ~n8427 ;
  assign n8429 = n8426 & ~n8427 ;
  assign n8430 = ~n8428 & ~n8429 ;
  assign n8431 = ~n6366 & n6499 ;
  assign n8432 = ~n6375 & n6495 ;
  assign n8433 = n6362 & n6497 ;
  assign n8434 = ~n8432 & ~n8433 ;
  assign n8435 = ~n8431 & n8434 ;
  assign n8436 = ~n6490 & n8435 ;
  assign n8437 = ~n6822 & n8435 ;
  assign n8438 = ~n8436 & ~n8437 ;
  assign n8439 = n4469 & ~n8438 ;
  assign n8440 = ~n4469 & n8438 ;
  assign n8441 = ~n8439 & ~n8440 ;
  assign n8442 = ~n8430 & n8441 ;
  assign n8443 = n8430 & ~n8441 ;
  assign n8444 = ~n8442 & ~n8443 ;
  assign n8445 = ~n8412 & n8444 ;
  assign n8446 = n8412 & ~n8444 ;
  assign n8447 = ~n8445 & ~n8446 ;
  assign n8448 = ~n8411 & n8447 ;
  assign n8449 = ~n8411 & ~n8448 ;
  assign n8450 = n8447 & ~n8448 ;
  assign n8451 = ~n8449 & ~n8450 ;
  assign n8452 = ~n8206 & ~n8212 ;
  assign n8453 = n8451 & n8452 ;
  assign n8454 = ~n8451 & ~n8452 ;
  assign n8455 = ~n8453 & ~n8454 ;
  assign n8456 = n4095 & n7550 ;
  assign n8457 = n6360 & n7072 ;
  assign n8458 = n6367 & ~n7428 ;
  assign n8459 = ~n8457 & ~n8458 ;
  assign n8460 = ~n8456 & n8459 ;
  assign n8461 = ~n6371 & n8460 ;
  assign n8462 = ~n7562 & n8460 ;
  assign n8463 = ~n8461 & ~n8462 ;
  assign n8464 = n4075 & ~n8463 ;
  assign n8465 = ~n4075 & n8463 ;
  assign n8466 = ~n8464 & ~n8465 ;
  assign n8467 = n8455 & n8466 ;
  assign n8468 = ~n8455 & ~n8466 ;
  assign n8469 = ~n8467 & ~n8468 ;
  assign n8470 = ~n8400 & n8469 ;
  assign n8471 = n8400 & ~n8469 ;
  assign n8472 = ~n8470 & ~n8471 ;
  assign n8473 = ~n8393 & n8472 ;
  assign n8474 = n8393 & ~n8472 ;
  assign n8475 = ~n8473 & ~n8474 ;
  assign n8476 = ~n8392 & n8475 ;
  assign n8477 = n8392 & ~n8475 ;
  assign n8478 = ~n8476 & ~n8477 ;
  assign n8479 = ~n8390 & n8478 ;
  assign n8480 = ~n8390 & ~n8479 ;
  assign n8481 = n8478 & ~n8479 ;
  assign n8482 = ~n8480 & ~n8481 ;
  assign n8483 = ~n8245 & ~n8482 ;
  assign n8484 = n8245 & ~n8481 ;
  assign n8485 = ~n8480 & n8484 ;
  assign n8486 = ~n8483 & ~n8485 ;
  assign n8487 = n8249 & n8486 ;
  assign n8488 = n8486 & ~n8487 ;
  assign n8489 = n8249 & ~n8487 ;
  assign n8490 = ~n8488 & ~n8489 ;
  assign n8491 = ~n8250 & n8251 ;
  assign n8492 = ~n7831 & ~n8491 ;
  assign n8493 = ~n8490 & n8492 ;
  assign n8494 = n8490 & ~n8492 ;
  assign n8495 = ~n8493 & ~n8494 ;
  assign n8498 = ~n8495 & ~x27 ;
  assign n8499 = ~n8497 & ~n8498 ;
  assign n8500 = ~n8361 & ~n8365 ;
  assign n8501 = n321 & n471 ;
  assign n8502 = n276 & n8501 ;
  assign n8503 = n2439 & n8502 ;
  assign n8504 = n950 & n8503 ;
  assign n8505 = n727 & n8504 ;
  assign n8506 = n619 & n8505 ;
  assign n8507 = n2393 & n8506 ;
  assign n8508 = ~n153 & n8507 ;
  assign n8509 = ~n169 & n8508 ;
  assign n8510 = ~n564 & n8509 ;
  assign n8511 = ~n8355 & ~n8358 ;
  assign n8512 = ~n8349 & ~n8352 ;
  assign n8513 = ~n8330 & ~n8336 ;
  assign n8514 = ~n8324 & ~n8327 ;
  assign n8515 = ~n2550 & n2643 ;
  assign n8516 = ~n2557 & n2751 ;
  assign n8517 = n2553 & n2641 ;
  assign n8518 = ~n8516 & ~n8517 ;
  assign n8519 = ~n8515 & n8518 ;
  assign n8520 = n2649 & n2964 ;
  assign n8521 = n8519 & ~n8520 ;
  assign n8522 = ~n500 & ~n8521 ;
  assign n8523 = ~n8521 & ~n8522 ;
  assign n8524 = ~n500 & ~n8522 ;
  assign n8525 = ~n8523 & ~n8524 ;
  assign n8526 = ~n266 & ~n500 ;
  assign n8527 = ~n2561 & n8526 ;
  assign n8528 = ~n266 & ~n8527 ;
  assign n8529 = ~n2561 & ~n8527 ;
  assign n8530 = ~n500 & n8529 ;
  assign n8531 = ~n8528 & ~n8530 ;
  assign n8532 = ~n8525 & ~n8531 ;
  assign n8533 = ~n8525 & ~n8532 ;
  assign n8534 = ~n8531 & ~n8532 ;
  assign n8535 = ~n8533 & ~n8534 ;
  assign n8536 = ~n500 & ~n2565 ;
  assign n8537 = n8304 & n8536 ;
  assign n8538 = ~n8309 & ~n8537 ;
  assign n8539 = n8535 & ~n8538 ;
  assign n8540 = ~n8535 & n8538 ;
  assign n8541 = ~n8539 & ~n8540 ;
  assign n8542 = ~n2529 & n2674 ;
  assign n8543 = n2537 & n2670 ;
  assign n8544 = ~n2541 & n2672 ;
  assign n8545 = ~n8543 & ~n8544 ;
  assign n8546 = ~n8542 & n8545 ;
  assign n8547 = n2627 & n2665 ;
  assign n8548 = n8546 & ~n8547 ;
  assign n8549 = ~n644 & ~n8548 ;
  assign n8550 = n644 & n8548 ;
  assign n8551 = ~n8549 & ~n8550 ;
  assign n8552 = ~n8541 & n8551 ;
  assign n8553 = ~n8541 & ~n8552 ;
  assign n8554 = n8551 & ~n8552 ;
  assign n8555 = ~n8553 & ~n8554 ;
  assign n8556 = ~n8514 & n8555 ;
  assign n8557 = n8514 & ~n8555 ;
  assign n8558 = ~n8556 & ~n8557 ;
  assign n8559 = n2777 & n3247 ;
  assign n8560 = n2783 & n3252 ;
  assign n8561 = n2785 & ~n3255 ;
  assign n8562 = ~n8560 & ~n8561 ;
  assign n8563 = ~n8559 & n8562 ;
  assign n8564 = n2792 & n3277 ;
  assign n8565 = n8563 & ~n8564 ;
  assign n8566 = ~n996 & ~n8565 ;
  assign n8567 = ~n996 & ~n8566 ;
  assign n8568 = ~n8565 & ~n8566 ;
  assign n8569 = ~n8567 & ~n8568 ;
  assign n8570 = ~n8558 & ~n8569 ;
  assign n8571 = n8558 & n8569 ;
  assign n8572 = ~n8570 & ~n8571 ;
  assign n8573 = ~n8513 & n8572 ;
  assign n8574 = n8513 & ~n8572 ;
  assign n8575 = ~n8573 & ~n8574 ;
  assign n8576 = n270 & n7700 ;
  assign n8577 = n2535 & ~n3603 ;
  assign n8578 = n2542 & n3725 ;
  assign n8579 = ~n8577 & ~n8578 ;
  assign n8580 = ~n8576 & n8579 ;
  assign n8581 = n2546 & n7712 ;
  assign n8582 = n8580 & ~n8581 ;
  assign n8583 = ~n250 & ~n8582 ;
  assign n8584 = n250 & n8582 ;
  assign n8585 = ~n8583 & ~n8584 ;
  assign n8586 = n8575 & n8585 ;
  assign n8587 = ~n8575 & ~n8585 ;
  assign n8588 = ~n8586 & ~n8587 ;
  assign n8589 = ~n8512 & n8588 ;
  assign n8590 = n8512 & ~n8588 ;
  assign n8591 = ~n8589 & ~n8590 ;
  assign n8592 = n8511 & ~n8591 ;
  assign n8593 = ~n8511 & n8591 ;
  assign n8594 = ~n8592 & ~n8593 ;
  assign n8595 = n8510 & ~n8594 ;
  assign n8596 = ~n8510 & n8594 ;
  assign n8597 = ~n8595 & ~n8596 ;
  assign n8598 = ~n8500 & n8597 ;
  assign n8599 = n8500 & ~n8597 ;
  assign n8600 = ~n8598 & ~n8599 ;
  assign n8601 = ~n8369 & ~n8600 ;
  assign n8602 = n8369 & n8600 ;
  assign n8603 = ~n8601 & ~n8602 ;
  assign n8604 = n8372 & n8373 ;
  assign n8605 = ~n7831 & ~n8604 ;
  assign n8606 = ~n8603 & n8605 ;
  assign n8607 = n8603 & ~n8605 ;
  assign n8608 = ~n8606 & ~n8607 ;
  assign n8719 = ~n8608 & x28 ;
  assign n8609 = ~n8479 & ~n8483 ;
  assign n8610 = n4146 & n4296 ;
  assign n8611 = n4101 & n8610 ;
  assign n8612 = n6264 & n8611 ;
  assign n8613 = n4775 & n8612 ;
  assign n8614 = n4552 & n8613 ;
  assign n8615 = n4444 & n8614 ;
  assign n8616 = n6218 & n8615 ;
  assign n8617 = ~n3978 & n8616 ;
  assign n8618 = ~n3994 & n8617 ;
  assign n8619 = ~n4389 & n8618 ;
  assign n8620 = ~n8473 & ~n8476 ;
  assign n8621 = ~n8467 & ~n8470 ;
  assign n8622 = ~n8448 & ~n8454 ;
  assign n8623 = ~n8442 & ~n8445 ;
  assign n8624 = ~n6375 & n6468 ;
  assign n8625 = ~n6382 & n6576 ;
  assign n8626 = n6378 & n6466 ;
  assign n8627 = ~n8625 & ~n8626 ;
  assign n8628 = ~n8624 & n8627 ;
  assign n8629 = n6474 & n6789 ;
  assign n8630 = n8628 & ~n8629 ;
  assign n8631 = ~n4325 & ~n8630 ;
  assign n8632 = ~n8630 & ~n8631 ;
  assign n8633 = ~n4325 & ~n8631 ;
  assign n8634 = ~n8632 & ~n8633 ;
  assign n8635 = ~n4091 & ~n4325 ;
  assign n8636 = ~n6386 & n8635 ;
  assign n8637 = ~n4091 & ~n8636 ;
  assign n8638 = ~n6386 & ~n8636 ;
  assign n8639 = ~n4325 & n8638 ;
  assign n8640 = ~n8637 & ~n8639 ;
  assign n8641 = ~n8634 & ~n8640 ;
  assign n8642 = ~n8634 & ~n8641 ;
  assign n8643 = ~n8640 & ~n8641 ;
  assign n8644 = ~n8642 & ~n8643 ;
  assign n8645 = ~n4325 & ~n6390 ;
  assign n8646 = n8422 & n8645 ;
  assign n8647 = ~n8427 & ~n8646 ;
  assign n8648 = n8644 & ~n8647 ;
  assign n8649 = ~n8644 & n8647 ;
  assign n8650 = ~n8648 & ~n8649 ;
  assign n8651 = ~n6354 & n6499 ;
  assign n8652 = n6362 & n6495 ;
  assign n8653 = ~n6366 & n6497 ;
  assign n8654 = ~n8652 & ~n8653 ;
  assign n8655 = ~n8651 & n8654 ;
  assign n8656 = n6452 & n6490 ;
  assign n8657 = n8655 & ~n8656 ;
  assign n8658 = ~n4469 & ~n8657 ;
  assign n8659 = n4469 & n8657 ;
  assign n8660 = ~n8658 & ~n8659 ;
  assign n8661 = ~n8650 & n8660 ;
  assign n8662 = ~n8650 & ~n8661 ;
  assign n8663 = n8660 & ~n8661 ;
  assign n8664 = ~n8662 & ~n8663 ;
  assign n8665 = ~n8623 & n8664 ;
  assign n8666 = n8623 & ~n8664 ;
  assign n8667 = ~n8665 & ~n8666 ;
  assign n8668 = n6602 & n7072 ;
  assign n8669 = n6608 & n7077 ;
  assign n8670 = n6610 & ~n7080 ;
  assign n8671 = ~n8669 & ~n8670 ;
  assign n8672 = ~n8668 & n8671 ;
  assign n8673 = n6617 & n7102 ;
  assign n8674 = n8672 & ~n8673 ;
  assign n8675 = ~n4821 & ~n8674 ;
  assign n8676 = ~n4821 & ~n8675 ;
  assign n8677 = ~n8674 & ~n8675 ;
  assign n8678 = ~n8676 & ~n8677 ;
  assign n8679 = ~n8667 & ~n8678 ;
  assign n8680 = n8667 & n8678 ;
  assign n8681 = ~n8679 & ~n8680 ;
  assign n8682 = ~n8622 & n8681 ;
  assign n8683 = n8622 & ~n8681 ;
  assign n8684 = ~n8682 & ~n8683 ;
  assign n8685 = n4095 & n7857 ;
  assign n8686 = n6360 & ~n7428 ;
  assign n8687 = n6367 & n7550 ;
  assign n8688 = ~n8686 & ~n8687 ;
  assign n8689 = ~n8685 & n8688 ;
  assign n8690 = n6371 & n7869 ;
  assign n8691 = n8689 & ~n8690 ;
  assign n8692 = ~n4075 & ~n8691 ;
  assign n8693 = n4075 & n8691 ;
  assign n8694 = ~n8692 & ~n8693 ;
  assign n8695 = n8684 & n8694 ;
  assign n8696 = ~n8684 & ~n8694 ;
  assign n8697 = ~n8695 & ~n8696 ;
  assign n8698 = ~n8621 & n8697 ;
  assign n8699 = n8621 & ~n8697 ;
  assign n8700 = ~n8698 & ~n8699 ;
  assign n8701 = n8620 & ~n8700 ;
  assign n8702 = ~n8620 & n8700 ;
  assign n8703 = ~n8701 & ~n8702 ;
  assign n8704 = n8619 & ~n8703 ;
  assign n8705 = ~n8619 & n8703 ;
  assign n8706 = ~n8704 & ~n8705 ;
  assign n8707 = ~n8609 & n8706 ;
  assign n8708 = n8609 & ~n8706 ;
  assign n8709 = ~n8707 & ~n8708 ;
  assign n8710 = ~n8487 & ~n8709 ;
  assign n8711 = n8487 & n8709 ;
  assign n8712 = ~n8710 & ~n8711 ;
  assign n8713 = n8490 & n8491 ;
  assign n8714 = ~n7831 & ~n8713 ;
  assign n8715 = ~n8712 & n8714 ;
  assign n8716 = n8712 & ~n8714 ;
  assign n8717 = ~n8715 & ~n8716 ;
  assign n8720 = n8717 & ~x28 ;
  assign n8721 = ~n8719 & ~n8720 ;
  assign n8722 = ~n8596 & ~n8598 ;
  assign n8723 = ~n292 & ~n334 ;
  assign n8724 = ~n447 & n8723 ;
  assign n8725 = n164 & n782 ;
  assign n8726 = n8724 & n8725 ;
  assign n8727 = n2292 & n8726 ;
  assign n8728 = n289 & n8727 ;
  assign n8729 = n7687 & n8728 ;
  assign n8730 = n3218 & n8729 ;
  assign n8731 = n7806 & n8730 ;
  assign n8732 = n344 & n8731 ;
  assign n8733 = ~n153 & n8732 ;
  assign n8734 = ~n392 & n8733 ;
  assign n8735 = ~n274 & n8734 ;
  assign n8736 = ~n212 & n8735 ;
  assign n8737 = ~n8589 & ~n8593 ;
  assign n8738 = ~n8573 & ~n8586 ;
  assign n8739 = ~n8514 & ~n8555 ;
  assign n8740 = ~n8570 & ~n8739 ;
  assign n8741 = n2777 & ~n3603 ;
  assign n8742 = n2783 & ~n3255 ;
  assign n8743 = n2785 & n3247 ;
  assign n8744 = ~n8742 & ~n8743 ;
  assign n8745 = ~n8741 & n8744 ;
  assign n8746 = n2792 & n3616 ;
  assign n8747 = n8745 & ~n8746 ;
  assign n8748 = ~n996 & ~n8747 ;
  assign n8749 = ~n8747 & ~n8748 ;
  assign n8750 = ~n996 & ~n8748 ;
  assign n8751 = ~n8749 & ~n8750 ;
  assign n8752 = ~n8535 & ~n8538 ;
  assign n8753 = ~n8552 & ~n8752 ;
  assign n8754 = ~n8527 & ~n8532 ;
  assign n8755 = ~n2557 & n8526 ;
  assign n8756 = ~n266 & ~n8755 ;
  assign n8757 = ~n2557 & ~n8755 ;
  assign n8758 = ~n500 & n8757 ;
  assign n8759 = ~n8756 & ~n8758 ;
  assign n8760 = ~n8754 & ~n8759 ;
  assign n8761 = ~n8754 & ~n8760 ;
  assign n8762 = ~n8759 & ~n8760 ;
  assign n8763 = ~n8761 & ~n8762 ;
  assign n8764 = n2537 & n2643 ;
  assign n8765 = n2553 & n2751 ;
  assign n8766 = ~n2550 & n2641 ;
  assign n8767 = ~n8765 & ~n8766 ;
  assign n8768 = ~n8764 & n8767 ;
  assign n8769 = ~n2649 & n8768 ;
  assign n8770 = ~n3017 & n8768 ;
  assign n8771 = ~n8769 & ~n8770 ;
  assign n8772 = n500 & ~n8771 ;
  assign n8773 = ~n500 & n8771 ;
  assign n8774 = ~n8772 & ~n8773 ;
  assign n8775 = ~n8763 & n8774 ;
  assign n8776 = ~n8763 & ~n8775 ;
  assign n8777 = n8774 & ~n8775 ;
  assign n8778 = ~n8776 & ~n8777 ;
  assign n8779 = n2674 & n3252 ;
  assign n8780 = ~n2541 & n2670 ;
  assign n8781 = ~n2529 & n2672 ;
  assign n8782 = ~n8780 & ~n8781 ;
  assign n8783 = ~n8779 & n8782 ;
  assign n8784 = n2665 & n3307 ;
  assign n8785 = n8783 & ~n8784 ;
  assign n8786 = ~n644 & ~n8785 ;
  assign n8787 = n644 & n8785 ;
  assign n8788 = ~n8786 & ~n8787 ;
  assign n8789 = ~n8778 & n8788 ;
  assign n8790 = ~n8777 & ~n8788 ;
  assign n8791 = ~n8776 & n8790 ;
  assign n8792 = ~n8789 & ~n8791 ;
  assign n8793 = ~n8753 & n8792 ;
  assign n8794 = ~n8753 & ~n8793 ;
  assign n8795 = n8792 & ~n8793 ;
  assign n8796 = ~n8794 & ~n8795 ;
  assign n8797 = ~n8751 & ~n8796 ;
  assign n8798 = n8751 & ~n8795 ;
  assign n8799 = ~n8794 & n8798 ;
  assign n8800 = ~n8797 & ~n8799 ;
  assign n8801 = ~n8740 & n8800 ;
  assign n8802 = ~n8740 & ~n8801 ;
  assign n8803 = n8800 & ~n8801 ;
  assign n8804 = ~n8802 & ~n8803 ;
  assign n8805 = n2535 & n3725 ;
  assign n8806 = n2542 & n7700 ;
  assign n8807 = ~n8805 & ~n8806 ;
  assign n8808 = n2546 & n8018 ;
  assign n8809 = n8807 & ~n8808 ;
  assign n8810 = ~n250 & ~n8809 ;
  assign n8811 = n250 & n8809 ;
  assign n8812 = ~n8810 & ~n8811 ;
  assign n8813 = ~n8804 & n8812 ;
  assign n8814 = ~n8803 & ~n8812 ;
  assign n8815 = ~n8802 & n8814 ;
  assign n8816 = ~n8813 & ~n8815 ;
  assign n8817 = ~n8738 & n8816 ;
  assign n8818 = n8738 & ~n8816 ;
  assign n8819 = ~n8817 & ~n8818 ;
  assign n8820 = ~n8737 & n8819 ;
  assign n8821 = n8737 & ~n8819 ;
  assign n8822 = ~n8820 & ~n8821 ;
  assign n8823 = n8736 & ~n8822 ;
  assign n8824 = ~n8736 & n8822 ;
  assign n8825 = ~n8823 & ~n8824 ;
  assign n8826 = ~n8722 & n8825 ;
  assign n8827 = n8722 & ~n8825 ;
  assign n8828 = ~n8826 & ~n8827 ;
  assign n8829 = ~n8602 & ~n8828 ;
  assign n8830 = n8602 & n8828 ;
  assign n8831 = ~n8829 & ~n8830 ;
  assign n8832 = ~n8603 & n8604 ;
  assign n8833 = ~n7831 & ~n8832 ;
  assign n8834 = ~n8831 & n8833 ;
  assign n8835 = n8831 & ~n8833 ;
  assign n8836 = ~n8834 & ~n8835 ;
  assign n8953 = ~n8836 & x29 ;
  assign n8837 = ~n8705 & ~n8707 ;
  assign n8838 = ~n4117 & ~n4159 ;
  assign n8839 = ~n4272 & n8838 ;
  assign n8840 = n3989 & n4607 ;
  assign n8841 = n8839 & n8840 ;
  assign n8842 = n6117 & n8841 ;
  assign n8843 = n4114 & n8842 ;
  assign n8844 = n7844 & n8843 ;
  assign n8845 = n7043 & n8844 ;
  assign n8846 = n7963 & n8845 ;
  assign n8847 = n4169 & n8846 ;
  assign n8848 = ~n3978 & n8847 ;
  assign n8849 = ~n4217 & n8848 ;
  assign n8850 = ~n4099 & n8849 ;
  assign n8851 = ~n4037 & n8850 ;
  assign n8852 = ~n8698 & ~n8702 ;
  assign n8853 = ~n8682 & ~n8695 ;
  assign n8854 = ~n8623 & ~n8664 ;
  assign n8855 = ~n8679 & ~n8854 ;
  assign n8856 = n6602 & ~n7428 ;
  assign n8857 = n6608 & ~n7080 ;
  assign n8858 = n6610 & n7072 ;
  assign n8859 = ~n8857 & ~n8858 ;
  assign n8860 = ~n8856 & n8859 ;
  assign n8861 = n6617 & n7441 ;
  assign n8862 = n8860 & ~n8861 ;
  assign n8863 = ~n4821 & ~n8862 ;
  assign n8864 = ~n8862 & ~n8863 ;
  assign n8865 = ~n4821 & ~n8863 ;
  assign n8866 = ~n8864 & ~n8865 ;
  assign n8867 = ~n8644 & ~n8647 ;
  assign n8868 = ~n8661 & ~n8867 ;
  assign n8869 = ~n8636 & ~n8641 ;
  assign n8870 = ~n6382 & n8635 ;
  assign n8871 = ~n4091 & ~n8870 ;
  assign n8872 = ~n6382 & ~n8870 ;
  assign n8873 = ~n4325 & n8872 ;
  assign n8874 = ~n8871 & ~n8873 ;
  assign n8875 = ~n8869 & ~n8874 ;
  assign n8876 = ~n8869 & ~n8875 ;
  assign n8877 = ~n8874 & ~n8875 ;
  assign n8878 = ~n8876 & ~n8877 ;
  assign n8879 = n6362 & n6468 ;
  assign n8880 = n6378 & n6576 ;
  assign n8881 = ~n6375 & n6466 ;
  assign n8882 = ~n8880 & ~n8881 ;
  assign n8883 = ~n8879 & n8882 ;
  assign n8884 = ~n6474 & n8883 ;
  assign n8885 = ~n6842 & n8883 ;
  assign n8886 = ~n8884 & ~n8885 ;
  assign n8887 = n4325 & ~n8886 ;
  assign n8888 = ~n4325 & n8886 ;
  assign n8889 = ~n8887 & ~n8888 ;
  assign n8890 = ~n8878 & n8889 ;
  assign n8891 = ~n8878 & ~n8890 ;
  assign n8892 = n8889 & ~n8890 ;
  assign n8893 = ~n8891 & ~n8892 ;
  assign n8894 = n6499 & n7077 ;
  assign n8895 = ~n6366 & n6495 ;
  assign n8896 = ~n6354 & n6497 ;
  assign n8897 = ~n8895 & ~n8896 ;
  assign n8898 = ~n8894 & n8897 ;
  assign n8899 = n6490 & n7132 ;
  assign n8900 = n8898 & ~n8899 ;
  assign n8901 = ~n4469 & ~n8900 ;
  assign n8902 = n4469 & n8900 ;
  assign n8903 = ~n8901 & ~n8902 ;
  assign n8904 = ~n8893 & n8903 ;
  assign n8905 = ~n8892 & ~n8903 ;
  assign n8906 = ~n8891 & n8905 ;
  assign n8907 = ~n8904 & ~n8906 ;
  assign n8908 = ~n8868 & n8907 ;
  assign n8909 = ~n8868 & ~n8908 ;
  assign n8910 = n8907 & ~n8908 ;
  assign n8911 = ~n8909 & ~n8910 ;
  assign n8912 = ~n8866 & ~n8911 ;
  assign n8913 = n8866 & ~n8910 ;
  assign n8914 = ~n8909 & n8913 ;
  assign n8915 = ~n8912 & ~n8914 ;
  assign n8916 = ~n8855 & n8915 ;
  assign n8917 = ~n8855 & ~n8916 ;
  assign n8918 = n8915 & ~n8916 ;
  assign n8919 = ~n8917 & ~n8918 ;
  assign n8920 = n6360 & n7550 ;
  assign n8921 = n6367 & n7857 ;
  assign n8922 = ~n8920 & ~n8921 ;
  assign n8923 = n6371 & n8149 ;
  assign n8924 = n8922 & ~n8923 ;
  assign n8925 = ~n4075 & ~n8924 ;
  assign n8926 = n4075 & n8924 ;
  assign n8927 = ~n8925 & ~n8926 ;
  assign n8928 = ~n8919 & n8927 ;
  assign n8929 = ~n8918 & ~n8927 ;
  assign n8930 = ~n8917 & n8929 ;
  assign n8931 = ~n8928 & ~n8930 ;
  assign n8932 = ~n8853 & n8931 ;
  assign n8933 = n8853 & ~n8931 ;
  assign n8934 = ~n8932 & ~n8933 ;
  assign n8935 = ~n8852 & n8934 ;
  assign n8936 = n8852 & ~n8934 ;
  assign n8937 = ~n8935 & ~n8936 ;
  assign n8938 = n8851 & ~n8937 ;
  assign n8939 = ~n8851 & n8937 ;
  assign n8940 = ~n8938 & ~n8939 ;
  assign n8941 = ~n8837 & n8940 ;
  assign n8942 = n8837 & ~n8940 ;
  assign n8943 = ~n8941 & ~n8942 ;
  assign n8944 = ~n8711 & ~n8943 ;
  assign n8945 = n8711 & n8943 ;
  assign n8946 = ~n8944 & ~n8945 ;
  assign n8947 = ~n8712 & n8713 ;
  assign n8948 = ~n7831 & ~n8947 ;
  assign n8949 = ~n8946 & n8948 ;
  assign n8950 = n8946 & ~n8948 ;
  assign n8951 = ~n8949 & ~n8950 ;
  assign n8954 = n8951 & ~x29 ;
  assign n8955 = ~n8953 & ~n8954 ;
  assign n8956 = ~n8824 & ~n8826 ;
  assign n8957 = n291 & n1092 ;
  assign n8958 = n561 & n8957 ;
  assign n8959 = n2396 & n8958 ;
  assign n8960 = n2315 & n8959 ;
  assign n8961 = n131 & n8960 ;
  assign n8962 = n344 & n8961 ;
  assign n8963 = n951 & n8962 ;
  assign n8964 = ~n332 & n8963 ;
  assign n8965 = n228 & n945 ;
  assign n8966 = n2433 & n8965 ;
  assign n8967 = n3234 & n8966 ;
  assign n8968 = n8964 & n8967 ;
  assign n8969 = ~n312 & n8968 ;
  assign n8970 = ~n125 & n8969 ;
  assign n8971 = ~n147 & n8970 ;
  assign n8972 = ~n144 & n8971 ;
  assign n8973 = ~n422 & n8972 ;
  assign n8974 = ~n123 & n8973 ;
  assign n8975 = ~n8817 & ~n8820 ;
  assign n8976 = ~n8801 & ~n8813 ;
  assign n8977 = ~n8793 & ~n8797 ;
  assign n8978 = n2535 & n7700 ;
  assign n8979 = n2546 & n8016 ;
  assign n8980 = ~n8978 & ~n8979 ;
  assign n8981 = n250 & ~n8980 ;
  assign n8982 = ~n250 & n8980 ;
  assign n8983 = ~n8981 & ~n8982 ;
  assign n8984 = ~n8977 & ~n8983 ;
  assign n8985 = n8977 & n8983 ;
  assign n8986 = ~n8984 & ~n8985 ;
  assign n8987 = n2777 & n3725 ;
  assign n8988 = n2783 & n3247 ;
  assign n8989 = n2785 & ~n3603 ;
  assign n8990 = ~n8988 & ~n8989 ;
  assign n8991 = ~n8987 & n8990 ;
  assign n8992 = n2792 & n3737 ;
  assign n8993 = n8991 & ~n8992 ;
  assign n8994 = ~n996 & ~n8993 ;
  assign n8995 = ~n8993 & ~n8994 ;
  assign n8996 = ~n996 & ~n8994 ;
  assign n8997 = ~n8995 & ~n8996 ;
  assign n8998 = ~n8775 & ~n8789 ;
  assign n8999 = ~n8755 & ~n8760 ;
  assign n9000 = n2553 & n8526 ;
  assign n9001 = ~n266 & ~n9000 ;
  assign n9002 = n2553 & ~n9000 ;
  assign n9003 = ~n500 & n9002 ;
  assign n9004 = ~n9001 & ~n9003 ;
  assign n9005 = ~n8999 & ~n9004 ;
  assign n9006 = ~n8999 & ~n9005 ;
  assign n9007 = ~n9004 & ~n9005 ;
  assign n9008 = ~n9006 & ~n9007 ;
  assign n9009 = ~n2541 & n2643 ;
  assign n9010 = ~n2550 & n2751 ;
  assign n9011 = n2537 & n2641 ;
  assign n9012 = ~n9010 & ~n9011 ;
  assign n9013 = ~n9009 & n9012 ;
  assign n9014 = ~n2649 & n9013 ;
  assign n9015 = ~n2997 & n9013 ;
  assign n9016 = ~n9014 & ~n9015 ;
  assign n9017 = n500 & ~n9016 ;
  assign n9018 = ~n500 & n9016 ;
  assign n9019 = ~n9017 & ~n9018 ;
  assign n9020 = ~n9008 & n9019 ;
  assign n9021 = ~n9008 & ~n9020 ;
  assign n9022 = n9019 & ~n9020 ;
  assign n9023 = ~n9021 & ~n9022 ;
  assign n9024 = n2674 & ~n3255 ;
  assign n9025 = ~n2529 & n2670 ;
  assign n9026 = n2672 & n3252 ;
  assign n9027 = ~n9025 & ~n9026 ;
  assign n9028 = ~n9024 & n9027 ;
  assign n9029 = n2665 & n3293 ;
  assign n9030 = n9028 & ~n9029 ;
  assign n9031 = ~n644 & ~n9030 ;
  assign n9032 = n644 & n9030 ;
  assign n9033 = ~n9031 & ~n9032 ;
  assign n9034 = ~n9023 & n9033 ;
  assign n9035 = ~n9022 & ~n9033 ;
  assign n9036 = ~n9021 & n9035 ;
  assign n9037 = ~n9034 & ~n9036 ;
  assign n9038 = ~n8998 & n9037 ;
  assign n9039 = ~n8998 & ~n9038 ;
  assign n9040 = n9037 & ~n9038 ;
  assign n9041 = ~n9039 & ~n9040 ;
  assign n9042 = ~n8997 & ~n9041 ;
  assign n9043 = n8997 & ~n9040 ;
  assign n9044 = ~n9039 & n9043 ;
  assign n9045 = ~n9042 & ~n9044 ;
  assign n9046 = n8986 & n9045 ;
  assign n9047 = ~n8986 & ~n9045 ;
  assign n9048 = ~n9046 & ~n9047 ;
  assign n9049 = ~n8976 & n9048 ;
  assign n9050 = n8976 & ~n9048 ;
  assign n9051 = ~n9049 & ~n9050 ;
  assign n9052 = ~n8975 & n9051 ;
  assign n9053 = n8975 & ~n9051 ;
  assign n9054 = ~n9052 & ~n9053 ;
  assign n9055 = n8974 & ~n9054 ;
  assign n9056 = ~n8974 & n9054 ;
  assign n9057 = ~n9055 & ~n9056 ;
  assign n9058 = ~n8956 & n9057 ;
  assign n9059 = n8956 & ~n9057 ;
  assign n9060 = ~n9058 & ~n9059 ;
  assign n9061 = ~n8830 & ~n9060 ;
  assign n9062 = n8830 & n9060 ;
  assign n9063 = ~n9061 & ~n9062 ;
  assign n9064 = ~n8831 & n8832 ;
  assign n9065 = ~n7831 & ~n9064 ;
  assign n9066 = ~n9063 & n9065 ;
  assign n9067 = n9063 & ~n9065 ;
  assign n9068 = ~n9066 & ~n9067 ;
  assign n9183 = ~n9068 & x30 ;
  assign n9069 = ~n8939 & ~n8941 ;
  assign n9070 = n4116 & n4917 ;
  assign n9071 = n4386 & n9070 ;
  assign n9072 = n6221 & n9071 ;
  assign n9073 = n6140 & n9072 ;
  assign n9074 = n3956 & n9073 ;
  assign n9075 = n4169 & n9074 ;
  assign n9076 = n4776 & n9075 ;
  assign n9077 = ~n4157 & n9076 ;
  assign n9078 = n4053 & n4770 ;
  assign n9079 = n6258 & n9078 ;
  assign n9080 = n7059 & n9079 ;
  assign n9081 = n9077 & n9080 ;
  assign n9082 = ~n4137 & n9081 ;
  assign n9083 = ~n3950 & n9082 ;
  assign n9084 = ~n3972 & n9083 ;
  assign n9085 = ~n3969 & n9084 ;
  assign n9086 = ~n4247 & n9085 ;
  assign n9087 = ~n3948 & n9086 ;
  assign n9088 = ~n8932 & ~n8935 ;
  assign n9089 = ~n8916 & ~n8928 ;
  assign n9090 = ~n8908 & ~n8912 ;
  assign n9091 = n6360 & n7857 ;
  assign n9092 = n6371 & n8147 ;
  assign n9093 = ~n9091 & ~n9092 ;
  assign n9094 = n4075 & ~n9093 ;
  assign n9095 = ~n4075 & n9093 ;
  assign n9096 = ~n9094 & ~n9095 ;
  assign n9097 = ~n9090 & ~n9096 ;
  assign n9098 = n9090 & n9096 ;
  assign n9099 = ~n9097 & ~n9098 ;
  assign n9100 = n6602 & n7550 ;
  assign n9101 = n6608 & n7072 ;
  assign n9102 = n6610 & ~n7428 ;
  assign n9103 = ~n9101 & ~n9102 ;
  assign n9104 = ~n9100 & n9103 ;
  assign n9105 = n6617 & n7562 ;
  assign n9106 = n9104 & ~n9105 ;
  assign n9107 = ~n4821 & ~n9106 ;
  assign n9108 = ~n9106 & ~n9107 ;
  assign n9109 = ~n4821 & ~n9107 ;
  assign n9110 = ~n9108 & ~n9109 ;
  assign n9111 = ~n8890 & ~n8904 ;
  assign n9112 = ~n8870 & ~n8875 ;
  assign n9113 = n6378 & n8635 ;
  assign n9114 = ~n4091 & ~n9113 ;
  assign n9115 = n6378 & ~n9113 ;
  assign n9116 = ~n4325 & n9115 ;
  assign n9117 = ~n9114 & ~n9116 ;
  assign n9118 = ~n9112 & ~n9117 ;
  assign n9119 = ~n9112 & ~n9118 ;
  assign n9120 = ~n9117 & ~n9118 ;
  assign n9121 = ~n9119 & ~n9120 ;
  assign n9122 = ~n6366 & n6468 ;
  assign n9123 = ~n6375 & n6576 ;
  assign n9124 = n6362 & n6466 ;
  assign n9125 = ~n9123 & ~n9124 ;
  assign n9126 = ~n9122 & n9125 ;
  assign n9127 = ~n6474 & n9126 ;
  assign n9128 = ~n6822 & n9126 ;
  assign n9129 = ~n9127 & ~n9128 ;
  assign n9130 = n4325 & ~n9129 ;
  assign n9131 = ~n4325 & n9129 ;
  assign n9132 = ~n9130 & ~n9131 ;
  assign n9133 = ~n9121 & n9132 ;
  assign n9134 = ~n9121 & ~n9133 ;
  assign n9135 = n9132 & ~n9133 ;
  assign n9136 = ~n9134 & ~n9135 ;
  assign n9137 = n6499 & ~n7080 ;
  assign n9138 = ~n6354 & n6495 ;
  assign n9139 = n6497 & n7077 ;
  assign n9140 = ~n9138 & ~n9139 ;
  assign n9141 = ~n9137 & n9140 ;
  assign n9142 = n6490 & n7118 ;
  assign n9143 = n9141 & ~n9142 ;
  assign n9144 = ~n4469 & ~n9143 ;
  assign n9145 = n4469 & n9143 ;
  assign n9146 = ~n9144 & ~n9145 ;
  assign n9147 = ~n9136 & n9146 ;
  assign n9148 = ~n9135 & ~n9146 ;
  assign n9149 = ~n9134 & n9148 ;
  assign n9150 = ~n9147 & ~n9149 ;
  assign n9151 = ~n9111 & n9150 ;
  assign n9152 = ~n9111 & ~n9151 ;
  assign n9153 = n9150 & ~n9151 ;
  assign n9154 = ~n9152 & ~n9153 ;
  assign n9155 = ~n9110 & ~n9154 ;
  assign n9156 = n9110 & ~n9153 ;
  assign n9157 = ~n9152 & n9156 ;
  assign n9158 = ~n9155 & ~n9157 ;
  assign n9159 = n9099 & n9158 ;
  assign n9160 = ~n9099 & ~n9158 ;
  assign n9161 = ~n9159 & ~n9160 ;
  assign n9162 = ~n9089 & n9161 ;
  assign n9163 = n9089 & ~n9161 ;
  assign n9164 = ~n9162 & ~n9163 ;
  assign n9165 = ~n9088 & n9164 ;
  assign n9166 = n9088 & ~n9164 ;
  assign n9167 = ~n9165 & ~n9166 ;
  assign n9168 = n9087 & ~n9167 ;
  assign n9169 = ~n9087 & n9167 ;
  assign n9170 = ~n9168 & ~n9169 ;
  assign n9171 = ~n9069 & n9170 ;
  assign n9172 = n9069 & ~n9170 ;
  assign n9173 = ~n9171 & ~n9172 ;
  assign n9174 = ~n8945 & ~n9173 ;
  assign n9175 = n8945 & n9173 ;
  assign n9176 = ~n9174 & ~n9175 ;
  assign n9177 = ~n8946 & n8947 ;
  assign n9178 = ~n7831 & ~n9177 ;
  assign n9179 = ~n9176 & n9178 ;
  assign n9180 = n9176 & ~n9178 ;
  assign n9181 = ~n9179 & ~n9180 ;
  assign n9184 = n9181 & ~x30 ;
  assign n9185 = ~n9183 & ~n9184 ;
  assign n9186 = ~n9056 & ~n9058 ;
  assign n9187 = ~n8984 & ~n9046 ;
  assign n9188 = ~n9038 & ~n9042 ;
  assign n9189 = n2777 & n7700 ;
  assign n9190 = n2783 & ~n3603 ;
  assign n9191 = n2785 & n3725 ;
  assign n9192 = ~n9190 & ~n9191 ;
  assign n9193 = ~n9189 & n9192 ;
  assign n9194 = ~n7712 & n9193 ;
  assign n9195 = ~n2792 & n9193 ;
  assign n9196 = ~n9194 & ~n9195 ;
  assign n9197 = n996 & ~n9196 ;
  assign n9198 = ~n996 & n9196 ;
  assign n9199 = ~n9197 & ~n9198 ;
  assign n9200 = ~n9188 & n9199 ;
  assign n9201 = n9188 & ~n9199 ;
  assign n9202 = ~n9200 & ~n9201 ;
  assign n9203 = ~n9020 & ~n9034 ;
  assign n9204 = ~n9000 & ~n9005 ;
  assign n9205 = ~n2529 & n2643 ;
  assign n9206 = n2537 & n2751 ;
  assign n9207 = ~n2541 & n2641 ;
  assign n9208 = ~n9206 & ~n9207 ;
  assign n9209 = ~n9205 & n9208 ;
  assign n9210 = n2627 & n2649 ;
  assign n9211 = n9209 & ~n9210 ;
  assign n9212 = ~n500 & ~n9211 ;
  assign n9213 = ~n9211 & ~n9212 ;
  assign n9214 = ~n500 & ~n9212 ;
  assign n9215 = ~n9213 & ~n9214 ;
  assign n9216 = ~n500 & ~n2550 ;
  assign n9217 = n250 & n266 ;
  assign n9218 = ~n250 & ~n266 ;
  assign n9219 = ~n9217 & ~n9218 ;
  assign n9220 = n9216 & n9219 ;
  assign n9221 = ~n9216 & ~n9219 ;
  assign n9222 = ~n9220 & ~n9221 ;
  assign n9223 = ~n9215 & n9222 ;
  assign n9224 = ~n9215 & ~n9223 ;
  assign n9225 = n9222 & ~n9223 ;
  assign n9226 = ~n9224 & ~n9225 ;
  assign n9227 = ~n9204 & n9226 ;
  assign n9228 = n9204 & ~n9226 ;
  assign n9229 = ~n9227 & ~n9228 ;
  assign n9230 = n2674 & n3247 ;
  assign n9231 = n2670 & n3252 ;
  assign n9232 = n2672 & ~n3255 ;
  assign n9233 = ~n9231 & ~n9232 ;
  assign n9234 = ~n9230 & n9233 ;
  assign n9235 = ~n2665 & n9234 ;
  assign n9236 = ~n3277 & n9234 ;
  assign n9237 = ~n9235 & ~n9236 ;
  assign n9238 = n644 & ~n9237 ;
  assign n9239 = ~n644 & n9237 ;
  assign n9240 = ~n9238 & ~n9239 ;
  assign n9241 = ~n9229 & n9240 ;
  assign n9242 = ~n9229 & ~n9241 ;
  assign n9243 = n9240 & ~n9241 ;
  assign n9244 = ~n9242 & ~n9243 ;
  assign n9245 = ~n9203 & ~n9244 ;
  assign n9246 = ~n9203 & ~n9245 ;
  assign n9247 = ~n9244 & ~n9245 ;
  assign n9248 = ~n9246 & ~n9247 ;
  assign n9249 = n9202 & ~n9248 ;
  assign n9250 = n9202 & ~n9249 ;
  assign n9251 = ~n9248 & ~n9249 ;
  assign n9252 = ~n9250 & ~n9251 ;
  assign n9253 = ~n9187 & n9252 ;
  assign n9254 = n9187 & ~n9252 ;
  assign n9255 = ~n9253 & ~n9254 ;
  assign n9256 = ~n9049 & ~n9052 ;
  assign n9257 = n9255 & n9256 ;
  assign n9258 = ~n9255 & ~n9256 ;
  assign n9259 = ~n9257 & ~n9258 ;
  assign n9260 = n906 & n2256 ;
  assign n9261 = n8724 & n9260 ;
  assign n9262 = n784 & n9261 ;
  assign n9263 = n8964 & n9262 ;
  assign n9264 = ~n104 & n9263 ;
  assign n9265 = ~n169 & n9264 ;
  assign n9266 = ~n112 & n9265 ;
  assign n9267 = ~n193 & n9266 ;
  assign n9268 = n1065 & n9267 ;
  assign n9269 = ~n143 & n9268 ;
  assign n9270 = ~n420 & n9269 ;
  assign n9271 = n9259 & ~n9270 ;
  assign n9272 = ~n9259 & n9270 ;
  assign n9273 = ~n9271 & ~n9272 ;
  assign n9274 = ~n9186 & n9273 ;
  assign n9275 = n9186 & ~n9273 ;
  assign n9276 = ~n9274 & ~n9275 ;
  assign n9277 = n9062 & n9276 ;
  assign n9278 = ~n9062 & ~n9276 ;
  assign n9279 = ~n9277 & ~n9278 ;
  assign n9280 = ~n9063 & n9064 ;
  assign n9281 = ~n7831 & ~n9280 ;
  assign n9282 = ~n9279 & n9281 ;
  assign n9283 = n9279 & ~n9281 ;
  assign n9284 = ~n9282 & ~n9283 ;
  assign n9385 = ~n9284 & x31 ;
  assign n9285 = ~n9169 & ~n9171 ;
  assign n9286 = ~n9097 & ~n9159 ;
  assign n9287 = ~n9151 & ~n9155 ;
  assign n9288 = n6602 & n7857 ;
  assign n9289 = n6608 & ~n7428 ;
  assign n9290 = n6610 & n7550 ;
  assign n9291 = ~n9289 & ~n9290 ;
  assign n9292 = ~n9288 & n9291 ;
  assign n9293 = ~n7869 & n9292 ;
  assign n9294 = ~n6617 & n9292 ;
  assign n9295 = ~n9293 & ~n9294 ;
  assign n9296 = n4821 & ~n9295 ;
  assign n9297 = ~n4821 & n9295 ;
  assign n9298 = ~n9296 & ~n9297 ;
  assign n9299 = ~n9287 & n9298 ;
  assign n9300 = n9287 & ~n9298 ;
  assign n9301 = ~n9299 & ~n9300 ;
  assign n9302 = ~n9133 & ~n9147 ;
  assign n9303 = ~n9113 & ~n9118 ;
  assign n9304 = ~n6354 & n6468 ;
  assign n9305 = n6362 & n6576 ;
  assign n9306 = ~n6366 & n6466 ;
  assign n9307 = ~n9305 & ~n9306 ;
  assign n9308 = ~n9304 & n9307 ;
  assign n9309 = n6452 & n6474 ;
  assign n9310 = n9308 & ~n9309 ;
  assign n9311 = ~n4325 & ~n9310 ;
  assign n9312 = ~n9310 & ~n9311 ;
  assign n9313 = ~n4325 & ~n9311 ;
  assign n9314 = ~n9312 & ~n9313 ;
  assign n9315 = ~n4325 & ~n6375 ;
  assign n9316 = n4075 & n4091 ;
  assign n9317 = ~n4075 & ~n4091 ;
  assign n9318 = ~n9316 & ~n9317 ;
  assign n9319 = n9315 & n9318 ;
  assign n9320 = ~n9315 & ~n9318 ;
  assign n9321 = ~n9319 & ~n9320 ;
  assign n9322 = ~n9314 & n9321 ;
  assign n9323 = ~n9314 & ~n9322 ;
  assign n9324 = n9321 & ~n9322 ;
  assign n9325 = ~n9323 & ~n9324 ;
  assign n9326 = ~n9303 & n9325 ;
  assign n9327 = n9303 & ~n9325 ;
  assign n9328 = ~n9326 & ~n9327 ;
  assign n9329 = n6499 & n7072 ;
  assign n9330 = n6495 & n7077 ;
  assign n9331 = n6497 & ~n7080 ;
  assign n9332 = ~n9330 & ~n9331 ;
  assign n9333 = ~n9329 & n9332 ;
  assign n9334 = ~n6490 & n9333 ;
  assign n9335 = ~n7102 & n9333 ;
  assign n9336 = ~n9334 & ~n9335 ;
  assign n9337 = n4469 & ~n9336 ;
  assign n9338 = ~n4469 & n9336 ;
  assign n9339 = ~n9337 & ~n9338 ;
  assign n9340 = ~n9328 & n9339 ;
  assign n9341 = ~n9328 & ~n9340 ;
  assign n9342 = n9339 & ~n9340 ;
  assign n9343 = ~n9341 & ~n9342 ;
  assign n9344 = ~n9302 & ~n9343 ;
  assign n9345 = ~n9302 & ~n9344 ;
  assign n9346 = ~n9343 & ~n9344 ;
  assign n9347 = ~n9345 & ~n9346 ;
  assign n9348 = n9301 & ~n9347 ;
  assign n9349 = n9301 & ~n9348 ;
  assign n9350 = ~n9347 & ~n9348 ;
  assign n9351 = ~n9349 & ~n9350 ;
  assign n9352 = ~n9286 & n9351 ;
  assign n9353 = n9286 & ~n9351 ;
  assign n9354 = ~n9352 & ~n9353 ;
  assign n9355 = ~n9162 & ~n9165 ;
  assign n9356 = n9354 & n9355 ;
  assign n9357 = ~n9354 & ~n9355 ;
  assign n9358 = ~n9356 & ~n9357 ;
  assign n9359 = n4731 & n6081 ;
  assign n9360 = n8839 & n9359 ;
  assign n9361 = n4609 & n9360 ;
  assign n9362 = n9077 & n9361 ;
  assign n9363 = ~n3929 & n9362 ;
  assign n9364 = ~n3994 & n9363 ;
  assign n9365 = ~n3937 & n9364 ;
  assign n9366 = ~n4018 & n9365 ;
  assign n9367 = n4890 & n9366 ;
  assign n9368 = ~n3968 & n9367 ;
  assign n9369 = ~n4245 & n9368 ;
  assign n9370 = n9358 & ~n9369 ;
  assign n9371 = ~n9358 & n9369 ;
  assign n9372 = ~n9370 & ~n9371 ;
  assign n9373 = ~n9285 & n9372 ;
  assign n9374 = n9285 & ~n9372 ;
  assign n9375 = ~n9373 & ~n9374 ;
  assign n9376 = n9175 & n9375 ;
  assign n9377 = ~n9175 & ~n9375 ;
  assign n9378 = ~n9376 & ~n9377 ;
  assign n9379 = ~n9176 & n9177 ;
  assign n9380 = ~n7831 & ~n9379 ;
  assign n9381 = ~n9378 & n9380 ;
  assign n9382 = n9378 & ~n9380 ;
  assign n9383 = ~n9381 & ~n9382 ;
  assign n9386 = n9383 & ~x31 ;
  assign n9387 = ~n9385 & ~n9386 ;
  assign n9388 = ~n9271 & ~n9274 ;
  assign n9389 = n584 & n2156 ;
  assign n9390 = n140 & n9389 ;
  assign n9391 = ~n196 & n9390 ;
  assign n9392 = ~n194 & n9391 ;
  assign n9393 = ~n142 & n9392 ;
  assign n9394 = ~n200 & n9393 ;
  assign n9395 = ~n421 & n9394 ;
  assign n9396 = ~n86 & n9395 ;
  assign n9397 = ~n186 & n9396 ;
  assign n9398 = n936 & n2317 ;
  assign n9399 = n954 & n9398 ;
  assign n9400 = n3653 & n9399 ;
  assign n9401 = n9397 & n9400 ;
  assign n9402 = ~n383 & n9401 ;
  assign n9403 = ~n232 & n9402 ;
  assign n9404 = ~n182 & n9403 ;
  assign n9405 = ~n336 & n9404 ;
  assign n9406 = ~n199 & n9405 ;
  assign n9407 = ~n301 & n9406 ;
  assign n9408 = ~n444 & n9407 ;
  assign n9409 = ~n9187 & ~n9252 ;
  assign n9410 = ~n9258 & ~n9409 ;
  assign n9411 = ~n9200 & ~n9249 ;
  assign n9412 = n2783 & n3725 ;
  assign n9413 = n2785 & n7700 ;
  assign n9414 = ~n9412 & ~n9413 ;
  assign n9415 = n2792 & n8018 ;
  assign n9416 = n9414 & ~n9415 ;
  assign n9417 = ~n996 & ~n9416 ;
  assign n9418 = ~n9416 & ~n9417 ;
  assign n9419 = ~n996 & ~n9417 ;
  assign n9420 = ~n9418 & ~n9419 ;
  assign n9421 = ~n9241 & ~n9245 ;
  assign n9422 = ~n9204 & ~n9226 ;
  assign n9423 = ~n9223 & ~n9422 ;
  assign n9424 = ~n500 & n2537 ;
  assign n9425 = ~n9217 & ~n9220 ;
  assign n9426 = ~n9424 & ~n9425 ;
  assign n9427 = ~n9424 & ~n9426 ;
  assign n9428 = ~n9425 & ~n9426 ;
  assign n9429 = ~n9427 & ~n9428 ;
  assign n9430 = n2643 & n3252 ;
  assign n9431 = ~n2541 & n2751 ;
  assign n9432 = ~n2529 & n2641 ;
  assign n9433 = ~n9431 & ~n9432 ;
  assign n9434 = ~n9430 & n9433 ;
  assign n9435 = ~n2649 & n9434 ;
  assign n9436 = ~n3307 & n9434 ;
  assign n9437 = ~n9435 & ~n9436 ;
  assign n9438 = n500 & ~n9437 ;
  assign n9439 = ~n500 & n9437 ;
  assign n9440 = ~n9438 & ~n9439 ;
  assign n9441 = ~n9429 & n9440 ;
  assign n9442 = n9429 & ~n9440 ;
  assign n9443 = ~n9441 & ~n9442 ;
  assign n9444 = ~n9423 & n9443 ;
  assign n9445 = ~n9423 & ~n9444 ;
  assign n9446 = n9443 & ~n9444 ;
  assign n9447 = ~n9445 & ~n9446 ;
  assign n9448 = n2674 & ~n3603 ;
  assign n9449 = n2670 & ~n3255 ;
  assign n9450 = n2672 & n3247 ;
  assign n9451 = ~n9449 & ~n9450 ;
  assign n9452 = ~n9448 & n9451 ;
  assign n9453 = n2665 & n3616 ;
  assign n9454 = n9452 & ~n9453 ;
  assign n9455 = ~n644 & ~n9454 ;
  assign n9456 = n644 & n9454 ;
  assign n9457 = ~n9455 & ~n9456 ;
  assign n9458 = ~n9447 & n9457 ;
  assign n9459 = ~n9446 & ~n9457 ;
  assign n9460 = ~n9445 & n9459 ;
  assign n9461 = ~n9458 & ~n9460 ;
  assign n9462 = ~n9421 & n9461 ;
  assign n9463 = n9421 & ~n9461 ;
  assign n9464 = ~n9462 & ~n9463 ;
  assign n9465 = ~n9420 & n9464 ;
  assign n9466 = n9420 & ~n9464 ;
  assign n9467 = ~n9465 & ~n9466 ;
  assign n9468 = ~n9411 & n9467 ;
  assign n9469 = n9411 & ~n9467 ;
  assign n9470 = ~n9468 & ~n9469 ;
  assign n9471 = ~n9410 & n9470 ;
  assign n9472 = n9410 & ~n9470 ;
  assign n9473 = ~n9471 & ~n9472 ;
  assign n9474 = n9408 & ~n9473 ;
  assign n9475 = ~n9408 & n9473 ;
  assign n9476 = ~n9474 & ~n9475 ;
  assign n9477 = ~n9388 & n9476 ;
  assign n9478 = n9388 & ~n9476 ;
  assign n9479 = ~n9477 & ~n9478 ;
  assign n9480 = ~n9277 & ~n9479 ;
  assign n9481 = n9277 & n9479 ;
  assign n9482 = ~n9480 & ~n9481 ;
  assign n9483 = ~n9279 & n9280 ;
  assign n9484 = ~n7831 & ~n9483 ;
  assign n9485 = ~n9482 & n9484 ;
  assign n9486 = n9482 & ~n9484 ;
  assign n9487 = ~n9485 & ~n9486 ;
  assign n9589 = ~n9487 & x32 ;
  assign n9488 = ~n9370 & ~n9373 ;
  assign n9489 = n4409 & n5981 ;
  assign n9490 = n3965 & n9489 ;
  assign n9491 = ~n4021 & n9490 ;
  assign n9492 = ~n4019 & n9491 ;
  assign n9493 = ~n3967 & n9492 ;
  assign n9494 = ~n4025 & n9493 ;
  assign n9495 = ~n4246 & n9494 ;
  assign n9496 = ~n3911 & n9495 ;
  assign n9497 = ~n4011 & n9496 ;
  assign n9498 = n4761 & n6142 ;
  assign n9499 = n4779 & n9498 ;
  assign n9500 = n7478 & n9499 ;
  assign n9501 = n9497 & n9500 ;
  assign n9502 = ~n4208 & n9501 ;
  assign n9503 = ~n4057 & n9502 ;
  assign n9504 = ~n4007 & n9503 ;
  assign n9505 = ~n4161 & n9504 ;
  assign n9506 = ~n4024 & n9505 ;
  assign n9507 = ~n4126 & n9506 ;
  assign n9508 = ~n4269 & n9507 ;
  assign n9509 = ~n9286 & ~n9351 ;
  assign n9510 = ~n9357 & ~n9509 ;
  assign n9511 = ~n9299 & ~n9348 ;
  assign n9512 = n6608 & n7550 ;
  assign n9513 = n6610 & n7857 ;
  assign n9514 = ~n9512 & ~n9513 ;
  assign n9515 = n6617 & n8149 ;
  assign n9516 = n9514 & ~n9515 ;
  assign n9517 = ~n4821 & ~n9516 ;
  assign n9518 = ~n9516 & ~n9517 ;
  assign n9519 = ~n4821 & ~n9517 ;
  assign n9520 = ~n9518 & ~n9519 ;
  assign n9521 = ~n9340 & ~n9344 ;
  assign n9522 = ~n9303 & ~n9325 ;
  assign n9523 = ~n9322 & ~n9522 ;
  assign n9524 = ~n4325 & n6362 ;
  assign n9525 = ~n9316 & ~n9319 ;
  assign n9526 = ~n9524 & ~n9525 ;
  assign n9527 = ~n9524 & ~n9526 ;
  assign n9528 = ~n9525 & ~n9526 ;
  assign n9529 = ~n9527 & ~n9528 ;
  assign n9530 = n6468 & n7077 ;
  assign n9531 = ~n6366 & n6576 ;
  assign n9532 = ~n6354 & n6466 ;
  assign n9533 = ~n9531 & ~n9532 ;
  assign n9534 = ~n9530 & n9533 ;
  assign n9535 = ~n6474 & n9534 ;
  assign n9536 = ~n7132 & n9534 ;
  assign n9537 = ~n9535 & ~n9536 ;
  assign n9538 = n4325 & ~n9537 ;
  assign n9539 = ~n4325 & n9537 ;
  assign n9540 = ~n9538 & ~n9539 ;
  assign n9541 = ~n9529 & n9540 ;
  assign n9542 = n9529 & ~n9540 ;
  assign n9543 = ~n9541 & ~n9542 ;
  assign n9544 = ~n9523 & n9543 ;
  assign n9545 = ~n9523 & ~n9544 ;
  assign n9546 = n9543 & ~n9544 ;
  assign n9547 = ~n9545 & ~n9546 ;
  assign n9548 = n6499 & ~n7428 ;
  assign n9549 = n6495 & ~n7080 ;
  assign n9550 = n6497 & n7072 ;
  assign n9551 = ~n9549 & ~n9550 ;
  assign n9552 = ~n9548 & n9551 ;
  assign n9553 = n6490 & n7441 ;
  assign n9554 = n9552 & ~n9553 ;
  assign n9555 = ~n4469 & ~n9554 ;
  assign n9556 = n4469 & n9554 ;
  assign n9557 = ~n9555 & ~n9556 ;
  assign n9558 = ~n9547 & n9557 ;
  assign n9559 = ~n9546 & ~n9557 ;
  assign n9560 = ~n9545 & n9559 ;
  assign n9561 = ~n9558 & ~n9560 ;
  assign n9562 = ~n9521 & n9561 ;
  assign n9563 = n9521 & ~n9561 ;
  assign n9564 = ~n9562 & ~n9563 ;
  assign n9565 = ~n9520 & n9564 ;
  assign n9566 = n9520 & ~n9564 ;
  assign n9567 = ~n9565 & ~n9566 ;
  assign n9568 = ~n9511 & n9567 ;
  assign n9569 = n9511 & ~n9567 ;
  assign n9570 = ~n9568 & ~n9569 ;
  assign n9571 = ~n9510 & n9570 ;
  assign n9572 = n9510 & ~n9570 ;
  assign n9573 = ~n9571 & ~n9572 ;
  assign n9574 = n9508 & ~n9573 ;
  assign n9575 = ~n9508 & n9573 ;
  assign n9576 = ~n9574 & ~n9575 ;
  assign n9577 = ~n9488 & n9576 ;
  assign n9578 = n9488 & ~n9576 ;
  assign n9579 = ~n9577 & ~n9578 ;
  assign n9580 = ~n9376 & ~n9579 ;
  assign n9581 = n9376 & n9579 ;
  assign n9582 = ~n9580 & ~n9581 ;
  assign n9583 = ~n9378 & n9379 ;
  assign n9584 = ~n7831 & ~n9583 ;
  assign n9585 = ~n9582 & n9584 ;
  assign n9586 = n9582 & ~n9584 ;
  assign n9587 = ~n9585 & ~n9586 ;
  assign n9590 = n9587 & ~x32 ;
  assign n9591 = ~n9589 & ~n9590 ;
  assign n9592 = ~n9475 & ~n9477 ;
  assign n9593 = n732 & n784 ;
  assign n9594 = n179 & n9593 ;
  assign n9595 = n3206 & n9594 ;
  assign n9596 = n2407 & n9595 ;
  assign n9597 = n3234 & n9596 ;
  assign n9598 = ~n312 & n9597 ;
  assign n9599 = ~n302 & n9598 ;
  assign n9600 = ~n200 & n9599 ;
  assign n9601 = ~n108 & n9600 ;
  assign n9602 = ~n209 & n9601 ;
  assign n9603 = ~n331 & n9602 ;
  assign n9604 = ~n191 & n9603 ;
  assign n9605 = ~n9462 & ~n9465 ;
  assign n9606 = ~n9426 & ~n9441 ;
  assign n9607 = n2643 & ~n3255 ;
  assign n9608 = ~n2529 & n2751 ;
  assign n9609 = n2641 & n3252 ;
  assign n9610 = ~n9608 & ~n9609 ;
  assign n9611 = ~n9607 & n9610 ;
  assign n9612 = n2649 & n3293 ;
  assign n9613 = n9611 & ~n9612 ;
  assign n9614 = ~n500 & ~n9613 ;
  assign n9615 = ~n9613 & ~n9614 ;
  assign n9616 = ~n500 & ~n9614 ;
  assign n9617 = ~n9615 & ~n9616 ;
  assign n9618 = ~n500 & n2619 ;
  assign n9619 = ~n9617 & ~n9618 ;
  assign n9620 = ~n9617 & ~n9619 ;
  assign n9621 = ~n9618 & ~n9619 ;
  assign n9622 = ~n9620 & ~n9621 ;
  assign n9623 = ~n9606 & n9622 ;
  assign n9624 = n9606 & ~n9622 ;
  assign n9625 = ~n9623 & ~n9624 ;
  assign n9626 = n2674 & n3725 ;
  assign n9627 = n2670 & n3247 ;
  assign n9628 = n2672 & ~n3603 ;
  assign n9629 = ~n9627 & ~n9628 ;
  assign n9630 = ~n9626 & n9629 ;
  assign n9631 = n2665 & n3737 ;
  assign n9632 = n9630 & ~n9631 ;
  assign n9633 = ~n644 & ~n9632 ;
  assign n9634 = n644 & n9632 ;
  assign n9635 = ~n9633 & ~n9634 ;
  assign n9636 = ~n9625 & n9635 ;
  assign n9637 = ~n9625 & ~n9636 ;
  assign n9638 = n9635 & ~n9636 ;
  assign n9639 = ~n9637 & ~n9638 ;
  assign n9640 = ~n9444 & ~n9458 ;
  assign n9641 = n2783 & n7700 ;
  assign n9642 = n2792 & n8016 ;
  assign n9643 = ~n9641 & ~n9642 ;
  assign n9644 = ~n996 & n9643 ;
  assign n9645 = n996 & ~n9643 ;
  assign n9646 = ~n9644 & ~n9645 ;
  assign n9647 = ~n9640 & ~n9646 ;
  assign n9648 = n9640 & n9646 ;
  assign n9649 = ~n9647 & ~n9648 ;
  assign n9650 = ~n9639 & n9649 ;
  assign n9651 = ~n9639 & ~n9650 ;
  assign n9652 = n9649 & ~n9650 ;
  assign n9653 = ~n9651 & ~n9652 ;
  assign n9654 = ~n9605 & n9653 ;
  assign n9655 = n9605 & ~n9653 ;
  assign n9656 = ~n9654 & ~n9655 ;
  assign n9657 = ~n9468 & ~n9471 ;
  assign n9658 = n9656 & n9657 ;
  assign n9659 = ~n9656 & ~n9657 ;
  assign n9660 = ~n9658 & ~n9659 ;
  assign n9661 = n9604 & ~n9660 ;
  assign n9662 = ~n9604 & n9660 ;
  assign n9663 = ~n9661 & ~n9662 ;
  assign n9664 = ~n9592 & n9663 ;
  assign n9665 = n9592 & ~n9663 ;
  assign n9666 = ~n9664 & ~n9665 ;
  assign n9667 = ~n9481 & ~n9666 ;
  assign n9668 = n9481 & n9666 ;
  assign n9669 = ~n9667 & ~n9668 ;
  assign n9670 = ~n9482 & n9483 ;
  assign n9671 = ~n7831 & ~n9670 ;
  assign n9672 = ~n9669 & n9671 ;
  assign n9673 = n9669 & ~n9671 ;
  assign n9674 = ~n9672 & ~n9673 ;
  assign n9759 = ~n9674 & x33 ;
  assign n9675 = ~n9575 & ~n9577 ;
  assign n9676 = n4557 & n4609 ;
  assign n9677 = n4004 & n9676 ;
  assign n9678 = n7031 & n9677 ;
  assign n9679 = n6232 & n9678 ;
  assign n9680 = n7059 & n9679 ;
  assign n9681 = ~n4137 & n9680 ;
  assign n9682 = ~n4127 & n9681 ;
  assign n9683 = ~n4025 & n9682 ;
  assign n9684 = ~n3933 & n9683 ;
  assign n9685 = ~n4034 & n9684 ;
  assign n9686 = ~n4156 & n9685 ;
  assign n9687 = ~n4016 & n9686 ;
  assign n9688 = ~n9562 & ~n9565 ;
  assign n9689 = ~n9526 & ~n9541 ;
  assign n9690 = n6468 & ~n7080 ;
  assign n9691 = ~n6354 & n6576 ;
  assign n9692 = n6466 & n7077 ;
  assign n9693 = ~n9691 & ~n9692 ;
  assign n9694 = ~n9690 & n9693 ;
  assign n9695 = n6474 & n7118 ;
  assign n9696 = n9694 & ~n9695 ;
  assign n9697 = ~n4325 & ~n9696 ;
  assign n9698 = ~n9696 & ~n9697 ;
  assign n9699 = ~n4325 & ~n9697 ;
  assign n9700 = ~n9698 & ~n9699 ;
  assign n9701 = ~n4325 & n6444 ;
  assign n9702 = ~n9700 & ~n9701 ;
  assign n9703 = ~n9700 & ~n9702 ;
  assign n9704 = ~n9701 & ~n9702 ;
  assign n9705 = ~n9703 & ~n9704 ;
  assign n9706 = ~n9689 & n9705 ;
  assign n9707 = n9689 & ~n9705 ;
  assign n9708 = ~n9706 & ~n9707 ;
  assign n9709 = n6499 & n7550 ;
  assign n9710 = n6495 & n7072 ;
  assign n9711 = n6497 & ~n7428 ;
  assign n9712 = ~n9710 & ~n9711 ;
  assign n9713 = ~n9709 & n9712 ;
  assign n9714 = n6490 & n7562 ;
  assign n9715 = n9713 & ~n9714 ;
  assign n9716 = ~n4469 & ~n9715 ;
  assign n9717 = n4469 & n9715 ;
  assign n9718 = ~n9716 & ~n9717 ;
  assign n9719 = ~n9708 & n9718 ;
  assign n9720 = ~n9708 & ~n9719 ;
  assign n9721 = n9718 & ~n9719 ;
  assign n9722 = ~n9720 & ~n9721 ;
  assign n9723 = ~n9544 & ~n9558 ;
  assign n9724 = n6608 & n7857 ;
  assign n9725 = n6617 & n8147 ;
  assign n9726 = ~n9724 & ~n9725 ;
  assign n9727 = ~n4821 & n9726 ;
  assign n9728 = n4821 & ~n9726 ;
  assign n9729 = ~n9727 & ~n9728 ;
  assign n9730 = ~n9723 & ~n9729 ;
  assign n9731 = n9723 & n9729 ;
  assign n9732 = ~n9730 & ~n9731 ;
  assign n9733 = ~n9722 & n9732 ;
  assign n9734 = ~n9722 & ~n9733 ;
  assign n9735 = n9732 & ~n9733 ;
  assign n9736 = ~n9734 & ~n9735 ;
  assign n9737 = ~n9688 & n9736 ;
  assign n9738 = n9688 & ~n9736 ;
  assign n9739 = ~n9737 & ~n9738 ;
  assign n9740 = ~n9568 & ~n9571 ;
  assign n9741 = n9739 & n9740 ;
  assign n9742 = ~n9739 & ~n9740 ;
  assign n9743 = ~n9741 & ~n9742 ;
  assign n9744 = n9687 & ~n9743 ;
  assign n9745 = ~n9687 & n9743 ;
  assign n9746 = ~n9744 & ~n9745 ;
  assign n9747 = ~n9675 & n9746 ;
  assign n9748 = n9675 & ~n9746 ;
  assign n9749 = ~n9747 & ~n9748 ;
  assign n9750 = ~n9581 & ~n9749 ;
  assign n9751 = n9581 & n9749 ;
  assign n9752 = ~n9750 & ~n9751 ;
  assign n9753 = ~n9582 & n9583 ;
  assign n9754 = ~n7831 & ~n9753 ;
  assign n9755 = ~n9752 & n9754 ;
  assign n9756 = n9752 & ~n9754 ;
  assign n9757 = ~n9755 & ~n9756 ;
  assign n9760 = n9757 & ~x33 ;
  assign n9761 = ~n9759 & ~n9760 ;
  assign n9762 = ~n9662 & ~n9664 ;
  assign n9763 = n234 & n630 ;
  assign n9764 = n451 & n9763 ;
  assign n9765 = n480 & n9764 ;
  assign n9766 = n185 & n9765 ;
  assign n9767 = n3641 & n9766 ;
  assign n9768 = n1079 & n9767 ;
  assign n9769 = n3234 & n9768 ;
  assign n9770 = n952 & n9769 ;
  assign n9771 = ~n287 & n9770 ;
  assign n9772 = ~n167 & n9771 ;
  assign n9773 = ~n290 & n9772 ;
  assign n9774 = ~n9605 & ~n9653 ;
  assign n9775 = ~n9659 & ~n9774 ;
  assign n9776 = ~n9647 & ~n9650 ;
  assign n9777 = ~n2541 & ~n9424 ;
  assign n9778 = ~n500 & n9777 ;
  assign n9779 = ~n9619 & ~n9778 ;
  assign n9780 = ~n500 & ~n2529 ;
  assign n9781 = ~n996 & ~n9780 ;
  assign n9782 = n996 & n9780 ;
  assign n9783 = n9424 & ~n9782 ;
  assign n9784 = ~n9781 & n9783 ;
  assign n9785 = n9424 & ~n9784 ;
  assign n9786 = ~n9782 & ~n9784 ;
  assign n9787 = ~n9781 & n9786 ;
  assign n9788 = ~n9785 & ~n9787 ;
  assign n9789 = ~n9779 & ~n9788 ;
  assign n9790 = ~n9779 & ~n9789 ;
  assign n9791 = ~n9788 & ~n9789 ;
  assign n9792 = ~n9790 & ~n9791 ;
  assign n9793 = n2643 & n3247 ;
  assign n9794 = n2751 & n3252 ;
  assign n9795 = n2641 & ~n3255 ;
  assign n9796 = ~n9794 & ~n9795 ;
  assign n9797 = ~n9793 & n9796 ;
  assign n9798 = n2649 & n3277 ;
  assign n9799 = n9797 & ~n9798 ;
  assign n9800 = ~n500 & ~n9799 ;
  assign n9801 = ~n500 & ~n9800 ;
  assign n9802 = ~n9799 & ~n9800 ;
  assign n9803 = ~n9801 & ~n9802 ;
  assign n9804 = ~n9792 & ~n9803 ;
  assign n9805 = ~n9792 & ~n9804 ;
  assign n9806 = ~n9803 & ~n9804 ;
  assign n9807 = ~n9805 & ~n9806 ;
  assign n9808 = ~n9606 & ~n9622 ;
  assign n9809 = ~n9636 & ~n9808 ;
  assign n9810 = n2674 & n7700 ;
  assign n9811 = n2670 & ~n3603 ;
  assign n9812 = n2672 & n3725 ;
  assign n9813 = ~n9811 & ~n9812 ;
  assign n9814 = ~n9810 & n9813 ;
  assign n9815 = ~n2665 & n9814 ;
  assign n9816 = ~n7712 & n9814 ;
  assign n9817 = ~n9815 & ~n9816 ;
  assign n9818 = n644 & ~n9817 ;
  assign n9819 = ~n644 & n9817 ;
  assign n9820 = ~n9818 & ~n9819 ;
  assign n9821 = ~n9809 & n9820 ;
  assign n9822 = ~n9809 & ~n9821 ;
  assign n9823 = n9820 & ~n9821 ;
  assign n9824 = ~n9822 & ~n9823 ;
  assign n9825 = ~n9807 & ~n9824 ;
  assign n9826 = n9807 & ~n9823 ;
  assign n9827 = ~n9822 & n9826 ;
  assign n9828 = ~n9825 & ~n9827 ;
  assign n9829 = ~n9776 & n9828 ;
  assign n9830 = n9776 & ~n9828 ;
  assign n9831 = ~n9829 & ~n9830 ;
  assign n9832 = ~n9775 & n9831 ;
  assign n9833 = n9775 & ~n9831 ;
  assign n9834 = ~n9832 & ~n9833 ;
  assign n9835 = n9773 & ~n9834 ;
  assign n9836 = ~n9773 & n9834 ;
  assign n9837 = ~n9835 & ~n9836 ;
  assign n9838 = ~n9762 & n9837 ;
  assign n9839 = n9762 & ~n9837 ;
  assign n9840 = ~n9838 & ~n9839 ;
  assign n9841 = ~n9668 & ~n9840 ;
  assign n9842 = n9668 & n9840 ;
  assign n9843 = ~n9841 & ~n9842 ;
  assign n9844 = ~n9669 & n9670 ;
  assign n9845 = ~n7831 & ~n9844 ;
  assign n9846 = ~n9843 & n9845 ;
  assign n9847 = n9843 & ~n9845 ;
  assign n9848 = ~n9846 & ~n9847 ;
  assign n9937 = ~n9848 & x34 ;
  assign n9849 = ~n9745 & ~n9747 ;
  assign n9850 = n4059 & n4455 ;
  assign n9851 = n4276 & n9850 ;
  assign n9852 = n4305 & n9851 ;
  assign n9853 = n4010 & n9852 ;
  assign n9854 = n7466 & n9853 ;
  assign n9855 = n4904 & n9854 ;
  assign n9856 = n7059 & n9855 ;
  assign n9857 = n4777 & n9856 ;
  assign n9858 = ~n4112 & n9857 ;
  assign n9859 = ~n3992 & n9858 ;
  assign n9860 = ~n4115 & n9859 ;
  assign n9861 = ~n9688 & ~n9736 ;
  assign n9862 = ~n9742 & ~n9861 ;
  assign n9863 = ~n9730 & ~n9733 ;
  assign n9864 = ~n6366 & ~n9524 ;
  assign n9865 = ~n4325 & n9864 ;
  assign n9866 = ~n9702 & ~n9865 ;
  assign n9867 = ~n4325 & ~n6354 ;
  assign n9868 = ~n4821 & ~n9867 ;
  assign n9869 = n4821 & n9867 ;
  assign n9870 = n9524 & ~n9869 ;
  assign n9871 = ~n9868 & n9870 ;
  assign n9872 = n9524 & ~n9871 ;
  assign n9873 = ~n9869 & ~n9871 ;
  assign n9874 = ~n9868 & n9873 ;
  assign n9875 = ~n9872 & ~n9874 ;
  assign n9876 = ~n9866 & ~n9875 ;
  assign n9877 = ~n9866 & ~n9876 ;
  assign n9878 = ~n9875 & ~n9876 ;
  assign n9879 = ~n9877 & ~n9878 ;
  assign n9880 = n6468 & n7072 ;
  assign n9881 = n6576 & n7077 ;
  assign n9882 = n6466 & ~n7080 ;
  assign n9883 = ~n9881 & ~n9882 ;
  assign n9884 = ~n9880 & n9883 ;
  assign n9885 = n6474 & n7102 ;
  assign n9886 = n9884 & ~n9885 ;
  assign n9887 = ~n4325 & ~n9886 ;
  assign n9888 = ~n4325 & ~n9887 ;
  assign n9889 = ~n9886 & ~n9887 ;
  assign n9890 = ~n9888 & ~n9889 ;
  assign n9891 = ~n9879 & ~n9890 ;
  assign n9892 = ~n9879 & ~n9891 ;
  assign n9893 = ~n9890 & ~n9891 ;
  assign n9894 = ~n9892 & ~n9893 ;
  assign n9895 = ~n9689 & ~n9705 ;
  assign n9896 = ~n9719 & ~n9895 ;
  assign n9897 = n6499 & n7857 ;
  assign n9898 = n6495 & ~n7428 ;
  assign n9899 = n6497 & n7550 ;
  assign n9900 = ~n9898 & ~n9899 ;
  assign n9901 = ~n9897 & n9900 ;
  assign n9902 = ~n6490 & n9901 ;
  assign n9903 = ~n7869 & n9901 ;
  assign n9904 = ~n9902 & ~n9903 ;
  assign n9905 = n4469 & ~n9904 ;
  assign n9906 = ~n4469 & n9904 ;
  assign n9907 = ~n9905 & ~n9906 ;
  assign n9908 = ~n9896 & n9907 ;
  assign n9909 = ~n9896 & ~n9908 ;
  assign n9910 = n9907 & ~n9908 ;
  assign n9911 = ~n9909 & ~n9910 ;
  assign n9912 = ~n9894 & ~n9911 ;
  assign n9913 = n9894 & ~n9910 ;
  assign n9914 = ~n9909 & n9913 ;
  assign n9915 = ~n9912 & ~n9914 ;
  assign n9916 = ~n9863 & n9915 ;
  assign n9917 = n9863 & ~n9915 ;
  assign n9918 = ~n9916 & ~n9917 ;
  assign n9919 = ~n9862 & n9918 ;
  assign n9920 = n9862 & ~n9918 ;
  assign n9921 = ~n9919 & ~n9920 ;
  assign n9922 = n9860 & ~n9921 ;
  assign n9923 = ~n9860 & n9921 ;
  assign n9924 = ~n9922 & ~n9923 ;
  assign n9925 = ~n9849 & n9924 ;
  assign n9926 = n9849 & ~n9924 ;
  assign n9927 = ~n9925 & ~n9926 ;
  assign n9928 = ~n9751 & ~n9927 ;
  assign n9929 = n9751 & n9927 ;
  assign n9930 = ~n9928 & ~n9929 ;
  assign n9931 = ~n9752 & n9753 ;
  assign n9932 = ~n7831 & ~n9931 ;
  assign n9933 = ~n9930 & n9932 ;
  assign n9934 = n9930 & ~n9932 ;
  assign n9935 = ~n9933 & ~n9934 ;
  assign n9938 = n9935 & ~x34 ;
  assign n9939 = ~n9937 & ~n9938 ;
  assign n9940 = ~n9836 & ~n9838 ;
  assign n9941 = n886 & n944 ;
  assign n9942 = n474 & n9941 ;
  assign n9943 = n3709 & n9942 ;
  assign n9944 = n611 & n9943 ;
  assign n9945 = n428 & n9944 ;
  assign n9946 = ~n311 & n9945 ;
  assign n9947 = ~n9829 & ~n9832 ;
  assign n9948 = ~n9821 & ~n9825 ;
  assign n9949 = ~n9789 & ~n9804 ;
  assign n9950 = ~n500 & n3252 ;
  assign n9951 = ~n9786 & n9950 ;
  assign n9952 = n9786 & ~n9950 ;
  assign n9953 = ~n9951 & ~n9952 ;
  assign n9954 = n2643 & ~n3603 ;
  assign n9955 = n2751 & ~n3255 ;
  assign n9956 = n2641 & n3247 ;
  assign n9957 = ~n9955 & ~n9956 ;
  assign n9958 = ~n9954 & n9957 ;
  assign n9959 = ~n2649 & n9958 ;
  assign n9960 = ~n3616 & n9958 ;
  assign n9961 = ~n9959 & ~n9960 ;
  assign n9962 = n500 & ~n9961 ;
  assign n9963 = ~n500 & n9961 ;
  assign n9964 = ~n9962 & ~n9963 ;
  assign n9965 = ~n9953 & n9964 ;
  assign n9966 = n9953 & ~n9964 ;
  assign n9967 = ~n9965 & ~n9966 ;
  assign n9968 = ~n9949 & n9967 ;
  assign n9969 = ~n9949 & ~n9968 ;
  assign n9970 = n9967 & ~n9968 ;
  assign n9971 = ~n9969 & ~n9970 ;
  assign n9972 = n2670 & n3725 ;
  assign n9973 = n2672 & n7700 ;
  assign n9974 = ~n9972 & ~n9973 ;
  assign n9975 = n2665 & n8018 ;
  assign n9976 = n9974 & ~n9975 ;
  assign n9977 = ~n644 & ~n9976 ;
  assign n9978 = n644 & n9976 ;
  assign n9979 = ~n9977 & ~n9978 ;
  assign n9980 = ~n9971 & n9979 ;
  assign n9981 = ~n9970 & ~n9979 ;
  assign n9982 = ~n9969 & n9981 ;
  assign n9983 = ~n9980 & ~n9982 ;
  assign n9984 = ~n9948 & n9983 ;
  assign n9985 = n9948 & ~n9983 ;
  assign n9986 = ~n9984 & ~n9985 ;
  assign n9987 = ~n9947 & n9986 ;
  assign n9988 = n9947 & ~n9986 ;
  assign n9989 = ~n9987 & ~n9988 ;
  assign n9990 = n9946 & ~n9989 ;
  assign n9991 = ~n9946 & n9989 ;
  assign n9992 = ~n9990 & ~n9991 ;
  assign n9993 = ~n9940 & n9992 ;
  assign n9994 = n9940 & ~n9992 ;
  assign n9995 = ~n9993 & ~n9994 ;
  assign n9996 = ~n9842 & ~n9995 ;
  assign n9997 = n9842 & n9995 ;
  assign n9998 = ~n9996 & ~n9997 ;
  assign n9999 = ~n9843 & n9844 ;
  assign n10000 = ~n7831 & ~n9999 ;
  assign n10001 = ~n9998 & n10000 ;
  assign n10002 = n9998 & ~n10000 ;
  assign n10003 = ~n10001 & ~n10002 ;
  assign n10069 = ~n10003 & x35 ;
  assign n10004 = ~n9923 & ~n9925 ;
  assign n10005 = n4711 & n4769 ;
  assign n10006 = n4299 & n10005 ;
  assign n10007 = n7534 & n10006 ;
  assign n10008 = n4436 & n10007 ;
  assign n10009 = n4253 & n10008 ;
  assign n10010 = ~n4136 & n10009 ;
  assign n10011 = ~n9916 & ~n9919 ;
  assign n10012 = ~n9908 & ~n9912 ;
  assign n10013 = ~n9876 & ~n9891 ;
  assign n10014 = ~n4325 & n7077 ;
  assign n10015 = ~n9873 & n10014 ;
  assign n10016 = n9873 & ~n10014 ;
  assign n10017 = ~n10015 & ~n10016 ;
  assign n10018 = n6468 & ~n7428 ;
  assign n10019 = n6576 & ~n7080 ;
  assign n10020 = n6466 & n7072 ;
  assign n10021 = ~n10019 & ~n10020 ;
  assign n10022 = ~n10018 & n10021 ;
  assign n10023 = ~n6474 & n10022 ;
  assign n10024 = ~n7441 & n10022 ;
  assign n10025 = ~n10023 & ~n10024 ;
  assign n10026 = n4325 & ~n10025 ;
  assign n10027 = ~n4325 & n10025 ;
  assign n10028 = ~n10026 & ~n10027 ;
  assign n10029 = ~n10017 & n10028 ;
  assign n10030 = n10017 & ~n10028 ;
  assign n10031 = ~n10029 & ~n10030 ;
  assign n10032 = ~n10013 & n10031 ;
  assign n10033 = ~n10013 & ~n10032 ;
  assign n10034 = n10031 & ~n10032 ;
  assign n10035 = ~n10033 & ~n10034 ;
  assign n10036 = n6495 & n7550 ;
  assign n10037 = n6497 & n7857 ;
  assign n10038 = ~n10036 & ~n10037 ;
  assign n10039 = n6490 & n8149 ;
  assign n10040 = n10038 & ~n10039 ;
  assign n10041 = ~n4469 & ~n10040 ;
  assign n10042 = n4469 & n10040 ;
  assign n10043 = ~n10041 & ~n10042 ;
  assign n10044 = ~n10035 & n10043 ;
  assign n10045 = ~n10034 & ~n10043 ;
  assign n10046 = ~n10033 & n10045 ;
  assign n10047 = ~n10044 & ~n10046 ;
  assign n10048 = ~n10012 & n10047 ;
  assign n10049 = n10012 & ~n10047 ;
  assign n10050 = ~n10048 & ~n10049 ;
  assign n10051 = ~n10011 & n10050 ;
  assign n10052 = n10011 & ~n10050 ;
  assign n10053 = ~n10051 & ~n10052 ;
  assign n10054 = n10010 & ~n10053 ;
  assign n10055 = ~n10010 & n10053 ;
  assign n10056 = ~n10054 & ~n10055 ;
  assign n10057 = ~n10004 & n10056 ;
  assign n10058 = n10004 & ~n10056 ;
  assign n10059 = ~n10057 & ~n10058 ;
  assign n10060 = ~n9929 & ~n10059 ;
  assign n10061 = n9929 & n10059 ;
  assign n10062 = ~n10060 & ~n10061 ;
  assign n10063 = ~n9930 & n9931 ;
  assign n10064 = ~n7831 & ~n10063 ;
  assign n10065 = ~n10062 & n10064 ;
  assign n10066 = n10062 & ~n10064 ;
  assign n10067 = ~n10065 & ~n10066 ;
  assign n10070 = n10067 & ~x35 ;
  assign n10071 = ~n10069 & ~n10070 ;
  assign n10072 = ~n9991 & ~n9993 ;
  assign n10073 = ~n152 & ~n161 ;
  assign n10074 = ~n182 & n10073 ;
  assign n10075 = ~n209 & n10074 ;
  assign n10076 = ~n310 & n10075 ;
  assign n10077 = n2342 & n10076 ;
  assign n10078 = n921 & n10077 ;
  assign n10079 = n7999 & n10078 ;
  assign n10080 = n2225 & n10079 ;
  assign n10081 = n355 & n10080 ;
  assign n10082 = ~n114 & n10081 ;
  assign n10083 = ~n109 & n10082 ;
  assign n10084 = ~n186 & n10083 ;
  assign n10085 = ~n9984 & ~n9987 ;
  assign n10086 = ~n9968 & ~n9980 ;
  assign n10087 = n2670 & n7700 ;
  assign n10088 = n2665 & n8016 ;
  assign n10089 = ~n10087 & ~n10088 ;
  assign n10090 = ~n644 & ~n10089 ;
  assign n10091 = n644 & n10089 ;
  assign n10092 = ~n10090 & ~n10091 ;
  assign n10093 = n2643 & n3725 ;
  assign n10094 = n2751 & n3247 ;
  assign n10095 = n2641 & ~n3603 ;
  assign n10096 = ~n10094 & ~n10095 ;
  assign n10097 = ~n10093 & n10096 ;
  assign n10098 = n2649 & n3737 ;
  assign n10099 = n10097 & ~n10098 ;
  assign n10100 = ~n500 & ~n10099 ;
  assign n10101 = ~n500 & ~n10100 ;
  assign n10102 = ~n10099 & ~n10100 ;
  assign n10103 = ~n10101 & ~n10102 ;
  assign n10104 = n10092 & ~n10103 ;
  assign n10105 = n10092 & ~n10104 ;
  assign n10106 = ~n10103 & ~n10104 ;
  assign n10107 = ~n10105 & ~n10106 ;
  assign n10108 = ~n9786 & ~n9950 ;
  assign n10109 = ~n9965 & ~n10108 ;
  assign n10110 = ~n500 & ~n3255 ;
  assign n10111 = ~n9950 & n10110 ;
  assign n10112 = n9950 & ~n10110 ;
  assign n10113 = ~n10109 & ~n10112 ;
  assign n10114 = ~n10111 & n10113 ;
  assign n10115 = ~n10109 & ~n10114 ;
  assign n10116 = ~n10112 & ~n10114 ;
  assign n10117 = ~n10111 & n10116 ;
  assign n10118 = ~n10115 & ~n10117 ;
  assign n10119 = ~n10107 & n10118 ;
  assign n10120 = n10107 & ~n10118 ;
  assign n10121 = ~n10119 & ~n10120 ;
  assign n10122 = ~n10086 & ~n10121 ;
  assign n10123 = n10086 & n10121 ;
  assign n10124 = ~n10122 & ~n10123 ;
  assign n10125 = ~n10085 & n10124 ;
  assign n10126 = n10085 & ~n10124 ;
  assign n10127 = ~n10125 & ~n10126 ;
  assign n10128 = n10084 & ~n10127 ;
  assign n10129 = ~n10084 & n10127 ;
  assign n10130 = ~n10128 & ~n10129 ;
  assign n10131 = ~n10072 & n10130 ;
  assign n10132 = n10072 & ~n10130 ;
  assign n10133 = ~n10131 & ~n10132 ;
  assign n10134 = ~n9997 & ~n10133 ;
  assign n10135 = n9997 & n10133 ;
  assign n10136 = ~n10134 & ~n10135 ;
  assign n10137 = ~n9998 & n9999 ;
  assign n10138 = ~n7831 & ~n10137 ;
  assign n10139 = ~n10136 & n10138 ;
  assign n10140 = n10136 & ~n10138 ;
  assign n10141 = ~n10139 & ~n10140 ;
  assign n10213 = ~n10141 & x36 ;
  assign n10142 = ~n10055 & ~n10057 ;
  assign n10143 = ~n3977 & ~n3986 ;
  assign n10144 = ~n4007 & n10143 ;
  assign n10145 = ~n4034 & n10144 ;
  assign n10146 = ~n4135 & n10145 ;
  assign n10147 = n6167 & n10146 ;
  assign n10148 = n4746 & n10147 ;
  assign n10149 = n8130 & n10148 ;
  assign n10150 = n6050 & n10149 ;
  assign n10151 = n4180 & n10150 ;
  assign n10152 = ~n3939 & n10151 ;
  assign n10153 = ~n3934 & n10152 ;
  assign n10154 = ~n4011 & n10153 ;
  assign n10155 = ~n10048 & ~n10051 ;
  assign n10156 = ~n10032 & ~n10044 ;
  assign n10157 = n6495 & n7857 ;
  assign n10158 = n6490 & n8147 ;
  assign n10159 = ~n10157 & ~n10158 ;
  assign n10160 = ~n4469 & ~n10159 ;
  assign n10161 = n4469 & n10159 ;
  assign n10162 = ~n10160 & ~n10161 ;
  assign n10163 = n6468 & n7550 ;
  assign n10164 = n6576 & n7072 ;
  assign n10165 = n6466 & ~n7428 ;
  assign n10166 = ~n10164 & ~n10165 ;
  assign n10167 = ~n10163 & n10166 ;
  assign n10168 = n6474 & n7562 ;
  assign n10169 = n10167 & ~n10168 ;
  assign n10170 = ~n4325 & ~n10169 ;
  assign n10171 = ~n4325 & ~n10170 ;
  assign n10172 = ~n10169 & ~n10170 ;
  assign n10173 = ~n10171 & ~n10172 ;
  assign n10174 = n10162 & ~n10173 ;
  assign n10175 = n10162 & ~n10174 ;
  assign n10176 = ~n10173 & ~n10174 ;
  assign n10177 = ~n10175 & ~n10176 ;
  assign n10178 = ~n9873 & ~n10014 ;
  assign n10179 = ~n10029 & ~n10178 ;
  assign n10180 = ~n4325 & ~n7080 ;
  assign n10181 = ~n10014 & n10180 ;
  assign n10182 = n10014 & ~n10180 ;
  assign n10183 = ~n10179 & ~n10182 ;
  assign n10184 = ~n10181 & n10183 ;
  assign n10185 = ~n10179 & ~n10184 ;
  assign n10186 = ~n10182 & ~n10184 ;
  assign n10187 = ~n10181 & n10186 ;
  assign n10188 = ~n10185 & ~n10187 ;
  assign n10189 = ~n10177 & n10188 ;
  assign n10190 = n10177 & ~n10188 ;
  assign n10191 = ~n10189 & ~n10190 ;
  assign n10192 = ~n10156 & ~n10191 ;
  assign n10193 = n10156 & n10191 ;
  assign n10194 = ~n10192 & ~n10193 ;
  assign n10195 = ~n10155 & n10194 ;
  assign n10196 = n10155 & ~n10194 ;
  assign n10197 = ~n10195 & ~n10196 ;
  assign n10198 = n10154 & ~n10197 ;
  assign n10199 = ~n10154 & n10197 ;
  assign n10200 = ~n10198 & ~n10199 ;
  assign n10201 = ~n10142 & n10200 ;
  assign n10202 = n10142 & ~n10200 ;
  assign n10203 = ~n10201 & ~n10202 ;
  assign n10204 = ~n10061 & ~n10203 ;
  assign n10205 = n10061 & n10203 ;
  assign n10206 = ~n10204 & ~n10205 ;
  assign n10207 = ~n10062 & n10063 ;
  assign n10208 = ~n7831 & ~n10207 ;
  assign n10209 = ~n10206 & n10208 ;
  assign n10210 = n10206 & ~n10208 ;
  assign n10211 = ~n10209 & ~n10210 ;
  assign n10214 = n10211 & ~x36 ;
  assign n10215 = ~n10213 & ~n10214 ;
  assign n10216 = ~n10129 & ~n10131 ;
  assign n10217 = ~n169 & ~n369 ;
  assign n10218 = ~n230 & n10217 ;
  assign n10219 = ~n335 & n10218 ;
  assign n10220 = ~n93 & n10219 ;
  assign n10221 = n131 & n10220 ;
  assign n10222 = n7806 & n10221 ;
  assign n10223 = n286 & n10222 ;
  assign n10224 = n2153 & n10223 ;
  assign n10225 = n955 & n10224 ;
  assign n10226 = n3674 & n10225 ;
  assign n10227 = ~n171 & n10226 ;
  assign n10228 = ~n318 & n10227 ;
  assign n10229 = ~n232 & n10228 ;
  assign n10230 = ~n144 & n10229 ;
  assign n10231 = ~n117 & n10230 ;
  assign n10232 = ~n445 & n10231 ;
  assign n10233 = ~n326 & n10232 ;
  assign n10234 = ~n10122 & ~n10125 ;
  assign n10235 = n2643 & n7700 ;
  assign n10236 = n2751 & ~n3603 ;
  assign n10237 = n2641 & n3725 ;
  assign n10238 = ~n10236 & ~n10237 ;
  assign n10239 = ~n10235 & n10238 ;
  assign n10240 = n2649 & n7712 ;
  assign n10241 = n10239 & ~n10240 ;
  assign n10242 = ~n500 & ~n10241 ;
  assign n10243 = ~n10241 & ~n10242 ;
  assign n10244 = ~n500 & ~n10242 ;
  assign n10245 = ~n10243 & ~n10244 ;
  assign n10246 = n644 & n10110 ;
  assign n10247 = ~n644 & ~n10110 ;
  assign n10248 = ~n10246 & ~n10247 ;
  assign n10249 = ~n500 & n3247 ;
  assign n10250 = n10248 & n10249 ;
  assign n10251 = ~n10248 & ~n10249 ;
  assign n10252 = ~n10250 & ~n10251 ;
  assign n10253 = ~n10245 & n10252 ;
  assign n10254 = ~n10245 & ~n10253 ;
  assign n10255 = n10252 & ~n10253 ;
  assign n10256 = ~n10254 & ~n10255 ;
  assign n10257 = ~n10116 & n10256 ;
  assign n10258 = n10116 & ~n10256 ;
  assign n10259 = ~n10257 & ~n10258 ;
  assign n10260 = ~n10107 & ~n10118 ;
  assign n10261 = ~n10104 & ~n10260 ;
  assign n10262 = ~n10259 & ~n10261 ;
  assign n10263 = n10259 & n10261 ;
  assign n10264 = ~n10262 & ~n10263 ;
  assign n10265 = ~n10234 & n10264 ;
  assign n10266 = n10234 & ~n10264 ;
  assign n10267 = ~n10265 & ~n10266 ;
  assign n10268 = ~n10233 & n10267 ;
  assign n10269 = n10233 & ~n10267 ;
  assign n10270 = ~n10216 & ~n10269 ;
  assign n10271 = ~n10268 & n10270 ;
  assign n10272 = ~n10216 & ~n10271 ;
  assign n10273 = ~n10268 & ~n10271 ;
  assign n10274 = ~n10269 & n10273 ;
  assign n10275 = ~n10272 & ~n10274 ;
  assign n10276 = ~n10135 & n10275 ;
  assign n10277 = n10135 & ~n10275 ;
  assign n10278 = ~n10276 & ~n10277 ;
  assign n10279 = ~n10136 & n10137 ;
  assign n10280 = ~n7831 & ~n10279 ;
  assign n10281 = ~n10278 & n10280 ;
  assign n10282 = n10278 & ~n10280 ;
  assign n10283 = ~n10281 & ~n10282 ;
  assign n10353 = ~n10283 & x37 ;
  assign n10284 = ~n10199 & ~n10201 ;
  assign n10285 = ~n3994 & ~n4194 ;
  assign n10286 = ~n4055 & n10285 ;
  assign n10287 = ~n4160 & n10286 ;
  assign n10288 = ~n3918 & n10287 ;
  assign n10289 = n3956 & n10288 ;
  assign n10290 = n7963 & n10289 ;
  assign n10291 = n4111 & n10290 ;
  assign n10292 = n5978 & n10291 ;
  assign n10293 = n4780 & n10292 ;
  assign n10294 = n7499 & n10293 ;
  assign n10295 = ~n3996 & n10294 ;
  assign n10296 = ~n4143 & n10295 ;
  assign n10297 = ~n4057 & n10296 ;
  assign n10298 = ~n3969 & n10297 ;
  assign n10299 = ~n3942 & n10298 ;
  assign n10300 = ~n4270 & n10299 ;
  assign n10301 = ~n4151 & n10300 ;
  assign n10302 = ~n10192 & ~n10195 ;
  assign n10303 = n6468 & n7857 ;
  assign n10304 = n6576 & ~n7428 ;
  assign n10305 = n6466 & n7550 ;
  assign n10306 = ~n10304 & ~n10305 ;
  assign n10307 = ~n10303 & n10306 ;
  assign n10308 = n6474 & n7869 ;
  assign n10309 = n10307 & ~n10308 ;
  assign n10310 = ~n4325 & ~n10309 ;
  assign n10311 = ~n10309 & ~n10310 ;
  assign n10312 = ~n4325 & ~n10310 ;
  assign n10313 = ~n10311 & ~n10312 ;
  assign n10314 = n4469 & n10180 ;
  assign n10315 = ~n4469 & ~n10180 ;
  assign n10316 = ~n10314 & ~n10315 ;
  assign n10317 = ~n4325 & n7072 ;
  assign n10318 = n10316 & n10317 ;
  assign n10319 = ~n10316 & ~n10317 ;
  assign n10320 = ~n10318 & ~n10319 ;
  assign n10321 = ~n10313 & n10320 ;
  assign n10322 = ~n10313 & ~n10321 ;
  assign n10323 = n10320 & ~n10321 ;
  assign n10324 = ~n10322 & ~n10323 ;
  assign n10325 = ~n10186 & n10324 ;
  assign n10326 = n10186 & ~n10324 ;
  assign n10327 = ~n10325 & ~n10326 ;
  assign n10328 = ~n10177 & ~n10188 ;
  assign n10329 = ~n10174 & ~n10328 ;
  assign n10330 = ~n10327 & ~n10329 ;
  assign n10331 = n10327 & n10329 ;
  assign n10332 = ~n10330 & ~n10331 ;
  assign n10333 = ~n10302 & n10332 ;
  assign n10334 = n10302 & ~n10332 ;
  assign n10335 = ~n10333 & ~n10334 ;
  assign n10336 = ~n10301 & n10335 ;
  assign n10337 = n10301 & ~n10335 ;
  assign n10338 = ~n10284 & ~n10337 ;
  assign n10339 = ~n10336 & n10338 ;
  assign n10340 = ~n10284 & ~n10339 ;
  assign n10341 = ~n10336 & ~n10339 ;
  assign n10342 = ~n10337 & n10341 ;
  assign n10343 = ~n10340 & ~n10342 ;
  assign n10344 = ~n10205 & n10343 ;
  assign n10345 = n10205 & ~n10343 ;
  assign n10346 = ~n10344 & ~n10345 ;
  assign n10347 = ~n10206 & n10207 ;
  assign n10348 = ~n7831 & ~n10347 ;
  assign n10349 = ~n10346 & n10348 ;
  assign n10350 = n10346 & ~n10348 ;
  assign n10351 = ~n10349 & ~n10350 ;
  assign n10354 = n10351 & ~x37 ;
  assign n10355 = ~n10353 & ~n10354 ;
  assign n10356 = n2342 & n2408 ;
  assign n10357 = n448 & n10356 ;
  assign n10358 = n942 & n10357 ;
  assign n10359 = n2165 & n10358 ;
  assign n10360 = n1432 & n10359 ;
  assign n10361 = n958 & n10360 ;
  assign n10362 = n3234 & n10361 ;
  assign n10363 = ~n113 & n10362 ;
  assign n10364 = ~n151 & n10363 ;
  assign n10365 = ~n102 & n10364 ;
  assign n10366 = ~n318 & n10365 ;
  assign n10367 = ~n345 & n10366 ;
  assign n10368 = ~n311 & n10367 ;
  assign n10369 = ~n481 & n10368 ;
  assign n10370 = ~n10262 & ~n10265 ;
  assign n10371 = ~n10116 & ~n10256 ;
  assign n10372 = ~n10253 & ~n10371 ;
  assign n10373 = ~n500 & ~n3603 ;
  assign n10374 = ~n10246 & ~n10250 ;
  assign n10375 = ~n10373 & ~n10374 ;
  assign n10376 = ~n10373 & ~n10375 ;
  assign n10377 = ~n10374 & ~n10375 ;
  assign n10378 = ~n10376 & ~n10377 ;
  assign n10379 = n2751 & n3725 ;
  assign n10380 = n2641 & n7700 ;
  assign n10381 = ~n10379 & ~n10380 ;
  assign n10382 = ~n2649 & n10381 ;
  assign n10383 = ~n8018 & n10381 ;
  assign n10384 = ~n10382 & ~n10383 ;
  assign n10385 = n500 & ~n10384 ;
  assign n10386 = ~n500 & n10384 ;
  assign n10387 = ~n10385 & ~n10386 ;
  assign n10388 = ~n10378 & n10387 ;
  assign n10389 = n10378 & ~n10387 ;
  assign n10390 = ~n10388 & ~n10389 ;
  assign n10391 = ~n10372 & n10390 ;
  assign n10392 = n10372 & ~n10390 ;
  assign n10393 = ~n10391 & ~n10392 ;
  assign n10394 = ~n10370 & n10393 ;
  assign n10395 = n10370 & ~n10393 ;
  assign n10396 = ~n10394 & ~n10395 ;
  assign n10397 = n10369 & ~n10396 ;
  assign n10398 = ~n10369 & n10396 ;
  assign n10399 = ~n10397 & ~n10398 ;
  assign n10400 = ~n10273 & n10399 ;
  assign n10401 = n10273 & ~n10399 ;
  assign n10402 = ~n10400 & ~n10401 ;
  assign n10403 = ~n10277 & ~n10402 ;
  assign n10404 = n10277 & n10402 ;
  assign n10405 = ~n10403 & ~n10404 ;
  assign n10406 = ~n10278 & n10279 ;
  assign n10407 = ~n7831 & ~n10406 ;
  assign n10408 = ~n10405 & n10407 ;
  assign n10409 = n10405 & ~n10407 ;
  assign n10410 = ~n10408 & ~n10409 ;
  assign n10467 = ~n10410 & x38 ;
  assign n10411 = n6167 & n6233 ;
  assign n10412 = n4273 & n10411 ;
  assign n10413 = n4767 & n10412 ;
  assign n10414 = n5990 & n10413 ;
  assign n10415 = n5257 & n10414 ;
  assign n10416 = n4783 & n10415 ;
  assign n10417 = n7059 & n10416 ;
  assign n10418 = ~n3938 & n10417 ;
  assign n10419 = ~n3976 & n10418 ;
  assign n10420 = ~n3927 & n10419 ;
  assign n10421 = ~n4143 & n10420 ;
  assign n10422 = ~n4170 & n10421 ;
  assign n10423 = ~n4136 & n10422 ;
  assign n10424 = ~n4306 & n10423 ;
  assign n10425 = ~n10330 & ~n10333 ;
  assign n10426 = ~n10186 & ~n10324 ;
  assign n10427 = ~n10321 & ~n10426 ;
  assign n10428 = ~n4325 & ~n7428 ;
  assign n10429 = ~n10314 & ~n10318 ;
  assign n10430 = ~n10428 & ~n10429 ;
  assign n10431 = ~n10428 & ~n10430 ;
  assign n10432 = ~n10429 & ~n10430 ;
  assign n10433 = ~n10431 & ~n10432 ;
  assign n10434 = n6576 & n7550 ;
  assign n10435 = n6466 & n7857 ;
  assign n10436 = ~n10434 & ~n10435 ;
  assign n10437 = ~n6474 & n10436 ;
  assign n10438 = ~n8149 & n10436 ;
  assign n10439 = ~n10437 & ~n10438 ;
  assign n10440 = n4325 & ~n10439 ;
  assign n10441 = ~n4325 & n10439 ;
  assign n10442 = ~n10440 & ~n10441 ;
  assign n10443 = ~n10433 & n10442 ;
  assign n10444 = n10433 & ~n10442 ;
  assign n10445 = ~n10443 & ~n10444 ;
  assign n10446 = ~n10427 & n10445 ;
  assign n10447 = n10427 & ~n10445 ;
  assign n10448 = ~n10446 & ~n10447 ;
  assign n10449 = ~n10425 & n10448 ;
  assign n10450 = n10425 & ~n10448 ;
  assign n10451 = ~n10449 & ~n10450 ;
  assign n10452 = n10424 & ~n10451 ;
  assign n10453 = ~n10424 & n10451 ;
  assign n10454 = ~n10452 & ~n10453 ;
  assign n10455 = ~n10341 & n10454 ;
  assign n10456 = n10341 & ~n10454 ;
  assign n10457 = ~n10455 & ~n10456 ;
  assign n10458 = ~n10345 & ~n10457 ;
  assign n10459 = n10345 & n10457 ;
  assign n10460 = ~n10458 & ~n10459 ;
  assign n10461 = ~n10346 & n10347 ;
  assign n10462 = ~n7831 & ~n10461 ;
  assign n10463 = ~n10460 & n10462 ;
  assign n10464 = n10460 & ~n10462 ;
  assign n10465 = ~n10463 & ~n10464 ;
  assign n10468 = n10465 & ~x38 ;
  assign n10469 = ~n10467 & ~n10468 ;
  assign n10470 = ~n10398 & ~n10400 ;
  assign n10471 = ~n312 & n1120 ;
  assign n10472 = ~n303 & n10471 ;
  assign n10473 = ~n229 & n10472 ;
  assign n10474 = n945 & n10473 ;
  assign n10475 = n319 & n10474 ;
  assign n10476 = n10076 & n10475 ;
  assign n10477 = n2350 & n10476 ;
  assign n10478 = n1090 & n10477 ;
  assign n10479 = ~n102 & n10478 ;
  assign n10480 = ~n201 & n10479 ;
  assign n10481 = ~n192 & n10480 ;
  assign n10482 = ~n331 & n10481 ;
  assign n10483 = ~n481 & n10482 ;
  assign n10484 = ~n711 & n10483 ;
  assign n10485 = n2751 & n7700 ;
  assign n10486 = n2649 & n8016 ;
  assign n10487 = ~n10485 & ~n10486 ;
  assign n10488 = ~n500 & ~n10487 ;
  assign n10489 = ~n10487 & ~n10488 ;
  assign n10490 = ~n500 & ~n10488 ;
  assign n10491 = ~n10489 & ~n10490 ;
  assign n10492 = ~n500 & n3734 ;
  assign n10493 = ~n10491 & ~n10492 ;
  assign n10494 = ~n10491 & ~n10493 ;
  assign n10495 = ~n10492 & ~n10493 ;
  assign n10496 = ~n10494 & ~n10495 ;
  assign n10497 = ~n10375 & ~n10388 ;
  assign n10498 = n10496 & n10497 ;
  assign n10499 = ~n10496 & ~n10497 ;
  assign n10500 = ~n10498 & ~n10499 ;
  assign n10501 = ~n10391 & ~n10394 ;
  assign n10502 = ~n10500 & n10501 ;
  assign n10503 = n10500 & ~n10501 ;
  assign n10504 = ~n10502 & ~n10503 ;
  assign n10505 = ~n10484 & n10504 ;
  assign n10506 = n10484 & ~n10504 ;
  assign n10507 = ~n10470 & ~n10506 ;
  assign n10508 = ~n10505 & n10507 ;
  assign n10509 = ~n10470 & ~n10508 ;
  assign n10510 = ~n10505 & ~n10508 ;
  assign n10511 = ~n10506 & n10510 ;
  assign n10512 = ~n10509 & ~n10511 ;
  assign n10513 = ~n10404 & n10512 ;
  assign n10514 = n10404 & ~n10512 ;
  assign n10515 = ~n10513 & ~n10514 ;
  assign n10516 = ~n10405 & n10406 ;
  assign n10517 = ~n7831 & ~n10516 ;
  assign n10518 = ~n10515 & n10517 ;
  assign n10519 = n10515 & ~n10517 ;
  assign n10520 = ~n10518 & ~n10519 ;
  assign n10573 = ~n10520 & x39 ;
  assign n10521 = ~n10453 & ~n10455 ;
  assign n10522 = ~n4137 & n4945 ;
  assign n10523 = ~n4128 & n10522 ;
  assign n10524 = ~n4054 & n10523 ;
  assign n10525 = n4770 & n10524 ;
  assign n10526 = n4144 & n10525 ;
  assign n10527 = n10146 & n10526 ;
  assign n10528 = n6175 & n10527 ;
  assign n10529 = n4915 & n10528 ;
  assign n10530 = ~n3927 & n10529 ;
  assign n10531 = ~n4026 & n10530 ;
  assign n10532 = ~n4017 & n10531 ;
  assign n10533 = ~n4156 & n10532 ;
  assign n10534 = ~n4306 & n10533 ;
  assign n10535 = ~n4536 & n10534 ;
  assign n10536 = n6576 & n7857 ;
  assign n10537 = n6474 & n8147 ;
  assign n10538 = ~n10536 & ~n10537 ;
  assign n10539 = ~n4325 & ~n10538 ;
  assign n10540 = ~n10538 & ~n10539 ;
  assign n10541 = ~n4325 & ~n10539 ;
  assign n10542 = ~n10540 & ~n10541 ;
  assign n10543 = ~n4325 & n7559 ;
  assign n10544 = ~n10542 & ~n10543 ;
  assign n10545 = ~n10542 & ~n10544 ;
  assign n10546 = ~n10543 & ~n10544 ;
  assign n10547 = ~n10545 & ~n10546 ;
  assign n10548 = ~n10430 & ~n10443 ;
  assign n10549 = n10547 & n10548 ;
  assign n10550 = ~n10547 & ~n10548 ;
  assign n10551 = ~n10549 & ~n10550 ;
  assign n10552 = ~n10446 & ~n10449 ;
  assign n10553 = ~n10551 & n10552 ;
  assign n10554 = n10551 & ~n10552 ;
  assign n10555 = ~n10553 & ~n10554 ;
  assign n10556 = ~n10535 & n10555 ;
  assign n10557 = n10535 & ~n10555 ;
  assign n10558 = ~n10521 & ~n10557 ;
  assign n10559 = ~n10556 & n10558 ;
  assign n10560 = ~n10521 & ~n10559 ;
  assign n10561 = ~n10556 & ~n10559 ;
  assign n10562 = ~n10557 & n10561 ;
  assign n10563 = ~n10560 & ~n10562 ;
  assign n10564 = ~n10459 & n10563 ;
  assign n10565 = n10459 & ~n10563 ;
  assign n10566 = ~n10564 & ~n10565 ;
  assign n10567 = ~n10460 & n10461 ;
  assign n10568 = ~n7831 & ~n10567 ;
  assign n10569 = ~n10566 & n10568 ;
  assign n10570 = n10566 & ~n10568 ;
  assign n10571 = ~n10569 & ~n10570 ;
  assign n10574 = n10571 & ~x39 ;
  assign n10575 = ~n10573 & ~n10574 ;
  assign n10576 = n613 & n2288 ;
  assign n10577 = n2227 & n10576 ;
  assign n10578 = n10220 & n10577 ;
  assign n10579 = n208 & n10578 ;
  assign n10580 = n450 & n10579 ;
  assign n10581 = n3677 & n10580 ;
  assign n10582 = ~n183 & n10581 ;
  assign n10583 = ~n422 & n10582 ;
  assign n10584 = ~n452 & n10583 ;
  assign n10585 = ~n10499 & ~n10503 ;
  assign n10586 = n3725 & ~n10373 ;
  assign n10587 = ~n500 & n10586 ;
  assign n10588 = ~n10493 & ~n10587 ;
  assign n10589 = ~n10585 & n10588 ;
  assign n10590 = n10585 & ~n10588 ;
  assign n10591 = ~n10589 & ~n10590 ;
  assign n10592 = n7700 & ~n10373 ;
  assign n10593 = ~n7700 & n10373 ;
  assign n10594 = ~n10592 & ~n10593 ;
  assign n10595 = ~n500 & n10594 ;
  assign n10596 = n10591 & ~n10595 ;
  assign n10597 = ~n10591 & n10595 ;
  assign n10598 = ~n10596 & ~n10597 ;
  assign n10599 = ~n10584 & ~n10598 ;
  assign n10600 = n10584 & n10598 ;
  assign n10601 = ~n10510 & ~n10600 ;
  assign n10602 = ~n10599 & n10601 ;
  assign n10603 = ~n10510 & ~n10602 ;
  assign n10604 = ~n10599 & ~n10602 ;
  assign n10605 = ~n10600 & n10604 ;
  assign n10606 = ~n10603 & ~n10605 ;
  assign n10607 = ~n10514 & n10606 ;
  assign n10608 = n10514 & ~n10606 ;
  assign n10609 = ~n10607 & ~n10608 ;
  assign n10610 = ~n10515 & n10516 ;
  assign n10611 = ~n7831 & ~n10610 ;
  assign n10612 = ~n10609 & n10611 ;
  assign n10613 = n10609 & ~n10611 ;
  assign n10614 = ~n10612 & ~n10613 ;
  assign n10655 = ~n10614 & x40 ;
  assign n10615 = n4438 & n6113 ;
  assign n10616 = n6052 & n10615 ;
  assign n10617 = n10288 & n10616 ;
  assign n10618 = n4033 & n10617 ;
  assign n10619 = n4275 & n10618 ;
  assign n10620 = n7502 & n10619 ;
  assign n10621 = ~n4008 & n10620 ;
  assign n10622 = ~n4247 & n10621 ;
  assign n10623 = ~n4277 & n10622 ;
  assign n10624 = ~n10550 & ~n10554 ;
  assign n10625 = n7550 & ~n10428 ;
  assign n10626 = ~n4325 & n10625 ;
  assign n10627 = ~n10544 & ~n10626 ;
  assign n10628 = ~n10624 & n10627 ;
  assign n10629 = n10624 & ~n10627 ;
  assign n10630 = ~n10628 & ~n10629 ;
  assign n10631 = n7857 & ~n10428 ;
  assign n10632 = ~n7857 & n10428 ;
  assign n10633 = ~n10631 & ~n10632 ;
  assign n10634 = ~n4325 & n10633 ;
  assign n10635 = n10630 & ~n10634 ;
  assign n10636 = ~n10630 & n10634 ;
  assign n10637 = ~n10635 & ~n10636 ;
  assign n10638 = ~n10623 & ~n10637 ;
  assign n10639 = n10623 & n10637 ;
  assign n10640 = ~n10561 & ~n10639 ;
  assign n10641 = ~n10638 & n10640 ;
  assign n10642 = ~n10561 & ~n10641 ;
  assign n10643 = ~n10638 & ~n10641 ;
  assign n10644 = ~n10639 & n10643 ;
  assign n10645 = ~n10642 & ~n10644 ;
  assign n10646 = ~n10565 & n10645 ;
  assign n10647 = n10565 & ~n10645 ;
  assign n10648 = ~n10646 & ~n10647 ;
  assign n10649 = ~n10566 & n10567 ;
  assign n10650 = ~n7831 & ~n10649 ;
  assign n10651 = ~n10648 & n10650 ;
  assign n10652 = n10648 & ~n10650 ;
  assign n10653 = ~n10651 & ~n10652 ;
  assign n10656 = n10653 & ~x40 ;
  assign n10657 = ~n10655 & ~n10656 ;
  assign n10658 = n133 & n750 ;
  assign n10659 = n881 & n10658 ;
  assign n10660 = n234 & n10659 ;
  assign n10661 = n3218 & n10660 ;
  assign n10662 = n546 & n10661 ;
  assign n10663 = n955 & n10662 ;
  assign n10664 = ~n114 & n10663 ;
  assign n10665 = ~n182 & n10664 ;
  assign n10666 = ~n272 & n10665 ;
  assign n10667 = ~n343 & n10666 ;
  assign n10668 = ~n190 & n10667 ;
  assign n10669 = ~n10604 & ~n10668 ;
  assign n10670 = n10604 & n10668 ;
  assign n10671 = ~n10669 & ~n10670 ;
  assign n10672 = ~n10608 & n10671 ;
  assign n10673 = n10608 & ~n10671 ;
  assign n10674 = ~n10672 & ~n10673 ;
  assign n10675 = ~n10609 & n10610 ;
  assign n10676 = ~n7831 & ~n10675 ;
  assign n10677 = ~n10674 & n10676 ;
  assign n10678 = n10674 & ~n10676 ;
  assign n10679 = ~n10677 & ~n10678 ;
  assign n10703 = n10679 & x41 ;
  assign n10680 = n3958 & n4575 ;
  assign n10681 = n4706 & n10680 ;
  assign n10682 = n4059 & n10681 ;
  assign n10683 = n7043 & n10682 ;
  assign n10684 = n4371 & n10683 ;
  assign n10685 = n4780 & n10684 ;
  assign n10686 = ~n3939 & n10685 ;
  assign n10687 = ~n4007 & n10686 ;
  assign n10688 = ~n4097 & n10687 ;
  assign n10689 = ~n4168 & n10688 ;
  assign n10690 = ~n4015 & n10689 ;
  assign n10691 = ~n10643 & ~n10690 ;
  assign n10692 = n10643 & n10690 ;
  assign n10693 = ~n10691 & ~n10692 ;
  assign n10694 = ~n10647 & n10693 ;
  assign n10695 = n10647 & ~n10693 ;
  assign n10696 = ~n10694 & ~n10695 ;
  assign n10697 = ~n10648 & n10649 ;
  assign n10698 = ~n7831 & ~n10697 ;
  assign n10699 = ~n10696 & n10698 ;
  assign n10700 = n10696 & ~n10698 ;
  assign n10701 = ~n10699 & ~n10700 ;
  assign n10704 = ~n10701 & ~x41 ;
  assign n10705 = ~n10703 & ~n10704 ;
  assign n10706 = n10608 & n10671 ;
  assign n10707 = n563 & n2145 ;
  assign n10708 = n583 & n10707 ;
  assign n10709 = n1127 & n10708 ;
  assign n10710 = n1083 & n10709 ;
  assign n10711 = n961 & n10710 ;
  assign n10712 = n3650 & n10711 ;
  assign n10713 = ~n151 & n10712 ;
  assign n10714 = ~n202 & n10713 ;
  assign n10715 = ~n182 & n10714 ;
  assign n10716 = ~n332 & n10715 ;
  assign n10717 = ~n213 & n10716 ;
  assign n10718 = n10669 & ~n10717 ;
  assign n10719 = ~n10669 & n10717 ;
  assign n10720 = ~n10718 & ~n10719 ;
  assign n10721 = ~n10706 & ~n10720 ;
  assign n10722 = n10706 & ~n10719 ;
  assign n10723 = ~n10721 & ~n10722 ;
  assign n10724 = n10674 & n10675 ;
  assign n10725 = ~n7831 & ~n10724 ;
  assign n10726 = ~n10723 & n10725 ;
  assign n10727 = n10723 & ~n10725 ;
  assign n10728 = ~n10726 & ~n10727 ;
  assign n10753 = ~n10728 & x42 ;
  assign n10729 = n10647 & n10693 ;
  assign n10730 = n4388 & n5970 ;
  assign n10731 = n4408 & n10730 ;
  assign n10732 = n4952 & n10731 ;
  assign n10733 = n4908 & n10732 ;
  assign n10734 = n4786 & n10733 ;
  assign n10735 = n7475 & n10734 ;
  assign n10736 = ~n3976 & n10735 ;
  assign n10737 = ~n4027 & n10736 ;
  assign n10738 = ~n4007 & n10737 ;
  assign n10739 = ~n4157 & n10738 ;
  assign n10740 = ~n4038 & n10739 ;
  assign n10741 = n10691 & ~n10740 ;
  assign n10742 = ~n10691 & n10740 ;
  assign n10743 = ~n10741 & ~n10742 ;
  assign n10744 = ~n10729 & ~n10743 ;
  assign n10745 = n10729 & ~n10742 ;
  assign n10746 = ~n10744 & ~n10745 ;
  assign n10747 = n10696 & n10697 ;
  assign n10748 = ~n7831 & ~n10747 ;
  assign n10749 = ~n10746 & n10748 ;
  assign n10750 = n10746 & ~n10748 ;
  assign n10751 = ~n10749 & ~n10750 ;
  assign n10754 = n10751 & ~x42 ;
  assign n10755 = ~n10753 & ~n10754 ;
  assign n10756 = n8724 & n10473 ;
  assign n10757 = n348 & n10756 ;
  assign n10758 = n2515 & n10757 ;
  assign n10759 = n913 & n10758 ;
  assign n10760 = ~n119 & n10759 ;
  assign n10761 = ~n127 & n10760 ;
  assign n10762 = ~n183 & n10761 ;
  assign n10763 = ~n115 & n10762 ;
  assign n10764 = ~n421 & n10763 ;
  assign n10765 = ~n273 & n10764 ;
  assign n10766 = ~n181 & n10765 ;
  assign n10767 = ~n10718 & n10766 ;
  assign n10768 = n10718 & ~n10766 ;
  assign n10769 = ~n10767 & ~n10768 ;
  assign n10770 = ~n10722 & ~n10769 ;
  assign n10771 = n10722 & n10769 ;
  assign n10772 = ~n10770 & ~n10771 ;
  assign n10773 = ~n10723 & n10724 ;
  assign n10774 = ~n7831 & ~n10773 ;
  assign n10775 = ~n10772 & n10774 ;
  assign n10776 = n10772 & ~n10774 ;
  assign n10777 = ~n10775 & ~n10776 ;
  assign n10801 = ~n10777 & x43 ;
  assign n10778 = n8839 & n10524 ;
  assign n10779 = n4173 & n10778 ;
  assign n10780 = n6340 & n10779 ;
  assign n10781 = n4738 & n10780 ;
  assign n10782 = ~n3944 & n10781 ;
  assign n10783 = ~n3952 & n10782 ;
  assign n10784 = ~n4008 & n10783 ;
  assign n10785 = ~n3940 & n10784 ;
  assign n10786 = ~n4246 & n10785 ;
  assign n10787 = ~n4098 & n10786 ;
  assign n10788 = ~n4006 & n10787 ;
  assign n10789 = ~n10741 & n10788 ;
  assign n10790 = n10741 & ~n10788 ;
  assign n10791 = ~n10789 & ~n10790 ;
  assign n10792 = ~n10745 & ~n10791 ;
  assign n10793 = n10745 & n10791 ;
  assign n10794 = ~n10792 & ~n10793 ;
  assign n10795 = ~n10746 & n10747 ;
  assign n10796 = ~n7831 & ~n10795 ;
  assign n10797 = ~n10794 & n10796 ;
  assign n10798 = n10794 & ~n10796 ;
  assign n10799 = ~n10797 & ~n10798 ;
  assign n10802 = n10799 & ~x43 ;
  assign n10803 = ~n10801 & ~n10802 ;
  assign n10804 = n164 & n434 ;
  assign n10805 = n974 & n10804 ;
  assign n10806 = n477 & n10805 ;
  assign n10807 = n9397 & n10806 ;
  assign n10808 = n344 & n10807 ;
  assign n10809 = ~n169 & n10808 ;
  assign n10810 = ~n202 & n10809 ;
  assign n10811 = ~n287 & n10810 ;
  assign n10812 = ~n193 & n10811 ;
  assign n10813 = ~n188 & n10812 ;
  assign n10814 = ~n187 & n10813 ;
  assign n10815 = ~n529 & n10814 ;
  assign n10816 = n10768 & ~n10815 ;
  assign n10817 = ~n10768 & n10815 ;
  assign n10818 = ~n10816 & ~n10817 ;
  assign n10819 = ~n10771 & ~n10818 ;
  assign n10820 = n10771 & ~n10817 ;
  assign n10821 = ~n10819 & ~n10820 ;
  assign n10822 = ~n10772 & n10773 ;
  assign n10823 = ~n7831 & ~n10822 ;
  assign n10824 = ~n10821 & n10823 ;
  assign n10825 = n10821 & ~n10823 ;
  assign n10826 = ~n10824 & ~n10825 ;
  assign n10851 = ~n10826 & x44 ;
  assign n10827 = n3989 & n4259 ;
  assign n10828 = n4799 & n10827 ;
  assign n10829 = n4302 & n10828 ;
  assign n10830 = n9497 & n10829 ;
  assign n10831 = n4169 & n10830 ;
  assign n10832 = ~n3994 & n10831 ;
  assign n10833 = ~n4027 & n10832 ;
  assign n10834 = ~n4112 & n10833 ;
  assign n10835 = ~n4018 & n10834 ;
  assign n10836 = ~n4013 & n10835 ;
  assign n10837 = ~n4012 & n10836 ;
  assign n10838 = ~n4354 & n10837 ;
  assign n10839 = n10790 & ~n10838 ;
  assign n10840 = ~n10790 & n10838 ;
  assign n10841 = ~n10839 & ~n10840 ;
  assign n10842 = ~n10793 & ~n10841 ;
  assign n10843 = n10793 & ~n10840 ;
  assign n10844 = ~n10842 & ~n10843 ;
  assign n10845 = ~n10794 & n10795 ;
  assign n10846 = ~n7831 & ~n10845 ;
  assign n10847 = ~n10844 & n10846 ;
  assign n10848 = n10844 & ~n10846 ;
  assign n10849 = ~n10847 & ~n10848 ;
  assign n10852 = n10849 & ~x44 ;
  assign n10853 = ~n10851 & ~n10852 ;
  assign n10854 = n464 & n3592 ;
  assign n10855 = n419 & n10854 ;
  assign n10856 = ~n318 & n10855 ;
  assign n10857 = ~n335 & n10856 ;
  assign n10858 = ~n10816 & n10857 ;
  assign n10859 = n10816 & ~n10857 ;
  assign n10860 = ~n10858 & ~n10859 ;
  assign n10861 = ~n10820 & ~n10860 ;
  assign n10862 = n10820 & n10860 ;
  assign n10863 = ~n10861 & ~n10862 ;
  assign n10864 = ~n10821 & n10822 ;
  assign n10865 = ~n7831 & ~n10864 ;
  assign n10866 = ~n10863 & n10865 ;
  assign n10867 = n10863 & ~n10865 ;
  assign n10868 = ~n10866 & ~n10867 ;
  assign n10885 = ~n10868 & x45 ;
  assign n10869 = n4289 & n7417 ;
  assign n10870 = n4244 & n10869 ;
  assign n10871 = ~n4143 & n10870 ;
  assign n10872 = ~n4160 & n10871 ;
  assign n10873 = ~n10839 & n10872 ;
  assign n10874 = n10839 & ~n10872 ;
  assign n10875 = ~n10873 & ~n10874 ;
  assign n10876 = ~n10843 & ~n10875 ;
  assign n10877 = n10843 & n10875 ;
  assign n10878 = ~n10876 & ~n10877 ;
  assign n10879 = ~n10844 & n10845 ;
  assign n10880 = ~n7831 & ~n10879 ;
  assign n10881 = ~n10878 & n10880 ;
  assign n10882 = n10878 & ~n10880 ;
  assign n10883 = ~n10881 & ~n10882 ;
  assign n10886 = n10883 & ~x45 ;
  assign n10887 = ~n10885 & ~n10886 ;
  assign n10888 = n419 & n492 ;
  assign n10889 = n10859 & ~n10888 ;
  assign n10890 = ~n10859 & n10888 ;
  assign n10891 = ~n10889 & ~n10890 ;
  assign n10892 = ~n10862 & ~n10891 ;
  assign n10893 = n10862 & ~n10890 ;
  assign n10894 = ~n10892 & ~n10893 ;
  assign n10895 = ~n10863 & n10864 ;
  assign n10896 = ~n7831 & ~n10895 ;
  assign n10897 = ~n10894 & n10896 ;
  assign n10898 = n10894 & ~n10896 ;
  assign n10899 = ~n10897 & ~n10898 ;
  assign n10913 = ~n10899 & x46 ;
  assign n10900 = n4244 & n4317 ;
  assign n10901 = n10874 & ~n10900 ;
  assign n10902 = ~n10874 & n10900 ;
  assign n10903 = ~n10901 & ~n10902 ;
  assign n10904 = ~n10877 & ~n10903 ;
  assign n10905 = n10877 & ~n10902 ;
  assign n10906 = ~n10904 & ~n10905 ;
  assign n10907 = ~n10878 & n10879 ;
  assign n10908 = ~n7831 & ~n10907 ;
  assign n10909 = ~n10906 & n10908 ;
  assign n10910 = n10906 & ~n10908 ;
  assign n10911 = ~n10909 & ~n10910 ;
  assign n10914 = n10911 & ~x46 ;
  assign n10915 = ~n10913 & ~n10914 ;
  assign n10916 = ~x22 & n46 ;
  assign n10917 = ~n10889 & ~n10893 ;
  assign n10918 = n10889 & n10893 ;
  assign n10919 = ~n10917 & ~n10918 ;
  assign n10920 = ~n10894 & n10895 ;
  assign n10921 = ~n7831 & ~n10920 ;
  assign n10922 = n10919 & ~n10921 ;
  assign n10923 = ~n10919 & n10921 ;
  assign n10924 = ~n10922 & ~n10923 ;
  assign n10925 = ~n10916 & n10924 ;
  assign n10937 = ~n10925 & x47 ;
  assign n10926 = x22 & n3871 ;
  assign n10927 = ~n10901 & ~n10905 ;
  assign n10928 = n10901 & n10905 ;
  assign n10929 = ~n10927 & ~n10928 ;
  assign n10930 = ~n10906 & n10907 ;
  assign n10931 = ~n7831 & ~n10930 ;
  assign n10932 = n10929 & ~n10931 ;
  assign n10933 = ~n10929 & n10931 ;
  assign n10934 = ~n10932 & ~n10933 ;
  assign n10935 = ~n10926 & n10934 ;
  assign n10938 = n10935 & ~x47 ;
  assign n10939 = ~n10937 & ~n10938 ;
  assign n10940 = ~n10917 & n10920 ;
  assign n10941 = ~n10918 & ~n10920 ;
  assign n10942 = ~n10940 & ~n10941 ;
  assign n10943 = ~n10916 & n10942 ;
  assign n10944 = ~n7831 & ~n10943 ;
  assign n10951 = n10944 & x48 ;
  assign n10945 = ~n10927 & n10930 ;
  assign n10946 = ~n10928 & ~n10930 ;
  assign n10947 = ~n10945 & ~n10946 ;
  assign n10948 = ~n10926 & n10947 ;
  assign n10949 = ~n7831 & ~n10948 ;
  assign n10952 = ~n10949 & ~x48 ;
  assign n10953 = ~n10951 & ~n10952 ;
  assign y0 = ~n7678 ;
  assign y1 = ~n7993 ;
  assign y2 = ~n8259 ;
  assign y3 = ~n8499 ;
  assign y4 = ~n8721 ;
  assign y5 = ~n8955 ;
  assign y6 = ~n9185 ;
  assign y7 = ~n9387 ;
  assign y8 = ~n9591 ;
  assign y9 = ~n9761 ;
  assign y10 = ~n9939 ;
  assign y11 = ~n10071 ;
  assign y12 = ~n10215 ;
  assign y13 = ~n10355 ;
  assign y14 = ~n10469 ;
  assign y15 = ~n10575 ;
  assign y16 = ~n10657 ;
  assign y17 = ~n10705 ;
  assign y18 = ~n10755 ;
  assign y19 = ~n10803 ;
  assign y20 = ~n10853 ;
  assign y21 = ~n10887 ;
  assign y22 = ~n10915 ;
  assign y23 = ~n10939 ;
  assign y24 = ~n10953 ;
endmodule
