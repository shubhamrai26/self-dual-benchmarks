module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 , y256 , y257 , y258 , y259 , y260 , y261 , y262 , y263 , y264 , y265 , y266 , y267 , y268 , y269 , y270 , y271 , y272 , y273 , y274 , y275 , y276 , y277 , y278 , y279 , y280 , y281 , y282 , y283 , y284 , y285 , y286 , y287 , y288 , y289 , y290 , y291 , y292 , y293 , y294 , y295 , y296 , y297 , y298 , y299 , y300 , y301 , y302 , y303 , y304 , y305 , y306 , y307 , y308 , y309 , y310 , y311 , y312 , y313 , y314 , y315 , y316 , y317 , y318 , y319 , y320 , y321 , y322 , y323 , y324 , y325 , y326 , y327 , y328 , y329 , y330 , y331 , y332 , y333 , y334 , y335 , y336 , y337 , y338 , y339 , y340 , y341 , y342 , y343 , y344 , y345 , y346 , y347 , y348 , y349 , y350 , y351 , y352 , y353 , y354 , y355 , y356 , y357 , y358 , y359 , y360 , y361 , y362 , y363 , y364 , y365 , y366 , y367 , y368 , y369 , y370 , y371 , y372 , y373 , y374 , y375 , y376 , y377 , y378 , y379 , y380 , y381 , y382 , y383 , y384 , y385 , y386 , y387 , y388 , y389 , y390 , y391 , y392 , y393 , y394 , y395 , y396 , y397 , y398 , y399 , y400 , y401 , y402 , y403 , y404 , y405 , y406 , y407 , y408 , y409 , y410 , y411 , y412 , y413 , y414 , y415 , y416 , y417 , y418 , y419 , y420 , y421 , y422 , y423 , y424 , y425 , y426 , y427 , y428 , y429 , y430 , y431 , y432 , y433 , y434 , y435 , y436 , y437 , y438 , y439 , y440 , y441 , y442 , y443 , y444 , y445 , y446 , y447 , y448 , y449 , y450 , y451 , y452 , y453 , y454 , y455 , y456 , y457 , y458 , y459 , y460 , y461 , y462 , y463 , y464 , y465 , y466 , y467 , y468 , y469 , y470 , y471 , y472 , y473 , y474 , y475 , y476 , y477 , y478 , y479 , y480 , y481 , y482 , y483 , y484 , y485 , y486 , y487 , y488 , y489 , y490 , y491 , y492 , y493 , y494 , y495 , y496 , y497 , y498 , y499 , y500 , y501 , y502 , y503 , y504 , y505 , y506 , y507 , y508 , y509 , y510 , y511 , y512 , y513 , y514 , y515 , y516 , y517 , y518 , y519 , y520 , y521 , y522 , y523 , y524 , y525 , y526 , y527 , y528 , y529 , y530 , y531 , y532 , y533 , y534 , y535 , y536 , y537 , y538 , y539 , y540 , y541 , y542 , y543 , y544 , y545 , y546 , y547 , y548 , y549 , y550 , y551 , y552 , y553 , y554 , y555 , y556 , y557 , y558 , y559 , y560 , y561 , y562 , y563 , y564 , y565 , y566 , y567 , y568 , y569 , y570 , y571 , y572 , y573 , y574 , y575 , y576 , y577 , y578 , y579 , y580 , y581 , y582 , y583 , y584 , y585 , y586 , y587 , y588 , y589 , y590 , y591 , y592 , y593 , y594 , y595 , y596 , y597 , y598 , y599 , y600 , y601 , y602 , y603 , y604 , y605 , y606 , y607 , y608 , y609 , y610 , y611 , y612 , y613 , y614 , y615 , y616 , y617 , y618 , y619 , y620 , y621 , y622 , y623 , y624 , y625 , y626 , y627 , y628 , y629 , y630 , y631 , y632 , y633 , y634 , y635 , y636 , y637 , y638 , y639 , y640 , y641 , y642 , y643 , y644 , y645 , y646 , y647 , y648 , y649 , y650 , y651 , y652 , y653 , y654 , y655 , y656 , y657 , y658 , y659 , y660 , y661 , y662 , y663 , y664 , y665 , y666 , y667 , y668 , y669 , y670 , y671 , y672 , y673 , y674 , y675 , y676 , y677 , y678 , y679 , y680 , y681 , y682 , y683 , y684 , y685 , y686 , y687 , y688 , y689 , y690 , y691 , y692 , y693 , y694 , y695 , y696 , y697 , y698 , y699 , y700 , y701 , y702 , y703 , y704 , y705 , y706 , y707 , y708 , y709 , y710 , y711 , y712 , y713 , y714 , y715 , y716 , y717 , y718 , y719 , y720 , y721 , y722 , y723 , y724 , y725 , y726 , y727 , y728 , y729 , y730 , y731 , y732 , y733 , y734 , y735 , y736 , y737 , y738 , y739 , y740 , y741 , y742 , y743 , y744 , y745 , y746 , y747 , y748 , y749 , y750 , y751 , y752 , y753 , y754 , y755 , y756 , y757 , y758 , y759 , y760 , y761 , y762 , y763 , y764 , y765 , y766 , y767 , y768 , y769 , y770 , y771 , y772 , y773 , y774 , y775 , y776 , y777 , y778 , y779 , y780 , y781 , y782 , y783 , y784 , y785 , y786 , y787 , y788 , y789 , y790 , y791 , y792 , y793 , y794 , y795 , y796 , y797 , y798 , y799 , y800 , y801 , y802 , y803 , y804 , y805 , y806 , y807 , y808 , y809 , y810 , y811 , y812 , y813 , y814 , y815 , y816 , y817 , y818 , y819 , y820 , y821 , y822 , y823 , y824 , y825 , y826 , y827 , y828 , y829 , y830 , y831 , y832 , y833 , y834 , y835 , y836 , y837 , y838 , y839 , y840 , y841 , y842 , y843 , y844 , y845 , y846 , y847 , y848 , y849 , y850 , y851 , y852 , y853 , y854 , y855 , y856 , y857 , y858 , y859 , y860 , y861 , y862 , y863 , y864 , y865 , y866 , y867 , y868 , y869 , y870 , y871 , y872 , y873 , y874 , y875 , y876 , y877 , y878 , y879 , y880 , y881 , y882 , y883 , y884 , y885 , y886 , y887 , y888 , y889 , y890 , y891 , y892 , y893 , y894 , y895 , y896 , y897 , y898 , y899 , y900 , y901 , y902 , y903 , y904 , y905 , y906 , y907 , y908 , y909 , y910 , y911 , y912 , y913 , y914 , y915 , y916 , y917 , y918 , y919 , y920 , y921 , y922 , y923 , y924 , y925 , y926 , y927 , y928 , y929 , y930 , y931 , y932 , y933 , y934 , y935 , y936 , y937 , y938 , y939 , y940 , y941 , y942 , y943 , y944 , y945 , y946 , y947 , y948 , y949 , y950 , y951 , y952 , y953 , y954 , y955 , y956 , y957 , y958 , y959 , y960 , y961 , y962 , y963 , y964 , y965 , y966 , y967 , y968 , y969 , y970 , y971 , y972 , y973 , y974 , y975 , y976 , y977 , y978 , y979 , y980 , y981 , y982 , y983 , y984 , y985 , y986 , y987 , y988 , y989 , y990 , y991 , y992 , y993 , y994 , y995 , y996 , y997 , y998 , y999 , y1000 , y1001 , y1002 , y1003 , y1004 , y1005 , y1006 , y1007 , y1008 , y1009 , y1010 , y1011 , y1012 , y1013 , y1014 , y1015 , y1016 , y1017 , y1018 , y1019 , y1020 , y1021 , y1022 , y1023 , y1024 , y1025 , y1026 , y1027 , y1028 , y1029 , y1030 , y1031 , y1032 , y1033 , y1034 , y1035 , y1036 , y1037 , y1038 , y1039 , y1040 , y1041 , y1042 , y1043 , y1044 , y1045 , y1046 , y1047 , y1048 , y1049 , y1050 , y1051 , y1052 , y1053 , y1054 , y1055 , y1056 , y1057 , y1058 , y1059 , y1060 , y1061 , y1062 , y1063 , y1064 , y1065 , y1066 , y1067 , y1068 , y1069 , y1070 , y1071 , y1072 , y1073 , y1074 , y1075 , y1076 , y1077 , y1078 , y1079 , y1080 , y1081 , y1082 , y1083 , y1084 , y1085 , y1086 , y1087 , y1088 , y1089 , y1090 , y1091 , y1092 , y1093 , y1094 , y1095 , y1096 , y1097 , y1098 , y1099 , y1100 , y1101 , y1102 , y1103 , y1104 , y1105 , y1106 , y1107 , y1108 , y1109 , y1110 , y1111 , y1112 , y1113 , y1114 , y1115 , y1116 , y1117 , y1118 , y1119 , y1120 , y1121 , y1122 , y1123 , y1124 , y1125 , y1126 , y1127 , y1128 , y1129 , y1130 , y1131 , y1132 , y1133 , y1134 , y1135 , y1136 , y1137 , y1138 , y1139 , y1140 , y1141 , y1142 , y1143 , y1144 , y1145 , y1146 , y1147 , y1148 , y1149 , y1150 , y1151 , y1152 , y1153 , y1154 , y1155 , y1156 , y1157 , y1158 , y1159 , y1160 , y1161 , y1162 , y1163 , y1164 , y1165 , y1166 , y1167 , y1168 , y1169 , y1170 , y1171 , y1172 , y1173 , y1174 , y1175 , y1176 , y1177 , y1178 , y1179 , y1180 , y1181 , y1182 , y1183 , y1184 , y1185 , y1186 , y1187 , y1188 , y1189 , y1190 , y1191 , y1192 , y1193 , y1194 , y1195 , y1196 , y1197 , y1198 , y1199 , y1200 , y1201 , y1202 , y1203 , y1204 , y1205 , y1206 , y1207 , y1208 , y1209 , y1210 , y1211 , y1212 , y1213 , y1214 , y1215 , y1216 , y1217 , y1218 , y1219 , y1220 , y1221 , y1222 , y1223 , y1224 , y1225 , y1226 , y1227 , y1228 , y1229 , y1230 , y1231 , y1232 , y1233 , y1234 , y1235 , y1236 , y1237 , y1238 , y1239 , y1240 , y1241 , y1242 , y1243 , y1244 , y1245 , y1246 , y1247 , y1248 , y1249 , y1250 , y1251 , y1252 , y1253 , y1254 , y1255 , y1256 , y1257 , y1258 , y1259 , y1260 , y1261 , y1262 , y1263 , y1264 , y1265 , y1266 , y1267 , y1268 , y1269 , y1270 , y1271 , y1272 , y1273 , y1274 , y1275 , y1276 , y1277 , y1278 , y1279 , y1280 , y1281 , y1282 , y1283 , y1284 , y1285 , y1286 , y1287 , y1288 , y1289 , y1290 , y1291 , y1292 , y1293 , y1294 , y1295 , y1296 , y1297 , y1298 , y1299 , y1300 , y1301 , y1302 , y1303 , y1304 , y1305 , y1306 , y1307 , y1308 , y1309 , y1310 , y1311 , y1312 , y1313 , y1314 , y1315 , y1316 , y1317 , y1318 , y1319 , y1320 , y1321 , y1322 , y1323 , y1324 , y1325 , y1326 , y1327 , y1328 , y1329 , y1330 , y1331 , y1332 , y1333 , y1334 , y1335 , y1336 , y1337 , y1338 , y1339 , y1340 , y1341 , y1342 , y1343 , y1344 , y1345 , y1346 , y1347 , y1348 , y1349 , y1350 , y1351 , y1352 , y1353 , y1354 , y1355 , y1356 , y1357 , y1358 , y1359 , y1360 , y1361 , y1362 , y1363 , y1364 , y1365 , y1366 , y1367 , y1368 , y1369 , y1370 , y1371 , y1372 , y1373 , y1374 , y1375 , y1376 , y1377 , y1378 , y1379 , y1380 , y1381 , y1382 , y1383 , y1384 , y1385 , y1386 , y1387 , y1388 , y1389 , y1390 , y1391 , y1392 , y1393 , y1394 , y1395 , y1396 , y1397 , y1398 , y1399 , y1400 , y1401 , y1402 , y1403 , y1404 , y1405 , y1406 , y1407 , y1408 , y1409 , y1410 , y1411 , y1412 , y1413 , y1414 , y1415 , y1416 , y1417 , y1418 , y1419 , y1420 , y1421 , y1422 , y1423 , y1424 , y1425 , y1426 , y1427 , y1428 , y1429 , y1430 , y1431 , y1432 , y1433 , y1434 , y1435 , y1436 , y1437 , y1438 , y1439 , y1440 , y1441 , y1442 , y1443 , y1444 , y1445 , y1446 , y1447 , y1448 , y1449 , y1450 , y1451 , y1452 , y1453 , y1454 , y1455 , y1456 , y1457 , y1458 , y1459 , y1460 , y1461 , y1462 , y1463 , y1464 , y1465 , y1466 , y1467 , y1468 , y1469 , y1470 , y1471 , y1472 , y1473 , y1474 , y1475 , y1476 , y1477 , y1478 , y1479 , y1480 , y1481 , y1482 , y1483 , y1484 , y1485 , y1486 , y1487 , y1488 , y1489 , y1490 , y1491 , y1492 , y1493 , y1494 , y1495 , y1496 , y1497 , y1498 , y1499 , y1500 , y1501 , y1502 , y1503 , y1504 , y1505 , y1506 , y1507 , y1508 , y1509 , y1510 , y1511 , y1512 , y1513 , y1514 , y1515 , y1516 , y1517 , y1518 , y1519 , y1520 , y1521 , y1522 , y1523 , y1524 , y1525 , y1526 , y1527 , y1528 , y1529 , y1530 , y1531 , y1532 , y1533 , y1534 , y1535 , y1536 , y1537 , y1538 , y1539 , y1540 , y1541 , y1542 , y1543 , y1544 , y1545 , y1546 , y1547 , y1548 , y1549 , y1550 , y1551 , y1552 , y1553 , y1554 , y1555 , y1556 , y1557 , y1558 , y1559 , y1560 , y1561 , y1562 , y1563 , y1564 , y1565 , y1566 , y1567 , y1568 , y1569 , y1570 , y1571 , y1572 , y1573 , y1574 , y1575 , y1576 , y1577 , y1578 , y1579 , y1580 , y1581 , y1582 , y1583 , y1584 , y1585 , y1586 , y1587 , y1588 , y1589 , y1590 , y1591 , y1592 , y1593 , y1594 , y1595 , y1596 , y1597 , y1598 , y1599 , y1600 , y1601 , y1602 , y1603 , y1604 , y1605 , y1606 , y1607 , y1608 , y1609 , y1610 , y1611 , y1612 , y1613 , y1614 , y1615 , y1616 , y1617 , y1618 , y1619 , y1620 , y1621 , y1622 , y1623 , y1624 , y1625 , y1626 , y1627 , y1628 , y1629 , y1630 , y1631 , y1632 , y1633 , y1634 , y1635 , y1636 , y1637 , y1638 , y1639 , y1640 , y1641 , y1642 , y1643 , y1644 , y1645 , y1646 , y1647 , y1648 , y1649 , y1650 , y1651 , y1652 , y1653 , y1654 , y1655 , y1656 , y1657 , y1658 , y1659 , y1660 , y1661 , y1662 , y1663 , y1664 , y1665 , y1666 , y1667 , y1668 , y1669 , y1670 , y1671 , y1672 , y1673 , y1674 , y1675 , y1676 , y1677 , y1678 , y1679 , y1680 , y1681 , y1682 , y1683 , y1684 , y1685 , y1686 , y1687 , y1688 , y1689 , y1690 , y1691 , y1692 , y1693 , y1694 , y1695 , y1696 , y1697 , y1698 , y1699 , y1700 , y1701 , y1702 , y1703 , y1704 , y1705 , y1706 , y1707 , y1708 , y1709 , y1710 , y1711 , y1712 , y1713 , y1714 , y1715 , y1716 , y1717 , y1718 , y1719 , y1720 , y1721 , y1722 , y1723 , y1724 , y1725 , y1726 , y1727 , y1728 , y1729 , y1730 , y1731 , y1732 , y1733 , y1734 , y1735 , y1736 , y1737 , y1738 , y1739 , y1740 , y1741 , y1742 , y1743 , y1744 , y1745 , y1746 , y1747 , y1748 , y1749 , y1750 , y1751 , y1752 , y1753 , y1754 , y1755 , y1756 , y1757 , y1758 , y1759 , y1760 , y1761 , y1762 , y1763 , y1764 , y1765 , y1766 , y1767 , y1768 , y1769 , y1770 , y1771 , y1772 , y1773 , y1774 , y1775 , y1776 , y1777 , y1778 , y1779 , y1780 , y1781 , y1782 , y1783 , y1784 , y1785 , y1786 , y1787 , y1788 , y1789 , y1790 , y1791 , y1792 , y1793 , y1794 , y1795 , y1796 , y1797 , y1798 , y1799 , y1800 , y1801 , y1802 , y1803 , y1804 , y1805 , y1806 , y1807 , y1808 , y1809 , y1810 , y1811 , y1812 , y1813 , y1814 , y1815 , y1816 , y1817 , y1818 , y1819 , y1820 , y1821 , y1822 , y1823 , y1824 , y1825 , y1826 , y1827 , y1828 , y1829 , y1830 , y1831 , y1832 , y1833 , y1834 , y1835 , y1836 , y1837 , y1838 , y1839 , y1840 , y1841 , y1842 , y1843 , y1844 , y1845 , y1846 , y1847 , y1848 , y1849 , y1850 , y1851 , y1852 , y1853 , y1854 , y1855 , y1856 , y1857 , y1858 , y1859 , y1860 , y1861 , y1862 , y1863 , y1864 , y1865 , y1866 , y1867 , y1868 , y1869 , y1870 , y1871 , y1872 , y1873 , y1874 , y1875 , y1876 , y1877 , y1878 , y1879 , y1880 , y1881 , y1882 , y1883 , y1884 , y1885 , y1886 , y1887 , y1888 , y1889 , y1890 , y1891 , y1892 , y1893 , y1894 , y1895 , y1896 , y1897 , y1898 , y1899 , y1900 , y1901 , y1902 , y1903 , y1904 , y1905 , y1906 , y1907 , y1908 , y1909 , y1910 , y1911 , y1912 , y1913 , y1914 , y1915 , y1916 , y1917 , y1918 , y1919 , y1920 , y1921 , y1922 , y1923 , y1924 , y1925 , y1926 , y1927 , y1928 , y1929 , y1930 , y1931 , y1932 , y1933 , y1934 , y1935 , y1936 , y1937 , y1938 , y1939 , y1940 , y1941 , y1942 , y1943 , y1944 , y1945 , y1946 , y1947 , y1948 , y1949 , y1950 , y1951 , y1952 , y1953 , y1954 , y1955 , y1956 , y1957 , y1958 , y1959 , y1960 , y1961 , y1962 , y1963 , y1964 , y1965 , y1966 , y1967 , y1968 , y1969 , y1970 , y1971 , y1972 , y1973 , y1974 , y1975 , y1976 , y1977 , y1978 , y1979 , y1980 , y1981 , y1982 , y1983 , y1984 , y1985 , y1986 , y1987 , y1988 , y1989 , y1990 , y1991 , y1992 , y1993 , y1994 , y1995 , y1996 , y1997 , y1998 , y1999 , y2000 , y2001 , y2002 , y2003 , y2004 , y2005 , y2006 , y2007 , y2008 , y2009 , y2010 , y2011 , y2012 , y2013 , y2014 , y2015 , y2016 , y2017 , y2018 , y2019 , y2020 , y2021 , y2022 , y2023 , y2024 , y2025 , y2026 , y2027 , y2028 , y2029 , y2030 , y2031 , y2032 , y2033 , y2034 , y2035 , y2036 , y2037 , y2038 , y2039 , y2040 , y2041 , y2042 , y2043 , y2044 , y2045 , y2046 , y2047 , y2048 , y2049 , y2050 , y2051 , y2052 , y2053 , y2054 , y2055 , y2056 , y2057 , y2058 , y2059 , y2060 , y2061 , y2062 , y2063 , y2064 , y2065 , y2066 , y2067 , y2068 , y2069 , y2070 , y2071 , y2072 , y2073 , y2074 , y2075 , y2076 , y2077 , y2078 , y2079 , y2080 , y2081 , y2082 , y2083 , y2084 , y2085 , y2086 , y2087 , y2088 , y2089 , y2090 , y2091 , y2092 , y2093 , y2094 , y2095 , y2096 , y2097 , y2098 , y2099 , y2100 , y2101 , y2102 , y2103 , y2104 , y2105 , y2106 , y2107 , y2108 , y2109 , y2110 , y2111 , y2112 , y2113 , y2114 , y2115 , y2116 , y2117 , y2118 , y2119 , y2120 , y2121 , y2122 , y2123 , y2124 , y2125 , y2126 , y2127 , y2128 , y2129 , y2130 , y2131 , y2132 , y2133 , y2134 , y2135 , y2136 , y2137 , y2138 , y2139 , y2140 , y2141 , y2142 , y2143 , y2144 , y2145 , y2146 , y2147 , y2148 , y2149 , y2150 , y2151 , y2152 , y2153 , y2154 , y2155 , y2156 , y2157 , y2158 , y2159 , y2160 , y2161 , y2162 , y2163 , y2164 , y2165 , y2166 , y2167 , y2168 , y2169 , y2170 , y2171 , y2172 , y2173 , y2174 , y2175 , y2176 , y2177 , y2178 , y2179 , y2180 , y2181 , y2182 , y2183 , y2184 , y2185 , y2186 , y2187 , y2188 , y2189 , y2190 , y2191 , y2192 , y2193 , y2194 , y2195 , y2196 , y2197 , y2198 , y2199 , y2200 , y2201 , y2202 , y2203 , y2204 , y2205 , y2206 , y2207 , y2208 , y2209 , y2210 , y2211 , y2212 , y2213 , y2214 , y2215 , y2216 , y2217 , y2218 , y2219 , y2220 , y2221 , y2222 , y2223 , y2224 , y2225 , y2226 , y2227 , y2228 , y2229 , y2230 , y2231 , y2232 , y2233 , y2234 , y2235 , y2236 , y2237 , y2238 , y2239 , y2240 , y2241 , y2242 , y2243 , y2244 , y2245 , y2246 , y2247 , y2248 , y2249 , y2250 , y2251 , y2252 , y2253 , y2254 , y2255 , y2256 , y2257 , y2258 , y2259 , y2260 , y2261 , y2262 , y2263 , y2264 , y2265 , y2266 , y2267 , y2268 , y2269 , y2270 , y2271 , y2272 , y2273 , y2274 , y2275 , y2276 , y2277 , y2278 , y2279 , y2280 , y2281 , y2282 , y2283 , y2284 , y2285 , y2286 , y2287 , y2288 , y2289 , y2290 , y2291 , y2292 , y2293 , y2294 , y2295 , y2296 , y2297 , y2298 , y2299 , y2300 , y2301 , y2302 , y2303 , y2304 , y2305 , y2306 , y2307 , y2308 , y2309 , y2310 , y2311 , y2312 , y2313 , y2314 , y2315 , y2316 , y2317 , y2318 , y2319 , y2320 , y2321 , y2322 , y2323 , y2324 , y2325 , y2326 , y2327 , y2328 , y2329 , y2330 , y2331 , y2332 , y2333 , y2334 , y2335 , y2336 , y2337 , y2338 , y2339 , y2340 , y2341 , y2342 , y2343 , y2344 , y2345 , y2346 , y2347 , y2348 , y2349 , y2350 , y2351 , y2352 , y2353 , y2354 , y2355 , y2356 , y2357 , y2358 , y2359 , y2360 , y2361 , y2362 , y2363 , y2364 , y2365 , y2366 , y2367 , y2368 , y2369 , y2370 , y2371 , y2372 , y2373 , y2374 , y2375 , y2376 , y2377 , y2378 , y2379 , y2380 , y2381 , y2382 , y2383 , y2384 , y2385 , y2386 , y2387 , y2388 , y2389 , y2390 , y2391 , y2392 , y2393 , y2394 , y2395 , y2396 , y2397 , y2398 , y2399 , y2400 , y2401 , y2402 , y2403 , y2404 , y2405 , y2406 , y2407 , y2408 , y2409 , y2410 , y2411 , y2412 , y2413 , y2414 , y2415 , y2416 , y2417 , y2418 , y2419 , y2420 , y2421 , y2422 , y2423 , y2424 , y2425 , y2426 , y2427 , y2428 , y2429 , y2430 , y2431 , y2432 , y2433 , y2434 , y2435 , y2436 , y2437 , y2438 , y2439 , y2440 , y2441 , y2442 , y2443 , y2444 , y2445 , y2446 , y2447 , y2448 , y2449 , y2450 , y2451 , y2452 , y2453 , y2454 , y2455 , y2456 , y2457 , y2458 , y2459 , y2460 , y2461 , y2462 , y2463 , y2464 , y2465 , y2466 , y2467 , y2468 , y2469 , y2470 , y2471 , y2472 , y2473 , y2474 , y2475 , y2476 , y2477 , y2478 , y2479 , y2480 , y2481 , y2482 , y2483 , y2484 , y2485 , y2486 , y2487 , y2488 , y2489 , y2490 , y2491 , y2492 , y2493 , y2494 , y2495 , y2496 , y2497 , y2498 , y2499 , y2500 , y2501 , y2502 , y2503 , y2504 , y2505 , y2506 , y2507 , y2508 , y2509 , y2510 , y2511 , y2512 , y2513 , y2514 , y2515 , y2516 , y2517 , y2518 , y2519 , y2520 , y2521 , y2522 , y2523 , y2524 , y2525 , y2526 , y2527 , y2528 , y2529 , y2530 , y2531 , y2532 , y2533 , y2534 , y2535 , y2536 , y2537 , y2538 , y2539 , y2540 , y2541 , y2542 , y2543 , y2544 , y2545 , y2546 , y2547 , y2548 , y2549 , y2550 , y2551 , y2552 , y2553 , y2554 , y2555 , y2556 , y2557 , y2558 , y2559 , y2560 , y2561 , y2562 , y2563 , y2564 , y2565 , y2566 , y2567 , y2568 , y2569 , y2570 , y2571 , y2572 , y2573 , y2574 , y2575 , y2576 , y2577 , y2578 , y2579 , y2580 , y2581 , y2582 , y2583 , y2584 , y2585 , y2586 , y2587 , y2588 , y2589 , y2590 , y2591 , y2592 , y2593 , y2594 , y2595 , y2596 , y2597 , y2598 , y2599 , y2600 , y2601 , y2602 , y2603 , y2604 , y2605 , y2606 , y2607 , y2608 , y2609 , y2610 , y2611 , y2612 , y2613 , y2614 , y2615 , y2616 , y2617 , y2618 , y2619 , y2620 , y2621 , y2622 , y2623 , y2624 , y2625 , y2626 , y2627 , y2628 , y2629 , y2630 , y2631 , y2632 , y2633 , y2634 , y2635 , y2636 , y2637 , y2638 , y2639 , y2640 , y2641 , y2642 , y2643 , y2644 , y2645 , y2646 , y2647 , y2648 , y2649 , y2650 , y2651 , y2652 , y2653 , y2654 , y2655 , y2656 , y2657 , y2658 , y2659 , y2660 , y2661 , y2662 , y2663 , y2664 , y2665 , y2666 , y2667 , y2668 , y2669 , y2670 , y2671 , y2672 , y2673 , y2674 , y2675 , y2676 , y2677 , y2678 , y2679 , y2680 , y2681 , y2682 , y2683 , y2684 , y2685 , y2686 , y2687 , y2688 , y2689 , y2690 , y2691 , y2692 , y2693 , y2694 , y2695 , y2696 , y2697 , y2698 , y2699 , y2700 , y2701 , y2702 , y2703 , y2704 , y2705 , y2706 , y2707 , y2708 , y2709 , y2710 , y2711 , y2712 , y2713 , y2714 , y2715 , y2716 , y2717 , y2718 , y2719 , y2720 , y2721 , y2722 , y2723 , y2724 , y2725 , y2726 , y2727 , y2728 , y2729 , y2730 , y2731 , y2732 , y2733 , y2734 , y2735 , y2736 , y2737 , y2738 , y2739 , y2740 , y2741 , y2742 , y2743 , y2744 , y2745 , y2746 , y2747 , y2748 , y2749 , y2750 , y2751 , y2752 , y2753 , y2754 , y2755 , y2756 , y2757 , y2758 , y2759 , y2760 , y2761 , y2762 , y2763 , y2764 , y2765 , y2766 , y2767 , y2768 , y2769 , y2770 , y2771 , y2772 , y2773 , y2774 , y2775 , y2776 , y2777 , y2778 , y2779 , y2780 , y2781 , y2782 , y2783 , y2784 , y2785 , y2786 , y2787 , y2788 , y2789 , y2790 , y2791 , y2792 , y2793 , y2794 , y2795 , y2796 , y2797 , y2798 , y2799 , y2800 , y2801 , y2802 , y2803 , y2804 , y2805 , y2806 , y2807 , y2808 , y2809 , y2810 , y2811 , y2812 , y2813 , y2814 , y2815 , y2816 , y2817 , y2818 , y2819 , y2820 , y2821 , y2822 , y2823 , y2824 , y2825 , y2826 , y2827 , y2828 , y2829 , y2830 , y2831 , y2832 , y2833 , y2834 , y2835 , y2836 , y2837 , y2838 , y2839 , y2840 , y2841 , y2842 , y2843 , y2844 , y2845 , y2846 , y2847 , y2848 , y2849 , y2850 , y2851 , y2852 , y2853 , y2854 , y2855 , y2856 , y2857 , y2858 , y2859 , y2860 , y2861 , y2862 , y2863 , y2864 , y2865 , y2866 , y2867 , y2868 , y2869 , y2870 , y2871 , y2872 , y2873 , y2874 , y2875 , y2876 , y2877 , y2878 , y2879 , y2880 , y2881 , y2882 , y2883 , y2884 , y2885 , y2886 , y2887 , y2888 , y2889 , y2890 , y2891 , y2892 , y2893 , y2894 , y2895 , y2896 , y2897 , y2898 , y2899 , y2900 , y2901 , y2902 , y2903 , y2904 , y2905 , y2906 , y2907 , y2908 , y2909 , y2910 , y2911 , y2912 , y2913 , y2914 , y2915 , y2916 , y2917 , y2918 , y2919 , y2920 , y2921 , y2922 , y2923 , y2924 , y2925 , y2926 , y2927 , y2928 , y2929 , y2930 , y2931 , y2932 , y2933 , y2934 , y2935 , y2936 , y2937 , y2938 , y2939 , y2940 , y2941 , y2942 , y2943 , y2944 , y2945 , y2946 , y2947 , y2948 , y2949 , y2950 , y2951 , y2952 , y2953 , y2954 , y2955 , y2956 , y2957 , y2958 , y2959 , y2960 , y2961 , y2962 , y2963 , y2964 , y2965 , y2966 , y2967 , y2968 , y2969 , y2970 , y2971 , y2972 , y2973 , y2974 , y2975 , y2976 , y2977 , y2978 , y2979 , y2980 , y2981 , y2982 , y2983 , y2984 , y2985 , y2986 , y2987 , y2988 , y2989 , y2990 , y2991 , y2992 , y2993 , y2994 , y2995 , y2996 , y2997 , y2998 , y2999 , y3000 , y3001 , y3002 , y3003 , y3004 , y3005 , y3006 , y3007 , y3008 , y3009 , y3010 , y3011 , y3012 , y3013 , y3014 , y3015 , y3016 , y3017 , y3018 , y3019 , y3020 , y3021 , y3022 , y3023 , y3024 , y3025 , y3026 , y3027 , y3028 , y3029 , y3030 , y3031 , y3032 , y3033 , y3034 , y3035 , y3036 , y3037 , y3038 , y3039 , y3040 , y3041 , y3042 , y3043 , y3044 , y3045 , y3046 , y3047 , y3048 , y3049 , y3050 , y3051 , y3052 , y3053 , y3054 , y3055 , y3056 , y3057 , y3058 , y3059 , y3060 , y3061 , y3062 , y3063 , y3064 , y3065 , y3066 , y3067 , y3068 , y3069 , y3070 , y3071 , y3072 , y3073 , y3074 , y3075 , y3076 , y3077 , y3078 , y3079 , y3080 , y3081 , y3082 , y3083 , y3084 , y3085 , y3086 , y3087 , y3088 , y3089 , y3090 , y3091 , y3092 , y3093 , y3094 , y3095 , y3096 , y3097 , y3098 , y3099 , y3100 , y3101 , y3102 , y3103 , y3104 , y3105 , y3106 , y3107 , y3108 , y3109 , y3110 , y3111 , y3112 , y3113 , y3114 , y3115 , y3116 , y3117 , y3118 , y3119 , y3120 , y3121 , y3122 , y3123 , y3124 , y3125 , y3126 , y3127 , y3128 , y3129 , y3130 , y3131 , y3132 , y3133 , y3134 , y3135 , y3136 , y3137 , y3138 , y3139 , y3140 , y3141 , y3142 , y3143 , y3144 , y3145 , y3146 , y3147 , y3148 , y3149 , y3150 , y3151 , y3152 , y3153 , y3154 , y3155 , y3156 , y3157 , y3158 , y3159 , y3160 , y3161 , y3162 , y3163 , y3164 , y3165 , y3166 , y3167 , y3168 , y3169 , y3170 , y3171 , y3172 , y3173 , y3174 , y3175 , y3176 , y3177 , y3178 , y3179 , y3180 , y3181 , y3182 , y3183 , y3184 , y3185 , y3186 , y3187 , y3188 , y3189 , y3190 , y3191 , y3192 , y3193 , y3194 , y3195 , y3196 , y3197 , y3198 , y3199 , y3200 , y3201 , y3202 , y3203 , y3204 , y3205 , y3206 , y3207 , y3208 , y3209 , y3210 , y3211 , y3212 , y3213 , y3214 , y3215 , y3216 , y3217 , y3218 , y3219 , y3220 , y3221 , y3222 , y3223 , y3224 , y3225 , y3226 , y3227 , y3228 , y3229 , y3230 , y3231 , y3232 , y3233 , y3234 , y3235 , y3236 , y3237 , y3238 , y3239 , y3240 , y3241 , y3242 , y3243 , y3244 , y3245 , y3246 , y3247 , y3248 , y3249 , y3250 , y3251 , y3252 , y3253 , y3254 , y3255 , y3256 , y3257 , y3258 , y3259 , y3260 , y3261 , y3262 , y3263 , y3264 , y3265 , y3266 , y3267 , y3268 , y3269 , y3270 , y3271 , y3272 , y3273 , y3274 , y3275 , y3276 , y3277 , y3278 , y3279 , y3280 , y3281 , y3282 , y3283 , y3284 , y3285 , y3286 , y3287 , y3288 , y3289 , y3290 , y3291 , y3292 , y3293 , y3294 , y3295 , y3296 , y3297 , y3298 , y3299 , y3300 , y3301 , y3302 , y3303 , y3304 , y3305 , y3306 , y3307 , y3308 , y3309 , y3310 , y3311 , y3312 , y3313 , y3314 , y3315 , y3316 , y3317 , y3318 , y3319 , y3320 , y3321 , y3322 , y3323 , y3324 , y3325 , y3326 , y3327 , y3328 , y3329 , y3330 , y3331 , y3332 , y3333 , y3334 , y3335 , y3336 , y3337 , y3338 , y3339 , y3340 , y3341 , y3342 , y3343 , y3344 , y3345 , y3346 , y3347 , y3348 , y3349 , y3350 , y3351 , y3352 , y3353 , y3354 , y3355 , y3356 , y3357 , y3358 , y3359 , y3360 , y3361 , y3362 , y3363 , y3364 , y3365 , y3366 , y3367 , y3368 , y3369 , y3370 , y3371 , y3372 , y3373 , y3374 , y3375 , y3376 , y3377 , y3378 , y3379 , y3380 , y3381 , y3382 , y3383 , y3384 , y3385 , y3386 , y3387 , y3388 , y3389 , y3390 , y3391 , y3392 , y3393 , y3394 , y3395 , y3396 , y3397 , y3398 , y3399 , y3400 , y3401 , y3402 , y3403 , y3404 , y3405 , y3406 , y3407 , y3408 , y3409 , y3410 , y3411 , y3412 , y3413 , y3414 , y3415 , y3416 , y3417 , y3418 , y3419 , y3420 , y3421 , y3422 , y3423 , y3424 , y3425 , y3426 , y3427 , y3428 , y3429 , y3430 , y3431 , y3432 , y3433 , y3434 , y3435 , y3436 , y3437 , y3438 , y3439 , y3440 , y3441 , y3442 , y3443 , y3444 , y3445 , y3446 , y3447 , y3448 , y3449 , y3450 , y3451 , y3452 , y3453 , y3454 , y3455 , y3456 , y3457 , y3458 , y3459 , y3460 , y3461 , y3462 , y3463 , y3464 , y3465 , y3466 , y3467 , y3468 , y3469 , y3470 , y3471 , y3472 , y3473 , y3474 , y3475 , y3476 , y3477 , y3478 , y3479 , y3480 , y3481 , y3482 , y3483 , y3484 , y3485 , y3486 , y3487 , y3488 , y3489 , y3490 , y3491 , y3492 , y3493 , y3494 , y3495 , y3496 , y3497 , y3498 , y3499 , y3500 , y3501 , y3502 , y3503 , y3504 , y3505 , y3506 , y3507 , y3508 , y3509 , y3510 , y3511 , y3512 , y3513 , y3514 , y3515 , y3516 , y3517 , y3518 , y3519 , y3520 , y3521 , y3522 , y3523 , y3524 , y3525 , y3526 , y3527 , y3528 , y3529 , y3530 , y3531 , y3532 , y3533 , y3534 , y3535 , y3536 , y3537 , y3538 , y3539 , y3540 , y3541 , y3542 , y3543 , y3544 , y3545 , y3546 , y3547 , y3548 , y3549 , y3550 , y3551 , y3552 , y3553 , y3554 , y3555 , y3556 , y3557 , y3558 , y3559 , y3560 , y3561 , y3562 , y3563 , y3564 , y3565 , y3566 , y3567 , y3568 , y3569 , y3570 , y3571 , y3572 , y3573 , y3574 , y3575 , y3576 , y3577 , y3578 , y3579 , y3580 , y3581 , y3582 , y3583 , y3584 , y3585 , y3586 , y3587 , y3588 , y3589 , y3590 , y3591 , y3592 , y3593 , y3594 , y3595 , y3596 , y3597 , y3598 , y3599 , y3600 , y3601 , y3602 , y3603 , y3604 , y3605 , y3606 , y3607 , y3608 , y3609 , y3610 , y3611 , y3612 , y3613 , y3614 , y3615 , y3616 , y3617 , y3618 , y3619 , y3620 , y3621 , y3622 , y3623 , y3624 , y3625 , y3626 , y3627 , y3628 , y3629 , y3630 , y3631 , y3632 , y3633 , y3634 , y3635 , y3636 , y3637 , y3638 , y3639 , y3640 , y3641 , y3642 , y3643 , y3644 , y3645 , y3646 , y3647 , y3648 , y3649 , y3650 , y3651 , y3652 , y3653 , y3654 , y3655 , y3656 , y3657 , y3658 , y3659 , y3660 , y3661 , y3662 , y3663 , y3664 , y3665 , y3666 , y3667 , y3668 , y3669 , y3670 , y3671 , y3672 , y3673 , y3674 , y3675 , y3676 , y3677 , y3678 , y3679 , y3680 , y3681 , y3682 , y3683 , y3684 , y3685 , y3686 , y3687 , y3688 , y3689 , y3690 , y3691 , y3692 , y3693 , y3694 , y3695 , y3696 , y3697 , y3698 , y3699 , y3700 , y3701 , y3702 , y3703 , y3704 , y3705 , y3706 , y3707 , y3708 , y3709 , y3710 , y3711 , y3712 , y3713 , y3714 , y3715 , y3716 , y3717 , y3718 , y3719 , y3720 , y3721 , y3722 , y3723 , y3724 , y3725 , y3726 , y3727 , y3728 , y3729 , y3730 , y3731 , y3732 , y3733 , y3734 , y3735 , y3736 , y3737 , y3738 , y3739 , y3740 , y3741 , y3742 , y3743 , y3744 , y3745 , y3746 , y3747 , y3748 , y3749 , y3750 , y3751 , y3752 , y3753 , y3754 , y3755 , y3756 , y3757 , y3758 , y3759 , y3760 , y3761 , y3762 , y3763 , y3764 , y3765 , y3766 , y3767 , y3768 , y3769 , y3770 , y3771 , y3772 , y3773 , y3774 , y3775 , y3776 , y3777 , y3778 , y3779 , y3780 , y3781 , y3782 , y3783 , y3784 , y3785 , y3786 , y3787 , y3788 , y3789 , y3790 , y3791 , y3792 , y3793 , y3794 , y3795 , y3796 , y3797 , y3798 , y3799 , y3800 , y3801 , y3802 , y3803 , y3804 , y3805 , y3806 , y3807 , y3808 , y3809 , y3810 , y3811 , y3812 , y3813 , y3814 , y3815 , y3816 , y3817 , y3818 , y3819 , y3820 , y3821 , y3822 , y3823 , y3824 , y3825 , y3826 , y3827 , y3828 , y3829 , y3830 , y3831 , y3832 , y3833 , y3834 , y3835 , y3836 , y3837 , y3838 , y3839 , y3840 , y3841 , y3842 , y3843 , y3844 , y3845 , y3846 , y3847 , y3848 , y3849 , y3850 , y3851 , y3852 , y3853 , y3854 , y3855 , y3856 , y3857 , y3858 , y3859 , y3860 , y3861 , y3862 , y3863 , y3864 , y3865 , y3866 , y3867 , y3868 , y3869 , y3870 , y3871 , y3872 , y3873 , y3874 , y3875 , y3876 , y3877 , y3878 , y3879 , y3880 , y3881 , y3882 , y3883 , y3884 , y3885 , y3886 , y3887 , y3888 , y3889 , y3890 , y3891 , y3892 , y3893 , y3894 , y3895 , y3896 , y3897 , y3898 , y3899 , y3900 , y3901 , y3902 , y3903 , y3904 , y3905 , y3906 , y3907 , y3908 , y3909 , y3910 , y3911 , y3912 , y3913 , y3914 , y3915 , y3916 , y3917 , y3918 , y3919 , y3920 , y3921 , y3922 , y3923 , y3924 , y3925 , y3926 , y3927 , y3928 , y3929 , y3930 , y3931 , y3932 , y3933 , y3934 , y3935 , y3936 , y3937 , y3938 , y3939 , y3940 , y3941 , y3942 , y3943 , y3944 , y3945 , y3946 , y3947 , y3948 , y3949 , y3950 , y3951 , y3952 , y3953 , y3954 , y3955 , y3956 , y3957 , y3958 , y3959 , y3960 , y3961 , y3962 , y3963 , y3964 , y3965 , y3966 , y3967 , y3968 , y3969 , y3970 , y3971 , y3972 , y3973 , y3974 , y3975 , y3976 , y3977 , y3978 , y3979 , y3980 , y3981 , y3982 , y3983 , y3984 , y3985 , y3986 , y3987 , y3988 , y3989 , y3990 , y3991 , y3992 , y3993 , y3994 , y3995 , y3996 , y3997 , y3998 , y3999 , y4000 , y4001 , y4002 , y4003 , y4004 , y4005 , y4006 , y4007 , y4008 , y4009 , y4010 , y4011 , y4012 , y4013 , y4014 , y4015 , y4016 , y4017 , y4018 , y4019 , y4020 , y4021 , y4022 , y4023 , y4024 , y4025 , y4026 , y4027 , y4028 , y4029 , y4030 , y4031 , y4032 , y4033 , y4034 , y4035 , y4036 , y4037 , y4038 , y4039 , y4040 , y4041 , y4042 , y4043 , y4044 , y4045 , y4046 , y4047 , y4048 , y4049 , y4050 , y4051 , y4052 , y4053 , y4054 , y4055 , y4056 , y4057 , y4058 , y4059 , y4060 , y4061 , y4062 , y4063 , y4064 , y4065 , y4066 , y4067 , y4068 , y4069 , y4070 , y4071 , y4072 , y4073 , y4074 , y4075 , y4076 , y4077 , y4078 , y4079 , y4080 , y4081 , y4082 , y4083 , y4084 , y4085 , y4086 , y4087 , y4088 , y4089 , y4090 , y4091 , y4092 , y4093 , y4094 , y4095 , y4096 , y4097 , y4098 , y4099 , y4100 , y4101 , y4102 , y4103 , y4104 , y4105 , y4106 , y4107 , y4108 , y4109 , y4110 , y4111 , y4112 , y4113 , y4114 , y4115 , y4116 , y4117 , y4118 , y4119 , y4120 , y4121 , y4122 , y4123 , y4124 , y4125 , y4126 , y4127 , y4128 , y4129 , y4130 , y4131 , y4132 , y4133 , y4134 , y4135 , y4136 , y4137 , y4138 , y4139 , y4140 , y4141 , y4142 , y4143 , y4144 , y4145 , y4146 , y4147 , y4148 , y4149 , y4150 , y4151 , y4152 , y4153 , y4154 , y4155 , y4156 , y4157 , y4158 , y4159 , y4160 , y4161 , y4162 , y4163 , y4164 , y4165 , y4166 , y4167 , y4168 , y4169 , y4170 , y4171 , y4172 , y4173 , y4174 , y4175 , y4176 , y4177 , y4178 , y4179 , y4180 , y4181 , y4182 , y4183 , y4184 , y4185 , y4186 , y4187 , y4188 , y4189 , y4190 , y4191 , y4192 , y4193 , y4194 , y4195 , y4196 , y4197 , y4198 , y4199 , y4200 , y4201 , y4202 , y4203 , y4204 , y4205 , y4206 , y4207 , y4208 , y4209 , y4210 , y4211 , y4212 , y4213 , y4214 , y4215 , y4216 , y4217 , y4218 , y4219 , y4220 , y4221 , y4222 , y4223 , y4224 , y4225 , y4226 , y4227 , y4228 , y4229 , y4230 , y4231 , y4232 , y4233 , y4234 , y4235 , y4236 , y4237 , y4238 , y4239 , y4240 , y4241 , y4242 , y4243 , y4244 , y4245 , y4246 , y4247 , y4248 , y4249 , y4250 , y4251 , y4252 , y4253 , y4254 , y4255 , y4256 , y4257 , y4258 , y4259 , y4260 , y4261 , y4262 , y4263 , y4264 , y4265 , y4266 , y4267 , y4268 , y4269 , y4270 , y4271 , y4272 , y4273 , y4274 , y4275 , y4276 , y4277 , y4278 , y4279 , y4280 , y4281 , y4282 , y4283 , y4284 , y4285 , y4286 , y4287 , y4288 , y4289 , y4290 , y4291 , y4292 , y4293 , y4294 , y4295 , y4296 , y4297 , y4298 , y4299 , y4300 , y4301 , y4302 , y4303 , y4304 , y4305 , y4306 , y4307 , y4308 , y4309 , y4310 , y4311 , y4312 , y4313 , y4314 , y4315 , y4316 , y4317 , y4318 , y4319 , y4320 , y4321 , y4322 , y4323 , y4324 , y4325 , y4326 , y4327 , y4328 , y4329 , y4330 , y4331 , y4332 , y4333 , y4334 , y4335 , y4336 , y4337 , y4338 , y4339 , y4340 , y4341 , y4342 , y4343 , y4344 , y4345 , y4346 , y4347 , y4348 , y4349 , y4350 , y4351 , y4352 , y4353 , y4354 , y4355 , y4356 , y4357 , y4358 , y4359 , y4360 , y4361 , y4362 , y4363 , y4364 , y4365 , y4366 , y4367 , y4368 , y4369 , y4370 , y4371 , y4372 , y4373 , y4374 , y4375 , y4376 , y4377 , y4378 , y4379 , y4380 , y4381 , y4382 , y4383 , y4384 , y4385 , y4386 , y4387 , y4388 , y4389 , y4390 , y4391 , y4392 , y4393 , y4394 , y4395 , y4396 , y4397 , y4398 , y4399 , y4400 , y4401 , y4402 , y4403 , y4404 , y4405 , y4406 , y4407 , y4408 , y4409 , y4410 , y4411 , y4412 , y4413 , y4414 , y4415 , y4416 , y4417 , y4418 , y4419 , y4420 , y4421 , y4422 , y4423 , y4424 , y4425 , y4426 , y4427 , y4428 , y4429 , y4430 , y4431 , y4432 , y4433 , y4434 , y4435 , y4436 , y4437 , y4438 , y4439 , y4440 , y4441 , y4442 , y4443 , y4444 , y4445 , y4446 , y4447 , y4448 , y4449 , y4450 , y4451 , y4452 , y4453 , y4454 , y4455 , y4456 , y4457 , y4458 , y4459 , y4460 , y4461 , y4462 , y4463 , y4464 , y4465 , y4466 , y4467 , y4468 , y4469 , y4470 , y4471 , y4472 , y4473 , y4474 , y4475 , y4476 , y4477 , y4478 , y4479 , y4480 , y4481 , y4482 , y4483 , y4484 , y4485 , y4486 , y4487 , y4488 , y4489 , y4490 , y4491 , y4492 , y4493 , y4494 , y4495 , y4496 , y4497 , y4498 , y4499 , y4500 , y4501 , y4502 , y4503 , y4504 , y4505 , y4506 , y4507 , y4508 , y4509 , y4510 , y4511 , y4512 , y4513 , y4514 , y4515 , y4516 , y4517 , y4518 , y4519 , y4520 , y4521 , y4522 , y4523 , y4524 , y4525 , y4526 , y4527 , y4528 , y4529 , y4530 , y4531 , y4532 , y4533 , y4534 , y4535 , y4536 , y4537 , y4538 , y4539 , y4540 , y4541 , y4542 , y4543 , y4544 , y4545 , y4546 , y4547 , y4548 , y4549 , y4550 , y4551 , y4552 , y4553 , y4554 , y4555 , y4556 , y4557 , y4558 , y4559 , y4560 , y4561 , y4562 , y4563 , y4564 , y4565 , y4566 , y4567 , y4568 , y4569 , y4570 , y4571 , y4572 , y4573 , y4574 , y4575 , y4576 , y4577 , y4578 , y4579 , y4580 , y4581 , y4582 , y4583 , y4584 , y4585 , y4586 , y4587 , y4588 , y4589 , y4590 , y4591 , y4592 , y4593 , y4594 , y4595 , y4596 , y4597 , y4598 , y4599 , y4600 , y4601 , y4602 , y4603 , y4604 , y4605 , y4606 , y4607 , y4608 , y4609 , y4610 , y4611 , y4612 , y4613 , y4614 , y4615 , y4616 , y4617 , y4618 , y4619 , y4620 , y4621 , y4622 , y4623 , y4624 , y4625 , y4626 , y4627 , y4628 , y4629 , y4630 , y4631 , y4632 , y4633 , y4634 , y4635 , y4636 , y4637 , y4638 , y4639 , y4640 , y4641 , y4642 , y4643 , y4644 , y4645 , y4646 , y4647 , y4648 , y4649 , y4650 , y4651 , y4652 , y4653 , y4654 , y4655 , y4656 , y4657 , y4658 , y4659 , y4660 , y4661 , y4662 , y4663 , y4664 , y4665 , y4666 , y4667 , y4668 , y4669 , y4670 , y4671 , y4672 , y4673 , y4674 , y4675 , y4676 , y4677 , y4678 , y4679 , y4680 , y4681 , y4682 , y4683 , y4684 , y4685 , y4686 , y4687 , y4688 , y4689 , y4690 , y4691 , y4692 , y4693 , y4694 , y4695 , y4696 , y4697 , y4698 , y4699 , y4700 , y4701 , y4702 , y4703 , y4704 , y4705 , y4706 , y4707 , y4708 , y4709 , y4710 , y4711 , y4712 , y4713 , y4714 , y4715 , y4716 , y4717 , y4718 , y4719 , y4720 , y4721 , y4722 , y4723 , y4724 , y4725 , y4726 , y4727 , y4728 , y4729 , y4730 , y4731 , y4732 , y4733 , y4734 , y4735 , y4736 , y4737 , y4738 , y4739 , y4740 , y4741 , y4742 , y4743 , y4744 , y4745 , y4746 , y4747 , y4748 , y4749 , y4750 , y4751 , y4752 , y4753 , y4754 , y4755 , y4756 , y4757 , y4758 , y4759 , y4760 , y4761 , y4762 , y4763 , y4764 , y4765 , y4766 , y4767 , y4768 , y4769 , y4770 , y4771 , y4772 , y4773 , y4774 , y4775 , y4776 , y4777 , y4778 , y4779 , y4780 , y4781 , y4782 , y4783 , y4784 , y4785 , y4786 , y4787 , y4788 , y4789 , y4790 , y4791 , y4792 , y4793 , y4794 , y4795 , y4796 , y4797 , y4798 , y4799 , y4800 , y4801 , y4802 , y4803 , y4804 , y4805 , y4806 , y4807 , y4808 , y4809 , y4810 , y4811 , y4812 , y4813 , y4814 , y4815 , y4816 , y4817 , y4818 , y4819 , y4820 , y4821 , y4822 , y4823 , y4824 , y4825 , y4826 , y4827 , y4828 , y4829 , y4830 , y4831 , y4832 , y4833 , y4834 , y4835 , y4836 , y4837 , y4838 , y4839 , y4840 , y4841 , y4842 , y4843 , y4844 , y4845 , y4846 , y4847 , y4848 , y4849 , y4850 , y4851 , y4852 , y4853 , y4854 , y4855 , y4856 , y4857 , y4858 , y4859 , y4860 , y4861 , y4862 , y4863 , y4864 , y4865 , y4866 , y4867 , y4868 , y4869 , y4870 , y4871 , y4872 , y4873 , y4874 , y4875 , y4876 , y4877 , y4878 , y4879 , y4880 , y4881 , y4882 , y4883 , y4884 , y4885 , y4886 , y4887 , y4888 , y4889 , y4890 , y4891 , y4892 , y4893 , y4894 , y4895 , y4896 , y4897 , y4898 , y4899 , y4900 , y4901 , y4902 , y4903 , y4904 , y4905 , y4906 , y4907 , y4908 , y4909 , y4910 , y4911 , y4912 , y4913 , y4914 , y4915 , y4916 , y4917 , y4918 , y4919 , y4920 , y4921 , y4922 , y4923 , y4924 , y4925 , y4926 , y4927 , y4928 , y4929 , y4930 , y4931 , y4932 , y4933 , y4934 , y4935 , y4936 , y4937 , y4938 , y4939 , y4940 , y4941 , y4942 , y4943 , y4944 , y4945 , y4946 , y4947 , y4948 , y4949 , y4950 , y4951 , y4952 , y4953 , y4954 , y4955 , y4956 , y4957 , y4958 , y4959 , y4960 , y4961 , y4962 , y4963 , y4964 , y4965 , y4966 , y4967 , y4968 , y4969 , y4970 , y4971 , y4972 , y4973 , y4974 , y4975 , y4976 , y4977 , y4978 , y4979 , y4980 , y4981 , y4982 , y4983 , y4984 , y4985 , y4986 , y4987 , y4988 , y4989 , y4990 , y4991 , y4992 , y4993 , y4994 , y4995 , y4996 , y4997 , y4998 , y4999 , y5000 , y5001 , y5002 , y5003 , y5004 , y5005 , y5006 , y5007 , y5008 , y5009 , y5010 , y5011 , y5012 , y5013 , y5014 , y5015 , y5016 , y5017 , y5018 , y5019 , y5020 , y5021 , y5022 , y5023 , y5024 , y5025 , y5026 , y5027 , y5028 , y5029 , y5030 , y5031 , y5032 , y5033 , y5034 , y5035 , y5036 , y5037 , y5038 , y5039 , y5040 , y5041 , y5042 , y5043 , y5044 , y5045 , y5046 , y5047 , y5048 , y5049 , y5050 , y5051 , y5052 , y5053 , y5054 , y5055 , y5056 , y5057 , y5058 , y5059 , y5060 , y5061 , y5062 , y5063 , y5064 , y5065 , y5066 , y5067 , y5068 , y5069 , y5070 , y5071 , y5072 , y5073 , y5074 , y5075 , y5076 , y5077 , y5078 , y5079 , y5080 , y5081 , y5082 , y5083 , y5084 , y5085 , y5086 , y5087 , y5088 , y5089 , y5090 , y5091 , y5092 , y5093 , y5094 , y5095 , y5096 , y5097 , y5098 , y5099 , y5100 , y5101 , y5102 , y5103 , y5104 , y5105 , y5106 , y5107 , y5108 , y5109 , y5110 , y5111 , y5112 , y5113 , y5114 , y5115 , y5116 , y5117 , y5118 , y5119 , y5120 , y5121 , y5122 , y5123 , y5124 , y5125 , y5126 , y5127 , y5128 , y5129 , y5130 , y5131 , y5132 , y5133 , y5134 , y5135 , y5136 , y5137 , y5138 , y5139 , y5140 , y5141 , y5142 , y5143 , y5144 , y5145 , y5146 , y5147 , y5148 , y5149 , y5150 , y5151 , y5152 , y5153 , y5154 , y5155 , y5156 , y5157 , y5158 , y5159 , y5160 , y5161 , y5162 , y5163 , y5164 , y5165 , y5166 , y5167 , y5168 , y5169 , y5170 , y5171 , y5172 , y5173 , y5174 , y5175 , y5176 , y5177 , y5178 , y5179 , y5180 , y5181 , y5182 , y5183 , y5184 , y5185 , y5186 , y5187 , y5188 , y5189 , y5190 , y5191 , y5192 , y5193 , y5194 , y5195 , y5196 , y5197 , y5198 , y5199 , y5200 , y5201 , y5202 , y5203 , y5204 , y5205 , y5206 , y5207 , y5208 , y5209 , y5210 , y5211 , y5212 , y5213 , y5214 , y5215 , y5216 , y5217 , y5218 , y5219 , y5220 , y5221 , y5222 , y5223 , y5224 , y5225 , y5226 , y5227 , y5228 , y5229 , y5230 , y5231 , y5232 , y5233 , y5234 , y5235 , y5236 , y5237 , y5238 , y5239 , y5240 , y5241 , y5242 , y5243 , y5244 , y5245 , y5246 , y5247 , y5248 , y5249 , y5250 , y5251 , y5252 , y5253 , y5254 , y5255 , y5256 , y5257 , y5258 , y5259 , y5260 , y5261 , y5262 , y5263 , y5264 , y5265 , y5266 , y5267 , y5268 , y5269 , y5270 , y5271 , y5272 , y5273 , y5274 , y5275 , y5276 , y5277 , y5278 , y5279 , y5280 , y5281 , y5282 , y5283 , y5284 , y5285 , y5286 , y5287 , y5288 , y5289 , y5290 , y5291 , y5292 , y5293 , y5294 , y5295 , y5296 , y5297 , y5298 , y5299 , y5300 , y5301 , y5302 , y5303 , y5304 , y5305 , y5306 , y5307 , y5308 , y5309 , y5310 , y5311 , y5312 , y5313 , y5314 , y5315 , y5316 , y5317 , y5318 , y5319 , y5320 , y5321 , y5322 , y5323 , y5324 , y5325 , y5326 , y5327 , y5328 , y5329 , y5330 , y5331 , y5332 , y5333 , y5334 , y5335 , y5336 , y5337 , y5338 , y5339 , y5340 , y5341 , y5342 , y5343 , y5344 , y5345 , y5346 , y5347 , y5348 , y5349 , y5350 , y5351 , y5352 , y5353 , y5354 , y5355 , y5356 , y5357 , y5358 , y5359 , y5360 , y5361 , y5362 , y5363 , y5364 , y5365 , y5366 , y5367 , y5368 , y5369 , y5370 , y5371 , y5372 , y5373 , y5374 , y5375 , y5376 , y5377 , y5378 , y5379 , y5380 , y5381 , y5382 , y5383 , y5384 , y5385 , y5386 , y5387 , y5388 , y5389 , y5390 , y5391 , y5392 , y5393 , y5394 , y5395 , y5396 , y5397 , y5398 , y5399 , y5400 , y5401 , y5402 , y5403 , y5404 , y5405 , y5406 , y5407 , y5408 , y5409 , y5410 , y5411 , y5412 , y5413 , y5414 , y5415 , y5416 , y5417 , y5418 , y5419 , y5420 , y5421 , y5422 , y5423 , y5424 , y5425 , y5426 , y5427 , y5428 , y5429 , y5430 , y5431 , y5432 , y5433 , y5434 , y5435 , y5436 , y5437 , y5438 , y5439 , y5440 , y5441 , y5442 , y5443 , y5444 , y5445 , y5446 , y5447 , y5448 , y5449 , y5450 , y5451 , y5452 , y5453 , y5454 , y5455 , y5456 , y5457 , y5458 , y5459 , y5460 , y5461 , y5462 , y5463 , y5464 , y5465 , y5466 , y5467 , y5468 , y5469 , y5470 , y5471 , y5472 , y5473 , y5474 , y5475 , y5476 , y5477 , y5478 , y5479 , y5480 , y5481 , y5482 , y5483 , y5484 , y5485 , y5486 , y5487 , y5488 , y5489 , y5490 , y5491 , y5492 , y5493 , y5494 , y5495 , y5496 , y5497 , y5498 , y5499 , y5500 , y5501 , y5502 , y5503 , y5504 , y5505 , y5506 , y5507 , y5508 , y5509 , y5510 , y5511 , y5512 , y5513 , y5514 , y5515 , y5516 , y5517 , y5518 , y5519 , y5520 , y5521 , y5522 , y5523 , y5524 , y5525 , y5526 , y5527 , y5528 , y5529 , y5530 , y5531 , y5532 , y5533 , y5534 , y5535 , y5536 , y5537 , y5538 , y5539 , y5540 , y5541 , y5542 , y5543 , y5544 , y5545 , y5546 , y5547 , y5548 , y5549 , y5550 , y5551 , y5552 , y5553 , y5554 , y5555 , y5556 , y5557 , y5558 , y5559 , y5560 , y5561 , y5562 , y5563 , y5564 , y5565 , y5566 , y5567 , y5568 , y5569 , y5570 , y5571 , y5572 , y5573 , y5574 , y5575 , y5576 , y5577 , y5578 , y5579 , y5580 , y5581 , y5582 , y5583 , y5584 , y5585 , y5586 , y5587 , y5588 , y5589 , y5590 , y5591 , y5592 , y5593 , y5594 , y5595 , y5596 , y5597 , y5598 , y5599 , y5600 , y5601 , y5602 , y5603 , y5604 , y5605 , y5606 , y5607 , y5608 , y5609 , y5610 , y5611 , y5612 , y5613 , y5614 , y5615 , y5616 , y5617 , y5618 , y5619 , y5620 , y5621 , y5622 , y5623 , y5624 , y5625 , y5626 , y5627 , y5628 , y5629 , y5630 , y5631 , y5632 , y5633 , y5634 , y5635 , y5636 , y5637 , y5638 , y5639 , y5640 , y5641 , y5642 , y5643 , y5644 , y5645 , y5646 , y5647 , y5648 , y5649 , y5650 , y5651 , y5652 , y5653 , y5654 , y5655 , y5656 , y5657 , y5658 , y5659 , y5660 , y5661 , y5662 , y5663 , y5664 , y5665 , y5666 , y5667 , y5668 , y5669 , y5670 , y5671 , y5672 , y5673 , y5674 , y5675 , y5676 , y5677 , y5678 , y5679 , y5680 , y5681 , y5682 , y5683 , y5684 , y5685 , y5686 , y5687 , y5688 , y5689 , y5690 , y5691 , y5692 , y5693 , y5694 , y5695 , y5696 , y5697 , y5698 , y5699 , y5700 , y5701 , y5702 , y5703 , y5704 , y5705 , y5706 , y5707 , y5708 , y5709 , y5710 , y5711 , y5712 , y5713 , y5714 , y5715 , y5716 , y5717 , y5718 , y5719 , y5720 , y5721 , y5722 , y5723 , y5724 , y5725 , y5726 , y5727 , y5728 , y5729 , y5730 , y5731 , y5732 , y5733 , y5734 , y5735 , y5736 , y5737 , y5738 , y5739 , y5740 , y5741 , y5742 , y5743 , y5744 , y5745 , y5746 , y5747 , y5748 , y5749 , y5750 , y5751 , y5752 , y5753 , y5754 , y5755 , y5756 , y5757 , y5758 , y5759 , y5760 , y5761 , y5762 , y5763 , y5764 , y5765 , y5766 , y5767 , y5768 , y5769 , y5770 , y5771 , y5772 , y5773 , y5774 , y5775 , y5776 , y5777 , y5778 , y5779 , y5780 , y5781 , y5782 , y5783 , y5784 , y5785 , y5786 , y5787 , y5788 , y5789 , y5790 , y5791 , y5792 , y5793 , y5794 , y5795 , y5796 , y5797 , y5798 , y5799 , y5800 , y5801 , y5802 , y5803 , y5804 , y5805 , y5806 , y5807 , y5808 , y5809 , y5810 , y5811 , y5812 , y5813 , y5814 , y5815 , y5816 , y5817 , y5818 , y5819 , y5820 , y5821 , y5822 , y5823 , y5824 , y5825 , y5826 , y5827 , y5828 , y5829 , y5830 , y5831 , y5832 , y5833 , y5834 , y5835 , y5836 , y5837 , y5838 , y5839 , y5840 , y5841 , y5842 , y5843 , y5844 , y5845 , y5846 , y5847 , y5848 , y5849 , y5850 , y5851 , y5852 , y5853 , y5854 , y5855 , y5856 , y5857 , y5858 , y5859 , y5860 , y5861 , y5862 , y5863 , y5864 , y5865 , y5866 , y5867 , y5868 , y5869 , y5870 , y5871 , y5872 , y5873 , y5874 , y5875 , y5876 , y5877 , y5878 , y5879 , y5880 , y5881 , y5882 , y5883 , y5884 , y5885 , y5886 , y5887 , y5888 , y5889 , y5890 , y5891 , y5892 , y5893 , y5894 , y5895 , y5896 , y5897 , y5898 , y5899 , y5900 , y5901 , y5902 , y5903 , y5904 , y5905 , y5906 , y5907 , y5908 , y5909 , y5910 , y5911 , y5912 , y5913 , y5914 , y5915 , y5916 , y5917 , y5918 , y5919 , y5920 , y5921 , y5922 , y5923 , y5924 , y5925 , y5926 , y5927 , y5928 , y5929 , y5930 , y5931 , y5932 , y5933 , y5934 , y5935 , y5936 , y5937 , y5938 , y5939 , y5940 , y5941 , y5942 , y5943 , y5944 , y5945 , y5946 , y5947 , y5948 , y5949 , y5950 , y5951 , y5952 , y5953 , y5954 , y5955 , y5956 , y5957 , y5958 , y5959 , y5960 , y5961 , y5962 , y5963 , y5964 , y5965 , y5966 , y5967 , y5968 , y5969 , y5970 , y5971 , y5972 , y5973 , y5974 , y5975 , y5976 , y5977 , y5978 , y5979 , y5980 , y5981 , y5982 , y5983 , y5984 , y5985 , y5986 , y5987 , y5988 , y5989 , y5990 , y5991 , y5992 , y5993 , y5994 , y5995 , y5996 , y5997 , y5998 , y5999 , y6000 , y6001 , y6002 , y6003 , y6004 , y6005 , y6006 , y6007 , y6008 , y6009 , y6010 , y6011 , y6012 , y6013 , y6014 , y6015 , y6016 , y6017 , y6018 , y6019 , y6020 , y6021 , y6022 , y6023 , y6024 , y6025 , y6026 , y6027 , y6028 , y6029 , y6030 , y6031 , y6032 , y6033 , y6034 , y6035 , y6036 , y6037 , y6038 , y6039 , y6040 , y6041 , y6042 , y6043 , y6044 , y6045 , y6046 , y6047 , y6048 , y6049 , y6050 , y6051 , y6052 , y6053 , y6054 , y6055 , y6056 , y6057 , y6058 , y6059 , y6060 , y6061 , y6062 , y6063 , y6064 , y6065 , y6066 , y6067 , y6068 , y6069 , y6070 , y6071 , y6072 , y6073 , y6074 , y6075 , y6076 , y6077 , y6078 , y6079 , y6080 , y6081 , y6082 , y6083 , y6084 , y6085 , y6086 , y6087 , y6088 , y6089 , y6090 , y6091 , y6092 , y6093 , y6094 , y6095 , y6096 , y6097 , y6098 , y6099 , y6100 , y6101 , y6102 , y6103 , y6104 , y6105 , y6106 , y6107 , y6108 , y6109 , y6110 , y6111 , y6112 , y6113 , y6114 , y6115 , y6116 , y6117 , y6118 , y6119 , y6120 , y6121 , y6122 , y6123 , y6124 , y6125 , y6126 , y6127 , y6128 , y6129 , y6130 , y6131 , y6132 , y6133 , y6134 , y6135 , y6136 , y6137 , y6138 , y6139 , y6140 , y6141 , y6142 , y6143 , y6144 , y6145 , y6146 , y6147 , y6148 , y6149 , y6150 , y6151 , y6152 , y6153 , y6154 , y6155 , y6156 , y6157 , y6158 , y6159 , y6160 , y6161 , y6162 , y6163 , y6164 , y6165 , y6166 , y6167 , y6168 , y6169 , y6170 , y6171 , y6172 , y6173 , y6174 , y6175 , y6176 , y6177 , y6178 , y6179 , y6180 , y6181 , y6182 , y6183 , y6184 , y6185 , y6186 , y6187 , y6188 , y6189 , y6190 , y6191 , y6192 , y6193 , y6194 , y6195 , y6196 , y6197 , y6198 , y6199 , y6200 , y6201 , y6202 , y6203 , y6204 , y6205 , y6206 , y6207 , y6208 , y6209 , y6210 , y6211 , y6212 , y6213 , y6214 , y6215 , y6216 , y6217 , y6218 , y6219 , y6220 , y6221 , y6222 , y6223 , y6224 , y6225 , y6226 , y6227 , y6228 , y6229 , y6230 , y6231 , y6232 , y6233 , y6234 , y6235 , y6236 , y6237 , y6238 , y6239 , y6240 , y6241 , y6242 , y6243 , y6244 , y6245 , y6246 , y6247 , y6248 , y6249 , y6250 , y6251 , y6252 , y6253 , y6254 , y6255 , y6256 , y6257 , y6258 , y6259 , y6260 , y6261 , y6262 , y6263 , y6264 , y6265 , y6266 , y6267 , y6268 , y6269 , y6270 , y6271 , y6272 , y6273 , y6274 , y6275 , y6276 , y6277 , y6278 , y6279 , y6280 , y6281 , y6282 , y6283 , y6284 , y6285 , y6286 , y6287 , y6288 , y6289 , y6290 , y6291 , y6292 , y6293 , y6294 , y6295 , y6296 , y6297 , y6298 , y6299 , y6300 , y6301 , y6302 , y6303 , y6304 , y6305 , y6306 , y6307 , y6308 , y6309 , y6310 , y6311 , y6312 , y6313 , y6314 , y6315 , y6316 , y6317 , y6318 , y6319 , y6320 , y6321 , y6322 , y6323 , y6324 , y6325 , y6326 , y6327 , y6328 , y6329 , y6330 , y6331 , y6332 , y6333 , y6334 , y6335 , y6336 , y6337 , y6338 , y6339 , y6340 , y6341 , y6342 , y6343 , y6344 , y6345 , y6346 , y6347 , y6348 , y6349 , y6350 , y6351 , y6352 , y6353 , y6354 , y6355 , y6356 , y6357 , y6358 , y6359 , y6360 , y6361 , y6362 , y6363 , y6364 , y6365 , y6366 , y6367 , y6368 , y6369 , y6370 , y6371 , y6372 , y6373 , y6374 , y6375 , y6376 , y6377 , y6378 , y6379 , y6380 , y6381 , y6382 , y6383 , y6384 , y6385 , y6386 , y6387 , y6388 , y6389 , y6390 , y6391 , y6392 , y6393 , y6394 , y6395 , y6396 , y6397 , y6398 , y6399 , y6400 , y6401 , y6402 , y6403 , y6404 , y6405 , y6406 , y6407 , y6408 , y6409 , y6410 , y6411 , y6412 , y6413 , y6414 , y6415 , y6416 , y6417 , y6418 , y6419 , y6420 , y6421 , y6422 , y6423 , y6424 , y6425 , y6426 , y6427 , y6428 , y6429 , y6430 , y6431 , y6432 , y6433 , y6434 , y6435 , y6436 , y6437 , y6438 , y6439 , y6440 , y6441 , y6442 , y6443 , y6444 , y6445 , y6446 , y6447 , y6448 , y6449 , y6450 , y6451 , y6452 , y6453 , y6454 , y6455 , y6456 , y6457 , y6458 , y6459 , y6460 , y6461 , y6462 , y6463 , y6464 , y6465 , y6466 , y6467 , y6468 , y6469 , y6470 , y6471 , y6472 , y6473 , y6474 , y6475 , y6476 , y6477 , y6478 , y6479 , y6480 , y6481 , y6482 , y6483 , y6484 , y6485 , y6486 , y6487 , y6488 , y6489 , y6490 , y6491 , y6492 , y6493 , y6494 , y6495 , y6496 , y6497 , y6498 , y6499 , y6500 , y6501 , y6502 , y6503 , y6504 , y6505 , y6506 , y6507 , y6508 , y6509 , y6510 , y6511 , y6512 , y6513 , y6514 , y6515 , y6516 , y6517 , y6518 , y6519 , y6520 , y6521 , y6522 , y6523 , y6524 , y6525 , y6526 , y6527 , y6528 , y6529 , y6530 , y6531 , y6532 , y6533 , y6534 , y6535 , y6536 , y6537 , y6538 , y6539 , y6540 , y6541 , y6542 , y6543 , y6544 , y6545 , y6546 , y6547 , y6548 , y6549 , y6550 , y6551 , y6552 , y6553 , y6554 , y6555 , y6556 , y6557 , y6558 , y6559 , y6560 , y6561 , y6562 , y6563 , y6564 , y6565 , y6566 , y6567 , y6568 , y6569 , y6570 , y6571 , y6572 , y6573 , y6574 , y6575 , y6576 , y6577 , y6578 , y6579 , y6580 , y6581 , y6582 , y6583 , y6584 , y6585 , y6586 , y6587 , y6588 , y6589 , y6590 , y6591 , y6592 , y6593 , y6594 , y6595 , y6596 , y6597 , y6598 , y6599 , y6600 , y6601 , y6602 , y6603 , y6604 , y6605 , y6606 , y6607 , y6608 , y6609 , y6610 , y6611 , y6612 , y6613 , y6614 , y6615 , y6616 , y6617 , y6618 , y6619 , y6620 , y6621 , y6622 , y6623 , y6624 , y6625 , y6626 , y6627 , y6628 , y6629 , y6630 , y6631 , y6632 , y6633 , y6634 , y6635 , y6636 , y6637 , y6638 , y6639 , y6640 , y6641 , y6642 , y6643 , y6644 , y6645 , y6646 , y6647 , y6648 , y6649 , y6650 , y6651 , y6652 , y6653 , y6654 , y6655 , y6656 , y6657 , y6658 , y6659 , y6660 , y6661 , y6662 , y6663 , y6664 , y6665 , y6666 , y6667 , y6668 , y6669 , y6670 , y6671 , y6672 , y6673 , y6674 , y6675 , y6676 , y6677 , y6678 , y6679 , y6680 , y6681 , y6682 , y6683 , y6684 , y6685 , y6686 , y6687 , y6688 , y6689 , y6690 , y6691 , y6692 , y6693 , y6694 , y6695 , y6696 , y6697 , y6698 , y6699 , y6700 , y6701 , y6702 , y6703 , y6704 , y6705 , y6706 , y6707 , y6708 , y6709 , y6710 , y6711 , y6712 , y6713 , y6714 , y6715 , y6716 , y6717 , y6718 , y6719 , y6720 , y6721 , y6722 , y6723 , y6724 , y6725 , y6726 , y6727 , y6728 , y6729 , y6730 , y6731 , y6732 , y6733 , y6734 , y6735 , y6736 , y6737 , y6738 , y6739 , y6740 , y6741 , y6742 , y6743 , y6744 , y6745 , y6746 , y6747 , y6748 , y6749 , y6750 , y6751 , y6752 , y6753 , y6754 , y6755 , y6756 , y6757 , y6758 , y6759 , y6760 , y6761 , y6762 , y6763 , y6764 , y6765 , y6766 , y6767 , y6768 , y6769 , y6770 , y6771 , y6772 , y6773 , y6774 , y6775 , y6776 , y6777 , y6778 , y6779 , y6780 , y6781 , y6782 , y6783 , y6784 , y6785 , y6786 , y6787 , y6788 , y6789 , y6790 , y6791 , y6792 , y6793 , y6794 , y6795 , y6796 , y6797 , y6798 , y6799 , y6800 , y6801 , y6802 , y6803 , y6804 , y6805 , y6806 , y6807 , y6808 , y6809 , y6810 , y6811 , y6812 , y6813 , y6814 , y6815 , y6816 , y6817 , y6818 , y6819 , y6820 , y6821 , y6822 , y6823 , y6824 , y6825 , y6826 , y6827 , y6828 , y6829 , y6830 , y6831 , y6832 , y6833 , y6834 , y6835 , y6836 , y6837 , y6838 , y6839 , y6840 , y6841 , y6842 , y6843 , y6844 , y6845 , y6846 , y6847 , y6848 , y6849 , y6850 , y6851 , y6852 , y6853 , y6854 , y6855 , y6856 , y6857 , y6858 , y6859 , y6860 , y6861 , y6862 , y6863 , y6864 , y6865 , y6866 , y6867 , y6868 , y6869 , y6870 , y6871 , y6872 , y6873 , y6874 , y6875 , y6876 , y6877 , y6878 , y6879 , y6880 , y6881 , y6882 , y6883 , y6884 , y6885 , y6886 , y6887 , y6888 , y6889 , y6890 , y6891 , y6892 , y6893 , y6894 , y6895 , y6896 , y6897 , y6898 , y6899 , y6900 , y6901 , y6902 , y6903 , y6904 , y6905 , y6906 , y6907 , y6908 , y6909 , y6910 , y6911 , y6912 , y6913 , y6914 , y6915 , y6916 , y6917 , y6918 , y6919 , y6920 , y6921 , y6922 , y6923 , y6924 , y6925 , y6926 , y6927 , y6928 , y6929 , y6930 , y6931 , y6932 , y6933 , y6934 , y6935 , y6936 , y6937 , y6938 , y6939 , y6940 , y6941 , y6942 , y6943 , y6944 , y6945 , y6946 , y6947 , y6948 , y6949 , y6950 , y6951 , y6952 , y6953 , y6954 , y6955 , y6956 , y6957 , y6958 , y6959 , y6960 , y6961 , y6962 , y6963 , y6964 , y6965 , y6966 , y6967 , y6968 , y6969 , y6970 , y6971 , y6972 , y6973 , y6974 , y6975 , y6976 , y6977 , y6978 , y6979 , y6980 , y6981 , y6982 , y6983 , y6984 , y6985 , y6986 , y6987 , y6988 , y6989 , y6990 , y6991 , y6992 , y6993 , y6994 , y6995 , y6996 , y6997 , y6998 , y6999 , y7000 , y7001 , y7002 , y7003 , y7004 , y7005 , y7006 , y7007 , y7008 , y7009 , y7010 , y7011 , y7012 , y7013 , y7014 , y7015 , y7016 , y7017 , y7018 , y7019 , y7020 , y7021 , y7022 , y7023 , y7024 , y7025 , y7026 , y7027 , y7028 , y7029 , y7030 , y7031 , y7032 , y7033 , y7034 , y7035 , y7036 , y7037 , y7038 , y7039 , y7040 , y7041 , y7042 , y7043 , y7044 , y7045 , y7046 , y7047 , y7048 , y7049 , y7050 , y7051 , y7052 , y7053 , y7054 , y7055 , y7056 , y7057 , y7058 , y7059 , y7060 , y7061 , y7062 , y7063 , y7064 , y7065 , y7066 , y7067 , y7068 , y7069 , y7070 , y7071 , y7072 , y7073 , y7074 , y7075 , y7076 , y7077 , y7078 , y7079 , y7080 , y7081 , y7082 , y7083 , y7084 , y7085 , y7086 , y7087 , y7088 , y7089 , y7090 , y7091 , y7092 , y7093 , y7094 , y7095 , y7096 , y7097 , y7098 , y7099 , y7100 , y7101 , y7102 , y7103 , y7104 , y7105 , y7106 , y7107 , y7108 , y7109 , y7110 , y7111 , y7112 , y7113 , y7114 , y7115 , y7116 , y7117 , y7118 , y7119 , y7120 , y7121 , y7122 , y7123 , y7124 , y7125 , y7126 , y7127 , y7128 , y7129 , y7130 , y7131 , y7132 , y7133 , y7134 , y7135 , y7136 , y7137 , y7138 , y7139 , y7140 , y7141 , y7142 , y7143 , y7144 , y7145 , y7146 , y7147 , y7148 , y7149 , y7150 , y7151 , y7152 , y7153 , y7154 , y7155 , y7156 , y7157 , y7158 , y7159 , y7160 , y7161 , y7162 , y7163 , y7164 , y7165 , y7166 , y7167 , y7168 , y7169 , y7170 , y7171 , y7172 , y7173 , y7174 , y7175 , y7176 , y7177 , y7178 , y7179 , y7180 , y7181 , y7182 , y7183 , y7184 , y7185 , y7186 , y7187 , y7188 , y7189 , y7190 , y7191 , y7192 , y7193 , y7194 , y7195 , y7196 , y7197 , y7198 , y7199 , y7200 , y7201 , y7202 , y7203 , y7204 , y7205 , y7206 , y7207 , y7208 , y7209 , y7210 , y7211 , y7212 , y7213 , y7214 , y7215 , y7216 , y7217 , y7218 , y7219 , y7220 , y7221 , y7222 , y7223 , y7224 , y7225 , y7226 , y7227 , y7228 , y7229 , y7230 , y7231 , y7232 , y7233 , y7234 , y7235 , y7236 , y7237 , y7238 , y7239 , y7240 , y7241 , y7242 , y7243 , y7244 , y7245 , y7246 , y7247 , y7248 , y7249 , y7250 , y7251 , y7252 , y7253 , y7254 , y7255 , y7256 , y7257 , y7258 , y7259 , y7260 , y7261 , y7262 , y7263 , y7264 , y7265 , y7266 , y7267 , y7268 , y7269 , y7270 , y7271 , y7272 , y7273 , y7274 , y7275 , y7276 , y7277 , y7278 , y7279 , y7280 , y7281 , y7282 , y7283 , y7284 , y7285 , y7286 , y7287 , y7288 , y7289 , y7290 , y7291 , y7292 , y7293 , y7294 , y7295 , y7296 , y7297 , y7298 , y7299 , y7300 , y7301 , y7302 , y7303 , y7304 , y7305 , y7306 , y7307 , y7308 , y7309 , y7310 , y7311 , y7312 , y7313 , y7314 , y7315 , y7316 , y7317 , y7318 , y7319 , y7320 , y7321 , y7322 , y7323 , y7324 , y7325 , y7326 , y7327 , y7328 , y7329 , y7330 , y7331 , y7332 , y7333 , y7334 , y7335 , y7336 , y7337 , y7338 , y7339 , y7340 , y7341 , y7342 , y7343 , y7344 , y7345 , y7346 , y7347 , y7348 , y7349 , y7350 , y7351 , y7352 , y7353 , y7354 , y7355 , y7356 , y7357 , y7358 , y7359 , y7360 , y7361 , y7362 , y7363 , y7364 , y7365 , y7366 , y7367 , y7368 , y7369 , y7370 , y7371 , y7372 , y7373 , y7374 , y7375 , y7376 , y7377 , y7378 , y7379 , y7380 , y7381 , y7382 , y7383 , y7384 , y7385 , y7386 , y7387 , y7388 , y7389 , y7390 , y7391 , y7392 , y7393 , y7394 , y7395 , y7396 , y7397 , y7398 , y7399 , y7400 , y7401 , y7402 , y7403 , y7404 , y7405 , y7406 , y7407 , y7408 , y7409 , y7410 , y7411 , y7412 , y7413 , y7414 , y7415 , y7416 , y7417 , y7418 , y7419 , y7420 , y7421 , y7422 , y7423 , y7424 , y7425 , y7426 , y7427 , y7428 , y7429 , y7430 , y7431 , y7432 , y7433 , y7434 , y7435 , y7436 , y7437 , y7438 , y7439 , y7440 , y7441 , y7442 , y7443 , y7444 , y7445 , y7446 , y7447 , y7448 , y7449 , y7450 , y7451 , y7452 , y7453 , y7454 , y7455 , y7456 , y7457 , y7458 , y7459 , y7460 , y7461 , y7462 , y7463 , y7464 , y7465 , y7466 , y7467 , y7468 , y7469 , y7470 , y7471 , y7472 , y7473 , y7474 , y7475 , y7476 , y7477 , y7478 , y7479 , y7480 , y7481 , y7482 , y7483 , y7484 , y7485 , y7486 , y7487 , y7488 , y7489 , y7490 , y7491 , y7492 , y7493 , y7494 , y7495 , y7496 , y7497 , y7498 , y7499 , y7500 , y7501 , y7502 , y7503 , y7504 , y7505 , y7506 , y7507 , y7508 , y7509 , y7510 , y7511 , y7512 , y7513 , y7514 , y7515 , y7516 , y7517 , y7518 , y7519 , y7520 , y7521 , y7522 , y7523 , y7524 , y7525 , y7526 , y7527 , y7528 , y7529 , y7530 , y7531 , y7532 , y7533 , y7534 , y7535 , y7536 , y7537 , y7538 , y7539 , y7540 , y7541 , y7542 , y7543 , y7544 , y7545 , y7546 , y7547 , y7548 , y7549 , y7550 , y7551 , y7552 , y7553 , y7554 , y7555 , y7556 , y7557 , y7558 , y7559 , y7560 , y7561 , y7562 , y7563 , y7564 , y7565 , y7566 , y7567 , y7568 , y7569 , y7570 , y7571 , y7572 , y7573 , y7574 , y7575 , y7576 , y7577 , y7578 , y7579 , y7580 , y7581 , y7582 , y7583 , y7584 , y7585 , y7586 , y7587 , y7588 , y7589 , y7590 , y7591 , y7592 , y7593 , y7594 , y7595 , y7596 , y7597 , y7598 , y7599 , y7600 , y7601 , y7602 , y7603 , y7604 , y7605 , y7606 , y7607 , y7608 , y7609 , y7610 , y7611 , y7612 , y7613 , y7614 , y7615 , y7616 , y7617 , y7618 , y7619 , y7620 , y7621 , y7622 , y7623 , y7624 , y7625 , y7626 , y7627 , y7628 , y7629 , y7630 , y7631 , y7632 , y7633 , y7634 , y7635 , y7636 , y7637 , y7638 , y7639 , y7640 , y7641 , y7642 , y7643 , y7644 , y7645 , y7646 , y7647 , y7648 , y7649 , y7650 , y7651 , y7652 , y7653 , y7654 , y7655 , y7656 , y7657 , y7658 , y7659 , y7660 , y7661 , y7662 , y7663 , y7664 , y7665 , y7666 , y7667 , y7668 , y7669 , y7670 , y7671 , y7672 , y7673 , y7674 , y7675 , y7676 , y7677 , y7678 , y7679 , y7680 , y7681 , y7682 , y7683 , y7684 , y7685 , y7686 , y7687 , y7688 , y7689 , y7690 , y7691 , y7692 , y7693 , y7694 , y7695 , y7696 , y7697 , y7698 , y7699 , y7700 , y7701 , y7702 , y7703 , y7704 , y7705 , y7706 , y7707 , y7708 , y7709 , y7710 , y7711 , y7712 , y7713 , y7714 , y7715 , y7716 , y7717 , y7718 , y7719 , y7720 , y7721 , y7722 , y7723 , y7724 , y7725 , y7726 , y7727 , y7728 , y7729 , y7730 , y7731 , y7732 , y7733 , y7734 , y7735 , y7736 , y7737 , y7738 , y7739 , y7740 , y7741 , y7742 , y7743 , y7744 , y7745 , y7746 , y7747 , y7748 , y7749 , y7750 , y7751 , y7752 , y7753 , y7754 , y7755 , y7756 , y7757 , y7758 , y7759 , y7760 , y7761 , y7762 , y7763 , y7764 , y7765 , y7766 , y7767 , y7768 , y7769 , y7770 , y7771 , y7772 , y7773 , y7774 , y7775 , y7776 , y7777 , y7778 , y7779 , y7780 , y7781 , y7782 , y7783 , y7784 , y7785 , y7786 , y7787 , y7788 , y7789 , y7790 , y7791 , y7792 , y7793 , y7794 , y7795 , y7796 , y7797 , y7798 , y7799 , y7800 , y7801 , y7802 , y7803 , y7804 , y7805 , y7806 , y7807 , y7808 , y7809 , y7810 , y7811 , y7812 , y7813 , y7814 , y7815 , y7816 , y7817 , y7818 , y7819 , y7820 , y7821 , y7822 , y7823 , y7824 , y7825 , y7826 , y7827 , y7828 , y7829 , y7830 , y7831 , y7832 , y7833 , y7834 , y7835 , y7836 , y7837 , y7838 , y7839 , y7840 , y7841 , y7842 , y7843 , y7844 , y7845 , y7846 , y7847 , y7848 , y7849 , y7850 , y7851 , y7852 , y7853 , y7854 , y7855 , y7856 , y7857 , y7858 , y7859 , y7860 , y7861 , y7862 , y7863 , y7864 , y7865 , y7866 , y7867 , y7868 , y7869 , y7870 , y7871 , y7872 , y7873 , y7874 , y7875 , y7876 , y7877 , y7878 , y7879 , y7880 , y7881 , y7882 , y7883 , y7884 , y7885 , y7886 , y7887 , y7888 , y7889 , y7890 , y7891 , y7892 , y7893 , y7894 , y7895 , y7896 , y7897 , y7898 , y7899 , y7900 , y7901 , y7902 , y7903 , y7904 , y7905 , y7906 , y7907 , y7908 , y7909 , y7910 , y7911 , y7912 , y7913 , y7914 , y7915 , y7916 , y7917 , y7918 , y7919 , y7920 , y7921 , y7922 , y7923 , y7924 , y7925 , y7926 , y7927 , y7928 , y7929 , y7930 , y7931 , y7932 , y7933 , y7934 , y7935 , y7936 , y7937 , y7938 , y7939 , y7940 , y7941 , y7942 , y7943 , y7944 , y7945 , y7946 , y7947 , y7948 , y7949 , y7950 , y7951 , y7952 , y7953 , y7954 , y7955 , y7956 , y7957 , y7958 , y7959 , y7960 , y7961 , y7962 , y7963 , y7964 , y7965 , y7966 , y7967 , y7968 , y7969 , y7970 , y7971 , y7972 , y7973 , y7974 , y7975 , y7976 , y7977 , y7978 , y7979 , y7980 , y7981 , y7982 , y7983 , y7984 , y7985 , y7986 , y7987 , y7988 , y7989 , y7990 , y7991 , y7992 , y7993 , y7994 , y7995 , y7996 , y7997 , y7998 , y7999 , y8000 , y8001 , y8002 , y8003 , y8004 , y8005 , y8006 , y8007 , y8008 , y8009 , y8010 , y8011 , y8012 , y8013 , y8014 , y8015 , y8016 , y8017 , y8018 , y8019 , y8020 , y8021 , y8022 , y8023 , y8024 , y8025 , y8026 , y8027 , y8028 , y8029 , y8030 , y8031 , y8032 , y8033 , y8034 , y8035 , y8036 , y8037 , y8038 , y8039 , y8040 , y8041 , y8042 , y8043 , y8044 , y8045 , y8046 , y8047 , y8048 , y8049 , y8050 , y8051 , y8052 , y8053 , y8054 , y8055 , y8056 , y8057 , y8058 , y8059 , y8060 , y8061 , y8062 , y8063 , y8064 , y8065 , y8066 , y8067 , y8068 , y8069 , y8070 , y8071 , y8072 , y8073 , y8074 , y8075 , y8076 , y8077 , y8078 , y8079 , y8080 , y8081 , y8082 , y8083 , y8084 , y8085 , y8086 , y8087 , y8088 , y8089 , y8090 , y8091 , y8092 , y8093 , y8094 , y8095 , y8096 , y8097 , y8098 , y8099 , y8100 , y8101 , y8102 , y8103 , y8104 , y8105 , y8106 , y8107 , y8108 , y8109 , y8110 , y8111 , y8112 , y8113 , y8114 , y8115 , y8116 , y8117 , y8118 , y8119 , y8120 , y8121 , y8122 , y8123 , y8124 , y8125 , y8126 , y8127 , y8128 , y8129 , y8130 , y8131 , y8132 , y8133 , y8134 , y8135 , y8136 , y8137 , y8138 , y8139 , y8140 , y8141 , y8142 , y8143 , y8144 , y8145 , y8146 , y8147 , y8148 , y8149 , y8150 , y8151 , y8152 , y8153 , y8154 , y8155 , y8156 , y8157 , y8158 , y8159 , y8160 , y8161 , y8162 , y8163 , y8164 , y8165 , y8166 , y8167 , y8168 , y8169 , y8170 , y8171 , y8172 , y8173 , y8174 , y8175 , y8176 , y8177 , y8178 , y8179 , y8180 , y8181 , y8182 , y8183 , y8184 , y8185 , y8186 , y8187 , y8188 , y8189 , y8190 , y8191 , y8192 , y8193 , y8194 , y8195 , y8196 , y8197 , y8198 , y8199 , y8200 , y8201 , y8202 , y8203 , y8204 , y8205 , y8206 , y8207 , y8208 , y8209 , y8210 , y8211 , y8212 , y8213 , y8214 , y8215 , y8216 , y8217 , y8218 , y8219 , y8220 , y8221 , y8222 , y8223 , y8224 , y8225 , y8226 , y8227 , y8228 , y8229 , y8230 , y8231 , y8232 , y8233 , y8234 , y8235 , y8236 , y8237 , y8238 , y8239 , y8240 , y8241 , y8242 , y8243 , y8244 , y8245 , y8246 , y8247 , y8248 , y8249 , y8250 , y8251 , y8252 , y8253 , y8254 , y8255 , y8256 , y8257 , y8258 , y8259 , y8260 , y8261 , y8262 , y8263 , y8264 , y8265 , y8266 , y8267 , y8268 , y8269 , y8270 , y8271 , y8272 , y8273 , y8274 , y8275 , y8276 , y8277 , y8278 , y8279 , y8280 , y8281 , y8282 , y8283 , y8284 , y8285 , y8286 , y8287 , y8288 , y8289 , y8290 , y8291 , y8292 , y8293 , y8294 , y8295 , y8296 , y8297 , y8298 , y8299 , y8300 , y8301 , y8302 , y8303 , y8304 , y8305 , y8306 , y8307 , y8308 , y8309 , y8310 , y8311 , y8312 , y8313 , y8314 , y8315 , y8316 , y8317 , y8318 , y8319 , y8320 , y8321 , y8322 , y8323 , y8324 , y8325 , y8326 , y8327 , y8328 , y8329 , y8330 , y8331 , y8332 , y8333 , y8334 , y8335 , y8336 , y8337 , y8338 , y8339 , y8340 , y8341 , y8342 , y8343 , y8344 , y8345 , y8346 , y8347 , y8348 , y8349 , y8350 , y8351 , y8352 , y8353 , y8354 , y8355 , y8356 , y8357 , y8358 , y8359 , y8360 , y8361 , y8362 , y8363 , y8364 , y8365 , y8366 , y8367 , y8368 , y8369 , y8370 , y8371 , y8372 , y8373 , y8374 , y8375 , y8376 , y8377 , y8378 , y8379 , y8380 , y8381 , y8382 , y8383 , y8384 , y8385 , y8386 , y8387 , y8388 , y8389 , y8390 , y8391 , y8392 , y8393 , y8394 , y8395 , y8396 , y8397 , y8398 , y8399 , y8400 , y8401 , y8402 , y8403 , y8404 , y8405 , y8406 , y8407 , y8408 , y8409 , y8410 , y8411 , y8412 , y8413 , y8414 , y8415 , y8416 , y8417 , y8418 , y8419 , y8420 , y8421 , y8422 , y8423 , y8424 , y8425 , y8426 , y8427 , y8428 , y8429 , y8430 , y8431 , y8432 , y8433 , y8434 , y8435 , y8436 , y8437 , y8438 , y8439 , y8440 , y8441 , y8442 , y8443 , y8444 , y8445 , y8446 , y8447 , y8448 , y8449 , y8450 , y8451 , y8452 , y8453 , y8454 , y8455 , y8456 , y8457 , y8458 , y8459 , y8460 , y8461 , y8462 , y8463 , y8464 , y8465 , y8466 , y8467 , y8468 , y8469 , y8470 , y8471 , y8472 , y8473 , y8474 , y8475 , y8476 , y8477 , y8478 , y8479 , y8480 , y8481 , y8482 , y8483 , y8484 , y8485 , y8486 , y8487 , y8488 , y8489 , y8490 , y8491 , y8492 , y8493 , y8494 , y8495 , y8496 , y8497 , y8498 , y8499 , y8500 , y8501 , y8502 , y8503 , y8504 , y8505 , y8506 , y8507 , y8508 , y8509 , y8510 , y8511 , y8512 , y8513 , y8514 , y8515 , y8516 , y8517 , y8518 , y8519 , y8520 , y8521 , y8522 , y8523 , y8524 , y8525 , y8526 , y8527 , y8528 , y8529 , y8530 , y8531 , y8532 , y8533 , y8534 , y8535 , y8536 , y8537 , y8538 , y8539 , y8540 , y8541 , y8542 , y8543 , y8544 , y8545 , y8546 , y8547 , y8548 , y8549 , y8550 , y8551 , y8552 , y8553 , y8554 , y8555 , y8556 , y8557 , y8558 , y8559 , y8560 , y8561 , y8562 , y8563 , y8564 , y8565 , y8566 , y8567 , y8568 , y8569 , y8570 , y8571 , y8572 , y8573 , y8574 , y8575 , y8576 , y8577 , y8578 , y8579 , y8580 , y8581 , y8582 , y8583 , y8584 , y8585 , y8586 , y8587 , y8588 , y8589 , y8590 , y8591 , y8592 , y8593 , y8594 , y8595 , y8596 , y8597 , y8598 , y8599 , y8600 , y8601 , y8602 , y8603 , y8604 , y8605 , y8606 , y8607 , y8608 , y8609 , y8610 , y8611 , y8612 , y8613 , y8614 , y8615 , y8616 , y8617 , y8618 , y8619 , y8620 , y8621 , y8622 , y8623 , y8624 , y8625 , y8626 , y8627 , y8628 , y8629 , y8630 , y8631 , y8632 , y8633 , y8634 , y8635 , y8636 , y8637 , y8638 , y8639 , y8640 , y8641 , y8642 , y8643 , y8644 , y8645 , y8646 , y8647 , y8648 , y8649 , y8650 , y8651 , y8652 , y8653 , y8654 , y8655 , y8656 , y8657 , y8658 , y8659 , y8660 , y8661 , y8662 , y8663 , y8664 , y8665 , y8666 , y8667 , y8668 , y8669 , y8670 , y8671 , y8672 , y8673 , y8674 , y8675 , y8676 , y8677 , y8678 , y8679 , y8680 , y8681 , y8682 , y8683 , y8684 , y8685 , y8686 , y8687 , y8688 , y8689 , y8690 , y8691 , y8692 , y8693 , y8694 , y8695 , y8696 , y8697 , y8698 , y8699 , y8700 , y8701 , y8702 , y8703 , y8704 , y8705 , y8706 , y8707 , y8708 , y8709 , y8710 , y8711 , y8712 , y8713 , y8714 , y8715 , y8716 , y8717 , y8718 , y8719 , y8720 , y8721 , y8722 , y8723 , y8724 , y8725 , y8726 , y8727 , y8728 , y8729 , y8730 , y8731 , y8732 , y8733 , y8734 , y8735 , y8736 , y8737 , y8738 , y8739 , y8740 , y8741 , y8742 , y8743 , y8744 , y8745 , y8746 , y8747 , y8748 , y8749 , y8750 , y8751 , y8752 , y8753 , y8754 , y8755 , y8756 , y8757 , y8758 , y8759 , y8760 , y8761 , y8762 , y8763 , y8764 , y8765 , y8766 , y8767 , y8768 , y8769 , y8770 , y8771 , y8772 , y8773 , y8774 , y8775 , y8776 , y8777 , y8778 , y8779 , y8780 , y8781 , y8782 , y8783 , y8784 , y8785 , y8786 , y8787 , y8788 , y8789 , y8790 , y8791 , y8792 , y8793 , y8794 , y8795 , y8796 , y8797 , y8798 , y8799 , y8800 , y8801 , y8802 , y8803 , y8804 , y8805 , y8806 , y8807 , y8808 , y8809 , y8810 , y8811 , y8812 , y8813 , y8814 , y8815 , y8816 , y8817 , y8818 , y8819 , y8820 , y8821 , y8822 , y8823 , y8824 , y8825 , y8826 , y8827 , y8828 , y8829 , y8830 , y8831 , y8832 , y8833 , y8834 , y8835 , y8836 , y8837 , y8838 , y8839 , y8840 , y8841 , y8842 , y8843 , y8844 , y8845 , y8846 , y8847 , y8848 , y8849 , y8850 , y8851 , y8852 , y8853 , y8854 , y8855 , y8856 , y8857 , y8858 , y8859 , y8860 , y8861 , y8862 , y8863 , y8864 , y8865 , y8866 , y8867 , y8868 , y8869 , y8870 , y8871 , y8872 , y8873 , y8874 , y8875 , y8876 , y8877 , y8878 , y8879 , y8880 , y8881 , y8882 , y8883 , y8884 , y8885 , y8886 , y8887 , y8888 , y8889 , y8890 , y8891 , y8892 , y8893 , y8894 , y8895 , y8896 , y8897 , y8898 , y8899 , y8900 , y8901 , y8902 , y8903 , y8904 , y8905 , y8906 , y8907 , y8908 , y8909 , y8910 , y8911 , y8912 , y8913 , y8914 , y8915 , y8916 , y8917 , y8918 , y8919 , y8920 , y8921 , y8922 , y8923 , y8924 , y8925 , y8926 , y8927 , y8928 , y8929 , y8930 , y8931 , y8932 , y8933 , y8934 , y8935 , y8936 , y8937 , y8938 , y8939 , y8940 , y8941 , y8942 , y8943 , y8944 , y8945 , y8946 , y8947 , y8948 , y8949 , y8950 , y8951 , y8952 , y8953 , y8954 , y8955 , y8956 , y8957 , y8958 , y8959 , y8960 , y8961 , y8962 , y8963 , y8964 , y8965 , y8966 , y8967 , y8968 , y8969 , y8970 , y8971 , y8972 , y8973 , y8974 , y8975 , y8976 , y8977 , y8978 , y8979 , y8980 , y8981 , y8982 , y8983 , y8984 , y8985 , y8986 , y8987 , y8988 , y8989 , y8990 , y8991 , y8992 , y8993 , y8994 , y8995 , y8996 , y8997 , y8998 , y8999 , y9000 , y9001 , y9002 , y9003 , y9004 , y9005 , y9006 , y9007 , y9008 , y9009 , y9010 , y9011 , y9012 , y9013 , y9014 , y9015 , y9016 , y9017 , y9018 , y9019 , y9020 , y9021 , y9022 , y9023 , y9024 , y9025 , y9026 , y9027 , y9028 , y9029 , y9030 , y9031 , y9032 , y9033 , y9034 , y9035 , y9036 , y9037 , y9038 , y9039 , y9040 , y9041 , y9042 , y9043 , y9044 , y9045 , y9046 , y9047 , y9048 , y9049 , y9050 , y9051 , y9052 , y9053 , y9054 , y9055 , y9056 , y9057 , y9058 , y9059 , y9060 , y9061 , y9062 , y9063 , y9064 , y9065 , y9066 , y9067 , y9068 , y9069 , y9070 , y9071 , y9072 , y9073 , y9074 , y9075 , y9076 , y9077 , y9078 , y9079 , y9080 , y9081 , y9082 , y9083 , y9084 , y9085 , y9086 , y9087 , y9088 , y9089 , y9090 , y9091 , y9092 , y9093 , y9094 , y9095 , y9096 , y9097 , y9098 , y9099 , y9100 , y9101 , y9102 , y9103 , y9104 , y9105 , y9106 , y9107 , y9108 , y9109 , y9110 , y9111 , y9112 , y9113 , y9114 , y9115 , y9116 , y9117 , y9118 , y9119 , y9120 , y9121 , y9122 , y9123 , y9124 , y9125 , y9126 , y9127 , y9128 , y9129 , y9130 , y9131 , y9132 , y9133 , y9134 , y9135 , y9136 , y9137 , y9138 , y9139 , y9140 , y9141 , y9142 , y9143 , y9144 , y9145 , y9146 , y9147 , y9148 , y9149 , y9150 , y9151 , y9152 , y9153 , y9154 , y9155 , y9156 , y9157 , y9158 , y9159 , y9160 , y9161 , y9162 , y9163 , y9164 , y9165 , y9166 , y9167 , y9168 , y9169 , y9170 , y9171 , y9172 , y9173 , y9174 , y9175 , y9176 , y9177 , y9178 , y9179 , y9180 , y9181 , y9182 , y9183 , y9184 , y9185 , y9186 , y9187 , y9188 , y9189 , y9190 , y9191 , y9192 , y9193 , y9194 , y9195 , y9196 , y9197 , y9198 , y9199 , y9200 , y9201 , y9202 , y9203 , y9204 , y9205 , y9206 , y9207 , y9208 , y9209 , y9210 , y9211 , y9212 , y9213 , y9214 , y9215 , y9216 , y9217 , y9218 , y9219 , y9220 , y9221 , y9222 , y9223 , y9224 , y9225 , y9226 , y9227 , y9228 , y9229 , y9230 , y9231 , y9232 , y9233 , y9234 , y9235 , y9236 , y9237 , y9238 , y9239 , y9240 , y9241 , y9242 , y9243 , y9244 , y9245 , y9246 , y9247 , y9248 , y9249 , y9250 , y9251 , y9252 , y9253 , y9254 , y9255 , y9256 , y9257 , y9258 , y9259 , y9260 , y9261 , y9262 , y9263 , y9264 , y9265 , y9266 , y9267 , y9268 , y9269 , y9270 , y9271 , y9272 , y9273 , y9274 , y9275 , y9276 , y9277 , y9278 , y9279 , y9280 , y9281 , y9282 , y9283 , y9284 , y9285 , y9286 , y9287 , y9288 , y9289 , y9290 , y9291 , y9292 , y9293 , y9294 , y9295 , y9296 , y9297 , y9298 , y9299 , y9300 , y9301 , y9302 , y9303 , y9304 , y9305 , y9306 , y9307 , y9308 , y9309 , y9310 , y9311 , y9312 , y9313 , y9314 , y9315 , y9316 , y9317 , y9318 , y9319 , y9320 , y9321 , y9322 , y9323 , y9324 , y9325 , y9326 , y9327 , y9328 , y9329 , y9330 , y9331 , y9332 , y9333 , y9334 , y9335 , y9336 , y9337 , y9338 , y9339 , y9340 , y9341 , y9342 , y9343 , y9344 , y9345 , y9346 , y9347 , y9348 , y9349 , y9350 , y9351 , y9352 , y9353 , y9354 , y9355 , y9356 , y9357 , y9358 , y9359 , y9360 , y9361 , y9362 , y9363 , y9364 , y9365 , y9366 , y9367 , y9368 , y9369 , y9370 , y9371 , y9372 , y9373 , y9374 , y9375 , y9376 , y9377 , y9378 , y9379 , y9380 , y9381 , y9382 , y9383 , y9384 , y9385 , y9386 , y9387 , y9388 , y9389 , y9390 , y9391 , y9392 , y9393 , y9394 , y9395 , y9396 , y9397 , y9398 , y9399 , y9400 , y9401 , y9402 , y9403 , y9404 , y9405 , y9406 , y9407 , y9408 , y9409 , y9410 , y9411 , y9412 , y9413 , y9414 , y9415 , y9416 , y9417 , y9418 , y9419 , y9420 , y9421 , y9422 , y9423 , y9424 , y9425 , y9426 , y9427 , y9428 , y9429 , y9430 , y9431 , y9432 , y9433 , y9434 , y9435 , y9436 , y9437 , y9438 , y9439 , y9440 , y9441 , y9442 , y9443 , y9444 , y9445 , y9446 , y9447 , y9448 , y9449 , y9450 , y9451 , y9452 , y9453 , y9454 , y9455 , y9456 , y9457 , y9458 , y9459 , y9460 , y9461 , y9462 , y9463 , y9464 , y9465 , y9466 , y9467 , y9468 , y9469 , y9470 , y9471 , y9472 , y9473 , y9474 , y9475 , y9476 , y9477 , y9478 , y9479 , y9480 , y9481 , y9482 , y9483 , y9484 , y9485 , y9486 , y9487 , y9488 , y9489 , y9490 , y9491 , y9492 , y9493 , y9494 , y9495 , y9496 , y9497 , y9498 , y9499 , y9500 , y9501 , y9502 , y9503 , y9504 , y9505 , y9506 , y9507 , y9508 , y9509 , y9510 , y9511 , y9512 , y9513 , y9514 , y9515 , y9516 , y9517 , y9518 , y9519 , y9520 , y9521 , y9522 , y9523 , y9524 , y9525 , y9526 , y9527 , y9528 , y9529 , y9530 , y9531 , y9532 , y9533 , y9534 , y9535 , y9536 , y9537 , y9538 , y9539 , y9540 , y9541 , y9542 , y9543 , y9544 , y9545 , y9546 , y9547 , y9548 , y9549 , y9550 , y9551 , y9552 , y9553 , y9554 , y9555 , y9556 , y9557 , y9558 , y9559 , y9560 , y9561 , y9562 , y9563 , y9564 , y9565 , y9566 , y9567 , y9568 , y9569 , y9570 , y9571 , y9572 , y9573 , y9574 , y9575 , y9576 , y9577 , y9578 , y9579 , y9580 , y9581 , y9582 , y9583 , y9584 , y9585 , y9586 , y9587 , y9588 , y9589 , y9590 , y9591 , y9592 , y9593 , y9594 , y9595 , y9596 , y9597 , y9598 , y9599 , y9600 , y9601 , y9602 , y9603 , y9604 , y9605 , y9606 , y9607 , y9608 , y9609 , y9610 , y9611 , y9612 , y9613 , y9614 , y9615 , y9616 , y9617 , y9618 , y9619 , y9620 , y9621 , y9622 , y9623 , y9624 , y9625 , y9626 , y9627 , y9628 , y9629 , y9630 , y9631 , y9632 , y9633 , y9634 , y9635 , y9636 , y9637 , y9638 , y9639 , y9640 , y9641 , y9642 , y9643 , y9644 , y9645 , y9646 , y9647 , y9648 , y9649 , y9650 , y9651 , y9652 , y9653 , y9654 , y9655 , y9656 , y9657 , y9658 , y9659 , y9660 , y9661 , y9662 , y9663 , y9664 , y9665 , y9666 , y9667 , y9668 , y9669 , y9670 , y9671 , y9672 , y9673 , y9674 , y9675 , y9676 , y9677 , y9678 , y9679 , y9680 , y9681 , y9682 , y9683 , y9684 , y9685 , y9686 , y9687 , y9688 , y9689 , y9690 , y9691 , y9692 , y9693 , y9694 , y9695 , y9696 , y9697 , y9698 , y9699 , y9700 , y9701 , y9702 , y9703 , y9704 , y9705 , y9706 , y9707 , y9708 , y9709 , y9710 , y9711 , y9712 , y9713 , y9714 , y9715 , y9716 , y9717 , y9718 , y9719 , y9720 , y9721 , y9722 , y9723 , y9724 , y9725 , y9726 , y9727 , y9728 , y9729 , y9730 , y9731 , y9732 , y9733 , y9734 , y9735 , y9736 , y9737 , y9738 , y9739 , y9740 , y9741 , y9742 , y9743 , y9744 , y9745 , y9746 , y9747 , y9748 , y9749 , y9750 , y9751 , y9752 , y9753 , y9754 , y9755 , y9756 , y9757 , y9758 , y9759 , y9760 , y9761 , y9762 , y9763 , y9764 , y9765 , y9766 , y9767 , y9768 , y9769 , y9770 , y9771 , y9772 , y9773 , y9774 , y9775 , y9776 , y9777 , y9778 , y9779 , y9780 , y9781 , y9782 , y9783 , y9784 , y9785 , y9786 , y9787 , y9788 , y9789 , y9790 , y9791 , y9792 , y9793 , y9794 , y9795 , y9796 , y9797 , y9798 , y9799 , y9800 , y9801 , y9802 , y9803 , y9804 , y9805 , y9806 , y9807 , y9808 , y9809 , y9810 , y9811 , y9812 , y9813 , y9814 , y9815 , y9816 , y9817 , y9818 , y9819 , y9820 , y9821 , y9822 , y9823 , y9824 , y9825 , y9826 , y9827 , y9828 , y9829 , y9830 , y9831 , y9832 , y9833 , y9834 , y9835 , y9836 , y9837 , y9838 , y9839 , y9840 , y9841 , y9842 , y9843 , y9844 , y9845 , y9846 , y9847 , y9848 , y9849 , y9850 , y9851 , y9852 , y9853 , y9854 , y9855 , y9856 , y9857 , y9858 , y9859 , y9860 , y9861 , y9862 , y9863 , y9864 , y9865 , y9866 , y9867 , y9868 , y9869 , y9870 , y9871 , y9872 , y9873 , y9874 , y9875 , y9876 , y9877 , y9878 , y9879 , y9880 , y9881 , y9882 , y9883 , y9884 , y9885 , y9886 , y9887 , y9888 , y9889 , y9890 , y9891 , y9892 , y9893 , y9894 , y9895 , y9896 , y9897 , y9898 , y9899 , y9900 , y9901 , y9902 , y9903 , y9904 , y9905 , y9906 , y9907 , y9908 , y9909 , y9910 , y9911 , y9912 , y9913 , y9914 , y9915 , y9916 , y9917 , y9918 , y9919 , y9920 , y9921 , y9922 , y9923 , y9924 , y9925 , y9926 , y9927 , y9928 , y9929 , y9930 , y9931 , y9932 , y9933 , y9934 , y9935 , y9936 , y9937 , y9938 , y9939 , y9940 , y9941 , y9942 , y9943 , y9944 , y9945 , y9946 , y9947 , y9948 , y9949 , y9950 , y9951 , y9952 , y9953 , y9954 , y9955 , y9956 , y9957 , y9958 , y9959 , y9960 , y9961 , y9962 , y9963 , y9964 , y9965 , y9966 , y9967 , y9968 , y9969 , y9970 , y9971 , y9972 , y9973 , y9974 , y9975 , y9976 , y9977 , y9978 , y9979 , y9980 , y9981 , y9982 , y9983 , y9984 , y9985 , y9986 , y9987 , y9988 , y9989 , y9990 , y9991 , y9992 , y9993 , y9994 , y9995 , y9996 , y9997 , y9998 , y9999 , y10000 , y10001 , y10002 , y10003 , y10004 , y10005 , y10006 , y10007 , y10008 , y10009 , y10010 , y10011 , y10012 , y10013 , y10014 , y10015 , y10016 , y10017 , y10018 , y10019 , y10020 , y10021 , y10022 , y10023 , y10024 , y10025 , y10026 , y10027 , y10028 , y10029 , y10030 , y10031 , y10032 , y10033 , y10034 , y10035 , y10036 , y10037 , y10038 , y10039 , y10040 , y10041 , y10042 , y10043 , y10044 , y10045 , y10046 , y10047 , y10048 , y10049 , y10050 , y10051 , y10052 , y10053 , y10054 , y10055 , y10056 , y10057 , y10058 , y10059 , y10060 , y10061 , y10062 , y10063 , y10064 , y10065 , y10066 , y10067 , y10068 , y10069 , y10070 , y10071 , y10072 , y10073 , y10074 , y10075 , y10076 , y10077 , y10078 , y10079 , y10080 , y10081 , y10082 , y10083 , y10084 , y10085 , y10086 , y10087 , y10088 , y10089 , y10090 , y10091 , y10092 , y10093 , y10094 , y10095 , y10096 , y10097 , y10098 , y10099 , y10100 , y10101 , y10102 , y10103 , y10104 , y10105 , y10106 , y10107 , y10108 , y10109 , y10110 , y10111 , y10112 , y10113 , y10114 , y10115 , y10116 , y10117 , y10118 , y10119 , y10120 , y10121 , y10122 , y10123 , y10124 , y10125 , y10126 , y10127 , y10128 , y10129 , y10130 , y10131 , y10132 , y10133 , y10134 , y10135 , y10136 , y10137 , y10138 , y10139 , y10140 , y10141 , y10142 , y10143 , y10144 , y10145 , y10146 , y10147 , y10148 , y10149 , y10150 , y10151 , y10152 , y10153 , y10154 , y10155 , y10156 , y10157 , y10158 , y10159 , y10160 , y10161 , y10162 , y10163 , y10164 , y10165 , y10166 , y10167 , y10168 , y10169 , y10170 , y10171 , y10172 , y10173 , y10174 , y10175 , y10176 , y10177 , y10178 , y10179 , y10180 , y10181 , y10182 , y10183 , y10184 , y10185 , y10186 , y10187 , y10188 , y10189 , y10190 , y10191 , y10192 , y10193 , y10194 , y10195 , y10196 , y10197 , y10198 , y10199 , y10200 , y10201 , y10202 , y10203 , y10204 , y10205 , y10206 , y10207 , y10208 , y10209 , y10210 , y10211 , y10212 , y10213 , y10214 , y10215 , y10216 , y10217 , y10218 , y10219 , y10220 , y10221 , y10222 , y10223 , y10224 , y10225 , y10226 , y10227 , y10228 , y10229 , y10230 , y10231 , y10232 , y10233 , y10234 , y10235 , y10236 , y10237 , y10238 , y10239 , y10240 , y10241 , y10242 , y10243 , y10244 , y10245 , y10246 , y10247 , y10248 , y10249 , y10250 , y10251 , y10252 , y10253 , y10254 , y10255 , y10256 , y10257 , y10258 , y10259 , y10260 , y10261 , y10262 , y10263 , y10264 , y10265 , y10266 , y10267 , y10268 , y10269 , y10270 , y10271 , y10272 , y10273 , y10274 , y10275 , y10276 , y10277 , y10278 , y10279 , y10280 , y10281 , y10282 , y10283 , y10284 , y10285 , y10286 , y10287 , y10288 , y10289 , y10290 , y10291 , y10292 , y10293 , y10294 , y10295 , y10296 , y10297 , y10298 , y10299 , y10300 , y10301 , y10302 , y10303 , y10304 , y10305 , y10306 , y10307 , y10308 , y10309 , y10310 , y10311 , y10312 , y10313 , y10314 , y10315 , y10316 , y10317 , y10318 , y10319 , y10320 , y10321 , y10322 , y10323 , y10324 , y10325 , y10326 , y10327 , y10328 , y10329 , y10330 , y10331 , y10332 , y10333 , y10334 , y10335 , y10336 , y10337 , y10338 , y10339 , y10340 , y10341 , y10342 , y10343 , y10344 , y10345 , y10346 , y10347 , y10348 , y10349 , y10350 , y10351 , y10352 , y10353 , y10354 , y10355 , y10356 , y10357 , y10358 , y10359 , y10360 , y10361 , y10362 , y10363 , y10364 , y10365 , y10366 , y10367 , y10368 , y10369 , y10370 , y10371 , y10372 , y10373 , y10374 , y10375 , y10376 , y10377 , y10378 , y10379 , y10380 , y10381 , y10382 , y10383 , y10384 , y10385 , y10386 , y10387 , y10388 , y10389 , y10390 , y10391 , y10392 , y10393 , y10394 , y10395 , y10396 , y10397 , y10398 , y10399 , y10400 , y10401 , y10402 , y10403 , y10404 , y10405 , y10406 , y10407 , y10408 , y10409 , y10410 , y10411 , y10412 , y10413 , y10414 , y10415 , y10416 , y10417 , y10418 , y10419 , y10420 , y10421 , y10422 , y10423 , y10424 , y10425 , y10426 , y10427 , y10428 , y10429 , y10430 , y10431 , y10432 , y10433 , y10434 , y10435 , y10436 , y10437 , y10438 , y10439 , y10440 , y10441 , y10442 , y10443 , y10444 , y10445 , y10446 , y10447 , y10448 , y10449 , y10450 , y10451 , y10452 , y10453 , y10454 , y10455 , y10456 , y10457 , y10458 , y10459 , y10460 , y10461 , y10462 , y10463 , y10464 , y10465 , y10466 , y10467 , y10468 , y10469 , y10470 , y10471 , y10472 , y10473 , y10474 , y10475 , y10476 , y10477 , y10478 , y10479 , y10480 , y10481 , y10482 , y10483 , y10484 , y10485 , y10486 , y10487 , y10488 , y10489 , y10490 , y10491 , y10492 , y10493 , y10494 , y10495 , y10496 , y10497 , y10498 , y10499 , y10500 , y10501 , y10502 , y10503 , y10504 , y10505 , y10506 , y10507 , y10508 , y10509 , y10510 , y10511 , y10512 , y10513 , y10514 , y10515 , y10516 , y10517 , y10518 , y10519 , y10520 , y10521 , y10522 , y10523 , y10524 , y10525 , y10526 , y10527 , y10528 , y10529 , y10530 , y10531 , y10532 , y10533 , y10534 , y10535 , y10536 , y10537 , y10538 , y10539 , y10540 , y10541 , y10542 , y10543 , y10544 , y10545 , y10546 , y10547 , y10548 , y10549 , y10550 , y10551 , y10552 , y10553 , y10554 , y10555 , y10556 , y10557 , y10558 , y10559 , y10560 , y10561 , y10562 , y10563 , y10564 , y10565 , y10566 , y10567 , y10568 , y10569 , y10570 , y10571 , y10572 , y10573 , y10574 , y10575 , y10576 , y10577 , y10578 , y10579 , y10580 , y10581 , y10582 , y10583 , y10584 , y10585 , y10586 , y10587 , y10588 , y10589 , y10590 , y10591 , y10592 , y10593 , y10594 , y10595 , y10596 , y10597 , y10598 , y10599 , y10600 , y10601 , y10602 , y10603 , y10604 , y10605 , y10606 , y10607 , y10608 , y10609 , y10610 , y10611 , y10612 , y10613 , y10614 , y10615 , y10616 , y10617 , y10618 , y10619 , y10620 , y10621 , y10622 , y10623 , y10624 , y10625 , y10626 , y10627 , y10628 , y10629 , y10630 , y10631 , y10632 , y10633 , y10634 , y10635 , y10636 , y10637 , y10638 , y10639 , y10640 , y10641 , y10642 , y10643 , y10644 , y10645 , y10646 , y10647 , y10648 , y10649 , y10650 , y10651 , y10652 , y10653 , y10654 , y10655 , y10656 , y10657 , y10658 , y10659 , y10660 , y10661 , y10662 , y10663 , y10664 , y10665 , y10666 , y10667 , y10668 , y10669 , y10670 , y10671 , y10672 , y10673 , y10674 , y10675 , y10676 , y10677 , y10678 , y10679 , y10680 , y10681 , y10682 , y10683 , y10684 , y10685 , y10686 , y10687 , y10688 , y10689 , y10690 , y10691 , y10692 , y10693 , y10694 , y10695 , y10696 , y10697 , y10698 , y10699 , y10700 , y10701 , y10702 , y10703 , y10704 , y10705 , y10706 , y10707 , y10708 , y10709 , y10710 , y10711 , y10712 , y10713 , y10714 , y10715 , y10716 , y10717 , y10718 , y10719 , y10720 , y10721 , y10722 , y10723 , y10724 , y10725 , y10726 , y10727 , y10728 , y10729 , y10730 , y10731 , y10732 , y10733 , y10734 , y10735 , y10736 , y10737 , y10738 , y10739 , y10740 , y10741 , y10742 , y10743 , y10744 , y10745 , y10746 , y10747 , y10748 , y10749 , y10750 , y10751 , y10752 , y10753 , y10754 , y10755 , y10756 , y10757 , y10758 , y10759 , y10760 , y10761 , y10762 , y10763 , y10764 , y10765 , y10766 , y10767 , y10768 , y10769 , y10770 , y10771 , y10772 , y10773 , y10774 , y10775 , y10776 , y10777 , y10778 , y10779 , y10780 , y10781 , y10782 , y10783 , y10784 , y10785 , y10786 , y10787 , y10788 , y10789 , y10790 , y10791 , y10792 , y10793 , y10794 , y10795 , y10796 , y10797 , y10798 , y10799 , y10800 , y10801 , y10802 , y10803 , y10804 , y10805 , y10806 , y10807 , y10808 , y10809 , y10810 , y10811 , y10812 , y10813 , y10814 , y10815 , y10816 , y10817 , y10818 , y10819 , y10820 , y10821 , y10822 , y10823 , y10824 , y10825 , y10826 , y10827 , y10828 , y10829 , y10830 , y10831 , y10832 , y10833 , y10834 , y10835 , y10836 , y10837 , y10838 , y10839 , y10840 , y10841 , y10842 , y10843 , y10844 , y10845 , y10846 , y10847 , y10848 , y10849 , y10850 , y10851 , y10852 , y10853 , y10854 , y10855 , y10856 , y10857 , y10858 , y10859 , y10860 , y10861 , y10862 , y10863 , y10864 , y10865 , y10866 , y10867 , y10868 , y10869 , y10870 , y10871 , y10872 , y10873 , y10874 , y10875 , y10876 , y10877 , y10878 , y10879 , y10880 , y10881 , y10882 , y10883 , y10884 , y10885 , y10886 , y10887 , y10888 , y10889 , y10890 , y10891 , y10892 , y10893 , y10894 , y10895 , y10896 , y10897 , y10898 , y10899 , y10900 , y10901 , y10902 , y10903 , y10904 , y10905 , y10906 , y10907 , y10908 , y10909 , y10910 , y10911 , y10912 , y10913 , y10914 , y10915 , y10916 , y10917 , y10918 , y10919 , y10920 , y10921 , y10922 , y10923 , y10924 , y10925 , y10926 , y10927 , y10928 , y10929 , y10930 , y10931 , y10932 , y10933 , y10934 , y10935 , y10936 , y10937 , y10938 , y10939 , y10940 , y10941 , y10942 , y10943 , y10944 , y10945 , y10946 , y10947 , y10948 , y10949 , y10950 , y10951 , y10952 , y10953 , y10954 , y10955 , y10956 , y10957 , y10958 , y10959 , y10960 , y10961 , y10962 , y10963 , y10964 , y10965 , y10966 , y10967 , y10968 , y10969 , y10970 , y10971 , y10972 , y10973 , y10974 , y10975 , y10976 , y10977 , y10978 , y10979 , y10980 , y10981 , y10982 , y10983 , y10984 , y10985 , y10986 , y10987 , y10988 , y10989 , y10990 , y10991 , y10992 , y10993 , y10994 , y10995 , y10996 , y10997 , y10998 , y10999 , y11000 , y11001 , y11002 , y11003 , y11004 , y11005 , y11006 , y11007 , y11008 , y11009 , y11010 , y11011 , y11012 , y11013 , y11014 , y11015 , y11016 , y11017 , y11018 , y11019 , y11020 , y11021 , y11022 , y11023 , y11024 , y11025 , y11026 , y11027 , y11028 , y11029 , y11030 , y11031 , y11032 , y11033 , y11034 , y11035 , y11036 , y11037 , y11038 , y11039 , y11040 , y11041 , y11042 , y11043 , y11044 , y11045 , y11046 , y11047 , y11048 , y11049 , y11050 , y11051 , y11052 , y11053 , y11054 , y11055 , y11056 , y11057 , y11058 , y11059 , y11060 , y11061 , y11062 , y11063 , y11064 , y11065 , y11066 , y11067 , y11068 , y11069 , y11070 , y11071 , y11072 , y11073 , y11074 , y11075 , y11076 , y11077 , y11078 , y11079 , y11080 , y11081 , y11082 , y11083 , y11084 , y11085 , y11086 , y11087 , y11088 , y11089 , y11090 , y11091 , y11092 , y11093 , y11094 , y11095 , y11096 , y11097 , y11098 , y11099 , y11100 , y11101 , y11102 , y11103 , y11104 , y11105 , y11106 , y11107 , y11108 , y11109 , y11110 , y11111 , y11112 , y11113 , y11114 , y11115 , y11116 , y11117 , y11118 , y11119 , y11120 , y11121 , y11122 , y11123 , y11124 , y11125 , y11126 , y11127 , y11128 , y11129 , y11130 , y11131 , y11132 , y11133 , y11134 , y11135 , y11136 , y11137 , y11138 , y11139 , y11140 , y11141 , y11142 , y11143 , y11144 , y11145 , y11146 , y11147 , y11148 , y11149 , y11150 , y11151 , y11152 , y11153 , y11154 , y11155 , y11156 , y11157 , y11158 , y11159 , y11160 , y11161 , y11162 , y11163 , y11164 , y11165 , y11166 , y11167 , y11168 , y11169 , y11170 , y11171 , y11172 , y11173 , y11174 , y11175 , y11176 , y11177 , y11178 , y11179 , y11180 , y11181 , y11182 , y11183 , y11184 , y11185 , y11186 , y11187 , y11188 , y11189 , y11190 , y11191 , y11192 , y11193 , y11194 , y11195 , y11196 , y11197 , y11198 , y11199 , y11200 , y11201 , y11202 , y11203 , y11204 , y11205 , y11206 , y11207 , y11208 , y11209 , y11210 , y11211 , y11212 , y11213 , y11214 , y11215 , y11216 , y11217 , y11218 , y11219 , y11220 , y11221 , y11222 , y11223 , y11224 , y11225 , y11226 , y11227 , y11228 , y11229 , y11230 , y11231 , y11232 , y11233 , y11234 , y11235 , y11236 , y11237 , y11238 , y11239 , y11240 , y11241 , y11242 , y11243 , y11244 , y11245 , y11246 , y11247 , y11248 , y11249 , y11250 , y11251 , y11252 , y11253 , y11254 , y11255 , y11256 , y11257 , y11258 , y11259 , y11260 , y11261 , y11262 , y11263 , y11264 , y11265 , y11266 , y11267 , y11268 , y11269 , y11270 , y11271 , y11272 , y11273 , y11274 , y11275 , y11276 , y11277 , y11278 , y11279 , y11280 , y11281 , y11282 , y11283 , y11284 , y11285 , y11286 , y11287 , y11288 , y11289 , y11290 , y11291 , y11292 , y11293 , y11294 , y11295 , y11296 , y11297 , y11298 , y11299 , y11300 , y11301 , y11302 , y11303 , y11304 , y11305 , y11306 , y11307 , y11308 , y11309 , y11310 , y11311 , y11312 , y11313 , y11314 , y11315 , y11316 , y11317 , y11318 , y11319 , y11320 , y11321 , y11322 , y11323 , y11324 , y11325 , y11326 , y11327 , y11328 , y11329 , y11330 , y11331 , y11332 , y11333 , y11334 , y11335 , y11336 , y11337 , y11338 , y11339 , y11340 , y11341 , y11342 , y11343 , y11344 , y11345 , y11346 , y11347 , y11348 , y11349 , y11350 , y11351 , y11352 , y11353 , y11354 , y11355 , y11356 , y11357 , y11358 , y11359 , y11360 , y11361 , y11362 , y11363 , y11364 , y11365 , y11366 , y11367 , y11368 , y11369 , y11370 , y11371 , y11372 , y11373 , y11374 , y11375 , y11376 , y11377 , y11378 , y11379 , y11380 , y11381 , y11382 , y11383 , y11384 , y11385 , y11386 , y11387 , y11388 , y11389 , y11390 , y11391 , y11392 , y11393 , y11394 , y11395 , y11396 , y11397 , y11398 , y11399 , y11400 , y11401 , y11402 , y11403 , y11404 , y11405 , y11406 , y11407 , y11408 , y11409 , y11410 , y11411 , y11412 , y11413 , y11414 , y11415 , y11416 , y11417 , y11418 , y11419 , y11420 , y11421 , y11422 , y11423 , y11424 , y11425 , y11426 , y11427 , y11428 , y11429 , y11430 , y11431 , y11432 , y11433 , y11434 , y11435 , y11436 , y11437 , y11438 , y11439 , y11440 , y11441 , y11442 , y11443 , y11444 , y11445 , y11446 , y11447 , y11448 , y11449 , y11450 , y11451 , y11452 , y11453 , y11454 , y11455 , y11456 , y11457 , y11458 , y11459 , y11460 , y11461 , y11462 , y11463 , y11464 , y11465 , y11466 , y11467 , y11468 , y11469 , y11470 , y11471 , y11472 , y11473 , y11474 , y11475 , y11476 , y11477 , y11478 , y11479 , y11480 , y11481 , y11482 , y11483 , y11484 , y11485 , y11486 , y11487 , y11488 , y11489 , y11490 , y11491 , y11492 , y11493 , y11494 , y11495 , y11496 , y11497 , y11498 , y11499 , y11500 , y11501 , y11502 , y11503 , y11504 , y11505 , y11506 , y11507 , y11508 , y11509 , y11510 , y11511 , y11512 , y11513 , y11514 , y11515 , y11516 , y11517 , y11518 , y11519 , y11520 , y11521 , y11522 , y11523 , y11524 , y11525 , y11526 , y11527 , y11528 , y11529 , y11530 , y11531 , y11532 , y11533 , y11534 , y11535 , y11536 , y11537 , y11538 , y11539 , y11540 , y11541 , y11542 , y11543 , y11544 , y11545 , y11546 , y11547 , y11548 , y11549 , y11550 , y11551 , y11552 , y11553 , y11554 , y11555 , y11556 , y11557 , y11558 , y11559 , y11560 , y11561 , y11562 , y11563 , y11564 , y11565 , y11566 , y11567 , y11568 , y11569 , y11570 , y11571 , y11572 , y11573 , y11574 , y11575 , y11576 , y11577 , y11578 , y11579 , y11580 , y11581 , y11582 , y11583 , y11584 , y11585 , y11586 , y11587 , y11588 , y11589 , y11590 , y11591 , y11592 , y11593 , y11594 , y11595 , y11596 , y11597 , y11598 , y11599 , y11600 , y11601 , y11602 , y11603 , y11604 , y11605 , y11606 , y11607 , y11608 , y11609 , y11610 , y11611 , y11612 , y11613 , y11614 , y11615 , y11616 , y11617 , y11618 , y11619 , y11620 , y11621 , y11622 , y11623 , y11624 , y11625 , y11626 , y11627 , y11628 , y11629 , y11630 , y11631 , y11632 , y11633 , y11634 , y11635 , y11636 , y11637 , y11638 , y11639 , y11640 , y11641 , y11642 , y11643 , y11644 , y11645 , y11646 , y11647 , y11648 , y11649 , y11650 , y11651 , y11652 , y11653 , y11654 , y11655 , y11656 , y11657 , y11658 , y11659 , y11660 , y11661 , y11662 , y11663 , y11664 , y11665 , y11666 , y11667 , y11668 , y11669 , y11670 , y11671 , y11672 , y11673 , y11674 , y11675 , y11676 , y11677 , y11678 , y11679 , y11680 , y11681 , y11682 , y11683 , y11684 , y11685 , y11686 , y11687 , y11688 , y11689 , y11690 , y11691 , y11692 , y11693 , y11694 , y11695 , y11696 , y11697 , y11698 , y11699 , y11700 , y11701 , y11702 , y11703 , y11704 , y11705 , y11706 , y11707 , y11708 , y11709 , y11710 , y11711 , y11712 , y11713 , y11714 , y11715 , y11716 , y11717 , y11718 , y11719 , y11720 , y11721 , y11722 , y11723 , y11724 , y11725 , y11726 , y11727 , y11728 , y11729 , y11730 , y11731 , y11732 , y11733 , y11734 , y11735 , y11736 , y11737 , y11738 , y11739 , y11740 , y11741 , y11742 , y11743 , y11744 , y11745 , y11746 , y11747 , y11748 , y11749 , y11750 , y11751 , y11752 , y11753 , y11754 , y11755 , y11756 , y11757 , y11758 , y11759 , y11760 , y11761 , y11762 , y11763 , y11764 , y11765 , y11766 , y11767 , y11768 , y11769 , y11770 , y11771 , y11772 , y11773 , y11774 , y11775 , y11776 , y11777 , y11778 , y11779 , y11780 , y11781 , y11782 , y11783 , y11784 , y11785 , y11786 , y11787 , y11788 , y11789 , y11790 , y11791 , y11792 , y11793 , y11794 , y11795 , y11796 , y11797 , y11798 , y11799 , y11800 , y11801 , y11802 , y11803 , y11804 , y11805 , y11806 , y11807 , y11808 , y11809 , y11810 , y11811 , y11812 , y11813 , y11814 , y11815 , y11816 , y11817 , y11818 , y11819 , y11820 , y11821 , y11822 , y11823 , y11824 , y11825 , y11826 , y11827 , y11828 , y11829 , y11830 , y11831 , y11832 , y11833 , y11834 , y11835 , y11836 , y11837 , y11838 , y11839 , y11840 , y11841 , y11842 , y11843 , y11844 , y11845 , y11846 , y11847 , y11848 , y11849 , y11850 , y11851 , y11852 , y11853 , y11854 , y11855 , y11856 , y11857 , y11858 , y11859 , y11860 , y11861 , y11862 , y11863 , y11864 , y11865 , y11866 , y11867 , y11868 , y11869 , y11870 , y11871 , y11872 , y11873 , y11874 , y11875 , y11876 , y11877 , y11878 , y11879 , y11880 , y11881 , y11882 , y11883 , y11884 , y11885 , y11886 , y11887 , y11888 , y11889 , y11890 , y11891 , y11892 , y11893 , y11894 , y11895 , y11896 , y11897 , y11898 , y11899 , y11900 , y11901 , y11902 , y11903 , y11904 , y11905 , y11906 , y11907 , y11908 , y11909 , y11910 , y11911 , y11912 , y11913 , y11914 , y11915 , y11916 , y11917 , y11918 , y11919 , y11920 , y11921 , y11922 , y11923 , y11924 , y11925 , y11926 , y11927 , y11928 , y11929 , y11930 , y11931 , y11932 , y11933 , y11934 , y11935 , y11936 , y11937 , y11938 , y11939 , y11940 , y11941 , y11942 , y11943 , y11944 , y11945 , y11946 , y11947 , y11948 , y11949 , y11950 , y11951 , y11952 , y11953 , y11954 , y11955 , y11956 , y11957 , y11958 , y11959 , y11960 , y11961 , y11962 , y11963 , y11964 , y11965 , y11966 , y11967 , y11968 , y11969 , y11970 , y11971 , y11972 , y11973 , y11974 , y11975 , y11976 , y11977 , y11978 , y11979 , y11980 , y11981 , y11982 , y11983 , y11984 , y11985 , y11986 , y11987 , y11988 , y11989 , y11990 , y11991 , y11992 , y11993 , y11994 , y11995 , y11996 , y11997 , y11998 , y11999 , y12000 , y12001 , y12002 , y12003 , y12004 , y12005 , y12006 , y12007 , y12008 , y12009 , y12010 , y12011 , y12012 , y12013 , y12014 , y12015 , y12016 , y12017 , y12018 , y12019 , y12020 , y12021 , y12022 , y12023 , y12024 , y12025 , y12026 , y12027 , y12028 , y12029 , y12030 , y12031 , y12032 , y12033 , y12034 , y12035 , y12036 , y12037 , y12038 , y12039 , y12040 , y12041 , y12042 , y12043 , y12044 , y12045 , y12046 , y12047 , y12048 , y12049 , y12050 , y12051 , y12052 , y12053 , y12054 , y12055 , y12056 , y12057 , y12058 , y12059 , y12060 , y12061 , y12062 , y12063 , y12064 , y12065 , y12066 , y12067 , y12068 , y12069 , y12070 , y12071 , y12072 , y12073 , y12074 , y12075 , y12076 , y12077 , y12078 , y12079 , y12080 , y12081 , y12082 , y12083 , y12084 , y12085 , y12086 , y12087 , y12088 , y12089 , y12090 , y12091 , y12092 , y12093 , y12094 , y12095 , y12096 , y12097 , y12098 , y12099 , y12100 , y12101 , y12102 , y12103 , y12104 , y12105 , y12106 , y12107 , y12108 , y12109 , y12110 , y12111 , y12112 , y12113 , y12114 , y12115 , y12116 , y12117 , y12118 , y12119 , y12120 , y12121 , y12122 , y12123 , y12124 , y12125 , y12126 , y12127 , y12128 , y12129 , y12130 , y12131 , y12132 , y12133 , y12134 , y12135 , y12136 , y12137 , y12138 , y12139 , y12140 , y12141 , y12142 , y12143 , y12144 , y12145 , y12146 , y12147 , y12148 , y12149 , y12150 , y12151 , y12152 , y12153 , y12154 , y12155 , y12156 , y12157 , y12158 , y12159 , y12160 , y12161 , y12162 , y12163 , y12164 , y12165 , y12166 , y12167 , y12168 , y12169 , y12170 , y12171 , y12172 , y12173 , y12174 , y12175 , y12176 , y12177 , y12178 , y12179 , y12180 , y12181 , y12182 , y12183 , y12184 , y12185 , y12186 , y12187 , y12188 , y12189 , y12190 , y12191 , y12192 , y12193 , y12194 , y12195 , y12196 , y12197 , y12198 , y12199 , y12200 , y12201 , y12202 , y12203 , y12204 , y12205 , y12206 , y12207 , y12208 , y12209 , y12210 , y12211 , y12212 , y12213 , y12214 , y12215 , y12216 , y12217 , y12218 , y12219 , y12220 , y12221 , y12222 , y12223 , y12224 , y12225 , y12226 , y12227 , y12228 , y12229 , y12230 , y12231 , y12232 , y12233 , y12234 , y12235 , y12236 , y12237 , y12238 , y12239 , y12240 , y12241 , y12242 , y12243 , y12244 , y12245 , y12246 , y12247 , y12248 , y12249 , y12250 , y12251 , y12252 , y12253 , y12254 , y12255 , y12256 , y12257 , y12258 , y12259 , y12260 , y12261 , y12262 , y12263 , y12264 , y12265 , y12266 , y12267 , y12268 , y12269 , y12270 , y12271 , y12272 , y12273 , y12274 , y12275 , y12276 , y12277 , y12278 , y12279 , y12280 , y12281 , y12282 , y12283 , y12284 , y12285 , y12286 , y12287 , y12288 , y12289 , y12290 , y12291 , y12292 , y12293 , y12294 , y12295 , y12296 , y12297 , y12298 , y12299 , y12300 , y12301 , y12302 , y12303 , y12304 , y12305 , y12306 , y12307 , y12308 , y12309 , y12310 , y12311 , y12312 , y12313 , y12314 , y12315 , y12316 , y12317 , y12318 , y12319 , y12320 , y12321 , y12322 , y12323 , y12324 , y12325 , y12326 , y12327 , y12328 , y12329 , y12330 , y12331 , y12332 , y12333 , y12334 , y12335 , y12336 , y12337 , y12338 , y12339 , y12340 , y12341 , y12342 , y12343 , y12344 , y12345 , y12346 , y12347 , y12348 , y12349 , y12350 , y12351 , y12352 , y12353 , y12354 , y12355 , y12356 , y12357 , y12358 , y12359 , y12360 , y12361 , y12362 , y12363 , y12364 , y12365 , y12366 , y12367 , y12368 , y12369 , y12370 , y12371 , y12372 , y12373 , y12374 , y12375 , y12376 , y12377 , y12378 , y12379 , y12380 , y12381 , y12382 , y12383 , y12384 , y12385 , y12386 , y12387 , y12388 , y12389 , y12390 , y12391 , y12392 , y12393 , y12394 , y12395 , y12396 , y12397 , y12398 , y12399 , y12400 , y12401 , y12402 , y12403 , y12404 , y12405 , y12406 , y12407 , y12408 , y12409 , y12410 , y12411 , y12412 , y12413 , y12414 , y12415 , y12416 , y12417 , y12418 , y12419 , y12420 , y12421 , y12422 , y12423 , y12424 , y12425 , y12426 , y12427 , y12428 , y12429 , y12430 , y12431 , y12432 , y12433 , y12434 , y12435 , y12436 , y12437 , y12438 , y12439 , y12440 , y12441 , y12442 , y12443 , y12444 , y12445 , y12446 , y12447 , y12448 , y12449 , y12450 , y12451 , y12452 , y12453 , y12454 , y12455 , y12456 , y12457 , y12458 , y12459 , y12460 , y12461 , y12462 , y12463 , y12464 , y12465 , y12466 , y12467 , y12468 , y12469 , y12470 , y12471 , y12472 , y12473 , y12474 , y12475 , y12476 , y12477 , y12478 , y12479 , y12480 , y12481 , y12482 , y12483 , y12484 , y12485 , y12486 , y12487 , y12488 , y12489 , y12490 , y12491 , y12492 , y12493 , y12494 , y12495 , y12496 , y12497 , y12498 , y12499 , y12500 , y12501 , y12502 , y12503 , y12504 , y12505 , y12506 , y12507 , y12508 , y12509 , y12510 , y12511 , y12512 , y12513 , y12514 , y12515 , y12516 , y12517 , y12518 , y12519 , y12520 , y12521 , y12522 , y12523 , y12524 , y12525 , y12526 , y12527 , y12528 , y12529 , y12530 , y12531 , y12532 , y12533 , y12534 , y12535 , y12536 , y12537 , y12538 , y12539 , y12540 , y12541 , y12542 , y12543 , y12544 , y12545 , y12546 , y12547 , y12548 , y12549 , y12550 , y12551 , y12552 , y12553 , y12554 , y12555 , y12556 , y12557 , y12558 , y12559 , y12560 , y12561 , y12562 , y12563 , y12564 , y12565 , y12566 , y12567 , y12568 , y12569 , y12570 , y12571 , y12572 , y12573 , y12574 , y12575 , y12576 , y12577 , y12578 , y12579 , y12580 , y12581 , y12582 , y12583 , y12584 , y12585 , y12586 , y12587 , y12588 , y12589 , y12590 , y12591 , y12592 , y12593 , y12594 , y12595 , y12596 , y12597 , y12598 , y12599 , y12600 , y12601 , y12602 , y12603 , y12604 , y12605 , y12606 , y12607 , y12608 , y12609 , y12610 , y12611 , y12612 , y12613 , y12614 , y12615 , y12616 , y12617 , y12618 , y12619 , y12620 , y12621 , y12622 , y12623 , y12624 , y12625 , y12626 , y12627 , y12628 , y12629 , y12630 , y12631 , y12632 , y12633 , y12634 , y12635 , y12636 , y12637 , y12638 , y12639 , y12640 , y12641 , y12642 , y12643 , y12644 , y12645 , y12646 , y12647 , y12648 , y12649 , y12650 , y12651 , y12652 , y12653 , y12654 , y12655 , y12656 , y12657 , y12658 , y12659 , y12660 , y12661 , y12662 , y12663 , y12664 , y12665 , y12666 , y12667 , y12668 , y12669 , y12670 , y12671 , y12672 , y12673 , y12674 , y12675 , y12676 , y12677 , y12678 , y12679 , y12680 , y12681 , y12682 , y12683 , y12684 , y12685 , y12686 , y12687 , y12688 , y12689 , y12690 , y12691 , y12692 , y12693 , y12694 , y12695 , y12696 , y12697 , y12698 , y12699 , y12700 , y12701 , y12702 , y12703 , y12704 , y12705 , y12706 , y12707 , y12708 , y12709 , y12710 , y12711 , y12712 , y12713 , y12714 , y12715 , y12716 , y12717 , y12718 , y12719 , y12720 , y12721 , y12722 , y12723 , y12724 , y12725 , y12726 , y12727 , y12728 , y12729 , y12730 , y12731 , y12732 , y12733 , y12734 , y12735 , y12736 , y12737 , y12738 , y12739 , y12740 , y12741 , y12742 , y12743 , y12744 , y12745 , y12746 , y12747 , y12748 , y12749 , y12750 , y12751 , y12752 , y12753 , y12754 , y12755 , y12756 , y12757 , y12758 , y12759 , y12760 , y12761 , y12762 , y12763 , y12764 , y12765 , y12766 , y12767 , y12768 , y12769 , y12770 , y12771 , y12772 , y12773 , y12774 , y12775 , y12776 , y12777 , y12778 , y12779 , y12780 , y12781 , y12782 , y12783 , y12784 , y12785 , y12786 , y12787 , y12788 , y12789 , y12790 , y12791 , y12792 , y12793 , y12794 , y12795 , y12796 , y12797 , y12798 , y12799 , y12800 , y12801 , y12802 , y12803 , y12804 , y12805 , y12806 , y12807 , y12808 , y12809 , y12810 , y12811 , y12812 , y12813 , y12814 , y12815 , y12816 , y12817 , y12818 , y12819 , y12820 , y12821 , y12822 , y12823 , y12824 , y12825 , y12826 , y12827 , y12828 , y12829 , y12830 , y12831 , y12832 , y12833 , y12834 , y12835 , y12836 , y12837 , y12838 , y12839 , y12840 , y12841 , y12842 , y12843 , y12844 , y12845 , y12846 , y12847 , y12848 , y12849 , y12850 , y12851 , y12852 , y12853 , y12854 , y12855 , y12856 , y12857 , y12858 , y12859 , y12860 , y12861 , y12862 , y12863 , y12864 , y12865 , y12866 , y12867 , y12868 , y12869 , y12870 , y12871 , y12872 , y12873 , y12874 , y12875 , y12876 , y12877 , y12878 , y12879 , y12880 , y12881 , y12882 , y12883 , y12884 , y12885 , y12886 , y12887 , y12888 , y12889 , y12890 , y12891 , y12892 , y12893 , y12894 , y12895 , y12896 , y12897 , y12898 , y12899 , y12900 , y12901 , y12902 , y12903 , y12904 , y12905 , y12906 , y12907 , y12908 , y12909 , y12910 , y12911 , y12912 , y12913 , y12914 , y12915 , y12916 , y12917 , y12918 , y12919 , y12920 , y12921 , y12922 , y12923 , y12924 , y12925 , y12926 , y12927 , y12928 , y12929 , y12930 , y12931 , y12932 , y12933 , y12934 , y12935 , y12936 , y12937 , y12938 , y12939 , y12940 , y12941 , y12942 , y12943 , y12944 , y12945 , y12946 , y12947 , y12948 , y12949 , y12950 , y12951 , y12952 , y12953 , y12954 , y12955 , y12956 , y12957 , y12958 , y12959 , y12960 , y12961 , y12962 , y12963 , y12964 , y12965 , y12966 , y12967 , y12968 , y12969 , y12970 , y12971 , y12972 , y12973 , y12974 , y12975 , y12976 , y12977 , y12978 , y12979 , y12980 , y12981 , y12982 , y12983 , y12984 , y12985 , y12986 , y12987 , y12988 , y12989 , y12990 , y12991 , y12992 , y12993 , y12994 , y12995 , y12996 , y12997 , y12998 , y12999 , y13000 , y13001 , y13002 , y13003 , y13004 , y13005 , y13006 , y13007 , y13008 , y13009 , y13010 , y13011 , y13012 , y13013 , y13014 , y13015 , y13016 , y13017 , y13018 , y13019 , y13020 , y13021 , y13022 , y13023 , y13024 , y13025 , y13026 , y13027 , y13028 , y13029 , y13030 , y13031 , y13032 , y13033 , y13034 , y13035 , y13036 , y13037 , y13038 , y13039 , y13040 , y13041 , y13042 , y13043 , y13044 , y13045 , y13046 , y13047 , y13048 , y13049 , y13050 , y13051 , y13052 , y13053 , y13054 , y13055 , y13056 , y13057 , y13058 , y13059 , y13060 , y13061 , y13062 , y13063 , y13064 , y13065 , y13066 , y13067 , y13068 , y13069 , y13070 , y13071 , y13072 , y13073 , y13074 , y13075 , y13076 , y13077 , y13078 , y13079 , y13080 , y13081 , y13082 , y13083 , y13084 , y13085 , y13086 , y13087 , y13088 , y13089 , y13090 , y13091 , y13092 , y13093 , y13094 , y13095 , y13096 , y13097 , y13098 , y13099 , y13100 , y13101 , y13102 , y13103 , y13104 , y13105 , y13106 , y13107 , y13108 , y13109 , y13110 , y13111 , y13112 , y13113 , y13114 , y13115 , y13116 , y13117 , y13118 , y13119 , y13120 , y13121 , y13122 , y13123 , y13124 , y13125 , y13126 , y13127 , y13128 , y13129 , y13130 , y13131 , y13132 , y13133 , y13134 , y13135 , y13136 , y13137 , y13138 , y13139 , y13140 , y13141 , y13142 , y13143 , y13144 , y13145 , y13146 , y13147 , y13148 , y13149 , y13150 , y13151 , y13152 , y13153 , y13154 , y13155 , y13156 , y13157 , y13158 , y13159 , y13160 , y13161 , y13162 , y13163 , y13164 , y13165 , y13166 , y13167 , y13168 , y13169 , y13170 , y13171 , y13172 , y13173 , y13174 , y13175 , y13176 , y13177 , y13178 , y13179 , y13180 , y13181 , y13182 , y13183 , y13184 , y13185 , y13186 , y13187 , y13188 , y13189 , y13190 , y13191 , y13192 , y13193 , y13194 , y13195 , y13196 , y13197 , y13198 , y13199 , y13200 , y13201 , y13202 , y13203 , y13204 , y13205 , y13206 , y13207 , y13208 , y13209 , y13210 , y13211 , y13212 , y13213 , y13214 , y13215 , y13216 , y13217 , y13218 , y13219 , y13220 , y13221 , y13222 , y13223 , y13224 , y13225 , y13226 , y13227 , y13228 , y13229 , y13230 , y13231 , y13232 , y13233 , y13234 , y13235 , y13236 , y13237 , y13238 , y13239 , y13240 , y13241 , y13242 , y13243 , y13244 , y13245 , y13246 , y13247 , y13248 , y13249 , y13250 , y13251 , y13252 , y13253 , y13254 , y13255 , y13256 , y13257 , y13258 , y13259 , y13260 , y13261 , y13262 , y13263 , y13264 , y13265 , y13266 , y13267 , y13268 , y13269 , y13270 , y13271 , y13272 , y13273 , y13274 , y13275 , y13276 , y13277 , y13278 , y13279 , y13280 , y13281 , y13282 , y13283 , y13284 , y13285 , y13286 , y13287 , y13288 , y13289 , y13290 , y13291 , y13292 , y13293 , y13294 , y13295 , y13296 , y13297 , y13298 , y13299 , y13300 , y13301 , y13302 , y13303 , y13304 , y13305 , y13306 , y13307 , y13308 , y13309 , y13310 , y13311 , y13312 , y13313 , y13314 , y13315 , y13316 , y13317 , y13318 , y13319 , y13320 , y13321 , y13322 , y13323 , y13324 , y13325 , y13326 , y13327 , y13328 , y13329 , y13330 , y13331 , y13332 , y13333 , y13334 , y13335 , y13336 , y13337 , y13338 , y13339 , y13340 , y13341 , y13342 , y13343 , y13344 , y13345 , y13346 , y13347 , y13348 , y13349 , y13350 , y13351 , y13352 , y13353 , y13354 , y13355 , y13356 , y13357 , y13358 , y13359 , y13360 , y13361 , y13362 , y13363 , y13364 , y13365 , y13366 , y13367 , y13368 , y13369 , y13370 , y13371 , y13372 , y13373 , y13374 , y13375 , y13376 , y13377 , y13378 , y13379 , y13380 , y13381 , y13382 , y13383 , y13384 , y13385 , y13386 , y13387 , y13388 , y13389 , y13390 , y13391 , y13392 , y13393 , y13394 , y13395 , y13396 , y13397 , y13398 , y13399 , y13400 , y13401 , y13402 , y13403 , y13404 , y13405 , y13406 , y13407 , y13408 , y13409 , y13410 , y13411 , y13412 , y13413 , y13414 , y13415 , y13416 , y13417 , y13418 , y13419 , y13420 , y13421 , y13422 , y13423 , y13424 , y13425 , y13426 , y13427 , y13428 , y13429 , y13430 , y13431 , y13432 , y13433 , y13434 , y13435 , y13436 , y13437 , y13438 , y13439 , y13440 , y13441 , y13442 , y13443 , y13444 , y13445 , y13446 , y13447 , y13448 , y13449 , y13450 , y13451 , y13452 , y13453 , y13454 , y13455 , y13456 , y13457 , y13458 , y13459 , y13460 , y13461 , y13462 , y13463 , y13464 , y13465 , y13466 , y13467 , y13468 , y13469 , y13470 , y13471 , y13472 , y13473 , y13474 , y13475 , y13476 , y13477 , y13478 , y13479 , y13480 , y13481 , y13482 , y13483 , y13484 , y13485 , y13486 , y13487 , y13488 , y13489 , y13490 , y13491 , y13492 , y13493 , y13494 , y13495 , y13496 , y13497 , y13498 , y13499 , y13500 , y13501 , y13502 , y13503 , y13504 , y13505 , y13506 , y13507 , y13508 , y13509 , y13510 , y13511 , y13512 , y13513 , y13514 , y13515 , y13516 , y13517 , y13518 , y13519 , y13520 , y13521 , y13522 , y13523 , y13524 , y13525 , y13526 , y13527 , y13528 , y13529 , y13530 , y13531 , y13532 , y13533 , y13534 , y13535 , y13536 , y13537 , y13538 , y13539 , y13540 , y13541 , y13542 , y13543 , y13544 , y13545 , y13546 , y13547 , y13548 , y13549 , y13550 , y13551 , y13552 , y13553 , y13554 , y13555 , y13556 , y13557 , y13558 , y13559 , y13560 , y13561 , y13562 , y13563 , y13564 , y13565 , y13566 , y13567 , y13568 , y13569 , y13570 , y13571 , y13572 , y13573 , y13574 , y13575 , y13576 , y13577 , y13578 , y13579 , y13580 , y13581 , y13582 , y13583 , y13584 , y13585 , y13586 , y13587 , y13588 , y13589 , y13590 , y13591 , y13592 , y13593 , y13594 , y13595 , y13596 , y13597 , y13598 , y13599 , y13600 , y13601 , y13602 , y13603 , y13604 , y13605 , y13606 , y13607 , y13608 , y13609 , y13610 , y13611 , y13612 , y13613 , y13614 , y13615 , y13616 , y13617 , y13618 , y13619 , y13620 , y13621 , y13622 , y13623 , y13624 , y13625 , y13626 , y13627 , y13628 , y13629 , y13630 , y13631 , y13632 , y13633 , y13634 , y13635 , y13636 , y13637 , y13638 , y13639 , y13640 , y13641 , y13642 , y13643 , y13644 , y13645 , y13646 , y13647 , y13648 , y13649 , y13650 , y13651 , y13652 , y13653 , y13654 , y13655 , y13656 , y13657 , y13658 , y13659 , y13660 , y13661 , y13662 , y13663 , y13664 , y13665 , y13666 , y13667 , y13668 , y13669 , y13670 , y13671 , y13672 , y13673 , y13674 , y13675 , y13676 , y13677 , y13678 , y13679 , y13680 , y13681 , y13682 , y13683 , y13684 , y13685 , y13686 , y13687 , y13688 , y13689 , y13690 , y13691 , y13692 , y13693 , y13694 , y13695 , y13696 , y13697 , y13698 , y13699 , y13700 , y13701 , y13702 , y13703 , y13704 , y13705 , y13706 , y13707 , y13708 , y13709 , y13710 , y13711 , y13712 , y13713 , y13714 , y13715 , y13716 , y13717 , y13718 , y13719 , y13720 , y13721 , y13722 , y13723 , y13724 , y13725 , y13726 , y13727 , y13728 , y13729 , y13730 , y13731 , y13732 , y13733 , y13734 , y13735 , y13736 , y13737 , y13738 , y13739 , y13740 , y13741 , y13742 , y13743 , y13744 , y13745 , y13746 , y13747 , y13748 , y13749 , y13750 , y13751 , y13752 , y13753 , y13754 , y13755 , y13756 , y13757 , y13758 , y13759 , y13760 , y13761 , y13762 , y13763 , y13764 , y13765 , y13766 , y13767 , y13768 , y13769 , y13770 , y13771 , y13772 , y13773 , y13774 , y13775 , y13776 , y13777 , y13778 , y13779 , y13780 , y13781 , y13782 , y13783 , y13784 , y13785 , y13786 , y13787 , y13788 , y13789 , y13790 , y13791 , y13792 , y13793 , y13794 , y13795 , y13796 , y13797 , y13798 , y13799 , y13800 , y13801 , y13802 , y13803 , y13804 , y13805 , y13806 , y13807 , y13808 , y13809 , y13810 , y13811 , y13812 , y13813 , y13814 , y13815 , y13816 , y13817 , y13818 , y13819 , y13820 , y13821 , y13822 , y13823 , y13824 , y13825 , y13826 , y13827 , y13828 , y13829 , y13830 , y13831 , y13832 , y13833 , y13834 , y13835 , y13836 , y13837 , y13838 , y13839 , y13840 , y13841 , y13842 , y13843 , y13844 , y13845 , y13846 , y13847 , y13848 , y13849 , y13850 , y13851 , y13852 , y13853 , y13854 , y13855 , y13856 , y13857 , y13858 , y13859 , y13860 , y13861 , y13862 , y13863 , y13864 , y13865 , y13866 , y13867 , y13868 , y13869 , y13870 , y13871 , y13872 , y13873 , y13874 , y13875 , y13876 , y13877 , y13878 , y13879 , y13880 , y13881 , y13882 , y13883 , y13884 , y13885 , y13886 , y13887 , y13888 , y13889 , y13890 , y13891 , y13892 , y13893 , y13894 , y13895 , y13896 , y13897 , y13898 , y13899 , y13900 , y13901 , y13902 , y13903 , y13904 , y13905 , y13906 , y13907 , y13908 , y13909 , y13910 , y13911 , y13912 , y13913 , y13914 , y13915 , y13916 , y13917 , y13918 , y13919 , y13920 , y13921 , y13922 , y13923 , y13924 , y13925 , y13926 , y13927 , y13928 , y13929 , y13930 , y13931 , y13932 , y13933 , y13934 , y13935 , y13936 , y13937 , y13938 , y13939 , y13940 , y13941 , y13942 , y13943 , y13944 , y13945 , y13946 , y13947 , y13948 , y13949 , y13950 , y13951 , y13952 , y13953 , y13954 , y13955 , y13956 , y13957 , y13958 , y13959 , y13960 , y13961 , y13962 , y13963 , y13964 , y13965 , y13966 , y13967 , y13968 , y13969 , y13970 , y13971 , y13972 , y13973 , y13974 , y13975 , y13976 , y13977 , y13978 , y13979 , y13980 , y13981 , y13982 , y13983 , y13984 , y13985 , y13986 , y13987 , y13988 , y13989 , y13990 , y13991 , y13992 , y13993 , y13994 , y13995 , y13996 , y13997 , y13998 , y13999 , y14000 , y14001 , y14002 , y14003 , y14004 , y14005 , y14006 , y14007 , y14008 , y14009 , y14010 , y14011 , y14012 , y14013 , y14014 , y14015 , y14016 , y14017 , y14018 , y14019 , y14020 , y14021 , y14022 , y14023 , y14024 , y14025 , y14026 , y14027 , y14028 , y14029 , y14030 , y14031 , y14032 , y14033 , y14034 , y14035 , y14036 , y14037 , y14038 , y14039 , y14040 , y14041 , y14042 , y14043 , y14044 , y14045 , y14046 , y14047 , y14048 , y14049 , y14050 , y14051 , y14052 , y14053 , y14054 , y14055 , y14056 , y14057 , y14058 , y14059 , y14060 , y14061 , y14062 , y14063 , y14064 , y14065 , y14066 , y14067 , y14068 , y14069 , y14070 , y14071 , y14072 , y14073 , y14074 , y14075 , y14076 , y14077 , y14078 , y14079 , y14080 , y14081 , y14082 , y14083 , y14084 , y14085 , y14086 , y14087 , y14088 , y14089 , y14090 , y14091 , y14092 , y14093 , y14094 , y14095 , y14096 , y14097 , y14098 , y14099 , y14100 , y14101 , y14102 , y14103 , y14104 , y14105 , y14106 , y14107 , y14108 , y14109 , y14110 , y14111 , y14112 , y14113 , y14114 , y14115 , y14116 , y14117 , y14118 , y14119 , y14120 , y14121 , y14122 , y14123 , y14124 , y14125 , y14126 , y14127 , y14128 , y14129 , y14130 , y14131 , y14132 , y14133 , y14134 , y14135 , y14136 , y14137 , y14138 , y14139 , y14140 , y14141 , y14142 , y14143 , y14144 , y14145 , y14146 , y14147 , y14148 , y14149 , y14150 , y14151 , y14152 , y14153 , y14154 , y14155 , y14156 , y14157 , y14158 , y14159 , y14160 , y14161 , y14162 , y14163 , y14164 , y14165 , y14166 , y14167 , y14168 , y14169 , y14170 , y14171 , y14172 , y14173 , y14174 , y14175 , y14176 , y14177 , y14178 , y14179 , y14180 , y14181 , y14182 , y14183 , y14184 , y14185 , y14186 , y14187 , y14188 , y14189 , y14190 , y14191 , y14192 , y14193 , y14194 , y14195 , y14196 , y14197 , y14198 , y14199 , y14200 , y14201 , y14202 , y14203 , y14204 , y14205 , y14206 , y14207 , y14208 , y14209 , y14210 , y14211 , y14212 , y14213 , y14214 , y14215 , y14216 , y14217 , y14218 , y14219 , y14220 , y14221 , y14222 , y14223 , y14224 , y14225 , y14226 , y14227 , y14228 , y14229 , y14230 , y14231 , y14232 , y14233 , y14234 , y14235 , y14236 , y14237 , y14238 , y14239 , y14240 , y14241 , y14242 , y14243 , y14244 , y14245 , y14246 , y14247 , y14248 , y14249 , y14250 , y14251 , y14252 , y14253 , y14254 , y14255 , y14256 , y14257 , y14258 , y14259 , y14260 , y14261 , y14262 , y14263 , y14264 , y14265 , y14266 , y14267 , y14268 , y14269 , y14270 , y14271 , y14272 , y14273 , y14274 , y14275 , y14276 , y14277 , y14278 , y14279 , y14280 , y14281 , y14282 , y14283 , y14284 , y14285 , y14286 , y14287 , y14288 , y14289 , y14290 , y14291 , y14292 , y14293 , y14294 , y14295 , y14296 , y14297 , y14298 , y14299 , y14300 , y14301 , y14302 , y14303 , y14304 , y14305 , y14306 , y14307 , y14308 , y14309 , y14310 , y14311 , y14312 , y14313 , y14314 , y14315 , y14316 , y14317 , y14318 , y14319 , y14320 , y14321 , y14322 , y14323 , y14324 , y14325 , y14326 , y14327 , y14328 , y14329 , y14330 , y14331 , y14332 , y14333 , y14334 , y14335 , y14336 , y14337 , y14338 , y14339 , y14340 , y14341 , y14342 , y14343 , y14344 , y14345 , y14346 , y14347 , y14348 , y14349 , y14350 , y14351 , y14352 , y14353 , y14354 , y14355 , y14356 , y14357 , y14358 , y14359 , y14360 , y14361 , y14362 , y14363 , y14364 , y14365 , y14366 , y14367 , y14368 , y14369 , y14370 , y14371 , y14372 , y14373 , y14374 , y14375 , y14376 , y14377 , y14378 , y14379 , y14380 , y14381 , y14382 , y14383 , y14384 , y14385 , y14386 , y14387 , y14388 , y14389 , y14390 , y14391 , y14392 , y14393 , y14394 , y14395 , y14396 , y14397 , y14398 , y14399 , y14400 , y14401 , y14402 , y14403 , y14404 , y14405 , y14406 , y14407 , y14408 , y14409 , y14410 , y14411 , y14412 , y14413 , y14414 , y14415 , y14416 , y14417 , y14418 , y14419 , y14420 , y14421 , y14422 , y14423 , y14424 , y14425 , y14426 , y14427 , y14428 , y14429 , y14430 , y14431 , y14432 , y14433 , y14434 , y14435 , y14436 , y14437 , y14438 , y14439 , y14440 , y14441 , y14442 , y14443 , y14444 , y14445 , y14446 , y14447 , y14448 , y14449 , y14450 , y14451 , y14452 , y14453 , y14454 , y14455 , y14456 , y14457 , y14458 , y14459 , y14460 , y14461 , y14462 , y14463 , y14464 , y14465 , y14466 , y14467 , y14468 , y14469 , y14470 , y14471 , y14472 , y14473 , y14474 , y14475 , y14476 , y14477 , y14478 , y14479 , y14480 , y14481 , y14482 , y14483 , y14484 , y14485 , y14486 , y14487 , y14488 , y14489 , y14490 , y14491 , y14492 , y14493 , y14494 , y14495 , y14496 , y14497 , y14498 , y14499 , y14500 , y14501 , y14502 , y14503 , y14504 , y14505 , y14506 , y14507 , y14508 , y14509 , y14510 , y14511 , y14512 , y14513 , y14514 , y14515 , y14516 , y14517 , y14518 , y14519 , y14520 , y14521 , y14522 , y14523 , y14524 , y14525 , y14526 , y14527 , y14528 , y14529 , y14530 , y14531 , y14532 , y14533 , y14534 , y14535 , y14536 , y14537 , y14538 , y14539 , y14540 , y14541 , y14542 , y14543 , y14544 , y14545 , y14546 , y14547 , y14548 , y14549 , y14550 , y14551 , y14552 , y14553 , y14554 , y14555 , y14556 , y14557 , y14558 , y14559 , y14560 , y14561 , y14562 , y14563 , y14564 , y14565 , y14566 , y14567 , y14568 , y14569 , y14570 , y14571 , y14572 , y14573 , y14574 , y14575 , y14576 , y14577 , y14578 , y14579 , y14580 , y14581 , y14582 , y14583 , y14584 , y14585 , y14586 , y14587 , y14588 , y14589 , y14590 , y14591 , y14592 , y14593 , y14594 , y14595 , y14596 , y14597 , y14598 , y14599 , y14600 , y14601 , y14602 , y14603 , y14604 , y14605 , y14606 , y14607 , y14608 , y14609 , y14610 , y14611 , y14612 , y14613 , y14614 , y14615 , y14616 , y14617 , y14618 , y14619 , y14620 , y14621 , y14622 , y14623 , y14624 , y14625 , y14626 , y14627 , y14628 , y14629 , y14630 , y14631 , y14632 , y14633 , y14634 , y14635 , y14636 , y14637 , y14638 , y14639 , y14640 , y14641 , y14642 , y14643 , y14644 , y14645 , y14646 , y14647 , y14648 , y14649 , y14650 , y14651 , y14652 , y14653 , y14654 , y14655 , y14656 , y14657 , y14658 , y14659 , y14660 , y14661 , y14662 , y14663 , y14664 , y14665 , y14666 , y14667 , y14668 , y14669 , y14670 , y14671 , y14672 , y14673 , y14674 , y14675 , y14676 , y14677 , y14678 , y14679 , y14680 , y14681 , y14682 , y14683 , y14684 , y14685 , y14686 , y14687 , y14688 , y14689 , y14690 , y14691 , y14692 , y14693 , y14694 , y14695 , y14696 , y14697 , y14698 , y14699 , y14700 , y14701 , y14702 , y14703 , y14704 , y14705 , y14706 , y14707 , y14708 , y14709 , y14710 , y14711 , y14712 , y14713 , y14714 , y14715 , y14716 , y14717 , y14718 , y14719 , y14720 , y14721 , y14722 , y14723 , y14724 , y14725 , y14726 , y14727 , y14728 , y14729 , y14730 , y14731 , y14732 , y14733 , y14734 , y14735 , y14736 , y14737 , y14738 , y14739 , y14740 , y14741 , y14742 , y14743 , y14744 , y14745 , y14746 , y14747 , y14748 , y14749 , y14750 , y14751 , y14752 , y14753 , y14754 , y14755 , y14756 , y14757 , y14758 , y14759 , y14760 , y14761 , y14762 , y14763 , y14764 , y14765 , y14766 , y14767 , y14768 , y14769 , y14770 , y14771 , y14772 , y14773 , y14774 , y14775 , y14776 , y14777 , y14778 , y14779 , y14780 , y14781 , y14782 , y14783 , y14784 , y14785 , y14786 , y14787 , y14788 , y14789 , y14790 , y14791 , y14792 , y14793 , y14794 , y14795 , y14796 , y14797 , y14798 , y14799 , y14800 , y14801 , y14802 , y14803 , y14804 , y14805 , y14806 , y14807 , y14808 , y14809 , y14810 , y14811 , y14812 , y14813 , y14814 , y14815 , y14816 , y14817 , y14818 , y14819 , y14820 , y14821 , y14822 , y14823 , y14824 , y14825 , y14826 , y14827 , y14828 , y14829 , y14830 , y14831 , y14832 , y14833 , y14834 , y14835 , y14836 , y14837 , y14838 , y14839 , y14840 , y14841 , y14842 , y14843 , y14844 , y14845 , y14846 , y14847 , y14848 , y14849 , y14850 , y14851 , y14852 , y14853 , y14854 , y14855 , y14856 , y14857 , y14858 , y14859 , y14860 , y14861 , y14862 , y14863 , y14864 , y14865 , y14866 , y14867 , y14868 , y14869 , y14870 , y14871 , y14872 , y14873 , y14874 , y14875 , y14876 , y14877 , y14878 , y14879 , y14880 , y14881 , y14882 , y14883 , y14884 , y14885 , y14886 , y14887 , y14888 , y14889 , y14890 , y14891 , y14892 , y14893 , y14894 , y14895 , y14896 , y14897 , y14898 , y14899 , y14900 , y14901 , y14902 , y14903 , y14904 , y14905 , y14906 , y14907 , y14908 , y14909 , y14910 , y14911 , y14912 , y14913 , y14914 , y14915 , y14916 , y14917 , y14918 , y14919 , y14920 , y14921 , y14922 , y14923 , y14924 , y14925 , y14926 , y14927 , y14928 , y14929 , y14930 , y14931 , y14932 , y14933 , y14934 , y14935 , y14936 , y14937 , y14938 , y14939 , y14940 , y14941 , y14942 , y14943 , y14944 , y14945 , y14946 , y14947 , y14948 , y14949 , y14950 , y14951 , y14952 , y14953 , y14954 , y14955 , y14956 , y14957 , y14958 , y14959 , y14960 , y14961 , y14962 , y14963 , y14964 , y14965 , y14966 , y14967 , y14968 , y14969 , y14970 , y14971 , y14972 , y14973 , y14974 , y14975 , y14976 , y14977 , y14978 , y14979 , y14980 , y14981 , y14982 , y14983 , y14984 , y14985 , y14986 , y14987 , y14988 , y14989 , y14990 , y14991 , y14992 , y14993 , y14994 , y14995 , y14996 , y14997 , y14998 , y14999 , y15000 , y15001 , y15002 , y15003 , y15004 , y15005 , y15006 , y15007 , y15008 , y15009 , y15010 , y15011 , y15012 , y15013 , y15014 , y15015 , y15016 , y15017 , y15018 , y15019 , y15020 , y15021 , y15022 , y15023 , y15024 , y15025 , y15026 , y15027 , y15028 , y15029 , y15030 , y15031 , y15032 , y15033 , y15034 , y15035 , y15036 , y15037 , y15038 , y15039 , y15040 , y15041 , y15042 , y15043 , y15044 , y15045 , y15046 , y15047 , y15048 , y15049 , y15050 , y15051 , y15052 , y15053 , y15054 , y15055 , y15056 , y15057 , y15058 , y15059 , y15060 , y15061 , y15062 , y15063 , y15064 , y15065 , y15066 , y15067 , y15068 , y15069 , y15070 , y15071 , y15072 , y15073 , y15074 , y15075 , y15076 , y15077 , y15078 , y15079 , y15080 , y15081 , y15082 , y15083 , y15084 , y15085 , y15086 , y15087 , y15088 , y15089 , y15090 , y15091 , y15092 , y15093 , y15094 , y15095 , y15096 , y15097 , y15098 , y15099 , y15100 , y15101 , y15102 , y15103 , y15104 , y15105 , y15106 , y15107 , y15108 , y15109 , y15110 , y15111 , y15112 , y15113 , y15114 , y15115 , y15116 , y15117 , y15118 , y15119 , y15120 , y15121 , y15122 , y15123 , y15124 , y15125 , y15126 , y15127 , y15128 , y15129 , y15130 , y15131 , y15132 , y15133 , y15134 , y15135 , y15136 , y15137 , y15138 , y15139 , y15140 , y15141 , y15142 , y15143 , y15144 , y15145 , y15146 , y15147 , y15148 , y15149 , y15150 , y15151 , y15152 , y15153 , y15154 , y15155 , y15156 , y15157 , y15158 , y15159 , y15160 , y15161 , y15162 , y15163 , y15164 , y15165 , y15166 , y15167 , y15168 , y15169 , y15170 , y15171 , y15172 , y15173 , y15174 , y15175 , y15176 , y15177 , y15178 , y15179 , y15180 , y15181 , y15182 , y15183 , y15184 , y15185 , y15186 , y15187 , y15188 , y15189 , y15190 , y15191 , y15192 , y15193 , y15194 , y15195 , y15196 , y15197 , y15198 , y15199 , y15200 , y15201 , y15202 , y15203 , y15204 , y15205 , y15206 , y15207 , y15208 , y15209 , y15210 , y15211 , y15212 , y15213 , y15214 , y15215 , y15216 , y15217 , y15218 , y15219 , y15220 , y15221 , y15222 , y15223 , y15224 , y15225 , y15226 , y15227 , y15228 , y15229 , y15230 , y15231 , y15232 , y15233 , y15234 , y15235 , y15236 , y15237 , y15238 , y15239 , y15240 , y15241 , y15242 , y15243 , y15244 , y15245 , y15246 , y15247 , y15248 , y15249 , y15250 , y15251 , y15252 , y15253 , y15254 , y15255 , y15256 , y15257 , y15258 , y15259 , y15260 , y15261 , y15262 , y15263 , y15264 , y15265 , y15266 , y15267 , y15268 , y15269 , y15270 , y15271 , y15272 , y15273 , y15274 , y15275 , y15276 , y15277 , y15278 , y15279 , y15280 , y15281 , y15282 , y15283 , y15284 , y15285 , y15286 , y15287 , y15288 , y15289 , y15290 , y15291 , y15292 , y15293 , y15294 , y15295 , y15296 , y15297 , y15298 , y15299 , y15300 , y15301 , y15302 , y15303 , y15304 , y15305 , y15306 , y15307 , y15308 , y15309 , y15310 , y15311 , y15312 , y15313 , y15314 , y15315 , y15316 , y15317 , y15318 , y15319 , y15320 , y15321 , y15322 , y15323 , y15324 , y15325 , y15326 , y15327 , y15328 , y15329 , y15330 , y15331 , y15332 , y15333 , y15334 , y15335 , y15336 , y15337 , y15338 , y15339 , y15340 , y15341 , y15342 , y15343 , y15344 , y15345 , y15346 , y15347 , y15348 , y15349 , y15350 , y15351 , y15352 , y15353 , y15354 , y15355 , y15356 , y15357 , y15358 , y15359 , y15360 , y15361 , y15362 , y15363 , y15364 , y15365 , y15366 , y15367 , y15368 , y15369 , y15370 , y15371 , y15372 , y15373 , y15374 , y15375 , y15376 , y15377 , y15378 , y15379 , y15380 , y15381 , y15382 , y15383 , y15384 , y15385 , y15386 , y15387 , y15388 , y15389 , y15390 , y15391 , y15392 , y15393 , y15394 , y15395 , y15396 , y15397 , y15398 , y15399 , y15400 , y15401 , y15402 , y15403 , y15404 , y15405 , y15406 , y15407 , y15408 , y15409 , y15410 , y15411 , y15412 , y15413 , y15414 , y15415 , y15416 , y15417 , y15418 , y15419 , y15420 , y15421 , y15422 , y15423 , y15424 , y15425 , y15426 , y15427 , y15428 , y15429 , y15430 , y15431 , y15432 , y15433 , y15434 , y15435 , y15436 , y15437 , y15438 , y15439 , y15440 , y15441 , y15442 , y15443 , y15444 , y15445 , y15446 , y15447 , y15448 , y15449 , y15450 , y15451 , y15452 , y15453 , y15454 , y15455 , y15456 , y15457 , y15458 , y15459 , y15460 , y15461 , y15462 , y15463 , y15464 , y15465 , y15466 , y15467 , y15468 , y15469 , y15470 , y15471 , y15472 , y15473 , y15474 , y15475 , y15476 , y15477 , y15478 , y15479 , y15480 , y15481 , y15482 , y15483 , y15484 , y15485 , y15486 , y15487 , y15488 , y15489 , y15490 , y15491 , y15492 , y15493 , y15494 , y15495 , y15496 , y15497 , y15498 , y15499 , y15500 , y15501 , y15502 , y15503 , y15504 , y15505 , y15506 , y15507 , y15508 , y15509 , y15510 , y15511 , y15512 , y15513 , y15514 , y15515 , y15516 , y15517 , y15518 , y15519 , y15520 , y15521 , y15522 , y15523 , y15524 , y15525 , y15526 , y15527 , y15528 , y15529 , y15530 , y15531 , y15532 , y15533 , y15534 , y15535 , y15536 , y15537 , y15538 , y15539 , y15540 , y15541 , y15542 , y15543 , y15544 , y15545 , y15546 , y15547 , y15548 , y15549 , y15550 , y15551 , y15552 , y15553 , y15554 , y15555 , y15556 , y15557 , y15558 , y15559 , y15560 , y15561 , y15562 , y15563 , y15564 , y15565 , y15566 , y15567 , y15568 , y15569 , y15570 , y15571 , y15572 , y15573 , y15574 , y15575 , y15576 , y15577 , y15578 , y15579 , y15580 , y15581 , y15582 , y15583 , y15584 , y15585 , y15586 , y15587 , y15588 , y15589 , y15590 , y15591 , y15592 , y15593 , y15594 , y15595 , y15596 , y15597 , y15598 , y15599 , y15600 , y15601 , y15602 , y15603 , y15604 , y15605 , y15606 , y15607 , y15608 , y15609 , y15610 , y15611 , y15612 , y15613 , y15614 , y15615 , y15616 , y15617 , y15618 , y15619 , y15620 , y15621 , y15622 , y15623 , y15624 , y15625 , y15626 , y15627 , y15628 , y15629 , y15630 , y15631 , y15632 , y15633 , y15634 , y15635 , y15636 , y15637 , y15638 , y15639 , y15640 , y15641 , y15642 , y15643 , y15644 , y15645 , y15646 , y15647 , y15648 , y15649 , y15650 , y15651 , y15652 , y15653 , y15654 , y15655 , y15656 , y15657 , y15658 , y15659 , y15660 , y15661 , y15662 , y15663 , y15664 , y15665 , y15666 , y15667 , y15668 , y15669 , y15670 , y15671 , y15672 , y15673 , y15674 , y15675 , y15676 , y15677 , y15678 , y15679 , y15680 , y15681 , y15682 , y15683 , y15684 , y15685 , y15686 , y15687 , y15688 , y15689 , y15690 , y15691 , y15692 , y15693 , y15694 , y15695 , y15696 , y15697 , y15698 , y15699 , y15700 , y15701 , y15702 , y15703 , y15704 , y15705 , y15706 , y15707 , y15708 , y15709 , y15710 , y15711 , y15712 , y15713 , y15714 , y15715 , y15716 , y15717 , y15718 , y15719 , y15720 , y15721 , y15722 , y15723 , y15724 , y15725 , y15726 , y15727 , y15728 , y15729 , y15730 , y15731 , y15732 , y15733 , y15734 , y15735 , y15736 , y15737 , y15738 , y15739 , y15740 , y15741 , y15742 , y15743 , y15744 , y15745 , y15746 , y15747 , y15748 , y15749 , y15750 , y15751 , y15752 , y15753 , y15754 , y15755 , y15756 , y15757 , y15758 , y15759 , y15760 , y15761 , y15762 , y15763 , y15764 , y15765 , y15766 , y15767 , y15768 , y15769 , y15770 , y15771 , y15772 , y15773 , y15774 , y15775 , y15776 , y15777 , y15778 , y15779 , y15780 , y15781 , y15782 , y15783 , y15784 , y15785 , y15786 , y15787 , y15788 , y15789 , y15790 , y15791 , y15792 , y15793 , y15794 , y15795 , y15796 , y15797 , y15798 , y15799 , y15800 , y15801 , y15802 , y15803 , y15804 , y15805 , y15806 , y15807 , y15808 , y15809 , y15810 , y15811 , y15812 , y15813 , y15814 , y15815 , y15816 , y15817 , y15818 , y15819 , y15820 , y15821 , y15822 , y15823 , y15824 , y15825 , y15826 , y15827 , y15828 , y15829 , y15830 , y15831 , y15832 , y15833 , y15834 , y15835 , y15836 , y15837 , y15838 , y15839 , y15840 , y15841 , y15842 , y15843 , y15844 , y15845 , y15846 , y15847 , y15848 , y15849 , y15850 , y15851 , y15852 , y15853 , y15854 , y15855 , y15856 , y15857 , y15858 , y15859 , y15860 , y15861 , y15862 , y15863 , y15864 , y15865 , y15866 , y15867 , y15868 , y15869 , y15870 , y15871 , y15872 , y15873 , y15874 , y15875 , y15876 , y15877 , y15878 , y15879 , y15880 , y15881 , y15882 , y15883 , y15884 , y15885 , y15886 , y15887 , y15888 , y15889 , y15890 , y15891 , y15892 , y15893 , y15894 , y15895 , y15896 , y15897 , y15898 , y15899 , y15900 , y15901 , y15902 , y15903 , y15904 , y15905 , y15906 , y15907 , y15908 , y15909 , y15910 , y15911 , y15912 , y15913 , y15914 , y15915 , y15916 , y15917 , y15918 , y15919 , y15920 , y15921 , y15922 , y15923 , y15924 , y15925 , y15926 , y15927 , y15928 , y15929 , y15930 , y15931 , y15932 , y15933 , y15934 , y15935 , y15936 , y15937 , y15938 , y15939 , y15940 , y15941 , y15942 , y15943 , y15944 , y15945 , y15946 , y15947 , y15948 , y15949 , y15950 , y15951 , y15952 , y15953 , y15954 , y15955 , y15956 , y15957 , y15958 , y15959 , y15960 , y15961 , y15962 , y15963 , y15964 , y15965 , y15966 , y15967 , y15968 , y15969 , y15970 , y15971 , y15972 , y15973 , y15974 , y15975 , y15976 , y15977 , y15978 , y15979 , y15980 , y15981 , y15982 , y15983 , y15984 , y15985 , y15986 , y15987 , y15988 , y15989 , y15990 , y15991 , y15992 , y15993 , y15994 , y15995 , y15996 , y15997 , y15998 , y15999 , y16000 , y16001 , y16002 , y16003 , y16004 , y16005 , y16006 , y16007 , y16008 , y16009 , y16010 , y16011 , y16012 , y16013 , y16014 , y16015 , y16016 , y16017 , y16018 , y16019 , y16020 , y16021 , y16022 , y16023 , y16024 , y16025 , y16026 , y16027 , y16028 , y16029 , y16030 , y16031 , y16032 , y16033 , y16034 , y16035 , y16036 , y16037 , y16038 , y16039 , y16040 , y16041 , y16042 , y16043 , y16044 , y16045 , y16046 , y16047 , y16048 , y16049 , y16050 , y16051 , y16052 , y16053 , y16054 , y16055 , y16056 , y16057 , y16058 , y16059 , y16060 , y16061 , y16062 , y16063 , y16064 , y16065 , y16066 , y16067 , y16068 , y16069 , y16070 , y16071 , y16072 , y16073 , y16074 , y16075 , y16076 , y16077 , y16078 , y16079 , y16080 , y16081 , y16082 , y16083 , y16084 , y16085 , y16086 , y16087 , y16088 , y16089 , y16090 , y16091 , y16092 , y16093 , y16094 , y16095 , y16096 , y16097 , y16098 , y16099 , y16100 , y16101 , y16102 , y16103 , y16104 , y16105 , y16106 , y16107 , y16108 , y16109 , y16110 , y16111 , y16112 , y16113 , y16114 , y16115 , y16116 , y16117 , y16118 , y16119 , y16120 , y16121 , y16122 , y16123 , y16124 , y16125 , y16126 , y16127 , y16128 , y16129 , y16130 , y16131 , y16132 , y16133 , y16134 , y16135 , y16136 , y16137 , y16138 , y16139 , y16140 , y16141 , y16142 , y16143 , y16144 , y16145 , y16146 , y16147 , y16148 , y16149 , y16150 , y16151 , y16152 , y16153 , y16154 , y16155 , y16156 , y16157 , y16158 , y16159 , y16160 , y16161 , y16162 , y16163 , y16164 , y16165 , y16166 , y16167 , y16168 , y16169 , y16170 , y16171 , y16172 , y16173 , y16174 , y16175 , y16176 , y16177 , y16178 , y16179 , y16180 , y16181 , y16182 , y16183 , y16184 , y16185 , y16186 , y16187 , y16188 , y16189 , y16190 , y16191 , y16192 , y16193 , y16194 , y16195 , y16196 , y16197 , y16198 , y16199 , y16200 , y16201 , y16202 , y16203 , y16204 , y16205 , y16206 , y16207 , y16208 , y16209 , y16210 , y16211 , y16212 , y16213 , y16214 , y16215 , y16216 , y16217 , y16218 , y16219 , y16220 , y16221 , y16222 , y16223 , y16224 , y16225 , y16226 , y16227 , y16228 , y16229 , y16230 , y16231 , y16232 , y16233 , y16234 , y16235 , y16236 , y16237 , y16238 , y16239 , y16240 , y16241 , y16242 , y16243 , y16244 , y16245 , y16246 , y16247 , y16248 , y16249 , y16250 , y16251 , y16252 , y16253 , y16254 , y16255 , y16256 , y16257 , y16258 , y16259 , y16260 , y16261 , y16262 , y16263 , y16264 , y16265 , y16266 , y16267 , y16268 , y16269 , y16270 , y16271 , y16272 , y16273 , y16274 , y16275 , y16276 , y16277 , y16278 , y16279 , y16280 , y16281 , y16282 , y16283 , y16284 , y16285 , y16286 , y16287 , y16288 , y16289 , y16290 , y16291 , y16292 , y16293 , y16294 , y16295 , y16296 , y16297 , y16298 , y16299 , y16300 , y16301 , y16302 , y16303 , y16304 , y16305 , y16306 , y16307 , y16308 , y16309 , y16310 , y16311 , y16312 , y16313 , y16314 , y16315 , y16316 , y16317 , y16318 , y16319 , y16320 , y16321 , y16322 , y16323 , y16324 , y16325 , y16326 , y16327 , y16328 , y16329 , y16330 , y16331 , y16332 , y16333 , y16334 , y16335 , y16336 , y16337 , y16338 , y16339 , y16340 , y16341 , y16342 , y16343 , y16344 , y16345 , y16346 , y16347 , y16348 , y16349 , y16350 , y16351 , y16352 , y16353 , y16354 , y16355 , y16356 , y16357 , y16358 , y16359 , y16360 , y16361 , y16362 , y16363 , y16364 , y16365 , y16366 , y16367 , y16368 , y16369 , y16370 , y16371 , y16372 , y16373 , y16374 , y16375 , y16376 , y16377 , y16378 , y16379 , y16380 , y16381 , y16382 , y16383 , y16384 , y16385 , y16386 , y16387 , y16388 , y16389 , y16390 , y16391 , y16392 , y16393 , y16394 , y16395 , y16396 , y16397 , y16398 , y16399 , y16400 , y16401 , y16402 , y16403 , y16404 , y16405 , y16406 , y16407 , y16408 , y16409 , y16410 , y16411 , y16412 , y16413 , y16414 , y16415 , y16416 , y16417 , y16418 , y16419 , y16420 , y16421 , y16422 , y16423 , y16424 , y16425 , y16426 , y16427 , y16428 , y16429 , y16430 , y16431 , y16432 , y16433 , y16434 , y16435 , y16436 , y16437 , y16438 , y16439 , y16440 , y16441 , y16442 , y16443 , y16444 , y16445 , y16446 , y16447 , y16448 , y16449 , y16450 , y16451 , y16452 , y16453 , y16454 , y16455 , y16456 , y16457 , y16458 , y16459 , y16460 , y16461 , y16462 , y16463 , y16464 , y16465 , y16466 , y16467 , y16468 , y16469 , y16470 , y16471 , y16472 , y16473 , y16474 , y16475 , y16476 , y16477 , y16478 , y16479 , y16480 , y16481 , y16482 , y16483 , y16484 , y16485 , y16486 , y16487 , y16488 , y16489 , y16490 , y16491 , y16492 , y16493 , y16494 , y16495 , y16496 , y16497 , y16498 , y16499 , y16500 , y16501 , y16502 , y16503 , y16504 , y16505 , y16506 , y16507 , y16508 , y16509 , y16510 , y16511 , y16512 , y16513 , y16514 , y16515 , y16516 , y16517 , y16518 , y16519 , y16520 , y16521 , y16522 , y16523 , y16524 , y16525 , y16526 , y16527 , y16528 , y16529 , y16530 , y16531 , y16532 , y16533 , y16534 , y16535 , y16536 , y16537 , y16538 , y16539 , y16540 , y16541 , y16542 , y16543 , y16544 , y16545 , y16546 , y16547 , y16548 , y16549 , y16550 , y16551 , y16552 , y16553 , y16554 , y16555 , y16556 , y16557 , y16558 , y16559 , y16560 , y16561 , y16562 , y16563 , y16564 , y16565 , y16566 , y16567 , y16568 , y16569 , y16570 , y16571 , y16572 , y16573 , y16574 , y16575 , y16576 , y16577 , y16578 , y16579 , y16580 , y16581 , y16582 , y16583 , y16584 , y16585 , y16586 , y16587 , y16588 , y16589 , y16590 , y16591 , y16592 , y16593 , y16594 , y16595 , y16596 , y16597 , y16598 , y16599 , y16600 , y16601 , y16602 , y16603 , y16604 , y16605 , y16606 , y16607 , y16608 , y16609 , y16610 , y16611 , y16612 , y16613 , y16614 , y16615 , y16616 , y16617 , y16618 , y16619 , y16620 , y16621 , y16622 , y16623 , y16624 , y16625 , y16626 , y16627 , y16628 , y16629 , y16630 , y16631 , y16632 , y16633 , y16634 , y16635 , y16636 , y16637 , y16638 , y16639 , y16640 , y16641 , y16642 , y16643 , y16644 , y16645 , y16646 , y16647 , y16648 , y16649 , y16650 , y16651 , y16652 , y16653 , y16654 , y16655 , y16656 , y16657 , y16658 , y16659 , y16660 , y16661 , y16662 , y16663 , y16664 , y16665 , y16666 , y16667 , y16668 , y16669 , y16670 , y16671 , y16672 , y16673 , y16674 , y16675 , y16676 , y16677 , y16678 , y16679 , y16680 , y16681 , y16682 , y16683 , y16684 , y16685 , y16686 , y16687 , y16688 , y16689 , y16690 , y16691 , y16692 , y16693 , y16694 , y16695 , y16696 , y16697 , y16698 , y16699 , y16700 , y16701 , y16702 , y16703 , y16704 , y16705 , y16706 , y16707 , y16708 , y16709 , y16710 , y16711 , y16712 , y16713 , y16714 , y16715 , y16716 , y16717 , y16718 , y16719 , y16720 , y16721 , y16722 , y16723 , y16724 , y16725 , y16726 , y16727 , y16728 , y16729 , y16730 , y16731 , y16732 , y16733 , y16734 , y16735 , y16736 , y16737 , y16738 , y16739 , y16740 , y16741 , y16742 , y16743 , y16744 , y16745 , y16746 , y16747 , y16748 , y16749 , y16750 , y16751 , y16752 , y16753 , y16754 , y16755 , y16756 , y16757 , y16758 , y16759 , y16760 , y16761 , y16762 , y16763 , y16764 , y16765 , y16766 , y16767 , y16768 , y16769 , y16770 , y16771 , y16772 , y16773 , y16774 , y16775 , y16776 , y16777 , y16778 , y16779 , y16780 , y16781 , y16782 , y16783 , y16784 , y16785 , y16786 , y16787 , y16788 , y16789 , y16790 , y16791 , y16792 , y16793 , y16794 , y16795 , y16796 , y16797 , y16798 , y16799 , y16800 , y16801 , y16802 , y16803 , y16804 , y16805 , y16806 , y16807 , y16808 , y16809 , y16810 , y16811 , y16812 , y16813 , y16814 , y16815 , y16816 , y16817 , y16818 , y16819 , y16820 , y16821 , y16822 , y16823 , y16824 , y16825 , y16826 , y16827 , y16828 , y16829 , y16830 , y16831 , y16832 , y16833 , y16834 , y16835 , y16836 , y16837 , y16838 , y16839 , y16840 , y16841 , y16842 , y16843 , y16844 , y16845 , y16846 , y16847 , y16848 , y16849 , y16850 , y16851 , y16852 , y16853 , y16854 , y16855 , y16856 , y16857 , y16858 , y16859 , y16860 , y16861 , y16862 , y16863 , y16864 , y16865 , y16866 , y16867 , y16868 , y16869 , y16870 , y16871 , y16872 , y16873 , y16874 , y16875 , y16876 , y16877 , y16878 , y16879 , y16880 , y16881 , y16882 , y16883 , y16884 , y16885 , y16886 , y16887 , y16888 , y16889 , y16890 , y16891 , y16892 , y16893 , y16894 , y16895 , y16896 , y16897 , y16898 , y16899 , y16900 , y16901 , y16902 , y16903 , y16904 , y16905 , y16906 , y16907 , y16908 , y16909 , y16910 , y16911 , y16912 , y16913 , y16914 , y16915 , y16916 , y16917 , y16918 , y16919 , y16920 , y16921 , y16922 , y16923 , y16924 , y16925 , y16926 , y16927 , y16928 , y16929 , y16930 , y16931 , y16932 , y16933 , y16934 , y16935 , y16936 , y16937 , y16938 , y16939 , y16940 , y16941 , y16942 , y16943 , y16944 , y16945 , y16946 , y16947 , y16948 , y16949 , y16950 , y16951 , y16952 , y16953 , y16954 , y16955 , y16956 , y16957 , y16958 , y16959 , y16960 , y16961 , y16962 , y16963 , y16964 , y16965 , y16966 , y16967 , y16968 , y16969 , y16970 , y16971 , y16972 , y16973 , y16974 , y16975 , y16976 , y16977 , y16978 , y16979 , y16980 , y16981 , y16982 , y16983 , y16984 , y16985 , y16986 , y16987 , y16988 , y16989 , y16990 , y16991 , y16992 , y16993 , y16994 , y16995 , y16996 , y16997 , y16998 , y16999 , y17000 , y17001 , y17002 , y17003 , y17004 , y17005 , y17006 , y17007 , y17008 , y17009 , y17010 , y17011 , y17012 , y17013 , y17014 , y17015 , y17016 , y17017 , y17018 , y17019 , y17020 , y17021 , y17022 , y17023 , y17024 , y17025 , y17026 , y17027 , y17028 , y17029 , y17030 , y17031 , y17032 , y17033 , y17034 , y17035 , y17036 , y17037 , y17038 , y17039 , y17040 , y17041 , y17042 , y17043 , y17044 , y17045 , y17046 , y17047 , y17048 , y17049 , y17050 , y17051 , y17052 , y17053 , y17054 , y17055 , y17056 , y17057 , y17058 , y17059 , y17060 , y17061 , y17062 , y17063 , y17064 , y17065 , y17066 , y17067 , y17068 , y17069 , y17070 , y17071 , y17072 , y17073 , y17074 , y17075 , y17076 , y17077 , y17078 , y17079 , y17080 , y17081 , y17082 , y17083 , y17084 , y17085 , y17086 , y17087 , y17088 , y17089 , y17090 , y17091 , y17092 , y17093 , y17094 , y17095 , y17096 , y17097 , y17098 , y17099 , y17100 , y17101 , y17102 , y17103 , y17104 , y17105 , y17106 , y17107 , y17108 , y17109 , y17110 , y17111 , y17112 , y17113 , y17114 , y17115 , y17116 , y17117 , y17118 , y17119 , y17120 , y17121 , y17122 , y17123 , y17124 , y17125 , y17126 , y17127 , y17128 , y17129 , y17130 , y17131 , y17132 , y17133 , y17134 , y17135 , y17136 , y17137 , y17138 , y17139 , y17140 , y17141 , y17142 , y17143 , y17144 , y17145 , y17146 , y17147 , y17148 , y17149 , y17150 , y17151 , y17152 , y17153 , y17154 , y17155 , y17156 , y17157 , y17158 , y17159 , y17160 , y17161 , y17162 , y17163 , y17164 , y17165 , y17166 , y17167 , y17168 , y17169 , y17170 , y17171 , y17172 , y17173 , y17174 , y17175 , y17176 , y17177 , y17178 , y17179 , y17180 , y17181 , y17182 , y17183 , y17184 , y17185 , y17186 , y17187 , y17188 , y17189 , y17190 , y17191 , y17192 , y17193 , y17194 , y17195 , y17196 , y17197 , y17198 , y17199 , y17200 , y17201 , y17202 , y17203 , y17204 , y17205 , y17206 , y17207 , y17208 , y17209 , y17210 , y17211 , y17212 , y17213 , y17214 , y17215 , y17216 , y17217 , y17218 , y17219 , y17220 , y17221 , y17222 , y17223 , y17224 , y17225 , y17226 , y17227 , y17228 , y17229 , y17230 , y17231 , y17232 , y17233 , y17234 , y17235 , y17236 , y17237 , y17238 , y17239 , y17240 , y17241 , y17242 , y17243 , y17244 , y17245 , y17246 , y17247 , y17248 , y17249 , y17250 , y17251 , y17252 , y17253 , y17254 , y17255 , y17256 , y17257 , y17258 , y17259 , y17260 , y17261 , y17262 , y17263 , y17264 , y17265 , y17266 , y17267 , y17268 , y17269 , y17270 , y17271 , y17272 , y17273 , y17274 , y17275 , y17276 , y17277 , y17278 , y17279 , y17280 , y17281 , y17282 , y17283 , y17284 , y17285 , y17286 , y17287 , y17288 , y17289 , y17290 , y17291 , y17292 , y17293 , y17294 , y17295 , y17296 , y17297 , y17298 , y17299 , y17300 , y17301 , y17302 , y17303 , y17304 , y17305 , y17306 , y17307 , y17308 , y17309 , y17310 , y17311 , y17312 , y17313 , y17314 , y17315 , y17316 , y17317 , y17318 , y17319 , y17320 , y17321 , y17322 , y17323 , y17324 , y17325 , y17326 , y17327 , y17328 , y17329 , y17330 , y17331 , y17332 , y17333 , y17334 , y17335 , y17336 , y17337 , y17338 , y17339 , y17340 , y17341 , y17342 , y17343 , y17344 , y17345 , y17346 , y17347 , y17348 , y17349 , y17350 , y17351 , y17352 , y17353 , y17354 , y17355 , y17356 , y17357 , y17358 , y17359 , y17360 , y17361 , y17362 , y17363 , y17364 , y17365 , y17366 , y17367 , y17368 , y17369 , y17370 , y17371 , y17372 , y17373 , y17374 , y17375 , y17376 , y17377 , y17378 , y17379 , y17380 , y17381 , y17382 , y17383 , y17384 , y17385 , y17386 , y17387 , y17388 , y17389 , y17390 , y17391 , y17392 , y17393 , y17394 , y17395 , y17396 , y17397 , y17398 , y17399 , y17400 , y17401 , y17402 , y17403 , y17404 , y17405 , y17406 , y17407 , y17408 , y17409 , y17410 , y17411 , y17412 , y17413 , y17414 , y17415 , y17416 , y17417 , y17418 , y17419 , y17420 , y17421 , y17422 , y17423 , y17424 , y17425 , y17426 , y17427 , y17428 , y17429 , y17430 , y17431 , y17432 , y17433 , y17434 , y17435 , y17436 , y17437 , y17438 , y17439 , y17440 , y17441 , y17442 , y17443 , y17444 , y17445 , y17446 , y17447 , y17448 , y17449 , y17450 , y17451 , y17452 , y17453 , y17454 , y17455 , y17456 , y17457 , y17458 , y17459 , y17460 , y17461 , y17462 , y17463 , y17464 , y17465 , y17466 , y17467 , y17468 , y17469 , y17470 , y17471 , y17472 , y17473 , y17474 , y17475 , y17476 , y17477 , y17478 , y17479 , y17480 , y17481 , y17482 , y17483 , y17484 , y17485 , y17486 , y17487 , y17488 , y17489 , y17490 , y17491 , y17492 , y17493 , y17494 , y17495 , y17496 , y17497 , y17498 , y17499 , y17500 , y17501 , y17502 , y17503 , y17504 , y17505 , y17506 , y17507 , y17508 , y17509 , y17510 , y17511 , y17512 , y17513 , y17514 , y17515 , y17516 , y17517 , y17518 , y17519 , y17520 , y17521 , y17522 , y17523 , y17524 , y17525 , y17526 , y17527 , y17528 , y17529 , y17530 , y17531 , y17532 , y17533 , y17534 , y17535 , y17536 , y17537 , y17538 , y17539 , y17540 , y17541 , y17542 , y17543 , y17544 , y17545 , y17546 , y17547 , y17548 , y17549 , y17550 , y17551 , y17552 , y17553 , y17554 , y17555 , y17556 , y17557 , y17558 , y17559 , y17560 , y17561 , y17562 , y17563 , y17564 , y17565 , y17566 , y17567 , y17568 , y17569 , y17570 , y17571 , y17572 , y17573 , y17574 , y17575 , y17576 , y17577 , y17578 , y17579 , y17580 , y17581 , y17582 , y17583 , y17584 , y17585 , y17586 , y17587 , y17588 , y17589 , y17590 , y17591 , y17592 , y17593 , y17594 , y17595 , y17596 , y17597 , y17598 , y17599 , y17600 , y17601 , y17602 , y17603 , y17604 , y17605 , y17606 , y17607 , y17608 , y17609 , y17610 , y17611 , y17612 , y17613 , y17614 , y17615 , y17616 , y17617 , y17618 , y17619 , y17620 , y17621 , y17622 , y17623 , y17624 , y17625 , y17626 , y17627 , y17628 , y17629 , y17630 , y17631 , y17632 , y17633 , y17634 , y17635 , y17636 , y17637 , y17638 , y17639 , y17640 , y17641 , y17642 , y17643 , y17644 , y17645 , y17646 , y17647 , y17648 , y17649 , y17650 , y17651 , y17652 , y17653 , y17654 , y17655 , y17656 , y17657 , y17658 , y17659 , y17660 , y17661 , y17662 , y17663 , y17664 , y17665 , y17666 , y17667 , y17668 , y17669 , y17670 , y17671 , y17672 , y17673 , y17674 , y17675 , y17676 , y17677 , y17678 , y17679 , y17680 , y17681 , y17682 , y17683 , y17684 , y17685 , y17686 , y17687 , y17688 , y17689 , y17690 , y17691 , y17692 , y17693 , y17694 , y17695 , y17696 , y17697 , y17698 , y17699 , y17700 , y17701 , y17702 , y17703 , y17704 , y17705 , y17706 , y17707 , y17708 , y17709 , y17710 , y17711 , y17712 , y17713 , y17714 , y17715 , y17716 , y17717 , y17718 , y17719 , y17720 , y17721 , y17722 , y17723 , y17724 , y17725 , y17726 , y17727 , y17728 , y17729 , y17730 , y17731 , y17732 , y17733 , y17734 , y17735 , y17736 , y17737 , y17738 , y17739 , y17740 , y17741 , y17742 , y17743 , y17744 , y17745 , y17746 , y17747 , y17748 , y17749 , y17750 , y17751 , y17752 , y17753 , y17754 , y17755 , y17756 , y17757 , y17758 , y17759 , y17760 , y17761 , y17762 , y17763 , y17764 , y17765 , y17766 , y17767 , y17768 , y17769 , y17770 , y17771 , y17772 , y17773 , y17774 , y17775 , y17776 , y17777 , y17778 , y17779 , y17780 , y17781 , y17782 , y17783 , y17784 , y17785 , y17786 , y17787 , y17788 , y17789 , y17790 , y17791 , y17792 , y17793 , y17794 , y17795 , y17796 , y17797 , y17798 , y17799 , y17800 , y17801 , y17802 , y17803 , y17804 , y17805 , y17806 , y17807 , y17808 , y17809 , y17810 , y17811 , y17812 , y17813 , y17814 , y17815 , y17816 , y17817 , y17818 , y17819 , y17820 , y17821 , y17822 , y17823 , y17824 , y17825 , y17826 , y17827 , y17828 , y17829 , y17830 , y17831 , y17832 , y17833 , y17834 , y17835 , y17836 , y17837 , y17838 , y17839 , y17840 , y17841 , y17842 , y17843 , y17844 , y17845 , y17846 , y17847 , y17848 , y17849 , y17850 , y17851 , y17852 , y17853 , y17854 , y17855 , y17856 , y17857 , y17858 , y17859 , y17860 , y17861 , y17862 , y17863 , y17864 , y17865 , y17866 , y17867 , y17868 , y17869 , y17870 , y17871 , y17872 , y17873 , y17874 , y17875 , y17876 , y17877 , y17878 , y17879 , y17880 , y17881 , y17882 , y17883 , y17884 , y17885 , y17886 , y17887 , y17888 , y17889 , y17890 , y17891 , y17892 , y17893 , y17894 , y17895 , y17896 , y17897 , y17898 , y17899 , y17900 , y17901 , y17902 , y17903 , y17904 , y17905 , y17906 , y17907 , y17908 , y17909 , y17910 , y17911 , y17912 , y17913 , y17914 , y17915 , y17916 , y17917 , y17918 , y17919 , y17920 , y17921 , y17922 , y17923 , y17924 , y17925 , y17926 , y17927 , y17928 , y17929 , y17930 , y17931 , y17932 , y17933 , y17934 , y17935 , y17936 , y17937 , y17938 , y17939 , y17940 , y17941 , y17942 , y17943 , y17944 , y17945 , y17946 , y17947 , y17948 , y17949 , y17950 , y17951 , y17952 , y17953 , y17954 , y17955 , y17956 , y17957 , y17958 , y17959 , y17960 , y17961 , y17962 , y17963 , y17964 , y17965 , y17966 , y17967 , y17968 , y17969 , y17970 , y17971 , y17972 , y17973 , y17974 , y17975 , y17976 , y17977 , y17978 , y17979 , y17980 , y17981 , y17982 , y17983 , y17984 , y17985 , y17986 , y17987 , y17988 , y17989 , y17990 , y17991 , y17992 , y17993 , y17994 , y17995 , y17996 , y17997 , y17998 , y17999 , y18000 , y18001 , y18002 , y18003 , y18004 , y18005 , y18006 , y18007 , y18008 , y18009 , y18010 , y18011 , y18012 , y18013 , y18014 , y18015 , y18016 , y18017 , y18018 , y18019 , y18020 , y18021 , y18022 , y18023 , y18024 , y18025 , y18026 , y18027 , y18028 , y18029 , y18030 , y18031 , y18032 , y18033 , y18034 , y18035 , y18036 , y18037 , y18038 , y18039 , y18040 , y18041 , y18042 , y18043 , y18044 , y18045 , y18046 , y18047 , y18048 , y18049 , y18050 , y18051 , y18052 , y18053 , y18054 , y18055 , y18056 , y18057 , y18058 , y18059 , y18060 , y18061 , y18062 , y18063 , y18064 , y18065 , y18066 , y18067 , y18068 , y18069 , y18070 , y18071 , y18072 , y18073 , y18074 , y18075 , y18076 , y18077 , y18078 , y18079 , y18080 , y18081 , y18082 , y18083 , y18084 , y18085 , y18086 , y18087 , y18088 , y18089 , y18090 , y18091 , y18092 , y18093 , y18094 , y18095 , y18096 , y18097 , y18098 , y18099 , y18100 , y18101 , y18102 , y18103 , y18104 , y18105 , y18106 , y18107 , y18108 , y18109 , y18110 , y18111 , y18112 , y18113 , y18114 , y18115 , y18116 , y18117 , y18118 , y18119 , y18120 , y18121 , y18122 , y18123 , y18124 , y18125 , y18126 , y18127 , y18128 , y18129 , y18130 , y18131 , y18132 , y18133 , y18134 , y18135 , y18136 , y18137 , y18138 , y18139 , y18140 , y18141 , y18142 , y18143 , y18144 , y18145 , y18146 , y18147 , y18148 , y18149 , y18150 , y18151 , y18152 , y18153 , y18154 , y18155 , y18156 , y18157 , y18158 , y18159 , y18160 , y18161 , y18162 , y18163 , y18164 , y18165 , y18166 , y18167 , y18168 , y18169 , y18170 , y18171 , y18172 , y18173 , y18174 , y18175 , y18176 , y18177 , y18178 , y18179 , y18180 , y18181 , y18182 , y18183 , y18184 , y18185 , y18186 , y18187 , y18188 , y18189 , y18190 , y18191 , y18192 , y18193 , y18194 , y18195 , y18196 , y18197 , y18198 , y18199 , y18200 , y18201 , y18202 , y18203 , y18204 , y18205 , y18206 , y18207 , y18208 , y18209 , y18210 , y18211 , y18212 , y18213 , y18214 , y18215 , y18216 , y18217 , y18218 , y18219 , y18220 , y18221 , y18222 , y18223 , y18224 , y18225 , y18226 , y18227 , y18228 , y18229 , y18230 , y18231 , y18232 , y18233 , y18234 , y18235 , y18236 , y18237 , y18238 , y18239 , y18240 , y18241 , y18242 , y18243 , y18244 , y18245 , y18246 , y18247 , y18248 , y18249 , y18250 , y18251 , y18252 , y18253 , y18254 , y18255 , y18256 , y18257 , y18258 , y18259 , y18260 , y18261 , y18262 , y18263 , y18264 , y18265 , y18266 , y18267 , y18268 , y18269 , y18270 , y18271 , y18272 , y18273 , y18274 , y18275 , y18276 , y18277 , y18278 , y18279 , y18280 , y18281 , y18282 , y18283 , y18284 , y18285 , y18286 , y18287 , y18288 , y18289 , y18290 , y18291 , y18292 , y18293 , y18294 , y18295 , y18296 , y18297 , y18298 , y18299 , y18300 , y18301 , y18302 , y18303 , y18304 , y18305 , y18306 , y18307 , y18308 , y18309 , y18310 , y18311 , y18312 , y18313 , y18314 , y18315 , y18316 , y18317 , y18318 , y18319 , y18320 , y18321 , y18322 , y18323 , y18324 , y18325 , y18326 , y18327 , y18328 , y18329 , y18330 , y18331 , y18332 , y18333 , y18334 , y18335 , y18336 , y18337 , y18338 , y18339 , y18340 , y18341 , y18342 , y18343 , y18344 , y18345 , y18346 , y18347 , y18348 , y18349 , y18350 , y18351 , y18352 , y18353 , y18354 , y18355 , y18356 , y18357 , y18358 , y18359 , y18360 , y18361 , y18362 , y18363 , y18364 , y18365 , y18366 , y18367 , y18368 , y18369 , y18370 , y18371 , y18372 , y18373 , y18374 , y18375 , y18376 , y18377 , y18378 , y18379 , y18380 , y18381 , y18382 , y18383 , y18384 , y18385 , y18386 , y18387 , y18388 , y18389 , y18390 , y18391 , y18392 , y18393 , y18394 , y18395 , y18396 , y18397 , y18398 , y18399 , y18400 , y18401 , y18402 , y18403 , y18404 , y18405 , y18406 , y18407 , y18408 , y18409 , y18410 , y18411 , y18412 , y18413 , y18414 , y18415 , y18416 , y18417 , y18418 , y18419 , y18420 , y18421 , y18422 , y18423 , y18424 , y18425 , y18426 , y18427 , y18428 , y18429 , y18430 , y18431 , y18432 , y18433 , y18434 , y18435 , y18436 , y18437 , y18438 , y18439 , y18440 , y18441 , y18442 , y18443 , y18444 , y18445 , y18446 , y18447 , y18448 , y18449 , y18450 , y18451 , y18452 , y18453 , y18454 , y18455 , y18456 , y18457 , y18458 , y18459 , y18460 , y18461 , y18462 , y18463 , y18464 , y18465 , y18466 , y18467 , y18468 , y18469 , y18470 , y18471 , y18472 , y18473 , y18474 , y18475 , y18476 , y18477 , y18478 , y18479 , y18480 , y18481 , y18482 , y18483 , y18484 , y18485 , y18486 , y18487 , y18488 , y18489 , y18490 , y18491 , y18492 , y18493 , y18494 , y18495 , y18496 , y18497 , y18498 , y18499 , y18500 , y18501 , y18502 , y18503 , y18504 , y18505 , y18506 , y18507 , y18508 , y18509 , y18510 , y18511 , y18512 , y18513 , y18514 , y18515 , y18516 , y18517 , y18518 , y18519 , y18520 , y18521 , y18522 , y18523 , y18524 , y18525 , y18526 , y18527 , y18528 , y18529 , y18530 , y18531 , y18532 , y18533 , y18534 , y18535 , y18536 , y18537 , y18538 , y18539 , y18540 , y18541 , y18542 , y18543 , y18544 , y18545 , y18546 , y18547 , y18548 , y18549 , y18550 , y18551 , y18552 , y18553 , y18554 , y18555 , y18556 , y18557 , y18558 , y18559 , y18560 , y18561 , y18562 , y18563 , y18564 , y18565 , y18566 , y18567 , y18568 , y18569 , y18570 , y18571 , y18572 , y18573 , y18574 , y18575 , y18576 , y18577 , y18578 , y18579 , y18580 , y18581 , y18582 , y18583 , y18584 , y18585 , y18586 , y18587 , y18588 , y18589 , y18590 , y18591 , y18592 , y18593 , y18594 , y18595 , y18596 , y18597 , y18598 , y18599 , y18600 , y18601 , y18602 , y18603 , y18604 , y18605 , y18606 , y18607 , y18608 , y18609 , y18610 , y18611 , y18612 , y18613 , y18614 , y18615 , y18616 , y18617 , y18618 , y18619 , y18620 , y18621 , y18622 , y18623 , y18624 , y18625 , y18626 , y18627 , y18628 , y18629 , y18630 , y18631 , y18632 , y18633 , y18634 , y18635 , y18636 , y18637 , y18638 , y18639 , y18640 , y18641 , y18642 , y18643 , y18644 , y18645 , y18646 , y18647 , y18648 , y18649 , y18650 , y18651 , y18652 , y18653 , y18654 , y18655 , y18656 , y18657 , y18658 , y18659 , y18660 , y18661 , y18662 , y18663 , y18664 , y18665 , y18666 , y18667 , y18668 , y18669 , y18670 , y18671 , y18672 , y18673 , y18674 , y18675 , y18676 , y18677 , y18678 , y18679 , y18680 , y18681 , y18682 , y18683 , y18684 , y18685 , y18686 , y18687 , y18688 , y18689 , y18690 , y18691 , y18692 , y18693 , y18694 , y18695 , y18696 , y18697 , y18698 , y18699 , y18700 , y18701 , y18702 , y18703 , y18704 , y18705 , y18706 , y18707 , y18708 , y18709 , y18710 , y18711 , y18712 , y18713 , y18714 , y18715 , y18716 , y18717 , y18718 , y18719 , y18720 , y18721 , y18722 , y18723 , y18724 , y18725 , y18726 , y18727 , y18728 , y18729 , y18730 , y18731 , y18732 , y18733 , y18734 , y18735 , y18736 , y18737 , y18738 , y18739 , y18740 , y18741 , y18742 , y18743 , y18744 , y18745 , y18746 , y18747 , y18748 , y18749 , y18750 , y18751 , y18752 , y18753 , y18754 , y18755 , y18756 , y18757 , y18758 , y18759 , y18760 , y18761 , y18762 , y18763 , y18764 , y18765 , y18766 , y18767 , y18768 , y18769 , y18770 , y18771 , y18772 , y18773 , y18774 , y18775 , y18776 , y18777 , y18778 , y18779 , y18780 , y18781 , y18782 , y18783 , y18784 , y18785 , y18786 , y18787 , y18788 , y18789 , y18790 , y18791 , y18792 , y18793 , y18794 , y18795 , y18796 , y18797 , y18798 , y18799 , y18800 , y18801 , y18802 , y18803 , y18804 , y18805 , y18806 , y18807 , y18808 , y18809 , y18810 , y18811 , y18812 , y18813 , y18814 , y18815 , y18816 , y18817 , y18818 , y18819 , y18820 , y18821 , y18822 , y18823 , y18824 , y18825 , y18826 , y18827 , y18828 , y18829 , y18830 , y18831 , y18832 , y18833 , y18834 , y18835 , y18836 , y18837 , y18838 , y18839 , y18840 , y18841 , y18842 , y18843 , y18844 , y18845 , y18846 , y18847 , y18848 , y18849 , y18850 , y18851 , y18852 , y18853 , y18854 , y18855 , y18856 , y18857 , y18858 , y18859 , y18860 , y18861 , y18862 , y18863 , y18864 , y18865 , y18866 , y18867 , y18868 , y18869 , y18870 , y18871 , y18872 , y18873 , y18874 , y18875 , y18876 , y18877 , y18878 , y18879 , y18880 , y18881 , y18882 , y18883 , y18884 , y18885 , y18886 , y18887 , y18888 , y18889 , y18890 , y18891 , y18892 , y18893 , y18894 , y18895 , y18896 , y18897 , y18898 , y18899 , y18900 , y18901 , y18902 , y18903 , y18904 , y18905 , y18906 , y18907 , y18908 , y18909 , y18910 , y18911 , y18912 , y18913 , y18914 , y18915 , y18916 , y18917 , y18918 , y18919 , y18920 , y18921 , y18922 , y18923 , y18924 , y18925 , y18926 , y18927 , y18928 , y18929 , y18930 , y18931 , y18932 , y18933 , y18934 , y18935 , y18936 , y18937 , y18938 , y18939 , y18940 , y18941 , y18942 , y18943 , y18944 , y18945 , y18946 , y18947 , y18948 , y18949 , y18950 , y18951 , y18952 , y18953 , y18954 , y18955 , y18956 , y18957 , y18958 , y18959 , y18960 , y18961 , y18962 , y18963 , y18964 , y18965 , y18966 , y18967 , y18968 , y18969 , y18970 , y18971 , y18972 , y18973 , y18974 , y18975 , y18976 , y18977 , y18978 , y18979 , y18980 , y18981 , y18982 , y18983 , y18984 , y18985 , y18986 , y18987 , y18988 , y18989 , y18990 , y18991 , y18992 , y18993 , y18994 , y18995 , y18996 , y18997 , y18998 , y18999 , y19000 , y19001 , y19002 , y19003 , y19004 , y19005 , y19006 , y19007 , y19008 , y19009 , y19010 , y19011 , y19012 , y19013 , y19014 , y19015 , y19016 , y19017 , y19018 , y19019 , y19020 , y19021 , y19022 , y19023 , y19024 , y19025 , y19026 , y19027 , y19028 , y19029 , y19030 , y19031 , y19032 , y19033 , y19034 , y19035 , y19036 , y19037 , y19038 , y19039 , y19040 , y19041 , y19042 , y19043 , y19044 , y19045 , y19046 , y19047 , y19048 , y19049 , y19050 , y19051 , y19052 , y19053 , y19054 , y19055 , y19056 , y19057 , y19058 , y19059 , y19060 , y19061 , y19062 , y19063 , y19064 , y19065 , y19066 , y19067 , y19068 , y19069 , y19070 , y19071 , y19072 , y19073 , y19074 , y19075 , y19076 , y19077 , y19078 , y19079 , y19080 , y19081 , y19082 , y19083 , y19084 , y19085 , y19086 , y19087 , y19088 , y19089 , y19090 , y19091 , y19092 , y19093 , y19094 , y19095 , y19096 , y19097 , y19098 , y19099 , y19100 , y19101 , y19102 , y19103 , y19104 , y19105 , y19106 , y19107 , y19108 , y19109 , y19110 , y19111 , y19112 , y19113 , y19114 , y19115 , y19116 , y19117 , y19118 , y19119 , y19120 , y19121 , y19122 , y19123 , y19124 , y19125 , y19126 , y19127 , y19128 , y19129 , y19130 , y19131 , y19132 , y19133 , y19134 , y19135 , y19136 , y19137 , y19138 , y19139 , y19140 , y19141 , y19142 , y19143 , y19144 , y19145 , y19146 , y19147 , y19148 , y19149 , y19150 , y19151 , y19152 , y19153 , y19154 , y19155 , y19156 , y19157 , y19158 , y19159 , y19160 , y19161 , y19162 , y19163 , y19164 , y19165 , y19166 , y19167 , y19168 , y19169 , y19170 , y19171 , y19172 , y19173 , y19174 , y19175 , y19176 , y19177 , y19178 , y19179 , y19180 , y19181 , y19182 , y19183 , y19184 , y19185 , y19186 , y19187 , y19188 , y19189 , y19190 , y19191 , y19192 , y19193 , y19194 , y19195 , y19196 , y19197 , y19198 , y19199 , y19200 , y19201 , y19202 , y19203 , y19204 , y19205 , y19206 , y19207 , y19208 , y19209 , y19210 , y19211 , y19212 , y19213 , y19214 , y19215 , y19216 , y19217 , y19218 , y19219 , y19220 , y19221 , y19222 , y19223 , y19224 , y19225 , y19226 , y19227 , y19228 , y19229 , y19230 , y19231 , y19232 , y19233 , y19234 , y19235 , y19236 , y19237 , y19238 , y19239 , y19240 , y19241 , y19242 , y19243 , y19244 , y19245 , y19246 , y19247 , y19248 , y19249 , y19250 , y19251 , y19252 , y19253 , y19254 , y19255 , y19256 , y19257 , y19258 , y19259 , y19260 , y19261 , y19262 , y19263 , y19264 , y19265 , y19266 , y19267 , y19268 , y19269 , y19270 , y19271 , y19272 , y19273 , y19274 , y19275 , y19276 , y19277 , y19278 , y19279 , y19280 , y19281 , y19282 , y19283 , y19284 , y19285 , y19286 , y19287 , y19288 , y19289 , y19290 , y19291 , y19292 , y19293 , y19294 , y19295 , y19296 , y19297 , y19298 , y19299 , y19300 , y19301 , y19302 , y19303 , y19304 , y19305 , y19306 , y19307 , y19308 , y19309 , y19310 , y19311 , y19312 , y19313 , y19314 , y19315 , y19316 , y19317 , y19318 , y19319 , y19320 , y19321 , y19322 , y19323 , y19324 , y19325 , y19326 , y19327 , y19328 , y19329 , y19330 , y19331 , y19332 , y19333 , y19334 , y19335 , y19336 , y19337 , y19338 , y19339 , y19340 , y19341 , y19342 , y19343 , y19344 , y19345 , y19346 , y19347 , y19348 , y19349 , y19350 , y19351 , y19352 , y19353 , y19354 , y19355 , y19356 , y19357 , y19358 , y19359 , y19360 , y19361 , y19362 , y19363 , y19364 , y19365 , y19366 , y19367 , y19368 , y19369 , y19370 , y19371 , y19372 , y19373 , y19374 , y19375 , y19376 , y19377 , y19378 , y19379 , y19380 , y19381 , y19382 , y19383 , y19384 , y19385 , y19386 , y19387 , y19388 , y19389 , y19390 , y19391 , y19392 , y19393 , y19394 , y19395 , y19396 , y19397 , y19398 , y19399 , y19400 , y19401 , y19402 , y19403 , y19404 , y19405 , y19406 , y19407 , y19408 , y19409 , y19410 , y19411 , y19412 , y19413 , y19414 , y19415 , y19416 , y19417 , y19418 , y19419 , y19420 , y19421 , y19422 , y19423 , y19424 , y19425 , y19426 , y19427 , y19428 , y19429 , y19430 , y19431 , y19432 , y19433 , y19434 , y19435 , y19436 , y19437 , y19438 , y19439 , y19440 , y19441 , y19442 , y19443 , y19444 , y19445 , y19446 , y19447 , y19448 , y19449 , y19450 , y19451 , y19452 , y19453 , y19454 , y19455 , y19456 , y19457 , y19458 , y19459 , y19460 , y19461 , y19462 , y19463 , y19464 , y19465 , y19466 , y19467 , y19468 , y19469 , y19470 , y19471 , y19472 , y19473 , y19474 , y19475 , y19476 , y19477 , y19478 , y19479 , y19480 , y19481 , y19482 , y19483 , y19484 , y19485 , y19486 , y19487 , y19488 , y19489 , y19490 , y19491 , y19492 , y19493 , y19494 , y19495 , y19496 , y19497 , y19498 , y19499 , y19500 , y19501 , y19502 , y19503 , y19504 , y19505 , y19506 , y19507 , y19508 , y19509 , y19510 , y19511 , y19512 , y19513 , y19514 , y19515 , y19516 , y19517 , y19518 , y19519 , y19520 , y19521 , y19522 , y19523 , y19524 , y19525 , y19526 , y19527 , y19528 , y19529 , y19530 , y19531 , y19532 , y19533 , y19534 , y19535 , y19536 , y19537 , y19538 , y19539 , y19540 , y19541 , y19542 , y19543 , y19544 , y19545 , y19546 , y19547 , y19548 , y19549 , y19550 , y19551 , y19552 , y19553 , y19554 , y19555 , y19556 , y19557 , y19558 , y19559 , y19560 , y19561 , y19562 , y19563 , y19564 , y19565 , y19566 , y19567 , y19568 , y19569 , y19570 , y19571 , y19572 , y19573 , y19574 , y19575 , y19576 , y19577 , y19578 , y19579 , y19580 , y19581 , y19582 , y19583 , y19584 , y19585 , y19586 , y19587 , y19588 , y19589 , y19590 , y19591 , y19592 , y19593 , y19594 , y19595 , y19596 , y19597 , y19598 , y19599 , y19600 , y19601 , y19602 , y19603 , y19604 , y19605 , y19606 , y19607 , y19608 , y19609 , y19610 , y19611 , y19612 , y19613 , y19614 , y19615 , y19616 , y19617 , y19618 , y19619 , y19620 , y19621 , y19622 , y19623 , y19624 , y19625 , y19626 , y19627 , y19628 , y19629 , y19630 , y19631 , y19632 , y19633 , y19634 , y19635 , y19636 , y19637 , y19638 , y19639 , y19640 , y19641 , y19642 , y19643 , y19644 , y19645 , y19646 , y19647 , y19648 , y19649 , y19650 , y19651 , y19652 , y19653 , y19654 , y19655 , y19656 , y19657 , y19658 , y19659 , y19660 , y19661 , y19662 , y19663 , y19664 , y19665 , y19666 , y19667 , y19668 , y19669 , y19670 , y19671 , y19672 , y19673 , y19674 , y19675 , y19676 , y19677 , y19678 , y19679 , y19680 , y19681 , y19682 , y19683 , y19684 , y19685 , y19686 , y19687 , y19688 , y19689 , y19690 , y19691 , y19692 , y19693 , y19694 , y19695 , y19696 , y19697 , y19698 , y19699 , y19700 , y19701 , y19702 , y19703 , y19704 , y19705 , y19706 , y19707 , y19708 , y19709 , y19710 , y19711 , y19712 , y19713 , y19714 , y19715 , y19716 , y19717 , y19718 , y19719 , y19720 , y19721 , y19722 , y19723 , y19724 , y19725 , y19726 , y19727 , y19728 , y19729 , y19730 , y19731 , y19732 , y19733 , y19734 , y19735 , y19736 , y19737 , y19738 , y19739 , y19740 , y19741 , y19742 , y19743 , y19744 , y19745 , y19746 , y19747 , y19748 , y19749 , y19750 , y19751 , y19752 , y19753 , y19754 , y19755 , y19756 , y19757 , y19758 , y19759 , y19760 , y19761 , y19762 , y19763 , y19764 , y19765 , y19766 , y19767 , y19768 , y19769 , y19770 , y19771 , y19772 , y19773 , y19774 , y19775 , y19776 , y19777 , y19778 , y19779 , y19780 , y19781 , y19782 , y19783 , y19784 , y19785 , y19786 , y19787 , y19788 , y19789 , y19790 , y19791 , y19792 , y19793 , y19794 , y19795 , y19796 , y19797 , y19798 , y19799 , y19800 , y19801 , y19802 , y19803 , y19804 , y19805 , y19806 , y19807 , y19808 , y19809 , y19810 , y19811 , y19812 , y19813 , y19814 , y19815 , y19816 , y19817 , y19818 , y19819 , y19820 , y19821 , y19822 , y19823 , y19824 , y19825 , y19826 , y19827 , y19828 , y19829 , y19830 , y19831 , y19832 , y19833 , y19834 , y19835 , y19836 , y19837 , y19838 , y19839 , y19840 , y19841 , y19842 , y19843 , y19844 , y19845 , y19846 , y19847 , y19848 , y19849 , y19850 , y19851 , y19852 , y19853 , y19854 , y19855 , y19856 , y19857 , y19858 , y19859 , y19860 , y19861 , y19862 , y19863 , y19864 , y19865 , y19866 , y19867 , y19868 , y19869 , y19870 , y19871 , y19872 , y19873 , y19874 , y19875 , y19876 , y19877 , y19878 , y19879 , y19880 , y19881 , y19882 , y19883 , y19884 , y19885 , y19886 , y19887 , y19888 , y19889 , y19890 , y19891 , y19892 , y19893 , y19894 , y19895 , y19896 , y19897 , y19898 , y19899 , y19900 , y19901 , y19902 , y19903 , y19904 , y19905 , y19906 , y19907 , y19908 , y19909 , y19910 , y19911 , y19912 , y19913 , y19914 , y19915 , y19916 , y19917 , y19918 , y19919 , y19920 , y19921 , y19922 , y19923 , y19924 , y19925 , y19926 , y19927 , y19928 , y19929 , y19930 , y19931 , y19932 , y19933 , y19934 , y19935 , y19936 , y19937 , y19938 , y19939 , y19940 , y19941 , y19942 , y19943 , y19944 , y19945 , y19946 , y19947 , y19948 , y19949 , y19950 , y19951 , y19952 , y19953 , y19954 , y19955 , y19956 , y19957 , y19958 , y19959 , y19960 , y19961 , y19962 , y19963 , y19964 , y19965 , y19966 , y19967 , y19968 , y19969 , y19970 , y19971 , y19972 , y19973 , y19974 , y19975 , y19976 , y19977 , y19978 , y19979 , y19980 , y19981 , y19982 , y19983 , y19984 , y19985 , y19986 , y19987 , y19988 , y19989 , y19990 , y19991 , y19992 , y19993 , y19994 , y19995 , y19996 , y19997 , y19998 , y19999 , y20000 , y20001 , y20002 , y20003 , y20004 , y20005 , y20006 , y20007 , y20008 , y20009 , y20010 , y20011 , y20012 , y20013 , y20014 , y20015 , y20016 , y20017 , y20018 , y20019 , y20020 , y20021 , y20022 , y20023 , y20024 , y20025 , y20026 , y20027 , y20028 , y20029 , y20030 , y20031 , y20032 , y20033 , y20034 , y20035 , y20036 , y20037 , y20038 , y20039 , y20040 , y20041 , y20042 , y20043 , y20044 , y20045 , y20046 , y20047 , y20048 , y20049 , y20050 , y20051 , y20052 , y20053 , y20054 , y20055 , y20056 , y20057 , y20058 , y20059 , y20060 , y20061 , y20062 , y20063 , y20064 , y20065 , y20066 , y20067 , y20068 , y20069 , y20070 , y20071 , y20072 , y20073 , y20074 , y20075 , y20076 , y20077 , y20078 , y20079 , y20080 , y20081 , y20082 , y20083 , y20084 , y20085 , y20086 , y20087 , y20088 , y20089 , y20090 , y20091 , y20092 , y20093 , y20094 , y20095 , y20096 , y20097 , y20098 , y20099 , y20100 , y20101 , y20102 , y20103 , y20104 , y20105 , y20106 , y20107 , y20108 , y20109 , y20110 , y20111 , y20112 , y20113 , y20114 , y20115 , y20116 , y20117 , y20118 , y20119 , y20120 , y20121 , y20122 , y20123 , y20124 , y20125 , y20126 , y20127 , y20128 , y20129 , y20130 , y20131 , y20132 , y20133 , y20134 , y20135 , y20136 , y20137 , y20138 , y20139 , y20140 , y20141 , y20142 , y20143 , y20144 , y20145 , y20146 , y20147 , y20148 , y20149 , y20150 , y20151 , y20152 , y20153 , y20154 , y20155 , y20156 , y20157 , y20158 , y20159 , y20160 , y20161 , y20162 , y20163 , y20164 , y20165 , y20166 , y20167 , y20168 , y20169 , y20170 , y20171 , y20172 , y20173 , y20174 , y20175 , y20176 , y20177 , y20178 , y20179 , y20180 , y20181 , y20182 , y20183 , y20184 , y20185 , y20186 , y20187 , y20188 , y20189 , y20190 , y20191 , y20192 , y20193 , y20194 , y20195 , y20196 , y20197 , y20198 , y20199 , y20200 , y20201 , y20202 , y20203 , y20204 , y20205 , y20206 , y20207 , y20208 , y20209 , y20210 , y20211 , y20212 , y20213 , y20214 , y20215 , y20216 , y20217 , y20218 , y20219 , y20220 , y20221 , y20222 , y20223 , y20224 , y20225 , y20226 , y20227 , y20228 , y20229 , y20230 , y20231 , y20232 , y20233 , y20234 , y20235 , y20236 , y20237 , y20238 , y20239 , y20240 , y20241 , y20242 , y20243 , y20244 , y20245 , y20246 , y20247 , y20248 , y20249 , y20250 , y20251 , y20252 , y20253 , y20254 , y20255 , y20256 , y20257 , y20258 , y20259 , y20260 , y20261 , y20262 , y20263 , y20264 , y20265 , y20266 , y20267 , y20268 , y20269 , y20270 , y20271 , y20272 , y20273 , y20274 , y20275 , y20276 , y20277 , y20278 , y20279 , y20280 , y20281 , y20282 , y20283 , y20284 , y20285 , y20286 , y20287 , y20288 , y20289 , y20290 , y20291 , y20292 , y20293 , y20294 , y20295 , y20296 , y20297 , y20298 , y20299 , y20300 , y20301 , y20302 , y20303 , y20304 , y20305 , y20306 , y20307 , y20308 , y20309 , y20310 , y20311 , y20312 , y20313 , y20314 , y20315 , y20316 , y20317 , y20318 , y20319 , y20320 , y20321 , y20322 , y20323 , y20324 , y20325 , y20326 , y20327 , y20328 , y20329 , y20330 , y20331 , y20332 , y20333 , y20334 , y20335 , y20336 , y20337 , y20338 , y20339 , y20340 , y20341 , y20342 , y20343 , y20344 , y20345 , y20346 , y20347 , y20348 , y20349 , y20350 , y20351 , y20352 , y20353 , y20354 , y20355 , y20356 , y20357 , y20358 , y20359 , y20360 , y20361 , y20362 , y20363 , y20364 , y20365 , y20366 , y20367 , y20368 , y20369 , y20370 , y20371 , y20372 , y20373 , y20374 , y20375 , y20376 , y20377 , y20378 , y20379 , y20380 , y20381 , y20382 , y20383 , y20384 , y20385 , y20386 , y20387 , y20388 , y20389 , y20390 , y20391 , y20392 , y20393 , y20394 , y20395 , y20396 , y20397 , y20398 , y20399 , y20400 , y20401 , y20402 , y20403 , y20404 , y20405 , y20406 , y20407 , y20408 , y20409 , y20410 , y20411 , y20412 , y20413 , y20414 , y20415 , y20416 , y20417 , y20418 , y20419 , y20420 , y20421 , y20422 , y20423 , y20424 , y20425 , y20426 , y20427 , y20428 , y20429 , y20430 , y20431 , y20432 , y20433 , y20434 , y20435 , y20436 , y20437 , y20438 , y20439 , y20440 , y20441 , y20442 , y20443 , y20444 , y20445 , y20446 , y20447 , y20448 , y20449 , y20450 , y20451 , y20452 , y20453 , y20454 , y20455 , y20456 , y20457 , y20458 , y20459 , y20460 , y20461 , y20462 , y20463 , y20464 , y20465 , y20466 , y20467 , y20468 , y20469 , y20470 , y20471 , y20472 , y20473 , y20474 , y20475 , y20476 , y20477 , y20478 , y20479 , y20480 , y20481 , y20482 , y20483 , y20484 , y20485 , y20486 , y20487 , y20488 , y20489 , y20490 , y20491 , y20492 , y20493 , y20494 , y20495 , y20496 , y20497 , y20498 , y20499 , y20500 , y20501 , y20502 , y20503 , y20504 , y20505 , y20506 , y20507 , y20508 , y20509 , y20510 , y20511 , y20512 , y20513 , y20514 , y20515 , y20516 , y20517 , y20518 , y20519 , y20520 , y20521 , y20522 , y20523 , y20524 , y20525 , y20526 , y20527 , y20528 , y20529 , y20530 , y20531 , y20532 , y20533 , y20534 , y20535 , y20536 , y20537 , y20538 , y20539 , y20540 , y20541 , y20542 , y20543 , y20544 , y20545 , y20546 , y20547 , y20548 , y20549 , y20550 , y20551 , y20552 , y20553 , y20554 , y20555 , y20556 , y20557 , y20558 , y20559 , y20560 , y20561 , y20562 , y20563 , y20564 , y20565 , y20566 , y20567 , y20568 , y20569 , y20570 , y20571 , y20572 , y20573 , y20574 , y20575 , y20576 , y20577 , y20578 , y20579 , y20580 , y20581 , y20582 , y20583 , y20584 , y20585 , y20586 , y20587 , y20588 , y20589 , y20590 , y20591 , y20592 , y20593 , y20594 , y20595 , y20596 , y20597 , y20598 , y20599 , y20600 , y20601 , y20602 , y20603 , y20604 , y20605 , y20606 , y20607 , y20608 , y20609 , y20610 , y20611 , y20612 , y20613 , y20614 , y20615 , y20616 , y20617 , y20618 , y20619 , y20620 , y20621 , y20622 , y20623 , y20624 , y20625 , y20626 , y20627 , y20628 , y20629 , y20630 , y20631 , y20632 , y20633 , y20634 , y20635 , y20636 , y20637 , y20638 , y20639 , y20640 , y20641 , y20642 , y20643 , y20644 , y20645 , y20646 , y20647 , y20648 , y20649 , y20650 , y20651 , y20652 , y20653 , y20654 , y20655 , y20656 , y20657 , y20658 , y20659 , y20660 , y20661 , y20662 , y20663 , y20664 , y20665 , y20666 , y20667 , y20668 , y20669 , y20670 , y20671 , y20672 , y20673 , y20674 , y20675 , y20676 , y20677 , y20678 , y20679 , y20680 , y20681 , y20682 , y20683 , y20684 , y20685 , y20686 , y20687 , y20688 , y20689 , y20690 , y20691 , y20692 , y20693 , y20694 , y20695 , y20696 , y20697 , y20698 , y20699 , y20700 , y20701 , y20702 , y20703 , y20704 , y20705 , y20706 , y20707 , y20708 , y20709 , y20710 , y20711 , y20712 , y20713 , y20714 , y20715 , y20716 , y20717 , y20718 , y20719 , y20720 , y20721 , y20722 , y20723 , y20724 , y20725 , y20726 , y20727 , y20728 , y20729 , y20730 , y20731 , y20732 , y20733 , y20734 , y20735 , y20736 , y20737 , y20738 , y20739 , y20740 , y20741 , y20742 , y20743 , y20744 , y20745 , y20746 , y20747 , y20748 , y20749 , y20750 , y20751 , y20752 , y20753 , y20754 , y20755 , y20756 , y20757 , y20758 , y20759 , y20760 , y20761 , y20762 , y20763 , y20764 , y20765 , y20766 , y20767 , y20768 , y20769 , y20770 , y20771 , y20772 , y20773 , y20774 , y20775 , y20776 , y20777 , y20778 , y20779 , y20780 , y20781 , y20782 , y20783 , y20784 , y20785 , y20786 , y20787 , y20788 , y20789 , y20790 , y20791 , y20792 , y20793 , y20794 , y20795 , y20796 , y20797 , y20798 , y20799 , y20800 , y20801 , y20802 , y20803 , y20804 , y20805 , y20806 , y20807 , y20808 , y20809 , y20810 , y20811 , y20812 , y20813 , y20814 , y20815 , y20816 , y20817 , y20818 , y20819 , y20820 , y20821 , y20822 , y20823 , y20824 , y20825 , y20826 , y20827 , y20828 , y20829 , y20830 , y20831 , y20832 , y20833 , y20834 , y20835 , y20836 , y20837 , y20838 , y20839 , y20840 , y20841 , y20842 , y20843 , y20844 , y20845 , y20846 , y20847 , y20848 , y20849 , y20850 , y20851 , y20852 , y20853 , y20854 , y20855 , y20856 , y20857 , y20858 , y20859 , y20860 , y20861 , y20862 , y20863 , y20864 , y20865 , y20866 , y20867 , y20868 , y20869 , y20870 , y20871 , y20872 , y20873 , y20874 , y20875 , y20876 , y20877 , y20878 , y20879 , y20880 , y20881 , y20882 , y20883 , y20884 , y20885 , y20886 , y20887 , y20888 , y20889 , y20890 , y20891 , y20892 , y20893 , y20894 , y20895 , y20896 , y20897 , y20898 , y20899 , y20900 , y20901 , y20902 , y20903 , y20904 , y20905 , y20906 , y20907 , y20908 , y20909 , y20910 , y20911 , y20912 , y20913 , y20914 , y20915 , y20916 , y20917 , y20918 , y20919 , y20920 , y20921 , y20922 , y20923 , y20924 , y20925 , y20926 , y20927 , y20928 , y20929 , y20930 , y20931 , y20932 , y20933 , y20934 , y20935 , y20936 , y20937 , y20938 , y20939 , y20940 , y20941 , y20942 , y20943 , y20944 , y20945 , y20946 , y20947 , y20948 , y20949 , y20950 , y20951 , y20952 , y20953 , y20954 , y20955 , y20956 , y20957 , y20958 , y20959 , y20960 , y20961 , y20962 , y20963 , y20964 , y20965 , y20966 , y20967 , y20968 , y20969 , y20970 , y20971 , y20972 , y20973 , y20974 , y20975 , y20976 , y20977 , y20978 , y20979 , y20980 , y20981 , y20982 , y20983 , y20984 , y20985 , y20986 , y20987 , y20988 , y20989 , y20990 , y20991 , y20992 , y20993 , y20994 , y20995 , y20996 , y20997 , y20998 , y20999 , y21000 , y21001 , y21002 , y21003 , y21004 , y21005 , y21006 , y21007 , y21008 , y21009 , y21010 , y21011 , y21012 , y21013 , y21014 , y21015 , y21016 , y21017 , y21018 , y21019 , y21020 , y21021 , y21022 , y21023 , y21024 , y21025 , y21026 , y21027 , y21028 , y21029 , y21030 , y21031 , y21032 , y21033 , y21034 , y21035 , y21036 , y21037 , y21038 , y21039 , y21040 , y21041 , y21042 , y21043 , y21044 , y21045 , y21046 , y21047 , y21048 , y21049 , y21050 , y21051 , y21052 , y21053 , y21054 , y21055 , y21056 , y21057 , y21058 , y21059 , y21060 , y21061 , y21062 , y21063 , y21064 , y21065 , y21066 , y21067 , y21068 , y21069 , y21070 , y21071 , y21072 , y21073 , y21074 , y21075 , y21076 , y21077 , y21078 , y21079 , y21080 , y21081 , y21082 , y21083 , y21084 , y21085 , y21086 , y21087 , y21088 , y21089 , y21090 , y21091 , y21092 , y21093 , y21094 , y21095 , y21096 , y21097 , y21098 , y21099 , y21100 , y21101 , y21102 , y21103 , y21104 , y21105 , y21106 , y21107 , y21108 , y21109 , y21110 , y21111 , y21112 , y21113 , y21114 , y21115 , y21116 , y21117 , y21118 , y21119 , y21120 , y21121 , y21122 , y21123 , y21124 , y21125 , y21126 , y21127 , y21128 , y21129 , y21130 , y21131 , y21132 , y21133 , y21134 , y21135 , y21136 , y21137 , y21138 , y21139 , y21140 , y21141 , y21142 , y21143 , y21144 , y21145 , y21146 , y21147 , y21148 , y21149 , y21150 , y21151 , y21152 , y21153 , y21154 , y21155 , y21156 , y21157 , y21158 , y21159 , y21160 , y21161 , y21162 , y21163 , y21164 , y21165 , y21166 , y21167 , y21168 , y21169 , y21170 , y21171 , y21172 , y21173 , y21174 , y21175 , y21176 , y21177 , y21178 , y21179 , y21180 , y21181 , y21182 , y21183 , y21184 , y21185 , y21186 , y21187 , y21188 , y21189 , y21190 , y21191 , y21192 , y21193 , y21194 , y21195 , y21196 , y21197 , y21198 , y21199 , y21200 , y21201 , y21202 , y21203 , y21204 , y21205 , y21206 , y21207 , y21208 , y21209 , y21210 , y21211 , y21212 , y21213 , y21214 , y21215 , y21216 , y21217 , y21218 , y21219 , y21220 , y21221 , y21222 , y21223 , y21224 , y21225 , y21226 , y21227 , y21228 , y21229 , y21230 , y21231 , y21232 , y21233 , y21234 , y21235 , y21236 , y21237 , y21238 , y21239 , y21240 , y21241 , y21242 , y21243 , y21244 , y21245 , y21246 , y21247 , y21248 , y21249 , y21250 , y21251 , y21252 , y21253 , y21254 , y21255 , y21256 , y21257 , y21258 , y21259 , y21260 , y21261 , y21262 , y21263 , y21264 , y21265 , y21266 , y21267 , y21268 , y21269 , y21270 , y21271 , y21272 , y21273 , y21274 , y21275 , y21276 , y21277 , y21278 , y21279 , y21280 , y21281 , y21282 , y21283 , y21284 , y21285 , y21286 , y21287 , y21288 , y21289 , y21290 , y21291 , y21292 , y21293 , y21294 , y21295 , y21296 , y21297 , y21298 , y21299 , y21300 , y21301 , y21302 , y21303 , y21304 , y21305 , y21306 , y21307 , y21308 , y21309 , y21310 , y21311 , y21312 , y21313 , y21314 , y21315 , y21316 , y21317 , y21318 , y21319 , y21320 , y21321 , y21322 , y21323 , y21324 , y21325 , y21326 , y21327 , y21328 , y21329 , y21330 , y21331 , y21332 , y21333 , y21334 , y21335 , y21336 , y21337 , y21338 , y21339 , y21340 , y21341 , y21342 , y21343 , y21344 , y21345 , y21346 , y21347 , y21348 , y21349 , y21350 , y21351 , y21352 , y21353 , y21354 , y21355 , y21356 , y21357 , y21358 , y21359 , y21360 , y21361 , y21362 , y21363 , y21364 , y21365 , y21366 , y21367 , y21368 , y21369 , y21370 , y21371 , y21372 , y21373 , y21374 , y21375 , y21376 , y21377 , y21378 , y21379 , y21380 , y21381 , y21382 , y21383 , y21384 , y21385 , y21386 , y21387 , y21388 , y21389 , y21390 , y21391 , y21392 , y21393 , y21394 , y21395 , y21396 , y21397 , y21398 , y21399 , y21400 , y21401 , y21402 , y21403 , y21404 , y21405 , y21406 , y21407 , y21408 , y21409 , y21410 , y21411 , y21412 , y21413 , y21414 , y21415 , y21416 , y21417 , y21418 , y21419 , y21420 , y21421 , y21422 , y21423 , y21424 , y21425 , y21426 , y21427 , y21428 , y21429 , y21430 , y21431 , y21432 , y21433 , y21434 , y21435 , y21436 , y21437 , y21438 , y21439 , y21440 , y21441 , y21442 , y21443 , y21444 , y21445 , y21446 , y21447 , y21448 , y21449 , y21450 , y21451 , y21452 , y21453 , y21454 , y21455 , y21456 , y21457 , y21458 , y21459 , y21460 , y21461 , y21462 , y21463 , y21464 , y21465 , y21466 , y21467 , y21468 , y21469 , y21470 , y21471 , y21472 , y21473 , y21474 , y21475 , y21476 , y21477 , y21478 , y21479 , y21480 , y21481 , y21482 , y21483 , y21484 , y21485 , y21486 , y21487 , y21488 , y21489 , y21490 , y21491 , y21492 , y21493 , y21494 , y21495 , y21496 , y21497 , y21498 , y21499 , y21500 , y21501 , y21502 , y21503 , y21504 , y21505 , y21506 , y21507 , y21508 , y21509 , y21510 , y21511 , y21512 , y21513 , y21514 , y21515 , y21516 , y21517 , y21518 , y21519 , y21520 , y21521 , y21522 , y21523 , y21524 , y21525 , y21526 , y21527 , y21528 , y21529 , y21530 , y21531 , y21532 , y21533 , y21534 , y21535 , y21536 , y21537 , y21538 , y21539 , y21540 , y21541 , y21542 , y21543 , y21544 , y21545 , y21546 , y21547 , y21548 , y21549 , y21550 , y21551 , y21552 , y21553 , y21554 , y21555 , y21556 , y21557 , y21558 , y21559 , y21560 , y21561 , y21562 , y21563 , y21564 , y21565 , y21566 , y21567 , y21568 , y21569 , y21570 , y21571 , y21572 , y21573 , y21574 , y21575 , y21576 , y21577 , y21578 , y21579 , y21580 , y21581 , y21582 , y21583 , y21584 , y21585 , y21586 , y21587 , y21588 , y21589 , y21590 , y21591 , y21592 , y21593 , y21594 , y21595 , y21596 , y21597 , y21598 , y21599 , y21600 , y21601 , y21602 , y21603 , y21604 , y21605 , y21606 , y21607 , y21608 , y21609 , y21610 , y21611 , y21612 , y21613 , y21614 , y21615 , y21616 , y21617 , y21618 , y21619 , y21620 , y21621 , y21622 , y21623 , y21624 , y21625 , y21626 , y21627 , y21628 , y21629 , y21630 , y21631 , y21632 , y21633 , y21634 , y21635 , y21636 , y21637 , y21638 , y21639 , y21640 , y21641 , y21642 , y21643 , y21644 , y21645 , y21646 , y21647 , y21648 , y21649 , y21650 , y21651 , y21652 , y21653 , y21654 , y21655 , y21656 , y21657 , y21658 , y21659 , y21660 , y21661 , y21662 , y21663 , y21664 , y21665 , y21666 , y21667 , y21668 , y21669 , y21670 , y21671 , y21672 , y21673 , y21674 , y21675 , y21676 , y21677 , y21678 , y21679 , y21680 , y21681 , y21682 , y21683 , y21684 , y21685 , y21686 , y21687 , y21688 , y21689 , y21690 , y21691 , y21692 , y21693 , y21694 , y21695 , y21696 , y21697 , y21698 , y21699 , y21700 , y21701 , y21702 , y21703 , y21704 , y21705 , y21706 , y21707 , y21708 , y21709 , y21710 , y21711 , y21712 , y21713 , y21714 , y21715 , y21716 , y21717 , y21718 , y21719 , y21720 , y21721 , y21722 , y21723 , y21724 , y21725 , y21726 , y21727 , y21728 , y21729 , y21730 , y21731 , y21732 , y21733 , y21734 , y21735 , y21736 , y21737 , y21738 , y21739 , y21740 , y21741 , y21742 , y21743 , y21744 , y21745 , y21746 , y21747 , y21748 , y21749 , y21750 , y21751 , y21752 , y21753 , y21754 , y21755 , y21756 , y21757 , y21758 , y21759 , y21760 , y21761 , y21762 , y21763 , y21764 , y21765 , y21766 , y21767 , y21768 , y21769 , y21770 , y21771 , y21772 , y21773 , y21774 , y21775 , y21776 , y21777 , y21778 , y21779 , y21780 , y21781 , y21782 , y21783 , y21784 , y21785 , y21786 , y21787 , y21788 , y21789 , y21790 , y21791 , y21792 , y21793 , y21794 , y21795 , y21796 , y21797 , y21798 , y21799 , y21800 , y21801 , y21802 , y21803 , y21804 , y21805 , y21806 , y21807 , y21808 , y21809 , y21810 , y21811 , y21812 , y21813 , y21814 , y21815 , y21816 , y21817 , y21818 , y21819 , y21820 , y21821 , y21822 , y21823 , y21824 , y21825 , y21826 , y21827 , y21828 , y21829 , y21830 , y21831 , y21832 , y21833 , y21834 , y21835 , y21836 , y21837 , y21838 , y21839 , y21840 , y21841 , y21842 , y21843 , y21844 , y21845 , y21846 , y21847 , y21848 , y21849 , y21850 , y21851 , y21852 , y21853 , y21854 , y21855 , y21856 , y21857 , y21858 , y21859 , y21860 , y21861 , y21862 , y21863 , y21864 , y21865 , y21866 , y21867 , y21868 , y21869 , y21870 , y21871 , y21872 , y21873 , y21874 , y21875 , y21876 , y21877 , y21878 , y21879 , y21880 , y21881 , y21882 , y21883 , y21884 , y21885 , y21886 , y21887 , y21888 , y21889 , y21890 , y21891 , y21892 , y21893 , y21894 , y21895 , y21896 , y21897 , y21898 , y21899 , y21900 , y21901 , y21902 , y21903 , y21904 , y21905 , y21906 , y21907 , y21908 , y21909 , y21910 , y21911 , y21912 , y21913 , y21914 , y21915 , y21916 , y21917 , y21918 , y21919 , y21920 , y21921 , y21922 , y21923 , y21924 , y21925 , y21926 , y21927 , y21928 , y21929 , y21930 , y21931 , y21932 , y21933 , y21934 , y21935 , y21936 , y21937 , y21938 , y21939 , y21940 , y21941 , y21942 , y21943 , y21944 , y21945 , y21946 , y21947 , y21948 , y21949 , y21950 , y21951 , y21952 , y21953 , y21954 , y21955 , y21956 , y21957 , y21958 , y21959 , y21960 , y21961 , y21962 , y21963 , y21964 , y21965 , y21966 , y21967 , y21968 , y21969 , y21970 , y21971 , y21972 , y21973 , y21974 , y21975 , y21976 , y21977 , y21978 , y21979 , y21980 , y21981 , y21982 , y21983 , y21984 , y21985 , y21986 , y21987 , y21988 , y21989 , y21990 , y21991 , y21992 , y21993 , y21994 , y21995 , y21996 , y21997 , y21998 , y21999 , y22000 , y22001 , y22002 , y22003 , y22004 , y22005 , y22006 , y22007 , y22008 , y22009 , y22010 , y22011 , y22012 , y22013 , y22014 , y22015 , y22016 , y22017 , y22018 , y22019 , y22020 , y22021 , y22022 , y22023 , y22024 , y22025 , y22026 , y22027 , y22028 , y22029 , y22030 , y22031 , y22032 , y22033 , y22034 , y22035 , y22036 , y22037 , y22038 , y22039 , y22040 , y22041 , y22042 , y22043 , y22044 , y22045 , y22046 , y22047 , y22048 , y22049 , y22050 , y22051 , y22052 , y22053 , y22054 , y22055 , y22056 , y22057 , y22058 , y22059 , y22060 , y22061 , y22062 , y22063 , y22064 , y22065 , y22066 , y22067 , y22068 , y22069 , y22070 , y22071 , y22072 , y22073 , y22074 , y22075 , y22076 , y22077 , y22078 , y22079 , y22080 , y22081 , y22082 , y22083 , y22084 , y22085 , y22086 , y22087 , y22088 , y22089 , y22090 , y22091 , y22092 , y22093 , y22094 , y22095 , y22096 , y22097 , y22098 , y22099 , y22100 , y22101 , y22102 , y22103 , y22104 , y22105 , y22106 , y22107 , y22108 , y22109 , y22110 , y22111 , y22112 , y22113 , y22114 , y22115 , y22116 , y22117 , y22118 , y22119 , y22120 , y22121 , y22122 , y22123 , y22124 , y22125 , y22126 , y22127 , y22128 , y22129 , y22130 , y22131 , y22132 , y22133 , y22134 , y22135 , y22136 , y22137 , y22138 , y22139 , y22140 , y22141 , y22142 , y22143 , y22144 , y22145 , y22146 , y22147 , y22148 , y22149 , y22150 , y22151 , y22152 , y22153 , y22154 , y22155 , y22156 , y22157 , y22158 , y22159 , y22160 , y22161 , y22162 , y22163 , y22164 , y22165 , y22166 , y22167 , y22168 , y22169 , y22170 , y22171 , y22172 , y22173 , y22174 , y22175 , y22176 , y22177 , y22178 , y22179 , y22180 , y22181 , y22182 , y22183 , y22184 , y22185 , y22186 , y22187 , y22188 , y22189 , y22190 , y22191 , y22192 , y22193 , y22194 , y22195 , y22196 , y22197 , y22198 , y22199 , y22200 , y22201 , y22202 , y22203 , y22204 , y22205 , y22206 , y22207 , y22208 , y22209 , y22210 , y22211 , y22212 , y22213 , y22214 , y22215 , y22216 , y22217 , y22218 , y22219 , y22220 , y22221 , y22222 , y22223 , y22224 , y22225 , y22226 , y22227 , y22228 , y22229 , y22230 , y22231 , y22232 , y22233 , y22234 , y22235 , y22236 , y22237 , y22238 , y22239 , y22240 , y22241 , y22242 , y22243 , y22244 , y22245 , y22246 , y22247 , y22248 , y22249 , y22250 , y22251 , y22252 , y22253 , y22254 , y22255 , y22256 , y22257 , y22258 , y22259 , y22260 , y22261 , y22262 , y22263 , y22264 , y22265 , y22266 , y22267 , y22268 , y22269 , y22270 , y22271 , y22272 , y22273 , y22274 , y22275 , y22276 , y22277 , y22278 , y22279 , y22280 , y22281 , y22282 , y22283 , y22284 , y22285 , y22286 , y22287 , y22288 , y22289 , y22290 , y22291 , y22292 , y22293 , y22294 , y22295 , y22296 , y22297 , y22298 , y22299 , y22300 , y22301 , y22302 , y22303 , y22304 , y22305 , y22306 , y22307 , y22308 , y22309 , y22310 , y22311 , y22312 , y22313 , y22314 , y22315 , y22316 , y22317 , y22318 , y22319 , y22320 , y22321 , y22322 , y22323 , y22324 , y22325 , y22326 , y22327 , y22328 , y22329 , y22330 , y22331 , y22332 , y22333 , y22334 , y22335 , y22336 , y22337 , y22338 , y22339 , y22340 , y22341 , y22342 , y22343 , y22344 , y22345 , y22346 , y22347 , y22348 , y22349 , y22350 , y22351 , y22352 , y22353 , y22354 , y22355 , y22356 , y22357 , y22358 , y22359 , y22360 , y22361 , y22362 , y22363 , y22364 , y22365 , y22366 , y22367 , y22368 , y22369 , y22370 , y22371 , y22372 , y22373 , y22374 , y22375 , y22376 , y22377 , y22378 , y22379 , y22380 , y22381 , y22382 , y22383 , y22384 , y22385 , y22386 , y22387 , y22388 , y22389 , y22390 , y22391 , y22392 , y22393 , y22394 , y22395 , y22396 , y22397 , y22398 , y22399 , y22400 , y22401 , y22402 , y22403 , y22404 , y22405 , y22406 , y22407 , y22408 , y22409 , y22410 , y22411 , y22412 , y22413 , y22414 , y22415 , y22416 , y22417 , y22418 , y22419 , y22420 , y22421 , y22422 , y22423 , y22424 , y22425 , y22426 , y22427 , y22428 , y22429 , y22430 , y22431 , y22432 , y22433 , y22434 , y22435 , y22436 , y22437 , y22438 , y22439 , y22440 , y22441 , y22442 , y22443 , y22444 , y22445 , y22446 , y22447 , y22448 , y22449 , y22450 , y22451 , y22452 , y22453 , y22454 , y22455 , y22456 , y22457 , y22458 , y22459 , y22460 , y22461 , y22462 , y22463 , y22464 , y22465 , y22466 , y22467 , y22468 , y22469 , y22470 , y22471 , y22472 , y22473 , y22474 , y22475 , y22476 , y22477 , y22478 , y22479 , y22480 , y22481 , y22482 , y22483 , y22484 , y22485 , y22486 , y22487 , y22488 , y22489 , y22490 , y22491 , y22492 , y22493 , y22494 , y22495 , y22496 , y22497 , y22498 , y22499 , y22500 , y22501 , y22502 , y22503 , y22504 , y22505 , y22506 , y22507 , y22508 , y22509 , y22510 , y22511 , y22512 , y22513 , y22514 , y22515 , y22516 , y22517 , y22518 , y22519 , y22520 , y22521 , y22522 , y22523 , y22524 , y22525 , y22526 , y22527 , y22528 , y22529 , y22530 , y22531 , y22532 , y22533 , y22534 , y22535 , y22536 , y22537 , y22538 , y22539 , y22540 , y22541 , y22542 , y22543 , y22544 , y22545 , y22546 , y22547 , y22548 , y22549 , y22550 , y22551 , y22552 , y22553 , y22554 , y22555 , y22556 , y22557 , y22558 , y22559 , y22560 , y22561 , y22562 , y22563 , y22564 , y22565 , y22566 , y22567 , y22568 , y22569 , y22570 , y22571 , y22572 , y22573 , y22574 , y22575 , y22576 , y22577 , y22578 , y22579 , y22580 , y22581 , y22582 , y22583 , y22584 , y22585 , y22586 , y22587 , y22588 , y22589 , y22590 , y22591 , y22592 , y22593 , y22594 , y22595 , y22596 , y22597 , y22598 , y22599 , y22600 , y22601 , y22602 , y22603 , y22604 , y22605 , y22606 , y22607 , y22608 , y22609 , y22610 , y22611 , y22612 , y22613 , y22614 , y22615 , y22616 , y22617 , y22618 , y22619 , y22620 , y22621 , y22622 , y22623 , y22624 , y22625 , y22626 , y22627 , y22628 , y22629 , y22630 , y22631 , y22632 , y22633 , y22634 , y22635 , y22636 , y22637 , y22638 , y22639 , y22640 , y22641 , y22642 , y22643 , y22644 , y22645 , y22646 , y22647 , y22648 , y22649 , y22650 , y22651 , y22652 , y22653 , y22654 , y22655 , y22656 , y22657 , y22658 , y22659 , y22660 , y22661 , y22662 , y22663 , y22664 , y22665 , y22666 , y22667 , y22668 , y22669 , y22670 , y22671 , y22672 , y22673 , y22674 , y22675 , y22676 , y22677 , y22678 , y22679 , y22680 , y22681 , y22682 , y22683 , y22684 , y22685 , y22686 , y22687 , y22688 , y22689 , y22690 , y22691 , y22692 , y22693 , y22694 , y22695 , y22696 , y22697 , y22698 , y22699 , y22700 , y22701 , y22702 , y22703 , y22704 , y22705 , y22706 , y22707 , y22708 , y22709 , y22710 , y22711 , y22712 , y22713 , y22714 , y22715 , y22716 , y22717 , y22718 , y22719 , y22720 , y22721 , y22722 , y22723 , y22724 , y22725 , y22726 , y22727 , y22728 , y22729 , y22730 , y22731 , y22732 , y22733 , y22734 , y22735 , y22736 , y22737 , y22738 , y22739 , y22740 , y22741 , y22742 , y22743 , y22744 , y22745 , y22746 , y22747 , y22748 , y22749 , y22750 , y22751 , y22752 , y22753 , y22754 , y22755 , y22756 , y22757 , y22758 , y22759 , y22760 , y22761 , y22762 , y22763 , y22764 , y22765 , y22766 , y22767 , y22768 , y22769 , y22770 , y22771 , y22772 , y22773 , y22774 , y22775 , y22776 , y22777 , y22778 , y22779 , y22780 , y22781 , y22782 , y22783 , y22784 , y22785 , y22786 , y22787 , y22788 , y22789 , y22790 , y22791 , y22792 , y22793 , y22794 , y22795 , y22796 , y22797 , y22798 , y22799 , y22800 , y22801 , y22802 , y22803 , y22804 , y22805 , y22806 , y22807 , y22808 , y22809 , y22810 , y22811 , y22812 , y22813 , y22814 , y22815 , y22816 , y22817 , y22818 , y22819 , y22820 , y22821 , y22822 , y22823 , y22824 , y22825 , y22826 , y22827 , y22828 , y22829 , y22830 , y22831 , y22832 , y22833 , y22834 , y22835 , y22836 , y22837 , y22838 , y22839 , y22840 , y22841 , y22842 , y22843 , y22844 , y22845 , y22846 , y22847 , y22848 , y22849 , y22850 , y22851 , y22852 , y22853 , y22854 , y22855 , y22856 , y22857 , y22858 , y22859 , y22860 , y22861 , y22862 , y22863 , y22864 , y22865 , y22866 , y22867 , y22868 , y22869 , y22870 , y22871 , y22872 , y22873 , y22874 , y22875 , y22876 , y22877 , y22878 , y22879 , y22880 , y22881 , y22882 , y22883 , y22884 , y22885 , y22886 , y22887 , y22888 , y22889 , y22890 , y22891 , y22892 , y22893 , y22894 , y22895 , y22896 , y22897 , y22898 , y22899 , y22900 , y22901 , y22902 , y22903 , y22904 , y22905 , y22906 , y22907 , y22908 , y22909 , y22910 , y22911 , y22912 , y22913 , y22914 , y22915 , y22916 , y22917 , y22918 , y22919 , y22920 , y22921 , y22922 , y22923 , y22924 , y22925 , y22926 , y22927 , y22928 , y22929 , y22930 , y22931 , y22932 , y22933 , y22934 , y22935 , y22936 , y22937 , y22938 , y22939 , y22940 , y22941 , y22942 , y22943 , y22944 , y22945 , y22946 , y22947 , y22948 , y22949 , y22950 , y22951 , y22952 , y22953 , y22954 , y22955 , y22956 , y22957 , y22958 , y22959 , y22960 , y22961 , y22962 , y22963 , y22964 , y22965 , y22966 , y22967 , y22968 , y22969 , y22970 , y22971 , y22972 , y22973 , y22974 , y22975 , y22976 , y22977 , y22978 , y22979 , y22980 , y22981 , y22982 , y22983 , y22984 , y22985 , y22986 , y22987 , y22988 , y22989 , y22990 , y22991 , y22992 , y22993 , y22994 , y22995 , y22996 , y22997 , y22998 , y22999 , y23000 , y23001 , y23002 , y23003 , y23004 , y23005 , y23006 , y23007 , y23008 , y23009 , y23010 , y23011 , y23012 , y23013 , y23014 , y23015 , y23016 , y23017 , y23018 , y23019 , y23020 , y23021 , y23022 , y23023 , y23024 , y23025 , y23026 , y23027 , y23028 , y23029 , y23030 , y23031 , y23032 , y23033 , y23034 , y23035 , y23036 , y23037 , y23038 , y23039 , y23040 , y23041 , y23042 , y23043 , y23044 , y23045 , y23046 , y23047 , y23048 , y23049 , y23050 , y23051 , y23052 , y23053 , y23054 , y23055 , y23056 , y23057 , y23058 , y23059 , y23060 , y23061 , y23062 , y23063 , y23064 , y23065 , y23066 , y23067 , y23068 , y23069 , y23070 , y23071 , y23072 , y23073 , y23074 , y23075 , y23076 , y23077 , y23078 , y23079 , y23080 , y23081 , y23082 , y23083 , y23084 , y23085 , y23086 , y23087 , y23088 , y23089 , y23090 , y23091 , y23092 , y23093 , y23094 , y23095 , y23096 , y23097 , y23098 , y23099 , y23100 , y23101 , y23102 , y23103 , y23104 , y23105 , y23106 , y23107 , y23108 , y23109 , y23110 , y23111 , y23112 , y23113 , y23114 , y23115 , y23116 , y23117 , y23118 , y23119 , y23120 , y23121 , y23122 , y23123 , y23124 , y23125 , y23126 , y23127 , y23128 , y23129 , y23130 , y23131 , y23132 , y23133 , y23134 , y23135 , y23136 , y23137 , y23138 , y23139 , y23140 , y23141 , y23142 , y23143 , y23144 , y23145 , y23146 , y23147 , y23148 , y23149 , y23150 , y23151 , y23152 , y23153 , y23154 , y23155 , y23156 , y23157 , y23158 , y23159 , y23160 , y23161 , y23162 , y23163 , y23164 , y23165 , y23166 , y23167 , y23168 , y23169 , y23170 , y23171 , y23172 , y23173 , y23174 , y23175 , y23176 , y23177 , y23178 , y23179 , y23180 , y23181 , y23182 , y23183 , y23184 , y23185 , y23186 , y23187 , y23188 , y23189 , y23190 , y23191 , y23192 , y23193 , y23194 , y23195 , y23196 , y23197 , y23198 , y23199 , y23200 , y23201 , y23202 , y23203 , y23204 , y23205 , y23206 , y23207 , y23208 , y23209 , y23210 , y23211 , y23212 , y23213 , y23214 , y23215 , y23216 , y23217 , y23218 , y23219 , y23220 , y23221 , y23222 , y23223 , y23224 , y23225 , y23226 , y23227 , y23228 , y23229 , y23230 , y23231 , y23232 , y23233 , y23234 , y23235 , y23236 , y23237 , y23238 , y23239 , y23240 , y23241 , y23242 , y23243 , y23244 , y23245 , y23246 , y23247 , y23248 , y23249 , y23250 , y23251 , y23252 , y23253 , y23254 , y23255 , y23256 , y23257 , y23258 , y23259 , y23260 , y23261 , y23262 , y23263 , y23264 , y23265 , y23266 , y23267 , y23268 , y23269 , y23270 , y23271 , y23272 , y23273 , y23274 , y23275 , y23276 , y23277 , y23278 , y23279 , y23280 , y23281 , y23282 , y23283 , y23284 , y23285 , y23286 , y23287 , y23288 , y23289 , y23290 , y23291 , y23292 , y23293 , y23294 , y23295 , y23296 , y23297 , y23298 , y23299 , y23300 , y23301 , y23302 , y23303 , y23304 , y23305 , y23306 , y23307 , y23308 , y23309 , y23310 , y23311 , y23312 , y23313 , y23314 , y23315 , y23316 , y23317 , y23318 , y23319 , y23320 , y23321 , y23322 , y23323 , y23324 , y23325 , y23326 , y23327 , y23328 , y23329 , y23330 , y23331 , y23332 , y23333 , y23334 , y23335 , y23336 , y23337 , y23338 , y23339 , y23340 , y23341 , y23342 , y23343 , y23344 , y23345 , y23346 , y23347 , y23348 , y23349 , y23350 , y23351 , y23352 , y23353 , y23354 , y23355 , y23356 , y23357 , y23358 , y23359 , y23360 , y23361 , y23362 , y23363 , y23364 , y23365 , y23366 , y23367 , y23368 , y23369 , y23370 , y23371 , y23372 , y23373 , y23374 , y23375 , y23376 , y23377 , y23378 , y23379 , y23380 , y23381 , y23382 , y23383 , y23384 , y23385 , y23386 , y23387 , y23388 , y23389 , y23390 , y23391 , y23392 , y23393 , y23394 , y23395 , y23396 , y23397 , y23398 , y23399 , y23400 , y23401 , y23402 , y23403 , y23404 , y23405 , y23406 , y23407 , y23408 , y23409 , y23410 , y23411 , y23412 , y23413 , y23414 , y23415 , y23416 , y23417 , y23418 , y23419 , y23420 , y23421 , y23422 , y23423 , y23424 , y23425 , y23426 , y23427 , y23428 , y23429 , y23430 , y23431 , y23432 , y23433 , y23434 , y23435 , y23436 , y23437 , y23438 , y23439 , y23440 , y23441 , y23442 , y23443 , y23444 , y23445 , y23446 , y23447 , y23448 , y23449 , y23450 , y23451 , y23452 , y23453 , y23454 , y23455 , y23456 , y23457 , y23458 , y23459 , y23460 , y23461 , y23462 , y23463 , y23464 , y23465 , y23466 , y23467 , y23468 , y23469 , y23470 , y23471 , y23472 , y23473 , y23474 , y23475 , y23476 , y23477 , y23478 , y23479 , y23480 , y23481 , y23482 , y23483 , y23484 , y23485 , y23486 , y23487 , y23488 , y23489 , y23490 , y23491 , y23492 , y23493 , y23494 , y23495 , y23496 , y23497 , y23498 , y23499 , y23500 , y23501 , y23502 , y23503 , y23504 , y23505 , y23506 , y23507 , y23508 , y23509 , y23510 , y23511 , y23512 , y23513 , y23514 , y23515 , y23516 , y23517 , y23518 , y23519 , y23520 , y23521 , y23522 , y23523 , y23524 , y23525 , y23526 , y23527 , y23528 , y23529 , y23530 , y23531 , y23532 , y23533 , y23534 , y23535 , y23536 , y23537 , y23538 , y23539 , y23540 , y23541 , y23542 , y23543 , y23544 , y23545 , y23546 , y23547 , y23548 , y23549 , y23550 , y23551 , y23552 , y23553 , y23554 , y23555 , y23556 , y23557 , y23558 , y23559 , y23560 , y23561 , y23562 , y23563 , y23564 , y23565 , y23566 , y23567 , y23568 , y23569 , y23570 , y23571 , y23572 , y23573 , y23574 , y23575 , y23576 , y23577 , y23578 , y23579 , y23580 , y23581 , y23582 , y23583 , y23584 , y23585 , y23586 , y23587 , y23588 , y23589 , y23590 , y23591 , y23592 , y23593 , y23594 , y23595 , y23596 , y23597 , y23598 , y23599 , y23600 , y23601 , y23602 , y23603 , y23604 , y23605 , y23606 , y23607 , y23608 , y23609 , y23610 , y23611 , y23612 , y23613 , y23614 , y23615 , y23616 , y23617 , y23618 , y23619 , y23620 , y23621 , y23622 , y23623 , y23624 , y23625 , y23626 , y23627 , y23628 , y23629 , y23630 , y23631 , y23632 , y23633 , y23634 , y23635 , y23636 , y23637 , y23638 , y23639 , y23640 , y23641 , y23642 , y23643 , y23644 , y23645 , y23646 , y23647 , y23648 , y23649 , y23650 , y23651 , y23652 , y23653 , y23654 , y23655 , y23656 , y23657 , y23658 , y23659 , y23660 , y23661 , y23662 , y23663 , y23664 , y23665 , y23666 , y23667 , y23668 , y23669 , y23670 , y23671 , y23672 , y23673 , y23674 , y23675 , y23676 , y23677 , y23678 , y23679 , y23680 , y23681 , y23682 , y23683 , y23684 , y23685 , y23686 , y23687 , y23688 , y23689 , y23690 , y23691 , y23692 , y23693 , y23694 , y23695 , y23696 , y23697 , y23698 , y23699 , y23700 , y23701 , y23702 , y23703 , y23704 , y23705 , y23706 , y23707 , y23708 , y23709 , y23710 , y23711 , y23712 , y23713 , y23714 , y23715 , y23716 , y23717 , y23718 , y23719 , y23720 , y23721 , y23722 , y23723 , y23724 , y23725 , y23726 , y23727 , y23728 , y23729 , y23730 , y23731 , y23732 , y23733 , y23734 , y23735 , y23736 , y23737 , y23738 , y23739 , y23740 , y23741 , y23742 , y23743 , y23744 , y23745 , y23746 , y23747 , y23748 , y23749 , y23750 , y23751 , y23752 , y23753 , y23754 , y23755 , y23756 , y23757 , y23758 , y23759 , y23760 , y23761 , y23762 , y23763 , y23764 , y23765 , y23766 , y23767 , y23768 , y23769 , y23770 , y23771 , y23772 , y23773 , y23774 , y23775 , y23776 , y23777 , y23778 , y23779 , y23780 , y23781 , y23782 , y23783 , y23784 , y23785 , y23786 , y23787 , y23788 , y23789 , y23790 , y23791 , y23792 , y23793 , y23794 , y23795 , y23796 , y23797 , y23798 , y23799 , y23800 , y23801 , y23802 , y23803 , y23804 , y23805 , y23806 , y23807 , y23808 , y23809 , y23810 , y23811 , y23812 , y23813 , y23814 , y23815 , y23816 , y23817 , y23818 , y23819 , y23820 , y23821 , y23822 , y23823 , y23824 , y23825 , y23826 , y23827 , y23828 , y23829 , y23830 , y23831 , y23832 , y23833 , y23834 , y23835 , y23836 , y23837 , y23838 , y23839 , y23840 , y23841 , y23842 , y23843 , y23844 , y23845 , y23846 , y23847 , y23848 , y23849 , y23850 , y23851 , y23852 , y23853 , y23854 , y23855 , y23856 , y23857 , y23858 , y23859 , y23860 , y23861 , y23862 , y23863 , y23864 , y23865 , y23866 , y23867 , y23868 , y23869 , y23870 , y23871 , y23872 , y23873 , y23874 , y23875 , y23876 , y23877 , y23878 , y23879 , y23880 , y23881 , y23882 , y23883 , y23884 , y23885 , y23886 , y23887 , y23888 , y23889 , y23890 , y23891 , y23892 , y23893 , y23894 , y23895 , y23896 , y23897 , y23898 , y23899 , y23900 , y23901 , y23902 , y23903 , y23904 , y23905 , y23906 , y23907 , y23908 , y23909 , y23910 , y23911 , y23912 , y23913 , y23914 , y23915 , y23916 , y23917 , y23918 , y23919 , y23920 , y23921 , y23922 , y23923 , y23924 , y23925 , y23926 , y23927 , y23928 , y23929 , y23930 , y23931 , y23932 , y23933 , y23934 , y23935 , y23936 , y23937 , y23938 , y23939 , y23940 , y23941 , y23942 , y23943 , y23944 , y23945 , y23946 , y23947 , y23948 , y23949 , y23950 , y23951 , y23952 , y23953 , y23954 , y23955 , y23956 , y23957 , y23958 , y23959 , y23960 , y23961 , y23962 , y23963 , y23964 , y23965 , y23966 , y23967 , y23968 , y23969 , y23970 , y23971 , y23972 , y23973 , y23974 , y23975 , y23976 , y23977 , y23978 , y23979 , y23980 , y23981 , y23982 , y23983 , y23984 , y23985 , y23986 , y23987 , y23988 , y23989 , y23990 , y23991 , y23992 , y23993 , y23994 , y23995 , y23996 , y23997 , y23998 , y23999 , y24000 , y24001 , y24002 , y24003 , y24004 , y24005 , y24006 , y24007 , y24008 , y24009 , y24010 , y24011 , y24012 , y24013 , y24014 , y24015 , y24016 , y24017 , y24018 , y24019 , y24020 , y24021 , y24022 , y24023 , y24024 , y24025 , y24026 , y24027 , y24028 , y24029 , y24030 , y24031 , y24032 , y24033 , y24034 , y24035 , y24036 , y24037 , y24038 , y24039 , y24040 , y24041 , y24042 , y24043 , y24044 , y24045 , y24046 , y24047 , y24048 , y24049 , y24050 , y24051 , y24052 , y24053 , y24054 , y24055 , y24056 , y24057 , y24058 , y24059 , y24060 , y24061 , y24062 , y24063 , y24064 , y24065 , y24066 , y24067 , y24068 , y24069 , y24070 , y24071 , y24072 , y24073 , y24074 , y24075 , y24076 , y24077 , y24078 , y24079 , y24080 , y24081 , y24082 , y24083 , y24084 , y24085 , y24086 , y24087 , y24088 , y24089 , y24090 , y24091 , y24092 , y24093 , y24094 , y24095 , y24096 , y24097 , y24098 , y24099 , y24100 , y24101 , y24102 , y24103 , y24104 , y24105 , y24106 , y24107 , y24108 , y24109 , y24110 , y24111 , y24112 , y24113 , y24114 , y24115 , y24116 , y24117 , y24118 , y24119 , y24120 , y24121 , y24122 , y24123 , y24124 , y24125 , y24126 , y24127 , y24128 , y24129 , y24130 , y24131 , y24132 , y24133 , y24134 , y24135 , y24136 , y24137 , y24138 , y24139 , y24140 , y24141 , y24142 , y24143 , y24144 , y24145 , y24146 , y24147 , y24148 , y24149 , y24150 , y24151 , y24152 , y24153 , y24154 , y24155 , y24156 , y24157 , y24158 , y24159 , y24160 , y24161 , y24162 , y24163 , y24164 , y24165 , y24166 , y24167 , y24168 , y24169 , y24170 , y24171 , y24172 , y24173 , y24174 , y24175 , y24176 , y24177 , y24178 , y24179 , y24180 , y24181 , y24182 , y24183 , y24184 , y24185 , y24186 , y24187 , y24188 , y24189 , y24190 , y24191 , y24192 , y24193 , y24194 , y24195 , y24196 , y24197 , y24198 , y24199 , y24200 , y24201 , y24202 , y24203 , y24204 , y24205 , y24206 , y24207 , y24208 , y24209 , y24210 , y24211 , y24212 , y24213 , y24214 , y24215 , y24216 , y24217 , y24218 , y24219 , y24220 , y24221 , y24222 , y24223 , y24224 , y24225 , y24226 , y24227 , y24228 , y24229 , y24230 , y24231 , y24232 , y24233 , y24234 , y24235 , y24236 , y24237 , y24238 , y24239 , y24240 , y24241 , y24242 , y24243 , y24244 , y24245 , y24246 , y24247 , y24248 , y24249 , y24250 , y24251 , y24252 , y24253 , y24254 , y24255 , y24256 , y24257 , y24258 , y24259 , y24260 , y24261 , y24262 , y24263 , y24264 , y24265 , y24266 , y24267 , y24268 , y24269 , y24270 , y24271 , y24272 , y24273 , y24274 , y24275 , y24276 , y24277 , y24278 , y24279 , y24280 , y24281 , y24282 , y24283 , y24284 , y24285 , y24286 , y24287 , y24288 , y24289 , y24290 , y24291 , y24292 , y24293 , y24294 , y24295 , y24296 , y24297 , y24298 , y24299 , y24300 , y24301 , y24302 , y24303 , y24304 , y24305 , y24306 , y24307 , y24308 , y24309 , y24310 , y24311 , y24312 , y24313 , y24314 , y24315 , y24316 , y24317 , y24318 , y24319 , y24320 , y24321 , y24322 , y24323 , y24324 , y24325 , y24326 , y24327 , y24328 , y24329 , y24330 , y24331 , y24332 , y24333 , y24334 , y24335 , y24336 , y24337 , y24338 , y24339 , y24340 , y24341 , y24342 , y24343 , y24344 , y24345 , y24346 , y24347 , y24348 , y24349 , y24350 , y24351 , y24352 , y24353 , y24354 , y24355 , y24356 , y24357 , y24358 , y24359 , y24360 , y24361 , y24362 , y24363 , y24364 , y24365 , y24366 , y24367 , y24368 , y24369 , y24370 , y24371 , y24372 , y24373 , y24374 , y24375 , y24376 , y24377 , y24378 , y24379 , y24380 , y24381 , y24382 , y24383 , y24384 , y24385 , y24386 , y24387 , y24388 , y24389 , y24390 , y24391 , y24392 , y24393 , y24394 , y24395 , y24396 , y24397 , y24398 , y24399 , y24400 , y24401 , y24402 , y24403 , y24404 , y24405 , y24406 , y24407 , y24408 , y24409 , y24410 , y24411 , y24412 , y24413 , y24414 , y24415 , y24416 , y24417 , y24418 , y24419 , y24420 , y24421 , y24422 , y24423 , y24424 , y24425 , y24426 , y24427 , y24428 , y24429 , y24430 , y24431 , y24432 , y24433 , y24434 , y24435 , y24436 , y24437 , y24438 , y24439 , y24440 , y24441 , y24442 , y24443 , y24444 , y24445 , y24446 , y24447 , y24448 , y24449 , y24450 , y24451 , y24452 , y24453 , y24454 , y24455 , y24456 , y24457 , y24458 , y24459 , y24460 , y24461 , y24462 , y24463 , y24464 , y24465 , y24466 , y24467 , y24468 , y24469 , y24470 , y24471 , y24472 , y24473 , y24474 , y24475 , y24476 , y24477 , y24478 , y24479 , y24480 , y24481 , y24482 , y24483 , y24484 , y24485 , y24486 , y24487 , y24488 , y24489 , y24490 , y24491 , y24492 , y24493 , y24494 , y24495 , y24496 , y24497 , y24498 , y24499 , y24500 , y24501 , y24502 , y24503 , y24504 , y24505 , y24506 , y24507 , y24508 , y24509 , y24510 , y24511 , y24512 , y24513 , y24514 , y24515 , y24516 , y24517 , y24518 , y24519 , y24520 , y24521 , y24522 , y24523 , y24524 , y24525 , y24526 , y24527 , y24528 , y24529 , y24530 , y24531 , y24532 , y24533 , y24534 , y24535 , y24536 , y24537 , y24538 , y24539 , y24540 , y24541 , y24542 , y24543 , y24544 , y24545 , y24546 , y24547 , y24548 , y24549 , y24550 , y24551 , y24552 , y24553 , y24554 , y24555 , y24556 , y24557 , y24558 , y24559 , y24560 , y24561 , y24562 , y24563 , y24564 , y24565 , y24566 , y24567 , y24568 , y24569 , y24570 , y24571 , y24572 , y24573 , y24574 , y24575 , y24576 , y24577 , y24578 , y24579 , y24580 , y24581 , y24582 , y24583 , y24584 , y24585 , y24586 , y24587 , y24588 , y24589 , y24590 , y24591 , y24592 , y24593 , y24594 , y24595 , y24596 , y24597 , y24598 , y24599 , y24600 , y24601 , y24602 , y24603 , y24604 , y24605 , y24606 , y24607 , y24608 , y24609 , y24610 , y24611 , y24612 , y24613 , y24614 , y24615 , y24616 , y24617 , y24618 , y24619 , y24620 , y24621 , y24622 , y24623 , y24624 , y24625 , y24626 , y24627 , y24628 , y24629 , y24630 , y24631 , y24632 , y24633 , y24634 , y24635 , y24636 , y24637 , y24638 , y24639 , y24640 , y24641 , y24642 , y24643 , y24644 , y24645 , y24646 , y24647 , y24648 , y24649 , y24650 , y24651 , y24652 , y24653 , y24654 , y24655 , y24656 , y24657 , y24658 , y24659 , y24660 , y24661 , y24662 , y24663 , y24664 , y24665 , y24666 , y24667 , y24668 , y24669 , y24670 , y24671 , y24672 , y24673 , y24674 , y24675 , y24676 , y24677 , y24678 , y24679 , y24680 , y24681 , y24682 , y24683 , y24684 , y24685 , y24686 , y24687 , y24688 , y24689 , y24690 , y24691 , y24692 , y24693 , y24694 , y24695 , y24696 , y24697 , y24698 , y24699 , y24700 , y24701 , y24702 , y24703 , y24704 , y24705 , y24706 , y24707 , y24708 , y24709 , y24710 , y24711 , y24712 , y24713 , y24714 , y24715 , y24716 , y24717 , y24718 , y24719 , y24720 , y24721 , y24722 , y24723 , y24724 , y24725 , y24726 , y24727 , y24728 , y24729 , y24730 , y24731 , y24732 , y24733 , y24734 , y24735 , y24736 , y24737 , y24738 , y24739 , y24740 , y24741 , y24742 , y24743 , y24744 , y24745 , y24746 , y24747 , y24748 , y24749 , y24750 , y24751 , y24752 , y24753 , y24754 , y24755 , y24756 , y24757 , y24758 , y24759 , y24760 , y24761 , y24762 , y24763 , y24764 , y24765 , y24766 , y24767 , y24768 , y24769 , y24770 , y24771 , y24772 , y24773 , y24774 , y24775 , y24776 , y24777 , y24778 , y24779 , y24780 , y24781 , y24782 , y24783 , y24784 , y24785 , y24786 , y24787 , y24788 , y24789 , y24790 , y24791 , y24792 , y24793 , y24794 , y24795 , y24796 , y24797 , y24798 , y24799 , y24800 , y24801 , y24802 , y24803 , y24804 , y24805 , y24806 , y24807 , y24808 , y24809 , y24810 , y24811 , y24812 , y24813 , y24814 , y24815 , y24816 , y24817 , y24818 , y24819 , y24820 , y24821 , y24822 , y24823 , y24824 , y24825 , y24826 , y24827 , y24828 , y24829 , y24830 , y24831 , y24832 , y24833 , y24834 , y24835 , y24836 , y24837 , y24838 , y24839 , y24840 , y24841 , y24842 , y24843 , y24844 , y24845 , y24846 , y24847 , y24848 , y24849 , y24850 , y24851 , y24852 , y24853 , y24854 , y24855 , y24856 , y24857 , y24858 , y24859 , y24860 , y24861 , y24862 , y24863 , y24864 , y24865 , y24866 , y24867 , y24868 , y24869 , y24870 , y24871 , y24872 , y24873 , y24874 , y24875 , y24876 , y24877 , y24878 , y24879 , y24880 , y24881 , y24882 , y24883 , y24884 , y24885 , y24886 , y24887 , y24888 , y24889 , y24890 , y24891 , y24892 , y24893 , y24894 , y24895 , y24896 , y24897 , y24898 , y24899 , y24900 , y24901 , y24902 , y24903 , y24904 , y24905 , y24906 , y24907 , y24908 , y24909 , y24910 , y24911 , y24912 , y24913 , y24914 , y24915 , y24916 , y24917 , y24918 , y24919 , y24920 , y24921 , y24922 , y24923 , y24924 , y24925 , y24926 , y24927 , y24928 , y24929 , y24930 , y24931 , y24932 , y24933 , y24934 , y24935 , y24936 , y24937 , y24938 , y24939 , y24940 , y24941 , y24942 , y24943 , y24944 , y24945 , y24946 , y24947 , y24948 , y24949 , y24950 , y24951 , y24952 , y24953 , y24954 , y24955 , y24956 , y24957 , y24958 , y24959 , y24960 , y24961 , y24962 , y24963 , y24964 , y24965 , y24966 , y24967 , y24968 , y24969 , y24970 , y24971 , y24972 , y24973 , y24974 , y24975 , y24976 , y24977 , y24978 , y24979 , y24980 , y24981 , y24982 , y24983 , y24984 , y24985 , y24986 , y24987 , y24988 , y24989 , y24990 , y24991 , y24992 , y24993 , y24994 , y24995 , y24996 , y24997 , y24998 , y24999 , y25000 , y25001 , y25002 , y25003 , y25004 , y25005 , y25006 , y25007 , y25008 , y25009 , y25010 , y25011 , y25012 , y25013 , y25014 , y25015 , y25016 , y25017 , y25018 , y25019 , y25020 , y25021 , y25022 , y25023 , y25024 , y25025 , y25026 , y25027 , y25028 , y25029 , y25030 , y25031 , y25032 , y25033 , y25034 , y25035 , y25036 , y25037 , y25038 , y25039 , y25040 , y25041 , y25042 , y25043 , y25044 , y25045 , y25046 , y25047 , y25048 , y25049 , y25050 , y25051 , y25052 , y25053 , y25054 , y25055 , y25056 , y25057 , y25058 , y25059 , y25060 , y25061 , y25062 , y25063 , y25064 , y25065 , y25066 , y25067 , y25068 , y25069 , y25070 , y25071 , y25072 , y25073 , y25074 , y25075 , y25076 , y25077 , y25078 , y25079 , y25080 , y25081 , y25082 , y25083 , y25084 , y25085 , y25086 , y25087 , y25088 , y25089 , y25090 , y25091 , y25092 , y25093 , y25094 , y25095 , y25096 , y25097 , y25098 , y25099 , y25100 , y25101 , y25102 , y25103 , y25104 , y25105 , y25106 , y25107 , y25108 , y25109 , y25110 , y25111 , y25112 , y25113 , y25114 , y25115 , y25116 , y25117 , y25118 , y25119 , y25120 , y25121 , y25122 , y25123 , y25124 , y25125 , y25126 , y25127 , y25128 , y25129 , y25130 , y25131 , y25132 , y25133 , y25134 , y25135 , y25136 , y25137 , y25138 , y25139 , y25140 , y25141 , y25142 , y25143 , y25144 , y25145 , y25146 , y25147 , y25148 , y25149 , y25150 , y25151 , y25152 , y25153 , y25154 , y25155 , y25156 , y25157 , y25158 , y25159 , y25160 , y25161 , y25162 , y25163 , y25164 , y25165 , y25166 , y25167 , y25168 , y25169 , y25170 , y25171 , y25172 , y25173 , y25174 , y25175 , y25176 , y25177 , y25178 , y25179 , y25180 , y25181 , y25182 , y25183 , y25184 , y25185 , y25186 , y25187 , y25188 , y25189 , y25190 , y25191 , y25192 , y25193 , y25194 , y25195 , y25196 , y25197 , y25198 , y25199 , y25200 , y25201 , y25202 , y25203 , y25204 , y25205 , y25206 , y25207 , y25208 , y25209 , y25210 , y25211 , y25212 , y25213 , y25214 , y25215 , y25216 , y25217 , y25218 , y25219 , y25220 , y25221 , y25222 , y25223 , y25224 , y25225 , y25226 , y25227 , y25228 , y25229 , y25230 , y25231 , y25232 , y25233 , y25234 , y25235 , y25236 , y25237 , y25238 , y25239 , y25240 , y25241 , y25242 , y25243 , y25244 , y25245 , y25246 , y25247 , y25248 , y25249 , y25250 , y25251 , y25252 , y25253 , y25254 , y25255 , y25256 , y25257 , y25258 , y25259 , y25260 , y25261 , y25262 , y25263 , y25264 , y25265 , y25266 , y25267 , y25268 , y25269 , y25270 , y25271 , y25272 , y25273 , y25274 , y25275 , y25276 , y25277 , y25278 , y25279 , y25280 , y25281 , y25282 , y25283 , y25284 , y25285 , y25286 , y25287 , y25288 , y25289 , y25290 , y25291 , y25292 , y25293 , y25294 , y25295 , y25296 , y25297 , y25298 , y25299 , y25300 , y25301 , y25302 , y25303 , y25304 , y25305 , y25306 , y25307 , y25308 , y25309 , y25310 , y25311 , y25312 , y25313 , y25314 , y25315 , y25316 , y25317 , y25318 , y25319 , y25320 , y25321 , y25322 , y25323 , y25324 , y25325 , y25326 , y25327 , y25328 , y25329 , y25330 , y25331 , y25332 , y25333 , y25334 , y25335 , y25336 , y25337 , y25338 , y25339 , y25340 , y25341 , y25342 , y25343 , y25344 , y25345 , y25346 , y25347 , y25348 , y25349 , y25350 , y25351 , y25352 , y25353 , y25354 , y25355 , y25356 , y25357 , y25358 , y25359 , y25360 , y25361 , y25362 , y25363 , y25364 , y25365 , y25366 , y25367 , y25368 , y25369 , y25370 , y25371 , y25372 , y25373 , y25374 , y25375 , y25376 , y25377 , y25378 , y25379 , y25380 , y25381 , y25382 , y25383 , y25384 , y25385 , y25386 , y25387 , y25388 , y25389 , y25390 , y25391 , y25392 , y25393 , y25394 , y25395 , y25396 , y25397 , y25398 , y25399 , y25400 , y25401 , y25402 , y25403 , y25404 , y25405 , y25406 , y25407 , y25408 , y25409 , y25410 , y25411 , y25412 , y25413 , y25414 , y25415 , y25416 , y25417 , y25418 , y25419 , y25420 , y25421 , y25422 , y25423 , y25424 , y25425 , y25426 , y25427 , y25428 , y25429 , y25430 , y25431 , y25432 , y25433 , y25434 , y25435 , y25436 , y25437 , y25438 , y25439 , y25440 , y25441 , y25442 , y25443 , y25444 , y25445 , y25446 , y25447 , y25448 , y25449 , y25450 , y25451 , y25452 , y25453 , y25454 , y25455 , y25456 , y25457 , y25458 , y25459 , y25460 , y25461 , y25462 , y25463 , y25464 , y25465 , y25466 , y25467 , y25468 , y25469 , y25470 , y25471 , y25472 , y25473 , y25474 , y25475 , y25476 , y25477 , y25478 , y25479 , y25480 , y25481 , y25482 , y25483 , y25484 , y25485 , y25486 , y25487 , y25488 , y25489 , y25490 , y25491 , y25492 , y25493 , y25494 , y25495 , y25496 , y25497 , y25498 , y25499 , y25500 , y25501 , y25502 , y25503 , y25504 , y25505 , y25506 , y25507 , y25508 , y25509 , y25510 , y25511 , y25512 , y25513 , y25514 , y25515 , y25516 , y25517 , y25518 , y25519 , y25520 , y25521 , y25522 , y25523 , y25524 , y25525 , y25526 , y25527 , y25528 , y25529 , y25530 , y25531 , y25532 , y25533 , y25534 , y25535 , y25536 , y25537 , y25538 , y25539 , y25540 , y25541 , y25542 , y25543 , y25544 , y25545 , y25546 , y25547 , y25548 , y25549 , y25550 , y25551 , y25552 , y25553 , y25554 , y25555 , y25556 , y25557 , y25558 , y25559 , y25560 , y25561 , y25562 , y25563 , y25564 , y25565 , y25566 , y25567 , y25568 , y25569 , y25570 , y25571 , y25572 , y25573 , y25574 , y25575 , y25576 , y25577 , y25578 , y25579 , y25580 , y25581 , y25582 , y25583 , y25584 , y25585 , y25586 , y25587 , y25588 , y25589 , y25590 , y25591 , y25592 , y25593 , y25594 , y25595 , y25596 , y25597 , y25598 , y25599 , y25600 , y25601 , y25602 , y25603 , y25604 , y25605 , y25606 , y25607 , y25608 , y25609 , y25610 , y25611 , y25612 , y25613 , y25614 , y25615 , y25616 , y25617 , y25618 , y25619 , y25620 , y25621 , y25622 , y25623 , y25624 , y25625 , y25626 , y25627 , y25628 , y25629 , y25630 , y25631 , y25632 , y25633 , y25634 , y25635 , y25636 , y25637 , y25638 , y25639 , y25640 , y25641 , y25642 , y25643 , y25644 , y25645 , y25646 , y25647 , y25648 , y25649 , y25650 , y25651 , y25652 , y25653 , y25654 , y25655 , y25656 , y25657 , y25658 , y25659 , y25660 , y25661 , y25662 , y25663 , y25664 , y25665 , y25666 , y25667 , y25668 , y25669 , y25670 , y25671 , y25672 , y25673 , y25674 , y25675 , y25676 , y25677 , y25678 , y25679 , y25680 , y25681 , y25682 , y25683 , y25684 , y25685 , y25686 , y25687 , y25688 , y25689 , y25690 , y25691 , y25692 , y25693 , y25694 , y25695 , y25696 , y25697 , y25698 , y25699 , y25700 , y25701 , y25702 , y25703 , y25704 , y25705 , y25706 , y25707 , y25708 , y25709 , y25710 , y25711 , y25712 , y25713 , y25714 , y25715 , y25716 , y25717 , y25718 , y25719 , y25720 , y25721 , y25722 , y25723 , y25724 , y25725 , y25726 , y25727 , y25728 , y25729 , y25730 , y25731 , y25732 , y25733 , y25734 , y25735 , y25736 , y25737 , y25738 , y25739 , y25740 , y25741 , y25742 , y25743 , y25744 , y25745 , y25746 , y25747 , y25748 , y25749 , y25750 , y25751 , y25752 , y25753 , y25754 , y25755 , y25756 , y25757 , y25758 , y25759 , y25760 , y25761 , y25762 , y25763 , y25764 , y25765 , y25766 , y25767 , y25768 , y25769 , y25770 , y25771 , y25772 , y25773 , y25774 , y25775 , y25776 , y25777 , y25778 , y25779 , y25780 , y25781 , y25782 , y25783 , y25784 , y25785 , y25786 , y25787 , y25788 , y25789 , y25790 , y25791 , y25792 , y25793 , y25794 , y25795 , y25796 , y25797 , y25798 , y25799 , y25800 , y25801 , y25802 , y25803 , y25804 , y25805 , y25806 , y25807 , y25808 , y25809 , y25810 , y25811 , y25812 , y25813 , y25814 , y25815 , y25816 , y25817 , y25818 , y25819 , y25820 , y25821 , y25822 , y25823 , y25824 , y25825 , y25826 , y25827 , y25828 , y25829 , y25830 , y25831 , y25832 , y25833 , y25834 , y25835 , y25836 , y25837 , y25838 , y25839 , y25840 , y25841 , y25842 , y25843 , y25844 , y25845 , y25846 , y25847 , y25848 , y25849 , y25850 , y25851 , y25852 , y25853 , y25854 , y25855 , y25856 , y25857 , y25858 , y25859 , y25860 , y25861 , y25862 , y25863 , y25864 , y25865 , y25866 , y25867 , y25868 , y25869 , y25870 , y25871 , y25872 , y25873 , y25874 , y25875 , y25876 , y25877 , y25878 , y25879 , y25880 , y25881 , y25882 , y25883 , y25884 , y25885 , y25886 , y25887 , y25888 , y25889 , y25890 , y25891 , y25892 , y25893 , y25894 , y25895 , y25896 , y25897 , y25898 , y25899 , y25900 , y25901 , y25902 , y25903 , y25904 , y25905 , y25906 , y25907 , y25908 , y25909 , y25910 , y25911 , y25912 , y25913 , y25914 , y25915 , y25916 , y25917 , y25918 , y25919 , y25920 , y25921 , y25922 , y25923 , y25924 , y25925 , y25926 , y25927 , y25928 , y25929 , y25930 , y25931 , y25932 , y25933 , y25934 , y25935 , y25936 , y25937 , y25938 , y25939 , y25940 , y25941 , y25942 , y25943 , y25944 , y25945 , y25946 , y25947 , y25948 , y25949 , y25950 , y25951 , y25952 , y25953 , y25954 , y25955 , y25956 , y25957 , y25958 , y25959 , y25960 , y25961 , y25962 , y25963 , y25964 , y25965 , y25966 , y25967 , y25968 , y25969 , y25970 , y25971 , y25972 , y25973 , y25974 , y25975 , y25976 , y25977 , y25978 , y25979 , y25980 , y25981 , y25982 , y25983 , y25984 , y25985 , y25986 , y25987 , y25988 , y25989 , y25990 , y25991 , y25992 , y25993 , y25994 , y25995 , y25996 , y25997 , y25998 , y25999 , y26000 , y26001 , y26002 , y26003 , y26004 , y26005 , y26006 , y26007 , y26008 , y26009 , y26010 , y26011 , y26012 , y26013 , y26014 , y26015 , y26016 , y26017 , y26018 , y26019 , y26020 , y26021 , y26022 , y26023 , y26024 , y26025 , y26026 , y26027 , y26028 , y26029 , y26030 , y26031 , y26032 , y26033 , y26034 , y26035 , y26036 , y26037 , y26038 , y26039 , y26040 , y26041 , y26042 , y26043 , y26044 , y26045 , y26046 , y26047 , y26048 , y26049 , y26050 , y26051 , y26052 , y26053 , y26054 , y26055 , y26056 , y26057 , y26058 , y26059 , y26060 , y26061 , y26062 , y26063 , y26064 , y26065 , y26066 , y26067 , y26068 , y26069 , y26070 , y26071 , y26072 , y26073 , y26074 , y26075 , y26076 , y26077 , y26078 , y26079 , y26080 , y26081 , y26082 , y26083 , y26084 , y26085 , y26086 , y26087 , y26088 , y26089 , y26090 , y26091 , y26092 , y26093 , y26094 , y26095 , y26096 , y26097 , y26098 , y26099 , y26100 , y26101 , y26102 , y26103 , y26104 , y26105 , y26106 , y26107 , y26108 , y26109 , y26110 , y26111 , y26112 , y26113 , y26114 , y26115 , y26116 , y26117 , y26118 , y26119 , y26120 , y26121 , y26122 , y26123 , y26124 , y26125 , y26126 , y26127 , y26128 , y26129 , y26130 , y26131 , y26132 , y26133 , y26134 , y26135 , y26136 , y26137 , y26138 , y26139 , y26140 , y26141 , y26142 , y26143 , y26144 , y26145 , y26146 , y26147 , y26148 , y26149 , y26150 , y26151 , y26152 , y26153 , y26154 , y26155 , y26156 , y26157 , y26158 , y26159 , y26160 , y26161 , y26162 , y26163 , y26164 , y26165 , y26166 , y26167 , y26168 , y26169 , y26170 , y26171 , y26172 , y26173 , y26174 , y26175 , y26176 , y26177 , y26178 , y26179 , y26180 , y26181 , y26182 , y26183 , y26184 , y26185 , y26186 , y26187 , y26188 , y26189 , y26190 , y26191 , y26192 , y26193 , y26194 , y26195 , y26196 , y26197 , y26198 , y26199 , y26200 , y26201 , y26202 , y26203 , y26204 , y26205 , y26206 , y26207 , y26208 , y26209 , y26210 , y26211 , y26212 , y26213 , y26214 , y26215 , y26216 , y26217 , y26218 , y26219 , y26220 , y26221 , y26222 , y26223 , y26224 , y26225 , y26226 , y26227 , y26228 , y26229 , y26230 , y26231 , y26232 , y26233 , y26234 , y26235 , y26236 , y26237 , y26238 , y26239 , y26240 , y26241 , y26242 , y26243 , y26244 , y26245 , y26246 , y26247 , y26248 , y26249 , y26250 , y26251 , y26252 , y26253 , y26254 , y26255 , y26256 , y26257 , y26258 , y26259 , y26260 , y26261 , y26262 , y26263 , y26264 , y26265 , y26266 , y26267 , y26268 , y26269 , y26270 , y26271 , y26272 , y26273 , y26274 , y26275 , y26276 , y26277 , y26278 , y26279 , y26280 , y26281 , y26282 , y26283 , y26284 , y26285 , y26286 , y26287 , y26288 , y26289 , y26290 , y26291 , y26292 , y26293 , y26294 , y26295 , y26296 , y26297 , y26298 , y26299 , y26300 , y26301 , y26302 , y26303 , y26304 , y26305 , y26306 , y26307 , y26308 , y26309 , y26310 , y26311 , y26312 , y26313 , y26314 , y26315 , y26316 , y26317 , y26318 , y26319 , y26320 , y26321 , y26322 , y26323 , y26324 , y26325 , y26326 , y26327 , y26328 , y26329 , y26330 , y26331 , y26332 , y26333 , y26334 , y26335 , y26336 , y26337 , y26338 , y26339 , y26340 , y26341 , y26342 , y26343 , y26344 , y26345 , y26346 , y26347 , y26348 , y26349 , y26350 , y26351 , y26352 , y26353 , y26354 , y26355 , y26356 , y26357 , y26358 , y26359 , y26360 , y26361 , y26362 , y26363 , y26364 , y26365 , y26366 , y26367 , y26368 , y26369 , y26370 , y26371 , y26372 , y26373 , y26374 , y26375 , y26376 , y26377 , y26378 , y26379 , y26380 , y26381 , y26382 , y26383 , y26384 , y26385 , y26386 , y26387 , y26388 , y26389 , y26390 , y26391 , y26392 , y26393 , y26394 , y26395 , y26396 , y26397 , y26398 , y26399 , y26400 , y26401 , y26402 , y26403 , y26404 , y26405 , y26406 , y26407 , y26408 , y26409 , y26410 , y26411 , y26412 , y26413 , y26414 , y26415 , y26416 , y26417 , y26418 , y26419 , y26420 , y26421 , y26422 , y26423 , y26424 , y26425 , y26426 , y26427 , y26428 , y26429 , y26430 , y26431 , y26432 , y26433 , y26434 , y26435 , y26436 , y26437 , y26438 , y26439 , y26440 , y26441 , y26442 , y26443 , y26444 , y26445 , y26446 , y26447 , y26448 , y26449 , y26450 , y26451 , y26452 , y26453 , y26454 , y26455 , y26456 , y26457 , y26458 , y26459 , y26460 , y26461 , y26462 , y26463 , y26464 , y26465 , y26466 , y26467 , y26468 , y26469 , y26470 , y26471 , y26472 , y26473 , y26474 , y26475 , y26476 , y26477 , y26478 , y26479 , y26480 , y26481 , y26482 , y26483 , y26484 , y26485 , y26486 , y26487 , y26488 , y26489 , y26490 , y26491 , y26492 , y26493 , y26494 , y26495 , y26496 , y26497 , y26498 , y26499 , y26500 , y26501 , y26502 , y26503 , y26504 , y26505 , y26506 , y26507 , y26508 , y26509 , y26510 , y26511 , y26512 , y26513 , y26514 , y26515 , y26516 , y26517 , y26518 , y26519 , y26520 , y26521 , y26522 , y26523 , y26524 , y26525 , y26526 , y26527 , y26528 , y26529 , y26530 , y26531 , y26532 , y26533 , y26534 , y26535 , y26536 , y26537 , y26538 , y26539 , y26540 , y26541 , y26542 , y26543 , y26544 , y26545 , y26546 , y26547 , y26548 , y26549 , y26550 , y26551 , y26552 , y26553 , y26554 , y26555 , y26556 , y26557 , y26558 , y26559 , y26560 , y26561 , y26562 , y26563 , y26564 , y26565 , y26566 , y26567 , y26568 , y26569 , y26570 , y26571 , y26572 , y26573 , y26574 , y26575 , y26576 , y26577 , y26578 , y26579 , y26580 , y26581 , y26582 , y26583 , y26584 , y26585 , y26586 , y26587 , y26588 , y26589 , y26590 , y26591 , y26592 , y26593 , y26594 , y26595 , y26596 , y26597 , y26598 , y26599 , y26600 , y26601 , y26602 , y26603 , y26604 , y26605 , y26606 , y26607 , y26608 , y26609 , y26610 , y26611 , y26612 , y26613 , y26614 , y26615 , y26616 , y26617 , y26618 , y26619 , y26620 , y26621 , y26622 , y26623 , y26624 , y26625 , y26626 , y26627 , y26628 , y26629 , y26630 , y26631 , y26632 , y26633 , y26634 , y26635 , y26636 , y26637 , y26638 , y26639 , y26640 , y26641 , y26642 , y26643 , y26644 , y26645 , y26646 , y26647 , y26648 , y26649 , y26650 , y26651 , y26652 , y26653 , y26654 , y26655 , y26656 , y26657 , y26658 , y26659 , y26660 , y26661 , y26662 , y26663 , y26664 , y26665 , y26666 , y26667 , y26668 , y26669 , y26670 , y26671 , y26672 , y26673 , y26674 , y26675 , y26676 , y26677 , y26678 , y26679 , y26680 , y26681 , y26682 , y26683 , y26684 , y26685 , y26686 , y26687 , y26688 , y26689 , y26690 , y26691 , y26692 , y26693 , y26694 , y26695 , y26696 , y26697 , y26698 , y26699 , y26700 , y26701 , y26702 , y26703 , y26704 , y26705 , y26706 , y26707 , y26708 , y26709 , y26710 , y26711 , y26712 , y26713 , y26714 , y26715 , y26716 , y26717 , y26718 , y26719 , y26720 , y26721 , y26722 , y26723 , y26724 , y26725 , y26726 , y26727 , y26728 , y26729 , y26730 , y26731 , y26732 , y26733 , y26734 , y26735 , y26736 , y26737 , y26738 , y26739 , y26740 , y26741 , y26742 , y26743 , y26744 , y26745 , y26746 , y26747 , y26748 , y26749 , y26750 , y26751 , y26752 , y26753 , y26754 , y26755 , y26756 , y26757 , y26758 , y26759 , y26760 , y26761 , y26762 , y26763 , y26764 , y26765 , y26766 , y26767 , y26768 , y26769 , y26770 , y26771 , y26772 , y26773 , y26774 , y26775 , y26776 , y26777 , y26778 , y26779 , y26780 , y26781 , y26782 , y26783 , y26784 , y26785 , y26786 , y26787 , y26788 , y26789 , y26790 , y26791 , y26792 , y26793 , y26794 , y26795 , y26796 , y26797 , y26798 , y26799 , y26800 , y26801 , y26802 , y26803 , y26804 , y26805 , y26806 , y26807 , y26808 , y26809 , y26810 , y26811 , y26812 , y26813 , y26814 , y26815 , y26816 , y26817 , y26818 , y26819 , y26820 , y26821 , y26822 , y26823 , y26824 , y26825 , y26826 , y26827 , y26828 , y26829 , y26830 , y26831 , y26832 , y26833 , y26834 , y26835 , y26836 , y26837 , y26838 , y26839 , y26840 , y26841 , y26842 , y26843 , y26844 , y26845 , y26846 , y26847 , y26848 , y26849 , y26850 , y26851 , y26852 , y26853 , y26854 , y26855 , y26856 , y26857 , y26858 , y26859 , y26860 , y26861 , y26862 , y26863 , y26864 , y26865 , y26866 , y26867 , y26868 , y26869 , y26870 , y26871 , y26872 , y26873 , y26874 , y26875 , y26876 , y26877 , y26878 , y26879 , y26880 , y26881 , y26882 , y26883 , y26884 , y26885 , y26886 , y26887 , y26888 , y26889 , y26890 , y26891 , y26892 , y26893 , y26894 , y26895 , y26896 , y26897 , y26898 , y26899 , y26900 , y26901 , y26902 , y26903 , y26904 , y26905 , y26906 , y26907 , y26908 , y26909 , y26910 , y26911 , y26912 , y26913 , y26914 , y26915 , y26916 , y26917 , y26918 , y26919 , y26920 , y26921 , y26922 , y26923 , y26924 , y26925 , y26926 , y26927 , y26928 , y26929 , y26930 , y26931 , y26932 , y26933 , y26934 , y26935 , y26936 , y26937 , y26938 , y26939 , y26940 , y26941 , y26942 , y26943 , y26944 , y26945 , y26946 , y26947 , y26948 , y26949 , y26950 , y26951 , y26952 , y26953 , y26954 , y26955 , y26956 , y26957 , y26958 , y26959 , y26960 , y26961 , y26962 , y26963 , y26964 , y26965 , y26966 , y26967 , y26968 , y26969 , y26970 , y26971 , y26972 , y26973 , y26974 , y26975 , y26976 , y26977 , y26978 , y26979 , y26980 , y26981 , y26982 , y26983 , y26984 , y26985 , y26986 , y26987 , y26988 , y26989 , y26990 , y26991 , y26992 , y26993 , y26994 , y26995 , y26996 , y26997 , y26998 , y26999 , y27000 , y27001 , y27002 , y27003 , y27004 , y27005 , y27006 , y27007 , y27008 , y27009 , y27010 , y27011 , y27012 , y27013 , y27014 , y27015 , y27016 , y27017 , y27018 , y27019 , y27020 , y27021 , y27022 , y27023 , y27024 , y27025 , y27026 , y27027 , y27028 , y27029 , y27030 , y27031 , y27032 , y27033 , y27034 , y27035 , y27036 , y27037 , y27038 , y27039 , y27040 , y27041 , y27042 , y27043 , y27044 , y27045 , y27046 , y27047 , y27048 , y27049 , y27050 , y27051 , y27052 , y27053 , y27054 , y27055 , y27056 , y27057 , y27058 , y27059 , y27060 , y27061 , y27062 , y27063 , y27064 , y27065 , y27066 , y27067 , y27068 , y27069 , y27070 , y27071 , y27072 , y27073 , y27074 , y27075 , y27076 , y27077 , y27078 , y27079 , y27080 , y27081 , y27082 , y27083 , y27084 , y27085 , y27086 , y27087 , y27088 , y27089 , y27090 , y27091 , y27092 , y27093 , y27094 , y27095 , y27096 , y27097 , y27098 , y27099 , y27100 , y27101 , y27102 , y27103 , y27104 , y27105 , y27106 , y27107 , y27108 , y27109 , y27110 , y27111 , y27112 , y27113 , y27114 , y27115 , y27116 , y27117 , y27118 , y27119 , y27120 , y27121 , y27122 , y27123 , y27124 , y27125 , y27126 , y27127 , y27128 , y27129 , y27130 , y27131 , y27132 , y27133 , y27134 , y27135 , y27136 , y27137 , y27138 , y27139 , y27140 , y27141 , y27142 , y27143 , y27144 , y27145 , y27146 , y27147 , y27148 , y27149 , y27150 , y27151 , y27152 , y27153 , y27154 , y27155 , y27156 , y27157 , y27158 , y27159 , y27160 , y27161 , y27162 , y27163 , y27164 , y27165 , y27166 , y27167 , y27168 , y27169 , y27170 , y27171 , y27172 , y27173 , y27174 , y27175 , y27176 , y27177 , y27178 , y27179 , y27180 , y27181 , y27182 , y27183 , y27184 , y27185 , y27186 , y27187 , y27188 , y27189 , y27190 , y27191 , y27192 , y27193 , y27194 , y27195 , y27196 , y27197 , y27198 , y27199 , y27200 , y27201 , y27202 , y27203 , y27204 , y27205 , y27206 , y27207 , y27208 , y27209 , y27210 , y27211 , y27212 , y27213 , y27214 , y27215 , y27216 , y27217 , y27218 , y27219 , y27220 , y27221 , y27222 , y27223 , y27224 , y27225 , y27226 , y27227 , y27228 , y27229 , y27230 , y27231 , y27232 , y27233 , y27234 , y27235 , y27236 , y27237 , y27238 , y27239 , y27240 , y27241 , y27242 , y27243 , y27244 , y27245 , y27246 , y27247 , y27248 , y27249 , y27250 , y27251 , y27252 , y27253 , y27254 , y27255 , y27256 , y27257 , y27258 , y27259 , y27260 , y27261 , y27262 , y27263 , y27264 , y27265 , y27266 , y27267 , y27268 , y27269 , y27270 , y27271 , y27272 , y27273 , y27274 , y27275 , y27276 , y27277 , y27278 , y27279 , y27280 , y27281 , y27282 , y27283 , y27284 , y27285 , y27286 , y27287 , y27288 , y27289 , y27290 , y27291 , y27292 , y27293 , y27294 , y27295 , y27296 , y27297 , y27298 , y27299 , y27300 , y27301 , y27302 , y27303 , y27304 , y27305 , y27306 , y27307 , y27308 , y27309 , y27310 , y27311 , y27312 , y27313 , y27314 , y27315 , y27316 , y27317 , y27318 , y27319 , y27320 , y27321 , y27322 , y27323 , y27324 , y27325 , y27326 , y27327 , y27328 , y27329 , y27330 , y27331 , y27332 , y27333 , y27334 , y27335 , y27336 , y27337 , y27338 , y27339 , y27340 , y27341 , y27342 , y27343 , y27344 , y27345 , y27346 , y27347 , y27348 , y27349 , y27350 , y27351 , y27352 , y27353 , y27354 , y27355 , y27356 , y27357 , y27358 , y27359 , y27360 , y27361 , y27362 , y27363 , y27364 , y27365 , y27366 , y27367 , y27368 , y27369 , y27370 , y27371 , y27372 , y27373 , y27374 , y27375 , y27376 , y27377 , y27378 , y27379 , y27380 , y27381 , y27382 , y27383 , y27384 , y27385 , y27386 , y27387 , y27388 , y27389 , y27390 , y27391 , y27392 , y27393 , y27394 , y27395 , y27396 , y27397 , y27398 , y27399 , y27400 , y27401 , y27402 , y27403 , y27404 , y27405 , y27406 , y27407 , y27408 , y27409 , y27410 , y27411 , y27412 , y27413 , y27414 , y27415 , y27416 , y27417 , y27418 , y27419 , y27420 , y27421 , y27422 , y27423 , y27424 , y27425 , y27426 , y27427 , y27428 , y27429 , y27430 , y27431 , y27432 , y27433 , y27434 , y27435 , y27436 , y27437 , y27438 , y27439 , y27440 , y27441 , y27442 , y27443 , y27444 , y27445 , y27446 , y27447 , y27448 , y27449 , y27450 , y27451 , y27452 , y27453 , y27454 , y27455 , y27456 , y27457 , y27458 , y27459 , y27460 , y27461 , y27462 , y27463 , y27464 , y27465 , y27466 , y27467 , y27468 , y27469 , y27470 , y27471 , y27472 , y27473 , y27474 , y27475 , y27476 , y27477 , y27478 , y27479 , y27480 , y27481 , y27482 , y27483 , y27484 , y27485 , y27486 , y27487 , y27488 , y27489 , y27490 , y27491 , y27492 , y27493 , y27494 , y27495 , y27496 , y27497 , y27498 , y27499 , y27500 , y27501 , y27502 , y27503 , y27504 , y27505 , y27506 , y27507 , y27508 , y27509 , y27510 , y27511 , y27512 , y27513 , y27514 , y27515 , y27516 , y27517 , y27518 , y27519 , y27520 , y27521 , y27522 , y27523 , y27524 , y27525 , y27526 , y27527 , y27528 , y27529 , y27530 , y27531 , y27532 , y27533 , y27534 , y27535 , y27536 , y27537 , y27538 , y27539 , y27540 , y27541 , y27542 , y27543 , y27544 , y27545 , y27546 , y27547 , y27548 , y27549 , y27550 , y27551 , y27552 , y27553 , y27554 , y27555 , y27556 , y27557 , y27558 , y27559 , y27560 , y27561 , y27562 , y27563 , y27564 , y27565 , y27566 , y27567 , y27568 , y27569 , y27570 , y27571 , y27572 , y27573 , y27574 , y27575 , y27576 , y27577 , y27578 , y27579 , y27580 , y27581 , y27582 , y27583 , y27584 , y27585 , y27586 , y27587 , y27588 , y27589 , y27590 , y27591 , y27592 , y27593 , y27594 , y27595 , y27596 , y27597 , y27598 , y27599 , y27600 , y27601 , y27602 , y27603 , y27604 , y27605 , y27606 , y27607 , y27608 , y27609 , y27610 , y27611 , y27612 , y27613 , y27614 , y27615 , y27616 , y27617 , y27618 , y27619 , y27620 , y27621 , y27622 , y27623 , y27624 , y27625 , y27626 , y27627 , y27628 , y27629 , y27630 , y27631 , y27632 , y27633 , y27634 , y27635 , y27636 , y27637 , y27638 , y27639 , y27640 , y27641 , y27642 , y27643 , y27644 , y27645 , y27646 , y27647 , y27648 , y27649 , y27650 , y27651 , y27652 , y27653 , y27654 , y27655 , y27656 , y27657 , y27658 , y27659 , y27660 , y27661 , y27662 , y27663 , y27664 , y27665 , y27666 , y27667 , y27668 , y27669 , y27670 , y27671 , y27672 , y27673 , y27674 , y27675 , y27676 , y27677 , y27678 , y27679 , y27680 , y27681 , y27682 , y27683 , y27684 , y27685 , y27686 , y27687 , y27688 , y27689 , y27690 , y27691 , y27692 , y27693 , y27694 , y27695 , y27696 , y27697 , y27698 , y27699 , y27700 , y27701 , y27702 , y27703 , y27704 , y27705 , y27706 , y27707 , y27708 , y27709 , y27710 , y27711 , y27712 , y27713 , y27714 , y27715 , y27716 , y27717 , y27718 , y27719 , y27720 , y27721 , y27722 , y27723 , y27724 , y27725 , y27726 , y27727 , y27728 , y27729 , y27730 , y27731 , y27732 , y27733 , y27734 , y27735 , y27736 , y27737 , y27738 , y27739 , y27740 , y27741 , y27742 , y27743 , y27744 , y27745 , y27746 , y27747 , y27748 , y27749 , y27750 , y27751 , y27752 , y27753 , y27754 , y27755 , y27756 , y27757 , y27758 , y27759 , y27760 , y27761 , y27762 , y27763 , y27764 , y27765 , y27766 , y27767 , y27768 , y27769 , y27770 , y27771 , y27772 , y27773 , y27774 , y27775 , y27776 , y27777 , y27778 , y27779 , y27780 , y27781 , y27782 , y27783 , y27784 , y27785 , y27786 , y27787 , y27788 , y27789 , y27790 , y27791 , y27792 , y27793 , y27794 , y27795 , y27796 , y27797 , y27798 , y27799 , y27800 , y27801 , y27802 , y27803 , y27804 , y27805 , y27806 , y27807 , y27808 , y27809 , y27810 , y27811 , y27812 , y27813 , y27814 , y27815 , y27816 , y27817 , y27818 , y27819 , y27820 , y27821 , y27822 , y27823 , y27824 , y27825 , y27826 , y27827 , y27828 , y27829 , y27830 , y27831 , y27832 , y27833 , y27834 , y27835 , y27836 , y27837 , y27838 , y27839 , y27840 , y27841 , y27842 , y27843 , y27844 , y27845 , y27846 , y27847 , y27848 , y27849 , y27850 , y27851 , y27852 , y27853 , y27854 , y27855 , y27856 , y27857 , y27858 , y27859 , y27860 , y27861 , y27862 , y27863 , y27864 , y27865 , y27866 , y27867 , y27868 , y27869 , y27870 , y27871 , y27872 , y27873 , y27874 , y27875 , y27876 , y27877 , y27878 , y27879 , y27880 , y27881 , y27882 , y27883 , y27884 , y27885 , y27886 , y27887 , y27888 , y27889 , y27890 , y27891 , y27892 , y27893 , y27894 , y27895 , y27896 , y27897 , y27898 , y27899 , y27900 , y27901 , y27902 , y27903 , y27904 , y27905 , y27906 , y27907 , y27908 , y27909 , y27910 , y27911 , y27912 , y27913 , y27914 , y27915 , y27916 , y27917 , y27918 , y27919 , y27920 , y27921 , y27922 , y27923 , y27924 , y27925 , y27926 , y27927 , y27928 , y27929 , y27930 , y27931 , y27932 , y27933 , y27934 , y27935 , y27936 , y27937 , y27938 , y27939 , y27940 , y27941 , y27942 , y27943 , y27944 , y27945 , y27946 , y27947 , y27948 , y27949 , y27950 , y27951 , y27952 , y27953 , y27954 , y27955 , y27956 , y27957 , y27958 , y27959 , y27960 , y27961 , y27962 , y27963 , y27964 , y27965 , y27966 , y27967 , y27968 , y27969 , y27970 , y27971 , y27972 , y27973 , y27974 , y27975 , y27976 , y27977 , y27978 , y27979 , y27980 , y27981 , y27982 , y27983 , y27984 , y27985 , y27986 , y27987 , y27988 , y27989 , y27990 , y27991 , y27992 , y27993 , y27994 , y27995 , y27996 , y27997 , y27998 , y27999 , y28000 , y28001 , y28002 , y28003 , y28004 , y28005 , y28006 , y28007 , y28008 , y28009 , y28010 , y28011 , y28012 , y28013 , y28014 , y28015 , y28016 , y28017 , y28018 , y28019 , y28020 , y28021 , y28022 , y28023 , y28024 , y28025 , y28026 , y28027 , y28028 , y28029 , y28030 , y28031 , y28032 , y28033 , y28034 , y28035 , y28036 , y28037 , y28038 , y28039 , y28040 , y28041 , y28042 , y28043 , y28044 , y28045 , y28046 , y28047 , y28048 , y28049 , y28050 , y28051 , y28052 , y28053 , y28054 , y28055 , y28056 , y28057 , y28058 , y28059 , y28060 , y28061 , y28062 , y28063 , y28064 , y28065 , y28066 , y28067 , y28068 , y28069 , y28070 , y28071 , y28072 , y28073 , y28074 , y28075 , y28076 , y28077 , y28078 , y28079 , y28080 , y28081 , y28082 , y28083 , y28084 , y28085 , y28086 , y28087 , y28088 , y28089 , y28090 , y28091 , y28092 , y28093 , y28094 , y28095 , y28096 , y28097 , y28098 , y28099 , y28100 , y28101 , y28102 , y28103 , y28104 , y28105 , y28106 , y28107 , y28108 , y28109 , y28110 , y28111 , y28112 , y28113 , y28114 , y28115 , y28116 , y28117 , y28118 , y28119 , y28120 , y28121 , y28122 , y28123 , y28124 , y28125 , y28126 , y28127 , y28128 , y28129 , y28130 , y28131 , y28132 , y28133 , y28134 , y28135 , y28136 , y28137 , y28138 , y28139 , y28140 , y28141 , y28142 , y28143 , y28144 , y28145 , y28146 , y28147 , y28148 , y28149 , y28150 , y28151 , y28152 , y28153 , y28154 , y28155 , y28156 , y28157 , y28158 , y28159 , y28160 , y28161 , y28162 , y28163 , y28164 , y28165 , y28166 , y28167 , y28168 , y28169 , y28170 , y28171 , y28172 , y28173 , y28174 , y28175 , y28176 , y28177 , y28178 , y28179 , y28180 , y28181 , y28182 , y28183 , y28184 , y28185 , y28186 , y28187 , y28188 , y28189 , y28190 , y28191 , y28192 , y28193 , y28194 , y28195 , y28196 , y28197 , y28198 , y28199 , y28200 , y28201 , y28202 , y28203 , y28204 , y28205 , y28206 , y28207 , y28208 , y28209 , y28210 , y28211 , y28212 , y28213 , y28214 , y28215 , y28216 , y28217 , y28218 , y28219 , y28220 , y28221 , y28222 , y28223 , y28224 , y28225 , y28226 , y28227 , y28228 , y28229 , y28230 , y28231 , y28232 , y28233 , y28234 , y28235 , y28236 , y28237 , y28238 , y28239 , y28240 , y28241 , y28242 , y28243 , y28244 , y28245 , y28246 , y28247 , y28248 , y28249 , y28250 , y28251 , y28252 , y28253 , y28254 , y28255 , y28256 , y28257 , y28258 , y28259 , y28260 , y28261 , y28262 , y28263 , y28264 , y28265 , y28266 , y28267 , y28268 , y28269 , y28270 , y28271 , y28272 , y28273 , y28274 , y28275 , y28276 , y28277 , y28278 , y28279 , y28280 , y28281 , y28282 , y28283 , y28284 , y28285 , y28286 , y28287 , y28288 , y28289 , y28290 , y28291 , y28292 , y28293 , y28294 , y28295 , y28296 , y28297 , y28298 , y28299 , y28300 , y28301 , y28302 , y28303 , y28304 , y28305 , y28306 , y28307 , y28308 , y28309 , y28310 , y28311 , y28312 , y28313 , y28314 , y28315 , y28316 , y28317 , y28318 , y28319 , y28320 , y28321 , y28322 , y28323 , y28324 , y28325 , y28326 , y28327 , y28328 , y28329 , y28330 , y28331 , y28332 , y28333 , y28334 , y28335 , y28336 , y28337 , y28338 , y28339 , y28340 , y28341 , y28342 , y28343 , y28344 , y28345 , y28346 , y28347 , y28348 , y28349 , y28350 , y28351 , y28352 , y28353 , y28354 , y28355 , y28356 , y28357 , y28358 , y28359 , y28360 , y28361 , y28362 , y28363 , y28364 , y28365 , y28366 , y28367 , y28368 , y28369 , y28370 , y28371 , y28372 , y28373 , y28374 , y28375 , y28376 , y28377 , y28378 , y28379 , y28380 , y28381 , y28382 , y28383 , y28384 , y28385 , y28386 , y28387 , y28388 , y28389 , y28390 , y28391 , y28392 , y28393 , y28394 , y28395 , y28396 , y28397 , y28398 , y28399 , y28400 , y28401 , y28402 , y28403 , y28404 , y28405 , y28406 , y28407 , y28408 , y28409 , y28410 , y28411 , y28412 , y28413 , y28414 , y28415 , y28416 , y28417 , y28418 , y28419 , y28420 , y28421 , y28422 , y28423 , y28424 , y28425 , y28426 , y28427 , y28428 , y28429 , y28430 , y28431 , y28432 , y28433 , y28434 , y28435 , y28436 , y28437 , y28438 , y28439 , y28440 , y28441 , y28442 , y28443 , y28444 , y28445 , y28446 , y28447 , y28448 , y28449 , y28450 , y28451 , y28452 , y28453 , y28454 , y28455 , y28456 , y28457 , y28458 , y28459 , y28460 , y28461 , y28462 , y28463 , y28464 , y28465 , y28466 , y28467 , y28468 , y28469 , y28470 , y28471 , y28472 , y28473 , y28474 , y28475 , y28476 , y28477 , y28478 , y28479 , y28480 , y28481 , y28482 , y28483 , y28484 , y28485 , y28486 , y28487 , y28488 , y28489 , y28490 , y28491 , y28492 , y28493 , y28494 , y28495 , y28496 , y28497 , y28498 , y28499 , y28500 , y28501 , y28502 , y28503 , y28504 , y28505 , y28506 , y28507 , y28508 , y28509 , y28510 , y28511 , y28512 , y28513 , y28514 , y28515 , y28516 , y28517 , y28518 , y28519 , y28520 , y28521 , y28522 , y28523 , y28524 , y28525 , y28526 , y28527 , y28528 , y28529 , y28530 , y28531 , y28532 , y28533 , y28534 , y28535 , y28536 , y28537 , y28538 , y28539 , y28540 , y28541 , y28542 , y28543 , y28544 , y28545 , y28546 , y28547 , y28548 , y28549 , y28550 , y28551 , y28552 , y28553 , y28554 , y28555 , y28556 , y28557 , y28558 , y28559 , y28560 , y28561 , y28562 , y28563 , y28564 , y28565 , y28566 , y28567 , y28568 , y28569 , y28570 , y28571 , y28572 , y28573 , y28574 , y28575 , y28576 , y28577 , y28578 , y28579 , y28580 , y28581 , y28582 , y28583 , y28584 , y28585 , y28586 , y28587 , y28588 , y28589 , y28590 , y28591 , y28592 , y28593 , y28594 , y28595 , y28596 , y28597 , y28598 , y28599 , y28600 , y28601 , y28602 , y28603 , y28604 , y28605 , y28606 , y28607 , y28608 , y28609 , y28610 , y28611 , y28612 , y28613 , y28614 , y28615 , y28616 , y28617 , y28618 , y28619 , y28620 , y28621 , y28622 , y28623 , y28624 , y28625 , y28626 , y28627 , y28628 , y28629 , y28630 , y28631 , y28632 , y28633 , y28634 , y28635 , y28636 , y28637 , y28638 , y28639 , y28640 , y28641 , y28642 , y28643 , y28644 , y28645 , y28646 , y28647 , y28648 , y28649 , y28650 , y28651 , y28652 , y28653 , y28654 , y28655 , y28656 , y28657 , y28658 , y28659 , y28660 , y28661 , y28662 , y28663 , y28664 , y28665 , y28666 , y28667 , y28668 , y28669 , y28670 , y28671 , y28672 , y28673 , y28674 , y28675 , y28676 , y28677 , y28678 , y28679 , y28680 , y28681 , y28682 , y28683 , y28684 , y28685 , y28686 , y28687 , y28688 , y28689 , y28690 , y28691 , y28692 , y28693 , y28694 , y28695 , y28696 , y28697 , y28698 , y28699 , y28700 , y28701 , y28702 , y28703 , y28704 , y28705 , y28706 , y28707 , y28708 , y28709 , y28710 , y28711 , y28712 , y28713 , y28714 , y28715 , y28716 , y28717 , y28718 , y28719 , y28720 , y28721 , y28722 , y28723 , y28724 , y28725 , y28726 , y28727 , y28728 , y28729 , y28730 , y28731 , y28732 , y28733 , y28734 , y28735 , y28736 , y28737 , y28738 , y28739 , y28740 , y28741 , y28742 , y28743 , y28744 , y28745 , y28746 , y28747 , y28748 , y28749 , y28750 , y28751 , y28752 , y28753 , y28754 , y28755 , y28756 , y28757 , y28758 , y28759 , y28760 , y28761 , y28762 , y28763 , y28764 , y28765 , y28766 , y28767 , y28768 , y28769 , y28770 , y28771 , y28772 , y28773 , y28774 , y28775 , y28776 , y28777 , y28778 , y28779 , y28780 , y28781 , y28782 , y28783 , y28784 , y28785 , y28786 , y28787 , y28788 , y28789 , y28790 , y28791 , y28792 , y28793 , y28794 , y28795 , y28796 , y28797 , y28798 , y28799 , y28800 , y28801 , y28802 , y28803 , y28804 , y28805 , y28806 , y28807 , y28808 , y28809 , y28810 , y28811 , y28812 , y28813 , y28814 , y28815 , y28816 , y28817 , y28818 , y28819 , y28820 , y28821 , y28822 , y28823 , y28824 , y28825 , y28826 , y28827 , y28828 , y28829 , y28830 , y28831 , y28832 , y28833 , y28834 , y28835 , y28836 , y28837 , y28838 , y28839 , y28840 , y28841 , y28842 , y28843 , y28844 , y28845 , y28846 , y28847 , y28848 , y28849 , y28850 , y28851 , y28852 , y28853 , y28854 , y28855 , y28856 , y28857 , y28858 , y28859 , y28860 , y28861 , y28862 , y28863 , y28864 , y28865 , y28866 , y28867 , y28868 , y28869 , y28870 , y28871 , y28872 , y28873 , y28874 , y28875 , y28876 , y28877 , y28878 , y28879 , y28880 , y28881 , y28882 , y28883 , y28884 , y28885 , y28886 , y28887 , y28888 , y28889 , y28890 , y28891 , y28892 , y28893 , y28894 , y28895 , y28896 , y28897 , y28898 , y28899 , y28900 , y28901 , y28902 , y28903 , y28904 , y28905 , y28906 , y28907 , y28908 , y28909 , y28910 , y28911 , y28912 , y28913 , y28914 , y28915 , y28916 , y28917 , y28918 , y28919 , y28920 , y28921 , y28922 , y28923 , y28924 , y28925 , y28926 , y28927 , y28928 , y28929 , y28930 , y28931 , y28932 , y28933 , y28934 , y28935 , y28936 , y28937 , y28938 , y28939 , y28940 , y28941 , y28942 , y28943 , y28944 , y28945 , y28946 , y28947 , y28948 , y28949 , y28950 , y28951 , y28952 , y28953 , y28954 , y28955 , y28956 , y28957 , y28958 , y28959 , y28960 , y28961 , y28962 , y28963 , y28964 , y28965 , y28966 , y28967 , y28968 , y28969 , y28970 , y28971 , y28972 , y28973 , y28974 , y28975 , y28976 , y28977 , y28978 , y28979 , y28980 , y28981 , y28982 , y28983 , y28984 , y28985 , y28986 , y28987 , y28988 , y28989 , y28990 , y28991 , y28992 , y28993 , y28994 , y28995 , y28996 , y28997 , y28998 , y28999 , y29000 , y29001 , y29002 , y29003 , y29004 , y29005 , y29006 , y29007 , y29008 , y29009 , y29010 , y29011 , y29012 , y29013 , y29014 , y29015 , y29016 , y29017 , y29018 , y29019 , y29020 , y29021 , y29022 , y29023 , y29024 , y29025 , y29026 , y29027 , y29028 , y29029 , y29030 , y29031 , y29032 , y29033 , y29034 , y29035 , y29036 , y29037 , y29038 , y29039 , y29040 , y29041 , y29042 , y29043 , y29044 , y29045 , y29046 , y29047 , y29048 , y29049 , y29050 , y29051 , y29052 , y29053 , y29054 , y29055 , y29056 , y29057 , y29058 , y29059 , y29060 , y29061 , y29062 , y29063 , y29064 , y29065 , y29066 , y29067 , y29068 , y29069 , y29070 , y29071 , y29072 , y29073 , y29074 , y29075 , y29076 , y29077 , y29078 , y29079 , y29080 , y29081 , y29082 , y29083 , y29084 , y29085 , y29086 , y29087 , y29088 , y29089 , y29090 , y29091 , y29092 , y29093 , y29094 , y29095 , y29096 , y29097 , y29098 , y29099 , y29100 , y29101 , y29102 , y29103 , y29104 , y29105 , y29106 , y29107 , y29108 , y29109 , y29110 , y29111 , y29112 , y29113 , y29114 , y29115 , y29116 , y29117 , y29118 , y29119 , y29120 , y29121 , y29122 , y29123 , y29124 , y29125 , y29126 , y29127 , y29128 , y29129 , y29130 , y29131 , y29132 , y29133 , y29134 , y29135 , y29136 , y29137 , y29138 , y29139 , y29140 , y29141 , y29142 , y29143 , y29144 , y29145 , y29146 , y29147 , y29148 , y29149 , y29150 , y29151 , y29152 , y29153 , y29154 , y29155 , y29156 , y29157 , y29158 , y29159 , y29160 , y29161 , y29162 , y29163 , y29164 , y29165 , y29166 , y29167 , y29168 , y29169 , y29170 , y29171 , y29172 , y29173 , y29174 , y29175 , y29176 , y29177 , y29178 , y29179 , y29180 , y29181 , y29182 , y29183 , y29184 , y29185 , y29186 , y29187 , y29188 , y29189 , y29190 , y29191 , y29192 , y29193 , y29194 , y29195 , y29196 , y29197 , y29198 , y29199 , y29200 , y29201 , y29202 , y29203 , y29204 , y29205 , y29206 , y29207 , y29208 , y29209 , y29210 , y29211 , y29212 , y29213 , y29214 , y29215 , y29216 , y29217 , y29218 , y29219 , y29220 , y29221 , y29222 , y29223 , y29224 , y29225 , y29226 , y29227 , y29228 , y29229 , y29230 , y29231 , y29232 , y29233 , y29234 , y29235 , y29236 , y29237 , y29238 , y29239 , y29240 , y29241 , y29242 , y29243 , y29244 , y29245 , y29246 , y29247 , y29248 , y29249 , y29250 , y29251 , y29252 , y29253 , y29254 , y29255 , y29256 , y29257 , y29258 , y29259 , y29260 , y29261 , y29262 , y29263 , y29264 , y29265 , y29266 , y29267 , y29268 , y29269 , y29270 , y29271 , y29272 , y29273 , y29274 , y29275 , y29276 , y29277 , y29278 , y29279 , y29280 , y29281 , y29282 , y29283 , y29284 , y29285 , y29286 , y29287 , y29288 , y29289 , y29290 , y29291 , y29292 , y29293 , y29294 , y29295 , y29296 , y29297 , y29298 , y29299 , y29300 , y29301 , y29302 , y29303 , y29304 , y29305 , y29306 , y29307 , y29308 , y29309 , y29310 , y29311 , y29312 , y29313 , y29314 , y29315 , y29316 , y29317 , y29318 , y29319 , y29320 , y29321 , y29322 , y29323 , y29324 , y29325 , y29326 , y29327 , y29328 , y29329 , y29330 , y29331 , y29332 , y29333 , y29334 , y29335 , y29336 , y29337 , y29338 , y29339 , y29340 , y29341 , y29342 , y29343 , y29344 , y29345 , y29346 , y29347 , y29348 , y29349 , y29350 , y29351 , y29352 , y29353 , y29354 , y29355 , y29356 , y29357 , y29358 , y29359 , y29360 , y29361 , y29362 , y29363 , y29364 , y29365 , y29366 , y29367 , y29368 , y29369 , y29370 , y29371 , y29372 , y29373 , y29374 , y29375 , y29376 , y29377 , y29378 , y29379 , y29380 , y29381 , y29382 , y29383 , y29384 , y29385 , y29386 , y29387 , y29388 , y29389 , y29390 , y29391 , y29392 , y29393 , y29394 , y29395 , y29396 , y29397 , y29398 , y29399 , y29400 , y29401 , y29402 , y29403 , y29404 , y29405 , y29406 , y29407 , y29408 , y29409 , y29410 , y29411 , y29412 , y29413 , y29414 , y29415 , y29416 , y29417 , y29418 , y29419 , y29420 , y29421 , y29422 , y29423 , y29424 , y29425 , y29426 , y29427 , y29428 , y29429 , y29430 , y29431 , y29432 , y29433 , y29434 , y29435 , y29436 , y29437 , y29438 , y29439 , y29440 , y29441 , y29442 , y29443 , y29444 , y29445 , y29446 , y29447 , y29448 , y29449 , y29450 , y29451 , y29452 , y29453 , y29454 , y29455 , y29456 , y29457 , y29458 , y29459 , y29460 , y29461 , y29462 , y29463 , y29464 , y29465 , y29466 , y29467 , y29468 , y29469 , y29470 , y29471 , y29472 , y29473 , y29474 , y29475 , y29476 , y29477 , y29478 , y29479 , y29480 , y29481 , y29482 , y29483 , y29484 , y29485 , y29486 , y29487 , y29488 , y29489 , y29490 , y29491 , y29492 , y29493 , y29494 , y29495 , y29496 , y29497 , y29498 , y29499 , y29500 , y29501 , y29502 , y29503 , y29504 , y29505 , y29506 , y29507 , y29508 , y29509 , y29510 , y29511 , y29512 , y29513 , y29514 , y29515 , y29516 , y29517 , y29518 , y29519 , y29520 , y29521 , y29522 , y29523 , y29524 , y29525 , y29526 , y29527 , y29528 , y29529 , y29530 , y29531 , y29532 , y29533 , y29534 , y29535 , y29536 , y29537 , y29538 , y29539 , y29540 , y29541 , y29542 , y29543 , y29544 , y29545 , y29546 , y29547 , y29548 , y29549 , y29550 , y29551 , y29552 , y29553 , y29554 , y29555 , y29556 , y29557 , y29558 , y29559 , y29560 , y29561 , y29562 , y29563 , y29564 , y29565 , y29566 , y29567 , y29568 , y29569 , y29570 , y29571 , y29572 , y29573 , y29574 , y29575 , y29576 , y29577 , y29578 , y29579 , y29580 , y29581 , y29582 , y29583 , y29584 , y29585 , y29586 , y29587 , y29588 , y29589 , y29590 , y29591 , y29592 , y29593 , y29594 , y29595 , y29596 , y29597 , y29598 , y29599 , y29600 , y29601 , y29602 , y29603 , y29604 , y29605 , y29606 , y29607 , y29608 , y29609 , y29610 , y29611 , y29612 , y29613 , y29614 , y29615 , y29616 , y29617 , y29618 , y29619 , y29620 , y29621 , y29622 , y29623 , y29624 , y29625 , y29626 , y29627 , y29628 , y29629 , y29630 , y29631 , y29632 , y29633 , y29634 , y29635 , y29636 , y29637 , y29638 , y29639 , y29640 , y29641 , y29642 , y29643 , y29644 , y29645 , y29646 , y29647 , y29648 , y29649 , y29650 , y29651 , y29652 , y29653 , y29654 , y29655 , y29656 , y29657 , y29658 , y29659 , y29660 , y29661 , y29662 , y29663 , y29664 , y29665 , y29666 , y29667 , y29668 , y29669 , y29670 , y29671 , y29672 , y29673 , y29674 , y29675 , y29676 , y29677 , y29678 , y29679 , y29680 , y29681 , y29682 , y29683 , y29684 , y29685 , y29686 , y29687 , y29688 , y29689 , y29690 , y29691 , y29692 , y29693 , y29694 , y29695 , y29696 , y29697 , y29698 , y29699 , y29700 , y29701 , y29702 , y29703 , y29704 , y29705 , y29706 , y29707 , y29708 , y29709 , y29710 , y29711 , y29712 , y29713 , y29714 , y29715 , y29716 , y29717 , y29718 , y29719 , y29720 , y29721 , y29722 , y29723 , y29724 , y29725 , y29726 , y29727 , y29728 , y29729 , y29730 , y29731 , y29732 , y29733 , y29734 , y29735 , y29736 , y29737 , y29738 , y29739 , y29740 , y29741 , y29742 , y29743 , y29744 , y29745 , y29746 , y29747 , y29748 , y29749 , y29750 , y29751 , y29752 , y29753 , y29754 , y29755 , y29756 , y29757 , y29758 , y29759 , y29760 , y29761 , y29762 , y29763 , y29764 , y29765 , y29766 , y29767 , y29768 , y29769 , y29770 , y29771 , y29772 , y29773 , y29774 , y29775 , y29776 , y29777 , y29778 , y29779 , y29780 , y29781 , y29782 , y29783 , y29784 , y29785 , y29786 , y29787 , y29788 , y29789 , y29790 , y29791 , y29792 , y29793 , y29794 , y29795 , y29796 , y29797 , y29798 , y29799 , y29800 , y29801 , y29802 , y29803 , y29804 , y29805 , y29806 , y29807 , y29808 , y29809 , y29810 , y29811 , y29812 , y29813 , y29814 , y29815 , y29816 , y29817 , y29818 , y29819 , y29820 , y29821 , y29822 , y29823 , y29824 , y29825 , y29826 , y29827 , y29828 , y29829 , y29830 , y29831 , y29832 , y29833 , y29834 , y29835 , y29836 , y29837 , y29838 , y29839 , y29840 , y29841 , y29842 , y29843 , y29844 , y29845 , y29846 , y29847 , y29848 , y29849 , y29850 , y29851 , y29852 , y29853 , y29854 , y29855 , y29856 , y29857 , y29858 , y29859 , y29860 , y29861 , y29862 , y29863 , y29864 , y29865 , y29866 , y29867 , y29868 , y29869 , y29870 , y29871 , y29872 , y29873 , y29874 , y29875 , y29876 , y29877 , y29878 , y29879 , y29880 , y29881 , y29882 , y29883 , y29884 , y29885 , y29886 , y29887 , y29888 , y29889 , y29890 , y29891 , y29892 , y29893 , y29894 , y29895 , y29896 , y29897 , y29898 , y29899 , y29900 , y29901 , y29902 , y29903 , y29904 , y29905 , y29906 , y29907 , y29908 , y29909 , y29910 , y29911 , y29912 , y29913 , y29914 , y29915 , y29916 , y29917 , y29918 , y29919 , y29920 , y29921 , y29922 , y29923 , y29924 , y29925 , y29926 , y29927 , y29928 , y29929 , y29930 , y29931 , y29932 , y29933 , y29934 , y29935 , y29936 , y29937 , y29938 , y29939 , y29940 , y29941 , y29942 , y29943 , y29944 , y29945 , y29946 , y29947 , y29948 , y29949 , y29950 , y29951 , y29952 , y29953 , y29954 , y29955 , y29956 , y29957 , y29958 , y29959 , y29960 , y29961 , y29962 , y29963 , y29964 , y29965 , y29966 , y29967 , y29968 , y29969 , y29970 , y29971 , y29972 , y29973 , y29974 , y29975 , y29976 , y29977 , y29978 , y29979 , y29980 , y29981 , y29982 , y29983 , y29984 , y29985 , y29986 , y29987 , y29988 , y29989 , y29990 , y29991 , y29992 , y29993 , y29994 , y29995 , y29996 , y29997 , y29998 , y29999 , y30000 , y30001 , y30002 , y30003 , y30004 , y30005 , y30006 , y30007 , y30008 , y30009 , y30010 , y30011 , y30012 , y30013 , y30014 , y30015 , y30016 , y30017 , y30018 , y30019 , y30020 , y30021 , y30022 , y30023 , y30024 , y30025 , y30026 , y30027 , y30028 , y30029 , y30030 , y30031 , y30032 , y30033 , y30034 , y30035 , y30036 , y30037 , y30038 , y30039 , y30040 , y30041 , y30042 , y30043 , y30044 , y30045 , y30046 , y30047 , y30048 , y30049 , y30050 , y30051 , y30052 , y30053 , y30054 , y30055 , y30056 , y30057 , y30058 , y30059 , y30060 , y30061 , y30062 , y30063 , y30064 , y30065 , y30066 , y30067 , y30068 , y30069 , y30070 , y30071 , y30072 , y30073 , y30074 , y30075 , y30076 , y30077 , y30078 , y30079 , y30080 , y30081 , y30082 , y30083 , y30084 , y30085 , y30086 , y30087 , y30088 , y30089 , y30090 , y30091 , y30092 , y30093 , y30094 , y30095 , y30096 , y30097 , y30098 , y30099 , y30100 , y30101 , y30102 , y30103 , y30104 , y30105 , y30106 , y30107 , y30108 , y30109 , y30110 , y30111 , y30112 , y30113 , y30114 , y30115 , y30116 , y30117 , y30118 , y30119 , y30120 , y30121 , y30122 , y30123 , y30124 , y30125 , y30126 , y30127 , y30128 , y30129 , y30130 , y30131 , y30132 , y30133 , y30134 , y30135 , y30136 , y30137 , y30138 , y30139 , y30140 , y30141 , y30142 , y30143 , y30144 , y30145 , y30146 , y30147 , y30148 , y30149 , y30150 , y30151 , y30152 , y30153 , y30154 , y30155 , y30156 , y30157 , y30158 , y30159 , y30160 , y30161 , y30162 , y30163 , y30164 , y30165 , y30166 , y30167 , y30168 , y30169 , y30170 , y30171 , y30172 , y30173 , y30174 , y30175 , y30176 , y30177 , y30178 , y30179 , y30180 , y30181 , y30182 , y30183 , y30184 , y30185 , y30186 , y30187 , y30188 , y30189 , y30190 , y30191 , y30192 , y30193 , y30194 , y30195 , y30196 , y30197 , y30198 , y30199 , y30200 , y30201 , y30202 , y30203 , y30204 , y30205 , y30206 , y30207 , y30208 , y30209 , y30210 , y30211 , y30212 , y30213 , y30214 , y30215 , y30216 , y30217 , y30218 , y30219 , y30220 , y30221 , y30222 , y30223 , y30224 , y30225 , y30226 , y30227 , y30228 , y30229 , y30230 , y30231 , y30232 , y30233 , y30234 , y30235 , y30236 , y30237 , y30238 , y30239 , y30240 , y30241 , y30242 , y30243 , y30244 , y30245 , y30246 , y30247 , y30248 , y30249 , y30250 , y30251 , y30252 , y30253 , y30254 , y30255 , y30256 , y30257 , y30258 , y30259 , y30260 , y30261 , y30262 , y30263 , y30264 , y30265 , y30266 , y30267 , y30268 , y30269 , y30270 , y30271 , y30272 , y30273 , y30274 , y30275 , y30276 , y30277 , y30278 , y30279 , y30280 , y30281 , y30282 , y30283 , y30284 , y30285 , y30286 , y30287 , y30288 , y30289 , y30290 , y30291 , y30292 , y30293 , y30294 , y30295 , y30296 , y30297 , y30298 , y30299 , y30300 , y30301 , y30302 , y30303 , y30304 , y30305 , y30306 , y30307 , y30308 , y30309 , y30310 , y30311 , y30312 , y30313 , y30314 , y30315 , y30316 , y30317 , y30318 , y30319 , y30320 , y30321 , y30322 , y30323 , y30324 , y30325 , y30326 , y30327 , y30328 , y30329 , y30330 , y30331 , y30332 , y30333 , y30334 , y30335 , y30336 , y30337 , y30338 , y30339 , y30340 , y30341 , y30342 , y30343 , y30344 , y30345 , y30346 , y30347 , y30348 , y30349 , y30350 , y30351 , y30352 , y30353 , y30354 , y30355 , y30356 , y30357 , y30358 , y30359 , y30360 , y30361 , y30362 , y30363 , y30364 , y30365 , y30366 , y30367 , y30368 , y30369 , y30370 , y30371 , y30372 , y30373 , y30374 , y30375 , y30376 , y30377 , y30378 , y30379 , y30380 , y30381 , y30382 , y30383 , y30384 , y30385 , y30386 , y30387 , y30388 , y30389 , y30390 , y30391 , y30392 , y30393 , y30394 , y30395 , y30396 , y30397 , y30398 , y30399 , y30400 , y30401 , y30402 , y30403 , y30404 , y30405 , y30406 , y30407 , y30408 , y30409 , y30410 , y30411 , y30412 , y30413 , y30414 , y30415 , y30416 , y30417 , y30418 , y30419 , y30420 , y30421 , y30422 , y30423 , y30424 , y30425 , y30426 , y30427 , y30428 , y30429 , y30430 , y30431 , y30432 , y30433 , y30434 , y30435 , y30436 , y30437 , y30438 , y30439 , y30440 , y30441 , y30442 , y30443 , y30444 , y30445 , y30446 , y30447 , y30448 , y30449 , y30450 , y30451 , y30452 , y30453 , y30454 , y30455 , y30456 , y30457 , y30458 , y30459 , y30460 , y30461 , y30462 , y30463 , y30464 , y30465 , y30466 , y30467 , y30468 , y30469 , y30470 , y30471 , y30472 , y30473 , y30474 , y30475 , y30476 , y30477 , y30478 , y30479 , y30480 , y30481 , y30482 , y30483 , y30484 , y30485 , y30486 , y30487 , y30488 , y30489 , y30490 , y30491 , y30492 , y30493 , y30494 , y30495 , y30496 , y30497 , y30498 , y30499 , y30500 , y30501 , y30502 , y30503 , y30504 , y30505 , y30506 , y30507 , y30508 , y30509 , y30510 , y30511 , y30512 , y30513 , y30514 , y30515 , y30516 , y30517 , y30518 , y30519 , y30520 , y30521 , y30522 , y30523 , y30524 , y30525 , y30526 , y30527 , y30528 , y30529 , y30530 , y30531 , y30532 , y30533 , y30534 , y30535 , y30536 , y30537 , y30538 , y30539 , y30540 , y30541 , y30542 , y30543 , y30544 , y30545 , y30546 , y30547 , y30548 , y30549 , y30550 , y30551 , y30552 , y30553 , y30554 , y30555 , y30556 , y30557 , y30558 , y30559 , y30560 , y30561 , y30562 , y30563 , y30564 , y30565 , y30566 , y30567 , y30568 , y30569 , y30570 , y30571 , y30572 , y30573 , y30574 , y30575 , y30576 , y30577 , y30578 , y30579 , y30580 , y30581 , y30582 , y30583 , y30584 , y30585 , y30586 , y30587 , y30588 , y30589 , y30590 , y30591 , y30592 , y30593 , y30594 , y30595 , y30596 , y30597 , y30598 , y30599 , y30600 , y30601 , y30602 , y30603 , y30604 , y30605 , y30606 , y30607 , y30608 , y30609 , y30610 , y30611 , y30612 , y30613 , y30614 , y30615 , y30616 , y30617 , y30618 , y30619 , y30620 , y30621 , y30622 , y30623 , y30624 , y30625 , y30626 , y30627 , y30628 , y30629 , y30630 , y30631 , y30632 , y30633 , y30634 , y30635 , y30636 , y30637 , y30638 , y30639 , y30640 , y30641 , y30642 , y30643 , y30644 , y30645 , y30646 , y30647 , y30648 , y30649 , y30650 , y30651 , y30652 , y30653 , y30654 , y30655 , y30656 , y30657 , y30658 , y30659 , y30660 , y30661 , y30662 , y30663 , y30664 , y30665 , y30666 , y30667 , y30668 , y30669 , y30670 , y30671 , y30672 , y30673 , y30674 , y30675 , y30676 , y30677 , y30678 , y30679 , y30680 , y30681 , y30682 , y30683 , y30684 , y30685 , y30686 , y30687 , y30688 , y30689 , y30690 , y30691 , y30692 , y30693 , y30694 , y30695 , y30696 , y30697 , y30698 , y30699 , y30700 , y30701 , y30702 , y30703 , y30704 , y30705 , y30706 , y30707 , y30708 , y30709 , y30710 , y30711 , y30712 , y30713 , y30714 , y30715 , y30716 , y30717 , y30718 , y30719 , y30720 , y30721 , y30722 , y30723 , y30724 , y30725 , y30726 , y30727 , y30728 , y30729 , y30730 , y30731 , y30732 , y30733 , y30734 , y30735 , y30736 , y30737 , y30738 , y30739 , y30740 , y30741 , y30742 , y30743 , y30744 , y30745 , y30746 , y30747 , y30748 , y30749 , y30750 , y30751 , y30752 , y30753 , y30754 , y30755 , y30756 , y30757 , y30758 , y30759 , y30760 , y30761 , y30762 , y30763 , y30764 , y30765 , y30766 , y30767 , y30768 , y30769 , y30770 , y30771 , y30772 , y30773 , y30774 , y30775 , y30776 , y30777 , y30778 , y30779 , y30780 , y30781 , y30782 , y30783 , y30784 , y30785 , y30786 , y30787 , y30788 , y30789 , y30790 , y30791 , y30792 , y30793 , y30794 , y30795 , y30796 , y30797 , y30798 , y30799 , y30800 , y30801 , y30802 , y30803 , y30804 , y30805 , y30806 , y30807 , y30808 , y30809 , y30810 , y30811 , y30812 , y30813 , y30814 , y30815 , y30816 , y30817 , y30818 , y30819 , y30820 , y30821 , y30822 , y30823 , y30824 , y30825 , y30826 , y30827 , y30828 , y30829 , y30830 , y30831 , y30832 , y30833 , y30834 , y30835 , y30836 , y30837 , y30838 , y30839 , y30840 , y30841 , y30842 , y30843 , y30844 , y30845 , y30846 , y30847 , y30848 , y30849 , y30850 , y30851 , y30852 , y30853 , y30854 , y30855 , y30856 , y30857 , y30858 , y30859 , y30860 , y30861 , y30862 , y30863 , y30864 , y30865 , y30866 , y30867 , y30868 , y30869 , y30870 , y30871 , y30872 , y30873 , y30874 , y30875 , y30876 , y30877 , y30878 , y30879 , y30880 , y30881 , y30882 , y30883 , y30884 , y30885 , y30886 , y30887 , y30888 , y30889 , y30890 , y30891 , y30892 , y30893 , y30894 , y30895 , y30896 , y30897 , y30898 , y30899 , y30900 , y30901 , y30902 , y30903 , y30904 , y30905 , y30906 , y30907 , y30908 , y30909 , y30910 , y30911 , y30912 , y30913 , y30914 , y30915 , y30916 , y30917 , y30918 , y30919 , y30920 , y30921 , y30922 , y30923 , y30924 , y30925 , y30926 , y30927 , y30928 , y30929 , y30930 , y30931 , y30932 , y30933 , y30934 , y30935 , y30936 , y30937 , y30938 , y30939 , y30940 , y30941 , y30942 , y30943 , y30944 , y30945 , y30946 , y30947 , y30948 , y30949 , y30950 , y30951 , y30952 , y30953 , y30954 , y30955 , y30956 , y30957 , y30958 , y30959 , y30960 , y30961 , y30962 , y30963 , y30964 , y30965 , y30966 , y30967 , y30968 , y30969 , y30970 , y30971 , y30972 , y30973 , y30974 , y30975 , y30976 , y30977 , y30978 , y30979 , y30980 , y30981 , y30982 , y30983 , y30984 , y30985 , y30986 , y30987 , y30988 , y30989 , y30990 , y30991 , y30992 , y30993 , y30994 , y30995 , y30996 , y30997 , y30998 , y30999 , y31000 , y31001 , y31002 , y31003 , y31004 , y31005 , y31006 , y31007 , y31008 , y31009 , y31010 , y31011 , y31012 , y31013 , y31014 , y31015 , y31016 , y31017 , y31018 , y31019 , y31020 , y31021 , y31022 , y31023 , y31024 , y31025 , y31026 , y31027 , y31028 , y31029 , y31030 , y31031 , y31032 , y31033 , y31034 , y31035 , y31036 , y31037 , y31038 , y31039 , y31040 , y31041 , y31042 , y31043 , y31044 , y31045 , y31046 , y31047 , y31048 , y31049 , y31050 , y31051 , y31052 , y31053 , y31054 , y31055 , y31056 , y31057 , y31058 , y31059 , y31060 , y31061 , y31062 , y31063 , y31064 , y31065 , y31066 , y31067 , y31068 , y31069 , y31070 , y31071 , y31072 , y31073 , y31074 , y31075 , y31076 , y31077 , y31078 , y31079 , y31080 , y31081 , y31082 , y31083 , y31084 , y31085 , y31086 , y31087 , y31088 , y31089 , y31090 , y31091 , y31092 , y31093 , y31094 , y31095 , y31096 , y31097 , y31098 , y31099 , y31100 , y31101 , y31102 , y31103 , y31104 , y31105 , y31106 , y31107 , y31108 , y31109 , y31110 , y31111 , y31112 , y31113 , y31114 , y31115 , y31116 , y31117 , y31118 , y31119 , y31120 , y31121 , y31122 , y31123 , y31124 , y31125 , y31126 , y31127 , y31128 , y31129 , y31130 , y31131 , y31132 , y31133 , y31134 , y31135 , y31136 , y31137 , y31138 , y31139 , y31140 , y31141 , y31142 , y31143 , y31144 , y31145 , y31146 , y31147 , y31148 , y31149 , y31150 , y31151 , y31152 , y31153 , y31154 , y31155 , y31156 , y31157 , y31158 , y31159 , y31160 , y31161 , y31162 , y31163 , y31164 , y31165 , y31166 , y31167 , y31168 , y31169 , y31170 , y31171 , y31172 , y31173 , y31174 , y31175 , y31176 , y31177 , y31178 , y31179 , y31180 , y31181 , y31182 , y31183 , y31184 , y31185 , y31186 , y31187 , y31188 , y31189 , y31190 , y31191 , y31192 , y31193 , y31194 , y31195 , y31196 , y31197 , y31198 , y31199 , y31200 , y31201 , y31202 , y31203 , y31204 , y31205 , y31206 , y31207 , y31208 , y31209 , y31210 , y31211 , y31212 , y31213 , y31214 , y31215 , y31216 , y31217 , y31218 , y31219 , y31220 , y31221 , y31222 , y31223 , y31224 , y31225 , y31226 , y31227 , y31228 , y31229 , y31230 , y31231 , y31232 , y31233 , y31234 , y31235 , y31236 , y31237 , y31238 , y31239 , y31240 , y31241 , y31242 , y31243 , y31244 , y31245 , y31246 , y31247 , y31248 , y31249 , y31250 , y31251 , y31252 , y31253 , y31254 , y31255 , y31256 , y31257 , y31258 , y31259 , y31260 , y31261 , y31262 , y31263 , y31264 , y31265 , y31266 , y31267 , y31268 , y31269 , y31270 , y31271 , y31272 , y31273 , y31274 , y31275 , y31276 , y31277 , y31278 , y31279 , y31280 , y31281 , y31282 , y31283 , y31284 , y31285 , y31286 , y31287 , y31288 , y31289 , y31290 , y31291 , y31292 , y31293 , y31294 , y31295 , y31296 , y31297 , y31298 , y31299 , y31300 , y31301 , y31302 , y31303 , y31304 , y31305 , y31306 , y31307 , y31308 , y31309 , y31310 , y31311 , y31312 , y31313 , y31314 , y31315 , y31316 , y31317 , y31318 , y31319 , y31320 , y31321 , y31322 , y31323 , y31324 , y31325 , y31326 , y31327 , y31328 , y31329 , y31330 , y31331 , y31332 , y31333 , y31334 , y31335 , y31336 , y31337 , y31338 , y31339 , y31340 , y31341 , y31342 , y31343 , y31344 , y31345 , y31346 , y31347 , y31348 , y31349 , y31350 , y31351 , y31352 , y31353 , y31354 , y31355 , y31356 , y31357 , y31358 , y31359 , y31360 , y31361 , y31362 , y31363 , y31364 , y31365 , y31366 , y31367 , y31368 , y31369 , y31370 , y31371 , y31372 , y31373 , y31374 , y31375 , y31376 , y31377 , y31378 , y31379 , y31380 , y31381 , y31382 , y31383 , y31384 , y31385 , y31386 , y31387 , y31388 , y31389 , y31390 , y31391 , y31392 , y31393 , y31394 , y31395 , y31396 , y31397 , y31398 , y31399 , y31400 , y31401 , y31402 , y31403 , y31404 , y31405 , y31406 , y31407 , y31408 , y31409 , y31410 , y31411 , y31412 , y31413 , y31414 , y31415 , y31416 , y31417 , y31418 , y31419 , y31420 , y31421 , y31422 , y31423 , y31424 , y31425 , y31426 , y31427 , y31428 , y31429 , y31430 , y31431 , y31432 , y31433 , y31434 , y31435 , y31436 , y31437 , y31438 , y31439 , y31440 , y31441 , y31442 , y31443 , y31444 , y31445 , y31446 , y31447 , y31448 , y31449 , y31450 , y31451 , y31452 , y31453 , y31454 , y31455 , y31456 , y31457 , y31458 , y31459 , y31460 , y31461 , y31462 , y31463 , y31464 , y31465 , y31466 , y31467 , y31468 , y31469 , y31470 , y31471 , y31472 , y31473 , y31474 , y31475 , y31476 , y31477 , y31478 , y31479 , y31480 , y31481 , y31482 , y31483 , y31484 , y31485 , y31486 , y31487 , y31488 , y31489 , y31490 , y31491 , y31492 , y31493 , y31494 , y31495 , y31496 , y31497 , y31498 , y31499 , y31500 , y31501 , y31502 , y31503 , y31504 , y31505 , y31506 , y31507 , y31508 , y31509 , y31510 , y31511 , y31512 , y31513 , y31514 , y31515 , y31516 , y31517 , y31518 , y31519 , y31520 , y31521 , y31522 , y31523 , y31524 , y31525 , y31526 , y31527 , y31528 , y31529 , y31530 , y31531 , y31532 , y31533 , y31534 , y31535 , y31536 , y31537 , y31538 , y31539 , y31540 , y31541 , y31542 , y31543 , y31544 , y31545 , y31546 , y31547 , y31548 , y31549 , y31550 , y31551 , y31552 , y31553 , y31554 , y31555 , y31556 , y31557 , y31558 , y31559 , y31560 , y31561 , y31562 , y31563 , y31564 , y31565 , y31566 , y31567 , y31568 , y31569 , y31570 , y31571 , y31572 , y31573 , y31574 , y31575 , y31576 , y31577 , y31578 , y31579 , y31580 , y31581 , y31582 , y31583 , y31584 , y31585 , y31586 , y31587 , y31588 , y31589 , y31590 , y31591 , y31592 , y31593 , y31594 , y31595 , y31596 , y31597 , y31598 , y31599 , y31600 , y31601 , y31602 , y31603 , y31604 , y31605 , y31606 , y31607 , y31608 , y31609 , y31610 , y31611 , y31612 , y31613 , y31614 , y31615 , y31616 , y31617 , y31618 , y31619 , y31620 , y31621 , y31622 , y31623 , y31624 , y31625 , y31626 , y31627 , y31628 , y31629 , y31630 , y31631 , y31632 , y31633 , y31634 , y31635 , y31636 , y31637 , y31638 , y31639 , y31640 , y31641 , y31642 , y31643 , y31644 , y31645 , y31646 , y31647 , y31648 , y31649 , y31650 , y31651 , y31652 , y31653 , y31654 , y31655 , y31656 , y31657 , y31658 , y31659 , y31660 , y31661 , y31662 , y31663 , y31664 , y31665 , y31666 , y31667 , y31668 , y31669 , y31670 , y31671 , y31672 , y31673 , y31674 , y31675 , y31676 , y31677 , y31678 , y31679 , y31680 , y31681 , y31682 , y31683 , y31684 , y31685 , y31686 , y31687 , y31688 , y31689 , y31690 , y31691 , y31692 , y31693 , y31694 , y31695 , y31696 , y31697 , y31698 , y31699 , y31700 , y31701 , y31702 , y31703 , y31704 , y31705 , y31706 , y31707 , y31708 , y31709 , y31710 , y31711 , y31712 , y31713 , y31714 , y31715 , y31716 , y31717 , y31718 , y31719 , y31720 , y31721 , y31722 , y31723 , y31724 , y31725 , y31726 , y31727 , y31728 , y31729 , y31730 , y31731 , y31732 , y31733 , y31734 , y31735 , y31736 , y31737 , y31738 , y31739 , y31740 , y31741 , y31742 , y31743 , y31744 , y31745 , y31746 , y31747 , y31748 , y31749 , y31750 , y31751 , y31752 , y31753 , y31754 , y31755 , y31756 , y31757 , y31758 , y31759 , y31760 , y31761 , y31762 , y31763 , y31764 , y31765 , y31766 , y31767 , y31768 , y31769 , y31770 , y31771 , y31772 , y31773 , y31774 , y31775 , y31776 , y31777 , y31778 , y31779 , y31780 , y31781 , y31782 , y31783 , y31784 , y31785 , y31786 , y31787 , y31788 , y31789 , y31790 , y31791 , y31792 , y31793 , y31794 , y31795 , y31796 , y31797 , y31798 , y31799 , y31800 , y31801 , y31802 , y31803 , y31804 , y31805 , y31806 , y31807 , y31808 , y31809 , y31810 , y31811 , y31812 , y31813 , y31814 , y31815 , y31816 , y31817 , y31818 , y31819 , y31820 , y31821 , y31822 , y31823 , y31824 , y31825 , y31826 , y31827 , y31828 , y31829 , y31830 , y31831 , y31832 , y31833 , y31834 , y31835 , y31836 , y31837 , y31838 , y31839 , y31840 , y31841 , y31842 , y31843 , y31844 , y31845 , y31846 , y31847 , y31848 , y31849 , y31850 , y31851 , y31852 , y31853 , y31854 , y31855 , y31856 , y31857 , y31858 , y31859 , y31860 , y31861 , y31862 , y31863 , y31864 , y31865 , y31866 , y31867 , y31868 , y31869 , y31870 , y31871 , y31872 , y31873 , y31874 , y31875 , y31876 , y31877 , y31878 , y31879 , y31880 , y31881 , y31882 , y31883 , y31884 , y31885 , y31886 , y31887 , y31888 , y31889 , y31890 , y31891 , y31892 , y31893 , y31894 , y31895 , y31896 , y31897 , y31898 , y31899 , y31900 , y31901 , y31902 , y31903 , y31904 , y31905 , y31906 , y31907 , y31908 , y31909 , y31910 , y31911 , y31912 , y31913 , y31914 , y31915 , y31916 , y31917 , y31918 , y31919 , y31920 , y31921 , y31922 , y31923 , y31924 , y31925 , y31926 , y31927 , y31928 , y31929 , y31930 , y31931 , y31932 , y31933 , y31934 , y31935 , y31936 , y31937 , y31938 , y31939 , y31940 , y31941 , y31942 , y31943 , y31944 , y31945 , y31946 , y31947 , y31948 , y31949 , y31950 , y31951 , y31952 , y31953 , y31954 , y31955 , y31956 , y31957 , y31958 , y31959 , y31960 , y31961 , y31962 , y31963 , y31964 , y31965 , y31966 , y31967 , y31968 , y31969 , y31970 , y31971 , y31972 , y31973 , y31974 , y31975 , y31976 , y31977 , y31978 , y31979 , y31980 , y31981 , y31982 , y31983 , y31984 , y31985 , y31986 , y31987 , y31988 , y31989 , y31990 , y31991 , y31992 , y31993 , y31994 , y31995 , y31996 , y31997 , y31998 , y31999 , y32000 , y32001 , y32002 , y32003 , y32004 , y32005 , y32006 , y32007 , y32008 , y32009 , y32010 , y32011 , y32012 , y32013 , y32014 , y32015 , y32016 , y32017 , y32018 , y32019 , y32020 , y32021 , y32022 , y32023 , y32024 , y32025 , y32026 , y32027 , y32028 , y32029 , y32030 , y32031 , y32032 , y32033 , y32034 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 , y256 , y257 , y258 , y259 , y260 , y261 , y262 , y263 , y264 , y265 , y266 , y267 , y268 , y269 , y270 , y271 , y272 , y273 , y274 , y275 , y276 , y277 , y278 , y279 , y280 , y281 , y282 , y283 , y284 , y285 , y286 , y287 , y288 , y289 , y290 , y291 , y292 , y293 , y294 , y295 , y296 , y297 , y298 , y299 , y300 , y301 , y302 , y303 , y304 , y305 , y306 , y307 , y308 , y309 , y310 , y311 , y312 , y313 , y314 , y315 , y316 , y317 , y318 , y319 , y320 , y321 , y322 , y323 , y324 , y325 , y326 , y327 , y328 , y329 , y330 , y331 , y332 , y333 , y334 , y335 , y336 , y337 , y338 , y339 , y340 , y341 , y342 , y343 , y344 , y345 , y346 , y347 , y348 , y349 , y350 , y351 , y352 , y353 , y354 , y355 , y356 , y357 , y358 , y359 , y360 , y361 , y362 , y363 , y364 , y365 , y366 , y367 , y368 , y369 , y370 , y371 , y372 , y373 , y374 , y375 , y376 , y377 , y378 , y379 , y380 , y381 , y382 , y383 , y384 , y385 , y386 , y387 , y388 , y389 , y390 , y391 , y392 , y393 , y394 , y395 , y396 , y397 , y398 , y399 , y400 , y401 , y402 , y403 , y404 , y405 , y406 , y407 , y408 , y409 , y410 , y411 , y412 , y413 , y414 , y415 , y416 , y417 , y418 , y419 , y420 , y421 , y422 , y423 , y424 , y425 , y426 , y427 , y428 , y429 , y430 , y431 , y432 , y433 , y434 , y435 , y436 , y437 , y438 , y439 , y440 , y441 , y442 , y443 , y444 , y445 , y446 , y447 , y448 , y449 , y450 , y451 , y452 , y453 , y454 , y455 , y456 , y457 , y458 , y459 , y460 , y461 , y462 , y463 , y464 , y465 , y466 , y467 , y468 , y469 , y470 , y471 , y472 , y473 , y474 , y475 , y476 , y477 , y478 , y479 , y480 , y481 , y482 , y483 , y484 , y485 , y486 , y487 , y488 , y489 , y490 , y491 , y492 , y493 , y494 , y495 , y496 , y497 , y498 , y499 , y500 , y501 , y502 , y503 , y504 , y505 , y506 , y507 , y508 , y509 , y510 , y511 , y512 , y513 , y514 , y515 , y516 , y517 , y518 , y519 , y520 , y521 , y522 , y523 , y524 , y525 , y526 , y527 , y528 , y529 , y530 , y531 , y532 , y533 , y534 , y535 , y536 , y537 , y538 , y539 , y540 , y541 , y542 , y543 , y544 , y545 , y546 , y547 , y548 , y549 , y550 , y551 , y552 , y553 , y554 , y555 , y556 , y557 , y558 , y559 , y560 , y561 , y562 , y563 , y564 , y565 , y566 , y567 , y568 , y569 , y570 , y571 , y572 , y573 , y574 , y575 , y576 , y577 , y578 , y579 , y580 , y581 , y582 , y583 , y584 , y585 , y586 , y587 , y588 , y589 , y590 , y591 , y592 , y593 , y594 , y595 , y596 , y597 , y598 , y599 , y600 , y601 , y602 , y603 , y604 , y605 , y606 , y607 , y608 , y609 , y610 , y611 , y612 , y613 , y614 , y615 , y616 , y617 , y618 , y619 , y620 , y621 , y622 , y623 , y624 , y625 , y626 , y627 , y628 , y629 , y630 , y631 , y632 , y633 , y634 , y635 , y636 , y637 , y638 , y639 , y640 , y641 , y642 , y643 , y644 , y645 , y646 , y647 , y648 , y649 , y650 , y651 , y652 , y653 , y654 , y655 , y656 , y657 , y658 , y659 , y660 , y661 , y662 , y663 , y664 , y665 , y666 , y667 , y668 , y669 , y670 , y671 , y672 , y673 , y674 , y675 , y676 , y677 , y678 , y679 , y680 , y681 , y682 , y683 , y684 , y685 , y686 , y687 , y688 , y689 , y690 , y691 , y692 , y693 , y694 , y695 , y696 , y697 , y698 , y699 , y700 , y701 , y702 , y703 , y704 , y705 , y706 , y707 , y708 , y709 , y710 , y711 , y712 , y713 , y714 , y715 , y716 , y717 , y718 , y719 , y720 , y721 , y722 , y723 , y724 , y725 , y726 , y727 , y728 , y729 , y730 , y731 , y732 , y733 , y734 , y735 , y736 , y737 , y738 , y739 , y740 , y741 , y742 , y743 , y744 , y745 , y746 , y747 , y748 , y749 , y750 , y751 , y752 , y753 , y754 , y755 , y756 , y757 , y758 , y759 , y760 , y761 , y762 , y763 , y764 , y765 , y766 , y767 , y768 , y769 , y770 , y771 , y772 , y773 , y774 , y775 , y776 , y777 , y778 , y779 , y780 , y781 , y782 , y783 , y784 , y785 , y786 , y787 , y788 , y789 , y790 , y791 , y792 , y793 , y794 , y795 , y796 , y797 , y798 , y799 , y800 , y801 , y802 , y803 , y804 , y805 , y806 , y807 , y808 , y809 , y810 , y811 , y812 , y813 , y814 , y815 , y816 , y817 , y818 , y819 , y820 , y821 , y822 , y823 , y824 , y825 , y826 , y827 , y828 , y829 , y830 , y831 , y832 , y833 , y834 , y835 , y836 , y837 , y838 , y839 , y840 , y841 , y842 , y843 , y844 , y845 , y846 , y847 , y848 , y849 , y850 , y851 , y852 , y853 , y854 , y855 , y856 , y857 , y858 , y859 , y860 , y861 , y862 , y863 , y864 , y865 , y866 , y867 , y868 , y869 , y870 , y871 , y872 , y873 , y874 , y875 , y876 , y877 , y878 , y879 , y880 , y881 , y882 , y883 , y884 , y885 , y886 , y887 , y888 , y889 , y890 , y891 , y892 , y893 , y894 , y895 , y896 , y897 , y898 , y899 , y900 , y901 , y902 , y903 , y904 , y905 , y906 , y907 , y908 , y909 , y910 , y911 , y912 , y913 , y914 , y915 , y916 , y917 , y918 , y919 , y920 , y921 , y922 , y923 , y924 , y925 , y926 , y927 , y928 , y929 , y930 , y931 , y932 , y933 , y934 , y935 , y936 , y937 , y938 , y939 , y940 , y941 , y942 , y943 , y944 , y945 , y946 , y947 , y948 , y949 , y950 , y951 , y952 , y953 , y954 , y955 , y956 , y957 , y958 , y959 , y960 , y961 , y962 , y963 , y964 , y965 , y966 , y967 , y968 , y969 , y970 , y971 , y972 , y973 , y974 , y975 , y976 , y977 , y978 , y979 , y980 , y981 , y982 , y983 , y984 , y985 , y986 , y987 , y988 , y989 , y990 , y991 , y992 , y993 , y994 , y995 , y996 , y997 , y998 , y999 , y1000 , y1001 , y1002 , y1003 , y1004 , y1005 , y1006 , y1007 , y1008 , y1009 , y1010 , y1011 , y1012 , y1013 , y1014 , y1015 , y1016 , y1017 , y1018 , y1019 , y1020 , y1021 , y1022 , y1023 , y1024 , y1025 , y1026 , y1027 , y1028 , y1029 , y1030 , y1031 , y1032 , y1033 , y1034 , y1035 , y1036 , y1037 , y1038 , y1039 , y1040 , y1041 , y1042 , y1043 , y1044 , y1045 , y1046 , y1047 , y1048 , y1049 , y1050 , y1051 , y1052 , y1053 , y1054 , y1055 , y1056 , y1057 , y1058 , y1059 , y1060 , y1061 , y1062 , y1063 , y1064 , y1065 , y1066 , y1067 , y1068 , y1069 , y1070 , y1071 , y1072 , y1073 , y1074 , y1075 , y1076 , y1077 , y1078 , y1079 , y1080 , y1081 , y1082 , y1083 , y1084 , y1085 , y1086 , y1087 , y1088 , y1089 , y1090 , y1091 , y1092 , y1093 , y1094 , y1095 , y1096 , y1097 , y1098 , y1099 , y1100 , y1101 , y1102 , y1103 , y1104 , y1105 , y1106 , y1107 , y1108 , y1109 , y1110 , y1111 , y1112 , y1113 , y1114 , y1115 , y1116 , y1117 , y1118 , y1119 , y1120 , y1121 , y1122 , y1123 , y1124 , y1125 , y1126 , y1127 , y1128 , y1129 , y1130 , y1131 , y1132 , y1133 , y1134 , y1135 , y1136 , y1137 , y1138 , y1139 , y1140 , y1141 , y1142 , y1143 , y1144 , y1145 , y1146 , y1147 , y1148 , y1149 , y1150 , y1151 , y1152 , y1153 , y1154 , y1155 , y1156 , y1157 , y1158 , y1159 , y1160 , y1161 , y1162 , y1163 , y1164 , y1165 , y1166 , y1167 , y1168 , y1169 , y1170 , y1171 , y1172 , y1173 , y1174 , y1175 , y1176 , y1177 , y1178 , y1179 , y1180 , y1181 , y1182 , y1183 , y1184 , y1185 , y1186 , y1187 , y1188 , y1189 , y1190 , y1191 , y1192 , y1193 , y1194 , y1195 , y1196 , y1197 , y1198 , y1199 , y1200 , y1201 , y1202 , y1203 , y1204 , y1205 , y1206 , y1207 , y1208 , y1209 , y1210 , y1211 , y1212 , y1213 , y1214 , y1215 , y1216 , y1217 , y1218 , y1219 , y1220 , y1221 , y1222 , y1223 , y1224 , y1225 , y1226 , y1227 , y1228 , y1229 , y1230 , y1231 , y1232 , y1233 , y1234 , y1235 , y1236 , y1237 , y1238 , y1239 , y1240 , y1241 , y1242 , y1243 , y1244 , y1245 , y1246 , y1247 , y1248 , y1249 , y1250 , y1251 , y1252 , y1253 , y1254 , y1255 , y1256 , y1257 , y1258 , y1259 , y1260 , y1261 , y1262 , y1263 , y1264 , y1265 , y1266 , y1267 , y1268 , y1269 , y1270 , y1271 , y1272 , y1273 , y1274 , y1275 , y1276 , y1277 , y1278 , y1279 , y1280 , y1281 , y1282 , y1283 , y1284 , y1285 , y1286 , y1287 , y1288 , y1289 , y1290 , y1291 , y1292 , y1293 , y1294 , y1295 , y1296 , y1297 , y1298 , y1299 , y1300 , y1301 , y1302 , y1303 , y1304 , y1305 , y1306 , y1307 , y1308 , y1309 , y1310 , y1311 , y1312 , y1313 , y1314 , y1315 , y1316 , y1317 , y1318 , y1319 , y1320 , y1321 , y1322 , y1323 , y1324 , y1325 , y1326 , y1327 , y1328 , y1329 , y1330 , y1331 , y1332 , y1333 , y1334 , y1335 , y1336 , y1337 , y1338 , y1339 , y1340 , y1341 , y1342 , y1343 , y1344 , y1345 , y1346 , y1347 , y1348 , y1349 , y1350 , y1351 , y1352 , y1353 , y1354 , y1355 , y1356 , y1357 , y1358 , y1359 , y1360 , y1361 , y1362 , y1363 , y1364 , y1365 , y1366 , y1367 , y1368 , y1369 , y1370 , y1371 , y1372 , y1373 , y1374 , y1375 , y1376 , y1377 , y1378 , y1379 , y1380 , y1381 , y1382 , y1383 , y1384 , y1385 , y1386 , y1387 , y1388 , y1389 , y1390 , y1391 , y1392 , y1393 , y1394 , y1395 , y1396 , y1397 , y1398 , y1399 , y1400 , y1401 , y1402 , y1403 , y1404 , y1405 , y1406 , y1407 , y1408 , y1409 , y1410 , y1411 , y1412 , y1413 , y1414 , y1415 , y1416 , y1417 , y1418 , y1419 , y1420 , y1421 , y1422 , y1423 , y1424 , y1425 , y1426 , y1427 , y1428 , y1429 , y1430 , y1431 , y1432 , y1433 , y1434 , y1435 , y1436 , y1437 , y1438 , y1439 , y1440 , y1441 , y1442 , y1443 , y1444 , y1445 , y1446 , y1447 , y1448 , y1449 , y1450 , y1451 , y1452 , y1453 , y1454 , y1455 , y1456 , y1457 , y1458 , y1459 , y1460 , y1461 , y1462 , y1463 , y1464 , y1465 , y1466 , y1467 , y1468 , y1469 , y1470 , y1471 , y1472 , y1473 , y1474 , y1475 , y1476 , y1477 , y1478 , y1479 , y1480 , y1481 , y1482 , y1483 , y1484 , y1485 , y1486 , y1487 , y1488 , y1489 , y1490 , y1491 , y1492 , y1493 , y1494 , y1495 , y1496 , y1497 , y1498 , y1499 , y1500 , y1501 , y1502 , y1503 , y1504 , y1505 , y1506 , y1507 , y1508 , y1509 , y1510 , y1511 , y1512 , y1513 , y1514 , y1515 , y1516 , y1517 , y1518 , y1519 , y1520 , y1521 , y1522 , y1523 , y1524 , y1525 , y1526 , y1527 , y1528 , y1529 , y1530 , y1531 , y1532 , y1533 , y1534 , y1535 , y1536 , y1537 , y1538 , y1539 , y1540 , y1541 , y1542 , y1543 , y1544 , y1545 , y1546 , y1547 , y1548 , y1549 , y1550 , y1551 , y1552 , y1553 , y1554 , y1555 , y1556 , y1557 , y1558 , y1559 , y1560 , y1561 , y1562 , y1563 , y1564 , y1565 , y1566 , y1567 , y1568 , y1569 , y1570 , y1571 , y1572 , y1573 , y1574 , y1575 , y1576 , y1577 , y1578 , y1579 , y1580 , y1581 , y1582 , y1583 , y1584 , y1585 , y1586 , y1587 , y1588 , y1589 , y1590 , y1591 , y1592 , y1593 , y1594 , y1595 , y1596 , y1597 , y1598 , y1599 , y1600 , y1601 , y1602 , y1603 , y1604 , y1605 , y1606 , y1607 , y1608 , y1609 , y1610 , y1611 , y1612 , y1613 , y1614 , y1615 , y1616 , y1617 , y1618 , y1619 , y1620 , y1621 , y1622 , y1623 , y1624 , y1625 , y1626 , y1627 , y1628 , y1629 , y1630 , y1631 , y1632 , y1633 , y1634 , y1635 , y1636 , y1637 , y1638 , y1639 , y1640 , y1641 , y1642 , y1643 , y1644 , y1645 , y1646 , y1647 , y1648 , y1649 , y1650 , y1651 , y1652 , y1653 , y1654 , y1655 , y1656 , y1657 , y1658 , y1659 , y1660 , y1661 , y1662 , y1663 , y1664 , y1665 , y1666 , y1667 , y1668 , y1669 , y1670 , y1671 , y1672 , y1673 , y1674 , y1675 , y1676 , y1677 , y1678 , y1679 , y1680 , y1681 , y1682 , y1683 , y1684 , y1685 , y1686 , y1687 , y1688 , y1689 , y1690 , y1691 , y1692 , y1693 , y1694 , y1695 , y1696 , y1697 , y1698 , y1699 , y1700 , y1701 , y1702 , y1703 , y1704 , y1705 , y1706 , y1707 , y1708 , y1709 , y1710 , y1711 , y1712 , y1713 , y1714 , y1715 , y1716 , y1717 , y1718 , y1719 , y1720 , y1721 , y1722 , y1723 , y1724 , y1725 , y1726 , y1727 , y1728 , y1729 , y1730 , y1731 , y1732 , y1733 , y1734 , y1735 , y1736 , y1737 , y1738 , y1739 , y1740 , y1741 , y1742 , y1743 , y1744 , y1745 , y1746 , y1747 , y1748 , y1749 , y1750 , y1751 , y1752 , y1753 , y1754 , y1755 , y1756 , y1757 , y1758 , y1759 , y1760 , y1761 , y1762 , y1763 , y1764 , y1765 , y1766 , y1767 , y1768 , y1769 , y1770 , y1771 , y1772 , y1773 , y1774 , y1775 , y1776 , y1777 , y1778 , y1779 , y1780 , y1781 , y1782 , y1783 , y1784 , y1785 , y1786 , y1787 , y1788 , y1789 , y1790 , y1791 , y1792 , y1793 , y1794 , y1795 , y1796 , y1797 , y1798 , y1799 , y1800 , y1801 , y1802 , y1803 , y1804 , y1805 , y1806 , y1807 , y1808 , y1809 , y1810 , y1811 , y1812 , y1813 , y1814 , y1815 , y1816 , y1817 , y1818 , y1819 , y1820 , y1821 , y1822 , y1823 , y1824 , y1825 , y1826 , y1827 , y1828 , y1829 , y1830 , y1831 , y1832 , y1833 , y1834 , y1835 , y1836 , y1837 , y1838 , y1839 , y1840 , y1841 , y1842 , y1843 , y1844 , y1845 , y1846 , y1847 , y1848 , y1849 , y1850 , y1851 , y1852 , y1853 , y1854 , y1855 , y1856 , y1857 , y1858 , y1859 , y1860 , y1861 , y1862 , y1863 , y1864 , y1865 , y1866 , y1867 , y1868 , y1869 , y1870 , y1871 , y1872 , y1873 , y1874 , y1875 , y1876 , y1877 , y1878 , y1879 , y1880 , y1881 , y1882 , y1883 , y1884 , y1885 , y1886 , y1887 , y1888 , y1889 , y1890 , y1891 , y1892 , y1893 , y1894 , y1895 , y1896 , y1897 , y1898 , y1899 , y1900 , y1901 , y1902 , y1903 , y1904 , y1905 , y1906 , y1907 , y1908 , y1909 , y1910 , y1911 , y1912 , y1913 , y1914 , y1915 , y1916 , y1917 , y1918 , y1919 , y1920 , y1921 , y1922 , y1923 , y1924 , y1925 , y1926 , y1927 , y1928 , y1929 , y1930 , y1931 , y1932 , y1933 , y1934 , y1935 , y1936 , y1937 , y1938 , y1939 , y1940 , y1941 , y1942 , y1943 , y1944 , y1945 , y1946 , y1947 , y1948 , y1949 , y1950 , y1951 , y1952 , y1953 , y1954 , y1955 , y1956 , y1957 , y1958 , y1959 , y1960 , y1961 , y1962 , y1963 , y1964 , y1965 , y1966 , y1967 , y1968 , y1969 , y1970 , y1971 , y1972 , y1973 , y1974 , y1975 , y1976 , y1977 , y1978 , y1979 , y1980 , y1981 , y1982 , y1983 , y1984 , y1985 , y1986 , y1987 , y1988 , y1989 , y1990 , y1991 , y1992 , y1993 , y1994 , y1995 , y1996 , y1997 , y1998 , y1999 , y2000 , y2001 , y2002 , y2003 , y2004 , y2005 , y2006 , y2007 , y2008 , y2009 , y2010 , y2011 , y2012 , y2013 , y2014 , y2015 , y2016 , y2017 , y2018 , y2019 , y2020 , y2021 , y2022 , y2023 , y2024 , y2025 , y2026 , y2027 , y2028 , y2029 , y2030 , y2031 , y2032 , y2033 , y2034 , y2035 , y2036 , y2037 , y2038 , y2039 , y2040 , y2041 , y2042 , y2043 , y2044 , y2045 , y2046 , y2047 , y2048 , y2049 , y2050 , y2051 , y2052 , y2053 , y2054 , y2055 , y2056 , y2057 , y2058 , y2059 , y2060 , y2061 , y2062 , y2063 , y2064 , y2065 , y2066 , y2067 , y2068 , y2069 , y2070 , y2071 , y2072 , y2073 , y2074 , y2075 , y2076 , y2077 , y2078 , y2079 , y2080 , y2081 , y2082 , y2083 , y2084 , y2085 , y2086 , y2087 , y2088 , y2089 , y2090 , y2091 , y2092 , y2093 , y2094 , y2095 , y2096 , y2097 , y2098 , y2099 , y2100 , y2101 , y2102 , y2103 , y2104 , y2105 , y2106 , y2107 , y2108 , y2109 , y2110 , y2111 , y2112 , y2113 , y2114 , y2115 , y2116 , y2117 , y2118 , y2119 , y2120 , y2121 , y2122 , y2123 , y2124 , y2125 , y2126 , y2127 , y2128 , y2129 , y2130 , y2131 , y2132 , y2133 , y2134 , y2135 , y2136 , y2137 , y2138 , y2139 , y2140 , y2141 , y2142 , y2143 , y2144 , y2145 , y2146 , y2147 , y2148 , y2149 , y2150 , y2151 , y2152 , y2153 , y2154 , y2155 , y2156 , y2157 , y2158 , y2159 , y2160 , y2161 , y2162 , y2163 , y2164 , y2165 , y2166 , y2167 , y2168 , y2169 , y2170 , y2171 , y2172 , y2173 , y2174 , y2175 , y2176 , y2177 , y2178 , y2179 , y2180 , y2181 , y2182 , y2183 , y2184 , y2185 , y2186 , y2187 , y2188 , y2189 , y2190 , y2191 , y2192 , y2193 , y2194 , y2195 , y2196 , y2197 , y2198 , y2199 , y2200 , y2201 , y2202 , y2203 , y2204 , y2205 , y2206 , y2207 , y2208 , y2209 , y2210 , y2211 , y2212 , y2213 , y2214 , y2215 , y2216 , y2217 , y2218 , y2219 , y2220 , y2221 , y2222 , y2223 , y2224 , y2225 , y2226 , y2227 , y2228 , y2229 , y2230 , y2231 , y2232 , y2233 , y2234 , y2235 , y2236 , y2237 , y2238 , y2239 , y2240 , y2241 , y2242 , y2243 , y2244 , y2245 , y2246 , y2247 , y2248 , y2249 , y2250 , y2251 , y2252 , y2253 , y2254 , y2255 , y2256 , y2257 , y2258 , y2259 , y2260 , y2261 , y2262 , y2263 , y2264 , y2265 , y2266 , y2267 , y2268 , y2269 , y2270 , y2271 , y2272 , y2273 , y2274 , y2275 , y2276 , y2277 , y2278 , y2279 , y2280 , y2281 , y2282 , y2283 , y2284 , y2285 , y2286 , y2287 , y2288 , y2289 , y2290 , y2291 , y2292 , y2293 , y2294 , y2295 , y2296 , y2297 , y2298 , y2299 , y2300 , y2301 , y2302 , y2303 , y2304 , y2305 , y2306 , y2307 , y2308 , y2309 , y2310 , y2311 , y2312 , y2313 , y2314 , y2315 , y2316 , y2317 , y2318 , y2319 , y2320 , y2321 , y2322 , y2323 , y2324 , y2325 , y2326 , y2327 , y2328 , y2329 , y2330 , y2331 , y2332 , y2333 , y2334 , y2335 , y2336 , y2337 , y2338 , y2339 , y2340 , y2341 , y2342 , y2343 , y2344 , y2345 , y2346 , y2347 , y2348 , y2349 , y2350 , y2351 , y2352 , y2353 , y2354 , y2355 , y2356 , y2357 , y2358 , y2359 , y2360 , y2361 , y2362 , y2363 , y2364 , y2365 , y2366 , y2367 , y2368 , y2369 , y2370 , y2371 , y2372 , y2373 , y2374 , y2375 , y2376 , y2377 , y2378 , y2379 , y2380 , y2381 , y2382 , y2383 , y2384 , y2385 , y2386 , y2387 , y2388 , y2389 , y2390 , y2391 , y2392 , y2393 , y2394 , y2395 , y2396 , y2397 , y2398 , y2399 , y2400 , y2401 , y2402 , y2403 , y2404 , y2405 , y2406 , y2407 , y2408 , y2409 , y2410 , y2411 , y2412 , y2413 , y2414 , y2415 , y2416 , y2417 , y2418 , y2419 , y2420 , y2421 , y2422 , y2423 , y2424 , y2425 , y2426 , y2427 , y2428 , y2429 , y2430 , y2431 , y2432 , y2433 , y2434 , y2435 , y2436 , y2437 , y2438 , y2439 , y2440 , y2441 , y2442 , y2443 , y2444 , y2445 , y2446 , y2447 , y2448 , y2449 , y2450 , y2451 , y2452 , y2453 , y2454 , y2455 , y2456 , y2457 , y2458 , y2459 , y2460 , y2461 , y2462 , y2463 , y2464 , y2465 , y2466 , y2467 , y2468 , y2469 , y2470 , y2471 , y2472 , y2473 , y2474 , y2475 , y2476 , y2477 , y2478 , y2479 , y2480 , y2481 , y2482 , y2483 , y2484 , y2485 , y2486 , y2487 , y2488 , y2489 , y2490 , y2491 , y2492 , y2493 , y2494 , y2495 , y2496 , y2497 , y2498 , y2499 , y2500 , y2501 , y2502 , y2503 , y2504 , y2505 , y2506 , y2507 , y2508 , y2509 , y2510 , y2511 , y2512 , y2513 , y2514 , y2515 , y2516 , y2517 , y2518 , y2519 , y2520 , y2521 , y2522 , y2523 , y2524 , y2525 , y2526 , y2527 , y2528 , y2529 , y2530 , y2531 , y2532 , y2533 , y2534 , y2535 , y2536 , y2537 , y2538 , y2539 , y2540 , y2541 , y2542 , y2543 , y2544 , y2545 , y2546 , y2547 , y2548 , y2549 , y2550 , y2551 , y2552 , y2553 , y2554 , y2555 , y2556 , y2557 , y2558 , y2559 , y2560 , y2561 , y2562 , y2563 , y2564 , y2565 , y2566 , y2567 , y2568 , y2569 , y2570 , y2571 , y2572 , y2573 , y2574 , y2575 , y2576 , y2577 , y2578 , y2579 , y2580 , y2581 , y2582 , y2583 , y2584 , y2585 , y2586 , y2587 , y2588 , y2589 , y2590 , y2591 , y2592 , y2593 , y2594 , y2595 , y2596 , y2597 , y2598 , y2599 , y2600 , y2601 , y2602 , y2603 , y2604 , y2605 , y2606 , y2607 , y2608 , y2609 , y2610 , y2611 , y2612 , y2613 , y2614 , y2615 , y2616 , y2617 , y2618 , y2619 , y2620 , y2621 , y2622 , y2623 , y2624 , y2625 , y2626 , y2627 , y2628 , y2629 , y2630 , y2631 , y2632 , y2633 , y2634 , y2635 , y2636 , y2637 , y2638 , y2639 , y2640 , y2641 , y2642 , y2643 , y2644 , y2645 , y2646 , y2647 , y2648 , y2649 , y2650 , y2651 , y2652 , y2653 , y2654 , y2655 , y2656 , y2657 , y2658 , y2659 , y2660 , y2661 , y2662 , y2663 , y2664 , y2665 , y2666 , y2667 , y2668 , y2669 , y2670 , y2671 , y2672 , y2673 , y2674 , y2675 , y2676 , y2677 , y2678 , y2679 , y2680 , y2681 , y2682 , y2683 , y2684 , y2685 , y2686 , y2687 , y2688 , y2689 , y2690 , y2691 , y2692 , y2693 , y2694 , y2695 , y2696 , y2697 , y2698 , y2699 , y2700 , y2701 , y2702 , y2703 , y2704 , y2705 , y2706 , y2707 , y2708 , y2709 , y2710 , y2711 , y2712 , y2713 , y2714 , y2715 , y2716 , y2717 , y2718 , y2719 , y2720 , y2721 , y2722 , y2723 , y2724 , y2725 , y2726 , y2727 , y2728 , y2729 , y2730 , y2731 , y2732 , y2733 , y2734 , y2735 , y2736 , y2737 , y2738 , y2739 , y2740 , y2741 , y2742 , y2743 , y2744 , y2745 , y2746 , y2747 , y2748 , y2749 , y2750 , y2751 , y2752 , y2753 , y2754 , y2755 , y2756 , y2757 , y2758 , y2759 , y2760 , y2761 , y2762 , y2763 , y2764 , y2765 , y2766 , y2767 , y2768 , y2769 , y2770 , y2771 , y2772 , y2773 , y2774 , y2775 , y2776 , y2777 , y2778 , y2779 , y2780 , y2781 , y2782 , y2783 , y2784 , y2785 , y2786 , y2787 , y2788 , y2789 , y2790 , y2791 , y2792 , y2793 , y2794 , y2795 , y2796 , y2797 , y2798 , y2799 , y2800 , y2801 , y2802 , y2803 , y2804 , y2805 , y2806 , y2807 , y2808 , y2809 , y2810 , y2811 , y2812 , y2813 , y2814 , y2815 , y2816 , y2817 , y2818 , y2819 , y2820 , y2821 , y2822 , y2823 , y2824 , y2825 , y2826 , y2827 , y2828 , y2829 , y2830 , y2831 , y2832 , y2833 , y2834 , y2835 , y2836 , y2837 , y2838 , y2839 , y2840 , y2841 , y2842 , y2843 , y2844 , y2845 , y2846 , y2847 , y2848 , y2849 , y2850 , y2851 , y2852 , y2853 , y2854 , y2855 , y2856 , y2857 , y2858 , y2859 , y2860 , y2861 , y2862 , y2863 , y2864 , y2865 , y2866 , y2867 , y2868 , y2869 , y2870 , y2871 , y2872 , y2873 , y2874 , y2875 , y2876 , y2877 , y2878 , y2879 , y2880 , y2881 , y2882 , y2883 , y2884 , y2885 , y2886 , y2887 , y2888 , y2889 , y2890 , y2891 , y2892 , y2893 , y2894 , y2895 , y2896 , y2897 , y2898 , y2899 , y2900 , y2901 , y2902 , y2903 , y2904 , y2905 , y2906 , y2907 , y2908 , y2909 , y2910 , y2911 , y2912 , y2913 , y2914 , y2915 , y2916 , y2917 , y2918 , y2919 , y2920 , y2921 , y2922 , y2923 , y2924 , y2925 , y2926 , y2927 , y2928 , y2929 , y2930 , y2931 , y2932 , y2933 , y2934 , y2935 , y2936 , y2937 , y2938 , y2939 , y2940 , y2941 , y2942 , y2943 , y2944 , y2945 , y2946 , y2947 , y2948 , y2949 , y2950 , y2951 , y2952 , y2953 , y2954 , y2955 , y2956 , y2957 , y2958 , y2959 , y2960 , y2961 , y2962 , y2963 , y2964 , y2965 , y2966 , y2967 , y2968 , y2969 , y2970 , y2971 , y2972 , y2973 , y2974 , y2975 , y2976 , y2977 , y2978 , y2979 , y2980 , y2981 , y2982 , y2983 , y2984 , y2985 , y2986 , y2987 , y2988 , y2989 , y2990 , y2991 , y2992 , y2993 , y2994 , y2995 , y2996 , y2997 , y2998 , y2999 , y3000 , y3001 , y3002 , y3003 , y3004 , y3005 , y3006 , y3007 , y3008 , y3009 , y3010 , y3011 , y3012 , y3013 , y3014 , y3015 , y3016 , y3017 , y3018 , y3019 , y3020 , y3021 , y3022 , y3023 , y3024 , y3025 , y3026 , y3027 , y3028 , y3029 , y3030 , y3031 , y3032 , y3033 , y3034 , y3035 , y3036 , y3037 , y3038 , y3039 , y3040 , y3041 , y3042 , y3043 , y3044 , y3045 , y3046 , y3047 , y3048 , y3049 , y3050 , y3051 , y3052 , y3053 , y3054 , y3055 , y3056 , y3057 , y3058 , y3059 , y3060 , y3061 , y3062 , y3063 , y3064 , y3065 , y3066 , y3067 , y3068 , y3069 , y3070 , y3071 , y3072 , y3073 , y3074 , y3075 , y3076 , y3077 , y3078 , y3079 , y3080 , y3081 , y3082 , y3083 , y3084 , y3085 , y3086 , y3087 , y3088 , y3089 , y3090 , y3091 , y3092 , y3093 , y3094 , y3095 , y3096 , y3097 , y3098 , y3099 , y3100 , y3101 , y3102 , y3103 , y3104 , y3105 , y3106 , y3107 , y3108 , y3109 , y3110 , y3111 , y3112 , y3113 , y3114 , y3115 , y3116 , y3117 , y3118 , y3119 , y3120 , y3121 , y3122 , y3123 , y3124 , y3125 , y3126 , y3127 , y3128 , y3129 , y3130 , y3131 , y3132 , y3133 , y3134 , y3135 , y3136 , y3137 , y3138 , y3139 , y3140 , y3141 , y3142 , y3143 , y3144 , y3145 , y3146 , y3147 , y3148 , y3149 , y3150 , y3151 , y3152 , y3153 , y3154 , y3155 , y3156 , y3157 , y3158 , y3159 , y3160 , y3161 , y3162 , y3163 , y3164 , y3165 , y3166 , y3167 , y3168 , y3169 , y3170 , y3171 , y3172 , y3173 , y3174 , y3175 , y3176 , y3177 , y3178 , y3179 , y3180 , y3181 , y3182 , y3183 , y3184 , y3185 , y3186 , y3187 , y3188 , y3189 , y3190 , y3191 , y3192 , y3193 , y3194 , y3195 , y3196 , y3197 , y3198 , y3199 , y3200 , y3201 , y3202 , y3203 , y3204 , y3205 , y3206 , y3207 , y3208 , y3209 , y3210 , y3211 , y3212 , y3213 , y3214 , y3215 , y3216 , y3217 , y3218 , y3219 , y3220 , y3221 , y3222 , y3223 , y3224 , y3225 , y3226 , y3227 , y3228 , y3229 , y3230 , y3231 , y3232 , y3233 , y3234 , y3235 , y3236 , y3237 , y3238 , y3239 , y3240 , y3241 , y3242 , y3243 , y3244 , y3245 , y3246 , y3247 , y3248 , y3249 , y3250 , y3251 , y3252 , y3253 , y3254 , y3255 , y3256 , y3257 , y3258 , y3259 , y3260 , y3261 , y3262 , y3263 , y3264 , y3265 , y3266 , y3267 , y3268 , y3269 , y3270 , y3271 , y3272 , y3273 , y3274 , y3275 , y3276 , y3277 , y3278 , y3279 , y3280 , y3281 , y3282 , y3283 , y3284 , y3285 , y3286 , y3287 , y3288 , y3289 , y3290 , y3291 , y3292 , y3293 , y3294 , y3295 , y3296 , y3297 , y3298 , y3299 , y3300 , y3301 , y3302 , y3303 , y3304 , y3305 , y3306 , y3307 , y3308 , y3309 , y3310 , y3311 , y3312 , y3313 , y3314 , y3315 , y3316 , y3317 , y3318 , y3319 , y3320 , y3321 , y3322 , y3323 , y3324 , y3325 , y3326 , y3327 , y3328 , y3329 , y3330 , y3331 , y3332 , y3333 , y3334 , y3335 , y3336 , y3337 , y3338 , y3339 , y3340 , y3341 , y3342 , y3343 , y3344 , y3345 , y3346 , y3347 , y3348 , y3349 , y3350 , y3351 , y3352 , y3353 , y3354 , y3355 , y3356 , y3357 , y3358 , y3359 , y3360 , y3361 , y3362 , y3363 , y3364 , y3365 , y3366 , y3367 , y3368 , y3369 , y3370 , y3371 , y3372 , y3373 , y3374 , y3375 , y3376 , y3377 , y3378 , y3379 , y3380 , y3381 , y3382 , y3383 , y3384 , y3385 , y3386 , y3387 , y3388 , y3389 , y3390 , y3391 , y3392 , y3393 , y3394 , y3395 , y3396 , y3397 , y3398 , y3399 , y3400 , y3401 , y3402 , y3403 , y3404 , y3405 , y3406 , y3407 , y3408 , y3409 , y3410 , y3411 , y3412 , y3413 , y3414 , y3415 , y3416 , y3417 , y3418 , y3419 , y3420 , y3421 , y3422 , y3423 , y3424 , y3425 , y3426 , y3427 , y3428 , y3429 , y3430 , y3431 , y3432 , y3433 , y3434 , y3435 , y3436 , y3437 , y3438 , y3439 , y3440 , y3441 , y3442 , y3443 , y3444 , y3445 , y3446 , y3447 , y3448 , y3449 , y3450 , y3451 , y3452 , y3453 , y3454 , y3455 , y3456 , y3457 , y3458 , y3459 , y3460 , y3461 , y3462 , y3463 , y3464 , y3465 , y3466 , y3467 , y3468 , y3469 , y3470 , y3471 , y3472 , y3473 , y3474 , y3475 , y3476 , y3477 , y3478 , y3479 , y3480 , y3481 , y3482 , y3483 , y3484 , y3485 , y3486 , y3487 , y3488 , y3489 , y3490 , y3491 , y3492 , y3493 , y3494 , y3495 , y3496 , y3497 , y3498 , y3499 , y3500 , y3501 , y3502 , y3503 , y3504 , y3505 , y3506 , y3507 , y3508 , y3509 , y3510 , y3511 , y3512 , y3513 , y3514 , y3515 , y3516 , y3517 , y3518 , y3519 , y3520 , y3521 , y3522 , y3523 , y3524 , y3525 , y3526 , y3527 , y3528 , y3529 , y3530 , y3531 , y3532 , y3533 , y3534 , y3535 , y3536 , y3537 , y3538 , y3539 , y3540 , y3541 , y3542 , y3543 , y3544 , y3545 , y3546 , y3547 , y3548 , y3549 , y3550 , y3551 , y3552 , y3553 , y3554 , y3555 , y3556 , y3557 , y3558 , y3559 , y3560 , y3561 , y3562 , y3563 , y3564 , y3565 , y3566 , y3567 , y3568 , y3569 , y3570 , y3571 , y3572 , y3573 , y3574 , y3575 , y3576 , y3577 , y3578 , y3579 , y3580 , y3581 , y3582 , y3583 , y3584 , y3585 , y3586 , y3587 , y3588 , y3589 , y3590 , y3591 , y3592 , y3593 , y3594 , y3595 , y3596 , y3597 , y3598 , y3599 , y3600 , y3601 , y3602 , y3603 , y3604 , y3605 , y3606 , y3607 , y3608 , y3609 , y3610 , y3611 , y3612 , y3613 , y3614 , y3615 , y3616 , y3617 , y3618 , y3619 , y3620 , y3621 , y3622 , y3623 , y3624 , y3625 , y3626 , y3627 , y3628 , y3629 , y3630 , y3631 , y3632 , y3633 , y3634 , y3635 , y3636 , y3637 , y3638 , y3639 , y3640 , y3641 , y3642 , y3643 , y3644 , y3645 , y3646 , y3647 , y3648 , y3649 , y3650 , y3651 , y3652 , y3653 , y3654 , y3655 , y3656 , y3657 , y3658 , y3659 , y3660 , y3661 , y3662 , y3663 , y3664 , y3665 , y3666 , y3667 , y3668 , y3669 , y3670 , y3671 , y3672 , y3673 , y3674 , y3675 , y3676 , y3677 , y3678 , y3679 , y3680 , y3681 , y3682 , y3683 , y3684 , y3685 , y3686 , y3687 , y3688 , y3689 , y3690 , y3691 , y3692 , y3693 , y3694 , y3695 , y3696 , y3697 , y3698 , y3699 , y3700 , y3701 , y3702 , y3703 , y3704 , y3705 , y3706 , y3707 , y3708 , y3709 , y3710 , y3711 , y3712 , y3713 , y3714 , y3715 , y3716 , y3717 , y3718 , y3719 , y3720 , y3721 , y3722 , y3723 , y3724 , y3725 , y3726 , y3727 , y3728 , y3729 , y3730 , y3731 , y3732 , y3733 , y3734 , y3735 , y3736 , y3737 , y3738 , y3739 , y3740 , y3741 , y3742 , y3743 , y3744 , y3745 , y3746 , y3747 , y3748 , y3749 , y3750 , y3751 , y3752 , y3753 , y3754 , y3755 , y3756 , y3757 , y3758 , y3759 , y3760 , y3761 , y3762 , y3763 , y3764 , y3765 , y3766 , y3767 , y3768 , y3769 , y3770 , y3771 , y3772 , y3773 , y3774 , y3775 , y3776 , y3777 , y3778 , y3779 , y3780 , y3781 , y3782 , y3783 , y3784 , y3785 , y3786 , y3787 , y3788 , y3789 , y3790 , y3791 , y3792 , y3793 , y3794 , y3795 , y3796 , y3797 , y3798 , y3799 , y3800 , y3801 , y3802 , y3803 , y3804 , y3805 , y3806 , y3807 , y3808 , y3809 , y3810 , y3811 , y3812 , y3813 , y3814 , y3815 , y3816 , y3817 , y3818 , y3819 , y3820 , y3821 , y3822 , y3823 , y3824 , y3825 , y3826 , y3827 , y3828 , y3829 , y3830 , y3831 , y3832 , y3833 , y3834 , y3835 , y3836 , y3837 , y3838 , y3839 , y3840 , y3841 , y3842 , y3843 , y3844 , y3845 , y3846 , y3847 , y3848 , y3849 , y3850 , y3851 , y3852 , y3853 , y3854 , y3855 , y3856 , y3857 , y3858 , y3859 , y3860 , y3861 , y3862 , y3863 , y3864 , y3865 , y3866 , y3867 , y3868 , y3869 , y3870 , y3871 , y3872 , y3873 , y3874 , y3875 , y3876 , y3877 , y3878 , y3879 , y3880 , y3881 , y3882 , y3883 , y3884 , y3885 , y3886 , y3887 , y3888 , y3889 , y3890 , y3891 , y3892 , y3893 , y3894 , y3895 , y3896 , y3897 , y3898 , y3899 , y3900 , y3901 , y3902 , y3903 , y3904 , y3905 , y3906 , y3907 , y3908 , y3909 , y3910 , y3911 , y3912 , y3913 , y3914 , y3915 , y3916 , y3917 , y3918 , y3919 , y3920 , y3921 , y3922 , y3923 , y3924 , y3925 , y3926 , y3927 , y3928 , y3929 , y3930 , y3931 , y3932 , y3933 , y3934 , y3935 , y3936 , y3937 , y3938 , y3939 , y3940 , y3941 , y3942 , y3943 , y3944 , y3945 , y3946 , y3947 , y3948 , y3949 , y3950 , y3951 , y3952 , y3953 , y3954 , y3955 , y3956 , y3957 , y3958 , y3959 , y3960 , y3961 , y3962 , y3963 , y3964 , y3965 , y3966 , y3967 , y3968 , y3969 , y3970 , y3971 , y3972 , y3973 , y3974 , y3975 , y3976 , y3977 , y3978 , y3979 , y3980 , y3981 , y3982 , y3983 , y3984 , y3985 , y3986 , y3987 , y3988 , y3989 , y3990 , y3991 , y3992 , y3993 , y3994 , y3995 , y3996 , y3997 , y3998 , y3999 , y4000 , y4001 , y4002 , y4003 , y4004 , y4005 , y4006 , y4007 , y4008 , y4009 , y4010 , y4011 , y4012 , y4013 , y4014 , y4015 , y4016 , y4017 , y4018 , y4019 , y4020 , y4021 , y4022 , y4023 , y4024 , y4025 , y4026 , y4027 , y4028 , y4029 , y4030 , y4031 , y4032 , y4033 , y4034 , y4035 , y4036 , y4037 , y4038 , y4039 , y4040 , y4041 , y4042 , y4043 , y4044 , y4045 , y4046 , y4047 , y4048 , y4049 , y4050 , y4051 , y4052 , y4053 , y4054 , y4055 , y4056 , y4057 , y4058 , y4059 , y4060 , y4061 , y4062 , y4063 , y4064 , y4065 , y4066 , y4067 , y4068 , y4069 , y4070 , y4071 , y4072 , y4073 , y4074 , y4075 , y4076 , y4077 , y4078 , y4079 , y4080 , y4081 , y4082 , y4083 , y4084 , y4085 , y4086 , y4087 , y4088 , y4089 , y4090 , y4091 , y4092 , y4093 , y4094 , y4095 , y4096 , y4097 , y4098 , y4099 , y4100 , y4101 , y4102 , y4103 , y4104 , y4105 , y4106 , y4107 , y4108 , y4109 , y4110 , y4111 , y4112 , y4113 , y4114 , y4115 , y4116 , y4117 , y4118 , y4119 , y4120 , y4121 , y4122 , y4123 , y4124 , y4125 , y4126 , y4127 , y4128 , y4129 , y4130 , y4131 , y4132 , y4133 , y4134 , y4135 , y4136 , y4137 , y4138 , y4139 , y4140 , y4141 , y4142 , y4143 , y4144 , y4145 , y4146 , y4147 , y4148 , y4149 , y4150 , y4151 , y4152 , y4153 , y4154 , y4155 , y4156 , y4157 , y4158 , y4159 , y4160 , y4161 , y4162 , y4163 , y4164 , y4165 , y4166 , y4167 , y4168 , y4169 , y4170 , y4171 , y4172 , y4173 , y4174 , y4175 , y4176 , y4177 , y4178 , y4179 , y4180 , y4181 , y4182 , y4183 , y4184 , y4185 , y4186 , y4187 , y4188 , y4189 , y4190 , y4191 , y4192 , y4193 , y4194 , y4195 , y4196 , y4197 , y4198 , y4199 , y4200 , y4201 , y4202 , y4203 , y4204 , y4205 , y4206 , y4207 , y4208 , y4209 , y4210 , y4211 , y4212 , y4213 , y4214 , y4215 , y4216 , y4217 , y4218 , y4219 , y4220 , y4221 , y4222 , y4223 , y4224 , y4225 , y4226 , y4227 , y4228 , y4229 , y4230 , y4231 , y4232 , y4233 , y4234 , y4235 , y4236 , y4237 , y4238 , y4239 , y4240 , y4241 , y4242 , y4243 , y4244 , y4245 , y4246 , y4247 , y4248 , y4249 , y4250 , y4251 , y4252 , y4253 , y4254 , y4255 , y4256 , y4257 , y4258 , y4259 , y4260 , y4261 , y4262 , y4263 , y4264 , y4265 , y4266 , y4267 , y4268 , y4269 , y4270 , y4271 , y4272 , y4273 , y4274 , y4275 , y4276 , y4277 , y4278 , y4279 , y4280 , y4281 , y4282 , y4283 , y4284 , y4285 , y4286 , y4287 , y4288 , y4289 , y4290 , y4291 , y4292 , y4293 , y4294 , y4295 , y4296 , y4297 , y4298 , y4299 , y4300 , y4301 , y4302 , y4303 , y4304 , y4305 , y4306 , y4307 , y4308 , y4309 , y4310 , y4311 , y4312 , y4313 , y4314 , y4315 , y4316 , y4317 , y4318 , y4319 , y4320 , y4321 , y4322 , y4323 , y4324 , y4325 , y4326 , y4327 , y4328 , y4329 , y4330 , y4331 , y4332 , y4333 , y4334 , y4335 , y4336 , y4337 , y4338 , y4339 , y4340 , y4341 , y4342 , y4343 , y4344 , y4345 , y4346 , y4347 , y4348 , y4349 , y4350 , y4351 , y4352 , y4353 , y4354 , y4355 , y4356 , y4357 , y4358 , y4359 , y4360 , y4361 , y4362 , y4363 , y4364 , y4365 , y4366 , y4367 , y4368 , y4369 , y4370 , y4371 , y4372 , y4373 , y4374 , y4375 , y4376 , y4377 , y4378 , y4379 , y4380 , y4381 , y4382 , y4383 , y4384 , y4385 , y4386 , y4387 , y4388 , y4389 , y4390 , y4391 , y4392 , y4393 , y4394 , y4395 , y4396 , y4397 , y4398 , y4399 , y4400 , y4401 , y4402 , y4403 , y4404 , y4405 , y4406 , y4407 , y4408 , y4409 , y4410 , y4411 , y4412 , y4413 , y4414 , y4415 , y4416 , y4417 , y4418 , y4419 , y4420 , y4421 , y4422 , y4423 , y4424 , y4425 , y4426 , y4427 , y4428 , y4429 , y4430 , y4431 , y4432 , y4433 , y4434 , y4435 , y4436 , y4437 , y4438 , y4439 , y4440 , y4441 , y4442 , y4443 , y4444 , y4445 , y4446 , y4447 , y4448 , y4449 , y4450 , y4451 , y4452 , y4453 , y4454 , y4455 , y4456 , y4457 , y4458 , y4459 , y4460 , y4461 , y4462 , y4463 , y4464 , y4465 , y4466 , y4467 , y4468 , y4469 , y4470 , y4471 , y4472 , y4473 , y4474 , y4475 , y4476 , y4477 , y4478 , y4479 , y4480 , y4481 , y4482 , y4483 , y4484 , y4485 , y4486 , y4487 , y4488 , y4489 , y4490 , y4491 , y4492 , y4493 , y4494 , y4495 , y4496 , y4497 , y4498 , y4499 , y4500 , y4501 , y4502 , y4503 , y4504 , y4505 , y4506 , y4507 , y4508 , y4509 , y4510 , y4511 , y4512 , y4513 , y4514 , y4515 , y4516 , y4517 , y4518 , y4519 , y4520 , y4521 , y4522 , y4523 , y4524 , y4525 , y4526 , y4527 , y4528 , y4529 , y4530 , y4531 , y4532 , y4533 , y4534 , y4535 , y4536 , y4537 , y4538 , y4539 , y4540 , y4541 , y4542 , y4543 , y4544 , y4545 , y4546 , y4547 , y4548 , y4549 , y4550 , y4551 , y4552 , y4553 , y4554 , y4555 , y4556 , y4557 , y4558 , y4559 , y4560 , y4561 , y4562 , y4563 , y4564 , y4565 , y4566 , y4567 , y4568 , y4569 , y4570 , y4571 , y4572 , y4573 , y4574 , y4575 , y4576 , y4577 , y4578 , y4579 , y4580 , y4581 , y4582 , y4583 , y4584 , y4585 , y4586 , y4587 , y4588 , y4589 , y4590 , y4591 , y4592 , y4593 , y4594 , y4595 , y4596 , y4597 , y4598 , y4599 , y4600 , y4601 , y4602 , y4603 , y4604 , y4605 , y4606 , y4607 , y4608 , y4609 , y4610 , y4611 , y4612 , y4613 , y4614 , y4615 , y4616 , y4617 , y4618 , y4619 , y4620 , y4621 , y4622 , y4623 , y4624 , y4625 , y4626 , y4627 , y4628 , y4629 , y4630 , y4631 , y4632 , y4633 , y4634 , y4635 , y4636 , y4637 , y4638 , y4639 , y4640 , y4641 , y4642 , y4643 , y4644 , y4645 , y4646 , y4647 , y4648 , y4649 , y4650 , y4651 , y4652 , y4653 , y4654 , y4655 , y4656 , y4657 , y4658 , y4659 , y4660 , y4661 , y4662 , y4663 , y4664 , y4665 , y4666 , y4667 , y4668 , y4669 , y4670 , y4671 , y4672 , y4673 , y4674 , y4675 , y4676 , y4677 , y4678 , y4679 , y4680 , y4681 , y4682 , y4683 , y4684 , y4685 , y4686 , y4687 , y4688 , y4689 , y4690 , y4691 , y4692 , y4693 , y4694 , y4695 , y4696 , y4697 , y4698 , y4699 , y4700 , y4701 , y4702 , y4703 , y4704 , y4705 , y4706 , y4707 , y4708 , y4709 , y4710 , y4711 , y4712 , y4713 , y4714 , y4715 , y4716 , y4717 , y4718 , y4719 , y4720 , y4721 , y4722 , y4723 , y4724 , y4725 , y4726 , y4727 , y4728 , y4729 , y4730 , y4731 , y4732 , y4733 , y4734 , y4735 , y4736 , y4737 , y4738 , y4739 , y4740 , y4741 , y4742 , y4743 , y4744 , y4745 , y4746 , y4747 , y4748 , y4749 , y4750 , y4751 , y4752 , y4753 , y4754 , y4755 , y4756 , y4757 , y4758 , y4759 , y4760 , y4761 , y4762 , y4763 , y4764 , y4765 , y4766 , y4767 , y4768 , y4769 , y4770 , y4771 , y4772 , y4773 , y4774 , y4775 , y4776 , y4777 , y4778 , y4779 , y4780 , y4781 , y4782 , y4783 , y4784 , y4785 , y4786 , y4787 , y4788 , y4789 , y4790 , y4791 , y4792 , y4793 , y4794 , y4795 , y4796 , y4797 , y4798 , y4799 , y4800 , y4801 , y4802 , y4803 , y4804 , y4805 , y4806 , y4807 , y4808 , y4809 , y4810 , y4811 , y4812 , y4813 , y4814 , y4815 , y4816 , y4817 , y4818 , y4819 , y4820 , y4821 , y4822 , y4823 , y4824 , y4825 , y4826 , y4827 , y4828 , y4829 , y4830 , y4831 , y4832 , y4833 , y4834 , y4835 , y4836 , y4837 , y4838 , y4839 , y4840 , y4841 , y4842 , y4843 , y4844 , y4845 , y4846 , y4847 , y4848 , y4849 , y4850 , y4851 , y4852 , y4853 , y4854 , y4855 , y4856 , y4857 , y4858 , y4859 , y4860 , y4861 , y4862 , y4863 , y4864 , y4865 , y4866 , y4867 , y4868 , y4869 , y4870 , y4871 , y4872 , y4873 , y4874 , y4875 , y4876 , y4877 , y4878 , y4879 , y4880 , y4881 , y4882 , y4883 , y4884 , y4885 , y4886 , y4887 , y4888 , y4889 , y4890 , y4891 , y4892 , y4893 , y4894 , y4895 , y4896 , y4897 , y4898 , y4899 , y4900 , y4901 , y4902 , y4903 , y4904 , y4905 , y4906 , y4907 , y4908 , y4909 , y4910 , y4911 , y4912 , y4913 , y4914 , y4915 , y4916 , y4917 , y4918 , y4919 , y4920 , y4921 , y4922 , y4923 , y4924 , y4925 , y4926 , y4927 , y4928 , y4929 , y4930 , y4931 , y4932 , y4933 , y4934 , y4935 , y4936 , y4937 , y4938 , y4939 , y4940 , y4941 , y4942 , y4943 , y4944 , y4945 , y4946 , y4947 , y4948 , y4949 , y4950 , y4951 , y4952 , y4953 , y4954 , y4955 , y4956 , y4957 , y4958 , y4959 , y4960 , y4961 , y4962 , y4963 , y4964 , y4965 , y4966 , y4967 , y4968 , y4969 , y4970 , y4971 , y4972 , y4973 , y4974 , y4975 , y4976 , y4977 , y4978 , y4979 , y4980 , y4981 , y4982 , y4983 , y4984 , y4985 , y4986 , y4987 , y4988 , y4989 , y4990 , y4991 , y4992 , y4993 , y4994 , y4995 , y4996 , y4997 , y4998 , y4999 , y5000 , y5001 , y5002 , y5003 , y5004 , y5005 , y5006 , y5007 , y5008 , y5009 , y5010 , y5011 , y5012 , y5013 , y5014 , y5015 , y5016 , y5017 , y5018 , y5019 , y5020 , y5021 , y5022 , y5023 , y5024 , y5025 , y5026 , y5027 , y5028 , y5029 , y5030 , y5031 , y5032 , y5033 , y5034 , y5035 , y5036 , y5037 , y5038 , y5039 , y5040 , y5041 , y5042 , y5043 , y5044 , y5045 , y5046 , y5047 , y5048 , y5049 , y5050 , y5051 , y5052 , y5053 , y5054 , y5055 , y5056 , y5057 , y5058 , y5059 , y5060 , y5061 , y5062 , y5063 , y5064 , y5065 , y5066 , y5067 , y5068 , y5069 , y5070 , y5071 , y5072 , y5073 , y5074 , y5075 , y5076 , y5077 , y5078 , y5079 , y5080 , y5081 , y5082 , y5083 , y5084 , y5085 , y5086 , y5087 , y5088 , y5089 , y5090 , y5091 , y5092 , y5093 , y5094 , y5095 , y5096 , y5097 , y5098 , y5099 , y5100 , y5101 , y5102 , y5103 , y5104 , y5105 , y5106 , y5107 , y5108 , y5109 , y5110 , y5111 , y5112 , y5113 , y5114 , y5115 , y5116 , y5117 , y5118 , y5119 , y5120 , y5121 , y5122 , y5123 , y5124 , y5125 , y5126 , y5127 , y5128 , y5129 , y5130 , y5131 , y5132 , y5133 , y5134 , y5135 , y5136 , y5137 , y5138 , y5139 , y5140 , y5141 , y5142 , y5143 , y5144 , y5145 , y5146 , y5147 , y5148 , y5149 , y5150 , y5151 , y5152 , y5153 , y5154 , y5155 , y5156 , y5157 , y5158 , y5159 , y5160 , y5161 , y5162 , y5163 , y5164 , y5165 , y5166 , y5167 , y5168 , y5169 , y5170 , y5171 , y5172 , y5173 , y5174 , y5175 , y5176 , y5177 , y5178 , y5179 , y5180 , y5181 , y5182 , y5183 , y5184 , y5185 , y5186 , y5187 , y5188 , y5189 , y5190 , y5191 , y5192 , y5193 , y5194 , y5195 , y5196 , y5197 , y5198 , y5199 , y5200 , y5201 , y5202 , y5203 , y5204 , y5205 , y5206 , y5207 , y5208 , y5209 , y5210 , y5211 , y5212 , y5213 , y5214 , y5215 , y5216 , y5217 , y5218 , y5219 , y5220 , y5221 , y5222 , y5223 , y5224 , y5225 , y5226 , y5227 , y5228 , y5229 , y5230 , y5231 , y5232 , y5233 , y5234 , y5235 , y5236 , y5237 , y5238 , y5239 , y5240 , y5241 , y5242 , y5243 , y5244 , y5245 , y5246 , y5247 , y5248 , y5249 , y5250 , y5251 , y5252 , y5253 , y5254 , y5255 , y5256 , y5257 , y5258 , y5259 , y5260 , y5261 , y5262 , y5263 , y5264 , y5265 , y5266 , y5267 , y5268 , y5269 , y5270 , y5271 , y5272 , y5273 , y5274 , y5275 , y5276 , y5277 , y5278 , y5279 , y5280 , y5281 , y5282 , y5283 , y5284 , y5285 , y5286 , y5287 , y5288 , y5289 , y5290 , y5291 , y5292 , y5293 , y5294 , y5295 , y5296 , y5297 , y5298 , y5299 , y5300 , y5301 , y5302 , y5303 , y5304 , y5305 , y5306 , y5307 , y5308 , y5309 , y5310 , y5311 , y5312 , y5313 , y5314 , y5315 , y5316 , y5317 , y5318 , y5319 , y5320 , y5321 , y5322 , y5323 , y5324 , y5325 , y5326 , y5327 , y5328 , y5329 , y5330 , y5331 , y5332 , y5333 , y5334 , y5335 , y5336 , y5337 , y5338 , y5339 , y5340 , y5341 , y5342 , y5343 , y5344 , y5345 , y5346 , y5347 , y5348 , y5349 , y5350 , y5351 , y5352 , y5353 , y5354 , y5355 , y5356 , y5357 , y5358 , y5359 , y5360 , y5361 , y5362 , y5363 , y5364 , y5365 , y5366 , y5367 , y5368 , y5369 , y5370 , y5371 , y5372 , y5373 , y5374 , y5375 , y5376 , y5377 , y5378 , y5379 , y5380 , y5381 , y5382 , y5383 , y5384 , y5385 , y5386 , y5387 , y5388 , y5389 , y5390 , y5391 , y5392 , y5393 , y5394 , y5395 , y5396 , y5397 , y5398 , y5399 , y5400 , y5401 , y5402 , y5403 , y5404 , y5405 , y5406 , y5407 , y5408 , y5409 , y5410 , y5411 , y5412 , y5413 , y5414 , y5415 , y5416 , y5417 , y5418 , y5419 , y5420 , y5421 , y5422 , y5423 , y5424 , y5425 , y5426 , y5427 , y5428 , y5429 , y5430 , y5431 , y5432 , y5433 , y5434 , y5435 , y5436 , y5437 , y5438 , y5439 , y5440 , y5441 , y5442 , y5443 , y5444 , y5445 , y5446 , y5447 , y5448 , y5449 , y5450 , y5451 , y5452 , y5453 , y5454 , y5455 , y5456 , y5457 , y5458 , y5459 , y5460 , y5461 , y5462 , y5463 , y5464 , y5465 , y5466 , y5467 , y5468 , y5469 , y5470 , y5471 , y5472 , y5473 , y5474 , y5475 , y5476 , y5477 , y5478 , y5479 , y5480 , y5481 , y5482 , y5483 , y5484 , y5485 , y5486 , y5487 , y5488 , y5489 , y5490 , y5491 , y5492 , y5493 , y5494 , y5495 , y5496 , y5497 , y5498 , y5499 , y5500 , y5501 , y5502 , y5503 , y5504 , y5505 , y5506 , y5507 , y5508 , y5509 , y5510 , y5511 , y5512 , y5513 , y5514 , y5515 , y5516 , y5517 , y5518 , y5519 , y5520 , y5521 , y5522 , y5523 , y5524 , y5525 , y5526 , y5527 , y5528 , y5529 , y5530 , y5531 , y5532 , y5533 , y5534 , y5535 , y5536 , y5537 , y5538 , y5539 , y5540 , y5541 , y5542 , y5543 , y5544 , y5545 , y5546 , y5547 , y5548 , y5549 , y5550 , y5551 , y5552 , y5553 , y5554 , y5555 , y5556 , y5557 , y5558 , y5559 , y5560 , y5561 , y5562 , y5563 , y5564 , y5565 , y5566 , y5567 , y5568 , y5569 , y5570 , y5571 , y5572 , y5573 , y5574 , y5575 , y5576 , y5577 , y5578 , y5579 , y5580 , y5581 , y5582 , y5583 , y5584 , y5585 , y5586 , y5587 , y5588 , y5589 , y5590 , y5591 , y5592 , y5593 , y5594 , y5595 , y5596 , y5597 , y5598 , y5599 , y5600 , y5601 , y5602 , y5603 , y5604 , y5605 , y5606 , y5607 , y5608 , y5609 , y5610 , y5611 , y5612 , y5613 , y5614 , y5615 , y5616 , y5617 , y5618 , y5619 , y5620 , y5621 , y5622 , y5623 , y5624 , y5625 , y5626 , y5627 , y5628 , y5629 , y5630 , y5631 , y5632 , y5633 , y5634 , y5635 , y5636 , y5637 , y5638 , y5639 , y5640 , y5641 , y5642 , y5643 , y5644 , y5645 , y5646 , y5647 , y5648 , y5649 , y5650 , y5651 , y5652 , y5653 , y5654 , y5655 , y5656 , y5657 , y5658 , y5659 , y5660 , y5661 , y5662 , y5663 , y5664 , y5665 , y5666 , y5667 , y5668 , y5669 , y5670 , y5671 , y5672 , y5673 , y5674 , y5675 , y5676 , y5677 , y5678 , y5679 , y5680 , y5681 , y5682 , y5683 , y5684 , y5685 , y5686 , y5687 , y5688 , y5689 , y5690 , y5691 , y5692 , y5693 , y5694 , y5695 , y5696 , y5697 , y5698 , y5699 , y5700 , y5701 , y5702 , y5703 , y5704 , y5705 , y5706 , y5707 , y5708 , y5709 , y5710 , y5711 , y5712 , y5713 , y5714 , y5715 , y5716 , y5717 , y5718 , y5719 , y5720 , y5721 , y5722 , y5723 , y5724 , y5725 , y5726 , y5727 , y5728 , y5729 , y5730 , y5731 , y5732 , y5733 , y5734 , y5735 , y5736 , y5737 , y5738 , y5739 , y5740 , y5741 , y5742 , y5743 , y5744 , y5745 , y5746 , y5747 , y5748 , y5749 , y5750 , y5751 , y5752 , y5753 , y5754 , y5755 , y5756 , y5757 , y5758 , y5759 , y5760 , y5761 , y5762 , y5763 , y5764 , y5765 , y5766 , y5767 , y5768 , y5769 , y5770 , y5771 , y5772 , y5773 , y5774 , y5775 , y5776 , y5777 , y5778 , y5779 , y5780 , y5781 , y5782 , y5783 , y5784 , y5785 , y5786 , y5787 , y5788 , y5789 , y5790 , y5791 , y5792 , y5793 , y5794 , y5795 , y5796 , y5797 , y5798 , y5799 , y5800 , y5801 , y5802 , y5803 , y5804 , y5805 , y5806 , y5807 , y5808 , y5809 , y5810 , y5811 , y5812 , y5813 , y5814 , y5815 , y5816 , y5817 , y5818 , y5819 , y5820 , y5821 , y5822 , y5823 , y5824 , y5825 , y5826 , y5827 , y5828 , y5829 , y5830 , y5831 , y5832 , y5833 , y5834 , y5835 , y5836 , y5837 , y5838 , y5839 , y5840 , y5841 , y5842 , y5843 , y5844 , y5845 , y5846 , y5847 , y5848 , y5849 , y5850 , y5851 , y5852 , y5853 , y5854 , y5855 , y5856 , y5857 , y5858 , y5859 , y5860 , y5861 , y5862 , y5863 , y5864 , y5865 , y5866 , y5867 , y5868 , y5869 , y5870 , y5871 , y5872 , y5873 , y5874 , y5875 , y5876 , y5877 , y5878 , y5879 , y5880 , y5881 , y5882 , y5883 , y5884 , y5885 , y5886 , y5887 , y5888 , y5889 , y5890 , y5891 , y5892 , y5893 , y5894 , y5895 , y5896 , y5897 , y5898 , y5899 , y5900 , y5901 , y5902 , y5903 , y5904 , y5905 , y5906 , y5907 , y5908 , y5909 , y5910 , y5911 , y5912 , y5913 , y5914 , y5915 , y5916 , y5917 , y5918 , y5919 , y5920 , y5921 , y5922 , y5923 , y5924 , y5925 , y5926 , y5927 , y5928 , y5929 , y5930 , y5931 , y5932 , y5933 , y5934 , y5935 , y5936 , y5937 , y5938 , y5939 , y5940 , y5941 , y5942 , y5943 , y5944 , y5945 , y5946 , y5947 , y5948 , y5949 , y5950 , y5951 , y5952 , y5953 , y5954 , y5955 , y5956 , y5957 , y5958 , y5959 , y5960 , y5961 , y5962 , y5963 , y5964 , y5965 , y5966 , y5967 , y5968 , y5969 , y5970 , y5971 , y5972 , y5973 , y5974 , y5975 , y5976 , y5977 , y5978 , y5979 , y5980 , y5981 , y5982 , y5983 , y5984 , y5985 , y5986 , y5987 , y5988 , y5989 , y5990 , y5991 , y5992 , y5993 , y5994 , y5995 , y5996 , y5997 , y5998 , y5999 , y6000 , y6001 , y6002 , y6003 , y6004 , y6005 , y6006 , y6007 , y6008 , y6009 , y6010 , y6011 , y6012 , y6013 , y6014 , y6015 , y6016 , y6017 , y6018 , y6019 , y6020 , y6021 , y6022 , y6023 , y6024 , y6025 , y6026 , y6027 , y6028 , y6029 , y6030 , y6031 , y6032 , y6033 , y6034 , y6035 , y6036 , y6037 , y6038 , y6039 , y6040 , y6041 , y6042 , y6043 , y6044 , y6045 , y6046 , y6047 , y6048 , y6049 , y6050 , y6051 , y6052 , y6053 , y6054 , y6055 , y6056 , y6057 , y6058 , y6059 , y6060 , y6061 , y6062 , y6063 , y6064 , y6065 , y6066 , y6067 , y6068 , y6069 , y6070 , y6071 , y6072 , y6073 , y6074 , y6075 , y6076 , y6077 , y6078 , y6079 , y6080 , y6081 , y6082 , y6083 , y6084 , y6085 , y6086 , y6087 , y6088 , y6089 , y6090 , y6091 , y6092 , y6093 , y6094 , y6095 , y6096 , y6097 , y6098 , y6099 , y6100 , y6101 , y6102 , y6103 , y6104 , y6105 , y6106 , y6107 , y6108 , y6109 , y6110 , y6111 , y6112 , y6113 , y6114 , y6115 , y6116 , y6117 , y6118 , y6119 , y6120 , y6121 , y6122 , y6123 , y6124 , y6125 , y6126 , y6127 , y6128 , y6129 , y6130 , y6131 , y6132 , y6133 , y6134 , y6135 , y6136 , y6137 , y6138 , y6139 , y6140 , y6141 , y6142 , y6143 , y6144 , y6145 , y6146 , y6147 , y6148 , y6149 , y6150 , y6151 , y6152 , y6153 , y6154 , y6155 , y6156 , y6157 , y6158 , y6159 , y6160 , y6161 , y6162 , y6163 , y6164 , y6165 , y6166 , y6167 , y6168 , y6169 , y6170 , y6171 , y6172 , y6173 , y6174 , y6175 , y6176 , y6177 , y6178 , y6179 , y6180 , y6181 , y6182 , y6183 , y6184 , y6185 , y6186 , y6187 , y6188 , y6189 , y6190 , y6191 , y6192 , y6193 , y6194 , y6195 , y6196 , y6197 , y6198 , y6199 , y6200 , y6201 , y6202 , y6203 , y6204 , y6205 , y6206 , y6207 , y6208 , y6209 , y6210 , y6211 , y6212 , y6213 , y6214 , y6215 , y6216 , y6217 , y6218 , y6219 , y6220 , y6221 , y6222 , y6223 , y6224 , y6225 , y6226 , y6227 , y6228 , y6229 , y6230 , y6231 , y6232 , y6233 , y6234 , y6235 , y6236 , y6237 , y6238 , y6239 , y6240 , y6241 , y6242 , y6243 , y6244 , y6245 , y6246 , y6247 , y6248 , y6249 , y6250 , y6251 , y6252 , y6253 , y6254 , y6255 , y6256 , y6257 , y6258 , y6259 , y6260 , y6261 , y6262 , y6263 , y6264 , y6265 , y6266 , y6267 , y6268 , y6269 , y6270 , y6271 , y6272 , y6273 , y6274 , y6275 , y6276 , y6277 , y6278 , y6279 , y6280 , y6281 , y6282 , y6283 , y6284 , y6285 , y6286 , y6287 , y6288 , y6289 , y6290 , y6291 , y6292 , y6293 , y6294 , y6295 , y6296 , y6297 , y6298 , y6299 , y6300 , y6301 , y6302 , y6303 , y6304 , y6305 , y6306 , y6307 , y6308 , y6309 , y6310 , y6311 , y6312 , y6313 , y6314 , y6315 , y6316 , y6317 , y6318 , y6319 , y6320 , y6321 , y6322 , y6323 , y6324 , y6325 , y6326 , y6327 , y6328 , y6329 , y6330 , y6331 , y6332 , y6333 , y6334 , y6335 , y6336 , y6337 , y6338 , y6339 , y6340 , y6341 , y6342 , y6343 , y6344 , y6345 , y6346 , y6347 , y6348 , y6349 , y6350 , y6351 , y6352 , y6353 , y6354 , y6355 , y6356 , y6357 , y6358 , y6359 , y6360 , y6361 , y6362 , y6363 , y6364 , y6365 , y6366 , y6367 , y6368 , y6369 , y6370 , y6371 , y6372 , y6373 , y6374 , y6375 , y6376 , y6377 , y6378 , y6379 , y6380 , y6381 , y6382 , y6383 , y6384 , y6385 , y6386 , y6387 , y6388 , y6389 , y6390 , y6391 , y6392 , y6393 , y6394 , y6395 , y6396 , y6397 , y6398 , y6399 , y6400 , y6401 , y6402 , y6403 , y6404 , y6405 , y6406 , y6407 , y6408 , y6409 , y6410 , y6411 , y6412 , y6413 , y6414 , y6415 , y6416 , y6417 , y6418 , y6419 , y6420 , y6421 , y6422 , y6423 , y6424 , y6425 , y6426 , y6427 , y6428 , y6429 , y6430 , y6431 , y6432 , y6433 , y6434 , y6435 , y6436 , y6437 , y6438 , y6439 , y6440 , y6441 , y6442 , y6443 , y6444 , y6445 , y6446 , y6447 , y6448 , y6449 , y6450 , y6451 , y6452 , y6453 , y6454 , y6455 , y6456 , y6457 , y6458 , y6459 , y6460 , y6461 , y6462 , y6463 , y6464 , y6465 , y6466 , y6467 , y6468 , y6469 , y6470 , y6471 , y6472 , y6473 , y6474 , y6475 , y6476 , y6477 , y6478 , y6479 , y6480 , y6481 , y6482 , y6483 , y6484 , y6485 , y6486 , y6487 , y6488 , y6489 , y6490 , y6491 , y6492 , y6493 , y6494 , y6495 , y6496 , y6497 , y6498 , y6499 , y6500 , y6501 , y6502 , y6503 , y6504 , y6505 , y6506 , y6507 , y6508 , y6509 , y6510 , y6511 , y6512 , y6513 , y6514 , y6515 , y6516 , y6517 , y6518 , y6519 , y6520 , y6521 , y6522 , y6523 , y6524 , y6525 , y6526 , y6527 , y6528 , y6529 , y6530 , y6531 , y6532 , y6533 , y6534 , y6535 , y6536 , y6537 , y6538 , y6539 , y6540 , y6541 , y6542 , y6543 , y6544 , y6545 , y6546 , y6547 , y6548 , y6549 , y6550 , y6551 , y6552 , y6553 , y6554 , y6555 , y6556 , y6557 , y6558 , y6559 , y6560 , y6561 , y6562 , y6563 , y6564 , y6565 , y6566 , y6567 , y6568 , y6569 , y6570 , y6571 , y6572 , y6573 , y6574 , y6575 , y6576 , y6577 , y6578 , y6579 , y6580 , y6581 , y6582 , y6583 , y6584 , y6585 , y6586 , y6587 , y6588 , y6589 , y6590 , y6591 , y6592 , y6593 , y6594 , y6595 , y6596 , y6597 , y6598 , y6599 , y6600 , y6601 , y6602 , y6603 , y6604 , y6605 , y6606 , y6607 , y6608 , y6609 , y6610 , y6611 , y6612 , y6613 , y6614 , y6615 , y6616 , y6617 , y6618 , y6619 , y6620 , y6621 , y6622 , y6623 , y6624 , y6625 , y6626 , y6627 , y6628 , y6629 , y6630 , y6631 , y6632 , y6633 , y6634 , y6635 , y6636 , y6637 , y6638 , y6639 , y6640 , y6641 , y6642 , y6643 , y6644 , y6645 , y6646 , y6647 , y6648 , y6649 , y6650 , y6651 , y6652 , y6653 , y6654 , y6655 , y6656 , y6657 , y6658 , y6659 , y6660 , y6661 , y6662 , y6663 , y6664 , y6665 , y6666 , y6667 , y6668 , y6669 , y6670 , y6671 , y6672 , y6673 , y6674 , y6675 , y6676 , y6677 , y6678 , y6679 , y6680 , y6681 , y6682 , y6683 , y6684 , y6685 , y6686 , y6687 , y6688 , y6689 , y6690 , y6691 , y6692 , y6693 , y6694 , y6695 , y6696 , y6697 , y6698 , y6699 , y6700 , y6701 , y6702 , y6703 , y6704 , y6705 , y6706 , y6707 , y6708 , y6709 , y6710 , y6711 , y6712 , y6713 , y6714 , y6715 , y6716 , y6717 , y6718 , y6719 , y6720 , y6721 , y6722 , y6723 , y6724 , y6725 , y6726 , y6727 , y6728 , y6729 , y6730 , y6731 , y6732 , y6733 , y6734 , y6735 , y6736 , y6737 , y6738 , y6739 , y6740 , y6741 , y6742 , y6743 , y6744 , y6745 , y6746 , y6747 , y6748 , y6749 , y6750 , y6751 , y6752 , y6753 , y6754 , y6755 , y6756 , y6757 , y6758 , y6759 , y6760 , y6761 , y6762 , y6763 , y6764 , y6765 , y6766 , y6767 , y6768 , y6769 , y6770 , y6771 , y6772 , y6773 , y6774 , y6775 , y6776 , y6777 , y6778 , y6779 , y6780 , y6781 , y6782 , y6783 , y6784 , y6785 , y6786 , y6787 , y6788 , y6789 , y6790 , y6791 , y6792 , y6793 , y6794 , y6795 , y6796 , y6797 , y6798 , y6799 , y6800 , y6801 , y6802 , y6803 , y6804 , y6805 , y6806 , y6807 , y6808 , y6809 , y6810 , y6811 , y6812 , y6813 , y6814 , y6815 , y6816 , y6817 , y6818 , y6819 , y6820 , y6821 , y6822 , y6823 , y6824 , y6825 , y6826 , y6827 , y6828 , y6829 , y6830 , y6831 , y6832 , y6833 , y6834 , y6835 , y6836 , y6837 , y6838 , y6839 , y6840 , y6841 , y6842 , y6843 , y6844 , y6845 , y6846 , y6847 , y6848 , y6849 , y6850 , y6851 , y6852 , y6853 , y6854 , y6855 , y6856 , y6857 , y6858 , y6859 , y6860 , y6861 , y6862 , y6863 , y6864 , y6865 , y6866 , y6867 , y6868 , y6869 , y6870 , y6871 , y6872 , y6873 , y6874 , y6875 , y6876 , y6877 , y6878 , y6879 , y6880 , y6881 , y6882 , y6883 , y6884 , y6885 , y6886 , y6887 , y6888 , y6889 , y6890 , y6891 , y6892 , y6893 , y6894 , y6895 , y6896 , y6897 , y6898 , y6899 , y6900 , y6901 , y6902 , y6903 , y6904 , y6905 , y6906 , y6907 , y6908 , y6909 , y6910 , y6911 , y6912 , y6913 , y6914 , y6915 , y6916 , y6917 , y6918 , y6919 , y6920 , y6921 , y6922 , y6923 , y6924 , y6925 , y6926 , y6927 , y6928 , y6929 , y6930 , y6931 , y6932 , y6933 , y6934 , y6935 , y6936 , y6937 , y6938 , y6939 , y6940 , y6941 , y6942 , y6943 , y6944 , y6945 , y6946 , y6947 , y6948 , y6949 , y6950 , y6951 , y6952 , y6953 , y6954 , y6955 , y6956 , y6957 , y6958 , y6959 , y6960 , y6961 , y6962 , y6963 , y6964 , y6965 , y6966 , y6967 , y6968 , y6969 , y6970 , y6971 , y6972 , y6973 , y6974 , y6975 , y6976 , y6977 , y6978 , y6979 , y6980 , y6981 , y6982 , y6983 , y6984 , y6985 , y6986 , y6987 , y6988 , y6989 , y6990 , y6991 , y6992 , y6993 , y6994 , y6995 , y6996 , y6997 , y6998 , y6999 , y7000 , y7001 , y7002 , y7003 , y7004 , y7005 , y7006 , y7007 , y7008 , y7009 , y7010 , y7011 , y7012 , y7013 , y7014 , y7015 , y7016 , y7017 , y7018 , y7019 , y7020 , y7021 , y7022 , y7023 , y7024 , y7025 , y7026 , y7027 , y7028 , y7029 , y7030 , y7031 , y7032 , y7033 , y7034 , y7035 , y7036 , y7037 , y7038 , y7039 , y7040 , y7041 , y7042 , y7043 , y7044 , y7045 , y7046 , y7047 , y7048 , y7049 , y7050 , y7051 , y7052 , y7053 , y7054 , y7055 , y7056 , y7057 , y7058 , y7059 , y7060 , y7061 , y7062 , y7063 , y7064 , y7065 , y7066 , y7067 , y7068 , y7069 , y7070 , y7071 , y7072 , y7073 , y7074 , y7075 , y7076 , y7077 , y7078 , y7079 , y7080 , y7081 , y7082 , y7083 , y7084 , y7085 , y7086 , y7087 , y7088 , y7089 , y7090 , y7091 , y7092 , y7093 , y7094 , y7095 , y7096 , y7097 , y7098 , y7099 , y7100 , y7101 , y7102 , y7103 , y7104 , y7105 , y7106 , y7107 , y7108 , y7109 , y7110 , y7111 , y7112 , y7113 , y7114 , y7115 , y7116 , y7117 , y7118 , y7119 , y7120 , y7121 , y7122 , y7123 , y7124 , y7125 , y7126 , y7127 , y7128 , y7129 , y7130 , y7131 , y7132 , y7133 , y7134 , y7135 , y7136 , y7137 , y7138 , y7139 , y7140 , y7141 , y7142 , y7143 , y7144 , y7145 , y7146 , y7147 , y7148 , y7149 , y7150 , y7151 , y7152 , y7153 , y7154 , y7155 , y7156 , y7157 , y7158 , y7159 , y7160 , y7161 , y7162 , y7163 , y7164 , y7165 , y7166 , y7167 , y7168 , y7169 , y7170 , y7171 , y7172 , y7173 , y7174 , y7175 , y7176 , y7177 , y7178 , y7179 , y7180 , y7181 , y7182 , y7183 , y7184 , y7185 , y7186 , y7187 , y7188 , y7189 , y7190 , y7191 , y7192 , y7193 , y7194 , y7195 , y7196 , y7197 , y7198 , y7199 , y7200 , y7201 , y7202 , y7203 , y7204 , y7205 , y7206 , y7207 , y7208 , y7209 , y7210 , y7211 , y7212 , y7213 , y7214 , y7215 , y7216 , y7217 , y7218 , y7219 , y7220 , y7221 , y7222 , y7223 , y7224 , y7225 , y7226 , y7227 , y7228 , y7229 , y7230 , y7231 , y7232 , y7233 , y7234 , y7235 , y7236 , y7237 , y7238 , y7239 , y7240 , y7241 , y7242 , y7243 , y7244 , y7245 , y7246 , y7247 , y7248 , y7249 , y7250 , y7251 , y7252 , y7253 , y7254 , y7255 , y7256 , y7257 , y7258 , y7259 , y7260 , y7261 , y7262 , y7263 , y7264 , y7265 , y7266 , y7267 , y7268 , y7269 , y7270 , y7271 , y7272 , y7273 , y7274 , y7275 , y7276 , y7277 , y7278 , y7279 , y7280 , y7281 , y7282 , y7283 , y7284 , y7285 , y7286 , y7287 , y7288 , y7289 , y7290 , y7291 , y7292 , y7293 , y7294 , y7295 , y7296 , y7297 , y7298 , y7299 , y7300 , y7301 , y7302 , y7303 , y7304 , y7305 , y7306 , y7307 , y7308 , y7309 , y7310 , y7311 , y7312 , y7313 , y7314 , y7315 , y7316 , y7317 , y7318 , y7319 , y7320 , y7321 , y7322 , y7323 , y7324 , y7325 , y7326 , y7327 , y7328 , y7329 , y7330 , y7331 , y7332 , y7333 , y7334 , y7335 , y7336 , y7337 , y7338 , y7339 , y7340 , y7341 , y7342 , y7343 , y7344 , y7345 , y7346 , y7347 , y7348 , y7349 , y7350 , y7351 , y7352 , y7353 , y7354 , y7355 , y7356 , y7357 , y7358 , y7359 , y7360 , y7361 , y7362 , y7363 , y7364 , y7365 , y7366 , y7367 , y7368 , y7369 , y7370 , y7371 , y7372 , y7373 , y7374 , y7375 , y7376 , y7377 , y7378 , y7379 , y7380 , y7381 , y7382 , y7383 , y7384 , y7385 , y7386 , y7387 , y7388 , y7389 , y7390 , y7391 , y7392 , y7393 , y7394 , y7395 , y7396 , y7397 , y7398 , y7399 , y7400 , y7401 , y7402 , y7403 , y7404 , y7405 , y7406 , y7407 , y7408 , y7409 , y7410 , y7411 , y7412 , y7413 , y7414 , y7415 , y7416 , y7417 , y7418 , y7419 , y7420 , y7421 , y7422 , y7423 , y7424 , y7425 , y7426 , y7427 , y7428 , y7429 , y7430 , y7431 , y7432 , y7433 , y7434 , y7435 , y7436 , y7437 , y7438 , y7439 , y7440 , y7441 , y7442 , y7443 , y7444 , y7445 , y7446 , y7447 , y7448 , y7449 , y7450 , y7451 , y7452 , y7453 , y7454 , y7455 , y7456 , y7457 , y7458 , y7459 , y7460 , y7461 , y7462 , y7463 , y7464 , y7465 , y7466 , y7467 , y7468 , y7469 , y7470 , y7471 , y7472 , y7473 , y7474 , y7475 , y7476 , y7477 , y7478 , y7479 , y7480 , y7481 , y7482 , y7483 , y7484 , y7485 , y7486 , y7487 , y7488 , y7489 , y7490 , y7491 , y7492 , y7493 , y7494 , y7495 , y7496 , y7497 , y7498 , y7499 , y7500 , y7501 , y7502 , y7503 , y7504 , y7505 , y7506 , y7507 , y7508 , y7509 , y7510 , y7511 , y7512 , y7513 , y7514 , y7515 , y7516 , y7517 , y7518 , y7519 , y7520 , y7521 , y7522 , y7523 , y7524 , y7525 , y7526 , y7527 , y7528 , y7529 , y7530 , y7531 , y7532 , y7533 , y7534 , y7535 , y7536 , y7537 , y7538 , y7539 , y7540 , y7541 , y7542 , y7543 , y7544 , y7545 , y7546 , y7547 , y7548 , y7549 , y7550 , y7551 , y7552 , y7553 , y7554 , y7555 , y7556 , y7557 , y7558 , y7559 , y7560 , y7561 , y7562 , y7563 , y7564 , y7565 , y7566 , y7567 , y7568 , y7569 , y7570 , y7571 , y7572 , y7573 , y7574 , y7575 , y7576 , y7577 , y7578 , y7579 , y7580 , y7581 , y7582 , y7583 , y7584 , y7585 , y7586 , y7587 , y7588 , y7589 , y7590 , y7591 , y7592 , y7593 , y7594 , y7595 , y7596 , y7597 , y7598 , y7599 , y7600 , y7601 , y7602 , y7603 , y7604 , y7605 , y7606 , y7607 , y7608 , y7609 , y7610 , y7611 , y7612 , y7613 , y7614 , y7615 , y7616 , y7617 , y7618 , y7619 , y7620 , y7621 , y7622 , y7623 , y7624 , y7625 , y7626 , y7627 , y7628 , y7629 , y7630 , y7631 , y7632 , y7633 , y7634 , y7635 , y7636 , y7637 , y7638 , y7639 , y7640 , y7641 , y7642 , y7643 , y7644 , y7645 , y7646 , y7647 , y7648 , y7649 , y7650 , y7651 , y7652 , y7653 , y7654 , y7655 , y7656 , y7657 , y7658 , y7659 , y7660 , y7661 , y7662 , y7663 , y7664 , y7665 , y7666 , y7667 , y7668 , y7669 , y7670 , y7671 , y7672 , y7673 , y7674 , y7675 , y7676 , y7677 , y7678 , y7679 , y7680 , y7681 , y7682 , y7683 , y7684 , y7685 , y7686 , y7687 , y7688 , y7689 , y7690 , y7691 , y7692 , y7693 , y7694 , y7695 , y7696 , y7697 , y7698 , y7699 , y7700 , y7701 , y7702 , y7703 , y7704 , y7705 , y7706 , y7707 , y7708 , y7709 , y7710 , y7711 , y7712 , y7713 , y7714 , y7715 , y7716 , y7717 , y7718 , y7719 , y7720 , y7721 , y7722 , y7723 , y7724 , y7725 , y7726 , y7727 , y7728 , y7729 , y7730 , y7731 , y7732 , y7733 , y7734 , y7735 , y7736 , y7737 , y7738 , y7739 , y7740 , y7741 , y7742 , y7743 , y7744 , y7745 , y7746 , y7747 , y7748 , y7749 , y7750 , y7751 , y7752 , y7753 , y7754 , y7755 , y7756 , y7757 , y7758 , y7759 , y7760 , y7761 , y7762 , y7763 , y7764 , y7765 , y7766 , y7767 , y7768 , y7769 , y7770 , y7771 , y7772 , y7773 , y7774 , y7775 , y7776 , y7777 , y7778 , y7779 , y7780 , y7781 , y7782 , y7783 , y7784 , y7785 , y7786 , y7787 , y7788 , y7789 , y7790 , y7791 , y7792 , y7793 , y7794 , y7795 , y7796 , y7797 , y7798 , y7799 , y7800 , y7801 , y7802 , y7803 , y7804 , y7805 , y7806 , y7807 , y7808 , y7809 , y7810 , y7811 , y7812 , y7813 , y7814 , y7815 , y7816 , y7817 , y7818 , y7819 , y7820 , y7821 , y7822 , y7823 , y7824 , y7825 , y7826 , y7827 , y7828 , y7829 , y7830 , y7831 , y7832 , y7833 , y7834 , y7835 , y7836 , y7837 , y7838 , y7839 , y7840 , y7841 , y7842 , y7843 , y7844 , y7845 , y7846 , y7847 , y7848 , y7849 , y7850 , y7851 , y7852 , y7853 , y7854 , y7855 , y7856 , y7857 , y7858 , y7859 , y7860 , y7861 , y7862 , y7863 , y7864 , y7865 , y7866 , y7867 , y7868 , y7869 , y7870 , y7871 , y7872 , y7873 , y7874 , y7875 , y7876 , y7877 , y7878 , y7879 , y7880 , y7881 , y7882 , y7883 , y7884 , y7885 , y7886 , y7887 , y7888 , y7889 , y7890 , y7891 , y7892 , y7893 , y7894 , y7895 , y7896 , y7897 , y7898 , y7899 , y7900 , y7901 , y7902 , y7903 , y7904 , y7905 , y7906 , y7907 , y7908 , y7909 , y7910 , y7911 , y7912 , y7913 , y7914 , y7915 , y7916 , y7917 , y7918 , y7919 , y7920 , y7921 , y7922 , y7923 , y7924 , y7925 , y7926 , y7927 , y7928 , y7929 , y7930 , y7931 , y7932 , y7933 , y7934 , y7935 , y7936 , y7937 , y7938 , y7939 , y7940 , y7941 , y7942 , y7943 , y7944 , y7945 , y7946 , y7947 , y7948 , y7949 , y7950 , y7951 , y7952 , y7953 , y7954 , y7955 , y7956 , y7957 , y7958 , y7959 , y7960 , y7961 , y7962 , y7963 , y7964 , y7965 , y7966 , y7967 , y7968 , y7969 , y7970 , y7971 , y7972 , y7973 , y7974 , y7975 , y7976 , y7977 , y7978 , y7979 , y7980 , y7981 , y7982 , y7983 , y7984 , y7985 , y7986 , y7987 , y7988 , y7989 , y7990 , y7991 , y7992 , y7993 , y7994 , y7995 , y7996 , y7997 , y7998 , y7999 , y8000 , y8001 , y8002 , y8003 , y8004 , y8005 , y8006 , y8007 , y8008 , y8009 , y8010 , y8011 , y8012 , y8013 , y8014 , y8015 , y8016 , y8017 , y8018 , y8019 , y8020 , y8021 , y8022 , y8023 , y8024 , y8025 , y8026 , y8027 , y8028 , y8029 , y8030 , y8031 , y8032 , y8033 , y8034 , y8035 , y8036 , y8037 , y8038 , y8039 , y8040 , y8041 , y8042 , y8043 , y8044 , y8045 , y8046 , y8047 , y8048 , y8049 , y8050 , y8051 , y8052 , y8053 , y8054 , y8055 , y8056 , y8057 , y8058 , y8059 , y8060 , y8061 , y8062 , y8063 , y8064 , y8065 , y8066 , y8067 , y8068 , y8069 , y8070 , y8071 , y8072 , y8073 , y8074 , y8075 , y8076 , y8077 , y8078 , y8079 , y8080 , y8081 , y8082 , y8083 , y8084 , y8085 , y8086 , y8087 , y8088 , y8089 , y8090 , y8091 , y8092 , y8093 , y8094 , y8095 , y8096 , y8097 , y8098 , y8099 , y8100 , y8101 , y8102 , y8103 , y8104 , y8105 , y8106 , y8107 , y8108 , y8109 , y8110 , y8111 , y8112 , y8113 , y8114 , y8115 , y8116 , y8117 , y8118 , y8119 , y8120 , y8121 , y8122 , y8123 , y8124 , y8125 , y8126 , y8127 , y8128 , y8129 , y8130 , y8131 , y8132 , y8133 , y8134 , y8135 , y8136 , y8137 , y8138 , y8139 , y8140 , y8141 , y8142 , y8143 , y8144 , y8145 , y8146 , y8147 , y8148 , y8149 , y8150 , y8151 , y8152 , y8153 , y8154 , y8155 , y8156 , y8157 , y8158 , y8159 , y8160 , y8161 , y8162 , y8163 , y8164 , y8165 , y8166 , y8167 , y8168 , y8169 , y8170 , y8171 , y8172 , y8173 , y8174 , y8175 , y8176 , y8177 , y8178 , y8179 , y8180 , y8181 , y8182 , y8183 , y8184 , y8185 , y8186 , y8187 , y8188 , y8189 , y8190 , y8191 , y8192 , y8193 , y8194 , y8195 , y8196 , y8197 , y8198 , y8199 , y8200 , y8201 , y8202 , y8203 , y8204 , y8205 , y8206 , y8207 , y8208 , y8209 , y8210 , y8211 , y8212 , y8213 , y8214 , y8215 , y8216 , y8217 , y8218 , y8219 , y8220 , y8221 , y8222 , y8223 , y8224 , y8225 , y8226 , y8227 , y8228 , y8229 , y8230 , y8231 , y8232 , y8233 , y8234 , y8235 , y8236 , y8237 , y8238 , y8239 , y8240 , y8241 , y8242 , y8243 , y8244 , y8245 , y8246 , y8247 , y8248 , y8249 , y8250 , y8251 , y8252 , y8253 , y8254 , y8255 , y8256 , y8257 , y8258 , y8259 , y8260 , y8261 , y8262 , y8263 , y8264 , y8265 , y8266 , y8267 , y8268 , y8269 , y8270 , y8271 , y8272 , y8273 , y8274 , y8275 , y8276 , y8277 , y8278 , y8279 , y8280 , y8281 , y8282 , y8283 , y8284 , y8285 , y8286 , y8287 , y8288 , y8289 , y8290 , y8291 , y8292 , y8293 , y8294 , y8295 , y8296 , y8297 , y8298 , y8299 , y8300 , y8301 , y8302 , y8303 , y8304 , y8305 , y8306 , y8307 , y8308 , y8309 , y8310 , y8311 , y8312 , y8313 , y8314 , y8315 , y8316 , y8317 , y8318 , y8319 , y8320 , y8321 , y8322 , y8323 , y8324 , y8325 , y8326 , y8327 , y8328 , y8329 , y8330 , y8331 , y8332 , y8333 , y8334 , y8335 , y8336 , y8337 , y8338 , y8339 , y8340 , y8341 , y8342 , y8343 , y8344 , y8345 , y8346 , y8347 , y8348 , y8349 , y8350 , y8351 , y8352 , y8353 , y8354 , y8355 , y8356 , y8357 , y8358 , y8359 , y8360 , y8361 , y8362 , y8363 , y8364 , y8365 , y8366 , y8367 , y8368 , y8369 , y8370 , y8371 , y8372 , y8373 , y8374 , y8375 , y8376 , y8377 , y8378 , y8379 , y8380 , y8381 , y8382 , y8383 , y8384 , y8385 , y8386 , y8387 , y8388 , y8389 , y8390 , y8391 , y8392 , y8393 , y8394 , y8395 , y8396 , y8397 , y8398 , y8399 , y8400 , y8401 , y8402 , y8403 , y8404 , y8405 , y8406 , y8407 , y8408 , y8409 , y8410 , y8411 , y8412 , y8413 , y8414 , y8415 , y8416 , y8417 , y8418 , y8419 , y8420 , y8421 , y8422 , y8423 , y8424 , y8425 , y8426 , y8427 , y8428 , y8429 , y8430 , y8431 , y8432 , y8433 , y8434 , y8435 , y8436 , y8437 , y8438 , y8439 , y8440 , y8441 , y8442 , y8443 , y8444 , y8445 , y8446 , y8447 , y8448 , y8449 , y8450 , y8451 , y8452 , y8453 , y8454 , y8455 , y8456 , y8457 , y8458 , y8459 , y8460 , y8461 , y8462 , y8463 , y8464 , y8465 , y8466 , y8467 , y8468 , y8469 , y8470 , y8471 , y8472 , y8473 , y8474 , y8475 , y8476 , y8477 , y8478 , y8479 , y8480 , y8481 , y8482 , y8483 , y8484 , y8485 , y8486 , y8487 , y8488 , y8489 , y8490 , y8491 , y8492 , y8493 , y8494 , y8495 , y8496 , y8497 , y8498 , y8499 , y8500 , y8501 , y8502 , y8503 , y8504 , y8505 , y8506 , y8507 , y8508 , y8509 , y8510 , y8511 , y8512 , y8513 , y8514 , y8515 , y8516 , y8517 , y8518 , y8519 , y8520 , y8521 , y8522 , y8523 , y8524 , y8525 , y8526 , y8527 , y8528 , y8529 , y8530 , y8531 , y8532 , y8533 , y8534 , y8535 , y8536 , y8537 , y8538 , y8539 , y8540 , y8541 , y8542 , y8543 , y8544 , y8545 , y8546 , y8547 , y8548 , y8549 , y8550 , y8551 , y8552 , y8553 , y8554 , y8555 , y8556 , y8557 , y8558 , y8559 , y8560 , y8561 , y8562 , y8563 , y8564 , y8565 , y8566 , y8567 , y8568 , y8569 , y8570 , y8571 , y8572 , y8573 , y8574 , y8575 , y8576 , y8577 , y8578 , y8579 , y8580 , y8581 , y8582 , y8583 , y8584 , y8585 , y8586 , y8587 , y8588 , y8589 , y8590 , y8591 , y8592 , y8593 , y8594 , y8595 , y8596 , y8597 , y8598 , y8599 , y8600 , y8601 , y8602 , y8603 , y8604 , y8605 , y8606 , y8607 , y8608 , y8609 , y8610 , y8611 , y8612 , y8613 , y8614 , y8615 , y8616 , y8617 , y8618 , y8619 , y8620 , y8621 , y8622 , y8623 , y8624 , y8625 , y8626 , y8627 , y8628 , y8629 , y8630 , y8631 , y8632 , y8633 , y8634 , y8635 , y8636 , y8637 , y8638 , y8639 , y8640 , y8641 , y8642 , y8643 , y8644 , y8645 , y8646 , y8647 , y8648 , y8649 , y8650 , y8651 , y8652 , y8653 , y8654 , y8655 , y8656 , y8657 , y8658 , y8659 , y8660 , y8661 , y8662 , y8663 , y8664 , y8665 , y8666 , y8667 , y8668 , y8669 , y8670 , y8671 , y8672 , y8673 , y8674 , y8675 , y8676 , y8677 , y8678 , y8679 , y8680 , y8681 , y8682 , y8683 , y8684 , y8685 , y8686 , y8687 , y8688 , y8689 , y8690 , y8691 , y8692 , y8693 , y8694 , y8695 , y8696 , y8697 , y8698 , y8699 , y8700 , y8701 , y8702 , y8703 , y8704 , y8705 , y8706 , y8707 , y8708 , y8709 , y8710 , y8711 , y8712 , y8713 , y8714 , y8715 , y8716 , y8717 , y8718 , y8719 , y8720 , y8721 , y8722 , y8723 , y8724 , y8725 , y8726 , y8727 , y8728 , y8729 , y8730 , y8731 , y8732 , y8733 , y8734 , y8735 , y8736 , y8737 , y8738 , y8739 , y8740 , y8741 , y8742 , y8743 , y8744 , y8745 , y8746 , y8747 , y8748 , y8749 , y8750 , y8751 , y8752 , y8753 , y8754 , y8755 , y8756 , y8757 , y8758 , y8759 , y8760 , y8761 , y8762 , y8763 , y8764 , y8765 , y8766 , y8767 , y8768 , y8769 , y8770 , y8771 , y8772 , y8773 , y8774 , y8775 , y8776 , y8777 , y8778 , y8779 , y8780 , y8781 , y8782 , y8783 , y8784 , y8785 , y8786 , y8787 , y8788 , y8789 , y8790 , y8791 , y8792 , y8793 , y8794 , y8795 , y8796 , y8797 , y8798 , y8799 , y8800 , y8801 , y8802 , y8803 , y8804 , y8805 , y8806 , y8807 , y8808 , y8809 , y8810 , y8811 , y8812 , y8813 , y8814 , y8815 , y8816 , y8817 , y8818 , y8819 , y8820 , y8821 , y8822 , y8823 , y8824 , y8825 , y8826 , y8827 , y8828 , y8829 , y8830 , y8831 , y8832 , y8833 , y8834 , y8835 , y8836 , y8837 , y8838 , y8839 , y8840 , y8841 , y8842 , y8843 , y8844 , y8845 , y8846 , y8847 , y8848 , y8849 , y8850 , y8851 , y8852 , y8853 , y8854 , y8855 , y8856 , y8857 , y8858 , y8859 , y8860 , y8861 , y8862 , y8863 , y8864 , y8865 , y8866 , y8867 , y8868 , y8869 , y8870 , y8871 , y8872 , y8873 , y8874 , y8875 , y8876 , y8877 , y8878 , y8879 , y8880 , y8881 , y8882 , y8883 , y8884 , y8885 , y8886 , y8887 , y8888 , y8889 , y8890 , y8891 , y8892 , y8893 , y8894 , y8895 , y8896 , y8897 , y8898 , y8899 , y8900 , y8901 , y8902 , y8903 , y8904 , y8905 , y8906 , y8907 , y8908 , y8909 , y8910 , y8911 , y8912 , y8913 , y8914 , y8915 , y8916 , y8917 , y8918 , y8919 , y8920 , y8921 , y8922 , y8923 , y8924 , y8925 , y8926 , y8927 , y8928 , y8929 , y8930 , y8931 , y8932 , y8933 , y8934 , y8935 , y8936 , y8937 , y8938 , y8939 , y8940 , y8941 , y8942 , y8943 , y8944 , y8945 , y8946 , y8947 , y8948 , y8949 , y8950 , y8951 , y8952 , y8953 , y8954 , y8955 , y8956 , y8957 , y8958 , y8959 , y8960 , y8961 , y8962 , y8963 , y8964 , y8965 , y8966 , y8967 , y8968 , y8969 , y8970 , y8971 , y8972 , y8973 , y8974 , y8975 , y8976 , y8977 , y8978 , y8979 , y8980 , y8981 , y8982 , y8983 , y8984 , y8985 , y8986 , y8987 , y8988 , y8989 , y8990 , y8991 , y8992 , y8993 , y8994 , y8995 , y8996 , y8997 , y8998 , y8999 , y9000 , y9001 , y9002 , y9003 , y9004 , y9005 , y9006 , y9007 , y9008 , y9009 , y9010 , y9011 , y9012 , y9013 , y9014 , y9015 , y9016 , y9017 , y9018 , y9019 , y9020 , y9021 , y9022 , y9023 , y9024 , y9025 , y9026 , y9027 , y9028 , y9029 , y9030 , y9031 , y9032 , y9033 , y9034 , y9035 , y9036 , y9037 , y9038 , y9039 , y9040 , y9041 , y9042 , y9043 , y9044 , y9045 , y9046 , y9047 , y9048 , y9049 , y9050 , y9051 , y9052 , y9053 , y9054 , y9055 , y9056 , y9057 , y9058 , y9059 , y9060 , y9061 , y9062 , y9063 , y9064 , y9065 , y9066 , y9067 , y9068 , y9069 , y9070 , y9071 , y9072 , y9073 , y9074 , y9075 , y9076 , y9077 , y9078 , y9079 , y9080 , y9081 , y9082 , y9083 , y9084 , y9085 , y9086 , y9087 , y9088 , y9089 , y9090 , y9091 , y9092 , y9093 , y9094 , y9095 , y9096 , y9097 , y9098 , y9099 , y9100 , y9101 , y9102 , y9103 , y9104 , y9105 , y9106 , y9107 , y9108 , y9109 , y9110 , y9111 , y9112 , y9113 , y9114 , y9115 , y9116 , y9117 , y9118 , y9119 , y9120 , y9121 , y9122 , y9123 , y9124 , y9125 , y9126 , y9127 , y9128 , y9129 , y9130 , y9131 , y9132 , y9133 , y9134 , y9135 , y9136 , y9137 , y9138 , y9139 , y9140 , y9141 , y9142 , y9143 , y9144 , y9145 , y9146 , y9147 , y9148 , y9149 , y9150 , y9151 , y9152 , y9153 , y9154 , y9155 , y9156 , y9157 , y9158 , y9159 , y9160 , y9161 , y9162 , y9163 , y9164 , y9165 , y9166 , y9167 , y9168 , y9169 , y9170 , y9171 , y9172 , y9173 , y9174 , y9175 , y9176 , y9177 , y9178 , y9179 , y9180 , y9181 , y9182 , y9183 , y9184 , y9185 , y9186 , y9187 , y9188 , y9189 , y9190 , y9191 , y9192 , y9193 , y9194 , y9195 , y9196 , y9197 , y9198 , y9199 , y9200 , y9201 , y9202 , y9203 , y9204 , y9205 , y9206 , y9207 , y9208 , y9209 , y9210 , y9211 , y9212 , y9213 , y9214 , y9215 , y9216 , y9217 , y9218 , y9219 , y9220 , y9221 , y9222 , y9223 , y9224 , y9225 , y9226 , y9227 , y9228 , y9229 , y9230 , y9231 , y9232 , y9233 , y9234 , y9235 , y9236 , y9237 , y9238 , y9239 , y9240 , y9241 , y9242 , y9243 , y9244 , y9245 , y9246 , y9247 , y9248 , y9249 , y9250 , y9251 , y9252 , y9253 , y9254 , y9255 , y9256 , y9257 , y9258 , y9259 , y9260 , y9261 , y9262 , y9263 , y9264 , y9265 , y9266 , y9267 , y9268 , y9269 , y9270 , y9271 , y9272 , y9273 , y9274 , y9275 , y9276 , y9277 , y9278 , y9279 , y9280 , y9281 , y9282 , y9283 , y9284 , y9285 , y9286 , y9287 , y9288 , y9289 , y9290 , y9291 , y9292 , y9293 , y9294 , y9295 , y9296 , y9297 , y9298 , y9299 , y9300 , y9301 , y9302 , y9303 , y9304 , y9305 , y9306 , y9307 , y9308 , y9309 , y9310 , y9311 , y9312 , y9313 , y9314 , y9315 , y9316 , y9317 , y9318 , y9319 , y9320 , y9321 , y9322 , y9323 , y9324 , y9325 , y9326 , y9327 , y9328 , y9329 , y9330 , y9331 , y9332 , y9333 , y9334 , y9335 , y9336 , y9337 , y9338 , y9339 , y9340 , y9341 , y9342 , y9343 , y9344 , y9345 , y9346 , y9347 , y9348 , y9349 , y9350 , y9351 , y9352 , y9353 , y9354 , y9355 , y9356 , y9357 , y9358 , y9359 , y9360 , y9361 , y9362 , y9363 , y9364 , y9365 , y9366 , y9367 , y9368 , y9369 , y9370 , y9371 , y9372 , y9373 , y9374 , y9375 , y9376 , y9377 , y9378 , y9379 , y9380 , y9381 , y9382 , y9383 , y9384 , y9385 , y9386 , y9387 , y9388 , y9389 , y9390 , y9391 , y9392 , y9393 , y9394 , y9395 , y9396 , y9397 , y9398 , y9399 , y9400 , y9401 , y9402 , y9403 , y9404 , y9405 , y9406 , y9407 , y9408 , y9409 , y9410 , y9411 , y9412 , y9413 , y9414 , y9415 , y9416 , y9417 , y9418 , y9419 , y9420 , y9421 , y9422 , y9423 , y9424 , y9425 , y9426 , y9427 , y9428 , y9429 , y9430 , y9431 , y9432 , y9433 , y9434 , y9435 , y9436 , y9437 , y9438 , y9439 , y9440 , y9441 , y9442 , y9443 , y9444 , y9445 , y9446 , y9447 , y9448 , y9449 , y9450 , y9451 , y9452 , y9453 , y9454 , y9455 , y9456 , y9457 , y9458 , y9459 , y9460 , y9461 , y9462 , y9463 , y9464 , y9465 , y9466 , y9467 , y9468 , y9469 , y9470 , y9471 , y9472 , y9473 , y9474 , y9475 , y9476 , y9477 , y9478 , y9479 , y9480 , y9481 , y9482 , y9483 , y9484 , y9485 , y9486 , y9487 , y9488 , y9489 , y9490 , y9491 , y9492 , y9493 , y9494 , y9495 , y9496 , y9497 , y9498 , y9499 , y9500 , y9501 , y9502 , y9503 , y9504 , y9505 , y9506 , y9507 , y9508 , y9509 , y9510 , y9511 , y9512 , y9513 , y9514 , y9515 , y9516 , y9517 , y9518 , y9519 , y9520 , y9521 , y9522 , y9523 , y9524 , y9525 , y9526 , y9527 , y9528 , y9529 , y9530 , y9531 , y9532 , y9533 , y9534 , y9535 , y9536 , y9537 , y9538 , y9539 , y9540 , y9541 , y9542 , y9543 , y9544 , y9545 , y9546 , y9547 , y9548 , y9549 , y9550 , y9551 , y9552 , y9553 , y9554 , y9555 , y9556 , y9557 , y9558 , y9559 , y9560 , y9561 , y9562 , y9563 , y9564 , y9565 , y9566 , y9567 , y9568 , y9569 , y9570 , y9571 , y9572 , y9573 , y9574 , y9575 , y9576 , y9577 , y9578 , y9579 , y9580 , y9581 , y9582 , y9583 , y9584 , y9585 , y9586 , y9587 , y9588 , y9589 , y9590 , y9591 , y9592 , y9593 , y9594 , y9595 , y9596 , y9597 , y9598 , y9599 , y9600 , y9601 , y9602 , y9603 , y9604 , y9605 , y9606 , y9607 , y9608 , y9609 , y9610 , y9611 , y9612 , y9613 , y9614 , y9615 , y9616 , y9617 , y9618 , y9619 , y9620 , y9621 , y9622 , y9623 , y9624 , y9625 , y9626 , y9627 , y9628 , y9629 , y9630 , y9631 , y9632 , y9633 , y9634 , y9635 , y9636 , y9637 , y9638 , y9639 , y9640 , y9641 , y9642 , y9643 , y9644 , y9645 , y9646 , y9647 , y9648 , y9649 , y9650 , y9651 , y9652 , y9653 , y9654 , y9655 , y9656 , y9657 , y9658 , y9659 , y9660 , y9661 , y9662 , y9663 , y9664 , y9665 , y9666 , y9667 , y9668 , y9669 , y9670 , y9671 , y9672 , y9673 , y9674 , y9675 , y9676 , y9677 , y9678 , y9679 , y9680 , y9681 , y9682 , y9683 , y9684 , y9685 , y9686 , y9687 , y9688 , y9689 , y9690 , y9691 , y9692 , y9693 , y9694 , y9695 , y9696 , y9697 , y9698 , y9699 , y9700 , y9701 , y9702 , y9703 , y9704 , y9705 , y9706 , y9707 , y9708 , y9709 , y9710 , y9711 , y9712 , y9713 , y9714 , y9715 , y9716 , y9717 , y9718 , y9719 , y9720 , y9721 , y9722 , y9723 , y9724 , y9725 , y9726 , y9727 , y9728 , y9729 , y9730 , y9731 , y9732 , y9733 , y9734 , y9735 , y9736 , y9737 , y9738 , y9739 , y9740 , y9741 , y9742 , y9743 , y9744 , y9745 , y9746 , y9747 , y9748 , y9749 , y9750 , y9751 , y9752 , y9753 , y9754 , y9755 , y9756 , y9757 , y9758 , y9759 , y9760 , y9761 , y9762 , y9763 , y9764 , y9765 , y9766 , y9767 , y9768 , y9769 , y9770 , y9771 , y9772 , y9773 , y9774 , y9775 , y9776 , y9777 , y9778 , y9779 , y9780 , y9781 , y9782 , y9783 , y9784 , y9785 , y9786 , y9787 , y9788 , y9789 , y9790 , y9791 , y9792 , y9793 , y9794 , y9795 , y9796 , y9797 , y9798 , y9799 , y9800 , y9801 , y9802 , y9803 , y9804 , y9805 , y9806 , y9807 , y9808 , y9809 , y9810 , y9811 , y9812 , y9813 , y9814 , y9815 , y9816 , y9817 , y9818 , y9819 , y9820 , y9821 , y9822 , y9823 , y9824 , y9825 , y9826 , y9827 , y9828 , y9829 , y9830 , y9831 , y9832 , y9833 , y9834 , y9835 , y9836 , y9837 , y9838 , y9839 , y9840 , y9841 , y9842 , y9843 , y9844 , y9845 , y9846 , y9847 , y9848 , y9849 , y9850 , y9851 , y9852 , y9853 , y9854 , y9855 , y9856 , y9857 , y9858 , y9859 , y9860 , y9861 , y9862 , y9863 , y9864 , y9865 , y9866 , y9867 , y9868 , y9869 , y9870 , y9871 , y9872 , y9873 , y9874 , y9875 , y9876 , y9877 , y9878 , y9879 , y9880 , y9881 , y9882 , y9883 , y9884 , y9885 , y9886 , y9887 , y9888 , y9889 , y9890 , y9891 , y9892 , y9893 , y9894 , y9895 , y9896 , y9897 , y9898 , y9899 , y9900 , y9901 , y9902 , y9903 , y9904 , y9905 , y9906 , y9907 , y9908 , y9909 , y9910 , y9911 , y9912 , y9913 , y9914 , y9915 , y9916 , y9917 , y9918 , y9919 , y9920 , y9921 , y9922 , y9923 , y9924 , y9925 , y9926 , y9927 , y9928 , y9929 , y9930 , y9931 , y9932 , y9933 , y9934 , y9935 , y9936 , y9937 , y9938 , y9939 , y9940 , y9941 , y9942 , y9943 , y9944 , y9945 , y9946 , y9947 , y9948 , y9949 , y9950 , y9951 , y9952 , y9953 , y9954 , y9955 , y9956 , y9957 , y9958 , y9959 , y9960 , y9961 , y9962 , y9963 , y9964 , y9965 , y9966 , y9967 , y9968 , y9969 , y9970 , y9971 , y9972 , y9973 , y9974 , y9975 , y9976 , y9977 , y9978 , y9979 , y9980 , y9981 , y9982 , y9983 , y9984 , y9985 , y9986 , y9987 , y9988 , y9989 , y9990 , y9991 , y9992 , y9993 , y9994 , y9995 , y9996 , y9997 , y9998 , y9999 , y10000 , y10001 , y10002 , y10003 , y10004 , y10005 , y10006 , y10007 , y10008 , y10009 , y10010 , y10011 , y10012 , y10013 , y10014 , y10015 , y10016 , y10017 , y10018 , y10019 , y10020 , y10021 , y10022 , y10023 , y10024 , y10025 , y10026 , y10027 , y10028 , y10029 , y10030 , y10031 , y10032 , y10033 , y10034 , y10035 , y10036 , y10037 , y10038 , y10039 , y10040 , y10041 , y10042 , y10043 , y10044 , y10045 , y10046 , y10047 , y10048 , y10049 , y10050 , y10051 , y10052 , y10053 , y10054 , y10055 , y10056 , y10057 , y10058 , y10059 , y10060 , y10061 , y10062 , y10063 , y10064 , y10065 , y10066 , y10067 , y10068 , y10069 , y10070 , y10071 , y10072 , y10073 , y10074 , y10075 , y10076 , y10077 , y10078 , y10079 , y10080 , y10081 , y10082 , y10083 , y10084 , y10085 , y10086 , y10087 , y10088 , y10089 , y10090 , y10091 , y10092 , y10093 , y10094 , y10095 , y10096 , y10097 , y10098 , y10099 , y10100 , y10101 , y10102 , y10103 , y10104 , y10105 , y10106 , y10107 , y10108 , y10109 , y10110 , y10111 , y10112 , y10113 , y10114 , y10115 , y10116 , y10117 , y10118 , y10119 , y10120 , y10121 , y10122 , y10123 , y10124 , y10125 , y10126 , y10127 , y10128 , y10129 , y10130 , y10131 , y10132 , y10133 , y10134 , y10135 , y10136 , y10137 , y10138 , y10139 , y10140 , y10141 , y10142 , y10143 , y10144 , y10145 , y10146 , y10147 , y10148 , y10149 , y10150 , y10151 , y10152 , y10153 , y10154 , y10155 , y10156 , y10157 , y10158 , y10159 , y10160 , y10161 , y10162 , y10163 , y10164 , y10165 , y10166 , y10167 , y10168 , y10169 , y10170 , y10171 , y10172 , y10173 , y10174 , y10175 , y10176 , y10177 , y10178 , y10179 , y10180 , y10181 , y10182 , y10183 , y10184 , y10185 , y10186 , y10187 , y10188 , y10189 , y10190 , y10191 , y10192 , y10193 , y10194 , y10195 , y10196 , y10197 , y10198 , y10199 , y10200 , y10201 , y10202 , y10203 , y10204 , y10205 , y10206 , y10207 , y10208 , y10209 , y10210 , y10211 , y10212 , y10213 , y10214 , y10215 , y10216 , y10217 , y10218 , y10219 , y10220 , y10221 , y10222 , y10223 , y10224 , y10225 , y10226 , y10227 , y10228 , y10229 , y10230 , y10231 , y10232 , y10233 , y10234 , y10235 , y10236 , y10237 , y10238 , y10239 , y10240 , y10241 , y10242 , y10243 , y10244 , y10245 , y10246 , y10247 , y10248 , y10249 , y10250 , y10251 , y10252 , y10253 , y10254 , y10255 , y10256 , y10257 , y10258 , y10259 , y10260 , y10261 , y10262 , y10263 , y10264 , y10265 , y10266 , y10267 , y10268 , y10269 , y10270 , y10271 , y10272 , y10273 , y10274 , y10275 , y10276 , y10277 , y10278 , y10279 , y10280 , y10281 , y10282 , y10283 , y10284 , y10285 , y10286 , y10287 , y10288 , y10289 , y10290 , y10291 , y10292 , y10293 , y10294 , y10295 , y10296 , y10297 , y10298 , y10299 , y10300 , y10301 , y10302 , y10303 , y10304 , y10305 , y10306 , y10307 , y10308 , y10309 , y10310 , y10311 , y10312 , y10313 , y10314 , y10315 , y10316 , y10317 , y10318 , y10319 , y10320 , y10321 , y10322 , y10323 , y10324 , y10325 , y10326 , y10327 , y10328 , y10329 , y10330 , y10331 , y10332 , y10333 , y10334 , y10335 , y10336 , y10337 , y10338 , y10339 , y10340 , y10341 , y10342 , y10343 , y10344 , y10345 , y10346 , y10347 , y10348 , y10349 , y10350 , y10351 , y10352 , y10353 , y10354 , y10355 , y10356 , y10357 , y10358 , y10359 , y10360 , y10361 , y10362 , y10363 , y10364 , y10365 , y10366 , y10367 , y10368 , y10369 , y10370 , y10371 , y10372 , y10373 , y10374 , y10375 , y10376 , y10377 , y10378 , y10379 , y10380 , y10381 , y10382 , y10383 , y10384 , y10385 , y10386 , y10387 , y10388 , y10389 , y10390 , y10391 , y10392 , y10393 , y10394 , y10395 , y10396 , y10397 , y10398 , y10399 , y10400 , y10401 , y10402 , y10403 , y10404 , y10405 , y10406 , y10407 , y10408 , y10409 , y10410 , y10411 , y10412 , y10413 , y10414 , y10415 , y10416 , y10417 , y10418 , y10419 , y10420 , y10421 , y10422 , y10423 , y10424 , y10425 , y10426 , y10427 , y10428 , y10429 , y10430 , y10431 , y10432 , y10433 , y10434 , y10435 , y10436 , y10437 , y10438 , y10439 , y10440 , y10441 , y10442 , y10443 , y10444 , y10445 , y10446 , y10447 , y10448 , y10449 , y10450 , y10451 , y10452 , y10453 , y10454 , y10455 , y10456 , y10457 , y10458 , y10459 , y10460 , y10461 , y10462 , y10463 , y10464 , y10465 , y10466 , y10467 , y10468 , y10469 , y10470 , y10471 , y10472 , y10473 , y10474 , y10475 , y10476 , y10477 , y10478 , y10479 , y10480 , y10481 , y10482 , y10483 , y10484 , y10485 , y10486 , y10487 , y10488 , y10489 , y10490 , y10491 , y10492 , y10493 , y10494 , y10495 , y10496 , y10497 , y10498 , y10499 , y10500 , y10501 , y10502 , y10503 , y10504 , y10505 , y10506 , y10507 , y10508 , y10509 , y10510 , y10511 , y10512 , y10513 , y10514 , y10515 , y10516 , y10517 , y10518 , y10519 , y10520 , y10521 , y10522 , y10523 , y10524 , y10525 , y10526 , y10527 , y10528 , y10529 , y10530 , y10531 , y10532 , y10533 , y10534 , y10535 , y10536 , y10537 , y10538 , y10539 , y10540 , y10541 , y10542 , y10543 , y10544 , y10545 , y10546 , y10547 , y10548 , y10549 , y10550 , y10551 , y10552 , y10553 , y10554 , y10555 , y10556 , y10557 , y10558 , y10559 , y10560 , y10561 , y10562 , y10563 , y10564 , y10565 , y10566 , y10567 , y10568 , y10569 , y10570 , y10571 , y10572 , y10573 , y10574 , y10575 , y10576 , y10577 , y10578 , y10579 , y10580 , y10581 , y10582 , y10583 , y10584 , y10585 , y10586 , y10587 , y10588 , y10589 , y10590 , y10591 , y10592 , y10593 , y10594 , y10595 , y10596 , y10597 , y10598 , y10599 , y10600 , y10601 , y10602 , y10603 , y10604 , y10605 , y10606 , y10607 , y10608 , y10609 , y10610 , y10611 , y10612 , y10613 , y10614 , y10615 , y10616 , y10617 , y10618 , y10619 , y10620 , y10621 , y10622 , y10623 , y10624 , y10625 , y10626 , y10627 , y10628 , y10629 , y10630 , y10631 , y10632 , y10633 , y10634 , y10635 , y10636 , y10637 , y10638 , y10639 , y10640 , y10641 , y10642 , y10643 , y10644 , y10645 , y10646 , y10647 , y10648 , y10649 , y10650 , y10651 , y10652 , y10653 , y10654 , y10655 , y10656 , y10657 , y10658 , y10659 , y10660 , y10661 , y10662 , y10663 , y10664 , y10665 , y10666 , y10667 , y10668 , y10669 , y10670 , y10671 , y10672 , y10673 , y10674 , y10675 , y10676 , y10677 , y10678 , y10679 , y10680 , y10681 , y10682 , y10683 , y10684 , y10685 , y10686 , y10687 , y10688 , y10689 , y10690 , y10691 , y10692 , y10693 , y10694 , y10695 , y10696 , y10697 , y10698 , y10699 , y10700 , y10701 , y10702 , y10703 , y10704 , y10705 , y10706 , y10707 , y10708 , y10709 , y10710 , y10711 , y10712 , y10713 , y10714 , y10715 , y10716 , y10717 , y10718 , y10719 , y10720 , y10721 , y10722 , y10723 , y10724 , y10725 , y10726 , y10727 , y10728 , y10729 , y10730 , y10731 , y10732 , y10733 , y10734 , y10735 , y10736 , y10737 , y10738 , y10739 , y10740 , y10741 , y10742 , y10743 , y10744 , y10745 , y10746 , y10747 , y10748 , y10749 , y10750 , y10751 , y10752 , y10753 , y10754 , y10755 , y10756 , y10757 , y10758 , y10759 , y10760 , y10761 , y10762 , y10763 , y10764 , y10765 , y10766 , y10767 , y10768 , y10769 , y10770 , y10771 , y10772 , y10773 , y10774 , y10775 , y10776 , y10777 , y10778 , y10779 , y10780 , y10781 , y10782 , y10783 , y10784 , y10785 , y10786 , y10787 , y10788 , y10789 , y10790 , y10791 , y10792 , y10793 , y10794 , y10795 , y10796 , y10797 , y10798 , y10799 , y10800 , y10801 , y10802 , y10803 , y10804 , y10805 , y10806 , y10807 , y10808 , y10809 , y10810 , y10811 , y10812 , y10813 , y10814 , y10815 , y10816 , y10817 , y10818 , y10819 , y10820 , y10821 , y10822 , y10823 , y10824 , y10825 , y10826 , y10827 , y10828 , y10829 , y10830 , y10831 , y10832 , y10833 , y10834 , y10835 , y10836 , y10837 , y10838 , y10839 , y10840 , y10841 , y10842 , y10843 , y10844 , y10845 , y10846 , y10847 , y10848 , y10849 , y10850 , y10851 , y10852 , y10853 , y10854 , y10855 , y10856 , y10857 , y10858 , y10859 , y10860 , y10861 , y10862 , y10863 , y10864 , y10865 , y10866 , y10867 , y10868 , y10869 , y10870 , y10871 , y10872 , y10873 , y10874 , y10875 , y10876 , y10877 , y10878 , y10879 , y10880 , y10881 , y10882 , y10883 , y10884 , y10885 , y10886 , y10887 , y10888 , y10889 , y10890 , y10891 , y10892 , y10893 , y10894 , y10895 , y10896 , y10897 , y10898 , y10899 , y10900 , y10901 , y10902 , y10903 , y10904 , y10905 , y10906 , y10907 , y10908 , y10909 , y10910 , y10911 , y10912 , y10913 , y10914 , y10915 , y10916 , y10917 , y10918 , y10919 , y10920 , y10921 , y10922 , y10923 , y10924 , y10925 , y10926 , y10927 , y10928 , y10929 , y10930 , y10931 , y10932 , y10933 , y10934 , y10935 , y10936 , y10937 , y10938 , y10939 , y10940 , y10941 , y10942 , y10943 , y10944 , y10945 , y10946 , y10947 , y10948 , y10949 , y10950 , y10951 , y10952 , y10953 , y10954 , y10955 , y10956 , y10957 , y10958 , y10959 , y10960 , y10961 , y10962 , y10963 , y10964 , y10965 , y10966 , y10967 , y10968 , y10969 , y10970 , y10971 , y10972 , y10973 , y10974 , y10975 , y10976 , y10977 , y10978 , y10979 , y10980 , y10981 , y10982 , y10983 , y10984 , y10985 , y10986 , y10987 , y10988 , y10989 , y10990 , y10991 , y10992 , y10993 , y10994 , y10995 , y10996 , y10997 , y10998 , y10999 , y11000 , y11001 , y11002 , y11003 , y11004 , y11005 , y11006 , y11007 , y11008 , y11009 , y11010 , y11011 , y11012 , y11013 , y11014 , y11015 , y11016 , y11017 , y11018 , y11019 , y11020 , y11021 , y11022 , y11023 , y11024 , y11025 , y11026 , y11027 , y11028 , y11029 , y11030 , y11031 , y11032 , y11033 , y11034 , y11035 , y11036 , y11037 , y11038 , y11039 , y11040 , y11041 , y11042 , y11043 , y11044 , y11045 , y11046 , y11047 , y11048 , y11049 , y11050 , y11051 , y11052 , y11053 , y11054 , y11055 , y11056 , y11057 , y11058 , y11059 , y11060 , y11061 , y11062 , y11063 , y11064 , y11065 , y11066 , y11067 , y11068 , y11069 , y11070 , y11071 , y11072 , y11073 , y11074 , y11075 , y11076 , y11077 , y11078 , y11079 , y11080 , y11081 , y11082 , y11083 , y11084 , y11085 , y11086 , y11087 , y11088 , y11089 , y11090 , y11091 , y11092 , y11093 , y11094 , y11095 , y11096 , y11097 , y11098 , y11099 , y11100 , y11101 , y11102 , y11103 , y11104 , y11105 , y11106 , y11107 , y11108 , y11109 , y11110 , y11111 , y11112 , y11113 , y11114 , y11115 , y11116 , y11117 , y11118 , y11119 , y11120 , y11121 , y11122 , y11123 , y11124 , y11125 , y11126 , y11127 , y11128 , y11129 , y11130 , y11131 , y11132 , y11133 , y11134 , y11135 , y11136 , y11137 , y11138 , y11139 , y11140 , y11141 , y11142 , y11143 , y11144 , y11145 , y11146 , y11147 , y11148 , y11149 , y11150 , y11151 , y11152 , y11153 , y11154 , y11155 , y11156 , y11157 , y11158 , y11159 , y11160 , y11161 , y11162 , y11163 , y11164 , y11165 , y11166 , y11167 , y11168 , y11169 , y11170 , y11171 , y11172 , y11173 , y11174 , y11175 , y11176 , y11177 , y11178 , y11179 , y11180 , y11181 , y11182 , y11183 , y11184 , y11185 , y11186 , y11187 , y11188 , y11189 , y11190 , y11191 , y11192 , y11193 , y11194 , y11195 , y11196 , y11197 , y11198 , y11199 , y11200 , y11201 , y11202 , y11203 , y11204 , y11205 , y11206 , y11207 , y11208 , y11209 , y11210 , y11211 , y11212 , y11213 , y11214 , y11215 , y11216 , y11217 , y11218 , y11219 , y11220 , y11221 , y11222 , y11223 , y11224 , y11225 , y11226 , y11227 , y11228 , y11229 , y11230 , y11231 , y11232 , y11233 , y11234 , y11235 , y11236 , y11237 , y11238 , y11239 , y11240 , y11241 , y11242 , y11243 , y11244 , y11245 , y11246 , y11247 , y11248 , y11249 , y11250 , y11251 , y11252 , y11253 , y11254 , y11255 , y11256 , y11257 , y11258 , y11259 , y11260 , y11261 , y11262 , y11263 , y11264 , y11265 , y11266 , y11267 , y11268 , y11269 , y11270 , y11271 , y11272 , y11273 , y11274 , y11275 , y11276 , y11277 , y11278 , y11279 , y11280 , y11281 , y11282 , y11283 , y11284 , y11285 , y11286 , y11287 , y11288 , y11289 , y11290 , y11291 , y11292 , y11293 , y11294 , y11295 , y11296 , y11297 , y11298 , y11299 , y11300 , y11301 , y11302 , y11303 , y11304 , y11305 , y11306 , y11307 , y11308 , y11309 , y11310 , y11311 , y11312 , y11313 , y11314 , y11315 , y11316 , y11317 , y11318 , y11319 , y11320 , y11321 , y11322 , y11323 , y11324 , y11325 , y11326 , y11327 , y11328 , y11329 , y11330 , y11331 , y11332 , y11333 , y11334 , y11335 , y11336 , y11337 , y11338 , y11339 , y11340 , y11341 , y11342 , y11343 , y11344 , y11345 , y11346 , y11347 , y11348 , y11349 , y11350 , y11351 , y11352 , y11353 , y11354 , y11355 , y11356 , y11357 , y11358 , y11359 , y11360 , y11361 , y11362 , y11363 , y11364 , y11365 , y11366 , y11367 , y11368 , y11369 , y11370 , y11371 , y11372 , y11373 , y11374 , y11375 , y11376 , y11377 , y11378 , y11379 , y11380 , y11381 , y11382 , y11383 , y11384 , y11385 , y11386 , y11387 , y11388 , y11389 , y11390 , y11391 , y11392 , y11393 , y11394 , y11395 , y11396 , y11397 , y11398 , y11399 , y11400 , y11401 , y11402 , y11403 , y11404 , y11405 , y11406 , y11407 , y11408 , y11409 , y11410 , y11411 , y11412 , y11413 , y11414 , y11415 , y11416 , y11417 , y11418 , y11419 , y11420 , y11421 , y11422 , y11423 , y11424 , y11425 , y11426 , y11427 , y11428 , y11429 , y11430 , y11431 , y11432 , y11433 , y11434 , y11435 , y11436 , y11437 , y11438 , y11439 , y11440 , y11441 , y11442 , y11443 , y11444 , y11445 , y11446 , y11447 , y11448 , y11449 , y11450 , y11451 , y11452 , y11453 , y11454 , y11455 , y11456 , y11457 , y11458 , y11459 , y11460 , y11461 , y11462 , y11463 , y11464 , y11465 , y11466 , y11467 , y11468 , y11469 , y11470 , y11471 , y11472 , y11473 , y11474 , y11475 , y11476 , y11477 , y11478 , y11479 , y11480 , y11481 , y11482 , y11483 , y11484 , y11485 , y11486 , y11487 , y11488 , y11489 , y11490 , y11491 , y11492 , y11493 , y11494 , y11495 , y11496 , y11497 , y11498 , y11499 , y11500 , y11501 , y11502 , y11503 , y11504 , y11505 , y11506 , y11507 , y11508 , y11509 , y11510 , y11511 , y11512 , y11513 , y11514 , y11515 , y11516 , y11517 , y11518 , y11519 , y11520 , y11521 , y11522 , y11523 , y11524 , y11525 , y11526 , y11527 , y11528 , y11529 , y11530 , y11531 , y11532 , y11533 , y11534 , y11535 , y11536 , y11537 , y11538 , y11539 , y11540 , y11541 , y11542 , y11543 , y11544 , y11545 , y11546 , y11547 , y11548 , y11549 , y11550 , y11551 , y11552 , y11553 , y11554 , y11555 , y11556 , y11557 , y11558 , y11559 , y11560 , y11561 , y11562 , y11563 , y11564 , y11565 , y11566 , y11567 , y11568 , y11569 , y11570 , y11571 , y11572 , y11573 , y11574 , y11575 , y11576 , y11577 , y11578 , y11579 , y11580 , y11581 , y11582 , y11583 , y11584 , y11585 , y11586 , y11587 , y11588 , y11589 , y11590 , y11591 , y11592 , y11593 , y11594 , y11595 , y11596 , y11597 , y11598 , y11599 , y11600 , y11601 , y11602 , y11603 , y11604 , y11605 , y11606 , y11607 , y11608 , y11609 , y11610 , y11611 , y11612 , y11613 , y11614 , y11615 , y11616 , y11617 , y11618 , y11619 , y11620 , y11621 , y11622 , y11623 , y11624 , y11625 , y11626 , y11627 , y11628 , y11629 , y11630 , y11631 , y11632 , y11633 , y11634 , y11635 , y11636 , y11637 , y11638 , y11639 , y11640 , y11641 , y11642 , y11643 , y11644 , y11645 , y11646 , y11647 , y11648 , y11649 , y11650 , y11651 , y11652 , y11653 , y11654 , y11655 , y11656 , y11657 , y11658 , y11659 , y11660 , y11661 , y11662 , y11663 , y11664 , y11665 , y11666 , y11667 , y11668 , y11669 , y11670 , y11671 , y11672 , y11673 , y11674 , y11675 , y11676 , y11677 , y11678 , y11679 , y11680 , y11681 , y11682 , y11683 , y11684 , y11685 , y11686 , y11687 , y11688 , y11689 , y11690 , y11691 , y11692 , y11693 , y11694 , y11695 , y11696 , y11697 , y11698 , y11699 , y11700 , y11701 , y11702 , y11703 , y11704 , y11705 , y11706 , y11707 , y11708 , y11709 , y11710 , y11711 , y11712 , y11713 , y11714 , y11715 , y11716 , y11717 , y11718 , y11719 , y11720 , y11721 , y11722 , y11723 , y11724 , y11725 , y11726 , y11727 , y11728 , y11729 , y11730 , y11731 , y11732 , y11733 , y11734 , y11735 , y11736 , y11737 , y11738 , y11739 , y11740 , y11741 , y11742 , y11743 , y11744 , y11745 , y11746 , y11747 , y11748 , y11749 , y11750 , y11751 , y11752 , y11753 , y11754 , y11755 , y11756 , y11757 , y11758 , y11759 , y11760 , y11761 , y11762 , y11763 , y11764 , y11765 , y11766 , y11767 , y11768 , y11769 , y11770 , y11771 , y11772 , y11773 , y11774 , y11775 , y11776 , y11777 , y11778 , y11779 , y11780 , y11781 , y11782 , y11783 , y11784 , y11785 , y11786 , y11787 , y11788 , y11789 , y11790 , y11791 , y11792 , y11793 , y11794 , y11795 , y11796 , y11797 , y11798 , y11799 , y11800 , y11801 , y11802 , y11803 , y11804 , y11805 , y11806 , y11807 , y11808 , y11809 , y11810 , y11811 , y11812 , y11813 , y11814 , y11815 , y11816 , y11817 , y11818 , y11819 , y11820 , y11821 , y11822 , y11823 , y11824 , y11825 , y11826 , y11827 , y11828 , y11829 , y11830 , y11831 , y11832 , y11833 , y11834 , y11835 , y11836 , y11837 , y11838 , y11839 , y11840 , y11841 , y11842 , y11843 , y11844 , y11845 , y11846 , y11847 , y11848 , y11849 , y11850 , y11851 , y11852 , y11853 , y11854 , y11855 , y11856 , y11857 , y11858 , y11859 , y11860 , y11861 , y11862 , y11863 , y11864 , y11865 , y11866 , y11867 , y11868 , y11869 , y11870 , y11871 , y11872 , y11873 , y11874 , y11875 , y11876 , y11877 , y11878 , y11879 , y11880 , y11881 , y11882 , y11883 , y11884 , y11885 , y11886 , y11887 , y11888 , y11889 , y11890 , y11891 , y11892 , y11893 , y11894 , y11895 , y11896 , y11897 , y11898 , y11899 , y11900 , y11901 , y11902 , y11903 , y11904 , y11905 , y11906 , y11907 , y11908 , y11909 , y11910 , y11911 , y11912 , y11913 , y11914 , y11915 , y11916 , y11917 , y11918 , y11919 , y11920 , y11921 , y11922 , y11923 , y11924 , y11925 , y11926 , y11927 , y11928 , y11929 , y11930 , y11931 , y11932 , y11933 , y11934 , y11935 , y11936 , y11937 , y11938 , y11939 , y11940 , y11941 , y11942 , y11943 , y11944 , y11945 , y11946 , y11947 , y11948 , y11949 , y11950 , y11951 , y11952 , y11953 , y11954 , y11955 , y11956 , y11957 , y11958 , y11959 , y11960 , y11961 , y11962 , y11963 , y11964 , y11965 , y11966 , y11967 , y11968 , y11969 , y11970 , y11971 , y11972 , y11973 , y11974 , y11975 , y11976 , y11977 , y11978 , y11979 , y11980 , y11981 , y11982 , y11983 , y11984 , y11985 , y11986 , y11987 , y11988 , y11989 , y11990 , y11991 , y11992 , y11993 , y11994 , y11995 , y11996 , y11997 , y11998 , y11999 , y12000 , y12001 , y12002 , y12003 , y12004 , y12005 , y12006 , y12007 , y12008 , y12009 , y12010 , y12011 , y12012 , y12013 , y12014 , y12015 , y12016 , y12017 , y12018 , y12019 , y12020 , y12021 , y12022 , y12023 , y12024 , y12025 , y12026 , y12027 , y12028 , y12029 , y12030 , y12031 , y12032 , y12033 , y12034 , y12035 , y12036 , y12037 , y12038 , y12039 , y12040 , y12041 , y12042 , y12043 , y12044 , y12045 , y12046 , y12047 , y12048 , y12049 , y12050 , y12051 , y12052 , y12053 , y12054 , y12055 , y12056 , y12057 , y12058 , y12059 , y12060 , y12061 , y12062 , y12063 , y12064 , y12065 , y12066 , y12067 , y12068 , y12069 , y12070 , y12071 , y12072 , y12073 , y12074 , y12075 , y12076 , y12077 , y12078 , y12079 , y12080 , y12081 , y12082 , y12083 , y12084 , y12085 , y12086 , y12087 , y12088 , y12089 , y12090 , y12091 , y12092 , y12093 , y12094 , y12095 , y12096 , y12097 , y12098 , y12099 , y12100 , y12101 , y12102 , y12103 , y12104 , y12105 , y12106 , y12107 , y12108 , y12109 , y12110 , y12111 , y12112 , y12113 , y12114 , y12115 , y12116 , y12117 , y12118 , y12119 , y12120 , y12121 , y12122 , y12123 , y12124 , y12125 , y12126 , y12127 , y12128 , y12129 , y12130 , y12131 , y12132 , y12133 , y12134 , y12135 , y12136 , y12137 , y12138 , y12139 , y12140 , y12141 , y12142 , y12143 , y12144 , y12145 , y12146 , y12147 , y12148 , y12149 , y12150 , y12151 , y12152 , y12153 , y12154 , y12155 , y12156 , y12157 , y12158 , y12159 , y12160 , y12161 , y12162 , y12163 , y12164 , y12165 , y12166 , y12167 , y12168 , y12169 , y12170 , y12171 , y12172 , y12173 , y12174 , y12175 , y12176 , y12177 , y12178 , y12179 , y12180 , y12181 , y12182 , y12183 , y12184 , y12185 , y12186 , y12187 , y12188 , y12189 , y12190 , y12191 , y12192 , y12193 , y12194 , y12195 , y12196 , y12197 , y12198 , y12199 , y12200 , y12201 , y12202 , y12203 , y12204 , y12205 , y12206 , y12207 , y12208 , y12209 , y12210 , y12211 , y12212 , y12213 , y12214 , y12215 , y12216 , y12217 , y12218 , y12219 , y12220 , y12221 , y12222 , y12223 , y12224 , y12225 , y12226 , y12227 , y12228 , y12229 , y12230 , y12231 , y12232 , y12233 , y12234 , y12235 , y12236 , y12237 , y12238 , y12239 , y12240 , y12241 , y12242 , y12243 , y12244 , y12245 , y12246 , y12247 , y12248 , y12249 , y12250 , y12251 , y12252 , y12253 , y12254 , y12255 , y12256 , y12257 , y12258 , y12259 , y12260 , y12261 , y12262 , y12263 , y12264 , y12265 , y12266 , y12267 , y12268 , y12269 , y12270 , y12271 , y12272 , y12273 , y12274 , y12275 , y12276 , y12277 , y12278 , y12279 , y12280 , y12281 , y12282 , y12283 , y12284 , y12285 , y12286 , y12287 , y12288 , y12289 , y12290 , y12291 , y12292 , y12293 , y12294 , y12295 , y12296 , y12297 , y12298 , y12299 , y12300 , y12301 , y12302 , y12303 , y12304 , y12305 , y12306 , y12307 , y12308 , y12309 , y12310 , y12311 , y12312 , y12313 , y12314 , y12315 , y12316 , y12317 , y12318 , y12319 , y12320 , y12321 , y12322 , y12323 , y12324 , y12325 , y12326 , y12327 , y12328 , y12329 , y12330 , y12331 , y12332 , y12333 , y12334 , y12335 , y12336 , y12337 , y12338 , y12339 , y12340 , y12341 , y12342 , y12343 , y12344 , y12345 , y12346 , y12347 , y12348 , y12349 , y12350 , y12351 , y12352 , y12353 , y12354 , y12355 , y12356 , y12357 , y12358 , y12359 , y12360 , y12361 , y12362 , y12363 , y12364 , y12365 , y12366 , y12367 , y12368 , y12369 , y12370 , y12371 , y12372 , y12373 , y12374 , y12375 , y12376 , y12377 , y12378 , y12379 , y12380 , y12381 , y12382 , y12383 , y12384 , y12385 , y12386 , y12387 , y12388 , y12389 , y12390 , y12391 , y12392 , y12393 , y12394 , y12395 , y12396 , y12397 , y12398 , y12399 , y12400 , y12401 , y12402 , y12403 , y12404 , y12405 , y12406 , y12407 , y12408 , y12409 , y12410 , y12411 , y12412 , y12413 , y12414 , y12415 , y12416 , y12417 , y12418 , y12419 , y12420 , y12421 , y12422 , y12423 , y12424 , y12425 , y12426 , y12427 , y12428 , y12429 , y12430 , y12431 , y12432 , y12433 , y12434 , y12435 , y12436 , y12437 , y12438 , y12439 , y12440 , y12441 , y12442 , y12443 , y12444 , y12445 , y12446 , y12447 , y12448 , y12449 , y12450 , y12451 , y12452 , y12453 , y12454 , y12455 , y12456 , y12457 , y12458 , y12459 , y12460 , y12461 , y12462 , y12463 , y12464 , y12465 , y12466 , y12467 , y12468 , y12469 , y12470 , y12471 , y12472 , y12473 , y12474 , y12475 , y12476 , y12477 , y12478 , y12479 , y12480 , y12481 , y12482 , y12483 , y12484 , y12485 , y12486 , y12487 , y12488 , y12489 , y12490 , y12491 , y12492 , y12493 , y12494 , y12495 , y12496 , y12497 , y12498 , y12499 , y12500 , y12501 , y12502 , y12503 , y12504 , y12505 , y12506 , y12507 , y12508 , y12509 , y12510 , y12511 , y12512 , y12513 , y12514 , y12515 , y12516 , y12517 , y12518 , y12519 , y12520 , y12521 , y12522 , y12523 , y12524 , y12525 , y12526 , y12527 , y12528 , y12529 , y12530 , y12531 , y12532 , y12533 , y12534 , y12535 , y12536 , y12537 , y12538 , y12539 , y12540 , y12541 , y12542 , y12543 , y12544 , y12545 , y12546 , y12547 , y12548 , y12549 , y12550 , y12551 , y12552 , y12553 , y12554 , y12555 , y12556 , y12557 , y12558 , y12559 , y12560 , y12561 , y12562 , y12563 , y12564 , y12565 , y12566 , y12567 , y12568 , y12569 , y12570 , y12571 , y12572 , y12573 , y12574 , y12575 , y12576 , y12577 , y12578 , y12579 , y12580 , y12581 , y12582 , y12583 , y12584 , y12585 , y12586 , y12587 , y12588 , y12589 , y12590 , y12591 , y12592 , y12593 , y12594 , y12595 , y12596 , y12597 , y12598 , y12599 , y12600 , y12601 , y12602 , y12603 , y12604 , y12605 , y12606 , y12607 , y12608 , y12609 , y12610 , y12611 , y12612 , y12613 , y12614 , y12615 , y12616 , y12617 , y12618 , y12619 , y12620 , y12621 , y12622 , y12623 , y12624 , y12625 , y12626 , y12627 , y12628 , y12629 , y12630 , y12631 , y12632 , y12633 , y12634 , y12635 , y12636 , y12637 , y12638 , y12639 , y12640 , y12641 , y12642 , y12643 , y12644 , y12645 , y12646 , y12647 , y12648 , y12649 , y12650 , y12651 , y12652 , y12653 , y12654 , y12655 , y12656 , y12657 , y12658 , y12659 , y12660 , y12661 , y12662 , y12663 , y12664 , y12665 , y12666 , y12667 , y12668 , y12669 , y12670 , y12671 , y12672 , y12673 , y12674 , y12675 , y12676 , y12677 , y12678 , y12679 , y12680 , y12681 , y12682 , y12683 , y12684 , y12685 , y12686 , y12687 , y12688 , y12689 , y12690 , y12691 , y12692 , y12693 , y12694 , y12695 , y12696 , y12697 , y12698 , y12699 , y12700 , y12701 , y12702 , y12703 , y12704 , y12705 , y12706 , y12707 , y12708 , y12709 , y12710 , y12711 , y12712 , y12713 , y12714 , y12715 , y12716 , y12717 , y12718 , y12719 , y12720 , y12721 , y12722 , y12723 , y12724 , y12725 , y12726 , y12727 , y12728 , y12729 , y12730 , y12731 , y12732 , y12733 , y12734 , y12735 , y12736 , y12737 , y12738 , y12739 , y12740 , y12741 , y12742 , y12743 , y12744 , y12745 , y12746 , y12747 , y12748 , y12749 , y12750 , y12751 , y12752 , y12753 , y12754 , y12755 , y12756 , y12757 , y12758 , y12759 , y12760 , y12761 , y12762 , y12763 , y12764 , y12765 , y12766 , y12767 , y12768 , y12769 , y12770 , y12771 , y12772 , y12773 , y12774 , y12775 , y12776 , y12777 , y12778 , y12779 , y12780 , y12781 , y12782 , y12783 , y12784 , y12785 , y12786 , y12787 , y12788 , y12789 , y12790 , y12791 , y12792 , y12793 , y12794 , y12795 , y12796 , y12797 , y12798 , y12799 , y12800 , y12801 , y12802 , y12803 , y12804 , y12805 , y12806 , y12807 , y12808 , y12809 , y12810 , y12811 , y12812 , y12813 , y12814 , y12815 , y12816 , y12817 , y12818 , y12819 , y12820 , y12821 , y12822 , y12823 , y12824 , y12825 , y12826 , y12827 , y12828 , y12829 , y12830 , y12831 , y12832 , y12833 , y12834 , y12835 , y12836 , y12837 , y12838 , y12839 , y12840 , y12841 , y12842 , y12843 , y12844 , y12845 , y12846 , y12847 , y12848 , y12849 , y12850 , y12851 , y12852 , y12853 , y12854 , y12855 , y12856 , y12857 , y12858 , y12859 , y12860 , y12861 , y12862 , y12863 , y12864 , y12865 , y12866 , y12867 , y12868 , y12869 , y12870 , y12871 , y12872 , y12873 , y12874 , y12875 , y12876 , y12877 , y12878 , y12879 , y12880 , y12881 , y12882 , y12883 , y12884 , y12885 , y12886 , y12887 , y12888 , y12889 , y12890 , y12891 , y12892 , y12893 , y12894 , y12895 , y12896 , y12897 , y12898 , y12899 , y12900 , y12901 , y12902 , y12903 , y12904 , y12905 , y12906 , y12907 , y12908 , y12909 , y12910 , y12911 , y12912 , y12913 , y12914 , y12915 , y12916 , y12917 , y12918 , y12919 , y12920 , y12921 , y12922 , y12923 , y12924 , y12925 , y12926 , y12927 , y12928 , y12929 , y12930 , y12931 , y12932 , y12933 , y12934 , y12935 , y12936 , y12937 , y12938 , y12939 , y12940 , y12941 , y12942 , y12943 , y12944 , y12945 , y12946 , y12947 , y12948 , y12949 , y12950 , y12951 , y12952 , y12953 , y12954 , y12955 , y12956 , y12957 , y12958 , y12959 , y12960 , y12961 , y12962 , y12963 , y12964 , y12965 , y12966 , y12967 , y12968 , y12969 , y12970 , y12971 , y12972 , y12973 , y12974 , y12975 , y12976 , y12977 , y12978 , y12979 , y12980 , y12981 , y12982 , y12983 , y12984 , y12985 , y12986 , y12987 , y12988 , y12989 , y12990 , y12991 , y12992 , y12993 , y12994 , y12995 , y12996 , y12997 , y12998 , y12999 , y13000 , y13001 , y13002 , y13003 , y13004 , y13005 , y13006 , y13007 , y13008 , y13009 , y13010 , y13011 , y13012 , y13013 , y13014 , y13015 , y13016 , y13017 , y13018 , y13019 , y13020 , y13021 , y13022 , y13023 , y13024 , y13025 , y13026 , y13027 , y13028 , y13029 , y13030 , y13031 , y13032 , y13033 , y13034 , y13035 , y13036 , y13037 , y13038 , y13039 , y13040 , y13041 , y13042 , y13043 , y13044 , y13045 , y13046 , y13047 , y13048 , y13049 , y13050 , y13051 , y13052 , y13053 , y13054 , y13055 , y13056 , y13057 , y13058 , y13059 , y13060 , y13061 , y13062 , y13063 , y13064 , y13065 , y13066 , y13067 , y13068 , y13069 , y13070 , y13071 , y13072 , y13073 , y13074 , y13075 , y13076 , y13077 , y13078 , y13079 , y13080 , y13081 , y13082 , y13083 , y13084 , y13085 , y13086 , y13087 , y13088 , y13089 , y13090 , y13091 , y13092 , y13093 , y13094 , y13095 , y13096 , y13097 , y13098 , y13099 , y13100 , y13101 , y13102 , y13103 , y13104 , y13105 , y13106 , y13107 , y13108 , y13109 , y13110 , y13111 , y13112 , y13113 , y13114 , y13115 , y13116 , y13117 , y13118 , y13119 , y13120 , y13121 , y13122 , y13123 , y13124 , y13125 , y13126 , y13127 , y13128 , y13129 , y13130 , y13131 , y13132 , y13133 , y13134 , y13135 , y13136 , y13137 , y13138 , y13139 , y13140 , y13141 , y13142 , y13143 , y13144 , y13145 , y13146 , y13147 , y13148 , y13149 , y13150 , y13151 , y13152 , y13153 , y13154 , y13155 , y13156 , y13157 , y13158 , y13159 , y13160 , y13161 , y13162 , y13163 , y13164 , y13165 , y13166 , y13167 , y13168 , y13169 , y13170 , y13171 , y13172 , y13173 , y13174 , y13175 , y13176 , y13177 , y13178 , y13179 , y13180 , y13181 , y13182 , y13183 , y13184 , y13185 , y13186 , y13187 , y13188 , y13189 , y13190 , y13191 , y13192 , y13193 , y13194 , y13195 , y13196 , y13197 , y13198 , y13199 , y13200 , y13201 , y13202 , y13203 , y13204 , y13205 , y13206 , y13207 , y13208 , y13209 , y13210 , y13211 , y13212 , y13213 , y13214 , y13215 , y13216 , y13217 , y13218 , y13219 , y13220 , y13221 , y13222 , y13223 , y13224 , y13225 , y13226 , y13227 , y13228 , y13229 , y13230 , y13231 , y13232 , y13233 , y13234 , y13235 , y13236 , y13237 , y13238 , y13239 , y13240 , y13241 , y13242 , y13243 , y13244 , y13245 , y13246 , y13247 , y13248 , y13249 , y13250 , y13251 , y13252 , y13253 , y13254 , y13255 , y13256 , y13257 , y13258 , y13259 , y13260 , y13261 , y13262 , y13263 , y13264 , y13265 , y13266 , y13267 , y13268 , y13269 , y13270 , y13271 , y13272 , y13273 , y13274 , y13275 , y13276 , y13277 , y13278 , y13279 , y13280 , y13281 , y13282 , y13283 , y13284 , y13285 , y13286 , y13287 , y13288 , y13289 , y13290 , y13291 , y13292 , y13293 , y13294 , y13295 , y13296 , y13297 , y13298 , y13299 , y13300 , y13301 , y13302 , y13303 , y13304 , y13305 , y13306 , y13307 , y13308 , y13309 , y13310 , y13311 , y13312 , y13313 , y13314 , y13315 , y13316 , y13317 , y13318 , y13319 , y13320 , y13321 , y13322 , y13323 , y13324 , y13325 , y13326 , y13327 , y13328 , y13329 , y13330 , y13331 , y13332 , y13333 , y13334 , y13335 , y13336 , y13337 , y13338 , y13339 , y13340 , y13341 , y13342 , y13343 , y13344 , y13345 , y13346 , y13347 , y13348 , y13349 , y13350 , y13351 , y13352 , y13353 , y13354 , y13355 , y13356 , y13357 , y13358 , y13359 , y13360 , y13361 , y13362 , y13363 , y13364 , y13365 , y13366 , y13367 , y13368 , y13369 , y13370 , y13371 , y13372 , y13373 , y13374 , y13375 , y13376 , y13377 , y13378 , y13379 , y13380 , y13381 , y13382 , y13383 , y13384 , y13385 , y13386 , y13387 , y13388 , y13389 , y13390 , y13391 , y13392 , y13393 , y13394 , y13395 , y13396 , y13397 , y13398 , y13399 , y13400 , y13401 , y13402 , y13403 , y13404 , y13405 , y13406 , y13407 , y13408 , y13409 , y13410 , y13411 , y13412 , y13413 , y13414 , y13415 , y13416 , y13417 , y13418 , y13419 , y13420 , y13421 , y13422 , y13423 , y13424 , y13425 , y13426 , y13427 , y13428 , y13429 , y13430 , y13431 , y13432 , y13433 , y13434 , y13435 , y13436 , y13437 , y13438 , y13439 , y13440 , y13441 , y13442 , y13443 , y13444 , y13445 , y13446 , y13447 , y13448 , y13449 , y13450 , y13451 , y13452 , y13453 , y13454 , y13455 , y13456 , y13457 , y13458 , y13459 , y13460 , y13461 , y13462 , y13463 , y13464 , y13465 , y13466 , y13467 , y13468 , y13469 , y13470 , y13471 , y13472 , y13473 , y13474 , y13475 , y13476 , y13477 , y13478 , y13479 , y13480 , y13481 , y13482 , y13483 , y13484 , y13485 , y13486 , y13487 , y13488 , y13489 , y13490 , y13491 , y13492 , y13493 , y13494 , y13495 , y13496 , y13497 , y13498 , y13499 , y13500 , y13501 , y13502 , y13503 , y13504 , y13505 , y13506 , y13507 , y13508 , y13509 , y13510 , y13511 , y13512 , y13513 , y13514 , y13515 , y13516 , y13517 , y13518 , y13519 , y13520 , y13521 , y13522 , y13523 , y13524 , y13525 , y13526 , y13527 , y13528 , y13529 , y13530 , y13531 , y13532 , y13533 , y13534 , y13535 , y13536 , y13537 , y13538 , y13539 , y13540 , y13541 , y13542 , y13543 , y13544 , y13545 , y13546 , y13547 , y13548 , y13549 , y13550 , y13551 , y13552 , y13553 , y13554 , y13555 , y13556 , y13557 , y13558 , y13559 , y13560 , y13561 , y13562 , y13563 , y13564 , y13565 , y13566 , y13567 , y13568 , y13569 , y13570 , y13571 , y13572 , y13573 , y13574 , y13575 , y13576 , y13577 , y13578 , y13579 , y13580 , y13581 , y13582 , y13583 , y13584 , y13585 , y13586 , y13587 , y13588 , y13589 , y13590 , y13591 , y13592 , y13593 , y13594 , y13595 , y13596 , y13597 , y13598 , y13599 , y13600 , y13601 , y13602 , y13603 , y13604 , y13605 , y13606 , y13607 , y13608 , y13609 , y13610 , y13611 , y13612 , y13613 , y13614 , y13615 , y13616 , y13617 , y13618 , y13619 , y13620 , y13621 , y13622 , y13623 , y13624 , y13625 , y13626 , y13627 , y13628 , y13629 , y13630 , y13631 , y13632 , y13633 , y13634 , y13635 , y13636 , y13637 , y13638 , y13639 , y13640 , y13641 , y13642 , y13643 , y13644 , y13645 , y13646 , y13647 , y13648 , y13649 , y13650 , y13651 , y13652 , y13653 , y13654 , y13655 , y13656 , y13657 , y13658 , y13659 , y13660 , y13661 , y13662 , y13663 , y13664 , y13665 , y13666 , y13667 , y13668 , y13669 , y13670 , y13671 , y13672 , y13673 , y13674 , y13675 , y13676 , y13677 , y13678 , y13679 , y13680 , y13681 , y13682 , y13683 , y13684 , y13685 , y13686 , y13687 , y13688 , y13689 , y13690 , y13691 , y13692 , y13693 , y13694 , y13695 , y13696 , y13697 , y13698 , y13699 , y13700 , y13701 , y13702 , y13703 , y13704 , y13705 , y13706 , y13707 , y13708 , y13709 , y13710 , y13711 , y13712 , y13713 , y13714 , y13715 , y13716 , y13717 , y13718 , y13719 , y13720 , y13721 , y13722 , y13723 , y13724 , y13725 , y13726 , y13727 , y13728 , y13729 , y13730 , y13731 , y13732 , y13733 , y13734 , y13735 , y13736 , y13737 , y13738 , y13739 , y13740 , y13741 , y13742 , y13743 , y13744 , y13745 , y13746 , y13747 , y13748 , y13749 , y13750 , y13751 , y13752 , y13753 , y13754 , y13755 , y13756 , y13757 , y13758 , y13759 , y13760 , y13761 , y13762 , y13763 , y13764 , y13765 , y13766 , y13767 , y13768 , y13769 , y13770 , y13771 , y13772 , y13773 , y13774 , y13775 , y13776 , y13777 , y13778 , y13779 , y13780 , y13781 , y13782 , y13783 , y13784 , y13785 , y13786 , y13787 , y13788 , y13789 , y13790 , y13791 , y13792 , y13793 , y13794 , y13795 , y13796 , y13797 , y13798 , y13799 , y13800 , y13801 , y13802 , y13803 , y13804 , y13805 , y13806 , y13807 , y13808 , y13809 , y13810 , y13811 , y13812 , y13813 , y13814 , y13815 , y13816 , y13817 , y13818 , y13819 , y13820 , y13821 , y13822 , y13823 , y13824 , y13825 , y13826 , y13827 , y13828 , y13829 , y13830 , y13831 , y13832 , y13833 , y13834 , y13835 , y13836 , y13837 , y13838 , y13839 , y13840 , y13841 , y13842 , y13843 , y13844 , y13845 , y13846 , y13847 , y13848 , y13849 , y13850 , y13851 , y13852 , y13853 , y13854 , y13855 , y13856 , y13857 , y13858 , y13859 , y13860 , y13861 , y13862 , y13863 , y13864 , y13865 , y13866 , y13867 , y13868 , y13869 , y13870 , y13871 , y13872 , y13873 , y13874 , y13875 , y13876 , y13877 , y13878 , y13879 , y13880 , y13881 , y13882 , y13883 , y13884 , y13885 , y13886 , y13887 , y13888 , y13889 , y13890 , y13891 , y13892 , y13893 , y13894 , y13895 , y13896 , y13897 , y13898 , y13899 , y13900 , y13901 , y13902 , y13903 , y13904 , y13905 , y13906 , y13907 , y13908 , y13909 , y13910 , y13911 , y13912 , y13913 , y13914 , y13915 , y13916 , y13917 , y13918 , y13919 , y13920 , y13921 , y13922 , y13923 , y13924 , y13925 , y13926 , y13927 , y13928 , y13929 , y13930 , y13931 , y13932 , y13933 , y13934 , y13935 , y13936 , y13937 , y13938 , y13939 , y13940 , y13941 , y13942 , y13943 , y13944 , y13945 , y13946 , y13947 , y13948 , y13949 , y13950 , y13951 , y13952 , y13953 , y13954 , y13955 , y13956 , y13957 , y13958 , y13959 , y13960 , y13961 , y13962 , y13963 , y13964 , y13965 , y13966 , y13967 , y13968 , y13969 , y13970 , y13971 , y13972 , y13973 , y13974 , y13975 , y13976 , y13977 , y13978 , y13979 , y13980 , y13981 , y13982 , y13983 , y13984 , y13985 , y13986 , y13987 , y13988 , y13989 , y13990 , y13991 , y13992 , y13993 , y13994 , y13995 , y13996 , y13997 , y13998 , y13999 , y14000 , y14001 , y14002 , y14003 , y14004 , y14005 , y14006 , y14007 , y14008 , y14009 , y14010 , y14011 , y14012 , y14013 , y14014 , y14015 , y14016 , y14017 , y14018 , y14019 , y14020 , y14021 , y14022 , y14023 , y14024 , y14025 , y14026 , y14027 , y14028 , y14029 , y14030 , y14031 , y14032 , y14033 , y14034 , y14035 , y14036 , y14037 , y14038 , y14039 , y14040 , y14041 , y14042 , y14043 , y14044 , y14045 , y14046 , y14047 , y14048 , y14049 , y14050 , y14051 , y14052 , y14053 , y14054 , y14055 , y14056 , y14057 , y14058 , y14059 , y14060 , y14061 , y14062 , y14063 , y14064 , y14065 , y14066 , y14067 , y14068 , y14069 , y14070 , y14071 , y14072 , y14073 , y14074 , y14075 , y14076 , y14077 , y14078 , y14079 , y14080 , y14081 , y14082 , y14083 , y14084 , y14085 , y14086 , y14087 , y14088 , y14089 , y14090 , y14091 , y14092 , y14093 , y14094 , y14095 , y14096 , y14097 , y14098 , y14099 , y14100 , y14101 , y14102 , y14103 , y14104 , y14105 , y14106 , y14107 , y14108 , y14109 , y14110 , y14111 , y14112 , y14113 , y14114 , y14115 , y14116 , y14117 , y14118 , y14119 , y14120 , y14121 , y14122 , y14123 , y14124 , y14125 , y14126 , y14127 , y14128 , y14129 , y14130 , y14131 , y14132 , y14133 , y14134 , y14135 , y14136 , y14137 , y14138 , y14139 , y14140 , y14141 , y14142 , y14143 , y14144 , y14145 , y14146 , y14147 , y14148 , y14149 , y14150 , y14151 , y14152 , y14153 , y14154 , y14155 , y14156 , y14157 , y14158 , y14159 , y14160 , y14161 , y14162 , y14163 , y14164 , y14165 , y14166 , y14167 , y14168 , y14169 , y14170 , y14171 , y14172 , y14173 , y14174 , y14175 , y14176 , y14177 , y14178 , y14179 , y14180 , y14181 , y14182 , y14183 , y14184 , y14185 , y14186 , y14187 , y14188 , y14189 , y14190 , y14191 , y14192 , y14193 , y14194 , y14195 , y14196 , y14197 , y14198 , y14199 , y14200 , y14201 , y14202 , y14203 , y14204 , y14205 , y14206 , y14207 , y14208 , y14209 , y14210 , y14211 , y14212 , y14213 , y14214 , y14215 , y14216 , y14217 , y14218 , y14219 , y14220 , y14221 , y14222 , y14223 , y14224 , y14225 , y14226 , y14227 , y14228 , y14229 , y14230 , y14231 , y14232 , y14233 , y14234 , y14235 , y14236 , y14237 , y14238 , y14239 , y14240 , y14241 , y14242 , y14243 , y14244 , y14245 , y14246 , y14247 , y14248 , y14249 , y14250 , y14251 , y14252 , y14253 , y14254 , y14255 , y14256 , y14257 , y14258 , y14259 , y14260 , y14261 , y14262 , y14263 , y14264 , y14265 , y14266 , y14267 , y14268 , y14269 , y14270 , y14271 , y14272 , y14273 , y14274 , y14275 , y14276 , y14277 , y14278 , y14279 , y14280 , y14281 , y14282 , y14283 , y14284 , y14285 , y14286 , y14287 , y14288 , y14289 , y14290 , y14291 , y14292 , y14293 , y14294 , y14295 , y14296 , y14297 , y14298 , y14299 , y14300 , y14301 , y14302 , y14303 , y14304 , y14305 , y14306 , y14307 , y14308 , y14309 , y14310 , y14311 , y14312 , y14313 , y14314 , y14315 , y14316 , y14317 , y14318 , y14319 , y14320 , y14321 , y14322 , y14323 , y14324 , y14325 , y14326 , y14327 , y14328 , y14329 , y14330 , y14331 , y14332 , y14333 , y14334 , y14335 , y14336 , y14337 , y14338 , y14339 , y14340 , y14341 , y14342 , y14343 , y14344 , y14345 , y14346 , y14347 , y14348 , y14349 , y14350 , y14351 , y14352 , y14353 , y14354 , y14355 , y14356 , y14357 , y14358 , y14359 , y14360 , y14361 , y14362 , y14363 , y14364 , y14365 , y14366 , y14367 , y14368 , y14369 , y14370 , y14371 , y14372 , y14373 , y14374 , y14375 , y14376 , y14377 , y14378 , y14379 , y14380 , y14381 , y14382 , y14383 , y14384 , y14385 , y14386 , y14387 , y14388 , y14389 , y14390 , y14391 , y14392 , y14393 , y14394 , y14395 , y14396 , y14397 , y14398 , y14399 , y14400 , y14401 , y14402 , y14403 , y14404 , y14405 , y14406 , y14407 , y14408 , y14409 , y14410 , y14411 , y14412 , y14413 , y14414 , y14415 , y14416 , y14417 , y14418 , y14419 , y14420 , y14421 , y14422 , y14423 , y14424 , y14425 , y14426 , y14427 , y14428 , y14429 , y14430 , y14431 , y14432 , y14433 , y14434 , y14435 , y14436 , y14437 , y14438 , y14439 , y14440 , y14441 , y14442 , y14443 , y14444 , y14445 , y14446 , y14447 , y14448 , y14449 , y14450 , y14451 , y14452 , y14453 , y14454 , y14455 , y14456 , y14457 , y14458 , y14459 , y14460 , y14461 , y14462 , y14463 , y14464 , y14465 , y14466 , y14467 , y14468 , y14469 , y14470 , y14471 , y14472 , y14473 , y14474 , y14475 , y14476 , y14477 , y14478 , y14479 , y14480 , y14481 , y14482 , y14483 , y14484 , y14485 , y14486 , y14487 , y14488 , y14489 , y14490 , y14491 , y14492 , y14493 , y14494 , y14495 , y14496 , y14497 , y14498 , y14499 , y14500 , y14501 , y14502 , y14503 , y14504 , y14505 , y14506 , y14507 , y14508 , y14509 , y14510 , y14511 , y14512 , y14513 , y14514 , y14515 , y14516 , y14517 , y14518 , y14519 , y14520 , y14521 , y14522 , y14523 , y14524 , y14525 , y14526 , y14527 , y14528 , y14529 , y14530 , y14531 , y14532 , y14533 , y14534 , y14535 , y14536 , y14537 , y14538 , y14539 , y14540 , y14541 , y14542 , y14543 , y14544 , y14545 , y14546 , y14547 , y14548 , y14549 , y14550 , y14551 , y14552 , y14553 , y14554 , y14555 , y14556 , y14557 , y14558 , y14559 , y14560 , y14561 , y14562 , y14563 , y14564 , y14565 , y14566 , y14567 , y14568 , y14569 , y14570 , y14571 , y14572 , y14573 , y14574 , y14575 , y14576 , y14577 , y14578 , y14579 , y14580 , y14581 , y14582 , y14583 , y14584 , y14585 , y14586 , y14587 , y14588 , y14589 , y14590 , y14591 , y14592 , y14593 , y14594 , y14595 , y14596 , y14597 , y14598 , y14599 , y14600 , y14601 , y14602 , y14603 , y14604 , y14605 , y14606 , y14607 , y14608 , y14609 , y14610 , y14611 , y14612 , y14613 , y14614 , y14615 , y14616 , y14617 , y14618 , y14619 , y14620 , y14621 , y14622 , y14623 , y14624 , y14625 , y14626 , y14627 , y14628 , y14629 , y14630 , y14631 , y14632 , y14633 , y14634 , y14635 , y14636 , y14637 , y14638 , y14639 , y14640 , y14641 , y14642 , y14643 , y14644 , y14645 , y14646 , y14647 , y14648 , y14649 , y14650 , y14651 , y14652 , y14653 , y14654 , y14655 , y14656 , y14657 , y14658 , y14659 , y14660 , y14661 , y14662 , y14663 , y14664 , y14665 , y14666 , y14667 , y14668 , y14669 , y14670 , y14671 , y14672 , y14673 , y14674 , y14675 , y14676 , y14677 , y14678 , y14679 , y14680 , y14681 , y14682 , y14683 , y14684 , y14685 , y14686 , y14687 , y14688 , y14689 , y14690 , y14691 , y14692 , y14693 , y14694 , y14695 , y14696 , y14697 , y14698 , y14699 , y14700 , y14701 , y14702 , y14703 , y14704 , y14705 , y14706 , y14707 , y14708 , y14709 , y14710 , y14711 , y14712 , y14713 , y14714 , y14715 , y14716 , y14717 , y14718 , y14719 , y14720 , y14721 , y14722 , y14723 , y14724 , y14725 , y14726 , y14727 , y14728 , y14729 , y14730 , y14731 , y14732 , y14733 , y14734 , y14735 , y14736 , y14737 , y14738 , y14739 , y14740 , y14741 , y14742 , y14743 , y14744 , y14745 , y14746 , y14747 , y14748 , y14749 , y14750 , y14751 , y14752 , y14753 , y14754 , y14755 , y14756 , y14757 , y14758 , y14759 , y14760 , y14761 , y14762 , y14763 , y14764 , y14765 , y14766 , y14767 , y14768 , y14769 , y14770 , y14771 , y14772 , y14773 , y14774 , y14775 , y14776 , y14777 , y14778 , y14779 , y14780 , y14781 , y14782 , y14783 , y14784 , y14785 , y14786 , y14787 , y14788 , y14789 , y14790 , y14791 , y14792 , y14793 , y14794 , y14795 , y14796 , y14797 , y14798 , y14799 , y14800 , y14801 , y14802 , y14803 , y14804 , y14805 , y14806 , y14807 , y14808 , y14809 , y14810 , y14811 , y14812 , y14813 , y14814 , y14815 , y14816 , y14817 , y14818 , y14819 , y14820 , y14821 , y14822 , y14823 , y14824 , y14825 , y14826 , y14827 , y14828 , y14829 , y14830 , y14831 , y14832 , y14833 , y14834 , y14835 , y14836 , y14837 , y14838 , y14839 , y14840 , y14841 , y14842 , y14843 , y14844 , y14845 , y14846 , y14847 , y14848 , y14849 , y14850 , y14851 , y14852 , y14853 , y14854 , y14855 , y14856 , y14857 , y14858 , y14859 , y14860 , y14861 , y14862 , y14863 , y14864 , y14865 , y14866 , y14867 , y14868 , y14869 , y14870 , y14871 , y14872 , y14873 , y14874 , y14875 , y14876 , y14877 , y14878 , y14879 , y14880 , y14881 , y14882 , y14883 , y14884 , y14885 , y14886 , y14887 , y14888 , y14889 , y14890 , y14891 , y14892 , y14893 , y14894 , y14895 , y14896 , y14897 , y14898 , y14899 , y14900 , y14901 , y14902 , y14903 , y14904 , y14905 , y14906 , y14907 , y14908 , y14909 , y14910 , y14911 , y14912 , y14913 , y14914 , y14915 , y14916 , y14917 , y14918 , y14919 , y14920 , y14921 , y14922 , y14923 , y14924 , y14925 , y14926 , y14927 , y14928 , y14929 , y14930 , y14931 , y14932 , y14933 , y14934 , y14935 , y14936 , y14937 , y14938 , y14939 , y14940 , y14941 , y14942 , y14943 , y14944 , y14945 , y14946 , y14947 , y14948 , y14949 , y14950 , y14951 , y14952 , y14953 , y14954 , y14955 , y14956 , y14957 , y14958 , y14959 , y14960 , y14961 , y14962 , y14963 , y14964 , y14965 , y14966 , y14967 , y14968 , y14969 , y14970 , y14971 , y14972 , y14973 , y14974 , y14975 , y14976 , y14977 , y14978 , y14979 , y14980 , y14981 , y14982 , y14983 , y14984 , y14985 , y14986 , y14987 , y14988 , y14989 , y14990 , y14991 , y14992 , y14993 , y14994 , y14995 , y14996 , y14997 , y14998 , y14999 , y15000 , y15001 , y15002 , y15003 , y15004 , y15005 , y15006 , y15007 , y15008 , y15009 , y15010 , y15011 , y15012 , y15013 , y15014 , y15015 , y15016 , y15017 , y15018 , y15019 , y15020 , y15021 , y15022 , y15023 , y15024 , y15025 , y15026 , y15027 , y15028 , y15029 , y15030 , y15031 , y15032 , y15033 , y15034 , y15035 , y15036 , y15037 , y15038 , y15039 , y15040 , y15041 , y15042 , y15043 , y15044 , y15045 , y15046 , y15047 , y15048 , y15049 , y15050 , y15051 , y15052 , y15053 , y15054 , y15055 , y15056 , y15057 , y15058 , y15059 , y15060 , y15061 , y15062 , y15063 , y15064 , y15065 , y15066 , y15067 , y15068 , y15069 , y15070 , y15071 , y15072 , y15073 , y15074 , y15075 , y15076 , y15077 , y15078 , y15079 , y15080 , y15081 , y15082 , y15083 , y15084 , y15085 , y15086 , y15087 , y15088 , y15089 , y15090 , y15091 , y15092 , y15093 , y15094 , y15095 , y15096 , y15097 , y15098 , y15099 , y15100 , y15101 , y15102 , y15103 , y15104 , y15105 , y15106 , y15107 , y15108 , y15109 , y15110 , y15111 , y15112 , y15113 , y15114 , y15115 , y15116 , y15117 , y15118 , y15119 , y15120 , y15121 , y15122 , y15123 , y15124 , y15125 , y15126 , y15127 , y15128 , y15129 , y15130 , y15131 , y15132 , y15133 , y15134 , y15135 , y15136 , y15137 , y15138 , y15139 , y15140 , y15141 , y15142 , y15143 , y15144 , y15145 , y15146 , y15147 , y15148 , y15149 , y15150 , y15151 , y15152 , y15153 , y15154 , y15155 , y15156 , y15157 , y15158 , y15159 , y15160 , y15161 , y15162 , y15163 , y15164 , y15165 , y15166 , y15167 , y15168 , y15169 , y15170 , y15171 , y15172 , y15173 , y15174 , y15175 , y15176 , y15177 , y15178 , y15179 , y15180 , y15181 , y15182 , y15183 , y15184 , y15185 , y15186 , y15187 , y15188 , y15189 , y15190 , y15191 , y15192 , y15193 , y15194 , y15195 , y15196 , y15197 , y15198 , y15199 , y15200 , y15201 , y15202 , y15203 , y15204 , y15205 , y15206 , y15207 , y15208 , y15209 , y15210 , y15211 , y15212 , y15213 , y15214 , y15215 , y15216 , y15217 , y15218 , y15219 , y15220 , y15221 , y15222 , y15223 , y15224 , y15225 , y15226 , y15227 , y15228 , y15229 , y15230 , y15231 , y15232 , y15233 , y15234 , y15235 , y15236 , y15237 , y15238 , y15239 , y15240 , y15241 , y15242 , y15243 , y15244 , y15245 , y15246 , y15247 , y15248 , y15249 , y15250 , y15251 , y15252 , y15253 , y15254 , y15255 , y15256 , y15257 , y15258 , y15259 , y15260 , y15261 , y15262 , y15263 , y15264 , y15265 , y15266 , y15267 , y15268 , y15269 , y15270 , y15271 , y15272 , y15273 , y15274 , y15275 , y15276 , y15277 , y15278 , y15279 , y15280 , y15281 , y15282 , y15283 , y15284 , y15285 , y15286 , y15287 , y15288 , y15289 , y15290 , y15291 , y15292 , y15293 , y15294 , y15295 , y15296 , y15297 , y15298 , y15299 , y15300 , y15301 , y15302 , y15303 , y15304 , y15305 , y15306 , y15307 , y15308 , y15309 , y15310 , y15311 , y15312 , y15313 , y15314 , y15315 , y15316 , y15317 , y15318 , y15319 , y15320 , y15321 , y15322 , y15323 , y15324 , y15325 , y15326 , y15327 , y15328 , y15329 , y15330 , y15331 , y15332 , y15333 , y15334 , y15335 , y15336 , y15337 , y15338 , y15339 , y15340 , y15341 , y15342 , y15343 , y15344 , y15345 , y15346 , y15347 , y15348 , y15349 , y15350 , y15351 , y15352 , y15353 , y15354 , y15355 , y15356 , y15357 , y15358 , y15359 , y15360 , y15361 , y15362 , y15363 , y15364 , y15365 , y15366 , y15367 , y15368 , y15369 , y15370 , y15371 , y15372 , y15373 , y15374 , y15375 , y15376 , y15377 , y15378 , y15379 , y15380 , y15381 , y15382 , y15383 , y15384 , y15385 , y15386 , y15387 , y15388 , y15389 , y15390 , y15391 , y15392 , y15393 , y15394 , y15395 , y15396 , y15397 , y15398 , y15399 , y15400 , y15401 , y15402 , y15403 , y15404 , y15405 , y15406 , y15407 , y15408 , y15409 , y15410 , y15411 , y15412 , y15413 , y15414 , y15415 , y15416 , y15417 , y15418 , y15419 , y15420 , y15421 , y15422 , y15423 , y15424 , y15425 , y15426 , y15427 , y15428 , y15429 , y15430 , y15431 , y15432 , y15433 , y15434 , y15435 , y15436 , y15437 , y15438 , y15439 , y15440 , y15441 , y15442 , y15443 , y15444 , y15445 , y15446 , y15447 , y15448 , y15449 , y15450 , y15451 , y15452 , y15453 , y15454 , y15455 , y15456 , y15457 , y15458 , y15459 , y15460 , y15461 , y15462 , y15463 , y15464 , y15465 , y15466 , y15467 , y15468 , y15469 , y15470 , y15471 , y15472 , y15473 , y15474 , y15475 , y15476 , y15477 , y15478 , y15479 , y15480 , y15481 , y15482 , y15483 , y15484 , y15485 , y15486 , y15487 , y15488 , y15489 , y15490 , y15491 , y15492 , y15493 , y15494 , y15495 , y15496 , y15497 , y15498 , y15499 , y15500 , y15501 , y15502 , y15503 , y15504 , y15505 , y15506 , y15507 , y15508 , y15509 , y15510 , y15511 , y15512 , y15513 , y15514 , y15515 , y15516 , y15517 , y15518 , y15519 , y15520 , y15521 , y15522 , y15523 , y15524 , y15525 , y15526 , y15527 , y15528 , y15529 , y15530 , y15531 , y15532 , y15533 , y15534 , y15535 , y15536 , y15537 , y15538 , y15539 , y15540 , y15541 , y15542 , y15543 , y15544 , y15545 , y15546 , y15547 , y15548 , y15549 , y15550 , y15551 , y15552 , y15553 , y15554 , y15555 , y15556 , y15557 , y15558 , y15559 , y15560 , y15561 , y15562 , y15563 , y15564 , y15565 , y15566 , y15567 , y15568 , y15569 , y15570 , y15571 , y15572 , y15573 , y15574 , y15575 , y15576 , y15577 , y15578 , y15579 , y15580 , y15581 , y15582 , y15583 , y15584 , y15585 , y15586 , y15587 , y15588 , y15589 , y15590 , y15591 , y15592 , y15593 , y15594 , y15595 , y15596 , y15597 , y15598 , y15599 , y15600 , y15601 , y15602 , y15603 , y15604 , y15605 , y15606 , y15607 , y15608 , y15609 , y15610 , y15611 , y15612 , y15613 , y15614 , y15615 , y15616 , y15617 , y15618 , y15619 , y15620 , y15621 , y15622 , y15623 , y15624 , y15625 , y15626 , y15627 , y15628 , y15629 , y15630 , y15631 , y15632 , y15633 , y15634 , y15635 , y15636 , y15637 , y15638 , y15639 , y15640 , y15641 , y15642 , y15643 , y15644 , y15645 , y15646 , y15647 , y15648 , y15649 , y15650 , y15651 , y15652 , y15653 , y15654 , y15655 , y15656 , y15657 , y15658 , y15659 , y15660 , y15661 , y15662 , y15663 , y15664 , y15665 , y15666 , y15667 , y15668 , y15669 , y15670 , y15671 , y15672 , y15673 , y15674 , y15675 , y15676 , y15677 , y15678 , y15679 , y15680 , y15681 , y15682 , y15683 , y15684 , y15685 , y15686 , y15687 , y15688 , y15689 , y15690 , y15691 , y15692 , y15693 , y15694 , y15695 , y15696 , y15697 , y15698 , y15699 , y15700 , y15701 , y15702 , y15703 , y15704 , y15705 , y15706 , y15707 , y15708 , y15709 , y15710 , y15711 , y15712 , y15713 , y15714 , y15715 , y15716 , y15717 , y15718 , y15719 , y15720 , y15721 , y15722 , y15723 , y15724 , y15725 , y15726 , y15727 , y15728 , y15729 , y15730 , y15731 , y15732 , y15733 , y15734 , y15735 , y15736 , y15737 , y15738 , y15739 , y15740 , y15741 , y15742 , y15743 , y15744 , y15745 , y15746 , y15747 , y15748 , y15749 , y15750 , y15751 , y15752 , y15753 , y15754 , y15755 , y15756 , y15757 , y15758 , y15759 , y15760 , y15761 , y15762 , y15763 , y15764 , y15765 , y15766 , y15767 , y15768 , y15769 , y15770 , y15771 , y15772 , y15773 , y15774 , y15775 , y15776 , y15777 , y15778 , y15779 , y15780 , y15781 , y15782 , y15783 , y15784 , y15785 , y15786 , y15787 , y15788 , y15789 , y15790 , y15791 , y15792 , y15793 , y15794 , y15795 , y15796 , y15797 , y15798 , y15799 , y15800 , y15801 , y15802 , y15803 , y15804 , y15805 , y15806 , y15807 , y15808 , y15809 , y15810 , y15811 , y15812 , y15813 , y15814 , y15815 , y15816 , y15817 , y15818 , y15819 , y15820 , y15821 , y15822 , y15823 , y15824 , y15825 , y15826 , y15827 , y15828 , y15829 , y15830 , y15831 , y15832 , y15833 , y15834 , y15835 , y15836 , y15837 , y15838 , y15839 , y15840 , y15841 , y15842 , y15843 , y15844 , y15845 , y15846 , y15847 , y15848 , y15849 , y15850 , y15851 , y15852 , y15853 , y15854 , y15855 , y15856 , y15857 , y15858 , y15859 , y15860 , y15861 , y15862 , y15863 , y15864 , y15865 , y15866 , y15867 , y15868 , y15869 , y15870 , y15871 , y15872 , y15873 , y15874 , y15875 , y15876 , y15877 , y15878 , y15879 , y15880 , y15881 , y15882 , y15883 , y15884 , y15885 , y15886 , y15887 , y15888 , y15889 , y15890 , y15891 , y15892 , y15893 , y15894 , y15895 , y15896 , y15897 , y15898 , y15899 , y15900 , y15901 , y15902 , y15903 , y15904 , y15905 , y15906 , y15907 , y15908 , y15909 , y15910 , y15911 , y15912 , y15913 , y15914 , y15915 , y15916 , y15917 , y15918 , y15919 , y15920 , y15921 , y15922 , y15923 , y15924 , y15925 , y15926 , y15927 , y15928 , y15929 , y15930 , y15931 , y15932 , y15933 , y15934 , y15935 , y15936 , y15937 , y15938 , y15939 , y15940 , y15941 , y15942 , y15943 , y15944 , y15945 , y15946 , y15947 , y15948 , y15949 , y15950 , y15951 , y15952 , y15953 , y15954 , y15955 , y15956 , y15957 , y15958 , y15959 , y15960 , y15961 , y15962 , y15963 , y15964 , y15965 , y15966 , y15967 , y15968 , y15969 , y15970 , y15971 , y15972 , y15973 , y15974 , y15975 , y15976 , y15977 , y15978 , y15979 , y15980 , y15981 , y15982 , y15983 , y15984 , y15985 , y15986 , y15987 , y15988 , y15989 , y15990 , y15991 , y15992 , y15993 , y15994 , y15995 , y15996 , y15997 , y15998 , y15999 , y16000 , y16001 , y16002 , y16003 , y16004 , y16005 , y16006 , y16007 , y16008 , y16009 , y16010 , y16011 , y16012 , y16013 , y16014 , y16015 , y16016 , y16017 , y16018 , y16019 , y16020 , y16021 , y16022 , y16023 , y16024 , y16025 , y16026 , y16027 , y16028 , y16029 , y16030 , y16031 , y16032 , y16033 , y16034 , y16035 , y16036 , y16037 , y16038 , y16039 , y16040 , y16041 , y16042 , y16043 , y16044 , y16045 , y16046 , y16047 , y16048 , y16049 , y16050 , y16051 , y16052 , y16053 , y16054 , y16055 , y16056 , y16057 , y16058 , y16059 , y16060 , y16061 , y16062 , y16063 , y16064 , y16065 , y16066 , y16067 , y16068 , y16069 , y16070 , y16071 , y16072 , y16073 , y16074 , y16075 , y16076 , y16077 , y16078 , y16079 , y16080 , y16081 , y16082 , y16083 , y16084 , y16085 , y16086 , y16087 , y16088 , y16089 , y16090 , y16091 , y16092 , y16093 , y16094 , y16095 , y16096 , y16097 , y16098 , y16099 , y16100 , y16101 , y16102 , y16103 , y16104 , y16105 , y16106 , y16107 , y16108 , y16109 , y16110 , y16111 , y16112 , y16113 , y16114 , y16115 , y16116 , y16117 , y16118 , y16119 , y16120 , y16121 , y16122 , y16123 , y16124 , y16125 , y16126 , y16127 , y16128 , y16129 , y16130 , y16131 , y16132 , y16133 , y16134 , y16135 , y16136 , y16137 , y16138 , y16139 , y16140 , y16141 , y16142 , y16143 , y16144 , y16145 , y16146 , y16147 , y16148 , y16149 , y16150 , y16151 , y16152 , y16153 , y16154 , y16155 , y16156 , y16157 , y16158 , y16159 , y16160 , y16161 , y16162 , y16163 , y16164 , y16165 , y16166 , y16167 , y16168 , y16169 , y16170 , y16171 , y16172 , y16173 , y16174 , y16175 , y16176 , y16177 , y16178 , y16179 , y16180 , y16181 , y16182 , y16183 , y16184 , y16185 , y16186 , y16187 , y16188 , y16189 , y16190 , y16191 , y16192 , y16193 , y16194 , y16195 , y16196 , y16197 , y16198 , y16199 , y16200 , y16201 , y16202 , y16203 , y16204 , y16205 , y16206 , y16207 , y16208 , y16209 , y16210 , y16211 , y16212 , y16213 , y16214 , y16215 , y16216 , y16217 , y16218 , y16219 , y16220 , y16221 , y16222 , y16223 , y16224 , y16225 , y16226 , y16227 , y16228 , y16229 , y16230 , y16231 , y16232 , y16233 , y16234 , y16235 , y16236 , y16237 , y16238 , y16239 , y16240 , y16241 , y16242 , y16243 , y16244 , y16245 , y16246 , y16247 , y16248 , y16249 , y16250 , y16251 , y16252 , y16253 , y16254 , y16255 , y16256 , y16257 , y16258 , y16259 , y16260 , y16261 , y16262 , y16263 , y16264 , y16265 , y16266 , y16267 , y16268 , y16269 , y16270 , y16271 , y16272 , y16273 , y16274 , y16275 , y16276 , y16277 , y16278 , y16279 , y16280 , y16281 , y16282 , y16283 , y16284 , y16285 , y16286 , y16287 , y16288 , y16289 , y16290 , y16291 , y16292 , y16293 , y16294 , y16295 , y16296 , y16297 , y16298 , y16299 , y16300 , y16301 , y16302 , y16303 , y16304 , y16305 , y16306 , y16307 , y16308 , y16309 , y16310 , y16311 , y16312 , y16313 , y16314 , y16315 , y16316 , y16317 , y16318 , y16319 , y16320 , y16321 , y16322 , y16323 , y16324 , y16325 , y16326 , y16327 , y16328 , y16329 , y16330 , y16331 , y16332 , y16333 , y16334 , y16335 , y16336 , y16337 , y16338 , y16339 , y16340 , y16341 , y16342 , y16343 , y16344 , y16345 , y16346 , y16347 , y16348 , y16349 , y16350 , y16351 , y16352 , y16353 , y16354 , y16355 , y16356 , y16357 , y16358 , y16359 , y16360 , y16361 , y16362 , y16363 , y16364 , y16365 , y16366 , y16367 , y16368 , y16369 , y16370 , y16371 , y16372 , y16373 , y16374 , y16375 , y16376 , y16377 , y16378 , y16379 , y16380 , y16381 , y16382 , y16383 , y16384 , y16385 , y16386 , y16387 , y16388 , y16389 , y16390 , y16391 , y16392 , y16393 , y16394 , y16395 , y16396 , y16397 , y16398 , y16399 , y16400 , y16401 , y16402 , y16403 , y16404 , y16405 , y16406 , y16407 , y16408 , y16409 , y16410 , y16411 , y16412 , y16413 , y16414 , y16415 , y16416 , y16417 , y16418 , y16419 , y16420 , y16421 , y16422 , y16423 , y16424 , y16425 , y16426 , y16427 , y16428 , y16429 , y16430 , y16431 , y16432 , y16433 , y16434 , y16435 , y16436 , y16437 , y16438 , y16439 , y16440 , y16441 , y16442 , y16443 , y16444 , y16445 , y16446 , y16447 , y16448 , y16449 , y16450 , y16451 , y16452 , y16453 , y16454 , y16455 , y16456 , y16457 , y16458 , y16459 , y16460 , y16461 , y16462 , y16463 , y16464 , y16465 , y16466 , y16467 , y16468 , y16469 , y16470 , y16471 , y16472 , y16473 , y16474 , y16475 , y16476 , y16477 , y16478 , y16479 , y16480 , y16481 , y16482 , y16483 , y16484 , y16485 , y16486 , y16487 , y16488 , y16489 , y16490 , y16491 , y16492 , y16493 , y16494 , y16495 , y16496 , y16497 , y16498 , y16499 , y16500 , y16501 , y16502 , y16503 , y16504 , y16505 , y16506 , y16507 , y16508 , y16509 , y16510 , y16511 , y16512 , y16513 , y16514 , y16515 , y16516 , y16517 , y16518 , y16519 , y16520 , y16521 , y16522 , y16523 , y16524 , y16525 , y16526 , y16527 , y16528 , y16529 , y16530 , y16531 , y16532 , y16533 , y16534 , y16535 , y16536 , y16537 , y16538 , y16539 , y16540 , y16541 , y16542 , y16543 , y16544 , y16545 , y16546 , y16547 , y16548 , y16549 , y16550 , y16551 , y16552 , y16553 , y16554 , y16555 , y16556 , y16557 , y16558 , y16559 , y16560 , y16561 , y16562 , y16563 , y16564 , y16565 , y16566 , y16567 , y16568 , y16569 , y16570 , y16571 , y16572 , y16573 , y16574 , y16575 , y16576 , y16577 , y16578 , y16579 , y16580 , y16581 , y16582 , y16583 , y16584 , y16585 , y16586 , y16587 , y16588 , y16589 , y16590 , y16591 , y16592 , y16593 , y16594 , y16595 , y16596 , y16597 , y16598 , y16599 , y16600 , y16601 , y16602 , y16603 , y16604 , y16605 , y16606 , y16607 , y16608 , y16609 , y16610 , y16611 , y16612 , y16613 , y16614 , y16615 , y16616 , y16617 , y16618 , y16619 , y16620 , y16621 , y16622 , y16623 , y16624 , y16625 , y16626 , y16627 , y16628 , y16629 , y16630 , y16631 , y16632 , y16633 , y16634 , y16635 , y16636 , y16637 , y16638 , y16639 , y16640 , y16641 , y16642 , y16643 , y16644 , y16645 , y16646 , y16647 , y16648 , y16649 , y16650 , y16651 , y16652 , y16653 , y16654 , y16655 , y16656 , y16657 , y16658 , y16659 , y16660 , y16661 , y16662 , y16663 , y16664 , y16665 , y16666 , y16667 , y16668 , y16669 , y16670 , y16671 , y16672 , y16673 , y16674 , y16675 , y16676 , y16677 , y16678 , y16679 , y16680 , y16681 , y16682 , y16683 , y16684 , y16685 , y16686 , y16687 , y16688 , y16689 , y16690 , y16691 , y16692 , y16693 , y16694 , y16695 , y16696 , y16697 , y16698 , y16699 , y16700 , y16701 , y16702 , y16703 , y16704 , y16705 , y16706 , y16707 , y16708 , y16709 , y16710 , y16711 , y16712 , y16713 , y16714 , y16715 , y16716 , y16717 , y16718 , y16719 , y16720 , y16721 , y16722 , y16723 , y16724 , y16725 , y16726 , y16727 , y16728 , y16729 , y16730 , y16731 , y16732 , y16733 , y16734 , y16735 , y16736 , y16737 , y16738 , y16739 , y16740 , y16741 , y16742 , y16743 , y16744 , y16745 , y16746 , y16747 , y16748 , y16749 , y16750 , y16751 , y16752 , y16753 , y16754 , y16755 , y16756 , y16757 , y16758 , y16759 , y16760 , y16761 , y16762 , y16763 , y16764 , y16765 , y16766 , y16767 , y16768 , y16769 , y16770 , y16771 , y16772 , y16773 , y16774 , y16775 , y16776 , y16777 , y16778 , y16779 , y16780 , y16781 , y16782 , y16783 , y16784 , y16785 , y16786 , y16787 , y16788 , y16789 , y16790 , y16791 , y16792 , y16793 , y16794 , y16795 , y16796 , y16797 , y16798 , y16799 , y16800 , y16801 , y16802 , y16803 , y16804 , y16805 , y16806 , y16807 , y16808 , y16809 , y16810 , y16811 , y16812 , y16813 , y16814 , y16815 , y16816 , y16817 , y16818 , y16819 , y16820 , y16821 , y16822 , y16823 , y16824 , y16825 , y16826 , y16827 , y16828 , y16829 , y16830 , y16831 , y16832 , y16833 , y16834 , y16835 , y16836 , y16837 , y16838 , y16839 , y16840 , y16841 , y16842 , y16843 , y16844 , y16845 , y16846 , y16847 , y16848 , y16849 , y16850 , y16851 , y16852 , y16853 , y16854 , y16855 , y16856 , y16857 , y16858 , y16859 , y16860 , y16861 , y16862 , y16863 , y16864 , y16865 , y16866 , y16867 , y16868 , y16869 , y16870 , y16871 , y16872 , y16873 , y16874 , y16875 , y16876 , y16877 , y16878 , y16879 , y16880 , y16881 , y16882 , y16883 , y16884 , y16885 , y16886 , y16887 , y16888 , y16889 , y16890 , y16891 , y16892 , y16893 , y16894 , y16895 , y16896 , y16897 , y16898 , y16899 , y16900 , y16901 , y16902 , y16903 , y16904 , y16905 , y16906 , y16907 , y16908 , y16909 , y16910 , y16911 , y16912 , y16913 , y16914 , y16915 , y16916 , y16917 , y16918 , y16919 , y16920 , y16921 , y16922 , y16923 , y16924 , y16925 , y16926 , y16927 , y16928 , y16929 , y16930 , y16931 , y16932 , y16933 , y16934 , y16935 , y16936 , y16937 , y16938 , y16939 , y16940 , y16941 , y16942 , y16943 , y16944 , y16945 , y16946 , y16947 , y16948 , y16949 , y16950 , y16951 , y16952 , y16953 , y16954 , y16955 , y16956 , y16957 , y16958 , y16959 , y16960 , y16961 , y16962 , y16963 , y16964 , y16965 , y16966 , y16967 , y16968 , y16969 , y16970 , y16971 , y16972 , y16973 , y16974 , y16975 , y16976 , y16977 , y16978 , y16979 , y16980 , y16981 , y16982 , y16983 , y16984 , y16985 , y16986 , y16987 , y16988 , y16989 , y16990 , y16991 , y16992 , y16993 , y16994 , y16995 , y16996 , y16997 , y16998 , y16999 , y17000 , y17001 , y17002 , y17003 , y17004 , y17005 , y17006 , y17007 , y17008 , y17009 , y17010 , y17011 , y17012 , y17013 , y17014 , y17015 , y17016 , y17017 , y17018 , y17019 , y17020 , y17021 , y17022 , y17023 , y17024 , y17025 , y17026 , y17027 , y17028 , y17029 , y17030 , y17031 , y17032 , y17033 , y17034 , y17035 , y17036 , y17037 , y17038 , y17039 , y17040 , y17041 , y17042 , y17043 , y17044 , y17045 , y17046 , y17047 , y17048 , y17049 , y17050 , y17051 , y17052 , y17053 , y17054 , y17055 , y17056 , y17057 , y17058 , y17059 , y17060 , y17061 , y17062 , y17063 , y17064 , y17065 , y17066 , y17067 , y17068 , y17069 , y17070 , y17071 , y17072 , y17073 , y17074 , y17075 , y17076 , y17077 , y17078 , y17079 , y17080 , y17081 , y17082 , y17083 , y17084 , y17085 , y17086 , y17087 , y17088 , y17089 , y17090 , y17091 , y17092 , y17093 , y17094 , y17095 , y17096 , y17097 , y17098 , y17099 , y17100 , y17101 , y17102 , y17103 , y17104 , y17105 , y17106 , y17107 , y17108 , y17109 , y17110 , y17111 , y17112 , y17113 , y17114 , y17115 , y17116 , y17117 , y17118 , y17119 , y17120 , y17121 , y17122 , y17123 , y17124 , y17125 , y17126 , y17127 , y17128 , y17129 , y17130 , y17131 , y17132 , y17133 , y17134 , y17135 , y17136 , y17137 , y17138 , y17139 , y17140 , y17141 , y17142 , y17143 , y17144 , y17145 , y17146 , y17147 , y17148 , y17149 , y17150 , y17151 , y17152 , y17153 , y17154 , y17155 , y17156 , y17157 , y17158 , y17159 , y17160 , y17161 , y17162 , y17163 , y17164 , y17165 , y17166 , y17167 , y17168 , y17169 , y17170 , y17171 , y17172 , y17173 , y17174 , y17175 , y17176 , y17177 , y17178 , y17179 , y17180 , y17181 , y17182 , y17183 , y17184 , y17185 , y17186 , y17187 , y17188 , y17189 , y17190 , y17191 , y17192 , y17193 , y17194 , y17195 , y17196 , y17197 , y17198 , y17199 , y17200 , y17201 , y17202 , y17203 , y17204 , y17205 , y17206 , y17207 , y17208 , y17209 , y17210 , y17211 , y17212 , y17213 , y17214 , y17215 , y17216 , y17217 , y17218 , y17219 , y17220 , y17221 , y17222 , y17223 , y17224 , y17225 , y17226 , y17227 , y17228 , y17229 , y17230 , y17231 , y17232 , y17233 , y17234 , y17235 , y17236 , y17237 , y17238 , y17239 , y17240 , y17241 , y17242 , y17243 , y17244 , y17245 , y17246 , y17247 , y17248 , y17249 , y17250 , y17251 , y17252 , y17253 , y17254 , y17255 , y17256 , y17257 , y17258 , y17259 , y17260 , y17261 , y17262 , y17263 , y17264 , y17265 , y17266 , y17267 , y17268 , y17269 , y17270 , y17271 , y17272 , y17273 , y17274 , y17275 , y17276 , y17277 , y17278 , y17279 , y17280 , y17281 , y17282 , y17283 , y17284 , y17285 , y17286 , y17287 , y17288 , y17289 , y17290 , y17291 , y17292 , y17293 , y17294 , y17295 , y17296 , y17297 , y17298 , y17299 , y17300 , y17301 , y17302 , y17303 , y17304 , y17305 , y17306 , y17307 , y17308 , y17309 , y17310 , y17311 , y17312 , y17313 , y17314 , y17315 , y17316 , y17317 , y17318 , y17319 , y17320 , y17321 , y17322 , y17323 , y17324 , y17325 , y17326 , y17327 , y17328 , y17329 , y17330 , y17331 , y17332 , y17333 , y17334 , y17335 , y17336 , y17337 , y17338 , y17339 , y17340 , y17341 , y17342 , y17343 , y17344 , y17345 , y17346 , y17347 , y17348 , y17349 , y17350 , y17351 , y17352 , y17353 , y17354 , y17355 , y17356 , y17357 , y17358 , y17359 , y17360 , y17361 , y17362 , y17363 , y17364 , y17365 , y17366 , y17367 , y17368 , y17369 , y17370 , y17371 , y17372 , y17373 , y17374 , y17375 , y17376 , y17377 , y17378 , y17379 , y17380 , y17381 , y17382 , y17383 , y17384 , y17385 , y17386 , y17387 , y17388 , y17389 , y17390 , y17391 , y17392 , y17393 , y17394 , y17395 , y17396 , y17397 , y17398 , y17399 , y17400 , y17401 , y17402 , y17403 , y17404 , y17405 , y17406 , y17407 , y17408 , y17409 , y17410 , y17411 , y17412 , y17413 , y17414 , y17415 , y17416 , y17417 , y17418 , y17419 , y17420 , y17421 , y17422 , y17423 , y17424 , y17425 , y17426 , y17427 , y17428 , y17429 , y17430 , y17431 , y17432 , y17433 , y17434 , y17435 , y17436 , y17437 , y17438 , y17439 , y17440 , y17441 , y17442 , y17443 , y17444 , y17445 , y17446 , y17447 , y17448 , y17449 , y17450 , y17451 , y17452 , y17453 , y17454 , y17455 , y17456 , y17457 , y17458 , y17459 , y17460 , y17461 , y17462 , y17463 , y17464 , y17465 , y17466 , y17467 , y17468 , y17469 , y17470 , y17471 , y17472 , y17473 , y17474 , y17475 , y17476 , y17477 , y17478 , y17479 , y17480 , y17481 , y17482 , y17483 , y17484 , y17485 , y17486 , y17487 , y17488 , y17489 , y17490 , y17491 , y17492 , y17493 , y17494 , y17495 , y17496 , y17497 , y17498 , y17499 , y17500 , y17501 , y17502 , y17503 , y17504 , y17505 , y17506 , y17507 , y17508 , y17509 , y17510 , y17511 , y17512 , y17513 , y17514 , y17515 , y17516 , y17517 , y17518 , y17519 , y17520 , y17521 , y17522 , y17523 , y17524 , y17525 , y17526 , y17527 , y17528 , y17529 , y17530 , y17531 , y17532 , y17533 , y17534 , y17535 , y17536 , y17537 , y17538 , y17539 , y17540 , y17541 , y17542 , y17543 , y17544 , y17545 , y17546 , y17547 , y17548 , y17549 , y17550 , y17551 , y17552 , y17553 , y17554 , y17555 , y17556 , y17557 , y17558 , y17559 , y17560 , y17561 , y17562 , y17563 , y17564 , y17565 , y17566 , y17567 , y17568 , y17569 , y17570 , y17571 , y17572 , y17573 , y17574 , y17575 , y17576 , y17577 , y17578 , y17579 , y17580 , y17581 , y17582 , y17583 , y17584 , y17585 , y17586 , y17587 , y17588 , y17589 , y17590 , y17591 , y17592 , y17593 , y17594 , y17595 , y17596 , y17597 , y17598 , y17599 , y17600 , y17601 , y17602 , y17603 , y17604 , y17605 , y17606 , y17607 , y17608 , y17609 , y17610 , y17611 , y17612 , y17613 , y17614 , y17615 , y17616 , y17617 , y17618 , y17619 , y17620 , y17621 , y17622 , y17623 , y17624 , y17625 , y17626 , y17627 , y17628 , y17629 , y17630 , y17631 , y17632 , y17633 , y17634 , y17635 , y17636 , y17637 , y17638 , y17639 , y17640 , y17641 , y17642 , y17643 , y17644 , y17645 , y17646 , y17647 , y17648 , y17649 , y17650 , y17651 , y17652 , y17653 , y17654 , y17655 , y17656 , y17657 , y17658 , y17659 , y17660 , y17661 , y17662 , y17663 , y17664 , y17665 , y17666 , y17667 , y17668 , y17669 , y17670 , y17671 , y17672 , y17673 , y17674 , y17675 , y17676 , y17677 , y17678 , y17679 , y17680 , y17681 , y17682 , y17683 , y17684 , y17685 , y17686 , y17687 , y17688 , y17689 , y17690 , y17691 , y17692 , y17693 , y17694 , y17695 , y17696 , y17697 , y17698 , y17699 , y17700 , y17701 , y17702 , y17703 , y17704 , y17705 , y17706 , y17707 , y17708 , y17709 , y17710 , y17711 , y17712 , y17713 , y17714 , y17715 , y17716 , y17717 , y17718 , y17719 , y17720 , y17721 , y17722 , y17723 , y17724 , y17725 , y17726 , y17727 , y17728 , y17729 , y17730 , y17731 , y17732 , y17733 , y17734 , y17735 , y17736 , y17737 , y17738 , y17739 , y17740 , y17741 , y17742 , y17743 , y17744 , y17745 , y17746 , y17747 , y17748 , y17749 , y17750 , y17751 , y17752 , y17753 , y17754 , y17755 , y17756 , y17757 , y17758 , y17759 , y17760 , y17761 , y17762 , y17763 , y17764 , y17765 , y17766 , y17767 , y17768 , y17769 , y17770 , y17771 , y17772 , y17773 , y17774 , y17775 , y17776 , y17777 , y17778 , y17779 , y17780 , y17781 , y17782 , y17783 , y17784 , y17785 , y17786 , y17787 , y17788 , y17789 , y17790 , y17791 , y17792 , y17793 , y17794 , y17795 , y17796 , y17797 , y17798 , y17799 , y17800 , y17801 , y17802 , y17803 , y17804 , y17805 , y17806 , y17807 , y17808 , y17809 , y17810 , y17811 , y17812 , y17813 , y17814 , y17815 , y17816 , y17817 , y17818 , y17819 , y17820 , y17821 , y17822 , y17823 , y17824 , y17825 , y17826 , y17827 , y17828 , y17829 , y17830 , y17831 , y17832 , y17833 , y17834 , y17835 , y17836 , y17837 , y17838 , y17839 , y17840 , y17841 , y17842 , y17843 , y17844 , y17845 , y17846 , y17847 , y17848 , y17849 , y17850 , y17851 , y17852 , y17853 , y17854 , y17855 , y17856 , y17857 , y17858 , y17859 , y17860 , y17861 , y17862 , y17863 , y17864 , y17865 , y17866 , y17867 , y17868 , y17869 , y17870 , y17871 , y17872 , y17873 , y17874 , y17875 , y17876 , y17877 , y17878 , y17879 , y17880 , y17881 , y17882 , y17883 , y17884 , y17885 , y17886 , y17887 , y17888 , y17889 , y17890 , y17891 , y17892 , y17893 , y17894 , y17895 , y17896 , y17897 , y17898 , y17899 , y17900 , y17901 , y17902 , y17903 , y17904 , y17905 , y17906 , y17907 , y17908 , y17909 , y17910 , y17911 , y17912 , y17913 , y17914 , y17915 , y17916 , y17917 , y17918 , y17919 , y17920 , y17921 , y17922 , y17923 , y17924 , y17925 , y17926 , y17927 , y17928 , y17929 , y17930 , y17931 , y17932 , y17933 , y17934 , y17935 , y17936 , y17937 , y17938 , y17939 , y17940 , y17941 , y17942 , y17943 , y17944 , y17945 , y17946 , y17947 , y17948 , y17949 , y17950 , y17951 , y17952 , y17953 , y17954 , y17955 , y17956 , y17957 , y17958 , y17959 , y17960 , y17961 , y17962 , y17963 , y17964 , y17965 , y17966 , y17967 , y17968 , y17969 , y17970 , y17971 , y17972 , y17973 , y17974 , y17975 , y17976 , y17977 , y17978 , y17979 , y17980 , y17981 , y17982 , y17983 , y17984 , y17985 , y17986 , y17987 , y17988 , y17989 , y17990 , y17991 , y17992 , y17993 , y17994 , y17995 , y17996 , y17997 , y17998 , y17999 , y18000 , y18001 , y18002 , y18003 , y18004 , y18005 , y18006 , y18007 , y18008 , y18009 , y18010 , y18011 , y18012 , y18013 , y18014 , y18015 , y18016 , y18017 , y18018 , y18019 , y18020 , y18021 , y18022 , y18023 , y18024 , y18025 , y18026 , y18027 , y18028 , y18029 , y18030 , y18031 , y18032 , y18033 , y18034 , y18035 , y18036 , y18037 , y18038 , y18039 , y18040 , y18041 , y18042 , y18043 , y18044 , y18045 , y18046 , y18047 , y18048 , y18049 , y18050 , y18051 , y18052 , y18053 , y18054 , y18055 , y18056 , y18057 , y18058 , y18059 , y18060 , y18061 , y18062 , y18063 , y18064 , y18065 , y18066 , y18067 , y18068 , y18069 , y18070 , y18071 , y18072 , y18073 , y18074 , y18075 , y18076 , y18077 , y18078 , y18079 , y18080 , y18081 , y18082 , y18083 , y18084 , y18085 , y18086 , y18087 , y18088 , y18089 , y18090 , y18091 , y18092 , y18093 , y18094 , y18095 , y18096 , y18097 , y18098 , y18099 , y18100 , y18101 , y18102 , y18103 , y18104 , y18105 , y18106 , y18107 , y18108 , y18109 , y18110 , y18111 , y18112 , y18113 , y18114 , y18115 , y18116 , y18117 , y18118 , y18119 , y18120 , y18121 , y18122 , y18123 , y18124 , y18125 , y18126 , y18127 , y18128 , y18129 , y18130 , y18131 , y18132 , y18133 , y18134 , y18135 , y18136 , y18137 , y18138 , y18139 , y18140 , y18141 , y18142 , y18143 , y18144 , y18145 , y18146 , y18147 , y18148 , y18149 , y18150 , y18151 , y18152 , y18153 , y18154 , y18155 , y18156 , y18157 , y18158 , y18159 , y18160 , y18161 , y18162 , y18163 , y18164 , y18165 , y18166 , y18167 , y18168 , y18169 , y18170 , y18171 , y18172 , y18173 , y18174 , y18175 , y18176 , y18177 , y18178 , y18179 , y18180 , y18181 , y18182 , y18183 , y18184 , y18185 , y18186 , y18187 , y18188 , y18189 , y18190 , y18191 , y18192 , y18193 , y18194 , y18195 , y18196 , y18197 , y18198 , y18199 , y18200 , y18201 , y18202 , y18203 , y18204 , y18205 , y18206 , y18207 , y18208 , y18209 , y18210 , y18211 , y18212 , y18213 , y18214 , y18215 , y18216 , y18217 , y18218 , y18219 , y18220 , y18221 , y18222 , y18223 , y18224 , y18225 , y18226 , y18227 , y18228 , y18229 , y18230 , y18231 , y18232 , y18233 , y18234 , y18235 , y18236 , y18237 , y18238 , y18239 , y18240 , y18241 , y18242 , y18243 , y18244 , y18245 , y18246 , y18247 , y18248 , y18249 , y18250 , y18251 , y18252 , y18253 , y18254 , y18255 , y18256 , y18257 , y18258 , y18259 , y18260 , y18261 , y18262 , y18263 , y18264 , y18265 , y18266 , y18267 , y18268 , y18269 , y18270 , y18271 , y18272 , y18273 , y18274 , y18275 , y18276 , y18277 , y18278 , y18279 , y18280 , y18281 , y18282 , y18283 , y18284 , y18285 , y18286 , y18287 , y18288 , y18289 , y18290 , y18291 , y18292 , y18293 , y18294 , y18295 , y18296 , y18297 , y18298 , y18299 , y18300 , y18301 , y18302 , y18303 , y18304 , y18305 , y18306 , y18307 , y18308 , y18309 , y18310 , y18311 , y18312 , y18313 , y18314 , y18315 , y18316 , y18317 , y18318 , y18319 , y18320 , y18321 , y18322 , y18323 , y18324 , y18325 , y18326 , y18327 , y18328 , y18329 , y18330 , y18331 , y18332 , y18333 , y18334 , y18335 , y18336 , y18337 , y18338 , y18339 , y18340 , y18341 , y18342 , y18343 , y18344 , y18345 , y18346 , y18347 , y18348 , y18349 , y18350 , y18351 , y18352 , y18353 , y18354 , y18355 , y18356 , y18357 , y18358 , y18359 , y18360 , y18361 , y18362 , y18363 , y18364 , y18365 , y18366 , y18367 , y18368 , y18369 , y18370 , y18371 , y18372 , y18373 , y18374 , y18375 , y18376 , y18377 , y18378 , y18379 , y18380 , y18381 , y18382 , y18383 , y18384 , y18385 , y18386 , y18387 , y18388 , y18389 , y18390 , y18391 , y18392 , y18393 , y18394 , y18395 , y18396 , y18397 , y18398 , y18399 , y18400 , y18401 , y18402 , y18403 , y18404 , y18405 , y18406 , y18407 , y18408 , y18409 , y18410 , y18411 , y18412 , y18413 , y18414 , y18415 , y18416 , y18417 , y18418 , y18419 , y18420 , y18421 , y18422 , y18423 , y18424 , y18425 , y18426 , y18427 , y18428 , y18429 , y18430 , y18431 , y18432 , y18433 , y18434 , y18435 , y18436 , y18437 , y18438 , y18439 , y18440 , y18441 , y18442 , y18443 , y18444 , y18445 , y18446 , y18447 , y18448 , y18449 , y18450 , y18451 , y18452 , y18453 , y18454 , y18455 , y18456 , y18457 , y18458 , y18459 , y18460 , y18461 , y18462 , y18463 , y18464 , y18465 , y18466 , y18467 , y18468 , y18469 , y18470 , y18471 , y18472 , y18473 , y18474 , y18475 , y18476 , y18477 , y18478 , y18479 , y18480 , y18481 , y18482 , y18483 , y18484 , y18485 , y18486 , y18487 , y18488 , y18489 , y18490 , y18491 , y18492 , y18493 , y18494 , y18495 , y18496 , y18497 , y18498 , y18499 , y18500 , y18501 , y18502 , y18503 , y18504 , y18505 , y18506 , y18507 , y18508 , y18509 , y18510 , y18511 , y18512 , y18513 , y18514 , y18515 , y18516 , y18517 , y18518 , y18519 , y18520 , y18521 , y18522 , y18523 , y18524 , y18525 , y18526 , y18527 , y18528 , y18529 , y18530 , y18531 , y18532 , y18533 , y18534 , y18535 , y18536 , y18537 , y18538 , y18539 , y18540 , y18541 , y18542 , y18543 , y18544 , y18545 , y18546 , y18547 , y18548 , y18549 , y18550 , y18551 , y18552 , y18553 , y18554 , y18555 , y18556 , y18557 , y18558 , y18559 , y18560 , y18561 , y18562 , y18563 , y18564 , y18565 , y18566 , y18567 , y18568 , y18569 , y18570 , y18571 , y18572 , y18573 , y18574 , y18575 , y18576 , y18577 , y18578 , y18579 , y18580 , y18581 , y18582 , y18583 , y18584 , y18585 , y18586 , y18587 , y18588 , y18589 , y18590 , y18591 , y18592 , y18593 , y18594 , y18595 , y18596 , y18597 , y18598 , y18599 , y18600 , y18601 , y18602 , y18603 , y18604 , y18605 , y18606 , y18607 , y18608 , y18609 , y18610 , y18611 , y18612 , y18613 , y18614 , y18615 , y18616 , y18617 , y18618 , y18619 , y18620 , y18621 , y18622 , y18623 , y18624 , y18625 , y18626 , y18627 , y18628 , y18629 , y18630 , y18631 , y18632 , y18633 , y18634 , y18635 , y18636 , y18637 , y18638 , y18639 , y18640 , y18641 , y18642 , y18643 , y18644 , y18645 , y18646 , y18647 , y18648 , y18649 , y18650 , y18651 , y18652 , y18653 , y18654 , y18655 , y18656 , y18657 , y18658 , y18659 , y18660 , y18661 , y18662 , y18663 , y18664 , y18665 , y18666 , y18667 , y18668 , y18669 , y18670 , y18671 , y18672 , y18673 , y18674 , y18675 , y18676 , y18677 , y18678 , y18679 , y18680 , y18681 , y18682 , y18683 , y18684 , y18685 , y18686 , y18687 , y18688 , y18689 , y18690 , y18691 , y18692 , y18693 , y18694 , y18695 , y18696 , y18697 , y18698 , y18699 , y18700 , y18701 , y18702 , y18703 , y18704 , y18705 , y18706 , y18707 , y18708 , y18709 , y18710 , y18711 , y18712 , y18713 , y18714 , y18715 , y18716 , y18717 , y18718 , y18719 , y18720 , y18721 , y18722 , y18723 , y18724 , y18725 , y18726 , y18727 , y18728 , y18729 , y18730 , y18731 , y18732 , y18733 , y18734 , y18735 , y18736 , y18737 , y18738 , y18739 , y18740 , y18741 , y18742 , y18743 , y18744 , y18745 , y18746 , y18747 , y18748 , y18749 , y18750 , y18751 , y18752 , y18753 , y18754 , y18755 , y18756 , y18757 , y18758 , y18759 , y18760 , y18761 , y18762 , y18763 , y18764 , y18765 , y18766 , y18767 , y18768 , y18769 , y18770 , y18771 , y18772 , y18773 , y18774 , y18775 , y18776 , y18777 , y18778 , y18779 , y18780 , y18781 , y18782 , y18783 , y18784 , y18785 , y18786 , y18787 , y18788 , y18789 , y18790 , y18791 , y18792 , y18793 , y18794 , y18795 , y18796 , y18797 , y18798 , y18799 , y18800 , y18801 , y18802 , y18803 , y18804 , y18805 , y18806 , y18807 , y18808 , y18809 , y18810 , y18811 , y18812 , y18813 , y18814 , y18815 , y18816 , y18817 , y18818 , y18819 , y18820 , y18821 , y18822 , y18823 , y18824 , y18825 , y18826 , y18827 , y18828 , y18829 , y18830 , y18831 , y18832 , y18833 , y18834 , y18835 , y18836 , y18837 , y18838 , y18839 , y18840 , y18841 , y18842 , y18843 , y18844 , y18845 , y18846 , y18847 , y18848 , y18849 , y18850 , y18851 , y18852 , y18853 , y18854 , y18855 , y18856 , y18857 , y18858 , y18859 , y18860 , y18861 , y18862 , y18863 , y18864 , y18865 , y18866 , y18867 , y18868 , y18869 , y18870 , y18871 , y18872 , y18873 , y18874 , y18875 , y18876 , y18877 , y18878 , y18879 , y18880 , y18881 , y18882 , y18883 , y18884 , y18885 , y18886 , y18887 , y18888 , y18889 , y18890 , y18891 , y18892 , y18893 , y18894 , y18895 , y18896 , y18897 , y18898 , y18899 , y18900 , y18901 , y18902 , y18903 , y18904 , y18905 , y18906 , y18907 , y18908 , y18909 , y18910 , y18911 , y18912 , y18913 , y18914 , y18915 , y18916 , y18917 , y18918 , y18919 , y18920 , y18921 , y18922 , y18923 , y18924 , y18925 , y18926 , y18927 , y18928 , y18929 , y18930 , y18931 , y18932 , y18933 , y18934 , y18935 , y18936 , y18937 , y18938 , y18939 , y18940 , y18941 , y18942 , y18943 , y18944 , y18945 , y18946 , y18947 , y18948 , y18949 , y18950 , y18951 , y18952 , y18953 , y18954 , y18955 , y18956 , y18957 , y18958 , y18959 , y18960 , y18961 , y18962 , y18963 , y18964 , y18965 , y18966 , y18967 , y18968 , y18969 , y18970 , y18971 , y18972 , y18973 , y18974 , y18975 , y18976 , y18977 , y18978 , y18979 , y18980 , y18981 , y18982 , y18983 , y18984 , y18985 , y18986 , y18987 , y18988 , y18989 , y18990 , y18991 , y18992 , y18993 , y18994 , y18995 , y18996 , y18997 , y18998 , y18999 , y19000 , y19001 , y19002 , y19003 , y19004 , y19005 , y19006 , y19007 , y19008 , y19009 , y19010 , y19011 , y19012 , y19013 , y19014 , y19015 , y19016 , y19017 , y19018 , y19019 , y19020 , y19021 , y19022 , y19023 , y19024 , y19025 , y19026 , y19027 , y19028 , y19029 , y19030 , y19031 , y19032 , y19033 , y19034 , y19035 , y19036 , y19037 , y19038 , y19039 , y19040 , y19041 , y19042 , y19043 , y19044 , y19045 , y19046 , y19047 , y19048 , y19049 , y19050 , y19051 , y19052 , y19053 , y19054 , y19055 , y19056 , y19057 , y19058 , y19059 , y19060 , y19061 , y19062 , y19063 , y19064 , y19065 , y19066 , y19067 , y19068 , y19069 , y19070 , y19071 , y19072 , y19073 , y19074 , y19075 , y19076 , y19077 , y19078 , y19079 , y19080 , y19081 , y19082 , y19083 , y19084 , y19085 , y19086 , y19087 , y19088 , y19089 , y19090 , y19091 , y19092 , y19093 , y19094 , y19095 , y19096 , y19097 , y19098 , y19099 , y19100 , y19101 , y19102 , y19103 , y19104 , y19105 , y19106 , y19107 , y19108 , y19109 , y19110 , y19111 , y19112 , y19113 , y19114 , y19115 , y19116 , y19117 , y19118 , y19119 , y19120 , y19121 , y19122 , y19123 , y19124 , y19125 , y19126 , y19127 , y19128 , y19129 , y19130 , y19131 , y19132 , y19133 , y19134 , y19135 , y19136 , y19137 , y19138 , y19139 , y19140 , y19141 , y19142 , y19143 , y19144 , y19145 , y19146 , y19147 , y19148 , y19149 , y19150 , y19151 , y19152 , y19153 , y19154 , y19155 , y19156 , y19157 , y19158 , y19159 , y19160 , y19161 , y19162 , y19163 , y19164 , y19165 , y19166 , y19167 , y19168 , y19169 , y19170 , y19171 , y19172 , y19173 , y19174 , y19175 , y19176 , y19177 , y19178 , y19179 , y19180 , y19181 , y19182 , y19183 , y19184 , y19185 , y19186 , y19187 , y19188 , y19189 , y19190 , y19191 , y19192 , y19193 , y19194 , y19195 , y19196 , y19197 , y19198 , y19199 , y19200 , y19201 , y19202 , y19203 , y19204 , y19205 , y19206 , y19207 , y19208 , y19209 , y19210 , y19211 , y19212 , y19213 , y19214 , y19215 , y19216 , y19217 , y19218 , y19219 , y19220 , y19221 , y19222 , y19223 , y19224 , y19225 , y19226 , y19227 , y19228 , y19229 , y19230 , y19231 , y19232 , y19233 , y19234 , y19235 , y19236 , y19237 , y19238 , y19239 , y19240 , y19241 , y19242 , y19243 , y19244 , y19245 , y19246 , y19247 , y19248 , y19249 , y19250 , y19251 , y19252 , y19253 , y19254 , y19255 , y19256 , y19257 , y19258 , y19259 , y19260 , y19261 , y19262 , y19263 , y19264 , y19265 , y19266 , y19267 , y19268 , y19269 , y19270 , y19271 , y19272 , y19273 , y19274 , y19275 , y19276 , y19277 , y19278 , y19279 , y19280 , y19281 , y19282 , y19283 , y19284 , y19285 , y19286 , y19287 , y19288 , y19289 , y19290 , y19291 , y19292 , y19293 , y19294 , y19295 , y19296 , y19297 , y19298 , y19299 , y19300 , y19301 , y19302 , y19303 , y19304 , y19305 , y19306 , y19307 , y19308 , y19309 , y19310 , y19311 , y19312 , y19313 , y19314 , y19315 , y19316 , y19317 , y19318 , y19319 , y19320 , y19321 , y19322 , y19323 , y19324 , y19325 , y19326 , y19327 , y19328 , y19329 , y19330 , y19331 , y19332 , y19333 , y19334 , y19335 , y19336 , y19337 , y19338 , y19339 , y19340 , y19341 , y19342 , y19343 , y19344 , y19345 , y19346 , y19347 , y19348 , y19349 , y19350 , y19351 , y19352 , y19353 , y19354 , y19355 , y19356 , y19357 , y19358 , y19359 , y19360 , y19361 , y19362 , y19363 , y19364 , y19365 , y19366 , y19367 , y19368 , y19369 , y19370 , y19371 , y19372 , y19373 , y19374 , y19375 , y19376 , y19377 , y19378 , y19379 , y19380 , y19381 , y19382 , y19383 , y19384 , y19385 , y19386 , y19387 , y19388 , y19389 , y19390 , y19391 , y19392 , y19393 , y19394 , y19395 , y19396 , y19397 , y19398 , y19399 , y19400 , y19401 , y19402 , y19403 , y19404 , y19405 , y19406 , y19407 , y19408 , y19409 , y19410 , y19411 , y19412 , y19413 , y19414 , y19415 , y19416 , y19417 , y19418 , y19419 , y19420 , y19421 , y19422 , y19423 , y19424 , y19425 , y19426 , y19427 , y19428 , y19429 , y19430 , y19431 , y19432 , y19433 , y19434 , y19435 , y19436 , y19437 , y19438 , y19439 , y19440 , y19441 , y19442 , y19443 , y19444 , y19445 , y19446 , y19447 , y19448 , y19449 , y19450 , y19451 , y19452 , y19453 , y19454 , y19455 , y19456 , y19457 , y19458 , y19459 , y19460 , y19461 , y19462 , y19463 , y19464 , y19465 , y19466 , y19467 , y19468 , y19469 , y19470 , y19471 , y19472 , y19473 , y19474 , y19475 , y19476 , y19477 , y19478 , y19479 , y19480 , y19481 , y19482 , y19483 , y19484 , y19485 , y19486 , y19487 , y19488 , y19489 , y19490 , y19491 , y19492 , y19493 , y19494 , y19495 , y19496 , y19497 , y19498 , y19499 , y19500 , y19501 , y19502 , y19503 , y19504 , y19505 , y19506 , y19507 , y19508 , y19509 , y19510 , y19511 , y19512 , y19513 , y19514 , y19515 , y19516 , y19517 , y19518 , y19519 , y19520 , y19521 , y19522 , y19523 , y19524 , y19525 , y19526 , y19527 , y19528 , y19529 , y19530 , y19531 , y19532 , y19533 , y19534 , y19535 , y19536 , y19537 , y19538 , y19539 , y19540 , y19541 , y19542 , y19543 , y19544 , y19545 , y19546 , y19547 , y19548 , y19549 , y19550 , y19551 , y19552 , y19553 , y19554 , y19555 , y19556 , y19557 , y19558 , y19559 , y19560 , y19561 , y19562 , y19563 , y19564 , y19565 , y19566 , y19567 , y19568 , y19569 , y19570 , y19571 , y19572 , y19573 , y19574 , y19575 , y19576 , y19577 , y19578 , y19579 , y19580 , y19581 , y19582 , y19583 , y19584 , y19585 , y19586 , y19587 , y19588 , y19589 , y19590 , y19591 , y19592 , y19593 , y19594 , y19595 , y19596 , y19597 , y19598 , y19599 , y19600 , y19601 , y19602 , y19603 , y19604 , y19605 , y19606 , y19607 , y19608 , y19609 , y19610 , y19611 , y19612 , y19613 , y19614 , y19615 , y19616 , y19617 , y19618 , y19619 , y19620 , y19621 , y19622 , y19623 , y19624 , y19625 , y19626 , y19627 , y19628 , y19629 , y19630 , y19631 , y19632 , y19633 , y19634 , y19635 , y19636 , y19637 , y19638 , y19639 , y19640 , y19641 , y19642 , y19643 , y19644 , y19645 , y19646 , y19647 , y19648 , y19649 , y19650 , y19651 , y19652 , y19653 , y19654 , y19655 , y19656 , y19657 , y19658 , y19659 , y19660 , y19661 , y19662 , y19663 , y19664 , y19665 , y19666 , y19667 , y19668 , y19669 , y19670 , y19671 , y19672 , y19673 , y19674 , y19675 , y19676 , y19677 , y19678 , y19679 , y19680 , y19681 , y19682 , y19683 , y19684 , y19685 , y19686 , y19687 , y19688 , y19689 , y19690 , y19691 , y19692 , y19693 , y19694 , y19695 , y19696 , y19697 , y19698 , y19699 , y19700 , y19701 , y19702 , y19703 , y19704 , y19705 , y19706 , y19707 , y19708 , y19709 , y19710 , y19711 , y19712 , y19713 , y19714 , y19715 , y19716 , y19717 , y19718 , y19719 , y19720 , y19721 , y19722 , y19723 , y19724 , y19725 , y19726 , y19727 , y19728 , y19729 , y19730 , y19731 , y19732 , y19733 , y19734 , y19735 , y19736 , y19737 , y19738 , y19739 , y19740 , y19741 , y19742 , y19743 , y19744 , y19745 , y19746 , y19747 , y19748 , y19749 , y19750 , y19751 , y19752 , y19753 , y19754 , y19755 , y19756 , y19757 , y19758 , y19759 , y19760 , y19761 , y19762 , y19763 , y19764 , y19765 , y19766 , y19767 , y19768 , y19769 , y19770 , y19771 , y19772 , y19773 , y19774 , y19775 , y19776 , y19777 , y19778 , y19779 , y19780 , y19781 , y19782 , y19783 , y19784 , y19785 , y19786 , y19787 , y19788 , y19789 , y19790 , y19791 , y19792 , y19793 , y19794 , y19795 , y19796 , y19797 , y19798 , y19799 , y19800 , y19801 , y19802 , y19803 , y19804 , y19805 , y19806 , y19807 , y19808 , y19809 , y19810 , y19811 , y19812 , y19813 , y19814 , y19815 , y19816 , y19817 , y19818 , y19819 , y19820 , y19821 , y19822 , y19823 , y19824 , y19825 , y19826 , y19827 , y19828 , y19829 , y19830 , y19831 , y19832 , y19833 , y19834 , y19835 , y19836 , y19837 , y19838 , y19839 , y19840 , y19841 , y19842 , y19843 , y19844 , y19845 , y19846 , y19847 , y19848 , y19849 , y19850 , y19851 , y19852 , y19853 , y19854 , y19855 , y19856 , y19857 , y19858 , y19859 , y19860 , y19861 , y19862 , y19863 , y19864 , y19865 , y19866 , y19867 , y19868 , y19869 , y19870 , y19871 , y19872 , y19873 , y19874 , y19875 , y19876 , y19877 , y19878 , y19879 , y19880 , y19881 , y19882 , y19883 , y19884 , y19885 , y19886 , y19887 , y19888 , y19889 , y19890 , y19891 , y19892 , y19893 , y19894 , y19895 , y19896 , y19897 , y19898 , y19899 , y19900 , y19901 , y19902 , y19903 , y19904 , y19905 , y19906 , y19907 , y19908 , y19909 , y19910 , y19911 , y19912 , y19913 , y19914 , y19915 , y19916 , y19917 , y19918 , y19919 , y19920 , y19921 , y19922 , y19923 , y19924 , y19925 , y19926 , y19927 , y19928 , y19929 , y19930 , y19931 , y19932 , y19933 , y19934 , y19935 , y19936 , y19937 , y19938 , y19939 , y19940 , y19941 , y19942 , y19943 , y19944 , y19945 , y19946 , y19947 , y19948 , y19949 , y19950 , y19951 , y19952 , y19953 , y19954 , y19955 , y19956 , y19957 , y19958 , y19959 , y19960 , y19961 , y19962 , y19963 , y19964 , y19965 , y19966 , y19967 , y19968 , y19969 , y19970 , y19971 , y19972 , y19973 , y19974 , y19975 , y19976 , y19977 , y19978 , y19979 , y19980 , y19981 , y19982 , y19983 , y19984 , y19985 , y19986 , y19987 , y19988 , y19989 , y19990 , y19991 , y19992 , y19993 , y19994 , y19995 , y19996 , y19997 , y19998 , y19999 , y20000 , y20001 , y20002 , y20003 , y20004 , y20005 , y20006 , y20007 , y20008 , y20009 , y20010 , y20011 , y20012 , y20013 , y20014 , y20015 , y20016 , y20017 , y20018 , y20019 , y20020 , y20021 , y20022 , y20023 , y20024 , y20025 , y20026 , y20027 , y20028 , y20029 , y20030 , y20031 , y20032 , y20033 , y20034 , y20035 , y20036 , y20037 , y20038 , y20039 , y20040 , y20041 , y20042 , y20043 , y20044 , y20045 , y20046 , y20047 , y20048 , y20049 , y20050 , y20051 , y20052 , y20053 , y20054 , y20055 , y20056 , y20057 , y20058 , y20059 , y20060 , y20061 , y20062 , y20063 , y20064 , y20065 , y20066 , y20067 , y20068 , y20069 , y20070 , y20071 , y20072 , y20073 , y20074 , y20075 , y20076 , y20077 , y20078 , y20079 , y20080 , y20081 , y20082 , y20083 , y20084 , y20085 , y20086 , y20087 , y20088 , y20089 , y20090 , y20091 , y20092 , y20093 , y20094 , y20095 , y20096 , y20097 , y20098 , y20099 , y20100 , y20101 , y20102 , y20103 , y20104 , y20105 , y20106 , y20107 , y20108 , y20109 , y20110 , y20111 , y20112 , y20113 , y20114 , y20115 , y20116 , y20117 , y20118 , y20119 , y20120 , y20121 , y20122 , y20123 , y20124 , y20125 , y20126 , y20127 , y20128 , y20129 , y20130 , y20131 , y20132 , y20133 , y20134 , y20135 , y20136 , y20137 , y20138 , y20139 , y20140 , y20141 , y20142 , y20143 , y20144 , y20145 , y20146 , y20147 , y20148 , y20149 , y20150 , y20151 , y20152 , y20153 , y20154 , y20155 , y20156 , y20157 , y20158 , y20159 , y20160 , y20161 , y20162 , y20163 , y20164 , y20165 , y20166 , y20167 , y20168 , y20169 , y20170 , y20171 , y20172 , y20173 , y20174 , y20175 , y20176 , y20177 , y20178 , y20179 , y20180 , y20181 , y20182 , y20183 , y20184 , y20185 , y20186 , y20187 , y20188 , y20189 , y20190 , y20191 , y20192 , y20193 , y20194 , y20195 , y20196 , y20197 , y20198 , y20199 , y20200 , y20201 , y20202 , y20203 , y20204 , y20205 , y20206 , y20207 , y20208 , y20209 , y20210 , y20211 , y20212 , y20213 , y20214 , y20215 , y20216 , y20217 , y20218 , y20219 , y20220 , y20221 , y20222 , y20223 , y20224 , y20225 , y20226 , y20227 , y20228 , y20229 , y20230 , y20231 , y20232 , y20233 , y20234 , y20235 , y20236 , y20237 , y20238 , y20239 , y20240 , y20241 , y20242 , y20243 , y20244 , y20245 , y20246 , y20247 , y20248 , y20249 , y20250 , y20251 , y20252 , y20253 , y20254 , y20255 , y20256 , y20257 , y20258 , y20259 , y20260 , y20261 , y20262 , y20263 , y20264 , y20265 , y20266 , y20267 , y20268 , y20269 , y20270 , y20271 , y20272 , y20273 , y20274 , y20275 , y20276 , y20277 , y20278 , y20279 , y20280 , y20281 , y20282 , y20283 , y20284 , y20285 , y20286 , y20287 , y20288 , y20289 , y20290 , y20291 , y20292 , y20293 , y20294 , y20295 , y20296 , y20297 , y20298 , y20299 , y20300 , y20301 , y20302 , y20303 , y20304 , y20305 , y20306 , y20307 , y20308 , y20309 , y20310 , y20311 , y20312 , y20313 , y20314 , y20315 , y20316 , y20317 , y20318 , y20319 , y20320 , y20321 , y20322 , y20323 , y20324 , y20325 , y20326 , y20327 , y20328 , y20329 , y20330 , y20331 , y20332 , y20333 , y20334 , y20335 , y20336 , y20337 , y20338 , y20339 , y20340 , y20341 , y20342 , y20343 , y20344 , y20345 , y20346 , y20347 , y20348 , y20349 , y20350 , y20351 , y20352 , y20353 , y20354 , y20355 , y20356 , y20357 , y20358 , y20359 , y20360 , y20361 , y20362 , y20363 , y20364 , y20365 , y20366 , y20367 , y20368 , y20369 , y20370 , y20371 , y20372 , y20373 , y20374 , y20375 , y20376 , y20377 , y20378 , y20379 , y20380 , y20381 , y20382 , y20383 , y20384 , y20385 , y20386 , y20387 , y20388 , y20389 , y20390 , y20391 , y20392 , y20393 , y20394 , y20395 , y20396 , y20397 , y20398 , y20399 , y20400 , y20401 , y20402 , y20403 , y20404 , y20405 , y20406 , y20407 , y20408 , y20409 , y20410 , y20411 , y20412 , y20413 , y20414 , y20415 , y20416 , y20417 , y20418 , y20419 , y20420 , y20421 , y20422 , y20423 , y20424 , y20425 , y20426 , y20427 , y20428 , y20429 , y20430 , y20431 , y20432 , y20433 , y20434 , y20435 , y20436 , y20437 , y20438 , y20439 , y20440 , y20441 , y20442 , y20443 , y20444 , y20445 , y20446 , y20447 , y20448 , y20449 , y20450 , y20451 , y20452 , y20453 , y20454 , y20455 , y20456 , y20457 , y20458 , y20459 , y20460 , y20461 , y20462 , y20463 , y20464 , y20465 , y20466 , y20467 , y20468 , y20469 , y20470 , y20471 , y20472 , y20473 , y20474 , y20475 , y20476 , y20477 , y20478 , y20479 , y20480 , y20481 , y20482 , y20483 , y20484 , y20485 , y20486 , y20487 , y20488 , y20489 , y20490 , y20491 , y20492 , y20493 , y20494 , y20495 , y20496 , y20497 , y20498 , y20499 , y20500 , y20501 , y20502 , y20503 , y20504 , y20505 , y20506 , y20507 , y20508 , y20509 , y20510 , y20511 , y20512 , y20513 , y20514 , y20515 , y20516 , y20517 , y20518 , y20519 , y20520 , y20521 , y20522 , y20523 , y20524 , y20525 , y20526 , y20527 , y20528 , y20529 , y20530 , y20531 , y20532 , y20533 , y20534 , y20535 , y20536 , y20537 , y20538 , y20539 , y20540 , y20541 , y20542 , y20543 , y20544 , y20545 , y20546 , y20547 , y20548 , y20549 , y20550 , y20551 , y20552 , y20553 , y20554 , y20555 , y20556 , y20557 , y20558 , y20559 , y20560 , y20561 , y20562 , y20563 , y20564 , y20565 , y20566 , y20567 , y20568 , y20569 , y20570 , y20571 , y20572 , y20573 , y20574 , y20575 , y20576 , y20577 , y20578 , y20579 , y20580 , y20581 , y20582 , y20583 , y20584 , y20585 , y20586 , y20587 , y20588 , y20589 , y20590 , y20591 , y20592 , y20593 , y20594 , y20595 , y20596 , y20597 , y20598 , y20599 , y20600 , y20601 , y20602 , y20603 , y20604 , y20605 , y20606 , y20607 , y20608 , y20609 , y20610 , y20611 , y20612 , y20613 , y20614 , y20615 , y20616 , y20617 , y20618 , y20619 , y20620 , y20621 , y20622 , y20623 , y20624 , y20625 , y20626 , y20627 , y20628 , y20629 , y20630 , y20631 , y20632 , y20633 , y20634 , y20635 , y20636 , y20637 , y20638 , y20639 , y20640 , y20641 , y20642 , y20643 , y20644 , y20645 , y20646 , y20647 , y20648 , y20649 , y20650 , y20651 , y20652 , y20653 , y20654 , y20655 , y20656 , y20657 , y20658 , y20659 , y20660 , y20661 , y20662 , y20663 , y20664 , y20665 , y20666 , y20667 , y20668 , y20669 , y20670 , y20671 , y20672 , y20673 , y20674 , y20675 , y20676 , y20677 , y20678 , y20679 , y20680 , y20681 , y20682 , y20683 , y20684 , y20685 , y20686 , y20687 , y20688 , y20689 , y20690 , y20691 , y20692 , y20693 , y20694 , y20695 , y20696 , y20697 , y20698 , y20699 , y20700 , y20701 , y20702 , y20703 , y20704 , y20705 , y20706 , y20707 , y20708 , y20709 , y20710 , y20711 , y20712 , y20713 , y20714 , y20715 , y20716 , y20717 , y20718 , y20719 , y20720 , y20721 , y20722 , y20723 , y20724 , y20725 , y20726 , y20727 , y20728 , y20729 , y20730 , y20731 , y20732 , y20733 , y20734 , y20735 , y20736 , y20737 , y20738 , y20739 , y20740 , y20741 , y20742 , y20743 , y20744 , y20745 , y20746 , y20747 , y20748 , y20749 , y20750 , y20751 , y20752 , y20753 , y20754 , y20755 , y20756 , y20757 , y20758 , y20759 , y20760 , y20761 , y20762 , y20763 , y20764 , y20765 , y20766 , y20767 , y20768 , y20769 , y20770 , y20771 , y20772 , y20773 , y20774 , y20775 , y20776 , y20777 , y20778 , y20779 , y20780 , y20781 , y20782 , y20783 , y20784 , y20785 , y20786 , y20787 , y20788 , y20789 , y20790 , y20791 , y20792 , y20793 , y20794 , y20795 , y20796 , y20797 , y20798 , y20799 , y20800 , y20801 , y20802 , y20803 , y20804 , y20805 , y20806 , y20807 , y20808 , y20809 , y20810 , y20811 , y20812 , y20813 , y20814 , y20815 , y20816 , y20817 , y20818 , y20819 , y20820 , y20821 , y20822 , y20823 , y20824 , y20825 , y20826 , y20827 , y20828 , y20829 , y20830 , y20831 , y20832 , y20833 , y20834 , y20835 , y20836 , y20837 , y20838 , y20839 , y20840 , y20841 , y20842 , y20843 , y20844 , y20845 , y20846 , y20847 , y20848 , y20849 , y20850 , y20851 , y20852 , y20853 , y20854 , y20855 , y20856 , y20857 , y20858 , y20859 , y20860 , y20861 , y20862 , y20863 , y20864 , y20865 , y20866 , y20867 , y20868 , y20869 , y20870 , y20871 , y20872 , y20873 , y20874 , y20875 , y20876 , y20877 , y20878 , y20879 , y20880 , y20881 , y20882 , y20883 , y20884 , y20885 , y20886 , y20887 , y20888 , y20889 , y20890 , y20891 , y20892 , y20893 , y20894 , y20895 , y20896 , y20897 , y20898 , y20899 , y20900 , y20901 , y20902 , y20903 , y20904 , y20905 , y20906 , y20907 , y20908 , y20909 , y20910 , y20911 , y20912 , y20913 , y20914 , y20915 , y20916 , y20917 , y20918 , y20919 , y20920 , y20921 , y20922 , y20923 , y20924 , y20925 , y20926 , y20927 , y20928 , y20929 , y20930 , y20931 , y20932 , y20933 , y20934 , y20935 , y20936 , y20937 , y20938 , y20939 , y20940 , y20941 , y20942 , y20943 , y20944 , y20945 , y20946 , y20947 , y20948 , y20949 , y20950 , y20951 , y20952 , y20953 , y20954 , y20955 , y20956 , y20957 , y20958 , y20959 , y20960 , y20961 , y20962 , y20963 , y20964 , y20965 , y20966 , y20967 , y20968 , y20969 , y20970 , y20971 , y20972 , y20973 , y20974 , y20975 , y20976 , y20977 , y20978 , y20979 , y20980 , y20981 , y20982 , y20983 , y20984 , y20985 , y20986 , y20987 , y20988 , y20989 , y20990 , y20991 , y20992 , y20993 , y20994 , y20995 , y20996 , y20997 , y20998 , y20999 , y21000 , y21001 , y21002 , y21003 , y21004 , y21005 , y21006 , y21007 , y21008 , y21009 , y21010 , y21011 , y21012 , y21013 , y21014 , y21015 , y21016 , y21017 , y21018 , y21019 , y21020 , y21021 , y21022 , y21023 , y21024 , y21025 , y21026 , y21027 , y21028 , y21029 , y21030 , y21031 , y21032 , y21033 , y21034 , y21035 , y21036 , y21037 , y21038 , y21039 , y21040 , y21041 , y21042 , y21043 , y21044 , y21045 , y21046 , y21047 , y21048 , y21049 , y21050 , y21051 , y21052 , y21053 , y21054 , y21055 , y21056 , y21057 , y21058 , y21059 , y21060 , y21061 , y21062 , y21063 , y21064 , y21065 , y21066 , y21067 , y21068 , y21069 , y21070 , y21071 , y21072 , y21073 , y21074 , y21075 , y21076 , y21077 , y21078 , y21079 , y21080 , y21081 , y21082 , y21083 , y21084 , y21085 , y21086 , y21087 , y21088 , y21089 , y21090 , y21091 , y21092 , y21093 , y21094 , y21095 , y21096 , y21097 , y21098 , y21099 , y21100 , y21101 , y21102 , y21103 , y21104 , y21105 , y21106 , y21107 , y21108 , y21109 , y21110 , y21111 , y21112 , y21113 , y21114 , y21115 , y21116 , y21117 , y21118 , y21119 , y21120 , y21121 , y21122 , y21123 , y21124 , y21125 , y21126 , y21127 , y21128 , y21129 , y21130 , y21131 , y21132 , y21133 , y21134 , y21135 , y21136 , y21137 , y21138 , y21139 , y21140 , y21141 , y21142 , y21143 , y21144 , y21145 , y21146 , y21147 , y21148 , y21149 , y21150 , y21151 , y21152 , y21153 , y21154 , y21155 , y21156 , y21157 , y21158 , y21159 , y21160 , y21161 , y21162 , y21163 , y21164 , y21165 , y21166 , y21167 , y21168 , y21169 , y21170 , y21171 , y21172 , y21173 , y21174 , y21175 , y21176 , y21177 , y21178 , y21179 , y21180 , y21181 , y21182 , y21183 , y21184 , y21185 , y21186 , y21187 , y21188 , y21189 , y21190 , y21191 , y21192 , y21193 , y21194 , y21195 , y21196 , y21197 , y21198 , y21199 , y21200 , y21201 , y21202 , y21203 , y21204 , y21205 , y21206 , y21207 , y21208 , y21209 , y21210 , y21211 , y21212 , y21213 , y21214 , y21215 , y21216 , y21217 , y21218 , y21219 , y21220 , y21221 , y21222 , y21223 , y21224 , y21225 , y21226 , y21227 , y21228 , y21229 , y21230 , y21231 , y21232 , y21233 , y21234 , y21235 , y21236 , y21237 , y21238 , y21239 , y21240 , y21241 , y21242 , y21243 , y21244 , y21245 , y21246 , y21247 , y21248 , y21249 , y21250 , y21251 , y21252 , y21253 , y21254 , y21255 , y21256 , y21257 , y21258 , y21259 , y21260 , y21261 , y21262 , y21263 , y21264 , y21265 , y21266 , y21267 , y21268 , y21269 , y21270 , y21271 , y21272 , y21273 , y21274 , y21275 , y21276 , y21277 , y21278 , y21279 , y21280 , y21281 , y21282 , y21283 , y21284 , y21285 , y21286 , y21287 , y21288 , y21289 , y21290 , y21291 , y21292 , y21293 , y21294 , y21295 , y21296 , y21297 , y21298 , y21299 , y21300 , y21301 , y21302 , y21303 , y21304 , y21305 , y21306 , y21307 , y21308 , y21309 , y21310 , y21311 , y21312 , y21313 , y21314 , y21315 , y21316 , y21317 , y21318 , y21319 , y21320 , y21321 , y21322 , y21323 , y21324 , y21325 , y21326 , y21327 , y21328 , y21329 , y21330 , y21331 , y21332 , y21333 , y21334 , y21335 , y21336 , y21337 , y21338 , y21339 , y21340 , y21341 , y21342 , y21343 , y21344 , y21345 , y21346 , y21347 , y21348 , y21349 , y21350 , y21351 , y21352 , y21353 , y21354 , y21355 , y21356 , y21357 , y21358 , y21359 , y21360 , y21361 , y21362 , y21363 , y21364 , y21365 , y21366 , y21367 , y21368 , y21369 , y21370 , y21371 , y21372 , y21373 , y21374 , y21375 , y21376 , y21377 , y21378 , y21379 , y21380 , y21381 , y21382 , y21383 , y21384 , y21385 , y21386 , y21387 , y21388 , y21389 , y21390 , y21391 , y21392 , y21393 , y21394 , y21395 , y21396 , y21397 , y21398 , y21399 , y21400 , y21401 , y21402 , y21403 , y21404 , y21405 , y21406 , y21407 , y21408 , y21409 , y21410 , y21411 , y21412 , y21413 , y21414 , y21415 , y21416 , y21417 , y21418 , y21419 , y21420 , y21421 , y21422 , y21423 , y21424 , y21425 , y21426 , y21427 , y21428 , y21429 , y21430 , y21431 , y21432 , y21433 , y21434 , y21435 , y21436 , y21437 , y21438 , y21439 , y21440 , y21441 , y21442 , y21443 , y21444 , y21445 , y21446 , y21447 , y21448 , y21449 , y21450 , y21451 , y21452 , y21453 , y21454 , y21455 , y21456 , y21457 , y21458 , y21459 , y21460 , y21461 , y21462 , y21463 , y21464 , y21465 , y21466 , y21467 , y21468 , y21469 , y21470 , y21471 , y21472 , y21473 , y21474 , y21475 , y21476 , y21477 , y21478 , y21479 , y21480 , y21481 , y21482 , y21483 , y21484 , y21485 , y21486 , y21487 , y21488 , y21489 , y21490 , y21491 , y21492 , y21493 , y21494 , y21495 , y21496 , y21497 , y21498 , y21499 , y21500 , y21501 , y21502 , y21503 , y21504 , y21505 , y21506 , y21507 , y21508 , y21509 , y21510 , y21511 , y21512 , y21513 , y21514 , y21515 , y21516 , y21517 , y21518 , y21519 , y21520 , y21521 , y21522 , y21523 , y21524 , y21525 , y21526 , y21527 , y21528 , y21529 , y21530 , y21531 , y21532 , y21533 , y21534 , y21535 , y21536 , y21537 , y21538 , y21539 , y21540 , y21541 , y21542 , y21543 , y21544 , y21545 , y21546 , y21547 , y21548 , y21549 , y21550 , y21551 , y21552 , y21553 , y21554 , y21555 , y21556 , y21557 , y21558 , y21559 , y21560 , y21561 , y21562 , y21563 , y21564 , y21565 , y21566 , y21567 , y21568 , y21569 , y21570 , y21571 , y21572 , y21573 , y21574 , y21575 , y21576 , y21577 , y21578 , y21579 , y21580 , y21581 , y21582 , y21583 , y21584 , y21585 , y21586 , y21587 , y21588 , y21589 , y21590 , y21591 , y21592 , y21593 , y21594 , y21595 , y21596 , y21597 , y21598 , y21599 , y21600 , y21601 , y21602 , y21603 , y21604 , y21605 , y21606 , y21607 , y21608 , y21609 , y21610 , y21611 , y21612 , y21613 , y21614 , y21615 , y21616 , y21617 , y21618 , y21619 , y21620 , y21621 , y21622 , y21623 , y21624 , y21625 , y21626 , y21627 , y21628 , y21629 , y21630 , y21631 , y21632 , y21633 , y21634 , y21635 , y21636 , y21637 , y21638 , y21639 , y21640 , y21641 , y21642 , y21643 , y21644 , y21645 , y21646 , y21647 , y21648 , y21649 , y21650 , y21651 , y21652 , y21653 , y21654 , y21655 , y21656 , y21657 , y21658 , y21659 , y21660 , y21661 , y21662 , y21663 , y21664 , y21665 , y21666 , y21667 , y21668 , y21669 , y21670 , y21671 , y21672 , y21673 , y21674 , y21675 , y21676 , y21677 , y21678 , y21679 , y21680 , y21681 , y21682 , y21683 , y21684 , y21685 , y21686 , y21687 , y21688 , y21689 , y21690 , y21691 , y21692 , y21693 , y21694 , y21695 , y21696 , y21697 , y21698 , y21699 , y21700 , y21701 , y21702 , y21703 , y21704 , y21705 , y21706 , y21707 , y21708 , y21709 , y21710 , y21711 , y21712 , y21713 , y21714 , y21715 , y21716 , y21717 , y21718 , y21719 , y21720 , y21721 , y21722 , y21723 , y21724 , y21725 , y21726 , y21727 , y21728 , y21729 , y21730 , y21731 , y21732 , y21733 , y21734 , y21735 , y21736 , y21737 , y21738 , y21739 , y21740 , y21741 , y21742 , y21743 , y21744 , y21745 , y21746 , y21747 , y21748 , y21749 , y21750 , y21751 , y21752 , y21753 , y21754 , y21755 , y21756 , y21757 , y21758 , y21759 , y21760 , y21761 , y21762 , y21763 , y21764 , y21765 , y21766 , y21767 , y21768 , y21769 , y21770 , y21771 , y21772 , y21773 , y21774 , y21775 , y21776 , y21777 , y21778 , y21779 , y21780 , y21781 , y21782 , y21783 , y21784 , y21785 , y21786 , y21787 , y21788 , y21789 , y21790 , y21791 , y21792 , y21793 , y21794 , y21795 , y21796 , y21797 , y21798 , y21799 , y21800 , y21801 , y21802 , y21803 , y21804 , y21805 , y21806 , y21807 , y21808 , y21809 , y21810 , y21811 , y21812 , y21813 , y21814 , y21815 , y21816 , y21817 , y21818 , y21819 , y21820 , y21821 , y21822 , y21823 , y21824 , y21825 , y21826 , y21827 , y21828 , y21829 , y21830 , y21831 , y21832 , y21833 , y21834 , y21835 , y21836 , y21837 , y21838 , y21839 , y21840 , y21841 , y21842 , y21843 , y21844 , y21845 , y21846 , y21847 , y21848 , y21849 , y21850 , y21851 , y21852 , y21853 , y21854 , y21855 , y21856 , y21857 , y21858 , y21859 , y21860 , y21861 , y21862 , y21863 , y21864 , y21865 , y21866 , y21867 , y21868 , y21869 , y21870 , y21871 , y21872 , y21873 , y21874 , y21875 , y21876 , y21877 , y21878 , y21879 , y21880 , y21881 , y21882 , y21883 , y21884 , y21885 , y21886 , y21887 , y21888 , y21889 , y21890 , y21891 , y21892 , y21893 , y21894 , y21895 , y21896 , y21897 , y21898 , y21899 , y21900 , y21901 , y21902 , y21903 , y21904 , y21905 , y21906 , y21907 , y21908 , y21909 , y21910 , y21911 , y21912 , y21913 , y21914 , y21915 , y21916 , y21917 , y21918 , y21919 , y21920 , y21921 , y21922 , y21923 , y21924 , y21925 , y21926 , y21927 , y21928 , y21929 , y21930 , y21931 , y21932 , y21933 , y21934 , y21935 , y21936 , y21937 , y21938 , y21939 , y21940 , y21941 , y21942 , y21943 , y21944 , y21945 , y21946 , y21947 , y21948 , y21949 , y21950 , y21951 , y21952 , y21953 , y21954 , y21955 , y21956 , y21957 , y21958 , y21959 , y21960 , y21961 , y21962 , y21963 , y21964 , y21965 , y21966 , y21967 , y21968 , y21969 , y21970 , y21971 , y21972 , y21973 , y21974 , y21975 , y21976 , y21977 , y21978 , y21979 , y21980 , y21981 , y21982 , y21983 , y21984 , y21985 , y21986 , y21987 , y21988 , y21989 , y21990 , y21991 , y21992 , y21993 , y21994 , y21995 , y21996 , y21997 , y21998 , y21999 , y22000 , y22001 , y22002 , y22003 , y22004 , y22005 , y22006 , y22007 , y22008 , y22009 , y22010 , y22011 , y22012 , y22013 , y22014 , y22015 , y22016 , y22017 , y22018 , y22019 , y22020 , y22021 , y22022 , y22023 , y22024 , y22025 , y22026 , y22027 , y22028 , y22029 , y22030 , y22031 , y22032 , y22033 , y22034 , y22035 , y22036 , y22037 , y22038 , y22039 , y22040 , y22041 , y22042 , y22043 , y22044 , y22045 , y22046 , y22047 , y22048 , y22049 , y22050 , y22051 , y22052 , y22053 , y22054 , y22055 , y22056 , y22057 , y22058 , y22059 , y22060 , y22061 , y22062 , y22063 , y22064 , y22065 , y22066 , y22067 , y22068 , y22069 , y22070 , y22071 , y22072 , y22073 , y22074 , y22075 , y22076 , y22077 , y22078 , y22079 , y22080 , y22081 , y22082 , y22083 , y22084 , y22085 , y22086 , y22087 , y22088 , y22089 , y22090 , y22091 , y22092 , y22093 , y22094 , y22095 , y22096 , y22097 , y22098 , y22099 , y22100 , y22101 , y22102 , y22103 , y22104 , y22105 , y22106 , y22107 , y22108 , y22109 , y22110 , y22111 , y22112 , y22113 , y22114 , y22115 , y22116 , y22117 , y22118 , y22119 , y22120 , y22121 , y22122 , y22123 , y22124 , y22125 , y22126 , y22127 , y22128 , y22129 , y22130 , y22131 , y22132 , y22133 , y22134 , y22135 , y22136 , y22137 , y22138 , y22139 , y22140 , y22141 , y22142 , y22143 , y22144 , y22145 , y22146 , y22147 , y22148 , y22149 , y22150 , y22151 , y22152 , y22153 , y22154 , y22155 , y22156 , y22157 , y22158 , y22159 , y22160 , y22161 , y22162 , y22163 , y22164 , y22165 , y22166 , y22167 , y22168 , y22169 , y22170 , y22171 , y22172 , y22173 , y22174 , y22175 , y22176 , y22177 , y22178 , y22179 , y22180 , y22181 , y22182 , y22183 , y22184 , y22185 , y22186 , y22187 , y22188 , y22189 , y22190 , y22191 , y22192 , y22193 , y22194 , y22195 , y22196 , y22197 , y22198 , y22199 , y22200 , y22201 , y22202 , y22203 , y22204 , y22205 , y22206 , y22207 , y22208 , y22209 , y22210 , y22211 , y22212 , y22213 , y22214 , y22215 , y22216 , y22217 , y22218 , y22219 , y22220 , y22221 , y22222 , y22223 , y22224 , y22225 , y22226 , y22227 , y22228 , y22229 , y22230 , y22231 , y22232 , y22233 , y22234 , y22235 , y22236 , y22237 , y22238 , y22239 , y22240 , y22241 , y22242 , y22243 , y22244 , y22245 , y22246 , y22247 , y22248 , y22249 , y22250 , y22251 , y22252 , y22253 , y22254 , y22255 , y22256 , y22257 , y22258 , y22259 , y22260 , y22261 , y22262 , y22263 , y22264 , y22265 , y22266 , y22267 , y22268 , y22269 , y22270 , y22271 , y22272 , y22273 , y22274 , y22275 , y22276 , y22277 , y22278 , y22279 , y22280 , y22281 , y22282 , y22283 , y22284 , y22285 , y22286 , y22287 , y22288 , y22289 , y22290 , y22291 , y22292 , y22293 , y22294 , y22295 , y22296 , y22297 , y22298 , y22299 , y22300 , y22301 , y22302 , y22303 , y22304 , y22305 , y22306 , y22307 , y22308 , y22309 , y22310 , y22311 , y22312 , y22313 , y22314 , y22315 , y22316 , y22317 , y22318 , y22319 , y22320 , y22321 , y22322 , y22323 , y22324 , y22325 , y22326 , y22327 , y22328 , y22329 , y22330 , y22331 , y22332 , y22333 , y22334 , y22335 , y22336 , y22337 , y22338 , y22339 , y22340 , y22341 , y22342 , y22343 , y22344 , y22345 , y22346 , y22347 , y22348 , y22349 , y22350 , y22351 , y22352 , y22353 , y22354 , y22355 , y22356 , y22357 , y22358 , y22359 , y22360 , y22361 , y22362 , y22363 , y22364 , y22365 , y22366 , y22367 , y22368 , y22369 , y22370 , y22371 , y22372 , y22373 , y22374 , y22375 , y22376 , y22377 , y22378 , y22379 , y22380 , y22381 , y22382 , y22383 , y22384 , y22385 , y22386 , y22387 , y22388 , y22389 , y22390 , y22391 , y22392 , y22393 , y22394 , y22395 , y22396 , y22397 , y22398 , y22399 , y22400 , y22401 , y22402 , y22403 , y22404 , y22405 , y22406 , y22407 , y22408 , y22409 , y22410 , y22411 , y22412 , y22413 , y22414 , y22415 , y22416 , y22417 , y22418 , y22419 , y22420 , y22421 , y22422 , y22423 , y22424 , y22425 , y22426 , y22427 , y22428 , y22429 , y22430 , y22431 , y22432 , y22433 , y22434 , y22435 , y22436 , y22437 , y22438 , y22439 , y22440 , y22441 , y22442 , y22443 , y22444 , y22445 , y22446 , y22447 , y22448 , y22449 , y22450 , y22451 , y22452 , y22453 , y22454 , y22455 , y22456 , y22457 , y22458 , y22459 , y22460 , y22461 , y22462 , y22463 , y22464 , y22465 , y22466 , y22467 , y22468 , y22469 , y22470 , y22471 , y22472 , y22473 , y22474 , y22475 , y22476 , y22477 , y22478 , y22479 , y22480 , y22481 , y22482 , y22483 , y22484 , y22485 , y22486 , y22487 , y22488 , y22489 , y22490 , y22491 , y22492 , y22493 , y22494 , y22495 , y22496 , y22497 , y22498 , y22499 , y22500 , y22501 , y22502 , y22503 , y22504 , y22505 , y22506 , y22507 , y22508 , y22509 , y22510 , y22511 , y22512 , y22513 , y22514 , y22515 , y22516 , y22517 , y22518 , y22519 , y22520 , y22521 , y22522 , y22523 , y22524 , y22525 , y22526 , y22527 , y22528 , y22529 , y22530 , y22531 , y22532 , y22533 , y22534 , y22535 , y22536 , y22537 , y22538 , y22539 , y22540 , y22541 , y22542 , y22543 , y22544 , y22545 , y22546 , y22547 , y22548 , y22549 , y22550 , y22551 , y22552 , y22553 , y22554 , y22555 , y22556 , y22557 , y22558 , y22559 , y22560 , y22561 , y22562 , y22563 , y22564 , y22565 , y22566 , y22567 , y22568 , y22569 , y22570 , y22571 , y22572 , y22573 , y22574 , y22575 , y22576 , y22577 , y22578 , y22579 , y22580 , y22581 , y22582 , y22583 , y22584 , y22585 , y22586 , y22587 , y22588 , y22589 , y22590 , y22591 , y22592 , y22593 , y22594 , y22595 , y22596 , y22597 , y22598 , y22599 , y22600 , y22601 , y22602 , y22603 , y22604 , y22605 , y22606 , y22607 , y22608 , y22609 , y22610 , y22611 , y22612 , y22613 , y22614 , y22615 , y22616 , y22617 , y22618 , y22619 , y22620 , y22621 , y22622 , y22623 , y22624 , y22625 , y22626 , y22627 , y22628 , y22629 , y22630 , y22631 , y22632 , y22633 , y22634 , y22635 , y22636 , y22637 , y22638 , y22639 , y22640 , y22641 , y22642 , y22643 , y22644 , y22645 , y22646 , y22647 , y22648 , y22649 , y22650 , y22651 , y22652 , y22653 , y22654 , y22655 , y22656 , y22657 , y22658 , y22659 , y22660 , y22661 , y22662 , y22663 , y22664 , y22665 , y22666 , y22667 , y22668 , y22669 , y22670 , y22671 , y22672 , y22673 , y22674 , y22675 , y22676 , y22677 , y22678 , y22679 , y22680 , y22681 , y22682 , y22683 , y22684 , y22685 , y22686 , y22687 , y22688 , y22689 , y22690 , y22691 , y22692 , y22693 , y22694 , y22695 , y22696 , y22697 , y22698 , y22699 , y22700 , y22701 , y22702 , y22703 , y22704 , y22705 , y22706 , y22707 , y22708 , y22709 , y22710 , y22711 , y22712 , y22713 , y22714 , y22715 , y22716 , y22717 , y22718 , y22719 , y22720 , y22721 , y22722 , y22723 , y22724 , y22725 , y22726 , y22727 , y22728 , y22729 , y22730 , y22731 , y22732 , y22733 , y22734 , y22735 , y22736 , y22737 , y22738 , y22739 , y22740 , y22741 , y22742 , y22743 , y22744 , y22745 , y22746 , y22747 , y22748 , y22749 , y22750 , y22751 , y22752 , y22753 , y22754 , y22755 , y22756 , y22757 , y22758 , y22759 , y22760 , y22761 , y22762 , y22763 , y22764 , y22765 , y22766 , y22767 , y22768 , y22769 , y22770 , y22771 , y22772 , y22773 , y22774 , y22775 , y22776 , y22777 , y22778 , y22779 , y22780 , y22781 , y22782 , y22783 , y22784 , y22785 , y22786 , y22787 , y22788 , y22789 , y22790 , y22791 , y22792 , y22793 , y22794 , y22795 , y22796 , y22797 , y22798 , y22799 , y22800 , y22801 , y22802 , y22803 , y22804 , y22805 , y22806 , y22807 , y22808 , y22809 , y22810 , y22811 , y22812 , y22813 , y22814 , y22815 , y22816 , y22817 , y22818 , y22819 , y22820 , y22821 , y22822 , y22823 , y22824 , y22825 , y22826 , y22827 , y22828 , y22829 , y22830 , y22831 , y22832 , y22833 , y22834 , y22835 , y22836 , y22837 , y22838 , y22839 , y22840 , y22841 , y22842 , y22843 , y22844 , y22845 , y22846 , y22847 , y22848 , y22849 , y22850 , y22851 , y22852 , y22853 , y22854 , y22855 , y22856 , y22857 , y22858 , y22859 , y22860 , y22861 , y22862 , y22863 , y22864 , y22865 , y22866 , y22867 , y22868 , y22869 , y22870 , y22871 , y22872 , y22873 , y22874 , y22875 , y22876 , y22877 , y22878 , y22879 , y22880 , y22881 , y22882 , y22883 , y22884 , y22885 , y22886 , y22887 , y22888 , y22889 , y22890 , y22891 , y22892 , y22893 , y22894 , y22895 , y22896 , y22897 , y22898 , y22899 , y22900 , y22901 , y22902 , y22903 , y22904 , y22905 , y22906 , y22907 , y22908 , y22909 , y22910 , y22911 , y22912 , y22913 , y22914 , y22915 , y22916 , y22917 , y22918 , y22919 , y22920 , y22921 , y22922 , y22923 , y22924 , y22925 , y22926 , y22927 , y22928 , y22929 , y22930 , y22931 , y22932 , y22933 , y22934 , y22935 , y22936 , y22937 , y22938 , y22939 , y22940 , y22941 , y22942 , y22943 , y22944 , y22945 , y22946 , y22947 , y22948 , y22949 , y22950 , y22951 , y22952 , y22953 , y22954 , y22955 , y22956 , y22957 , y22958 , y22959 , y22960 , y22961 , y22962 , y22963 , y22964 , y22965 , y22966 , y22967 , y22968 , y22969 , y22970 , y22971 , y22972 , y22973 , y22974 , y22975 , y22976 , y22977 , y22978 , y22979 , y22980 , y22981 , y22982 , y22983 , y22984 , y22985 , y22986 , y22987 , y22988 , y22989 , y22990 , y22991 , y22992 , y22993 , y22994 , y22995 , y22996 , y22997 , y22998 , y22999 , y23000 , y23001 , y23002 , y23003 , y23004 , y23005 , y23006 , y23007 , y23008 , y23009 , y23010 , y23011 , y23012 , y23013 , y23014 , y23015 , y23016 , y23017 , y23018 , y23019 , y23020 , y23021 , y23022 , y23023 , y23024 , y23025 , y23026 , y23027 , y23028 , y23029 , y23030 , y23031 , y23032 , y23033 , y23034 , y23035 , y23036 , y23037 , y23038 , y23039 , y23040 , y23041 , y23042 , y23043 , y23044 , y23045 , y23046 , y23047 , y23048 , y23049 , y23050 , y23051 , y23052 , y23053 , y23054 , y23055 , y23056 , y23057 , y23058 , y23059 , y23060 , y23061 , y23062 , y23063 , y23064 , y23065 , y23066 , y23067 , y23068 , y23069 , y23070 , y23071 , y23072 , y23073 , y23074 , y23075 , y23076 , y23077 , y23078 , y23079 , y23080 , y23081 , y23082 , y23083 , y23084 , y23085 , y23086 , y23087 , y23088 , y23089 , y23090 , y23091 , y23092 , y23093 , y23094 , y23095 , y23096 , y23097 , y23098 , y23099 , y23100 , y23101 , y23102 , y23103 , y23104 , y23105 , y23106 , y23107 , y23108 , y23109 , y23110 , y23111 , y23112 , y23113 , y23114 , y23115 , y23116 , y23117 , y23118 , y23119 , y23120 , y23121 , y23122 , y23123 , y23124 , y23125 , y23126 , y23127 , y23128 , y23129 , y23130 , y23131 , y23132 , y23133 , y23134 , y23135 , y23136 , y23137 , y23138 , y23139 , y23140 , y23141 , y23142 , y23143 , y23144 , y23145 , y23146 , y23147 , y23148 , y23149 , y23150 , y23151 , y23152 , y23153 , y23154 , y23155 , y23156 , y23157 , y23158 , y23159 , y23160 , y23161 , y23162 , y23163 , y23164 , y23165 , y23166 , y23167 , y23168 , y23169 , y23170 , y23171 , y23172 , y23173 , y23174 , y23175 , y23176 , y23177 , y23178 , y23179 , y23180 , y23181 , y23182 , y23183 , y23184 , y23185 , y23186 , y23187 , y23188 , y23189 , y23190 , y23191 , y23192 , y23193 , y23194 , y23195 , y23196 , y23197 , y23198 , y23199 , y23200 , y23201 , y23202 , y23203 , y23204 , y23205 , y23206 , y23207 , y23208 , y23209 , y23210 , y23211 , y23212 , y23213 , y23214 , y23215 , y23216 , y23217 , y23218 , y23219 , y23220 , y23221 , y23222 , y23223 , y23224 , y23225 , y23226 , y23227 , y23228 , y23229 , y23230 , y23231 , y23232 , y23233 , y23234 , y23235 , y23236 , y23237 , y23238 , y23239 , y23240 , y23241 , y23242 , y23243 , y23244 , y23245 , y23246 , y23247 , y23248 , y23249 , y23250 , y23251 , y23252 , y23253 , y23254 , y23255 , y23256 , y23257 , y23258 , y23259 , y23260 , y23261 , y23262 , y23263 , y23264 , y23265 , y23266 , y23267 , y23268 , y23269 , y23270 , y23271 , y23272 , y23273 , y23274 , y23275 , y23276 , y23277 , y23278 , y23279 , y23280 , y23281 , y23282 , y23283 , y23284 , y23285 , y23286 , y23287 , y23288 , y23289 , y23290 , y23291 , y23292 , y23293 , y23294 , y23295 , y23296 , y23297 , y23298 , y23299 , y23300 , y23301 , y23302 , y23303 , y23304 , y23305 , y23306 , y23307 , y23308 , y23309 , y23310 , y23311 , y23312 , y23313 , y23314 , y23315 , y23316 , y23317 , y23318 , y23319 , y23320 , y23321 , y23322 , y23323 , y23324 , y23325 , y23326 , y23327 , y23328 , y23329 , y23330 , y23331 , y23332 , y23333 , y23334 , y23335 , y23336 , y23337 , y23338 , y23339 , y23340 , y23341 , y23342 , y23343 , y23344 , y23345 , y23346 , y23347 , y23348 , y23349 , y23350 , y23351 , y23352 , y23353 , y23354 , y23355 , y23356 , y23357 , y23358 , y23359 , y23360 , y23361 , y23362 , y23363 , y23364 , y23365 , y23366 , y23367 , y23368 , y23369 , y23370 , y23371 , y23372 , y23373 , y23374 , y23375 , y23376 , y23377 , y23378 , y23379 , y23380 , y23381 , y23382 , y23383 , y23384 , y23385 , y23386 , y23387 , y23388 , y23389 , y23390 , y23391 , y23392 , y23393 , y23394 , y23395 , y23396 , y23397 , y23398 , y23399 , y23400 , y23401 , y23402 , y23403 , y23404 , y23405 , y23406 , y23407 , y23408 , y23409 , y23410 , y23411 , y23412 , y23413 , y23414 , y23415 , y23416 , y23417 , y23418 , y23419 , y23420 , y23421 , y23422 , y23423 , y23424 , y23425 , y23426 , y23427 , y23428 , y23429 , y23430 , y23431 , y23432 , y23433 , y23434 , y23435 , y23436 , y23437 , y23438 , y23439 , y23440 , y23441 , y23442 , y23443 , y23444 , y23445 , y23446 , y23447 , y23448 , y23449 , y23450 , y23451 , y23452 , y23453 , y23454 , y23455 , y23456 , y23457 , y23458 , y23459 , y23460 , y23461 , y23462 , y23463 , y23464 , y23465 , y23466 , y23467 , y23468 , y23469 , y23470 , y23471 , y23472 , y23473 , y23474 , y23475 , y23476 , y23477 , y23478 , y23479 , y23480 , y23481 , y23482 , y23483 , y23484 , y23485 , y23486 , y23487 , y23488 , y23489 , y23490 , y23491 , y23492 , y23493 , y23494 , y23495 , y23496 , y23497 , y23498 , y23499 , y23500 , y23501 , y23502 , y23503 , y23504 , y23505 , y23506 , y23507 , y23508 , y23509 , y23510 , y23511 , y23512 , y23513 , y23514 , y23515 , y23516 , y23517 , y23518 , y23519 , y23520 , y23521 , y23522 , y23523 , y23524 , y23525 , y23526 , y23527 , y23528 , y23529 , y23530 , y23531 , y23532 , y23533 , y23534 , y23535 , y23536 , y23537 , y23538 , y23539 , y23540 , y23541 , y23542 , y23543 , y23544 , y23545 , y23546 , y23547 , y23548 , y23549 , y23550 , y23551 , y23552 , y23553 , y23554 , y23555 , y23556 , y23557 , y23558 , y23559 , y23560 , y23561 , y23562 , y23563 , y23564 , y23565 , y23566 , y23567 , y23568 , y23569 , y23570 , y23571 , y23572 , y23573 , y23574 , y23575 , y23576 , y23577 , y23578 , y23579 , y23580 , y23581 , y23582 , y23583 , y23584 , y23585 , y23586 , y23587 , y23588 , y23589 , y23590 , y23591 , y23592 , y23593 , y23594 , y23595 , y23596 , y23597 , y23598 , y23599 , y23600 , y23601 , y23602 , y23603 , y23604 , y23605 , y23606 , y23607 , y23608 , y23609 , y23610 , y23611 , y23612 , y23613 , y23614 , y23615 , y23616 , y23617 , y23618 , y23619 , y23620 , y23621 , y23622 , y23623 , y23624 , y23625 , y23626 , y23627 , y23628 , y23629 , y23630 , y23631 , y23632 , y23633 , y23634 , y23635 , y23636 , y23637 , y23638 , y23639 , y23640 , y23641 , y23642 , y23643 , y23644 , y23645 , y23646 , y23647 , y23648 , y23649 , y23650 , y23651 , y23652 , y23653 , y23654 , y23655 , y23656 , y23657 , y23658 , y23659 , y23660 , y23661 , y23662 , y23663 , y23664 , y23665 , y23666 , y23667 , y23668 , y23669 , y23670 , y23671 , y23672 , y23673 , y23674 , y23675 , y23676 , y23677 , y23678 , y23679 , y23680 , y23681 , y23682 , y23683 , y23684 , y23685 , y23686 , y23687 , y23688 , y23689 , y23690 , y23691 , y23692 , y23693 , y23694 , y23695 , y23696 , y23697 , y23698 , y23699 , y23700 , y23701 , y23702 , y23703 , y23704 , y23705 , y23706 , y23707 , y23708 , y23709 , y23710 , y23711 , y23712 , y23713 , y23714 , y23715 , y23716 , y23717 , y23718 , y23719 , y23720 , y23721 , y23722 , y23723 , y23724 , y23725 , y23726 , y23727 , y23728 , y23729 , y23730 , y23731 , y23732 , y23733 , y23734 , y23735 , y23736 , y23737 , y23738 , y23739 , y23740 , y23741 , y23742 , y23743 , y23744 , y23745 , y23746 , y23747 , y23748 , y23749 , y23750 , y23751 , y23752 , y23753 , y23754 , y23755 , y23756 , y23757 , y23758 , y23759 , y23760 , y23761 , y23762 , y23763 , y23764 , y23765 , y23766 , y23767 , y23768 , y23769 , y23770 , y23771 , y23772 , y23773 , y23774 , y23775 , y23776 , y23777 , y23778 , y23779 , y23780 , y23781 , y23782 , y23783 , y23784 , y23785 , y23786 , y23787 , y23788 , y23789 , y23790 , y23791 , y23792 , y23793 , y23794 , y23795 , y23796 , y23797 , y23798 , y23799 , y23800 , y23801 , y23802 , y23803 , y23804 , y23805 , y23806 , y23807 , y23808 , y23809 , y23810 , y23811 , y23812 , y23813 , y23814 , y23815 , y23816 , y23817 , y23818 , y23819 , y23820 , y23821 , y23822 , y23823 , y23824 , y23825 , y23826 , y23827 , y23828 , y23829 , y23830 , y23831 , y23832 , y23833 , y23834 , y23835 , y23836 , y23837 , y23838 , y23839 , y23840 , y23841 , y23842 , y23843 , y23844 , y23845 , y23846 , y23847 , y23848 , y23849 , y23850 , y23851 , y23852 , y23853 , y23854 , y23855 , y23856 , y23857 , y23858 , y23859 , y23860 , y23861 , y23862 , y23863 , y23864 , y23865 , y23866 , y23867 , y23868 , y23869 , y23870 , y23871 , y23872 , y23873 , y23874 , y23875 , y23876 , y23877 , y23878 , y23879 , y23880 , y23881 , y23882 , y23883 , y23884 , y23885 , y23886 , y23887 , y23888 , y23889 , y23890 , y23891 , y23892 , y23893 , y23894 , y23895 , y23896 , y23897 , y23898 , y23899 , y23900 , y23901 , y23902 , y23903 , y23904 , y23905 , y23906 , y23907 , y23908 , y23909 , y23910 , y23911 , y23912 , y23913 , y23914 , y23915 , y23916 , y23917 , y23918 , y23919 , y23920 , y23921 , y23922 , y23923 , y23924 , y23925 , y23926 , y23927 , y23928 , y23929 , y23930 , y23931 , y23932 , y23933 , y23934 , y23935 , y23936 , y23937 , y23938 , y23939 , y23940 , y23941 , y23942 , y23943 , y23944 , y23945 , y23946 , y23947 , y23948 , y23949 , y23950 , y23951 , y23952 , y23953 , y23954 , y23955 , y23956 , y23957 , y23958 , y23959 , y23960 , y23961 , y23962 , y23963 , y23964 , y23965 , y23966 , y23967 , y23968 , y23969 , y23970 , y23971 , y23972 , y23973 , y23974 , y23975 , y23976 , y23977 , y23978 , y23979 , y23980 , y23981 , y23982 , y23983 , y23984 , y23985 , y23986 , y23987 , y23988 , y23989 , y23990 , y23991 , y23992 , y23993 , y23994 , y23995 , y23996 , y23997 , y23998 , y23999 , y24000 , y24001 , y24002 , y24003 , y24004 , y24005 , y24006 , y24007 , y24008 , y24009 , y24010 , y24011 , y24012 , y24013 , y24014 , y24015 , y24016 , y24017 , y24018 , y24019 , y24020 , y24021 , y24022 , y24023 , y24024 , y24025 , y24026 , y24027 , y24028 , y24029 , y24030 , y24031 , y24032 , y24033 , y24034 , y24035 , y24036 , y24037 , y24038 , y24039 , y24040 , y24041 , y24042 , y24043 , y24044 , y24045 , y24046 , y24047 , y24048 , y24049 , y24050 , y24051 , y24052 , y24053 , y24054 , y24055 , y24056 , y24057 , y24058 , y24059 , y24060 , y24061 , y24062 , y24063 , y24064 , y24065 , y24066 , y24067 , y24068 , y24069 , y24070 , y24071 , y24072 , y24073 , y24074 , y24075 , y24076 , y24077 , y24078 , y24079 , y24080 , y24081 , y24082 , y24083 , y24084 , y24085 , y24086 , y24087 , y24088 , y24089 , y24090 , y24091 , y24092 , y24093 , y24094 , y24095 , y24096 , y24097 , y24098 , y24099 , y24100 , y24101 , y24102 , y24103 , y24104 , y24105 , y24106 , y24107 , y24108 , y24109 , y24110 , y24111 , y24112 , y24113 , y24114 , y24115 , y24116 , y24117 , y24118 , y24119 , y24120 , y24121 , y24122 , y24123 , y24124 , y24125 , y24126 , y24127 , y24128 , y24129 , y24130 , y24131 , y24132 , y24133 , y24134 , y24135 , y24136 , y24137 , y24138 , y24139 , y24140 , y24141 , y24142 , y24143 , y24144 , y24145 , y24146 , y24147 , y24148 , y24149 , y24150 , y24151 , y24152 , y24153 , y24154 , y24155 , y24156 , y24157 , y24158 , y24159 , y24160 , y24161 , y24162 , y24163 , y24164 , y24165 , y24166 , y24167 , y24168 , y24169 , y24170 , y24171 , y24172 , y24173 , y24174 , y24175 , y24176 , y24177 , y24178 , y24179 , y24180 , y24181 , y24182 , y24183 , y24184 , y24185 , y24186 , y24187 , y24188 , y24189 , y24190 , y24191 , y24192 , y24193 , y24194 , y24195 , y24196 , y24197 , y24198 , y24199 , y24200 , y24201 , y24202 , y24203 , y24204 , y24205 , y24206 , y24207 , y24208 , y24209 , y24210 , y24211 , y24212 , y24213 , y24214 , y24215 , y24216 , y24217 , y24218 , y24219 , y24220 , y24221 , y24222 , y24223 , y24224 , y24225 , y24226 , y24227 , y24228 , y24229 , y24230 , y24231 , y24232 , y24233 , y24234 , y24235 , y24236 , y24237 , y24238 , y24239 , y24240 , y24241 , y24242 , y24243 , y24244 , y24245 , y24246 , y24247 , y24248 , y24249 , y24250 , y24251 , y24252 , y24253 , y24254 , y24255 , y24256 , y24257 , y24258 , y24259 , y24260 , y24261 , y24262 , y24263 , y24264 , y24265 , y24266 , y24267 , y24268 , y24269 , y24270 , y24271 , y24272 , y24273 , y24274 , y24275 , y24276 , y24277 , y24278 , y24279 , y24280 , y24281 , y24282 , y24283 , y24284 , y24285 , y24286 , y24287 , y24288 , y24289 , y24290 , y24291 , y24292 , y24293 , y24294 , y24295 , y24296 , y24297 , y24298 , y24299 , y24300 , y24301 , y24302 , y24303 , y24304 , y24305 , y24306 , y24307 , y24308 , y24309 , y24310 , y24311 , y24312 , y24313 , y24314 , y24315 , y24316 , y24317 , y24318 , y24319 , y24320 , y24321 , y24322 , y24323 , y24324 , y24325 , y24326 , y24327 , y24328 , y24329 , y24330 , y24331 , y24332 , y24333 , y24334 , y24335 , y24336 , y24337 , y24338 , y24339 , y24340 , y24341 , y24342 , y24343 , y24344 , y24345 , y24346 , y24347 , y24348 , y24349 , y24350 , y24351 , y24352 , y24353 , y24354 , y24355 , y24356 , y24357 , y24358 , y24359 , y24360 , y24361 , y24362 , y24363 , y24364 , y24365 , y24366 , y24367 , y24368 , y24369 , y24370 , y24371 , y24372 , y24373 , y24374 , y24375 , y24376 , y24377 , y24378 , y24379 , y24380 , y24381 , y24382 , y24383 , y24384 , y24385 , y24386 , y24387 , y24388 , y24389 , y24390 , y24391 , y24392 , y24393 , y24394 , y24395 , y24396 , y24397 , y24398 , y24399 , y24400 , y24401 , y24402 , y24403 , y24404 , y24405 , y24406 , y24407 , y24408 , y24409 , y24410 , y24411 , y24412 , y24413 , y24414 , y24415 , y24416 , y24417 , y24418 , y24419 , y24420 , y24421 , y24422 , y24423 , y24424 , y24425 , y24426 , y24427 , y24428 , y24429 , y24430 , y24431 , y24432 , y24433 , y24434 , y24435 , y24436 , y24437 , y24438 , y24439 , y24440 , y24441 , y24442 , y24443 , y24444 , y24445 , y24446 , y24447 , y24448 , y24449 , y24450 , y24451 , y24452 , y24453 , y24454 , y24455 , y24456 , y24457 , y24458 , y24459 , y24460 , y24461 , y24462 , y24463 , y24464 , y24465 , y24466 , y24467 , y24468 , y24469 , y24470 , y24471 , y24472 , y24473 , y24474 , y24475 , y24476 , y24477 , y24478 , y24479 , y24480 , y24481 , y24482 , y24483 , y24484 , y24485 , y24486 , y24487 , y24488 , y24489 , y24490 , y24491 , y24492 , y24493 , y24494 , y24495 , y24496 , y24497 , y24498 , y24499 , y24500 , y24501 , y24502 , y24503 , y24504 , y24505 , y24506 , y24507 , y24508 , y24509 , y24510 , y24511 , y24512 , y24513 , y24514 , y24515 , y24516 , y24517 , y24518 , y24519 , y24520 , y24521 , y24522 , y24523 , y24524 , y24525 , y24526 , y24527 , y24528 , y24529 , y24530 , y24531 , y24532 , y24533 , y24534 , y24535 , y24536 , y24537 , y24538 , y24539 , y24540 , y24541 , y24542 , y24543 , y24544 , y24545 , y24546 , y24547 , y24548 , y24549 , y24550 , y24551 , y24552 , y24553 , y24554 , y24555 , y24556 , y24557 , y24558 , y24559 , y24560 , y24561 , y24562 , y24563 , y24564 , y24565 , y24566 , y24567 , y24568 , y24569 , y24570 , y24571 , y24572 , y24573 , y24574 , y24575 , y24576 , y24577 , y24578 , y24579 , y24580 , y24581 , y24582 , y24583 , y24584 , y24585 , y24586 , y24587 , y24588 , y24589 , y24590 , y24591 , y24592 , y24593 , y24594 , y24595 , y24596 , y24597 , y24598 , y24599 , y24600 , y24601 , y24602 , y24603 , y24604 , y24605 , y24606 , y24607 , y24608 , y24609 , y24610 , y24611 , y24612 , y24613 , y24614 , y24615 , y24616 , y24617 , y24618 , y24619 , y24620 , y24621 , y24622 , y24623 , y24624 , y24625 , y24626 , y24627 , y24628 , y24629 , y24630 , y24631 , y24632 , y24633 , y24634 , y24635 , y24636 , y24637 , y24638 , y24639 , y24640 , y24641 , y24642 , y24643 , y24644 , y24645 , y24646 , y24647 , y24648 , y24649 , y24650 , y24651 , y24652 , y24653 , y24654 , y24655 , y24656 , y24657 , y24658 , y24659 , y24660 , y24661 , y24662 , y24663 , y24664 , y24665 , y24666 , y24667 , y24668 , y24669 , y24670 , y24671 , y24672 , y24673 , y24674 , y24675 , y24676 , y24677 , y24678 , y24679 , y24680 , y24681 , y24682 , y24683 , y24684 , y24685 , y24686 , y24687 , y24688 , y24689 , y24690 , y24691 , y24692 , y24693 , y24694 , y24695 , y24696 , y24697 , y24698 , y24699 , y24700 , y24701 , y24702 , y24703 , y24704 , y24705 , y24706 , y24707 , y24708 , y24709 , y24710 , y24711 , y24712 , y24713 , y24714 , y24715 , y24716 , y24717 , y24718 , y24719 , y24720 , y24721 , y24722 , y24723 , y24724 , y24725 , y24726 , y24727 , y24728 , y24729 , y24730 , y24731 , y24732 , y24733 , y24734 , y24735 , y24736 , y24737 , y24738 , y24739 , y24740 , y24741 , y24742 , y24743 , y24744 , y24745 , y24746 , y24747 , y24748 , y24749 , y24750 , y24751 , y24752 , y24753 , y24754 , y24755 , y24756 , y24757 , y24758 , y24759 , y24760 , y24761 , y24762 , y24763 , y24764 , y24765 , y24766 , y24767 , y24768 , y24769 , y24770 , y24771 , y24772 , y24773 , y24774 , y24775 , y24776 , y24777 , y24778 , y24779 , y24780 , y24781 , y24782 , y24783 , y24784 , y24785 , y24786 , y24787 , y24788 , y24789 , y24790 , y24791 , y24792 , y24793 , y24794 , y24795 , y24796 , y24797 , y24798 , y24799 , y24800 , y24801 , y24802 , y24803 , y24804 , y24805 , y24806 , y24807 , y24808 , y24809 , y24810 , y24811 , y24812 , y24813 , y24814 , y24815 , y24816 , y24817 , y24818 , y24819 , y24820 , y24821 , y24822 , y24823 , y24824 , y24825 , y24826 , y24827 , y24828 , y24829 , y24830 , y24831 , y24832 , y24833 , y24834 , y24835 , y24836 , y24837 , y24838 , y24839 , y24840 , y24841 , y24842 , y24843 , y24844 , y24845 , y24846 , y24847 , y24848 , y24849 , y24850 , y24851 , y24852 , y24853 , y24854 , y24855 , y24856 , y24857 , y24858 , y24859 , y24860 , y24861 , y24862 , y24863 , y24864 , y24865 , y24866 , y24867 , y24868 , y24869 , y24870 , y24871 , y24872 , y24873 , y24874 , y24875 , y24876 , y24877 , y24878 , y24879 , y24880 , y24881 , y24882 , y24883 , y24884 , y24885 , y24886 , y24887 , y24888 , y24889 , y24890 , y24891 , y24892 , y24893 , y24894 , y24895 , y24896 , y24897 , y24898 , y24899 , y24900 , y24901 , y24902 , y24903 , y24904 , y24905 , y24906 , y24907 , y24908 , y24909 , y24910 , y24911 , y24912 , y24913 , y24914 , y24915 , y24916 , y24917 , y24918 , y24919 , y24920 , y24921 , y24922 , y24923 , y24924 , y24925 , y24926 , y24927 , y24928 , y24929 , y24930 , y24931 , y24932 , y24933 , y24934 , y24935 , y24936 , y24937 , y24938 , y24939 , y24940 , y24941 , y24942 , y24943 , y24944 , y24945 , y24946 , y24947 , y24948 , y24949 , y24950 , y24951 , y24952 , y24953 , y24954 , y24955 , y24956 , y24957 , y24958 , y24959 , y24960 , y24961 , y24962 , y24963 , y24964 , y24965 , y24966 , y24967 , y24968 , y24969 , y24970 , y24971 , y24972 , y24973 , y24974 , y24975 , y24976 , y24977 , y24978 , y24979 , y24980 , y24981 , y24982 , y24983 , y24984 , y24985 , y24986 , y24987 , y24988 , y24989 , y24990 , y24991 , y24992 , y24993 , y24994 , y24995 , y24996 , y24997 , y24998 , y24999 , y25000 , y25001 , y25002 , y25003 , y25004 , y25005 , y25006 , y25007 , y25008 , y25009 , y25010 , y25011 , y25012 , y25013 , y25014 , y25015 , y25016 , y25017 , y25018 , y25019 , y25020 , y25021 , y25022 , y25023 , y25024 , y25025 , y25026 , y25027 , y25028 , y25029 , y25030 , y25031 , y25032 , y25033 , y25034 , y25035 , y25036 , y25037 , y25038 , y25039 , y25040 , y25041 , y25042 , y25043 , y25044 , y25045 , y25046 , y25047 , y25048 , y25049 , y25050 , y25051 , y25052 , y25053 , y25054 , y25055 , y25056 , y25057 , y25058 , y25059 , y25060 , y25061 , y25062 , y25063 , y25064 , y25065 , y25066 , y25067 , y25068 , y25069 , y25070 , y25071 , y25072 , y25073 , y25074 , y25075 , y25076 , y25077 , y25078 , y25079 , y25080 , y25081 , y25082 , y25083 , y25084 , y25085 , y25086 , y25087 , y25088 , y25089 , y25090 , y25091 , y25092 , y25093 , y25094 , y25095 , y25096 , y25097 , y25098 , y25099 , y25100 , y25101 , y25102 , y25103 , y25104 , y25105 , y25106 , y25107 , y25108 , y25109 , y25110 , y25111 , y25112 , y25113 , y25114 , y25115 , y25116 , y25117 , y25118 , y25119 , y25120 , y25121 , y25122 , y25123 , y25124 , y25125 , y25126 , y25127 , y25128 , y25129 , y25130 , y25131 , y25132 , y25133 , y25134 , y25135 , y25136 , y25137 , y25138 , y25139 , y25140 , y25141 , y25142 , y25143 , y25144 , y25145 , y25146 , y25147 , y25148 , y25149 , y25150 , y25151 , y25152 , y25153 , y25154 , y25155 , y25156 , y25157 , y25158 , y25159 , y25160 , y25161 , y25162 , y25163 , y25164 , y25165 , y25166 , y25167 , y25168 , y25169 , y25170 , y25171 , y25172 , y25173 , y25174 , y25175 , y25176 , y25177 , y25178 , y25179 , y25180 , y25181 , y25182 , y25183 , y25184 , y25185 , y25186 , y25187 , y25188 , y25189 , y25190 , y25191 , y25192 , y25193 , y25194 , y25195 , y25196 , y25197 , y25198 , y25199 , y25200 , y25201 , y25202 , y25203 , y25204 , y25205 , y25206 , y25207 , y25208 , y25209 , y25210 , y25211 , y25212 , y25213 , y25214 , y25215 , y25216 , y25217 , y25218 , y25219 , y25220 , y25221 , y25222 , y25223 , y25224 , y25225 , y25226 , y25227 , y25228 , y25229 , y25230 , y25231 , y25232 , y25233 , y25234 , y25235 , y25236 , y25237 , y25238 , y25239 , y25240 , y25241 , y25242 , y25243 , y25244 , y25245 , y25246 , y25247 , y25248 , y25249 , y25250 , y25251 , y25252 , y25253 , y25254 , y25255 , y25256 , y25257 , y25258 , y25259 , y25260 , y25261 , y25262 , y25263 , y25264 , y25265 , y25266 , y25267 , y25268 , y25269 , y25270 , y25271 , y25272 , y25273 , y25274 , y25275 , y25276 , y25277 , y25278 , y25279 , y25280 , y25281 , y25282 , y25283 , y25284 , y25285 , y25286 , y25287 , y25288 , y25289 , y25290 , y25291 , y25292 , y25293 , y25294 , y25295 , y25296 , y25297 , y25298 , y25299 , y25300 , y25301 , y25302 , y25303 , y25304 , y25305 , y25306 , y25307 , y25308 , y25309 , y25310 , y25311 , y25312 , y25313 , y25314 , y25315 , y25316 , y25317 , y25318 , y25319 , y25320 , y25321 , y25322 , y25323 , y25324 , y25325 , y25326 , y25327 , y25328 , y25329 , y25330 , y25331 , y25332 , y25333 , y25334 , y25335 , y25336 , y25337 , y25338 , y25339 , y25340 , y25341 , y25342 , y25343 , y25344 , y25345 , y25346 , y25347 , y25348 , y25349 , y25350 , y25351 , y25352 , y25353 , y25354 , y25355 , y25356 , y25357 , y25358 , y25359 , y25360 , y25361 , y25362 , y25363 , y25364 , y25365 , y25366 , y25367 , y25368 , y25369 , y25370 , y25371 , y25372 , y25373 , y25374 , y25375 , y25376 , y25377 , y25378 , y25379 , y25380 , y25381 , y25382 , y25383 , y25384 , y25385 , y25386 , y25387 , y25388 , y25389 , y25390 , y25391 , y25392 , y25393 , y25394 , y25395 , y25396 , y25397 , y25398 , y25399 , y25400 , y25401 , y25402 , y25403 , y25404 , y25405 , y25406 , y25407 , y25408 , y25409 , y25410 , y25411 , y25412 , y25413 , y25414 , y25415 , y25416 , y25417 , y25418 , y25419 , y25420 , y25421 , y25422 , y25423 , y25424 , y25425 , y25426 , y25427 , y25428 , y25429 , y25430 , y25431 , y25432 , y25433 , y25434 , y25435 , y25436 , y25437 , y25438 , y25439 , y25440 , y25441 , y25442 , y25443 , y25444 , y25445 , y25446 , y25447 , y25448 , y25449 , y25450 , y25451 , y25452 , y25453 , y25454 , y25455 , y25456 , y25457 , y25458 , y25459 , y25460 , y25461 , y25462 , y25463 , y25464 , y25465 , y25466 , y25467 , y25468 , y25469 , y25470 , y25471 , y25472 , y25473 , y25474 , y25475 , y25476 , y25477 , y25478 , y25479 , y25480 , y25481 , y25482 , y25483 , y25484 , y25485 , y25486 , y25487 , y25488 , y25489 , y25490 , y25491 , y25492 , y25493 , y25494 , y25495 , y25496 , y25497 , y25498 , y25499 , y25500 , y25501 , y25502 , y25503 , y25504 , y25505 , y25506 , y25507 , y25508 , y25509 , y25510 , y25511 , y25512 , y25513 , y25514 , y25515 , y25516 , y25517 , y25518 , y25519 , y25520 , y25521 , y25522 , y25523 , y25524 , y25525 , y25526 , y25527 , y25528 , y25529 , y25530 , y25531 , y25532 , y25533 , y25534 , y25535 , y25536 , y25537 , y25538 , y25539 , y25540 , y25541 , y25542 , y25543 , y25544 , y25545 , y25546 , y25547 , y25548 , y25549 , y25550 , y25551 , y25552 , y25553 , y25554 , y25555 , y25556 , y25557 , y25558 , y25559 , y25560 , y25561 , y25562 , y25563 , y25564 , y25565 , y25566 , y25567 , y25568 , y25569 , y25570 , y25571 , y25572 , y25573 , y25574 , y25575 , y25576 , y25577 , y25578 , y25579 , y25580 , y25581 , y25582 , y25583 , y25584 , y25585 , y25586 , y25587 , y25588 , y25589 , y25590 , y25591 , y25592 , y25593 , y25594 , y25595 , y25596 , y25597 , y25598 , y25599 , y25600 , y25601 , y25602 , y25603 , y25604 , y25605 , y25606 , y25607 , y25608 , y25609 , y25610 , y25611 , y25612 , y25613 , y25614 , y25615 , y25616 , y25617 , y25618 , y25619 , y25620 , y25621 , y25622 , y25623 , y25624 , y25625 , y25626 , y25627 , y25628 , y25629 , y25630 , y25631 , y25632 , y25633 , y25634 , y25635 , y25636 , y25637 , y25638 , y25639 , y25640 , y25641 , y25642 , y25643 , y25644 , y25645 , y25646 , y25647 , y25648 , y25649 , y25650 , y25651 , y25652 , y25653 , y25654 , y25655 , y25656 , y25657 , y25658 , y25659 , y25660 , y25661 , y25662 , y25663 , y25664 , y25665 , y25666 , y25667 , y25668 , y25669 , y25670 , y25671 , y25672 , y25673 , y25674 , y25675 , y25676 , y25677 , y25678 , y25679 , y25680 , y25681 , y25682 , y25683 , y25684 , y25685 , y25686 , y25687 , y25688 , y25689 , y25690 , y25691 , y25692 , y25693 , y25694 , y25695 , y25696 , y25697 , y25698 , y25699 , y25700 , y25701 , y25702 , y25703 , y25704 , y25705 , y25706 , y25707 , y25708 , y25709 , y25710 , y25711 , y25712 , y25713 , y25714 , y25715 , y25716 , y25717 , y25718 , y25719 , y25720 , y25721 , y25722 , y25723 , y25724 , y25725 , y25726 , y25727 , y25728 , y25729 , y25730 , y25731 , y25732 , y25733 , y25734 , y25735 , y25736 , y25737 , y25738 , y25739 , y25740 , y25741 , y25742 , y25743 , y25744 , y25745 , y25746 , y25747 , y25748 , y25749 , y25750 , y25751 , y25752 , y25753 , y25754 , y25755 , y25756 , y25757 , y25758 , y25759 , y25760 , y25761 , y25762 , y25763 , y25764 , y25765 , y25766 , y25767 , y25768 , y25769 , y25770 , y25771 , y25772 , y25773 , y25774 , y25775 , y25776 , y25777 , y25778 , y25779 , y25780 , y25781 , y25782 , y25783 , y25784 , y25785 , y25786 , y25787 , y25788 , y25789 , y25790 , y25791 , y25792 , y25793 , y25794 , y25795 , y25796 , y25797 , y25798 , y25799 , y25800 , y25801 , y25802 , y25803 , y25804 , y25805 , y25806 , y25807 , y25808 , y25809 , y25810 , y25811 , y25812 , y25813 , y25814 , y25815 , y25816 , y25817 , y25818 , y25819 , y25820 , y25821 , y25822 , y25823 , y25824 , y25825 , y25826 , y25827 , y25828 , y25829 , y25830 , y25831 , y25832 , y25833 , y25834 , y25835 , y25836 , y25837 , y25838 , y25839 , y25840 , y25841 , y25842 , y25843 , y25844 , y25845 , y25846 , y25847 , y25848 , y25849 , y25850 , y25851 , y25852 , y25853 , y25854 , y25855 , y25856 , y25857 , y25858 , y25859 , y25860 , y25861 , y25862 , y25863 , y25864 , y25865 , y25866 , y25867 , y25868 , y25869 , y25870 , y25871 , y25872 , y25873 , y25874 , y25875 , y25876 , y25877 , y25878 , y25879 , y25880 , y25881 , y25882 , y25883 , y25884 , y25885 , y25886 , y25887 , y25888 , y25889 , y25890 , y25891 , y25892 , y25893 , y25894 , y25895 , y25896 , y25897 , y25898 , y25899 , y25900 , y25901 , y25902 , y25903 , y25904 , y25905 , y25906 , y25907 , y25908 , y25909 , y25910 , y25911 , y25912 , y25913 , y25914 , y25915 , y25916 , y25917 , y25918 , y25919 , y25920 , y25921 , y25922 , y25923 , y25924 , y25925 , y25926 , y25927 , y25928 , y25929 , y25930 , y25931 , y25932 , y25933 , y25934 , y25935 , y25936 , y25937 , y25938 , y25939 , y25940 , y25941 , y25942 , y25943 , y25944 , y25945 , y25946 , y25947 , y25948 , y25949 , y25950 , y25951 , y25952 , y25953 , y25954 , y25955 , y25956 , y25957 , y25958 , y25959 , y25960 , y25961 , y25962 , y25963 , y25964 , y25965 , y25966 , y25967 , y25968 , y25969 , y25970 , y25971 , y25972 , y25973 , y25974 , y25975 , y25976 , y25977 , y25978 , y25979 , y25980 , y25981 , y25982 , y25983 , y25984 , y25985 , y25986 , y25987 , y25988 , y25989 , y25990 , y25991 , y25992 , y25993 , y25994 , y25995 , y25996 , y25997 , y25998 , y25999 , y26000 , y26001 , y26002 , y26003 , y26004 , y26005 , y26006 , y26007 , y26008 , y26009 , y26010 , y26011 , y26012 , y26013 , y26014 , y26015 , y26016 , y26017 , y26018 , y26019 , y26020 , y26021 , y26022 , y26023 , y26024 , y26025 , y26026 , y26027 , y26028 , y26029 , y26030 , y26031 , y26032 , y26033 , y26034 , y26035 , y26036 , y26037 , y26038 , y26039 , y26040 , y26041 , y26042 , y26043 , y26044 , y26045 , y26046 , y26047 , y26048 , y26049 , y26050 , y26051 , y26052 , y26053 , y26054 , y26055 , y26056 , y26057 , y26058 , y26059 , y26060 , y26061 , y26062 , y26063 , y26064 , y26065 , y26066 , y26067 , y26068 , y26069 , y26070 , y26071 , y26072 , y26073 , y26074 , y26075 , y26076 , y26077 , y26078 , y26079 , y26080 , y26081 , y26082 , y26083 , y26084 , y26085 , y26086 , y26087 , y26088 , y26089 , y26090 , y26091 , y26092 , y26093 , y26094 , y26095 , y26096 , y26097 , y26098 , y26099 , y26100 , y26101 , y26102 , y26103 , y26104 , y26105 , y26106 , y26107 , y26108 , y26109 , y26110 , y26111 , y26112 , y26113 , y26114 , y26115 , y26116 , y26117 , y26118 , y26119 , y26120 , y26121 , y26122 , y26123 , y26124 , y26125 , y26126 , y26127 , y26128 , y26129 , y26130 , y26131 , y26132 , y26133 , y26134 , y26135 , y26136 , y26137 , y26138 , y26139 , y26140 , y26141 , y26142 , y26143 , y26144 , y26145 , y26146 , y26147 , y26148 , y26149 , y26150 , y26151 , y26152 , y26153 , y26154 , y26155 , y26156 , y26157 , y26158 , y26159 , y26160 , y26161 , y26162 , y26163 , y26164 , y26165 , y26166 , y26167 , y26168 , y26169 , y26170 , y26171 , y26172 , y26173 , y26174 , y26175 , y26176 , y26177 , y26178 , y26179 , y26180 , y26181 , y26182 , y26183 , y26184 , y26185 , y26186 , y26187 , y26188 , y26189 , y26190 , y26191 , y26192 , y26193 , y26194 , y26195 , y26196 , y26197 , y26198 , y26199 , y26200 , y26201 , y26202 , y26203 , y26204 , y26205 , y26206 , y26207 , y26208 , y26209 , y26210 , y26211 , y26212 , y26213 , y26214 , y26215 , y26216 , y26217 , y26218 , y26219 , y26220 , y26221 , y26222 , y26223 , y26224 , y26225 , y26226 , y26227 , y26228 , y26229 , y26230 , y26231 , y26232 , y26233 , y26234 , y26235 , y26236 , y26237 , y26238 , y26239 , y26240 , y26241 , y26242 , y26243 , y26244 , y26245 , y26246 , y26247 , y26248 , y26249 , y26250 , y26251 , y26252 , y26253 , y26254 , y26255 , y26256 , y26257 , y26258 , y26259 , y26260 , y26261 , y26262 , y26263 , y26264 , y26265 , y26266 , y26267 , y26268 , y26269 , y26270 , y26271 , y26272 , y26273 , y26274 , y26275 , y26276 , y26277 , y26278 , y26279 , y26280 , y26281 , y26282 , y26283 , y26284 , y26285 , y26286 , y26287 , y26288 , y26289 , y26290 , y26291 , y26292 , y26293 , y26294 , y26295 , y26296 , y26297 , y26298 , y26299 , y26300 , y26301 , y26302 , y26303 , y26304 , y26305 , y26306 , y26307 , y26308 , y26309 , y26310 , y26311 , y26312 , y26313 , y26314 , y26315 , y26316 , y26317 , y26318 , y26319 , y26320 , y26321 , y26322 , y26323 , y26324 , y26325 , y26326 , y26327 , y26328 , y26329 , y26330 , y26331 , y26332 , y26333 , y26334 , y26335 , y26336 , y26337 , y26338 , y26339 , y26340 , y26341 , y26342 , y26343 , y26344 , y26345 , y26346 , y26347 , y26348 , y26349 , y26350 , y26351 , y26352 , y26353 , y26354 , y26355 , y26356 , y26357 , y26358 , y26359 , y26360 , y26361 , y26362 , y26363 , y26364 , y26365 , y26366 , y26367 , y26368 , y26369 , y26370 , y26371 , y26372 , y26373 , y26374 , y26375 , y26376 , y26377 , y26378 , y26379 , y26380 , y26381 , y26382 , y26383 , y26384 , y26385 , y26386 , y26387 , y26388 , y26389 , y26390 , y26391 , y26392 , y26393 , y26394 , y26395 , y26396 , y26397 , y26398 , y26399 , y26400 , y26401 , y26402 , y26403 , y26404 , y26405 , y26406 , y26407 , y26408 , y26409 , y26410 , y26411 , y26412 , y26413 , y26414 , y26415 , y26416 , y26417 , y26418 , y26419 , y26420 , y26421 , y26422 , y26423 , y26424 , y26425 , y26426 , y26427 , y26428 , y26429 , y26430 , y26431 , y26432 , y26433 , y26434 , y26435 , y26436 , y26437 , y26438 , y26439 , y26440 , y26441 , y26442 , y26443 , y26444 , y26445 , y26446 , y26447 , y26448 , y26449 , y26450 , y26451 , y26452 , y26453 , y26454 , y26455 , y26456 , y26457 , y26458 , y26459 , y26460 , y26461 , y26462 , y26463 , y26464 , y26465 , y26466 , y26467 , y26468 , y26469 , y26470 , y26471 , y26472 , y26473 , y26474 , y26475 , y26476 , y26477 , y26478 , y26479 , y26480 , y26481 , y26482 , y26483 , y26484 , y26485 , y26486 , y26487 , y26488 , y26489 , y26490 , y26491 , y26492 , y26493 , y26494 , y26495 , y26496 , y26497 , y26498 , y26499 , y26500 , y26501 , y26502 , y26503 , y26504 , y26505 , y26506 , y26507 , y26508 , y26509 , y26510 , y26511 , y26512 , y26513 , y26514 , y26515 , y26516 , y26517 , y26518 , y26519 , y26520 , y26521 , y26522 , y26523 , y26524 , y26525 , y26526 , y26527 , y26528 , y26529 , y26530 , y26531 , y26532 , y26533 , y26534 , y26535 , y26536 , y26537 , y26538 , y26539 , y26540 , y26541 , y26542 , y26543 , y26544 , y26545 , y26546 , y26547 , y26548 , y26549 , y26550 , y26551 , y26552 , y26553 , y26554 , y26555 , y26556 , y26557 , y26558 , y26559 , y26560 , y26561 , y26562 , y26563 , y26564 , y26565 , y26566 , y26567 , y26568 , y26569 , y26570 , y26571 , y26572 , y26573 , y26574 , y26575 , y26576 , y26577 , y26578 , y26579 , y26580 , y26581 , y26582 , y26583 , y26584 , y26585 , y26586 , y26587 , y26588 , y26589 , y26590 , y26591 , y26592 , y26593 , y26594 , y26595 , y26596 , y26597 , y26598 , y26599 , y26600 , y26601 , y26602 , y26603 , y26604 , y26605 , y26606 , y26607 , y26608 , y26609 , y26610 , y26611 , y26612 , y26613 , y26614 , y26615 , y26616 , y26617 , y26618 , y26619 , y26620 , y26621 , y26622 , y26623 , y26624 , y26625 , y26626 , y26627 , y26628 , y26629 , y26630 , y26631 , y26632 , y26633 , y26634 , y26635 , y26636 , y26637 , y26638 , y26639 , y26640 , y26641 , y26642 , y26643 , y26644 , y26645 , y26646 , y26647 , y26648 , y26649 , y26650 , y26651 , y26652 , y26653 , y26654 , y26655 , y26656 , y26657 , y26658 , y26659 , y26660 , y26661 , y26662 , y26663 , y26664 , y26665 , y26666 , y26667 , y26668 , y26669 , y26670 , y26671 , y26672 , y26673 , y26674 , y26675 , y26676 , y26677 , y26678 , y26679 , y26680 , y26681 , y26682 , y26683 , y26684 , y26685 , y26686 , y26687 , y26688 , y26689 , y26690 , y26691 , y26692 , y26693 , y26694 , y26695 , y26696 , y26697 , y26698 , y26699 , y26700 , y26701 , y26702 , y26703 , y26704 , y26705 , y26706 , y26707 , y26708 , y26709 , y26710 , y26711 , y26712 , y26713 , y26714 , y26715 , y26716 , y26717 , y26718 , y26719 , y26720 , y26721 , y26722 , y26723 , y26724 , y26725 , y26726 , y26727 , y26728 , y26729 , y26730 , y26731 , y26732 , y26733 , y26734 , y26735 , y26736 , y26737 , y26738 , y26739 , y26740 , y26741 , y26742 , y26743 , y26744 , y26745 , y26746 , y26747 , y26748 , y26749 , y26750 , y26751 , y26752 , y26753 , y26754 , y26755 , y26756 , y26757 , y26758 , y26759 , y26760 , y26761 , y26762 , y26763 , y26764 , y26765 , y26766 , y26767 , y26768 , y26769 , y26770 , y26771 , y26772 , y26773 , y26774 , y26775 , y26776 , y26777 , y26778 , y26779 , y26780 , y26781 , y26782 , y26783 , y26784 , y26785 , y26786 , y26787 , y26788 , y26789 , y26790 , y26791 , y26792 , y26793 , y26794 , y26795 , y26796 , y26797 , y26798 , y26799 , y26800 , y26801 , y26802 , y26803 , y26804 , y26805 , y26806 , y26807 , y26808 , y26809 , y26810 , y26811 , y26812 , y26813 , y26814 , y26815 , y26816 , y26817 , y26818 , y26819 , y26820 , y26821 , y26822 , y26823 , y26824 , y26825 , y26826 , y26827 , y26828 , y26829 , y26830 , y26831 , y26832 , y26833 , y26834 , y26835 , y26836 , y26837 , y26838 , y26839 , y26840 , y26841 , y26842 , y26843 , y26844 , y26845 , y26846 , y26847 , y26848 , y26849 , y26850 , y26851 , y26852 , y26853 , y26854 , y26855 , y26856 , y26857 , y26858 , y26859 , y26860 , y26861 , y26862 , y26863 , y26864 , y26865 , y26866 , y26867 , y26868 , y26869 , y26870 , y26871 , y26872 , y26873 , y26874 , y26875 , y26876 , y26877 , y26878 , y26879 , y26880 , y26881 , y26882 , y26883 , y26884 , y26885 , y26886 , y26887 , y26888 , y26889 , y26890 , y26891 , y26892 , y26893 , y26894 , y26895 , y26896 , y26897 , y26898 , y26899 , y26900 , y26901 , y26902 , y26903 , y26904 , y26905 , y26906 , y26907 , y26908 , y26909 , y26910 , y26911 , y26912 , y26913 , y26914 , y26915 , y26916 , y26917 , y26918 , y26919 , y26920 , y26921 , y26922 , y26923 , y26924 , y26925 , y26926 , y26927 , y26928 , y26929 , y26930 , y26931 , y26932 , y26933 , y26934 , y26935 , y26936 , y26937 , y26938 , y26939 , y26940 , y26941 , y26942 , y26943 , y26944 , y26945 , y26946 , y26947 , y26948 , y26949 , y26950 , y26951 , y26952 , y26953 , y26954 , y26955 , y26956 , y26957 , y26958 , y26959 , y26960 , y26961 , y26962 , y26963 , y26964 , y26965 , y26966 , y26967 , y26968 , y26969 , y26970 , y26971 , y26972 , y26973 , y26974 , y26975 , y26976 , y26977 , y26978 , y26979 , y26980 , y26981 , y26982 , y26983 , y26984 , y26985 , y26986 , y26987 , y26988 , y26989 , y26990 , y26991 , y26992 , y26993 , y26994 , y26995 , y26996 , y26997 , y26998 , y26999 , y27000 , y27001 , y27002 , y27003 , y27004 , y27005 , y27006 , y27007 , y27008 , y27009 , y27010 , y27011 , y27012 , y27013 , y27014 , y27015 , y27016 , y27017 , y27018 , y27019 , y27020 , y27021 , y27022 , y27023 , y27024 , y27025 , y27026 , y27027 , y27028 , y27029 , y27030 , y27031 , y27032 , y27033 , y27034 , y27035 , y27036 , y27037 , y27038 , y27039 , y27040 , y27041 , y27042 , y27043 , y27044 , y27045 , y27046 , y27047 , y27048 , y27049 , y27050 , y27051 , y27052 , y27053 , y27054 , y27055 , y27056 , y27057 , y27058 , y27059 , y27060 , y27061 , y27062 , y27063 , y27064 , y27065 , y27066 , y27067 , y27068 , y27069 , y27070 , y27071 , y27072 , y27073 , y27074 , y27075 , y27076 , y27077 , y27078 , y27079 , y27080 , y27081 , y27082 , y27083 , y27084 , y27085 , y27086 , y27087 , y27088 , y27089 , y27090 , y27091 , y27092 , y27093 , y27094 , y27095 , y27096 , y27097 , y27098 , y27099 , y27100 , y27101 , y27102 , y27103 , y27104 , y27105 , y27106 , y27107 , y27108 , y27109 , y27110 , y27111 , y27112 , y27113 , y27114 , y27115 , y27116 , y27117 , y27118 , y27119 , y27120 , y27121 , y27122 , y27123 , y27124 , y27125 , y27126 , y27127 , y27128 , y27129 , y27130 , y27131 , y27132 , y27133 , y27134 , y27135 , y27136 , y27137 , y27138 , y27139 , y27140 , y27141 , y27142 , y27143 , y27144 , y27145 , y27146 , y27147 , y27148 , y27149 , y27150 , y27151 , y27152 , y27153 , y27154 , y27155 , y27156 , y27157 , y27158 , y27159 , y27160 , y27161 , y27162 , y27163 , y27164 , y27165 , y27166 , y27167 , y27168 , y27169 , y27170 , y27171 , y27172 , y27173 , y27174 , y27175 , y27176 , y27177 , y27178 , y27179 , y27180 , y27181 , y27182 , y27183 , y27184 , y27185 , y27186 , y27187 , y27188 , y27189 , y27190 , y27191 , y27192 , y27193 , y27194 , y27195 , y27196 , y27197 , y27198 , y27199 , y27200 , y27201 , y27202 , y27203 , y27204 , y27205 , y27206 , y27207 , y27208 , y27209 , y27210 , y27211 , y27212 , y27213 , y27214 , y27215 , y27216 , y27217 , y27218 , y27219 , y27220 , y27221 , y27222 , y27223 , y27224 , y27225 , y27226 , y27227 , y27228 , y27229 , y27230 , y27231 , y27232 , y27233 , y27234 , y27235 , y27236 , y27237 , y27238 , y27239 , y27240 , y27241 , y27242 , y27243 , y27244 , y27245 , y27246 , y27247 , y27248 , y27249 , y27250 , y27251 , y27252 , y27253 , y27254 , y27255 , y27256 , y27257 , y27258 , y27259 , y27260 , y27261 , y27262 , y27263 , y27264 , y27265 , y27266 , y27267 , y27268 , y27269 , y27270 , y27271 , y27272 , y27273 , y27274 , y27275 , y27276 , y27277 , y27278 , y27279 , y27280 , y27281 , y27282 , y27283 , y27284 , y27285 , y27286 , y27287 , y27288 , y27289 , y27290 , y27291 , y27292 , y27293 , y27294 , y27295 , y27296 , y27297 , y27298 , y27299 , y27300 , y27301 , y27302 , y27303 , y27304 , y27305 , y27306 , y27307 , y27308 , y27309 , y27310 , y27311 , y27312 , y27313 , y27314 , y27315 , y27316 , y27317 , y27318 , y27319 , y27320 , y27321 , y27322 , y27323 , y27324 , y27325 , y27326 , y27327 , y27328 , y27329 , y27330 , y27331 , y27332 , y27333 , y27334 , y27335 , y27336 , y27337 , y27338 , y27339 , y27340 , y27341 , y27342 , y27343 , y27344 , y27345 , y27346 , y27347 , y27348 , y27349 , y27350 , y27351 , y27352 , y27353 , y27354 , y27355 , y27356 , y27357 , y27358 , y27359 , y27360 , y27361 , y27362 , y27363 , y27364 , y27365 , y27366 , y27367 , y27368 , y27369 , y27370 , y27371 , y27372 , y27373 , y27374 , y27375 , y27376 , y27377 , y27378 , y27379 , y27380 , y27381 , y27382 , y27383 , y27384 , y27385 , y27386 , y27387 , y27388 , y27389 , y27390 , y27391 , y27392 , y27393 , y27394 , y27395 , y27396 , y27397 , y27398 , y27399 , y27400 , y27401 , y27402 , y27403 , y27404 , y27405 , y27406 , y27407 , y27408 , y27409 , y27410 , y27411 , y27412 , y27413 , y27414 , y27415 , y27416 , y27417 , y27418 , y27419 , y27420 , y27421 , y27422 , y27423 , y27424 , y27425 , y27426 , y27427 , y27428 , y27429 , y27430 , y27431 , y27432 , y27433 , y27434 , y27435 , y27436 , y27437 , y27438 , y27439 , y27440 , y27441 , y27442 , y27443 , y27444 , y27445 , y27446 , y27447 , y27448 , y27449 , y27450 , y27451 , y27452 , y27453 , y27454 , y27455 , y27456 , y27457 , y27458 , y27459 , y27460 , y27461 , y27462 , y27463 , y27464 , y27465 , y27466 , y27467 , y27468 , y27469 , y27470 , y27471 , y27472 , y27473 , y27474 , y27475 , y27476 , y27477 , y27478 , y27479 , y27480 , y27481 , y27482 , y27483 , y27484 , y27485 , y27486 , y27487 , y27488 , y27489 , y27490 , y27491 , y27492 , y27493 , y27494 , y27495 , y27496 , y27497 , y27498 , y27499 , y27500 , y27501 , y27502 , y27503 , y27504 , y27505 , y27506 , y27507 , y27508 , y27509 , y27510 , y27511 , y27512 , y27513 , y27514 , y27515 , y27516 , y27517 , y27518 , y27519 , y27520 , y27521 , y27522 , y27523 , y27524 , y27525 , y27526 , y27527 , y27528 , y27529 , y27530 , y27531 , y27532 , y27533 , y27534 , y27535 , y27536 , y27537 , y27538 , y27539 , y27540 , y27541 , y27542 , y27543 , y27544 , y27545 , y27546 , y27547 , y27548 , y27549 , y27550 , y27551 , y27552 , y27553 , y27554 , y27555 , y27556 , y27557 , y27558 , y27559 , y27560 , y27561 , y27562 , y27563 , y27564 , y27565 , y27566 , y27567 , y27568 , y27569 , y27570 , y27571 , y27572 , y27573 , y27574 , y27575 , y27576 , y27577 , y27578 , y27579 , y27580 , y27581 , y27582 , y27583 , y27584 , y27585 , y27586 , y27587 , y27588 , y27589 , y27590 , y27591 , y27592 , y27593 , y27594 , y27595 , y27596 , y27597 , y27598 , y27599 , y27600 , y27601 , y27602 , y27603 , y27604 , y27605 , y27606 , y27607 , y27608 , y27609 , y27610 , y27611 , y27612 , y27613 , y27614 , y27615 , y27616 , y27617 , y27618 , y27619 , y27620 , y27621 , y27622 , y27623 , y27624 , y27625 , y27626 , y27627 , y27628 , y27629 , y27630 , y27631 , y27632 , y27633 , y27634 , y27635 , y27636 , y27637 , y27638 , y27639 , y27640 , y27641 , y27642 , y27643 , y27644 , y27645 , y27646 , y27647 , y27648 , y27649 , y27650 , y27651 , y27652 , y27653 , y27654 , y27655 , y27656 , y27657 , y27658 , y27659 , y27660 , y27661 , y27662 , y27663 , y27664 , y27665 , y27666 , y27667 , y27668 , y27669 , y27670 , y27671 , y27672 , y27673 , y27674 , y27675 , y27676 , y27677 , y27678 , y27679 , y27680 , y27681 , y27682 , y27683 , y27684 , y27685 , y27686 , y27687 , y27688 , y27689 , y27690 , y27691 , y27692 , y27693 , y27694 , y27695 , y27696 , y27697 , y27698 , y27699 , y27700 , y27701 , y27702 , y27703 , y27704 , y27705 , y27706 , y27707 , y27708 , y27709 , y27710 , y27711 , y27712 , y27713 , y27714 , y27715 , y27716 , y27717 , y27718 , y27719 , y27720 , y27721 , y27722 , y27723 , y27724 , y27725 , y27726 , y27727 , y27728 , y27729 , y27730 , y27731 , y27732 , y27733 , y27734 , y27735 , y27736 , y27737 , y27738 , y27739 , y27740 , y27741 , y27742 , y27743 , y27744 , y27745 , y27746 , y27747 , y27748 , y27749 , y27750 , y27751 , y27752 , y27753 , y27754 , y27755 , y27756 , y27757 , y27758 , y27759 , y27760 , y27761 , y27762 , y27763 , y27764 , y27765 , y27766 , y27767 , y27768 , y27769 , y27770 , y27771 , y27772 , y27773 , y27774 , y27775 , y27776 , y27777 , y27778 , y27779 , y27780 , y27781 , y27782 , y27783 , y27784 , y27785 , y27786 , y27787 , y27788 , y27789 , y27790 , y27791 , y27792 , y27793 , y27794 , y27795 , y27796 , y27797 , y27798 , y27799 , y27800 , y27801 , y27802 , y27803 , y27804 , y27805 , y27806 , y27807 , y27808 , y27809 , y27810 , y27811 , y27812 , y27813 , y27814 , y27815 , y27816 , y27817 , y27818 , y27819 , y27820 , y27821 , y27822 , y27823 , y27824 , y27825 , y27826 , y27827 , y27828 , y27829 , y27830 , y27831 , y27832 , y27833 , y27834 , y27835 , y27836 , y27837 , y27838 , y27839 , y27840 , y27841 , y27842 , y27843 , y27844 , y27845 , y27846 , y27847 , y27848 , y27849 , y27850 , y27851 , y27852 , y27853 , y27854 , y27855 , y27856 , y27857 , y27858 , y27859 , y27860 , y27861 , y27862 , y27863 , y27864 , y27865 , y27866 , y27867 , y27868 , y27869 , y27870 , y27871 , y27872 , y27873 , y27874 , y27875 , y27876 , y27877 , y27878 , y27879 , y27880 , y27881 , y27882 , y27883 , y27884 , y27885 , y27886 , y27887 , y27888 , y27889 , y27890 , y27891 , y27892 , y27893 , y27894 , y27895 , y27896 , y27897 , y27898 , y27899 , y27900 , y27901 , y27902 , y27903 , y27904 , y27905 , y27906 , y27907 , y27908 , y27909 , y27910 , y27911 , y27912 , y27913 , y27914 , y27915 , y27916 , y27917 , y27918 , y27919 , y27920 , y27921 , y27922 , y27923 , y27924 , y27925 , y27926 , y27927 , y27928 , y27929 , y27930 , y27931 , y27932 , y27933 , y27934 , y27935 , y27936 , y27937 , y27938 , y27939 , y27940 , y27941 , y27942 , y27943 , y27944 , y27945 , y27946 , y27947 , y27948 , y27949 , y27950 , y27951 , y27952 , y27953 , y27954 , y27955 , y27956 , y27957 , y27958 , y27959 , y27960 , y27961 , y27962 , y27963 , y27964 , y27965 , y27966 , y27967 , y27968 , y27969 , y27970 , y27971 , y27972 , y27973 , y27974 , y27975 , y27976 , y27977 , y27978 , y27979 , y27980 , y27981 , y27982 , y27983 , y27984 , y27985 , y27986 , y27987 , y27988 , y27989 , y27990 , y27991 , y27992 , y27993 , y27994 , y27995 , y27996 , y27997 , y27998 , y27999 , y28000 , y28001 , y28002 , y28003 , y28004 , y28005 , y28006 , y28007 , y28008 , y28009 , y28010 , y28011 , y28012 , y28013 , y28014 , y28015 , y28016 , y28017 , y28018 , y28019 , y28020 , y28021 , y28022 , y28023 , y28024 , y28025 , y28026 , y28027 , y28028 , y28029 , y28030 , y28031 , y28032 , y28033 , y28034 , y28035 , y28036 , y28037 , y28038 , y28039 , y28040 , y28041 , y28042 , y28043 , y28044 , y28045 , y28046 , y28047 , y28048 , y28049 , y28050 , y28051 , y28052 , y28053 , y28054 , y28055 , y28056 , y28057 , y28058 , y28059 , y28060 , y28061 , y28062 , y28063 , y28064 , y28065 , y28066 , y28067 , y28068 , y28069 , y28070 , y28071 , y28072 , y28073 , y28074 , y28075 , y28076 , y28077 , y28078 , y28079 , y28080 , y28081 , y28082 , y28083 , y28084 , y28085 , y28086 , y28087 , y28088 , y28089 , y28090 , y28091 , y28092 , y28093 , y28094 , y28095 , y28096 , y28097 , y28098 , y28099 , y28100 , y28101 , y28102 , y28103 , y28104 , y28105 , y28106 , y28107 , y28108 , y28109 , y28110 , y28111 , y28112 , y28113 , y28114 , y28115 , y28116 , y28117 , y28118 , y28119 , y28120 , y28121 , y28122 , y28123 , y28124 , y28125 , y28126 , y28127 , y28128 , y28129 , y28130 , y28131 , y28132 , y28133 , y28134 , y28135 , y28136 , y28137 , y28138 , y28139 , y28140 , y28141 , y28142 , y28143 , y28144 , y28145 , y28146 , y28147 , y28148 , y28149 , y28150 , y28151 , y28152 , y28153 , y28154 , y28155 , y28156 , y28157 , y28158 , y28159 , y28160 , y28161 , y28162 , y28163 , y28164 , y28165 , y28166 , y28167 , y28168 , y28169 , y28170 , y28171 , y28172 , y28173 , y28174 , y28175 , y28176 , y28177 , y28178 , y28179 , y28180 , y28181 , y28182 , y28183 , y28184 , y28185 , y28186 , y28187 , y28188 , y28189 , y28190 , y28191 , y28192 , y28193 , y28194 , y28195 , y28196 , y28197 , y28198 , y28199 , y28200 , y28201 , y28202 , y28203 , y28204 , y28205 , y28206 , y28207 , y28208 , y28209 , y28210 , y28211 , y28212 , y28213 , y28214 , y28215 , y28216 , y28217 , y28218 , y28219 , y28220 , y28221 , y28222 , y28223 , y28224 , y28225 , y28226 , y28227 , y28228 , y28229 , y28230 , y28231 , y28232 , y28233 , y28234 , y28235 , y28236 , y28237 , y28238 , y28239 , y28240 , y28241 , y28242 , y28243 , y28244 , y28245 , y28246 , y28247 , y28248 , y28249 , y28250 , y28251 , y28252 , y28253 , y28254 , y28255 , y28256 , y28257 , y28258 , y28259 , y28260 , y28261 , y28262 , y28263 , y28264 , y28265 , y28266 , y28267 , y28268 , y28269 , y28270 , y28271 , y28272 , y28273 , y28274 , y28275 , y28276 , y28277 , y28278 , y28279 , y28280 , y28281 , y28282 , y28283 , y28284 , y28285 , y28286 , y28287 , y28288 , y28289 , y28290 , y28291 , y28292 , y28293 , y28294 , y28295 , y28296 , y28297 , y28298 , y28299 , y28300 , y28301 , y28302 , y28303 , y28304 , y28305 , y28306 , y28307 , y28308 , y28309 , y28310 , y28311 , y28312 , y28313 , y28314 , y28315 , y28316 , y28317 , y28318 , y28319 , y28320 , y28321 , y28322 , y28323 , y28324 , y28325 , y28326 , y28327 , y28328 , y28329 , y28330 , y28331 , y28332 , y28333 , y28334 , y28335 , y28336 , y28337 , y28338 , y28339 , y28340 , y28341 , y28342 , y28343 , y28344 , y28345 , y28346 , y28347 , y28348 , y28349 , y28350 , y28351 , y28352 , y28353 , y28354 , y28355 , y28356 , y28357 , y28358 , y28359 , y28360 , y28361 , y28362 , y28363 , y28364 , y28365 , y28366 , y28367 , y28368 , y28369 , y28370 , y28371 , y28372 , y28373 , y28374 , y28375 , y28376 , y28377 , y28378 , y28379 , y28380 , y28381 , y28382 , y28383 , y28384 , y28385 , y28386 , y28387 , y28388 , y28389 , y28390 , y28391 , y28392 , y28393 , y28394 , y28395 , y28396 , y28397 , y28398 , y28399 , y28400 , y28401 , y28402 , y28403 , y28404 , y28405 , y28406 , y28407 , y28408 , y28409 , y28410 , y28411 , y28412 , y28413 , y28414 , y28415 , y28416 , y28417 , y28418 , y28419 , y28420 , y28421 , y28422 , y28423 , y28424 , y28425 , y28426 , y28427 , y28428 , y28429 , y28430 , y28431 , y28432 , y28433 , y28434 , y28435 , y28436 , y28437 , y28438 , y28439 , y28440 , y28441 , y28442 , y28443 , y28444 , y28445 , y28446 , y28447 , y28448 , y28449 , y28450 , y28451 , y28452 , y28453 , y28454 , y28455 , y28456 , y28457 , y28458 , y28459 , y28460 , y28461 , y28462 , y28463 , y28464 , y28465 , y28466 , y28467 , y28468 , y28469 , y28470 , y28471 , y28472 , y28473 , y28474 , y28475 , y28476 , y28477 , y28478 , y28479 , y28480 , y28481 , y28482 , y28483 , y28484 , y28485 , y28486 , y28487 , y28488 , y28489 , y28490 , y28491 , y28492 , y28493 , y28494 , y28495 , y28496 , y28497 , y28498 , y28499 , y28500 , y28501 , y28502 , y28503 , y28504 , y28505 , y28506 , y28507 , y28508 , y28509 , y28510 , y28511 , y28512 , y28513 , y28514 , y28515 , y28516 , y28517 , y28518 , y28519 , y28520 , y28521 , y28522 , y28523 , y28524 , y28525 , y28526 , y28527 , y28528 , y28529 , y28530 , y28531 , y28532 , y28533 , y28534 , y28535 , y28536 , y28537 , y28538 , y28539 , y28540 , y28541 , y28542 , y28543 , y28544 , y28545 , y28546 , y28547 , y28548 , y28549 , y28550 , y28551 , y28552 , y28553 , y28554 , y28555 , y28556 , y28557 , y28558 , y28559 , y28560 , y28561 , y28562 , y28563 , y28564 , y28565 , y28566 , y28567 , y28568 , y28569 , y28570 , y28571 , y28572 , y28573 , y28574 , y28575 , y28576 , y28577 , y28578 , y28579 , y28580 , y28581 , y28582 , y28583 , y28584 , y28585 , y28586 , y28587 , y28588 , y28589 , y28590 , y28591 , y28592 , y28593 , y28594 , y28595 , y28596 , y28597 , y28598 , y28599 , y28600 , y28601 , y28602 , y28603 , y28604 , y28605 , y28606 , y28607 , y28608 , y28609 , y28610 , y28611 , y28612 , y28613 , y28614 , y28615 , y28616 , y28617 , y28618 , y28619 , y28620 , y28621 , y28622 , y28623 , y28624 , y28625 , y28626 , y28627 , y28628 , y28629 , y28630 , y28631 , y28632 , y28633 , y28634 , y28635 , y28636 , y28637 , y28638 , y28639 , y28640 , y28641 , y28642 , y28643 , y28644 , y28645 , y28646 , y28647 , y28648 , y28649 , y28650 , y28651 , y28652 , y28653 , y28654 , y28655 , y28656 , y28657 , y28658 , y28659 , y28660 , y28661 , y28662 , y28663 , y28664 , y28665 , y28666 , y28667 , y28668 , y28669 , y28670 , y28671 , y28672 , y28673 , y28674 , y28675 , y28676 , y28677 , y28678 , y28679 , y28680 , y28681 , y28682 , y28683 , y28684 , y28685 , y28686 , y28687 , y28688 , y28689 , y28690 , y28691 , y28692 , y28693 , y28694 , y28695 , y28696 , y28697 , y28698 , y28699 , y28700 , y28701 , y28702 , y28703 , y28704 , y28705 , y28706 , y28707 , y28708 , y28709 , y28710 , y28711 , y28712 , y28713 , y28714 , y28715 , y28716 , y28717 , y28718 , y28719 , y28720 , y28721 , y28722 , y28723 , y28724 , y28725 , y28726 , y28727 , y28728 , y28729 , y28730 , y28731 , y28732 , y28733 , y28734 , y28735 , y28736 , y28737 , y28738 , y28739 , y28740 , y28741 , y28742 , y28743 , y28744 , y28745 , y28746 , y28747 , y28748 , y28749 , y28750 , y28751 , y28752 , y28753 , y28754 , y28755 , y28756 , y28757 , y28758 , y28759 , y28760 , y28761 , y28762 , y28763 , y28764 , y28765 , y28766 , y28767 , y28768 , y28769 , y28770 , y28771 , y28772 , y28773 , y28774 , y28775 , y28776 , y28777 , y28778 , y28779 , y28780 , y28781 , y28782 , y28783 , y28784 , y28785 , y28786 , y28787 , y28788 , y28789 , y28790 , y28791 , y28792 , y28793 , y28794 , y28795 , y28796 , y28797 , y28798 , y28799 , y28800 , y28801 , y28802 , y28803 , y28804 , y28805 , y28806 , y28807 , y28808 , y28809 , y28810 , y28811 , y28812 , y28813 , y28814 , y28815 , y28816 , y28817 , y28818 , y28819 , y28820 , y28821 , y28822 , y28823 , y28824 , y28825 , y28826 , y28827 , y28828 , y28829 , y28830 , y28831 , y28832 , y28833 , y28834 , y28835 , y28836 , y28837 , y28838 , y28839 , y28840 , y28841 , y28842 , y28843 , y28844 , y28845 , y28846 , y28847 , y28848 , y28849 , y28850 , y28851 , y28852 , y28853 , y28854 , y28855 , y28856 , y28857 , y28858 , y28859 , y28860 , y28861 , y28862 , y28863 , y28864 , y28865 , y28866 , y28867 , y28868 , y28869 , y28870 , y28871 , y28872 , y28873 , y28874 , y28875 , y28876 , y28877 , y28878 , y28879 , y28880 , y28881 , y28882 , y28883 , y28884 , y28885 , y28886 , y28887 , y28888 , y28889 , y28890 , y28891 , y28892 , y28893 , y28894 , y28895 , y28896 , y28897 , y28898 , y28899 , y28900 , y28901 , y28902 , y28903 , y28904 , y28905 , y28906 , y28907 , y28908 , y28909 , y28910 , y28911 , y28912 , y28913 , y28914 , y28915 , y28916 , y28917 , y28918 , y28919 , y28920 , y28921 , y28922 , y28923 , y28924 , y28925 , y28926 , y28927 , y28928 , y28929 , y28930 , y28931 , y28932 , y28933 , y28934 , y28935 , y28936 , y28937 , y28938 , y28939 , y28940 , y28941 , y28942 , y28943 , y28944 , y28945 , y28946 , y28947 , y28948 , y28949 , y28950 , y28951 , y28952 , y28953 , y28954 , y28955 , y28956 , y28957 , y28958 , y28959 , y28960 , y28961 , y28962 , y28963 , y28964 , y28965 , y28966 , y28967 , y28968 , y28969 , y28970 , y28971 , y28972 , y28973 , y28974 , y28975 , y28976 , y28977 , y28978 , y28979 , y28980 , y28981 , y28982 , y28983 , y28984 , y28985 , y28986 , y28987 , y28988 , y28989 , y28990 , y28991 , y28992 , y28993 , y28994 , y28995 , y28996 , y28997 , y28998 , y28999 , y29000 , y29001 , y29002 , y29003 , y29004 , y29005 , y29006 , y29007 , y29008 , y29009 , y29010 , y29011 , y29012 , y29013 , y29014 , y29015 , y29016 , y29017 , y29018 , y29019 , y29020 , y29021 , y29022 , y29023 , y29024 , y29025 , y29026 , y29027 , y29028 , y29029 , y29030 , y29031 , y29032 , y29033 , y29034 , y29035 , y29036 , y29037 , y29038 , y29039 , y29040 , y29041 , y29042 , y29043 , y29044 , y29045 , y29046 , y29047 , y29048 , y29049 , y29050 , y29051 , y29052 , y29053 , y29054 , y29055 , y29056 , y29057 , y29058 , y29059 , y29060 , y29061 , y29062 , y29063 , y29064 , y29065 , y29066 , y29067 , y29068 , y29069 , y29070 , y29071 , y29072 , y29073 , y29074 , y29075 , y29076 , y29077 , y29078 , y29079 , y29080 , y29081 , y29082 , y29083 , y29084 , y29085 , y29086 , y29087 , y29088 , y29089 , y29090 , y29091 , y29092 , y29093 , y29094 , y29095 , y29096 , y29097 , y29098 , y29099 , y29100 , y29101 , y29102 , y29103 , y29104 , y29105 , y29106 , y29107 , y29108 , y29109 , y29110 , y29111 , y29112 , y29113 , y29114 , y29115 , y29116 , y29117 , y29118 , y29119 , y29120 , y29121 , y29122 , y29123 , y29124 , y29125 , y29126 , y29127 , y29128 , y29129 , y29130 , y29131 , y29132 , y29133 , y29134 , y29135 , y29136 , y29137 , y29138 , y29139 , y29140 , y29141 , y29142 , y29143 , y29144 , y29145 , y29146 , y29147 , y29148 , y29149 , y29150 , y29151 , y29152 , y29153 , y29154 , y29155 , y29156 , y29157 , y29158 , y29159 , y29160 , y29161 , y29162 , y29163 , y29164 , y29165 , y29166 , y29167 , y29168 , y29169 , y29170 , y29171 , y29172 , y29173 , y29174 , y29175 , y29176 , y29177 , y29178 , y29179 , y29180 , y29181 , y29182 , y29183 , y29184 , y29185 , y29186 , y29187 , y29188 , y29189 , y29190 , y29191 , y29192 , y29193 , y29194 , y29195 , y29196 , y29197 , y29198 , y29199 , y29200 , y29201 , y29202 , y29203 , y29204 , y29205 , y29206 , y29207 , y29208 , y29209 , y29210 , y29211 , y29212 , y29213 , y29214 , y29215 , y29216 , y29217 , y29218 , y29219 , y29220 , y29221 , y29222 , y29223 , y29224 , y29225 , y29226 , y29227 , y29228 , y29229 , y29230 , y29231 , y29232 , y29233 , y29234 , y29235 , y29236 , y29237 , y29238 , y29239 , y29240 , y29241 , y29242 , y29243 , y29244 , y29245 , y29246 , y29247 , y29248 , y29249 , y29250 , y29251 , y29252 , y29253 , y29254 , y29255 , y29256 , y29257 , y29258 , y29259 , y29260 , y29261 , y29262 , y29263 , y29264 , y29265 , y29266 , y29267 , y29268 , y29269 , y29270 , y29271 , y29272 , y29273 , y29274 , y29275 , y29276 , y29277 , y29278 , y29279 , y29280 , y29281 , y29282 , y29283 , y29284 , y29285 , y29286 , y29287 , y29288 , y29289 , y29290 , y29291 , y29292 , y29293 , y29294 , y29295 , y29296 , y29297 , y29298 , y29299 , y29300 , y29301 , y29302 , y29303 , y29304 , y29305 , y29306 , y29307 , y29308 , y29309 , y29310 , y29311 , y29312 , y29313 , y29314 , y29315 , y29316 , y29317 , y29318 , y29319 , y29320 , y29321 , y29322 , y29323 , y29324 , y29325 , y29326 , y29327 , y29328 , y29329 , y29330 , y29331 , y29332 , y29333 , y29334 , y29335 , y29336 , y29337 , y29338 , y29339 , y29340 , y29341 , y29342 , y29343 , y29344 , y29345 , y29346 , y29347 , y29348 , y29349 , y29350 , y29351 , y29352 , y29353 , y29354 , y29355 , y29356 , y29357 , y29358 , y29359 , y29360 , y29361 , y29362 , y29363 , y29364 , y29365 , y29366 , y29367 , y29368 , y29369 , y29370 , y29371 , y29372 , y29373 , y29374 , y29375 , y29376 , y29377 , y29378 , y29379 , y29380 , y29381 , y29382 , y29383 , y29384 , y29385 , y29386 , y29387 , y29388 , y29389 , y29390 , y29391 , y29392 , y29393 , y29394 , y29395 , y29396 , y29397 , y29398 , y29399 , y29400 , y29401 , y29402 , y29403 , y29404 , y29405 , y29406 , y29407 , y29408 , y29409 , y29410 , y29411 , y29412 , y29413 , y29414 , y29415 , y29416 , y29417 , y29418 , y29419 , y29420 , y29421 , y29422 , y29423 , y29424 , y29425 , y29426 , y29427 , y29428 , y29429 , y29430 , y29431 , y29432 , y29433 , y29434 , y29435 , y29436 , y29437 , y29438 , y29439 , y29440 , y29441 , y29442 , y29443 , y29444 , y29445 , y29446 , y29447 , y29448 , y29449 , y29450 , y29451 , y29452 , y29453 , y29454 , y29455 , y29456 , y29457 , y29458 , y29459 , y29460 , y29461 , y29462 , y29463 , y29464 , y29465 , y29466 , y29467 , y29468 , y29469 , y29470 , y29471 , y29472 , y29473 , y29474 , y29475 , y29476 , y29477 , y29478 , y29479 , y29480 , y29481 , y29482 , y29483 , y29484 , y29485 , y29486 , y29487 , y29488 , y29489 , y29490 , y29491 , y29492 , y29493 , y29494 , y29495 , y29496 , y29497 , y29498 , y29499 , y29500 , y29501 , y29502 , y29503 , y29504 , y29505 , y29506 , y29507 , y29508 , y29509 , y29510 , y29511 , y29512 , y29513 , y29514 , y29515 , y29516 , y29517 , y29518 , y29519 , y29520 , y29521 , y29522 , y29523 , y29524 , y29525 , y29526 , y29527 , y29528 , y29529 , y29530 , y29531 , y29532 , y29533 , y29534 , y29535 , y29536 , y29537 , y29538 , y29539 , y29540 , y29541 , y29542 , y29543 , y29544 , y29545 , y29546 , y29547 , y29548 , y29549 , y29550 , y29551 , y29552 , y29553 , y29554 , y29555 , y29556 , y29557 , y29558 , y29559 , y29560 , y29561 , y29562 , y29563 , y29564 , y29565 , y29566 , y29567 , y29568 , y29569 , y29570 , y29571 , y29572 , y29573 , y29574 , y29575 , y29576 , y29577 , y29578 , y29579 , y29580 , y29581 , y29582 , y29583 , y29584 , y29585 , y29586 , y29587 , y29588 , y29589 , y29590 , y29591 , y29592 , y29593 , y29594 , y29595 , y29596 , y29597 , y29598 , y29599 , y29600 , y29601 , y29602 , y29603 , y29604 , y29605 , y29606 , y29607 , y29608 , y29609 , y29610 , y29611 , y29612 , y29613 , y29614 , y29615 , y29616 , y29617 , y29618 , y29619 , y29620 , y29621 , y29622 , y29623 , y29624 , y29625 , y29626 , y29627 , y29628 , y29629 , y29630 , y29631 , y29632 , y29633 , y29634 , y29635 , y29636 , y29637 , y29638 , y29639 , y29640 , y29641 , y29642 , y29643 , y29644 , y29645 , y29646 , y29647 , y29648 , y29649 , y29650 , y29651 , y29652 , y29653 , y29654 , y29655 , y29656 , y29657 , y29658 , y29659 , y29660 , y29661 , y29662 , y29663 , y29664 , y29665 , y29666 , y29667 , y29668 , y29669 , y29670 , y29671 , y29672 , y29673 , y29674 , y29675 , y29676 , y29677 , y29678 , y29679 , y29680 , y29681 , y29682 , y29683 , y29684 , y29685 , y29686 , y29687 , y29688 , y29689 , y29690 , y29691 , y29692 , y29693 , y29694 , y29695 , y29696 , y29697 , y29698 , y29699 , y29700 , y29701 , y29702 , y29703 , y29704 , y29705 , y29706 , y29707 , y29708 , y29709 , y29710 , y29711 , y29712 , y29713 , y29714 , y29715 , y29716 , y29717 , y29718 , y29719 , y29720 , y29721 , y29722 , y29723 , y29724 , y29725 , y29726 , y29727 , y29728 , y29729 , y29730 , y29731 , y29732 , y29733 , y29734 , y29735 , y29736 , y29737 , y29738 , y29739 , y29740 , y29741 , y29742 , y29743 , y29744 , y29745 , y29746 , y29747 , y29748 , y29749 , y29750 , y29751 , y29752 , y29753 , y29754 , y29755 , y29756 , y29757 , y29758 , y29759 , y29760 , y29761 , y29762 , y29763 , y29764 , y29765 , y29766 , y29767 , y29768 , y29769 , y29770 , y29771 , y29772 , y29773 , y29774 , y29775 , y29776 , y29777 , y29778 , y29779 , y29780 , y29781 , y29782 , y29783 , y29784 , y29785 , y29786 , y29787 , y29788 , y29789 , y29790 , y29791 , y29792 , y29793 , y29794 , y29795 , y29796 , y29797 , y29798 , y29799 , y29800 , y29801 , y29802 , y29803 , y29804 , y29805 , y29806 , y29807 , y29808 , y29809 , y29810 , y29811 , y29812 , y29813 , y29814 , y29815 , y29816 , y29817 , y29818 , y29819 , y29820 , y29821 , y29822 , y29823 , y29824 , y29825 , y29826 , y29827 , y29828 , y29829 , y29830 , y29831 , y29832 , y29833 , y29834 , y29835 , y29836 , y29837 , y29838 , y29839 , y29840 , y29841 , y29842 , y29843 , y29844 , y29845 , y29846 , y29847 , y29848 , y29849 , y29850 , y29851 , y29852 , y29853 , y29854 , y29855 , y29856 , y29857 , y29858 , y29859 , y29860 , y29861 , y29862 , y29863 , y29864 , y29865 , y29866 , y29867 , y29868 , y29869 , y29870 , y29871 , y29872 , y29873 , y29874 , y29875 , y29876 , y29877 , y29878 , y29879 , y29880 , y29881 , y29882 , y29883 , y29884 , y29885 , y29886 , y29887 , y29888 , y29889 , y29890 , y29891 , y29892 , y29893 , y29894 , y29895 , y29896 , y29897 , y29898 , y29899 , y29900 , y29901 , y29902 , y29903 , y29904 , y29905 , y29906 , y29907 , y29908 , y29909 , y29910 , y29911 , y29912 , y29913 , y29914 , y29915 , y29916 , y29917 , y29918 , y29919 , y29920 , y29921 , y29922 , y29923 , y29924 , y29925 , y29926 , y29927 , y29928 , y29929 , y29930 , y29931 , y29932 , y29933 , y29934 , y29935 , y29936 , y29937 , y29938 , y29939 , y29940 , y29941 , y29942 , y29943 , y29944 , y29945 , y29946 , y29947 , y29948 , y29949 , y29950 , y29951 , y29952 , y29953 , y29954 , y29955 , y29956 , y29957 , y29958 , y29959 , y29960 , y29961 , y29962 , y29963 , y29964 , y29965 , y29966 , y29967 , y29968 , y29969 , y29970 , y29971 , y29972 , y29973 , y29974 , y29975 , y29976 , y29977 , y29978 , y29979 , y29980 , y29981 , y29982 , y29983 , y29984 , y29985 , y29986 , y29987 , y29988 , y29989 , y29990 , y29991 , y29992 , y29993 , y29994 , y29995 , y29996 , y29997 , y29998 , y29999 , y30000 , y30001 , y30002 , y30003 , y30004 , y30005 , y30006 , y30007 , y30008 , y30009 , y30010 , y30011 , y30012 , y30013 , y30014 , y30015 , y30016 , y30017 , y30018 , y30019 , y30020 , y30021 , y30022 , y30023 , y30024 , y30025 , y30026 , y30027 , y30028 , y30029 , y30030 , y30031 , y30032 , y30033 , y30034 , y30035 , y30036 , y30037 , y30038 , y30039 , y30040 , y30041 , y30042 , y30043 , y30044 , y30045 , y30046 , y30047 , y30048 , y30049 , y30050 , y30051 , y30052 , y30053 , y30054 , y30055 , y30056 , y30057 , y30058 , y30059 , y30060 , y30061 , y30062 , y30063 , y30064 , y30065 , y30066 , y30067 , y30068 , y30069 , y30070 , y30071 , y30072 , y30073 , y30074 , y30075 , y30076 , y30077 , y30078 , y30079 , y30080 , y30081 , y30082 , y30083 , y30084 , y30085 , y30086 , y30087 , y30088 , y30089 , y30090 , y30091 , y30092 , y30093 , y30094 , y30095 , y30096 , y30097 , y30098 , y30099 , y30100 , y30101 , y30102 , y30103 , y30104 , y30105 , y30106 , y30107 , y30108 , y30109 , y30110 , y30111 , y30112 , y30113 , y30114 , y30115 , y30116 , y30117 , y30118 , y30119 , y30120 , y30121 , y30122 , y30123 , y30124 , y30125 , y30126 , y30127 , y30128 , y30129 , y30130 , y30131 , y30132 , y30133 , y30134 , y30135 , y30136 , y30137 , y30138 , y30139 , y30140 , y30141 , y30142 , y30143 , y30144 , y30145 , y30146 , y30147 , y30148 , y30149 , y30150 , y30151 , y30152 , y30153 , y30154 , y30155 , y30156 , y30157 , y30158 , y30159 , y30160 , y30161 , y30162 , y30163 , y30164 , y30165 , y30166 , y30167 , y30168 , y30169 , y30170 , y30171 , y30172 , y30173 , y30174 , y30175 , y30176 , y30177 , y30178 , y30179 , y30180 , y30181 , y30182 , y30183 , y30184 , y30185 , y30186 , y30187 , y30188 , y30189 , y30190 , y30191 , y30192 , y30193 , y30194 , y30195 , y30196 , y30197 , y30198 , y30199 , y30200 , y30201 , y30202 , y30203 , y30204 , y30205 , y30206 , y30207 , y30208 , y30209 , y30210 , y30211 , y30212 , y30213 , y30214 , y30215 , y30216 , y30217 , y30218 , y30219 , y30220 , y30221 , y30222 , y30223 , y30224 , y30225 , y30226 , y30227 , y30228 , y30229 , y30230 , y30231 , y30232 , y30233 , y30234 , y30235 , y30236 , y30237 , y30238 , y30239 , y30240 , y30241 , y30242 , y30243 , y30244 , y30245 , y30246 , y30247 , y30248 , y30249 , y30250 , y30251 , y30252 , y30253 , y30254 , y30255 , y30256 , y30257 , y30258 , y30259 , y30260 , y30261 , y30262 , y30263 , y30264 , y30265 , y30266 , y30267 , y30268 , y30269 , y30270 , y30271 , y30272 , y30273 , y30274 , y30275 , y30276 , y30277 , y30278 , y30279 , y30280 , y30281 , y30282 , y30283 , y30284 , y30285 , y30286 , y30287 , y30288 , y30289 , y30290 , y30291 , y30292 , y30293 , y30294 , y30295 , y30296 , y30297 , y30298 , y30299 , y30300 , y30301 , y30302 , y30303 , y30304 , y30305 , y30306 , y30307 , y30308 , y30309 , y30310 , y30311 , y30312 , y30313 , y30314 , y30315 , y30316 , y30317 , y30318 , y30319 , y30320 , y30321 , y30322 , y30323 , y30324 , y30325 , y30326 , y30327 , y30328 , y30329 , y30330 , y30331 , y30332 , y30333 , y30334 , y30335 , y30336 , y30337 , y30338 , y30339 , y30340 , y30341 , y30342 , y30343 , y30344 , y30345 , y30346 , y30347 , y30348 , y30349 , y30350 , y30351 , y30352 , y30353 , y30354 , y30355 , y30356 , y30357 , y30358 , y30359 , y30360 , y30361 , y30362 , y30363 , y30364 , y30365 , y30366 , y30367 , y30368 , y30369 , y30370 , y30371 , y30372 , y30373 , y30374 , y30375 , y30376 , y30377 , y30378 , y30379 , y30380 , y30381 , y30382 , y30383 , y30384 , y30385 , y30386 , y30387 , y30388 , y30389 , y30390 , y30391 , y30392 , y30393 , y30394 , y30395 , y30396 , y30397 , y30398 , y30399 , y30400 , y30401 , y30402 , y30403 , y30404 , y30405 , y30406 , y30407 , y30408 , y30409 , y30410 , y30411 , y30412 , y30413 , y30414 , y30415 , y30416 , y30417 , y30418 , y30419 , y30420 , y30421 , y30422 , y30423 , y30424 , y30425 , y30426 , y30427 , y30428 , y30429 , y30430 , y30431 , y30432 , y30433 , y30434 , y30435 , y30436 , y30437 , y30438 , y30439 , y30440 , y30441 , y30442 , y30443 , y30444 , y30445 , y30446 , y30447 , y30448 , y30449 , y30450 , y30451 , y30452 , y30453 , y30454 , y30455 , y30456 , y30457 , y30458 , y30459 , y30460 , y30461 , y30462 , y30463 , y30464 , y30465 , y30466 , y30467 , y30468 , y30469 , y30470 , y30471 , y30472 , y30473 , y30474 , y30475 , y30476 , y30477 , y30478 , y30479 , y30480 , y30481 , y30482 , y30483 , y30484 , y30485 , y30486 , y30487 , y30488 , y30489 , y30490 , y30491 , y30492 , y30493 , y30494 , y30495 , y30496 , y30497 , y30498 , y30499 , y30500 , y30501 , y30502 , y30503 , y30504 , y30505 , y30506 , y30507 , y30508 , y30509 , y30510 , y30511 , y30512 , y30513 , y30514 , y30515 , y30516 , y30517 , y30518 , y30519 , y30520 , y30521 , y30522 , y30523 , y30524 , y30525 , y30526 , y30527 , y30528 , y30529 , y30530 , y30531 , y30532 , y30533 , y30534 , y30535 , y30536 , y30537 , y30538 , y30539 , y30540 , y30541 , y30542 , y30543 , y30544 , y30545 , y30546 , y30547 , y30548 , y30549 , y30550 , y30551 , y30552 , y30553 , y30554 , y30555 , y30556 , y30557 , y30558 , y30559 , y30560 , y30561 , y30562 , y30563 , y30564 , y30565 , y30566 , y30567 , y30568 , y30569 , y30570 , y30571 , y30572 , y30573 , y30574 , y30575 , y30576 , y30577 , y30578 , y30579 , y30580 , y30581 , y30582 , y30583 , y30584 , y30585 , y30586 , y30587 , y30588 , y30589 , y30590 , y30591 , y30592 , y30593 , y30594 , y30595 , y30596 , y30597 , y30598 , y30599 , y30600 , y30601 , y30602 , y30603 , y30604 , y30605 , y30606 , y30607 , y30608 , y30609 , y30610 , y30611 , y30612 , y30613 , y30614 , y30615 , y30616 , y30617 , y30618 , y30619 , y30620 , y30621 , y30622 , y30623 , y30624 , y30625 , y30626 , y30627 , y30628 , y30629 , y30630 , y30631 , y30632 , y30633 , y30634 , y30635 , y30636 , y30637 , y30638 , y30639 , y30640 , y30641 , y30642 , y30643 , y30644 , y30645 , y30646 , y30647 , y30648 , y30649 , y30650 , y30651 , y30652 , y30653 , y30654 , y30655 , y30656 , y30657 , y30658 , y30659 , y30660 , y30661 , y30662 , y30663 , y30664 , y30665 , y30666 , y30667 , y30668 , y30669 , y30670 , y30671 , y30672 , y30673 , y30674 , y30675 , y30676 , y30677 , y30678 , y30679 , y30680 , y30681 , y30682 , y30683 , y30684 , y30685 , y30686 , y30687 , y30688 , y30689 , y30690 , y30691 , y30692 , y30693 , y30694 , y30695 , y30696 , y30697 , y30698 , y30699 , y30700 , y30701 , y30702 , y30703 , y30704 , y30705 , y30706 , y30707 , y30708 , y30709 , y30710 , y30711 , y30712 , y30713 , y30714 , y30715 , y30716 , y30717 , y30718 , y30719 , y30720 , y30721 , y30722 , y30723 , y30724 , y30725 , y30726 , y30727 , y30728 , y30729 , y30730 , y30731 , y30732 , y30733 , y30734 , y30735 , y30736 , y30737 , y30738 , y30739 , y30740 , y30741 , y30742 , y30743 , y30744 , y30745 , y30746 , y30747 , y30748 , y30749 , y30750 , y30751 , y30752 , y30753 , y30754 , y30755 , y30756 , y30757 , y30758 , y30759 , y30760 , y30761 , y30762 , y30763 , y30764 , y30765 , y30766 , y30767 , y30768 , y30769 , y30770 , y30771 , y30772 , y30773 , y30774 , y30775 , y30776 , y30777 , y30778 , y30779 , y30780 , y30781 , y30782 , y30783 , y30784 , y30785 , y30786 , y30787 , y30788 , y30789 , y30790 , y30791 , y30792 , y30793 , y30794 , y30795 , y30796 , y30797 , y30798 , y30799 , y30800 , y30801 , y30802 , y30803 , y30804 , y30805 , y30806 , y30807 , y30808 , y30809 , y30810 , y30811 , y30812 , y30813 , y30814 , y30815 , y30816 , y30817 , y30818 , y30819 , y30820 , y30821 , y30822 , y30823 , y30824 , y30825 , y30826 , y30827 , y30828 , y30829 , y30830 , y30831 , y30832 , y30833 , y30834 , y30835 , y30836 , y30837 , y30838 , y30839 , y30840 , y30841 , y30842 , y30843 , y30844 , y30845 , y30846 , y30847 , y30848 , y30849 , y30850 , y30851 , y30852 , y30853 , y30854 , y30855 , y30856 , y30857 , y30858 , y30859 , y30860 , y30861 , y30862 , y30863 , y30864 , y30865 , y30866 , y30867 , y30868 , y30869 , y30870 , y30871 , y30872 , y30873 , y30874 , y30875 , y30876 , y30877 , y30878 , y30879 , y30880 , y30881 , y30882 , y30883 , y30884 , y30885 , y30886 , y30887 , y30888 , y30889 , y30890 , y30891 , y30892 , y30893 , y30894 , y30895 , y30896 , y30897 , y30898 , y30899 , y30900 , y30901 , y30902 , y30903 , y30904 , y30905 , y30906 , y30907 , y30908 , y30909 , y30910 , y30911 , y30912 , y30913 , y30914 , y30915 , y30916 , y30917 , y30918 , y30919 , y30920 , y30921 , y30922 , y30923 , y30924 , y30925 , y30926 , y30927 , y30928 , y30929 , y30930 , y30931 , y30932 , y30933 , y30934 , y30935 , y30936 , y30937 , y30938 , y30939 , y30940 , y30941 , y30942 , y30943 , y30944 , y30945 , y30946 , y30947 , y30948 , y30949 , y30950 , y30951 , y30952 , y30953 , y30954 , y30955 , y30956 , y30957 , y30958 , y30959 , y30960 , y30961 , y30962 , y30963 , y30964 , y30965 , y30966 , y30967 , y30968 , y30969 , y30970 , y30971 , y30972 , y30973 , y30974 , y30975 , y30976 , y30977 , y30978 , y30979 , y30980 , y30981 , y30982 , y30983 , y30984 , y30985 , y30986 , y30987 , y30988 , y30989 , y30990 , y30991 , y30992 , y30993 , y30994 , y30995 , y30996 , y30997 , y30998 , y30999 , y31000 , y31001 , y31002 , y31003 , y31004 , y31005 , y31006 , y31007 , y31008 , y31009 , y31010 , y31011 , y31012 , y31013 , y31014 , y31015 , y31016 , y31017 , y31018 , y31019 , y31020 , y31021 , y31022 , y31023 , y31024 , y31025 , y31026 , y31027 , y31028 , y31029 , y31030 , y31031 , y31032 , y31033 , y31034 , y31035 , y31036 , y31037 , y31038 , y31039 , y31040 , y31041 , y31042 , y31043 , y31044 , y31045 , y31046 , y31047 , y31048 , y31049 , y31050 , y31051 , y31052 , y31053 , y31054 , y31055 , y31056 , y31057 , y31058 , y31059 , y31060 , y31061 , y31062 , y31063 , y31064 , y31065 , y31066 , y31067 , y31068 , y31069 , y31070 , y31071 , y31072 , y31073 , y31074 , y31075 , y31076 , y31077 , y31078 , y31079 , y31080 , y31081 , y31082 , y31083 , y31084 , y31085 , y31086 , y31087 , y31088 , y31089 , y31090 , y31091 , y31092 , y31093 , y31094 , y31095 , y31096 , y31097 , y31098 , y31099 , y31100 , y31101 , y31102 , y31103 , y31104 , y31105 , y31106 , y31107 , y31108 , y31109 , y31110 , y31111 , y31112 , y31113 , y31114 , y31115 , y31116 , y31117 , y31118 , y31119 , y31120 , y31121 , y31122 , y31123 , y31124 , y31125 , y31126 , y31127 , y31128 , y31129 , y31130 , y31131 , y31132 , y31133 , y31134 , y31135 , y31136 , y31137 , y31138 , y31139 , y31140 , y31141 , y31142 , y31143 , y31144 , y31145 , y31146 , y31147 , y31148 , y31149 , y31150 , y31151 , y31152 , y31153 , y31154 , y31155 , y31156 , y31157 , y31158 , y31159 , y31160 , y31161 , y31162 , y31163 , y31164 , y31165 , y31166 , y31167 , y31168 , y31169 , y31170 , y31171 , y31172 , y31173 , y31174 , y31175 , y31176 , y31177 , y31178 , y31179 , y31180 , y31181 , y31182 , y31183 , y31184 , y31185 , y31186 , y31187 , y31188 , y31189 , y31190 , y31191 , y31192 , y31193 , y31194 , y31195 , y31196 , y31197 , y31198 , y31199 , y31200 , y31201 , y31202 , y31203 , y31204 , y31205 , y31206 , y31207 , y31208 , y31209 , y31210 , y31211 , y31212 , y31213 , y31214 , y31215 , y31216 , y31217 , y31218 , y31219 , y31220 , y31221 , y31222 , y31223 , y31224 , y31225 , y31226 , y31227 , y31228 , y31229 , y31230 , y31231 , y31232 , y31233 , y31234 , y31235 , y31236 , y31237 , y31238 , y31239 , y31240 , y31241 , y31242 , y31243 , y31244 , y31245 , y31246 , y31247 , y31248 , y31249 , y31250 , y31251 , y31252 , y31253 , y31254 , y31255 , y31256 , y31257 , y31258 , y31259 , y31260 , y31261 , y31262 , y31263 , y31264 , y31265 , y31266 , y31267 , y31268 , y31269 , y31270 , y31271 , y31272 , y31273 , y31274 , y31275 , y31276 , y31277 , y31278 , y31279 , y31280 , y31281 , y31282 , y31283 , y31284 , y31285 , y31286 , y31287 , y31288 , y31289 , y31290 , y31291 , y31292 , y31293 , y31294 , y31295 , y31296 , y31297 , y31298 , y31299 , y31300 , y31301 , y31302 , y31303 , y31304 , y31305 , y31306 , y31307 , y31308 , y31309 , y31310 , y31311 , y31312 , y31313 , y31314 , y31315 , y31316 , y31317 , y31318 , y31319 , y31320 , y31321 , y31322 , y31323 , y31324 , y31325 , y31326 , y31327 , y31328 , y31329 , y31330 , y31331 , y31332 , y31333 , y31334 , y31335 , y31336 , y31337 , y31338 , y31339 , y31340 , y31341 , y31342 , y31343 , y31344 , y31345 , y31346 , y31347 , y31348 , y31349 , y31350 , y31351 , y31352 , y31353 , y31354 , y31355 , y31356 , y31357 , y31358 , y31359 , y31360 , y31361 , y31362 , y31363 , y31364 , y31365 , y31366 , y31367 , y31368 , y31369 , y31370 , y31371 , y31372 , y31373 , y31374 , y31375 , y31376 , y31377 , y31378 , y31379 , y31380 , y31381 , y31382 , y31383 , y31384 , y31385 , y31386 , y31387 , y31388 , y31389 , y31390 , y31391 , y31392 , y31393 , y31394 , y31395 , y31396 , y31397 , y31398 , y31399 , y31400 , y31401 , y31402 , y31403 , y31404 , y31405 , y31406 , y31407 , y31408 , y31409 , y31410 , y31411 , y31412 , y31413 , y31414 , y31415 , y31416 , y31417 , y31418 , y31419 , y31420 , y31421 , y31422 , y31423 , y31424 , y31425 , y31426 , y31427 , y31428 , y31429 , y31430 , y31431 , y31432 , y31433 , y31434 , y31435 , y31436 , y31437 , y31438 , y31439 , y31440 , y31441 , y31442 , y31443 , y31444 , y31445 , y31446 , y31447 , y31448 , y31449 , y31450 , y31451 , y31452 , y31453 , y31454 , y31455 , y31456 , y31457 , y31458 , y31459 , y31460 , y31461 , y31462 , y31463 , y31464 , y31465 , y31466 , y31467 , y31468 , y31469 , y31470 , y31471 , y31472 , y31473 , y31474 , y31475 , y31476 , y31477 , y31478 , y31479 , y31480 , y31481 , y31482 , y31483 , y31484 , y31485 , y31486 , y31487 , y31488 , y31489 , y31490 , y31491 , y31492 , y31493 , y31494 , y31495 , y31496 , y31497 , y31498 , y31499 , y31500 , y31501 , y31502 , y31503 , y31504 , y31505 , y31506 , y31507 , y31508 , y31509 , y31510 , y31511 , y31512 , y31513 , y31514 , y31515 , y31516 , y31517 , y31518 , y31519 , y31520 , y31521 , y31522 , y31523 , y31524 , y31525 , y31526 , y31527 , y31528 , y31529 , y31530 , y31531 , y31532 , y31533 , y31534 , y31535 , y31536 , y31537 , y31538 , y31539 , y31540 , y31541 , y31542 , y31543 , y31544 , y31545 , y31546 , y31547 , y31548 , y31549 , y31550 , y31551 , y31552 , y31553 , y31554 , y31555 , y31556 , y31557 , y31558 , y31559 , y31560 , y31561 , y31562 , y31563 , y31564 , y31565 , y31566 , y31567 , y31568 , y31569 , y31570 , y31571 , y31572 , y31573 , y31574 , y31575 , y31576 , y31577 , y31578 , y31579 , y31580 , y31581 , y31582 , y31583 , y31584 , y31585 , y31586 , y31587 , y31588 , y31589 , y31590 , y31591 , y31592 , y31593 , y31594 , y31595 , y31596 , y31597 , y31598 , y31599 , y31600 , y31601 , y31602 , y31603 , y31604 , y31605 , y31606 , y31607 , y31608 , y31609 , y31610 , y31611 , y31612 , y31613 , y31614 , y31615 , y31616 , y31617 , y31618 , y31619 , y31620 , y31621 , y31622 , y31623 , y31624 , y31625 , y31626 , y31627 , y31628 , y31629 , y31630 , y31631 , y31632 , y31633 , y31634 , y31635 , y31636 , y31637 , y31638 , y31639 , y31640 , y31641 , y31642 , y31643 , y31644 , y31645 , y31646 , y31647 , y31648 , y31649 , y31650 , y31651 , y31652 , y31653 , y31654 , y31655 , y31656 , y31657 , y31658 , y31659 , y31660 , y31661 , y31662 , y31663 , y31664 , y31665 , y31666 , y31667 , y31668 , y31669 , y31670 , y31671 , y31672 , y31673 , y31674 , y31675 , y31676 , y31677 , y31678 , y31679 , y31680 , y31681 , y31682 , y31683 , y31684 , y31685 , y31686 , y31687 , y31688 , y31689 , y31690 , y31691 , y31692 , y31693 , y31694 , y31695 , y31696 , y31697 , y31698 , y31699 , y31700 , y31701 , y31702 , y31703 , y31704 , y31705 , y31706 , y31707 , y31708 , y31709 , y31710 , y31711 , y31712 , y31713 , y31714 , y31715 , y31716 , y31717 , y31718 , y31719 , y31720 , y31721 , y31722 , y31723 , y31724 , y31725 , y31726 , y31727 , y31728 , y31729 , y31730 , y31731 , y31732 , y31733 , y31734 , y31735 , y31736 , y31737 , y31738 , y31739 , y31740 , y31741 , y31742 , y31743 , y31744 , y31745 , y31746 , y31747 , y31748 , y31749 , y31750 , y31751 , y31752 , y31753 , y31754 , y31755 , y31756 , y31757 , y31758 , y31759 , y31760 , y31761 , y31762 , y31763 , y31764 , y31765 , y31766 , y31767 , y31768 , y31769 , y31770 , y31771 , y31772 , y31773 , y31774 , y31775 , y31776 , y31777 , y31778 , y31779 , y31780 , y31781 , y31782 , y31783 , y31784 , y31785 , y31786 , y31787 , y31788 , y31789 , y31790 , y31791 , y31792 , y31793 , y31794 , y31795 , y31796 , y31797 , y31798 , y31799 , y31800 , y31801 , y31802 , y31803 , y31804 , y31805 , y31806 , y31807 , y31808 , y31809 , y31810 , y31811 , y31812 , y31813 , y31814 , y31815 , y31816 , y31817 , y31818 , y31819 , y31820 , y31821 , y31822 , y31823 , y31824 , y31825 , y31826 , y31827 , y31828 , y31829 , y31830 , y31831 , y31832 , y31833 , y31834 , y31835 , y31836 , y31837 , y31838 , y31839 , y31840 , y31841 , y31842 , y31843 , y31844 , y31845 , y31846 , y31847 , y31848 , y31849 , y31850 , y31851 , y31852 , y31853 , y31854 , y31855 , y31856 , y31857 , y31858 , y31859 , y31860 , y31861 , y31862 , y31863 , y31864 , y31865 , y31866 , y31867 , y31868 , y31869 , y31870 , y31871 , y31872 , y31873 , y31874 , y31875 , y31876 , y31877 , y31878 , y31879 , y31880 , y31881 , y31882 , y31883 , y31884 , y31885 , y31886 , y31887 , y31888 , y31889 , y31890 , y31891 , y31892 , y31893 , y31894 , y31895 , y31896 , y31897 , y31898 , y31899 , y31900 , y31901 , y31902 , y31903 , y31904 , y31905 , y31906 , y31907 , y31908 , y31909 , y31910 , y31911 , y31912 , y31913 , y31914 , y31915 , y31916 , y31917 , y31918 , y31919 , y31920 , y31921 , y31922 , y31923 , y31924 , y31925 , y31926 , y31927 , y31928 , y31929 , y31930 , y31931 , y31932 , y31933 , y31934 , y31935 , y31936 , y31937 , y31938 , y31939 , y31940 , y31941 , y31942 , y31943 , y31944 , y31945 , y31946 , y31947 , y31948 , y31949 , y31950 , y31951 , y31952 , y31953 , y31954 , y31955 , y31956 , y31957 , y31958 , y31959 , y31960 , y31961 , y31962 , y31963 , y31964 , y31965 , y31966 , y31967 , y31968 , y31969 , y31970 , y31971 , y31972 , y31973 , y31974 , y31975 , y31976 , y31977 , y31978 , y31979 , y31980 , y31981 , y31982 , y31983 , y31984 , y31985 , y31986 , y31987 , y31988 , y31989 , y31990 , y31991 , y31992 , y31993 , y31994 , y31995 , y31996 , y31997 , y31998 , y31999 , y32000 , y32001 , y32002 , y32003 , y32004 , y32005 , y32006 , y32007 , y32008 , y32009 , y32010 , y32011 , y32012 , y32013 , y32014 , y32015 , y32016 , y32017 , y32018 , y32019 , y32020 , y32021 , y32022 , y32023 , y32024 , y32025 , y32026 , y32027 , y32028 , y32029 , y32030 , y32031 , y32032 , y32033 , y32034 ;
  wire n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , n18511 , n18512 , n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , n18679 , n18680 , n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , n18709 , n18710 , n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , n18841 , n18842 , n18843 , n18844 , n18845 , n18846 , n18847 , n18848 , n18849 , n18850 , n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , n18870 , n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , n18891 , n18892 , n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , n18910 , n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , n18921 , n18922 , n18923 , n18924 , n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , n18969 , n18970 , n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , n18977 , n18978 , n18979 , n18980 , n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , n18989 , n18990 , n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , n18999 , n19000 , n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , n19017 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , n19029 , n19030 , n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , n19037 , n19038 , n19039 , n19040 , n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , n19049 , n19050 , n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , n19060 , n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , n19067 , n19068 , n19069 , n19070 , n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , n19079 , n19080 , n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , n19089 , n19090 , n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , n19099 , n19100 , n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , n19137 , n19138 , n19139 , n19140 , n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , n19157 , n19158 , n19159 , n19160 , n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , n19167 , n19168 , n19169 , n19170 , n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , n19179 , n19180 , n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , n19189 , n19190 , n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , n19198 , n19199 , n19200 , n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , n19210 , n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , n19217 , n19218 , n19219 , n19220 , n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , n19229 , n19230 , n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , n19239 , n19240 , n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , n19249 , n19250 , n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , n19259 , n19260 , n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , n19279 , n19280 , n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , n19287 , n19288 , n19289 , n19290 , n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , n19297 , n19298 , n19299 , n19300 , n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , n19309 , n19310 , n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , n19319 , n19320 , n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , n19329 , n19330 , n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , n19339 , n19340 , n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , n19359 , n19360 , n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , n19369 , n19370 , n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , n19379 , n19380 , n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19387 , n19388 , n19389 , n19390 , n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , n19400 , n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , n19410 , n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , n19417 , n19418 , n19419 , n19420 , n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , n19440 , n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , n19450 , n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , n19459 , n19460 , n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , n19470 , n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , n19529 , n19530 , n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , n19550 , n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , n19567 , n19568 , n19569 , n19570 , n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , n19587 , n19588 , n19589 , n19590 , n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , n19619 , n19620 , n19621 , n19622 , n19623 , n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , n19670 , n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , n19711 , n19712 , n19713 , n19714 , n19715 , n19716 , n19717 , n19718 , n19719 , n19720 , n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , n19737 , n19738 , n19739 , n19740 , n19741 , n19742 , n19743 , n19744 , n19745 , n19746 , n19747 , n19748 , n19749 , n19750 , n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , n19757 , n19758 , n19759 , n19760 , n19761 , n19762 , n19763 , n19764 , n19765 , n19766 , n19767 , n19768 , n19769 , n19770 , n19771 , n19772 , n19773 , n19774 , n19775 , n19776 , n19777 , n19778 , n19779 , n19780 , n19781 , n19782 , n19783 , n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , n19791 , n19792 , n19793 , n19794 , n19795 , n19796 , n19797 , n19798 , n19799 , n19800 , n19801 , n19802 , n19803 , n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , n19811 , n19812 , n19813 , n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , n19821 , n19822 , n19823 , n19824 , n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , n19831 , n19832 , n19833 , n19834 , n19835 , n19836 , n19837 , n19838 , n19839 , n19840 , n19841 , n19842 , n19843 , n19844 , n19845 , n19846 , n19847 , n19848 , n19849 , n19850 , n19851 , n19852 , n19853 , n19854 , n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , n19861 , n19862 , n19863 , n19864 , n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , n19871 , n19872 , n19873 , n19874 , n19875 , n19876 , n19877 , n19878 , n19879 , n19880 , n19881 , n19882 , n19883 , n19884 , n19885 , n19886 , n19887 , n19888 , n19889 , n19890 , n19891 , n19892 , n19893 , n19894 , n19895 , n19896 , n19897 , n19898 , n19899 , n19900 , n19901 , n19902 , n19903 , n19904 , n19905 , n19906 , n19907 , n19908 , n19909 , n19910 , n19911 , n19912 , n19913 , n19914 , n19915 , n19916 , n19917 , n19918 , n19919 , n19920 , n19921 , n19922 , n19923 , n19924 , n19925 , n19926 , n19927 , n19928 , n19929 , n19930 , n19931 , n19932 , n19933 , n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , n19940 , n19941 , n19942 , n19943 , n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , n19951 , n19952 , n19953 , n19954 , n19955 , n19956 , n19957 , n19958 , n19959 , n19960 , n19961 , n19962 , n19963 , n19964 , n19965 , n19966 , n19967 , n19968 , n19969 , n19970 , n19971 , n19972 , n19973 , n19974 , n19975 , n19976 , n19977 , n19978 , n19979 , n19980 , n19981 , n19982 , n19983 , n19984 , n19985 , n19986 , n19987 , n19988 , n19989 , n19990 , n19991 , n19992 , n19993 , n19994 , n19995 , n19996 , n19997 , n19998 , n19999 , n20000 , n20001 , n20002 , n20003 , n20004 , n20005 , n20006 , n20007 , n20008 , n20009 , n20010 , n20011 , n20012 , n20013 , n20014 , n20015 , n20016 , n20017 , n20018 , n20019 , n20020 , n20021 , n20022 , n20023 , n20024 , n20025 , n20026 , n20027 , n20028 , n20029 , n20030 , n20031 , n20032 , n20033 , n20034 , n20035 , n20036 , n20037 , n20038 , n20039 , n20040 , n20041 , n20042 , n20043 , n20044 , n20045 , n20046 , n20047 , n20048 , n20049 , n20050 , n20051 , n20052 , n20053 , n20054 , n20055 , n20056 , n20057 , n20058 , n20059 , n20060 , n20061 , n20062 , n20063 , n20064 , n20065 , n20066 , n20067 , n20068 , n20069 , n20070 , n20071 , n20072 , n20073 , n20074 , n20075 , n20076 , n20077 , n20078 , n20079 , n20080 , n20081 , n20082 , n20083 , n20084 , n20085 , n20086 , n20087 , n20088 , n20089 , n20090 , n20091 , n20092 , n20093 , n20094 , n20095 , n20096 , n20097 , n20098 , n20099 , n20100 , n20101 , n20102 , n20103 , n20104 , n20105 , n20106 , n20107 , n20108 , n20109 , n20110 , n20111 , n20112 , n20113 , n20114 , n20115 , n20116 , n20117 , n20118 , n20119 , n20120 , n20121 , n20122 , n20123 , n20124 , n20125 , n20126 , n20127 , n20128 , n20129 , n20130 , n20131 , n20132 , n20133 , n20134 , n20135 , n20136 , n20137 , n20138 , n20139 , n20140 , n20141 , n20142 , n20143 , n20144 , n20145 , n20146 , n20147 , n20148 , n20149 , n20150 , n20151 , n20152 , n20153 , n20154 , n20155 , n20156 , n20157 , n20158 , n20159 , n20160 , n20161 , n20162 , n20163 , n20164 , n20165 , n20166 , n20167 , n20168 , n20169 , n20170 , n20171 , n20172 , n20173 , n20174 , n20175 , n20176 , n20177 , n20178 , n20179 , n20180 , n20181 , n20182 , n20183 , n20184 , n20185 , n20186 , n20187 , n20188 , n20189 , n20190 , n20191 , n20192 , n20193 , n20194 , n20195 , n20196 , n20197 , n20198 , n20199 , n20200 , n20201 , n20202 , n20203 , n20204 , n20205 , n20206 , n20207 , n20208 , n20209 , n20210 , n20211 , n20212 , n20213 , n20214 , n20215 , n20216 , n20217 , n20218 , n20219 , n20220 , n20221 , n20222 , n20223 , n20224 , n20225 , n20226 , n20227 , n20228 , n20229 , n20230 , n20231 , n20232 , n20233 , n20234 , n20235 , n20236 , n20237 , n20238 , n20239 , n20240 , n20241 , n20242 , n20243 , n20244 , n20245 , n20246 , n20247 , n20248 , n20249 , n20250 , n20251 , n20252 , n20253 , n20254 , n20255 , n20256 , n20257 , n20258 , n20259 , n20260 , n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , n20267 , n20268 , n20269 , n20270 , n20271 , n20272 , n20273 , n20274 , n20275 , n20276 , n20277 , n20278 , n20279 , n20280 , n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , n20287 , n20288 , n20289 , n20290 , n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , n20297 , n20298 , n20299 , n20300 , n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , n20307 , n20308 , n20309 , n20310 , n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , n20317 , n20318 , n20319 , n20320 , n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , n20327 , n20328 , n20329 , n20330 , n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , n20337 , n20338 , n20339 , n20340 , n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , n20347 , n20348 , n20349 , n20350 , n20351 , n20352 , n20353 , n20354 , n20355 , n20356 , n20357 , n20358 , n20359 , n20360 , n20361 , n20362 , n20363 , n20364 , n20365 , n20366 , n20367 , n20368 , n20369 , n20370 , n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , n20377 , n20378 , n20379 , n20380 , n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , n20389 , n20390 , n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , n20397 , n20398 , n20399 , n20400 , n20401 , n20402 , n20403 , n20404 , n20405 , n20406 , n20407 , n20408 , n20409 , n20410 , n20411 , n20412 , n20413 , n20414 , n20415 , n20416 , n20417 , n20418 , n20419 , n20420 , n20421 , n20422 , n20423 , n20424 , n20425 , n20426 , n20427 , n20428 , n20429 , n20430 , n20431 , n20432 , n20433 , n20434 , n20435 , n20436 , n20437 , n20438 , n20439 , n20440 , n20441 , n20442 , n20443 , n20444 , n20445 , n20446 , n20447 , n20448 , n20449 , n20450 , n20451 , n20452 , n20453 , n20454 , n20455 , n20456 , n20457 , n20458 , n20459 , n20460 , n20461 , n20462 , n20463 , n20464 , n20465 , n20466 , n20467 , n20468 , n20469 , n20470 , n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , n20477 , n20478 , n20479 , n20480 , n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , n20487 , n20488 , n20489 , n20490 , n20491 , n20492 , n20493 , n20494 , n20495 , n20496 , n20497 , n20498 , n20499 , n20500 , n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , n20507 , n20508 , n20509 , n20510 , n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , n20519 , n20520 , n20521 , n20522 , n20523 , n20524 , n20525 , n20526 , n20527 , n20528 , n20529 , n20530 , n20531 , n20532 , n20533 , n20534 , n20535 , n20536 , n20537 , n20538 , n20539 , n20540 , n20541 , n20542 , n20543 , n20544 , n20545 , n20546 , n20547 , n20548 , n20549 , n20550 , n20551 , n20552 , n20553 , n20554 , n20555 , n20556 , n20557 , n20558 , n20559 , n20560 , n20561 , n20562 , n20563 , n20564 , n20565 , n20566 , n20567 , n20568 , n20569 , n20570 , n20571 , n20572 , n20573 , n20574 , n20575 , n20576 , n20577 , n20578 , n20579 , n20580 , n20581 , n20582 , n20583 , n20584 , n20585 , n20586 , n20587 , n20588 , n20589 , n20590 , n20591 , n20592 , n20593 , n20594 , n20595 , n20596 , n20597 , n20598 , n20599 , n20600 , n20601 , n20602 , n20603 , n20604 , n20605 , n20606 , n20607 , n20608 , n20609 , n20610 , n20611 , n20612 , n20613 , n20614 , n20615 , n20616 , n20617 , n20618 , n20619 , n20620 , n20621 , n20622 , n20623 , n20624 , n20625 , n20626 , n20627 , n20628 , n20629 , n20630 , n20631 , n20632 , n20633 , n20634 , n20635 , n20636 , n20637 , n20638 , n20639 , n20640 , n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , n20647 , n20648 , n20649 , n20650 , n20651 , n20652 , n20653 , n20654 , n20655 , n20656 , n20657 , n20658 , n20659 , n20660 , n20661 , n20662 , n20663 , n20664 , n20665 , n20666 , n20667 , n20668 , n20669 , n20670 , n20671 , n20672 , n20673 , n20674 , n20675 , n20676 , n20677 , n20678 , n20679 , n20680 , n20681 , n20682 , n20683 , n20684 , n20685 , n20686 , n20687 , n20688 , n20689 , n20690 , n20691 , n20692 , n20693 , n20694 , n20695 , n20696 , n20697 , n20698 , n20699 , n20700 , n20701 , n20702 , n20703 , n20704 , n20705 , n20706 , n20707 , n20708 , n20709 , n20710 , n20711 , n20712 , n20713 , n20714 , n20715 , n20716 , n20717 , n20718 , n20719 , n20720 , n20721 , n20722 , n20723 , n20724 , n20725 , n20726 , n20727 , n20728 , n20729 , n20730 , n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , n20737 , n20738 , n20739 , n20740 , n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , n20747 , n20748 , n20749 , n20750 , n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , n20757 , n20758 , n20759 , n20760 , n20761 , n20762 , n20763 , n20764 , n20765 , n20766 , n20767 , n20768 , n20769 , n20770 , n20771 , n20772 , n20773 , n20774 , n20775 , n20776 , n20777 , n20778 , n20779 , n20780 , n20781 , n20782 , n20783 , n20784 , n20785 , n20786 , n20787 , n20788 , n20789 , n20790 , n20791 , n20792 , n20793 , n20794 , n20795 , n20796 , n20797 , n20798 , n20799 , n20800 , n20801 , n20802 , n20803 , n20804 , n20805 , n20806 , n20807 , n20808 , n20809 , n20810 , n20811 , n20812 , n20813 , n20814 , n20815 , n20816 , n20817 , n20818 , n20819 , n20820 , n20821 , n20822 , n20823 , n20824 , n20825 , n20826 , n20827 , n20828 , n20829 , n20830 , n20831 , n20832 , n20833 , n20834 , n20835 , n20836 , n20837 , n20838 , n20839 , n20840 , n20841 , n20842 , n20843 , n20844 , n20845 , n20846 , n20847 , n20848 , n20849 , n20850 , n20851 , n20852 , n20853 , n20854 , n20855 , n20856 , n20857 , n20858 , n20859 , n20860 , n20861 , n20862 , n20863 , n20864 , n20865 , n20866 , n20867 , n20868 , n20869 , n20870 , n20871 , n20872 , n20873 , n20874 , n20875 , n20876 , n20877 , n20878 , n20879 , n20880 , n20881 , n20882 , n20883 , n20884 , n20885 , n20886 , n20887 , n20888 , n20889 , n20890 , n20891 , n20892 , n20893 , n20894 , n20895 , n20896 , n20897 , n20898 , n20899 , n20900 , n20901 , n20902 , n20903 , n20904 , n20905 , n20906 , n20907 , n20908 , n20909 , n20910 , n20911 , n20912 , n20913 , n20914 , n20915 , n20916 , n20917 , n20918 , n20919 , n20920 , n20921 , n20922 , n20923 , n20924 , n20925 , n20926 , n20927 , n20928 , n20929 , n20930 , n20931 , n20932 , n20933 , n20934 , n20935 , n20936 , n20937 , n20938 , n20939 , n20940 , n20941 , n20942 , n20943 , n20944 , n20945 , n20946 , n20947 , n20948 , n20949 , n20950 , n20951 , n20952 , n20953 , n20954 , n20955 , n20956 , n20957 , n20958 , n20959 , n20960 , n20961 , n20962 , n20963 , n20964 , n20965 , n20966 , n20967 , n20968 , n20969 , n20970 , n20971 , n20972 , n20973 , n20974 , n20975 , n20976 , n20977 , n20978 , n20979 , n20980 , n20981 , n20982 , n20983 , n20984 , n20985 , n20986 , n20987 , n20988 , n20989 , n20990 , n20991 , n20992 , n20993 , n20994 , n20995 , n20996 , n20997 , n20998 , n20999 , n21000 , n21001 , n21002 , n21003 , n21004 , n21005 , n21006 , n21007 , n21008 , n21009 , n21010 , n21011 , n21012 , n21013 , n21014 , n21015 , n21016 , n21017 , n21018 , n21019 , n21020 , n21021 , n21022 , n21023 , n21024 , n21025 , n21026 , n21027 , n21028 , n21029 , n21030 , n21031 , n21032 , n21033 , n21034 , n21035 , n21036 , n21037 , n21038 , n21039 , n21040 , n21041 , n21042 , n21043 , n21044 , n21045 , n21046 , n21047 , n21048 , n21049 , n21050 , n21051 , n21052 , n21053 , n21054 , n21055 , n21056 , n21057 , n21058 , n21059 , n21060 , n21061 , n21062 , n21063 , n21064 , n21065 , n21066 , n21067 , n21068 , n21069 , n21070 , n21071 , n21072 , n21073 , n21074 , n21075 , n21076 , n21077 , n21078 , n21079 , n21080 , n21081 , n21082 , n21083 , n21084 , n21085 , n21086 , n21087 , n21088 , n21089 , n21090 , n21091 , n21092 , n21093 , n21094 , n21095 , n21096 , n21097 , n21098 , n21099 , n21100 , n21101 , n21102 , n21103 , n21104 , n21105 , n21106 , n21107 , n21108 , n21109 , n21110 , n21111 , n21112 , n21113 , n21114 , n21115 , n21116 , n21117 , n21118 , n21119 , n21120 , n21121 , n21122 , n21123 , n21124 , n21125 , n21126 , n21127 , n21128 , n21129 , n21130 , n21131 , n21132 , n21133 , n21134 , n21135 , n21136 , n21137 , n21138 , n21139 , n21140 , n21141 , n21142 , n21143 , n21144 , n21145 , n21146 , n21147 , n21148 , n21149 , n21150 , n21151 , n21152 , n21153 , n21154 , n21155 , n21156 , n21157 , n21158 , n21159 , n21160 , n21161 , n21162 , n21163 , n21164 , n21165 , n21166 , n21167 , n21168 , n21169 , n21170 , n21171 , n21172 , n21173 , n21174 , n21175 , n21176 , n21177 , n21178 , n21179 , n21180 , n21181 , n21182 , n21183 , n21184 , n21185 , n21186 , n21187 , n21188 , n21189 , n21190 , n21191 , n21192 , n21193 , n21194 , n21195 , n21196 , n21197 , n21198 , n21199 , n21200 , n21201 , n21202 , n21203 , n21204 , n21205 , n21206 , n21207 , n21208 , n21209 , n21210 , n21211 , n21212 , n21213 , n21214 , n21215 , n21216 , n21217 , n21218 , n21219 , n21220 , n21221 , n21222 , n21223 , n21224 , n21225 , n21226 , n21227 , n21228 , n21229 , n21230 , n21231 , n21232 , n21233 , n21234 , n21235 , n21236 , n21237 , n21238 , n21239 , n21240 , n21241 , n21242 , n21243 , n21244 , n21245 , n21246 , n21247 , n21248 , n21249 , n21250 , n21251 , n21252 , n21253 , n21254 , n21255 , n21256 , n21257 , n21258 , n21259 , n21260 , n21261 , n21262 , n21263 , n21264 , n21265 , n21266 , n21267 , n21268 , n21269 , n21270 , n21271 , n21272 , n21273 , n21274 , n21275 , n21276 , n21277 , n21278 , n21279 , n21280 , n21281 , n21282 , n21283 , n21284 , n21285 , n21286 , n21287 , n21288 , n21289 , n21290 , n21291 , n21292 , n21293 , n21294 , n21295 , n21296 , n21297 , n21298 , n21299 , n21300 , n21301 , n21302 , n21303 , n21304 , n21305 , n21306 , n21307 , n21308 , n21309 , n21310 , n21311 , n21312 , n21313 , n21314 , n21315 , n21316 , n21317 , n21318 , n21319 , n21320 , n21321 , n21322 , n21323 , n21324 , n21325 , n21326 , n21327 , n21328 , n21329 , n21330 , n21331 , n21332 , n21333 , n21334 , n21335 , n21336 , n21337 , n21338 , n21339 , n21340 , n21341 , n21342 , n21343 , n21344 , n21345 , n21346 , n21347 , n21348 , n21349 , n21350 , n21351 , n21352 , n21353 , n21354 , n21355 , n21356 , n21357 , n21358 , n21359 , n21360 , n21361 , n21362 , n21363 , n21364 , n21365 , n21366 , n21367 , n21368 , n21369 , n21370 , n21371 , n21372 , n21373 , n21374 , n21375 , n21376 , n21377 , n21378 , n21379 , n21380 , n21381 , n21382 , n21383 , n21384 , n21385 , n21386 , n21387 , n21388 , n21389 , n21390 , n21391 , n21392 , n21393 , n21394 , n21395 , n21396 , n21397 , n21398 , n21399 , n21400 , n21401 , n21402 , n21403 , n21404 , n21405 , n21406 , n21407 , n21408 , n21409 , n21410 , n21411 , n21412 , n21413 , n21414 , n21415 , n21416 , n21417 , n21418 , n21419 , n21420 , n21421 , n21422 , n21423 , n21424 , n21425 , n21426 , n21427 , n21428 , n21429 , n21430 , n21431 , n21432 , n21433 , n21434 , n21435 , n21436 , n21437 , n21438 , n21439 , n21440 , n21441 , n21442 , n21443 , n21444 , n21445 , n21446 , n21447 , n21448 , n21449 , n21450 , n21451 , n21452 , n21453 , n21454 , n21455 , n21456 , n21457 , n21458 , n21459 , n21460 , n21461 , n21462 , n21463 , n21464 , n21465 , n21466 , n21467 , n21468 , n21469 , n21470 , n21471 , n21472 , n21473 , n21474 , n21475 , n21476 , n21477 , n21478 , n21479 , n21480 , n21481 , n21482 , n21483 , n21484 , n21485 , n21486 , n21487 , n21488 , n21489 , n21490 , n21491 , n21492 , n21493 , n21494 , n21495 , n21496 , n21497 , n21498 , n21499 , n21500 , n21501 , n21502 , n21503 , n21504 , n21505 , n21506 , n21507 , n21508 , n21509 , n21510 , n21511 , n21512 , n21513 , n21514 , n21515 , n21516 , n21517 , n21518 , n21519 , n21520 , n21521 , n21522 , n21523 , n21524 , n21525 , n21526 , n21527 , n21528 , n21529 , n21530 , n21531 , n21532 , n21533 , n21534 , n21535 , n21536 , n21537 , n21538 , n21539 , n21540 , n21541 , n21542 , n21543 , n21544 , n21545 , n21546 , n21547 , n21548 , n21549 , n21550 , n21551 , n21552 , n21553 , n21554 , n21555 , n21556 , n21557 , n21558 , n21559 , n21560 , n21561 , n21562 , n21563 , n21564 , n21565 , n21566 , n21567 , n21568 , n21569 , n21570 , n21571 , n21572 , n21573 , n21574 , n21575 , n21576 , n21577 , n21578 , n21579 , n21580 , n21581 , n21582 , n21583 , n21584 , n21585 , n21586 , n21587 , n21588 , n21589 , n21590 , n21591 , n21592 , n21593 , n21594 , n21595 , n21596 , n21597 , n21598 , n21599 , n21600 , n21601 , n21602 , n21603 , n21604 , n21605 , n21606 , n21607 , n21608 , n21609 , n21610 , n21611 , n21612 , n21613 , n21614 , n21615 , n21616 , n21617 , n21618 , n21619 , n21620 , n21621 , n21622 , n21623 , n21624 , n21625 , n21626 , n21627 , n21628 , n21629 , n21630 , n21631 , n21632 , n21633 , n21634 , n21635 , n21636 , n21637 , n21638 , n21639 , n21640 , n21641 , n21642 , n21643 , n21644 , n21645 , n21646 , n21647 , n21648 , n21649 , n21650 , n21651 , n21652 , n21653 , n21654 , n21655 , n21656 , n21657 , n21658 , n21659 , n21660 , n21661 , n21662 , n21663 , n21664 , n21665 , n21666 , n21667 , n21668 , n21669 , n21670 , n21671 , n21672 , n21673 , n21674 , n21675 , n21676 , n21677 , n21678 , n21679 , n21680 , n21681 , n21682 , n21683 , n21684 , n21685 , n21686 , n21687 , n21688 , n21689 , n21690 , n21691 , n21692 , n21693 , n21694 , n21695 , n21696 , n21697 , n21698 , n21699 , n21700 , n21701 , n21702 , n21703 , n21704 , n21705 , n21706 , n21707 , n21708 , n21709 , n21710 , n21711 , n21712 , n21713 , n21714 , n21715 , n21716 , n21717 , n21718 , n21719 , n21720 , n21721 , n21722 , n21723 , n21724 , n21725 , n21726 , n21727 , n21728 , n21729 , n21730 , n21731 , n21732 , n21733 , n21734 , n21735 , n21736 , n21737 , n21738 , n21739 , n21740 , n21741 , n21742 , n21743 , n21744 , n21745 , n21746 , n21747 , n21748 , n21749 , n21750 , n21751 , n21752 , n21753 , n21754 , n21755 , n21756 , n21757 , n21758 , n21759 , n21760 , n21761 , n21762 , n21763 , n21764 , n21765 , n21766 , n21767 , n21768 , n21769 , n21770 , n21771 , n21772 , n21773 , n21774 , n21775 , n21776 , n21777 , n21778 , n21779 , n21780 , n21781 , n21782 , n21783 , n21784 , n21785 , n21786 , n21787 , n21788 , n21789 , n21790 , n21791 , n21792 , n21793 , n21794 , n21795 , n21796 , n21797 , n21798 , n21799 , n21800 , n21801 , n21802 , n21803 , n21804 , n21805 , n21806 , n21807 , n21808 , n21809 , n21810 , n21811 , n21812 , n21813 , n21814 , n21815 , n21816 , n21817 , n21818 , n21819 , n21820 , n21821 , n21822 , n21823 , n21824 , n21825 , n21826 , n21827 , n21828 , n21829 , n21830 , n21831 , n21832 , n21833 , n21834 , n21835 , n21836 , n21837 , n21838 , n21839 , n21840 , n21841 , n21842 , n21843 , n21844 , n21845 , n21846 , n21847 , n21848 , n21849 , n21850 , n21851 , n21852 , n21853 , n21854 , n21855 , n21856 , n21857 , n21858 , n21859 , n21860 , n21861 , n21862 , n21863 , n21864 , n21865 , n21866 , n21867 , n21868 , n21869 , n21870 , n21871 , n21872 , n21873 , n21874 , n21875 , n21876 , n21877 , n21878 , n21879 , n21880 , n21881 , n21882 , n21883 , n21884 , n21885 , n21886 , n21887 , n21888 , n21889 , n21890 , n21891 , n21892 , n21893 , n21894 , n21895 , n21896 , n21897 , n21898 , n21899 , n21900 , n21901 , n21902 , n21903 , n21904 , n21905 , n21906 , n21907 , n21908 , n21909 , n21910 , n21911 , n21912 , n21913 , n21914 , n21915 , n21916 , n21917 , n21918 , n21919 , n21920 , n21921 , n21922 , n21923 , n21924 , n21925 , n21926 , n21927 , n21928 , n21929 , n21930 , n21931 , n21932 , n21933 , n21934 , n21935 , n21936 , n21937 , n21938 , n21939 , n21940 , n21941 , n21942 , n21943 , n21944 , n21945 , n21946 , n21947 , n21948 , n21949 , n21950 , n21951 , n21952 , n21953 , n21954 , n21955 , n21956 , n21957 , n21958 , n21959 , n21960 , n21961 , n21962 , n21963 , n21964 , n21965 , n21966 , n21967 , n21968 , n21969 , n21970 , n21971 , n21972 , n21973 , n21974 , n21975 , n21976 , n21977 , n21978 , n21979 , n21980 , n21981 , n21982 , n21983 , n21984 , n21985 , n21986 , n21987 , n21988 , n21989 , n21990 , n21991 , n21992 , n21993 , n21994 , n21995 , n21996 , n21997 , n21998 , n21999 , n22000 , n22001 , n22002 , n22003 , n22004 , n22005 , n22006 , n22007 , n22008 , n22009 , n22010 , n22011 , n22012 , n22013 , n22014 , n22015 , n22016 , n22017 , n22018 , n22019 , n22020 , n22021 , n22022 , n22023 , n22024 , n22025 , n22026 , n22027 , n22028 , n22029 , n22030 , n22031 , n22032 , n22033 , n22034 , n22035 , n22036 , n22037 , n22038 , n22039 , n22040 , n22041 , n22042 , n22043 , n22044 , n22045 , n22046 , n22047 , n22048 , n22049 , n22050 , n22051 , n22052 , n22053 , n22054 , n22055 , n22056 , n22057 , n22058 , n22059 , n22060 , n22061 , n22062 , n22063 , n22064 , n22065 , n22066 , n22067 , n22068 , n22069 , n22070 , n22071 , n22072 , n22073 , n22074 , n22075 , n22076 , n22077 , n22078 , n22079 , n22080 , n22081 , n22082 , n22083 , n22084 , n22085 , n22086 , n22087 , n22088 , n22089 , n22090 , n22091 , n22092 , n22093 , n22094 , n22095 , n22096 , n22097 , n22098 , n22099 , n22100 , n22101 , n22102 , n22103 , n22104 , n22105 , n22106 , n22107 , n22108 , n22109 , n22110 , n22111 , n22112 , n22113 , n22114 , n22115 , n22116 , n22117 , n22118 , n22119 , n22120 , n22121 , n22122 , n22123 , n22124 , n22125 , n22126 , n22127 , n22128 , n22129 , n22130 , n22131 , n22132 , n22133 , n22134 , n22135 , n22136 , n22137 , n22138 , n22139 , n22140 , n22141 , n22142 , n22143 , n22144 , n22145 , n22146 , n22147 , n22148 , n22149 , n22150 , n22151 , n22152 , n22153 , n22154 , n22155 , n22156 , n22157 , n22158 , n22159 , n22160 , n22161 , n22162 , n22163 , n22164 , n22165 , n22166 , n22167 , n22168 , n22169 , n22170 , n22171 , n22172 , n22173 , n22174 , n22175 , n22176 , n22177 , n22178 , n22179 , n22180 , n22181 , n22182 , n22183 , n22184 , n22185 , n22186 , n22187 , n22188 , n22189 , n22190 , n22191 , n22192 , n22193 , n22194 , n22195 , n22196 , n22197 , n22198 , n22199 , n22200 , n22201 , n22202 , n22203 , n22204 , n22205 , n22206 , n22207 , n22208 , n22209 , n22210 , n22211 , n22212 , n22213 , n22214 , n22215 , n22216 , n22217 , n22218 , n22219 , n22220 , n22221 , n22222 , n22223 , n22224 , n22225 , n22226 , n22227 , n22228 , n22229 , n22230 , n22231 , n22232 , n22233 , n22234 , n22235 , n22236 , n22237 , n22238 , n22239 , n22240 , n22241 , n22242 , n22243 , n22244 , n22245 , n22246 , n22247 , n22248 , n22249 , n22250 , n22251 , n22252 , n22253 , n22254 , n22255 , n22256 , n22257 , n22258 , n22259 , n22260 , n22261 , n22262 , n22263 , n22264 , n22265 , n22266 , n22267 , n22268 , n22269 , n22270 , n22271 , n22272 , n22273 , n22274 , n22275 , n22276 , n22277 , n22278 , n22279 , n22280 , n22281 , n22282 , n22283 , n22284 , n22285 , n22286 , n22287 , n22288 , n22289 , n22290 , n22291 , n22292 , n22293 , n22294 , n22295 , n22296 , n22297 , n22298 , n22299 , n22300 , n22301 , n22302 , n22303 , n22304 , n22305 , n22306 , n22307 , n22308 , n22309 , n22310 , n22311 , n22312 , n22313 , n22314 , n22315 , n22316 , n22317 , n22318 , n22319 , n22320 , n22321 , n22322 , n22323 , n22324 , n22325 , n22326 , n22327 , n22328 , n22329 , n22330 , n22331 , n22332 , n22333 , n22334 , n22335 , n22336 , n22337 , n22338 , n22339 , n22340 , n22341 , n22342 , n22343 , n22344 , n22345 , n22346 , n22347 , n22348 , n22349 , n22350 , n22351 , n22352 , n22353 , n22354 , n22355 , n22356 , n22357 , n22358 , n22359 , n22360 , n22361 , n22362 , n22363 , n22364 , n22365 , n22366 , n22367 , n22368 , n22369 , n22370 , n22371 , n22372 , n22373 , n22374 , n22375 , n22376 , n22377 , n22378 , n22379 , n22380 , n22381 , n22382 , n22383 , n22384 , n22385 , n22386 , n22387 , n22388 , n22389 , n22390 , n22391 , n22392 , n22393 , n22394 , n22395 , n22396 , n22397 , n22398 , n22399 , n22400 , n22401 , n22402 , n22403 , n22404 , n22405 , n22406 , n22407 , n22408 , n22409 , n22410 , n22411 , n22412 , n22413 , n22414 , n22415 , n22416 , n22417 , n22418 , n22419 , n22420 , n22421 , n22422 , n22423 , n22424 , n22425 , n22426 , n22427 , n22428 , n22429 , n22430 , n22431 , n22432 , n22433 , n22434 , n22435 , n22436 , n22437 , n22438 , n22439 , n22440 , n22441 , n22442 , n22443 , n22444 , n22445 , n22446 , n22447 , n22448 , n22449 , n22450 , n22451 , n22452 , n22453 , n22454 , n22455 , n22456 , n22457 , n22458 , n22459 , n22460 , n22461 , n22462 , n22463 , n22464 , n22465 , n22466 , n22467 , n22468 , n22469 , n22470 , n22471 , n22472 , n22473 , n22474 , n22475 , n22476 , n22477 , n22478 , n22479 , n22480 , n22481 , n22482 , n22483 , n22484 , n22485 , n22486 , n22487 , n22488 , n22489 , n22490 , n22491 , n22492 , n22493 , n22494 , n22495 , n22496 , n22497 , n22498 , n22499 , n22500 , n22501 , n22502 , n22503 , n22504 , n22505 , n22506 , n22507 , n22508 , n22509 , n22510 , n22511 , n22512 , n22513 , n22514 , n22515 , n22516 , n22517 , n22518 , n22519 , n22520 , n22521 , n22522 , n22523 , n22524 , n22525 , n22526 , n22527 , n22528 , n22529 , n22530 , n22531 , n22532 , n22533 , n22534 , n22535 , n22536 , n22537 , n22538 , n22539 , n22540 , n22541 , n22542 , n22543 , n22544 , n22545 , n22546 , n22547 , n22548 , n22549 , n22550 , n22551 , n22552 , n22553 , n22554 , n22555 , n22556 , n22557 , n22558 , n22559 , n22560 , n22561 , n22562 , n22563 , n22564 , n22565 , n22566 , n22567 , n22568 , n22569 , n22570 , n22571 , n22572 , n22573 , n22574 , n22575 , n22576 , n22577 , n22578 , n22579 , n22580 , n22581 , n22582 , n22583 , n22584 , n22585 , n22586 , n22587 , n22588 , n22589 , n22590 , n22591 , n22592 , n22593 , n22594 , n22595 , n22596 , n22597 , n22598 , n22599 , n22600 , n22601 , n22602 , n22603 , n22604 , n22605 , n22606 , n22607 , n22608 , n22609 , n22610 , n22611 , n22612 , n22613 , n22614 , n22615 , n22616 , n22617 , n22618 , n22619 , n22620 , n22621 , n22622 , n22623 , n22624 , n22625 , n22626 , n22627 , n22628 , n22629 , n22630 , n22631 , n22632 , n22633 , n22634 , n22635 , n22636 , n22637 , n22638 , n22639 , n22640 , n22641 , n22642 , n22643 , n22644 , n22645 , n22646 , n22647 , n22648 , n22649 , n22650 , n22651 , n22652 , n22653 , n22654 , n22655 , n22656 , n22657 , n22658 , n22659 , n22660 , n22661 , n22662 , n22663 , n22664 , n22665 , n22666 , n22667 , n22668 , n22669 , n22670 , n22671 , n22672 , n22673 , n22674 , n22675 , n22676 , n22677 , n22678 , n22679 , n22680 , n22681 , n22682 , n22683 , n22684 , n22685 , n22686 , n22687 , n22688 , n22689 , n22690 , n22691 , n22692 , n22693 , n22694 , n22695 , n22696 , n22697 , n22698 , n22699 , n22700 , n22701 , n22702 , n22703 , n22704 , n22705 , n22706 , n22707 , n22708 , n22709 , n22710 , n22711 , n22712 , n22713 , n22714 , n22715 , n22716 , n22717 , n22718 , n22719 , n22720 , n22721 , n22722 , n22723 , n22724 , n22725 , n22726 , n22727 , n22728 , n22729 , n22730 , n22731 , n22732 , n22733 , n22734 , n22735 , n22736 , n22737 , n22738 , n22739 , n22740 , n22741 , n22742 , n22743 , n22744 , n22745 , n22746 , n22747 , n22748 , n22749 , n22750 , n22751 , n22752 , n22753 , n22754 , n22755 , n22756 , n22757 , n22758 , n22759 , n22760 , n22761 , n22762 , n22763 , n22764 , n22765 , n22766 , n22767 , n22768 , n22769 , n22770 , n22771 , n22772 , n22773 , n22774 , n22775 , n22776 , n22777 , n22778 , n22779 , n22780 , n22781 , n22782 , n22783 , n22784 , n22785 , n22786 , n22787 , n22788 , n22789 , n22790 , n22791 , n22792 , n22793 , n22794 , n22795 , n22796 , n22797 , n22798 , n22799 , n22800 , n22801 , n22802 , n22803 , n22804 , n22805 , n22806 , n22807 , n22808 , n22809 , n22810 , n22811 , n22812 , n22813 , n22814 , n22815 , n22816 , n22817 , n22818 , n22819 , n22820 , n22821 , n22822 , n22823 , n22824 , n22825 , n22826 , n22827 , n22828 , n22829 , n22830 , n22831 , n22832 , n22833 , n22834 , n22835 , n22836 , n22837 , n22838 , n22839 , n22840 , n22841 , n22842 , n22843 , n22844 , n22845 , n22846 , n22847 , n22848 , n22849 , n22850 , n22851 , n22852 , n22853 , n22854 , n22855 , n22856 , n22857 , n22858 , n22859 , n22860 , n22861 , n22862 , n22863 , n22864 , n22865 , n22866 , n22867 , n22868 , n22869 , n22870 , n22871 , n22872 , n22873 , n22874 , n22875 , n22876 , n22877 , n22878 , n22879 , n22880 , n22881 , n22882 , n22883 , n22884 , n22885 , n22886 , n22887 , n22888 , n22889 , n22890 , n22891 , n22892 , n22893 , n22894 , n22895 , n22896 , n22897 , n22898 , n22899 , n22900 , n22901 , n22902 , n22903 , n22904 , n22905 , n22906 , n22907 , n22908 , n22909 , n22910 , n22911 , n22912 , n22913 , n22914 , n22915 , n22916 , n22917 , n22918 , n22919 , n22920 , n22921 , n22922 , n22923 , n22924 , n22925 , n22926 , n22927 , n22928 , n22929 , n22930 , n22931 , n22932 , n22933 , n22934 , n22935 , n22936 , n22937 , n22938 , n22939 , n22940 , n22941 , n22942 , n22943 , n22944 , n22945 , n22946 , n22947 , n22948 , n22949 , n22950 , n22951 , n22952 , n22953 , n22954 , n22955 , n22956 , n22957 , n22958 , n22959 , n22960 , n22961 , n22962 , n22963 , n22964 , n22965 , n22966 , n22967 , n22968 , n22969 , n22970 , n22971 , n22972 , n22973 , n22974 , n22975 , n22976 , n22977 , n22978 , n22979 , n22980 , n22981 , n22982 , n22983 , n22984 , n22985 , n22986 , n22987 , n22988 , n22989 , n22990 , n22991 , n22992 , n22993 , n22994 , n22995 , n22996 , n22997 , n22998 , n22999 , n23000 , n23001 , n23002 , n23003 , n23004 , n23005 , n23006 , n23007 , n23008 , n23009 , n23010 , n23011 , n23012 , n23013 , n23014 , n23015 , n23016 , n23017 , n23018 , n23019 , n23020 , n23021 , n23022 , n23023 , n23024 , n23025 , n23026 , n23027 , n23028 , n23029 , n23030 , n23031 , n23032 , n23033 , n23034 , n23035 , n23036 , n23037 , n23038 , n23039 , n23040 , n23041 , n23042 , n23043 , n23044 , n23045 , n23046 , n23047 , n23048 , n23049 , n23050 , n23051 , n23052 , n23053 , n23054 , n23055 , n23056 , n23057 , n23058 , n23059 , n23060 , n23061 , n23062 , n23063 , n23064 , n23065 , n23066 , n23067 , n23068 , n23069 , n23070 , n23071 , n23072 , n23073 , n23074 , n23075 , n23076 , n23077 , n23078 , n23079 , n23080 , n23081 , n23082 , n23083 , n23084 , n23085 , n23086 , n23087 , n23088 , n23089 , n23090 , n23091 , n23092 , n23093 , n23094 , n23095 , n23096 , n23097 , n23098 , n23099 , n23100 , n23101 , n23102 , n23103 , n23104 , n23105 , n23106 , n23107 , n23108 , n23109 , n23110 , n23111 , n23112 , n23113 , n23114 , n23115 , n23116 , n23117 , n23118 , n23119 , n23120 , n23121 , n23122 , n23123 , n23124 , n23125 , n23126 , n23127 , n23128 , n23129 , n23130 , n23131 , n23132 , n23133 , n23134 , n23135 , n23136 , n23137 , n23138 , n23139 , n23140 , n23141 , n23142 , n23143 , n23144 , n23145 , n23146 , n23147 , n23148 , n23149 , n23150 , n23151 , n23152 , n23153 , n23154 , n23155 , n23156 , n23157 , n23158 , n23159 , n23160 , n23161 , n23162 , n23163 , n23164 , n23165 , n23166 , n23167 , n23168 , n23169 , n23170 , n23171 , n23172 , n23173 , n23174 , n23175 , n23176 , n23177 , n23178 , n23179 , n23180 , n23181 , n23182 , n23183 , n23184 , n23185 , n23186 , n23187 , n23188 , n23189 , n23190 , n23191 , n23192 , n23193 , n23194 , n23195 , n23196 , n23197 , n23198 , n23199 , n23200 , n23201 , n23202 , n23203 , n23204 , n23205 , n23206 , n23207 , n23208 , n23209 , n23210 , n23211 , n23212 , n23213 , n23214 , n23215 , n23216 , n23217 , n23218 , n23219 , n23220 , n23221 , n23222 , n23223 , n23224 , n23225 , n23226 , n23227 , n23228 , n23229 , n23230 , n23231 , n23232 , n23233 , n23234 , n23235 , n23236 , n23237 , n23238 , n23239 , n23240 , n23241 , n23242 , n23243 , n23244 , n23245 , n23246 , n23247 , n23248 , n23249 , n23250 , n23251 , n23252 , n23253 , n23254 , n23255 , n23256 , n23257 , n23258 , n23259 , n23260 , n23261 , n23262 , n23263 , n23264 , n23265 , n23266 , n23267 , n23268 , n23269 , n23270 , n23271 , n23272 , n23273 , n23274 , n23275 , n23276 , n23277 , n23278 , n23279 , n23280 , n23281 , n23282 , n23283 , n23284 , n23285 , n23286 , n23287 , n23288 , n23289 , n23290 , n23291 , n23292 , n23293 , n23294 , n23295 , n23296 , n23297 , n23298 , n23299 , n23300 , n23301 , n23302 , n23303 , n23304 , n23305 , n23306 , n23307 , n23308 , n23309 , n23310 , n23311 , n23312 , n23313 , n23314 , n23315 , n23316 , n23317 , n23318 , n23319 , n23320 , n23321 , n23322 , n23323 , n23324 , n23325 , n23326 , n23327 , n23328 , n23329 , n23330 , n23331 , n23332 , n23333 , n23334 , n23335 , n23336 , n23337 , n23338 , n23339 , n23340 , n23341 , n23342 , n23343 , n23344 , n23345 , n23346 , n23347 , n23348 , n23349 , n23350 , n23351 , n23352 , n23353 , n23354 , n23355 , n23356 , n23357 , n23358 , n23359 , n23360 , n23361 , n23362 , n23363 , n23364 , n23365 , n23366 , n23367 , n23368 , n23369 , n23370 , n23371 , n23372 , n23373 , n23374 , n23375 , n23376 , n23377 , n23378 , n23379 , n23380 , n23381 , n23382 , n23383 , n23384 , n23385 , n23386 , n23387 , n23388 , n23389 , n23390 , n23391 , n23392 , n23393 , n23394 , n23395 , n23396 , n23397 , n23398 , n23399 , n23400 , n23401 , n23402 , n23403 , n23404 , n23405 , n23406 , n23407 , n23408 , n23409 , n23410 , n23411 , n23412 , n23413 , n23414 , n23415 , n23416 , n23417 , n23418 , n23419 , n23420 , n23421 , n23422 , n23423 , n23424 , n23425 , n23426 , n23427 , n23428 , n23429 , n23430 , n23431 , n23432 , n23433 , n23434 , n23435 , n23436 , n23437 , n23438 , n23439 , n23440 , n23441 , n23442 , n23443 , n23444 , n23445 , n23446 , n23447 , n23448 , n23449 , n23450 , n23451 , n23452 , n23453 , n23454 , n23455 , n23456 , n23457 , n23458 , n23459 , n23460 , n23461 , n23462 , n23463 , n23464 , n23465 , n23466 , n23467 , n23468 , n23469 , n23470 , n23471 , n23472 , n23473 , n23474 , n23475 , n23476 , n23477 , n23478 , n23479 , n23480 , n23481 , n23482 , n23483 , n23484 , n23485 , n23486 , n23487 , n23488 , n23489 , n23490 , n23491 , n23492 , n23493 , n23494 , n23495 , n23496 , n23497 , n23498 , n23499 , n23500 , n23501 , n23502 , n23503 , n23504 , n23505 , n23506 , n23507 , n23508 , n23509 , n23510 , n23511 , n23512 , n23513 , n23514 , n23515 , n23516 , n23517 , n23518 , n23519 , n23520 , n23521 , n23522 , n23523 , n23524 , n23525 , n23526 , n23527 , n23528 , n23529 , n23530 , n23531 , n23532 , n23533 , n23534 , n23535 , n23536 , n23537 , n23538 , n23539 , n23540 , n23541 , n23542 , n23543 , n23544 , n23545 , n23546 , n23547 , n23548 , n23549 , n23550 , n23551 , n23552 , n23553 , n23554 , n23555 , n23556 , n23557 , n23558 , n23559 , n23560 , n23561 , n23562 , n23563 , n23564 , n23565 , n23566 , n23567 , n23568 , n23569 , n23570 , n23571 , n23572 , n23573 , n23574 , n23575 , n23576 , n23577 , n23578 , n23579 , n23580 , n23581 , n23582 , n23583 , n23584 , n23585 , n23586 , n23587 , n23588 , n23589 , n23590 , n23591 , n23592 , n23593 , n23594 , n23595 , n23596 , n23597 , n23598 , n23599 , n23600 , n23601 , n23602 , n23603 , n23604 , n23605 , n23606 , n23607 , n23608 , n23609 , n23610 , n23611 , n23612 , n23613 , n23614 , n23615 , n23616 , n23617 , n23618 , n23619 , n23620 , n23621 , n23622 , n23623 , n23624 , n23625 , n23626 , n23627 , n23628 , n23629 , n23630 , n23631 , n23632 , n23633 , n23634 , n23635 , n23636 , n23637 , n23638 , n23639 , n23640 , n23641 , n23642 , n23643 , n23644 , n23645 , n23646 , n23647 , n23648 , n23649 , n23650 , n23651 , n23652 , n23653 , n23654 , n23655 , n23656 , n23657 , n23658 , n23659 , n23660 , n23661 , n23662 , n23663 , n23664 , n23665 , n23666 , n23667 , n23668 , n23669 , n23670 , n23671 , n23672 , n23673 , n23674 , n23675 , n23676 , n23677 , n23678 , n23679 , n23680 , n23681 , n23682 , n23683 , n23684 , n23685 , n23686 , n23687 , n23688 , n23689 , n23690 , n23691 , n23692 , n23693 , n23694 , n23695 , n23696 , n23697 , n23698 , n23699 , n23700 , n23701 , n23702 , n23703 , n23704 , n23705 , n23706 , n23707 , n23708 , n23709 , n23710 , n23711 , n23712 , n23713 , n23714 , n23715 , n23716 , n23717 , n23718 , n23719 , n23720 , n23721 , n23722 , n23723 , n23724 , n23725 , n23726 , n23727 , n23728 , n23729 , n23730 , n23731 , n23732 , n23733 , n23734 , n23735 , n23736 , n23737 , n23738 , n23739 , n23740 , n23741 , n23742 , n23743 , n23744 , n23745 , n23746 , n23747 , n23748 , n23749 , n23750 , n23751 , n23752 , n23753 , n23754 , n23755 , n23756 , n23757 , n23758 , n23759 , n23760 , n23761 , n23762 , n23763 , n23764 , n23765 , n23766 , n23767 , n23768 , n23769 , n23770 , n23771 , n23772 , n23773 , n23774 , n23775 , n23776 , n23777 , n23778 , n23779 , n23780 , n23781 , n23782 , n23783 , n23784 , n23785 , n23786 , n23787 , n23788 , n23789 , n23790 , n23791 , n23792 , n23793 , n23794 , n23795 , n23796 , n23797 , n23798 , n23799 , n23800 , n23801 , n23802 , n23803 , n23804 , n23805 , n23806 , n23807 , n23808 , n23809 , n23810 , n23811 , n23812 , n23813 , n23814 , n23815 , n23816 , n23817 , n23818 , n23819 , n23820 , n23821 , n23822 , n23823 , n23824 , n23825 , n23826 , n23827 , n23828 , n23829 , n23830 , n23831 , n23832 , n23833 , n23834 , n23835 , n23836 , n23837 , n23838 , n23839 , n23840 , n23841 , n23842 , n23843 , n23844 , n23845 , n23846 , n23847 , n23848 , n23849 , n23850 , n23851 , n23852 , n23853 , n23854 , n23855 , n23856 , n23857 , n23858 , n23859 , n23860 , n23861 , n23862 , n23863 , n23864 , n23865 , n23866 , n23867 , n23868 , n23869 , n23870 , n23871 , n23872 , n23873 , n23874 , n23875 , n23876 , n23877 , n23878 , n23879 , n23880 , n23881 , n23882 , n23883 , n23884 , n23885 , n23886 , n23887 , n23888 , n23889 , n23890 , n23891 , n23892 , n23893 , n23894 , n23895 , n23896 , n23897 , n23898 , n23899 , n23900 , n23901 , n23902 , n23903 , n23904 , n23905 , n23906 , n23907 , n23908 , n23909 , n23910 , n23911 , n23912 , n23913 , n23914 , n23915 , n23916 , n23917 , n23918 , n23919 , n23920 , n23921 , n23922 , n23923 , n23924 , n23925 , n23926 , n23927 , n23928 , n23929 , n23930 , n23931 , n23932 , n23933 , n23934 , n23935 , n23936 , n23937 , n23938 , n23939 , n23940 , n23941 , n23942 , n23943 , n23944 , n23945 , n23946 , n23947 , n23948 , n23949 , n23950 , n23951 , n23952 , n23953 , n23954 , n23955 , n23956 , n23957 , n23958 , n23959 , n23960 , n23961 , n23962 , n23963 , n23964 , n23965 , n23966 , n23967 , n23968 , n23969 , n23970 , n23971 , n23972 , n23973 , n23974 , n23975 , n23976 , n23977 , n23978 , n23979 , n23980 , n23981 , n23982 , n23983 , n23984 , n23985 , n23986 , n23987 , n23988 , n23989 , n23990 , n23991 , n23992 , n23993 , n23994 , n23995 , n23996 , n23997 , n23998 , n23999 , n24000 , n24001 , n24002 , n24003 , n24004 , n24005 , n24006 , n24007 , n24008 , n24009 , n24010 , n24011 , n24012 , n24013 , n24014 , n24015 , n24016 , n24017 , n24018 , n24019 , n24020 , n24021 , n24022 , n24023 , n24024 , n24025 , n24026 , n24027 , n24028 , n24029 , n24030 , n24031 , n24032 , n24033 , n24034 , n24035 , n24036 , n24037 , n24038 , n24039 , n24040 , n24041 , n24042 , n24043 , n24044 , n24045 , n24046 , n24047 , n24048 , n24049 , n24050 , n24051 , n24052 , n24053 , n24054 , n24055 , n24056 , n24057 , n24058 , n24059 , n24060 , n24061 , n24062 , n24063 , n24064 , n24065 , n24066 , n24067 , n24068 , n24069 , n24070 , n24071 , n24072 , n24073 , n24074 , n24075 , n24076 , n24077 , n24078 , n24079 , n24080 , n24081 , n24082 , n24083 , n24084 , n24085 , n24086 , n24087 , n24088 , n24089 , n24090 , n24091 , n24092 , n24093 , n24094 , n24095 , n24096 , n24097 , n24098 , n24099 , n24100 , n24101 , n24102 , n24103 , n24104 , n24105 , n24106 , n24107 , n24108 , n24109 , n24110 , n24111 , n24112 , n24113 , n24114 , n24115 , n24116 , n24117 , n24118 , n24119 , n24120 , n24121 , n24122 , n24123 , n24124 , n24125 , n24126 , n24127 , n24128 , n24129 , n24130 , n24131 , n24132 , n24133 , n24134 , n24135 , n24136 , n24137 , n24138 , n24139 , n24140 , n24141 , n24142 , n24143 , n24144 , n24145 , n24146 , n24147 , n24148 , n24149 , n24150 , n24151 , n24152 , n24153 , n24154 , n24155 , n24156 , n24157 , n24158 , n24159 , n24160 , n24161 , n24162 , n24163 , n24164 , n24165 , n24166 , n24167 , n24168 , n24169 , n24170 , n24171 , n24172 , n24173 , n24174 , n24175 , n24176 , n24177 , n24178 , n24179 , n24180 , n24181 , n24182 , n24183 , n24184 , n24185 , n24186 , n24187 , n24188 , n24189 , n24190 , n24191 , n24192 , n24193 , n24194 , n24195 , n24196 , n24197 , n24198 , n24199 , n24200 , n24201 , n24202 , n24203 , n24204 , n24205 , n24206 , n24207 , n24208 , n24209 , n24210 , n24211 , n24212 , n24213 , n24214 , n24215 , n24216 , n24217 , n24218 , n24219 , n24220 , n24221 , n24222 , n24223 , n24224 , n24225 , n24226 , n24227 , n24228 , n24229 , n24230 , n24231 , n24232 , n24233 , n24234 , n24235 , n24236 , n24237 , n24238 , n24239 , n24240 , n24241 , n24242 , n24243 , n24244 , n24245 , n24246 , n24247 , n24248 , n24249 , n24250 , n24251 , n24252 , n24253 , n24254 , n24255 , n24256 , n24257 , n24258 , n24259 , n24260 , n24261 , n24262 , n24263 , n24264 , n24265 , n24266 , n24267 , n24268 , n24269 , n24270 , n24271 , n24272 , n24273 , n24274 , n24275 , n24276 , n24277 , n24278 , n24279 , n24280 , n24281 , n24282 , n24283 , n24284 , n24285 , n24286 , n24287 , n24288 , n24289 , n24290 , n24291 , n24292 , n24293 , n24294 , n24295 , n24296 , n24297 , n24298 , n24299 , n24300 , n24301 , n24302 , n24303 , n24304 , n24305 , n24306 , n24307 , n24308 , n24309 , n24310 , n24311 , n24312 , n24313 , n24314 , n24315 , n24316 , n24317 , n24318 , n24319 , n24320 , n24321 , n24322 , n24323 , n24324 , n24325 , n24326 , n24327 , n24328 , n24329 , n24330 , n24331 , n24332 , n24333 , n24334 , n24335 , n24336 , n24337 , n24338 , n24339 , n24340 , n24341 , n24342 , n24343 , n24344 , n24345 , n24346 , n24347 , n24348 , n24349 , n24350 , n24351 , n24352 , n24353 , n24354 , n24355 , n24356 , n24357 , n24358 , n24359 , n24360 , n24361 , n24362 , n24363 , n24364 , n24365 , n24366 , n24367 , n24368 , n24369 , n24370 , n24371 , n24372 , n24373 , n24374 , n24375 , n24376 , n24377 , n24378 , n24379 , n24380 , n24381 , n24382 , n24383 , n24384 , n24385 , n24386 , n24387 , n24388 , n24389 , n24390 , n24391 , n24392 , n24393 , n24394 , n24395 , n24396 , n24397 , n24398 , n24399 , n24400 , n24401 , n24402 , n24403 , n24404 , n24405 , n24406 , n24407 , n24408 , n24409 , n24410 , n24411 , n24412 , n24413 , n24414 , n24415 , n24416 , n24417 , n24418 , n24419 , n24420 , n24421 , n24422 , n24423 , n24424 , n24425 , n24426 , n24427 , n24428 , n24429 , n24430 , n24431 , n24432 , n24433 , n24434 , n24435 , n24436 , n24437 , n24438 , n24439 , n24440 , n24441 , n24442 , n24443 , n24444 , n24445 , n24446 , n24447 , n24448 , n24449 , n24450 , n24451 , n24452 , n24453 , n24454 , n24455 , n24456 , n24457 , n24458 , n24459 , n24460 , n24461 , n24462 , n24463 , n24464 , n24465 , n24466 , n24467 , n24468 , n24469 , n24470 , n24471 , n24472 , n24473 , n24474 , n24475 , n24476 , n24477 , n24478 , n24479 , n24480 , n24481 , n24482 , n24483 , n24484 , n24485 , n24486 , n24487 , n24488 , n24489 , n24490 , n24491 , n24492 , n24493 , n24494 , n24495 , n24496 , n24497 , n24498 , n24499 , n24500 , n24501 , n24502 , n24503 , n24504 , n24505 , n24506 , n24507 , n24508 , n24509 , n24510 , n24511 , n24512 , n24513 , n24514 , n24515 , n24516 , n24517 , n24518 , n24519 , n24520 , n24521 , n24522 , n24523 , n24524 , n24525 , n24526 , n24527 , n24528 , n24529 , n24530 , n24531 , n24532 , n24533 , n24534 , n24535 , n24536 , n24537 , n24538 , n24539 , n24540 , n24541 , n24542 , n24543 , n24544 , n24545 , n24546 , n24547 , n24548 , n24549 , n24550 , n24551 , n24552 , n24553 , n24554 , n24555 , n24556 , n24557 , n24558 , n24559 , n24560 , n24561 , n24562 , n24563 , n24564 , n24565 , n24566 , n24567 , n24568 , n24569 , n24570 , n24571 , n24572 , n24573 , n24574 , n24575 , n24576 , n24577 , n24578 , n24579 , n24580 , n24581 , n24582 , n24583 , n24584 , n24585 , n24586 , n24587 , n24588 , n24589 , n24590 , n24591 , n24592 , n24593 , n24594 , n24595 , n24596 , n24597 , n24598 , n24599 , n24600 , n24601 , n24602 , n24603 , n24604 , n24605 , n24606 , n24607 , n24608 , n24609 , n24610 , n24611 , n24612 , n24613 , n24614 , n24615 , n24616 , n24617 , n24618 , n24619 , n24620 , n24621 , n24622 , n24623 , n24624 , n24625 , n24626 , n24627 , n24628 , n24629 , n24630 , n24631 , n24632 , n24633 , n24634 , n24635 , n24636 , n24637 , n24638 , n24639 , n24640 , n24641 , n24642 , n24643 , n24644 , n24645 , n24646 , n24647 , n24648 , n24649 , n24650 , n24651 , n24652 , n24653 , n24654 , n24655 , n24656 , n24657 , n24658 , n24659 , n24660 , n24661 , n24662 , n24663 , n24664 , n24665 , n24666 , n24667 , n24668 , n24669 , n24670 , n24671 , n24672 , n24673 , n24674 , n24675 , n24676 , n24677 , n24678 , n24679 , n24680 , n24681 , n24682 , n24683 , n24684 , n24685 , n24686 , n24687 , n24688 , n24689 , n24690 , n24691 , n24692 , n24693 , n24694 , n24695 , n24696 , n24697 , n24698 , n24699 , n24700 , n24701 , n24702 , n24703 , n24704 , n24705 , n24706 , n24707 , n24708 , n24709 , n24710 , n24711 , n24712 , n24713 , n24714 , n24715 , n24716 , n24717 , n24718 , n24719 , n24720 , n24721 , n24722 , n24723 , n24724 , n24725 , n24726 , n24727 , n24728 , n24729 , n24730 , n24731 , n24732 , n24733 , n24734 , n24735 , n24736 , n24737 , n24738 , n24739 , n24740 , n24741 , n24742 , n24743 , n24744 , n24745 , n24746 , n24747 , n24748 , n24749 , n24750 , n24751 , n24752 , n24753 , n24754 , n24755 , n24756 , n24757 , n24758 , n24759 , n24760 , n24761 , n24762 , n24763 , n24764 , n24765 , n24766 , n24767 , n24768 , n24769 , n24770 , n24771 , n24772 , n24773 , n24774 , n24775 , n24776 , n24777 , n24778 , n24779 , n24780 , n24781 , n24782 , n24783 , n24784 , n24785 , n24786 , n24787 , n24788 , n24789 , n24790 , n24791 , n24792 , n24793 , n24794 , n24795 , n24796 , n24797 , n24798 , n24799 , n24800 , n24801 , n24802 , n24803 , n24804 , n24805 , n24806 , n24807 , n24808 , n24809 , n24810 , n24811 , n24812 , n24813 , n24814 , n24815 , n24816 , n24817 , n24818 , n24819 , n24820 , n24821 , n24822 , n24823 , n24824 , n24825 , n24826 , n24827 , n24828 , n24829 , n24830 , n24831 , n24832 , n24833 , n24834 , n24835 , n24836 , n24837 , n24838 , n24839 , n24840 , n24841 , n24842 , n24843 , n24844 , n24845 , n24846 , n24847 , n24848 , n24849 , n24850 , n24851 , n24852 , n24853 , n24854 , n24855 , n24856 , n24857 , n24858 , n24859 , n24860 , n24861 , n24862 , n24863 , n24864 , n24865 , n24866 , n24867 , n24868 , n24869 , n24870 , n24871 , n24872 , n24873 , n24874 , n24875 , n24876 , n24877 , n24878 , n24879 , n24880 , n24881 , n24882 , n24883 , n24884 , n24885 , n24886 , n24887 , n24888 , n24889 , n24890 , n24891 , n24892 , n24893 , n24894 , n24895 , n24896 , n24897 , n24898 , n24899 , n24900 , n24901 , n24902 , n24903 , n24904 , n24905 , n24906 , n24907 , n24908 , n24909 , n24910 , n24911 , n24912 , n24913 , n24914 , n24915 , n24916 , n24917 , n24918 , n24919 , n24920 , n24921 , n24922 , n24923 , n24924 , n24925 , n24926 , n24927 , n24928 , n24929 , n24930 , n24931 , n24932 , n24933 , n24934 , n24935 , n24936 , n24937 , n24938 , n24939 , n24940 , n24941 , n24942 , n24943 , n24944 , n24945 , n24946 , n24947 , n24948 , n24949 , n24950 , n24951 , n24952 , n24953 , n24954 , n24955 , n24956 , n24957 , n24958 , n24959 , n24960 , n24961 , n24962 , n24963 , n24964 , n24965 , n24966 , n24967 , n24968 , n24969 , n24970 , n24971 , n24972 , n24973 , n24974 , n24975 , n24976 , n24977 , n24978 , n24979 , n24980 , n24981 , n24982 , n24983 , n24984 , n24985 , n24986 , n24987 , n24988 , n24989 , n24990 , n24991 , n24992 , n24993 , n24994 , n24995 , n24996 , n24997 , n24998 , n24999 , n25000 , n25001 , n25002 , n25003 , n25004 , n25005 , n25006 , n25007 , n25008 , n25009 , n25010 , n25011 , n25012 , n25013 , n25014 , n25015 , n25016 , n25017 , n25018 , n25019 , n25020 , n25021 , n25022 , n25023 , n25024 , n25025 , n25026 , n25027 , n25028 , n25029 , n25030 , n25031 , n25032 , n25033 , n25034 , n25035 , n25036 , n25037 , n25038 , n25039 , n25040 , n25041 , n25042 , n25043 , n25044 , n25045 , n25046 , n25047 , n25048 , n25049 , n25050 , n25051 , n25052 , n25053 , n25054 , n25055 , n25056 , n25057 , n25058 , n25059 , n25060 , n25061 , n25062 , n25063 , n25064 , n25065 , n25066 , n25067 , n25068 , n25069 , n25070 , n25071 , n25072 , n25073 , n25074 , n25075 , n25076 , n25077 , n25078 , n25079 , n25080 , n25081 , n25082 , n25083 , n25084 , n25085 , n25086 , n25087 , n25088 , n25089 , n25090 , n25091 , n25092 , n25093 , n25094 , n25095 , n25096 , n25097 , n25098 , n25099 , n25100 , n25101 , n25102 , n25103 , n25104 , n25105 , n25106 , n25107 , n25108 , n25109 , n25110 , n25111 , n25112 , n25113 , n25114 , n25115 , n25116 , n25117 , n25118 , n25119 , n25120 , n25121 , n25122 , n25123 , n25124 , n25125 , n25126 , n25127 , n25128 , n25129 , n25130 , n25131 , n25132 , n25133 , n25134 , n25135 , n25136 , n25137 , n25138 , n25139 , n25140 , n25141 , n25142 , n25143 , n25144 , n25145 , n25146 , n25147 , n25148 , n25149 , n25150 , n25151 , n25152 , n25153 , n25154 , n25155 , n25156 , n25157 , n25158 , n25159 , n25160 , n25161 , n25162 , n25163 , n25164 , n25165 , n25166 , n25167 , n25168 , n25169 , n25170 , n25171 , n25172 , n25173 , n25174 , n25175 , n25176 , n25177 , n25178 , n25179 , n25180 , n25181 , n25182 , n25183 , n25184 , n25185 , n25186 , n25187 , n25188 , n25189 , n25190 , n25191 , n25192 , n25193 , n25194 , n25195 , n25196 , n25197 , n25198 , n25199 , n25200 , n25201 , n25202 , n25203 , n25204 , n25205 , n25206 , n25207 , n25208 , n25209 , n25210 , n25211 , n25212 , n25213 , n25214 , n25215 , n25216 , n25217 , n25218 , n25219 , n25220 , n25221 , n25222 , n25223 , n25224 , n25225 , n25226 , n25227 , n25228 , n25229 , n25230 , n25231 , n25232 , n25233 , n25234 , n25235 , n25236 , n25237 , n25238 , n25239 , n25240 , n25241 , n25242 , n25243 , n25244 , n25245 , n25246 , n25247 , n25248 , n25249 , n25250 , n25251 , n25252 , n25253 , n25254 , n25255 , n25256 , n25257 , n25258 , n25259 , n25260 , n25261 , n25262 , n25263 , n25264 , n25265 , n25266 , n25267 , n25268 , n25269 , n25270 , n25271 , n25272 , n25273 , n25274 , n25275 , n25276 , n25277 , n25278 , n25279 , n25280 , n25281 , n25282 , n25283 , n25284 , n25285 , n25286 , n25287 , n25288 , n25289 , n25290 , n25291 , n25292 , n25293 , n25294 , n25295 , n25296 , n25297 , n25298 , n25299 , n25300 , n25301 , n25302 , n25303 , n25304 , n25305 , n25306 , n25307 , n25308 , n25309 , n25310 , n25311 , n25312 , n25313 , n25314 , n25315 , n25316 , n25317 , n25318 , n25319 , n25320 , n25321 , n25322 , n25323 , n25324 , n25325 , n25326 , n25327 , n25328 , n25329 , n25330 , n25331 , n25332 , n25333 , n25334 , n25335 , n25336 , n25337 , n25338 , n25339 , n25340 , n25341 , n25342 , n25343 , n25344 , n25345 , n25346 , n25347 , n25348 , n25349 , n25350 , n25351 , n25352 , n25353 , n25354 , n25355 , n25356 , n25357 , n25358 , n25359 , n25360 , n25361 , n25362 , n25363 , n25364 , n25365 , n25366 , n25367 , n25368 , n25369 , n25370 , n25371 , n25372 , n25373 , n25374 , n25375 , n25376 , n25377 , n25378 , n25379 , n25380 , n25381 , n25382 , n25383 , n25384 , n25385 , n25386 , n25387 , n25388 , n25389 , n25390 , n25391 , n25392 , n25393 , n25394 , n25395 , n25396 , n25397 , n25398 , n25399 , n25400 , n25401 , n25402 , n25403 , n25404 , n25405 , n25406 , n25407 , n25408 , n25409 , n25410 , n25411 , n25412 , n25413 , n25414 , n25415 , n25416 , n25417 , n25418 , n25419 , n25420 , n25421 , n25422 , n25423 , n25424 , n25425 , n25426 , n25427 , n25428 , n25429 , n25430 , n25431 , n25432 , n25433 , n25434 , n25435 , n25436 , n25437 , n25438 , n25439 , n25440 , n25441 , n25442 , n25443 , n25444 , n25445 , n25446 , n25447 , n25448 , n25449 , n25450 , n25451 , n25452 , n25453 , n25454 , n25455 , n25456 , n25457 , n25458 , n25459 , n25460 , n25461 , n25462 , n25463 , n25464 , n25465 , n25466 , n25467 , n25468 , n25469 , n25470 , n25471 , n25472 , n25473 , n25474 , n25475 , n25476 , n25477 , n25478 , n25479 , n25480 , n25481 , n25482 , n25483 , n25484 , n25485 , n25486 , n25487 , n25488 , n25489 , n25490 , n25491 , n25492 , n25493 , n25494 , n25495 , n25496 , n25497 , n25498 , n25499 , n25500 , n25501 , n25502 , n25503 , n25504 , n25505 , n25506 , n25507 , n25508 , n25509 , n25510 , n25511 , n25512 , n25513 , n25514 , n25515 , n25516 , n25517 , n25518 , n25519 , n25520 , n25521 , n25522 , n25523 , n25524 , n25525 , n25526 , n25527 , n25528 , n25529 , n25530 , n25531 , n25532 , n25533 , n25534 , n25535 , n25536 , n25537 , n25538 , n25539 , n25540 , n25541 , n25542 , n25543 , n25544 , n25545 , n25546 , n25547 , n25548 , n25549 , n25550 , n25551 , n25552 , n25553 , n25554 , n25555 , n25556 , n25557 , n25558 , n25559 , n25560 , n25561 , n25562 , n25563 , n25564 , n25565 , n25566 , n25567 , n25568 , n25569 , n25570 , n25571 , n25572 , n25573 , n25574 , n25575 , n25576 , n25577 , n25578 , n25579 , n25580 , n25581 , n25582 , n25583 , n25584 , n25585 , n25586 , n25587 , n25588 , n25589 , n25590 , n25591 , n25592 , n25593 , n25594 , n25595 , n25596 , n25597 , n25598 , n25599 , n25600 , n25601 , n25602 , n25603 , n25604 , n25605 , n25606 , n25607 , n25608 , n25609 , n25610 , n25611 , n25612 , n25613 , n25614 , n25615 , n25616 , n25617 , n25618 , n25619 , n25620 , n25621 , n25622 , n25623 , n25624 , n25625 , n25626 , n25627 , n25628 , n25629 , n25630 , n25631 , n25632 , n25633 , n25634 , n25635 , n25636 , n25637 , n25638 , n25639 , n25640 , n25641 , n25642 , n25643 , n25644 , n25645 , n25646 , n25647 , n25648 , n25649 , n25650 , n25651 , n25652 , n25653 , n25654 , n25655 , n25656 , n25657 , n25658 , n25659 , n25660 , n25661 , n25662 , n25663 , n25664 , n25665 , n25666 , n25667 , n25668 , n25669 , n25670 , n25671 , n25672 , n25673 , n25674 , n25675 , n25676 , n25677 , n25678 , n25679 , n25680 , n25681 , n25682 , n25683 , n25684 , n25685 , n25686 , n25687 , n25688 , n25689 , n25690 , n25691 , n25692 , n25693 , n25694 , n25695 , n25696 , n25697 , n25698 , n25699 , n25700 , n25701 , n25702 , n25703 , n25704 , n25705 , n25706 , n25707 , n25708 , n25709 , n25710 , n25711 , n25712 , n25713 , n25714 , n25715 , n25716 , n25717 , n25718 , n25719 , n25720 , n25721 , n25722 , n25723 , n25724 , n25725 , n25726 , n25727 , n25728 , n25729 , n25730 , n25731 , n25732 , n25733 , n25734 , n25735 , n25736 , n25737 , n25738 , n25739 , n25740 , n25741 , n25742 , n25743 , n25744 , n25745 , n25746 , n25747 , n25748 , n25749 , n25750 , n25751 , n25752 , n25753 , n25754 , n25755 , n25756 , n25757 , n25758 , n25759 , n25760 , n25761 , n25762 , n25763 , n25764 , n25765 , n25766 , n25767 , n25768 , n25769 , n25770 , n25771 , n25772 , n25773 , n25774 , n25775 , n25776 , n25777 , n25778 , n25779 , n25780 , n25781 , n25782 , n25783 , n25784 , n25785 , n25786 , n25787 , n25788 , n25789 , n25790 , n25791 , n25792 , n25793 , n25794 , n25795 , n25796 , n25797 , n25798 , n25799 , n25800 , n25801 , n25802 , n25803 , n25804 , n25805 , n25806 , n25807 , n25808 , n25809 , n25810 , n25811 , n25812 , n25813 , n25814 , n25815 , n25816 , n25817 , n25818 , n25819 , n25820 , n25821 , n25822 , n25823 , n25824 , n25825 , n25826 , n25827 , n25828 , n25829 , n25830 , n25831 , n25832 , n25833 , n25834 , n25835 , n25836 , n25837 , n25838 , n25839 , n25840 , n25841 , n25842 , n25843 , n25844 , n25845 , n25846 , n25847 , n25848 , n25849 , n25850 , n25851 , n25852 , n25853 , n25854 , n25855 , n25856 , n25857 , n25858 , n25859 , n25860 , n25861 , n25862 , n25863 , n25864 , n25865 , n25866 , n25867 , n25868 , n25869 , n25870 , n25871 , n25872 , n25873 , n25874 , n25875 , n25876 , n25877 , n25878 , n25879 , n25880 , n25881 , n25882 , n25883 , n25884 , n25885 , n25886 , n25887 , n25888 , n25889 , n25890 , n25891 , n25892 , n25893 , n25894 , n25895 , n25896 , n25897 , n25898 , n25899 , n25900 , n25901 , n25902 , n25903 , n25904 , n25905 , n25906 , n25907 , n25908 , n25909 , n25910 , n25911 , n25912 , n25913 , n25914 , n25915 , n25916 , n25917 , n25918 , n25919 , n25920 , n25921 , n25922 , n25923 , n25924 , n25925 , n25926 , n25927 , n25928 , n25929 , n25930 , n25931 , n25932 , n25933 , n25934 , n25935 , n25936 , n25937 , n25938 , n25939 , n25940 , n25941 , n25942 , n25943 , n25944 , n25945 , n25946 , n25947 , n25948 , n25949 , n25950 , n25951 , n25952 , n25953 , n25954 , n25955 , n25956 , n25957 , n25958 , n25959 , n25960 , n25961 , n25962 , n25963 , n25964 , n25965 , n25966 , n25967 , n25968 , n25969 , n25970 , n25971 , n25972 , n25973 , n25974 , n25975 , n25976 , n25977 , n25978 , n25979 , n25980 , n25981 , n25982 , n25983 , n25984 , n25985 , n25986 , n25987 , n25988 , n25989 , n25990 , n25991 , n25992 , n25993 , n25994 , n25995 , n25996 , n25997 , n25998 , n25999 , n26000 , n26001 , n26002 , n26003 , n26004 , n26005 , n26006 , n26007 , n26008 , n26009 , n26010 , n26011 , n26012 , n26013 , n26014 , n26015 , n26016 , n26017 , n26018 , n26019 , n26020 , n26021 , n26022 , n26023 , n26024 , n26025 , n26026 , n26027 , n26028 , n26029 , n26030 , n26031 , n26032 , n26033 , n26034 , n26035 , n26036 , n26037 , n26038 , n26039 , n26040 , n26041 , n26042 , n26043 , n26044 , n26045 , n26046 , n26047 , n26048 , n26049 , n26050 , n26051 , n26052 , n26053 , n26054 , n26055 , n26056 , n26057 , n26058 , n26059 , n26060 , n26061 , n26062 , n26063 , n26064 , n26065 , n26066 , n26067 , n26068 , n26069 , n26070 , n26071 , n26072 , n26073 , n26074 , n26075 , n26076 , n26077 , n26078 , n26079 , n26080 , n26081 , n26082 , n26083 , n26084 , n26085 , n26086 , n26087 , n26088 , n26089 , n26090 , n26091 , n26092 , n26093 , n26094 , n26095 , n26096 , n26097 , n26098 , n26099 , n26100 , n26101 , n26102 , n26103 , n26104 , n26105 , n26106 , n26107 , n26108 , n26109 , n26110 , n26111 , n26112 , n26113 , n26114 , n26115 , n26116 , n26117 , n26118 , n26119 , n26120 , n26121 , n26122 , n26123 , n26124 , n26125 , n26126 , n26127 , n26128 , n26129 , n26130 , n26131 , n26132 , n26133 , n26134 , n26135 , n26136 , n26137 , n26138 , n26139 , n26140 , n26141 , n26142 , n26143 , n26144 , n26145 , n26146 , n26147 , n26148 , n26149 , n26150 , n26151 , n26152 , n26153 , n26154 , n26155 , n26156 , n26157 , n26158 , n26159 , n26160 , n26161 , n26162 , n26163 , n26164 , n26165 , n26166 , n26167 , n26168 , n26169 , n26170 , n26171 , n26172 , n26173 , n26174 , n26175 , n26176 , n26177 , n26178 , n26179 , n26180 , n26181 , n26182 , n26183 , n26184 , n26185 , n26186 , n26187 , n26188 , n26189 , n26190 , n26191 , n26192 , n26193 , n26194 , n26195 , n26196 , n26197 , n26198 , n26199 , n26200 , n26201 , n26202 , n26203 , n26204 , n26205 , n26206 , n26207 , n26208 , n26209 , n26210 , n26211 , n26212 , n26213 , n26214 , n26215 , n26216 , n26217 , n26218 , n26219 , n26220 , n26221 , n26222 , n26223 , n26224 , n26225 , n26226 , n26227 , n26228 , n26229 , n26230 , n26231 , n26232 , n26233 , n26234 , n26235 , n26236 , n26237 , n26238 , n26239 , n26240 , n26241 , n26242 , n26243 , n26244 , n26245 , n26246 , n26247 , n26248 , n26249 , n26250 , n26251 , n26252 , n26253 , n26254 , n26255 , n26256 , n26257 , n26258 , n26259 , n26260 , n26261 , n26262 , n26263 , n26264 , n26265 , n26266 , n26267 , n26268 , n26269 , n26270 , n26271 , n26272 , n26273 , n26274 , n26275 , n26276 , n26277 , n26278 , n26279 , n26280 , n26281 , n26282 , n26283 , n26284 , n26285 , n26286 , n26287 , n26288 , n26289 , n26290 , n26291 , n26292 , n26293 , n26294 , n26295 , n26296 , n26297 , n26298 , n26299 , n26300 , n26301 , n26302 , n26303 , n26304 , n26305 , n26306 , n26307 , n26308 , n26309 , n26310 , n26311 , n26312 , n26313 , n26314 , n26315 , n26316 , n26317 , n26318 , n26319 , n26320 , n26321 , n26322 , n26323 , n26324 , n26325 , n26326 , n26327 , n26328 , n26329 , n26330 , n26331 , n26332 , n26333 , n26334 , n26335 , n26336 , n26337 , n26338 , n26339 , n26340 , n26341 , n26342 , n26343 , n26344 , n26345 , n26346 , n26347 , n26348 , n26349 , n26350 , n26351 , n26352 , n26353 , n26354 , n26355 , n26356 , n26357 , n26358 , n26359 , n26360 , n26361 , n26362 , n26363 , n26364 , n26365 , n26366 , n26367 , n26368 , n26369 , n26370 , n26371 , n26372 , n26373 , n26374 , n26375 , n26376 , n26377 , n26378 , n26379 , n26380 , n26381 , n26382 , n26383 , n26384 , n26385 , n26386 , n26387 , n26388 , n26389 , n26390 , n26391 , n26392 , n26393 , n26394 , n26395 , n26396 , n26397 , n26398 , n26399 , n26400 , n26401 , n26402 , n26403 , n26404 , n26405 , n26406 , n26407 , n26408 , n26409 , n26410 , n26411 , n26412 , n26413 , n26414 , n26415 , n26416 , n26417 , n26418 , n26419 , n26420 , n26421 , n26422 , n26423 , n26424 , n26425 , n26426 , n26427 , n26428 , n26429 , n26430 , n26431 , n26432 , n26433 , n26434 , n26435 , n26436 , n26437 , n26438 , n26439 , n26440 , n26441 , n26442 , n26443 , n26444 , n26445 , n26446 , n26447 , n26448 , n26449 , n26450 , n26451 , n26452 , n26453 , n26454 , n26455 , n26456 , n26457 , n26458 , n26459 , n26460 , n26461 , n26462 , n26463 , n26464 , n26465 , n26466 , n26467 , n26468 , n26469 , n26470 , n26471 , n26472 , n26473 , n26474 , n26475 , n26476 , n26477 , n26478 , n26479 , n26480 , n26481 , n26482 , n26483 , n26484 , n26485 , n26486 , n26487 , n26488 , n26489 , n26490 , n26491 , n26492 , n26493 , n26494 , n26495 , n26496 , n26497 , n26498 , n26499 , n26500 , n26501 , n26502 , n26503 , n26504 , n26505 , n26506 , n26507 , n26508 , n26509 , n26510 , n26511 , n26512 , n26513 , n26514 , n26515 , n26516 , n26517 , n26518 , n26519 , n26520 , n26521 , n26522 , n26523 , n26524 , n26525 , n26526 , n26527 , n26528 , n26529 , n26530 , n26531 , n26532 , n26533 , n26534 , n26535 , n26536 , n26537 , n26538 , n26539 , n26540 , n26541 , n26542 , n26543 , n26544 , n26545 , n26546 , n26547 , n26548 , n26549 , n26550 , n26551 , n26552 , n26553 , n26554 , n26555 , n26556 , n26557 , n26558 , n26559 , n26560 , n26561 , n26562 , n26563 , n26564 , n26565 , n26566 , n26567 , n26568 , n26569 , n26570 , n26571 , n26572 , n26573 , n26574 , n26575 , n26576 , n26577 , n26578 , n26579 , n26580 , n26581 , n26582 , n26583 , n26584 , n26585 , n26586 , n26587 , n26588 , n26589 , n26590 , n26591 , n26592 , n26593 , n26594 , n26595 , n26596 , n26597 , n26598 , n26599 , n26600 , n26601 , n26602 , n26603 , n26604 , n26605 , n26606 , n26607 , n26608 , n26609 , n26610 , n26611 , n26612 , n26613 , n26614 , n26615 , n26616 , n26617 , n26618 , n26619 , n26620 , n26621 , n26622 , n26623 , n26624 , n26625 , n26626 , n26627 , n26628 , n26629 , n26630 , n26631 , n26632 , n26633 , n26634 , n26635 , n26636 , n26637 , n26638 , n26639 , n26640 , n26641 , n26642 , n26643 , n26644 , n26645 , n26646 , n26647 , n26648 , n26649 , n26650 , n26651 , n26652 , n26653 , n26654 , n26655 , n26656 , n26657 , n26658 , n26659 , n26660 , n26661 , n26662 , n26663 , n26664 , n26665 , n26666 , n26667 , n26668 , n26669 , n26670 , n26671 , n26672 , n26673 , n26674 , n26675 , n26676 , n26677 , n26678 , n26679 , n26680 , n26681 , n26682 , n26683 , n26684 , n26685 , n26686 , n26687 , n26688 , n26689 , n26690 , n26691 , n26692 , n26693 , n26694 , n26695 , n26696 , n26697 , n26698 , n26699 , n26700 , n26701 , n26702 , n26703 , n26704 , n26705 , n26706 , n26707 , n26708 , n26709 , n26710 , n26711 , n26712 , n26713 , n26714 , n26715 , n26716 , n26717 , n26718 , n26719 , n26720 , n26721 , n26722 , n26723 , n26724 , n26725 , n26726 , n26727 , n26728 , n26729 , n26730 , n26731 , n26732 , n26733 , n26734 , n26735 , n26736 , n26737 , n26738 , n26739 , n26740 , n26741 , n26742 , n26743 , n26744 , n26745 , n26746 , n26747 , n26748 , n26749 , n26750 , n26751 , n26752 , n26753 , n26754 , n26755 , n26756 , n26757 , n26758 , n26759 , n26760 , n26761 , n26762 , n26763 , n26764 , n26765 , n26766 , n26767 , n26768 , n26769 , n26770 , n26771 , n26772 , n26773 , n26774 , n26775 , n26776 , n26777 , n26778 , n26779 , n26780 , n26781 , n26782 , n26783 , n26784 , n26785 , n26786 , n26787 , n26788 , n26789 , n26790 , n26791 , n26792 , n26793 , n26794 , n26795 , n26796 , n26797 , n26798 , n26799 , n26800 , n26801 , n26802 , n26803 , n26804 , n26805 , n26806 , n26807 , n26808 , n26809 , n26810 , n26811 , n26812 , n26813 , n26814 , n26815 , n26816 , n26817 , n26818 , n26819 , n26820 , n26821 , n26822 , n26823 , n26824 , n26825 , n26826 , n26827 , n26828 , n26829 , n26830 , n26831 , n26832 , n26833 , n26834 , n26835 , n26836 , n26837 , n26838 , n26839 , n26840 , n26841 , n26842 , n26843 , n26844 , n26845 , n26846 , n26847 , n26848 , n26849 , n26850 , n26851 , n26852 , n26853 , n26854 , n26855 , n26856 , n26857 , n26858 , n26859 , n26860 , n26861 , n26862 , n26863 , n26864 , n26865 , n26866 , n26867 , n26868 , n26869 , n26870 , n26871 , n26872 , n26873 , n26874 , n26875 , n26876 , n26877 , n26878 , n26879 , n26880 , n26881 , n26882 , n26883 , n26884 , n26885 , n26886 , n26887 , n26888 , n26889 , n26890 , n26891 , n26892 , n26893 , n26894 , n26895 , n26896 , n26897 , n26898 , n26899 , n26900 , n26901 , n26902 , n26903 , n26904 , n26905 , n26906 , n26907 , n26908 , n26909 , n26910 , n26911 , n26912 , n26913 , n26914 , n26915 , n26916 , n26917 , n26918 , n26919 , n26920 , n26921 , n26922 , n26923 , n26924 , n26925 , n26926 , n26927 , n26928 , n26929 , n26930 , n26931 , n26932 , n26933 , n26934 , n26935 , n26936 , n26937 , n26938 , n26939 , n26940 , n26941 , n26942 , n26943 , n26944 , n26945 , n26946 , n26947 , n26948 , n26949 , n26950 , n26951 , n26952 , n26953 , n26954 , n26955 , n26956 , n26957 , n26958 , n26959 , n26960 , n26961 , n26962 , n26963 , n26964 , n26965 , n26966 , n26967 , n26968 , n26969 , n26970 , n26971 , n26972 , n26973 , n26974 , n26975 , n26976 , n26977 , n26978 , n26979 , n26980 , n26981 , n26982 , n26983 , n26984 , n26985 , n26986 , n26987 , n26988 , n26989 , n26990 , n26991 , n26992 , n26993 , n26994 , n26995 , n26996 , n26997 , n26998 , n26999 , n27000 , n27001 , n27002 , n27003 , n27004 , n27005 , n27006 , n27007 , n27008 , n27009 , n27010 , n27011 , n27012 , n27013 , n27014 , n27015 , n27016 , n27017 , n27018 , n27019 , n27020 , n27021 , n27022 , n27023 , n27024 , n27025 , n27026 , n27027 , n27028 , n27029 , n27030 , n27031 , n27032 , n27033 , n27034 , n27035 , n27036 , n27037 , n27038 , n27039 , n27040 , n27041 , n27042 , n27043 , n27044 , n27045 , n27046 , n27047 , n27048 , n27049 , n27050 , n27051 , n27052 , n27053 , n27054 , n27055 , n27056 , n27057 , n27058 , n27059 , n27060 , n27061 , n27062 , n27063 , n27064 , n27065 , n27066 , n27067 , n27068 , n27069 , n27070 , n27071 , n27072 , n27073 , n27074 , n27075 , n27076 , n27077 , n27078 , n27079 , n27080 , n27081 , n27082 , n27083 , n27084 , n27085 , n27086 , n27087 , n27088 , n27089 , n27090 , n27091 , n27092 , n27093 , n27094 , n27095 , n27096 , n27097 , n27098 , n27099 , n27100 , n27101 , n27102 , n27103 , n27104 , n27105 , n27106 , n27107 , n27108 , n27109 , n27110 , n27111 , n27112 , n27113 , n27114 , n27115 , n27116 , n27117 , n27118 , n27119 , n27120 , n27121 , n27122 , n27123 , n27124 , n27125 , n27126 , n27127 , n27128 , n27129 , n27130 , n27131 , n27132 , n27133 , n27134 , n27135 , n27136 , n27137 , n27138 , n27139 , n27140 , n27141 , n27142 , n27143 , n27144 , n27145 , n27146 , n27147 , n27148 , n27149 , n27150 , n27151 , n27152 , n27153 , n27154 , n27155 , n27156 , n27157 , n27158 , n27159 , n27160 , n27161 , n27162 , n27163 , n27164 , n27165 , n27166 , n27167 , n27168 , n27169 , n27170 , n27171 , n27172 , n27173 , n27174 , n27175 , n27176 , n27177 , n27178 , n27179 , n27180 , n27181 , n27182 , n27183 , n27184 , n27185 , n27186 , n27187 , n27188 , n27189 , n27190 , n27191 , n27192 , n27193 , n27194 , n27195 , n27196 , n27197 , n27198 , n27199 , n27200 , n27201 , n27202 , n27203 , n27204 , n27205 , n27206 , n27207 , n27208 , n27209 , n27210 , n27211 , n27212 , n27213 , n27214 , n27215 , n27216 , n27217 , n27218 , n27219 , n27220 , n27221 , n27222 , n27223 , n27224 , n27225 , n27226 , n27227 , n27228 , n27229 , n27230 , n27231 , n27232 , n27233 , n27234 , n27235 , n27236 , n27237 , n27238 , n27239 , n27240 , n27241 , n27242 , n27243 , n27244 , n27245 , n27246 , n27247 , n27248 , n27249 , n27250 , n27251 , n27252 , n27253 , n27254 , n27255 , n27256 , n27257 , n27258 , n27259 , n27260 , n27261 , n27262 , n27263 , n27264 , n27265 , n27266 , n27267 , n27268 , n27269 , n27270 , n27271 , n27272 , n27273 , n27274 , n27275 , n27276 , n27277 , n27278 , n27279 , n27280 , n27281 , n27282 , n27283 , n27284 , n27285 , n27286 , n27287 , n27288 , n27289 , n27290 , n27291 , n27292 , n27293 , n27294 , n27295 , n27296 , n27297 , n27298 , n27299 , n27300 , n27301 , n27302 , n27303 , n27304 , n27305 , n27306 , n27307 , n27308 , n27309 , n27310 , n27311 , n27312 , n27313 , n27314 , n27315 , n27316 , n27317 , n27318 , n27319 , n27320 , n27321 , n27322 , n27323 , n27324 , n27325 , n27326 , n27327 , n27328 , n27329 , n27330 , n27331 , n27332 , n27333 , n27334 , n27335 , n27336 , n27337 , n27338 , n27339 , n27340 , n27341 , n27342 , n27343 , n27344 , n27345 , n27346 , n27347 , n27348 , n27349 , n27350 , n27351 , n27352 , n27353 , n27354 , n27355 , n27356 , n27357 , n27358 , n27359 , n27360 , n27361 , n27362 , n27363 , n27364 , n27365 , n27366 , n27367 , n27368 , n27369 , n27370 , n27371 , n27372 , n27373 , n27374 , n27375 , n27376 , n27377 , n27378 , n27379 , n27380 , n27381 , n27382 , n27383 , n27384 , n27385 , n27386 , n27387 , n27388 , n27389 , n27390 , n27391 , n27392 , n27393 , n27394 , n27395 , n27396 , n27397 , n27398 , n27399 , n27400 , n27401 , n27402 , n27403 , n27404 , n27405 , n27406 , n27407 , n27408 , n27409 , n27410 , n27411 , n27412 , n27413 , n27414 , n27415 , n27416 , n27417 , n27418 , n27419 , n27420 , n27421 , n27422 , n27423 , n27424 , n27425 , n27426 , n27427 , n27428 , n27429 , n27430 , n27431 , n27432 , n27433 , n27434 , n27435 , n27436 , n27437 , n27438 , n27439 , n27440 , n27441 , n27442 , n27443 , n27444 , n27445 , n27446 , n27447 , n27448 , n27449 , n27450 , n27451 , n27452 , n27453 , n27454 , n27455 , n27456 , n27457 , n27458 , n27459 , n27460 , n27461 , n27462 , n27463 , n27464 , n27465 , n27466 , n27467 , n27468 , n27469 , n27470 , n27471 , n27472 , n27473 , n27474 , n27475 , n27476 , n27477 , n27478 , n27479 , n27480 , n27481 , n27482 , n27483 , n27484 , n27485 , n27486 , n27487 , n27488 , n27489 , n27490 , n27491 , n27492 , n27493 , n27494 , n27495 , n27496 , n27497 , n27498 , n27499 , n27500 , n27501 , n27502 , n27503 , n27504 , n27505 , n27506 , n27507 , n27508 , n27509 , n27510 , n27511 , n27512 , n27513 , n27514 , n27515 , n27516 , n27517 , n27518 , n27519 , n27520 , n27521 , n27522 , n27523 , n27524 , n27525 , n27526 , n27527 , n27528 , n27529 , n27530 , n27531 , n27532 , n27533 , n27534 , n27535 , n27536 , n27537 , n27538 , n27539 , n27540 , n27541 , n27542 , n27543 , n27544 , n27545 , n27546 , n27547 , n27548 , n27549 , n27550 , n27551 , n27552 , n27553 , n27554 , n27555 , n27556 , n27557 , n27558 , n27559 , n27560 , n27561 , n27562 , n27563 , n27564 , n27565 , n27566 , n27567 , n27568 , n27569 , n27570 , n27571 , n27572 , n27573 , n27574 , n27575 , n27576 , n27577 , n27578 , n27579 , n27580 , n27581 , n27582 , n27583 , n27584 , n27585 , n27586 , n27587 , n27588 , n27589 , n27590 , n27591 , n27592 , n27593 , n27594 , n27595 , n27596 , n27597 , n27598 , n27599 , n27600 , n27601 , n27602 , n27603 , n27604 , n27605 , n27606 , n27607 , n27608 , n27609 , n27610 , n27611 , n27612 , n27613 , n27614 , n27615 , n27616 , n27617 , n27618 , n27619 , n27620 , n27621 , n27622 , n27623 , n27624 , n27625 , n27626 , n27627 , n27628 , n27629 , n27630 , n27631 , n27632 , n27633 , n27634 , n27635 , n27636 , n27637 , n27638 , n27639 , n27640 , n27641 , n27642 , n27643 , n27644 , n27645 , n27646 , n27647 , n27648 , n27649 , n27650 , n27651 , n27652 , n27653 , n27654 , n27655 , n27656 , n27657 , n27658 , n27659 , n27660 , n27661 , n27662 , n27663 , n27664 , n27665 , n27666 , n27667 , n27668 , n27669 , n27670 , n27671 , n27672 , n27673 , n27674 , n27675 , n27676 , n27677 , n27678 , n27679 , n27680 , n27681 , n27682 , n27683 , n27684 , n27685 , n27686 , n27687 , n27688 , n27689 , n27690 , n27691 , n27692 , n27693 , n27694 , n27695 , n27696 , n27697 , n27698 , n27699 , n27700 , n27701 , n27702 , n27703 , n27704 , n27705 , n27706 , n27707 , n27708 , n27709 , n27710 , n27711 , n27712 , n27713 , n27714 , n27715 , n27716 , n27717 , n27718 , n27719 , n27720 , n27721 , n27722 , n27723 , n27724 , n27725 , n27726 , n27727 , n27728 , n27729 , n27730 , n27731 , n27732 , n27733 , n27734 , n27735 , n27736 , n27737 , n27738 , n27739 , n27740 , n27741 , n27742 , n27743 , n27744 , n27745 , n27746 , n27747 , n27748 , n27749 , n27750 , n27751 , n27752 , n27753 , n27754 , n27755 , n27756 , n27757 , n27758 , n27759 , n27760 , n27761 , n27762 , n27763 , n27764 , n27765 , n27766 , n27767 , n27768 , n27769 , n27770 , n27771 , n27772 , n27773 , n27774 , n27775 , n27776 , n27777 , n27778 , n27779 , n27780 , n27781 , n27782 , n27783 , n27784 , n27785 , n27786 , n27787 , n27788 , n27789 , n27790 , n27791 , n27792 , n27793 , n27794 , n27795 , n27796 , n27797 , n27798 , n27799 , n27800 , n27801 , n27802 , n27803 , n27804 , n27805 , n27806 , n27807 , n27808 , n27809 , n27810 , n27811 , n27812 , n27813 , n27814 , n27815 , n27816 , n27817 , n27818 , n27819 , n27820 , n27821 , n27822 , n27823 , n27824 , n27825 , n27826 , n27827 , n27828 , n27829 , n27830 , n27831 , n27832 , n27833 , n27834 , n27835 , n27836 , n27837 , n27838 , n27839 , n27840 , n27841 , n27842 , n27843 , n27844 , n27845 , n27846 , n27847 , n27848 , n27849 , n27850 , n27851 , n27852 , n27853 , n27854 , n27855 , n27856 , n27857 , n27858 , n27859 , n27860 , n27861 , n27862 , n27863 , n27864 , n27865 , n27866 , n27867 , n27868 , n27869 , n27870 , n27871 , n27872 , n27873 , n27874 , n27875 , n27876 , n27877 , n27878 , n27879 , n27880 , n27881 , n27882 , n27883 , n27884 , n27885 , n27886 , n27887 , n27888 , n27889 , n27890 , n27891 , n27892 , n27893 , n27894 , n27895 , n27896 , n27897 , n27898 , n27899 , n27900 , n27901 , n27902 , n27903 , n27904 , n27905 , n27906 , n27907 , n27908 , n27909 , n27910 , n27911 , n27912 , n27913 , n27914 , n27915 , n27916 , n27917 , n27918 , n27919 , n27920 , n27921 , n27922 , n27923 , n27924 , n27925 , n27926 , n27927 , n27928 , n27929 , n27930 , n27931 , n27932 , n27933 , n27934 , n27935 , n27936 , n27937 , n27938 , n27939 , n27940 , n27941 , n27942 , n27943 , n27944 , n27945 , n27946 , n27947 , n27948 , n27949 , n27950 , n27951 , n27952 , n27953 , n27954 , n27955 , n27956 , n27957 , n27958 , n27959 , n27960 , n27961 , n27962 , n27963 , n27964 , n27965 , n27966 , n27967 , n27968 , n27969 , n27970 , n27971 , n27972 , n27973 , n27974 , n27975 , n27976 , n27977 , n27978 , n27979 , n27980 , n27981 , n27982 , n27983 , n27984 , n27985 , n27986 , n27987 , n27988 , n27989 , n27990 , n27991 , n27992 , n27993 , n27994 , n27995 , n27996 , n27997 , n27998 , n27999 , n28000 , n28001 , n28002 , n28003 , n28004 , n28005 , n28006 , n28007 , n28008 , n28009 , n28010 , n28011 , n28012 , n28013 , n28014 , n28015 , n28016 , n28017 , n28018 , n28019 , n28020 , n28021 , n28022 , n28023 , n28024 , n28025 , n28026 , n28027 , n28028 , n28029 , n28030 , n28031 , n28032 , n28033 , n28034 , n28035 , n28036 , n28037 , n28038 , n28039 , n28040 , n28041 , n28042 , n28043 , n28044 , n28045 , n28046 , n28047 , n28048 , n28049 , n28050 , n28051 , n28052 , n28053 , n28054 , n28055 , n28056 , n28057 , n28058 , n28059 , n28060 , n28061 , n28062 , n28063 , n28064 , n28065 , n28066 , n28067 , n28068 , n28069 , n28070 , n28071 , n28072 , n28073 , n28074 , n28075 , n28076 , n28077 , n28078 , n28079 , n28080 , n28081 , n28082 , n28083 , n28084 , n28085 , n28086 , n28087 , n28088 , n28089 , n28090 , n28091 , n28092 , n28093 , n28094 , n28095 , n28096 , n28097 , n28098 , n28099 , n28100 , n28101 , n28102 , n28103 , n28104 , n28105 , n28106 , n28107 , n28108 , n28109 , n28110 , n28111 , n28112 , n28113 , n28114 , n28115 , n28116 , n28117 , n28118 , n28119 , n28120 , n28121 , n28122 , n28123 , n28124 , n28125 , n28126 , n28127 , n28128 , n28129 , n28130 , n28131 , n28132 , n28133 , n28134 , n28135 , n28136 , n28137 , n28138 , n28139 , n28140 , n28141 , n28142 , n28143 , n28144 , n28145 , n28146 , n28147 , n28148 , n28149 , n28150 , n28151 , n28152 , n28153 , n28154 , n28155 , n28156 , n28157 , n28158 , n28159 , n28160 , n28161 , n28162 , n28163 , n28164 , n28165 , n28166 , n28167 , n28168 , n28169 , n28170 , n28171 , n28172 , n28173 , n28174 , n28175 , n28176 , n28177 , n28178 , n28179 , n28180 , n28181 , n28182 , n28183 , n28184 , n28185 , n28186 , n28187 , n28188 , n28189 , n28190 , n28191 , n28192 , n28193 , n28194 , n28195 , n28196 , n28197 , n28198 , n28199 , n28200 , n28201 , n28202 , n28203 , n28204 , n28205 , n28206 , n28207 , n28208 , n28209 , n28210 , n28211 , n28212 , n28213 , n28214 , n28215 , n28216 , n28217 , n28218 , n28219 , n28220 , n28221 , n28222 , n28223 , n28224 , n28225 , n28226 , n28227 , n28228 , n28229 , n28230 , n28231 , n28232 , n28233 , n28234 , n28235 , n28236 , n28237 , n28238 , n28239 , n28240 , n28241 , n28242 , n28243 , n28244 , n28245 , n28246 , n28247 , n28248 , n28249 , n28250 , n28251 , n28252 , n28253 , n28254 , n28255 , n28256 , n28257 , n28258 , n28259 , n28260 , n28261 , n28262 , n28263 , n28264 , n28265 , n28266 , n28267 , n28268 , n28269 , n28270 , n28271 , n28272 , n28273 , n28274 , n28275 , n28276 , n28277 , n28278 , n28279 , n28280 , n28281 , n28282 , n28283 , n28284 , n28285 , n28286 , n28287 , n28288 , n28289 , n28290 , n28291 , n28292 , n28293 , n28294 , n28295 , n28296 , n28297 , n28298 , n28299 , n28300 , n28301 , n28302 , n28303 , n28304 , n28305 , n28306 , n28307 , n28308 , n28309 , n28310 , n28311 , n28312 , n28313 , n28314 , n28315 , n28316 , n28317 , n28318 , n28319 , n28320 , n28321 , n28322 , n28323 , n28324 , n28325 , n28326 , n28327 , n28328 , n28329 , n28330 , n28331 , n28332 , n28333 , n28334 , n28335 , n28336 , n28337 , n28338 , n28339 , n28340 , n28341 , n28342 , n28343 , n28344 , n28345 , n28346 , n28347 , n28348 , n28349 , n28350 , n28351 , n28352 , n28353 , n28354 , n28355 , n28356 , n28357 , n28358 , n28359 , n28360 , n28361 , n28362 , n28363 , n28364 , n28365 , n28366 , n28367 , n28368 , n28369 , n28370 , n28371 , n28372 , n28373 , n28374 , n28375 , n28376 , n28377 , n28378 , n28379 , n28380 , n28381 , n28382 , n28383 , n28384 , n28385 , n28386 , n28387 , n28388 , n28389 , n28390 , n28391 , n28392 , n28393 , n28394 , n28395 , n28396 , n28397 , n28398 , n28399 , n28400 , n28401 , n28402 , n28403 , n28404 , n28405 , n28406 , n28407 , n28408 , n28409 , n28410 , n28411 , n28412 , n28413 , n28414 , n28415 , n28416 , n28417 , n28418 , n28419 , n28420 , n28421 , n28422 , n28423 , n28424 , n28425 , n28426 , n28427 , n28428 , n28429 , n28430 , n28431 , n28432 , n28433 , n28434 , n28435 , n28436 , n28437 , n28438 , n28439 , n28440 , n28441 , n28442 , n28443 , n28444 , n28445 , n28446 , n28447 , n28448 , n28449 , n28450 , n28451 , n28452 , n28453 , n28454 , n28455 , n28456 , n28457 , n28458 , n28459 , n28460 , n28461 , n28462 , n28463 , n28464 , n28465 , n28466 , n28467 , n28468 , n28469 , n28470 , n28471 , n28472 , n28473 , n28474 , n28475 , n28476 , n28477 , n28478 , n28479 , n28480 , n28481 , n28482 , n28483 , n28484 , n28485 , n28486 , n28487 , n28488 , n28489 , n28490 , n28491 , n28492 , n28493 , n28494 , n28495 , n28496 , n28497 , n28498 , n28499 , n28500 , n28501 , n28502 , n28503 , n28504 , n28505 , n28506 , n28507 , n28508 , n28509 , n28510 , n28511 , n28512 , n28513 , n28514 , n28515 , n28516 , n28517 , n28518 , n28519 , n28520 , n28521 , n28522 , n28523 , n28524 , n28525 , n28526 , n28527 , n28528 , n28529 , n28530 , n28531 , n28532 , n28533 , n28534 , n28535 , n28536 , n28537 , n28538 , n28539 , n28540 , n28541 , n28542 , n28543 , n28544 , n28545 , n28546 , n28547 , n28548 , n28549 , n28550 , n28551 , n28552 , n28553 , n28554 , n28555 , n28556 , n28557 , n28558 , n28559 , n28560 , n28561 , n28562 , n28563 , n28564 , n28565 , n28566 , n28567 , n28568 , n28569 , n28570 , n28571 , n28572 , n28573 , n28574 , n28575 , n28576 , n28577 , n28578 , n28579 , n28580 , n28581 , n28582 , n28583 , n28584 , n28585 , n28586 , n28587 , n28588 , n28589 , n28590 , n28591 , n28592 , n28593 , n28594 , n28595 , n28596 , n28597 , n28598 , n28599 , n28600 , n28601 , n28602 , n28603 , n28604 , n28605 , n28606 , n28607 , n28608 , n28609 , n28610 , n28611 , n28612 , n28613 , n28614 , n28615 , n28616 , n28617 , n28618 , n28619 , n28620 , n28621 , n28622 , n28623 , n28624 , n28625 , n28626 , n28627 , n28628 , n28629 , n28630 , n28631 , n28632 , n28633 , n28634 , n28635 , n28636 , n28637 , n28638 , n28639 , n28640 , n28641 , n28642 , n28643 , n28644 , n28645 , n28646 , n28647 , n28648 , n28649 , n28650 , n28651 , n28652 , n28653 , n28654 , n28655 , n28656 , n28657 , n28658 , n28659 , n28660 , n28661 , n28662 , n28663 , n28664 , n28665 , n28666 , n28667 , n28668 , n28669 , n28670 , n28671 , n28672 , n28673 , n28674 , n28675 , n28676 , n28677 , n28678 , n28679 , n28680 , n28681 , n28682 , n28683 , n28684 , n28685 , n28686 , n28687 , n28688 , n28689 , n28690 , n28691 , n28692 , n28693 , n28694 , n28695 , n28696 , n28697 , n28698 , n28699 , n28700 , n28701 , n28702 , n28703 , n28704 , n28705 , n28706 , n28707 , n28708 , n28709 , n28710 , n28711 , n28712 , n28713 , n28714 , n28715 , n28716 , n28717 , n28718 , n28719 , n28720 , n28721 , n28722 , n28723 , n28724 , n28725 , n28726 , n28727 , n28728 , n28729 , n28730 , n28731 , n28732 , n28733 , n28734 , n28735 , n28736 , n28737 , n28738 , n28739 , n28740 , n28741 , n28742 , n28743 , n28744 , n28745 , n28746 , n28747 , n28748 , n28749 , n28750 , n28751 , n28752 , n28753 , n28754 , n28755 , n28756 , n28757 , n28758 , n28759 , n28760 , n28761 , n28762 , n28763 , n28764 , n28765 , n28766 , n28767 , n28768 , n28769 , n28770 , n28771 , n28772 , n28773 , n28774 , n28775 , n28776 , n28777 , n28778 , n28779 , n28780 , n28781 , n28782 , n28783 , n28784 , n28785 , n28786 , n28787 , n28788 , n28789 , n28790 , n28791 , n28792 , n28793 , n28794 , n28795 , n28796 , n28797 , n28798 , n28799 , n28800 , n28801 , n28802 , n28803 , n28804 , n28805 , n28806 , n28807 , n28808 , n28809 , n28810 , n28811 , n28812 , n28813 , n28814 , n28815 , n28816 , n28817 , n28818 , n28819 , n28820 , n28821 , n28822 , n28823 , n28824 , n28825 , n28826 , n28827 , n28828 , n28829 , n28830 , n28831 , n28832 , n28833 , n28834 , n28835 , n28836 , n28837 , n28838 , n28839 , n28840 , n28841 , n28842 , n28843 , n28844 , n28845 , n28846 , n28847 , n28848 , n28849 , n28850 , n28851 , n28852 , n28853 , n28854 , n28855 , n28856 , n28857 , n28858 , n28859 , n28860 , n28861 , n28862 , n28863 , n28864 , n28865 , n28866 , n28867 , n28868 , n28869 , n28870 , n28871 , n28872 , n28873 , n28874 , n28875 , n28876 , n28877 , n28878 , n28879 , n28880 , n28881 , n28882 , n28883 , n28884 , n28885 , n28886 , n28887 , n28888 , n28889 , n28890 , n28891 , n28892 , n28893 , n28894 , n28895 , n28896 , n28897 , n28898 , n28899 , n28900 , n28901 , n28902 , n28903 , n28904 , n28905 , n28906 , n28907 , n28908 , n28909 , n28910 , n28911 , n28912 , n28913 , n28914 , n28915 , n28916 , n28917 , n28918 , n28919 , n28920 , n28921 , n28922 , n28923 , n28924 , n28925 , n28926 , n28927 , n28928 , n28929 , n28930 , n28931 , n28932 , n28933 , n28934 , n28935 , n28936 , n28937 , n28938 , n28939 , n28940 , n28941 , n28942 , n28943 , n28944 , n28945 , n28946 , n28947 , n28948 , n28949 , n28950 , n28951 , n28952 , n28953 , n28954 , n28955 , n28956 , n28957 , n28958 , n28959 , n28960 , n28961 , n28962 , n28963 , n28964 , n28965 , n28966 , n28967 , n28968 , n28969 , n28970 , n28971 , n28972 , n28973 , n28974 , n28975 , n28976 , n28977 , n28978 , n28979 , n28980 , n28981 , n28982 , n28983 , n28984 , n28985 , n28986 , n28987 , n28988 , n28989 , n28990 , n28991 , n28992 , n28993 , n28994 , n28995 , n28996 , n28997 , n28998 , n28999 , n29000 , n29001 , n29002 , n29003 , n29004 , n29005 , n29006 , n29007 , n29008 , n29009 , n29010 , n29011 , n29012 , n29013 , n29014 , n29015 , n29016 , n29017 , n29018 , n29019 , n29020 , n29021 , n29022 , n29023 , n29024 , n29025 , n29026 , n29027 , n29028 , n29029 , n29030 , n29031 , n29032 , n29033 , n29034 , n29035 , n29036 , n29037 , n29038 , n29039 , n29040 , n29041 , n29042 , n29043 , n29044 , n29045 , n29046 , n29047 , n29048 , n29049 , n29050 , n29051 , n29052 , n29053 , n29054 , n29055 , n29056 , n29057 , n29058 , n29059 , n29060 , n29061 , n29062 , n29063 , n29064 , n29065 , n29066 , n29067 , n29068 , n29069 , n29070 , n29071 , n29072 , n29073 , n29074 , n29075 , n29076 , n29077 , n29078 , n29079 , n29080 , n29081 , n29082 , n29083 , n29084 , n29085 , n29086 , n29087 , n29088 , n29089 , n29090 , n29091 , n29092 , n29093 , n29094 , n29095 , n29096 , n29097 , n29098 , n29099 , n29100 , n29101 , n29102 , n29103 , n29104 , n29105 , n29106 , n29107 , n29108 , n29109 , n29110 , n29111 , n29112 , n29113 , n29114 , n29115 , n29116 , n29117 , n29118 , n29119 , n29120 , n29121 , n29122 , n29123 , n29124 , n29125 , n29126 , n29127 , n29128 , n29129 , n29130 , n29131 , n29132 , n29133 , n29134 , n29135 , n29136 , n29137 , n29138 , n29139 , n29140 , n29141 , n29142 , n29143 , n29144 , n29145 , n29146 , n29147 , n29148 , n29149 , n29150 , n29151 , n29152 , n29153 , n29154 , n29155 , n29156 , n29157 , n29158 , n29159 , n29160 , n29161 , n29162 , n29163 , n29164 , n29165 , n29166 , n29167 , n29168 , n29169 , n29170 , n29171 , n29172 , n29173 , n29174 , n29175 , n29176 , n29177 , n29178 , n29179 , n29180 , n29181 , n29182 , n29183 , n29184 , n29185 , n29186 , n29187 , n29188 , n29189 , n29190 , n29191 , n29192 , n29193 , n29194 , n29195 , n29196 , n29197 , n29198 , n29199 , n29200 , n29201 , n29202 , n29203 , n29204 , n29205 , n29206 , n29207 , n29208 , n29209 , n29210 , n29211 , n29212 , n29213 , n29214 , n29215 , n29216 , n29217 , n29218 , n29219 , n29220 , n29221 , n29222 , n29223 , n29224 , n29225 , n29226 , n29227 , n29228 , n29229 , n29230 , n29231 , n29232 , n29233 , n29234 , n29235 , n29236 , n29237 , n29238 , n29239 , n29240 , n29241 , n29242 , n29243 , n29244 , n29245 , n29246 , n29247 , n29248 , n29249 , n29250 , n29251 , n29252 , n29253 , n29254 , n29255 , n29256 , n29257 , n29258 , n29259 , n29260 , n29261 , n29262 , n29263 , n29264 , n29265 , n29266 , n29267 , n29268 , n29269 , n29270 , n29271 , n29272 , n29273 , n29274 , n29275 , n29276 , n29277 , n29278 , n29279 , n29280 , n29281 , n29282 , n29283 , n29284 , n29285 , n29286 , n29287 , n29288 , n29289 , n29290 , n29291 , n29292 , n29293 , n29294 , n29295 , n29296 , n29297 , n29298 , n29299 , n29300 , n29301 , n29302 , n29303 , n29304 , n29305 , n29306 , n29307 , n29308 , n29309 , n29310 , n29311 , n29312 , n29313 , n29314 , n29315 , n29316 , n29317 , n29318 , n29319 , n29320 , n29321 , n29322 , n29323 , n29324 , n29325 , n29326 , n29327 , n29328 , n29329 , n29330 , n29331 , n29332 , n29333 , n29334 , n29335 , n29336 , n29337 , n29338 , n29339 , n29340 , n29341 , n29342 , n29343 , n29344 , n29345 , n29346 , n29347 , n29348 , n29349 , n29350 , n29351 , n29352 , n29353 , n29354 , n29355 , n29356 , n29357 , n29358 , n29359 , n29360 , n29361 , n29362 , n29363 , n29364 , n29365 , n29366 , n29367 , n29368 , n29369 , n29370 , n29371 , n29372 , n29373 , n29374 , n29375 , n29376 , n29377 , n29378 , n29379 , n29380 , n29381 , n29382 , n29383 , n29384 , n29385 , n29386 , n29387 , n29388 , n29389 , n29390 , n29391 , n29392 , n29393 , n29394 , n29395 , n29396 , n29397 , n29398 , n29399 , n29400 , n29401 , n29402 , n29403 , n29404 , n29405 , n29406 , n29407 , n29408 , n29409 , n29410 , n29411 , n29412 , n29413 , n29414 , n29415 , n29416 , n29417 , n29418 , n29419 , n29420 , n29421 , n29422 , n29423 , n29424 , n29425 , n29426 , n29427 , n29428 , n29429 , n29430 , n29431 , n29432 , n29433 , n29434 , n29435 , n29436 , n29437 , n29438 , n29439 , n29440 , n29441 , n29442 , n29443 , n29444 , n29445 , n29446 , n29447 , n29448 , n29449 , n29450 , n29451 , n29452 , n29453 , n29454 , n29455 , n29456 , n29457 , n29458 , n29459 , n29460 , n29461 , n29462 , n29463 , n29464 , n29465 , n29466 , n29467 , n29468 , n29469 , n29470 , n29471 , n29472 , n29473 , n29474 , n29475 , n29476 , n29477 , n29478 , n29479 , n29480 , n29481 , n29482 , n29483 , n29484 , n29485 , n29486 , n29487 , n29488 , n29489 , n29490 , n29491 , n29492 , n29493 , n29494 , n29495 , n29496 , n29497 , n29498 , n29499 , n29500 , n29501 , n29502 , n29503 , n29504 , n29505 , n29506 , n29507 , n29508 , n29509 , n29510 , n29511 , n29512 , n29513 , n29514 , n29515 , n29516 , n29517 , n29518 , n29519 , n29520 , n29521 , n29522 , n29523 , n29524 , n29525 , n29526 , n29527 , n29528 , n29529 , n29530 , n29531 , n29532 , n29533 , n29534 , n29535 , n29536 , n29537 , n29538 , n29539 , n29540 , n29541 , n29542 , n29543 , n29544 , n29545 , n29546 , n29547 , n29548 , n29549 , n29550 , n29551 , n29552 , n29553 , n29554 , n29555 , n29556 , n29557 , n29558 , n29559 , n29560 , n29561 , n29562 , n29563 , n29564 , n29565 , n29566 , n29567 , n29568 , n29569 , n29570 , n29571 , n29572 , n29573 , n29574 , n29575 , n29576 , n29577 , n29578 , n29579 , n29580 , n29581 , n29582 , n29583 , n29584 , n29585 , n29586 , n29587 , n29588 , n29589 , n29590 , n29591 , n29592 , n29593 , n29594 , n29595 , n29596 , n29597 , n29598 , n29599 , n29600 , n29601 , n29602 , n29603 , n29604 , n29605 , n29606 , n29607 , n29608 , n29609 , n29610 , n29611 , n29612 , n29613 , n29614 , n29615 , n29616 , n29617 , n29618 , n29619 , n29620 , n29621 , n29622 , n29623 , n29624 , n29625 , n29626 , n29627 , n29628 , n29629 , n29630 , n29631 , n29632 , n29633 , n29634 , n29635 , n29636 , n29637 , n29638 , n29639 , n29640 , n29641 , n29642 , n29643 , n29644 , n29645 , n29646 , n29647 , n29648 , n29649 , n29650 , n29651 , n29652 , n29653 , n29654 , n29655 , n29656 , n29657 , n29658 , n29659 , n29660 , n29661 , n29662 , n29663 , n29664 , n29665 , n29666 , n29667 , n29668 , n29669 , n29670 , n29671 , n29672 , n29673 , n29674 , n29675 , n29676 , n29677 , n29678 , n29679 , n29680 , n29681 , n29682 , n29683 , n29684 , n29685 , n29686 , n29687 , n29688 , n29689 , n29690 , n29691 , n29692 , n29693 , n29694 , n29695 , n29696 , n29697 , n29698 , n29699 , n29700 , n29701 , n29702 , n29703 , n29704 , n29705 , n29706 , n29707 , n29708 , n29709 , n29710 , n29711 , n29712 , n29713 , n29714 , n29715 , n29716 , n29717 , n29718 , n29719 , n29720 , n29721 , n29722 , n29723 , n29724 , n29725 , n29726 , n29727 , n29728 , n29729 , n29730 , n29731 , n29732 , n29733 , n29734 , n29735 , n29736 , n29737 , n29738 , n29739 , n29740 , n29741 , n29742 , n29743 , n29744 , n29745 , n29746 , n29747 , n29748 , n29749 , n29750 , n29751 , n29752 , n29753 , n29754 , n29755 , n29756 , n29757 , n29758 , n29759 , n29760 , n29761 , n29762 , n29763 , n29764 , n29765 , n29766 , n29767 , n29768 , n29769 , n29770 , n29771 , n29772 , n29773 , n29774 , n29775 , n29776 , n29777 , n29778 , n29779 , n29780 , n29781 , n29782 , n29783 , n29784 , n29785 , n29786 , n29787 , n29788 , n29789 , n29790 , n29791 , n29792 , n29793 , n29794 , n29795 , n29796 , n29797 , n29798 , n29799 , n29800 , n29801 , n29802 , n29803 , n29804 , n29805 , n29806 , n29807 , n29808 , n29809 , n29810 , n29811 , n29812 , n29813 , n29814 , n29815 , n29816 , n29817 , n29818 , n29819 , n29820 , n29821 , n29822 , n29823 , n29824 , n29825 , n29826 , n29827 , n29828 , n29829 , n29830 , n29831 , n29832 , n29833 , n29834 , n29835 , n29836 , n29837 , n29838 , n29839 , n29840 , n29841 , n29842 , n29843 , n29844 , n29845 , n29846 , n29847 , n29848 , n29849 , n29850 , n29851 , n29852 , n29853 , n29854 , n29855 , n29856 , n29857 , n29858 , n29859 , n29860 , n29861 , n29862 , n29863 , n29864 , n29865 , n29866 , n29867 , n29868 , n29869 , n29870 , n29871 , n29872 , n29873 , n29874 , n29875 , n29876 , n29877 , n29878 , n29879 , n29880 , n29881 , n29882 , n29883 , n29884 , n29885 , n29886 , n29887 , n29888 , n29889 , n29890 , n29891 , n29892 , n29893 , n29894 , n29895 , n29896 , n29897 , n29898 , n29899 , n29900 , n29901 , n29902 , n29903 , n29904 , n29905 , n29906 , n29907 , n29908 , n29909 , n29910 , n29911 , n29912 , n29913 , n29914 , n29915 , n29916 , n29917 , n29918 , n29919 , n29920 , n29921 , n29922 , n29923 , n29924 , n29925 , n29926 , n29927 , n29928 , n29929 , n29930 , n29931 , n29932 , n29933 , n29934 , n29935 , n29936 , n29937 , n29938 , n29939 , n29940 , n29941 , n29942 , n29943 , n29944 , n29945 , n29946 , n29947 , n29948 , n29949 , n29950 , n29951 , n29952 , n29953 , n29954 , n29955 , n29956 , n29957 , n29958 , n29959 , n29960 , n29961 , n29962 , n29963 , n29964 , n29965 , n29966 , n29967 , n29968 , n29969 , n29970 , n29971 , n29972 , n29973 , n29974 , n29975 , n29976 , n29977 , n29978 , n29979 , n29980 , n29981 , n29982 , n29983 , n29984 , n29985 , n29986 , n29987 , n29988 , n29989 , n29990 , n29991 , n29992 , n29993 , n29994 , n29995 , n29996 , n29997 , n29998 , n29999 , n30000 , n30001 , n30002 , n30003 , n30004 , n30005 , n30006 , n30007 , n30008 , n30009 , n30010 , n30011 , n30012 , n30013 , n30014 , n30015 , n30016 , n30017 , n30018 , n30019 , n30020 , n30021 , n30022 , n30023 , n30024 , n30025 , n30026 , n30027 , n30028 , n30029 , n30030 , n30031 , n30032 , n30033 , n30034 , n30035 , n30036 , n30037 , n30038 , n30039 , n30040 , n30041 , n30042 , n30043 , n30044 , n30045 , n30046 , n30047 , n30048 , n30049 , n30050 , n30051 , n30052 , n30053 , n30054 , n30055 , n30056 , n30057 , n30058 , n30059 , n30060 , n30061 , n30062 , n30063 , n30064 , n30065 , n30066 , n30067 , n30068 , n30069 , n30070 , n30071 , n30072 , n30073 , n30074 , n30075 , n30076 , n30077 , n30078 , n30079 , n30080 , n30081 , n30082 , n30083 , n30084 , n30085 , n30086 , n30087 , n30088 , n30089 , n30090 , n30091 , n30092 , n30093 , n30094 , n30095 , n30096 , n30097 , n30098 , n30099 , n30100 , n30101 , n30102 , n30103 , n30104 , n30105 , n30106 , n30107 , n30108 , n30109 , n30110 , n30111 , n30112 , n30113 , n30114 , n30115 , n30116 , n30117 , n30118 , n30119 , n30120 , n30121 , n30122 , n30123 , n30124 , n30125 , n30126 , n30127 , n30128 , n30129 , n30130 , n30131 , n30132 , n30133 , n30134 , n30135 , n30136 , n30137 , n30138 , n30139 , n30140 , n30141 , n30142 , n30143 , n30144 , n30145 , n30146 , n30147 , n30148 , n30149 , n30150 , n30151 , n30152 , n30153 , n30154 , n30155 , n30156 , n30157 , n30158 , n30159 , n30160 , n30161 , n30162 , n30163 , n30164 , n30165 , n30166 , n30167 , n30168 , n30169 , n30170 , n30171 , n30172 , n30173 , n30174 , n30175 , n30176 , n30177 , n30178 , n30179 , n30180 , n30181 , n30182 , n30183 , n30184 , n30185 , n30186 , n30187 , n30188 , n30189 , n30190 , n30191 , n30192 , n30193 , n30194 , n30195 , n30196 , n30197 , n30198 , n30199 , n30200 , n30201 , n30202 , n30203 , n30204 , n30205 , n30206 , n30207 , n30208 , n30209 , n30210 , n30211 , n30212 , n30213 , n30214 , n30215 , n30216 , n30217 , n30218 , n30219 , n30220 , n30221 , n30222 , n30223 , n30224 , n30225 , n30226 , n30227 , n30228 , n30229 , n30230 , n30231 , n30232 , n30233 , n30234 , n30235 , n30236 , n30237 , n30238 , n30239 , n30240 , n30241 , n30242 , n30243 , n30244 , n30245 , n30246 , n30247 , n30248 , n30249 , n30250 , n30251 , n30252 , n30253 , n30254 , n30255 , n30256 , n30257 , n30258 , n30259 , n30260 , n30261 , n30262 , n30263 , n30264 , n30265 , n30266 , n30267 , n30268 , n30269 , n30270 , n30271 , n30272 , n30273 , n30274 , n30275 , n30276 , n30277 , n30278 , n30279 , n30280 , n30281 , n30282 , n30283 , n30284 , n30285 , n30286 , n30287 , n30288 , n30289 , n30290 , n30291 , n30292 , n30293 , n30294 , n30295 , n30296 , n30297 , n30298 , n30299 , n30300 , n30301 , n30302 , n30303 , n30304 , n30305 , n30306 , n30307 , n30308 , n30309 , n30310 , n30311 , n30312 , n30313 , n30314 , n30315 , n30316 , n30317 , n30318 , n30319 , n30320 , n30321 , n30322 , n30323 , n30324 , n30325 , n30326 , n30327 , n30328 , n30329 , n30330 , n30331 , n30332 , n30333 , n30334 , n30335 , n30336 , n30337 , n30338 , n30339 , n30340 , n30341 , n30342 , n30343 , n30344 , n30345 , n30346 , n30347 , n30348 , n30349 , n30350 , n30351 , n30352 , n30353 , n30354 , n30355 , n30356 , n30357 , n30358 , n30359 , n30360 , n30361 , n30362 , n30363 , n30364 , n30365 , n30366 , n30367 , n30368 , n30369 , n30370 , n30371 , n30372 , n30373 , n30374 , n30375 , n30376 , n30377 , n30378 , n30379 , n30380 , n30381 , n30382 , n30383 , n30384 , n30385 , n30386 , n30387 , n30388 , n30389 , n30390 , n30391 , n30392 , n30393 , n30394 , n30395 , n30396 , n30397 , n30398 , n30399 , n30400 , n30401 , n30402 , n30403 , n30404 , n30405 , n30406 , n30407 , n30408 , n30409 , n30410 , n30411 , n30412 , n30413 , n30414 , n30415 , n30416 , n30417 , n30418 , n30419 , n30420 , n30421 , n30422 , n30423 , n30424 , n30425 , n30426 , n30427 , n30428 , n30429 , n30430 , n30431 , n30432 , n30433 , n30434 , n30435 , n30436 , n30437 , n30438 , n30439 , n30440 , n30441 , n30442 , n30443 , n30444 , n30445 , n30446 , n30447 , n30448 , n30449 , n30450 , n30451 , n30452 , n30453 , n30454 , n30455 , n30456 , n30457 , n30458 , n30459 , n30460 , n30461 , n30462 , n30463 , n30464 , n30465 , n30466 , n30467 , n30468 , n30469 , n30470 , n30471 , n30472 , n30473 , n30474 , n30475 , n30476 , n30477 , n30478 , n30479 , n30480 , n30481 , n30482 , n30483 , n30484 , n30485 , n30486 , n30487 , n30488 , n30489 , n30490 , n30491 , n30492 , n30493 , n30494 , n30495 , n30496 , n30497 , n30498 , n30499 , n30500 , n30501 , n30502 , n30503 , n30504 , n30505 , n30506 , n30507 , n30508 , n30509 , n30510 , n30511 , n30512 , n30513 , n30514 , n30515 , n30516 , n30517 , n30518 , n30519 , n30520 , n30521 , n30522 , n30523 , n30524 , n30525 , n30526 , n30527 , n30528 , n30529 , n30530 , n30531 , n30532 , n30533 , n30534 , n30535 , n30536 , n30537 , n30538 , n30539 , n30540 , n30541 , n30542 , n30543 , n30544 , n30545 , n30546 , n30547 , n30548 , n30549 , n30550 , n30551 , n30552 , n30553 , n30554 , n30555 , n30556 , n30557 , n30558 , n30559 , n30560 , n30561 , n30562 , n30563 , n30564 , n30565 , n30566 , n30567 , n30568 , n30569 , n30570 , n30571 , n30572 , n30573 , n30574 , n30575 , n30576 , n30577 , n30578 , n30579 , n30580 , n30581 , n30582 , n30583 , n30584 , n30585 , n30586 , n30587 , n30588 , n30589 , n30590 , n30591 , n30592 , n30593 , n30594 , n30595 , n30596 , n30597 , n30598 , n30599 , n30600 , n30601 , n30602 , n30603 , n30604 , n30605 , n30606 , n30607 , n30608 , n30609 , n30610 , n30611 , n30612 , n30613 , n30614 , n30615 , n30616 , n30617 , n30618 , n30619 , n30620 , n30621 , n30622 , n30623 , n30624 , n30625 , n30626 , n30627 , n30628 , n30629 , n30630 , n30631 , n30632 , n30633 , n30634 , n30635 , n30636 , n30637 , n30638 , n30639 , n30640 , n30641 , n30642 , n30643 , n30644 , n30645 , n30646 , n30647 , n30648 , n30649 , n30650 , n30651 , n30652 , n30653 , n30654 , n30655 , n30656 , n30657 , n30658 , n30659 , n30660 , n30661 , n30662 , n30663 , n30664 , n30665 , n30666 , n30667 , n30668 , n30669 , n30670 , n30671 , n30672 , n30673 , n30674 , n30675 , n30676 , n30677 , n30678 , n30679 , n30680 , n30681 , n30682 , n30683 , n30684 , n30685 , n30686 , n30687 , n30688 , n30689 , n30690 , n30691 , n30692 , n30693 , n30694 , n30695 , n30696 , n30697 , n30698 , n30699 , n30700 , n30701 , n30702 , n30703 , n30704 , n30705 , n30706 , n30707 , n30708 , n30709 , n30710 , n30711 , n30712 , n30713 , n30714 , n30715 , n30716 , n30717 , n30718 , n30719 , n30720 , n30721 , n30722 , n30723 , n30724 , n30725 , n30726 , n30727 , n30728 , n30729 , n30730 , n30731 , n30732 , n30733 , n30734 , n30735 , n30736 , n30737 , n30738 , n30739 , n30740 , n30741 , n30742 , n30743 , n30744 , n30745 , n30746 , n30747 , n30748 , n30749 , n30750 , n30751 , n30752 , n30753 , n30754 , n30755 , n30756 , n30757 , n30758 , n30759 , n30760 , n30761 , n30762 , n30763 , n30764 , n30765 , n30766 , n30767 , n30768 , n30769 , n30770 , n30771 , n30772 , n30773 , n30774 , n30775 , n30776 , n30777 , n30778 , n30779 , n30780 , n30781 , n30782 , n30783 , n30784 , n30785 , n30786 , n30787 , n30788 , n30789 , n30790 , n30791 , n30792 , n30793 , n30794 , n30795 , n30796 , n30797 , n30798 , n30799 , n30800 , n30801 , n30802 , n30803 , n30804 , n30805 , n30806 , n30807 , n30808 , n30809 , n30810 , n30811 , n30812 , n30813 , n30814 , n30815 , n30816 , n30817 , n30818 , n30819 , n30820 , n30821 , n30822 , n30823 , n30824 , n30825 , n30826 , n30827 , n30828 , n30829 , n30830 , n30831 , n30832 , n30833 , n30834 , n30835 , n30836 , n30837 , n30838 , n30839 , n30840 , n30841 , n30842 , n30843 , n30844 , n30845 , n30846 , n30847 , n30848 , n30849 , n30850 , n30851 , n30852 , n30853 , n30854 , n30855 , n30856 , n30857 , n30858 , n30859 , n30860 , n30861 , n30862 , n30863 , n30864 , n30865 , n30866 , n30867 , n30868 , n30869 , n30870 , n30871 , n30872 , n30873 , n30874 , n30875 , n30876 , n30877 , n30878 , n30879 , n30880 , n30881 , n30882 , n30883 , n30884 , n30885 , n30886 , n30887 , n30888 , n30889 , n30890 , n30891 , n30892 , n30893 , n30894 , n30895 , n30896 , n30897 , n30898 , n30899 , n30900 , n30901 , n30902 , n30903 , n30904 , n30905 , n30906 , n30907 , n30908 , n30909 , n30910 , n30911 , n30912 , n30913 , n30914 , n30915 , n30916 , n30917 , n30918 , n30919 , n30920 , n30921 , n30922 , n30923 , n30924 , n30925 , n30926 , n30927 , n30928 , n30929 , n30930 , n30931 , n30932 , n30933 , n30934 , n30935 , n30936 , n30937 , n30938 , n30939 , n30940 , n30941 , n30942 , n30943 , n30944 , n30945 , n30946 , n30947 , n30948 , n30949 , n30950 , n30951 , n30952 , n30953 , n30954 , n30955 , n30956 , n30957 , n30958 , n30959 , n30960 , n30961 , n30962 , n30963 , n30964 , n30965 , n30966 , n30967 , n30968 , n30969 , n30970 , n30971 , n30972 , n30973 , n30974 , n30975 , n30976 , n30977 , n30978 , n30979 , n30980 , n30981 , n30982 , n30983 , n30984 , n30985 , n30986 , n30987 , n30988 , n30989 , n30990 , n30991 , n30992 , n30993 , n30994 , n30995 , n30996 , n30997 , n30998 , n30999 , n31000 , n31001 , n31002 , n31003 , n31004 , n31005 , n31006 , n31007 , n31008 , n31009 , n31010 , n31011 , n31012 , n31013 , n31014 , n31015 , n31016 , n31017 , n31018 , n31019 , n31020 , n31021 , n31022 , n31023 , n31024 , n31025 , n31026 , n31027 , n31028 , n31029 , n31030 , n31031 , n31032 , n31033 , n31034 , n31035 , n31036 , n31037 , n31038 , n31039 , n31040 , n31041 , n31042 , n31043 , n31044 , n31045 , n31046 , n31047 , n31048 , n31049 , n31050 , n31051 , n31052 , n31053 , n31054 , n31055 , n31056 , n31057 , n31058 , n31059 , n31060 , n31061 , n31062 , n31063 , n31064 , n31065 , n31066 , n31067 , n31068 , n31069 , n31070 , n31071 , n31072 , n31073 , n31074 , n31075 , n31076 , n31077 , n31078 , n31079 , n31080 , n31081 , n31082 , n31083 , n31084 , n31085 , n31086 , n31087 , n31088 , n31089 , n31090 , n31091 , n31092 , n31093 , n31094 , n31095 , n31096 , n31097 , n31098 , n31099 , n31100 , n31101 , n31102 , n31103 , n31104 , n31105 , n31106 , n31107 , n31108 , n31109 , n31110 , n31111 , n31112 , n31113 , n31114 , n31115 , n31116 , n31117 , n31118 , n31119 , n31120 , n31121 , n31122 , n31123 , n31124 , n31125 , n31126 , n31127 , n31128 , n31129 , n31130 , n31131 , n31132 , n31133 , n31134 , n31135 , n31136 , n31137 , n31138 , n31139 , n31140 , n31141 , n31142 , n31143 , n31144 , n31145 , n31146 , n31147 , n31148 , n31149 , n31150 , n31151 , n31152 , n31153 , n31154 , n31155 , n31156 , n31157 , n31158 , n31159 , n31160 , n31161 , n31162 , n31163 , n31164 , n31165 , n31166 , n31167 , n31168 , n31169 , n31170 , n31171 , n31172 , n31173 , n31174 , n31175 , n31176 , n31177 , n31178 , n31179 , n31180 , n31181 , n31182 , n31183 , n31184 , n31185 , n31186 , n31187 , n31188 , n31189 , n31190 , n31191 , n31192 , n31193 , n31194 , n31195 , n31196 , n31197 , n31198 , n31199 , n31200 , n31201 , n31202 , n31203 , n31204 , n31205 , n31206 , n31207 , n31208 , n31209 , n31210 , n31211 , n31212 , n31213 , n31214 , n31215 , n31216 , n31217 , n31218 , n31219 , n31220 , n31221 , n31222 , n31223 , n31224 , n31225 , n31226 , n31227 , n31228 , n31229 , n31230 , n31231 , n31232 , n31233 , n31234 , n31235 , n31236 , n31237 , n31238 , n31239 , n31240 , n31241 , n31242 , n31243 , n31244 , n31245 , n31246 , n31247 , n31248 , n31249 , n31250 , n31251 , n31252 , n31253 , n31254 , n31255 , n31256 , n31257 , n31258 , n31259 , n31260 , n31261 , n31262 , n31263 , n31264 , n31265 , n31266 , n31267 , n31268 , n31269 , n31270 , n31271 , n31272 , n31273 , n31274 , n31275 , n31276 , n31277 , n31278 , n31279 , n31280 , n31281 , n31282 , n31283 , n31284 , n31285 , n31286 , n31287 , n31288 , n31289 , n31290 , n31291 , n31292 , n31293 , n31294 , n31295 , n31296 , n31297 , n31298 , n31299 , n31300 , n31301 , n31302 , n31303 , n31304 , n31305 , n31306 , n31307 , n31308 , n31309 , n31310 , n31311 , n31312 , n31313 , n31314 , n31315 , n31316 , n31317 , n31318 , n31319 , n31320 , n31321 , n31322 , n31323 , n31324 , n31325 , n31326 , n31327 , n31328 , n31329 , n31330 , n31331 , n31332 , n31333 , n31334 , n31335 , n31336 , n31337 , n31338 , n31339 , n31340 , n31341 , n31342 , n31343 , n31344 , n31345 , n31346 , n31347 , n31348 , n31349 , n31350 , n31351 , n31352 , n31353 , n31354 , n31355 , n31356 , n31357 , n31358 , n31359 , n31360 , n31361 , n31362 , n31363 , n31364 , n31365 , n31366 , n31367 , n31368 , n31369 , n31370 , n31371 , n31372 , n31373 , n31374 , n31375 , n31376 , n31377 , n31378 , n31379 , n31380 , n31381 , n31382 , n31383 , n31384 , n31385 , n31386 , n31387 , n31388 , n31389 , n31390 , n31391 , n31392 , n31393 , n31394 , n31395 , n31396 , n31397 , n31398 , n31399 , n31400 , n31401 , n31402 , n31403 , n31404 , n31405 , n31406 , n31407 , n31408 , n31409 , n31410 , n31411 , n31412 , n31413 , n31414 , n31415 , n31416 , n31417 , n31418 , n31419 , n31420 , n31421 , n31422 , n31423 , n31424 , n31425 , n31426 , n31427 , n31428 , n31429 , n31430 , n31431 , n31432 , n31433 , n31434 , n31435 , n31436 , n31437 , n31438 , n31439 , n31440 , n31441 , n31442 , n31443 , n31444 , n31445 , n31446 , n31447 , n31448 , n31449 , n31450 , n31451 , n31452 , n31453 , n31454 , n31455 , n31456 , n31457 , n31458 , n31459 , n31460 , n31461 , n31462 , n31463 , n31464 , n31465 , n31466 , n31467 , n31468 , n31469 , n31470 , n31471 , n31472 , n31473 , n31474 , n31475 , n31476 , n31477 , n31478 , n31479 , n31480 , n31481 , n31482 , n31483 , n31484 , n31485 , n31486 , n31487 , n31488 , n31489 , n31490 , n31491 , n31492 , n31493 , n31494 , n31495 , n31496 , n31497 , n31498 , n31499 , n31500 , n31501 , n31502 , n31503 , n31504 , n31505 , n31506 , n31507 , n31508 , n31509 , n31510 , n31511 , n31512 , n31513 , n31514 , n31515 , n31516 , n31517 , n31518 , n31519 , n31520 , n31521 , n31522 , n31523 , n31524 , n31525 , n31526 , n31527 , n31528 , n31529 , n31530 , n31531 , n31532 , n31533 , n31534 , n31535 , n31536 , n31537 , n31538 , n31539 , n31540 , n31541 , n31542 , n31543 , n31544 , n31545 , n31546 , n31547 , n31548 , n31549 , n31550 , n31551 , n31552 , n31553 , n31554 , n31555 , n31556 , n31557 , n31558 , n31559 , n31560 , n31561 , n31562 , n31563 , n31564 , n31565 , n31566 , n31567 , n31568 , n31569 , n31570 , n31571 , n31572 , n31573 , n31574 , n31575 , n31576 , n31577 , n31578 , n31579 , n31580 , n31581 , n31582 , n31583 , n31584 , n31585 , n31586 , n31587 , n31588 , n31589 , n31590 , n31591 , n31592 , n31593 , n31594 , n31595 , n31596 , n31597 , n31598 , n31599 , n31600 , n31601 , n31602 , n31603 , n31604 , n31605 , n31606 , n31607 , n31608 , n31609 , n31610 , n31611 , n31612 , n31613 , n31614 , n31615 , n31616 , n31617 , n31618 , n31619 , n31620 , n31621 , n31622 , n31623 , n31624 , n31625 , n31626 , n31627 , n31628 , n31629 , n31630 , n31631 , n31632 , n31633 , n31634 , n31635 , n31636 , n31637 , n31638 , n31639 , n31640 , n31641 , n31642 , n31643 , n31644 , n31645 , n31646 , n31647 , n31648 , n31649 , n31650 , n31651 , n31652 , n31653 , n31654 , n31655 , n31656 , n31657 , n31658 , n31659 , n31660 , n31661 , n31662 , n31663 , n31664 , n31665 , n31666 , n31667 , n31668 , n31669 , n31670 , n31671 , n31672 , n31673 , n31674 , n31675 , n31676 , n31677 , n31678 , n31679 , n31680 , n31681 , n31682 , n31683 , n31684 , n31685 , n31686 , n31687 , n31688 , n31689 , n31690 , n31691 , n31692 , n31693 , n31694 , n31695 , n31696 , n31697 , n31698 , n31699 , n31700 , n31701 , n31702 , n31703 , n31704 , n31705 , n31706 , n31707 , n31708 , n31709 , n31710 , n31711 , n31712 , n31713 , n31714 , n31715 , n31716 , n31717 , n31718 , n31719 , n31720 , n31721 , n31722 , n31723 , n31724 , n31725 , n31726 , n31727 , n31728 , n31729 , n31730 , n31731 , n31732 , n31733 , n31734 , n31735 , n31736 , n31737 , n31738 , n31739 , n31740 , n31741 , n31742 , n31743 , n31744 , n31745 , n31746 , n31747 , n31748 , n31749 , n31750 , n31751 , n31752 , n31753 , n31754 , n31755 , n31756 , n31757 , n31758 , n31759 , n31760 , n31761 , n31762 , n31763 , n31764 , n31765 , n31766 , n31767 , n31768 , n31769 , n31770 , n31771 , n31772 , n31773 , n31774 , n31775 , n31776 , n31777 , n31778 , n31779 , n31780 , n31781 , n31782 , n31783 , n31784 , n31785 , n31786 , n31787 , n31788 , n31789 , n31790 , n31791 , n31792 , n31793 , n31794 , n31795 , n31796 , n31797 , n31798 , n31799 , n31800 , n31801 , n31802 , n31803 , n31804 , n31805 , n31806 , n31807 , n31808 , n31809 , n31810 , n31811 , n31812 , n31813 , n31814 , n31815 , n31816 , n31817 , n31818 , n31819 , n31820 , n31821 , n31822 , n31823 , n31824 , n31825 , n31826 , n31827 , n31828 , n31829 , n31830 , n31831 , n31832 , n31833 , n31834 , n31835 , n31836 , n31837 , n31838 , n31839 , n31840 , n31841 , n31842 , n31843 , n31844 , n31845 , n31846 , n31847 , n31848 , n31849 , n31850 , n31851 , n31852 , n31853 , n31854 , n31855 , n31856 , n31857 , n31858 , n31859 , n31860 , n31861 , n31862 , n31863 , n31864 , n31865 , n31866 , n31867 , n31868 , n31869 , n31870 , n31871 , n31872 , n31873 , n31874 , n31875 , n31876 , n31877 , n31878 , n31879 , n31880 , n31881 , n31882 , n31883 , n31884 , n31885 , n31886 , n31887 , n31888 , n31889 , n31890 , n31891 , n31892 , n31893 , n31894 , n31895 , n31896 , n31897 , n31898 , n31899 , n31900 , n31901 , n31902 , n31903 , n31904 , n31905 , n31906 , n31907 , n31908 , n31909 , n31910 , n31911 , n31912 , n31913 , n31914 , n31915 , n31916 , n31917 , n31918 , n31919 , n31920 , n31921 , n31922 , n31923 , n31924 , n31925 , n31926 , n31927 , n31928 , n31929 , n31930 , n31931 , n31932 , n31933 , n31934 , n31935 , n31936 , n31937 , n31938 , n31939 , n31940 , n31941 , n31942 , n31943 , n31944 , n31945 , n31946 , n31947 , n31948 , n31949 , n31950 , n31951 , n31952 , n31953 , n31954 , n31955 , n31956 , n31957 , n31958 , n31959 , n31960 , n31961 , n31962 , n31963 , n31964 , n31965 , n31966 , n31967 , n31968 , n31969 , n31970 , n31971 , n31972 , n31973 , n31974 , n31975 , n31976 , n31977 , n31978 , n31979 , n31980 , n31981 , n31982 , n31983 , n31984 , n31985 , n31986 , n31987 , n31988 , n31989 , n31990 , n31991 , n31992 , n31993 , n31994 , n31995 , n31996 , n31997 , n31998 , n31999 , n32000 , n32001 , n32002 , n32003 , n32004 , n32005 , n32006 , n32007 , n32008 , n32009 , n32010 , n32011 , n32012 , n32013 , n32014 , n32015 , n32016 , n32017 , n32018 , n32019 , n32020 , n32021 , n32022 , n32023 , n32024 , n32025 , n32026 , n32027 , n32028 , n32029 , n32030 , n32031 , n32032 , n32033 , n32034 , n32035 , n32036 , n32037 , n32038 , n32039 , n32040 , n32041 , n32042 , n32043 , n32044 , n32045 , n32046 , n32047 , n32048 , n32049 , n32050 , n32051 , n32052 , n32053 , n32054 , n32055 , n32056 , n32057 , n32058 , n32059 , n32060 , n32061 , n32062 , n32063 , n32064 , n32065 , n32066 , n32067 , n32068 , n32069 , n32070 , n32071 , n32072 , n32073 , n32074 , n32075 , n32076 , n32077 , n32078 , n32079 , n32080 , n32081 , n32082 , n32083 , n32084 , n32085 , n32086 , n32087 , n32088 , n32089 , n32090 , n32091 , n32092 , n32093 , n32094 , n32095 , n32096 , n32097 , n32098 , n32099 , n32100 , n32101 , n32102 , n32103 , n32104 , n32105 , n32106 , n32107 , n32108 , n32109 , n32110 , n32111 , n32112 , n32113 , n32114 , n32115 , n32116 , n32117 , n32118 , n32119 , n32120 , n32121 , n32122 , n32123 , n32124 , n32125 , n32126 , n32127 , n32128 , n32129 , n32130 , n32131 , n32132 , n32133 , n32134 , n32135 , n32136 , n32137 , n32138 , n32139 , n32140 , n32141 , n32142 , n32143 , n32144 , n32145 , n32146 , n32147 , n32148 , n32149 , n32150 , n32151 , n32152 , n32153 , n32154 , n32155 , n32156 , n32157 , n32158 , n32159 , n32160 , n32161 , n32162 , n32163 , n32164 , n32165 , n32166 , n32167 , n32168 , n32169 , n32170 , n32171 , n32172 , n32173 , n32174 , n32175 , n32176 , n32177 , n32178 , n32179 , n32180 , n32181 , n32182 , n32183 , n32184 , n32185 , n32186 , n32187 , n32188 , n32189 , n32190 , n32191 , n32192 , n32193 , n32194 , n32195 , n32196 , n32197 , n32198 , n32199 , n32200 , n32201 , n32202 , n32203 , n32204 , n32205 , n32206 , n32207 , n32208 , n32209 , n32210 , n32211 , n32212 , n32213 , n32214 , n32215 , n32216 , n32217 , n32218 , n32219 , n32220 , n32221 , n32222 , n32223 , n32224 , n32225 , n32226 , n32227 , n32228 , n32229 , n32230 , n32231 , n32232 , n32233 , n32234 , n32235 , n32236 , n32237 , n32238 , n32239 , n32240 , n32241 , n32242 , n32243 , n32244 , n32245 , n32246 , n32247 , n32248 , n32249 , n32250 , n32251 , n32252 , n32253 , n32254 , n32255 , n32256 , n32257 , n32258 , n32259 , n32260 , n32261 , n32262 , n32263 , n32264 , n32265 , n32266 , n32267 , n32268 , n32269 , n32270 , n32271 , n32272 , n32273 , n32274 , n32275 , n32276 , n32277 , n32278 , n32279 , n32280 , n32281 , n32282 , n32283 , n32284 , n32285 , n32286 , n32287 , n32288 , n32289 , n32290 , n32291 , n32292 , n32293 , n32294 , n32295 , n32296 , n32297 , n32298 , n32299 , n32300 , n32301 , n32302 , n32303 , n32304 , n32305 , n32306 , n32307 , n32308 , n32309 , n32310 , n32311 , n32312 , n32313 , n32314 , n32315 , n32316 , n32317 , n32318 , n32319 , n32320 , n32321 , n32322 , n32323 , n32324 , n32325 , n32326 , n32327 , n32328 , n32329 , n32330 , n32331 , n32332 , n32333 , n32334 , n32335 , n32336 , n32337 , n32338 , n32339 , n32340 , n32341 , n32342 , n32343 , n32344 , n32345 , n32346 , n32347 , n32348 , n32349 , n32350 , n32351 , n32352 , n32353 , n32354 , n32355 , n32356 , n32357 , n32358 , n32359 , n32360 , n32361 , n32362 , n32363 , n32364 , n32365 , n32366 , n32367 , n32368 , n32369 , n32370 , n32371 , n32372 , n32373 , n32374 , n32375 , n32376 , n32377 , n32378 , n32379 , n32380 , n32381 , n32382 , n32383 , n32384 , n32385 , n32386 , n32387 , n32388 , n32389 , n32390 , n32391 , n32392 , n32393 , n32394 , n32395 , n32396 , n32397 , n32398 , n32399 , n32400 , n32401 , n32402 , n32403 , n32404 , n32405 , n32406 , n32407 , n32408 , n32409 , n32410 , n32411 , n32412 , n32413 , n32414 , n32415 , n32416 , n32417 , n32418 , n32419 , n32420 , n32421 , n32422 , n32423 , n32424 , n32425 , n32426 , n32427 , n32428 , n32429 , n32430 , n32431 , n32432 , n32433 , n32434 , n32435 , n32436 , n32437 , n32438 , n32439 , n32440 , n32441 , n32442 , n32443 , n32444 , n32445 , n32446 , n32447 , n32448 , n32449 , n32450 , n32451 , n32452 , n32453 , n32454 , n32455 , n32456 , n32457 , n32458 , n32459 , n32460 , n32461 , n32462 , n32463 , n32464 , n32465 , n32466 , n32467 , n32468 , n32469 , n32470 , n32471 , n32472 , n32473 , n32474 , n32475 , n32476 , n32477 , n32478 , n32479 , n32480 , n32481 , n32482 , n32483 , n32484 , n32485 , n32486 , n32487 , n32488 , n32489 , n32490 , n32491 , n32492 , n32493 , n32494 , n32495 , n32496 , n32497 , n32498 , n32499 , n32500 , n32501 , n32502 , n32503 , n32504 , n32505 , n32506 , n32507 , n32508 , n32509 , n32510 , n32511 , n32512 , n32513 , n32514 , n32515 , n32516 , n32517 , n32518 , n32519 , n32520 , n32521 , n32522 , n32523 , n32524 , n32525 , n32526 , n32527 , n32528 , n32529 , n32530 , n32531 , n32532 , n32533 , n32534 , n32535 , n32536 , n32537 , n32538 , n32539 , n32540 , n32541 , n32542 , n32543 , n32544 , n32545 , n32546 , n32547 , n32548 , n32549 , n32550 , n32551 , n32552 , n32553 , n32554 , n32555 , n32556 , n32557 , n32558 , n32559 , n32560 , n32561 , n32562 , n32563 , n32564 , n32565 , n32566 , n32567 , n32568 , n32569 , n32570 , n32571 , n32572 , n32573 , n32574 , n32575 , n32576 , n32577 , n32578 , n32579 , n32580 , n32581 , n32582 , n32583 , n32584 , n32585 , n32586 , n32587 , n32588 , n32589 , n32590 , n32591 , n32592 , n32593 , n32594 , n32595 , n32596 , n32597 , n32598 , n32599 , n32600 , n32601 , n32602 , n32603 , n32604 , n32605 , n32606 , n32607 , n32608 , n32609 , n32610 , n32611 , n32612 , n32613 , n32614 , n32615 , n32616 , n32617 , n32618 , n32619 , n32620 , n32621 , n32622 , n32623 , n32624 , n32625 , n32626 , n32627 , n32628 , n32629 , n32630 , n32631 , n32632 , n32633 , n32634 , n32635 , n32636 , n32637 , n32638 , n32639 , n32640 , n32641 , n32642 , n32643 , n32644 , n32645 , n32646 , n32647 , n32648 , n32649 , n32650 , n32651 , n32652 , n32653 , n32654 , n32655 , n32656 , n32657 , n32658 , n32659 , n32660 , n32661 , n32662 , n32663 , n32664 , n32665 , n32666 , n32667 , n32668 , n32669 , n32670 , n32671 , n32672 , n32673 , n32674 , n32675 , n32676 , n32677 , n32678 , n32679 , n32680 , n32681 , n32682 , n32683 , n32684 , n32685 , n32686 , n32687 , n32688 , n32689 , n32690 , n32691 , n32692 , n32693 , n32694 , n32695 , n32696 , n32697 , n32698 , n32699 , n32700 , n32701 , n32702 , n32703 , n32704 , n32705 , n32706 , n32707 , n32708 , n32709 , n32710 , n32711 , n32712 , n32713 , n32714 , n32715 , n32716 , n32717 , n32718 , n32719 , n32720 , n32721 , n32722 , n32723 , n32724 , n32725 , n32726 , n32727 , n32728 , n32729 , n32730 , n32731 , n32732 , n32733 , n32734 , n32735 , n32736 , n32737 , n32738 , n32739 , n32740 , n32741 , n32742 , n32743 , n32744 , n32745 , n32746 , n32747 , n32748 , n32749 , n32750 , n32751 , n32752 , n32753 , n32754 , n32755 , n32756 , n32757 , n32758 , n32759 , n32760 , n32761 , n32762 , n32763 , n32764 , n32765 , n32766 , n32767 , n32768 , n32769 , n32770 , n32771 , n32772 , n32773 , n32774 , n32775 , n32776 , n32777 , n32778 , n32779 , n32780 , n32781 , n32782 , n32783 , n32784 , n32785 , n32786 , n32787 , n32788 , n32789 , n32790 , n32791 , n32792 , n32793 , n32794 , n32795 , n32796 , n32797 , n32798 , n32799 , n32800 , n32801 , n32802 , n32803 , n32804 , n32805 , n32806 , n32807 , n32808 , n32809 , n32810 , n32811 , n32812 , n32813 , n32814 , n32815 , n32816 , n32817 , n32818 , n32819 , n32820 , n32821 , n32822 , n32823 , n32824 , n32825 , n32826 , n32827 , n32828 , n32829 , n32830 , n32831 , n32832 , n32833 , n32834 , n32835 , n32836 , n32837 , n32838 , n32839 , n32840 , n32841 , n32842 , n32843 , n32844 , n32845 , n32846 , n32847 , n32848 , n32849 , n32850 , n32851 , n32852 , n32853 , n32854 , n32855 , n32856 , n32857 , n32858 , n32859 , n32860 , n32861 , n32862 , n32863 , n32864 , n32865 , n32866 , n32867 , n32868 , n32869 , n32870 , n32871 , n32872 , n32873 , n32874 , n32875 , n32876 , n32877 , n32878 , n32879 , n32880 , n32881 , n32882 , n32883 , n32884 , n32885 , n32886 , n32887 , n32888 , n32889 , n32890 , n32891 , n32892 , n32893 , n32894 , n32895 , n32896 , n32897 , n32898 , n32899 , n32900 , n32901 , n32902 , n32903 , n32904 , n32905 , n32906 , n32907 , n32908 , n32909 , n32910 , n32911 , n32912 , n32913 , n32914 , n32915 , n32916 , n32917 , n32918 , n32919 , n32920 , n32921 , n32922 , n32923 , n32924 , n32925 , n32926 , n32927 , n32928 , n32929 , n32930 , n32931 , n32932 , n32933 , n32934 , n32935 , n32936 , n32937 , n32938 , n32939 , n32940 , n32941 , n32942 , n32943 , n32944 , n32945 , n32946 , n32947 , n32948 , n32949 , n32950 , n32951 , n32952 , n32953 , n32954 , n32955 , n32956 , n32957 , n32958 , n32959 , n32960 , n32961 , n32962 , n32963 , n32964 , n32965 , n32966 , n32967 , n32968 , n32969 , n32970 , n32971 , n32972 , n32973 , n32974 , n32975 , n32976 , n32977 , n32978 , n32979 , n32980 , n32981 , n32982 , n32983 , n32984 , n32985 , n32986 , n32987 , n32988 , n32989 , n32990 , n32991 , n32992 , n32993 , n32994 , n32995 , n32996 , n32997 , n32998 , n32999 , n33000 , n33001 , n33002 , n33003 , n33004 , n33005 , n33006 , n33007 , n33008 , n33009 , n33010 , n33011 , n33012 , n33013 , n33014 , n33015 , n33016 , n33017 , n33018 , n33019 , n33020 , n33021 , n33022 , n33023 , n33024 , n33025 , n33026 , n33027 , n33028 , n33029 , n33030 , n33031 , n33032 , n33033 , n33034 , n33035 , n33036 , n33037 , n33038 , n33039 , n33040 , n33041 , n33042 , n33043 , n33044 , n33045 , n33046 , n33047 , n33048 , n33049 , n33050 , n33051 , n33052 , n33053 , n33054 , n33055 , n33056 , n33057 , n33058 , n33059 , n33060 , n33061 , n33062 , n33063 , n33064 , n33065 , n33066 , n33067 , n33068 , n33069 , n33070 , n33071 , n33072 , n33073 , n33074 , n33075 , n33076 , n33077 , n33078 , n33079 , n33080 , n33081 , n33082 , n33083 , n33084 , n33085 , n33086 , n33087 , n33088 , n33089 , n33090 , n33091 , n33092 , n33093 , n33094 , n33095 , n33096 , n33097 , n33098 , n33099 , n33100 , n33101 , n33102 , n33103 , n33104 , n33105 , n33106 , n33107 , n33108 , n33109 , n33110 , n33111 , n33112 , n33113 , n33114 , n33115 , n33116 , n33117 , n33118 , n33119 , n33120 , n33121 , n33122 , n33123 , n33124 , n33125 , n33126 , n33127 , n33128 , n33129 , n33130 , n33131 , n33132 , n33133 , n33134 , n33135 , n33136 , n33137 , n33138 , n33139 , n33140 , n33141 , n33142 , n33143 , n33144 , n33145 , n33146 , n33147 , n33148 , n33149 , n33150 , n33151 , n33152 , n33153 , n33154 , n33155 , n33156 , n33157 , n33158 , n33159 , n33160 , n33161 , n33162 , n33163 , n33164 , n33165 , n33166 , n33167 , n33168 , n33169 , n33170 , n33171 , n33172 , n33173 , n33174 , n33175 , n33176 , n33177 , n33178 , n33179 , n33180 , n33181 , n33182 , n33183 , n33184 , n33185 , n33186 , n33187 , n33188 , n33189 , n33190 , n33191 , n33192 , n33193 , n33194 , n33195 , n33196 , n33197 , n33198 , n33199 , n33200 , n33201 , n33202 , n33203 , n33204 , n33205 , n33206 , n33207 , n33208 , n33209 , n33210 , n33211 , n33212 , n33213 , n33214 , n33215 , n33216 , n33217 , n33218 , n33219 , n33220 , n33221 , n33222 , n33223 , n33224 , n33225 , n33226 , n33227 , n33228 , n33229 , n33230 , n33231 , n33232 , n33233 , n33234 , n33235 , n33236 , n33237 , n33238 , n33239 , n33240 , n33241 , n33242 , n33243 , n33244 , n33245 , n33246 , n33247 , n33248 , n33249 , n33250 , n33251 , n33252 , n33253 , n33254 , n33255 , n33256 , n33257 , n33258 , n33259 , n33260 , n33261 , n33262 , n33263 , n33264 , n33265 , n33266 , n33267 , n33268 , n33269 , n33270 , n33271 , n33272 , n33273 , n33274 , n33275 , n33276 , n33277 , n33278 , n33279 , n33280 , n33281 , n33282 , n33283 , n33284 , n33285 , n33286 , n33287 , n33288 , n33289 , n33290 , n33291 , n33292 , n33293 , n33294 , n33295 , n33296 , n33297 , n33298 , n33299 , n33300 , n33301 , n33302 , n33303 , n33304 , n33305 , n33306 , n33307 , n33308 , n33309 , n33310 , n33311 , n33312 , n33313 , n33314 , n33315 , n33316 , n33317 , n33318 , n33319 , n33320 , n33321 , n33322 , n33323 , n33324 , n33325 , n33326 , n33327 , n33328 , n33329 , n33330 , n33331 , n33332 , n33333 , n33334 , n33335 , n33336 , n33337 , n33338 , n33339 , n33340 , n33341 , n33342 , n33343 , n33344 , n33345 , n33346 , n33347 , n33348 , n33349 , n33350 , n33351 , n33352 , n33353 , n33354 , n33355 , n33356 , n33357 , n33358 , n33359 , n33360 , n33361 , n33362 , n33363 , n33364 , n33365 , n33366 , n33367 , n33368 , n33369 , n33370 , n33371 , n33372 , n33373 , n33374 , n33375 , n33376 , n33377 , n33378 , n33379 , n33380 , n33381 , n33382 , n33383 , n33384 , n33385 , n33386 , n33387 , n33388 , n33389 , n33390 , n33391 , n33392 , n33393 , n33394 , n33395 , n33396 , n33397 , n33398 , n33399 , n33400 , n33401 , n33402 , n33403 , n33404 , n33405 , n33406 , n33407 , n33408 , n33409 , n33410 , n33411 , n33412 , n33413 , n33414 , n33415 , n33416 , n33417 , n33418 , n33419 , n33420 , n33421 , n33422 , n33423 , n33424 , n33425 , n33426 , n33427 , n33428 , n33429 , n33430 , n33431 , n33432 , n33433 , n33434 , n33435 , n33436 , n33437 , n33438 , n33439 , n33440 , n33441 , n33442 , n33443 , n33444 , n33445 , n33446 , n33447 , n33448 , n33449 , n33450 , n33451 , n33452 , n33453 , n33454 , n33455 , n33456 , n33457 , n33458 , n33459 , n33460 , n33461 , n33462 , n33463 , n33464 , n33465 , n33466 , n33467 , n33468 , n33469 , n33470 , n33471 , n33472 , n33473 , n33474 , n33475 , n33476 , n33477 , n33478 , n33479 , n33480 , n33481 , n33482 , n33483 , n33484 , n33485 , n33486 , n33487 , n33488 , n33489 , n33490 , n33491 , n33492 , n33493 , n33494 , n33495 , n33496 , n33497 , n33498 , n33499 , n33500 , n33501 , n33502 , n33503 , n33504 , n33505 , n33506 , n33507 , n33508 , n33509 , n33510 , n33511 , n33512 , n33513 , n33514 , n33515 , n33516 , n33517 , n33518 , n33519 , n33520 , n33521 , n33522 , n33523 , n33524 , n33525 , n33526 , n33527 , n33528 , n33529 , n33530 , n33531 , n33532 , n33533 , n33534 , n33535 , n33536 , n33537 , n33538 , n33539 , n33540 , n33541 , n33542 , n33543 , n33544 , n33545 , n33546 , n33547 , n33548 , n33549 , n33550 , n33551 , n33552 , n33553 , n33554 , n33555 , n33556 , n33557 , n33558 , n33559 , n33560 , n33561 , n33562 , n33563 , n33564 , n33565 , n33566 , n33567 , n33568 , n33569 , n33570 , n33571 , n33572 , n33573 , n33574 , n33575 , n33576 , n33577 , n33578 , n33579 , n33580 , n33581 , n33582 , n33583 , n33584 , n33585 , n33586 , n33587 , n33588 , n33589 , n33590 , n33591 , n33592 , n33593 , n33594 , n33595 , n33596 , n33597 , n33598 , n33599 , n33600 , n33601 , n33602 , n33603 , n33604 , n33605 , n33606 , n33607 , n33608 , n33609 , n33610 , n33611 , n33612 , n33613 , n33614 , n33615 , n33616 , n33617 , n33618 , n33619 , n33620 , n33621 , n33622 , n33623 , n33624 , n33625 , n33626 , n33627 , n33628 , n33629 , n33630 , n33631 , n33632 , n33633 , n33634 , n33635 , n33636 , n33637 , n33638 , n33639 , n33640 , n33641 , n33642 , n33643 , n33644 , n33645 , n33646 , n33647 , n33648 , n33649 , n33650 , n33651 , n33652 , n33653 , n33654 , n33655 , n33656 , n33657 , n33658 , n33659 , n33660 , n33661 , n33662 , n33663 , n33664 , n33665 , n33666 , n33667 , n33668 , n33669 , n33670 , n33671 , n33672 , n33673 , n33674 , n33675 , n33676 , n33677 , n33678 , n33679 , n33680 , n33681 , n33682 , n33683 , n33684 , n33685 , n33686 , n33687 , n33688 , n33689 , n33690 , n33691 , n33692 , n33693 , n33694 , n33695 , n33696 , n33697 , n33698 , n33699 , n33700 , n33701 , n33702 , n33703 , n33704 , n33705 , n33706 , n33707 , n33708 , n33709 , n33710 , n33711 , n33712 , n33713 , n33714 , n33715 , n33716 , n33717 , n33718 , n33719 , n33720 , n33721 , n33722 , n33723 , n33724 , n33725 , n33726 , n33727 , n33728 , n33729 , n33730 , n33731 , n33732 , n33733 , n33734 , n33735 , n33736 , n33737 , n33738 , n33739 , n33740 , n33741 , n33742 , n33743 , n33744 , n33745 , n33746 , n33747 , n33748 , n33749 , n33750 , n33751 , n33752 , n33753 , n33754 , n33755 , n33756 , n33757 , n33758 , n33759 , n33760 , n33761 , n33762 , n33763 , n33764 , n33765 , n33766 , n33767 , n33768 , n33769 , n33770 , n33771 , n33772 , n33773 , n33774 , n33775 , n33776 , n33777 , n33778 , n33779 , n33780 , n33781 , n33782 , n33783 , n33784 , n33785 , n33786 , n33787 , n33788 , n33789 , n33790 , n33791 , n33792 , n33793 , n33794 , n33795 , n33796 , n33797 , n33798 , n33799 , n33800 , n33801 , n33802 , n33803 , n33804 , n33805 , n33806 , n33807 , n33808 , n33809 , n33810 , n33811 , n33812 , n33813 , n33814 , n33815 , n33816 , n33817 , n33818 , n33819 , n33820 , n33821 , n33822 , n33823 , n33824 , n33825 , n33826 , n33827 , n33828 , n33829 , n33830 , n33831 , n33832 , n33833 , n33834 , n33835 , n33836 , n33837 , n33838 , n33839 , n33840 , n33841 , n33842 , n33843 , n33844 , n33845 , n33846 , n33847 , n33848 , n33849 , n33850 , n33851 , n33852 , n33853 , n33854 , n33855 , n33856 , n33857 , n33858 , n33859 , n33860 , n33861 , n33862 , n33863 , n33864 , n33865 , n33866 , n33867 , n33868 , n33869 , n33870 , n33871 , n33872 , n33873 , n33874 , n33875 , n33876 , n33877 , n33878 , n33879 , n33880 , n33881 , n33882 , n33883 , n33884 , n33885 , n33886 , n33887 , n33888 , n33889 , n33890 , n33891 , n33892 , n33893 , n33894 , n33895 , n33896 , n33897 , n33898 , n33899 , n33900 , n33901 , n33902 , n33903 , n33904 , n33905 , n33906 , n33907 , n33908 , n33909 , n33910 , n33911 , n33912 , n33913 , n33914 , n33915 , n33916 , n33917 , n33918 , n33919 , n33920 , n33921 , n33922 , n33923 , n33924 , n33925 , n33926 , n33927 , n33928 , n33929 , n33930 , n33931 , n33932 , n33933 , n33934 , n33935 , n33936 , n33937 , n33938 , n33939 , n33940 , n33941 , n33942 , n33943 , n33944 , n33945 , n33946 , n33947 , n33948 , n33949 , n33950 , n33951 , n33952 , n33953 , n33954 , n33955 , n33956 , n33957 , n33958 , n33959 , n33960 , n33961 , n33962 , n33963 , n33964 , n33965 , n33966 , n33967 , n33968 , n33969 , n33970 , n33971 , n33972 , n33973 , n33974 , n33975 , n33976 , n33977 , n33978 , n33979 , n33980 , n33981 , n33982 , n33983 , n33984 , n33985 , n33986 , n33987 , n33988 , n33989 , n33990 , n33991 , n33992 , n33993 , n33994 , n33995 , n33996 , n33997 , n33998 , n33999 , n34000 , n34001 , n34002 , n34003 , n34004 , n34005 , n34006 , n34007 , n34008 , n34009 , n34010 , n34011 , n34012 , n34013 , n34014 , n34015 , n34016 , n34017 , n34018 , n34019 , n34020 , n34021 , n34022 , n34023 , n34024 , n34025 , n34026 , n34027 , n34028 , n34029 , n34030 , n34031 , n34032 , n34033 , n34034 , n34035 , n34036 , n34037 , n34038 , n34039 , n34040 , n34041 , n34042 , n34043 , n34044 , n34045 , n34046 , n34047 , n34048 , n34049 , n34050 , n34051 , n34052 , n34053 , n34054 , n34055 , n34056 , n34057 , n34058 , n34059 , n34060 , n34061 , n34062 , n34063 , n34064 , n34065 , n34066 , n34067 , n34068 , n34069 , n34070 , n34071 , n34072 , n34073 , n34074 , n34075 , n34076 , n34077 , n34078 , n34079 , n34080 , n34081 , n34082 , n34083 , n34084 , n34085 , n34086 , n34087 , n34088 , n34089 , n34090 , n34091 , n34092 , n34093 , n34094 , n34095 , n34096 , n34097 , n34098 , n34099 , n34100 , n34101 , n34102 , n34103 , n34104 , n34105 , n34106 , n34107 , n34108 , n34109 , n34110 , n34111 , n34112 , n34113 , n34114 , n34115 , n34116 , n34117 , n34118 , n34119 , n34120 , n34121 , n34122 , n34123 , n34124 , n34125 , n34126 , n34127 , n34128 , n34129 , n34130 , n34131 , n34132 , n34133 , n34134 , n34135 , n34136 , n34137 , n34138 , n34139 , n34140 , n34141 , n34142 , n34143 , n34144 , n34145 , n34146 , n34147 , n34148 , n34149 , n34150 , n34151 , n34152 , n34153 , n34154 , n34155 , n34156 , n34157 , n34158 , n34159 , n34160 , n34161 , n34162 , n34163 , n34164 , n34165 , n34166 , n34167 , n34168 , n34169 , n34170 , n34171 , n34172 , n34173 , n34174 , n34175 , n34176 , n34177 , n34178 , n34179 , n34180 , n34181 , n34182 , n34183 , n34184 , n34185 , n34186 , n34187 , n34188 , n34189 , n34190 , n34191 , n34192 , n34193 , n34194 , n34195 , n34196 , n34197 , n34198 , n34199 , n34200 , n34201 , n34202 , n34203 , n34204 , n34205 , n34206 , n34207 , n34208 , n34209 , n34210 , n34211 , n34212 , n34213 , n34214 , n34215 , n34216 , n34217 , n34218 , n34219 , n34220 , n34221 , n34222 , n34223 , n34224 , n34225 , n34226 , n34227 , n34228 , n34229 , n34230 , n34231 , n34232 , n34233 , n34234 , n34235 , n34236 , n34237 , n34238 , n34239 , n34240 , n34241 , n34242 , n34243 , n34244 , n34245 , n34246 , n34247 , n34248 , n34249 , n34250 , n34251 , n34252 , n34253 , n34254 , n34255 , n34256 , n34257 , n34258 , n34259 , n34260 , n34261 , n34262 , n34263 , n34264 , n34265 , n34266 , n34267 , n34268 , n34269 , n34270 , n34271 , n34272 , n34273 , n34274 , n34275 , n34276 , n34277 , n34278 , n34279 , n34280 , n34281 , n34282 , n34283 , n34284 , n34285 , n34286 , n34287 , n34288 , n34289 , n34290 , n34291 , n34292 , n34293 , n34294 , n34295 , n34296 , n34297 , n34298 , n34299 , n34300 , n34301 , n34302 , n34303 , n34304 , n34305 , n34306 , n34307 , n34308 , n34309 , n34310 , n34311 , n34312 , n34313 , n34314 , n34315 , n34316 , n34317 , n34318 , n34319 , n34320 , n34321 , n34322 , n34323 , n34324 , n34325 , n34326 , n34327 , n34328 , n34329 , n34330 , n34331 , n34332 , n34333 , n34334 , n34335 , n34336 , n34337 , n34338 , n34339 , n34340 , n34341 , n34342 , n34343 , n34344 , n34345 , n34346 , n34347 , n34348 , n34349 , n34350 , n34351 , n34352 , n34353 , n34354 , n34355 , n34356 , n34357 , n34358 , n34359 , n34360 , n34361 , n34362 , n34363 , n34364 , n34365 , n34366 , n34367 , n34368 , n34369 , n34370 , n34371 , n34372 , n34373 , n34374 , n34375 , n34376 , n34377 , n34378 , n34379 , n34380 , n34381 , n34382 , n34383 , n34384 , n34385 , n34386 , n34387 , n34388 , n34389 , n34390 , n34391 , n34392 , n34393 , n34394 , n34395 , n34396 , n34397 , n34398 , n34399 , n34400 , n34401 , n34402 , n34403 , n34404 , n34405 , n34406 , n34407 , n34408 , n34409 , n34410 , n34411 , n34412 , n34413 , n34414 , n34415 , n34416 , n34417 , n34418 , n34419 , n34420 , n34421 , n34422 , n34423 , n34424 , n34425 , n34426 , n34427 , n34428 , n34429 , n34430 , n34431 , n34432 , n34433 , n34434 , n34435 , n34436 , n34437 , n34438 , n34439 , n34440 , n34441 , n34442 , n34443 , n34444 , n34445 , n34446 , n34447 , n34448 , n34449 , n34450 , n34451 , n34452 , n34453 , n34454 , n34455 , n34456 , n34457 , n34458 , n34459 , n34460 , n34461 , n34462 , n34463 , n34464 , n34465 , n34466 , n34467 , n34468 , n34469 , n34470 , n34471 , n34472 , n34473 , n34474 , n34475 , n34476 , n34477 , n34478 , n34479 , n34480 , n34481 , n34482 , n34483 , n34484 , n34485 , n34486 , n34487 , n34488 , n34489 , n34490 , n34491 , n34492 , n34493 , n34494 , n34495 , n34496 , n34497 , n34498 , n34499 , n34500 , n34501 , n34502 , n34503 , n34504 , n34505 , n34506 , n34507 , n34508 , n34509 , n34510 , n34511 , n34512 , n34513 , n34514 , n34515 , n34516 , n34517 , n34518 , n34519 , n34520 , n34521 , n34522 , n34523 , n34524 , n34525 , n34526 , n34527 , n34528 , n34529 , n34530 , n34531 , n34532 , n34533 , n34534 , n34535 , n34536 , n34537 , n34538 , n34539 , n34540 , n34541 , n34542 , n34543 , n34544 , n34545 , n34546 , n34547 , n34548 , n34549 , n34550 , n34551 , n34552 , n34553 , n34554 , n34555 , n34556 , n34557 , n34558 , n34559 , n34560 , n34561 , n34562 , n34563 , n34564 , n34565 , n34566 , n34567 , n34568 , n34569 , n34570 , n34571 , n34572 , n34573 , n34574 , n34575 , n34576 , n34577 , n34578 , n34579 , n34580 , n34581 , n34582 , n34583 , n34584 , n34585 , n34586 , n34587 , n34588 , n34589 , n34590 , n34591 , n34592 , n34593 , n34594 , n34595 , n34596 , n34597 , n34598 , n34599 , n34600 , n34601 , n34602 , n34603 , n34604 , n34605 , n34606 , n34607 , n34608 , n34609 , n34610 , n34611 , n34612 , n34613 , n34614 , n34615 , n34616 , n34617 , n34618 , n34619 , n34620 , n34621 , n34622 , n34623 , n34624 , n34625 , n34626 , n34627 , n34628 , n34629 , n34630 , n34631 , n34632 , n34633 , n34634 , n34635 , n34636 , n34637 , n34638 , n34639 , n34640 , n34641 , n34642 , n34643 , n34644 , n34645 , n34646 , n34647 , n34648 , n34649 , n34650 , n34651 , n34652 , n34653 , n34654 , n34655 , n34656 , n34657 , n34658 , n34659 , n34660 , n34661 , n34662 , n34663 , n34664 , n34665 , n34666 , n34667 , n34668 , n34669 , n34670 , n34671 , n34672 , n34673 , n34674 , n34675 , n34676 , n34677 , n34678 , n34679 , n34680 , n34681 , n34682 , n34683 , n34684 , n34685 , n34686 , n34687 , n34688 , n34689 , n34690 , n34691 , n34692 , n34693 , n34694 , n34695 , n34696 , n34697 , n34698 , n34699 , n34700 , n34701 , n34702 , n34703 , n34704 , n34705 , n34706 , n34707 , n34708 , n34709 , n34710 , n34711 , n34712 , n34713 , n34714 , n34715 , n34716 , n34717 , n34718 , n34719 , n34720 , n34721 , n34722 , n34723 , n34724 , n34725 , n34726 , n34727 , n34728 , n34729 , n34730 , n34731 , n34732 , n34733 , n34734 , n34735 , n34736 , n34737 , n34738 , n34739 , n34740 , n34741 , n34742 , n34743 , n34744 , n34745 , n34746 , n34747 , n34748 , n34749 , n34750 , n34751 , n34752 , n34753 , n34754 , n34755 , n34756 , n34757 , n34758 , n34759 , n34760 , n34761 , n34762 , n34763 , n34764 , n34765 , n34766 , n34767 , n34768 , n34769 , n34770 , n34771 , n34772 , n34773 , n34774 , n34775 , n34776 , n34777 , n34778 , n34779 , n34780 , n34781 , n34782 , n34783 , n34784 , n34785 , n34786 , n34787 , n34788 , n34789 , n34790 , n34791 , n34792 , n34793 , n34794 , n34795 , n34796 , n34797 , n34798 , n34799 , n34800 , n34801 , n34802 , n34803 , n34804 , n34805 , n34806 , n34807 , n34808 , n34809 , n34810 , n34811 , n34812 , n34813 , n34814 , n34815 , n34816 , n34817 , n34818 , n34819 , n34820 , n34821 , n34822 , n34823 , n34824 , n34825 , n34826 , n34827 , n34828 , n34829 , n34830 , n34831 , n34832 , n34833 , n34834 , n34835 , n34836 , n34837 , n34838 , n34839 , n34840 , n34841 , n34842 , n34843 , n34844 , n34845 , n34846 , n34847 , n34848 , n34849 , n34850 , n34851 , n34852 , n34853 , n34854 , n34855 , n34856 , n34857 , n34858 , n34859 , n34860 , n34861 , n34862 , n34863 , n34864 , n34865 , n34866 , n34867 , n34868 , n34869 , n34870 , n34871 , n34872 , n34873 , n34874 , n34875 , n34876 , n34877 , n34878 , n34879 , n34880 , n34881 , n34882 , n34883 , n34884 , n34885 , n34886 , n34887 , n34888 , n34889 , n34890 , n34891 , n34892 , n34893 , n34894 , n34895 , n34896 , n34897 , n34898 , n34899 , n34900 , n34901 , n34902 , n34903 , n34904 , n34905 , n34906 , n34907 , n34908 , n34909 , n34910 , n34911 , n34912 , n34913 , n34914 , n34915 , n34916 , n34917 , n34918 , n34919 , n34920 , n34921 , n34922 , n34923 , n34924 , n34925 , n34926 , n34927 , n34928 , n34929 , n34930 , n34931 , n34932 , n34933 , n34934 , n34935 , n34936 , n34937 , n34938 , n34939 , n34940 , n34941 , n34942 , n34943 , n34944 , n34945 , n34946 , n34947 , n34948 , n34949 , n34950 , n34951 , n34952 , n34953 , n34954 , n34955 , n34956 , n34957 , n34958 , n34959 , n34960 , n34961 , n34962 , n34963 , n34964 , n34965 , n34966 , n34967 , n34968 , n34969 , n34970 , n34971 , n34972 , n34973 , n34974 , n34975 , n34976 , n34977 , n34978 , n34979 , n34980 , n34981 , n34982 , n34983 , n34984 , n34985 , n34986 , n34987 , n34988 , n34989 , n34990 , n34991 , n34992 , n34993 , n34994 , n34995 , n34996 , n34997 , n34998 , n34999 , n35000 , n35001 , n35002 , n35003 , n35004 , n35005 , n35006 , n35007 , n35008 , n35009 , n35010 , n35011 , n35012 , n35013 , n35014 , n35015 , n35016 , n35017 , n35018 , n35019 , n35020 , n35021 , n35022 , n35023 , n35024 , n35025 , n35026 , n35027 , n35028 , n35029 , n35030 , n35031 , n35032 , n35033 , n35034 , n35035 , n35036 , n35037 , n35038 , n35039 , n35040 , n35041 , n35042 , n35043 , n35044 , n35045 , n35046 , n35047 , n35048 , n35049 , n35050 , n35051 , n35052 , n35053 , n35054 , n35055 , n35056 , n35057 , n35058 , n35059 , n35060 , n35061 , n35062 , n35063 , n35064 , n35065 , n35066 , n35067 , n35068 , n35069 , n35070 , n35071 , n35072 , n35073 , n35074 , n35075 , n35076 , n35077 , n35078 , n35079 , n35080 , n35081 , n35082 , n35083 , n35084 , n35085 , n35086 , n35087 , n35088 , n35089 , n35090 , n35091 , n35092 , n35093 , n35094 , n35095 , n35096 , n35097 , n35098 , n35099 , n35100 , n35101 , n35102 , n35103 , n35104 , n35105 , n35106 , n35107 , n35108 , n35109 , n35110 , n35111 , n35112 , n35113 , n35114 , n35115 , n35116 , n35117 , n35118 , n35119 , n35120 , n35121 , n35122 , n35123 , n35124 , n35125 , n35126 , n35127 , n35128 , n35129 , n35130 , n35131 , n35132 , n35133 , n35134 , n35135 , n35136 , n35137 , n35138 , n35139 , n35140 , n35141 , n35142 , n35143 , n35144 , n35145 , n35146 , n35147 , n35148 , n35149 , n35150 , n35151 , n35152 , n35153 , n35154 , n35155 , n35156 , n35157 , n35158 , n35159 , n35160 , n35161 , n35162 , n35163 , n35164 , n35165 , n35166 , n35167 , n35168 , n35169 , n35170 , n35171 , n35172 , n35173 , n35174 , n35175 , n35176 , n35177 , n35178 , n35179 , n35180 , n35181 , n35182 , n35183 , n35184 , n35185 , n35186 , n35187 , n35188 , n35189 , n35190 , n35191 , n35192 , n35193 , n35194 , n35195 , n35196 , n35197 , n35198 , n35199 , n35200 , n35201 , n35202 , n35203 , n35204 , n35205 , n35206 , n35207 , n35208 , n35209 , n35210 , n35211 , n35212 , n35213 , n35214 , n35215 , n35216 , n35217 , n35218 , n35219 , n35220 , n35221 , n35222 , n35223 , n35224 , n35225 , n35226 , n35227 , n35228 , n35229 , n35230 , n35231 , n35232 , n35233 , n35234 , n35235 , n35236 , n35237 , n35238 , n35239 , n35240 , n35241 , n35242 , n35243 , n35244 , n35245 , n35246 , n35247 , n35248 , n35249 , n35250 , n35251 , n35252 , n35253 , n35254 , n35255 , n35256 , n35257 , n35258 , n35259 , n35260 , n35261 , n35262 , n35263 , n35264 , n35265 , n35266 , n35267 , n35268 , n35269 , n35270 , n35271 , n35272 , n35273 , n35274 , n35275 , n35276 , n35277 , n35278 , n35279 , n35280 , n35281 , n35282 , n35283 , n35284 , n35285 , n35286 , n35287 , n35288 , n35289 , n35290 , n35291 , n35292 , n35293 , n35294 , n35295 , n35296 , n35297 , n35298 , n35299 , n35300 , n35301 , n35302 , n35303 , n35304 , n35305 , n35306 , n35307 , n35308 , n35309 , n35310 , n35311 , n35312 , n35313 , n35314 , n35315 , n35316 , n35317 , n35318 , n35319 , n35320 , n35321 , n35322 , n35323 , n35324 , n35325 , n35326 , n35327 , n35328 , n35329 , n35330 , n35331 , n35332 , n35333 , n35334 , n35335 , n35336 , n35337 , n35338 , n35339 , n35340 , n35341 , n35342 , n35343 , n35344 , n35345 , n35346 , n35347 , n35348 , n35349 , n35350 , n35351 , n35352 , n35353 , n35354 , n35355 , n35356 , n35357 , n35358 , n35359 , n35360 , n35361 , n35362 , n35363 , n35364 , n35365 , n35366 , n35367 , n35368 , n35369 , n35370 , n35371 , n35372 , n35373 , n35374 , n35375 , n35376 , n35377 , n35378 , n35379 , n35380 , n35381 , n35382 , n35383 , n35384 , n35385 , n35386 , n35387 , n35388 , n35389 , n35390 , n35391 , n35392 , n35393 , n35394 , n35395 , n35396 , n35397 , n35398 , n35399 , n35400 , n35401 , n35402 , n35403 , n35404 , n35405 , n35406 , n35407 , n35408 , n35409 , n35410 , n35411 , n35412 , n35413 , n35414 , n35415 , n35416 , n35417 , n35418 , n35419 , n35420 , n35421 , n35422 , n35423 , n35424 , n35425 , n35426 , n35427 , n35428 , n35429 , n35430 , n35431 , n35432 , n35433 , n35434 , n35435 , n35436 , n35437 , n35438 , n35439 , n35440 , n35441 , n35442 , n35443 , n35444 , n35445 , n35446 , n35447 , n35448 , n35449 , n35450 , n35451 , n35452 , n35453 , n35454 , n35455 , n35456 , n35457 , n35458 , n35459 , n35460 , n35461 , n35462 , n35463 , n35464 , n35465 , n35466 , n35467 , n35468 , n35469 , n35470 , n35471 , n35472 , n35473 , n35474 , n35475 , n35476 , n35477 , n35478 , n35479 , n35480 , n35481 , n35482 , n35483 , n35484 , n35485 , n35486 , n35487 , n35488 , n35489 , n35490 , n35491 , n35492 , n35493 , n35494 , n35495 , n35496 , n35497 , n35498 , n35499 , n35500 , n35501 , n35502 , n35503 , n35504 , n35505 , n35506 , n35507 , n35508 , n35509 , n35510 , n35511 , n35512 , n35513 , n35514 , n35515 , n35516 , n35517 , n35518 , n35519 , n35520 , n35521 , n35522 , n35523 , n35524 , n35525 , n35526 , n35527 , n35528 , n35529 , n35530 , n35531 , n35532 , n35533 , n35534 , n35535 , n35536 , n35537 , n35538 , n35539 , n35540 , n35541 , n35542 , n35543 , n35544 , n35545 , n35546 , n35547 , n35548 , n35549 , n35550 , n35551 , n35552 , n35553 , n35554 , n35555 , n35556 , n35557 , n35558 , n35559 , n35560 , n35561 , n35562 , n35563 , n35564 , n35565 , n35566 , n35567 , n35568 , n35569 , n35570 , n35571 , n35572 , n35573 , n35574 , n35575 , n35576 , n35577 , n35578 , n35579 , n35580 , n35581 , n35582 , n35583 , n35584 , n35585 , n35586 , n35587 , n35588 , n35589 , n35590 , n35591 , n35592 , n35593 , n35594 , n35595 , n35596 , n35597 , n35598 , n35599 , n35600 , n35601 , n35602 , n35603 , n35604 , n35605 , n35606 , n35607 , n35608 , n35609 , n35610 , n35611 , n35612 , n35613 , n35614 , n35615 , n35616 , n35617 , n35618 , n35619 , n35620 , n35621 , n35622 , n35623 , n35624 , n35625 , n35626 , n35627 , n35628 , n35629 , n35630 , n35631 , n35632 , n35633 , n35634 , n35635 , n35636 , n35637 , n35638 , n35639 , n35640 , n35641 , n35642 , n35643 , n35644 , n35645 , n35646 , n35647 , n35648 , n35649 , n35650 , n35651 , n35652 , n35653 , n35654 , n35655 , n35656 , n35657 , n35658 , n35659 , n35660 , n35661 , n35662 , n35663 , n35664 , n35665 , n35666 , n35667 , n35668 , n35669 , n35670 , n35671 , n35672 , n35673 , n35674 , n35675 , n35676 , n35677 , n35678 , n35679 , n35680 , n35681 , n35682 , n35683 , n35684 , n35685 , n35686 , n35687 , n35688 , n35689 , n35690 , n35691 , n35692 , n35693 , n35694 , n35695 , n35696 , n35697 , n35698 , n35699 , n35700 , n35701 , n35702 , n35703 , n35704 , n35705 , n35706 , n35707 , n35708 , n35709 , n35710 , n35711 , n35712 , n35713 , n35714 , n35715 , n35716 , n35717 , n35718 , n35719 , n35720 , n35721 , n35722 , n35723 , n35724 , n35725 , n35726 , n35727 , n35728 , n35729 , n35730 , n35731 , n35732 , n35733 , n35734 , n35735 , n35736 , n35737 , n35738 , n35739 , n35740 , n35741 , n35742 , n35743 , n35744 , n35745 , n35746 , n35747 , n35748 , n35749 , n35750 , n35751 , n35752 , n35753 , n35754 , n35755 , n35756 , n35757 , n35758 , n35759 , n35760 , n35761 , n35762 , n35763 , n35764 , n35765 , n35766 , n35767 , n35768 , n35769 , n35770 , n35771 , n35772 , n35773 , n35774 , n35775 , n35776 , n35777 , n35778 , n35779 , n35780 , n35781 , n35782 , n35783 , n35784 , n35785 , n35786 , n35787 , n35788 , n35789 , n35790 , n35791 , n35792 , n35793 , n35794 , n35795 , n35796 , n35797 , n35798 , n35799 , n35800 , n35801 , n35802 , n35803 , n35804 , n35805 , n35806 , n35807 , n35808 , n35809 , n35810 , n35811 , n35812 , n35813 , n35814 , n35815 , n35816 , n35817 , n35818 , n35819 , n35820 , n35821 , n35822 , n35823 , n35824 , n35825 , n35826 , n35827 , n35828 , n35829 , n35830 , n35831 , n35832 , n35833 , n35834 , n35835 , n35836 , n35837 , n35838 , n35839 , n35840 , n35841 , n35842 , n35843 , n35844 , n35845 , n35846 , n35847 , n35848 , n35849 , n35850 , n35851 , n35852 , n35853 , n35854 , n35855 , n35856 , n35857 , n35858 , n35859 , n35860 , n35861 , n35862 , n35863 , n35864 , n35865 , n35866 , n35867 , n35868 , n35869 , n35870 , n35871 , n35872 , n35873 , n35874 , n35875 , n35876 , n35877 , n35878 , n35879 , n35880 , n35881 , n35882 , n35883 , n35884 , n35885 , n35886 , n35887 , n35888 , n35889 , n35890 , n35891 , n35892 , n35893 , n35894 , n35895 , n35896 , n35897 , n35898 , n35899 , n35900 , n35901 , n35902 , n35903 , n35904 , n35905 , n35906 , n35907 , n35908 , n35909 , n35910 , n35911 , n35912 , n35913 , n35914 , n35915 , n35916 , n35917 , n35918 , n35919 , n35920 , n35921 , n35922 , n35923 , n35924 , n35925 , n35926 , n35927 , n35928 , n35929 , n35930 , n35931 , n35932 , n35933 , n35934 , n35935 , n35936 , n35937 , n35938 , n35939 , n35940 , n35941 , n35942 , n35943 , n35944 , n35945 , n35946 , n35947 , n35948 , n35949 , n35950 , n35951 , n35952 , n35953 , n35954 , n35955 , n35956 , n35957 , n35958 , n35959 , n35960 , n35961 , n35962 , n35963 , n35964 , n35965 , n35966 , n35967 , n35968 , n35969 , n35970 , n35971 , n35972 , n35973 , n35974 , n35975 , n35976 , n35977 , n35978 , n35979 , n35980 , n35981 , n35982 , n35983 , n35984 , n35985 , n35986 , n35987 , n35988 , n35989 , n35990 , n35991 , n35992 , n35993 , n35994 , n35995 , n35996 , n35997 , n35998 , n35999 , n36000 , n36001 , n36002 , n36003 , n36004 , n36005 , n36006 , n36007 , n36008 , n36009 , n36010 , n36011 , n36012 , n36013 , n36014 , n36015 , n36016 , n36017 , n36018 , n36019 , n36020 , n36021 , n36022 , n36023 , n36024 , n36025 , n36026 , n36027 , n36028 , n36029 , n36030 , n36031 , n36032 , n36033 , n36034 , n36035 , n36036 , n36037 , n36038 , n36039 , n36040 , n36041 , n36042 , n36043 , n36044 , n36045 , n36046 , n36047 , n36048 , n36049 , n36050 , n36051 , n36052 , n36053 , n36054 , n36055 , n36056 , n36057 , n36058 , n36059 , n36060 , n36061 , n36062 , n36063 , n36064 , n36065 , n36066 , n36067 , n36068 , n36069 , n36070 , n36071 , n36072 , n36073 , n36074 , n36075 , n36076 , n36077 , n36078 , n36079 , n36080 , n36081 , n36082 , n36083 , n36084 , n36085 , n36086 , n36087 , n36088 , n36089 , n36090 , n36091 , n36092 , n36093 , n36094 , n36095 , n36096 , n36097 , n36098 , n36099 , n36100 , n36101 , n36102 , n36103 , n36104 , n36105 , n36106 , n36107 , n36108 , n36109 , n36110 , n36111 , n36112 , n36113 , n36114 , n36115 , n36116 , n36117 , n36118 , n36119 , n36120 , n36121 , n36122 , n36123 , n36124 , n36125 , n36126 , n36127 , n36128 , n36129 , n36130 , n36131 , n36132 , n36133 , n36134 , n36135 , n36136 , n36137 , n36138 , n36139 , n36140 , n36141 , n36142 , n36143 , n36144 , n36145 , n36146 , n36147 , n36148 , n36149 , n36150 , n36151 , n36152 , n36153 , n36154 , n36155 , n36156 , n36157 , n36158 , n36159 , n36160 , n36161 , n36162 , n36163 , n36164 , n36165 , n36166 , n36167 , n36168 , n36169 , n36170 , n36171 , n36172 , n36173 , n36174 , n36175 , n36176 , n36177 , n36178 , n36179 , n36180 , n36181 , n36182 , n36183 , n36184 , n36185 , n36186 , n36187 , n36188 , n36189 , n36190 , n36191 , n36192 , n36193 , n36194 , n36195 , n36196 , n36197 , n36198 , n36199 , n36200 , n36201 , n36202 , n36203 , n36204 , n36205 , n36206 , n36207 , n36208 , n36209 , n36210 , n36211 , n36212 , n36213 , n36214 , n36215 , n36216 , n36217 , n36218 , n36219 , n36220 , n36221 , n36222 , n36223 , n36224 , n36225 , n36226 , n36227 , n36228 , n36229 , n36230 , n36231 , n36232 , n36233 , n36234 , n36235 , n36236 , n36237 , n36238 , n36239 , n36240 , n36241 , n36242 , n36243 , n36244 , n36245 , n36246 , n36247 , n36248 , n36249 , n36250 , n36251 , n36252 , n36253 , n36254 , n36255 , n36256 , n36257 , n36258 , n36259 , n36260 , n36261 , n36262 , n36263 , n36264 , n36265 , n36266 , n36267 , n36268 , n36269 , n36270 , n36271 , n36272 , n36273 , n36274 , n36275 , n36276 , n36277 , n36278 , n36279 , n36280 , n36281 , n36282 , n36283 , n36284 , n36285 , n36286 , n36287 , n36288 , n36289 , n36290 , n36291 , n36292 , n36293 , n36294 , n36295 , n36296 , n36297 , n36298 , n36299 , n36300 , n36301 , n36302 , n36303 , n36304 , n36305 , n36306 , n36307 , n36308 , n36309 , n36310 , n36311 , n36312 , n36313 , n36314 , n36315 , n36316 , n36317 , n36318 , n36319 , n36320 , n36321 , n36322 , n36323 , n36324 , n36325 , n36326 , n36327 , n36328 , n36329 , n36330 , n36331 , n36332 , n36333 , n36334 , n36335 , n36336 , n36337 , n36338 , n36339 , n36340 , n36341 , n36342 , n36343 , n36344 , n36345 , n36346 , n36347 , n36348 , n36349 , n36350 , n36351 , n36352 , n36353 , n36354 , n36355 , n36356 , n36357 , n36358 , n36359 , n36360 , n36361 , n36362 , n36363 , n36364 , n36365 , n36366 , n36367 , n36368 , n36369 , n36370 , n36371 , n36372 , n36373 , n36374 , n36375 , n36376 , n36377 , n36378 , n36379 , n36380 , n36381 , n36382 , n36383 , n36384 , n36385 , n36386 , n36387 , n36388 , n36389 , n36390 , n36391 , n36392 , n36393 , n36394 , n36395 , n36396 , n36397 , n36398 , n36399 , n36400 , n36401 , n36402 , n36403 , n36404 , n36405 , n36406 , n36407 , n36408 , n36409 , n36410 , n36411 , n36412 , n36413 , n36414 , n36415 , n36416 , n36417 , n36418 , n36419 , n36420 , n36421 , n36422 , n36423 , n36424 , n36425 , n36426 , n36427 , n36428 , n36429 , n36430 , n36431 , n36432 , n36433 , n36434 , n36435 , n36436 , n36437 , n36438 , n36439 , n36440 , n36441 , n36442 , n36443 , n36444 , n36445 , n36446 , n36447 , n36448 , n36449 , n36450 , n36451 , n36452 , n36453 , n36454 , n36455 , n36456 , n36457 , n36458 , n36459 , n36460 , n36461 , n36462 , n36463 , n36464 , n36465 , n36466 , n36467 , n36468 , n36469 , n36470 , n36471 , n36472 , n36473 , n36474 , n36475 , n36476 , n36477 , n36478 , n36479 , n36480 , n36481 , n36482 , n36483 , n36484 , n36485 , n36486 , n36487 , n36488 , n36489 , n36490 , n36491 , n36492 , n36493 , n36494 , n36495 , n36496 , n36497 , n36498 , n36499 , n36500 , n36501 , n36502 , n36503 , n36504 , n36505 , n36506 , n36507 , n36508 , n36509 , n36510 , n36511 , n36512 , n36513 , n36514 , n36515 , n36516 , n36517 , n36518 , n36519 , n36520 , n36521 , n36522 , n36523 , n36524 , n36525 , n36526 , n36527 , n36528 , n36529 , n36530 , n36531 , n36532 , n36533 , n36534 , n36535 , n36536 , n36537 , n36538 , n36539 , n36540 , n36541 , n36542 , n36543 , n36544 , n36545 , n36546 , n36547 , n36548 , n36549 , n36550 , n36551 , n36552 , n36553 , n36554 , n36555 , n36556 , n36557 , n36558 , n36559 , n36560 , n36561 , n36562 , n36563 , n36564 , n36565 , n36566 , n36567 , n36568 , n36569 , n36570 , n36571 , n36572 , n36573 , n36574 , n36575 , n36576 , n36577 , n36578 , n36579 , n36580 , n36581 , n36582 , n36583 , n36584 , n36585 , n36586 , n36587 , n36588 , n36589 , n36590 , n36591 , n36592 , n36593 , n36594 , n36595 , n36596 , n36597 , n36598 , n36599 , n36600 , n36601 , n36602 , n36603 , n36604 , n36605 , n36606 , n36607 , n36608 , n36609 , n36610 , n36611 , n36612 , n36613 , n36614 , n36615 , n36616 , n36617 , n36618 , n36619 , n36620 , n36621 , n36622 , n36623 , n36624 , n36625 , n36626 , n36627 , n36628 , n36629 , n36630 , n36631 , n36632 , n36633 , n36634 , n36635 , n36636 , n36637 , n36638 , n36639 , n36640 , n36641 , n36642 , n36643 , n36644 , n36645 , n36646 , n36647 , n36648 , n36649 , n36650 , n36651 , n36652 , n36653 , n36654 , n36655 , n36656 , n36657 , n36658 , n36659 , n36660 , n36661 , n36662 , n36663 , n36664 , n36665 , n36666 , n36667 , n36668 , n36669 , n36670 , n36671 , n36672 , n36673 , n36674 , n36675 , n36676 , n36677 , n36678 , n36679 , n36680 , n36681 , n36682 , n36683 , n36684 , n36685 , n36686 , n36687 , n36688 , n36689 , n36690 , n36691 , n36692 , n36693 , n36694 , n36695 , n36696 , n36697 , n36698 , n36699 , n36700 , n36701 , n36702 , n36703 , n36704 , n36705 , n36706 , n36707 , n36708 , n36709 , n36710 , n36711 , n36712 , n36713 , n36714 , n36715 , n36716 , n36717 , n36718 , n36719 , n36720 , n36721 , n36722 , n36723 , n36724 , n36725 , n36726 , n36727 , n36728 , n36729 , n36730 , n36731 , n36732 , n36733 , n36734 , n36735 , n36736 , n36737 , n36738 , n36739 , n36740 , n36741 , n36742 , n36743 , n36744 , n36745 , n36746 , n36747 , n36748 , n36749 , n36750 , n36751 , n36752 , n36753 , n36754 , n36755 , n36756 , n36757 , n36758 , n36759 , n36760 , n36761 , n36762 , n36763 , n36764 , n36765 , n36766 , n36767 , n36768 , n36769 , n36770 , n36771 , n36772 , n36773 , n36774 , n36775 , n36776 , n36777 , n36778 , n36779 , n36780 , n36781 , n36782 , n36783 , n36784 , n36785 , n36786 , n36787 , n36788 , n36789 , n36790 , n36791 , n36792 , n36793 , n36794 , n36795 , n36796 , n36797 , n36798 , n36799 , n36800 , n36801 , n36802 , n36803 , n36804 , n36805 , n36806 , n36807 , n36808 , n36809 , n36810 , n36811 , n36812 , n36813 , n36814 , n36815 , n36816 , n36817 , n36818 , n36819 , n36820 , n36821 , n36822 , n36823 , n36824 , n36825 , n36826 , n36827 , n36828 , n36829 , n36830 , n36831 , n36832 , n36833 , n36834 , n36835 , n36836 , n36837 , n36838 , n36839 , n36840 , n36841 , n36842 , n36843 , n36844 , n36845 , n36846 , n36847 , n36848 , n36849 , n36850 , n36851 , n36852 , n36853 , n36854 , n36855 , n36856 , n36857 , n36858 , n36859 , n36860 , n36861 , n36862 , n36863 , n36864 , n36865 , n36866 , n36867 , n36868 , n36869 , n36870 , n36871 , n36872 , n36873 , n36874 , n36875 , n36876 , n36877 , n36878 , n36879 , n36880 , n36881 , n36882 , n36883 , n36884 , n36885 , n36886 , n36887 , n36888 , n36889 , n36890 , n36891 , n36892 , n36893 , n36894 , n36895 , n36896 , n36897 , n36898 , n36899 , n36900 , n36901 , n36902 , n36903 , n36904 , n36905 , n36906 , n36907 , n36908 , n36909 , n36910 , n36911 , n36912 , n36913 , n36914 , n36915 , n36916 , n36917 , n36918 , n36919 , n36920 , n36921 , n36922 , n36923 , n36924 , n36925 , n36926 , n36927 , n36928 , n36929 , n36930 , n36931 , n36932 , n36933 , n36934 , n36935 , n36936 , n36937 , n36938 , n36939 , n36940 , n36941 , n36942 , n36943 , n36944 , n36945 , n36946 , n36947 , n36948 , n36949 , n36950 , n36951 , n36952 , n36953 , n36954 , n36955 , n36956 , n36957 , n36958 , n36959 , n36960 , n36961 , n36962 , n36963 , n36964 , n36965 , n36966 , n36967 , n36968 , n36969 , n36970 , n36971 , n36972 , n36973 , n36974 , n36975 , n36976 , n36977 , n36978 , n36979 , n36980 , n36981 , n36982 , n36983 , n36984 , n36985 , n36986 , n36987 , n36988 , n36989 , n36990 , n36991 , n36992 , n36993 , n36994 , n36995 , n36996 , n36997 , n36998 , n36999 , n37000 , n37001 , n37002 , n37003 , n37004 , n37005 , n37006 , n37007 , n37008 , n37009 , n37010 , n37011 , n37012 , n37013 , n37014 , n37015 , n37016 , n37017 , n37018 , n37019 , n37020 , n37021 , n37022 , n37023 , n37024 , n37025 , n37026 , n37027 , n37028 , n37029 , n37030 , n37031 , n37032 , n37033 , n37034 , n37035 , n37036 , n37037 , n37038 , n37039 , n37040 , n37041 , n37042 , n37043 , n37044 , n37045 , n37046 , n37047 , n37048 , n37049 , n37050 , n37051 , n37052 , n37053 , n37054 , n37055 , n37056 , n37057 , n37058 , n37059 , n37060 , n37061 , n37062 , n37063 , n37064 , n37065 , n37066 , n37067 , n37068 , n37069 , n37070 , n37071 , n37072 , n37073 , n37074 , n37075 , n37076 , n37077 , n37078 , n37079 , n37080 , n37081 , n37082 , n37083 , n37084 , n37085 , n37086 , n37087 , n37088 , n37089 , n37090 , n37091 , n37092 , n37093 , n37094 , n37095 , n37096 , n37097 , n37098 , n37099 , n37100 , n37101 , n37102 , n37103 , n37104 , n37105 , n37106 , n37107 , n37108 , n37109 , n37110 , n37111 , n37112 , n37113 , n37114 , n37115 , n37116 , n37117 , n37118 , n37119 , n37120 , n37121 , n37122 , n37123 , n37124 , n37125 , n37126 , n37127 , n37128 , n37129 , n37130 , n37131 , n37132 , n37133 , n37134 , n37135 , n37136 , n37137 , n37138 , n37139 , n37140 , n37141 , n37142 , n37143 , n37144 , n37145 , n37146 , n37147 , n37148 , n37149 , n37150 , n37151 , n37152 , n37153 , n37154 , n37155 , n37156 , n37157 , n37158 , n37159 , n37160 , n37161 , n37162 , n37163 , n37164 , n37165 , n37166 , n37167 , n37168 , n37169 , n37170 , n37171 , n37172 , n37173 , n37174 , n37175 , n37176 , n37177 , n37178 , n37179 , n37180 , n37181 , n37182 , n37183 , n37184 , n37185 , n37186 , n37187 , n37188 , n37189 , n37190 , n37191 , n37192 , n37193 , n37194 , n37195 , n37196 , n37197 , n37198 , n37199 , n37200 , n37201 , n37202 , n37203 , n37204 , n37205 , n37206 , n37207 , n37208 , n37209 , n37210 , n37211 , n37212 , n37213 , n37214 , n37215 , n37216 , n37217 , n37218 , n37219 , n37220 , n37221 , n37222 , n37223 , n37224 , n37225 , n37226 , n37227 , n37228 , n37229 , n37230 , n37231 , n37232 , n37233 , n37234 , n37235 , n37236 , n37237 , n37238 , n37239 , n37240 , n37241 , n37242 , n37243 , n37244 , n37245 , n37246 , n37247 , n37248 , n37249 , n37250 , n37251 , n37252 , n37253 , n37254 , n37255 , n37256 , n37257 , n37258 , n37259 , n37260 , n37261 , n37262 , n37263 , n37264 , n37265 , n37266 , n37267 , n37268 , n37269 , n37270 , n37271 , n37272 , n37273 , n37274 , n37275 , n37276 , n37277 , n37278 , n37279 , n37280 , n37281 , n37282 , n37283 , n37284 , n37285 , n37286 , n37287 , n37288 , n37289 , n37290 , n37291 , n37292 , n37293 , n37294 , n37295 , n37296 , n37297 , n37298 , n37299 , n37300 , n37301 , n37302 , n37303 , n37304 , n37305 , n37306 , n37307 , n37308 , n37309 , n37310 , n37311 , n37312 , n37313 , n37314 , n37315 , n37316 , n37317 , n37318 , n37319 , n37320 , n37321 , n37322 , n37323 , n37324 , n37325 , n37326 , n37327 , n37328 , n37329 , n37330 , n37331 , n37332 , n37333 , n37334 , n37335 , n37336 , n37337 , n37338 , n37339 , n37340 , n37341 , n37342 , n37343 , n37344 , n37345 , n37346 , n37347 , n37348 , n37349 , n37350 , n37351 , n37352 , n37353 , n37354 , n37355 , n37356 , n37357 , n37358 , n37359 , n37360 , n37361 , n37362 , n37363 , n37364 , n37365 , n37366 , n37367 , n37368 , n37369 , n37370 , n37371 , n37372 , n37373 , n37374 , n37375 , n37376 , n37377 , n37378 , n37379 , n37380 , n37381 , n37382 , n37383 , n37384 , n37385 , n37386 , n37387 , n37388 , n37389 , n37390 , n37391 , n37392 , n37393 , n37394 , n37395 , n37396 , n37397 , n37398 , n37399 , n37400 , n37401 , n37402 , n37403 , n37404 , n37405 , n37406 , n37407 , n37408 , n37409 , n37410 , n37411 , n37412 , n37413 , n37414 , n37415 , n37416 , n37417 , n37418 , n37419 , n37420 , n37421 , n37422 , n37423 , n37424 , n37425 , n37426 , n37427 , n37428 , n37429 , n37430 , n37431 , n37432 , n37433 , n37434 , n37435 , n37436 , n37437 , n37438 , n37439 , n37440 , n37441 , n37442 , n37443 , n37444 , n37445 , n37446 , n37447 , n37448 , n37449 , n37450 , n37451 , n37452 , n37453 , n37454 , n37455 , n37456 , n37457 , n37458 , n37459 , n37460 , n37461 , n37462 , n37463 , n37464 , n37465 , n37466 , n37467 , n37468 , n37469 , n37470 , n37471 , n37472 , n37473 , n37474 , n37475 , n37476 , n37477 , n37478 , n37479 , n37480 , n37481 , n37482 , n37483 , n37484 , n37485 , n37486 , n37487 , n37488 , n37489 , n37490 , n37491 , n37492 , n37493 , n37494 , n37495 , n37496 , n37497 , n37498 , n37499 , n37500 , n37501 , n37502 , n37503 , n37504 , n37505 , n37506 , n37507 , n37508 , n37509 , n37510 , n37511 , n37512 , n37513 , n37514 , n37515 , n37516 , n37517 , n37518 , n37519 , n37520 , n37521 , n37522 , n37523 , n37524 , n37525 , n37526 , n37527 , n37528 , n37529 , n37530 , n37531 , n37532 , n37533 , n37534 , n37535 , n37536 , n37537 , n37538 , n37539 , n37540 , n37541 , n37542 , n37543 , n37544 , n37545 , n37546 , n37547 , n37548 , n37549 , n37550 , n37551 , n37552 , n37553 , n37554 , n37555 , n37556 , n37557 , n37558 , n37559 , n37560 , n37561 , n37562 , n37563 , n37564 , n37565 , n37566 , n37567 , n37568 , n37569 , n37570 , n37571 , n37572 , n37573 , n37574 , n37575 , n37576 , n37577 , n37578 , n37579 , n37580 , n37581 , n37582 , n37583 , n37584 , n37585 , n37586 , n37587 , n37588 , n37589 , n37590 , n37591 , n37592 , n37593 , n37594 , n37595 , n37596 , n37597 , n37598 , n37599 , n37600 , n37601 , n37602 , n37603 , n37604 , n37605 , n37606 , n37607 , n37608 , n37609 , n37610 , n37611 , n37612 , n37613 , n37614 , n37615 , n37616 , n37617 , n37618 , n37619 , n37620 , n37621 , n37622 , n37623 , n37624 , n37625 , n37626 , n37627 , n37628 , n37629 , n37630 , n37631 , n37632 , n37633 , n37634 , n37635 , n37636 , n37637 , n37638 , n37639 , n37640 , n37641 , n37642 , n37643 , n37644 , n37645 , n37646 , n37647 , n37648 , n37649 , n37650 , n37651 , n37652 , n37653 , n37654 , n37655 , n37656 , n37657 , n37658 , n37659 , n37660 , n37661 , n37662 , n37663 , n37664 , n37665 , n37666 , n37667 , n37668 , n37669 , n37670 , n37671 , n37672 , n37673 , n37674 , n37675 , n37676 , n37677 , n37678 , n37679 , n37680 , n37681 , n37682 , n37683 , n37684 , n37685 , n37686 , n37687 , n37688 , n37689 , n37690 , n37691 , n37692 , n37693 , n37694 , n37695 , n37696 , n37697 , n37698 , n37699 , n37700 , n37701 , n37702 , n37703 , n37704 , n37705 , n37706 , n37707 , n37708 , n37709 , n37710 , n37711 , n37712 , n37713 , n37714 , n37715 , n37716 , n37717 , n37718 , n37719 , n37720 , n37721 , n37722 , n37723 , n37724 , n37725 , n37726 , n37727 , n37728 , n37729 , n37730 , n37731 , n37732 , n37733 , n37734 , n37735 , n37736 , n37737 , n37738 , n37739 , n37740 , n37741 , n37742 , n37743 , n37744 , n37745 , n37746 , n37747 , n37748 , n37749 , n37750 , n37751 , n37752 , n37753 , n37754 , n37755 , n37756 , n37757 , n37758 , n37759 , n37760 , n37761 , n37762 , n37763 , n37764 , n37765 , n37766 , n37767 , n37768 , n37769 , n37770 , n37771 , n37772 , n37773 , n37774 , n37775 , n37776 , n37777 , n37778 , n37779 , n37780 , n37781 , n37782 , n37783 , n37784 , n37785 , n37786 , n37787 , n37788 , n37789 , n37790 , n37791 , n37792 , n37793 , n37794 , n37795 , n37796 , n37797 , n37798 , n37799 , n37800 , n37801 , n37802 , n37803 , n37804 , n37805 , n37806 , n37807 , n37808 , n37809 , n37810 , n37811 , n37812 , n37813 , n37814 , n37815 , n37816 , n37817 , n37818 , n37819 , n37820 , n37821 , n37822 , n37823 , n37824 , n37825 , n37826 , n37827 , n37828 , n37829 , n37830 , n37831 , n37832 , n37833 , n37834 , n37835 , n37836 , n37837 , n37838 , n37839 , n37840 , n37841 , n37842 , n37843 , n37844 , n37845 , n37846 , n37847 , n37848 , n37849 , n37850 , n37851 , n37852 , n37853 , n37854 , n37855 , n37856 , n37857 , n37858 , n37859 , n37860 , n37861 , n37862 , n37863 , n37864 , n37865 , n37866 , n37867 , n37868 , n37869 , n37870 , n37871 , n37872 , n37873 , n37874 , n37875 , n37876 , n37877 , n37878 , n37879 , n37880 , n37881 , n37882 , n37883 , n37884 , n37885 , n37886 , n37887 , n37888 , n37889 , n37890 , n37891 , n37892 , n37893 , n37894 , n37895 , n37896 , n37897 , n37898 , n37899 , n37900 , n37901 , n37902 , n37903 , n37904 , n37905 , n37906 , n37907 , n37908 , n37909 , n37910 , n37911 , n37912 , n37913 , n37914 , n37915 , n37916 , n37917 , n37918 , n37919 , n37920 , n37921 , n37922 , n37923 , n37924 , n37925 , n37926 , n37927 , n37928 , n37929 , n37930 , n37931 , n37932 , n37933 , n37934 , n37935 , n37936 , n37937 , n37938 , n37939 , n37940 , n37941 , n37942 , n37943 , n37944 , n37945 , n37946 , n37947 , n37948 , n37949 , n37950 , n37951 , n37952 , n37953 , n37954 , n37955 , n37956 , n37957 , n37958 , n37959 , n37960 , n37961 , n37962 , n37963 , n37964 , n37965 , n37966 , n37967 , n37968 , n37969 , n37970 , n37971 , n37972 , n37973 , n37974 , n37975 , n37976 , n37977 , n37978 , n37979 , n37980 , n37981 , n37982 , n37983 , n37984 , n37985 , n37986 , n37987 , n37988 , n37989 , n37990 , n37991 , n37992 , n37993 , n37994 , n37995 , n37996 , n37997 , n37998 , n37999 , n38000 , n38001 , n38002 , n38003 , n38004 , n38005 , n38006 , n38007 , n38008 , n38009 , n38010 , n38011 , n38012 , n38013 , n38014 , n38015 , n38016 , n38017 , n38018 , n38019 , n38020 , n38021 , n38022 , n38023 , n38024 , n38025 , n38026 , n38027 , n38028 , n38029 , n38030 , n38031 , n38032 , n38033 , n38034 , n38035 , n38036 , n38037 , n38038 , n38039 , n38040 , n38041 , n38042 , n38043 , n38044 , n38045 , n38046 , n38047 , n38048 , n38049 , n38050 , n38051 , n38052 , n38053 , n38054 , n38055 , n38056 , n38057 , n38058 , n38059 , n38060 , n38061 , n38062 , n38063 , n38064 , n38065 , n38066 , n38067 , n38068 , n38069 , n38070 , n38071 , n38072 , n38073 , n38074 , n38075 , n38076 , n38077 , n38078 , n38079 , n38080 , n38081 , n38082 , n38083 , n38084 , n38085 , n38086 , n38087 , n38088 , n38089 , n38090 , n38091 , n38092 , n38093 , n38094 , n38095 , n38096 , n38097 , n38098 , n38099 , n38100 , n38101 , n38102 , n38103 , n38104 , n38105 , n38106 , n38107 , n38108 , n38109 , n38110 , n38111 , n38112 , n38113 , n38114 , n38115 , n38116 , n38117 , n38118 , n38119 , n38120 , n38121 , n38122 , n38123 , n38124 , n38125 , n38126 , n38127 , n38128 , n38129 , n38130 , n38131 , n38132 , n38133 , n38134 , n38135 , n38136 , n38137 , n38138 , n38139 , n38140 , n38141 , n38142 , n38143 , n38144 , n38145 , n38146 , n38147 , n38148 , n38149 , n38150 , n38151 , n38152 , n38153 , n38154 , n38155 , n38156 , n38157 , n38158 , n38159 , n38160 , n38161 , n38162 , n38163 , n38164 , n38165 , n38166 , n38167 , n38168 , n38169 , n38170 , n38171 , n38172 , n38173 , n38174 , n38175 , n38176 , n38177 , n38178 , n38179 , n38180 , n38181 , n38182 , n38183 , n38184 , n38185 , n38186 , n38187 , n38188 , n38189 , n38190 , n38191 , n38192 , n38193 , n38194 , n38195 , n38196 , n38197 , n38198 , n38199 , n38200 , n38201 , n38202 , n38203 , n38204 , n38205 , n38206 , n38207 , n38208 , n38209 , n38210 , n38211 , n38212 , n38213 , n38214 , n38215 , n38216 , n38217 , n38218 , n38219 , n38220 , n38221 , n38222 , n38223 , n38224 , n38225 , n38226 , n38227 , n38228 , n38229 , n38230 , n38231 , n38232 , n38233 , n38234 , n38235 , n38236 , n38237 , n38238 , n38239 , n38240 , n38241 , n38242 , n38243 , n38244 , n38245 , n38246 , n38247 , n38248 , n38249 , n38250 , n38251 , n38252 , n38253 , n38254 , n38255 , n38256 , n38257 , n38258 , n38259 , n38260 , n38261 , n38262 , n38263 , n38264 , n38265 , n38266 , n38267 , n38268 , n38269 , n38270 , n38271 , n38272 , n38273 , n38274 , n38275 , n38276 , n38277 , n38278 , n38279 , n38280 , n38281 , n38282 , n38283 , n38284 , n38285 , n38286 , n38287 , n38288 , n38289 , n38290 , n38291 , n38292 , n38293 , n38294 , n38295 , n38296 , n38297 , n38298 , n38299 , n38300 , n38301 , n38302 , n38303 , n38304 , n38305 , n38306 , n38307 , n38308 , n38309 , n38310 , n38311 , n38312 , n38313 , n38314 , n38315 , n38316 , n38317 , n38318 , n38319 , n38320 , n38321 , n38322 , n38323 , n38324 , n38325 , n38326 , n38327 , n38328 , n38329 , n38330 , n38331 , n38332 , n38333 , n38334 , n38335 , n38336 , n38337 , n38338 , n38339 , n38340 , n38341 , n38342 , n38343 , n38344 , n38345 , n38346 , n38347 , n38348 , n38349 , n38350 , n38351 , n38352 , n38353 , n38354 , n38355 , n38356 , n38357 , n38358 , n38359 , n38360 , n38361 , n38362 , n38363 , n38364 , n38365 , n38366 , n38367 , n38368 , n38369 , n38370 , n38371 , n38372 , n38373 , n38374 , n38375 , n38376 , n38377 , n38378 , n38379 , n38380 , n38381 , n38382 , n38383 , n38384 , n38385 , n38386 , n38387 , n38388 , n38389 , n38390 , n38391 , n38392 , n38393 , n38394 , n38395 , n38396 , n38397 , n38398 , n38399 , n38400 , n38401 , n38402 , n38403 , n38404 , n38405 , n38406 , n38407 , n38408 , n38409 , n38410 , n38411 , n38412 , n38413 , n38414 , n38415 , n38416 , n38417 , n38418 , n38419 , n38420 , n38421 , n38422 , n38423 , n38424 , n38425 , n38426 , n38427 , n38428 , n38429 , n38430 , n38431 , n38432 , n38433 , n38434 , n38435 , n38436 , n38437 , n38438 , n38439 , n38440 , n38441 , n38442 , n38443 , n38444 , n38445 , n38446 , n38447 , n38448 , n38449 , n38450 , n38451 , n38452 , n38453 , n38454 , n38455 , n38456 , n38457 , n38458 , n38459 , n38460 , n38461 , n38462 , n38463 , n38464 , n38465 , n38466 , n38467 , n38468 , n38469 , n38470 , n38471 , n38472 , n38473 , n38474 , n38475 , n38476 , n38477 , n38478 , n38479 , n38480 , n38481 , n38482 , n38483 , n38484 , n38485 , n38486 , n38487 , n38488 , n38489 , n38490 , n38491 , n38492 , n38493 , n38494 , n38495 , n38496 , n38497 , n38498 , n38499 , n38500 , n38501 , n38502 , n38503 , n38504 , n38505 , n38506 , n38507 , n38508 , n38509 , n38510 , n38511 , n38512 , n38513 , n38514 , n38515 , n38516 , n38517 , n38518 , n38519 , n38520 , n38521 , n38522 , n38523 , n38524 , n38525 , n38526 , n38527 , n38528 , n38529 , n38530 , n38531 , n38532 , n38533 , n38534 , n38535 , n38536 , n38537 , n38538 , n38539 , n38540 , n38541 , n38542 , n38543 , n38544 , n38545 , n38546 , n38547 , n38548 , n38549 , n38550 , n38551 , n38552 , n38553 , n38554 , n38555 , n38556 , n38557 , n38558 , n38559 , n38560 , n38561 , n38562 , n38563 , n38564 , n38565 , n38566 , n38567 , n38568 , n38569 , n38570 , n38571 , n38572 , n38573 , n38574 , n38575 , n38576 , n38577 , n38578 , n38579 , n38580 , n38581 , n38582 , n38583 , n38584 , n38585 , n38586 , n38587 , n38588 , n38589 , n38590 , n38591 , n38592 , n38593 , n38594 , n38595 , n38596 , n38597 , n38598 , n38599 , n38600 , n38601 , n38602 , n38603 , n38604 , n38605 , n38606 , n38607 , n38608 , n38609 , n38610 , n38611 , n38612 , n38613 , n38614 , n38615 , n38616 , n38617 , n38618 , n38619 , n38620 , n38621 , n38622 , n38623 , n38624 , n38625 , n38626 , n38627 , n38628 , n38629 , n38630 , n38631 , n38632 , n38633 , n38634 , n38635 , n38636 , n38637 , n38638 , n38639 , n38640 , n38641 , n38642 , n38643 , n38644 , n38645 , n38646 , n38647 , n38648 , n38649 , n38650 , n38651 , n38652 , n38653 , n38654 , n38655 , n38656 , n38657 , n38658 , n38659 , n38660 , n38661 , n38662 , n38663 , n38664 , n38665 , n38666 , n38667 , n38668 , n38669 , n38670 , n38671 , n38672 , n38673 , n38674 , n38675 , n38676 , n38677 , n38678 , n38679 , n38680 , n38681 , n38682 , n38683 , n38684 , n38685 , n38686 , n38687 , n38688 , n38689 , n38690 , n38691 , n38692 , n38693 , n38694 , n38695 , n38696 , n38697 , n38698 , n38699 , n38700 , n38701 , n38702 , n38703 , n38704 , n38705 , n38706 , n38707 , n38708 , n38709 , n38710 , n38711 , n38712 , n38713 , n38714 , n38715 , n38716 , n38717 , n38718 , n38719 , n38720 , n38721 , n38722 , n38723 , n38724 , n38725 , n38726 , n38727 , n38728 , n38729 , n38730 , n38731 , n38732 , n38733 , n38734 , n38735 , n38736 , n38737 , n38738 , n38739 , n38740 , n38741 , n38742 , n38743 , n38744 , n38745 , n38746 , n38747 , n38748 , n38749 , n38750 , n38751 , n38752 , n38753 , n38754 , n38755 , n38756 , n38757 , n38758 , n38759 , n38760 , n38761 , n38762 , n38763 , n38764 , n38765 , n38766 , n38767 , n38768 , n38769 , n38770 , n38771 , n38772 , n38773 , n38774 , n38775 , n38776 , n38777 , n38778 , n38779 , n38780 , n38781 , n38782 , n38783 , n38784 , n38785 , n38786 , n38787 , n38788 , n38789 , n38790 , n38791 , n38792 , n38793 , n38794 , n38795 , n38796 , n38797 , n38798 , n38799 , n38800 , n38801 , n38802 , n38803 , n38804 , n38805 , n38806 , n38807 , n38808 , n38809 , n38810 , n38811 , n38812 , n38813 , n38814 , n38815 , n38816 , n38817 , n38818 , n38819 , n38820 , n38821 , n38822 , n38823 , n38824 , n38825 , n38826 , n38827 , n38828 , n38829 , n38830 , n38831 , n38832 , n38833 , n38834 , n38835 , n38836 , n38837 , n38838 , n38839 , n38840 , n38841 , n38842 , n38843 , n38844 , n38845 , n38846 , n38847 , n38848 , n38849 , n38850 , n38851 , n38852 , n38853 , n38854 , n38855 , n38856 , n38857 , n38858 , n38859 , n38860 , n38861 , n38862 , n38863 , n38864 , n38865 , n38866 , n38867 , n38868 , n38869 , n38870 , n38871 , n38872 , n38873 , n38874 , n38875 , n38876 , n38877 , n38878 , n38879 , n38880 , n38881 , n38882 , n38883 , n38884 , n38885 , n38886 , n38887 , n38888 , n38889 , n38890 , n38891 , n38892 , n38893 , n38894 , n38895 , n38896 , n38897 , n38898 , n38899 , n38900 , n38901 , n38902 , n38903 , n38904 , n38905 , n38906 , n38907 , n38908 , n38909 , n38910 , n38911 , n38912 , n38913 , n38914 , n38915 , n38916 , n38917 , n38918 , n38919 , n38920 , n38921 , n38922 , n38923 , n38924 , n38925 , n38926 , n38927 , n38928 , n38929 , n38930 , n38931 , n38932 , n38933 , n38934 , n38935 , n38936 , n38937 , n38938 , n38939 , n38940 , n38941 , n38942 , n38943 , n38944 , n38945 , n38946 , n38947 , n38948 , n38949 , n38950 , n38951 , n38952 , n38953 , n38954 , n38955 , n38956 , n38957 , n38958 , n38959 , n38960 , n38961 , n38962 , n38963 , n38964 , n38965 , n38966 , n38967 , n38968 , n38969 , n38970 , n38971 , n38972 , n38973 , n38974 , n38975 , n38976 , n38977 , n38978 , n38979 , n38980 , n38981 , n38982 , n38983 , n38984 , n38985 , n38986 , n38987 , n38988 , n38989 , n38990 , n38991 , n38992 , n38993 , n38994 , n38995 , n38996 , n38997 , n38998 , n38999 , n39000 , n39001 , n39002 , n39003 , n39004 , n39005 , n39006 , n39007 , n39008 , n39009 , n39010 , n39011 , n39012 , n39013 , n39014 , n39015 , n39016 , n39017 , n39018 , n39019 , n39020 , n39021 , n39022 , n39023 , n39024 , n39025 , n39026 , n39027 , n39028 , n39029 , n39030 , n39031 , n39032 , n39033 , n39034 , n39035 , n39036 , n39037 , n39038 , n39039 , n39040 , n39041 , n39042 , n39043 , n39044 , n39045 , n39046 , n39047 , n39048 , n39049 , n39050 , n39051 , n39052 , n39053 , n39054 , n39055 , n39056 , n39057 , n39058 , n39059 , n39060 , n39061 , n39062 , n39063 , n39064 , n39065 , n39066 , n39067 , n39068 , n39069 , n39070 , n39071 , n39072 , n39073 , n39074 , n39075 , n39076 , n39077 , n39078 , n39079 , n39080 , n39081 , n39082 , n39083 , n39084 , n39085 , n39086 , n39087 , n39088 , n39089 , n39090 , n39091 , n39092 , n39093 , n39094 , n39095 , n39096 , n39097 , n39098 , n39099 , n39100 , n39101 , n39102 , n39103 , n39104 , n39105 , n39106 , n39107 , n39108 , n39109 , n39110 , n39111 , n39112 , n39113 , n39114 , n39115 , n39116 , n39117 , n39118 , n39119 , n39120 , n39121 , n39122 , n39123 , n39124 , n39125 , n39126 , n39127 , n39128 , n39129 , n39130 , n39131 , n39132 , n39133 , n39134 , n39135 , n39136 , n39137 , n39138 , n39139 , n39140 , n39141 , n39142 , n39143 , n39144 , n39145 , n39146 , n39147 , n39148 , n39149 , n39150 , n39151 , n39152 , n39153 , n39154 , n39155 , n39156 , n39157 , n39158 , n39159 , n39160 , n39161 , n39162 , n39163 , n39164 , n39165 , n39166 , n39167 , n39168 , n39169 , n39170 , n39171 , n39172 , n39173 , n39174 , n39175 , n39176 , n39177 , n39178 , n39179 , n39180 , n39181 , n39182 , n39183 , n39184 , n39185 , n39186 , n39187 , n39188 , n39189 , n39190 , n39191 , n39192 , n39193 , n39194 , n39195 , n39196 , n39197 , n39198 , n39199 , n39200 , n39201 , n39202 , n39203 , n39204 , n39205 , n39206 , n39207 , n39208 , n39209 , n39210 , n39211 , n39212 , n39213 , n39214 , n39215 , n39216 , n39217 , n39218 , n39219 , n39220 , n39221 , n39222 , n39223 , n39224 , n39225 , n39226 , n39227 , n39228 , n39229 , n39230 , n39231 , n39232 , n39233 , n39234 , n39235 , n39236 , n39237 , n39238 , n39239 , n39240 , n39241 , n39242 , n39243 , n39244 , n39245 , n39246 , n39247 , n39248 , n39249 , n39250 , n39251 , n39252 , n39253 , n39254 , n39255 , n39256 , n39257 , n39258 , n39259 , n39260 , n39261 , n39262 , n39263 , n39264 , n39265 , n39266 , n39267 , n39268 , n39269 , n39270 , n39271 , n39272 , n39273 , n39274 , n39275 , n39276 , n39277 , n39278 , n39279 , n39280 , n39281 , n39282 , n39283 , n39284 , n39285 , n39286 , n39287 , n39288 , n39289 , n39290 , n39291 , n39292 , n39293 , n39294 , n39295 , n39296 , n39297 , n39298 , n39299 , n39300 , n39301 , n39302 , n39303 , n39304 , n39305 , n39306 , n39307 , n39308 , n39309 , n39310 , n39311 , n39312 , n39313 , n39314 , n39315 , n39316 , n39317 , n39318 , n39319 , n39320 , n39321 , n39322 , n39323 , n39324 , n39325 , n39326 , n39327 , n39328 , n39329 , n39330 , n39331 , n39332 , n39333 , n39334 , n39335 , n39336 , n39337 , n39338 , n39339 , n39340 , n39341 , n39342 , n39343 , n39344 , n39345 , n39346 , n39347 , n39348 , n39349 , n39350 , n39351 , n39352 , n39353 , n39354 , n39355 , n39356 , n39357 , n39358 , n39359 , n39360 , n39361 , n39362 , n39363 , n39364 , n39365 , n39366 , n39367 , n39368 , n39369 , n39370 , n39371 , n39372 , n39373 , n39374 , n39375 , n39376 , n39377 , n39378 , n39379 , n39380 , n39381 , n39382 , n39383 , n39384 , n39385 , n39386 , n39387 , n39388 , n39389 , n39390 , n39391 , n39392 , n39393 , n39394 , n39395 , n39396 , n39397 , n39398 , n39399 , n39400 , n39401 , n39402 , n39403 , n39404 , n39405 , n39406 , n39407 , n39408 , n39409 , n39410 , n39411 , n39412 , n39413 , n39414 , n39415 , n39416 , n39417 , n39418 , n39419 , n39420 , n39421 , n39422 , n39423 , n39424 , n39425 , n39426 , n39427 , n39428 , n39429 , n39430 , n39431 , n39432 , n39433 , n39434 , n39435 , n39436 , n39437 , n39438 , n39439 , n39440 , n39441 , n39442 , n39443 , n39444 , n39445 , n39446 , n39447 , n39448 , n39449 , n39450 , n39451 , n39452 , n39453 , n39454 , n39455 , n39456 , n39457 , n39458 , n39459 , n39460 , n39461 , n39462 , n39463 , n39464 , n39465 , n39466 , n39467 , n39468 , n39469 , n39470 , n39471 , n39472 , n39473 , n39474 , n39475 , n39476 , n39477 , n39478 , n39479 , n39480 , n39481 , n39482 , n39483 , n39484 , n39485 , n39486 , n39487 , n39488 , n39489 , n39490 , n39491 , n39492 , n39493 , n39494 , n39495 , n39496 , n39497 , n39498 , n39499 , n39500 , n39501 , n39502 , n39503 , n39504 , n39505 , n39506 , n39507 , n39508 , n39509 , n39510 , n39511 , n39512 , n39513 , n39514 , n39515 , n39516 , n39517 , n39518 , n39519 , n39520 , n39521 , n39522 , n39523 , n39524 , n39525 , n39526 , n39527 , n39528 , n39529 , n39530 , n39531 , n39532 , n39533 , n39534 , n39535 , n39536 , n39537 , n39538 , n39539 , n39540 , n39541 , n39542 , n39543 , n39544 , n39545 , n39546 , n39547 , n39548 , n39549 , n39550 , n39551 , n39552 , n39553 , n39554 , n39555 , n39556 , n39557 , n39558 , n39559 , n39560 , n39561 , n39562 , n39563 , n39564 , n39565 , n39566 , n39567 , n39568 , n39569 , n39570 , n39571 , n39572 , n39573 , n39574 , n39575 , n39576 , n39577 , n39578 , n39579 , n39580 , n39581 , n39582 , n39583 , n39584 , n39585 , n39586 , n39587 , n39588 , n39589 , n39590 , n39591 , n39592 , n39593 , n39594 , n39595 , n39596 , n39597 , n39598 , n39599 , n39600 , n39601 , n39602 , n39603 , n39604 , n39605 , n39606 , n39607 , n39608 , n39609 , n39610 , n39611 , n39612 , n39613 , n39614 , n39615 , n39616 , n39617 , n39618 , n39619 , n39620 , n39621 , n39622 , n39623 , n39624 , n39625 , n39626 , n39627 , n39628 , n39629 , n39630 , n39631 , n39632 , n39633 , n39634 , n39635 , n39636 , n39637 , n39638 , n39639 , n39640 , n39641 , n39642 , n39643 , n39644 , n39645 , n39646 , n39647 , n39648 , n39649 , n39650 , n39651 , n39652 , n39653 , n39654 , n39655 , n39656 , n39657 , n39658 , n39659 , n39660 , n39661 , n39662 , n39663 , n39664 , n39665 , n39666 , n39667 , n39668 , n39669 , n39670 , n39671 , n39672 , n39673 , n39674 , n39675 , n39676 , n39677 , n39678 , n39679 , n39680 , n39681 , n39682 , n39683 , n39684 , n39685 , n39686 , n39687 , n39688 , n39689 , n39690 , n39691 , n39692 , n39693 , n39694 , n39695 , n39696 , n39697 , n39698 , n39699 , n39700 , n39701 , n39702 , n39703 , n39704 , n39705 , n39706 , n39707 , n39708 , n39709 , n39710 , n39711 , n39712 , n39713 , n39714 , n39715 , n39716 , n39717 , n39718 , n39719 , n39720 , n39721 , n39722 , n39723 , n39724 , n39725 , n39726 , n39727 , n39728 , n39729 , n39730 , n39731 , n39732 , n39733 , n39734 , n39735 , n39736 , n39737 , n39738 , n39739 , n39740 , n39741 , n39742 , n39743 , n39744 , n39745 , n39746 , n39747 , n39748 , n39749 , n39750 , n39751 , n39752 , n39753 , n39754 , n39755 , n39756 , n39757 , n39758 , n39759 , n39760 , n39761 , n39762 , n39763 , n39764 , n39765 , n39766 , n39767 , n39768 , n39769 , n39770 , n39771 , n39772 , n39773 , n39774 , n39775 , n39776 , n39777 , n39778 , n39779 , n39780 , n39781 , n39782 , n39783 , n39784 , n39785 , n39786 , n39787 , n39788 , n39789 , n39790 , n39791 , n39792 , n39793 , n39794 , n39795 , n39796 , n39797 , n39798 , n39799 , n39800 , n39801 , n39802 , n39803 , n39804 , n39805 , n39806 , n39807 , n39808 , n39809 , n39810 , n39811 , n39812 , n39813 , n39814 , n39815 , n39816 , n39817 , n39818 , n39819 , n39820 , n39821 , n39822 , n39823 , n39824 , n39825 , n39826 , n39827 , n39828 , n39829 , n39830 , n39831 , n39832 , n39833 , n39834 , n39835 , n39836 , n39837 , n39838 , n39839 , n39840 , n39841 , n39842 , n39843 , n39844 , n39845 , n39846 , n39847 , n39848 , n39849 , n39850 , n39851 , n39852 , n39853 , n39854 , n39855 , n39856 , n39857 , n39858 , n39859 , n39860 , n39861 , n39862 , n39863 , n39864 , n39865 , n39866 , n39867 , n39868 , n39869 , n39870 , n39871 , n39872 , n39873 , n39874 , n39875 , n39876 , n39877 , n39878 , n39879 , n39880 , n39881 , n39882 , n39883 , n39884 , n39885 , n39886 , n39887 , n39888 , n39889 , n39890 , n39891 , n39892 , n39893 , n39894 , n39895 , n39896 , n39897 , n39898 , n39899 , n39900 , n39901 , n39902 , n39903 , n39904 , n39905 , n39906 , n39907 , n39908 , n39909 , n39910 , n39911 , n39912 , n39913 , n39914 , n39915 , n39916 , n39917 , n39918 , n39919 , n39920 , n39921 , n39922 , n39923 , n39924 , n39925 , n39926 , n39927 , n39928 , n39929 , n39930 , n39931 , n39932 , n39933 , n39934 , n39935 , n39936 , n39937 , n39938 , n39939 , n39940 , n39941 , n39942 , n39943 , n39944 , n39945 , n39946 , n39947 , n39948 , n39949 , n39950 , n39951 , n39952 , n39953 , n39954 , n39955 , n39956 , n39957 , n39958 , n39959 , n39960 , n39961 , n39962 , n39963 , n39964 , n39965 , n39966 , n39967 , n39968 , n39969 , n39970 , n39971 , n39972 , n39973 , n39974 , n39975 , n39976 , n39977 , n39978 , n39979 , n39980 , n39981 , n39982 , n39983 , n39984 , n39985 , n39986 , n39987 , n39988 , n39989 , n39990 , n39991 , n39992 , n39993 , n39994 , n39995 , n39996 , n39997 , n39998 , n39999 , n40000 , n40001 , n40002 , n40003 , n40004 , n40005 , n40006 , n40007 , n40008 , n40009 , n40010 , n40011 , n40012 , n40013 , n40014 , n40015 , n40016 , n40017 , n40018 , n40019 , n40020 , n40021 , n40022 , n40023 , n40024 , n40025 , n40026 , n40027 , n40028 , n40029 , n40030 , n40031 , n40032 , n40033 , n40034 , n40035 , n40036 , n40037 , n40038 , n40039 , n40040 , n40041 , n40042 , n40043 , n40044 , n40045 , n40046 , n40047 , n40048 , n40049 , n40050 , n40051 , n40052 , n40053 , n40054 , n40055 , n40056 , n40057 , n40058 , n40059 , n40060 , n40061 , n40062 , n40063 , n40064 , n40065 , n40066 , n40067 , n40068 , n40069 , n40070 , n40071 , n40072 , n40073 , n40074 , n40075 , n40076 , n40077 , n40078 , n40079 , n40080 , n40081 , n40082 , n40083 , n40084 , n40085 , n40086 , n40087 , n40088 , n40089 , n40090 , n40091 , n40092 , n40093 , n40094 , n40095 , n40096 , n40097 , n40098 , n40099 , n40100 , n40101 , n40102 , n40103 , n40104 , n40105 , n40106 , n40107 , n40108 , n40109 , n40110 , n40111 , n40112 , n40113 , n40114 , n40115 , n40116 , n40117 , n40118 , n40119 , n40120 , n40121 , n40122 , n40123 , n40124 , n40125 , n40126 , n40127 , n40128 , n40129 , n40130 , n40131 , n40132 , n40133 , n40134 , n40135 , n40136 , n40137 , n40138 , n40139 , n40140 , n40141 , n40142 , n40143 , n40144 , n40145 , n40146 , n40147 , n40148 , n40149 , n40150 , n40151 , n40152 , n40153 , n40154 , n40155 , n40156 , n40157 , n40158 , n40159 , n40160 , n40161 , n40162 , n40163 , n40164 , n40165 , n40166 , n40167 , n40168 , n40169 , n40170 , n40171 , n40172 , n40173 , n40174 , n40175 , n40176 , n40177 , n40178 , n40179 , n40180 , n40181 , n40182 , n40183 , n40184 , n40185 , n40186 , n40187 , n40188 , n40189 , n40190 , n40191 , n40192 , n40193 , n40194 , n40195 , n40196 , n40197 , n40198 , n40199 , n40200 , n40201 , n40202 , n40203 , n40204 , n40205 , n40206 , n40207 , n40208 , n40209 , n40210 , n40211 , n40212 , n40213 , n40214 , n40215 , n40216 , n40217 , n40218 , n40219 , n40220 , n40221 , n40222 , n40223 , n40224 , n40225 , n40226 , n40227 , n40228 , n40229 , n40230 , n40231 , n40232 , n40233 , n40234 , n40235 , n40236 , n40237 , n40238 , n40239 , n40240 , n40241 , n40242 , n40243 , n40244 , n40245 , n40246 , n40247 , n40248 , n40249 , n40250 , n40251 , n40252 , n40253 , n40254 , n40255 , n40256 , n40257 , n40258 , n40259 , n40260 , n40261 , n40262 , n40263 , n40264 , n40265 , n40266 , n40267 , n40268 , n40269 , n40270 , n40271 , n40272 , n40273 , n40274 , n40275 , n40276 , n40277 , n40278 , n40279 , n40280 , n40281 , n40282 , n40283 , n40284 , n40285 , n40286 , n40287 , n40288 , n40289 , n40290 , n40291 , n40292 , n40293 , n40294 , n40295 , n40296 , n40297 , n40298 , n40299 , n40300 , n40301 , n40302 , n40303 , n40304 , n40305 , n40306 , n40307 , n40308 , n40309 , n40310 , n40311 , n40312 , n40313 , n40314 , n40315 , n40316 , n40317 , n40318 , n40319 , n40320 , n40321 , n40322 , n40323 , n40324 , n40325 , n40326 , n40327 , n40328 , n40329 , n40330 , n40331 , n40332 , n40333 , n40334 , n40335 , n40336 , n40337 , n40338 , n40339 , n40340 , n40341 , n40342 , n40343 , n40344 , n40345 , n40346 , n40347 , n40348 , n40349 , n40350 , n40351 , n40352 , n40353 , n40354 , n40355 , n40356 , n40357 , n40358 , n40359 , n40360 , n40361 , n40362 , n40363 , n40364 , n40365 , n40366 , n40367 , n40368 , n40369 , n40370 , n40371 , n40372 , n40373 , n40374 , n40375 , n40376 , n40377 , n40378 , n40379 , n40380 , n40381 , n40382 , n40383 , n40384 , n40385 , n40386 , n40387 , n40388 , n40389 , n40390 , n40391 , n40392 , n40393 , n40394 , n40395 , n40396 , n40397 , n40398 , n40399 , n40400 , n40401 , n40402 , n40403 , n40404 , n40405 , n40406 , n40407 , n40408 , n40409 , n40410 , n40411 , n40412 , n40413 , n40414 , n40415 , n40416 , n40417 , n40418 , n40419 , n40420 , n40421 , n40422 , n40423 , n40424 , n40425 , n40426 , n40427 , n40428 , n40429 , n40430 , n40431 , n40432 , n40433 , n40434 , n40435 , n40436 , n40437 , n40438 , n40439 , n40440 , n40441 , n40442 , n40443 , n40444 , n40445 , n40446 , n40447 , n40448 , n40449 , n40450 , n40451 , n40452 , n40453 , n40454 , n40455 , n40456 , n40457 , n40458 , n40459 , n40460 , n40461 , n40462 , n40463 , n40464 , n40465 , n40466 , n40467 , n40468 , n40469 , n40470 , n40471 , n40472 , n40473 , n40474 , n40475 , n40476 , n40477 , n40478 , n40479 , n40480 , n40481 , n40482 , n40483 , n40484 , n40485 , n40486 , n40487 , n40488 , n40489 , n40490 , n40491 , n40492 , n40493 , n40494 , n40495 , n40496 , n40497 , n40498 , n40499 , n40500 , n40501 , n40502 , n40503 , n40504 , n40505 , n40506 , n40507 , n40508 , n40509 , n40510 , n40511 , n40512 , n40513 , n40514 , n40515 , n40516 , n40517 , n40518 , n40519 , n40520 , n40521 , n40522 , n40523 , n40524 , n40525 , n40526 , n40527 , n40528 , n40529 , n40530 , n40531 , n40532 , n40533 , n40534 , n40535 , n40536 , n40537 , n40538 , n40539 , n40540 , n40541 , n40542 , n40543 , n40544 , n40545 , n40546 , n40547 , n40548 , n40549 , n40550 , n40551 , n40552 , n40553 , n40554 , n40555 , n40556 , n40557 , n40558 , n40559 , n40560 , n40561 , n40562 , n40563 , n40564 , n40565 , n40566 , n40567 , n40568 , n40569 , n40570 , n40571 , n40572 , n40573 , n40574 , n40575 , n40576 , n40577 , n40578 , n40579 , n40580 , n40581 , n40582 , n40583 , n40584 , n40585 , n40586 , n40587 , n40588 , n40589 , n40590 , n40591 , n40592 , n40593 , n40594 , n40595 , n40596 , n40597 , n40598 , n40599 , n40600 , n40601 , n40602 , n40603 , n40604 , n40605 , n40606 , n40607 , n40608 , n40609 , n40610 , n40611 , n40612 , n40613 , n40614 , n40615 , n40616 , n40617 , n40618 , n40619 , n40620 , n40621 , n40622 , n40623 , n40624 , n40625 , n40626 , n40627 , n40628 , n40629 , n40630 , n40631 , n40632 , n40633 , n40634 , n40635 , n40636 , n40637 , n40638 , n40639 , n40640 , n40641 , n40642 , n40643 , n40644 , n40645 , n40646 , n40647 , n40648 , n40649 , n40650 , n40651 , n40652 , n40653 , n40654 , n40655 , n40656 , n40657 , n40658 , n40659 , n40660 , n40661 , n40662 , n40663 , n40664 , n40665 , n40666 , n40667 , n40668 , n40669 , n40670 , n40671 , n40672 , n40673 , n40674 , n40675 , n40676 , n40677 , n40678 , n40679 , n40680 , n40681 , n40682 , n40683 , n40684 , n40685 , n40686 , n40687 , n40688 , n40689 , n40690 , n40691 , n40692 , n40693 , n40694 , n40695 , n40696 , n40697 , n40698 , n40699 , n40700 , n40701 , n40702 , n40703 , n40704 , n40705 , n40706 , n40707 , n40708 , n40709 , n40710 , n40711 , n40712 , n40713 , n40714 , n40715 , n40716 , n40717 , n40718 , n40719 , n40720 , n40721 , n40722 , n40723 , n40724 , n40725 , n40726 , n40727 , n40728 , n40729 , n40730 , n40731 , n40732 , n40733 , n40734 , n40735 , n40736 , n40737 , n40738 , n40739 , n40740 , n40741 , n40742 , n40743 , n40744 , n40745 , n40746 , n40747 , n40748 , n40749 , n40750 , n40751 , n40752 , n40753 , n40754 , n40755 , n40756 , n40757 , n40758 , n40759 , n40760 , n40761 , n40762 , n40763 , n40764 , n40765 , n40766 , n40767 , n40768 , n40769 , n40770 , n40771 , n40772 , n40773 , n40774 , n40775 , n40776 , n40777 , n40778 , n40779 , n40780 , n40781 , n40782 , n40783 , n40784 , n40785 , n40786 , n40787 , n40788 , n40789 , n40790 , n40791 , n40792 , n40793 , n40794 , n40795 , n40796 , n40797 , n40798 , n40799 , n40800 , n40801 , n40802 , n40803 , n40804 , n40805 , n40806 , n40807 , n40808 , n40809 , n40810 , n40811 , n40812 , n40813 , n40814 , n40815 , n40816 , n40817 , n40818 , n40819 , n40820 , n40821 , n40822 , n40823 , n40824 , n40825 , n40826 , n40827 , n40828 , n40829 , n40830 , n40831 , n40832 , n40833 , n40834 , n40835 , n40836 , n40837 , n40838 , n40839 , n40840 , n40841 , n40842 , n40843 , n40844 , n40845 , n40846 , n40847 , n40848 , n40849 , n40850 , n40851 , n40852 , n40853 , n40854 , n40855 , n40856 , n40857 , n40858 , n40859 , n40860 , n40861 , n40862 , n40863 , n40864 , n40865 , n40866 , n40867 , n40868 , n40869 , n40870 , n40871 , n40872 , n40873 , n40874 , n40875 , n40876 , n40877 , n40878 , n40879 , n40880 , n40881 , n40882 , n40883 , n40884 , n40885 , n40886 , n40887 , n40888 , n40889 , n40890 , n40891 , n40892 , n40893 , n40894 , n40895 , n40896 , n40897 , n40898 , n40899 , n40900 , n40901 , n40902 , n40903 , n40904 , n40905 , n40906 , n40907 , n40908 , n40909 , n40910 , n40911 , n40912 , n40913 , n40914 , n40915 , n40916 , n40917 , n40918 , n40919 , n40920 , n40921 , n40922 , n40923 , n40924 , n40925 , n40926 , n40927 , n40928 , n40929 , n40930 , n40931 , n40932 , n40933 , n40934 , n40935 , n40936 , n40937 , n40938 , n40939 , n40940 , n40941 , n40942 , n40943 , n40944 , n40945 , n40946 , n40947 , n40948 , n40949 , n40950 , n40951 , n40952 , n40953 , n40954 , n40955 , n40956 , n40957 , n40958 , n40959 , n40960 , n40961 , n40962 , n40963 , n40964 , n40965 , n40966 , n40967 , n40968 , n40969 , n40970 , n40971 , n40972 , n40973 , n40974 , n40975 , n40976 , n40977 , n40978 , n40979 , n40980 , n40981 , n40982 , n40983 , n40984 , n40985 , n40986 , n40987 , n40988 , n40989 , n40990 , n40991 , n40992 , n40993 , n40994 , n40995 , n40996 , n40997 , n40998 , n40999 , n41000 , n41001 , n41002 , n41003 , n41004 , n41005 , n41006 , n41007 , n41008 , n41009 , n41010 , n41011 , n41012 , n41013 , n41014 , n41015 , n41016 , n41017 , n41018 , n41019 , n41020 , n41021 , n41022 , n41023 , n41024 , n41025 , n41026 , n41027 , n41028 , n41029 , n41030 , n41031 , n41032 , n41033 , n41034 , n41035 , n41036 , n41037 , n41038 , n41039 , n41040 , n41041 , n41042 , n41043 , n41044 , n41045 , n41046 , n41047 , n41048 , n41049 , n41050 , n41051 , n41052 , n41053 , n41054 , n41055 , n41056 , n41057 , n41058 , n41059 , n41060 , n41061 , n41062 , n41063 , n41064 , n41065 , n41066 , n41067 , n41068 , n41069 , n41070 , n41071 , n41072 , n41073 , n41074 , n41075 , n41076 , n41077 , n41078 , n41079 , n41080 , n41081 , n41082 , n41083 , n41084 , n41085 , n41086 , n41087 , n41088 , n41089 , n41090 , n41091 , n41092 , n41093 , n41094 , n41095 , n41096 , n41097 , n41098 , n41099 , n41100 , n41101 , n41102 , n41103 , n41104 , n41105 , n41106 , n41107 , n41108 , n41109 , n41110 , n41111 , n41112 , n41113 , n41114 , n41115 , n41116 , n41117 , n41118 , n41119 , n41120 , n41121 , n41122 , n41123 , n41124 , n41125 , n41126 , n41127 , n41128 , n41129 , n41130 , n41131 , n41132 , n41133 , n41134 , n41135 , n41136 , n41137 , n41138 , n41139 , n41140 , n41141 , n41142 , n41143 , n41144 , n41145 , n41146 , n41147 , n41148 , n41149 , n41150 , n41151 , n41152 , n41153 , n41154 , n41155 , n41156 , n41157 , n41158 , n41159 , n41160 , n41161 , n41162 , n41163 , n41164 , n41165 , n41166 , n41167 , n41168 , n41169 , n41170 , n41171 , n41172 , n41173 , n41174 , n41175 , n41176 , n41177 , n41178 , n41179 , n41180 , n41181 , n41182 , n41183 , n41184 , n41185 , n41186 , n41187 , n41188 , n41189 , n41190 , n41191 , n41192 , n41193 , n41194 , n41195 , n41196 , n41197 , n41198 , n41199 , n41200 , n41201 , n41202 , n41203 , n41204 , n41205 , n41206 , n41207 , n41208 , n41209 , n41210 , n41211 , n41212 , n41213 , n41214 , n41215 , n41216 , n41217 , n41218 , n41219 , n41220 , n41221 , n41222 , n41223 , n41224 , n41225 , n41226 , n41227 , n41228 , n41229 , n41230 , n41231 , n41232 , n41233 , n41234 , n41235 , n41236 , n41237 , n41238 , n41239 , n41240 , n41241 , n41242 , n41243 , n41244 , n41245 , n41246 , n41247 , n41248 , n41249 , n41250 , n41251 , n41252 , n41253 , n41254 , n41255 , n41256 , n41257 , n41258 , n41259 , n41260 , n41261 , n41262 , n41263 , n41264 , n41265 , n41266 , n41267 , n41268 , n41269 , n41270 , n41271 , n41272 , n41273 , n41274 , n41275 , n41276 , n41277 , n41278 , n41279 , n41280 , n41281 , n41282 , n41283 , n41284 , n41285 , n41286 , n41287 , n41288 , n41289 , n41290 , n41291 , n41292 , n41293 , n41294 , n41295 , n41296 , n41297 , n41298 , n41299 , n41300 , n41301 , n41302 , n41303 , n41304 , n41305 , n41306 , n41307 , n41308 , n41309 , n41310 , n41311 , n41312 , n41313 , n41314 , n41315 , n41316 , n41317 , n41318 , n41319 , n41320 , n41321 , n41322 , n41323 , n41324 , n41325 , n41326 , n41327 , n41328 , n41329 , n41330 , n41331 , n41332 , n41333 , n41334 , n41335 , n41336 , n41337 , n41338 , n41339 , n41340 , n41341 , n41342 , n41343 , n41344 , n41345 , n41346 , n41347 , n41348 , n41349 , n41350 , n41351 , n41352 , n41353 , n41354 , n41355 , n41356 , n41357 , n41358 , n41359 , n41360 , n41361 , n41362 , n41363 , n41364 , n41365 , n41366 , n41367 , n41368 , n41369 , n41370 , n41371 , n41372 , n41373 , n41374 , n41375 , n41376 , n41377 , n41378 , n41379 , n41380 , n41381 , n41382 , n41383 , n41384 , n41385 , n41386 , n41387 , n41388 , n41389 , n41390 , n41391 , n41392 , n41393 , n41394 , n41395 , n41396 , n41397 , n41398 , n41399 , n41400 , n41401 , n41402 , n41403 , n41404 , n41405 , n41406 , n41407 , n41408 , n41409 , n41410 , n41411 , n41412 , n41413 , n41414 , n41415 , n41416 , n41417 , n41418 , n41419 , n41420 , n41421 , n41422 , n41423 , n41424 , n41425 , n41426 , n41427 , n41428 , n41429 , n41430 , n41431 , n41432 , n41433 , n41434 , n41435 , n41436 , n41437 , n41438 , n41439 , n41440 , n41441 , n41442 , n41443 , n41444 , n41445 , n41446 , n41447 , n41448 , n41449 , n41450 , n41451 , n41452 , n41453 , n41454 , n41455 , n41456 , n41457 , n41458 , n41459 , n41460 , n41461 , n41462 , n41463 , n41464 , n41465 , n41466 , n41467 , n41468 , n41469 , n41470 , n41471 , n41472 , n41473 , n41474 , n41475 , n41476 , n41477 , n41478 , n41479 , n41480 , n41481 , n41482 , n41483 , n41484 , n41485 , n41486 , n41487 , n41488 , n41489 , n41490 , n41491 , n41492 , n41493 , n41494 , n41495 , n41496 , n41497 , n41498 , n41499 , n41500 , n41501 , n41502 , n41503 , n41504 , n41505 , n41506 , n41507 , n41508 , n41509 , n41510 , n41511 , n41512 , n41513 , n41514 , n41515 , n41516 , n41517 , n41518 , n41519 , n41520 , n41521 , n41522 , n41523 , n41524 , n41525 , n41526 , n41527 , n41528 , n41529 , n41530 , n41531 , n41532 , n41533 , n41534 , n41535 , n41536 , n41537 , n41538 , n41539 , n41540 , n41541 , n41542 , n41543 , n41544 , n41545 , n41546 , n41547 , n41548 , n41549 , n41550 , n41551 , n41552 , n41553 , n41554 , n41555 , n41556 , n41557 , n41558 , n41559 , n41560 , n41561 , n41562 , n41563 , n41564 , n41565 , n41566 , n41567 , n41568 , n41569 , n41570 , n41571 , n41572 , n41573 , n41574 , n41575 , n41576 , n41577 , n41578 , n41579 , n41580 , n41581 , n41582 , n41583 , n41584 , n41585 , n41586 , n41587 , n41588 , n41589 , n41590 , n41591 , n41592 , n41593 , n41594 , n41595 , n41596 , n41597 , n41598 , n41599 , n41600 , n41601 , n41602 , n41603 , n41604 , n41605 , n41606 , n41607 , n41608 , n41609 , n41610 , n41611 , n41612 , n41613 , n41614 , n41615 , n41616 , n41617 , n41618 , n41619 , n41620 , n41621 , n41622 , n41623 , n41624 , n41625 , n41626 , n41627 , n41628 , n41629 , n41630 , n41631 , n41632 , n41633 , n41634 , n41635 , n41636 , n41637 , n41638 , n41639 , n41640 , n41641 , n41642 , n41643 , n41644 , n41645 , n41646 , n41647 , n41648 , n41649 , n41650 , n41651 , n41652 , n41653 , n41654 , n41655 , n41656 , n41657 , n41658 , n41659 , n41660 , n41661 , n41662 , n41663 , n41664 , n41665 , n41666 , n41667 , n41668 , n41669 , n41670 , n41671 , n41672 , n41673 , n41674 , n41675 , n41676 , n41677 , n41678 , n41679 , n41680 , n41681 , n41682 , n41683 , n41684 , n41685 , n41686 , n41687 , n41688 , n41689 , n41690 , n41691 , n41692 , n41693 , n41694 , n41695 , n41696 , n41697 , n41698 , n41699 , n41700 , n41701 , n41702 , n41703 , n41704 , n41705 , n41706 , n41707 , n41708 , n41709 , n41710 , n41711 , n41712 , n41713 , n41714 , n41715 , n41716 , n41717 , n41718 , n41719 , n41720 , n41721 , n41722 , n41723 , n41724 , n41725 , n41726 , n41727 , n41728 , n41729 , n41730 , n41731 , n41732 , n41733 , n41734 , n41735 , n41736 , n41737 , n41738 , n41739 , n41740 , n41741 , n41742 , n41743 ;
  assign n13 = x6 & x7 ;
  assign n14 = ~x2 & n13 ;
  assign n15 = ( x1 & x5 ) | ( x1 & ~x10 ) | ( x5 & ~x10 ) ;
  assign n16 = n15 ^ x10 ^ 1'b0 ;
  assign n17 = x9 & ~n16 ;
  assign n18 = x3 & ~n17 ;
  assign n19 = ~x8 & n18 ;
  assign n20 = x4 & n16 ;
  assign n21 = n20 ^ n19 ^ 1'b0 ;
  assign n22 = x7 & ~n17 ;
  assign n23 = n22 ^ x2 ^ 1'b0 ;
  assign n24 = n23 ^ x8 ^ 1'b0 ;
  assign n25 = ( ~x0 & n21 ) | ( ~x0 & n24 ) | ( n21 & n24 ) ;
  assign n26 = n17 ^ x4 ^ 1'b0 ;
  assign n27 = x7 & ~n26 ;
  assign n28 = x0 & ~n24 ;
  assign n30 = x7 ^ x6 ^ x5 ;
  assign n31 = x3 & x7 ;
  assign n32 = n31 ^ x5 ^ 1'b0 ;
  assign n33 = n30 | n32 ;
  assign n34 = n33 ^ x1 ^ 1'b0 ;
  assign n35 = x5 & n34 ;
  assign n29 = x9 & ~n24 ;
  assign n36 = n35 ^ n29 ^ 1'b0 ;
  assign n37 = x8 ^ x0 ^ 1'b0 ;
  assign n38 = ~n21 & n37 ;
  assign n39 = n38 ^ x7 ^ 1'b0 ;
  assign n40 = x11 & n39 ;
  assign n41 = ~n23 & n40 ;
  assign n42 = ~x2 & n41 ;
  assign n43 = x1 & n16 ;
  assign n44 = ~n32 & n43 ;
  assign n45 = n43 ^ n28 ^ 1'b0 ;
  assign n46 = x3 & n45 ;
  assign n47 = ~n16 & n40 ;
  assign n48 = n47 ^ n44 ^ 1'b0 ;
  assign n49 = n21 ^ x0 ^ 1'b0 ;
  assign n50 = n34 & n49 ;
  assign n51 = n50 ^ n14 ^ 1'b0 ;
  assign n52 = ~x5 & x8 ;
  assign n53 = ( n17 & n35 ) | ( n17 & n52 ) | ( n35 & n52 ) ;
  assign n54 = ~n17 & n34 ;
  assign n55 = n54 ^ n15 ^ 1'b0 ;
  assign n56 = x4 & x11 ;
  assign n57 = ~n23 & n56 ;
  assign n58 = n57 ^ n27 ^ 1'b0 ;
  assign n59 = x2 & ~n37 ;
  assign n60 = n59 ^ x3 ^ 1'b0 ;
  assign n61 = x1 & ~n60 ;
  assign n62 = n61 ^ x10 ^ 1'b0 ;
  assign n68 = n47 ^ n23 ^ 1'b0 ;
  assign n69 = n68 ^ n56 ^ 1'b0 ;
  assign n63 = ~n17 & n38 ;
  assign n64 = n25 & n63 ;
  assign n65 = n16 & ~n64 ;
  assign n66 = n65 ^ n21 ^ 1'b0 ;
  assign n67 = n24 | n66 ;
  assign n70 = n69 ^ n67 ^ 1'b0 ;
  assign n71 = n16 & ~n35 ;
  assign n72 = n71 ^ n25 ^ 1'b0 ;
  assign n73 = ~x0 & x8 ;
  assign n74 = ~x4 & n15 ;
  assign n75 = n74 ^ x4 ^ 1'b0 ;
  assign n76 = ( ~n40 & n73 ) | ( ~n40 & n75 ) | ( n73 & n75 ) ;
  assign n77 = n19 ^ x8 ^ 1'b0 ;
  assign n78 = n40 | n77 ;
  assign n79 = ~n62 & n78 ;
  assign n80 = ( ~x4 & x7 ) | ( ~x4 & n17 ) | ( x7 & n17 ) ;
  assign n81 = n46 & n80 ;
  assign n82 = x7 & ~n43 ;
  assign n83 = x2 & x4 ;
  assign n84 = n44 & n83 ;
  assign n85 = n84 ^ n83 ^ 1'b0 ;
  assign n86 = x3 | n80 ;
  assign n87 = ( x4 & ~n19 ) | ( x4 & n86 ) | ( ~n19 & n86 ) ;
  assign n90 = n19 & ~n32 ;
  assign n91 = x6 & ~n14 ;
  assign n92 = ~n21 & n91 ;
  assign n93 = n34 & ~n92 ;
  assign n94 = n90 & n93 ;
  assign n88 = n30 ^ n25 ^ 1'b0 ;
  assign n89 = n88 ^ n35 ^ 1'b0 ;
  assign n95 = n94 ^ n89 ^ 1'b0 ;
  assign n96 = n35 | n95 ;
  assign n97 = x10 & ~n37 ;
  assign n98 = ~n83 & n97 ;
  assign n99 = x9 & n37 ;
  assign n100 = ~n37 & n99 ;
  assign n101 = n56 & ~n100 ;
  assign n102 = n36 & ~n101 ;
  assign n103 = ~n92 & n102 ;
  assign n104 = n103 ^ n19 ^ 1'b0 ;
  assign n105 = n75 ^ n24 ^ 1'b0 ;
  assign n106 = n15 & ~n38 ;
  assign n107 = ~x7 & n34 ;
  assign n108 = n107 ^ x11 ^ 1'b0 ;
  assign n109 = n52 & ~n108 ;
  assign n110 = n55 | n106 ;
  assign n111 = n110 ^ n47 ^ 1'b0 ;
  assign n112 = n64 ^ x2 ^ 1'b0 ;
  assign n113 = n37 & ~n112 ;
  assign n114 = x9 & ~n55 ;
  assign n115 = ~n24 & n88 ;
  assign n116 = n115 ^ x3 ^ 1'b0 ;
  assign n117 = n40 ^ n25 ^ 1'b0 ;
  assign n118 = n15 & ~n19 ;
  assign n119 = n118 ^ n101 ^ 1'b0 ;
  assign n120 = ~n37 & n119 ;
  assign n121 = n15 & n43 ;
  assign n122 = ~n30 & n43 ;
  assign n123 = ( n55 & n121 ) | ( n55 & ~n122 ) | ( n121 & ~n122 ) ;
  assign n124 = n98 & n123 ;
  assign n125 = n124 ^ n81 ^ 1'b0 ;
  assign n127 = x0 & ~n69 ;
  assign n128 = ~n37 & n127 ;
  assign n126 = n82 & ~n116 ;
  assign n129 = n128 ^ n126 ^ 1'b0 ;
  assign n130 = n108 ^ n40 ^ 1'b0 ;
  assign n131 = x6 | n119 ;
  assign n132 = n28 & n55 ;
  assign n133 = n132 ^ x7 ^ 1'b0 ;
  assign n134 = n70 ^ x9 ^ 1'b0 ;
  assign n135 = n50 & ~n134 ;
  assign n136 = n135 ^ n44 ^ 1'b0 ;
  assign n137 = n105 & n136 ;
  assign n138 = n123 & n137 ;
  assign n139 = n138 ^ n27 ^ 1'b0 ;
  assign n140 = n90 ^ n89 ^ 1'b0 ;
  assign n141 = n37 | n140 ;
  assign n142 = ~n96 & n141 ;
  assign n143 = n73 & n129 ;
  assign n144 = n25 & n143 ;
  assign n145 = n106 | n144 ;
  assign n146 = n48 & ~n145 ;
  assign n147 = x0 & x9 ;
  assign n148 = n147 ^ n111 ^ 1'b0 ;
  assign n149 = n43 ^ n38 ^ 1'b0 ;
  assign n150 = ~n86 & n149 ;
  assign n151 = ~x2 & n150 ;
  assign n152 = n55 ^ n50 ^ 1'b0 ;
  assign n153 = n52 & ~n152 ;
  assign n154 = n151 | n153 ;
  assign n155 = n40 & ~n117 ;
  assign n156 = n15 & n141 ;
  assign n157 = ~n37 & n83 ;
  assign n158 = n135 ^ n87 ^ n56 ;
  assign n159 = n32 ^ n25 ^ 1'b0 ;
  assign n160 = x2 & n159 ;
  assign n161 = n160 ^ n32 ^ 1'b0 ;
  assign n162 = ~n32 & n161 ;
  assign n163 = ~x6 & n162 ;
  assign n164 = ( n85 & n123 ) | ( n85 & n163 ) | ( n123 & n163 ) ;
  assign n165 = n15 | n70 ;
  assign n166 = x8 & n87 ;
  assign n167 = n32 & n166 ;
  assign n168 = n81 ^ x0 ^ 1'b0 ;
  assign n169 = n17 & ~n69 ;
  assign n170 = n36 | n169 ;
  assign n171 = n117 | n141 ;
  assign n172 = x3 | n171 ;
  assign n173 = n135 & n172 ;
  assign n174 = ~n102 & n173 ;
  assign n175 = ~n30 & n146 ;
  assign n176 = ~n42 & n129 ;
  assign n177 = ~n37 & n176 ;
  assign n178 = n151 & ~n177 ;
  assign n179 = n17 | n130 ;
  assign n180 = n155 & n179 ;
  assign n181 = n72 & ~n89 ;
  assign n182 = n88 & n181 ;
  assign n183 = ~n77 & n117 ;
  assign n184 = n183 ^ n144 ^ n111 ;
  assign n185 = n184 ^ n178 ^ 1'b0 ;
  assign n186 = n170 ^ n135 ^ 1'b0 ;
  assign n187 = n183 ^ n101 ^ n90 ;
  assign n188 = n187 ^ n165 ^ 1'b0 ;
  assign n189 = n28 & ~n58 ;
  assign n190 = n60 & n189 ;
  assign n191 = x4 | n159 ;
  assign n192 = x9 & n191 ;
  assign n193 = x4 | n131 ;
  assign n194 = n106 ^ x6 ^ 1'b0 ;
  assign n195 = n194 ^ n157 ^ 1'b0 ;
  assign n196 = n195 ^ n190 ^ 1'b0 ;
  assign n197 = n153 & n188 ;
  assign n198 = n17 | n81 ;
  assign n202 = n172 ^ n125 ^ 1'b0 ;
  assign n203 = n72 & ~n202 ;
  assign n199 = n55 ^ n52 ^ 1'b0 ;
  assign n200 = n24 | n199 ;
  assign n201 = n131 | n200 ;
  assign n204 = n203 ^ n201 ^ 1'b0 ;
  assign n205 = ~n164 & n204 ;
  assign n206 = n81 & ~n101 ;
  assign n207 = n35 & ~n108 ;
  assign n208 = ( n80 & ~n106 ) | ( n80 & n207 ) | ( ~n106 & n207 ) ;
  assign n209 = n125 | n142 ;
  assign n210 = n209 ^ n190 ^ 1'b0 ;
  assign n211 = n14 | n200 ;
  assign n212 = n94 & ~n211 ;
  assign n213 = n139 ^ n86 ^ 1'b0 ;
  assign n214 = x7 & n213 ;
  assign n215 = n214 ^ x1 ^ 1'b0 ;
  assign n219 = n53 ^ n19 ^ 1'b0 ;
  assign n220 = n137 & n219 ;
  assign n225 = n15 & n220 ;
  assign n226 = n225 ^ n130 ^ 1'b0 ;
  assign n216 = n34 & n117 ;
  assign n217 = n37 | n120 ;
  assign n218 = n216 & ~n217 ;
  assign n221 = n218 ^ n14 ^ 1'b0 ;
  assign n222 = n221 ^ n64 ^ 1'b0 ;
  assign n223 = n220 & n222 ;
  assign n224 = ~n218 & n223 ;
  assign n227 = n226 ^ n224 ^ 1'b0 ;
  assign n228 = ~n75 & n80 ;
  assign n229 = n83 | n190 ;
  assign n230 = n55 & ~n141 ;
  assign n231 = n230 ^ n123 ^ 1'b0 ;
  assign n232 = n141 ^ n92 ^ n55 ;
  assign n233 = n72 & n232 ;
  assign n234 = n191 ^ n50 ^ 1'b0 ;
  assign n235 = n75 ^ x1 ^ 1'b0 ;
  assign n236 = n23 | n32 ;
  assign n237 = n17 | n200 ;
  assign n238 = n44 | n237 ;
  assign n239 = ~n236 & n238 ;
  assign n240 = x10 & ~n239 ;
  assign n241 = ~n104 & n240 ;
  assign n242 = ~n14 & n36 ;
  assign n243 = n239 & n242 ;
  assign n244 = n139 | n243 ;
  assign n245 = n195 ^ n19 ^ 1'b0 ;
  assign n246 = n119 | n245 ;
  assign n247 = n133 & n232 ;
  assign n250 = n55 ^ n28 ^ 1'b0 ;
  assign n248 = n40 & ~n200 ;
  assign n249 = n248 ^ n146 ^ 1'b0 ;
  assign n251 = n250 ^ n249 ^ 1'b0 ;
  assign n252 = n129 ^ n55 ^ 1'b0 ;
  assign n253 = n21 & ~n141 ;
  assign n254 = ~n234 & n252 ;
  assign n257 = n55 ^ n42 ^ 1'b0 ;
  assign n258 = n257 ^ n66 ^ 1'b0 ;
  assign n255 = ( n37 & n88 ) | ( n37 & ~n159 ) | ( n88 & ~n159 ) ;
  assign n256 = n37 & ~n255 ;
  assign n259 = n258 ^ n256 ^ 1'b0 ;
  assign n260 = n168 & ~n259 ;
  assign n261 = n35 & n260 ;
  assign n262 = n207 ^ n19 ^ 1'b0 ;
  assign n263 = n172 & ~n262 ;
  assign n264 = n192 ^ x0 ^ 1'b0 ;
  assign n265 = n263 & ~n264 ;
  assign n267 = n97 & n181 ;
  assign n268 = ~n113 & n267 ;
  assign n269 = n268 ^ n137 ^ 1'b0 ;
  assign n266 = n179 ^ n75 ^ 1'b0 ;
  assign n270 = n269 ^ n266 ^ n83 ;
  assign n271 = n116 & ~n241 ;
  assign n272 = n81 | n169 ;
  assign n273 = n77 ^ x7 ^ 1'b0 ;
  assign n274 = n135 | n179 ;
  assign n275 = n157 & ~n274 ;
  assign n276 = n275 ^ n177 ^ 1'b0 ;
  assign n277 = n276 ^ n210 ^ n19 ;
  assign n278 = n113 & n274 ;
  assign n279 = ~n72 & n153 ;
  assign n280 = n144 & ~n210 ;
  assign n281 = x6 | n280 ;
  assign n282 = ~n142 & n281 ;
  assign n283 = n282 ^ n55 ^ 1'b0 ;
  assign n284 = n216 ^ n37 ^ 1'b0 ;
  assign n285 = n81 & n98 ;
  assign n286 = n285 ^ n186 ^ 1'b0 ;
  assign n287 = n36 ^ x2 ^ 1'b0 ;
  assign n288 = n179 | n287 ;
  assign n289 = x8 & n83 ;
  assign n290 = n289 ^ n81 ^ 1'b0 ;
  assign n291 = n250 | n290 ;
  assign n292 = n42 & ~n77 ;
  assign n293 = n292 ^ n178 ^ n177 ;
  assign n294 = x0 & n86 ;
  assign n295 = n24 & n178 ;
  assign n296 = ~n182 & n287 ;
  assign n297 = n226 ^ n55 ^ 1'b0 ;
  assign n298 = n83 & n297 ;
  assign n299 = n298 ^ n131 ^ 1'b0 ;
  assign n300 = ~n296 & n299 ;
  assign n301 = n142 | n300 ;
  assign n302 = n301 ^ n284 ^ 1'b0 ;
  assign n307 = n114 & ~n137 ;
  assign n308 = n307 ^ n148 ^ 1'b0 ;
  assign n303 = n15 & ~n94 ;
  assign n304 = n131 & n303 ;
  assign n305 = n304 ^ n215 ^ 1'b0 ;
  assign n306 = n129 & n305 ;
  assign n309 = n308 ^ n306 ^ n204 ;
  assign n310 = n105 & ~n144 ;
  assign n311 = n205 ^ n175 ^ 1'b0 ;
  assign n312 = n229 & ~n270 ;
  assign n313 = n312 ^ n283 ^ 1'b0 ;
  assign n314 = n296 ^ n96 ^ 1'b0 ;
  assign n315 = ~n283 & n314 ;
  assign n316 = n268 ^ n177 ^ n168 ;
  assign n318 = n101 ^ n72 ^ 1'b0 ;
  assign n317 = ~n55 & n88 ;
  assign n319 = n318 ^ n317 ^ 1'b0 ;
  assign n320 = n319 ^ n47 ^ 1'b0 ;
  assign n321 = n196 & n320 ;
  assign n322 = n254 & ~n291 ;
  assign n323 = n47 ^ n19 ^ 1'b0 ;
  assign n324 = n148 ^ n19 ^ 1'b0 ;
  assign n325 = n294 ^ n178 ^ 1'b0 ;
  assign n326 = n324 | n325 ;
  assign n327 = n15 | n326 ;
  assign n328 = n258 & ~n323 ;
  assign n331 = ~n86 & n165 ;
  assign n332 = n331 ^ n323 ^ 1'b0 ;
  assign n329 = n47 & n55 ;
  assign n330 = n329 ^ x4 ^ 1'b0 ;
  assign n333 = n332 ^ n330 ^ 1'b0 ;
  assign n334 = n113 & ~n307 ;
  assign n335 = n334 ^ n75 ^ 1'b0 ;
  assign n336 = n268 | n330 ;
  assign n337 = n47 & ~n336 ;
  assign n338 = n216 ^ n196 ^ n182 ;
  assign n339 = n292 & n318 ;
  assign n340 = n62 | n243 ;
  assign n341 = n159 | n324 ;
  assign n342 = n297 | n341 ;
  assign n343 = n111 | n231 ;
  assign n344 = n338 ^ n58 ^ 1'b0 ;
  assign n345 = n175 | n344 ;
  assign n346 = n21 ^ x11 ^ 1'b0 ;
  assign n347 = n156 & n226 ;
  assign n348 = n347 ^ n55 ^ 1'b0 ;
  assign n349 = n348 ^ x3 ^ 1'b0 ;
  assign n350 = n346 & n349 ;
  assign n351 = n27 & ~n191 ;
  assign n352 = n351 ^ x3 ^ 1'b0 ;
  assign n353 = n139 & ~n194 ;
  assign n354 = n273 ^ n107 ^ 1'b0 ;
  assign n355 = n354 ^ n64 ^ 1'b0 ;
  assign n356 = ~n353 & n355 ;
  assign n357 = n92 ^ n74 ^ 1'b0 ;
  assign n358 = n357 ^ n226 ^ 1'b0 ;
  assign n359 = n356 & ~n358 ;
  assign n360 = n97 & ~n159 ;
  assign n361 = n360 ^ n268 ^ 1'b0 ;
  assign n362 = n270 & n315 ;
  assign n363 = ~x6 & n362 ;
  assign n364 = n226 | n363 ;
  assign n365 = x1 & ~n53 ;
  assign n366 = n365 ^ n265 ^ 1'b0 ;
  assign n367 = n83 ^ n25 ^ 1'b0 ;
  assign n368 = n183 ^ n181 ^ 1'b0 ;
  assign n369 = n232 & n368 ;
  assign n370 = ~n102 & n369 ;
  assign n371 = n370 ^ n278 ^ 1'b0 ;
  assign n372 = ~n131 & n223 ;
  assign n373 = n371 & ~n372 ;
  assign n374 = ~n367 & n373 ;
  assign n375 = ~n113 & n208 ;
  assign n376 = x8 & ~n195 ;
  assign n377 = n111 ^ n64 ^ 1'b0 ;
  assign n378 = n299 & ~n377 ;
  assign n379 = n203 ^ n86 ^ 1'b0 ;
  assign n380 = n266 | n379 ;
  assign n381 = n207 & n380 ;
  assign n384 = n274 ^ n117 ^ 1'b0 ;
  assign n382 = n23 | n92 ;
  assign n383 = n348 & ~n382 ;
  assign n385 = n384 ^ n383 ^ 1'b0 ;
  assign n386 = n255 ^ n159 ^ 1'b0 ;
  assign n387 = n346 & ~n386 ;
  assign n388 = n387 ^ n325 ^ 1'b0 ;
  assign n389 = n252 & ~n388 ;
  assign n390 = n109 ^ n88 ^ 1'b0 ;
  assign n391 = n390 ^ n79 ^ 1'b0 ;
  assign n392 = n391 ^ n180 ^ 1'b0 ;
  assign n393 = n392 ^ n47 ^ 1'b0 ;
  assign n394 = n390 ^ n172 ^ 1'b0 ;
  assign n395 = n163 | n394 ;
  assign n396 = n106 | n141 ;
  assign n397 = n114 | n396 ;
  assign n398 = ( n142 & n253 ) | ( n142 & n397 ) | ( n253 & n397 ) ;
  assign n399 = x10 & n15 ;
  assign n400 = n92 & n399 ;
  assign n401 = ~n307 & n387 ;
  assign n402 = n401 ^ n37 ^ 1'b0 ;
  assign n403 = ~x3 & n402 ;
  assign n404 = n281 | n403 ;
  assign n405 = n400 & ~n404 ;
  assign n406 = ( n184 & ~n190 ) | ( n184 & n236 ) | ( ~n190 & n236 ) ;
  assign n407 = ~n277 & n406 ;
  assign n408 = ~n263 & n407 ;
  assign n409 = n78 & n327 ;
  assign n410 = n409 ^ n272 ^ 1'b0 ;
  assign n411 = n290 ^ n266 ^ 1'b0 ;
  assign n412 = n292 & n411 ;
  assign n413 = n170 & n208 ;
  assign n414 = n413 ^ n200 ^ 1'b0 ;
  assign n415 = n270 & n414 ;
  assign n417 = n84 & ~n307 ;
  assign n416 = n27 & n328 ;
  assign n418 = n417 ^ n416 ^ 1'b0 ;
  assign n419 = n86 & n318 ;
  assign n420 = n108 ^ n37 ^ 1'b0 ;
  assign n421 = ~n234 & n420 ;
  assign n422 = n300 ^ n74 ^ 1'b0 ;
  assign n423 = ~x0 & n422 ;
  assign n424 = n17 & n423 ;
  assign n425 = ~n421 & n424 ;
  assign n426 = n55 | n79 ;
  assign n427 = n426 ^ n258 ^ 1'b0 ;
  assign n428 = n62 | n113 ;
  assign n429 = n334 ^ n24 ^ 1'b0 ;
  assign n430 = n92 | n429 ;
  assign n431 = n19 | n430 ;
  assign n432 = n133 & ~n431 ;
  assign n433 = n239 & n412 ;
  assign n434 = n177 ^ x8 ^ 1'b0 ;
  assign n435 = n158 ^ n86 ^ 1'b0 ;
  assign n436 = n284 ^ n114 ^ 1'b0 ;
  assign n437 = n37 & ~n436 ;
  assign n438 = x8 | n114 ;
  assign n439 = ~n235 & n438 ;
  assign n440 = n300 | n439 ;
  assign n441 = n440 ^ n130 ^ 1'b0 ;
  assign n442 = x8 | n258 ;
  assign n443 = n155 ^ n113 ^ 1'b0 ;
  assign n444 = n443 ^ n213 ^ 1'b0 ;
  assign n445 = ~n279 & n444 ;
  assign n446 = n231 & ~n302 ;
  assign n447 = n446 ^ n139 ^ 1'b0 ;
  assign n448 = n52 & ~n447 ;
  assign n449 = n185 ^ n19 ^ 1'b0 ;
  assign n450 = n356 & ~n449 ;
  assign n452 = x10 & n19 ;
  assign n453 = x1 & ~n68 ;
  assign n454 = ~n452 & n453 ;
  assign n451 = n34 | n336 ;
  assign n455 = n454 ^ n451 ^ 1'b0 ;
  assign n456 = n196 & n270 ;
  assign n457 = n55 & n456 ;
  assign n458 = n403 | n457 ;
  assign n459 = n294 ^ n38 ^ n19 ;
  assign n460 = n141 ^ x8 ^ 1'b0 ;
  assign n461 = n177 & ~n460 ;
  assign n462 = n434 ^ n42 ^ 1'b0 ;
  assign n464 = n19 | n163 ;
  assign n465 = n464 ^ n308 ^ 1'b0 ;
  assign n463 = n87 & n232 ;
  assign n466 = n465 ^ n463 ^ 1'b0 ;
  assign n467 = n178 ^ n72 ^ 1'b0 ;
  assign n468 = n191 & ~n467 ;
  assign n469 = n50 & ~n111 ;
  assign n470 = n469 ^ n216 ^ 1'b0 ;
  assign n471 = n382 | n470 ;
  assign n472 = n322 ^ n175 ^ n111 ;
  assign n473 = n426 & ~n472 ;
  assign n474 = n473 ^ n27 ^ 1'b0 ;
  assign n475 = ~n231 & n246 ;
  assign n476 = n426 ^ n89 ^ 1'b0 ;
  assign n477 = n476 ^ n378 ^ 1'b0 ;
  assign n478 = n388 ^ n234 ^ 1'b0 ;
  assign n479 = x10 | n234 ;
  assign n481 = n70 & n73 ;
  assign n480 = x7 & n426 ;
  assign n482 = n481 ^ n480 ^ 1'b0 ;
  assign n484 = n207 ^ n190 ^ 1'b0 ;
  assign n483 = n380 ^ n182 ^ 1'b0 ;
  assign n485 = n484 ^ n483 ^ 1'b0 ;
  assign n486 = n388 & ~n485 ;
  assign n487 = n284 & n486 ;
  assign n488 = n55 & ~n274 ;
  assign n489 = ~n259 & n488 ;
  assign n490 = n72 ^ x0 ^ 1'b0 ;
  assign n491 = ~n23 & n490 ;
  assign n492 = ~n278 & n491 ;
  assign n493 = n475 ^ n461 ^ 1'b0 ;
  assign n494 = n423 ^ n50 ^ 1'b0 ;
  assign n495 = ~n391 & n494 ;
  assign n496 = n86 & n438 ;
  assign n497 = n496 ^ n479 ^ 1'b0 ;
  assign n498 = ~n125 & n191 ;
  assign n499 = n498 ^ n129 ^ 1'b0 ;
  assign n500 = n499 ^ n218 ^ n196 ;
  assign n506 = n19 & n272 ;
  assign n507 = n148 & n506 ;
  assign n501 = ~n85 & n90 ;
  assign n502 = n501 ^ n128 ^ 1'b0 ;
  assign n503 = n195 & ~n502 ;
  assign n504 = n410 | n503 ;
  assign n505 = ~n179 & n504 ;
  assign n508 = n507 ^ n505 ^ 1'b0 ;
  assign n509 = n439 ^ n294 ^ 1'b0 ;
  assign n510 = ~n389 & n503 ;
  assign n511 = n200 ^ n25 ^ 1'b0 ;
  assign n512 = n51 & n511 ;
  assign n513 = n196 & n512 ;
  assign n514 = n107 & ~n513 ;
  assign n515 = n50 & ~n205 ;
  assign n516 = n141 | n353 ;
  assign n517 = n516 ^ n204 ^ 1'b0 ;
  assign n518 = n515 & n517 ;
  assign n519 = ( n205 & n328 ) | ( n205 & ~n517 ) | ( n328 & ~n517 ) ;
  assign n520 = ~n457 & n519 ;
  assign n521 = n419 | n469 ;
  assign n522 = n34 | n521 ;
  assign n523 = n522 ^ n384 ^ 1'b0 ;
  assign n524 = n55 & n523 ;
  assign n525 = n311 ^ n76 ^ 1'b0 ;
  assign n526 = n292 & ~n525 ;
  assign n527 = n129 & n220 ;
  assign n528 = n257 ^ n58 ^ 1'b0 ;
  assign n529 = n271 ^ n55 ^ 1'b0 ;
  assign n530 = n180 | n529 ;
  assign n531 = n376 | n530 ;
  assign n532 = n457 | n531 ;
  assign n533 = x8 & ~n203 ;
  assign n534 = n527 & ~n533 ;
  assign n535 = n459 ^ n241 ^ 1'b0 ;
  assign n536 = x4 | n23 ;
  assign n537 = n36 & ~n536 ;
  assign n538 = n537 ^ n532 ^ 1'b0 ;
  assign n539 = n338 ^ n79 ^ 1'b0 ;
  assign n540 = n249 ^ n121 ^ 1'b0 ;
  assign n541 = n273 | n408 ;
  assign n542 = n205 ^ n23 ^ 1'b0 ;
  assign n543 = n450 ^ n119 ^ 1'b0 ;
  assign n544 = n346 & ~n543 ;
  assign n545 = n179 ^ n114 ^ 1'b0 ;
  assign n546 = n495 ^ n120 ^ 1'b0 ;
  assign n547 = ( n14 & n185 ) | ( n14 & ~n397 ) | ( n185 & ~n397 ) ;
  assign n548 = n547 ^ n37 ^ 1'b0 ;
  assign n549 = ~n546 & n548 ;
  assign n550 = ~n292 & n549 ;
  assign n551 = n545 & n550 ;
  assign n552 = n392 ^ n62 ^ 1'b0 ;
  assign n553 = n545 ^ n78 ^ n38 ;
  assign n554 = n259 ^ n70 ^ 1'b0 ;
  assign n555 = n553 & n554 ;
  assign n556 = n270 & ~n318 ;
  assign n558 = n109 ^ n28 ^ 1'b0 ;
  assign n557 = n294 ^ n40 ^ 1'b0 ;
  assign n559 = n558 ^ n557 ^ 1'b0 ;
  assign n560 = n104 & ~n559 ;
  assign n561 = n556 & n560 ;
  assign n562 = n172 & ~n348 ;
  assign n563 = n221 ^ n47 ^ 1'b0 ;
  assign n564 = n378 & ~n563 ;
  assign n565 = n286 ^ n68 ^ 1'b0 ;
  assign n566 = n254 ^ n119 ^ 1'b0 ;
  assign n567 = ~n223 & n566 ;
  assign n568 = n205 ^ n204 ^ 1'b0 ;
  assign n569 = n174 | n515 ;
  assign n570 = n421 | n569 ;
  assign n571 = ~n153 & n259 ;
  assign n572 = n571 ^ n258 ^ 1'b0 ;
  assign n573 = n570 & n572 ;
  assign n574 = n546 ^ n204 ^ 1'b0 ;
  assign n575 = n340 | n574 ;
  assign n576 = ~n168 & n533 ;
  assign n578 = n227 & n392 ;
  assign n577 = n336 & ~n381 ;
  assign n579 = n578 ^ n577 ^ 1'b0 ;
  assign n580 = ~n528 & n579 ;
  assign n581 = x0 & n270 ;
  assign n582 = ~n239 & n581 ;
  assign n583 = n55 | n210 ;
  assign n584 = n249 | n583 ;
  assign n585 = n337 ^ n185 ^ 1'b0 ;
  assign n586 = n133 | n325 ;
  assign n587 = n586 ^ n510 ^ 1'b0 ;
  assign n588 = n587 ^ n512 ^ n235 ;
  assign n589 = x1 & n51 ;
  assign n590 = n589 ^ n491 ^ 1'b0 ;
  assign n591 = n328 & n590 ;
  assign n592 = n191 ^ n84 ^ 1'b0 ;
  assign n593 = n592 ^ n208 ^ 1'b0 ;
  assign n595 = n321 ^ n62 ^ 1'b0 ;
  assign n594 = n198 | n364 ;
  assign n596 = n595 ^ n594 ^ 1'b0 ;
  assign n597 = n46 ^ n32 ^ 1'b0 ;
  assign n598 = n104 & ~n597 ;
  assign n599 = ~n328 & n598 ;
  assign n600 = n336 ^ n208 ^ 1'b0 ;
  assign n601 = n599 | n600 ;
  assign n602 = ~n84 & n507 ;
  assign n603 = n477 ^ n274 ^ 1'b0 ;
  assign n604 = n85 & n327 ;
  assign n605 = n604 ^ n167 ^ 1'b0 ;
  assign n606 = n185 ^ x7 ^ 1'b0 ;
  assign n607 = ~n425 & n606 ;
  assign n608 = n605 & n607 ;
  assign n609 = n387 ^ n381 ^ 1'b0 ;
  assign n612 = x0 | n58 ;
  assign n613 = n612 ^ n270 ^ 1'b0 ;
  assign n614 = n182 & n613 ;
  assign n610 = n545 ^ n302 ^ 1'b0 ;
  assign n611 = ~n359 & n610 ;
  assign n615 = n614 ^ n611 ^ n46 ;
  assign n616 = n107 & ~n258 ;
  assign n617 = n440 | n616 ;
  assign n618 = n503 | n617 ;
  assign n619 = n618 ^ n322 ^ 1'b0 ;
  assign n620 = n75 | n605 ;
  assign n621 = n547 & ~n620 ;
  assign n622 = n567 ^ n261 ^ 1'b0 ;
  assign n623 = ~n236 & n513 ;
  assign n624 = n623 ^ n621 ^ 1'b0 ;
  assign n625 = ~n55 & n257 ;
  assign n626 = ~n273 & n625 ;
  assign n627 = n121 | n278 ;
  assign n628 = n226 ^ n141 ^ 1'b0 ;
  assign n629 = ~n108 & n506 ;
  assign n630 = n629 ^ n281 ^ 1'b0 ;
  assign n631 = ~n192 & n630 ;
  assign n632 = ~n628 & n631 ;
  assign n633 = n141 & ~n460 ;
  assign n634 = ( n86 & n558 ) | ( n86 & n633 ) | ( n558 & n633 ) ;
  assign n635 = n299 ^ n220 ^ 1'b0 ;
  assign n636 = n249 & n635 ;
  assign n637 = n384 & ~n636 ;
  assign n638 = ~n287 & n476 ;
  assign n639 = ~n37 & n564 ;
  assign n640 = n624 ^ n83 ^ 1'b0 ;
  assign n642 = ( x1 & n208 ) | ( x1 & n270 ) | ( n208 & n270 ) ;
  assign n641 = n588 ^ x8 ^ 1'b0 ;
  assign n643 = n642 ^ n641 ^ 1'b0 ;
  assign n644 = n37 | n122 ;
  assign n645 = ~n66 & n154 ;
  assign n646 = n83 ^ x3 ^ 1'b0 ;
  assign n647 = n645 | n646 ;
  assign n648 = n553 & ~n632 ;
  assign n649 = ~n34 & n648 ;
  assign n651 = n164 & n269 ;
  assign n652 = n286 & n651 ;
  assign n650 = n246 & ~n352 ;
  assign n653 = n652 ^ n650 ^ 1'b0 ;
  assign n654 = n481 ^ n318 ^ 1'b0 ;
  assign n655 = n336 & ~n654 ;
  assign n656 = n655 ^ n235 ^ 1'b0 ;
  assign n657 = n276 ^ n86 ^ 1'b0 ;
  assign n658 = n657 ^ n308 ^ 1'b0 ;
  assign n659 = ~n323 & n658 ;
  assign n660 = n213 & n361 ;
  assign n661 = n660 ^ n348 ^ 1'b0 ;
  assign n662 = n661 ^ n436 ^ 1'b0 ;
  assign n663 = n153 & ~n194 ;
  assign n664 = n236 & n328 ;
  assign n665 = n437 & n455 ;
  assign n666 = n410 ^ n21 ^ 1'b0 ;
  assign n667 = x7 & n666 ;
  assign n668 = n86 | n236 ;
  assign n669 = n278 & ~n668 ;
  assign n670 = n117 | n669 ;
  assign n671 = n76 ^ n75 ^ 1'b0 ;
  assign n672 = n450 ^ n191 ^ 1'b0 ;
  assign n673 = ~n444 & n672 ;
  assign n674 = n232 & n278 ;
  assign n675 = ~n596 & n674 ;
  assign n676 = n161 & n501 ;
  assign n677 = ~n185 & n676 ;
  assign n678 = n677 ^ n608 ^ 1'b0 ;
  assign n679 = n363 ^ n236 ^ 1'b0 ;
  assign n680 = n185 & n414 ;
  assign n681 = n680 ^ n157 ^ 1'b0 ;
  assign n682 = ~n302 & n481 ;
  assign n683 = n682 ^ x10 ^ 1'b0 ;
  assign n684 = n83 & n203 ;
  assign n685 = ~n510 & n684 ;
  assign n686 = n685 ^ n119 ^ 1'b0 ;
  assign n687 = n169 | n686 ;
  assign n688 = n687 ^ n339 ^ 1'b0 ;
  assign n689 = ~n400 & n599 ;
  assign n691 = n109 & ~n114 ;
  assign n690 = n75 & n139 ;
  assign n692 = n691 ^ n690 ^ 1'b0 ;
  assign n693 = n323 ^ n151 ^ 1'b0 ;
  assign n694 = n194 & n693 ;
  assign n695 = n436 | n694 ;
  assign n696 = n695 ^ n190 ^ 1'b0 ;
  assign n697 = ~n692 & n696 ;
  assign n698 = n165 | n678 ;
  assign n699 = n299 ^ n148 ^ 1'b0 ;
  assign n700 = n524 ^ n119 ^ 1'b0 ;
  assign n701 = n497 & ~n509 ;
  assign n702 = n701 ^ n425 ^ n149 ;
  assign n703 = n90 & n568 ;
  assign n704 = n212 ^ n148 ^ 1'b0 ;
  assign n705 = n500 ^ n233 ^ 1'b0 ;
  assign n706 = n191 ^ n159 ^ 1'b0 ;
  assign n707 = n392 & n706 ;
  assign n708 = ( ~n177 & n296 ) | ( ~n177 & n375 ) | ( n296 & n375 ) ;
  assign n709 = n633 ^ n520 ^ 1'b0 ;
  assign n710 = n88 & ~n610 ;
  assign n711 = n255 | n551 ;
  assign n712 = n711 ^ n547 ^ 1'b0 ;
  assign n713 = n388 ^ n194 ^ 1'b0 ;
  assign n714 = n21 & ~n555 ;
  assign n715 = n304 ^ n257 ^ 1'b0 ;
  assign n716 = ~n119 & n715 ;
  assign n717 = n716 ^ n652 ^ 1'b0 ;
  assign n718 = ~n296 & n717 ;
  assign n719 = n718 ^ n55 ^ 1'b0 ;
  assign n720 = n342 & ~n419 ;
  assign n721 = ~n719 & n720 ;
  assign n722 = n169 & n250 ;
  assign n723 = n284 ^ n50 ^ 1'b0 ;
  assign n724 = n268 & n354 ;
  assign n725 = n723 & ~n724 ;
  assign n726 = n725 ^ n375 ^ 1'b0 ;
  assign n727 = ~n102 & n726 ;
  assign n728 = n722 & n727 ;
  assign n729 = n721 & n728 ;
  assign n730 = n694 ^ n518 ^ 1'b0 ;
  assign n731 = ~n92 & n730 ;
  assign n732 = n731 ^ n721 ^ n412 ;
  assign n733 = n68 | n128 ;
  assign n734 = n733 ^ n284 ^ 1'b0 ;
  assign n735 = n55 ^ x2 ^ 1'b0 ;
  assign n736 = n475 & ~n735 ;
  assign n737 = ~n181 & n736 ;
  assign n738 = ( n156 & ~n436 ) | ( n156 & n737 ) | ( ~n436 & n737 ) ;
  assign n739 = n400 & n738 ;
  assign n740 = n734 & n739 ;
  assign n741 = n184 ^ n68 ^ 1'b0 ;
  assign n742 = n318 & ~n741 ;
  assign n743 = ~n336 & n742 ;
  assign n744 = x10 & ~n609 ;
  assign n745 = n47 & ~n310 ;
  assign n746 = n253 & n484 ;
  assign n747 = n745 & n746 ;
  assign n748 = n346 & n677 ;
  assign n749 = n82 ^ x2 ^ 1'b0 ;
  assign n750 = n749 ^ n426 ^ 1'b0 ;
  assign n751 = ( n144 & ~n748 ) | ( n144 & n750 ) | ( ~n748 & n750 ) ;
  assign n752 = ~n294 & n751 ;
  assign n753 = ~n426 & n752 ;
  assign n754 = n694 | n753 ;
  assign n755 = n159 ^ x9 ^ 1'b0 ;
  assign n756 = n129 | n755 ;
  assign n757 = ~n621 & n756 ;
  assign n758 = n191 | n460 ;
  assign n759 = n148 | n758 ;
  assign n760 = ~n294 & n759 ;
  assign n761 = n406 & ~n419 ;
  assign n762 = n761 ^ n412 ^ 1'b0 ;
  assign n763 = ~n384 & n762 ;
  assign n764 = n207 ^ n148 ^ 1'b0 ;
  assign n765 = n130 | n764 ;
  assign n766 = n618 & n764 ;
  assign n767 = n21 & ~n766 ;
  assign n768 = n178 ^ n44 ^ 1'b0 ;
  assign n769 = n557 ^ n393 ^ 1'b0 ;
  assign n770 = ~n768 & n769 ;
  assign n771 = n486 ^ n46 ^ 1'b0 ;
  assign n772 = ~n737 & n771 ;
  assign n773 = n722 ^ n292 ^ 1'b0 ;
  assign n774 = n141 & ~n390 ;
  assign n775 = n481 ^ n371 ^ 1'b0 ;
  assign n776 = ~n94 & n775 ;
  assign n777 = n149 & ~n353 ;
  assign n778 = n777 ^ n79 ^ 1'b0 ;
  assign n779 = n278 | n778 ;
  assign n780 = n170 & ~n779 ;
  assign n781 = n780 ^ n107 ^ 1'b0 ;
  assign n782 = n776 & n781 ;
  assign n783 = n327 & ~n338 ;
  assign n784 = n783 ^ n445 ^ 1'b0 ;
  assign n785 = n266 & n784 ;
  assign n786 = n323 ^ n92 ^ 1'b0 ;
  assign n787 = n194 & ~n786 ;
  assign n788 = n337 & n546 ;
  assign n789 = n310 & n318 ;
  assign n790 = n378 ^ n15 ^ 1'b0 ;
  assign n791 = ~n789 & n790 ;
  assign n792 = n788 & n791 ;
  assign n793 = ~n441 & n576 ;
  assign n794 = n793 ^ n342 ^ 1'b0 ;
  assign n795 = n250 & ~n274 ;
  assign n796 = n795 ^ n332 ^ 1'b0 ;
  assign n797 = n387 ^ x1 ^ 1'b0 ;
  assign n798 = ~n796 & n797 ;
  assign n799 = n404 & n715 ;
  assign n800 = ~n311 & n501 ;
  assign n801 = n142 & ~n654 ;
  assign n802 = ~n800 & n801 ;
  assign n803 = n802 ^ n161 ^ 1'b0 ;
  assign n804 = ~n128 & n803 ;
  assign n805 = n691 ^ n640 ^ 1'b0 ;
  assign n806 = n659 & ~n805 ;
  assign n807 = n781 | n799 ;
  assign n808 = n114 ^ n34 ^ 1'b0 ;
  assign n809 = n122 & n808 ;
  assign n810 = ( ~n69 & n284 ) | ( ~n69 & n809 ) | ( n284 & n809 ) ;
  assign n811 = n92 & n488 ;
  assign n812 = n508 | n811 ;
  assign n813 = n605 | n760 ;
  assign n814 = n144 & ~n164 ;
  assign n815 = n814 ^ n55 ^ 1'b0 ;
  assign n816 = n16 | n524 ;
  assign n817 = ~n296 & n816 ;
  assign n818 = n221 ^ n159 ^ 1'b0 ;
  assign n819 = n818 ^ n389 ^ 1'b0 ;
  assign n820 = n148 | n819 ;
  assign n821 = n540 ^ n313 ^ 1'b0 ;
  assign n822 = n417 | n821 ;
  assign n823 = ~n796 & n822 ;
  assign n824 = n518 & n823 ;
  assign n825 = n824 ^ n77 ^ 1'b0 ;
  assign n826 = ~n210 & n506 ;
  assign n827 = n826 ^ n745 ^ 1'b0 ;
  assign n828 = n306 & ~n827 ;
  assign n829 = n68 | n200 ;
  assign n830 = n829 ^ n182 ^ 1'b0 ;
  assign n831 = ~n310 & n327 ;
  assign n832 = n218 & n831 ;
  assign n833 = n832 ^ n384 ^ 1'b0 ;
  assign n834 = ~n68 & n191 ;
  assign n835 = n822 & n834 ;
  assign n836 = n768 ^ n630 ^ 1'b0 ;
  assign n837 = n835 & n836 ;
  assign n838 = x0 | n690 ;
  assign n839 = n837 & ~n838 ;
  assign n840 = n495 ^ n468 ^ 1'b0 ;
  assign n841 = n618 | n840 ;
  assign n842 = x0 & ~n89 ;
  assign n843 = ~n190 & n842 ;
  assign n844 = n40 & ~n461 ;
  assign n845 = n414 & ~n844 ;
  assign n846 = ~n46 & n845 ;
  assign n847 = n643 ^ n159 ^ 1'b0 ;
  assign n848 = ~n177 & n390 ;
  assign n849 = n141 | n848 ;
  assign n850 = ~n299 & n849 ;
  assign n851 = ( n24 & n47 ) | ( n24 & n154 ) | ( n47 & n154 ) ;
  assign n852 = n308 | n851 ;
  assign n853 = n850 | n852 ;
  assign n854 = ~n142 & n310 ;
  assign n855 = n94 & n854 ;
  assign n856 = n175 | n855 ;
  assign n857 = x1 & n30 ;
  assign n858 = n856 & ~n857 ;
  assign n859 = n278 & n858 ;
  assign n860 = ~n81 & n229 ;
  assign n861 = n310 & n860 ;
  assign n862 = n149 & ~n283 ;
  assign n867 = n604 ^ n215 ^ 1'b0 ;
  assign n865 = ( n40 & ~n220 ) | ( n40 & n842 ) | ( ~n220 & n842 ) ;
  assign n863 = ~n94 & n392 ;
  assign n864 = ~n139 & n863 ;
  assign n866 = n865 ^ n864 ^ 1'b0 ;
  assign n868 = n867 ^ n866 ^ 1'b0 ;
  assign n869 = n628 & n868 ;
  assign n870 = n843 ^ n258 ^ 1'b0 ;
  assign n871 = n498 ^ n417 ^ 1'b0 ;
  assign n872 = n356 & n871 ;
  assign n873 = n131 | n621 ;
  assign n874 = n872 & ~n873 ;
  assign n875 = n167 & n549 ;
  assign n876 = n875 ^ n767 ^ 1'b0 ;
  assign n877 = n653 ^ n534 ^ 1'b0 ;
  assign n878 = n342 & ~n877 ;
  assign n879 = n828 ^ n708 ^ 1'b0 ;
  assign n880 = n17 | n292 ;
  assign n881 = n410 | n880 ;
  assign n882 = n881 ^ n678 ^ 1'b0 ;
  assign n883 = n364 ^ n234 ^ 1'b0 ;
  assign n884 = ~n581 & n636 ;
  assign n885 = ~n221 & n227 ;
  assign n886 = ~n412 & n885 ;
  assign n887 = ~n330 & n434 ;
  assign n888 = n887 ^ n427 ^ 1'b0 ;
  assign n889 = n886 | n888 ;
  assign n890 = n884 & ~n889 ;
  assign n891 = n164 & n258 ;
  assign n892 = n618 & n891 ;
  assign n893 = n558 ^ n308 ^ 1'b0 ;
  assign n894 = ~n79 & n893 ;
  assign n895 = n372 ^ n352 ^ 1'b0 ;
  assign n896 = n895 ^ n844 ^ 1'b0 ;
  assign n897 = n388 & ~n403 ;
  assign n898 = ~n346 & n897 ;
  assign n899 = ~n243 & n898 ;
  assign n900 = n899 ^ n236 ^ 1'b0 ;
  assign n901 = n900 ^ n403 ^ 1'b0 ;
  assign n902 = n901 ^ n717 ^ 1'b0 ;
  assign n903 = n489 & n902 ;
  assign n904 = n903 ^ n493 ^ 1'b0 ;
  assign n905 = ~n512 & n629 ;
  assign n906 = n904 & ~n905 ;
  assign n907 = n608 ^ n352 ^ 1'b0 ;
  assign n908 = n567 ^ n73 ^ 1'b0 ;
  assign n909 = n184 & n384 ;
  assign n910 = ~n16 & n909 ;
  assign n911 = n114 & ~n769 ;
  assign n912 = n68 & n911 ;
  assign n913 = n354 & n587 ;
  assign n914 = n913 ^ n904 ^ 1'b0 ;
  assign n916 = ~n35 & n83 ;
  assign n917 = n916 ^ n72 ^ 1'b0 ;
  assign n918 = n625 ^ n122 ^ 1'b0 ;
  assign n919 = n917 | n918 ;
  assign n915 = n69 | n486 ;
  assign n920 = n919 ^ n915 ^ 1'b0 ;
  assign n921 = n364 & n920 ;
  assign n922 = n296 ^ n146 ^ 1'b0 ;
  assign n923 = ~n336 & n634 ;
  assign n924 = ~n922 & n923 ;
  assign n925 = n128 | n216 ;
  assign n926 = n925 ^ n300 ^ 1'b0 ;
  assign n927 = n675 & ~n926 ;
  assign n928 = n273 ^ n123 ^ 1'b0 ;
  assign n929 = ~x0 & n928 ;
  assign n931 = ~n500 & n690 ;
  assign n930 = n436 ^ n109 ^ 1'b0 ;
  assign n932 = n931 ^ n930 ^ 1'b0 ;
  assign n933 = n283 & ~n698 ;
  assign n934 = n933 ^ n512 ^ 1'b0 ;
  assign n935 = n678 ^ n599 ^ 1'b0 ;
  assign n936 = ~n102 & n438 ;
  assign n937 = ~n55 & n936 ;
  assign n938 = n457 ^ n55 ^ 1'b0 ;
  assign n939 = n938 ^ n185 ^ 1'b0 ;
  assign n940 = ~n937 & n939 ;
  assign n941 = n135 & ~n226 ;
  assign n942 = n941 ^ n205 ^ 1'b0 ;
  assign n943 = n942 ^ n860 ^ 1'b0 ;
  assign n944 = ~n479 & n943 ;
  assign n945 = ~n208 & n555 ;
  assign n946 = n627 ^ n255 ^ 1'b0 ;
  assign n947 = ~n374 & n946 ;
  assign n948 = n945 & n947 ;
  assign n949 = n948 ^ n244 ^ 1'b0 ;
  assign n950 = x9 & ~n378 ;
  assign n951 = n950 ^ n736 ^ 1'b0 ;
  assign n952 = ~n92 & n848 ;
  assign n953 = ~n381 & n952 ;
  assign n954 = n953 ^ n123 ^ 1'b0 ;
  assign n955 = n954 ^ n107 ^ 1'b0 ;
  assign n956 = n86 & ~n87 ;
  assign n957 = n743 & n848 ;
  assign n958 = n956 & n957 ;
  assign n959 = n754 ^ n146 ^ 1'b0 ;
  assign n960 = ~n310 & n959 ;
  assign n961 = ~n42 & n469 ;
  assign n962 = ~n220 & n697 ;
  assign n963 = n246 | n962 ;
  assign n964 = n957 ^ n614 ^ 1'b0 ;
  assign n965 = n475 ^ n159 ^ 1'b0 ;
  assign n966 = n965 ^ n734 ^ 1'b0 ;
  assign n967 = n381 | n698 ;
  assign n968 = n967 ^ n777 ^ 1'b0 ;
  assign n969 = n133 | n665 ;
  assign n970 = n969 ^ n361 ^ 1'b0 ;
  assign n971 = n968 & ~n970 ;
  assign n972 = n971 ^ n679 ^ 1'b0 ;
  assign n973 = n699 & n972 ;
  assign n974 = n170 & n853 ;
  assign n975 = n791 ^ n684 ^ 1'b0 ;
  assign n976 = n330 & ~n493 ;
  assign n977 = n503 & n976 ;
  assign n978 = n86 | n904 ;
  assign n979 = n81 | n978 ;
  assign n980 = ~n55 & n979 ;
  assign n981 = n161 & n709 ;
  assign n982 = n352 & n981 ;
  assign n983 = n681 | n982 ;
  assign n984 = n55 & n215 ;
  assign n985 = n244 ^ n142 ^ 1'b0 ;
  assign n986 = n84 & ~n985 ;
  assign n987 = ~n168 & n205 ;
  assign n988 = n390 | n987 ;
  assign n989 = n52 & ~n206 ;
  assign n990 = n236 | n989 ;
  assign n991 = n990 ^ n412 ^ 1'b0 ;
  assign n992 = n991 ^ n602 ^ 1'b0 ;
  assign n993 = n334 & n992 ;
  assign n995 = x1 & ~n168 ;
  assign n994 = ~n576 & n765 ;
  assign n996 = n995 ^ n994 ^ 1'b0 ;
  assign n997 = n850 & n996 ;
  assign n998 = n400 & ~n997 ;
  assign n999 = n761 ^ n117 ^ 1'b0 ;
  assign n1000 = n44 & ~n999 ;
  assign n1001 = n869 ^ n403 ^ n286 ;
  assign n1002 = n549 ^ n238 ^ 1'b0 ;
  assign n1003 = n607 ^ n452 ^ 1'b0 ;
  assign n1004 = n269 & n417 ;
  assign n1005 = n508 | n1004 ;
  assign n1007 = n257 ^ n151 ^ 1'b0 ;
  assign n1006 = x3 & n203 ;
  assign n1008 = n1007 ^ n1006 ^ 1'b0 ;
  assign n1009 = n792 ^ x0 ^ 1'b0 ;
  assign n1010 = n903 & ~n1009 ;
  assign n1011 = ( n294 & ~n295 ) | ( n294 & n857 ) | ( ~n295 & n857 ) ;
  assign n1012 = n599 | n1011 ;
  assign n1013 = n1010 | n1012 ;
  assign n1014 = ~n434 & n751 ;
  assign n1015 = ~n269 & n1014 ;
  assign n1016 = n841 ^ n715 ^ 1'b0 ;
  assign n1018 = n87 & ~n611 ;
  assign n1019 = n1018 ^ n56 ^ 1'b0 ;
  assign n1017 = ~n281 & n1010 ;
  assign n1020 = n1019 ^ n1017 ^ 1'b0 ;
  assign n1021 = n670 & ~n958 ;
  assign n1022 = n1021 ^ n139 ^ 1'b0 ;
  assign n1023 = n255 & ~n640 ;
  assign n1024 = n1023 ^ n384 ^ 1'b0 ;
  assign n1025 = n748 ^ n286 ^ 1'b0 ;
  assign n1026 = n181 ^ n55 ^ 1'b0 ;
  assign n1027 = n1026 ^ n339 ^ 1'b0 ;
  assign n1028 = n269 & n581 ;
  assign n1029 = n1027 & n1028 ;
  assign n1030 = n482 & ~n1029 ;
  assign n1031 = n1030 ^ n1023 ^ 1'b0 ;
  assign n1032 = n68 | n588 ;
  assign n1033 = n1032 ^ n258 ^ 1'b0 ;
  assign n1034 = n1033 ^ n491 ^ 1'b0 ;
  assign n1035 = n83 & ~n94 ;
  assign n1036 = n55 & n1035 ;
  assign n1037 = n251 & ~n553 ;
  assign n1038 = ~n751 & n1037 ;
  assign n1039 = n184 | n1038 ;
  assign n1040 = n849 ^ n281 ^ 1'b0 ;
  assign n1041 = n1040 ^ n912 ^ n342 ;
  assign n1042 = ~n316 & n564 ;
  assign n1043 = n708 & n1042 ;
  assign n1044 = n233 & ~n628 ;
  assign n1045 = n717 ^ n273 ^ 1'b0 ;
  assign n1046 = ~n1044 & n1045 ;
  assign n1047 = n1046 ^ n389 ^ 1'b0 ;
  assign n1048 = n161 & n732 ;
  assign n1049 = n875 ^ n806 ^ 1'b0 ;
  assign n1050 = n205 & ~n279 ;
  assign n1051 = ~n274 & n662 ;
  assign n1052 = n604 ^ n133 ^ 1'b0 ;
  assign n1053 = n80 | n542 ;
  assign n1054 = x0 & ~n130 ;
  assign n1055 = x4 & n1013 ;
  assign n1056 = n1055 ^ n111 ^ 1'b0 ;
  assign n1057 = n233 ^ n83 ^ 1'b0 ;
  assign n1058 = n55 & n1057 ;
  assign n1059 = ( ~n123 & n564 ) | ( ~n123 & n688 ) | ( n564 & n688 ) ;
  assign n1062 = n205 ^ n116 ^ 1'b0 ;
  assign n1063 = n476 & ~n1062 ;
  assign n1061 = ~n587 & n642 ;
  assign n1064 = n1063 ^ n1061 ^ 1'b0 ;
  assign n1060 = n278 ^ n238 ^ 1'b0 ;
  assign n1065 = n1064 ^ n1060 ^ 1'b0 ;
  assign n1066 = n459 & ~n1065 ;
  assign n1067 = n336 | n769 ;
  assign n1068 = n952 ^ n423 ^ 1'b0 ;
  assign n1069 = ~n958 & n1068 ;
  assign n1070 = ~n250 & n337 ;
  assign n1071 = n1070 ^ n704 ^ 1'b0 ;
  assign n1072 = ~n989 & n1071 ;
  assign n1073 = n685 ^ n325 ^ 1'b0 ;
  assign n1074 = n1073 ^ n239 ^ 1'b0 ;
  assign n1075 = n1072 & ~n1074 ;
  assign n1076 = n553 & n823 ;
  assign n1077 = ~n1075 & n1076 ;
  assign n1078 = ~n690 & n853 ;
  assign n1079 = ~n135 & n1040 ;
  assign n1080 = n120 ^ n50 ^ 1'b0 ;
  assign n1081 = n939 & n1080 ;
  assign n1082 = n215 & ~n799 ;
  assign n1083 = n1081 & ~n1082 ;
  assign n1084 = n993 ^ n653 ^ 1'b0 ;
  assign n1085 = n279 & n1084 ;
  assign n1086 = n1085 ^ n1047 ^ 1'b0 ;
  assign n1087 = n234 ^ n185 ^ 1'b0 ;
  assign n1088 = n1087 ^ n286 ^ 1'b0 ;
  assign n1089 = ~n530 & n811 ;
  assign n1094 = n184 ^ n94 ^ 1'b0 ;
  assign n1095 = n886 | n1094 ;
  assign n1090 = ( n16 & n68 ) | ( n16 & n350 ) | ( n68 & n350 ) ;
  assign n1091 = n512 & n1090 ;
  assign n1092 = ~n231 & n1091 ;
  assign n1093 = n1092 ^ n367 ^ 1'b0 ;
  assign n1096 = n1095 ^ n1093 ^ 1'b0 ;
  assign n1097 = n487 ^ n315 ^ 1'b0 ;
  assign n1098 = n34 & ~n713 ;
  assign n1102 = n79 | n107 ;
  assign n1099 = n758 ^ n607 ^ 1'b0 ;
  assign n1100 = x2 & ~n1099 ;
  assign n1101 = n527 & n1100 ;
  assign n1103 = n1102 ^ n1101 ^ 1'b0 ;
  assign n1104 = n206 ^ n114 ^ 1'b0 ;
  assign n1105 = n1104 ^ n182 ^ 1'b0 ;
  assign n1106 = n662 & ~n1105 ;
  assign n1107 = ~n612 & n659 ;
  assign n1108 = n1107 ^ n300 ^ 1'b0 ;
  assign n1109 = n1108 ^ n393 ^ 1'b0 ;
  assign n1110 = n878 ^ n139 ^ 1'b0 ;
  assign n1111 = n215 | n296 ;
  assign n1112 = n1111 ^ n273 ^ 1'b0 ;
  assign n1113 = ~n530 & n928 ;
  assign n1114 = n641 & ~n907 ;
  assign n1115 = n1114 ^ n102 ^ 1'b0 ;
  assign n1116 = ~n131 & n653 ;
  assign n1117 = ~n233 & n1116 ;
  assign n1118 = n787 ^ n294 ^ 1'b0 ;
  assign n1119 = ~n34 & n461 ;
  assign n1120 = n849 ^ n253 ^ 1'b0 ;
  assign n1121 = ~n694 & n1120 ;
  assign n1123 = n271 ^ n82 ^ 1'b0 ;
  assign n1124 = n111 & n1123 ;
  assign n1122 = n133 | n675 ;
  assign n1125 = n1124 ^ n1122 ^ 1'b0 ;
  assign n1126 = n457 & n1125 ;
  assign n1127 = n1126 ^ n142 ^ 1'b0 ;
  assign n1128 = ~n632 & n1127 ;
  assign n1129 = n1128 ^ n479 ^ 1'b0 ;
  assign n1130 = n694 ^ n200 ^ 1'b0 ;
  assign n1131 = n359 & ~n964 ;
  assign n1132 = ~n1057 & n1131 ;
  assign n1133 = n346 & ~n570 ;
  assign n1134 = n1133 ^ n208 ^ 1'b0 ;
  assign n1137 = n125 & ~n846 ;
  assign n1135 = n483 ^ n478 ^ 1'b0 ;
  assign n1136 = n590 | n1135 ;
  assign n1138 = n1137 ^ n1136 ^ 1'b0 ;
  assign n1139 = ~n87 & n185 ;
  assign n1140 = n292 & ~n859 ;
  assign n1141 = n191 | n1140 ;
  assign n1142 = n690 ^ n69 ^ 1'b0 ;
  assign n1143 = n1142 ^ n712 ^ 1'b0 ;
  assign n1144 = ~n23 & n643 ;
  assign n1145 = n400 ^ n330 ^ 1'b0 ;
  assign n1146 = n265 & n1145 ;
  assign n1147 = ~n274 & n1146 ;
  assign n1148 = n1147 ^ n466 ^ 1'b0 ;
  assign n1149 = n879 ^ n859 ^ n79 ;
  assign n1150 = n670 & n1149 ;
  assign n1151 = n1150 ^ n982 ^ 1'b0 ;
  assign n1152 = n1081 ^ n952 ^ 1'b0 ;
  assign n1153 = n450 & n501 ;
  assign n1154 = n307 & n1153 ;
  assign n1155 = n1154 ^ n295 ^ 1'b0 ;
  assign n1156 = ~n820 & n1155 ;
  assign n1157 = n1156 ^ n191 ^ 1'b0 ;
  assign n1158 = n107 ^ n55 ^ 1'b0 ;
  assign n1159 = n636 & n840 ;
  assign n1160 = n1159 ^ n701 ^ 1'b0 ;
  assign n1161 = n1158 & n1160 ;
  assign n1162 = n1104 ^ n584 ^ 1'b0 ;
  assign n1163 = n443 ^ n436 ^ 1'b0 ;
  assign n1164 = n427 & ~n670 ;
  assign n1165 = n246 ^ n105 ^ 1'b0 ;
  assign n1166 = ~n169 & n1165 ;
  assign n1167 = n32 ^ x10 ^ 1'b0 ;
  assign n1168 = n194 ^ n52 ^ 1'b0 ;
  assign n1169 = n161 & n1168 ;
  assign n1170 = n1167 & n1169 ;
  assign n1171 = n321 ^ n58 ^ 1'b0 ;
  assign n1172 = n257 & n1171 ;
  assign n1173 = ~n55 & n72 ;
  assign n1174 = n79 | n169 ;
  assign n1175 = n122 & ~n241 ;
  assign n1176 = ~n1174 & n1175 ;
  assign n1177 = ~n1173 & n1176 ;
  assign n1178 = n1172 & n1177 ;
  assign n1179 = n1178 ^ n280 ^ 1'b0 ;
  assign n1180 = ~n75 & n364 ;
  assign n1181 = n1180 ^ n931 ^ 1'b0 ;
  assign n1182 = n35 | n1181 ;
  assign n1183 = n1182 ^ n404 ^ 1'b0 ;
  assign n1184 = ( ~n244 & n643 ) | ( ~n244 & n646 ) | ( n643 & n646 ) ;
  assign n1185 = n177 ^ n113 ^ 1'b0 ;
  assign n1190 = n381 | n440 ;
  assign n1191 = n1190 ^ n62 ^ 1'b0 ;
  assign n1186 = n1168 ^ n292 ^ 1'b0 ;
  assign n1187 = n172 & ~n793 ;
  assign n1188 = ~n1186 & n1187 ;
  assign n1189 = n527 & ~n1188 ;
  assign n1192 = n1191 ^ n1189 ^ 1'b0 ;
  assign n1193 = n357 | n626 ;
  assign n1194 = ~n77 & n253 ;
  assign n1195 = n363 & n392 ;
  assign n1196 = n738 ^ x1 ^ 1'b0 ;
  assign n1197 = n1195 | n1196 ;
  assign n1198 = n43 & n777 ;
  assign n1199 = ~n474 & n1198 ;
  assign n1200 = ~n1103 & n1199 ;
  assign n1201 = ~n540 & n1200 ;
  assign n1202 = x2 & ~n35 ;
  assign n1204 = x5 & n194 ;
  assign n1205 = n79 & n1204 ;
  assign n1203 = n333 | n340 ;
  assign n1206 = n1205 ^ n1203 ^ 1'b0 ;
  assign n1207 = n1172 ^ n566 ^ 1'b0 ;
  assign n1208 = n210 | n1207 ;
  assign n1209 = n518 & n694 ;
  assign n1210 = ~n313 & n592 ;
  assign n1211 = ~n501 & n709 ;
  assign n1212 = ~n671 & n1211 ;
  assign n1213 = n435 & ~n662 ;
  assign n1214 = n971 ^ n781 ^ 1'b0 ;
  assign n1215 = ~x0 & n486 ;
  assign n1216 = n1215 ^ n745 ^ 1'b0 ;
  assign n1217 = n1216 ^ n643 ^ 1'b0 ;
  assign n1218 = n993 & ~n1217 ;
  assign n1219 = n432 & n756 ;
  assign n1220 = n1219 ^ n47 ^ 1'b0 ;
  assign n1221 = ~n236 & n1175 ;
  assign n1222 = n1221 ^ n857 ^ 1'b0 ;
  assign n1223 = n141 | n907 ;
  assign n1224 = n927 & ~n1154 ;
  assign n1225 = n423 ^ n274 ^ 1'b0 ;
  assign n1226 = n1225 ^ n323 ^ 1'b0 ;
  assign n1227 = n507 ^ n165 ^ 1'b0 ;
  assign n1228 = n1227 ^ n939 ^ 1'b0 ;
  assign n1229 = n241 | n1228 ;
  assign n1230 = n508 | n1102 ;
  assign n1231 = n619 ^ n446 ^ 1'b0 ;
  assign n1232 = n55 & ~n705 ;
  assign n1233 = n200 | n1169 ;
  assign n1234 = n47 | n1233 ;
  assign n1235 = n83 & n86 ;
  assign n1236 = n596 & ~n1235 ;
  assign n1237 = n1142 ^ n277 ^ 1'b0 ;
  assign n1238 = n1236 & n1237 ;
  assign n1239 = ~n1234 & n1238 ;
  assign n1240 = n226 & n388 ;
  assign n1241 = n1240 ^ n677 ^ 1'b0 ;
  assign n1242 = n94 ^ n43 ^ 1'b0 ;
  assign n1243 = n1241 & ~n1242 ;
  assign n1244 = n1243 ^ n390 ^ 1'b0 ;
  assign n1245 = n290 | n1244 ;
  assign n1246 = n1245 ^ x8 ^ 1'b0 ;
  assign n1247 = n302 ^ n218 ^ 1'b0 ;
  assign n1248 = n659 & n1247 ;
  assign n1249 = ( n659 & n986 ) | ( n659 & ~n1248 ) | ( n986 & ~n1248 ) ;
  assign n1250 = n643 ^ n328 ^ 1'b0 ;
  assign n1256 = n122 | n1064 ;
  assign n1253 = n297 & n309 ;
  assign n1254 = n1253 ^ n573 ^ 1'b0 ;
  assign n1251 = n164 & ~n1235 ;
  assign n1252 = n1251 ^ n400 ^ 1'b0 ;
  assign n1255 = n1254 ^ n1252 ^ n417 ;
  assign n1257 = n1256 ^ n1255 ^ n477 ;
  assign n1258 = n540 & ~n788 ;
  assign n1259 = ~n472 & n477 ;
  assign n1260 = n1258 & n1259 ;
  assign n1261 = n318 | n891 ;
  assign n1262 = n1048 & ~n1261 ;
  assign n1263 = n304 & n1100 ;
  assign n1264 = n1263 ^ x0 ^ 1'b0 ;
  assign n1265 = n738 & ~n989 ;
  assign n1266 = n900 & n1265 ;
  assign n1267 = n1013 | n1266 ;
  assign n1268 = n153 & ~n581 ;
  assign n1269 = n56 & ~n847 ;
  assign n1270 = ~n562 & n1269 ;
  assign n1271 = n722 ^ n641 ^ 1'b0 ;
  assign n1272 = n183 & n1271 ;
  assign n1273 = n1272 ^ n158 ^ 1'b0 ;
  assign n1274 = n374 & n1273 ;
  assign n1275 = n462 ^ n255 ^ 1'b0 ;
  assign n1276 = ~n1274 & n1275 ;
  assign n1277 = n1067 | n1080 ;
  assign n1278 = n665 ^ n181 ^ 1'b0 ;
  assign n1279 = n1278 ^ n613 ^ 1'b0 ;
  assign n1280 = ~n390 & n1279 ;
  assign n1281 = ~n23 & n52 ;
  assign n1282 = n1281 ^ n188 ^ 1'b0 ;
  assign n1283 = ~n546 & n1282 ;
  assign n1284 = n1280 & ~n1283 ;
  assign n1285 = n390 | n816 ;
  assign n1286 = ~n694 & n732 ;
  assign n1287 = n55 & n1286 ;
  assign n1288 = n113 & ~n393 ;
  assign n1289 = ~n566 & n1288 ;
  assign n1290 = n226 & n1214 ;
  assign n1291 = n1290 ^ n23 ^ 1'b0 ;
  assign n1292 = n1008 ^ n654 ^ 1'b0 ;
  assign n1293 = n412 ^ n216 ^ n168 ;
  assign n1294 = n185 & n309 ;
  assign n1295 = ~n1293 & n1294 ;
  assign n1296 = n613 ^ n475 ^ 1'b0 ;
  assign n1297 = n1295 | n1296 ;
  assign n1298 = n1280 ^ n357 ^ 1'b0 ;
  assign n1299 = n169 | n1154 ;
  assign n1300 = n1299 ^ n419 ^ 1'b0 ;
  assign n1301 = n1300 ^ n456 ^ 1'b0 ;
  assign n1302 = ~n228 & n1301 ;
  assign n1303 = n37 & n1295 ;
  assign n1304 = n86 & ~n137 ;
  assign n1305 = n475 | n1304 ;
  assign n1306 = n1305 ^ n621 ^ 1'b0 ;
  assign n1307 = n1306 ^ n849 ^ 1'b0 ;
  assign n1308 = n1132 ^ n75 ^ 1'b0 ;
  assign n1309 = n343 & n535 ;
  assign n1315 = n190 | n397 ;
  assign n1316 = n1093 & ~n1315 ;
  assign n1313 = ~n389 & n596 ;
  assign n1310 = n1283 ^ n654 ^ 1'b0 ;
  assign n1311 = n1144 ^ n117 ^ 1'b0 ;
  assign n1312 = n1310 & n1311 ;
  assign n1314 = n1313 ^ n1312 ^ 1'b0 ;
  assign n1317 = n1316 ^ n1314 ^ 1'b0 ;
  assign n1318 = n1309 | n1317 ;
  assign n1319 = ~n86 & n830 ;
  assign n1320 = n133 & n1319 ;
  assign n1321 = n121 & ~n1320 ;
  assign n1322 = n988 & n1321 ;
  assign n1324 = n1075 ^ n657 ^ 1'b0 ;
  assign n1323 = n354 ^ n276 ^ 1'b0 ;
  assign n1325 = n1324 ^ n1323 ^ 1'b0 ;
  assign n1326 = n252 ^ n153 ^ 1'b0 ;
  assign n1327 = n287 & ~n917 ;
  assign n1328 = n221 & n1327 ;
  assign n1329 = n1328 ^ n311 ^ 1'b0 ;
  assign n1330 = n32 | n903 ;
  assign n1331 = n547 | n1330 ;
  assign n1332 = n630 & ~n1085 ;
  assign n1333 = ~n85 & n208 ;
  assign n1334 = n1333 ^ n1170 ^ 1'b0 ;
  assign n1335 = n1004 & n1155 ;
  assign n1336 = n133 | n1295 ;
  assign n1337 = n86 & ~n1336 ;
  assign n1338 = n945 & ~n1070 ;
  assign n1339 = ~n513 & n1338 ;
  assign n1340 = n1339 ^ n404 ^ 1'b0 ;
  assign n1341 = n984 & n1340 ;
  assign n1342 = n169 & ~n724 ;
  assign n1343 = n43 | n68 ;
  assign n1344 = n1343 ^ n460 ^ 1'b0 ;
  assign n1345 = ~n1342 & n1344 ;
  assign n1346 = n330 ^ n116 ^ 1'b0 ;
  assign n1347 = n328 | n1058 ;
  assign n1348 = n856 ^ x0 ^ 1'b0 ;
  assign n1349 = n1007 | n1348 ;
  assign n1350 = n1077 ^ n556 ^ 1'b0 ;
  assign n1351 = n576 | n924 ;
  assign n1352 = n180 & ~n1351 ;
  assign n1353 = n1352 ^ n861 ^ 1'b0 ;
  assign n1354 = n1350 & ~n1353 ;
  assign n1355 = n1304 ^ n390 ^ 1'b0 ;
  assign n1356 = x0 & ~n702 ;
  assign n1357 = ~n1355 & n1356 ;
  assign n1358 = n582 ^ n196 ^ 1'b0 ;
  assign n1359 = n1315 | n1358 ;
  assign n1360 = n125 & n810 ;
  assign n1366 = n1184 ^ n980 ^ 1'b0 ;
  assign n1361 = ~n310 & n777 ;
  assign n1362 = n208 | n1361 ;
  assign n1363 = n481 ^ n461 ^ 1'b0 ;
  assign n1364 = n1181 & n1363 ;
  assign n1365 = n1362 & n1364 ;
  assign n1367 = n1366 ^ n1365 ^ 1'b0 ;
  assign n1368 = n279 & ~n698 ;
  assign n1369 = n851 ^ n83 ^ 1'b0 ;
  assign n1370 = n1369 ^ n1052 ^ 1'b0 ;
  assign n1371 = n426 ^ n365 ^ 1'b0 ;
  assign n1372 = n182 & n1371 ;
  assign n1373 = ~n898 & n1372 ;
  assign n1374 = ~n1056 & n1373 ;
  assign n1375 = n1374 ^ n1086 ^ 1'b0 ;
  assign n1376 = n1375 ^ n123 ^ 1'b0 ;
  assign n1377 = n1241 & n1376 ;
  assign n1378 = ~n17 & n977 ;
  assign n1379 = n1378 ^ n1368 ^ 1'b0 ;
  assign n1381 = n352 | n694 ;
  assign n1380 = n269 & n400 ;
  assign n1382 = n1381 ^ n1380 ^ n81 ;
  assign n1383 = n835 ^ n528 ^ 1'b0 ;
  assign n1384 = ~n1382 & n1383 ;
  assign n1385 = n775 & ~n926 ;
  assign n1386 = ~n68 & n1070 ;
  assign n1387 = n1386 ^ n812 ^ n291 ;
  assign n1388 = ~n608 & n1387 ;
  assign n1389 = n421 & n723 ;
  assign n1390 = ~n794 & n1389 ;
  assign n1391 = ~n23 & n238 ;
  assign n1392 = ~n1390 & n1391 ;
  assign n1393 = n288 ^ n284 ^ 1'b0 ;
  assign n1394 = n21 & n1393 ;
  assign n1395 = n1394 ^ n652 ^ 1'b0 ;
  assign n1396 = n299 & ~n1395 ;
  assign n1397 = ~n117 & n233 ;
  assign n1398 = ~n1396 & n1397 ;
  assign n1399 = n1143 | n1398 ;
  assign n1400 = n753 | n1399 ;
  assign n1401 = n989 & ~n1400 ;
  assign n1402 = n653 ^ n448 ^ 1'b0 ;
  assign n1403 = n323 & n1402 ;
  assign n1404 = x1 & n513 ;
  assign n1405 = n1404 ^ n417 ^ 1'b0 ;
  assign n1406 = n1403 & ~n1405 ;
  assign n1407 = ~n129 & n346 ;
  assign n1408 = n390 ^ n238 ^ 1'b0 ;
  assign n1409 = n250 & ~n1408 ;
  assign n1410 = ~n1407 & n1409 ;
  assign n1411 = n25 & ~n479 ;
  assign n1412 = n161 & n636 ;
  assign n1413 = n1118 ^ n113 ^ 1'b0 ;
  assign n1414 = n1412 & ~n1413 ;
  assign n1415 = n955 ^ n75 ^ 1'b0 ;
  assign n1416 = n1415 ^ n381 ^ 1'b0 ;
  assign n1417 = n23 & n337 ;
  assign n1418 = n553 | n1417 ;
  assign n1419 = n221 | n809 ;
  assign n1420 = ~n86 & n1419 ;
  assign n1421 = n1420 ^ n292 ^ 1'b0 ;
  assign n1422 = n1421 ^ n800 ^ 1'b0 ;
  assign n1423 = n465 | n1422 ;
  assign n1424 = n640 | n1423 ;
  assign n1425 = n901 | n1424 ;
  assign n1426 = n766 ^ n226 ^ 1'b0 ;
  assign n1427 = n1425 & n1426 ;
  assign n1428 = ~n468 & n1427 ;
  assign n1429 = n939 ^ n25 ^ 1'b0 ;
  assign n1430 = n215 ^ n123 ^ 1'b0 ;
  assign n1431 = n1407 & ~n1430 ;
  assign n1432 = n867 ^ n406 ^ 1'b0 ;
  assign n1433 = n15 & n310 ;
  assign n1434 = n1433 ^ n1154 ^ 1'b0 ;
  assign n1435 = ~n1432 & n1434 ;
  assign n1436 = ~n690 & n1435 ;
  assign n1437 = ~n51 & n1436 ;
  assign n1438 = n645 | n917 ;
  assign n1439 = n178 | n690 ;
  assign n1440 = n338 | n758 ;
  assign n1441 = n777 & ~n986 ;
  assign n1442 = n227 & n1441 ;
  assign n1443 = n927 & n1442 ;
  assign n1444 = ~n876 & n1443 ;
  assign n1445 = ~n144 & n1444 ;
  assign n1446 = n55 & ~n995 ;
  assign n1447 = n1446 ^ n1002 ^ 1'b0 ;
  assign n1448 = n182 | n771 ;
  assign n1449 = n1448 ^ n1165 ^ 1'b0 ;
  assign n1450 = n1449 ^ n816 ^ 1'b0 ;
  assign n1451 = ~n255 & n398 ;
  assign n1452 = ~n827 & n1451 ;
  assign n1453 = ~n837 & n1452 ;
  assign n1454 = n956 | n1440 ;
  assign n1455 = n1453 | n1454 ;
  assign n1456 = x4 & ~n281 ;
  assign n1457 = n852 ^ n206 ^ 1'b0 ;
  assign n1458 = n356 & n1457 ;
  assign n1459 = n1458 ^ n929 ^ 1'b0 ;
  assign n1460 = ~n1456 & n1459 ;
  assign n1461 = ~n1309 & n1460 ;
  assign n1462 = ~n288 & n1461 ;
  assign n1463 = n976 ^ n582 ^ n461 ;
  assign n1464 = n139 | n867 ;
  assign n1465 = n1084 ^ n144 ^ 1'b0 ;
  assign n1469 = n647 & ~n1010 ;
  assign n1470 = ~n1152 & n1469 ;
  assign n1466 = n313 ^ n23 ^ 1'b0 ;
  assign n1467 = n1466 ^ n585 ^ 1'b0 ;
  assign n1468 = ~n632 & n1467 ;
  assign n1471 = n1470 ^ n1468 ^ 1'b0 ;
  assign n1472 = n1471 ^ n614 ^ 1'b0 ;
  assign n1473 = n565 ^ n55 ^ 1'b0 ;
  assign n1474 = n1419 | n1473 ;
  assign n1475 = n1177 | n1474 ;
  assign n1476 = n1106 ^ n283 ^ 1'b0 ;
  assign n1477 = n1476 ^ n779 ^ 1'b0 ;
  assign n1478 = n787 & n886 ;
  assign n1479 = n510 ^ n169 ^ 1'b0 ;
  assign n1480 = n1479 ^ n1174 ^ 1'b0 ;
  assign n1481 = n440 ^ n44 ^ 1'b0 ;
  assign n1482 = n726 & ~n1481 ;
  assign n1483 = n1482 ^ n412 ^ 1'b0 ;
  assign n1484 = n1483 ^ n135 ^ 1'b0 ;
  assign n1485 = n114 & ~n382 ;
  assign n1486 = n1485 ^ n159 ^ 1'b0 ;
  assign n1487 = ~n1314 & n1486 ;
  assign n1488 = n512 ^ n48 ^ 1'b0 ;
  assign n1489 = n381 | n1488 ;
  assign n1490 = n294 & ~n1489 ;
  assign n1491 = n492 | n1490 ;
  assign n1492 = n1086 & ~n1491 ;
  assign n1493 = n75 | n1161 ;
  assign n1494 = n327 ^ x1 ^ 1'b0 ;
  assign n1495 = n292 & n1494 ;
  assign n1496 = n1495 ^ n585 ^ 1'b0 ;
  assign n1497 = n863 ^ n709 ^ n636 ;
  assign n1498 = n671 ^ n609 ^ 1'b0 ;
  assign n1499 = n191 & ~n989 ;
  assign n1500 = n734 ^ n596 ^ 1'b0 ;
  assign n1501 = ~n1499 & n1500 ;
  assign n1502 = n1501 ^ n474 ^ 1'b0 ;
  assign n1503 = n1502 ^ n1188 ^ 1'b0 ;
  assign n1504 = n1498 & ~n1503 ;
  assign n1505 = n306 ^ n263 ^ 1'b0 ;
  assign n1506 = ~n243 & n438 ;
  assign n1507 = ~n866 & n1506 ;
  assign n1508 = ~n503 & n1507 ;
  assign n1509 = n129 ^ n79 ^ 1'b0 ;
  assign n1510 = n1509 ^ n849 ^ 1'b0 ;
  assign n1511 = n280 | n1510 ;
  assign n1512 = n950 & ~n1235 ;
  assign n1513 = n1001 & n1313 ;
  assign n1514 = n714 & ~n1163 ;
  assign n1515 = n866 & n1514 ;
  assign n1516 = n540 & n1443 ;
  assign n1517 = n257 | n1198 ;
  assign n1518 = n1112 | n1517 ;
  assign n1519 = ( n190 & n755 ) | ( n190 & n764 ) | ( n755 & n764 ) ;
  assign n1520 = n55 & ~n191 ;
  assign n1521 = n1520 ^ n1329 ^ 1'b0 ;
  assign n1522 = n1521 ^ n86 ^ 1'b0 ;
  assign n1523 = n1522 ^ n1181 ^ 1'b0 ;
  assign n1524 = n247 & n392 ;
  assign n1525 = n1524 ^ n799 ^ 1'b0 ;
  assign n1526 = n846 | n1525 ;
  assign n1527 = n471 ^ x3 ^ 1'b0 ;
  assign n1528 = x7 | n596 ;
  assign n1529 = n249 & ~n1528 ;
  assign n1530 = x6 & ~n83 ;
  assign n1533 = n1466 ^ n556 ^ 1'b0 ;
  assign n1534 = n178 & n851 ;
  assign n1535 = ~n1533 & n1534 ;
  assign n1531 = ~n278 & n297 ;
  assign n1532 = n40 & ~n1531 ;
  assign n1536 = n1535 ^ n1532 ^ 1'b0 ;
  assign n1537 = n254 & ~n1536 ;
  assign n1538 = n512 | n1163 ;
  assign n1539 = n741 ^ n55 ^ 1'b0 ;
  assign n1540 = ~n888 & n1467 ;
  assign n1541 = n1540 ^ n19 ^ 1'b0 ;
  assign n1542 = n719 & n1425 ;
  assign n1543 = n1077 & n1542 ;
  assign n1544 = n206 | n1543 ;
  assign n1545 = n547 & ~n1544 ;
  assign n1546 = n114 & ~n194 ;
  assign n1547 = n592 | n865 ;
  assign n1548 = ~n1546 & n1547 ;
  assign n1549 = n1548 ^ n549 ^ 1'b0 ;
  assign n1550 = n1549 ^ n719 ^ 1'b0 ;
  assign n1551 = n388 & ~n1087 ;
  assign n1552 = n1551 ^ n1358 ^ 1'b0 ;
  assign n1554 = n350 & n647 ;
  assign n1555 = n353 & n1554 ;
  assign n1556 = n1555 ^ n86 ^ 1'b0 ;
  assign n1557 = n111 & n1520 ;
  assign n1558 = n1556 & n1557 ;
  assign n1553 = n895 | n908 ;
  assign n1559 = n1558 ^ n1553 ^ 1'b0 ;
  assign n1560 = n1361 ^ n799 ^ 1'b0 ;
  assign n1565 = n683 ^ n169 ^ 1'b0 ;
  assign n1561 = n346 ^ n19 ^ 1'b0 ;
  assign n1562 = n17 | n1561 ;
  assign n1563 = n715 & ~n1562 ;
  assign n1564 = n1563 ^ n1098 ^ 1'b0 ;
  assign n1566 = n1565 ^ n1564 ^ 1'b0 ;
  assign n1567 = n82 & n158 ;
  assign n1568 = n354 | n440 ;
  assign n1569 = n323 & ~n1568 ;
  assign n1570 = n1569 ^ n628 ^ 1'b0 ;
  assign n1571 = n1567 | n1570 ;
  assign n1572 = n715 & ~n865 ;
  assign n1573 = ~n133 & n1572 ;
  assign n1574 = n204 & n694 ;
  assign n1575 = n1574 ^ n233 ^ 1'b0 ;
  assign n1576 = n1573 | n1575 ;
  assign n1577 = n339 | n1576 ;
  assign n1578 = n1577 ^ n896 ^ 1'b0 ;
  assign n1579 = ~n198 & n1578 ;
  assign n1580 = n327 & ~n539 ;
  assign n1581 = n1580 ^ n1146 ^ 1'b0 ;
  assign n1582 = ~n1022 & n1276 ;
  assign n1584 = n456 ^ n142 ^ 1'b0 ;
  assign n1583 = n195 & ~n1016 ;
  assign n1585 = n1584 ^ n1583 ^ 1'b0 ;
  assign n1586 = n777 ^ n177 ^ 1'b0 ;
  assign n1587 = x8 & ~n1586 ;
  assign n1588 = ~n1585 & n1587 ;
  assign n1589 = ~n372 & n1226 ;
  assign n1590 = n1589 ^ n1183 ^ 1'b0 ;
  assign n1591 = ~x0 & n1590 ;
  assign n1592 = ( ~n153 & n1072 ) | ( ~n153 & n1399 ) | ( n1072 & n1399 ) ;
  assign n1593 = n931 & ~n1592 ;
  assign n1594 = n492 | n499 ;
  assign n1595 = n859 & ~n1594 ;
  assign n1596 = n448 & ~n1095 ;
  assign n1597 = n1595 & n1596 ;
  assign n1598 = n292 ^ n55 ^ 1'b0 ;
  assign n1599 = ~n616 & n1598 ;
  assign n1600 = ( ~n90 & n556 ) | ( ~n90 & n1486 ) | ( n556 & n1486 ) ;
  assign n1601 = ( n76 & n1004 ) | ( n76 & n1600 ) | ( n1004 & n1600 ) ;
  assign n1602 = ~n1056 & n1601 ;
  assign n1603 = n1283 | n1508 ;
  assign n1604 = x3 | n1603 ;
  assign n1608 = n359 & ~n1453 ;
  assign n1605 = n1487 ^ n861 ^ 1'b0 ;
  assign n1606 = ~n832 & n1605 ;
  assign n1607 = n987 & n1606 ;
  assign n1609 = n1608 ^ n1607 ^ 1'b0 ;
  assign n1610 = n1342 ^ n86 ^ 1'b0 ;
  assign n1611 = ~n479 & n1610 ;
  assign n1612 = n1611 ^ n34 ^ 1'b0 ;
  assign n1613 = ~n390 & n1612 ;
  assign n1614 = n900 ^ n690 ^ 1'b0 ;
  assign n1615 = n1613 & n1614 ;
  assign n1616 = n185 & ~n1007 ;
  assign n1617 = ~n1271 & n1616 ;
  assign n1619 = ( n102 & n313 ) | ( n102 & n592 ) | ( n313 & n592 ) ;
  assign n1618 = n108 | n175 ;
  assign n1620 = n1619 ^ n1618 ^ 1'b0 ;
  assign n1621 = n566 | n1620 ;
  assign n1622 = n1617 & ~n1621 ;
  assign n1623 = n976 ^ n501 ^ 1'b0 ;
  assign n1624 = n495 & n1623 ;
  assign n1625 = n753 ^ n185 ^ 1'b0 ;
  assign n1626 = n111 & ~n1625 ;
  assign n1627 = ~n86 & n365 ;
  assign n1628 = n37 & n323 ;
  assign n1629 = n391 & n1628 ;
  assign n1630 = n1519 ^ n697 ^ 1'b0 ;
  assign n1631 = n1185 ^ n701 ^ 1'b0 ;
  assign n1632 = n43 | n1325 ;
  assign n1633 = ( ~n257 & n788 ) | ( ~n257 & n878 ) | ( n788 & n878 ) ;
  assign n1634 = n257 & ~n1633 ;
  assign n1635 = n884 | n1066 ;
  assign n1636 = n164 & ~n432 ;
  assign n1637 = ~n775 & n1636 ;
  assign n1638 = ~n643 & n1637 ;
  assign n1639 = n1023 ^ n472 ^ 1'b0 ;
  assign n1640 = ~n1289 & n1639 ;
  assign n1641 = n459 | n934 ;
  assign n1642 = n178 | n1641 ;
  assign n1643 = n607 ^ n74 ^ 1'b0 ;
  assign n1644 = n1125 & ~n1643 ;
  assign n1645 = n1627 & ~n1644 ;
  assign n1647 = n419 & ~n802 ;
  assign n1648 = n782 & n1647 ;
  assign n1646 = ~n94 & n384 ;
  assign n1649 = n1648 ^ n1646 ^ 1'b0 ;
  assign n1650 = n318 | n1547 ;
  assign n1652 = ~n116 & n330 ;
  assign n1653 = n55 & ~n1652 ;
  assign n1651 = n378 & ~n1433 ;
  assign n1654 = n1653 ^ n1651 ^ 1'b0 ;
  assign n1655 = n673 & ~n1654 ;
  assign n1656 = n1526 | n1606 ;
  assign n1657 = n1178 ^ n613 ^ 1'b0 ;
  assign n1658 = n527 & n1657 ;
  assign n1659 = n107 & n458 ;
  assign n1660 = n1659 ^ n259 ^ 1'b0 ;
  assign n1662 = n654 ^ n226 ^ n208 ;
  assign n1661 = n178 & ~n274 ;
  assign n1663 = n1662 ^ n1661 ^ 1'b0 ;
  assign n1664 = n1433 & ~n1663 ;
  assign n1665 = n1075 ^ n666 ^ 1'b0 ;
  assign n1666 = n865 & n1665 ;
  assign n1667 = n16 & ~n1584 ;
  assign n1668 = n1667 ^ n833 ^ 1'b0 ;
  assign n1669 = ~n782 & n1668 ;
  assign n1670 = ~n280 & n596 ;
  assign n1671 = n1670 ^ n328 ^ 1'b0 ;
  assign n1672 = n348 & n1044 ;
  assign n1673 = n637 ^ n513 ^ 1'b0 ;
  assign n1674 = n1673 ^ n216 ^ 1'b0 ;
  assign n1675 = n1674 ^ n1194 ^ 1'b0 ;
  assign n1676 = n1672 | n1675 ;
  assign n1677 = ~n119 & n789 ;
  assign n1678 = n79 | n737 ;
  assign n1679 = n1677 | n1678 ;
  assign n1680 = n1679 ^ n1081 ^ 1'b0 ;
  assign n1681 = n229 & n1680 ;
  assign n1682 = n626 ^ n235 ^ 1'b0 ;
  assign n1683 = n539 | n1682 ;
  assign n1684 = n768 ^ n158 ^ 1'b0 ;
  assign n1685 = n541 & n1684 ;
  assign n1686 = n1685 ^ n1093 ^ 1'b0 ;
  assign n1687 = n1686 ^ n75 ^ 1'b0 ;
  assign n1688 = n671 & ~n1124 ;
  assign n1690 = n279 & n387 ;
  assign n1689 = n279 | n456 ;
  assign n1691 = n1690 ^ n1689 ^ 1'b0 ;
  assign n1692 = n1588 & ~n1602 ;
  assign n1693 = n629 ^ n158 ^ 1'b0 ;
  assign n1694 = n799 & ~n940 ;
  assign n1695 = n1694 ^ n811 ^ 1'b0 ;
  assign n1696 = ~n292 & n865 ;
  assign n1697 = n1696 ^ n932 ^ 1'b0 ;
  assign n1698 = n427 ^ x10 ^ 1'b0 ;
  assign n1699 = n908 & n1698 ;
  assign n1700 = n292 | n1052 ;
  assign n1701 = n288 | n1700 ;
  assign n1702 = n178 & n1203 ;
  assign n1703 = n513 & n883 ;
  assign n1704 = n1703 ^ n919 ^ 1'b0 ;
  assign n1705 = n354 & ~n1704 ;
  assign n1706 = x0 & n883 ;
  assign n1707 = n1706 ^ x3 ^ 1'b0 ;
  assign n1708 = n402 & ~n1707 ;
  assign n1709 = n847 ^ n457 ^ 1'b0 ;
  assign n1710 = n749 | n788 ;
  assign n1711 = n1600 ^ n1049 ^ 1'b0 ;
  assign n1712 = n770 & ~n950 ;
  assign n1713 = n580 & ~n703 ;
  assign n1714 = n921 | n956 ;
  assign n1715 = n1714 ^ x9 ^ 1'b0 ;
  assign n1718 = n253 ^ n101 ^ 1'b0 ;
  assign n1716 = n182 & ~n249 ;
  assign n1717 = ~n1260 & n1716 ;
  assign n1719 = n1718 ^ n1717 ^ 1'b0 ;
  assign n1720 = n1027 | n1719 ;
  assign n1721 = n1254 ^ x2 ^ 1'b0 ;
  assign n1722 = n619 ^ n308 ^ 1'b0 ;
  assign n1726 = n630 & n769 ;
  assign n1723 = n1499 ^ n944 ^ 1'b0 ;
  assign n1724 = n812 | n1723 ;
  assign n1725 = n493 & ~n1724 ;
  assign n1727 = n1726 ^ n1725 ^ 1'b0 ;
  assign n1728 = n271 & n1727 ;
  assign n1729 = n701 | n898 ;
  assign n1730 = n1168 & ~n1729 ;
  assign n1731 = n1081 ^ n481 ^ n319 ;
  assign n1732 = ~n1051 & n1731 ;
  assign n1733 = ~n907 & n1311 ;
  assign n1734 = n1733 ^ n70 ^ 1'b0 ;
  assign n1735 = n323 & n862 ;
  assign n1736 = n1735 ^ n542 ^ 1'b0 ;
  assign n1737 = n228 | n922 ;
  assign n1738 = ~n901 & n1226 ;
  assign n1739 = n1738 ^ n477 ^ 1'b0 ;
  assign n1740 = n1026 | n1739 ;
  assign n1741 = n788 ^ n108 ^ 1'b0 ;
  assign n1742 = ~n944 & n1741 ;
  assign n1743 = n847 & ~n1742 ;
  assign n1744 = ~n149 & n1079 ;
  assign n1745 = n34 | n1744 ;
  assign n1746 = n37 | n158 ;
  assign n1747 = n1210 | n1746 ;
  assign n1748 = n1412 ^ n330 ^ 1'b0 ;
  assign n1749 = n1388 ^ n777 ^ 1'b0 ;
  assign n1750 = n1748 & ~n1749 ;
  assign n1751 = n1504 ^ n1105 ^ 1'b0 ;
  assign n1754 = n1158 ^ n277 ^ 1'b0 ;
  assign n1752 = n94 | n927 ;
  assign n1753 = n656 & ~n1752 ;
  assign n1755 = n1754 ^ n1753 ^ 1'b0 ;
  assign n1756 = n328 & n1755 ;
  assign n1757 = n497 & ~n876 ;
  assign n1758 = n364 & n616 ;
  assign n1759 = n1758 ^ n283 ^ 1'b0 ;
  assign n1760 = n921 ^ n433 ^ 1'b0 ;
  assign n1761 = ~n64 & n1220 ;
  assign n1762 = n1761 ^ n1127 ^ 1'b0 ;
  assign n1763 = ~n1513 & n1762 ;
  assign n1764 = n1760 & n1763 ;
  assign n1765 = n89 & ~n963 ;
  assign n1766 = n906 ^ n191 ^ 1'b0 ;
  assign n1767 = n1000 & ~n1709 ;
  assign n1768 = n1767 ^ n228 ^ 1'b0 ;
  assign n1769 = n364 & ~n1313 ;
  assign n1770 = n1769 ^ n528 ^ 1'b0 ;
  assign n1771 = n339 & n737 ;
  assign n1772 = n55 | n1771 ;
  assign n1773 = n1772 ^ n876 ^ 1'b0 ;
  assign n1774 = ~n1499 & n1773 ;
  assign n1775 = n947 & ~n1064 ;
  assign n1776 = n390 | n737 ;
  assign n1777 = n849 | n1776 ;
  assign n1778 = n1777 ^ n666 ^ 1'b0 ;
  assign n1779 = n1775 | n1778 ;
  assign n1780 = n205 & ~n1329 ;
  assign n1781 = n1780 ^ n452 ^ 1'b0 ;
  assign n1782 = n191 | n1781 ;
  assign n1783 = ~n1262 & n1782 ;
  assign n1784 = n596 ^ n452 ^ 1'b0 ;
  assign n1785 = n1385 & n1784 ;
  assign n1786 = n1785 ^ n21 ^ 1'b0 ;
  assign n1788 = n619 ^ n340 ^ 1'b0 ;
  assign n1789 = n158 | n1788 ;
  assign n1787 = ~n454 & n1135 ;
  assign n1790 = n1789 ^ n1787 ^ 1'b0 ;
  assign n1791 = n380 | n470 ;
  assign n1792 = n487 ^ n86 ^ 1'b0 ;
  assign n1793 = n1386 ^ n73 ^ 1'b0 ;
  assign n1794 = n1793 ^ n53 ^ 1'b0 ;
  assign n1795 = ~n934 & n1061 ;
  assign n1796 = n1329 | n1795 ;
  assign n1797 = n1110 & ~n1796 ;
  assign n1798 = n1797 ^ n159 ^ 1'b0 ;
  assign n1799 = n1798 ^ n188 ^ 1'b0 ;
  assign n1800 = n618 & n1799 ;
  assign n1801 = n24 | n215 ;
  assign n1802 = n1801 ^ n172 ^ 1'b0 ;
  assign n1803 = ~n469 & n1458 ;
  assign n1804 = ~n257 & n1803 ;
  assign n1805 = n861 & ~n1804 ;
  assign n1806 = n479 & n1805 ;
  assign n1807 = ~n1348 & n1806 ;
  assign n1809 = n603 ^ n276 ^ 1'b0 ;
  assign n1810 = ~n1430 & n1809 ;
  assign n1808 = ~n1429 & n1598 ;
  assign n1811 = n1810 ^ n1808 ^ 1'b0 ;
  assign n1812 = n398 ^ n78 ^ 1'b0 ;
  assign n1813 = n1388 | n1812 ;
  assign n1814 = n1498 | n1813 ;
  assign n1815 = n1814 ^ n1330 ^ 1'b0 ;
  assign n1816 = ( n52 & n205 ) | ( n52 & ~n367 ) | ( n205 & ~n367 ) ;
  assign n1817 = n435 & ~n971 ;
  assign n1818 = n1164 & ~n1505 ;
  assign n1819 = n122 & n1707 ;
  assign n1820 = n1819 ^ n1478 ^ 1'b0 ;
  assign n1821 = n1595 ^ n1425 ^ n1157 ;
  assign n1822 = n622 ^ n336 ^ 1'b0 ;
  assign n1823 = ~n475 & n700 ;
  assign n1824 = n1823 ^ n731 ^ 1'b0 ;
  assign n1825 = n1822 | n1824 ;
  assign n1826 = n1825 ^ n616 ^ 1'b0 ;
  assign n1827 = n339 & ~n788 ;
  assign n1828 = n55 | n1217 ;
  assign n1829 = n1811 ^ n604 ^ 1'b0 ;
  assign n1830 = x0 & ~n1217 ;
  assign n1831 = n1830 ^ n612 ^ 1'b0 ;
  assign n1832 = n607 ^ n181 ^ 1'b0 ;
  assign n1833 = n793 ^ n210 ^ 1'b0 ;
  assign n1834 = n1358 ^ n83 ^ 1'b0 ;
  assign n1835 = n1834 ^ n1119 ^ 1'b0 ;
  assign n1836 = ~n55 & n732 ;
  assign n1837 = ~n1835 & n1836 ;
  assign n1838 = n1837 ^ n1115 ^ 1'b0 ;
  assign n1839 = n1159 | n1697 ;
  assign n1840 = n432 ^ n198 ^ 1'b0 ;
  assign n1841 = n83 & n1110 ;
  assign n1842 = n390 & ~n690 ;
  assign n1843 = n1227 | n1842 ;
  assign n1844 = n665 & ~n1843 ;
  assign n1845 = n500 & n1677 ;
  assign n1846 = n956 ^ n488 ^ 1'b0 ;
  assign n1847 = ~n55 & n1846 ;
  assign n1849 = n1439 & n1679 ;
  assign n1848 = n703 & n843 ;
  assign n1850 = n1849 ^ n1848 ^ 1'b0 ;
  assign n1851 = n204 & n1850 ;
  assign n1852 = ~n259 & n1165 ;
  assign n1853 = n318 ^ n114 ^ 1'b0 ;
  assign n1854 = n498 & ~n1853 ;
  assign n1855 = n1375 ^ n1063 ^ n82 ;
  assign n1856 = n1854 & ~n1855 ;
  assign n1857 = n1041 | n1165 ;
  assign n1858 = n493 ^ n290 ^ n213 ;
  assign n1859 = ~n649 & n1048 ;
  assign n1862 = n47 & n182 ;
  assign n1863 = ~n185 & n1862 ;
  assign n1860 = n1130 ^ n872 ^ 1'b0 ;
  assign n1861 = n325 | n1860 ;
  assign n1864 = n1863 ^ n1861 ^ 1'b0 ;
  assign n1865 = n582 | n1038 ;
  assign n1866 = n533 & ~n1865 ;
  assign n1867 = n736 & ~n1866 ;
  assign n1868 = n452 & ~n907 ;
  assign n1871 = n1134 & n1311 ;
  assign n1872 = n1871 ^ n80 ^ 1'b0 ;
  assign n1869 = n937 ^ n92 ^ 1'b0 ;
  assign n1870 = n1060 & n1869 ;
  assign n1873 = n1872 ^ n1870 ^ 1'b0 ;
  assign n1874 = n1745 ^ n1588 ^ 1'b0 ;
  assign n1875 = ~n532 & n1721 ;
  assign n1876 = n582 ^ n393 ^ 1'b0 ;
  assign n1877 = n44 | n1876 ;
  assign n1878 = n1877 ^ n323 ^ 1'b0 ;
  assign n1879 = n1179 ^ n155 ^ n17 ;
  assign n1880 = n1043 | n1879 ;
  assign n1881 = n216 & n1787 ;
  assign n1882 = n1270 | n1881 ;
  assign n1883 = n975 | n1882 ;
  assign n1884 = n21 & ~n488 ;
  assign n1885 = n1096 ^ n493 ^ 1'b0 ;
  assign n1886 = x2 & n798 ;
  assign n1887 = n883 & n1886 ;
  assign n1888 = n114 & ~n467 ;
  assign n1889 = ~n472 & n588 ;
  assign n1890 = n1491 ^ n702 ^ 1'b0 ;
  assign n1891 = ~n472 & n1890 ;
  assign n1892 = n1891 ^ n169 ^ 1'b0 ;
  assign n1893 = n1889 | n1892 ;
  assign n1894 = n168 & ~n1622 ;
  assign n1895 = n1894 ^ n749 ^ 1'b0 ;
  assign n1896 = n787 & ~n1166 ;
  assign n1897 = n279 & ~n1177 ;
  assign n1898 = ~n1896 & n1897 ;
  assign n1899 = ~n190 & n1898 ;
  assign n1900 = x7 & n643 ;
  assign n1901 = n1083 & n1900 ;
  assign n1902 = n1095 ^ n665 ^ 1'b0 ;
  assign n1903 = ( n38 & ~n156 ) | ( n38 & n1043 ) | ( ~n156 & n1043 ) ;
  assign n1904 = n1903 ^ n55 ^ 1'b0 ;
  assign n1905 = n573 & n618 ;
  assign n1906 = ~n1904 & n1905 ;
  assign n1907 = n753 | n1888 ;
  assign n1908 = n306 ^ n98 ^ 1'b0 ;
  assign n1909 = n1908 ^ n1789 ^ 1'b0 ;
  assign n1917 = n328 ^ n55 ^ 1'b0 ;
  assign n1910 = n501 & n1304 ;
  assign n1911 = n273 & n1910 ;
  assign n1912 = n1911 ^ n514 ^ 1'b0 ;
  assign n1913 = n1912 ^ n1011 ^ 1'b0 ;
  assign n1914 = n89 & n1283 ;
  assign n1915 = n1051 & n1914 ;
  assign n1916 = ~n1913 & n1915 ;
  assign n1918 = n1917 ^ n1916 ^ 1'b0 ;
  assign n1919 = n328 & n1125 ;
  assign n1920 = ~n184 & n1919 ;
  assign n1923 = n159 & ~n811 ;
  assign n1924 = n1923 ^ n906 ^ 1'b0 ;
  assign n1921 = n1235 ^ n161 ^ 1'b0 ;
  assign n1922 = n715 & n1921 ;
  assign n1925 = n1924 ^ n1922 ^ 1'b0 ;
  assign n1926 = n1920 | n1925 ;
  assign n1927 = n465 ^ x0 ^ 1'b0 ;
  assign n1928 = ~n1213 & n1638 ;
  assign n1929 = n154 | n318 ;
  assign n1930 = ~n246 & n1831 ;
  assign n1931 = ~n1929 & n1930 ;
  assign n1932 = n223 & ~n611 ;
  assign n1933 = n395 & n1380 ;
  assign n1934 = n931 & ~n1323 ;
  assign n1935 = n268 | n1934 ;
  assign n1936 = n1133 & n1379 ;
  assign n1937 = n1135 ^ n1040 ^ 1'b0 ;
  assign n1938 = n1207 & n1937 ;
  assign n1939 = ~n1157 & n1938 ;
  assign n1940 = n119 | n213 ;
  assign n1941 = ~n286 & n1000 ;
  assign n1942 = n1941 ^ n843 ^ 1'b0 ;
  assign n1943 = n641 & ~n1942 ;
  assign n1944 = n618 & n935 ;
  assign n1945 = n177 ^ n168 ^ 1'b0 ;
  assign n1946 = n1945 ^ n1855 ^ 1'b0 ;
  assign n1947 = n1264 & ~n1379 ;
  assign n1948 = n129 & ~n1909 ;
  assign n1949 = n1948 ^ n497 ^ 1'b0 ;
  assign n1950 = ~n128 & n1102 ;
  assign n1953 = n381 ^ n200 ^ 1'b0 ;
  assign n1951 = ~n25 & n102 ;
  assign n1952 = ~n1344 & n1951 ;
  assign n1954 = n1953 ^ n1952 ^ 1'b0 ;
  assign n1955 = ~n1361 & n1750 ;
  assign n1956 = n436 & n1955 ;
  assign n1957 = n438 | n1549 ;
  assign n1958 = n276 | n300 ;
  assign n1959 = n1786 & n1958 ;
  assign n1960 = n35 & n223 ;
  assign n1961 = n141 | n627 ;
  assign n1962 = n899 ^ n133 ^ 1'b0 ;
  assign n1963 = ~n1961 & n1962 ;
  assign n1964 = n233 ^ n158 ^ 1'b0 ;
  assign n1965 = ~n1276 & n1915 ;
  assign n1966 = n1965 ^ n229 ^ 1'b0 ;
  assign n1967 = n646 ^ n128 ^ 1'b0 ;
  assign n1968 = n1666 & n1967 ;
  assign n1969 = n1968 ^ n582 ^ 1'b0 ;
  assign n1970 = n1220 & n1969 ;
  assign n1971 = n547 & ~n1070 ;
  assign n1973 = ~n62 & n129 ;
  assign n1974 = n1973 ^ n291 ^ 1'b0 ;
  assign n1975 = n1974 ^ n1804 ^ 1'b0 ;
  assign n1972 = n535 & ~n867 ;
  assign n1976 = n1975 ^ n1972 ^ 1'b0 ;
  assign n1977 = ~n24 & n1273 ;
  assign n1982 = n492 ^ n486 ^ 1'b0 ;
  assign n1978 = ~n492 & n1495 ;
  assign n1979 = n1978 ^ n839 ^ 1'b0 ;
  assign n1980 = n1979 ^ n1255 ^ 1'b0 ;
  assign n1981 = n527 & ~n1980 ;
  assign n1983 = n1982 ^ n1981 ^ 1'b0 ;
  assign n1984 = n1977 & ~n1983 ;
  assign n1985 = n89 & ~n1676 ;
  assign n1986 = n1985 ^ n522 ^ 1'b0 ;
  assign n1987 = n1069 | n1227 ;
  assign n1988 = n304 ^ n105 ^ 1'b0 ;
  assign n1989 = n1988 ^ n812 ^ 1'b0 ;
  assign n1990 = ~n1987 & n1989 ;
  assign n1991 = ~x4 & n34 ;
  assign n1992 = n188 & ~n1991 ;
  assign n1993 = n483 | n1920 ;
  assign n1994 = n602 | n1993 ;
  assign n1995 = n81 & n1495 ;
  assign n1996 = n1995 ^ n1686 ^ 1'b0 ;
  assign n1997 = n1613 & ~n1996 ;
  assign n2000 = n403 ^ n14 ^ 1'b0 ;
  assign n2001 = ~n1569 & n2000 ;
  assign n2002 = n40 & n2001 ;
  assign n2003 = n23 & n2002 ;
  assign n1998 = n1369 ^ n79 ^ 1'b0 ;
  assign n1999 = n510 | n1998 ;
  assign n2004 = n2003 ^ n1999 ^ 1'b0 ;
  assign n2005 = n618 ^ n512 ^ 1'b0 ;
  assign n2006 = n898 | n1472 ;
  assign n2007 = n36 | n2006 ;
  assign n2008 = ~n1124 & n1412 ;
  assign n2009 = n874 & n2008 ;
  assign n2010 = n2009 ^ n321 ^ 1'b0 ;
  assign n2011 = n284 ^ n135 ^ 1'b0 ;
  assign n2012 = n78 | n873 ;
  assign n2013 = n567 & n636 ;
  assign n2014 = n755 & n2013 ;
  assign n2015 = n354 & ~n1023 ;
  assign n2016 = n2015 ^ n309 ^ 1'b0 ;
  assign n2017 = n356 | n2016 ;
  assign n2018 = n1205 ^ n671 ^ n596 ;
  assign n2019 = n37 & ~n323 ;
  assign n2020 = n294 & n2019 ;
  assign n2021 = n117 | n235 ;
  assign n2022 = n1089 & ~n2021 ;
  assign n2023 = n2020 | n2022 ;
  assign n2024 = n1550 ^ n193 ^ 1'b0 ;
  assign n2025 = ~n2023 & n2024 ;
  assign n2026 = n2025 ^ n713 ^ 1'b0 ;
  assign n2027 = n1541 & n2026 ;
  assign n2028 = n337 & n1690 ;
  assign n2029 = n2028 ^ n441 ^ 1'b0 ;
  assign n2030 = n87 & ~n390 ;
  assign n2031 = ~n2029 & n2030 ;
  assign n2032 = n299 | n880 ;
  assign n2033 = n1026 | n1304 ;
  assign n2034 = n883 | n2033 ;
  assign n2039 = n417 & ~n1430 ;
  assign n2040 = n2039 ^ n872 ^ 1'b0 ;
  assign n2035 = n524 & n738 ;
  assign n2036 = ~n799 & n2035 ;
  assign n2037 = n363 | n546 ;
  assign n2038 = n2036 & ~n2037 ;
  assign n2041 = n2040 ^ n2038 ^ 1'b0 ;
  assign n2042 = n83 & ~n261 ;
  assign n2043 = n2042 ^ x0 ^ 1'b0 ;
  assign n2044 = ~n566 & n2043 ;
  assign n2045 = n812 ^ n753 ^ 1'b0 ;
  assign n2046 = ~n68 & n2045 ;
  assign n2047 = ~n408 & n1325 ;
  assign n2048 = n2047 ^ n1642 ^ 1'b0 ;
  assign n2049 = n2046 & n2048 ;
  assign n2050 = n55 | n1471 ;
  assign n2051 = n337 & ~n458 ;
  assign n2052 = n458 & n2051 ;
  assign n2053 = ~n296 & n1600 ;
  assign n2054 = n296 & n2053 ;
  assign n2055 = n532 ^ n342 ^ 1'b0 ;
  assign n2056 = n2054 | n2055 ;
  assign n2057 = n2052 & ~n2056 ;
  assign n2058 = ( n253 & ~n1763 ) | ( n253 & n2057 ) | ( ~n1763 & n2057 ) ;
  assign n2059 = n269 ^ n62 ^ 1'b0 ;
  assign n2060 = n313 | n1060 ;
  assign n2061 = n296 | n1326 ;
  assign n2062 = n2061 ^ n641 ^ 1'b0 ;
  assign n2063 = n1026 ^ n876 ^ 1'b0 ;
  assign n2064 = n1262 | n1619 ;
  assign n2065 = n2064 ^ n1677 ^ n1250 ;
  assign n2066 = n96 | n1004 ;
  assign n2067 = n197 | n2066 ;
  assign n2070 = n616 | n758 ;
  assign n2068 = n632 & ~n1306 ;
  assign n2069 = n414 & n2068 ;
  assign n2071 = n2070 ^ n2069 ^ 1'b0 ;
  assign n2072 = ~n1029 & n2071 ;
  assign n2073 = ~n1236 & n1302 ;
  assign n2074 = n2073 ^ n353 ^ n292 ;
  assign n2075 = ~n1061 & n2074 ;
  assign n2076 = n159 | n1044 ;
  assign n2077 = n23 | n643 ;
  assign n2078 = n227 | n2077 ;
  assign n2079 = n2076 & n2078 ;
  assign n2080 = n2079 ^ n348 ^ 1'b0 ;
  assign n2081 = n1195 ^ n369 ^ 1'b0 ;
  assign n2082 = n715 & ~n2081 ;
  assign n2083 = n2080 | n2082 ;
  assign n2084 = n128 | n255 ;
  assign n2085 = n2084 ^ n908 ^ 1'b0 ;
  assign n2086 = n931 & ~n2085 ;
  assign n2087 = n1730 | n2086 ;
  assign n2088 = n265 & ~n1585 ;
  assign n2093 = n690 ^ n390 ^ 1'b0 ;
  assign n2089 = ~n608 & n645 ;
  assign n2090 = n2089 ^ n123 ^ 1'b0 ;
  assign n2091 = n551 | n2090 ;
  assign n2092 = n2091 ^ n624 ^ 1'b0 ;
  assign n2094 = n2093 ^ n2092 ^ 1'b0 ;
  assign n2095 = ~n891 & n2094 ;
  assign n2096 = n2088 & n2095 ;
  assign n2097 = n1449 & ~n1479 ;
  assign n2098 = n75 | n1303 ;
  assign n2099 = n2097 | n2098 ;
  assign n2100 = n954 | n2093 ;
  assign n2101 = ~n540 & n1965 ;
  assign n2102 = n2101 ^ n340 ^ 1'b0 ;
  assign n2103 = n1491 ^ n142 ^ 1'b0 ;
  assign n2104 = n1479 ^ n1198 ^ n388 ;
  assign n2105 = n37 & n659 ;
  assign n2106 = n2105 ^ n236 ^ 1'b0 ;
  assign n2107 = x4 & n1283 ;
  assign n2108 = ~n1638 & n2107 ;
  assign n2109 = n1798 ^ n798 ^ n133 ;
  assign n2110 = n195 ^ n92 ^ 1'b0 ;
  assign n2111 = n1859 ^ n284 ^ 1'b0 ;
  assign n2112 = n2110 & n2111 ;
  assign n2113 = n1527 ^ n1059 ^ 1'b0 ;
  assign n2114 = n899 | n2113 ;
  assign n2115 = ~n585 & n748 ;
  assign n2116 = n1095 & n2115 ;
  assign n2117 = ~n363 & n2116 ;
  assign n2118 = n581 | n2117 ;
  assign n2119 = n83 | n2118 ;
  assign n2120 = ~n259 & n856 ;
  assign n2121 = n327 & n2120 ;
  assign n2122 = n2011 & n2121 ;
  assign n2123 = n207 & ~n1015 ;
  assign n2124 = n2123 ^ n86 ^ 1'b0 ;
  assign n2125 = n221 & n448 ;
  assign n2126 = n338 & n2125 ;
  assign n2127 = n2126 ^ n113 ^ 1'b0 ;
  assign n2128 = n489 & n2127 ;
  assign n2129 = n380 & ~n995 ;
  assign n2130 = n288 & n2129 ;
  assign n2131 = n986 ^ n851 ^ 1'b0 ;
  assign n2132 = n929 & ~n1711 ;
  assign n2133 = n2132 ^ n1184 ^ 1'b0 ;
  assign n2134 = n369 & ~n1398 ;
  assign n2135 = n652 | n1004 ;
  assign n2136 = n397 & n649 ;
  assign n2137 = n903 ^ n161 ^ 1'b0 ;
  assign n2138 = ~n177 & n2137 ;
  assign n2139 = n266 | n2011 ;
  assign n2140 = n2138 & ~n2139 ;
  assign n2141 = n608 & ~n1165 ;
  assign n2142 = n1692 ^ n254 ^ 1'b0 ;
  assign n2144 = ~n164 & n251 ;
  assign n2143 = n769 & ~n878 ;
  assign n2145 = n2144 ^ n2143 ^ 1'b0 ;
  assign n2146 = n294 & n527 ;
  assign n2147 = n2146 ^ n745 ^ 1'b0 ;
  assign n2148 = n873 | n2147 ;
  assign n2149 = n1469 ^ n506 ^ 1'b0 ;
  assign n2150 = n2097 & ~n2149 ;
  assign n2151 = ~n468 & n1387 ;
  assign n2152 = n2017 & n2151 ;
  assign n2153 = n685 & n788 ;
  assign n2154 = n2153 ^ n1236 ^ 1'b0 ;
  assign n2155 = n2154 ^ n434 ^ 1'b0 ;
  assign n2156 = n802 | n1900 ;
  assign n2157 = n1025 & ~n1597 ;
  assign n2158 = n2156 | n2157 ;
  assign n2159 = n168 | n2158 ;
  assign n2160 = n1473 ^ n153 ^ 1'b0 ;
  assign n2161 = ~n161 & n357 ;
  assign n2162 = n2161 ^ n774 ^ 1'b0 ;
  assign n2163 = n861 | n2072 ;
  assign n2164 = ~n2012 & n2163 ;
  assign n2165 = n1234 ^ n55 ^ 1'b0 ;
  assign n2166 = n302 & n2165 ;
  assign n2167 = ~n1380 & n2166 ;
  assign n2168 = n986 | n1656 ;
  assign n2169 = n1283 | n2168 ;
  assign n2170 = n82 | n2169 ;
  assign n2171 = n1132 | n2117 ;
  assign n2172 = n2171 ^ n324 ^ 1'b0 ;
  assign n2173 = n1366 ^ n310 ^ 1'b0 ;
  assign n2174 = n359 | n1740 ;
  assign n2175 = n2173 & ~n2174 ;
  assign n2176 = n16 | n364 ;
  assign n2177 = ~n444 & n635 ;
  assign n2178 = n1034 & n2177 ;
  assign n2179 = n400 & n423 ;
  assign n2180 = ( n286 & ~n777 ) | ( n286 & n2179 ) | ( ~n777 & n2179 ) ;
  assign n2181 = n1367 ^ n188 ^ 1'b0 ;
  assign n2182 = n1430 ^ n612 ^ 1'b0 ;
  assign n2183 = ~n290 & n2182 ;
  assign n2184 = n83 & ~n385 ;
  assign n2185 = n200 & n2184 ;
  assign n2186 = n310 & ~n2185 ;
  assign n2187 = n637 ^ n632 ^ 1'b0 ;
  assign n2188 = ~n899 & n2187 ;
  assign n2189 = n191 & n515 ;
  assign n2195 = n284 | n547 ;
  assign n2196 = n292 & ~n2195 ;
  assign n2190 = n324 ^ n228 ^ 1'b0 ;
  assign n2191 = n1281 & n2190 ;
  assign n2192 = n2191 ^ n634 ^ 1'b0 ;
  assign n2193 = ~n520 & n2192 ;
  assign n2194 = n2193 ^ n1742 ^ 1'b0 ;
  assign n2197 = n2196 ^ n2194 ^ 1'b0 ;
  assign n2198 = n2189 & ~n2197 ;
  assign n2199 = n2198 ^ n1308 ^ 1'b0 ;
  assign n2200 = n622 | n642 ;
  assign n2201 = n1263 ^ n425 ^ 1'b0 ;
  assign n2202 = ~n753 & n2201 ;
  assign n2203 = n2202 ^ n1640 ^ 1'b0 ;
  assign n2204 = n241 & ~n557 ;
  assign n2205 = n2196 ^ n1500 ^ 1'b0 ;
  assign n2206 = n1283 ^ n434 ^ 1'b0 ;
  assign n2207 = n1380 & n2206 ;
  assign n2208 = n2205 & n2207 ;
  assign n2209 = n68 & n2208 ;
  assign n2210 = n799 | n1637 ;
  assign n2211 = ~n1170 & n1719 ;
  assign n2212 = n624 & n2211 ;
  assign n2213 = n1205 ^ n996 ^ 1'b0 ;
  assign n2214 = n1531 & n2213 ;
  assign n2215 = n2214 ^ n195 ^ 1'b0 ;
  assign n2216 = ~n2212 & n2215 ;
  assign n2217 = n293 | n1404 ;
  assign n2218 = n2217 ^ n109 ^ 1'b0 ;
  assign n2219 = ~n318 & n768 ;
  assign n2220 = n430 & ~n1562 ;
  assign n2221 = n626 ^ n593 ^ 1'b0 ;
  assign n2222 = ~n2155 & n2221 ;
  assign n2223 = n534 & n627 ;
  assign n2224 = n596 ^ n588 ^ 1'b0 ;
  assign n2225 = n784 & n2224 ;
  assign n2226 = n2225 ^ n1106 ^ 1'b0 ;
  assign n2227 = n2223 & n2226 ;
  assign n2228 = n278 | n549 ;
  assign n2229 = ~n216 & n233 ;
  assign n2230 = n2229 ^ n653 ^ 1'b0 ;
  assign n2231 = ~n1025 & n2230 ;
  assign n2232 = n427 & ~n880 ;
  assign n2233 = n2232 ^ n1105 ^ 1'b0 ;
  assign n2234 = n37 | n2233 ;
  assign n2235 = n1932 | n2234 ;
  assign n2236 = n251 & n279 ;
  assign n2237 = n1311 ^ n1254 ^ 1'b0 ;
  assign n2238 = n2236 & ~n2237 ;
  assign n2239 = n1433 & n1566 ;
  assign n2240 = n2150 ^ n1058 ^ 1'b0 ;
  assign n2241 = n859 | n963 ;
  assign n2242 = n2241 ^ n1971 ^ 1'b0 ;
  assign n2243 = n1880 ^ n196 ^ 1'b0 ;
  assign n2244 = n391 & ~n677 ;
  assign n2245 = n323 ^ n66 ^ 1'b0 ;
  assign n2246 = n1000 | n1219 ;
  assign n2247 = n621 ^ n287 ^ 1'b0 ;
  assign n2248 = n2246 & ~n2247 ;
  assign n2249 = n330 ^ n257 ^ 1'b0 ;
  assign n2250 = ~n284 & n2249 ;
  assign n2251 = n575 & n2250 ;
  assign n2252 = n2151 ^ n912 ^ 1'b0 ;
  assign n2253 = n1063 & n2120 ;
  assign n2254 = n403 & n2253 ;
  assign n2255 = n1024 & ~n2254 ;
  assign n2256 = ~n207 & n2255 ;
  assign n2257 = n2256 ^ n1807 ^ 1'b0 ;
  assign n2258 = n713 | n964 ;
  assign n2259 = n1718 | n2258 ;
  assign n2260 = n2259 ^ n656 ^ 1'b0 ;
  assign n2261 = n1518 | n2260 ;
  assign n2262 = n340 | n508 ;
  assign n2263 = n318 & ~n2262 ;
  assign n2264 = n662 | n2263 ;
  assign n2265 = n2229 & n2264 ;
  assign n2266 = n2265 ^ n701 ^ 1'b0 ;
  assign n2267 = n165 & ~n1330 ;
  assign n2268 = n375 | n556 ;
  assign n2269 = n2268 ^ n719 ^ n253 ;
  assign n2270 = n2269 ^ n1268 ^ 1'b0 ;
  assign n2271 = n567 ^ n456 ^ 1'b0 ;
  assign n2272 = n388 & n2271 ;
  assign n2273 = n1146 ^ n216 ^ 1'b0 ;
  assign n2274 = n859 | n2273 ;
  assign n2275 = n483 & ~n2274 ;
  assign n2276 = n2272 & ~n2275 ;
  assign n2277 = n2276 ^ n1248 ^ 1'b0 ;
  assign n2278 = n2046 ^ n323 ^ 1'b0 ;
  assign n2279 = n2278 ^ n510 ^ 1'b0 ;
  assign n2280 = ~n34 & n927 ;
  assign n2281 = n19 & n721 ;
  assign n2282 = n1091 ^ n853 ^ n683 ;
  assign n2283 = n1334 ^ n857 ^ 1'b0 ;
  assign n2284 = n1095 ^ n43 ^ 1'b0 ;
  assign n2285 = n1175 ^ n314 ^ 1'b0 ;
  assign n2286 = n2284 & n2285 ;
  assign n2287 = ~n744 & n2286 ;
  assign n2288 = n1431 & n2287 ;
  assign n2289 = n336 & n777 ;
  assign n2290 = n1372 & ~n1584 ;
  assign n2291 = n2290 ^ n125 ^ 1'b0 ;
  assign n2292 = ~n69 & n139 ;
  assign n2293 = n850 | n2292 ;
  assign n2294 = n2293 ^ n1854 ^ 1'b0 ;
  assign n2295 = n470 & ~n2294 ;
  assign n2296 = n46 & n297 ;
  assign n2297 = ~n2295 & n2296 ;
  assign n2298 = n1895 ^ n832 ^ 1'b0 ;
  assign n2299 = n2298 ^ n1360 ^ 1'b0 ;
  assign n2300 = n2297 | n2299 ;
  assign n2301 = ( n2289 & ~n2291 ) | ( n2289 & n2300 ) | ( ~n2291 & n2300 ) ;
  assign n2302 = n135 & ~n534 ;
  assign n2303 = n419 & n489 ;
  assign n2304 = ~n418 & n2277 ;
  assign n2305 = ~n336 & n894 ;
  assign n2306 = n1077 | n2305 ;
  assign n2307 = n665 & ~n2306 ;
  assign n2308 = n330 & n2193 ;
  assign n2309 = n408 ^ n37 ^ 1'b0 ;
  assign n2310 = n1531 & ~n2309 ;
  assign n2311 = ~n129 & n1841 ;
  assign n2312 = n1658 ^ n42 ^ 1'b0 ;
  assign n2313 = n2245 & n2312 ;
  assign n2315 = n867 ^ n68 ^ 1'b0 ;
  assign n2316 = n1508 & ~n2315 ;
  assign n2314 = n1974 ^ x6 ^ 1'b0 ;
  assign n2317 = n2316 ^ n2314 ^ 1'b0 ;
  assign n2318 = n2117 ^ n1144 ^ 1'b0 ;
  assign n2319 = n1782 | n2318 ;
  assign n2320 = n406 | n2319 ;
  assign n2321 = n2320 ^ n102 ^ 1'b0 ;
  assign n2322 = n1346 | n2321 ;
  assign n2323 = n402 & n1815 ;
  assign n2324 = ~n247 & n2323 ;
  assign n2325 = ~n321 & n1431 ;
  assign n2326 = ~n1207 & n2325 ;
  assign n2327 = ~n1705 & n2238 ;
  assign n2328 = n2326 & n2327 ;
  assign n2329 = n1113 | n2328 ;
  assign n2330 = n489 | n2329 ;
  assign n2331 = n290 | n2097 ;
  assign n2332 = n1506 ^ n1309 ^ n498 ;
  assign n2333 = n1233 ^ n1135 ^ 1'b0 ;
  assign n2334 = n1036 ^ n443 ^ 1'b0 ;
  assign n2335 = n2334 ^ n1097 ^ 1'b0 ;
  assign n2336 = ~n53 & n549 ;
  assign n2337 = n2336 ^ n1029 ^ 1'b0 ;
  assign n2338 = ~n131 & n2337 ;
  assign n2339 = ~n697 & n2338 ;
  assign n2340 = n1896 ^ n58 ^ 1'b0 ;
  assign n2341 = n1097 | n2340 ;
  assign n2342 = ~n2339 & n2341 ;
  assign n2343 = n609 ^ n161 ^ 1'b0 ;
  assign n2344 = n928 & ~n2343 ;
  assign n2347 = n1216 ^ n117 ^ 1'b0 ;
  assign n2345 = n151 ^ n23 ^ 1'b0 ;
  assign n2346 = ~n1417 & n2345 ;
  assign n2348 = n2347 ^ n2346 ^ 1'b0 ;
  assign n2349 = n1950 | n2070 ;
  assign n2350 = n673 ^ n363 ^ 1'b0 ;
  assign n2351 = n2239 & ~n2350 ;
  assign n2352 = n509 ^ n44 ^ 1'b0 ;
  assign n2353 = ~n1981 & n2352 ;
  assign n2354 = n492 ^ n207 ^ 1'b0 ;
  assign n2355 = n204 & n412 ;
  assign n2356 = ~n2354 & n2355 ;
  assign n2357 = n1001 ^ n553 ^ 1'b0 ;
  assign n2358 = n157 & ~n2357 ;
  assign n2359 = n2358 ^ n311 ^ 1'b0 ;
  assign n2360 = n809 & n2359 ;
  assign n2361 = n1230 ^ n910 ^ 1'b0 ;
  assign n2362 = n1441 ^ n159 ^ 1'b0 ;
  assign n2363 = n528 ^ n273 ^ 1'b0 ;
  assign n2364 = n980 & ~n2363 ;
  assign n2365 = n2364 ^ n678 ^ 1'b0 ;
  assign n2366 = n2362 | n2365 ;
  assign n2367 = n1626 & n1848 ;
  assign n2368 = n1731 & n2367 ;
  assign n2369 = n2368 ^ n338 ^ 1'b0 ;
  assign n2370 = n133 | n2110 ;
  assign n2371 = ~n64 & n1697 ;
  assign n2372 = n1498 ^ n313 ^ 1'b0 ;
  assign n2373 = n2371 & ~n2372 ;
  assign n2374 = n513 & n1664 ;
  assign n2375 = n2374 ^ n630 ^ 1'b0 ;
  assign n2376 = n758 ^ n479 ^ 1'b0 ;
  assign n2377 = n1523 & n2376 ;
  assign n2378 = n2242 & n2358 ;
  assign n2379 = n1887 ^ n769 ^ 1'b0 ;
  assign n2380 = n1345 & ~n2379 ;
  assign n2381 = n671 | n1781 ;
  assign n2382 = n934 & ~n2381 ;
  assign n2383 = n2324 ^ n2073 ^ 1'b0 ;
  assign n2384 = ~n608 & n2383 ;
  assign n2385 = n483 ^ n131 ^ x1 ;
  assign n2386 = ~n455 & n2385 ;
  assign n2390 = n1546 | n2154 ;
  assign n2391 = n722 | n2390 ;
  assign n2387 = n2076 ^ n545 ^ 1'b0 ;
  assign n2388 = n364 & ~n2387 ;
  assign n2389 = n461 & n2388 ;
  assign n2392 = n2391 ^ n2389 ^ 1'b0 ;
  assign n2393 = n204 & ~n2392 ;
  assign n2394 = n2393 ^ n456 ^ 1'b0 ;
  assign n2395 = n1069 & ~n1527 ;
  assign n2396 = n186 & n203 ;
  assign n2397 = n2396 ^ n169 ^ 1'b0 ;
  assign n2398 = n395 | n1113 ;
  assign n2399 = n2397 | n2398 ;
  assign n2400 = n1816 ^ n1414 ^ 1'b0 ;
  assign n2401 = n2400 ^ n812 ^ 1'b0 ;
  assign n2402 = n2362 ^ n553 ^ 1'b0 ;
  assign n2403 = n1024 & ~n2402 ;
  assign n2404 = ( n297 & ~n1511 ) | ( n297 & n1829 ) | ( ~n1511 & n1829 ) ;
  assign n2405 = n76 ^ n72 ^ 1'b0 ;
  assign n2406 = n300 | n2405 ;
  assign n2407 = n154 ^ n37 ^ 1'b0 ;
  assign n2408 = ~n37 & n2407 ;
  assign n2409 = n2408 ^ n996 ^ 1'b0 ;
  assign n2410 = n2406 & ~n2409 ;
  assign n2411 = n701 | n1198 ;
  assign n2412 = n1096 & ~n2411 ;
  assign n2413 = ~n120 & n238 ;
  assign n2414 = n2413 ^ n105 ^ 1'b0 ;
  assign n2415 = n2414 ^ n1227 ^ 1'b0 ;
  assign n2416 = n1339 ^ n649 ^ 1'b0 ;
  assign n2417 = n83 & n2416 ;
  assign n2418 = ~n184 & n2417 ;
  assign n2419 = n1205 ^ n1144 ^ n342 ;
  assign n2421 = ~n60 & n488 ;
  assign n2422 = ~n359 & n2421 ;
  assign n2420 = n76 & ~n177 ;
  assign n2423 = n2422 ^ n2420 ^ 1'b0 ;
  assign n2424 = ~n2065 & n2423 ;
  assign n2425 = n19 & ~n1388 ;
  assign n2427 = ~n546 & n930 ;
  assign n2428 = ~n84 & n2427 ;
  assign n2426 = n765 ^ n412 ^ 1'b0 ;
  assign n2429 = n2428 ^ n2426 ^ 1'b0 ;
  assign n2430 = ~n294 & n2429 ;
  assign n2431 = n1142 ^ n210 ^ 1'b0 ;
  assign n2432 = n512 & n1334 ;
  assign n2433 = n1416 ^ n153 ^ 1'b0 ;
  assign n2434 = n241 & n498 ;
  assign n2435 = n1999 & n2434 ;
  assign n2436 = n461 & n1232 ;
  assign n2437 = n541 | n609 ;
  assign n2438 = ~n323 & n2096 ;
  assign n2439 = ( ~n70 & n236 ) | ( ~n70 & n241 ) | ( n236 & n241 ) ;
  assign n2440 = n311 & ~n2439 ;
  assign n2441 = n2010 ^ n599 ^ 1'b0 ;
  assign n2442 = ~n128 & n2441 ;
  assign n2443 = n2442 ^ n671 ^ 1'b0 ;
  assign n2444 = ~n190 & n294 ;
  assign n2445 = n79 & n2444 ;
  assign n2446 = n2445 ^ n1165 ^ 1'b0 ;
  assign n2447 = n827 ^ n593 ^ 1'b0 ;
  assign n2448 = ~n1986 & n2447 ;
  assign n2449 = n1449 ^ n475 ^ 1'b0 ;
  assign n2450 = ~n192 & n2449 ;
  assign n2451 = n2450 ^ n122 ^ 1'b0 ;
  assign n2452 = n609 & n2451 ;
  assign n2453 = n339 & ~n1298 ;
  assign n2454 = n1142 | n2453 ;
  assign n2455 = n1677 & ~n2150 ;
  assign n2456 = n1441 ^ n659 ^ n74 ;
  assign n2457 = n1367 & n2456 ;
  assign n2458 = n546 & n2457 ;
  assign n2459 = n2458 ^ n2318 ^ 1'b0 ;
  assign n2460 = n1158 & ~n2459 ;
  assign n2461 = n457 & ~n1673 ;
  assign n2462 = n400 & ~n2461 ;
  assign n2463 = n311 & ~n423 ;
  assign n2464 = n912 | n2463 ;
  assign n2465 = n2462 & ~n2464 ;
  assign n2466 = n294 & n1151 ;
  assign n2467 = n2466 ^ n34 ^ 1'b0 ;
  assign n2468 = ~n390 & n714 ;
  assign n2469 = n520 & n2468 ;
  assign n2470 = n493 & ~n2469 ;
  assign n2471 = n2470 ^ n37 ^ 1'b0 ;
  assign n2472 = n2467 | n2471 ;
  assign n2476 = n1471 ^ n157 ^ 1'b0 ;
  assign n2473 = n1695 ^ n491 ^ 1'b0 ;
  assign n2474 = n238 & n2473 ;
  assign n2475 = ~n2470 & n2474 ;
  assign n2477 = n2476 ^ n2475 ^ 1'b0 ;
  assign n2478 = n479 | n745 ;
  assign n2479 = ( n841 & n1989 ) | ( n841 & ~n2478 ) | ( n1989 & ~n2478 ) ;
  assign n2480 = n2479 ^ n468 ^ 1'b0 ;
  assign n2481 = n2480 ^ n161 ^ 1'b0 ;
  assign n2482 = ~n372 & n891 ;
  assign n2483 = n1273 & ~n2482 ;
  assign n2484 = n722 ^ n102 ^ 1'b0 ;
  assign n2485 = n1880 ^ n302 ^ 1'b0 ;
  assign n2486 = n1300 & ~n2376 ;
  assign n2487 = n2136 | n2401 ;
  assign n2489 = n205 | n646 ;
  assign n2488 = n170 & ~n675 ;
  assign n2490 = n2489 ^ n2488 ^ 1'b0 ;
  assign n2491 = ~n83 & n2490 ;
  assign n2492 = n1163 | n1235 ;
  assign n2493 = n2491 | n2492 ;
  assign n2494 = n1352 & ~n2080 ;
  assign n2495 = n789 | n1212 ;
  assign n2496 = n666 ^ n79 ^ 1'b0 ;
  assign n2497 = ~n614 & n1549 ;
  assign n2498 = n2497 ^ n788 ^ 1'b0 ;
  assign n2499 = n1628 & n2498 ;
  assign n2500 = ~n188 & n498 ;
  assign n2501 = ~n866 & n2500 ;
  assign n2502 = n1506 ^ n86 ^ 1'b0 ;
  assign n2503 = n249 & ~n1007 ;
  assign n2504 = n2503 ^ n220 ^ 1'b0 ;
  assign n2505 = n2504 ^ n679 ^ 1'b0 ;
  assign n2506 = n1588 & ~n2505 ;
  assign n2507 = n1415 & n2027 ;
  assign n2508 = n2507 ^ n321 ^ 1'b0 ;
  assign n2509 = x6 | n807 ;
  assign n2510 = n1130 ^ n294 ^ 1'b0 ;
  assign n2511 = n184 & ~n1896 ;
  assign n2512 = n553 & ~n2511 ;
  assign n2513 = ( n227 & n1818 ) | ( n227 & ~n2512 ) | ( n1818 & ~n2512 ) ;
  assign n2514 = n2495 ^ n904 ^ 1'b0 ;
  assign n2515 = n727 & n2320 ;
  assign n2516 = ~n671 & n1158 ;
  assign n2517 = ~n2308 & n2516 ;
  assign n2518 = ~n546 & n825 ;
  assign n2519 = n2518 ^ n354 ^ 1'b0 ;
  assign n2520 = n314 & ~n2519 ;
  assign n2521 = n2520 ^ n129 ^ 1'b0 ;
  assign n2522 = n1001 | n2521 ;
  assign n2523 = n2522 ^ n758 ^ 1'b0 ;
  assign n2524 = n690 ^ n101 ^ 1'b0 ;
  assign n2525 = n2524 ^ n70 ^ 1'b0 ;
  assign n2526 = n1412 & ~n2525 ;
  assign n2527 = n83 & n1943 ;
  assign n2528 = n2527 ^ n272 ^ 1'b0 ;
  assign n2529 = n384 & ~n2528 ;
  assign n2531 = ~n665 & n796 ;
  assign n2532 = n2157 | n2531 ;
  assign n2530 = n488 & n1237 ;
  assign n2533 = n2532 ^ n2530 ^ 1'b0 ;
  assign n2534 = n313 & n1486 ;
  assign n2535 = n2534 ^ n753 ^ 1'b0 ;
  assign n2536 = n375 ^ n17 ^ 1'b0 ;
  assign n2537 = n2073 & ~n2536 ;
  assign n2538 = n512 ^ n417 ^ 1'b0 ;
  assign n2539 = n1154 ^ n1067 ^ 1'b0 ;
  assign n2540 = n2144 & n2539 ;
  assign n2541 = n2538 & n2540 ;
  assign n2542 = ~n723 & n1655 ;
  assign n2543 = ~n622 & n2542 ;
  assign n2544 = n359 & ~n441 ;
  assign n2545 = n546 & n2544 ;
  assign n2546 = ~n1844 & n2545 ;
  assign n2547 = n88 & n206 ;
  assign n2548 = n682 ^ x1 ^ 1'b0 ;
  assign n2549 = n2547 & ~n2548 ;
  assign n2550 = ~n1097 & n2366 ;
  assign n2551 = ~n159 & n2203 ;
  assign n2552 = n1027 & n1309 ;
  assign n2553 = n984 & n2552 ;
  assign n2554 = n500 | n1063 ;
  assign n2555 = n457 ^ n247 ^ 1'b0 ;
  assign n2556 = n2249 & n2555 ;
  assign n2557 = n1341 & n2556 ;
  assign n2558 = n2557 ^ n1034 ^ 1'b0 ;
  assign n2559 = n1891 & n2558 ;
  assign n2560 = ~n2554 & n2559 ;
  assign n2561 = ~n444 & n497 ;
  assign n2562 = n2561 ^ n1088 ^ 1'b0 ;
  assign n2563 = ~n1718 & n2562 ;
  assign n2564 = ~n1210 & n2563 ;
  assign n2565 = n2564 ^ n2135 ^ 1'b0 ;
  assign n2566 = n851 ^ n799 ^ 1'b0 ;
  assign n2567 = n883 ^ n164 ^ 1'b0 ;
  assign n2568 = n2567 ^ n2461 ^ 1'b0 ;
  assign n2569 = ~n1806 & n2491 ;
  assign n2570 = n1500 ^ n247 ^ 1'b0 ;
  assign n2571 = n1146 & ~n2570 ;
  assign n2572 = ~n652 & n2571 ;
  assign n2573 = n683 ^ n443 ^ 1'b0 ;
  assign n2574 = n254 & ~n666 ;
  assign n2575 = ~n2573 & n2574 ;
  assign n2576 = n1179 ^ n412 ^ 1'b0 ;
  assign n2577 = n1086 ^ n993 ^ n647 ;
  assign n2578 = n2577 ^ n1007 ^ 1'b0 ;
  assign n2579 = n364 & ~n1845 ;
  assign n2580 = n2138 & n2579 ;
  assign n2581 = ~n2463 & n2580 ;
  assign n2582 = n1095 ^ n710 ^ 1'b0 ;
  assign n2583 = n2526 & ~n2582 ;
  assign n2584 = n2583 ^ n1067 ^ 1'b0 ;
  assign n2585 = n1000 & n1113 ;
  assign n2586 = n404 ^ n243 ^ 1'b0 ;
  assign n2587 = n497 & n2586 ;
  assign n2591 = x11 | n781 ;
  assign n2592 = n287 & ~n591 ;
  assign n2593 = n2591 & n2592 ;
  assign n2588 = n102 & n332 ;
  assign n2589 = ~n1531 & n2588 ;
  assign n2590 = n905 | n2589 ;
  assign n2594 = n2593 ^ n2590 ^ 1'b0 ;
  assign n2595 = n2431 ^ n2129 ^ 1'b0 ;
  assign n2596 = n246 & n2060 ;
  assign n2597 = n2596 ^ n55 ^ 1'b0 ;
  assign n2598 = n302 | n2597 ;
  assign n2599 = n2129 | n2598 ;
  assign n2600 = n767 & n1777 ;
  assign n2601 = n2449 & n2600 ;
  assign n2602 = n508 ^ n254 ^ 1'b0 ;
  assign n2603 = n2117 | n2602 ;
  assign n2604 = n799 & ~n1785 ;
  assign n2605 = n2604 ^ n758 ^ 1'b0 ;
  assign n2606 = ~n2603 & n2605 ;
  assign n2607 = n646 ^ n608 ^ 1'b0 ;
  assign n2608 = n703 & n2607 ;
  assign n2609 = n1390 ^ n1054 ^ 1'b0 ;
  assign n2610 = n1388 | n2609 ;
  assign n2611 = n2610 ^ n322 ^ n177 ;
  assign n2612 = n356 | n1250 ;
  assign n2613 = n255 & n2571 ;
  assign n2614 = n125 | n961 ;
  assign n2615 = n1017 | n2614 ;
  assign n2616 = ~n77 & n2615 ;
  assign n2617 = ~n2613 & n2616 ;
  assign n2618 = n307 | n1250 ;
  assign n2620 = n1449 ^ n1278 ^ 1'b0 ;
  assign n2621 = n83 & ~n2620 ;
  assign n2619 = n2022 ^ n1267 ^ 1'b0 ;
  assign n2622 = n2621 ^ n2619 ^ 1'b0 ;
  assign n2623 = ~n1671 & n2622 ;
  assign n2624 = ~n92 & n1498 ;
  assign n2625 = x1 & n1207 ;
  assign n2626 = n1920 & n2625 ;
  assign n2627 = n2624 & ~n2626 ;
  assign n2628 = ~n956 & n1529 ;
  assign n2629 = n2628 ^ n288 ^ 1'b0 ;
  assign n2630 = n2629 ^ n1718 ^ 1'b0 ;
  assign n2631 = ~n804 & n984 ;
  assign n2632 = n194 & n1600 ;
  assign n2633 = n2632 ^ n346 ^ 1'b0 ;
  assign n2634 = n719 & n2633 ;
  assign n2635 = ~n2064 & n2634 ;
  assign n2636 = ~n1423 & n2635 ;
  assign n2637 = n2636 ^ n159 ^ 1'b0 ;
  assign n2638 = n1079 & ~n1833 ;
  assign n2639 = n2638 ^ n993 ^ 1'b0 ;
  assign n2640 = n292 | n510 ;
  assign n2641 = n699 & n2640 ;
  assign n2642 = n2641 ^ n1495 ^ 1'b0 ;
  assign n2643 = n2642 ^ n713 ^ 1'b0 ;
  assign n2644 = ~n94 & n2643 ;
  assign n2645 = ~n1323 & n2644 ;
  assign n2646 = ~n2642 & n2645 ;
  assign n2647 = n2646 ^ n2020 ^ 1'b0 ;
  assign n2649 = n297 | n1025 ;
  assign n2648 = ~n294 & n350 ;
  assign n2650 = n2649 ^ n2648 ^ 1'b0 ;
  assign n2651 = n709 & n2650 ;
  assign n2652 = n2651 ^ n2443 ^ 1'b0 ;
  assign n2653 = n549 & n914 ;
  assign n2654 = n2653 ^ n470 ^ 1'b0 ;
  assign n2655 = n2654 ^ n1144 ^ 1'b0 ;
  assign n2656 = n1246 ^ n236 ^ 1'b0 ;
  assign n2657 = n1304 & n2656 ;
  assign n2658 = ~n1206 & n2657 ;
  assign n2659 = ~x8 & n1721 ;
  assign n2660 = n750 ^ n279 ^ 1'b0 ;
  assign n2661 = n956 | n1501 ;
  assign n2662 = n2661 ^ n687 ^ 1'b0 ;
  assign n2663 = ~n745 & n1283 ;
  assign n2664 = n2663 ^ n1697 ^ 1'b0 ;
  assign n2665 = ~n461 & n2664 ;
  assign n2666 = n715 & ~n2258 ;
  assign n2667 = n2666 ^ n1077 ^ 1'b0 ;
  assign n2668 = n227 & n954 ;
  assign n2669 = n1143 | n2668 ;
  assign n2670 = n2669 ^ n530 ^ 1'b0 ;
  assign n2671 = n2061 & n2670 ;
  assign n2672 = ~n2667 & n2671 ;
  assign n2673 = n2672 ^ n2572 ^ 1'b0 ;
  assign n2674 = ~n2672 & n2673 ;
  assign n2675 = n198 | n1690 ;
  assign n2676 = n381 & ~n2675 ;
  assign n2677 = n390 ^ n206 ^ 1'b0 ;
  assign n2678 = n814 ^ x1 ^ 1'b0 ;
  assign n2679 = n1144 & n2678 ;
  assign n2680 = n191 | n293 ;
  assign n2681 = n2679 | n2680 ;
  assign n2682 = ~n83 & n2681 ;
  assign n2683 = n178 & ~n436 ;
  assign n2684 = n2683 ^ n800 ^ 1'b0 ;
  assign n2685 = n1668 ^ n1173 ^ 1'b0 ;
  assign n2686 = ~n2684 & n2685 ;
  assign n2687 = n1381 ^ n745 ^ 1'b0 ;
  assign n2688 = n2562 ^ n2071 ^ 1'b0 ;
  assign n2689 = ~n2687 & n2688 ;
  assign n2690 = n689 ^ n472 ^ 1'b0 ;
  assign n2692 = n1019 & n1531 ;
  assign n2691 = n34 | n907 ;
  assign n2693 = n2692 ^ n2691 ^ 1'b0 ;
  assign n2694 = n2693 ^ n1463 ^ 1'b0 ;
  assign n2695 = n2694 ^ n1015 ^ 1'b0 ;
  assign n2696 = n949 | n988 ;
  assign n2697 = n168 & n2696 ;
  assign n2698 = ~n646 & n2697 ;
  assign n2699 = n2698 ^ n2458 ^ 1'b0 ;
  assign n2700 = n365 ^ n361 ^ 1'b0 ;
  assign n2701 = n2700 ^ n2696 ^ 1'b0 ;
  assign n2702 = n1139 & n2701 ;
  assign n2703 = n1205 ^ n461 ^ 1'b0 ;
  assign n2704 = n208 & n2703 ;
  assign n2705 = n75 | n2704 ;
  assign n2706 = n86 | n139 ;
  assign n2707 = n2706 ^ n514 ^ 1'b0 ;
  assign n2708 = n43 & n1355 ;
  assign n2709 = n2708 ^ n815 ^ 1'b0 ;
  assign n2710 = n1075 & n1360 ;
  assign n2711 = ~n418 & n2710 ;
  assign n2712 = n2711 ^ n2036 ^ 1'b0 ;
  assign n2717 = ~n281 & n694 ;
  assign n2718 = n269 & ~n2717 ;
  assign n2719 = n2718 ^ n263 ^ 1'b0 ;
  assign n2713 = n486 & n703 ;
  assign n2714 = n2713 ^ n261 ^ 1'b0 ;
  assign n2715 = n2714 ^ n515 ^ 1'b0 ;
  assign n2716 = n346 & ~n2715 ;
  assign n2720 = n2719 ^ n2716 ^ 1'b0 ;
  assign n2721 = ~n2004 & n2720 ;
  assign n2722 = ~n454 & n1245 ;
  assign n2723 = n455 & ~n2500 ;
  assign n2724 = n616 ^ n614 ^ 1'b0 ;
  assign n2725 = n1049 & ~n2724 ;
  assign n2726 = n1441 & n2725 ;
  assign n2727 = n1663 ^ n354 ^ n86 ;
  assign n2728 = n2727 ^ n2135 ^ 1'b0 ;
  assign n2729 = n587 & n2364 ;
  assign n2730 = n840 & n2729 ;
  assign n2731 = ~n1404 & n2665 ;
  assign n2732 = n938 & n1031 ;
  assign n2733 = n2714 ^ n332 ^ 1'b0 ;
  assign n2734 = ~n1031 & n2733 ;
  assign n2735 = n2562 & n2734 ;
  assign n2736 = ~n37 & n454 ;
  assign n2738 = ~n325 & n986 ;
  assign n2737 = x3 & ~n169 ;
  assign n2739 = n2738 ^ n2737 ^ 1'b0 ;
  assign n2740 = ~n556 & n802 ;
  assign n2741 = n2739 | n2740 ;
  assign n2742 = ( ~n2480 & n2736 ) | ( ~n2480 & n2741 ) | ( n2736 & n2741 ) ;
  assign n2743 = n2735 | n2742 ;
  assign n2744 = n2732 | n2743 ;
  assign n2745 = ~n139 & n805 ;
  assign n2746 = ~n643 & n2196 ;
  assign n2747 = n2746 ^ n1104 ^ 1'b0 ;
  assign n2748 = ~x0 & n1151 ;
  assign n2749 = n2748 ^ n553 ^ 1'b0 ;
  assign n2750 = n2749 ^ n869 ^ 1'b0 ;
  assign n2751 = n1139 | n2750 ;
  assign n2752 = n2044 | n2751 ;
  assign n2753 = n133 & ~n2752 ;
  assign n2756 = n1409 & ~n1842 ;
  assign n2757 = n2756 ^ n438 ^ 1'b0 ;
  assign n2758 = n221 | n2757 ;
  assign n2759 = n2758 ^ n1588 ^ 1'b0 ;
  assign n2754 = n153 & n510 ;
  assign n2755 = n1904 & ~n2754 ;
  assign n2760 = n2759 ^ n2755 ^ 1'b0 ;
  assign n2761 = n1304 ^ n1112 ^ 1'b0 ;
  assign n2762 = n1525 ^ n284 ^ 1'b0 ;
  assign n2763 = n788 | n2762 ;
  assign n2764 = n2567 & ~n2763 ;
  assign n2766 = n310 & ~n799 ;
  assign n2765 = ~n1708 & n2166 ;
  assign n2767 = n2766 ^ n2765 ^ 1'b0 ;
  assign n2768 = n750 & ~n2767 ;
  assign n2769 = ~n1722 & n2768 ;
  assign n2770 = n1490 ^ n618 ^ 1'b0 ;
  assign n2771 = n75 & n694 ;
  assign n2772 = n1810 ^ n694 ^ 1'b0 ;
  assign n2773 = n1127 & n2772 ;
  assign n2774 = n763 | n1751 ;
  assign n2775 = n628 ^ n608 ^ 1'b0 ;
  assign n2776 = n662 & ~n2775 ;
  assign n2777 = n758 & n2776 ;
  assign n2778 = n2777 ^ n1709 ^ 1'b0 ;
  assign n2779 = ~n1462 & n2778 ;
  assign n2781 = n907 ^ n628 ^ 1'b0 ;
  assign n2782 = n2029 & ~n2781 ;
  assign n2780 = n2478 & ~n2543 ;
  assign n2783 = n2782 ^ n2780 ^ 1'b0 ;
  assign n2784 = ~n924 & n2783 ;
  assign n2785 = ~n229 & n1332 ;
  assign n2786 = n2245 ^ n848 ^ 1'b0 ;
  assign n2787 = n567 | n1241 ;
  assign n2788 = n1089 & n1860 ;
  assign n2789 = n221 | n984 ;
  assign n2794 = n2316 ^ n1645 ^ 1'b0 ;
  assign n2795 = n2110 & ~n2794 ;
  assign n2790 = n1870 ^ n1528 ^ 1'b0 ;
  assign n2791 = n1814 & n2222 ;
  assign n2792 = n2791 ^ n2272 ^ 1'b0 ;
  assign n2793 = n2790 | n2792 ;
  assign n2796 = n2795 ^ n2793 ^ 1'b0 ;
  assign n2797 = n458 | n2141 ;
  assign n2798 = n848 & ~n1206 ;
  assign n2799 = ~n618 & n2798 ;
  assign n2800 = n1857 ^ n1013 ^ 1'b0 ;
  assign n2801 = n1137 | n2800 ;
  assign n2802 = n1140 | n2801 ;
  assign n2803 = n812 | n1432 ;
  assign n2804 = n2803 ^ n1091 ^ 1'b0 ;
  assign n2805 = n1711 | n2804 ;
  assign n2807 = n773 ^ n514 ^ 1'b0 ;
  assign n2806 = n1093 | n2629 ;
  assign n2808 = n2807 ^ n2806 ^ 1'b0 ;
  assign n2809 = n2805 & n2808 ;
  assign n2810 = n1604 ^ n731 ^ 1'b0 ;
  assign n2811 = n1879 & n2613 ;
  assign n2812 = ~n708 & n1047 ;
  assign n2813 = ~n788 & n818 ;
  assign n2814 = n2812 & n2813 ;
  assign n2815 = n577 & n1053 ;
  assign n2816 = n2815 ^ n450 ^ 1'b0 ;
  assign n2817 = ( n629 & ~n1695 ) | ( n629 & n2816 ) | ( ~n1695 & n2816 ) ;
  assign n2818 = ~n2043 & n2681 ;
  assign n2819 = n1931 ^ n1895 ^ 1'b0 ;
  assign n2820 = n70 | n595 ;
  assign n2821 = n2820 ^ n619 ^ 1'b0 ;
  assign n2822 = n653 & n2821 ;
  assign n2825 = n338 ^ n69 ^ 1'b0 ;
  assign n2826 = n135 & ~n2825 ;
  assign n2823 = ~n284 & n639 ;
  assign n2824 = ~n1048 & n2823 ;
  assign n2827 = n2826 ^ n2824 ^ 1'b0 ;
  assign n2828 = n60 | n2827 ;
  assign n2829 = ~n2817 & n2828 ;
  assign n2830 = n359 | n2218 ;
  assign n2831 = n89 | n1854 ;
  assign n2832 = n2220 ^ n622 ^ 1'b0 ;
  assign n2833 = n883 & ~n2832 ;
  assign n2834 = n1195 & n2833 ;
  assign n2835 = n391 ^ n203 ^ 1'b0 ;
  assign n2836 = n513 & ~n2835 ;
  assign n2837 = n364 ^ n158 ^ 1'b0 ;
  assign n2838 = n719 ^ n258 ^ 1'b0 ;
  assign n2839 = ~n1184 & n2838 ;
  assign n2840 = n2839 ^ n1082 ^ 1'b0 ;
  assign n2841 = n861 ^ n28 ^ 1'b0 ;
  assign n2842 = n1185 ^ n582 ^ 1'b0 ;
  assign n2843 = n198 & ~n1876 ;
  assign n2844 = n2843 ^ n700 ^ 1'b0 ;
  assign n2845 = n1346 ^ n390 ^ 1'b0 ;
  assign n2846 = n787 & ~n2845 ;
  assign n2847 = n2846 ^ n2351 ^ 1'b0 ;
  assign n2848 = ~n130 & n445 ;
  assign n2849 = n532 & n1316 ;
  assign n2850 = n533 & ~n2849 ;
  assign n2851 = n542 & ~n964 ;
  assign n2852 = n2851 ^ n2022 ^ 1'b0 ;
  assign n2853 = n144 | n2852 ;
  assign n2854 = n759 & ~n2185 ;
  assign n2855 = ~n232 & n2854 ;
  assign n2856 = ~n284 & n568 ;
  assign n2857 = ~n130 & n2856 ;
  assign n2858 = n2857 ^ n1669 ^ 1'b0 ;
  assign n2859 = ~n158 & n2426 ;
  assign n2860 = n1642 | n2064 ;
  assign n2861 = n330 & ~n794 ;
  assign n2862 = n1884 ^ n1334 ^ 1'b0 ;
  assign n2863 = n55 | n1181 ;
  assign n2864 = n1198 & ~n2863 ;
  assign n2865 = n1287 ^ n1044 ^ 1'b0 ;
  assign n2866 = ~n2701 & n2865 ;
  assign n2867 = n601 ^ n517 ^ 1'b0 ;
  assign n2868 = n2261 ^ n139 ^ 1'b0 ;
  assign n2869 = n60 | n2868 ;
  assign n2870 = n1770 ^ n970 ^ 1'b0 ;
  assign n2871 = x6 & ~n1471 ;
  assign n2872 = n900 & n2871 ;
  assign n2873 = n226 ^ n167 ^ 1'b0 ;
  assign n2874 = n117 & n814 ;
  assign n2875 = n1143 ^ n619 ^ 1'b0 ;
  assign n2876 = n1084 ^ n167 ^ 1'b0 ;
  assign n2877 = n2875 | n2876 ;
  assign n2878 = n649 & ~n2877 ;
  assign n2879 = n688 & n2878 ;
  assign n2880 = n2874 & n2879 ;
  assign n2881 = n66 | n310 ;
  assign n2883 = n281 | n2321 ;
  assign n2882 = n525 | n1810 ;
  assign n2884 = n2883 ^ n2882 ^ 1'b0 ;
  assign n2887 = n1100 ^ n390 ^ 1'b0 ;
  assign n2888 = n2887 ^ n2194 ^ n323 ;
  assign n2885 = n741 ^ n339 ^ 1'b0 ;
  assign n2886 = n2453 | n2885 ;
  assign n2889 = n2888 ^ n2886 ^ 1'b0 ;
  assign n2890 = n2884 & ~n2889 ;
  assign n2891 = ~n2881 & n2890 ;
  assign n2892 = ~n135 & n810 ;
  assign n2893 = ~n2168 & n2892 ;
  assign n2894 = n546 & ~n2633 ;
  assign n2895 = n894 & ~n1067 ;
  assign n2896 = n1546 & n2895 ;
  assign n2897 = n2896 ^ n922 ^ 1'b0 ;
  assign n2898 = x5 | n2897 ;
  assign n2899 = n1278 ^ n741 ^ 1'b0 ;
  assign n2900 = ~n428 & n1463 ;
  assign n2901 = n497 & n1316 ;
  assign n2902 = n2901 ^ n310 ^ 1'b0 ;
  assign n2903 = n87 & n338 ;
  assign n2904 = n1158 | n1382 ;
  assign n2905 = n274 & ~n694 ;
  assign n2906 = n2904 & n2905 ;
  assign n2907 = n227 | n294 ;
  assign n2908 = n2386 ^ n427 ^ 1'b0 ;
  assign n2909 = n169 | n611 ;
  assign n2910 = n2909 ^ n2093 ^ 1'b0 ;
  assign n2911 = n1979 | n2076 ;
  assign n2912 = ( n489 & n1027 ) | ( n489 & n2127 ) | ( n1027 & n2127 ) ;
  assign n2913 = ~n539 & n2912 ;
  assign n2914 = n939 & ~n1720 ;
  assign n2915 = n2146 ^ n2059 ^ 1'b0 ;
  assign n2916 = n822 & ~n2726 ;
  assign n2917 = n1753 ^ n835 ^ 1'b0 ;
  assign n2918 = n1430 ^ n297 ^ 1'b0 ;
  assign n2919 = n66 | n2918 ;
  assign n2920 = n102 | n2919 ;
  assign n2921 = ~n161 & n2920 ;
  assign n2922 = ~n1845 & n2921 ;
  assign n2923 = n2922 ^ n2131 ^ 1'b0 ;
  assign n2924 = n1763 | n2633 ;
  assign n2925 = ~n441 & n1811 ;
  assign n2926 = n776 ^ n593 ^ 1'b0 ;
  assign n2927 = n2925 & ~n2926 ;
  assign n2928 = n2927 ^ n1323 ^ 1'b0 ;
  assign n2929 = ~n462 & n2928 ;
  assign n2930 = ~n233 & n2079 ;
  assign n2931 = n102 & ~n278 ;
  assign n2932 = n2931 ^ n1539 ^ n450 ;
  assign n2933 = ~n2930 & n2932 ;
  assign n2934 = n2724 ^ n400 ^ 1'b0 ;
  assign n2935 = n2347 & n2934 ;
  assign n2936 = n2935 ^ n1637 ^ 1'b0 ;
  assign n2937 = n108 | n1129 ;
  assign n2938 = n555 & n2937 ;
  assign n2939 = n630 | n1845 ;
  assign n2940 = n83 & n2939 ;
  assign n2941 = n2940 ^ n457 ^ 1'b0 ;
  assign n2942 = n2941 ^ n2417 ^ 1'b0 ;
  assign n2943 = n2942 ^ n186 ^ 1'b0 ;
  assign n2944 = n2733 & n2753 ;
  assign n2945 = ~n530 & n2944 ;
  assign n2946 = n2062 ^ n1721 ^ 1'b0 ;
  assign n2947 = n608 ^ n323 ^ 1'b0 ;
  assign n2948 = ~n325 & n1151 ;
  assign n2949 = n387 & n641 ;
  assign n2950 = n2949 ^ n236 ^ 1'b0 ;
  assign n2951 = n703 | n2950 ;
  assign n2952 = n2951 ^ n2825 ^ 1'b0 ;
  assign n2953 = n2948 & ~n2952 ;
  assign n2954 = n158 | n1660 ;
  assign n2955 = n995 & ~n2954 ;
  assign n2956 = n1167 & ~n2955 ;
  assign n2957 = n549 & ~n581 ;
  assign n2958 = n2957 ^ n1555 ^ 1'b0 ;
  assign n2959 = n2956 & n2958 ;
  assign n2960 = n825 & n1000 ;
  assign n2961 = n917 & n2960 ;
  assign n2962 = n385 & n506 ;
  assign n2963 = n2961 & n2962 ;
  assign n2964 = n618 & n1546 ;
  assign n2965 = n381 | n2964 ;
  assign n2966 = n2414 & ~n2965 ;
  assign n2967 = n1701 | n2966 ;
  assign n2968 = n792 & ~n1133 ;
  assign n2969 = n1273 ^ n300 ^ 1'b0 ;
  assign n2970 = n1192 & ~n2889 ;
  assign n2971 = n2970 ^ n1726 ^ 1'b0 ;
  assign n2972 = n1531 & ~n1611 ;
  assign n2973 = n1250 & ~n2972 ;
  assign n2974 = n1044 & n2910 ;
  assign n2975 = ( n24 & ~n2154 ) | ( n24 & n2974 ) | ( ~n2154 & n2974 ) ;
  assign n2976 = ~n1450 & n1873 ;
  assign n2977 = n2976 ^ n2150 ^ 1'b0 ;
  assign n2978 = x2 | n2977 ;
  assign n2979 = n2150 ^ n1229 ^ n1199 ;
  assign n2980 = ~n538 & n1245 ;
  assign n2981 = n2644 ^ n806 ^ 1'b0 ;
  assign n2982 = n2980 & n2981 ;
  assign n2983 = n172 & n1057 ;
  assign n2984 = n996 | n2154 ;
  assign n2985 = n2983 & n2984 ;
  assign n2986 = n2985 ^ n1435 ^ 1'b0 ;
  assign n2987 = n2018 ^ x0 ^ 1'b0 ;
  assign n2988 = n184 & ~n2987 ;
  assign n2989 = n2824 ^ n776 ^ 1'b0 ;
  assign n2990 = ~n1865 & n2989 ;
  assign n2991 = n1254 ^ n314 ^ 1'b0 ;
  assign n2998 = n1328 ^ n491 ^ 1'b0 ;
  assign n2992 = ~n139 & n866 ;
  assign n2993 = n487 & n704 ;
  assign n2994 = n2993 ^ n321 ^ 1'b0 ;
  assign n2995 = n2994 ^ n268 ^ 1'b0 ;
  assign n2996 = n2992 & n2995 ;
  assign n2997 = n2996 ^ n113 ^ 1'b0 ;
  assign n2999 = n2998 ^ n2997 ^ 1'b0 ;
  assign n3000 = n1929 ^ n582 ^ 1'b0 ;
  assign n3001 = n1234 & ~n3000 ;
  assign n3002 = n1089 ^ n536 ^ 1'b0 ;
  assign n3003 = n2105 ^ n1499 ^ 1'b0 ;
  assign n3004 = n278 & ~n3003 ;
  assign n3005 = n3004 ^ n294 ^ 1'b0 ;
  assign n3006 = n3005 ^ n235 ^ 1'b0 ;
  assign n3007 = n52 | n3006 ;
  assign n3008 = n155 & ~n507 ;
  assign n3009 = n3008 ^ n76 ^ 1'b0 ;
  assign n3010 = ~n1854 & n2261 ;
  assign n3012 = n1016 ^ n169 ^ 1'b0 ;
  assign n3013 = n3012 ^ n1044 ^ 1'b0 ;
  assign n3011 = n314 & ~n483 ;
  assign n3014 = n3013 ^ n3011 ^ 1'b0 ;
  assign n3021 = n1473 ^ n1163 ^ 1'b0 ;
  assign n3016 = n102 & ~n1766 ;
  assign n3017 = n1441 & n3016 ;
  assign n3015 = n694 & n1961 ;
  assign n3018 = n3017 ^ n3015 ^ 1'b0 ;
  assign n3019 = n1848 & n3018 ;
  assign n3020 = ~n246 & n3019 ;
  assign n3022 = n3021 ^ n3020 ^ 1'b0 ;
  assign n3023 = ~n2137 & n2891 ;
  assign n3024 = ~n1205 & n2640 ;
  assign n3025 = n129 ^ n21 ^ 1'b0 ;
  assign n3026 = n3025 ^ n713 ^ 1'b0 ;
  assign n3027 = ~n2568 & n3026 ;
  assign n3028 = ~n1100 & n1330 ;
  assign n3029 = ~n68 & n223 ;
  assign n3030 = ~n1166 & n3029 ;
  assign n3031 = n928 ^ n129 ^ 1'b0 ;
  assign n3032 = n170 & n3031 ;
  assign n3033 = n318 & n3032 ;
  assign n3034 = n653 & ~n927 ;
  assign n3035 = n3034 ^ n400 ^ 1'b0 ;
  assign n3036 = ~n3033 & n3035 ;
  assign n3037 = n3036 ^ n2674 ^ 1'b0 ;
  assign n3038 = n1764 | n2572 ;
  assign n3039 = n3038 ^ n2639 ^ 1'b0 ;
  assign n3040 = n2977 & ~n3039 ;
  assign n3041 = n1906 | n2788 ;
  assign n3042 = n3041 ^ n364 ^ 1'b0 ;
  assign n3043 = n2020 ^ n1104 ^ 1'b0 ;
  assign n3044 = ~n1880 & n3043 ;
  assign n3045 = n1573 ^ n1546 ^ 1'b0 ;
  assign n3046 = n2739 & n3045 ;
  assign n3047 = n818 & ~n3046 ;
  assign n3048 = n3047 ^ n1875 ^ 1'b0 ;
  assign n3049 = n2474 & ~n3048 ;
  assign n3050 = n458 ^ n425 ^ 1'b0 ;
  assign n3051 = ~n729 & n3023 ;
  assign n3052 = ~n322 & n2134 ;
  assign n3053 = n847 & n3052 ;
  assign n3054 = ~n1239 & n2142 ;
  assign n3055 = n135 & n2361 ;
  assign n3056 = n3055 ^ n827 ^ 1'b0 ;
  assign n3057 = n2220 ^ n701 ^ 1'b0 ;
  assign n3058 = ~n599 & n1929 ;
  assign n3059 = n3058 ^ n665 ^ 1'b0 ;
  assign n3060 = n412 & n3059 ;
  assign n3061 = n3060 ^ n737 ^ 1'b0 ;
  assign n3062 = n196 & n842 ;
  assign n3063 = n3062 ^ n626 ^ 1'b0 ;
  assign n3064 = n3063 ^ n1027 ^ 1'b0 ;
  assign n3065 = n2947 ^ n1751 ^ 1'b0 ;
  assign n3066 = n1223 & ~n3065 ;
  assign n3067 = ~n872 & n3066 ;
  assign n3068 = ~n2295 & n2939 ;
  assign n3069 = n694 & ~n3068 ;
  assign n3070 = n530 | n1205 ;
  assign n3071 = n690 & ~n3070 ;
  assign n3072 = ( n86 & n159 ) | ( n86 & ~n3071 ) | ( n159 & ~n3071 ) ;
  assign n3073 = n3072 ^ n570 ^ 1'b0 ;
  assign n3074 = n1165 | n3073 ;
  assign n3075 = n3074 ^ n461 ^ 1'b0 ;
  assign n3076 = n385 & n2384 ;
  assign n3077 = n3076 ^ n64 ^ 1'b0 ;
  assign n3078 = n139 & n869 ;
  assign n3079 = n78 & ~n2684 ;
  assign n3080 = n3079 ^ n512 ^ 1'b0 ;
  assign n3081 = n212 & ~n2591 ;
  assign n3082 = n2394 & ~n3081 ;
  assign n3083 = n3082 ^ n1090 ^ 1'b0 ;
  assign n3084 = n226 | n2292 ;
  assign n3085 = n2891 & ~n3084 ;
  assign n3086 = n717 ^ n85 ^ 1'b0 ;
  assign n3087 = n758 | n3086 ;
  assign n3088 = n3087 ^ n1845 ^ 1'b0 ;
  assign n3089 = n3088 ^ n832 ^ 1'b0 ;
  assign n3090 = n1173 & n1630 ;
  assign n3091 = n3090 ^ n2134 ^ 1'b0 ;
  assign n3092 = n1591 ^ n1538 ^ 1'b0 ;
  assign n3093 = ~n1906 & n3092 ;
  assign n3094 = ~n133 & n622 ;
  assign n3095 = n609 & n3094 ;
  assign n3096 = n1407 | n2179 ;
  assign n3097 = ~n3095 & n3096 ;
  assign n3098 = n3097 ^ n2934 ^ 1'b0 ;
  assign n3099 = n196 & n1895 ;
  assign n3100 = ~n337 & n787 ;
  assign n3101 = n3100 ^ n460 ^ 1'b0 ;
  assign n3102 = n3101 ^ n1965 ^ 1'b0 ;
  assign n3103 = n1493 | n3102 ;
  assign n3104 = n838 ^ x11 ^ 1'b0 ;
  assign n3105 = n291 & ~n1001 ;
  assign n3106 = n3105 ^ n2853 ^ 1'b0 ;
  assign n3107 = n724 | n2958 ;
  assign n3108 = n491 & n1676 ;
  assign n3109 = n405 | n3108 ;
  assign n3110 = ~n671 & n1224 ;
  assign n3111 = n1385 & n1668 ;
  assign n3112 = ~n3110 & n3111 ;
  assign n3113 = n3112 ^ n1193 ^ 1'b0 ;
  assign n3114 = ~n3109 & n3113 ;
  assign n3115 = n2283 ^ n681 ^ 1'b0 ;
  assign n3116 = n38 ^ n37 ^ 1'b0 ;
  assign n3117 = n205 & ~n1097 ;
  assign n3118 = ~n527 & n3117 ;
  assign n3119 = n133 & ~n3118 ;
  assign n3120 = n3119 ^ n880 ^ 1'b0 ;
  assign n3121 = n1224 | n2469 ;
  assign n3122 = n3121 ^ n1660 ^ 1'b0 ;
  assign n3123 = n1863 ^ n1552 ^ 1'b0 ;
  assign n3124 = n43 & n302 ;
  assign n3125 = n3124 ^ n1023 ^ 1'b0 ;
  assign n3126 = n3125 ^ n1325 ^ 1'b0 ;
  assign n3127 = n804 | n1903 ;
  assign n3128 = ~n1286 & n1527 ;
  assign n3129 = n2198 & ~n3128 ;
  assign n3130 = n3129 ^ n2704 ^ 1'b0 ;
  assign n3131 = n3130 ^ n1085 ^ 1'b0 ;
  assign n3132 = n81 & n624 ;
  assign n3133 = ~n577 & n3132 ;
  assign n3134 = n1455 | n3133 ;
  assign n3135 = n3134 ^ n581 ^ 1'b0 ;
  assign n3136 = n299 & n1820 ;
  assign n3137 = n3136 ^ n1143 ^ 1'b0 ;
  assign n3138 = n1945 ^ n129 ^ 1'b0 ;
  assign n3139 = n2717 ^ n108 ^ 1'b0 ;
  assign n3140 = n48 | n3139 ;
  assign n3141 = n3140 ^ n156 ^ 1'b0 ;
  assign n3142 = n3141 ^ n232 ^ 1'b0 ;
  assign n3143 = ~n665 & n3142 ;
  assign n3144 = n3143 ^ n158 ^ 1'b0 ;
  assign n3145 = n3138 & n3144 ;
  assign n3146 = n3145 ^ n310 ^ 1'b0 ;
  assign n3148 = ~n55 & n3007 ;
  assign n3149 = n3148 ^ n135 ^ 1'b0 ;
  assign n3147 = ~n678 & n1630 ;
  assign n3150 = n3149 ^ n3147 ^ 1'b0 ;
  assign n3151 = ~n2348 & n3150 ;
  assign n3152 = n3151 ^ n618 ^ 1'b0 ;
  assign n3153 = n1499 | n2531 ;
  assign n3154 = n412 | n3153 ;
  assign n3155 = n1567 | n3007 ;
  assign n3156 = n3155 ^ n2459 ^ 1'b0 ;
  assign n3157 = n215 ^ n170 ^ 1'b0 ;
  assign n3158 = n1538 | n3157 ;
  assign n3159 = n1910 ^ n638 ^ 1'b0 ;
  assign n3160 = ~n1922 & n3159 ;
  assign n3161 = n700 ^ n37 ^ 1'b0 ;
  assign n3162 = n2882 & n3161 ;
  assign n3163 = n694 | n1205 ;
  assign n3164 = n286 & ~n3163 ;
  assign n3165 = n3164 ^ n2188 ^ 1'b0 ;
  assign n3166 = n1541 & n3165 ;
  assign n3167 = n419 ^ x6 ^ 1'b0 ;
  assign n3168 = n252 | n912 ;
  assign n3169 = n3168 ^ n2223 ^ 1'b0 ;
  assign n3170 = n1874 ^ n520 ^ 1'b0 ;
  assign n3171 = n3169 & ~n3170 ;
  assign n3172 = n582 ^ n30 ^ 1'b0 ;
  assign n3173 = n3171 & ~n3172 ;
  assign n3174 = n1620 ^ n419 ^ 1'b0 ;
  assign n3175 = n602 & ~n3174 ;
  assign n3176 = n723 & ~n812 ;
  assign n3177 = n2514 & n3176 ;
  assign n3178 = n506 & ~n1539 ;
  assign n3179 = n3178 ^ n1224 ^ 1'b0 ;
  assign n3180 = n1538 | n1909 ;
  assign n3181 = n2187 | n3124 ;
  assign n3182 = n3181 ^ n83 ^ 1'b0 ;
  assign n3183 = n3182 ^ n1550 ^ 1'b0 ;
  assign n3184 = n2825 ^ n540 ^ 1'b0 ;
  assign n3185 = n3183 & n3184 ;
  assign n3186 = ~n585 & n2382 ;
  assign n3187 = ~n493 & n2939 ;
  assign n3188 = n313 & n3187 ;
  assign n3189 = n1233 & n3188 ;
  assign n3190 = n3189 ^ n2151 ^ 1'b0 ;
  assign n3191 = n1363 & ~n3190 ;
  assign n3192 = n2304 ^ n847 ^ 1'b0 ;
  assign n3193 = n982 & n1271 ;
  assign n3194 = n281 & n295 ;
  assign n3195 = n3194 ^ n459 ^ 1'b0 ;
  assign n3196 = ~n708 & n3195 ;
  assign n3197 = n1987 & n3196 ;
  assign n3198 = n51 & n52 ;
  assign n3199 = n2148 & n3198 ;
  assign n3200 = n2152 ^ n2114 ^ 1'b0 ;
  assign n3201 = ~n1935 & n3200 ;
  assign n3202 = ~n743 & n3201 ;
  assign n3203 = n1146 ^ n102 ^ 1'b0 ;
  assign n3204 = n1988 ^ n337 ^ 1'b0 ;
  assign n3205 = n1406 | n2148 ;
  assign n3206 = n3204 & ~n3205 ;
  assign n3207 = n310 | n3206 ;
  assign n3208 = n1848 & n2571 ;
  assign n3209 = n2964 ^ n1194 ^ 1'b0 ;
  assign n3210 = n3209 ^ n758 ^ 1'b0 ;
  assign n3211 = n3208 & n3210 ;
  assign n3212 = n903 ^ n200 ^ 1'b0 ;
  assign n3213 = n2667 ^ n323 ^ 1'b0 ;
  assign n3214 = n2647 & ~n3213 ;
  assign n3215 = ~n1348 & n2228 ;
  assign n3216 = n3025 & n3215 ;
  assign n3217 = ~n322 & n2281 ;
  assign n3218 = n2014 & ~n2693 ;
  assign n3219 = n1078 ^ n839 ^ 1'b0 ;
  assign n3220 = x11 | n567 ;
  assign n3221 = n1194 ^ n294 ^ 1'b0 ;
  assign n3222 = n1040 & n1566 ;
  assign n3223 = n1889 & n3222 ;
  assign n3224 = n332 & ~n3223 ;
  assign n3225 = n1581 | n3224 ;
  assign n3226 = n661 & ~n1672 ;
  assign n3227 = n1475 & n2751 ;
  assign n3228 = n1686 & n2426 ;
  assign n3229 = n75 | n1411 ;
  assign n3230 = n1010 & n1887 ;
  assign n3231 = ~n251 & n3230 ;
  assign n3232 = n1341 & ~n3012 ;
  assign n3233 = n588 & n3232 ;
  assign n3234 = n666 ^ n52 ^ 1'b0 ;
  assign n3235 = n98 & ~n3234 ;
  assign n3236 = ~n2318 & n3235 ;
  assign n3237 = n2273 & n3236 ;
  assign n3238 = n3237 ^ n2173 ^ 1'b0 ;
  assign n3239 = n551 & ~n2260 ;
  assign n3240 = ~n799 & n836 ;
  assign n3241 = n839 & ~n1044 ;
  assign n3242 = n3241 ^ n149 ^ 1'b0 ;
  assign n3243 = n340 ^ n151 ^ 1'b0 ;
  assign n3244 = n2604 ^ n1630 ^ 1'b0 ;
  assign n3245 = ~n1113 & n2829 ;
  assign n3246 = n630 & n1342 ;
  assign n3247 = n279 & n1629 ;
  assign n3248 = n3133 & ~n3247 ;
  assign n3249 = n1198 ^ n657 ^ 1'b0 ;
  assign n3250 = n241 & n2220 ;
  assign n3251 = ~n3249 & n3250 ;
  assign n3252 = n3251 ^ n917 ^ 1'b0 ;
  assign n3253 = ~n2973 & n3252 ;
  assign n3254 = n3253 ^ n627 ^ 1'b0 ;
  assign n3255 = ~n2136 & n2785 ;
  assign n3264 = n195 | n758 ;
  assign n3263 = n1198 ^ n807 ^ 1'b0 ;
  assign n3256 = ~n295 & n2700 ;
  assign n3257 = n1361 ^ n174 ^ 1'b0 ;
  assign n3258 = ~n3081 & n3257 ;
  assign n3259 = n2547 & n3258 ;
  assign n3260 = ~n3256 & n3259 ;
  assign n3261 = n2811 & ~n2812 ;
  assign n3262 = n3260 & n3261 ;
  assign n3265 = n3264 ^ n3263 ^ n3262 ;
  assign n3266 = n3191 ^ n2603 ^ 1'b0 ;
  assign n3267 = n476 & ~n1655 ;
  assign n3268 = n2337 ^ n662 ^ n16 ;
  assign n3269 = n1314 & n1385 ;
  assign n3270 = n46 & n1344 ;
  assign n3271 = n1387 | n3270 ;
  assign n3272 = n510 | n3271 ;
  assign n3273 = n3272 ^ n604 ^ 1'b0 ;
  assign n3274 = n380 | n3273 ;
  assign n3275 = ~n616 & n825 ;
  assign n3276 = n3275 ^ n1377 ^ 1'b0 ;
  assign n3277 = n1285 | n3276 ;
  assign n3278 = n2063 | n2959 ;
  assign n3279 = n622 & n804 ;
  assign n3280 = n157 & ~n3279 ;
  assign n3281 = n2494 ^ n2270 ^ 1'b0 ;
  assign n3282 = n322 & n3281 ;
  assign n3283 = n1233 ^ n939 ^ 1'b0 ;
  assign n3284 = n3283 ^ n1895 ^ 1'b0 ;
  assign n3285 = n2403 ^ n929 ^ n30 ;
  assign n3286 = n1504 & n2465 ;
  assign n3287 = ~n83 & n1142 ;
  assign n3288 = n1157 & n1827 ;
  assign n3289 = n3288 ^ n2932 ^ 1'b0 ;
  assign n3290 = n1719 ^ n793 ^ 1'b0 ;
  assign n3293 = n2239 ^ n323 ^ 1'b0 ;
  assign n3291 = n1134 | n2842 ;
  assign n3292 = n3291 ^ n2667 ^ 1'b0 ;
  assign n3294 = n3293 ^ n3292 ^ 1'b0 ;
  assign n3295 = n3290 & n3294 ;
  assign n3296 = n128 | n241 ;
  assign n3297 = x8 | n3296 ;
  assign n3298 = n359 & n3297 ;
  assign n3299 = n384 | n3298 ;
  assign n3300 = n448 & ~n1264 ;
  assign n3301 = ~n1231 & n3300 ;
  assign n3302 = x11 & ~n1676 ;
  assign n3303 = ~n3301 & n3302 ;
  assign n3304 = ~n1059 & n1630 ;
  assign n3305 = ~n1230 & n2322 ;
  assign n3306 = ( n748 & n823 ) | ( n748 & n2881 ) | ( n823 & n2881 ) ;
  assign n3307 = n1403 ^ n856 ^ 1'b0 ;
  assign n3308 = n2245 & n2677 ;
  assign n3309 = n3308 ^ n748 ^ 1'b0 ;
  assign n3311 = n1175 ^ n935 ^ 1'b0 ;
  assign n3310 = n806 & ~n1227 ;
  assign n3312 = n3311 ^ n3310 ^ 1'b0 ;
  assign n3313 = n2916 ^ n2200 ^ 1'b0 ;
  assign n3314 = n3312 | n3313 ;
  assign n3318 = n2431 & n2696 ;
  assign n3315 = n1433 ^ n938 ^ 1'b0 ;
  assign n3316 = n3315 ^ n3034 ^ 1'b0 ;
  assign n3317 = n194 & ~n3316 ;
  assign n3319 = n3318 ^ n3317 ^ 1'b0 ;
  assign n3320 = n671 & ~n3319 ;
  assign n3321 = n546 & n713 ;
  assign n3322 = n1867 | n3144 ;
  assign n3323 = n60 | n2459 ;
  assign n3324 = n3323 ^ x0 ^ 1'b0 ;
  assign n3325 = n3322 & ~n3324 ;
  assign n3326 = n1781 ^ n628 ^ 1'b0 ;
  assign n3327 = n2261 | n3326 ;
  assign n3328 = n1988 ^ n1931 ^ 1'b0 ;
  assign n3329 = n1017 & ~n3328 ;
  assign n3330 = n1172 ^ n34 ^ 1'b0 ;
  assign n3331 = n1207 & ~n3330 ;
  assign n3332 = n556 ^ n441 ^ 1'b0 ;
  assign n3333 = ~n1416 & n3332 ;
  assign n3334 = ( n2321 & ~n3331 ) | ( n2321 & n3333 ) | ( ~n3331 & n3333 ) ;
  assign n3335 = n1135 ^ n695 ^ 1'b0 ;
  assign n3336 = n979 & ~n1737 ;
  assign n3337 = ~n184 & n3336 ;
  assign n3338 = n2172 ^ n90 ^ 1'b0 ;
  assign n3339 = n290 & ~n598 ;
  assign n3340 = n789 & n1988 ;
  assign n3341 = ~n3339 & n3340 ;
  assign n3342 = n2414 ^ n1792 ^ 1'b0 ;
  assign n3343 = n833 ^ n636 ^ 1'b0 ;
  assign n3344 = n3343 ^ n938 ^ 1'b0 ;
  assign n3345 = n3342 & n3344 ;
  assign n3346 = n236 & n628 ;
  assign n3347 = n55 & n3346 ;
  assign n3348 = n1886 ^ n1205 ^ n495 ;
  assign n3350 = n133 & n629 ;
  assign n3351 = n3350 ^ n517 ^ 1'b0 ;
  assign n3352 = ~n683 & n3351 ;
  assign n3349 = n1013 & n2214 ;
  assign n3353 = n3352 ^ n3349 ^ n1080 ;
  assign n3354 = n879 & ~n2125 ;
  assign n3355 = n338 ^ n141 ^ 1'b0 ;
  assign n3356 = n626 | n789 ;
  assign n3357 = ( n218 & ~n294 ) | ( n218 & n1386 ) | ( ~n294 & n1386 ) ;
  assign n3358 = n3357 ^ n68 ^ 1'b0 ;
  assign n3359 = n78 | n3358 ;
  assign n3360 = n58 & ~n2339 ;
  assign n3361 = n1302 & n3360 ;
  assign n3362 = n283 & ~n2200 ;
  assign n3363 = n1219 | n3362 ;
  assign n3364 = n442 ^ x7 ^ 1'b0 ;
  assign n3365 = n1432 | n3364 ;
  assign n3366 = n3365 ^ n807 ^ n754 ;
  assign n3367 = n1015 & ~n3366 ;
  assign n3368 = n643 & ~n3367 ;
  assign n3369 = n1777 ^ n910 ^ 1'b0 ;
  assign n3370 = n3369 ^ n2108 ^ 1'b0 ;
  assign n3371 = n3370 ^ n66 ^ 1'b0 ;
  assign n3372 = ~x8 & n1520 ;
  assign n3373 = n3372 ^ n1744 ^ 1'b0 ;
  assign n3374 = n323 & ~n3373 ;
  assign n3375 = n2127 ^ n557 ^ 1'b0 ;
  assign n3376 = n791 & ~n3375 ;
  assign n3377 = x11 | n3376 ;
  assign n3378 = n3176 ^ n2986 ^ 1'b0 ;
  assign n3379 = ~n906 & n1476 ;
  assign n3380 = ~n1592 & n3379 ;
  assign n3381 = n976 ^ n205 ^ 1'b0 ;
  assign n3382 = n976 & n3381 ;
  assign n3383 = n2898 | n3342 ;
  assign n3384 = n3382 | n3383 ;
  assign n3385 = n1245 ^ n475 ^ 1'b0 ;
  assign n3386 = n963 & ~n3118 ;
  assign n3387 = n1346 ^ n1118 ^ 1'b0 ;
  assign n3388 = n3188 ^ n962 ^ 1'b0 ;
  assign n3389 = n3387 & n3388 ;
  assign n3390 = n2004 ^ n1366 ^ 1'b0 ;
  assign n3391 = n3098 ^ n2881 ^ 1'b0 ;
  assign n3392 = n70 | n3391 ;
  assign n3393 = n596 & ~n3312 ;
  assign n3394 = n3393 ^ n997 ^ 1'b0 ;
  assign n3395 = ~n52 & n423 ;
  assign n3396 = n1957 & ~n2953 ;
  assign n3397 = n690 | n3396 ;
  assign n3398 = n1668 | n3397 ;
  assign n3399 = ~n75 & n1048 ;
  assign n3400 = n83 & ~n1601 ;
  assign n3401 = n191 & n3400 ;
  assign n3402 = ~n135 & n475 ;
  assign n3403 = n36 & n2375 ;
  assign n3404 = n489 & n954 ;
  assign n3405 = n3404 ^ n1235 ^ 1'b0 ;
  assign n3406 = n2490 ^ n1462 ^ n330 ;
  assign n3407 = n3406 ^ n1316 ^ 1'b0 ;
  assign n3408 = n3364 ^ n750 ^ 1'b0 ;
  assign n3409 = n246 & n1619 ;
  assign n3410 = n252 & ~n3409 ;
  assign n3411 = n3408 & n3410 ;
  assign n3412 = ( n616 & n963 ) | ( n616 & n1250 ) | ( n963 & n1250 ) ;
  assign n3413 = ~n1056 & n2284 ;
  assign n3414 = n2430 & n3413 ;
  assign n3415 = n2661 ^ n616 ^ n465 ;
  assign n3416 = n3032 ^ n1659 ^ 1'b0 ;
  assign n3417 = n2611 ^ n1743 ^ 1'b0 ;
  assign n3418 = ( n185 & n3416 ) | ( n185 & n3417 ) | ( n3416 & n3417 ) ;
  assign n3419 = n1532 ^ n295 ^ 1'b0 ;
  assign n3420 = n1161 & ~n3419 ;
  assign n3421 = n3420 ^ n2497 ^ 1'b0 ;
  assign n3422 = n691 | n3421 ;
  assign n3423 = n1015 & n1653 ;
  assign n3424 = n3125 ^ n1022 ^ 1'b0 ;
  assign n3425 = n685 & n3424 ;
  assign n3426 = n3425 ^ n907 ^ 1'b0 ;
  assign n3427 = ~n570 & n2822 ;
  assign n3428 = n3098 ^ n2071 ^ 1'b0 ;
  assign n3429 = n1060 & n2842 ;
  assign n3430 = ~n690 & n1966 ;
  assign n3431 = n2122 & n3430 ;
  assign n3432 = n56 & ~n818 ;
  assign n3433 = n609 & n3432 ;
  assign n3434 = n3433 ^ n1057 ^ 1'b0 ;
  assign n3435 = n2513 & n3434 ;
  assign n3436 = n1817 ^ n223 ^ 1'b0 ;
  assign n3437 = n226 & ~n1791 ;
  assign n3438 = n3176 ^ n770 ^ 1'b0 ;
  assign n3439 = n3438 ^ n277 ^ 1'b0 ;
  assign n3440 = n2129 & ~n3439 ;
  assign n3441 = n855 ^ n545 ^ 1'b0 ;
  assign n3442 = ~n2059 & n3441 ;
  assign n3443 = n798 & n3442 ;
  assign n3444 = ~n3420 & n3443 ;
  assign n3445 = n278 & ~n754 ;
  assign n3446 = n3445 ^ n827 ^ 1'b0 ;
  assign n3447 = n1048 ^ n609 ^ n102 ;
  assign n3448 = n3447 ^ n190 ^ 1'b0 ;
  assign n3449 = n364 & n3448 ;
  assign n3450 = n1900 & n2121 ;
  assign n3451 = ~n1810 & n3450 ;
  assign n3452 = n1060 ^ n174 ^ 1'b0 ;
  assign n3453 = n1144 & n3452 ;
  assign n3454 = ~n715 & n3453 ;
  assign n3455 = n3451 | n3454 ;
  assign n3456 = n3449 | n3455 ;
  assign n3457 = ~n1038 & n1965 ;
  assign n3458 = n3423 ^ n2988 ^ 1'b0 ;
  assign n3459 = n87 | n912 ;
  assign n3460 = n3459 ^ n501 ^ 1'b0 ;
  assign n3461 = n184 & n3460 ;
  assign n3462 = n582 ^ n266 ^ 1'b0 ;
  assign n3463 = ~n587 & n1932 ;
  assign n3464 = n3462 & n3463 ;
  assign n3465 = ~n425 & n2186 ;
  assign n3466 = n2438 ^ n170 ^ 1'b0 ;
  assign n3467 = n492 & ~n1315 ;
  assign n3468 = n2438 & n2830 ;
  assign n3469 = n3467 & n3468 ;
  assign n3471 = n156 & n500 ;
  assign n3470 = n406 & n928 ;
  assign n3472 = n3471 ^ n3470 ^ 1'b0 ;
  assign n3473 = n2599 ^ n774 ^ 1'b0 ;
  assign n3474 = n1001 | n1479 ;
  assign n3475 = n2120 | n3474 ;
  assign n3476 = n1587 ^ n841 ^ 1'b0 ;
  assign n3477 = n3476 ^ n1003 ^ 1'b0 ;
  assign n3480 = n873 ^ n495 ^ 1'b0 ;
  assign n3478 = n2941 ^ n1065 ^ 1'b0 ;
  assign n3479 = n86 & n3478 ;
  assign n3481 = n3480 ^ n3479 ^ 1'b0 ;
  assign n3482 = n566 | n867 ;
  assign n3483 = n131 & ~n3482 ;
  assign n3484 = n2046 ^ n58 ^ 1'b0 ;
  assign n3485 = n688 & ~n1588 ;
  assign n3486 = n3485 ^ n2727 ^ 1'b0 ;
  assign n3487 = n3484 & ~n3486 ;
  assign n3488 = n1151 & n3408 ;
  assign n3489 = ~n1663 & n3488 ;
  assign n3490 = n403 | n2017 ;
  assign n3491 = ~n1229 & n1409 ;
  assign n3492 = n3491 ^ n2117 ^ 1'b0 ;
  assign n3493 = ~n1566 & n3492 ;
  assign n3494 = n907 | n1165 ;
  assign n3495 = n3494 ^ n133 ^ 1'b0 ;
  assign n3496 = ~n1078 & n2804 ;
  assign n3497 = n1726 & n3496 ;
  assign n3498 = n2142 & ~n3497 ;
  assign n3499 = n2591 ^ n1358 ^ 1'b0 ;
  assign n3500 = n3499 ^ n2032 ^ 1'b0 ;
  assign n3501 = ( ~n2209 & n2426 ) | ( ~n2209 & n3500 ) | ( n2426 & n3500 ) ;
  assign n3502 = ~n131 & n2205 ;
  assign n3503 = n3502 ^ n929 ^ 1'b0 ;
  assign n3505 = n497 & n1159 ;
  assign n3504 = n3229 ^ n1483 ^ 1'b0 ;
  assign n3506 = n3505 ^ n3504 ^ 1'b0 ;
  assign n3507 = n261 ^ n153 ^ 1'b0 ;
  assign n3508 = n3295 & ~n3507 ;
  assign n3509 = n1637 & n3508 ;
  assign n3510 = n2185 ^ n1113 ^ 1'b0 ;
  assign n3511 = n48 | n3510 ;
  assign n3512 = n3511 ^ n1332 ^ 1'b0 ;
  assign n3513 = n1908 ^ n532 ^ 1'b0 ;
  assign n3514 = n715 ^ n417 ^ 1'b0 ;
  assign n3515 = n1246 & ~n1392 ;
  assign n3516 = n3515 ^ n1445 ^ 1'b0 ;
  assign n3518 = n2196 ^ n128 ^ 1'b0 ;
  assign n3519 = ~n270 & n3518 ;
  assign n3520 = n1416 & n3519 ;
  assign n3517 = n419 & n714 ;
  assign n3521 = n3520 ^ n3517 ^ 1'b0 ;
  assign n3522 = n3521 ^ n1252 ^ 1'b0 ;
  assign n3523 = n1426 ^ n663 ^ 1'b0 ;
  assign n3524 = ~n459 & n1173 ;
  assign n3525 = n1469 & n2060 ;
  assign n3526 = ~n3524 & n3525 ;
  assign n3527 = n3523 & ~n3526 ;
  assign n3528 = n477 & n975 ;
  assign n3529 = n3528 ^ n273 ^ 1'b0 ;
  assign n3530 = n3529 ^ n1771 ^ 1'b0 ;
  assign n3531 = n637 | n962 ;
  assign n3532 = n3530 | n3531 ;
  assign n3533 = x11 | n2768 ;
  assign n3534 = n141 | n3023 ;
  assign n3535 = ~n185 & n1406 ;
  assign n3536 = n3535 ^ n800 ^ 1'b0 ;
  assign n3537 = ~n191 & n3536 ;
  assign n3538 = n302 | n2693 ;
  assign n3539 = n3538 ^ n1191 ^ 1'b0 ;
  assign n3540 = n3539 ^ n3030 ^ n129 ;
  assign n3541 = n1506 ^ n402 ^ 1'b0 ;
  assign n3542 = n1341 & n3541 ;
  assign n3544 = ~n492 & n878 ;
  assign n3545 = n3544 ^ n813 ^ 1'b0 ;
  assign n3543 = n398 & ~n1112 ;
  assign n3546 = n3545 ^ n3543 ^ 1'b0 ;
  assign n3547 = n1902 ^ n364 ^ 1'b0 ;
  assign n3548 = ~n2076 & n3547 ;
  assign n3551 = n472 | n927 ;
  assign n3552 = n750 | n3551 ;
  assign n3553 = n1293 & n3552 ;
  assign n3554 = n3553 ^ n984 ^ 1'b0 ;
  assign n3549 = n616 | n2949 ;
  assign n3550 = n2157 & ~n3549 ;
  assign n3555 = n3554 ^ n3550 ^ 1'b0 ;
  assign n3556 = n863 & ~n3555 ;
  assign n3558 = n310 & ~n1061 ;
  assign n3557 = n348 & ~n3344 ;
  assign n3559 = n3558 ^ n3557 ^ n284 ;
  assign n3560 = n804 ^ n553 ^ 1'b0 ;
  assign n3561 = n3560 ^ n448 ^ 1'b0 ;
  assign n3562 = n2550 ^ n2200 ^ 1'b0 ;
  assign n3563 = ~n2529 & n3562 ;
  assign n3564 = n3561 | n3563 ;
  assign n3565 = n3420 ^ n1912 ^ 1'b0 ;
  assign n3566 = n3116 | n3565 ;
  assign n3567 = n520 | n3566 ;
  assign n3569 = n163 | n764 ;
  assign n3568 = n278 | n1233 ;
  assign n3570 = n3569 ^ n3568 ^ 1'b0 ;
  assign n3571 = n3295 | n3570 ;
  assign n3572 = n325 & n1210 ;
  assign n3573 = n1224 & n3572 ;
  assign n3574 = n3573 ^ n1691 ^ 1'b0 ;
  assign n3575 = n1793 | n1924 ;
  assign n3576 = ~n227 & n3575 ;
  assign n3577 = n963 & n1441 ;
  assign n3578 = ~n404 & n1624 ;
  assign n3579 = n3578 ^ n878 ^ 1'b0 ;
  assign n3580 = n1588 ^ n649 ^ 1'b0 ;
  assign n3581 = n2360 & n2959 ;
  assign n3582 = n859 ^ n412 ^ 1'b0 ;
  assign n3583 = n117 | n3582 ;
  assign n3584 = n582 | n2932 ;
  assign n3585 = x11 & n310 ;
  assign n3586 = ~n106 & n1295 ;
  assign n3587 = n482 & ~n1754 ;
  assign n3588 = n3586 & n3587 ;
  assign n3589 = n3588 ^ n198 ^ 1'b0 ;
  assign n3590 = n2082 & ~n3589 ;
  assign n3591 = ~n457 & n3590 ;
  assign n3592 = n348 & ~n3591 ;
  assign n3593 = n3112 ^ n2418 ^ 1'b0 ;
  assign n3594 = n1001 ^ n415 ^ 1'b0 ;
  assign n3595 = n3594 ^ n904 ^ 1'b0 ;
  assign n3596 = n2065 & ~n3595 ;
  assign n3597 = n652 & n3596 ;
  assign n3598 = n1467 & n2426 ;
  assign n3599 = n161 | n3598 ;
  assign n3600 = ~n346 & n1241 ;
  assign n3602 = n338 | n657 ;
  assign n3601 = n2334 & ~n3150 ;
  assign n3603 = n3602 ^ n3601 ^ n2710 ;
  assign n3604 = n835 & ~n963 ;
  assign n3605 = n758 & ~n3051 ;
  assign n3606 = n3605 ^ n713 ^ 1'b0 ;
  assign n3607 = n342 & ~n941 ;
  assign n3608 = ~n1368 & n3607 ;
  assign n3612 = n539 & ~n3595 ;
  assign n3613 = n3612 ^ n971 ^ 1'b0 ;
  assign n3614 = n3613 ^ n2992 ^ 1'b0 ;
  assign n3609 = n315 & ~n1280 ;
  assign n3610 = n862 ^ n273 ^ 1'b0 ;
  assign n3611 = n3609 | n3610 ;
  assign n3615 = n3614 ^ n3611 ^ 1'b0 ;
  assign n3616 = n3608 | n3615 ;
  assign n3617 = n1965 | n2348 ;
  assign n3619 = n804 & ~n1407 ;
  assign n3620 = n3619 ^ n2043 ^ 1'b0 ;
  assign n3621 = n2415 & n3620 ;
  assign n3618 = n148 & n1426 ;
  assign n3622 = n3621 ^ n3618 ^ 1'b0 ;
  assign n3626 = ~n186 & n306 ;
  assign n3625 = n1961 & ~n2998 ;
  assign n3627 = n3626 ^ n3625 ^ 1'b0 ;
  assign n3628 = n758 ^ n364 ^ 1'b0 ;
  assign n3629 = n119 | n3628 ;
  assign n3630 = n3629 ^ n1745 ^ 1'b0 ;
  assign n3631 = n3627 & ~n3630 ;
  assign n3623 = n2112 & n3077 ;
  assign n3624 = n3623 ^ n161 ^ 1'b0 ;
  assign n3632 = n3631 ^ n3624 ^ n293 ;
  assign n3633 = n1874 & ~n1877 ;
  assign n3634 = n3633 ^ n1219 ^ 1'b0 ;
  assign n3635 = n142 & n3634 ;
  assign n3636 = n3034 & n3103 ;
  assign n3637 = n2144 ^ n1011 ^ 1'b0 ;
  assign n3638 = n1855 ^ n1335 ^ 1'b0 ;
  assign n3639 = n1300 ^ n359 ^ 1'b0 ;
  assign n3640 = n3638 | n3639 ;
  assign n3641 = n1573 & ~n2907 ;
  assign n3642 = n1328 ^ n1237 ^ 1'b0 ;
  assign n3643 = n3642 ^ n55 ^ 1'b0 ;
  assign n3644 = n738 ^ n359 ^ 1'b0 ;
  assign n3645 = ~n53 & n3644 ;
  assign n3646 = n3645 ^ n1083 ^ 1'b0 ;
  assign n3647 = ~n637 & n1519 ;
  assign n3648 = n3647 ^ n3640 ^ 1'b0 ;
  assign n3649 = n594 & ~n1771 ;
  assign n3650 = n271 & n3649 ;
  assign n3651 = n141 & n1073 ;
  assign n3652 = n3651 ^ n1807 ^ 1'b0 ;
  assign n3653 = n417 & ~n3652 ;
  assign n3654 = ~n135 & n3653 ;
  assign n3655 = n3654 ^ n2594 ^ 1'b0 ;
  assign n3656 = n83 & n236 ;
  assign n3657 = n3656 ^ n1368 ^ 1'b0 ;
  assign n3658 = ~n1067 & n3657 ;
  assign n3659 = n3658 ^ n3527 ^ 1'b0 ;
  assign n3660 = n1235 | n1802 ;
  assign n3661 = n1348 | n3660 ;
  assign n3662 = n3661 ^ n2833 ^ 1'b0 ;
  assign n3663 = n1239 ^ n715 ^ 1'b0 ;
  assign n3664 = n1129 | n3663 ;
  assign n3665 = n3662 | n3664 ;
  assign n3666 = n927 ^ n799 ^ 1'b0 ;
  assign n3667 = n3666 ^ n1271 ^ 1'b0 ;
  assign n3668 = n2634 & n3667 ;
  assign n3669 = n1655 & ~n3413 ;
  assign n3670 = n340 & ~n3669 ;
  assign n3671 = n3387 ^ n2822 ^ 1'b0 ;
  assign n3672 = n2065 ^ n52 ^ 1'b0 ;
  assign n3673 = n3672 ^ n1655 ^ 1'b0 ;
  assign n3674 = n3276 | n3673 ;
  assign n3675 = n2131 ^ n1370 ^ 1'b0 ;
  assign n3676 = ~n3674 & n3675 ;
  assign n3677 = n2388 ^ n1263 ^ 1'b0 ;
  assign n3678 = n148 | n3677 ;
  assign n3679 = n663 & n1304 ;
  assign n3680 = n3679 ^ n2360 ^ 1'b0 ;
  assign n3681 = n3059 & n3333 ;
  assign n3682 = n1870 ^ n89 ^ 1'b0 ;
  assign n3683 = n479 | n1392 ;
  assign n3684 = n1203 | n3683 ;
  assign n3685 = n3682 & n3684 ;
  assign n3686 = n3685 ^ n3684 ^ 1'b0 ;
  assign n3687 = n1243 & n3686 ;
  assign n3688 = n108 & n3687 ;
  assign n3689 = n1364 & ~n2593 ;
  assign n3690 = n1920 & n3689 ;
  assign n3691 = x6 & ~n3690 ;
  assign n3692 = ~n1142 & n3691 ;
  assign n3693 = n2534 ^ n741 ^ 1'b0 ;
  assign n3694 = n748 | n3693 ;
  assign n3695 = n1246 & n3694 ;
  assign n3696 = n3692 & n3695 ;
  assign n3697 = n2601 ^ n1525 ^ 1'b0 ;
  assign n3698 = n1210 & n3697 ;
  assign n3699 = n817 & ~n1472 ;
  assign n3700 = n3699 ^ n2905 ^ 1'b0 ;
  assign n3701 = ~n690 & n3700 ;
  assign n3702 = n1235 & n1663 ;
  assign n3703 = n372 | n3462 ;
  assign n3704 = n3703 ^ n2317 ^ 1'b0 ;
  assign n3705 = n1161 & ~n2814 ;
  assign n3706 = n3705 ^ n2011 ^ 1'b0 ;
  assign n3707 = n2162 ^ n835 ^ 1'b0 ;
  assign n3708 = n450 & ~n2872 ;
  assign n3709 = ~n1380 & n1932 ;
  assign n3717 = n68 | n567 ;
  assign n3710 = ( n934 & n2082 ) | ( n934 & ~n2204 ) | ( n2082 & ~n2204 ) ;
  assign n3711 = n175 | n311 ;
  assign n3712 = n2311 | n3711 ;
  assign n3713 = n195 | n3712 ;
  assign n3714 = ~n3710 & n3713 ;
  assign n3715 = n3714 ^ n3385 ^ 1'b0 ;
  assign n3716 = ~n796 & n3715 ;
  assign n3718 = n3717 ^ n3716 ^ 1'b0 ;
  assign n3719 = n2790 ^ n1354 ^ 1'b0 ;
  assign n3720 = ~n789 & n1886 ;
  assign n3721 = ~n2097 & n3720 ;
  assign n3722 = ~n3719 & n3721 ;
  assign n3723 = ~n2633 & n3722 ;
  assign n3724 = ~n3167 & n3723 ;
  assign n3725 = n595 & ~n1421 ;
  assign n3726 = n3725 ^ n1008 ^ 1'b0 ;
  assign n3727 = n3726 ^ n2839 ^ 1'b0 ;
  assign n3728 = n784 ^ n709 ^ 1'b0 ;
  assign n3729 = n1941 & n3728 ;
  assign n3730 = n58 | n2892 ;
  assign n3731 = n3729 & ~n3730 ;
  assign n3732 = ~n1121 & n3731 ;
  assign n3733 = n622 & n3413 ;
  assign n3734 = n3733 ^ n3707 ^ 1'b0 ;
  assign n3735 = n747 ^ n210 ^ 1'b0 ;
  assign n3736 = n3735 ^ n3078 ^ 1'b0 ;
  assign n3737 = n3734 & ~n3736 ;
  assign n3738 = n2824 ^ n2059 ^ 1'b0 ;
  assign n3739 = n104 & n1401 ;
  assign n3740 = n2939 & n3739 ;
  assign n3741 = n3740 ^ n175 ^ 1'b0 ;
  assign n3743 = x2 & n459 ;
  assign n3742 = ~n55 & n2106 ;
  assign n3744 = n3743 ^ n3742 ^ n2307 ;
  assign n3745 = n1502 ^ n515 ^ 1'b0 ;
  assign n3746 = n3640 & n3745 ;
  assign n3747 = n627 & n1469 ;
  assign n3748 = n3747 ^ n3685 ^ 1'b0 ;
  assign n3749 = n477 & n3069 ;
  assign n3750 = n683 | n1069 ;
  assign n3751 = n1683 ^ n191 ^ 1'b0 ;
  assign n3752 = n1236 & ~n3751 ;
  assign n3753 = n1011 ^ n16 ^ 1'b0 ;
  assign n3754 = n1415 & n2939 ;
  assign n3755 = n3754 ^ n2136 ^ 1'b0 ;
  assign n3756 = n501 & n3755 ;
  assign n3757 = n1854 ^ n1572 ^ 1'b0 ;
  assign n3758 = n3756 & ~n3757 ;
  assign n3759 = ~n428 & n850 ;
  assign n3760 = n3759 ^ n688 ^ 1'b0 ;
  assign n3761 = n1081 & n3760 ;
  assign n3762 = n356 & n582 ;
  assign n3763 = ~n870 & n1475 ;
  assign n3764 = n3763 ^ n246 ^ 1'b0 ;
  assign n3765 = n489 ^ n355 ^ n64 ;
  assign n3766 = n3523 & ~n3765 ;
  assign n3767 = n1079 & ~n1344 ;
  assign n3768 = n3767 ^ n1227 ^ 1'b0 ;
  assign n3769 = n2186 & n3768 ;
  assign n3770 = n862 | n1410 ;
  assign n3771 = n1831 | n3770 ;
  assign n3772 = n105 & n2067 ;
  assign n3773 = n3772 ^ n2925 ^ 1'b0 ;
  assign n3774 = n3637 & n3773 ;
  assign n3775 = ~n3771 & n3774 ;
  assign n3776 = n2105 ^ n1670 ^ 1'b0 ;
  assign n3777 = n3776 ^ n1015 ^ 1'b0 ;
  assign n3778 = n3100 ^ x8 ^ 1'b0 ;
  assign n3779 = ( ~n64 & n2367 ) | ( ~n64 & n2401 ) | ( n2367 & n2401 ) ;
  assign n3780 = n2342 ^ n2315 ^ 1'b0 ;
  assign n3781 = n1900 ^ n1106 ^ 1'b0 ;
  assign n3782 = n707 & ~n3173 ;
  assign n3783 = n53 & ~n1370 ;
  assign n3784 = n1268 & ~n3783 ;
  assign n3785 = ~n178 & n1027 ;
  assign n3786 = n2137 & ~n2435 ;
  assign n3787 = n1999 & ~n2270 ;
  assign n3788 = n807 ^ n73 ^ 1'b0 ;
  assign n3789 = n3787 | n3788 ;
  assign n3790 = n896 & n1759 ;
  assign n3791 = n3790 ^ n2931 ^ 1'b0 ;
  assign n3792 = n3755 ^ n356 ^ 1'b0 ;
  assign n3793 = n2514 ^ n2082 ^ 1'b0 ;
  assign n3794 = n2130 & n3793 ;
  assign n3795 = ~n965 & n3794 ;
  assign n3796 = n3795 ^ n310 ^ 1'b0 ;
  assign n3797 = n2079 & n2166 ;
  assign n3798 = n3126 | n3570 ;
  assign n3799 = ~n859 & n2594 ;
  assign n3800 = n159 & ~n3627 ;
  assign n3801 = ~n131 & n519 ;
  assign n3802 = n3801 ^ n2348 ^ 1'b0 ;
  assign n3803 = n149 ^ n68 ^ 1'b0 ;
  assign n3804 = n3378 & n3803 ;
  assign n3805 = ~n330 & n1500 ;
  assign n3806 = n2996 ^ n1254 ^ 1'b0 ;
  assign n3807 = n169 | n2511 ;
  assign n3808 = n3290 ^ n2880 ^ 1'b0 ;
  assign n3809 = n86 & ~n813 ;
  assign n3810 = n3809 ^ n76 ^ 1'b0 ;
  assign n3811 = n324 | n2963 ;
  assign n3812 = n3811 ^ n1250 ^ 1'b0 ;
  assign n3813 = n2500 | n3603 ;
  assign n3814 = n3265 ^ n2063 ^ 1'b0 ;
  assign n3815 = n2137 ^ n1241 ^ 1'b0 ;
  assign n3816 = n1345 & ~n3815 ;
  assign n3817 = ~n372 & n3816 ;
  assign n3818 = n1777 & n2771 ;
  assign n3819 = n2148 ^ n929 ^ 1'b0 ;
  assign n3820 = n1763 & ~n3819 ;
  assign n3821 = n3820 ^ n1191 ^ 1'b0 ;
  assign n3822 = n1205 ^ n277 ^ 1'b0 ;
  assign n3823 = ~n1104 & n3822 ;
  assign n3824 = n2937 ^ n458 ^ 1'b0 ;
  assign n3825 = n3620 & ~n3824 ;
  assign n3826 = n3825 ^ n1828 ^ 1'b0 ;
  assign n3827 = n1714 ^ n235 ^ 1'b0 ;
  assign n3828 = n271 & ~n3827 ;
  assign n3829 = n652 | n3663 ;
  assign n3830 = n1826 | n3829 ;
  assign n3831 = ~n1935 & n3830 ;
  assign n3832 = n3831 ^ n2097 ^ 1'b0 ;
  assign n3833 = n122 & ~n1315 ;
  assign n3834 = n1644 ^ n55 ^ 1'b0 ;
  assign n3835 = n3833 & ~n3834 ;
  assign n3836 = n2573 ^ n641 ^ 1'b0 ;
  assign n3837 = n348 | n1939 ;
  assign n3838 = n584 & ~n3837 ;
  assign n3839 = ~n364 & n3838 ;
  assign n3840 = n534 | n1118 ;
  assign n3841 = n1216 | n3840 ;
  assign n3842 = n246 & n2696 ;
  assign n3843 = ~n28 & n3842 ;
  assign n3844 = ~n135 & n2642 ;
  assign n3845 = n468 & n1630 ;
  assign n3846 = n398 & ~n1001 ;
  assign n3847 = ~n1601 & n3846 ;
  assign n3848 = n2859 & n3847 ;
  assign n3849 = n1252 ^ n1178 ^ 1'b0 ;
  assign n3850 = n3849 ^ n277 ^ 1'b0 ;
  assign n3851 = ~n2096 & n2826 ;
  assign n3852 = n1484 | n3139 ;
  assign n3853 = n375 | n3852 ;
  assign n3854 = n525 | n3853 ;
  assign n3855 = n1268 & ~n2723 ;
  assign n3856 = n3581 | n3855 ;
  assign n3857 = n398 & ~n3788 ;
  assign n3858 = ~n340 & n3857 ;
  assign n3859 = n520 ^ n310 ^ 1'b0 ;
  assign n3860 = n414 & ~n475 ;
  assign n3861 = n3860 ^ n307 ^ 1'b0 ;
  assign n3862 = n3861 ^ n3789 ^ 1'b0 ;
  assign n3863 = ~n212 & n249 ;
  assign n3864 = n1961 & n3863 ;
  assign n3865 = n3864 ^ n2771 ^ 1'b0 ;
  assign n3866 = n350 & n3865 ;
  assign n3867 = n1278 & ~n3008 ;
  assign n3868 = n3867 ^ n340 ^ 1'b0 ;
  assign n3869 = n2433 | n2888 ;
  assign n3870 = n2110 | n3869 ;
  assign n3871 = n635 | n3870 ;
  assign n3872 = n760 & ~n1493 ;
  assign n3873 = n3872 ^ n1072 ^ 1'b0 ;
  assign n3874 = n3873 ^ n97 ^ 1'b0 ;
  assign n3875 = n1040 & ~n2873 ;
  assign n3876 = n1330 & ~n3875 ;
  assign n3877 = ~n1177 & n3876 ;
  assign n3878 = n1304 & n3784 ;
  assign n3879 = ~n55 & n378 ;
  assign n3880 = n3879 ^ n359 ^ 1'b0 ;
  assign n3881 = n2055 | n3208 ;
  assign n3882 = n3880 | n3881 ;
  assign n3883 = n2312 & n2500 ;
  assign n3884 = n3883 ^ n2455 ^ 1'b0 ;
  assign n3885 = ~n3708 & n3884 ;
  assign n3886 = n3104 & ~n3454 ;
  assign n3887 = ~n55 & n2201 ;
  assign n3888 = n3301 & ~n3887 ;
  assign n3889 = n438 ^ n191 ^ 1'b0 ;
  assign n3890 = ~n1793 & n3889 ;
  assign n3891 = n979 & ~n2971 ;
  assign n3892 = n3574 ^ n3169 ^ 1'b0 ;
  assign n3893 = n2366 ^ n336 ^ 1'b0 ;
  assign n3894 = n83 & ~n481 ;
  assign n3895 = n2369 | n3894 ;
  assign n3896 = n3895 ^ n1558 ^ 1'b0 ;
  assign n3897 = n1474 & ~n3179 ;
  assign n3898 = n246 & n3897 ;
  assign n3899 = n3896 & n3898 ;
  assign n3900 = n1080 ^ n1003 ^ 1'b0 ;
  assign n3901 = ~n1193 & n3900 ;
  assign n3902 = n1599 & ~n2455 ;
  assign n3903 = n3902 ^ n2159 ^ 1'b0 ;
  assign n3904 = n3635 & ~n3903 ;
  assign n3905 = ~n3901 & n3904 ;
  assign n3907 = ~n1061 & n1770 ;
  assign n3906 = n535 & ~n624 ;
  assign n3908 = n3907 ^ n3906 ^ 1'b0 ;
  assign n3909 = n1695 & n2476 ;
  assign n3910 = n233 & n587 ;
  assign n3911 = ~n233 & n3910 ;
  assign n3912 = n2493 & ~n3911 ;
  assign n3913 = ~n2493 & n3912 ;
  assign n3914 = n3913 ^ n2539 ^ 1'b0 ;
  assign n3915 = n2535 ^ n443 ^ 1'b0 ;
  assign n3916 = ~n3329 & n3915 ;
  assign n3917 = n1515 | n3346 ;
  assign n3918 = ~n330 & n2830 ;
  assign n3919 = n3917 & n3918 ;
  assign n3920 = n2023 ^ n325 ^ 1'b0 ;
  assign n3921 = n159 & ~n3920 ;
  assign n3922 = n1426 ^ n1255 ^ n536 ;
  assign n3923 = n1355 ^ n491 ^ 1'b0 ;
  assign n3924 = n1412 & n3923 ;
  assign n3925 = n1031 ^ x4 ^ 1'b0 ;
  assign n3926 = n3924 | n3925 ;
  assign n3927 = n3922 & ~n3926 ;
  assign n3928 = n3927 ^ n974 ^ 1'b0 ;
  assign n3929 = n3014 ^ n675 ^ 1'b0 ;
  assign n3930 = ~n2140 & n2155 ;
  assign n3931 = n1165 & n3930 ;
  assign n3932 = n935 | n2031 ;
  assign n3933 = n3932 ^ n3755 ^ 1'b0 ;
  assign n3935 = n987 ^ n122 ^ 1'b0 ;
  assign n3934 = n78 & ~n1598 ;
  assign n3936 = n3935 ^ n3934 ^ 1'b0 ;
  assign n3937 = n576 | n2902 ;
  assign n3938 = n3936 | n3937 ;
  assign n3939 = n86 & n3938 ;
  assign n3940 = n3569 ^ n456 ^ 1'b0 ;
  assign n3941 = n3940 ^ n2144 ^ 1'b0 ;
  assign n3942 = n3160 ^ n1390 ^ 1'b0 ;
  assign n3943 = n945 & n3942 ;
  assign n3944 = n1498 & n3943 ;
  assign n3945 = ~n3583 & n3944 ;
  assign n3946 = n2225 | n2738 ;
  assign n3947 = ( ~n2067 & n3868 ) | ( ~n2067 & n3946 ) | ( n3868 & n3946 ) ;
  assign n3948 = n169 | n592 ;
  assign n3949 = n3948 ^ n3247 ^ 1'b0 ;
  assign n3950 = ~n28 & n2491 ;
  assign n3951 = n16 & ~n330 ;
  assign n3952 = n3950 | n3951 ;
  assign n3953 = x10 | n3952 ;
  assign n3954 = n2562 ^ n1635 ^ 1'b0 ;
  assign n3956 = n1048 | n1118 ;
  assign n3957 = n3956 ^ n1005 ^ 1'b0 ;
  assign n3958 = ~n1082 & n3957 ;
  assign n3959 = n257 & n3958 ;
  assign n3955 = ~n1748 & n2701 ;
  assign n3960 = n3959 ^ n3955 ^ 1'b0 ;
  assign n3961 = ~n2502 & n3960 ;
  assign n3962 = n3961 ^ n1274 ^ 1'b0 ;
  assign n3963 = n713 & n2571 ;
  assign n3964 = n3963 ^ n1194 ^ 1'b0 ;
  assign n3965 = n3789 ^ n1947 ^ 1'b0 ;
  assign n3966 = n2017 & n3697 ;
  assign n3967 = n993 | n2633 ;
  assign n3968 = n3967 ^ n2028 ^ 1'b0 ;
  assign n3969 = n3968 ^ n3339 ^ 1'b0 ;
  assign n3970 = ~n296 & n1273 ;
  assign n3971 = n2410 | n3970 ;
  assign n3972 = n465 | n1693 ;
  assign n3973 = n3929 | n3972 ;
  assign n3974 = n3973 ^ n2378 ^ 1'b0 ;
  assign n3975 = n364 & n1506 ;
  assign n3976 = n3975 ^ n1842 ^ 1'b0 ;
  assign n3977 = n798 & n3976 ;
  assign n3978 = n1931 & n3977 ;
  assign n3979 = n178 & n2155 ;
  assign n3980 = n3979 ^ n2331 ^ 1'b0 ;
  assign n3981 = ( ~n527 & n860 ) | ( ~n527 & n2994 ) | ( n860 & n2994 ) ;
  assign n3982 = n2229 & n3338 ;
  assign n3983 = n70 & n3982 ;
  assign n3984 = n135 & ~n375 ;
  assign n3985 = n3984 ^ n345 ^ 1'b0 ;
  assign n3986 = n1286 & n3985 ;
  assign n3987 = n1898 ^ n1759 ^ 1'b0 ;
  assign n3988 = n629 & ~n3987 ;
  assign n3989 = n3986 & ~n3988 ;
  assign n3990 = ~n1108 & n3989 ;
  assign n3991 = n621 | n3990 ;
  assign n3992 = n3991 ^ n1309 ^ 1'b0 ;
  assign n3993 = n1258 ^ n1216 ^ 1'b0 ;
  assign n3994 = n310 | n3993 ;
  assign n3995 = n3994 ^ n2261 ^ 1'b0 ;
  assign n3996 = n2911 ^ n820 ^ 1'b0 ;
  assign n3997 = ~n1007 & n3996 ;
  assign n3998 = n3995 & n3997 ;
  assign n3999 = n1608 | n1795 ;
  assign n4000 = n837 ^ n249 ^ 1'b0 ;
  assign n4001 = n1742 & n4000 ;
  assign n4002 = n2310 & ~n4001 ;
  assign n4003 = n4002 ^ n2582 ^ 1'b0 ;
  assign n4004 = n1741 ^ n641 ^ 1'b0 ;
  assign n4005 = n443 & ~n4004 ;
  assign n4006 = n2872 & n4005 ;
  assign n4007 = n2167 & ~n4006 ;
  assign n4008 = ~n1825 & n4007 ;
  assign n4009 = n2927 ^ n2601 ^ n595 ;
  assign n4010 = ~n986 & n2639 ;
  assign n4011 = n3345 & n3579 ;
  assign n4012 = n4011 ^ n322 ^ 1'b0 ;
  assign n4013 = n1316 & ~n2467 ;
  assign n4014 = n1313 ^ n855 ^ 1'b0 ;
  assign n4015 = n527 & ~n4014 ;
  assign n4016 = n4013 & ~n4015 ;
  assign n4017 = n1901 & n4016 ;
  assign n4018 = ~n3992 & n4017 ;
  assign n4019 = ~n779 & n1673 ;
  assign n4020 = n2210 & n4019 ;
  assign n4021 = n1633 ^ n1388 ^ 1'b0 ;
  assign n4022 = n704 ^ n517 ^ 1'b0 ;
  assign n4023 = n4022 ^ n1826 ^ 1'b0 ;
  assign n4024 = ~n164 & n3575 ;
  assign n4025 = ( n441 & n1399 ) | ( n441 & n4024 ) | ( n1399 & n4024 ) ;
  assign n4026 = n4025 ^ n3854 ^ n1330 ;
  assign n4027 = n665 ^ n205 ^ 1'b0 ;
  assign n4028 = n3467 | n3851 ;
  assign n4029 = n653 & ~n2910 ;
  assign n4030 = n4029 ^ n2814 ^ 1'b0 ;
  assign n4031 = n3059 & n4030 ;
  assign n4032 = n4031 ^ n1097 ^ 1'b0 ;
  assign n4033 = n4028 | n4032 ;
  assign n4034 = ~n228 & n263 ;
  assign n4035 = n4034 ^ n1786 ^ 1'b0 ;
  assign n4036 = n765 & n4035 ;
  assign n4037 = n4036 ^ n2062 ^ 1'b0 ;
  assign n4038 = n4037 ^ n601 ^ 1'b0 ;
  assign n4039 = ~n357 & n4038 ;
  assign n4040 = n712 ^ n295 ^ 1'b0 ;
  assign n4041 = n3679 & n4040 ;
  assign n4042 = ( n337 & n489 ) | ( n337 & ~n4041 ) | ( n489 & ~n4041 ) ;
  assign n4043 = n1452 & n3882 ;
  assign n4047 = n257 & ~n442 ;
  assign n4048 = ~n86 & n4047 ;
  assign n4044 = n497 & n1232 ;
  assign n4045 = n1845 ^ n1000 ^ 1'b0 ;
  assign n4046 = ~n4044 & n4045 ;
  assign n4049 = n4048 ^ n4046 ^ 1'b0 ;
  assign n4050 = n1944 & ~n3206 ;
  assign n4051 = n4050 ^ n2243 ^ 1'b0 ;
  assign n4052 = n2883 ^ n1518 ^ 1'b0 ;
  assign n4053 = n4052 ^ n1048 ^ 1'b0 ;
  assign n4054 = n468 ^ n228 ^ 1'b0 ;
  assign n4055 = n1328 ^ n69 ^ 1'b0 ;
  assign n4056 = n2792 | n4055 ;
  assign n4057 = n75 & ~n4056 ;
  assign n4058 = n1918 ^ n754 ^ 1'b0 ;
  assign n4059 = n2157 | n4058 ;
  assign n4060 = n3343 ^ n3318 ^ 1'b0 ;
  assign n4061 = n2103 ^ n1075 ^ 1'b0 ;
  assign n4062 = n958 & ~n2645 ;
  assign n4063 = n1320 | n1910 ;
  assign n4064 = n1463 & n4063 ;
  assign n4065 = n4062 & n4064 ;
  assign n4066 = n512 & n4065 ;
  assign n4067 = n2694 ^ n278 ^ 1'b0 ;
  assign n4068 = n4066 & n4067 ;
  assign n4069 = ( n274 & n499 ) | ( n274 & ~n596 ) | ( n499 & ~n596 ) ;
  assign n4070 = n241 & n2720 ;
  assign n4071 = n149 | n3803 ;
  assign n4072 = n4071 ^ n364 ^ 1'b0 ;
  assign n4073 = n2428 ^ n246 ^ 1'b0 ;
  assign n4074 = ~n4072 & n4073 ;
  assign n4075 = n27 & n4074 ;
  assign n4076 = n3622 ^ n1588 ^ n292 ;
  assign n4077 = n1790 ^ n766 ^ 1'b0 ;
  assign n4078 = n4077 ^ n2606 ^ 1'b0 ;
  assign n4079 = n822 ^ n415 ^ x5 ;
  assign n4080 = n191 & ~n1388 ;
  assign n4081 = ~n4079 & n4080 ;
  assign n4082 = n898 | n3516 ;
  assign n4083 = n2360 & n4082 ;
  assign n4084 = n4081 & n4083 ;
  assign n4086 = n1388 | n3258 ;
  assign n4087 = n4086 ^ n261 ^ 1'b0 ;
  assign n4085 = n1467 & ~n4044 ;
  assign n4088 = n4087 ^ n4085 ^ 1'b0 ;
  assign n4089 = n479 ^ n35 ^ 1'b0 ;
  assign n4090 = ~n3940 & n4089 ;
  assign n4091 = n3025 & n4090 ;
  assign n4092 = n3037 ^ n804 ^ 1'b0 ;
  assign n4093 = n2676 ^ n962 ^ 1'b0 ;
  assign n4094 = n2183 & n4093 ;
  assign n4095 = n4094 ^ n777 ^ 1'b0 ;
  assign n4096 = ~n75 & n1396 ;
  assign n4097 = n3617 ^ n2050 ^ n975 ;
  assign n4098 = n1027 ^ n553 ^ 1'b0 ;
  assign n4099 = n2945 | n4098 ;
  assign n4100 = n4099 ^ n3643 ^ 1'b0 ;
  assign n4101 = ~n1179 & n2686 ;
  assign n4102 = n4101 ^ n3360 ^ 1'b0 ;
  assign n4103 = n1029 | n3978 ;
  assign n4104 = n2122 | n4103 ;
  assign n4105 = ~n741 & n3638 ;
  assign n4106 = n753 | n2654 ;
  assign n4107 = n247 & n960 ;
  assign n4108 = n729 & n4107 ;
  assign n4109 = n475 ^ x5 ^ 1'b0 ;
  assign n4110 = ~n1315 & n3685 ;
  assign n4111 = n2155 & n4110 ;
  assign n4114 = ~n338 & n3154 ;
  assign n4112 = n1782 ^ n1513 ^ 1'b0 ;
  assign n4113 = ~n4111 & n4112 ;
  assign n4115 = n4114 ^ n4113 ^ 1'b0 ;
  assign n4116 = n740 & n1300 ;
  assign n4117 = ( n2373 & n2762 ) | ( n2373 & n4116 ) | ( n2762 & n4116 ) ;
  assign n4118 = ~n198 & n3756 ;
  assign n4119 = n986 ^ n859 ^ 1'b0 ;
  assign n4120 = ~n1491 & n4119 ;
  assign n4121 = n3178 ^ n1555 ^ 1'b0 ;
  assign n4122 = ~n2385 & n4121 ;
  assign n4123 = n4122 ^ n2186 ^ 1'b0 ;
  assign n4125 = n144 | n1170 ;
  assign n4126 = n3940 & n4125 ;
  assign n4124 = n1889 | n2575 ;
  assign n4127 = n4126 ^ n4124 ^ 1'b0 ;
  assign n4128 = n975 & ~n1015 ;
  assign n4129 = n2233 & n4128 ;
  assign n4130 = n1234 & ~n4129 ;
  assign n4131 = n924 & n4130 ;
  assign n4132 = n2008 | n4131 ;
  assign n4133 = n512 & n3034 ;
  assign n4134 = n348 & ~n472 ;
  assign n4135 = ~n1048 & n4134 ;
  assign n4136 = ~n75 & n2735 ;
  assign n4137 = n2855 | n4136 ;
  assign n4138 = n4135 | n4137 ;
  assign n4139 = n2945 & ~n4138 ;
  assign n4140 = n1326 ^ n712 ^ 1'b0 ;
  assign n4141 = ~n596 & n2547 ;
  assign n4142 = n596 & n4141 ;
  assign n4143 = n4142 ^ n622 ^ 1'b0 ;
  assign n4144 = n185 & ~n891 ;
  assign n4145 = ~n185 & n4144 ;
  assign n4146 = n1598 | n4145 ;
  assign n4147 = n4143 & ~n4146 ;
  assign n4148 = ~n1896 & n4147 ;
  assign n4149 = n1241 ^ n1203 ^ 1'b0 ;
  assign n4150 = n389 & n4149 ;
  assign n4151 = n4008 ^ n1693 ^ 1'b0 ;
  assign n4152 = n4150 & n4151 ;
  assign n4153 = n1900 & ~n2235 ;
  assign n4154 = n414 ^ n163 ^ 1'b0 ;
  assign n4155 = n3258 & ~n4154 ;
  assign n4156 = n1931 ^ n1133 ^ 1'b0 ;
  assign n4157 = n4155 & ~n4156 ;
  assign n4158 = n4157 ^ n2200 ^ n1060 ;
  assign n4159 = n2512 ^ n234 ^ 1'b0 ;
  assign n4160 = n48 | n4159 ;
  assign n4161 = n844 & ~n4160 ;
  assign n4162 = n515 | n2511 ;
  assign n4163 = n626 & ~n4162 ;
  assign n4164 = n1725 | n4163 ;
  assign n4165 = n4164 ^ n567 ^ 1'b0 ;
  assign n4166 = ~n123 & n161 ;
  assign n4167 = n1739 & n2185 ;
  assign n4168 = n227 | n1781 ;
  assign n4169 = n1396 | n4168 ;
  assign n4170 = n2308 & n4169 ;
  assign n4171 = n576 & n4170 ;
  assign n4172 = n1274 ^ n278 ^ 1'b0 ;
  assign n4173 = n1630 & ~n4172 ;
  assign n4174 = n3991 & n4173 ;
  assign n4175 = n1155 & n2438 ;
  assign n4176 = n621 & n4175 ;
  assign n4177 = n337 & ~n4176 ;
  assign n4178 = n4177 ^ n2979 ^ 1'b0 ;
  assign n4179 = n553 | n915 ;
  assign n4180 = ~n3007 & n4179 ;
  assign n4181 = n4180 ^ n520 ^ 1'b0 ;
  assign n4182 = ~n4178 & n4181 ;
  assign n4183 = n1960 & ~n3960 ;
  assign n4184 = n1295 ^ n788 ^ 1'b0 ;
  assign n4185 = n4183 & ~n4184 ;
  assign n4186 = n1533 & ~n3694 ;
  assign n4187 = ~n2726 & n4186 ;
  assign n4188 = n4187 ^ n2159 ^ 1'b0 ;
  assign n4189 = n4188 ^ n884 ^ 1'b0 ;
  assign n4190 = n1040 & ~n2263 ;
  assign n4191 = n4190 ^ n479 ^ 1'b0 ;
  assign n4192 = ~n2999 & n4191 ;
  assign n4193 = n1096 & ~n1690 ;
  assign n4194 = ~n2011 & n4193 ;
  assign n4195 = n2725 ^ n2110 ^ 1'b0 ;
  assign n4196 = n1243 ^ n1195 ^ 1'b0 ;
  assign n4197 = n2875 ^ n44 ^ 1'b0 ;
  assign n4198 = n2862 & ~n4197 ;
  assign n4199 = n1105 ^ n876 ^ 1'b0 ;
  assign n4200 = n973 & n4199 ;
  assign n4201 = n241 & n4200 ;
  assign n4202 = n3260 & ~n4201 ;
  assign n4203 = n968 ^ n56 ^ 1'b0 ;
  assign n4204 = n4203 ^ n3139 ^ 1'b0 ;
  assign n4205 = n1003 | n4204 ;
  assign n4206 = n4112 | n4205 ;
  assign n4207 = n4206 ^ n3922 ^ n1235 ;
  assign n4208 = n273 & ~n822 ;
  assign n4209 = ~n223 & n4208 ;
  assign n4210 = n914 | n4209 ;
  assign n4211 = n1197 ^ n671 ^ 1'b0 ;
  assign n4212 = n4211 ^ n200 ^ 1'b0 ;
  assign n4213 = n1300 ^ n185 ^ 1'b0 ;
  assign n4214 = ~n1197 & n4213 ;
  assign n4215 = n4214 ^ n509 ^ 1'b0 ;
  assign n4216 = ~n4207 & n4215 ;
  assign n4217 = n578 | n3663 ;
  assign n4218 = n1598 & ~n2943 ;
  assign n4219 = ~n4217 & n4218 ;
  assign n4220 = ~n1881 & n2542 ;
  assign n4221 = n475 & ~n4220 ;
  assign n4222 = n1888 ^ n1082 ^ 1'b0 ;
  assign n4223 = n4222 ^ n1559 ^ 1'b0 ;
  assign n4224 = ~n1423 & n2291 ;
  assign n4225 = n4224 ^ n3297 ^ 1'b0 ;
  assign n4226 = n3311 | n4225 ;
  assign n4227 = n929 | n4226 ;
  assign n4228 = n3114 & ~n4227 ;
  assign n4235 = n2736 ^ n775 ^ 1'b0 ;
  assign n4236 = n293 | n4235 ;
  assign n4229 = n47 & n3003 ;
  assign n4230 = n1070 ^ n827 ^ 1'b0 ;
  assign n4231 = n2316 & ~n4230 ;
  assign n4232 = n4231 ^ n4040 ^ 1'b0 ;
  assign n4233 = ~n4229 & n4232 ;
  assign n4234 = ~n255 & n4233 ;
  assign n4237 = n4236 ^ n4234 ^ 1'b0 ;
  assign n4238 = n1716 & n4237 ;
  assign n4239 = n4238 ^ n185 ^ 1'b0 ;
  assign n4240 = n1770 & ~n2931 ;
  assign n4241 = n273 & n806 ;
  assign n4242 = n4241 ^ n2384 ^ 1'b0 ;
  assign n4243 = n2222 & ~n4242 ;
  assign n4244 = n4243 ^ n178 ^ 1'b0 ;
  assign n4245 = n4240 & n4244 ;
  assign n4246 = ~n3280 & n4245 ;
  assign n4247 = n3484 ^ n1533 ^ n973 ;
  assign n4248 = n1162 ^ n888 ^ 1'b0 ;
  assign n4249 = n4247 & n4248 ;
  assign n4250 = n900 ^ n602 ^ 1'b0 ;
  assign n4251 = n4250 ^ n1660 ^ 1'b0 ;
  assign n4252 = x0 & ~n890 ;
  assign n4253 = ~n1951 & n4252 ;
  assign n4254 = n1202 | n4253 ;
  assign n4255 = ~n164 & n414 ;
  assign n4256 = n385 & n4255 ;
  assign n4257 = ~n294 & n3957 ;
  assign n4258 = n4256 & ~n4257 ;
  assign n4259 = n19 | n4258 ;
  assign n4260 = n4181 ^ n3001 ^ 1'b0 ;
  assign n4261 = n246 & n4260 ;
  assign n4262 = n3228 ^ n194 ^ 1'b0 ;
  assign n4263 = n951 | n4262 ;
  assign n4264 = n1683 ^ n1435 ^ 1'b0 ;
  assign n4265 = n188 & n1463 ;
  assign n4266 = n1315 & n4265 ;
  assign n4267 = n939 & ~n4266 ;
  assign n4268 = n636 | n4267 ;
  assign n4269 = n4217 | n4268 ;
  assign n4270 = n2010 | n2642 ;
  assign n4271 = n4270 ^ n1571 ^ x0 ;
  assign n4272 = ~n652 & n756 ;
  assign n4273 = n4272 ^ n272 ^ 1'b0 ;
  assign n4274 = n4273 ^ n255 ^ 1'b0 ;
  assign n4275 = n4274 ^ n4181 ^ 1'b0 ;
  assign n4276 = n2639 ^ n2400 ^ 1'b0 ;
  assign n4277 = ~n322 & n4276 ;
  assign n4278 = n1638 & n4277 ;
  assign n4279 = n3311 ^ n1710 ^ x1 ;
  assign n4280 = n204 & ~n1948 ;
  assign n4282 = ~n740 & n1822 ;
  assign n4283 = n4282 ^ n1946 ^ 1'b0 ;
  assign n4284 = ~n1914 & n4283 ;
  assign n4281 = n78 & n4215 ;
  assign n4285 = n4284 ^ n4281 ^ 1'b0 ;
  assign n4286 = n1910 & n3377 ;
  assign n4287 = n1406 ^ n798 ^ n178 ;
  assign n4288 = ~n191 & n4287 ;
  assign n4289 = ~n37 & n4288 ;
  assign n4290 = ~n2767 & n4289 ;
  assign n4291 = n4290 ^ n3556 ^ n930 ;
  assign n4292 = ~n1406 & n1418 ;
  assign n4293 = n2517 & ~n3483 ;
  assign n4294 = n1213 & n2093 ;
  assign n4295 = n4294 ^ n144 ^ 1'b0 ;
  assign n4296 = ~n1159 & n2655 ;
  assign n4297 = n498 ^ n354 ^ 1'b0 ;
  assign n4298 = n2303 & n4297 ;
  assign n4299 = n2191 ^ n86 ^ 1'b0 ;
  assign n4300 = n1081 | n3759 ;
  assign n4301 = ~n1162 & n1783 ;
  assign n4302 = n4301 ^ n3033 ^ 1'b0 ;
  assign n4303 = n532 & n4302 ;
  assign n4304 = n1719 ^ n1063 ^ 1'b0 ;
  assign n4305 = n4304 ^ n310 ^ 1'b0 ;
  assign n4306 = n1142 & ~n4305 ;
  assign n4307 = n1080 & n1775 ;
  assign n4308 = n4307 ^ n1054 ^ 1'b0 ;
  assign n4310 = n767 ^ n227 ^ 1'b0 ;
  assign n4311 = n294 & ~n4310 ;
  assign n4312 = n4311 ^ n229 ^ 1'b0 ;
  assign n4309 = n700 & ~n3708 ;
  assign n4313 = n4312 ^ n4309 ^ 1'b0 ;
  assign n4314 = n2157 & n4223 ;
  assign n4315 = n236 ^ n135 ^ 1'b0 ;
  assign n4316 = n4256 ^ n192 ^ 1'b0 ;
  assign n4317 = ~n4315 & n4316 ;
  assign n4318 = n375 & n2597 ;
  assign n4319 = ~n507 & n1155 ;
  assign n4320 = n2684 & ~n3373 ;
  assign n4321 = n842 | n4320 ;
  assign n4322 = n1216 & n2640 ;
  assign n4326 = n102 | n148 ;
  assign n4323 = ~n310 & n2061 ;
  assign n4324 = n4323 ^ n1600 ^ 1'b0 ;
  assign n4325 = n3315 | n4324 ;
  assign n4327 = n4326 ^ n4325 ^ 1'b0 ;
  assign n4328 = ~n4322 & n4327 ;
  assign n4329 = n1898 ^ n879 ^ n390 ;
  assign n4330 = n487 ^ n102 ^ x1 ;
  assign n4331 = n194 & ~n1304 ;
  assign n4332 = n2629 ^ n1929 ^ 1'b0 ;
  assign n4333 = n1795 ^ n1715 ^ 1'b0 ;
  assign n4334 = n50 & n4333 ;
  assign n4335 = n4334 ^ n2058 ^ 1'b0 ;
  assign n4336 = n4332 & n4335 ;
  assign n4337 = ~n4331 & n4336 ;
  assign n4338 = n1482 ^ n644 ^ 1'b0 ;
  assign n4339 = n540 | n4338 ;
  assign n4340 = n4339 ^ n470 ^ 1'b0 ;
  assign n4341 = ( n113 & ~n1015 ) | ( n113 & n4340 ) | ( ~n1015 & n4340 ) ;
  assign n4342 = n3087 | n4341 ;
  assign n4343 = n367 & n1256 ;
  assign n4344 = n4343 ^ n842 ^ 1'b0 ;
  assign n4345 = n4321 & ~n4344 ;
  assign n4346 = n4241 & n4345 ;
  assign n4347 = n2985 ^ n471 ^ 1'b0 ;
  assign n4348 = n800 ^ n590 ^ 1'b0 ;
  assign n4349 = n1626 ^ n405 ^ 1'b0 ;
  assign n4350 = n4349 ^ n2626 ^ 1'b0 ;
  assign n4351 = n4350 ^ n3417 ^ 1'b0 ;
  assign n4352 = n3348 & ~n4351 ;
  assign n4353 = n4352 ^ n512 ^ 1'b0 ;
  assign n4354 = n2348 & n4241 ;
  assign n4355 = n271 & n324 ;
  assign n4356 = ~n4273 & n4355 ;
  assign n4357 = n1899 & n3530 ;
  assign n4358 = n2358 | n2362 ;
  assign n4359 = ~n669 & n4358 ;
  assign n4360 = ~n4357 & n4359 ;
  assign n4361 = n155 | n418 ;
  assign n4362 = n2013 & n2480 ;
  assign n4363 = ~n4361 & n4362 ;
  assign n4364 = n1396 & n2987 ;
  assign n4365 = n880 & n4364 ;
  assign n4366 = n562 ^ n55 ^ 1'b0 ;
  assign n4367 = ~n4365 & n4366 ;
  assign n4368 = ~n1597 & n4367 ;
  assign n4369 = n191 & ~n1283 ;
  assign n4370 = n580 | n850 ;
  assign n4371 = n1366 | n4370 ;
  assign n4372 = n4371 ^ n261 ^ 1'b0 ;
  assign n4373 = n4372 ^ n722 ^ 1'b0 ;
  assign n4374 = n4373 ^ n2388 ^ 1'b0 ;
  assign n4375 = n633 ^ n509 ^ 1'b0 ;
  assign n4376 = n4375 ^ n4299 ^ 1'b0 ;
  assign n4377 = ~n1016 & n4376 ;
  assign n4378 = n879 & n4377 ;
  assign n4379 = n2209 ^ n120 ^ 1'b0 ;
  assign n4380 = n1940 & n3579 ;
  assign n4381 = ~n406 & n4380 ;
  assign n4382 = n299 ^ n129 ^ 1'b0 ;
  assign n4383 = ~n2257 & n4382 ;
  assign n4384 = n552 & ~n1328 ;
  assign n4385 = n4384 ^ n1085 ^ 1'b0 ;
  assign n4386 = n427 & ~n4385 ;
  assign n4387 = ~n272 & n4386 ;
  assign n4388 = n3613 | n4387 ;
  assign n4389 = n3659 & ~n4388 ;
  assign n4390 = n16 & ~n1361 ;
  assign n4391 = ~n604 & n4390 ;
  assign n4392 = ~n1849 & n4391 ;
  assign n4393 = n3859 ^ n2997 ^ 1'b0 ;
  assign n4394 = n2146 & n4393 ;
  assign n4395 = n318 | n3284 ;
  assign n4396 = n1582 | n2991 ;
  assign n4397 = n519 & ~n4285 ;
  assign n4398 = n3467 & n4397 ;
  assign n4399 = n869 | n1001 ;
  assign n4400 = n4399 ^ n2455 ^ 1'b0 ;
  assign n4401 = n1198 & ~n1811 ;
  assign n4402 = n970 & ~n2185 ;
  assign n4403 = n4402 ^ n2985 ^ 1'b0 ;
  assign n4404 = n42 | n3631 ;
  assign n4405 = n190 | n1399 ;
  assign n4406 = n4405 ^ n487 ^ 1'b0 ;
  assign n4407 = n1552 | n1588 ;
  assign n4408 = n595 ^ n169 ^ 1'b0 ;
  assign n4409 = n4407 | n4408 ;
  assign n4410 = n1737 ^ n1001 ^ 1'b0 ;
  assign n4411 = n1409 & n4410 ;
  assign n4412 = n3141 ^ n83 ^ 1'b0 ;
  assign n4413 = ~n583 & n872 ;
  assign n4414 = n4413 ^ n1080 ^ 1'b0 ;
  assign n4415 = n4414 ^ n1944 ^ 1'b0 ;
  assign n4416 = n37 & ~n4415 ;
  assign n4417 = ~n2531 & n4077 ;
  assign n4418 = n4417 ^ n1304 ^ 1'b0 ;
  assign n4419 = n3034 & ~n4418 ;
  assign n4420 = n1137 & n3962 ;
  assign n4421 = n2085 & n2501 ;
  assign n4422 = n1036 & n1254 ;
  assign n4423 = n685 & ~n4422 ;
  assign n4424 = ~n2913 & n4423 ;
  assign n4425 = n43 & ~n744 ;
  assign n4426 = n455 & n4425 ;
  assign n4427 = n767 | n4426 ;
  assign n4428 = n4427 ^ n1726 ^ 1'b0 ;
  assign n4429 = ( ~n2392 & n2472 ) | ( ~n2392 & n4428 ) | ( n2472 & n4428 ) ;
  assign n4430 = n4429 ^ n83 ^ 1'b0 ;
  assign n4431 = n1564 ^ n1138 ^ 1'b0 ;
  assign n4434 = n1901 & ~n3057 ;
  assign n4435 = n4434 ^ n3007 ^ 1'b0 ;
  assign n4432 = n158 ^ n66 ^ 1'b0 ;
  assign n4433 = n43 & n4432 ;
  assign n4436 = n4435 ^ n4433 ^ 1'b0 ;
  assign n4437 = ~n2018 & n3890 ;
  assign n4438 = ~n1751 & n3413 ;
  assign n4439 = n2483 & n4438 ;
  assign n4440 = ~n4437 & n4439 ;
  assign n4441 = n2280 ^ n747 ^ n47 ;
  assign n4442 = n694 & ~n1829 ;
  assign n4443 = n4442 ^ n1825 ^ 1'b0 ;
  assign n4444 = n2221 ^ n702 ^ 1'b0 ;
  assign n4445 = n157 & ~n4444 ;
  assign n4446 = n178 & n4445 ;
  assign n4447 = n1642 & ~n2702 ;
  assign n4448 = n4447 ^ n1067 ^ 1'b0 ;
  assign n4449 = n2425 & n4448 ;
  assign n4450 = ~n302 & n2356 ;
  assign n4451 = ~n2384 & n2542 ;
  assign n4452 = ~n974 & n1345 ;
  assign n4453 = ~n784 & n4452 ;
  assign n4454 = n1286 & ~n4453 ;
  assign n4455 = n4454 ^ n3104 ^ 1'b0 ;
  assign n4456 = n4455 ^ n1354 ^ 1'b0 ;
  assign n4457 = n101 & ~n3095 ;
  assign n4458 = n1143 & n4457 ;
  assign n4459 = n83 & ~n4458 ;
  assign n4460 = ~n4448 & n4459 ;
  assign n4461 = n4460 ^ n1863 ^ 1'b0 ;
  assign n4462 = ~n1325 & n4461 ;
  assign n4463 = n4462 ^ n1165 ^ 1'b0 ;
  assign n4464 = n3611 | n4269 ;
  assign n4465 = n1918 & ~n4464 ;
  assign n4466 = ~n1866 & n2998 ;
  assign n4467 = ~n934 & n2532 ;
  assign n4468 = n4467 ^ n4140 ^ 1'b0 ;
  assign n4469 = n46 & ~n4392 ;
  assign n4470 = n3472 & n4469 ;
  assign n4471 = n2702 & n4470 ;
  assign n4472 = n3648 ^ n75 ^ 1'b0 ;
  assign n4473 = n3458 & n4472 ;
  assign n4474 = n1509 ^ n418 ^ 1'b0 ;
  assign n4477 = n385 | n1404 ;
  assign n4478 = n4024 | n4477 ;
  assign n4475 = n814 ^ n205 ^ 1'b0 ;
  assign n4476 = n1771 | n4475 ;
  assign n4479 = n4478 ^ n4476 ^ 1'b0 ;
  assign n4480 = n566 ^ x8 ^ 1'b0 ;
  assign n4481 = ~n2332 & n4480 ;
  assign n4482 = n246 & n4322 ;
  assign n4483 = n2704 ^ n1664 ^ n793 ;
  assign n4484 = ~n690 & n4483 ;
  assign n4485 = n4484 ^ n838 ^ 1'b0 ;
  assign n4490 = n2633 ^ n1331 ^ 1'b0 ;
  assign n4491 = n302 | n4490 ;
  assign n4486 = n255 | n1225 ;
  assign n4487 = n157 | n4486 ;
  assign n4488 = n4487 ^ n873 ^ 1'b0 ;
  assign n4489 = n764 | n4488 ;
  assign n4492 = n4491 ^ n4489 ^ 1'b0 ;
  assign n4493 = n307 & ~n654 ;
  assign n4494 = n292 & n1192 ;
  assign n4495 = n4493 & n4494 ;
  assign n4496 = n1760 ^ n1550 ^ 1'b0 ;
  assign n4497 = n4495 | n4496 ;
  assign n4498 = n715 | n2073 ;
  assign n4499 = n4498 ^ n350 ^ 1'b0 ;
  assign n4500 = n133 | n989 ;
  assign n4501 = n1859 | n4500 ;
  assign n4502 = n1513 | n4326 ;
  assign n4503 = n4501 | n4502 ;
  assign n4504 = n4503 ^ n3631 ^ 1'b0 ;
  assign n4505 = n364 | n3346 ;
  assign n4506 = n4504 | n4505 ;
  assign n4507 = n624 & ~n794 ;
  assign n4508 = n16 & n4507 ;
  assign n4509 = ~n3679 & n4455 ;
  assign n4510 = n1278 ^ n758 ^ n272 ;
  assign n4511 = n1982 ^ n461 ^ 1'b0 ;
  assign n4512 = ~n2560 & n4511 ;
  assign n4513 = n4510 & n4512 ;
  assign n4514 = n1855 ^ n1528 ^ n36 ;
  assign n4515 = n4284 ^ n1287 ^ 1'b0 ;
  assign n4516 = ~n4514 & n4515 ;
  assign n4517 = n1096 | n3524 ;
  assign n4518 = ~n1562 & n1933 ;
  assign n4519 = n4517 & n4518 ;
  assign n4520 = n1968 & ~n2672 ;
  assign n4521 = n553 & n1465 ;
  assign n4522 = n4451 ^ n290 ^ 1'b0 ;
  assign n4523 = n181 ^ n86 ^ 1'b0 ;
  assign n4524 = n775 & n4523 ;
  assign n4525 = n4524 ^ n1829 ^ 1'b0 ;
  assign n4526 = ~n1960 & n4525 ;
  assign n4527 = n1856 ^ n1104 ^ 1'b0 ;
  assign n4528 = ~n1026 & n4527 ;
  assign n4531 = n350 | n1886 ;
  assign n4529 = n709 & n1686 ;
  assign n4530 = n1900 & n4529 ;
  assign n4532 = n4531 ^ n4530 ^ 1'b0 ;
  assign n4533 = n300 & ~n2439 ;
  assign n4534 = n1257 | n4533 ;
  assign n4535 = n88 | n4534 ;
  assign n4536 = n4535 ^ n3957 ^ 1'b0 ;
  assign n4537 = ~n4532 & n4536 ;
  assign n4538 = n3684 ^ n538 ^ 1'b0 ;
  assign n4539 = n83 & ~n4081 ;
  assign n4540 = n4539 ^ n3771 ^ 1'b0 ;
  assign n4541 = n1963 & ~n3907 ;
  assign n4542 = ~n2406 & n4112 ;
  assign n4543 = n215 & n4542 ;
  assign n4544 = n3164 ^ n1637 ^ 1'b0 ;
  assign n4545 = n471 | n2636 ;
  assign n4546 = n2799 & n4545 ;
  assign n4547 = n1546 & ~n2991 ;
  assign n4548 = n4547 ^ n3300 ^ 1'b0 ;
  assign n4549 = ~n474 & n963 ;
  assign n4550 = n2920 ^ n1185 ^ 1'b0 ;
  assign n4551 = n2610 & n4550 ;
  assign n4552 = n3504 | n3857 ;
  assign n4553 = n30 & ~n705 ;
  assign n4554 = n4553 ^ n2129 ^ 1'b0 ;
  assign n4555 = n536 | n4554 ;
  assign n4556 = n4555 ^ n3256 ^ 1'b0 ;
  assign n4557 = n1243 & n1543 ;
  assign n4562 = x1 & ~n141 ;
  assign n4563 = ~n1504 & n4562 ;
  assign n4564 = ~n1598 & n4563 ;
  assign n4558 = n678 ^ x2 ^ 1'b0 ;
  assign n4559 = n1824 | n4558 ;
  assign n4560 = n1644 & n2576 ;
  assign n4561 = ~n4559 & n4560 ;
  assign n4565 = n4564 ^ n4561 ^ 1'b0 ;
  assign n4566 = ~n3529 & n4197 ;
  assign n4567 = n4566 ^ n2956 ^ 1'b0 ;
  assign n4568 = n1968 ^ n477 ^ 1'b0 ;
  assign n4569 = ~n4404 & n4568 ;
  assign n4570 = n975 | n1133 ;
  assign n4572 = n419 & n767 ;
  assign n4571 = n798 & ~n901 ;
  assign n4573 = n4572 ^ n4571 ^ 1'b0 ;
  assign n4574 = n139 & n1849 ;
  assign n4575 = n1001 & n4574 ;
  assign n4576 = n4253 ^ n1848 ^ 1'b0 ;
  assign n4577 = n278 | n4576 ;
  assign n4578 = n461 & n1900 ;
  assign n4579 = n2648 & ~n4578 ;
  assign n4580 = n4577 & n4579 ;
  assign n4581 = n1203 & n4580 ;
  assign n4582 = n2264 & n4581 ;
  assign n4584 = n3138 | n4414 ;
  assign n4583 = n1316 & n4045 ;
  assign n4585 = n4584 ^ n4583 ^ 1'b0 ;
  assign n4586 = ~n1900 & n2122 ;
  assign n4587 = n549 & ~n4586 ;
  assign n4588 = n2907 & n4587 ;
  assign n4594 = n252 & n510 ;
  assign n4590 = n364 & n2179 ;
  assign n4589 = n384 & n1248 ;
  assign n4591 = n4590 ^ n4589 ^ 1'b0 ;
  assign n4592 = n2406 | n4591 ;
  assign n4593 = n216 | n4592 ;
  assign n4595 = n4594 ^ n4593 ^ 1'b0 ;
  assign n4596 = n4595 ^ x8 ^ 1'b0 ;
  assign n4597 = n3620 & n4596 ;
  assign n4598 = n2353 & ~n4448 ;
  assign n4599 = ~n4597 & n4598 ;
  assign n4600 = ~n3546 & n4599 ;
  assign n4601 = n113 & n323 ;
  assign n4602 = n2534 & n4601 ;
  assign n4603 = n4602 ^ n4485 ^ n4428 ;
  assign n4604 = n3049 & ~n4603 ;
  assign n4605 = ~n724 & n2225 ;
  assign n4606 = n4605 ^ n760 ^ 1'b0 ;
  assign n4607 = n1491 & n4284 ;
  assign n4608 = n4606 | n4607 ;
  assign n4609 = n2999 & ~n4608 ;
  assign n4610 = n272 & n1523 ;
  assign n4611 = n875 & n3694 ;
  assign n4612 = n2437 | n4611 ;
  assign n4613 = n2073 & ~n4612 ;
  assign n4614 = n4613 ^ n621 ^ 1'b0 ;
  assign n4615 = ~n37 & n4614 ;
  assign n4616 = n83 & n4615 ;
  assign n4617 = n3320 & ~n4616 ;
  assign n4618 = n721 & n4617 ;
  assign n4619 = n2040 ^ n846 ^ 1'b0 ;
  assign n4620 = n338 & ~n4304 ;
  assign n4621 = n35 & ~n3642 ;
  assign n4622 = ~n268 & n4621 ;
  assign n4623 = ( n3131 & n4049 ) | ( n3131 & n4622 ) | ( n4049 & n4622 ) ;
  assign n4626 = n122 & n1493 ;
  assign n4624 = n3139 | n3732 ;
  assign n4625 = n4624 ^ n1267 ^ 1'b0 ;
  assign n4627 = n4626 ^ n4625 ^ 1'b0 ;
  assign n4628 = n1358 & n4627 ;
  assign n4629 = n390 ^ n34 ^ 1'b0 ;
  assign n4630 = ~n2426 & n4629 ;
  assign n4631 = n632 & n4630 ;
  assign n4632 = n1613 & n4631 ;
  assign n4633 = n87 & ~n149 ;
  assign n4634 = n4632 & ~n4633 ;
  assign n4635 = ~n487 & n3627 ;
  assign n4636 = n4635 ^ n544 ^ 1'b0 ;
  assign n4637 = x3 & n1477 ;
  assign n4638 = n4637 ^ n52 ^ 1'b0 ;
  assign n4639 = n1329 & n2426 ;
  assign n4640 = n4639 ^ n2342 ^ 1'b0 ;
  assign n4641 = n4253 ^ n462 ^ 1'b0 ;
  assign n4642 = n208 & n4641 ;
  assign n4643 = ~n2478 & n4642 ;
  assign n4644 = n2973 ^ n70 ^ 1'b0 ;
  assign n4645 = n4644 ^ n1260 ^ 1'b0 ;
  assign n4646 = n2333 | n2800 ;
  assign n4647 = n1928 & ~n2665 ;
  assign n4650 = n1608 | n3177 ;
  assign n4648 = x0 | n1513 ;
  assign n4649 = n4648 ^ n1530 ^ 1'b0 ;
  assign n4651 = n4650 ^ n4649 ^ 1'b0 ;
  assign n4652 = n549 & n4651 ;
  assign n4653 = n3777 ^ n101 ^ 1'b0 ;
  assign n4654 = ~n4652 & n4653 ;
  assign n4655 = n2586 | n2991 ;
  assign n4656 = n2103 & n3353 ;
  assign n4657 = ~n1463 & n4656 ;
  assign n4658 = ~n627 & n1447 ;
  assign n4659 = n4658 ^ n931 ^ 1'b0 ;
  assign n4660 = n471 & n602 ;
  assign n4661 = n4660 ^ n458 ^ 1'b0 ;
  assign n4662 = n3364 ^ n1286 ^ 1'b0 ;
  assign n4663 = ~n206 & n2433 ;
  assign n4664 = n4663 ^ n4087 ^ 1'b0 ;
  assign n4665 = n3806 ^ n527 ^ 1'b0 ;
  assign n4666 = n3103 | n4665 ;
  assign n4667 = n4435 ^ n3995 ^ n2591 ;
  assign n4668 = n2378 ^ n984 ^ 1'b0 ;
  assign n4669 = ~n158 & n328 ;
  assign n4670 = n4669 ^ n512 ^ 1'b0 ;
  assign n4671 = ( ~n3356 & n3634 ) | ( ~n3356 & n4670 ) | ( n3634 & n4670 ) ;
  assign n4672 = ~n1061 & n2929 ;
  assign n4673 = n2742 & n4672 ;
  assign n4674 = n3282 ^ n157 ^ 1'b0 ;
  assign n4677 = n1227 ^ n592 ^ 1'b0 ;
  assign n4675 = n2916 | n4577 ;
  assign n4676 = n4675 ^ n290 ^ 1'b0 ;
  assign n4678 = n4677 ^ n4676 ^ 1'b0 ;
  assign n4679 = n4108 | n4678 ;
  assign n4682 = ~n324 & n452 ;
  assign n4683 = n956 & n4682 ;
  assign n4684 = n4683 ^ n1129 ^ 1'b0 ;
  assign n4685 = n2419 & ~n4684 ;
  assign n4686 = n4685 ^ n2385 ^ 1'b0 ;
  assign n4680 = n3692 ^ n694 ^ 1'b0 ;
  assign n4681 = n1010 & ~n4680 ;
  assign n4687 = n4686 ^ n4681 ^ 1'b0 ;
  assign n4689 = n68 & n178 ;
  assign n4688 = n3668 ^ n2595 ^ 1'b0 ;
  assign n4690 = n4689 ^ n4688 ^ 1'b0 ;
  assign n4691 = n430 | n2800 ;
  assign n4692 = n372 & ~n4691 ;
  assign n4693 = n4692 ^ n2172 ^ 1'b0 ;
  assign n4694 = n273 | n4693 ;
  assign n4695 = n3038 ^ n530 ^ 1'b0 ;
  assign n4697 = n1889 ^ n719 ^ 1'b0 ;
  assign n4696 = n2454 ^ n363 ^ 1'b0 ;
  assign n4698 = n4697 ^ n4696 ^ 1'b0 ;
  assign n4699 = n55 | n200 ;
  assign n4700 = n4594 & ~n4699 ;
  assign n4701 = n257 & ~n4668 ;
  assign n4702 = ~n2446 & n3537 ;
  assign n4703 = n4702 ^ n873 ^ 1'b0 ;
  assign n4704 = n2313 | n2418 ;
  assign n4705 = n1367 ^ n813 ^ 1'b0 ;
  assign n4706 = n667 & ~n4705 ;
  assign n4707 = n4054 ^ n768 ^ 1'b0 ;
  assign n4708 = ~n663 & n4707 ;
  assign n4709 = n2065 ^ n1652 ^ 1'b0 ;
  assign n4710 = n1552 | n4709 ;
  assign n4711 = n4710 ^ n309 ^ 1'b0 ;
  assign n4712 = n1902 & ~n4711 ;
  assign n4713 = n1063 & n1255 ;
  assign n4714 = n4713 ^ n2366 ^ 1'b0 ;
  assign n4715 = n37 & n3078 ;
  assign n4716 = n116 | n4715 ;
  assign n4717 = n1684 & n4520 ;
  assign n4718 = n612 & n4717 ;
  assign n4719 = n2027 & ~n2362 ;
  assign n4720 = n4719 ^ n163 ^ 1'b0 ;
  assign n4721 = n827 & n4720 ;
  assign n4722 = n4721 ^ n1686 ^ 1'b0 ;
  assign n4723 = n186 & n769 ;
  assign n4724 = n1601 & n4723 ;
  assign n4725 = n1143 | n1708 ;
  assign n4726 = n2107 | n4725 ;
  assign n4727 = n439 | n1490 ;
  assign n4728 = n2510 | n4727 ;
  assign n4729 = n4728 ^ n1851 ^ 1'b0 ;
  assign n4730 = n1266 ^ n212 ^ 1'b0 ;
  assign n4731 = n4674 | n4730 ;
  assign n4734 = n1001 ^ n530 ^ 1'b0 ;
  assign n4732 = ~n726 & n1491 ;
  assign n4733 = n812 | n4732 ;
  assign n4735 = n4734 ^ n4733 ^ 1'b0 ;
  assign n4736 = n246 & n3830 ;
  assign n4737 = ~n2843 & n4736 ;
  assign n4738 = n4737 ^ n1884 ^ 1'b0 ;
  assign n4739 = n944 & ~n4738 ;
  assign n4740 = n2388 & ~n4739 ;
  assign n4741 = n2604 | n3178 ;
  assign n4742 = n4741 ^ n1475 ^ 1'b0 ;
  assign n4743 = n2085 & ~n4081 ;
  assign n4744 = n161 & ~n200 ;
  assign n4745 = n692 & n4744 ;
  assign n4746 = n880 | n1364 ;
  assign n4747 = n4745 | n4746 ;
  assign n4749 = n168 & n311 ;
  assign n4748 = n193 & ~n1884 ;
  assign n4750 = n4749 ^ n4748 ^ 1'b0 ;
  assign n4751 = ~n2079 & n3833 ;
  assign n4752 = n929 & ~n2835 ;
  assign n4753 = n113 & n2172 ;
  assign n4754 = n1173 & n4753 ;
  assign n4755 = ~n506 & n3442 ;
  assign n4756 = n4755 ^ n1456 ^ 1'b0 ;
  assign n4757 = n564 & n995 ;
  assign n4758 = n4757 ^ n366 ^ 1'b0 ;
  assign n4759 = n2303 & n4758 ;
  assign n4760 = n3001 ^ n1619 ^ 1'b0 ;
  assign n4761 = n1707 ^ n290 ^ 1'b0 ;
  assign n4762 = n644 | n2835 ;
  assign n4763 = n761 | n4762 ;
  assign n4764 = n4763 ^ n4657 ^ 1'b0 ;
  assign n4765 = n2689 ^ n2594 ^ 1'b0 ;
  assign n4766 = n2800 ^ n506 ^ 1'b0 ;
  assign n4767 = n177 & ~n4766 ;
  assign n4768 = n3793 ^ n2079 ^ 1'b0 ;
  assign n4769 = n663 & n4768 ;
  assign n4770 = n4769 ^ n3345 ^ 1'b0 ;
  assign n4771 = n2185 ^ n439 ^ 1'b0 ;
  assign n4772 = n4503 & ~n4771 ;
  assign n4773 = n268 | n616 ;
  assign n4774 = n2446 | n4773 ;
  assign n4775 = n934 & n4774 ;
  assign n4776 = n1063 | n2414 ;
  assign n4777 = n2778 & ~n4523 ;
  assign n4778 = ~n1814 & n3472 ;
  assign n4779 = n330 & ~n2295 ;
  assign n4780 = ~n545 & n4779 ;
  assign n4781 = x1 & n395 ;
  assign n4782 = ( n123 & ~n325 ) | ( n123 & n2027 ) | ( ~n325 & n2027 ) ;
  assign n4783 = ~n284 & n4782 ;
  assign n4784 = n4606 & n4783 ;
  assign n4785 = n1202 & ~n2148 ;
  assign n4786 = n3664 | n4785 ;
  assign n4787 = n4786 ^ n2896 ^ 1'b0 ;
  assign n4788 = ~n1792 & n4495 ;
  assign n4789 = n142 & ~n3894 ;
  assign n4790 = n4789 ^ n356 ^ 1'b0 ;
  assign n4791 = n428 | n4790 ;
  assign n4792 = n578 ^ x1 ^ 1'b0 ;
  assign n4793 = ~n177 & n4792 ;
  assign n4794 = ~n2064 & n4793 ;
  assign n4795 = ~n4791 & n4794 ;
  assign n4796 = n489 & n4795 ;
  assign n4797 = ~n729 & n2469 ;
  assign n4798 = n610 | n4797 ;
  assign n4799 = n4312 ^ n1105 ^ 1'b0 ;
  assign n4800 = ~n2483 & n4799 ;
  assign n4801 = n1471 | n1653 ;
  assign n4802 = n3929 ^ n2920 ^ 1'b0 ;
  assign n4803 = n4801 | n4802 ;
  assign n4804 = ( ~n634 & n2121 ) | ( ~n634 & n3669 ) | ( n2121 & n3669 ) ;
  assign n4805 = n3125 ^ n1216 ^ 1'b0 ;
  assign n4806 = n4805 ^ n2542 ^ 1'b0 ;
  assign n4807 = n2067 & n4806 ;
  assign n4808 = n576 | n4807 ;
  assign n4809 = n4804 & ~n4808 ;
  assign n4810 = n46 & ~n833 ;
  assign n4811 = n4810 ^ n1479 ^ 1'b0 ;
  assign n4812 = n4811 ^ n770 ^ 1'b0 ;
  assign n4813 = n4812 ^ n417 ^ 1'b0 ;
  assign n4814 = n1458 & n2817 ;
  assign n4815 = n2849 ^ n2191 ^ 1'b0 ;
  assign n4816 = x0 & n4815 ;
  assign n4817 = ~n286 & n2348 ;
  assign n4818 = n1342 ^ n55 ^ 1'b0 ;
  assign n4819 = ~n591 & n4818 ;
  assign n4820 = ~n1061 & n4819 ;
  assign n4821 = n2604 & ~n4820 ;
  assign n4822 = n48 & n4821 ;
  assign n4823 = n4822 ^ n348 ^ 1'b0 ;
  assign n4824 = n4698 ^ n2774 ^ 1'b0 ;
  assign n4825 = ~n1072 & n3804 ;
  assign n4826 = n2027 & n4079 ;
  assign n4827 = ~n3693 & n4826 ;
  assign n4835 = n161 | n4225 ;
  assign n4829 = n546 ^ n34 ^ 1'b0 ;
  assign n4830 = n608 | n4829 ;
  assign n4831 = n616 | n4830 ;
  assign n4832 = n4831 ^ n1193 ^ 1'b0 ;
  assign n4828 = ~n469 & n2480 ;
  assign n4833 = n4832 ^ n4828 ^ 1'b0 ;
  assign n4834 = ~n551 & n4833 ;
  assign n4836 = n4835 ^ n4834 ^ 1'b0 ;
  assign n4837 = ~n278 & n630 ;
  assign n4838 = n1048 & n4837 ;
  assign n4839 = n2188 ^ n390 ^ 1'b0 ;
  assign n4840 = ~n4838 & n4839 ;
  assign n4841 = ~n3709 & n4840 ;
  assign n4842 = ~n2107 & n4841 ;
  assign n4843 = n191 | n4507 ;
  assign n4844 = n947 | n1283 ;
  assign n4845 = n517 & ~n1406 ;
  assign n4850 = ~n310 & n513 ;
  assign n4846 = ( n683 & n1075 ) | ( n683 & ~n2295 ) | ( n1075 & ~n2295 ) ;
  assign n4847 = ~n1229 & n2136 ;
  assign n4848 = n1245 & n4847 ;
  assign n4849 = ~n4846 & n4848 ;
  assign n4851 = n4850 ^ n4849 ^ 1'b0 ;
  assign n4852 = n2093 ^ n508 ^ 1'b0 ;
  assign n4853 = n1926 & n4852 ;
  assign n4854 = ~n23 & n2424 ;
  assign n4855 = n4854 ^ n294 ^ 1'b0 ;
  assign n4856 = n4855 ^ n2088 ^ 1'b0 ;
  assign n4857 = n456 | n3702 ;
  assign n4858 = ~n927 & n4857 ;
  assign n4859 = n478 & n4858 ;
  assign n4860 = n3900 ^ n1264 ^ 1'b0 ;
  assign n4861 = n391 | n3392 ;
  assign n4862 = n4860 | n4861 ;
  assign n4863 = n1747 & ~n3509 ;
  assign n4864 = ~n83 & n4863 ;
  assign n4865 = n2889 & ~n4864 ;
  assign n4866 = ~n982 & n3317 ;
  assign n4867 = n4866 ^ n3075 ^ 1'b0 ;
  assign n4868 = n3258 ^ n64 ^ 1'b0 ;
  assign n4869 = n1854 & ~n4868 ;
  assign n4870 = n2254 & n2486 ;
  assign n4871 = n4870 ^ n3649 ^ 1'b0 ;
  assign n4872 = ~n3724 & n4871 ;
  assign n4873 = n4872 ^ n2067 ^ n512 ;
  assign n4874 = n462 & ~n2834 ;
  assign n4875 = ~n1935 & n3853 ;
  assign n4876 = n3431 ^ n2951 ^ 1'b0 ;
  assign n4877 = ~n2150 & n4876 ;
  assign n4878 = n1389 & ~n1569 ;
  assign n4879 = n74 ^ n38 ^ 1'b0 ;
  assign n4880 = n4879 ^ n1774 ^ 1'b0 ;
  assign n4882 = n346 | n599 ;
  assign n4881 = n2289 & n4650 ;
  assign n4883 = n4882 ^ n4881 ^ 1'b0 ;
  assign n4884 = n3249 | n4883 ;
  assign n4885 = n1315 | n4286 ;
  assign n4886 = n3550 ^ n2704 ^ 1'b0 ;
  assign n4887 = ~n632 & n4886 ;
  assign n4888 = n627 & n1373 ;
  assign n4889 = ~n4589 & n4888 ;
  assign n4890 = n97 & n4889 ;
  assign n4891 = n4091 ^ n2128 ^ 1'b0 ;
  assign n4892 = n3348 ^ n2072 ^ 1'b0 ;
  assign n4893 = x11 & n4892 ;
  assign n4895 = n1606 & ~n3638 ;
  assign n4894 = n1863 & ~n4116 ;
  assign n4896 = n4895 ^ n4894 ^ 1'b0 ;
  assign n4897 = n2799 & n4896 ;
  assign n4898 = ~n274 & n3349 ;
  assign n4899 = n590 & ~n685 ;
  assign n4900 = n4856 ^ n982 ^ 1'b0 ;
  assign n4901 = ~n609 & n1169 ;
  assign n4902 = n4901 ^ n3087 ^ 1'b0 ;
  assign n4903 = ~n475 & n4902 ;
  assign n4904 = ( ~n191 & n782 ) | ( ~n191 & n4903 ) | ( n782 & n4903 ) ;
  assign n4905 = ~n1061 & n2408 ;
  assign n4906 = n4905 ^ n456 ^ 1'b0 ;
  assign n4907 = n4906 ^ n2307 ^ 1'b0 ;
  assign n4908 = n210 | n2547 ;
  assign n4909 = ( ~n2714 & n4455 ) | ( ~n2714 & n4908 ) | ( n4455 & n4908 ) ;
  assign n4910 = n2283 ^ n139 ^ 1'b0 ;
  assign n4911 = n2236 & ~n4910 ;
  assign n4912 = x0 & ~n3371 ;
  assign n4913 = n4912 ^ n191 ^ 1'b0 ;
  assign n4914 = n2599 ^ n488 ^ 1'b0 ;
  assign n4915 = n359 | n3822 ;
  assign n4916 = n4914 | n4915 ;
  assign n4917 = n294 & ~n2566 ;
  assign n4918 = n3077 ^ n233 ^ 1'b0 ;
  assign n4919 = n1360 | n4918 ;
  assign n4920 = n4919 ^ n619 ^ 1'b0 ;
  assign n4921 = n1741 & n4920 ;
  assign n4922 = n1521 ^ n1108 ^ 1'b0 ;
  assign n4923 = n1303 | n4922 ;
  assign n4924 = ~n613 & n767 ;
  assign n4925 = ~n2107 & n4639 ;
  assign n4926 = n3928 & ~n4925 ;
  assign n4927 = n1676 | n3109 ;
  assign n4928 = n520 | n3759 ;
  assign n4929 = n4927 & ~n4928 ;
  assign n4930 = n4024 ^ n165 ^ 1'b0 ;
  assign n4931 = n4930 ^ n1876 ^ 1'b0 ;
  assign n4932 = ~n452 & n1384 ;
  assign n4933 = n4932 ^ n1363 ^ 1'b0 ;
  assign n4934 = n1057 ^ n144 ^ 1'b0 ;
  assign n4935 = ~n293 & n2664 ;
  assign n4936 = n4934 & n4935 ;
  assign n4937 = n290 | n1280 ;
  assign n4938 = n4937 ^ n128 ^ 1'b0 ;
  assign n4939 = n1368 ^ n843 ^ 1'b0 ;
  assign n4940 = n4939 ^ n2185 ^ 1'b0 ;
  assign n4941 = n3991 | n4940 ;
  assign n4942 = n4941 ^ n4264 ^ 1'b0 ;
  assign n4943 = ~n977 & n1702 ;
  assign n4946 = n2458 & n2506 ;
  assign n4944 = ~n64 & n601 ;
  assign n4945 = n4482 & ~n4944 ;
  assign n4947 = n4946 ^ n4945 ^ 1'b0 ;
  assign n4948 = n3789 ^ n68 ^ 1'b0 ;
  assign n4949 = ~n963 & n4948 ;
  assign n4950 = n4949 ^ n461 ^ 1'b0 ;
  assign n4951 = n517 & ~n4950 ;
  assign n4952 = ( n105 & ~n984 ) | ( n105 & n2768 ) | ( ~n984 & n2768 ) ;
  assign n4953 = n4952 ^ n3688 ^ 1'b0 ;
  assign n4954 = n2264 & ~n4953 ;
  assign n4955 = ( n2690 & n3337 ) | ( n2690 & ~n4954 ) | ( n3337 & ~n4954 ) ;
  assign n4956 = n1555 ^ n60 ^ 1'b0 ;
  assign n4961 = n483 & n1040 ;
  assign n4962 = n137 & n4961 ;
  assign n4963 = ~n1096 & n4962 ;
  assign n4957 = n557 & n641 ;
  assign n4958 = ~n1286 & n4957 ;
  assign n4959 = n1795 ^ n1048 ^ 1'b0 ;
  assign n4960 = n4958 | n4959 ;
  assign n4964 = n4963 ^ n4960 ^ 1'b0 ;
  assign n4965 = n1044 | n4964 ;
  assign n4966 = ( ~n832 & n1129 ) | ( ~n832 & n3658 ) | ( n1129 & n3658 ) ;
  assign n4967 = n2450 & ~n4966 ;
  assign n4968 = n2645 & n2682 ;
  assign n4969 = n571 & ~n4968 ;
  assign n4970 = n3699 ^ n837 ^ 1'b0 ;
  assign n4971 = n4970 ^ n915 ^ 1'b0 ;
  assign n4972 = ~n327 & n4971 ;
  assign n4973 = n883 & ~n3887 ;
  assign n4974 = n2465 & n4973 ;
  assign n4975 = n1713 & ~n2385 ;
  assign n4976 = n270 & n4975 ;
  assign n4977 = n3602 ^ n3575 ^ 1'b0 ;
  assign n4978 = ~n1250 & n1364 ;
  assign n4979 = n1545 & n4978 ;
  assign n4980 = n1277 & n1763 ;
  assign n4981 = n4980 ^ n73 ^ 1'b0 ;
  assign n4982 = n1447 | n4981 ;
  assign n4983 = n4982 ^ n2311 ^ 1'b0 ;
  assign n4984 = n2291 | n4983 ;
  assign n4985 = n4979 | n4984 ;
  assign n4986 = n4985 ^ n3964 ^ 1'b0 ;
  assign n4987 = n3219 ^ n330 ^ 1'b0 ;
  assign n4988 = n2985 | n4987 ;
  assign n4989 = n315 & ~n1322 ;
  assign n4990 = ~n638 & n4989 ;
  assign n4991 = n4813 & ~n4990 ;
  assign n4992 = n1463 | n2116 ;
  assign n4993 = n2410 & ~n4992 ;
  assign n4994 = n1154 | n4161 ;
  assign n4995 = n4812 | n4994 ;
  assign n4996 = n3466 ^ n995 ^ 1'b0 ;
  assign n4997 = n1385 & n3443 ;
  assign n4998 = n4997 ^ n296 ^ 1'b0 ;
  assign n4999 = n1381 & ~n3624 ;
  assign n5000 = n436 & n4999 ;
  assign n5001 = ~n1712 & n1715 ;
  assign n5002 = n5001 ^ n190 ^ 1'b0 ;
  assign n5003 = n356 & ~n5002 ;
  assign n5004 = ~n1174 & n5003 ;
  assign n5005 = ~n1842 & n2092 ;
  assign n5006 = n346 & ~n1662 ;
  assign n5007 = n1031 & n5006 ;
  assign n5008 = ~n848 & n5007 ;
  assign n5009 = n567 & n2203 ;
  assign n5010 = n5009 ^ n481 ^ 1'b0 ;
  assign n5011 = n2726 | n5010 ;
  assign n5012 = n3475 ^ n1011 ^ n241 ;
  assign n5013 = n5012 ^ n249 ^ 1'b0 ;
  assign n5014 = n2604 | n4392 ;
  assign n5015 = n898 ^ n66 ^ 1'b0 ;
  assign n5016 = ~n1626 & n2170 ;
  assign n5017 = x1 | n5016 ;
  assign n5018 = n257 | n5017 ;
  assign n5019 = ~n5015 & n5018 ;
  assign n5020 = n5014 & n5019 ;
  assign n5021 = ~n66 & n1810 ;
  assign n5022 = ~n3277 & n5021 ;
  assign n5023 = n5020 & n5022 ;
  assign n5024 = n414 | n2257 ;
  assign n5025 = n533 & n5024 ;
  assign n5026 = ~n43 & n2218 ;
  assign n5027 = n2917 ^ n942 ^ 1'b0 ;
  assign n5028 = n1048 & ~n5027 ;
  assign n5029 = n4392 ^ n2029 ^ 1'b0 ;
  assign n5030 = ~x2 & n5029 ;
  assign n5031 = n2682 ^ n2249 ^ 1'b0 ;
  assign n5032 = n1609 & n1891 ;
  assign n5033 = n532 & ~n1097 ;
  assign n5034 = n2252 & n5033 ;
  assign n5035 = n907 | n2431 ;
  assign n5036 = n2431 & ~n5035 ;
  assign n5037 = n1097 | n5036 ;
  assign n5038 = n5036 & ~n5037 ;
  assign n5039 = ~n117 & n5038 ;
  assign n5040 = n568 & ~n2642 ;
  assign n5041 = ( ~n142 & n657 ) | ( ~n142 & n2020 ) | ( n657 & n2020 ) ;
  assign n5042 = n5040 & ~n5041 ;
  assign n5043 = n5042 ^ n3597 ^ 1'b0 ;
  assign n5044 = n614 | n1262 ;
  assign n5045 = n1495 | n5044 ;
  assign n5046 = n1875 | n5045 ;
  assign n5047 = n694 ^ n581 ^ 1'b0 ;
  assign n5048 = n2159 & ~n5047 ;
  assign n5049 = n19 | n2106 ;
  assign n5050 = n5048 & n5049 ;
  assign n5051 = ~n2512 & n3762 ;
  assign n5052 = n919 ^ n68 ^ 1'b0 ;
  assign n5053 = ~n832 & n5052 ;
  assign n5054 = n3059 ^ n1314 ^ 1'b0 ;
  assign n5055 = ~n1674 & n5054 ;
  assign n5056 = ~n1233 & n5055 ;
  assign n5057 = ~n1361 & n4850 ;
  assign n5058 = n4287 & ~n5057 ;
  assign n5059 = n974 & n5058 ;
  assign n5060 = n1931 ^ n666 ^ 1'b0 ;
  assign n5065 = x1 & ~n462 ;
  assign n5061 = n2058 & ~n2736 ;
  assign n5062 = n3969 & n5061 ;
  assign n5063 = n5062 ^ n3899 ^ 1'b0 ;
  assign n5064 = n1396 & n5063 ;
  assign n5066 = n5065 ^ n5064 ^ n1034 ;
  assign n5067 = ~n164 & n1078 ;
  assign n5068 = n3385 ^ x1 ^ 1'b0 ;
  assign n5069 = n619 & n976 ;
  assign n5070 = n5069 ^ n101 ^ 1'b0 ;
  assign n5071 = n5070 ^ n4889 ^ 1'b0 ;
  assign n5072 = ~n1181 & n5071 ;
  assign n5073 = ~n2281 & n5072 ;
  assign n5074 = n5073 ^ n1186 ^ 1'b0 ;
  assign n5075 = ~n1078 & n3682 ;
  assign n5076 = n1165 & n5075 ;
  assign n5077 = ~n515 & n1345 ;
  assign n5078 = n5077 ^ n1106 ^ 1'b0 ;
  assign n5083 = n1462 ^ n294 ^ 1'b0 ;
  assign n5079 = n1470 ^ n75 ^ 1'b0 ;
  assign n5080 = ~n701 & n5079 ;
  assign n5081 = n4636 ^ n363 ^ 1'b0 ;
  assign n5082 = n5080 & ~n5081 ;
  assign n5084 = n5083 ^ n5082 ^ 1'b0 ;
  assign n5085 = n1019 ^ n293 ^ 1'b0 ;
  assign n5086 = n799 & ~n5085 ;
  assign n5087 = ~n2027 & n5086 ;
  assign n5088 = ~n353 & n788 ;
  assign n5089 = n5088 ^ n905 ^ 1'b0 ;
  assign n5090 = n2444 & n3855 ;
  assign n5091 = n2556 & n5090 ;
  assign n5092 = n5091 ^ n322 ^ 1'b0 ;
  assign n5093 = n1036 | n5092 ;
  assign n5094 = n5089 | n5093 ;
  assign n5095 = n5087 | n5094 ;
  assign n5096 = n1741 & n2577 ;
  assign n5097 = n1716 ^ n1072 ^ 1'b0 ;
  assign n5098 = n2463 ^ n1285 ^ 1'b0 ;
  assign n5099 = n5097 & n5098 ;
  assign n5100 = n598 & n5099 ;
  assign n5101 = ~n5096 & n5100 ;
  assign n5102 = ~n2519 & n4951 ;
  assign n5103 = n2341 & n3143 ;
  assign n5104 = n427 & ~n4906 ;
  assign n5105 = n2068 & n2225 ;
  assign n5106 = n5105 ^ n4331 ^ 1'b0 ;
  assign n5107 = ~n3593 & n3752 ;
  assign n5108 = n5107 ^ n3054 ^ 1'b0 ;
  assign n5109 = ~n2477 & n2681 ;
  assign n5110 = n5108 & n5109 ;
  assign n5112 = n1795 ^ n270 ^ 1'b0 ;
  assign n5113 = n5112 ^ n4483 ^ 1'b0 ;
  assign n5114 = ~n2426 & n5113 ;
  assign n5115 = n5114 ^ n1205 ^ 1'b0 ;
  assign n5111 = n475 | n2947 ;
  assign n5116 = n5115 ^ n5111 ^ 1'b0 ;
  assign n5117 = ~n4320 & n4931 ;
  assign n5118 = n3231 & n5117 ;
  assign n5119 = n216 & n4540 ;
  assign n5120 = n713 | n4421 ;
  assign n5121 = n3757 & ~n5120 ;
  assign n5122 = n3993 ^ n1212 ^ 1'b0 ;
  assign n5123 = ( n2155 & n4582 ) | ( n2155 & n5122 ) | ( n4582 & n5122 ) ;
  assign n5124 = n506 & n3770 ;
  assign n5125 = n5124 ^ n2452 ^ 1'b0 ;
  assign n5126 = n3548 & n4701 ;
  assign n5127 = n461 & ~n4488 ;
  assign n5128 = n524 | n2148 ;
  assign n5129 = n3632 | n4594 ;
  assign n5130 = n66 | n5129 ;
  assign n5131 = n475 & ~n2424 ;
  assign n5132 = n5131 ^ n4565 ^ 1'b0 ;
  assign n5133 = n1688 | n5132 ;
  assign n5134 = n1081 & n3953 ;
  assign n5135 = n244 ^ n37 ^ 1'b0 ;
  assign n5136 = n2566 | n4077 ;
  assign n5137 = n3047 & ~n3520 ;
  assign n5138 = n1501 & n5137 ;
  assign n5139 = n2481 & ~n3444 ;
  assign n5140 = n5139 ^ n1739 ^ 1'b0 ;
  assign n5141 = n2567 & ~n3202 ;
  assign n5142 = n3939 & ~n4159 ;
  assign n5143 = n4590 ^ n2542 ^ 1'b0 ;
  assign n5144 = n619 & ~n1161 ;
  assign n5145 = n5144 ^ n942 ^ 1'b0 ;
  assign n5146 = n2741 & ~n3868 ;
  assign n5147 = n2417 | n2757 ;
  assign n5148 = n5147 ^ n1344 ^ 1'b0 ;
  assign n5149 = n5148 ^ n283 ^ 1'b0 ;
  assign n5150 = n1598 & ~n1793 ;
  assign n5151 = n5150 ^ n252 ^ 1'b0 ;
  assign n5152 = n1527 & n5151 ;
  assign n5153 = n497 & n3050 ;
  assign n5154 = n5153 ^ n4938 ^ 1'b0 ;
  assign n5155 = n1681 & ~n5053 ;
  assign n5156 = n2773 ^ n1900 ^ 1'b0 ;
  assign n5161 = n4772 ^ n3570 ^ 1'b0 ;
  assign n5157 = n84 & n3788 ;
  assign n5158 = ~n507 & n5157 ;
  assign n5159 = n772 | n5158 ;
  assign n5160 = n2436 & ~n5159 ;
  assign n5162 = n5161 ^ n5160 ^ 1'b0 ;
  assign n5163 = ~n3109 & n3363 ;
  assign n5164 = ~n4350 & n5163 ;
  assign n5165 = ( n274 & n734 ) | ( n274 & ~n3663 ) | ( n734 & ~n3663 ) ;
  assign n5166 = n2704 & ~n2834 ;
  assign n5167 = n5165 & n5166 ;
  assign n5168 = n681 | n2941 ;
  assign n5169 = n5168 ^ n546 ^ 1'b0 ;
  assign n5170 = n914 | n5169 ;
  assign n5171 = n1309 | n5170 ;
  assign n5172 = n5171 ^ n3614 ^ 1'b0 ;
  assign n5173 = n3793 ^ n506 ^ 1'b0 ;
  assign n5174 = ~n5122 & n5173 ;
  assign n5175 = n1745 & n2017 ;
  assign n5176 = ~x11 & n5175 ;
  assign n5177 = n3056 ^ n1774 ^ 1'b0 ;
  assign n5178 = n4851 & ~n5177 ;
  assign n5179 = n799 | n5095 ;
  assign n5180 = n1685 ^ n1283 ^ 1'b0 ;
  assign n5181 = n5180 ^ n3830 ^ 1'b0 ;
  assign n5182 = ~n1360 & n5181 ;
  assign n5183 = ~n757 & n5182 ;
  assign n5184 = n348 & ~n5078 ;
  assign n5185 = n3717 & n5184 ;
  assign n5186 = n715 & ~n3499 ;
  assign n5187 = ~n3340 & n5186 ;
  assign n5188 = n5187 ^ n3917 ^ 1'b0 ;
  assign n5189 = n5124 & n5188 ;
  assign n5190 = n2315 ^ n1105 ^ 1'b0 ;
  assign n5191 = n3003 | n5190 ;
  assign n5192 = n5189 | n5191 ;
  assign n5193 = n642 & ~n958 ;
  assign n5194 = n226 & ~n5193 ;
  assign n5195 = n157 & ~n472 ;
  assign n5196 = n5195 ^ n1934 ^ 1'b0 ;
  assign n5197 = n5196 ^ n1555 ^ 1'b0 ;
  assign n5198 = n799 & ~n5197 ;
  assign n5199 = n1198 & n5198 ;
  assign n5200 = ~n163 & n532 ;
  assign n5201 = n243 | n3374 ;
  assign n5202 = n1361 | n5201 ;
  assign n5203 = n5202 ^ n323 ^ 1'b0 ;
  assign n5204 = n5200 & ~n5203 ;
  assign n5205 = n2565 & ~n3126 ;
  assign n5206 = n414 ^ n191 ^ 1'b0 ;
  assign n5207 = n2055 | n5206 ;
  assign n5208 = ~n5205 & n5207 ;
  assign n5209 = n3750 ^ n1984 ^ 1'b0 ;
  assign n5210 = n459 & n1786 ;
  assign n5211 = n3803 ^ n3175 ^ 1'b0 ;
  assign n5212 = n5211 ^ n246 ^ 1'b0 ;
  assign n5213 = n4848 & n4964 ;
  assign n5214 = ~n4228 & n5213 ;
  assign n5215 = n691 ^ n161 ^ 1'b0 ;
  assign n5216 = ~n280 & n1411 ;
  assign n5217 = ~n2246 & n5216 ;
  assign n5218 = n1631 ^ n1138 ^ 1'b0 ;
  assign n5219 = n3329 ^ n2311 ^ 1'b0 ;
  assign n5220 = n311 ^ n40 ^ 1'b0 ;
  assign n5221 = x3 & n5220 ;
  assign n5222 = n1394 & ~n5221 ;
  assign n5223 = n2941 ^ n381 ^ 1'b0 ;
  assign n5224 = n4189 & ~n5223 ;
  assign n5225 = ~n5222 & n5224 ;
  assign n5226 = n281 & ~n2104 ;
  assign n5228 = ~n3649 & n4329 ;
  assign n5227 = n364 | n2018 ;
  assign n5229 = n5228 ^ n5227 ^ 1'b0 ;
  assign n5230 = ~n1889 & n5229 ;
  assign n5231 = n5230 ^ n2693 ^ 1'b0 ;
  assign n5232 = n507 & ~n1715 ;
  assign n5233 = n164 | n3839 ;
  assign n5234 = n1081 | n5233 ;
  assign n5235 = ~n785 & n4037 ;
  assign n5236 = n2665 ^ n2021 ^ 1'b0 ;
  assign n5237 = n2849 | n5236 ;
  assign n5238 = ~n1725 & n5180 ;
  assign n5239 = ( n2690 & n3223 ) | ( n2690 & n3561 ) | ( n3223 & n3561 ) ;
  assign n5240 = n308 | n4236 ;
  assign n5241 = n5240 ^ n1487 ^ 1'b0 ;
  assign n5242 = n313 | n4287 ;
  assign n5243 = ~n2945 & n3846 ;
  assign n5244 = ~n5242 & n5243 ;
  assign n5245 = n1070 ^ n235 ^ 1'b0 ;
  assign n5246 = n5245 ^ n2742 ^ 1'b0 ;
  assign n5247 = n5244 | n5246 ;
  assign n5248 = n4451 ^ n3940 ^ 1'b0 ;
  assign n5249 = n670 ^ n55 ^ 1'b0 ;
  assign n5250 = n108 | n5249 ;
  assign n5251 = n1693 | n5250 ;
  assign n5252 = ~n2885 & n5251 ;
  assign n5253 = ~n765 & n1255 ;
  assign n5254 = n5253 ^ n865 ^ 1'b0 ;
  assign n5255 = n1547 ^ n1192 ^ 1'b0 ;
  assign n5256 = n5254 & ~n5255 ;
  assign n5257 = n1685 & n3739 ;
  assign n5258 = ~n3088 & n5257 ;
  assign n5260 = ~n741 & n1109 ;
  assign n5261 = ~n1430 & n5260 ;
  assign n5262 = ~n375 & n5261 ;
  assign n5263 = ~n507 & n5262 ;
  assign n5259 = n679 & ~n2220 ;
  assign n5264 = n5263 ^ n5259 ^ 1'b0 ;
  assign n5265 = n2604 & n5264 ;
  assign n5266 = n3108 & n3297 ;
  assign n5267 = ~n79 & n5266 ;
  assign n5268 = n1342 | n2564 ;
  assign n5269 = n5268 ^ n19 ^ 1'b0 ;
  assign n5270 = n3571 ^ n2167 ^ 1'b0 ;
  assign n5271 = n3946 | n4498 ;
  assign n5272 = ~n1845 & n2061 ;
  assign n5273 = ~n2694 & n5272 ;
  assign n5274 = n5133 | n5273 ;
  assign n5275 = n5271 | n5274 ;
  assign n5276 = n4034 ^ n159 ^ 1'b0 ;
  assign n5277 = n4889 | n5276 ;
  assign n5278 = ~n1463 & n2245 ;
  assign n5279 = n4053 ^ n2321 ^ 1'b0 ;
  assign n5280 = n107 & ~n5279 ;
  assign n5281 = n345 ^ n330 ^ 1'b0 ;
  assign n5282 = n5281 ^ n1349 ^ 1'b0 ;
  assign n5283 = n4582 ^ n1054 ^ 1'b0 ;
  assign n5284 = n205 & n2155 ;
  assign n5285 = ~n832 & n1465 ;
  assign n5286 = ~n1546 & n5285 ;
  assign n5287 = n5286 ^ n252 ^ 1'b0 ;
  assign n5288 = n42 & ~n2435 ;
  assign n5289 = n5288 ^ n1174 ^ 1'b0 ;
  assign n5290 = n1662 & ~n4892 ;
  assign n5291 = n1300 & n3353 ;
  assign n5292 = n1409 & n5291 ;
  assign n5293 = n2460 & n5292 ;
  assign n5294 = n2577 & ~n3138 ;
  assign n5295 = n2818 ^ n520 ^ 1'b0 ;
  assign n5296 = n2587 & ~n4497 ;
  assign n5297 = n5296 ^ n1025 ^ 1'b0 ;
  assign n5298 = n1246 & n1704 ;
  assign n5299 = n5298 ^ n2932 ^ 1'b0 ;
  assign n5300 = n55 | n5299 ;
  assign n5301 = n2542 | n5300 ;
  assign n5302 = n5301 ^ n827 ^ 1'b0 ;
  assign n5308 = ~n1227 & n1790 ;
  assign n5303 = n250 & n2882 ;
  assign n5304 = n5303 ^ n1352 ^ 1'b0 ;
  assign n5305 = n5304 ^ n1961 ^ 1'b0 ;
  assign n5306 = n2584 & ~n5305 ;
  assign n5307 = ~n117 & n5306 ;
  assign n5309 = n5308 ^ n5307 ^ 1'b0 ;
  assign n5310 = ~n307 & n3690 ;
  assign n5311 = ~n663 & n1394 ;
  assign n5312 = n5310 & n5311 ;
  assign n5314 = n2684 ^ n2597 ^ 1'b0 ;
  assign n5313 = n3055 ^ n1549 ^ 1'b0 ;
  assign n5315 = n5314 ^ n5313 ^ 1'b0 ;
  assign n5316 = n2144 & ~n5315 ;
  assign n5317 = ( n850 & n3126 ) | ( n850 & n3917 ) | ( n3126 & n3917 ) ;
  assign n5318 = n4111 | n5317 ;
  assign n5319 = n5318 ^ n3177 ^ 1'b0 ;
  assign n5320 = n318 | n1162 ;
  assign n5321 = n5320 ^ n4536 ^ 1'b0 ;
  assign n5322 = n489 & n2994 ;
  assign n5323 = ~n307 & n5322 ;
  assign n5324 = n216 & n3366 ;
  assign n5325 = n632 ^ n367 ^ 1'b0 ;
  assign n5326 = n3254 ^ n1887 ^ 1'b0 ;
  assign n5327 = n5326 ^ n520 ^ 1'b0 ;
  assign n5328 = n738 & n2888 ;
  assign n5329 = n3835 & ~n4689 ;
  assign n5330 = n2187 & n5329 ;
  assign n5331 = n5156 ^ n1860 ^ 1'b0 ;
  assign n5332 = n2988 ^ n1671 ^ 1'b0 ;
  assign n5333 = n1264 ^ n624 ^ 1'b0 ;
  assign n5334 = ( n1430 & ~n1856 ) | ( n1430 & n5333 ) | ( ~n1856 & n5333 ) ;
  assign n5335 = n1198 ^ n497 ^ 1'b0 ;
  assign n5336 = n1471 & ~n2692 ;
  assign n5337 = x6 & n1644 ;
  assign n5338 = n5337 ^ n856 ^ 1'b0 ;
  assign n5339 = n5338 ^ n787 ^ 1'b0 ;
  assign n5340 = n2831 & ~n5339 ;
  assign n5342 = n1291 ^ n715 ^ 1'b0 ;
  assign n5341 = ~n1884 & n3704 ;
  assign n5343 = n5342 ^ n5341 ^ 1'b0 ;
  assign n5344 = n5340 & ~n5343 ;
  assign n5345 = n330 | n1870 ;
  assign n5346 = n4416 ^ n991 ^ 1'b0 ;
  assign n5347 = ~n2064 & n5346 ;
  assign n5348 = n2610 & ~n4114 ;
  assign n5349 = n811 ^ n83 ^ 1'b0 ;
  assign n5350 = ( n532 & n4194 ) | ( n532 & ~n5349 ) | ( n4194 & ~n5349 ) ;
  assign n5353 = n928 ^ n281 ^ 1'b0 ;
  assign n5354 = ~n748 & n5353 ;
  assign n5352 = n169 | n3507 ;
  assign n5355 = n5354 ^ n5352 ^ 1'b0 ;
  assign n5356 = n1960 & ~n5355 ;
  assign n5351 = x11 & ~n3454 ;
  assign n5357 = n5356 ^ n5351 ^ 1'b0 ;
  assign n5358 = n751 | n1452 ;
  assign n5359 = ~n2023 & n3315 ;
  assign n5360 = n348 & n5359 ;
  assign n5361 = n724 & n3413 ;
  assign n5362 = n598 ^ n229 ^ 1'b0 ;
  assign n5363 = n2582 | n5362 ;
  assign n5364 = n318 & n1234 ;
  assign n5365 = n5363 | n5364 ;
  assign n5366 = n1255 | n5365 ;
  assign n5367 = n4349 ^ n111 ^ 1'b0 ;
  assign n5368 = n4048 ^ n3395 ^ 1'b0 ;
  assign n5369 = n3807 | n4607 ;
  assign n5370 = n963 & n5369 ;
  assign n5371 = n764 | n3051 ;
  assign n5372 = n5371 ^ n2318 ^ 1'b0 ;
  assign n5373 = ~n1893 & n3177 ;
  assign n5374 = n2645 & n4499 ;
  assign n5375 = ~n2049 & n5374 ;
  assign n5376 = n2210 | n4025 ;
  assign n5377 = n5375 & ~n5376 ;
  assign n5378 = n3290 ^ n1572 ^ 1'b0 ;
  assign n5379 = n763 & n1304 ;
  assign n5380 = n5379 ^ n2983 ^ 1'b0 ;
  assign n5381 = ~n2512 & n5380 ;
  assign n5382 = ~n5378 & n5381 ;
  assign n5383 = n1932 | n5382 ;
  assign n5384 = n1756 & n5050 ;
  assign n5385 = ~n97 & n5384 ;
  assign n5386 = n1428 | n2880 ;
  assign n5387 = n5192 ^ n2835 ^ 1'b0 ;
  assign n5388 = n1318 ^ n318 ^ 1'b0 ;
  assign n5389 = n1444 & ~n5388 ;
  assign n5390 = n5389 ^ n97 ^ 1'b0 ;
  assign n5391 = n4485 & n5390 ;
  assign n5392 = n769 | n1499 ;
  assign n5393 = n5392 ^ n1874 ^ 1'b0 ;
  assign n5394 = n2104 ^ n823 ^ 1'b0 ;
  assign n5395 = n5393 & ~n5394 ;
  assign n5396 = n5395 ^ n619 ^ 1'b0 ;
  assign n5397 = n965 & ~n5396 ;
  assign n5398 = n148 & ~n859 ;
  assign n5399 = n5398 ^ n1069 ^ 1'b0 ;
  assign n5400 = n833 ^ n257 ^ 1'b0 ;
  assign n5401 = n5400 ^ n2542 ^ 1'b0 ;
  assign n5402 = n4254 ^ n996 ^ 1'b0 ;
  assign n5403 = n3706 ^ n2910 ^ 1'b0 ;
  assign n5404 = ~n3771 & n5403 ;
  assign n5405 = n2160 & n4180 ;
  assign n5406 = ~n1704 & n5405 ;
  assign n5407 = n4529 & ~n5406 ;
  assign n5408 = n4165 & n5407 ;
  assign n5409 = n573 & n4745 ;
  assign n5410 = ~n4191 & n5409 ;
  assign n5411 = n5410 ^ n1632 ^ 1'b0 ;
  assign n5412 = ~n1056 & n5411 ;
  assign n5413 = n81 & ~n5412 ;
  assign n5414 = n23 | n79 ;
  assign n5415 = n745 & ~n5414 ;
  assign n5416 = n5415 ^ n55 ^ 1'b0 ;
  assign n5417 = n330 & ~n4670 ;
  assign n5418 = ~n928 & n5417 ;
  assign n5419 = n311 | n2020 ;
  assign n5420 = n3928 ^ n1463 ^ 1'b0 ;
  assign n5421 = n2880 ^ n2569 ^ n2028 ;
  assign n5422 = n1719 & n3816 ;
  assign n5423 = n3080 & n3279 ;
  assign n5424 = n5422 & ~n5423 ;
  assign n5425 = ~n252 & n1243 ;
  assign n5426 = ~n561 & n955 ;
  assign n5427 = ~n5425 & n5426 ;
  assign n5428 = n848 ^ n518 ^ 1'b0 ;
  assign n5429 = n5428 ^ n758 ^ 1'b0 ;
  assign n5430 = n1795 | n5429 ;
  assign n5431 = n794 & ~n5430 ;
  assign n5432 = n2589 ^ n518 ^ 1'b0 ;
  assign n5433 = n5431 | n5432 ;
  assign n5434 = n4058 ^ n446 ^ n223 ;
  assign n5435 = n1555 | n3974 ;
  assign n5436 = n5434 & ~n5435 ;
  assign n5437 = n2055 & ~n5436 ;
  assign n5438 = n108 & n1658 ;
  assign n5439 = n5438 ^ n3882 ^ 1'b0 ;
  assign n5440 = n743 & ~n1034 ;
  assign n5441 = ~n3247 & n5440 ;
  assign n5442 = ~n388 & n5441 ;
  assign n5443 = n857 ^ n472 ^ 1'b0 ;
  assign n5444 = n58 | n616 ;
  assign n5445 = n688 & n1810 ;
  assign n5446 = ~n3088 & n4271 ;
  assign n5447 = n5446 ^ n2420 ^ 1'b0 ;
  assign n5448 = n5445 & n5447 ;
  assign n5449 = n5448 ^ n1863 ^ 1'b0 ;
  assign n5450 = n5449 ^ n1081 ^ 1'b0 ;
  assign n5451 = ~n5444 & n5450 ;
  assign n5452 = n549 & n1201 ;
  assign n5453 = n5452 ^ n269 ^ 1'b0 ;
  assign n5454 = n5453 ^ n216 ^ 1'b0 ;
  assign n5455 = n5454 ^ n4572 ^ n2364 ;
  assign n5456 = n2689 & n3627 ;
  assign n5457 = ~n2201 & n5456 ;
  assign n5458 = n1584 | n5457 ;
  assign n5459 = n754 | n4572 ;
  assign n5460 = ~n758 & n3457 ;
  assign n5461 = n5460 ^ n888 ^ 1'b0 ;
  assign n5462 = ( n1866 & n4507 ) | ( n1866 & n5461 ) | ( n4507 & n5461 ) ;
  assign n5463 = n5459 & n5462 ;
  assign n5464 = n5221 & ~n5326 ;
  assign n5465 = ~n715 & n5464 ;
  assign n5466 = ~n833 & n3099 ;
  assign n5467 = n1999 ^ n387 ^ 1'b0 ;
  assign n5468 = ~n1492 & n5467 ;
  assign n5469 = n5468 ^ n2751 ^ 1'b0 ;
  assign n5470 = ~n1170 & n1525 ;
  assign n5471 = n764 ^ n83 ^ 1'b0 ;
  assign n5472 = n3212 & n5440 ;
  assign n5473 = n5472 ^ n2196 ^ 1'b0 ;
  assign n5474 = n339 & n3297 ;
  assign n5475 = ~n339 & n5474 ;
  assign n5476 = n575 | n5475 ;
  assign n5477 = n5475 & ~n5476 ;
  assign n5478 = ~n17 & n5477 ;
  assign n5479 = n393 | n1025 ;
  assign n5480 = n1025 & ~n5479 ;
  assign n5481 = n4311 ^ n479 ^ 1'b0 ;
  assign n5482 = n5480 | n5481 ;
  assign n5483 = n5478 & ~n5482 ;
  assign n5484 = n2941 & ~n3005 ;
  assign n5485 = n2047 & n5484 ;
  assign n5486 = ~n2047 & n5485 ;
  assign n5487 = n2642 | n3271 ;
  assign n5488 = n3271 & ~n5487 ;
  assign n5489 = n5486 | n5488 ;
  assign n5490 = n5486 & ~n5489 ;
  assign n5491 = n5490 ^ n371 ^ 1'b0 ;
  assign n5492 = n5483 | n5491 ;
  assign n5493 = n1961 ^ n46 ^ 1'b0 ;
  assign n5494 = n549 & n1979 ;
  assign n5495 = ~n818 & n5494 ;
  assign n5496 = n1979 & n3173 ;
  assign n5497 = ~n1820 & n5496 ;
  assign n5498 = n3282 ^ n2975 ^ 1'b0 ;
  assign n5499 = n2984 | n5498 ;
  assign n5500 = n5497 | n5499 ;
  assign n5501 = n5495 | n5500 ;
  assign n5502 = n2980 ^ n1608 ^ 1'b0 ;
  assign n5503 = n1950 & ~n2420 ;
  assign n5504 = n330 & n5503 ;
  assign n5505 = n5502 & n5504 ;
  assign n5506 = ~n308 & n3046 ;
  assign n5508 = n37 | n1245 ;
  assign n5507 = n1130 | n2667 ;
  assign n5509 = n5508 ^ n5507 ^ 1'b0 ;
  assign n5510 = n5506 & ~n5509 ;
  assign n5511 = n5510 ^ n342 ^ 1'b0 ;
  assign n5512 = n15 & n5511 ;
  assign n5513 = ~n1768 & n5512 ;
  assign n5514 = n2577 & n3477 ;
  assign n5515 = n4964 ^ n1523 ^ 1'b0 ;
  assign n5516 = n86 & n5515 ;
  assign n5517 = ~n1428 & n5516 ;
  assign n5518 = n4448 ^ n3277 ^ 1'b0 ;
  assign n5519 = n4246 | n4812 ;
  assign n5520 = n5518 | n5519 ;
  assign n5521 = ~n604 & n3924 ;
  assign n5522 = n2156 & n5521 ;
  assign n5523 = n564 & n5522 ;
  assign n5524 = n641 & ~n5523 ;
  assign n5525 = n2249 ^ n1219 ^ 1'b0 ;
  assign n5526 = n5525 ^ n478 ^ 1'b0 ;
  assign n5527 = n3452 & ~n5526 ;
  assign n5528 = n327 & ~n1640 ;
  assign n5529 = n1437 & ~n5528 ;
  assign n5530 = n286 | n512 ;
  assign n5531 = n3169 & n5530 ;
  assign n5532 = n5531 ^ n1344 ^ 1'b0 ;
  assign n5533 = n2151 ^ n1961 ^ 1'b0 ;
  assign n5534 = n5533 ^ n319 ^ 1'b0 ;
  assign n5535 = ~n2301 & n5534 ;
  assign n5537 = n2586 ^ n607 ^ 1'b0 ;
  assign n5538 = n5537 ^ n3080 ^ 1'b0 ;
  assign n5536 = ~n142 & n700 ;
  assign n5539 = n5538 ^ n5536 ^ 1'b0 ;
  assign n5540 = n3853 ^ n3826 ^ 1'b0 ;
  assign n5541 = n2504 | n5540 ;
  assign n5542 = n294 | n657 ;
  assign n5543 = n94 | n5542 ;
  assign n5544 = ~n3854 & n4589 ;
  assign n5549 = ~n1090 & n3352 ;
  assign n5545 = ~n81 & n191 ;
  assign n5546 = ~n177 & n1205 ;
  assign n5547 = n5546 ^ n133 ^ 1'b0 ;
  assign n5548 = n5545 & n5547 ;
  assign n5550 = n5549 ^ n5548 ^ 1'b0 ;
  assign n5551 = n1113 | n1143 ;
  assign n5552 = ~n3629 & n5551 ;
  assign n5553 = n5552 ^ n294 ^ 1'b0 ;
  assign n5554 = ~n274 & n5553 ;
  assign n5555 = n685 | n4784 ;
  assign n5556 = n2539 ^ n328 ^ 1'b0 ;
  assign n5557 = n712 | n5556 ;
  assign n5558 = n3235 & n4799 ;
  assign n5559 = n5551 & n5558 ;
  assign n5560 = n1192 ^ n78 ^ 1'b0 ;
  assign n5561 = n172 | n1562 ;
  assign n5562 = n352 & ~n2521 ;
  assign n5563 = n5562 ^ n544 ^ 1'b0 ;
  assign n5564 = n2491 & n5563 ;
  assign n5565 = n1330 & n5466 ;
  assign n5566 = ~n1453 & n5565 ;
  assign n5567 = n626 & n1873 ;
  assign n5568 = n558 & ~n1165 ;
  assign n5569 = ~n1793 & n5301 ;
  assign n5570 = ( n5567 & n5568 ) | ( n5567 & ~n5569 ) | ( n5568 & ~n5569 ) ;
  assign n5571 = n236 | n2983 ;
  assign n5572 = n5541 ^ n2124 ^ 1'b0 ;
  assign n5573 = n4453 | n5572 ;
  assign n5574 = n19 | n258 ;
  assign n5575 = n187 & n5574 ;
  assign n5576 = n1075 & ~n5575 ;
  assign n5577 = ~n1075 & n5576 ;
  assign n5578 = n5577 ^ n5005 ^ 1'b0 ;
  assign n5579 = n1736 & ~n5578 ;
  assign n5580 = n3269 ^ n931 ^ 1'b0 ;
  assign n5581 = n2762 ^ n323 ^ 1'b0 ;
  assign n5582 = n4550 | n5581 ;
  assign n5583 = n5582 ^ n3529 ^ n860 ;
  assign n5584 = ( n478 & ~n958 ) | ( n478 & n3104 ) | ( ~n958 & n3104 ) ;
  assign n5585 = ~n5583 & n5584 ;
  assign n5586 = ~n5580 & n5585 ;
  assign n5587 = n1785 ^ n88 ^ 1'b0 ;
  assign n5588 = n233 & n5587 ;
  assign n5589 = n419 & n5588 ;
  assign n5590 = n5589 ^ n4586 ^ 1'b0 ;
  assign n5591 = ~n2610 & n5484 ;
  assign n5592 = n2610 & n5591 ;
  assign n5593 = n354 | n3561 ;
  assign n5594 = n3561 & ~n5593 ;
  assign n5595 = n268 & ~n3130 ;
  assign n5596 = n3130 & n5595 ;
  assign n5597 = n3424 ^ n1141 ^ 1'b0 ;
  assign n5598 = ~n5596 & n5597 ;
  assign n5599 = ~n5594 & n5598 ;
  assign n5600 = n5594 & n5599 ;
  assign n5601 = n5592 | n5600 ;
  assign n5602 = n1802 & n3093 ;
  assign n5603 = ~n815 & n5602 ;
  assign n5604 = n5603 ^ n1573 ^ 1'b0 ;
  assign n5605 = ~n5057 & n5604 ;
  assign n5606 = n4766 ^ n3324 ^ 1'b0 ;
  assign n5609 = n1379 | n3182 ;
  assign n5607 = n274 | n3346 ;
  assign n5608 = n832 & ~n5607 ;
  assign n5610 = n5609 ^ n5608 ^ 1'b0 ;
  assign n5611 = n461 | n4465 ;
  assign n5612 = n5611 ^ n567 ^ 1'b0 ;
  assign n5613 = ~n48 & n1041 ;
  assign n5614 = n5613 ^ n5099 ^ 1'b0 ;
  assign n5615 = ~n190 & n5614 ;
  assign n5616 = ~n3514 & n3866 ;
  assign n5617 = ~n4820 & n5616 ;
  assign n5618 = n816 & n1849 ;
  assign n5619 = ~n1108 & n5618 ;
  assign n5620 = n3072 ^ n823 ^ 1'b0 ;
  assign n5621 = ~n5619 & n5620 ;
  assign n5622 = n3638 | n5621 ;
  assign n5623 = n602 | n4072 ;
  assign n5624 = ~n2176 & n3247 ;
  assign n5625 = n323 ^ n148 ^ 1'b0 ;
  assign n5626 = ( ~n2828 & n4635 ) | ( ~n2828 & n5625 ) | ( n4635 & n5625 ) ;
  assign n5627 = ~n1231 & n5626 ;
  assign n5628 = n5627 ^ n1979 ^ 1'b0 ;
  assign n5629 = n1316 & n3061 ;
  assign n5630 = n2202 & ~n5629 ;
  assign n5631 = n1404 ^ n328 ^ 1'b0 ;
  assign n5632 = n1761 & ~n5631 ;
  assign n5633 = n5632 ^ n300 ^ 1'b0 ;
  assign n5634 = n564 & n5633 ;
  assign n5635 = ~n294 & n2613 ;
  assign n5636 = n622 & ~n5635 ;
  assign n5637 = ~n5634 & n5636 ;
  assign n5638 = n5637 ^ n1143 ^ 1'b0 ;
  assign n5639 = ~n2122 & n4862 ;
  assign n5640 = ~n901 & n2542 ;
  assign n5641 = n5097 ^ n4037 ^ 1'b0 ;
  assign n5642 = ~n5640 & n5641 ;
  assign n5643 = ~n5018 & n5642 ;
  assign n5644 = n2776 ^ n1848 ^ 1'b0 ;
  assign n5645 = n2842 & n5644 ;
  assign n5646 = n5645 ^ n3822 ^ 1'b0 ;
  assign n5647 = ~n827 & n5090 ;
  assign n5648 = n5647 ^ n334 ^ 1'b0 ;
  assign n5649 = n5646 & ~n5648 ;
  assign n5650 = n1840 | n4939 ;
  assign n5651 = n376 | n5650 ;
  assign n5652 = n5651 ^ n1464 ^ 1'b0 ;
  assign n5653 = n2932 & n4697 ;
  assign n5655 = n36 & ~n60 ;
  assign n5654 = n532 & n3457 ;
  assign n5656 = n5655 ^ n5654 ^ 1'b0 ;
  assign n5657 = n5653 & n5656 ;
  assign n5658 = n470 & ~n2742 ;
  assign n5659 = n986 & n5658 ;
  assign n5660 = n5580 ^ n549 ^ 1'b0 ;
  assign n5661 = n656 ^ n14 ^ 1'b0 ;
  assign n5662 = n2136 & ~n5661 ;
  assign n5663 = n1673 & n5662 ;
  assign n5664 = n820 | n1407 ;
  assign n5665 = n5664 ^ n4241 ^ 1'b0 ;
  assign n5666 = n332 & n605 ;
  assign n5667 = n5666 ^ n489 ^ 1'b0 ;
  assign n5668 = n5071 & n5667 ;
  assign n5670 = n2624 & n3160 ;
  assign n5671 = ~n135 & n5670 ;
  assign n5672 = ~n2749 & n5671 ;
  assign n5669 = n1043 | n3118 ;
  assign n5673 = n5672 ^ n5669 ^ 1'b0 ;
  assign n5674 = n178 & n756 ;
  assign n5675 = n5673 & n5674 ;
  assign n5676 = n3620 & ~n5675 ;
  assign n5677 = ~n144 & n5676 ;
  assign n5678 = n2146 & ~n4508 ;
  assign n5679 = n5678 ^ n3305 ^ 1'b0 ;
  assign n5680 = ~n86 & n973 ;
  assign n5681 = ~n5679 & n5680 ;
  assign n5682 = n827 ^ n353 ^ 1'b0 ;
  assign n5683 = n5682 ^ n2090 ^ 1'b0 ;
  assign n5684 = ~n2751 & n5683 ;
  assign n5687 = n322 | n743 ;
  assign n5688 = n5687 ^ n894 ^ 1'b0 ;
  assign n5685 = ~n19 & n995 ;
  assign n5686 = n1113 & ~n5685 ;
  assign n5689 = n5688 ^ n5686 ^ 1'b0 ;
  assign n5690 = n949 & ~n5689 ;
  assign n5691 = n621 | n939 ;
  assign n5692 = n1939 | n3645 ;
  assign n5693 = ~n5691 & n5692 ;
  assign n5694 = ~n183 & n5693 ;
  assign n5695 = n1878 | n4528 ;
  assign n5696 = n4022 | n5695 ;
  assign n5697 = n2142 ^ n185 ^ 1'b0 ;
  assign n5698 = n4211 & ~n5697 ;
  assign n5699 = n551 | n1440 ;
  assign n5700 = n1530 | n5699 ;
  assign n5701 = n1191 & n4003 ;
  assign n5702 = n5122 ^ n1363 ^ 1'b0 ;
  assign n5703 = n5702 ^ n5205 ^ 1'b0 ;
  assign n5704 = ~n5701 & n5703 ;
  assign n5705 = n1418 ^ n198 ^ 1'b0 ;
  assign n5706 = ~n2572 & n5705 ;
  assign n5707 = n2647 & n5706 ;
  assign n5708 = ~n412 & n616 ;
  assign n5710 = ~n284 & n342 ;
  assign n5709 = ~n19 & n5031 ;
  assign n5711 = n5710 ^ n5709 ^ 1'b0 ;
  assign n5712 = n1653 & n1944 ;
  assign n5713 = n5712 ^ n55 ^ 1'b0 ;
  assign n5714 = n3907 ^ n423 ^ 1'b0 ;
  assign n5715 = n40 & n2295 ;
  assign n5716 = n484 & n5715 ;
  assign n5717 = n5186 ^ n2298 ^ 1'b0 ;
  assign n5718 = n3880 & n5717 ;
  assign n5719 = ( n3560 & ~n4243 ) | ( n3560 & n5718 ) | ( ~n4243 & n5718 ) ;
  assign n5720 = n941 | n1341 ;
  assign n5721 = n1050 & ~n2904 ;
  assign n5722 = ~n4952 & n5508 ;
  assign n5723 = n3270 ^ n1768 ^ 1'b0 ;
  assign n5724 = ~n2321 & n3211 ;
  assign n5725 = n5723 & n5724 ;
  assign n5726 = n5429 ^ n104 ^ 1'b0 ;
  assign n5727 = n3887 ^ n567 ^ 1'b0 ;
  assign n5728 = n1173 & n5727 ;
  assign n5729 = n5728 ^ n66 ^ 1'b0 ;
  assign n5730 = n2210 ^ n2204 ^ n257 ;
  assign n5731 = n748 ^ n139 ^ 1'b0 ;
  assign n5732 = n743 & ~n5731 ;
  assign n5733 = n5534 ^ n532 ^ 1'b0 ;
  assign n5734 = ~n5732 & n5733 ;
  assign n5735 = n5734 ^ n4646 ^ 1'b0 ;
  assign n5736 = n77 & n5735 ;
  assign n5738 = n553 | n1066 ;
  assign n5739 = n294 & ~n5738 ;
  assign n5737 = n454 | n624 ;
  assign n5740 = n5739 ^ n5737 ^ 1'b0 ;
  assign n5741 = n1260 ^ n949 ^ 1'b0 ;
  assign n5742 = n1307 | n2593 ;
  assign n5743 = n5742 ^ n1082 ^ 1'b0 ;
  assign n5744 = ~n3021 & n5743 ;
  assign n5745 = ~n5741 & n5744 ;
  assign n5746 = n624 & n5745 ;
  assign n5747 = n52 | n2800 ;
  assign n5748 = n955 & n976 ;
  assign n5749 = n5748 ^ n1178 ^ 1'b0 ;
  assign n5750 = n1458 & ~n5749 ;
  assign n5751 = ~n2144 & n5750 ;
  assign n5752 = n1704 | n5751 ;
  assign n5753 = n2187 ^ x1 ^ 1'b0 ;
  assign n5754 = n2549 ^ n194 ^ 1'b0 ;
  assign n5755 = n997 | n4504 ;
  assign n5756 = n699 & n2040 ;
  assign n5757 = n5756 ^ n1588 ^ 1'b0 ;
  assign n5758 = n4178 & n5757 ;
  assign n5759 = n460 & n2298 ;
  assign n5760 = n5759 ^ n1432 ^ 1'b0 ;
  assign n5761 = n5760 ^ n4281 ^ 1'b0 ;
  assign n5762 = n4511 ^ n384 ^ 1'b0 ;
  assign n5763 = ~n470 & n1234 ;
  assign n5764 = ~n637 & n1437 ;
  assign n5765 = n5763 & n5764 ;
  assign n5766 = ~n5763 & n5765 ;
  assign n5767 = n5762 & ~n5766 ;
  assign n5768 = n5767 ^ n4278 ^ 1'b0 ;
  assign n5769 = n1202 | n2242 ;
  assign n5770 = n5769 ^ n1060 ^ 1'b0 ;
  assign n5771 = n1982 & ~n5770 ;
  assign n5772 = ~n4830 & n5677 ;
  assign n5773 = n582 & n5261 ;
  assign n5774 = n489 & n5773 ;
  assign n5775 = n1231 & n1795 ;
  assign n5776 = n1260 & ~n2254 ;
  assign n5777 = n5776 ^ n5155 ^ 1'b0 ;
  assign n5778 = n5775 | n5777 ;
  assign n5779 = n382 & ~n1233 ;
  assign n5780 = n5779 ^ n78 ^ 1'b0 ;
  assign n5781 = n5780 ^ n2107 ^ 1'b0 ;
  assign n5782 = n4358 & ~n5781 ;
  assign n5783 = n5616 ^ n1186 ^ 1'b0 ;
  assign n5784 = n4469 ^ n122 ^ 1'b0 ;
  assign n5785 = n1316 ^ n175 ^ 1'b0 ;
  assign n5786 = n471 | n741 ;
  assign n5787 = n1538 & ~n5786 ;
  assign n5788 = n3741 | n5787 ;
  assign n5789 = n5702 ^ n2577 ^ 1'b0 ;
  assign n5790 = n53 | n1800 ;
  assign n5791 = n3295 & n5790 ;
  assign n5792 = ~n5789 & n5791 ;
  assign n5793 = n2337 & n2695 ;
  assign n5794 = n1545 & n2615 ;
  assign n5795 = n5794 ^ n5412 ^ 1'b0 ;
  assign n5796 = n789 ^ n43 ^ 1'b0 ;
  assign n5797 = n159 | n5796 ;
  assign n5798 = n1065 & n2155 ;
  assign n5799 = n931 | n2762 ;
  assign n5800 = n2297 | n5799 ;
  assign n5801 = n1737 ^ n457 ^ 1'b0 ;
  assign n5806 = ( ~n192 & n246 ) | ( ~n192 & n524 ) | ( n246 & n524 ) ;
  assign n5802 = n3682 ^ n638 ^ n381 ;
  assign n5803 = ~n1528 & n5802 ;
  assign n5804 = ~n2701 & n5803 ;
  assign n5805 = ~n1471 & n5804 ;
  assign n5807 = n5806 ^ n5805 ^ 1'b0 ;
  assign n5808 = n5801 | n5807 ;
  assign n5809 = n1606 ^ n679 ^ 1'b0 ;
  assign n5810 = n3415 ^ n3033 ^ 1'b0 ;
  assign n5811 = n3449 & ~n5810 ;
  assign n5812 = n5811 ^ n1566 ^ 1'b0 ;
  assign n5813 = n5172 ^ n1263 ^ 1'b0 ;
  assign n5814 = n4361 ^ n3223 ^ 1'b0 ;
  assign n5815 = n1606 & ~n1664 ;
  assign n5816 = n5815 ^ n4580 ^ 1'b0 ;
  assign n5817 = n5814 | n5816 ;
  assign n5818 = n4330 & ~n4859 ;
  assign n5819 = n3283 ^ n3125 ^ 1'b0 ;
  assign n5820 = n2799 ^ n1691 ^ 1'b0 ;
  assign n5821 = n2701 | n4680 ;
  assign n5822 = n775 & ~n2209 ;
  assign n5823 = n5822 ^ n1464 ^ 1'b0 ;
  assign n5824 = ~n405 & n5823 ;
  assign n5825 = ~n37 & n5824 ;
  assign n5826 = n1235 & n3134 ;
  assign n5827 = n915 | n2687 ;
  assign n5828 = ( n1774 & ~n2170 ) | ( n1774 & n5827 ) | ( ~n2170 & n5827 ) ;
  assign n5829 = ~n3406 & n3420 ;
  assign n5830 = n5829 ^ n630 ^ 1'b0 ;
  assign n5831 = n5830 ^ n852 ^ 1'b0 ;
  assign n5832 = ( n564 & n963 ) | ( n564 & ~n5054 ) | ( n963 & ~n5054 ) ;
  assign n5833 = n2011 ^ n278 ^ 1'b0 ;
  assign n5834 = n5453 & ~n5833 ;
  assign n5835 = ~n1957 & n5834 ;
  assign n5836 = ~n603 & n1491 ;
  assign n5837 = n1041 & n5749 ;
  assign n5838 = n2020 | n5837 ;
  assign n5839 = n5838 ^ n3255 ^ 1'b0 ;
  assign n5840 = n3443 & n5839 ;
  assign n5841 = n3776 & n5840 ;
  assign n5842 = n5324 & n5625 ;
  assign n5843 = n1511 ^ n23 ^ 1'b0 ;
  assign n5844 = n1924 & n5843 ;
  assign n5845 = x11 & ~n5844 ;
  assign n5846 = n2796 ^ n2275 ^ 1'b0 ;
  assign n5847 = n4303 & n5846 ;
  assign n5848 = ~n5845 & n5847 ;
  assign n5849 = n5848 ^ n3546 ^ 1'b0 ;
  assign n5850 = n47 & ~n191 ;
  assign n5851 = n3005 | n4220 ;
  assign n5852 = n364 ^ n239 ^ 1'b0 ;
  assign n5853 = n939 | n5852 ;
  assign n5854 = n5853 ^ n5024 ^ n205 ;
  assign n5859 = n28 | n322 ;
  assign n5855 = n1300 & n1914 ;
  assign n5856 = n5855 ^ n1169 ^ 1'b0 ;
  assign n5857 = n615 ^ n184 ^ 1'b0 ;
  assign n5858 = ~n5856 & n5857 ;
  assign n5860 = n5859 ^ n5858 ^ 1'b0 ;
  assign n5861 = ~n757 & n1227 ;
  assign n5862 = ~n1089 & n5861 ;
  assign n5863 = n3181 ^ n2851 ^ 1'b0 ;
  assign n5864 = n1525 ^ n279 ^ 1'b0 ;
  assign n5866 = n3748 ^ n3466 ^ 1'b0 ;
  assign n5865 = n639 & ~n1008 ;
  assign n5867 = n5866 ^ n5865 ^ 1'b0 ;
  assign n5868 = n4778 | n5867 ;
  assign n5869 = n1814 & n2011 ;
  assign n5870 = n5869 ^ n88 ^ 1'b0 ;
  assign n5871 = n5870 ^ n1856 ^ 1'b0 ;
  assign n5872 = n1325 ^ n272 ^ 1'b0 ;
  assign n5873 = n1880 | n5872 ;
  assign n5874 = n1931 & ~n3237 ;
  assign n5875 = n2275 | n2847 ;
  assign n5876 = n5874 | n5875 ;
  assign n5877 = n5876 ^ n2252 ^ n2244 ;
  assign n5878 = n4801 ^ n3970 ^ n2575 ;
  assign n5879 = n3237 ^ n697 ^ 1'b0 ;
  assign n5880 = n5878 & ~n5879 ;
  assign n5881 = n817 & ~n1115 ;
  assign n5882 = n5881 ^ n1462 ^ 1'b0 ;
  assign n5883 = n1453 & ~n2178 ;
  assign n5884 = ~n5882 & n5883 ;
  assign n5885 = n5884 ^ n2104 ^ 1'b0 ;
  assign n5886 = x3 | n471 ;
  assign n5887 = n5886 ^ n60 ^ 1'b0 ;
  assign n5888 = n5887 ^ n4747 ^ 1'b0 ;
  assign n5889 = ~n1865 & n5888 ;
  assign n5890 = ~n1003 & n5731 ;
  assign n5891 = n1005 | n2233 ;
  assign n5892 = n2835 | n5891 ;
  assign n5893 = n2281 ^ n1005 ^ 1'b0 ;
  assign n5894 = ~n5892 & n5893 ;
  assign n5895 = n5894 ^ n1348 ^ 1'b0 ;
  assign n5896 = x1 & ~n1113 ;
  assign n5897 = n5896 ^ n68 ^ 1'b0 ;
  assign n5898 = n5897 ^ n5649 ^ 1'b0 ;
  assign n5899 = n3814 & ~n5898 ;
  assign n5900 = ( n2695 & ~n2948 ) | ( n2695 & n4602 ) | ( ~n2948 & n4602 ) ;
  assign n5901 = ~n1115 & n2542 ;
  assign n5902 = ~n4353 & n5901 ;
  assign n5903 = n4008 ^ n599 ^ 1'b0 ;
  assign n5904 = ~n169 & n1266 ;
  assign n5905 = n2450 & ~n5904 ;
  assign n5906 = n5148 ^ n632 ^ 1'b0 ;
  assign n5907 = n1883 & ~n5906 ;
  assign n5908 = n1097 | n4906 ;
  assign n5909 = n5908 ^ n1165 ^ 1'b0 ;
  assign n5910 = n1976 & ~n5238 ;
  assign n5911 = n142 & ~n2243 ;
  assign n5912 = n4913 & n5911 ;
  assign n5913 = n241 & ~n351 ;
  assign n5914 = n970 & ~n5913 ;
  assign n5915 = n246 & ~n1315 ;
  assign n5916 = n3859 & n4418 ;
  assign n5917 = ~n2209 & n5916 ;
  assign n5918 = n1856 & n2771 ;
  assign n5919 = n5918 ^ n4722 ^ 1'b0 ;
  assign n5920 = n4291 & n5919 ;
  assign n5921 = n758 | n4977 ;
  assign n5922 = n5921 ^ n1860 ^ 1'b0 ;
  assign n5923 = n1744 & ~n3329 ;
  assign n5924 = n5204 & n5808 ;
  assign n5926 = n503 & n1373 ;
  assign n5925 = n58 | n1117 ;
  assign n5927 = n5926 ^ n5925 ^ 1'b0 ;
  assign n5928 = n1855 & n5927 ;
  assign n5929 = n1110 & n5928 ;
  assign n5930 = n1546 ^ n319 ^ 1'b0 ;
  assign n5931 = n853 | n5930 ;
  assign n5932 = n5931 ^ n4052 ^ 1'b0 ;
  assign n5933 = n1829 | n5932 ;
  assign n5934 = ~n304 & n5933 ;
  assign n5935 = n804 & ~n880 ;
  assign n5936 = n5934 & n5935 ;
  assign n5937 = n2861 & ~n3711 ;
  assign n5938 = ~n1048 & n5937 ;
  assign n5939 = n5938 ^ n4176 ^ n1914 ;
  assign n5941 = n200 | n758 ;
  assign n5940 = n809 & n1685 ;
  assign n5942 = n5941 ^ n5940 ^ 1'b0 ;
  assign n5943 = ~n2849 & n3184 ;
  assign n5944 = n1412 & ~n5943 ;
  assign n5945 = n5944 ^ n5227 ^ 1'b0 ;
  assign n5946 = ~n310 & n3204 ;
  assign n5947 = ( n1112 & ~n3924 ) | ( n1112 & n5946 ) | ( ~n3924 & n5946 ) ;
  assign n5948 = n5947 ^ n4373 ^ 1'b0 ;
  assign n5949 = ~n180 & n4548 ;
  assign n5950 = n5632 ^ n484 ^ 1'b0 ;
  assign n5951 = n949 & n5950 ;
  assign n5952 = n3347 & n5951 ;
  assign n5953 = n820 & n1431 ;
  assign n5954 = n2934 & n3376 ;
  assign n5955 = ~n1075 & n5954 ;
  assign n5956 = n2257 ^ n241 ^ 1'b0 ;
  assign n5957 = n3188 | n4976 ;
  assign n5958 = n929 | n1662 ;
  assign n5959 = n813 ^ n340 ^ 1'b0 ;
  assign n5960 = n5959 ^ n302 ^ 1'b0 ;
  assign n5961 = n1547 & ~n5960 ;
  assign n5962 = n3311 ^ n1453 ^ n1007 ;
  assign n5963 = n878 & n5962 ;
  assign n5964 = n3139 ^ n669 ^ n278 ;
  assign n5965 = n3263 & n5964 ;
  assign n5966 = n5963 & ~n5965 ;
  assign n5967 = n5966 ^ n357 ^ 1'b0 ;
  assign n5968 = n603 & ~n4535 ;
  assign n5969 = n848 & n5968 ;
  assign n5970 = n5969 ^ n2292 ^ 1'b0 ;
  assign n5971 = ( n1874 & n4350 ) | ( n1874 & n4734 ) | ( n4350 & n4734 ) ;
  assign n5972 = n3182 ^ n3149 ^ 1'b0 ;
  assign n5973 = n228 & ~n4869 ;
  assign n5974 = n268 & n5973 ;
  assign n5975 = n5424 ^ n3221 ^ 1'b0 ;
  assign n5976 = n1744 & n3404 ;
  assign n5977 = n5976 ^ n1450 ^ 1'b0 ;
  assign n5978 = n1956 ^ n1742 ^ 1'b0 ;
  assign n5979 = ( n4575 & n5977 ) | ( n4575 & n5978 ) | ( n5977 & n5978 ) ;
  assign n5980 = n2964 ^ n1893 ^ 1'b0 ;
  assign n5981 = ~n3593 & n5980 ;
  assign n5982 = n28 & n584 ;
  assign n5983 = ( n1044 & n3446 ) | ( n1044 & ~n4241 ) | ( n3446 & ~n4241 ) ;
  assign n5984 = n5983 ^ n4677 ^ 1'b0 ;
  assign n5985 = n5984 ^ n5094 ^ n168 ;
  assign n5986 = ~n4787 & n5985 ;
  assign n5987 = n1170 ^ n193 ^ 1'b0 ;
  assign n5988 = n1488 | n5987 ;
  assign n5989 = ( n1255 & ~n3307 ) | ( n1255 & n5988 ) | ( ~n3307 & n5988 ) ;
  assign n5990 = n169 | n1232 ;
  assign n5991 = ~n694 & n5099 ;
  assign n5992 = n177 & n5991 ;
  assign n5993 = n5992 ^ n3466 ^ 1'b0 ;
  assign n5994 = n1416 | n5993 ;
  assign n5995 = ~n208 & n980 ;
  assign n5996 = n2754 ^ n1483 ^ 1'b0 ;
  assign n5997 = ~n591 & n2818 ;
  assign n5998 = ~n5440 & n5997 ;
  assign n5999 = n3789 & n5053 ;
  assign n6000 = n3036 ^ n900 ^ 1'b0 ;
  assign n6001 = n3498 & ~n6000 ;
  assign n6002 = n6001 ^ n3121 ^ 1'b0 ;
  assign n6003 = n3575 & ~n6002 ;
  assign n6004 = n4798 & n5932 ;
  assign n6005 = n6004 ^ x0 ^ 1'b0 ;
  assign n6006 = ~n5013 & n5147 ;
  assign n6007 = n842 & ~n2302 ;
  assign n6008 = n6007 ^ n1388 ^ 1'b0 ;
  assign n6009 = n443 & n6008 ;
  assign n6010 = n87 & n5634 ;
  assign n6011 = n2927 ^ n2861 ^ 1'b0 ;
  assign n6012 = n3278 & n6011 ;
  assign n6013 = n3002 & n6012 ;
  assign n6014 = n5609 & n6013 ;
  assign n6015 = n6014 ^ n5971 ^ 1'b0 ;
  assign n6016 = n506 & ~n2963 ;
  assign n6017 = n1143 ^ n37 ^ 1'b0 ;
  assign n6018 = n6017 ^ n1900 ^ 1'b0 ;
  assign n6019 = n250 & n6018 ;
  assign n6020 = n4508 & ~n5863 ;
  assign n6021 = n1986 & n6020 ;
  assign n6022 = n898 ^ n815 ^ 1'b0 ;
  assign n6023 = n2553 ^ n984 ^ n628 ;
  assign n6024 = n1419 | n6023 ;
  assign n6025 = n6024 ^ n963 ^ 1'b0 ;
  assign n6026 = n2073 ^ n158 ^ 1'b0 ;
  assign n6027 = ~n734 & n1912 ;
  assign n6028 = n5796 ^ n1822 ^ n184 ;
  assign n6029 = n4327 ^ n2524 ^ 1'b0 ;
  assign n6030 = n2455 & n6029 ;
  assign n6031 = n6030 ^ n4626 ^ 1'b0 ;
  assign n6032 = ~n532 & n4440 ;
  assign n6033 = n6032 ^ n954 ^ 1'b0 ;
  assign n6034 = n2882 ^ n231 ^ n227 ;
  assign n6035 = ~n4956 & n5588 ;
  assign n6036 = n6034 & n6035 ;
  assign n6037 = n475 & ~n1833 ;
  assign n6038 = n532 & ~n3931 ;
  assign n6039 = ~n6037 & n6038 ;
  assign n6040 = n2674 ^ n338 ^ 1'b0 ;
  assign n6041 = n4517 ^ n4241 ^ 1'b0 ;
  assign n6042 = n2509 & ~n5952 ;
  assign n6043 = n6042 ^ n1722 ^ 1'b0 ;
  assign n6044 = n3025 ^ n139 ^ 1'b0 ;
  assign n6045 = ~n2105 & n6044 ;
  assign n6046 = ~n1870 & n6045 ;
  assign n6047 = n168 & ~n5848 ;
  assign n6048 = n6047 ^ n1233 ^ 1'b0 ;
  assign n6049 = n627 & n4422 ;
  assign n6050 = ~n599 & n4586 ;
  assign n6051 = n323 & n2929 ;
  assign n6052 = n3594 ^ n190 ^ 1'b0 ;
  assign n6053 = ~n4197 & n6052 ;
  assign n6054 = n2395 & n6053 ;
  assign n6055 = n2124 & n3854 ;
  assign n6056 = n6054 | n6055 ;
  assign n6057 = n6056 ^ n102 ^ 1'b0 ;
  assign n6058 = n1453 | n5913 ;
  assign n6059 = n3037 & n3742 ;
  assign n6060 = n6058 & n6059 ;
  assign n6061 = ~n458 & n1546 ;
  assign n6063 = n4591 & ~n4963 ;
  assign n6064 = ~n1315 & n6063 ;
  assign n6065 = ~n2574 & n6064 ;
  assign n6066 = n3312 | n6065 ;
  assign n6067 = n6066 ^ n4603 ^ 1'b0 ;
  assign n6062 = n2931 ^ n1306 ^ 1'b0 ;
  assign n6068 = n6067 ^ n6062 ^ 1'b0 ;
  assign n6069 = n647 & n5241 ;
  assign n6070 = ~n2286 & n6069 ;
  assign n6071 = n5309 ^ n3366 ^ 1'b0 ;
  assign n6072 = ~n1185 & n4422 ;
  assign n6074 = ~n86 & n769 ;
  assign n6073 = n364 & n1841 ;
  assign n6075 = n6074 ^ n6073 ^ 1'b0 ;
  assign n6076 = n6072 | n6075 ;
  assign n6077 = n581 & ~n6076 ;
  assign n6078 = n1166 & ~n1522 ;
  assign n6079 = ~n562 & n6078 ;
  assign n6080 = n6079 ^ n602 ^ 1'b0 ;
  assign n6081 = ~n1732 & n2545 ;
  assign n6082 = n274 & ~n6081 ;
  assign n6083 = n5683 ^ n4449 ^ 1'b0 ;
  assign n6084 = n5097 & ~n6083 ;
  assign n6085 = n1656 & ~n1718 ;
  assign n6086 = n2938 & n6085 ;
  assign n6087 = ~n1350 & n6086 ;
  assign n6093 = n2021 ^ n60 ^ 1'b0 ;
  assign n6088 = n1887 ^ n47 ^ 1'b0 ;
  assign n6089 = ~n3883 & n6088 ;
  assign n6090 = n159 | n3985 ;
  assign n6091 = ~n6089 & n6090 ;
  assign n6092 = n4825 & ~n6091 ;
  assign n6094 = n6093 ^ n6092 ^ 1'b0 ;
  assign n6095 = n2426 ^ n38 ^ 1'b0 ;
  assign n6096 = n3799 ^ n1161 ^ n1080 ;
  assign n6097 = n634 | n1297 ;
  assign n6098 = n6097 ^ n385 ^ 1'b0 ;
  assign n6099 = n5484 & n6098 ;
  assign n6100 = n2020 | n2458 ;
  assign n6101 = ~n321 & n1520 ;
  assign n6102 = n6100 & n6101 ;
  assign n6103 = n2485 ^ n1245 ^ 1'b0 ;
  assign n6104 = ~n6102 & n6103 ;
  assign n6105 = n4582 ^ n1304 ^ 1'b0 ;
  assign n6106 = n2160 & ~n6105 ;
  assign n6107 = n4852 ^ n2941 ^ 1'b0 ;
  assign n6108 = n2728 | n6107 ;
  assign n6109 = n6106 | n6108 ;
  assign n6110 = n195 & ~n3633 ;
  assign n6111 = ~n2546 & n6110 ;
  assign n6112 = n1958 & ~n2454 ;
  assign n6113 = ~n1833 & n6112 ;
  assign n6114 = n6113 ^ n3341 ^ 1'b0 ;
  assign n6115 = n6114 ^ n425 ^ 1'b0 ;
  assign n6116 = n6115 ^ n392 ^ 1'b0 ;
  assign n6117 = n3947 | n6116 ;
  assign n6125 = n2924 & ~n4683 ;
  assign n6124 = ~n1015 & n4483 ;
  assign n6126 = n6125 ^ n6124 ^ 1'b0 ;
  assign n6123 = ~n1708 & n4063 ;
  assign n6127 = n6126 ^ n6123 ^ 1'b0 ;
  assign n6119 = n759 & ~n904 ;
  assign n6120 = n1608 & n6119 ;
  assign n6118 = n387 & n3793 ;
  assign n6121 = n6120 ^ n6118 ^ 1'b0 ;
  assign n6122 = ~n2943 & n6121 ;
  assign n6128 = n6127 ^ n6122 ^ 1'b0 ;
  assign n6129 = n122 ^ n79 ^ 1'b0 ;
  assign n6130 = n1987 & n3110 ;
  assign n6131 = n6129 & n6130 ;
  assign n6132 = n3071 ^ n760 ^ 1'b0 ;
  assign n6133 = n2068 & ~n6132 ;
  assign n6134 = n6133 ^ n875 ^ 1'b0 ;
  assign n6135 = n177 & n2097 ;
  assign n6136 = ~n1918 & n3679 ;
  assign n6137 = n1491 & ~n5688 ;
  assign n6138 = n1386 | n6137 ;
  assign n6139 = n6136 & ~n6138 ;
  assign n6140 = n310 | n1620 ;
  assign n6141 = n1065 & ~n6140 ;
  assign n6142 = n6141 ^ n1950 ^ n1632 ;
  assign n6143 = n784 | n6142 ;
  assign n6144 = ~n4121 & n5730 ;
  assign n6145 = n1112 ^ n333 ^ 1'b0 ;
  assign n6146 = n4903 ^ n2380 ^ 1'b0 ;
  assign n6147 = n4233 ^ n1488 ^ 1'b0 ;
  assign n6148 = n4241 & ~n6147 ;
  assign n6149 = n1227 ^ n133 ^ 1'b0 ;
  assign n6150 = n94 | n2067 ;
  assign n6151 = n6150 ^ n621 ^ 1'b0 ;
  assign n6152 = n1043 ^ n421 ^ 1'b0 ;
  assign n6155 = ~n23 & n1599 ;
  assign n6156 = n6155 ^ n2634 ^ 1'b0 ;
  assign n6153 = n4799 ^ n1008 ^ 1'b0 ;
  assign n6154 = ~n2907 & n6153 ;
  assign n6157 = n6156 ^ n6154 ^ n3512 ;
  assign n6158 = n6152 & n6157 ;
  assign n6159 = n6158 ^ n2185 ^ 1'b0 ;
  assign n6160 = n2220 ^ n1059 ^ 1'b0 ;
  assign n6161 = n1683 & ~n6160 ;
  assign n6162 = n1202 & n6161 ;
  assign n6163 = ~n3204 & n4737 ;
  assign n6164 = n1309 ^ n495 ^ 1'b0 ;
  assign n6165 = ~n6163 & n6164 ;
  assign n6166 = n4921 & ~n6165 ;
  assign n6167 = n1129 & n5928 ;
  assign n6168 = n1377 & n1410 ;
  assign n6169 = ~n5358 & n6168 ;
  assign n6170 = n2575 ^ n2463 ^ 1'b0 ;
  assign n6171 = n6170 ^ n1063 ^ 1'b0 ;
  assign n6172 = n6171 ^ n2807 ^ 1'b0 ;
  assign n6173 = n1394 & ~n3177 ;
  assign n6174 = n508 | n1958 ;
  assign n6175 = n736 | n6174 ;
  assign n6176 = n4451 | n6175 ;
  assign n6177 = n261 | n501 ;
  assign n6178 = n472 & ~n6177 ;
  assign n6179 = n190 | n6178 ;
  assign n6180 = n833 ^ n690 ^ 1'b0 ;
  assign n6181 = ~n284 & n6180 ;
  assign n6182 = n6181 ^ n4812 ^ 1'b0 ;
  assign n6183 = n3589 ^ n381 ^ 1'b0 ;
  assign n6184 = ~n5794 & n6183 ;
  assign n6185 = n2767 ^ n1142 ^ 1'b0 ;
  assign n6186 = ~n6184 & n6185 ;
  assign n6187 = n5416 ^ n4448 ^ n4381 ;
  assign n6188 = n308 | n1304 ;
  assign n6189 = ~n2913 & n6188 ;
  assign n6190 = n4011 ^ n3360 ^ 1'b0 ;
  assign n6191 = ~n359 & n4595 ;
  assign n6192 = n3516 ^ n1110 ^ 1'b0 ;
  assign n6193 = n5927 & ~n6192 ;
  assign n6194 = ~n1963 & n6193 ;
  assign n6195 = ~n772 & n6194 ;
  assign n6196 = ~n6191 & n6195 ;
  assign n6197 = n612 & ~n615 ;
  assign n6198 = n2647 ^ n183 ^ 1'b0 ;
  assign n6199 = n1142 & ~n1506 ;
  assign n6200 = n637 & n6199 ;
  assign n6201 = ~n1324 & n5946 ;
  assign n6202 = n6201 ^ n1207 ^ 1'b0 ;
  assign n6203 = n3828 | n6202 ;
  assign n6204 = n6200 & ~n6203 ;
  assign n6205 = n2567 & n6148 ;
  assign n6206 = ~n3801 & n6205 ;
  assign n6207 = n3420 & n5094 ;
  assign n6208 = n6207 ^ n2928 ^ 1'b0 ;
  assign n6209 = n1753 | n6208 ;
  assign n6210 = ~n796 & n1381 ;
  assign n6211 = ~n541 & n6210 ;
  assign n6212 = n169 & ~n3216 ;
  assign n6213 = n3459 | n6212 ;
  assign n6216 = ~n191 & n1064 ;
  assign n6217 = n6216 ^ n246 ^ 1'b0 ;
  assign n6214 = n1833 & ~n3540 ;
  assign n6215 = n6214 ^ n102 ^ 1'b0 ;
  assign n6218 = n6217 ^ n6215 ^ 1'b0 ;
  assign n6219 = ~n330 & n3311 ;
  assign n6220 = ~n1191 & n6219 ;
  assign n6221 = n6220 ^ n984 ^ 1'b0 ;
  assign n6222 = n2499 & ~n6221 ;
  assign n6223 = n549 ^ n236 ^ 1'b0 ;
  assign n6224 = n2973 | n6223 ;
  assign n6225 = ~n178 & n4653 ;
  assign n6226 = n4132 ^ n1655 ^ 1'b0 ;
  assign n6227 = n129 | n3908 ;
  assign n6228 = n6227 ^ n512 ^ 1'b0 ;
  assign n6230 = n5273 ^ n2409 ^ 1'b0 ;
  assign n6229 = n1152 & ~n1802 ;
  assign n6231 = n6230 ^ n6229 ^ 1'b0 ;
  assign n6232 = n4192 & ~n6231 ;
  assign n6233 = n6232 ^ n2322 ^ 1'b0 ;
  assign n6234 = ~n5827 & n6233 ;
  assign n6235 = n1246 ^ n528 ^ 1'b0 ;
  assign n6236 = n4577 ^ n4098 ^ 1'b0 ;
  assign n6237 = n4404 & ~n5259 ;
  assign n6238 = n6237 ^ n622 ^ 1'b0 ;
  assign n6239 = n55 | n5092 ;
  assign n6240 = n3345 | n6239 ;
  assign n6244 = n618 ^ n384 ^ 1'b0 ;
  assign n6241 = n2476 ^ n555 ^ 1'b0 ;
  assign n6242 = n1053 & n6241 ;
  assign n6243 = n3266 & n6242 ;
  assign n6245 = n6244 ^ n6243 ^ 1'b0 ;
  assign n6246 = n47 & ~n1404 ;
  assign n6247 = n6246 ^ n4838 ^ 1'b0 ;
  assign n6248 = n470 & ~n6247 ;
  assign n6249 = ~n5409 & n6248 ;
  assign n6250 = n841 ^ n75 ^ 1'b0 ;
  assign n6251 = n6250 ^ n102 ^ 1'b0 ;
  assign n6252 = n6251 ^ n938 ^ 1'b0 ;
  assign n6253 = n287 & n6252 ;
  assign n6254 = n777 | n4029 ;
  assign n6255 = ~n2762 & n6254 ;
  assign n6256 = n6255 ^ n799 ^ 1'b0 ;
  assign n6257 = n568 & ~n4195 ;
  assign n6258 = n5635 & n6257 ;
  assign n6259 = ~n1559 & n1772 ;
  assign n6260 = n1315 & n6259 ;
  assign n6261 = n6260 ^ n977 ^ 1'b0 ;
  assign n6262 = n894 & ~n6261 ;
  assign n6263 = n1487 & ~n6262 ;
  assign n6266 = n670 ^ n52 ^ 1'b0 ;
  assign n6267 = n3725 & ~n6266 ;
  assign n6268 = n1705 & n6267 ;
  assign n6264 = n1416 ^ n169 ^ 1'b0 ;
  assign n6265 = ~n1399 & n6264 ;
  assign n6269 = n6268 ^ n6265 ^ n2482 ;
  assign n6270 = n196 & ~n6269 ;
  assign n6271 = n2733 ^ n1225 ^ 1'b0 ;
  assign n6272 = n3946 | n6271 ;
  assign n6273 = n4195 | n4379 ;
  assign n6274 = n6273 ^ n1885 ^ 1'b0 ;
  assign n6277 = n1252 ^ n428 ^ 1'b0 ;
  assign n6275 = n477 & n1430 ;
  assign n6276 = n5467 & ~n6275 ;
  assign n6278 = n6277 ^ n6276 ^ 1'b0 ;
  assign n6279 = n4959 | n5074 ;
  assign n6280 = n958 | n2898 ;
  assign n6281 = ~n5774 & n6280 ;
  assign n6284 = ~n3271 & n5682 ;
  assign n6282 = ~n1310 & n1363 ;
  assign n6283 = ~n469 & n6282 ;
  assign n6285 = n6284 ^ n6283 ^ 1'b0 ;
  assign n6286 = n2349 ^ n288 ^ 1'b0 ;
  assign n6287 = n4737 ^ n1106 ^ 1'b0 ;
  assign n6288 = n520 | n5985 ;
  assign n6289 = n3317 | n6288 ;
  assign n6290 = n1946 ^ n456 ^ 1'b0 ;
  assign n6291 = ( n286 & n1960 ) | ( n286 & ~n3869 ) | ( n1960 & ~n3869 ) ;
  assign n6292 = n2681 | n4563 ;
  assign n6293 = ~n1771 & n2696 ;
  assign n6294 = n6293 ^ n2001 ^ 1'b0 ;
  assign n6295 = ~n562 & n6294 ;
  assign n6296 = n618 ^ n216 ^ n56 ;
  assign n6297 = ~n1761 & n4739 ;
  assign n6298 = ( x0 & n6296 ) | ( x0 & n6297 ) | ( n6296 & n6297 ) ;
  assign n6299 = n185 & n2705 ;
  assign n6300 = ~n52 & n6299 ;
  assign n6301 = n5013 ^ n252 ^ 1'b0 ;
  assign n6302 = n2283 ^ n294 ^ 1'b0 ;
  assign n6303 = ~n652 & n6302 ;
  assign n6304 = n1572 & n2562 ;
  assign n6305 = n310 | n592 ;
  assign n6306 = n1264 ^ n1170 ^ 1'b0 ;
  assign n6307 = n6305 | n6306 ;
  assign n6308 = n4091 | n6307 ;
  assign n6309 = n292 & ~n567 ;
  assign n6310 = ~n292 & n6309 ;
  assign n6311 = n1560 & ~n6310 ;
  assign n6312 = n5561 | n6311 ;
  assign n6313 = n6312 ^ n1256 ^ 1'b0 ;
  assign n6314 = n6204 ^ n64 ^ 1'b0 ;
  assign n6315 = ~n2303 & n6314 ;
  assign n6316 = n2933 & ~n3601 ;
  assign n6317 = n1306 | n2810 ;
  assign n6318 = n6316 | n6317 ;
  assign n6319 = n254 & n273 ;
  assign n6320 = ~n581 & n6319 ;
  assign n6321 = n6320 ^ n977 ^ 1'b0 ;
  assign n6322 = n2824 ^ n2455 ^ 1'b0 ;
  assign n6323 = n3782 ^ n114 ^ 1'b0 ;
  assign n6324 = n4223 & ~n6017 ;
  assign n6325 = n958 & n6324 ;
  assign n6326 = ~n2386 & n4193 ;
  assign n6327 = n6325 & n6326 ;
  assign n6329 = n28 & ~n252 ;
  assign n6330 = n2674 | n3660 ;
  assign n6331 = ~n6329 & n6330 ;
  assign n6328 = n1087 & n1354 ;
  assign n6332 = n6331 ^ n6328 ^ 1'b0 ;
  assign n6333 = n3373 | n4000 ;
  assign n6334 = ~n5180 & n6333 ;
  assign n6335 = n6334 ^ n5619 ^ n1920 ;
  assign n6336 = n6335 ^ n5467 ^ n665 ;
  assign n6337 = n4667 ^ n3858 ^ 1'b0 ;
  assign n6338 = n3226 ^ n1944 ^ n52 ;
  assign n6339 = ~n549 & n1075 ;
  assign n6340 = n690 | n5915 ;
  assign n6341 = n883 & n6307 ;
  assign n6342 = n3796 & ~n6341 ;
  assign n6343 = n6342 ^ n1307 ^ 1'b0 ;
  assign n6344 = ~n3999 & n6343 ;
  assign n6345 = n1754 & n6344 ;
  assign n6346 = n359 | n3722 ;
  assign n6347 = n4590 ^ n1227 ^ 1'b0 ;
  assign n6348 = ~n1025 & n6347 ;
  assign n6349 = n290 & n6348 ;
  assign n6350 = ~n822 & n6349 ;
  assign n6351 = ~n6346 & n6350 ;
  assign n6352 = n2549 & n5206 ;
  assign n6353 = n6352 ^ n4529 ^ 1'b0 ;
  assign n6354 = n621 | n1304 ;
  assign n6355 = n6353 & ~n6354 ;
  assign n6356 = n1314 & n2546 ;
  assign n6357 = ~n1044 & n6356 ;
  assign n6358 = n1366 | n5873 ;
  assign n6359 = n2117 & ~n6358 ;
  assign n6360 = n671 & ~n1761 ;
  assign n6361 = n4078 ^ n2228 ^ 1'b0 ;
  assign n6362 = n128 | n6361 ;
  assign n6363 = n6360 & ~n6362 ;
  assign n6364 = n1452 | n3254 ;
  assign n6365 = n6364 ^ n5549 ^ 1'b0 ;
  assign n6366 = n254 & ~n4269 ;
  assign n6367 = n2639 ^ n2040 ^ 1'b0 ;
  assign n6368 = n102 & n6367 ;
  assign n6369 = n323 & n1277 ;
  assign n6370 = n792 & n6369 ;
  assign n6371 = ~n1620 & n6168 ;
  assign n6372 = ~n6370 & n6371 ;
  assign n6373 = n6368 & n6372 ;
  assign n6374 = n1083 & ~n2266 ;
  assign n6375 = ~n2330 & n6374 ;
  assign n6376 = n404 | n4055 ;
  assign n6377 = n2437 ^ n1191 ^ 1'b0 ;
  assign n6378 = n4227 ^ n263 ^ 1'b0 ;
  assign n6379 = n1086 & ~n2060 ;
  assign n6380 = n872 & ~n2751 ;
  assign n6381 = ~n2414 & n6380 ;
  assign n6382 = n3480 ^ n2347 ^ 1'b0 ;
  assign n6383 = n203 & ~n6382 ;
  assign n6384 = ~n587 & n6383 ;
  assign n6385 = n4465 ^ n528 ^ 1'b0 ;
  assign n6386 = n497 & ~n4379 ;
  assign n6387 = n6385 & n6386 ;
  assign n6388 = n2995 ^ n633 ^ 1'b0 ;
  assign n6389 = n6388 ^ n1766 ^ 1'b0 ;
  assign n6390 = ~n963 & n6389 ;
  assign n6391 = n1936 ^ n1887 ^ 1'b0 ;
  assign n6392 = n83 | n6391 ;
  assign n6393 = n4220 ^ n2242 ^ 1'b0 ;
  assign n6394 = n5760 & n6393 ;
  assign n6395 = n6394 ^ n1480 ^ 1'b0 ;
  assign n6398 = n1845 ^ n741 ^ 1'b0 ;
  assign n6396 = n879 & n2509 ;
  assign n6397 = n6396 ^ n3376 ^ 1'b0 ;
  assign n6399 = n6398 ^ n6397 ^ 1'b0 ;
  assign n6400 = n3580 ^ n2433 ^ 1'b0 ;
  assign n6401 = ( n1624 & n6399 ) | ( n1624 & ~n6400 ) | ( n6399 & ~n6400 ) ;
  assign n6402 = n806 & n1423 ;
  assign n6403 = n2034 & ~n4941 ;
  assign n6404 = n1527 & ~n1979 ;
  assign n6405 = n789 & n6404 ;
  assign n6406 = n2284 | n6405 ;
  assign n6407 = n6113 ^ n1152 ^ 1'b0 ;
  assign n6408 = n2948 ^ n280 ^ 1'b0 ;
  assign n6409 = n6408 ^ n414 ^ 1'b0 ;
  assign n6410 = ~n3577 & n6409 ;
  assign n6411 = ~n161 & n6410 ;
  assign n6412 = n2438 & n3776 ;
  assign n6413 = n323 | n2834 ;
  assign n6414 = n3164 & ~n6413 ;
  assign n6416 = n683 | n1368 ;
  assign n6415 = n1103 | n2038 ;
  assign n6417 = n6416 ^ n6415 ^ 1'b0 ;
  assign n6418 = n3603 | n6417 ;
  assign n6419 = n6418 ^ n123 ^ 1'b0 ;
  assign n6420 = n1928 & ~n4024 ;
  assign n6421 = n552 & ~n3567 ;
  assign n6422 = n1469 ^ n977 ^ 1'b0 ;
  assign n6423 = n947 & ~n2676 ;
  assign n6424 = n6423 ^ n800 ^ 1'b0 ;
  assign n6425 = n880 | n6424 ;
  assign n6426 = n1112 & ~n6425 ;
  assign n6427 = n6426 ^ n3817 ^ 1'b0 ;
  assign n6428 = n3769 ^ n471 ^ 1'b0 ;
  assign n6429 = n6428 ^ n5907 ^ 1'b0 ;
  assign n6430 = n6003 ^ n573 ^ 1'b0 ;
  assign n6432 = ~n3008 & n4214 ;
  assign n6431 = n4689 ^ n175 ^ 1'b0 ;
  assign n6433 = n6432 ^ n6431 ^ n2577 ;
  assign n6435 = n2977 ^ n276 ^ 1'b0 ;
  assign n6436 = ~n1309 & n6435 ;
  assign n6437 = n6436 ^ n286 ^ 1'b0 ;
  assign n6438 = n2332 & ~n6437 ;
  assign n6434 = n5830 ^ n4879 ^ 1'b0 ;
  assign n6439 = n6438 ^ n6434 ^ 1'b0 ;
  assign n6440 = n190 & ~n596 ;
  assign n6441 = n514 & n1047 ;
  assign n6442 = n2846 ^ n544 ^ 1'b0 ;
  assign n6443 = n3514 | n6442 ;
  assign n6444 = n2027 & ~n4347 ;
  assign n6445 = ~n330 & n1073 ;
  assign n6446 = n2294 & ~n2642 ;
  assign n6447 = n6446 ^ n2059 ^ 1'b0 ;
  assign n6448 = n5314 & n6447 ;
  assign n6449 = n6445 & n6448 ;
  assign n6450 = ~n3719 & n6449 ;
  assign n6451 = n635 & ~n5012 ;
  assign n6452 = n2939 ^ n51 ^ 1'b0 ;
  assign n6453 = n4629 & n6452 ;
  assign n6454 = n6453 ^ n4531 ^ 1'b0 ;
  assign n6455 = n123 & n5749 ;
  assign n6456 = n6455 ^ n5256 ^ 1'b0 ;
  assign n6457 = n3220 ^ n2900 ^ 1'b0 ;
  assign n6458 = n142 | n6457 ;
  assign n6459 = ~n1096 & n6458 ;
  assign n6460 = ~n1473 & n4296 ;
  assign n6461 = n382 & n6460 ;
  assign n6462 = ~n1324 & n6162 ;
  assign n6463 = n5941 ^ n2735 ^ 1'b0 ;
  assign n6468 = n4136 ^ n985 ^ 1'b0 ;
  assign n6464 = n6142 ^ n5095 ^ 1'b0 ;
  assign n6465 = n1719 ^ n164 ^ 1'b0 ;
  assign n6466 = n6464 & n6465 ;
  assign n6467 = ~n4990 & n6466 ;
  assign n6469 = n6468 ^ n6467 ^ 1'b0 ;
  assign n6470 = n74 | n133 ;
  assign n6471 = n6470 ^ n2476 ^ 1'b0 ;
  assign n6472 = ( ~n98 & n1581 ) | ( ~n98 & n6471 ) | ( n1581 & n6471 ) ;
  assign n6473 = n2486 ^ n1940 ^ 1'b0 ;
  assign n6474 = n3186 & n6473 ;
  assign n6475 = ( n246 & n1220 ) | ( n246 & ~n6474 ) | ( n1220 & ~n6474 ) ;
  assign n6476 = n4589 & n6475 ;
  assign n6477 = ( ~n3158 & n5288 ) | ( ~n3158 & n5684 ) | ( n5288 & n5684 ) ;
  assign n6478 = x0 & ~n2059 ;
  assign n6479 = ~n5125 & n6478 ;
  assign n6480 = ~n1174 & n4482 ;
  assign n6481 = n6480 ^ n6444 ^ 1'b0 ;
  assign n6482 = n1867 ^ n1304 ^ 1'b0 ;
  assign n6484 = n2109 & ~n2303 ;
  assign n6483 = ~n1855 & n6127 ;
  assign n6485 = n6484 ^ n6483 ^ 1'b0 ;
  assign n6486 = n1693 & n3068 ;
  assign n6487 = n1431 ^ n226 ^ 1'b0 ;
  assign n6488 = n1884 & n6487 ;
  assign n6489 = ~n1812 & n1845 ;
  assign n6490 = n729 ^ n673 ^ n322 ;
  assign n6491 = ~n1339 & n6490 ;
  assign n6492 = n6489 & n6491 ;
  assign n6495 = n1944 & ~n6054 ;
  assign n6496 = n5135 & n6495 ;
  assign n6497 = n880 ^ n741 ^ 1'b0 ;
  assign n6498 = n276 & n6497 ;
  assign n6499 = ~n1398 & n6498 ;
  assign n6500 = n6496 & n6499 ;
  assign n6501 = n191 & ~n6500 ;
  assign n6493 = n1399 & ~n5831 ;
  assign n6494 = n5547 & n6493 ;
  assign n6502 = n6501 ^ n6494 ^ 1'b0 ;
  assign n6503 = n4166 ^ n879 ^ 1'b0 ;
  assign n6504 = n4600 & ~n6503 ;
  assign n6505 = ~n585 & n1924 ;
  assign n6506 = ~n929 & n6505 ;
  assign n6507 = n3533 | n6506 ;
  assign n6508 = n4100 | n6507 ;
  assign n6509 = n604 & ~n608 ;
  assign n6510 = n295 | n5612 ;
  assign n6511 = ~n216 & n323 ;
  assign n6512 = ~n5355 & n6511 ;
  assign n6513 = n1690 | n3929 ;
  assign n6514 = n6512 & ~n6513 ;
  assign n6515 = n4256 | n4924 ;
  assign n6516 = n2279 & ~n3602 ;
  assign n6517 = ~n2279 & n6516 ;
  assign n6518 = ~n5164 & n6517 ;
  assign n6519 = n2369 | n3462 ;
  assign n6520 = n1975 & ~n4933 ;
  assign n6521 = n6520 ^ n1474 ^ 1'b0 ;
  assign n6522 = n757 | n6521 ;
  assign n6523 = n3845 & ~n6522 ;
  assign n6524 = n985 & ~n1994 ;
  assign n6525 = ~n1970 & n6524 ;
  assign n6526 = n3284 & n4251 ;
  assign n6527 = n1415 & ~n3162 ;
  assign n6528 = n5533 & ~n6527 ;
  assign n6529 = n690 & n6528 ;
  assign n6530 = n3532 & ~n6501 ;
  assign n6531 = n539 ^ n484 ^ 1'b0 ;
  assign n6532 = ~n958 & n6079 ;
  assign n6533 = ~n544 & n6532 ;
  assign n6534 = n638 & n2436 ;
  assign n6535 = n3342 ^ n2236 ^ 1'b0 ;
  assign n6536 = n6534 & ~n6535 ;
  assign n6537 = n1271 & ~n3883 ;
  assign n6538 = ~n79 & n582 ;
  assign n6539 = n6538 ^ n3286 ^ 1'b0 ;
  assign n6540 = n6045 & n6400 ;
  assign n6541 = n1658 | n4044 ;
  assign n6542 = n816 ^ n122 ^ 1'b0 ;
  assign n6543 = n6541 | n6542 ;
  assign n6544 = n5269 ^ n2341 ^ 1'b0 ;
  assign n6545 = n6544 ^ n319 ^ 1'b0 ;
  assign n6546 = ~n1158 & n6545 ;
  assign n6547 = ~n5404 & n5733 ;
  assign n6548 = n1331 & ~n4114 ;
  assign n6549 = n6548 ^ n5096 ^ 1'b0 ;
  assign n6550 = n6549 ^ n348 ^ 1'b0 ;
  assign n6551 = n3345 & ~n6550 ;
  assign n6552 = ~n601 & n5968 ;
  assign n6562 = n1754 & ~n3549 ;
  assign n6561 = n857 | n2999 ;
  assign n6563 = n6562 ^ n6561 ^ 1'b0 ;
  assign n6553 = n1048 & ~n2700 ;
  assign n6554 = n4673 ^ n381 ^ 1'b0 ;
  assign n6555 = ~n6553 & n6554 ;
  assign n6556 = n1229 | n3570 ;
  assign n6557 = n1010 | n6556 ;
  assign n6558 = n3935 & n6557 ;
  assign n6559 = n6558 ^ n4683 ^ 1'b0 ;
  assign n6560 = n6555 & n6559 ;
  assign n6564 = n6563 ^ n6560 ^ 1'b0 ;
  assign n6565 = n6552 & ~n6564 ;
  assign n6566 = n2933 | n5760 ;
  assign n6567 = n2238 | n2294 ;
  assign n6568 = ~n200 & n501 ;
  assign n6569 = n6568 ^ n684 ^ 1'b0 ;
  assign n6570 = n1250 ^ n758 ^ 1'b0 ;
  assign n6571 = n274 | n6570 ;
  assign n6572 = n2478 | n3184 ;
  assign n6573 = n6572 ^ n1254 ^ 1'b0 ;
  assign n6574 = ~n6571 & n6573 ;
  assign n6575 = n6574 ^ n1308 ^ 1'b0 ;
  assign n6576 = n861 & ~n3449 ;
  assign n6577 = ~n6575 & n6576 ;
  assign n6578 = n6577 ^ n3318 ^ 1'b0 ;
  assign n6579 = n3264 ^ n3194 ^ 1'b0 ;
  assign n6580 = n6248 & ~n6579 ;
  assign n6581 = ~n290 & n1144 ;
  assign n6582 = n2142 & n6581 ;
  assign n6583 = ~n6580 & n6582 ;
  assign n6584 = n4126 ^ n3707 ^ 1'b0 ;
  assign n6586 = n1495 ^ n109 ^ 1'b0 ;
  assign n6585 = n3929 ^ n2188 ^ 1'b0 ;
  assign n6587 = n6586 ^ n6585 ^ 1'b0 ;
  assign n6588 = n6271 ^ n5377 ^ 1'b0 ;
  assign n6589 = n1659 | n4877 ;
  assign n6590 = n1760 | n3699 ;
  assign n6591 = ~n5023 & n6590 ;
  assign n6592 = ~n6589 & n6591 ;
  assign n6593 = n3228 ^ n1506 ^ 1'b0 ;
  assign n6594 = n2456 & n6593 ;
  assign n6595 = n6594 ^ n161 ^ 1'b0 ;
  assign n6596 = n766 ^ n536 ^ 1'b0 ;
  assign n6597 = ~n117 & n6596 ;
  assign n6598 = ~n2925 & n6597 ;
  assign n6599 = n6598 ^ n4197 ^ 1'b0 ;
  assign n6600 = n6599 ^ n2100 ^ 1'b0 ;
  assign n6601 = ~n2428 & n6600 ;
  assign n6602 = n2410 ^ n641 ^ 1'b0 ;
  assign n6603 = n6602 ^ n5180 ^ 1'b0 ;
  assign n6604 = n799 & ~n6603 ;
  assign n6605 = ~n4434 & n6604 ;
  assign n6606 = ~n3247 & n3265 ;
  assign n6607 = n6606 ^ n4606 ^ 1'b0 ;
  assign n6608 = ~n1655 & n3552 ;
  assign n6609 = n6608 ^ n1512 ^ 1'b0 ;
  assign n6610 = n2966 & n6609 ;
  assign n6611 = n2850 & ~n3877 ;
  assign n6612 = n2277 | n6611 ;
  assign n6613 = n3221 & ~n6612 ;
  assign n6614 = n6260 | n6613 ;
  assign n6615 = n6614 ^ n1732 ^ 1'b0 ;
  assign n6616 = n6615 ^ n2608 ^ 1'b0 ;
  assign n6617 = n369 & ~n1368 ;
  assign n6618 = n4449 ^ n866 ^ 1'b0 ;
  assign n6619 = n1260 & ~n6618 ;
  assign n6620 = n2700 ^ n265 ^ 1'b0 ;
  assign n6621 = n2568 ^ n164 ^ 1'b0 ;
  assign n6622 = n6620 & ~n6621 ;
  assign n6623 = ~n1227 & n6622 ;
  assign n6625 = n2436 ^ n1308 ^ 1'b0 ;
  assign n6626 = ~n1001 & n6625 ;
  assign n6624 = ~n692 & n6179 ;
  assign n6627 = n6626 ^ n6624 ^ 1'b0 ;
  assign n6628 = n5724 ^ n2243 ^ 1'b0 ;
  assign n6629 = n6628 ^ n2484 ^ 1'b0 ;
  assign n6638 = n1774 & n4487 ;
  assign n6639 = ~n4487 & n6638 ;
  assign n6630 = n37 | n2201 ;
  assign n6631 = n6630 ^ n713 ^ 1'b0 ;
  assign n6632 = n2256 | n6631 ;
  assign n6633 = n446 & ~n6632 ;
  assign n6634 = n1300 ^ n37 ^ 1'b0 ;
  assign n6635 = ~n6633 & n6634 ;
  assign n6636 = ~n155 & n6635 ;
  assign n6637 = n6300 | n6636 ;
  assign n6640 = n6639 ^ n6637 ^ 1'b0 ;
  assign n6641 = n2316 | n3141 ;
  assign n6642 = n4869 | n6641 ;
  assign n6643 = n6642 ^ n1555 ^ 1'b0 ;
  assign n6644 = n389 & n709 ;
  assign n6645 = ~n1270 & n2591 ;
  assign n6646 = ~n1039 & n6645 ;
  assign n6647 = n270 | n997 ;
  assign n6650 = n2065 | n4392 ;
  assign n6651 = n6650 ^ n290 ^ 1'b0 ;
  assign n6648 = n4088 ^ n709 ^ 1'b0 ;
  assign n6649 = n2482 & ~n6648 ;
  assign n6652 = n6651 ^ n6649 ^ 1'b0 ;
  assign n6653 = n6647 & ~n6652 ;
  assign n6654 = n1864 ^ n624 ^ 1'b0 ;
  assign n6655 = n4079 & n6654 ;
  assign n6656 = n6655 ^ n4706 ^ 1'b0 ;
  assign n6657 = n3360 & ~n4517 ;
  assign n6658 = ~n3477 & n6657 ;
  assign n6659 = n107 & ~n446 ;
  assign n6660 = n6659 ^ n3185 ^ 1'b0 ;
  assign n6661 = n963 | n2963 ;
  assign n6662 = n1492 | n6661 ;
  assign n6663 = n5532 | n6662 ;
  assign n6664 = n158 & ~n1920 ;
  assign n6665 = n1550 & n6664 ;
  assign n6666 = n231 & n6503 ;
  assign n6667 = n6666 ^ n75 ^ 1'b0 ;
  assign n6668 = n811 & ~n1691 ;
  assign n6669 = n6668 ^ n2951 ^ 1'b0 ;
  assign n6670 = n5853 & n6669 ;
  assign n6671 = ( n2431 & n4892 ) | ( n2431 & n6670 ) | ( n4892 & n6670 ) ;
  assign n6672 = n135 | n1219 ;
  assign n6673 = ( n641 & ~n5823 ) | ( n641 & n5974 ) | ( ~n5823 & n5974 ) ;
  assign n6674 = n365 & n4074 ;
  assign n6675 = n5382 ^ n4453 ^ 1'b0 ;
  assign n6676 = ~n4117 & n6675 ;
  assign n6677 = n584 & ~n3292 ;
  assign n6678 = n507 & n5512 ;
  assign n6679 = n6678 ^ n2759 ^ 1'b0 ;
  assign n6680 = n5493 | n6679 ;
  assign n6681 = n6680 ^ n5900 ^ 1'b0 ;
  assign n6682 = ( n2025 & ~n2222 ) | ( n2025 & n3830 ) | ( ~n2222 & n3830 ) ;
  assign n6683 = n2910 & ~n4349 ;
  assign n6684 = n3221 & ~n3350 ;
  assign n6685 = n3719 & n6684 ;
  assign n6686 = n4815 & ~n6685 ;
  assign n6687 = n6686 ^ n5655 ^ 1'b0 ;
  assign n6688 = n159 ^ n142 ^ 1'b0 ;
  assign n6689 = n2011 & ~n6688 ;
  assign n6690 = n6689 ^ n880 ^ 1'b0 ;
  assign n6691 = n6031 | n6690 ;
  assign n6693 = ~n1878 & n5180 ;
  assign n6694 = ~n4042 & n6693 ;
  assign n6692 = ~n4254 & n5367 ;
  assign n6695 = n6694 ^ n6692 ^ 1'b0 ;
  assign n6696 = n6695 ^ n4269 ^ 1'b0 ;
  assign n6697 = n1463 & ~n6696 ;
  assign n6698 = n5431 ^ n4195 ^ 1'b0 ;
  assign n6699 = n1961 ^ n618 ^ 1'b0 ;
  assign n6700 = ~n471 & n6699 ;
  assign n6701 = ~n454 & n6700 ;
  assign n6702 = n6701 ^ n5831 ^ 1'b0 ;
  assign n6703 = ~n1683 & n2637 ;
  assign n6704 = n2282 ^ n1450 ^ 1'b0 ;
  assign n6705 = ~n6703 & n6704 ;
  assign n6706 = n1721 ^ n159 ^ 1'b0 ;
  assign n6707 = n962 & n6706 ;
  assign n6708 = ~n79 & n1520 ;
  assign n6709 = n6708 ^ n154 ^ 1'b0 ;
  assign n6710 = ~n1015 & n6709 ;
  assign n6711 = n2695 & ~n5190 ;
  assign n6712 = n177 & n6711 ;
  assign n6713 = n378 & ~n951 ;
  assign n6714 = n6713 ^ n1093 ^ 1'b0 ;
  assign n6715 = n6712 & n6714 ;
  assign n6718 = n1674 | n3374 ;
  assign n6716 = n1693 ^ n1683 ^ 1'b0 ;
  assign n6717 = n1756 & ~n6716 ;
  assign n6719 = n6718 ^ n6717 ^ 1'b0 ;
  assign n6720 = n3398 & ~n3823 ;
  assign n6721 = n1798 & ~n3191 ;
  assign n6722 = n6721 ^ n2347 ^ 1'b0 ;
  assign n6723 = ~n2025 & n6722 ;
  assign n6724 = n1106 ^ n741 ^ 1'b0 ;
  assign n6725 = n2191 & ~n6724 ;
  assign n6726 = n6725 ^ n1693 ^ 1'b0 ;
  assign n6727 = n2906 ^ n229 ^ 1'b0 ;
  assign n6728 = n527 & n6727 ;
  assign n6729 = n4536 ^ n853 ^ 1'b0 ;
  assign n6730 = n931 | n1769 ;
  assign n6731 = n128 & ~n1039 ;
  assign n6732 = ~n6730 & n6731 ;
  assign n6733 = n5735 ^ n497 ^ 1'b0 ;
  assign n6734 = ~n5428 & n6733 ;
  assign n6735 = n6730 ^ n6392 ^ 1'b0 ;
  assign n6736 = n3251 | n3940 ;
  assign n6737 = n6736 ^ n1081 ^ 1'b0 ;
  assign n6738 = n6737 ^ n2577 ^ 1'b0 ;
  assign n6739 = n6735 & n6738 ;
  assign n6742 = n2531 ^ n1615 ^ 1'b0 ;
  assign n6740 = n1125 ^ n591 ^ 1'b0 ;
  assign n6741 = n3433 | n6740 ;
  assign n6743 = n6742 ^ n6741 ^ 1'b0 ;
  assign n6748 = n2150 ^ n1649 ^ n857 ;
  assign n6744 = n350 & ~n705 ;
  assign n6745 = n6744 ^ n608 ^ 1'b0 ;
  assign n6746 = ( ~n1224 & n3475 ) | ( ~n1224 & n4732 ) | ( n3475 & n4732 ) ;
  assign n6747 = n6745 & ~n6746 ;
  assign n6749 = n6748 ^ n6747 ^ 1'b0 ;
  assign n6750 = n928 & n5909 ;
  assign n6751 = n387 & n1188 ;
  assign n6752 = n6751 ^ n1044 ^ 1'b0 ;
  assign n6753 = n2693 ^ n1500 ^ 1'b0 ;
  assign n6754 = ~n2727 & n3475 ;
  assign n6755 = n6753 & n6754 ;
  assign n6756 = n6752 | n6755 ;
  assign n6757 = n6750 & ~n6756 ;
  assign n6760 = ~n844 & n3476 ;
  assign n6761 = ~n369 & n6760 ;
  assign n6758 = n83 | n6714 ;
  assign n6759 = n4136 | n6758 ;
  assign n6762 = n6761 ^ n6759 ^ n5431 ;
  assign n6763 = n1325 & ~n5269 ;
  assign n6764 = n6763 ^ n2973 ^ 1'b0 ;
  assign n6765 = n236 | n846 ;
  assign n6766 = n2116 & ~n6765 ;
  assign n6767 = n514 & n1235 ;
  assign n6768 = n6767 ^ n1323 ^ 1'b0 ;
  assign n6769 = ~n3599 & n6768 ;
  assign n6770 = n3756 | n6769 ;
  assign n6771 = n5574 & n6770 ;
  assign n6772 = n3181 | n4944 ;
  assign n6773 = n767 & n823 ;
  assign n6774 = ~n1268 & n5256 ;
  assign n6775 = n2807 & n6774 ;
  assign n6776 = n3694 | n6198 ;
  assign n6779 = n1205 & n3687 ;
  assign n6777 = n1552 | n5606 ;
  assign n6778 = n1082 | n6777 ;
  assign n6780 = n6779 ^ n6778 ^ 1'b0 ;
  assign n6781 = n3632 ^ n3502 ^ 1'b0 ;
  assign n6782 = n6781 ^ n6725 ^ 1'b0 ;
  assign n6783 = n226 & n6782 ;
  assign n6784 = ( n167 & n335 ) | ( n167 & ~n1591 ) | ( n335 & ~n1591 ) ;
  assign n6785 = ~n3887 & n5556 ;
  assign n6786 = n869 & n5161 ;
  assign n6787 = n1933 | n6527 ;
  assign n6788 = n2679 & ~n6787 ;
  assign n6789 = n4450 ^ n843 ^ 1'b0 ;
  assign n6790 = n299 & ~n1004 ;
  assign n6791 = ~n299 & n6790 ;
  assign n6792 = n390 | n6791 ;
  assign n6793 = n390 & ~n6792 ;
  assign n6794 = n116 | n304 ;
  assign n6795 = n116 & ~n6794 ;
  assign n6796 = n6795 ^ n4024 ^ 1'b0 ;
  assign n6797 = n6793 & n6796 ;
  assign n6802 = n97 & ~n304 ;
  assign n6803 = ~n97 & n6802 ;
  assign n6798 = x6 & ~n64 ;
  assign n6799 = ~x6 & n6798 ;
  assign n6800 = n278 & n6799 ;
  assign n6801 = n896 & n6800 ;
  assign n6804 = n6803 ^ n6801 ^ 1'b0 ;
  assign n6805 = n6797 & n6804 ;
  assign n6806 = ~n6797 & n6805 ;
  assign n6807 = n3745 ^ n1759 ^ 1'b0 ;
  assign n6808 = ~n2996 & n6807 ;
  assign n6809 = n258 | n857 ;
  assign n6810 = ~n1982 & n3579 ;
  assign n6811 = n489 & n3505 ;
  assign n6812 = ~n1388 & n6811 ;
  assign n6813 = n6810 & ~n6812 ;
  assign n6814 = n6809 & n6813 ;
  assign n6815 = n3903 ^ n1199 ^ 1'b0 ;
  assign n6816 = n458 | n6815 ;
  assign n6817 = ~n239 & n476 ;
  assign n6821 = n1552 ^ n671 ^ 1'b0 ;
  assign n6822 = n1655 & ~n6821 ;
  assign n6818 = n781 ^ n158 ^ 1'b0 ;
  assign n6819 = n5133 & ~n6818 ;
  assign n6820 = n532 & n6819 ;
  assign n6823 = n6822 ^ n6820 ^ 1'b0 ;
  assign n6824 = ~n747 & n2700 ;
  assign n6825 = n4268 & n6824 ;
  assign n6826 = n2476 & n6825 ;
  assign n6827 = n2919 ^ n114 ^ 1'b0 ;
  assign n6828 = n4025 & ~n6827 ;
  assign n6830 = n3369 & n3993 ;
  assign n6831 = n556 | n1227 ;
  assign n6832 = n3314 | n6831 ;
  assign n6833 = n6830 & ~n6832 ;
  assign n6829 = ~n52 & n3317 ;
  assign n6834 = n6833 ^ n6829 ^ 1'b0 ;
  assign n6835 = n3008 & n4756 ;
  assign n6836 = n1887 & n5025 ;
  assign n6837 = n6836 ^ n5882 ^ 1'b0 ;
  assign n6838 = n6837 ^ n3583 ^ 1'b0 ;
  assign n6839 = ~n6835 & n6838 ;
  assign n6840 = n4564 ^ n1425 ^ 1'b0 ;
  assign n6841 = ~n547 & n6840 ;
  assign n6842 = n1064 ^ n667 ^ 1'b0 ;
  assign n6843 = n6841 & ~n6842 ;
  assign n6844 = n2882 | n6071 ;
  assign n6845 = n5377 & ~n6844 ;
  assign n6846 = n3459 ^ n3290 ^ n484 ;
  assign n6847 = n1775 & ~n4679 ;
  assign n6852 = ~n986 & n6275 ;
  assign n6848 = n771 | n2896 ;
  assign n6849 = n866 & ~n6848 ;
  assign n6850 = n6849 ^ n3427 ^ 1'b0 ;
  assign n6851 = ~n4664 & n6850 ;
  assign n6853 = n6852 ^ n6851 ^ 1'b0 ;
  assign n6854 = n892 ^ n857 ^ 1'b0 ;
  assign n6855 = ~n1003 & n6854 ;
  assign n6856 = ~n4120 & n6855 ;
  assign n6857 = n6856 ^ n4812 ^ 1'b0 ;
  assign n6858 = ~n699 & n1331 ;
  assign n6859 = n1072 & n1287 ;
  assign n6860 = n6858 & n6859 ;
  assign n6862 = n4842 & n6367 ;
  assign n6861 = n1851 | n1909 ;
  assign n6863 = n6862 ^ n6861 ^ 1'b0 ;
  assign n6864 = n1007 ^ x0 ^ 1'b0 ;
  assign n6866 = n3357 ^ n3191 ^ 1'b0 ;
  assign n6865 = n2618 ^ n338 ^ 1'b0 ;
  assign n6867 = n6866 ^ n6865 ^ 1'b0 ;
  assign n6868 = ~n6174 & n6867 ;
  assign n6869 = n6864 & n6868 ;
  assign n6870 = n6869 ^ n1086 ^ 1'b0 ;
  assign n6871 = n4446 & n5582 ;
  assign n6872 = ~n2400 & n4668 ;
  assign n6873 = n6151 & n6872 ;
  assign n6874 = n3557 ^ n2060 ^ 1'b0 ;
  assign n6875 = n2205 & ~n6874 ;
  assign n6876 = ~n161 & n3348 ;
  assign n6877 = n1043 | n3305 ;
  assign n6878 = n6877 ^ n5158 ^ 1'b0 ;
  assign n6879 = ~n6876 & n6878 ;
  assign n6880 = n6879 ^ n3990 ^ 1'b0 ;
  assign n6881 = n60 | n6880 ;
  assign n6882 = n1802 & n2134 ;
  assign n6883 = n4204 ^ n3940 ^ 1'b0 ;
  assign n6884 = n6882 & n6883 ;
  assign n6885 = n6763 ^ n1659 ^ 1'b0 ;
  assign n6886 = n3220 ^ n2894 ^ 1'b0 ;
  assign n6889 = n2459 & n4866 ;
  assign n6887 = n191 & ~n460 ;
  assign n6888 = ~n5067 & n6887 ;
  assign n6890 = n6889 ^ n6888 ^ 1'b0 ;
  assign n6891 = n4653 & ~n5000 ;
  assign n6892 = n6891 ^ n4416 ^ 1'b0 ;
  assign n6893 = n2086 & n3327 ;
  assign n6894 = n3481 & n6893 ;
  assign n6895 = n5289 | n6894 ;
  assign n6896 = n4728 | n6895 ;
  assign n6897 = n899 ^ n284 ^ 1'b0 ;
  assign n6898 = n2022 | n6626 ;
  assign n6899 = n6897 | n6898 ;
  assign n6900 = n4884 ^ n4430 ^ 1'b0 ;
  assign n6901 = n246 & n445 ;
  assign n6902 = n3579 ^ n740 ^ 1'b0 ;
  assign n6903 = n268 & n1499 ;
  assign n6904 = n6903 ^ n6194 ^ 1'b0 ;
  assign n6908 = n1598 ^ n1533 ^ 1'b0 ;
  assign n6909 = n328 & ~n6908 ;
  assign n6910 = n1909 & n6909 ;
  assign n6905 = n35 | n1705 ;
  assign n6906 = n3013 & ~n6905 ;
  assign n6907 = n6906 ^ n6742 ^ 1'b0 ;
  assign n6911 = n6910 ^ n6907 ^ n5848 ;
  assign n6912 = n1979 & n5065 ;
  assign n6913 = ~x2 & n1080 ;
  assign n6914 = ~n3199 & n3329 ;
  assign n6915 = ~n6913 & n6914 ;
  assign n6916 = n354 & n1565 ;
  assign n6917 = n2707 & ~n3803 ;
  assign n6918 = n6916 & n6917 ;
  assign n6919 = n6051 | n6918 ;
  assign n6920 = ~n1608 & n1714 ;
  assign n6921 = n318 & ~n1178 ;
  assign n6922 = n2316 ^ n549 ^ 1'b0 ;
  assign n6923 = n1758 & ~n4537 ;
  assign n6924 = n4125 ^ n2825 ^ n96 ;
  assign n6928 = ~n68 & n1141 ;
  assign n6929 = n2243 & n6928 ;
  assign n6930 = n6929 ^ n5287 ^ n652 ;
  assign n6925 = n966 & n4838 ;
  assign n6926 = n6925 ^ n1409 ^ 1'b0 ;
  assign n6927 = ~n2460 & n6926 ;
  assign n6931 = n6930 ^ n6927 ^ 1'b0 ;
  assign n6932 = ~n129 & n6931 ;
  assign n6933 = n2068 ^ n2064 ^ n1439 ;
  assign n6934 = n4788 & n6896 ;
  assign n6935 = n5255 & n6934 ;
  assign n6936 = n3074 ^ n1325 ^ 1'b0 ;
  assign n6937 = n6936 ^ n4552 ^ 1'b0 ;
  assign n6938 = ~n1500 & n1880 ;
  assign n6939 = n596 & ~n6615 ;
  assign n6940 = ~n5056 & n6547 ;
  assign n6941 = n5513 ^ n4781 ^ 1'b0 ;
  assign n6942 = n793 | n6941 ;
  assign n6943 = ~n705 & n6037 ;
  assign n6944 = n6943 ^ n168 ^ 1'b0 ;
  assign n6945 = n6944 ^ n3405 ^ 1'b0 ;
  assign n6946 = n4257 | n6945 ;
  assign n6947 = n2526 & n6946 ;
  assign n6948 = n6947 ^ n4746 ^ 1'b0 ;
  assign n6949 = n1730 | n6080 ;
  assign n6950 = n75 | n4048 ;
  assign n6951 = n460 | n6950 ;
  assign n6952 = n6951 ^ n727 ^ 1'b0 ;
  assign n6953 = n6272 & ~n6952 ;
  assign n6954 = ~n182 & n6377 ;
  assign n6955 = n6953 & n6954 ;
  assign n6956 = n3270 ^ n442 ^ 1'b0 ;
  assign n6957 = ~n6779 & n6956 ;
  assign n6958 = n777 & ~n1943 ;
  assign n6964 = n2500 ^ n1127 ^ 1'b0 ;
  assign n6960 = n55 & ~n1479 ;
  assign n6961 = n759 & n6960 ;
  assign n6962 = n6961 ^ n507 ^ 1'b0 ;
  assign n6963 = n2059 & ~n6962 ;
  assign n6959 = n372 & ~n3756 ;
  assign n6965 = n6964 ^ n6963 ^ n6959 ;
  assign n6966 = n2315 ^ n2187 ^ n1931 ;
  assign n6967 = n6966 ^ n2039 ^ 1'b0 ;
  assign n6968 = n556 ^ n375 ^ 1'b0 ;
  assign n6969 = n6967 | n6968 ;
  assign n6970 = n6969 ^ n2899 ^ 1'b0 ;
  assign n6971 = n6207 ^ n5386 ^ 1'b0 ;
  assign n6972 = n5749 ^ n4361 ^ n3936 ;
  assign n6973 = n1523 & n1810 ;
  assign n6974 = ( n423 & ~n2936 ) | ( n423 & n6586 ) | ( ~n2936 & n6586 ) ;
  assign n6975 = n86 | n2422 ;
  assign n6976 = n6975 ^ n1480 ^ 1'b0 ;
  assign n6977 = n6976 ^ n1944 ^ 1'b0 ;
  assign n6978 = n6048 & n6977 ;
  assign n6979 = n6974 & n6978 ;
  assign n6980 = n313 | n2604 ;
  assign n6981 = n6980 ^ n6150 ^ 1'b0 ;
  assign n6982 = n4227 ^ n3069 ^ 1'b0 ;
  assign n6983 = n6981 & ~n6982 ;
  assign n6984 = n949 & ~n3178 ;
  assign n6985 = ~n2107 & n6984 ;
  assign n6986 = ~n1431 & n6985 ;
  assign n6988 = n1138 ^ n928 ^ 1'b0 ;
  assign n6989 = n1328 | n6988 ;
  assign n6987 = ~n652 & n1502 ;
  assign n6990 = n6989 ^ n6987 ^ 1'b0 ;
  assign n6991 = n5988 & n6990 ;
  assign n6992 = ~n1345 & n6991 ;
  assign n6993 = n6992 ^ n2459 ^ 1'b0 ;
  assign n6994 = n4422 | n6993 ;
  assign n6995 = n6553 ^ n4902 ^ 1'b0 ;
  assign n6996 = n6995 ^ n5225 ^ 1'b0 ;
  assign n6997 = n5054 & ~n6996 ;
  assign n6998 = n6994 | n6997 ;
  assign n7000 = n4903 ^ n926 ^ 1'b0 ;
  assign n7001 = ~n605 & n7000 ;
  assign n6999 = n804 | n1254 ;
  assign n7002 = n7001 ^ n6999 ^ 1'b0 ;
  assign n7003 = n2201 | n7002 ;
  assign n7004 = n3188 ^ n300 ^ 1'b0 ;
  assign n7005 = ~n7003 & n7004 ;
  assign n7006 = n2422 & n5718 ;
  assign n7007 = n32 & n2694 ;
  assign n7008 = n6773 & ~n7007 ;
  assign n7009 = n2189 & n4984 ;
  assign n7010 = n7007 ^ n5853 ^ 1'b0 ;
  assign n7011 = ~n7009 & n7010 ;
  assign n7012 = n1888 | n4618 ;
  assign n7013 = n7011 | n7012 ;
  assign n7014 = n6185 ^ n2836 ^ 1'b0 ;
  assign n7015 = n3258 & n7014 ;
  assign n7016 = ~n1492 & n2430 ;
  assign n7017 = ~n7015 & n7016 ;
  assign n7018 = n4793 ^ n3100 ^ 1'b0 ;
  assign n7019 = ~n7017 & n7018 ;
  assign n7020 = n7019 ^ n1161 ^ 1'b0 ;
  assign n7021 = ~n6228 & n7020 ;
  assign n7022 = n4193 ^ n3679 ^ 1'b0 ;
  assign n7023 = n1537 & ~n7022 ;
  assign n7024 = ~n322 & n4976 ;
  assign n7025 = n6291 & n7021 ;
  assign n7026 = n7025 ^ n3355 ^ 1'b0 ;
  assign n7031 = n931 ^ n875 ^ 1'b0 ;
  assign n7028 = n1252 & n3440 ;
  assign n7029 = n7028 ^ n5802 ^ 1'b0 ;
  assign n7027 = ~n2141 & n4115 ;
  assign n7030 = n7029 ^ n7027 ^ 1'b0 ;
  assign n7032 = n7031 ^ n7030 ^ 1'b0 ;
  assign n7033 = n6781 ^ n5401 ^ 1'b0 ;
  assign n7037 = ~n3088 & n4024 ;
  assign n7038 = n7037 ^ n1394 ^ 1'b0 ;
  assign n7036 = n300 & n2433 ;
  assign n7039 = n7038 ^ n7036 ^ 1'b0 ;
  assign n7034 = n1174 & n2850 ;
  assign n7035 = n4192 & ~n7034 ;
  assign n7040 = n7039 ^ n7035 ^ 1'b0 ;
  assign n7041 = n3068 & ~n4180 ;
  assign n7042 = n2476 & n2694 ;
  assign n7043 = n7042 ^ n1234 ^ 1'b0 ;
  assign n7044 = n7043 ^ n6028 ^ 1'b0 ;
  assign n7045 = n5545 & n7044 ;
  assign n7046 = n2934 & n7045 ;
  assign n7047 = ~n587 & n5985 ;
  assign n7048 = n2097 ^ n216 ^ 1'b0 ;
  assign n7049 = n7048 ^ n3663 ^ 1'b0 ;
  assign n7050 = n4704 & ~n4742 ;
  assign n7051 = n7050 ^ n2714 ^ 1'b0 ;
  assign n7052 = n1473 & n1820 ;
  assign n7053 = ~n3354 & n5134 ;
  assign n7054 = n4976 ^ n2441 ^ 1'b0 ;
  assign n7055 = n627 & n3560 ;
  assign n7056 = n664 ^ n659 ^ 1'b0 ;
  assign n7057 = n6672 ^ n759 ^ 1'b0 ;
  assign n7060 = n547 | n2210 ;
  assign n7061 = n7060 ^ n3204 ^ 1'b0 ;
  assign n7058 = n3702 & n5425 ;
  assign n7059 = n7058 ^ n6097 ^ 1'b0 ;
  assign n7062 = n7061 ^ n7059 ^ 1'b0 ;
  assign n7063 = n5222 & ~n7062 ;
  assign n7065 = n25 & ~n4536 ;
  assign n7066 = n7065 ^ n2096 ^ 1'b0 ;
  assign n7064 = n3093 & n5454 ;
  assign n7067 = n7066 ^ n7064 ^ 1'b0 ;
  assign n7069 = ~n216 & n2326 ;
  assign n7068 = n4599 | n5978 ;
  assign n7070 = n7069 ^ n7068 ^ 1'b0 ;
  assign n7071 = n170 & ~n5856 ;
  assign n7072 = n1163 ^ n1139 ^ 1'b0 ;
  assign n7074 = n4840 ^ n2597 ^ 1'b0 ;
  assign n7073 = n987 | n6325 ;
  assign n7075 = n7074 ^ n7073 ^ 1'b0 ;
  assign n7076 = ~n1324 & n2849 ;
  assign n7077 = n7076 ^ n6912 ^ 1'b0 ;
  assign n7078 = n4093 ^ n1926 ^ 1'b0 ;
  assign n7079 = n5431 | n7078 ;
  assign n7080 = ~n128 & n3301 ;
  assign n7081 = ~n2603 & n4853 ;
  assign n7082 = n4845 ^ n4104 ^ 1'b0 ;
  assign n7083 = n2535 | n3504 ;
  assign n7084 = n6420 ^ n3244 ^ 1'b0 ;
  assign n7085 = n6175 & ~n7084 ;
  assign n7086 = ~n64 & n804 ;
  assign n7087 = n7086 ^ n3120 ^ 1'b0 ;
  assign n7088 = n7087 ^ n2107 ^ 1'b0 ;
  assign n7089 = n1325 | n7088 ;
  assign n7090 = n7089 ^ n390 ^ 1'b0 ;
  assign n7091 = n1227 ^ n418 ^ 1'b0 ;
  assign n7092 = n7091 ^ n1152 ^ 1'b0 ;
  assign n7093 = n2254 | n7092 ;
  assign n7094 = n489 & n759 ;
  assign n7095 = ~n1008 & n7094 ;
  assign n7096 = n177 & ~n7095 ;
  assign n7097 = n1216 & n7096 ;
  assign n7098 = n7093 & n7097 ;
  assign n7099 = n1630 & n4140 ;
  assign n7100 = n6753 & n7099 ;
  assign n7101 = n2175 & n4966 ;
  assign n7102 = n1763 & ~n5688 ;
  assign n7103 = n1431 | n7102 ;
  assign n7104 = n952 | n1183 ;
  assign n7105 = ~n7103 & n7104 ;
  assign n7106 = n3331 ^ n1928 ^ 1'b0 ;
  assign n7107 = ~n216 & n1396 ;
  assign n7108 = ~n7106 & n7107 ;
  assign n7109 = n154 & ~n1205 ;
  assign n7110 = n6040 ^ n2998 ^ 1'b0 ;
  assign n7111 = ~n216 & n3037 ;
  assign n7112 = n2623 & n4199 ;
  assign n7113 = ~n186 & n7112 ;
  assign n7114 = n832 ^ n622 ^ 1'b0 ;
  assign n7115 = n7019 ^ n6537 ^ 1'b0 ;
  assign n7116 = ~n1056 & n2137 ;
  assign n7117 = n1142 & n7116 ;
  assign n7118 = n7117 ^ n86 ^ 1'b0 ;
  assign n7119 = n1484 ^ n1230 ^ 1'b0 ;
  assign n7120 = ( n114 & ~n775 ) | ( n114 & n3210 ) | ( ~n775 & n3210 ) ;
  assign n7121 = n4666 | n7120 ;
  assign n7122 = n96 ^ x0 ^ 1'b0 ;
  assign n7123 = n178 & ~n1668 ;
  assign n7124 = n4436 | n5217 ;
  assign n7128 = n1522 | n2267 ;
  assign n7125 = n984 & n2489 ;
  assign n7126 = n4225 & n7125 ;
  assign n7127 = n1188 | n7126 ;
  assign n7129 = n7128 ^ n7127 ^ 1'b0 ;
  assign n7130 = n273 | n7129 ;
  assign n7131 = n2495 | n3314 ;
  assign n7132 = n7131 ^ n5793 ^ 1'b0 ;
  assign n7133 = n2141 ^ n1396 ^ 1'b0 ;
  assign n7134 = n6185 & ~n7133 ;
  assign n7135 = ~n4331 & n6519 ;
  assign n7136 = n2566 ^ n178 ^ 1'b0 ;
  assign n7137 = n2988 | n7136 ;
  assign n7138 = n1956 ^ n1166 ^ 1'b0 ;
  assign n7139 = n7138 ^ n3074 ^ 1'b0 ;
  assign n7140 = n6063 ^ n2640 ^ 1'b0 ;
  assign n7141 = n4956 & ~n5004 ;
  assign n7142 = n3263 & n7141 ;
  assign n7143 = n2513 & ~n7142 ;
  assign n7144 = n3180 & n4264 ;
  assign n7145 = n1036 & n5724 ;
  assign n7146 = n748 & ~n4171 ;
  assign n7147 = n5995 ^ n5723 ^ 1'b0 ;
  assign n7148 = n741 & ~n3561 ;
  assign n7149 = n5808 ^ n58 ^ 1'b0 ;
  assign n7150 = n4209 | n7106 ;
  assign n7151 = n291 | n7150 ;
  assign n7152 = ~n2178 & n7151 ;
  assign n7153 = n6764 & n7152 ;
  assign n7154 = ~n2193 & n3144 ;
  assign n7155 = ~n194 & n4779 ;
  assign n7156 = ~n5336 & n7155 ;
  assign n7157 = n185 & ~n5238 ;
  assign n7158 = n3068 ^ n1879 ^ 1'b0 ;
  assign n7159 = ~n7157 & n7158 ;
  assign n7160 = ~n3581 & n4869 ;
  assign n7166 = n291 & n540 ;
  assign n7167 = ~n540 & n7166 ;
  assign n7168 = n290 | n7167 ;
  assign n7169 = n7167 & ~n7168 ;
  assign n7172 = ~n212 & n359 ;
  assign n7173 = ~n359 & n7172 ;
  assign n7170 = n43 & n153 ;
  assign n7171 = ~n43 & n7170 ;
  assign n7174 = n7173 ^ n7171 ^ 1'b0 ;
  assign n7175 = n7169 & n7174 ;
  assign n7161 = n280 & n292 ;
  assign n7162 = ~n499 & n629 ;
  assign n7163 = ~n629 & n7162 ;
  assign n7164 = n7161 | n7163 ;
  assign n7165 = n7161 & ~n7164 ;
  assign n7176 = n7175 ^ n7165 ^ 1'b0 ;
  assign n7177 = n7176 ^ n3789 ^ 1'b0 ;
  assign n7178 = n7160 & n7177 ;
  assign n7179 = ( n175 & ~n2695 ) | ( n175 & n4412 ) | ( ~n2695 & n4412 ) ;
  assign n7180 = n4409 & ~n7179 ;
  assign n7181 = n878 ^ n354 ^ 1'b0 ;
  assign n7182 = n4374 ^ n924 ^ 1'b0 ;
  assign n7183 = n7182 ^ n4253 ^ n1227 ;
  assign n7184 = ~n1452 & n3063 ;
  assign n7185 = n7184 ^ n6498 ^ 1'b0 ;
  assign n7186 = n488 | n6826 ;
  assign n7187 = n800 & n804 ;
  assign n7188 = n1826 & ~n7187 ;
  assign n7189 = n7188 ^ n4767 ^ 1'b0 ;
  assign n7190 = n323 & ~n7189 ;
  assign n7191 = ~n1914 & n7190 ;
  assign n7195 = n157 & ~n4745 ;
  assign n7192 = n1573 ^ n1045 ^ 1'b0 ;
  assign n7193 = n6055 | n7192 ;
  assign n7194 = ~n2930 & n7193 ;
  assign n7196 = n7195 ^ n7194 ^ 1'b0 ;
  assign n7197 = n4591 | n7196 ;
  assign n7198 = n55 | n3178 ;
  assign n7199 = n2480 | n7198 ;
  assign n7200 = n6160 & n7199 ;
  assign n7201 = ~n6966 & n7200 ;
  assign n7202 = n7201 ^ n5971 ^ 1'b0 ;
  assign n7203 = n461 | n7202 ;
  assign n7208 = n3169 ^ n673 ^ 1'b0 ;
  assign n7209 = n7208 ^ n2769 ^ 1'b0 ;
  assign n7210 = n2637 & ~n7209 ;
  assign n7204 = n1377 & n2142 ;
  assign n7205 = n7204 ^ n3459 ^ 1'b0 ;
  assign n7206 = n7205 ^ n128 ^ 1'b0 ;
  assign n7207 = n3137 & ~n7206 ;
  assign n7211 = n7210 ^ n7207 ^ 1'b0 ;
  assign n7212 = n6165 & n7211 ;
  assign n7213 = n6277 & n7212 ;
  assign n7214 = n7213 ^ n927 ^ 1'b0 ;
  assign n7218 = n3412 | n3781 ;
  assign n7219 = n3412 & ~n7218 ;
  assign n7215 = ~n96 & n2707 ;
  assign n7216 = ~n3343 & n7215 ;
  assign n7217 = n7216 ^ n4098 ^ 1'b0 ;
  assign n7220 = n7219 ^ n7217 ^ 1'b0 ;
  assign n7221 = n153 & ~n3406 ;
  assign n7222 = n7220 | n7221 ;
  assign n7223 = n3985 ^ n1567 ^ 1'b0 ;
  assign n7224 = n1372 ^ n506 ^ 1'b0 ;
  assign n7225 = n3560 & ~n7224 ;
  assign n7226 = n3939 & n7225 ;
  assign n7227 = ~n7223 & n7226 ;
  assign n7228 = n7227 ^ n1125 ^ 1'b0 ;
  assign n7229 = n1162 | n7228 ;
  assign n7230 = x2 & n476 ;
  assign n7231 = n7230 ^ n3054 ^ 1'b0 ;
  assign n7232 = n364 & n894 ;
  assign n7233 = n7231 & n7232 ;
  assign n7234 = n1169 ^ n128 ^ 1'b0 ;
  assign n7235 = n5269 | n6509 ;
  assign n7236 = n92 & ~n7235 ;
  assign n7237 = n1425 ^ n1267 ^ 1'b0 ;
  assign n7238 = ~n2012 & n7237 ;
  assign n7239 = n7238 ^ n4267 ^ 1'b0 ;
  assign n7240 = n6766 ^ n3490 ^ 1'b0 ;
  assign n7241 = ~n384 & n1950 ;
  assign n7243 = x0 | n1839 ;
  assign n7244 = n7243 ^ n2690 ^ 1'b0 ;
  assign n7242 = n556 | n4254 ;
  assign n7245 = n7244 ^ n7242 ^ 1'b0 ;
  assign n7246 = n7245 ^ n194 ^ 1'b0 ;
  assign n7247 = ~n7241 & n7246 ;
  assign n7248 = n3005 ^ n671 ^ 1'b0 ;
  assign n7249 = n236 | n7248 ;
  assign n7250 = n184 & ~n7249 ;
  assign n7254 = n2185 ^ n950 ^ 1'b0 ;
  assign n7255 = ~n2751 & n7254 ;
  assign n7256 = n468 & n7255 ;
  assign n7257 = n3635 & ~n7256 ;
  assign n7258 = n7257 ^ n5462 ^ 1'b0 ;
  assign n7251 = n247 | n1348 ;
  assign n7252 = ~n663 & n7251 ;
  assign n7253 = n117 & n7252 ;
  assign n7259 = n7258 ^ n7253 ^ 1'b0 ;
  assign n7260 = n4045 ^ n205 ^ 1'b0 ;
  assign n7261 = ~n2514 & n5199 ;
  assign n7262 = n2127 | n6818 ;
  assign n7263 = n191 | n7262 ;
  assign n7264 = n7263 ^ n4392 ^ 1'b0 ;
  assign n7265 = n765 ^ n732 ^ 1'b0 ;
  assign n7266 = n7265 ^ n1345 ^ 1'b0 ;
  assign n7267 = n698 & ~n7266 ;
  assign n7268 = n528 ^ n448 ^ 1'b0 ;
  assign n7269 = n7268 ^ n2322 ^ n495 ;
  assign n7270 = n7269 ^ n5706 ^ 1'b0 ;
  assign n7271 = n4267 & ~n7270 ;
  assign n7272 = ~n2316 & n7271 ;
  assign n7273 = n4488 ^ n1183 ^ 1'b0 ;
  assign n7274 = n7273 ^ n5133 ^ 1'b0 ;
  assign n7275 = n5174 & ~n7274 ;
  assign n7277 = n768 ^ n364 ^ 1'b0 ;
  assign n7276 = ~x0 & n863 ;
  assign n7278 = n7277 ^ n7276 ^ 1'b0 ;
  assign n7279 = n2510 & ~n6206 ;
  assign n7280 = ~x1 & n2537 ;
  assign n7281 = n7280 ^ n5973 ^ 1'b0 ;
  assign n7282 = ~n2003 & n5716 ;
  assign n7283 = n2203 ^ x1 ^ 1'b0 ;
  assign n7284 = n1624 & n2476 ;
  assign n7285 = n1479 ^ n263 ^ 1'b0 ;
  assign n7286 = ~n1709 & n2724 ;
  assign n7287 = n7286 ^ n4680 ^ 1'b0 ;
  assign n7288 = n7285 & ~n7287 ;
  assign n7291 = n2649 ^ n2027 ^ 1'b0 ;
  assign n7292 = n789 | n7291 ;
  assign n7293 = n3005 ^ n34 ^ 1'b0 ;
  assign n7294 = ~n7292 & n7293 ;
  assign n7289 = n1315 & n1914 ;
  assign n7290 = n7289 ^ n1363 ^ 1'b0 ;
  assign n7295 = n7294 ^ n7290 ^ 1'b0 ;
  assign n7296 = n5443 & ~n7295 ;
  assign n7297 = n1900 ^ n1250 ^ 1'b0 ;
  assign n7298 = n378 & n7297 ;
  assign n7299 = n7298 ^ n1431 ^ 1'b0 ;
  assign n7300 = n7299 ^ n1838 ^ 1'b0 ;
  assign n7301 = n3103 | n4987 ;
  assign n7302 = ~n788 & n2210 ;
  assign n7303 = ~n3762 & n7302 ;
  assign n7304 = ~n3211 & n4095 ;
  assign n7305 = n2067 & ~n7146 ;
  assign n7306 = n5444 | n6198 ;
  assign n7307 = n501 & ~n7306 ;
  assign n7308 = n1499 ^ n55 ^ 1'b0 ;
  assign n7309 = n869 & ~n7308 ;
  assign n7310 = n4710 & n7309 ;
  assign n7311 = ~n5681 & n7310 ;
  assign n7312 = n4217 & ~n5629 ;
  assign n7313 = n7312 ^ n5252 ^ 1'b0 ;
  assign n7314 = n906 | n3007 ;
  assign n7315 = n3945 & ~n7314 ;
  assign n7316 = n2500 | n7315 ;
  assign n7317 = n1968 ^ n471 ^ 1'b0 ;
  assign n7318 = n7317 ^ n4473 ^ 1'b0 ;
  assign n7319 = n713 | n7318 ;
  assign n7320 = n7319 ^ n5473 ^ 1'b0 ;
  assign n7321 = ~n1875 & n7320 ;
  assign n7322 = n870 & n7321 ;
  assign n7323 = n748 | n6865 ;
  assign n7324 = n581 & ~n4135 ;
  assign n7325 = n7324 ^ n2974 ^ 1'b0 ;
  assign n7326 = n675 & ~n7325 ;
  assign n7327 = n2307 | n7326 ;
  assign n7328 = n7282 ^ n466 ^ 1'b0 ;
  assign n7329 = n1466 ^ n19 ^ 1'b0 ;
  assign n7330 = n2499 & ~n7329 ;
  assign n7331 = n7330 ^ n6990 ^ 1'b0 ;
  assign n7332 = n391 | n2043 ;
  assign n7333 = n7332 ^ n3557 ^ 1'b0 ;
  assign n7334 = n404 ^ n218 ^ 1'b0 ;
  assign n7335 = n1252 & n7334 ;
  assign n7336 = n7335 ^ n226 ^ 1'b0 ;
  assign n7337 = n1367 & ~n1864 ;
  assign n7338 = ~n1745 & n7337 ;
  assign n7339 = n5837 | n7338 ;
  assign n7340 = n7339 ^ n1932 ^ 1'b0 ;
  assign n7341 = ~n3014 & n7340 ;
  assign n7342 = ~n3940 & n5584 ;
  assign n7343 = n6224 & n7342 ;
  assign n7344 = n665 | n6607 ;
  assign n7345 = n3131 & n7344 ;
  assign n7346 = n48 & n2987 ;
  assign n7347 = n3327 & n7346 ;
  assign n7348 = n7347 ^ n1386 ^ 1'b0 ;
  assign n7349 = n461 | n927 ;
  assign n7350 = n290 & ~n7349 ;
  assign n7351 = n3687 & ~n5334 ;
  assign n7352 = ~n6992 & n7351 ;
  assign n7353 = ( n5138 & ~n7350 ) | ( n5138 & n7352 ) | ( ~n7350 & n7352 ) ;
  assign n7354 = n229 ^ n169 ^ 1'b0 ;
  assign n7355 = x1 & ~n7354 ;
  assign n7356 = n290 & ~n5085 ;
  assign n7357 = n7356 ^ n296 ^ 1'b0 ;
  assign n7358 = ( n3469 & n7157 ) | ( n3469 & n7357 ) | ( n7157 & n7357 ) ;
  assign n7359 = n1631 & ~n5821 ;
  assign n7360 = n6174 & n7359 ;
  assign n7361 = n4274 ^ n3156 ^ 1'b0 ;
  assign n7362 = n6079 & n7361 ;
  assign n7363 = ~n6839 & n7362 ;
  assign n7364 = n1048 ^ n938 ^ 1'b0 ;
  assign n7365 = n2235 & n3632 ;
  assign n7366 = n445 & ~n2348 ;
  assign n7367 = n7366 ^ n1174 ^ 1'b0 ;
  assign n7368 = n7365 & n7367 ;
  assign n7369 = n5355 ^ n3570 ^ 1'b0 ;
  assign n7370 = n1945 & n2768 ;
  assign n7371 = n7310 & n7370 ;
  assign n7372 = n1674 ^ n665 ^ 1'b0 ;
  assign n7373 = n3100 & n7372 ;
  assign n7374 = n4250 & ~n7373 ;
  assign n7375 = n483 & ~n5975 ;
  assign n7376 = n1100 & ~n6773 ;
  assign n7377 = n737 & n3627 ;
  assign n7380 = ~n2850 & n5152 ;
  assign n7378 = n2446 | n7155 ;
  assign n7379 = n2988 & n7378 ;
  assign n7381 = n7380 ^ n7379 ^ 1'b0 ;
  assign n7382 = n4462 ^ n4437 ^ 1'b0 ;
  assign n7383 = n4670 | n7382 ;
  assign n7387 = n1695 & ~n7201 ;
  assign n7388 = n7387 ^ n83 ^ 1'b0 ;
  assign n7384 = n6552 ^ n4106 ^ n2148 ;
  assign n7385 = n7384 ^ n1836 ^ 1'b0 ;
  assign n7386 = n185 | n7385 ;
  assign n7389 = n7388 ^ n7386 ^ 1'b0 ;
  assign n7390 = n2704 & n7389 ;
  assign n7391 = n573 & n2426 ;
  assign n7392 = n1676 & n7391 ;
  assign n7393 = n7083 ^ n5465 ^ 1'b0 ;
  assign n7394 = ~n2948 & n7393 ;
  assign n7395 = n319 | n3602 ;
  assign n7396 = n16 & ~n390 ;
  assign n7397 = n7396 ^ n257 ^ 1'b0 ;
  assign n7398 = n3284 ^ n1203 ^ 1'b0 ;
  assign n7399 = n6903 & ~n7398 ;
  assign n7400 = n7399 ^ n7126 ^ 1'b0 ;
  assign n7404 = n3244 & ~n5549 ;
  assign n7405 = n1407 | n7404 ;
  assign n7406 = n7405 ^ n3203 ^ 1'b0 ;
  assign n7401 = n2034 | n3355 ;
  assign n7402 = ~n5336 & n7401 ;
  assign n7403 = n7402 ^ n2041 ^ 1'b0 ;
  assign n7407 = n7406 ^ n7403 ^ 1'b0 ;
  assign n7408 = ~n497 & n3044 ;
  assign n7409 = n1155 & ~n1447 ;
  assign n7410 = n7409 ^ n553 ^ 1'b0 ;
  assign n7411 = n2681 ^ n2542 ^ 1'b0 ;
  assign n7412 = n234 & ~n5607 ;
  assign n7413 = n3767 & ~n7412 ;
  assign n7414 = n5192 ^ n949 ^ 1'b0 ;
  assign n7415 = ~n316 & n7414 ;
  assign n7416 = ~n246 & n727 ;
  assign n7417 = ( n64 & ~n402 ) | ( n64 & n7416 ) | ( ~n402 & n7416 ) ;
  assign n7418 = ~n274 & n5700 ;
  assign n7419 = n731 & ~n1630 ;
  assign n7420 = n7251 | n7419 ;
  assign n7421 = ~n2167 & n7420 ;
  assign n7424 = n3186 ^ n2010 ^ 1'b0 ;
  assign n7422 = n5024 ^ n419 ^ n161 ;
  assign n7423 = n2425 & ~n7422 ;
  assign n7425 = n7424 ^ n7423 ^ 1'b0 ;
  assign n7426 = ~n7421 & n7425 ;
  assign n7427 = n2194 & n7426 ;
  assign n7428 = n697 & ~n2736 ;
  assign n7429 = n7428 ^ n2201 ^ n1793 ;
  assign n7430 = n1538 | n3504 ;
  assign n7431 = n107 & ~n7111 ;
  assign n7432 = n5900 ^ n1437 ^ 1'b0 ;
  assign n7433 = n1529 & n2426 ;
  assign n7434 = ~n5653 & n7433 ;
  assign n7435 = ~n5145 & n7434 ;
  assign n7436 = ~n4563 & n7435 ;
  assign n7437 = n928 ^ n726 ^ 1'b0 ;
  assign n7438 = n7436 | n7437 ;
  assign n7439 = n1772 ^ n1192 ^ 1'b0 ;
  assign n7440 = n6742 ^ n599 ^ 1'b0 ;
  assign n7441 = n5014 ^ n1234 ^ 1'b0 ;
  assign n7442 = n1638 | n7441 ;
  assign n7443 = n1051 ^ n294 ^ 1'b0 ;
  assign n7444 = n1964 | n2080 ;
  assign n7445 = n4357 ^ n685 ^ 1'b0 ;
  assign n7446 = n7445 ^ n246 ^ 1'b0 ;
  assign n7447 = n7444 & ~n7446 ;
  assign n7448 = n837 | n7447 ;
  assign n7449 = ~n4004 & n5833 ;
  assign n7450 = n1533 & ~n2316 ;
  assign n7451 = ( n1086 & n7449 ) | ( n1086 & ~n7450 ) | ( n7449 & ~n7450 ) ;
  assign n7452 = n7451 ^ n2835 ^ 1'b0 ;
  assign n7453 = n4243 ^ n2873 ^ 1'b0 ;
  assign n7454 = n7300 | n7453 ;
  assign n7455 = ~n1464 & n2491 ;
  assign n7456 = ~n3120 & n7455 ;
  assign n7457 = n580 & ~n1426 ;
  assign n7458 = ( n406 & n1404 ) | ( n406 & ~n7457 ) | ( n1404 & ~n7457 ) ;
  assign n7459 = n7458 ^ n2244 ^ 1'b0 ;
  assign n7460 = n3591 | n4407 ;
  assign n7461 = n7460 ^ n75 ^ 1'b0 ;
  assign n7462 = n159 & n2808 ;
  assign n7463 = n6099 ^ n246 ^ 1'b0 ;
  assign n7464 = n3846 & ~n7463 ;
  assign n7465 = n6074 ^ n926 ^ 1'b0 ;
  assign n7466 = n1976 ^ n997 ^ 1'b0 ;
  assign n7467 = n1060 | n7444 ;
  assign n7468 = n137 | n7467 ;
  assign n7469 = n7435 & n7468 ;
  assign n7470 = ~n7466 & n7469 ;
  assign n7471 = n7470 ^ n3621 ^ 1'b0 ;
  assign n7472 = n1662 | n6598 ;
  assign n7474 = ~n1065 & n1640 ;
  assign n7475 = n811 & n7474 ;
  assign n7473 = n691 | n5928 ;
  assign n7476 = n7475 ^ n7473 ^ 1'b0 ;
  assign n7477 = n7476 ^ n4166 ^ 1'b0 ;
  assign n7478 = n6376 ^ n4647 ^ 1'b0 ;
  assign n7479 = n7289 | n7478 ;
  assign n7480 = n475 & n1631 ;
  assign n7481 = n6014 | n7480 ;
  assign n7482 = n4155 & ~n6419 ;
  assign n7483 = n7481 & n7482 ;
  assign n7484 = n5922 ^ n1372 ^ 1'b0 ;
  assign n7485 = n2260 | n7484 ;
  assign n7486 = n7485 ^ n1472 ^ 1'b0 ;
  assign n7487 = ( n252 & ~n468 ) | ( n252 & n3314 ) | ( ~n468 & n3314 ) ;
  assign n7488 = n1645 | n5808 ;
  assign n7489 = n3579 | n4772 ;
  assign n7490 = n448 & ~n5445 ;
  assign n7491 = n7490 ^ n6370 ^ 1'b0 ;
  assign n7492 = n495 & n1825 ;
  assign n7493 = n1668 & n2254 ;
  assign n7494 = n7493 ^ n3532 ^ 1'b0 ;
  assign n7495 = n7494 ^ n3223 ^ n1212 ;
  assign n7496 = n6146 | n7495 ;
  assign n7497 = n7492 & ~n7496 ;
  assign n7498 = n5382 ^ n1250 ^ 1'b0 ;
  assign n7499 = n1358 & n7498 ;
  assign n7500 = n3980 & n7499 ;
  assign n7501 = n622 & ~n5338 ;
  assign n7502 = n1934 & ~n2068 ;
  assign n7510 = n295 | n1002 ;
  assign n7503 = n5856 ^ n4383 ^ 1'b0 ;
  assign n7506 = n1571 | n3883 ;
  assign n7504 = n2431 ^ n1033 ^ 1'b0 ;
  assign n7505 = n2062 & ~n7504 ;
  assign n7507 = n7506 ^ n7505 ^ 1'b0 ;
  assign n7508 = ~n7503 & n7507 ;
  assign n7509 = n553 & n7508 ;
  assign n7511 = n7510 ^ n7509 ^ 1'b0 ;
  assign n7512 = n4085 ^ n1800 ^ 1'b0 ;
  assign n7513 = n7511 & n7512 ;
  assign n7514 = ~n3211 & n7513 ;
  assign n7515 = n78 & ~n1796 ;
  assign n7516 = n7515 ^ n1530 ^ 1'b0 ;
  assign n7517 = n7516 ^ n6950 ^ 1'b0 ;
  assign n7518 = n632 & n7517 ;
  assign n7519 = n5049 & n7518 ;
  assign n7520 = n7519 ^ n7225 ^ 1'b0 ;
  assign n7521 = n3152 ^ n592 ^ 1'b0 ;
  assign n7522 = n4680 | n7521 ;
  assign n7527 = n3985 & n6408 ;
  assign n7528 = ~n2779 & n7527 ;
  assign n7529 = n3270 & ~n7528 ;
  assign n7523 = n6809 ^ n6447 ^ 1'b0 ;
  assign n7524 = n6398 & n7523 ;
  assign n7525 = x1 & n7524 ;
  assign n7526 = n5330 & n7525 ;
  assign n7530 = n7529 ^ n7526 ^ 1'b0 ;
  assign n7531 = ~n7522 & n7530 ;
  assign n7532 = n3853 ^ n381 ^ 1'b0 ;
  assign n7533 = n1151 ^ n55 ^ 1'b0 ;
  assign n7534 = n637 | n7533 ;
  assign n7535 = n7534 ^ n6489 ^ 1'b0 ;
  assign n7536 = n3211 ^ n2067 ^ 1'b0 ;
  assign n7537 = n1880 | n7536 ;
  assign n7539 = n2805 ^ n2298 ^ 1'b0 ;
  assign n7540 = n7539 ^ n6154 ^ n4643 ;
  assign n7538 = ~n3104 & n5005 ;
  assign n7541 = n7540 ^ n7538 ^ 1'b0 ;
  assign n7542 = n7537 | n7541 ;
  assign n7543 = n3001 ^ n2284 ^ 1'b0 ;
  assign n7544 = n3192 & n5235 ;
  assign n7545 = n7544 ^ n3245 ^ 1'b0 ;
  assign n7546 = n169 & n1844 ;
  assign n7547 = n1161 & ~n1569 ;
  assign n7548 = n7547 ^ n1751 ^ 1'b0 ;
  assign n7549 = n1928 & n7548 ;
  assign n7550 = n7549 ^ n3361 ^ 1'b0 ;
  assign n7551 = n3110 ^ n2159 ^ n168 ;
  assign n7552 = n3688 & ~n7551 ;
  assign n7553 = n1816 ^ n1368 ^ 1'b0 ;
  assign n7554 = ~n1100 & n7357 ;
  assign n7555 = n7553 & ~n7554 ;
  assign n7560 = n938 & ~n5661 ;
  assign n7561 = ~n938 & n7560 ;
  assign n7556 = ~x5 & n666 ;
  assign n7557 = ~n666 & n7556 ;
  assign n7558 = n423 & n7557 ;
  assign n7559 = n6634 & n7558 ;
  assign n7562 = n7561 ^ n7559 ^ 1'b0 ;
  assign n7563 = n3559 & n6046 ;
  assign n7564 = n3476 ^ n1038 ^ 1'b0 ;
  assign n7565 = n257 & ~n3469 ;
  assign n7566 = n7565 ^ n352 ^ 1'b0 ;
  assign n7567 = n4203 & ~n5011 ;
  assign n7568 = ~n1194 & n7567 ;
  assign n7569 = n2958 ^ n694 ^ 1'b0 ;
  assign n7570 = n7569 ^ n4712 ^ 1'b0 ;
  assign n7571 = n1132 | n4990 ;
  assign n7572 = n4119 | n7571 ;
  assign n7573 = n7572 ^ n5559 ^ n1584 ;
  assign n7574 = n1355 | n7573 ;
  assign n7575 = n2966 ^ n2282 ^ 1'b0 ;
  assign n7576 = n7574 & n7575 ;
  assign n7577 = n1070 & ~n1629 ;
  assign n7578 = n4334 & n7577 ;
  assign n7579 = ~n390 & n526 ;
  assign n7580 = n1708 & n1878 ;
  assign n7581 = n4540 | n6944 ;
  assign n7582 = ~n1100 & n7581 ;
  assign n7583 = n489 & n5439 ;
  assign n7584 = n4004 & n7583 ;
  assign n7585 = n2279 & n6065 ;
  assign n7586 = n7585 ^ n1958 ^ 1'b0 ;
  assign n7587 = n1072 & ~n4443 ;
  assign n7588 = n6901 & n7587 ;
  assign n7589 = n5692 ^ n508 ^ 1'b0 ;
  assign n7590 = ~n1329 & n2131 ;
  assign n7591 = n7590 ^ n2865 ^ 1'b0 ;
  assign n7592 = n1358 & n7591 ;
  assign n7593 = n1192 & n7592 ;
  assign n7594 = n2873 ^ n98 ^ 1'b0 ;
  assign n7595 = n2462 | n2751 ;
  assign n7596 = n917 & ~n7595 ;
  assign n7597 = ~x2 & n7596 ;
  assign n7598 = n2637 ^ n1207 ^ 1'b0 ;
  assign n7599 = ~n7597 & n7598 ;
  assign n7600 = ~n4439 & n7599 ;
  assign n7601 = n2426 & n7600 ;
  assign n7602 = n2218 & n2461 ;
  assign n7603 = ~n475 & n7602 ;
  assign n7604 = n6916 ^ n3669 ^ 1'b0 ;
  assign n7605 = n3585 ^ n1763 ^ 1'b0 ;
  assign n7606 = n929 & n7431 ;
  assign n7607 = n7047 ^ n616 ^ 1'b0 ;
  assign n7608 = n565 & n4805 ;
  assign n7609 = n7608 ^ n1802 ^ 1'b0 ;
  assign n7610 = n817 ^ n86 ^ 1'b0 ;
  assign n7611 = n6194 & n7610 ;
  assign n7612 = n311 ^ n309 ^ 1'b0 ;
  assign n7613 = n4193 & n7612 ;
  assign n7614 = n7611 & n7613 ;
  assign n7615 = n3422 ^ n608 ^ 1'b0 ;
  assign n7616 = n6125 & ~n7615 ;
  assign n7617 = n3394 & n5123 ;
  assign n7618 = n3466 ^ n2435 ^ 1'b0 ;
  assign n7619 = n1005 & n7618 ;
  assign n7620 = n1060 & n6960 ;
  assign n7621 = n7197 & n7620 ;
  assign n7622 = n7421 ^ n1736 ^ 1'b0 ;
  assign n7623 = n3442 ^ n1968 ^ 1'b0 ;
  assign n7624 = n2633 & n6990 ;
  assign n7625 = n1127 & ~n7624 ;
  assign n7626 = n1206 | n4623 ;
  assign n7627 = ~n117 & n7626 ;
  assign n7628 = n4618 | n7586 ;
  assign n7629 = ~n1020 & n5920 ;
  assign n7630 = ~n5710 & n7629 ;
  assign n7631 = n2166 & ~n2388 ;
  assign n7632 = n7631 ^ n4281 ^ 1'b0 ;
  assign n7633 = ~n4718 & n4740 ;
  assign n7634 = n7633 ^ n4550 ^ 1'b0 ;
  assign n7635 = n2027 & n7634 ;
  assign n7636 = n3940 & n7635 ;
  assign n7637 = n1926 & n6722 ;
  assign n7638 = n2038 | n2569 ;
  assign n7639 = n4495 & ~n7638 ;
  assign n7640 = n3521 ^ n2730 ^ 1'b0 ;
  assign n7641 = n374 | n7640 ;
  assign n7642 = n27 & n4355 ;
  assign n7643 = n3492 ^ n238 ^ 1'b0 ;
  assign n7644 = n7642 & n7643 ;
  assign n7645 = n769 & n7644 ;
  assign n7646 = ~n3074 & n7645 ;
  assign n7647 = n1943 ^ n1192 ^ 1'b0 ;
  assign n7648 = n210 & ~n7647 ;
  assign n7649 = n2307 | n4424 ;
  assign n7650 = n7649 ^ n792 ^ 1'b0 ;
  assign n7651 = n894 & ~n1543 ;
  assign n7652 = n310 & n7651 ;
  assign n7653 = n4483 & ~n7652 ;
  assign n7654 = n7653 ^ n3519 ^ 1'b0 ;
  assign n7655 = n7654 ^ n1480 ^ 1'b0 ;
  assign n7656 = n1684 & ~n3046 ;
  assign n7657 = ~n2717 & n7656 ;
  assign n7658 = n1572 ^ n36 ^ 1'b0 ;
  assign n7665 = n6129 ^ n2607 ^ 1'b0 ;
  assign n7659 = n323 & ~n4426 ;
  assign n7660 = n3143 ^ n2096 ^ 1'b0 ;
  assign n7661 = n364 & ~n7660 ;
  assign n7662 = n7661 ^ n310 ^ 1'b0 ;
  assign n7663 = n3804 | n7662 ;
  assign n7664 = n7659 | n7663 ;
  assign n7666 = n7665 ^ n7664 ^ n2068 ;
  assign n7667 = n1541 ^ n793 ^ 1'b0 ;
  assign n7668 = n257 ^ n246 ^ 1'b0 ;
  assign n7669 = n119 | n2696 ;
  assign n7670 = n27 & ~n6575 ;
  assign n7671 = n5629 ^ n2008 ^ n791 ;
  assign n7672 = ~n5938 & n7671 ;
  assign n7673 = n5953 & n7672 ;
  assign n7674 = n2105 ^ n328 ^ 1'b0 ;
  assign n7677 = n2594 | n3464 ;
  assign n7678 = n17 & ~n7677 ;
  assign n7675 = n1388 ^ n1273 ^ 1'b0 ;
  assign n7676 = n1280 | n7675 ;
  assign n7679 = n7678 ^ n7676 ^ n788 ;
  assign n7680 = n710 & ~n754 ;
  assign n7681 = n7680 ^ n705 ^ 1'b0 ;
  assign n7682 = n2377 & n7681 ;
  assign n7683 = n7682 ^ n190 ^ 1'b0 ;
  assign n7684 = n3742 | n7683 ;
  assign n7685 = n1350 & n4549 ;
  assign n7686 = n4667 | n7685 ;
  assign n7687 = n7401 ^ n116 ^ 1'b0 ;
  assign n7688 = n7687 ^ n7285 ^ 1'b0 ;
  assign n7689 = n6562 & ~n7088 ;
  assign n7690 = ~n4657 & n5083 ;
  assign n7691 = n7690 ^ n736 ^ 1'b0 ;
  assign n7692 = n1585 & n3374 ;
  assign n7693 = n7692 ^ n2187 ^ 1'b0 ;
  assign n7694 = n7693 ^ n3423 ^ 1'b0 ;
  assign n7695 = n456 ^ n19 ^ 1'b0 ;
  assign n7696 = n1267 & n7695 ;
  assign n7697 = n6900 & n7696 ;
  assign n7698 = n3826 & ~n4326 ;
  assign n7699 = n6698 ^ n468 ^ 1'b0 ;
  assign n7700 = n7375 ^ n2932 ^ 1'b0 ;
  assign n7701 = n3101 ^ n3064 ^ 1'b0 ;
  assign n7702 = n1684 & n2022 ;
  assign n7703 = n55 & n4865 ;
  assign n7704 = n7703 ^ n3709 ^ 1'b0 ;
  assign n7705 = ~n2485 & n5119 ;
  assign n7706 = ~n7704 & n7705 ;
  assign n7707 = n3545 | n7706 ;
  assign n7708 = n1051 & ~n2080 ;
  assign n7709 = n1315 & n7708 ;
  assign n7710 = n1227 & n1802 ;
  assign n7711 = n7710 ^ n205 ^ 1'b0 ;
  assign n7712 = n7711 ^ n1476 ^ 1'b0 ;
  assign n7713 = n592 | n7712 ;
  assign n7714 = n557 & ~n7713 ;
  assign n7715 = n3405 & n6626 ;
  assign n7716 = n3746 ^ n1501 ^ 1'b0 ;
  assign n7717 = n4377 & ~n7716 ;
  assign n7718 = n227 & ~n7717 ;
  assign n7719 = n5222 & ~n7442 ;
  assign n7720 = n4268 & n7719 ;
  assign n7721 = n736 & n4927 ;
  assign n7722 = n7721 ^ n7088 ^ n6775 ;
  assign n7723 = n1587 & n5562 ;
  assign n7724 = n7723 ^ n7214 ^ 1'b0 ;
  assign n7725 = n419 & ~n4606 ;
  assign n7726 = n7725 ^ n3576 ^ 1'b0 ;
  assign n7727 = n5018 & ~n7726 ;
  assign n7728 = ~n862 & n7727 ;
  assign n7729 = n7192 ^ n141 ^ 1'b0 ;
  assign n7730 = n7592 & ~n7729 ;
  assign n7733 = n932 ^ n928 ^ 1'b0 ;
  assign n7734 = ~n1130 & n7733 ;
  assign n7735 = n7734 ^ n3732 ^ 1'b0 ;
  assign n7736 = n508 & ~n7735 ;
  assign n7737 = n3857 ^ n2437 ^ 1'b0 ;
  assign n7738 = n6914 & ~n7737 ;
  assign n7739 = n7736 & n7738 ;
  assign n7731 = n120 & ~n4979 ;
  assign n7732 = ~n5701 & n7731 ;
  assign n7740 = n7739 ^ n7732 ^ n5065 ;
  assign n7741 = ( n989 & n3816 ) | ( n989 & ~n6768 ) | ( n3816 & ~n6768 ) ;
  assign n7742 = n4106 ^ n721 ^ 1'b0 ;
  assign n7743 = n6433 | n7742 ;
  assign n7744 = n7741 & ~n7743 ;
  assign n7745 = n2239 ^ n1216 ^ 1'b0 ;
  assign n7746 = n2122 & ~n4478 ;
  assign n7747 = n366 & n2114 ;
  assign n7748 = ~n3287 & n7747 ;
  assign n7749 = ~n7746 & n7748 ;
  assign n7750 = n2509 ^ n1347 ^ 1'b0 ;
  assign n7751 = n5445 ^ n2432 ^ 1'b0 ;
  assign n7752 = n68 | n522 ;
  assign n7753 = n541 ^ n419 ^ 1'b0 ;
  assign n7754 = n2288 ^ n233 ^ 1'b0 ;
  assign n7755 = n7754 ^ n4873 ^ n3104 ;
  assign n7756 = n7753 | n7755 ;
  assign n7757 = n7752 & ~n7756 ;
  assign n7758 = n119 | n757 ;
  assign n7759 = n7758 ^ n3194 ^ 1'b0 ;
  assign n7760 = ~n200 & n7759 ;
  assign n7761 = n7757 & n7760 ;
  assign n7762 = n7751 & ~n7761 ;
  assign n7763 = n7750 & n7762 ;
  assign n7764 = n7749 & ~n7763 ;
  assign n7765 = ~n539 & n630 ;
  assign n7766 = n7124 & n7765 ;
  assign n7767 = n83 & n1771 ;
  assign n7768 = n7767 ^ n6464 ^ 1'b0 ;
  assign n7769 = n5180 & n7768 ;
  assign n7770 = n6249 ^ n291 ^ 1'b0 ;
  assign n7771 = n5856 ^ n151 ^ 1'b0 ;
  assign n7772 = ~n938 & n3886 ;
  assign n7773 = ~n7771 & n7772 ;
  assign n7774 = n7061 ^ n5123 ^ 1'b0 ;
  assign n7775 = n1431 & ~n7774 ;
  assign n7776 = n7775 ^ n6955 ^ 1'b0 ;
  assign n7777 = ~n3967 & n7776 ;
  assign n7778 = n3833 ^ n3620 ^ 1'b0 ;
  assign n7779 = ~n520 & n7778 ;
  assign n7780 = ~n75 & n1695 ;
  assign n7781 = n419 & ~n3207 ;
  assign n7782 = ~n7780 & n7781 ;
  assign n7783 = ~n7596 & n7782 ;
  assign n7784 = n7612 ^ n4740 ^ 1'b0 ;
  assign n7785 = n3697 & n5467 ;
  assign n7786 = ~n4799 & n7785 ;
  assign n7787 = n2107 | n7786 ;
  assign n7788 = n200 & n7787 ;
  assign n7789 = ~n2122 & n7788 ;
  assign n7792 = n2874 ^ n566 ^ 1'b0 ;
  assign n7790 = n37 & n527 ;
  assign n7791 = ~n5089 & n7790 ;
  assign n7793 = n7792 ^ n7791 ^ 1'b0 ;
  assign n7794 = n7789 | n7793 ;
  assign n7795 = n3325 & ~n7794 ;
  assign n7796 = n2733 ^ n142 ^ 1'b0 ;
  assign n7797 = n7796 ^ n430 ^ 1'b0 ;
  assign n7798 = n7797 ^ n2222 ^ 1'b0 ;
  assign n7799 = n7126 ^ n1571 ^ n129 ;
  assign n7800 = n6916 ^ n1559 ^ 1'b0 ;
  assign n7801 = n2064 | n3189 ;
  assign n7802 = n3748 | n7801 ;
  assign n7803 = n3396 ^ n2484 ^ 1'b0 ;
  assign n7804 = n1358 & n7803 ;
  assign n7805 = ~n979 & n7804 ;
  assign n7806 = ~n5041 & n7553 ;
  assign n7807 = n5706 ^ n4519 ^ 1'b0 ;
  assign n7808 = n161 & ~n2203 ;
  assign n7809 = n1003 ^ n583 ^ 1'b0 ;
  assign n7810 = n434 & n7809 ;
  assign n7811 = n311 | n1067 ;
  assign n7812 = n4529 & ~n7811 ;
  assign n7814 = n504 | n626 ;
  assign n7813 = n1280 & n4061 ;
  assign n7815 = n7814 ^ n7813 ^ 1'b0 ;
  assign n7816 = n785 | n7752 ;
  assign n7817 = n6260 & ~n7816 ;
  assign n7818 = n113 & ~n7817 ;
  assign n7819 = n4370 & n7818 ;
  assign n7820 = n2388 | n3138 ;
  assign n7821 = n7820 ^ n4488 ^ 1'b0 ;
  assign n7822 = n2769 & n2906 ;
  assign n7823 = n4098 | n7822 ;
  assign n7824 = n7821 & ~n7823 ;
  assign n7825 = n4098 ^ n384 ^ 1'b0 ;
  assign n7826 = n7825 ^ n3861 ^ 1'b0 ;
  assign n7827 = n4439 | n7826 ;
  assign n7828 = ~n117 & n156 ;
  assign n7829 = n117 & n7828 ;
  assign n7830 = ~n69 & n7829 ;
  assign n7831 = ~n212 & n7830 ;
  assign n7832 = n121 & n7831 ;
  assign n7833 = n80 & n7832 ;
  assign n7834 = n3187 & n7833 ;
  assign n7835 = n337 & n354 ;
  assign n7836 = ~n337 & n7835 ;
  assign n7837 = n7834 | n7836 ;
  assign n7838 = n32 | n318 ;
  assign n7839 = n32 & ~n7838 ;
  assign n7840 = n1186 & n7839 ;
  assign n7841 = n7840 ^ n540 ^ 1'b0 ;
  assign n7842 = n7841 ^ n404 ^ 1'b0 ;
  assign n7843 = n7837 & ~n7842 ;
  assign n7844 = ~n2303 & n3626 ;
  assign n7845 = n7654 ^ n744 ^ 1'b0 ;
  assign n7846 = n4468 ^ n1794 ^ 1'b0 ;
  assign n7847 = n7846 ^ n6150 ^ 1'b0 ;
  assign n7848 = n3744 & n7847 ;
  assign n7849 = n3985 ^ n1731 ^ 1'b0 ;
  assign n7850 = n7848 & n7849 ;
  assign n7851 = ~n7845 & n7850 ;
  assign n7852 = n196 & ~n640 ;
  assign n7853 = n92 & n7852 ;
  assign n7854 = n294 | n7853 ;
  assign n7855 = n7854 ^ n139 ^ 1'b0 ;
  assign n7856 = n2724 & n4955 ;
  assign n7857 = n117 & n3560 ;
  assign n7858 = n971 | n1329 ;
  assign n7860 = n400 | n2260 ;
  assign n7859 = n3978 ^ n2850 ^ 1'b0 ;
  assign n7861 = n7860 ^ n7859 ^ 1'b0 ;
  assign n7862 = n7858 & n7861 ;
  assign n7863 = n6655 ^ n97 ^ 1'b0 ;
  assign n7864 = n6619 & n6776 ;
  assign n7865 = n2996 ^ n758 ^ 1'b0 ;
  assign n7866 = n7865 ^ n1597 ^ 1'b0 ;
  assign n7867 = ( ~n5456 & n6971 ) | ( ~n5456 & n7866 ) | ( n6971 & n7866 ) ;
  assign n7868 = ~n755 & n966 ;
  assign n7869 = ~n2552 & n7868 ;
  assign n7870 = ~n2721 & n7869 ;
  assign n7872 = ( n754 & n787 ) | ( n754 & ~n2887 ) | ( n787 & ~n2887 ) ;
  assign n7871 = ~n2911 & n3887 ;
  assign n7873 = n7872 ^ n7871 ^ 1'b0 ;
  assign n7874 = n6023 ^ n810 ^ 1'b0 ;
  assign n7875 = n7873 | n7874 ;
  assign n7876 = n4169 & n6626 ;
  assign n7877 = n713 & n7876 ;
  assign n7878 = n310 & n7877 ;
  assign n7879 = n3806 ^ n3389 ^ 1'b0 ;
  assign n7880 = n7879 ^ n2835 ^ 1'b0 ;
  assign n7881 = ~n1835 & n2380 ;
  assign n7882 = ~n1989 & n7881 ;
  assign n7883 = ~n2349 & n5772 ;
  assign n7884 = n7882 & n7883 ;
  assign n7886 = n2067 ^ n1966 ^ n935 ;
  assign n7885 = ~n1781 & n1825 ;
  assign n7887 = n7886 ^ n7885 ^ 1'b0 ;
  assign n7888 = n3868 ^ n16 ^ 1'b0 ;
  assign n7889 = n1664 & n7888 ;
  assign n7890 = ~n1368 & n7889 ;
  assign n7901 = n3662 & ~n4622 ;
  assign n7898 = n2109 ^ n1629 ^ 1'b0 ;
  assign n7899 = n7898 ^ n3001 ^ 1'b0 ;
  assign n7893 = ~n3433 & n6277 ;
  assign n7894 = n7893 ^ n5787 ^ 1'b0 ;
  assign n7895 = n5787 | n7894 ;
  assign n7891 = ~n1907 & n2085 ;
  assign n7892 = n7891 ^ n2417 ^ 1'b0 ;
  assign n7896 = n7895 ^ n7892 ^ 1'b0 ;
  assign n7897 = n2082 & n7896 ;
  assign n7900 = n7899 ^ n7897 ^ 1'b0 ;
  assign n7902 = n7901 ^ n7900 ^ 1'b0 ;
  assign n7903 = n7902 ^ n2762 ^ 1'b0 ;
  assign n7904 = n1488 | n7903 ;
  assign n7905 = n417 & n2198 ;
  assign n7906 = n7905 ^ n3983 ^ 1'b0 ;
  assign n7907 = n6316 & ~n7906 ;
  assign n7908 = ( n562 & n1737 ) | ( n562 & n5394 ) | ( n1737 & n5394 ) ;
  assign n7909 = ~n333 & n7908 ;
  assign n7910 = ~n56 & n3810 ;
  assign n7911 = n6927 ^ n713 ^ 1'b0 ;
  assign n7912 = n3382 & n7911 ;
  assign n7913 = ~n2686 & n7912 ;
  assign n7914 = n284 & ~n7913 ;
  assign n7915 = n3621 & ~n7118 ;
  assign n7916 = ~n681 & n2058 ;
  assign n7917 = n7916 ^ n5507 ^ 1'b0 ;
  assign n7918 = n7917 ^ n934 ^ 1'b0 ;
  assign n7919 = n1394 & ~n1673 ;
  assign n7920 = n7919 ^ n4446 ^ 1'b0 ;
  assign n7921 = n1027 & ~n5866 ;
  assign n7922 = n608 | n1213 ;
  assign n7923 = n4746 ^ n645 ^ 1'b0 ;
  assign n7924 = n7923 ^ n975 ^ 1'b0 ;
  assign n7925 = ~n465 & n5425 ;
  assign n7926 = n5135 & n7925 ;
  assign n7927 = ( n715 & n2076 ) | ( n715 & n3013 ) | ( n2076 & n3013 ) ;
  assign n7928 = ~n6876 & n7927 ;
  assign n7929 = n764 & ~n1672 ;
  assign n7930 = ~n1658 & n7929 ;
  assign n7931 = n599 | n7930 ;
  assign n7932 = n7931 ^ n3993 ^ 1'b0 ;
  assign n7933 = n7932 ^ n7596 ^ 1'b0 ;
  assign n7934 = n7933 ^ n279 ^ 1'b0 ;
  assign n7935 = n2637 & n3154 ;
  assign n7936 = n180 & n476 ;
  assign n7937 = n7936 ^ n2550 ^ 1'b0 ;
  assign n7938 = n4458 | n7937 ;
  assign n7939 = n2244 & ~n2843 ;
  assign n7940 = n7938 & n7939 ;
  assign n7941 = n1026 ^ n216 ^ 1'b0 ;
  assign n7942 = ~n144 & n7941 ;
  assign n7943 = ~n5045 & n7942 ;
  assign n7944 = n1656 & ~n2567 ;
  assign n7945 = n385 & ~n1227 ;
  assign n7946 = n7945 ^ n322 ^ 1'b0 ;
  assign n7947 = n7944 | n7946 ;
  assign n7948 = n1135 | n1486 ;
  assign n7949 = ~n1560 & n1898 ;
  assign n7950 = n3192 & n7628 ;
  assign n7951 = ~n7949 & n7950 ;
  assign n7952 = n7524 ^ n4181 ^ 1'b0 ;
  assign n7953 = n506 | n2136 ;
  assign n7954 = n7953 ^ n3443 ^ 1'b0 ;
  assign n7955 = n2125 | n2288 ;
  assign n7956 = ~n221 & n4214 ;
  assign n7957 = n7956 ^ n43 ^ 1'b0 ;
  assign n7958 = n7955 & n7957 ;
  assign n7959 = ~n461 & n4395 ;
  assign n7960 = n69 & ~n3609 ;
  assign n7961 = n5357 ^ n205 ^ 1'b0 ;
  assign n7962 = n7960 & ~n7961 ;
  assign n7963 = n4639 ^ n2320 ^ 1'b0 ;
  assign n7964 = n7962 & n7963 ;
  assign n7965 = n7964 ^ n3512 ^ 1'b0 ;
  assign n7966 = n7416 ^ n4210 ^ 1'b0 ;
  assign n7967 = n6977 & n7966 ;
  assign n7968 = n5932 ^ n1492 ^ 1'b0 ;
  assign n7969 = n3693 ^ n2754 ^ 1'b0 ;
  assign n7970 = ~n857 & n6948 ;
  assign n7971 = n2269 ^ n2217 ^ 1'b0 ;
  assign n7972 = n6197 | n7971 ;
  assign n7973 = n7972 ^ n4869 ^ n83 ;
  assign n7974 = n5032 ^ n3669 ^ 1'b0 ;
  assign n7975 = n1106 | n7974 ;
  assign n7976 = ~n1479 & n3941 ;
  assign n7977 = ~n975 & n7976 ;
  assign n7978 = n1250 | n7977 ;
  assign n7979 = ~n1790 & n3214 ;
  assign n7980 = n7979 ^ n743 ^ 1'b0 ;
  assign n7981 = n4136 ^ n354 ^ 1'b0 ;
  assign n7982 = n688 & n1982 ;
  assign n7983 = n7982 ^ n1329 ^ 1'b0 ;
  assign n7984 = n1599 & n4981 ;
  assign n7985 = ~n2987 & n7871 ;
  assign n7986 = n7985 ^ n439 ^ 1'b0 ;
  assign n7987 = n2219 ^ n695 ^ 1'b0 ;
  assign n7988 = ~n646 & n1900 ;
  assign n7989 = n3325 & ~n7988 ;
  assign n7990 = n7989 ^ n30 ^ 1'b0 ;
  assign n7991 = n6787 ^ n2506 ^ 1'b0 ;
  assign n7992 = n1496 & n7779 ;
  assign n7993 = n4642 ^ n624 ^ 1'b0 ;
  assign n7994 = n1335 & ~n7993 ;
  assign n7995 = n3179 | n7994 ;
  assign n7996 = n1302 ^ n419 ^ 1'b0 ;
  assign n7997 = n3766 | n5638 ;
  assign n7998 = ~n4428 & n7997 ;
  assign n7999 = n3606 & n7251 ;
  assign n8000 = n7999 ^ n3392 ^ 1'b0 ;
  assign n8001 = n2732 ^ n448 ^ 1'b0 ;
  assign n8002 = n385 & ~n4422 ;
  assign n8003 = n1155 & n3858 ;
  assign n8004 = n8003 ^ n6434 ^ 1'b0 ;
  assign n8005 = n3707 ^ n1685 ^ 1'b0 ;
  assign n8006 = n1447 ^ n338 ^ 1'b0 ;
  assign n8007 = n1112 | n8006 ;
  assign n8008 = n6445 & ~n8007 ;
  assign n8009 = n8005 & ~n8008 ;
  assign n8010 = n3509 & n8009 ;
  assign n8011 = n2994 & ~n4421 ;
  assign n8012 = n592 & ~n5085 ;
  assign n8013 = n5790 | n8012 ;
  assign n8014 = n1730 | n8013 ;
  assign n8015 = n1550 | n8014 ;
  assign n8016 = n1977 & n2205 ;
  assign n8017 = n7573 ^ n6399 ^ 1'b0 ;
  assign n8018 = n8016 & ~n8017 ;
  assign n8019 = ~n125 & n539 ;
  assign n8020 = n862 & ~n6740 ;
  assign n8021 = ~n4574 & n8020 ;
  assign n8022 = n8021 ^ n5761 ^ 1'b0 ;
  assign n8023 = x9 & n1737 ;
  assign n8024 = n8023 ^ n527 ^ 1'b0 ;
  assign n8025 = n38 & n3284 ;
  assign n8026 = n8025 ^ n5823 ^ 1'b0 ;
  assign n8027 = ~n8024 & n8026 ;
  assign n8028 = ~n3167 & n8027 ;
  assign n8029 = n1491 & ~n3617 ;
  assign n8030 = n8029 ^ n5285 ^ 1'b0 ;
  assign n8031 = n4590 ^ n1902 ^ 1'b0 ;
  assign n8032 = n423 & n5926 ;
  assign n8033 = ~n2573 & n8032 ;
  assign n8034 = n2394 & ~n8033 ;
  assign n8035 = ~n880 & n3078 ;
  assign n8036 = n8035 ^ n7669 ^ 1'b0 ;
  assign n8037 = ~n627 & n6438 ;
  assign n8038 = n3803 ^ n1602 ^ 1'b0 ;
  assign n8039 = n5986 & n8038 ;
  assign n8040 = n4754 ^ n75 ^ 1'b0 ;
  assign n8041 = n1771 ^ n309 ^ 1'b0 ;
  assign n8042 = n8041 ^ n7254 ^ 1'b0 ;
  assign n8043 = n2116 ^ n1757 ^ 1'b0 ;
  assign n8044 = n8042 | n8043 ;
  assign n8045 = ~n4491 & n6125 ;
  assign n8046 = ~n6907 & n8045 ;
  assign n8047 = n4207 | n8046 ;
  assign n8048 = n1310 ^ n1266 ^ 1'b0 ;
  assign n8049 = n3504 | n8048 ;
  assign n8050 = ~n6645 & n8049 ;
  assign n8051 = n5025 ^ n2236 ^ 1'b0 ;
  assign n8052 = n622 & n8051 ;
  assign n8053 = n532 & ~n8052 ;
  assign n8054 = ~n60 & n6411 ;
  assign n8055 = ~n907 & n2513 ;
  assign n8056 = n8055 ^ n1360 ^ 1'b0 ;
  assign n8057 = n8056 ^ n599 ^ 1'b0 ;
  assign n8058 = n1613 & n2974 ;
  assign n8059 = n4641 & n8058 ;
  assign n8060 = ~n2302 & n7780 ;
  assign n8061 = ~n1737 & n8060 ;
  assign n8062 = n1093 & n2542 ;
  assign n8063 = ~n8061 & n8062 ;
  assign n8064 = n8063 ^ n2136 ^ 1'b0 ;
  assign n8065 = n380 & ~n2467 ;
  assign n8066 = n8065 ^ n4662 ^ 1'b0 ;
  assign n8067 = ~n2288 & n4508 ;
  assign n8068 = n6546 ^ n5231 ^ 1'b0 ;
  assign n8069 = n5784 ^ n30 ^ 1'b0 ;
  assign n8070 = n666 | n2080 ;
  assign n8072 = n703 & n799 ;
  assign n8071 = n987 & n1976 ;
  assign n8073 = n8072 ^ n8071 ^ 1'b0 ;
  assign n8074 = n3477 ^ n2825 ^ 1'b0 ;
  assign n8075 = ~n4784 & n8074 ;
  assign n8076 = n207 & ~n1620 ;
  assign n8077 = n8076 ^ n5418 ^ n1458 ;
  assign n8078 = n384 & ~n852 ;
  assign n8079 = ~n1220 & n8078 ;
  assign n8080 = n278 & n3354 ;
  assign n8081 = n8079 & ~n8080 ;
  assign n8082 = n5158 ^ n3091 ^ 1'b0 ;
  assign n8083 = n4884 ^ n2478 ^ 1'b0 ;
  assign n8084 = n2551 & ~n8083 ;
  assign n8085 = n458 | n4197 ;
  assign n8086 = n8085 ^ n782 ^ 1'b0 ;
  assign n8087 = n1359 ^ n66 ^ 1'b0 ;
  assign n8088 = n2229 & ~n8087 ;
  assign n8089 = ~n1560 & n8088 ;
  assign n8090 = n8089 ^ n1900 ^ 1'b0 ;
  assign n8091 = n1330 | n1549 ;
  assign n8092 = n5860 ^ n993 ^ 1'b0 ;
  assign n8093 = n713 | n1608 ;
  assign n8094 = n1984 & ~n8093 ;
  assign n8095 = n241 & n8094 ;
  assign n8096 = n1748 | n3293 ;
  assign n8097 = n8096 ^ n7524 ^ 1'b0 ;
  assign n8098 = n58 | n8097 ;
  assign n8099 = ~n4570 & n8098 ;
  assign n8100 = n7251 ^ n3254 ^ 1'b0 ;
  assign n8101 = n4327 & n8100 ;
  assign n8102 = n3221 ^ n1598 ^ 1'b0 ;
  assign n8103 = n8102 ^ n5856 ^ 1'b0 ;
  assign n8104 = n5894 & ~n8103 ;
  assign n8105 = n6194 | n6442 ;
  assign n8106 = n2347 & n4791 ;
  assign n8107 = n5534 ^ n1274 ^ 1'b0 ;
  assign n8108 = n1034 | n7628 ;
  assign n8109 = n1040 ^ n715 ^ 1'b0 ;
  assign n8110 = n2316 | n3561 ;
  assign n8111 = n4029 ^ n1891 ^ 1'b0 ;
  assign n8112 = n5932 | n8111 ;
  assign n8113 = n6628 & ~n8112 ;
  assign n8114 = ~n2799 & n8113 ;
  assign n8115 = n2569 ^ n2243 ^ 1'b0 ;
  assign n8116 = n4186 | n5322 ;
  assign n8117 = n8065 ^ n499 ^ 1'b0 ;
  assign n8118 = n8019 ^ n7657 ^ 1'b0 ;
  assign n8119 = n4722 & n8118 ;
  assign n8120 = n385 & n7936 ;
  assign n8121 = ~n5308 & n8120 ;
  assign n8122 = n8121 ^ n4155 ^ 1'b0 ;
  assign n8124 = ~n86 & n1130 ;
  assign n8125 = n1437 & n8124 ;
  assign n8123 = n3063 & n5021 ;
  assign n8126 = n8125 ^ n8123 ^ 1'b0 ;
  assign n8127 = n7438 | n8126 ;
  assign n8128 = n7597 ^ n6598 ^ 1'b0 ;
  assign n8129 = n3533 & n5517 ;
  assign n8130 = n941 ^ n382 ^ 1'b0 ;
  assign n8131 = n3061 & ~n8130 ;
  assign n8132 = n6388 & n8131 ;
  assign n8133 = n5401 | n8132 ;
  assign n8134 = ~n384 & n8133 ;
  assign n8135 = n6225 ^ n509 ^ 1'b0 ;
  assign n8136 = n7440 ^ n2235 ^ 1'b0 ;
  assign n8137 = n4322 | n8136 ;
  assign n8138 = n607 & ~n726 ;
  assign n8139 = n198 | n2055 ;
  assign n8140 = n8139 ^ n3787 ^ 1'b0 ;
  assign n8141 = n6818 ^ n4747 ^ 1'b0 ;
  assign n8142 = n8141 ^ n274 ^ 1'b0 ;
  assign n8143 = n6703 & ~n8142 ;
  assign n8144 = n517 & ~n4513 ;
  assign n8145 = n4549 ^ n2964 ^ 1'b0 ;
  assign n8146 = n3825 & ~n3849 ;
  assign n8147 = n8146 ^ n495 ^ 1'b0 ;
  assign n8148 = n8145 & ~n8147 ;
  assign n8149 = n251 & n2014 ;
  assign n8150 = n6079 & n8149 ;
  assign n8151 = ~n3567 & n8150 ;
  assign n8152 = n2086 & n4191 ;
  assign n8153 = n8152 ^ n310 ^ 1'b0 ;
  assign n8154 = n8153 ^ n5355 ^ 1'b0 ;
  assign n8155 = n272 & n8154 ;
  assign n8156 = ~n456 & n2294 ;
  assign n8157 = n5953 | n7110 ;
  assign n8158 = n3719 & ~n8157 ;
  assign n8159 = ~n5362 & n6394 ;
  assign n8160 = n8159 ^ n405 ^ 1'b0 ;
  assign n8161 = ~n3880 & n4639 ;
  assign n8162 = n4288 & ~n8161 ;
  assign n8163 = n769 | n1922 ;
  assign n8165 = n83 | n474 ;
  assign n8164 = n6426 | n7555 ;
  assign n8166 = n8165 ^ n8164 ^ 1'b0 ;
  assign n8167 = n4730 ^ n2519 ^ 1'b0 ;
  assign n8168 = n8167 ^ n5532 ^ 1'b0 ;
  assign n8169 = n6275 | n8168 ;
  assign n8170 = n2790 ^ n111 ^ 1'b0 ;
  assign n8171 = n8170 ^ n2916 ^ 1'b0 ;
  assign n8172 = n4812 ^ n3603 ^ 1'b0 ;
  assign n8173 = n3927 | n4990 ;
  assign n8174 = n630 & n2302 ;
  assign n8175 = ~n8173 & n8174 ;
  assign n8176 = n5310 ^ n1441 ^ 1'b0 ;
  assign n8177 = n5962 | n8176 ;
  assign n8178 = n8175 | n8177 ;
  assign n8179 = n7625 & ~n8178 ;
  assign n8180 = ~n310 & n1565 ;
  assign n8181 = n8180 ^ n1692 ^ 1'b0 ;
  assign n8182 = ~n2138 & n8181 ;
  assign n8183 = n148 & n8182 ;
  assign n8184 = n8183 ^ n4908 ^ 1'b0 ;
  assign n8185 = ~n5282 & n5301 ;
  assign n8186 = ~n782 & n3532 ;
  assign n8188 = n2086 ^ n1412 ^ 1'b0 ;
  assign n8187 = n1976 | n7520 ;
  assign n8189 = n8188 ^ n8187 ^ 1'b0 ;
  assign n8190 = n8189 ^ n5835 ^ 1'b0 ;
  assign n8191 = ~n246 & n8190 ;
  assign n8192 = n1241 & ~n3483 ;
  assign n8193 = n5169 | n5283 ;
  assign n8194 = n8193 ^ n278 ^ 1'b0 ;
  assign n8195 = n7895 & n8194 ;
  assign n8196 = n7264 ^ n688 ^ 1'b0 ;
  assign n8197 = ~n3764 & n8196 ;
  assign n8198 = ~n5189 & n8197 ;
  assign n8199 = n158 & n3803 ;
  assign n8200 = n414 & ~n3311 ;
  assign n8201 = n1164 & n8200 ;
  assign n8202 = n375 & n8201 ;
  assign n8203 = n3106 ^ n607 ^ 1'b0 ;
  assign n8204 = n1433 | n2027 ;
  assign n8205 = n8203 & ~n8204 ;
  assign n8206 = n1274 ^ n1080 ^ 1'b0 ;
  assign n8207 = n6196 ^ n2313 ^ 1'b0 ;
  assign n8208 = n177 | n3108 ;
  assign n8209 = n8208 ^ n615 ^ 1'b0 ;
  assign n8210 = n804 & n3626 ;
  assign n8211 = n8210 ^ n7655 ^ 1'b0 ;
  assign n8212 = ~n8209 & n8211 ;
  assign n8213 = ~n1058 & n6468 ;
  assign n8214 = n8213 ^ n5241 ^ 1'b0 ;
  assign n8215 = n4969 ^ n832 ^ 1'b0 ;
  assign n8216 = n8215 ^ n812 ^ 1'b0 ;
  assign n8217 = n3404 ^ n3226 ^ 1'b0 ;
  assign n8218 = n3139 & ~n6835 ;
  assign n8219 = n3154 & ~n5201 ;
  assign n8220 = ~n4361 & n6810 ;
  assign n8221 = n3670 ^ n678 ^ 1'b0 ;
  assign n8222 = n8221 ^ n23 ^ 1'b0 ;
  assign n8223 = ~n591 & n8222 ;
  assign n8224 = n5659 & ~n6876 ;
  assign n8225 = ~n7589 & n8158 ;
  assign n8226 = n5550 | n6689 ;
  assign n8227 = n8226 ^ n8185 ^ n300 ;
  assign n8228 = n7180 ^ n592 ^ 1'b0 ;
  assign n8229 = n3905 | n8228 ;
  assign n8230 = n3774 & ~n6197 ;
  assign n8231 = n7388 ^ n3156 ^ 1'b0 ;
  assign n8232 = n7264 ^ n7124 ^ n3801 ;
  assign n8238 = n6960 ^ n69 ^ 1'b0 ;
  assign n8233 = n4353 ^ n862 ^ 1'b0 ;
  assign n8234 = n987 & n1271 ;
  assign n8235 = ~n6510 & n8234 ;
  assign n8236 = n3642 & n8235 ;
  assign n8237 = n8233 | n8236 ;
  assign n8239 = n8238 ^ n8237 ^ 1'b0 ;
  assign n8240 = n6761 ^ n1782 ^ 1'b0 ;
  assign n8241 = ~n488 & n8240 ;
  assign n8242 = n8241 ^ n6492 ^ 1'b0 ;
  assign n8243 = ~n5675 & n7717 ;
  assign n8244 = ~n2611 & n8243 ;
  assign n8245 = n255 & n1870 ;
  assign n8246 = n5794 | n8245 ;
  assign n8247 = n8246 ^ n5836 ^ 1'b0 ;
  assign n8248 = n5408 & n7612 ;
  assign n8249 = n7763 ^ n3449 ^ 1'b0 ;
  assign n8250 = n200 & ~n2463 ;
  assign n8251 = n5096 & n8250 ;
  assign n8252 = n3012 | n8251 ;
  assign n8253 = n8252 ^ n3820 ^ 1'b0 ;
  assign n8254 = n1447 & n1662 ;
  assign n8255 = n5647 ^ n5336 ^ 1'b0 ;
  assign n8256 = n8254 & n8255 ;
  assign n8257 = ~n2012 & n2076 ;
  assign n8258 = ~n111 & n580 ;
  assign n8259 = n1891 & ~n8258 ;
  assign n8260 = n1194 & n8259 ;
  assign n8261 = ~n8257 & n8260 ;
  assign n8262 = n3532 ^ n3221 ^ 1'b0 ;
  assign n8263 = n1260 | n2576 ;
  assign n8264 = n8263 ^ n192 ^ 1'b0 ;
  assign n8265 = ( n158 & n1207 ) | ( n158 & ~n1944 ) | ( n1207 & ~n1944 ) ;
  assign n8266 = n8265 ^ n3579 ^ 1'b0 ;
  assign n8270 = ~n1471 & n2220 ;
  assign n8271 = n5666 & n8270 ;
  assign n8267 = n346 & ~n915 ;
  assign n8268 = n8267 ^ n592 ^ 1'b0 ;
  assign n8269 = n8268 ^ n6160 ^ n1141 ;
  assign n8272 = n8271 ^ n8269 ^ 1'b0 ;
  assign n8273 = n8272 ^ n2148 ^ 1'b0 ;
  assign n8274 = ~n5860 & n8273 ;
  assign n8275 = n785 & n4311 ;
  assign n8276 = n4081 ^ n3046 ^ n847 ;
  assign n8277 = ~n591 & n8276 ;
  assign n8278 = n197 & n8277 ;
  assign n8279 = n2799 | n7087 ;
  assign n8280 = ~n55 & n8279 ;
  assign n8281 = n8044 ^ n545 ^ 1'b0 ;
  assign n8282 = n3112 ^ n515 ^ 1'b0 ;
  assign n8283 = n989 & n1411 ;
  assign n8284 = n8283 ^ n2869 ^ 1'b0 ;
  assign n8285 = n6334 & n8284 ;
  assign n8286 = ~n130 & n788 ;
  assign n8287 = n8286 ^ n3522 ^ 1'b0 ;
  assign n8288 = n319 & n8287 ;
  assign n8289 = n1166 ^ n1069 ^ 1'b0 ;
  assign n8290 = n8289 ^ n1814 ^ 1'b0 ;
  assign n8291 = n3116 | n4088 ;
  assign n8292 = n8291 ^ n2558 ^ 1'b0 ;
  assign n8293 = n2302 ^ n307 ^ 1'b0 ;
  assign n8294 = n2964 & ~n8293 ;
  assign n8295 = n843 & ~n1575 ;
  assign n8296 = n8295 ^ n457 ^ 1'b0 ;
  assign n8297 = n5704 ^ n5187 ^ 1'b0 ;
  assign n8298 = n8296 & ~n8297 ;
  assign n8299 = ~n3033 & n4219 ;
  assign n8300 = n6476 ^ n903 ^ 1'b0 ;
  assign n8301 = n984 & ~n7119 ;
  assign n8302 = n8301 ^ n2549 ^ 1'b0 ;
  assign n8303 = n8300 & ~n8302 ;
  assign n8304 = n8303 ^ n719 ^ 1'b0 ;
  assign n8305 = n4327 & ~n7424 ;
  assign n8306 = n1739 | n4961 ;
  assign n8307 = n4594 ^ n252 ^ 1'b0 ;
  assign n8308 = n8306 & n8307 ;
  assign n8309 = n8308 ^ n7330 ^ 1'b0 ;
  assign n8310 = n8309 ^ n5067 ^ n2933 ;
  assign n8311 = ~n6277 & n8310 ;
  assign n8312 = n1963 & n2828 ;
  assign n8313 = ~n1130 & n4626 ;
  assign n8314 = ~n8312 & n8313 ;
  assign n8315 = ~n1759 & n4100 ;
  assign n8316 = n8315 ^ n153 ^ 1'b0 ;
  assign n8317 = n4320 ^ n3276 ^ 1'b0 ;
  assign n8318 = n8317 ^ n79 ^ 1'b0 ;
  assign n8319 = n220 & n1105 ;
  assign n8320 = n3567 & ~n8319 ;
  assign n8321 = n1344 ^ n227 ^ 1'b0 ;
  assign n8322 = ~n2799 & n8321 ;
  assign n8323 = n2665 ^ n869 ^ 1'b0 ;
  assign n8324 = n294 & ~n8217 ;
  assign n8325 = n475 | n4919 ;
  assign n8326 = n6677 ^ n2714 ^ 1'b0 ;
  assign n8327 = n8325 & n8326 ;
  assign n8328 = n3037 & ~n5232 ;
  assign n8329 = n8328 ^ n5525 ^ 1'b0 ;
  assign n8330 = n754 & ~n8329 ;
  assign n8331 = n2136 ^ n1506 ^ 1'b0 ;
  assign n8332 = n3890 ^ n1453 ^ 1'b0 ;
  assign n8333 = ~n8331 & n8332 ;
  assign n8334 = n856 & ~n2414 ;
  assign n8335 = ~n856 & n8334 ;
  assign n8336 = ~n246 & n8335 ;
  assign n8337 = ~n1304 & n8336 ;
  assign n8338 = n4860 & ~n8337 ;
  assign n8339 = ~n4860 & n8338 ;
  assign n8343 = ~n1348 & n6585 ;
  assign n8344 = ~n6585 & n8343 ;
  assign n8340 = n7573 ^ n2927 ^ 1'b0 ;
  assign n8341 = n234 | n8340 ;
  assign n8342 = n4197 | n8341 ;
  assign n8345 = n8344 ^ n8342 ^ 1'b0 ;
  assign n8346 = n8339 | n8345 ;
  assign n8347 = n4327 ^ n1263 ^ n599 ;
  assign n8348 = n1106 & ~n3787 ;
  assign n8349 = n7794 & n8348 ;
  assign n8350 = n7715 & ~n8349 ;
  assign n8351 = n698 ^ n385 ^ 1'b0 ;
  assign n8353 = n5123 & ~n7106 ;
  assign n8354 = n8353 ^ n4336 ^ 1'b0 ;
  assign n8352 = ~n2280 & n3833 ;
  assign n8355 = n8354 ^ n8352 ^ 1'b0 ;
  assign n8356 = n1880 | n6220 ;
  assign n8357 = n8356 ^ n6090 ^ 1'b0 ;
  assign n8358 = n3025 & ~n8357 ;
  assign n8359 = n387 & ~n792 ;
  assign n8360 = n8359 ^ n1441 ^ 1'b0 ;
  assign n8361 = n423 & ~n1509 ;
  assign n8362 = ~n8360 & n8361 ;
  assign n8363 = n1437 ^ n748 ^ 1'b0 ;
  assign n8364 = n4229 ^ n588 ^ 1'b0 ;
  assign n8365 = ~n8363 & n8364 ;
  assign n8366 = n793 | n8365 ;
  assign n8367 = ~n3743 & n8366 ;
  assign n8368 = n8367 ^ n7599 ^ 1'b0 ;
  assign n8369 = n5020 | n7668 ;
  assign n8370 = n1532 | n8369 ;
  assign n8371 = ~n4455 & n5131 ;
  assign n8372 = n255 & n8371 ;
  assign n8373 = n1273 & ~n2728 ;
  assign n8374 = n699 & n2017 ;
  assign n8375 = n8374 ^ n3228 ^ 1'b0 ;
  assign n8376 = n5162 & n8375 ;
  assign n8377 = n8376 ^ n726 ^ 1'b0 ;
  assign n8378 = n876 | n3497 ;
  assign n8379 = n8378 ^ n1054 ^ 1'b0 ;
  assign n8380 = n8379 ^ n2531 ^ 1'b0 ;
  assign n8381 = n8380 ^ n927 ^ 1'b0 ;
  assign n8382 = ~n5891 & n6468 ;
  assign n8383 = n8382 ^ n776 ^ 1'b0 ;
  assign n8384 = n5957 | n8383 ;
  assign n8385 = n1672 | n2235 ;
  assign n8386 = n3606 & ~n8385 ;
  assign n8387 = ~n348 & n8386 ;
  assign n8388 = n1745 ^ n608 ^ n216 ;
  assign n8389 = ~n3520 & n6655 ;
  assign n8390 = n5090 & ~n8389 ;
  assign n8391 = ~n570 & n8390 ;
  assign n8392 = n21 & ~n60 ;
  assign n8393 = n1937 & n8392 ;
  assign n8394 = n732 ^ n280 ^ 1'b0 ;
  assign n8395 = n8393 | n8394 ;
  assign n8396 = n5201 & n7383 ;
  assign n8397 = n3444 ^ n2826 ^ 1'b0 ;
  assign n8398 = n1254 & n7696 ;
  assign n8399 = n1886 & ~n8398 ;
  assign n8401 = ~n694 & n1203 ;
  assign n8400 = ~n3074 & n8310 ;
  assign n8402 = n8401 ^ n8400 ^ 1'b0 ;
  assign n8403 = n3158 & ~n6200 ;
  assign n8405 = n186 & n2696 ;
  assign n8404 = ~n1070 & n5946 ;
  assign n8406 = n8405 ^ n8404 ^ 1'b0 ;
  assign n8407 = n284 & ~n450 ;
  assign n8408 = n4114 ^ n3408 ^ 1'b0 ;
  assign n8409 = n361 & n8408 ;
  assign n8410 = n1293 & n8409 ;
  assign n8411 = n4217 ^ n2014 ^ 1'b0 ;
  assign n8412 = n1149 ^ n286 ^ 1'b0 ;
  assign n8413 = n1947 | n8412 ;
  assign n8414 = n8411 | n8413 ;
  assign n8415 = n5706 ^ n5255 ^ 1'b0 ;
  assign n8416 = ~n3037 & n4857 ;
  assign n8417 = n7192 ^ n2312 ^ 1'b0 ;
  assign n8418 = n6966 & ~n8417 ;
  assign n8419 = n246 | n8418 ;
  assign n8420 = n1458 ^ n364 ^ 1'b0 ;
  assign n8421 = n5076 & ~n8420 ;
  assign n8422 = n8269 ^ n6090 ^ 1'b0 ;
  assign n8423 = n6977 & n7751 ;
  assign n8424 = n167 & n8423 ;
  assign n8425 = ~n611 & n3167 ;
  assign n8426 = ~n7391 & n8425 ;
  assign n8427 = n3908 & ~n3965 ;
  assign n8428 = n8427 ^ n5060 ^ 1'b0 ;
  assign n8429 = n178 & ~n8428 ;
  assign n8430 = n3064 & n7279 ;
  assign n8431 = n2719 ^ n1979 ^ 1'b0 ;
  assign n8432 = n3804 | n8431 ;
  assign n8433 = n4797 & ~n6989 ;
  assign n8434 = n3925 | n4514 ;
  assign n8435 = n8434 ^ n4303 ^ 1'b0 ;
  assign n8436 = n8433 & n8435 ;
  assign n8437 = n1622 & n8436 ;
  assign n8438 = n784 & n6335 ;
  assign n8439 = n8438 ^ n6918 ^ 1'b0 ;
  assign n8440 = ~n164 & n8439 ;
  assign n8441 = n8440 ^ n3399 ^ 1'b0 ;
  assign n8442 = n3780 & n6782 ;
  assign n8443 = n8442 ^ n3154 ^ 1'b0 ;
  assign n8444 = n5309 & ~n8443 ;
  assign n8445 = n6161 | n8329 ;
  assign n8446 = ~n357 & n418 ;
  assign n8447 = n6079 & ~n7006 ;
  assign n8448 = n8446 & n8447 ;
  assign n8449 = n2841 & ~n4156 ;
  assign n8450 = n161 & n8449 ;
  assign n8451 = n865 | n8450 ;
  assign n8452 = n4965 ^ n899 ^ 1'b0 ;
  assign n8453 = n1611 & ~n3427 ;
  assign n8454 = ~n691 & n8453 ;
  assign n8455 = ~n3097 & n8454 ;
  assign n8456 = n3638 ^ n615 ^ 1'b0 ;
  assign n8457 = ~n8455 & n8456 ;
  assign n8458 = n1237 | n8342 ;
  assign n8459 = n1786 & n4180 ;
  assign n8460 = n55 & n553 ;
  assign n8461 = n8460 ^ n3759 ^ 1'b0 ;
  assign n8462 = n1831 & ~n8387 ;
  assign n8463 = n8462 ^ n53 ^ 1'b0 ;
  assign n8464 = ( n818 & n1833 ) | ( n818 & ~n7812 ) | ( n1833 & ~n7812 ) ;
  assign n8465 = n2997 ^ n90 ^ 1'b0 ;
  assign n8466 = n3334 & ~n8465 ;
  assign n8467 = n4924 & n8466 ;
  assign n8468 = n4437 | n7810 ;
  assign n8469 = n8468 ^ n8451 ^ 1'b0 ;
  assign n8470 = ~n1349 & n1966 ;
  assign n8471 = n2120 & ~n4212 ;
  assign n8472 = n8471 ^ n1519 ^ 1'b0 ;
  assign n8473 = n3743 | n3916 ;
  assign n8474 = ~n390 & n8473 ;
  assign n8475 = n3219 & n8474 ;
  assign n8476 = n5597 & ~n5957 ;
  assign n8477 = ~n1733 & n8476 ;
  assign n8478 = ~n5917 & n7123 ;
  assign n8479 = n6090 & n8478 ;
  assign n8480 = n6849 ^ n4774 ^ 1'b0 ;
  assign n8481 = ~n142 & n2388 ;
  assign n8482 = ~n2189 & n8481 ;
  assign n8484 = n4349 & n4639 ;
  assign n8485 = n8484 ^ n1385 ^ 1'b0 ;
  assign n8486 = n7516 & ~n8485 ;
  assign n8483 = n4645 | n7067 ;
  assign n8487 = n8486 ^ n8483 ^ 1'b0 ;
  assign n8488 = n4874 ^ n137 ^ 1'b0 ;
  assign n8489 = n8488 ^ n1177 ^ 1'b0 ;
  assign n8490 = n5090 & ~n6651 ;
  assign n8491 = n5812 ^ n1926 ^ 1'b0 ;
  assign n8492 = n1256 & n3089 ;
  assign n8493 = n7487 & n8492 ;
  assign n8494 = n3387 & n7221 ;
  assign n8495 = n724 ^ n51 ^ 1'b0 ;
  assign n8496 = ~n6633 & n8495 ;
  assign n8497 = n1794 & n8496 ;
  assign n8498 = n3144 & ~n8497 ;
  assign n8499 = n532 & n8498 ;
  assign n8500 = n380 & n3376 ;
  assign n8501 = n1499 | n8500 ;
  assign n8502 = n1937 | n8501 ;
  assign n8503 = n1710 | n8502 ;
  assign n8508 = n6573 ^ n4623 ^ 1'b0 ;
  assign n8504 = n907 ^ n261 ^ 1'b0 ;
  assign n8505 = n2553 ^ n1091 ^ 1'b0 ;
  assign n8506 = n8504 | n8505 ;
  assign n8507 = n8506 ^ n1740 ^ 1'b0 ;
  assign n8509 = n8508 ^ n8507 ^ 1'b0 ;
  assign n8510 = n6041 | n8509 ;
  assign n8511 = n787 & ~n3743 ;
  assign n8512 = n8511 ^ n1069 ^ 1'b0 ;
  assign n8513 = ~n200 & n2731 ;
  assign n8514 = n5897 & n8513 ;
  assign n8515 = n703 & n8183 ;
  assign n8516 = n744 | n8515 ;
  assign n8517 = n8514 | n8516 ;
  assign n8518 = n35 & ~n2813 ;
  assign n8519 = n8518 ^ n4404 ^ 1'b0 ;
  assign n8520 = ~n216 & n8519 ;
  assign n8521 = ~n4780 & n8520 ;
  assign n8522 = n387 & n1777 ;
  assign n8523 = n8522 ^ n259 ^ 1'b0 ;
  assign n8524 = ~n68 & n8523 ;
  assign n8525 = n1829 ^ n781 ^ 1'b0 ;
  assign n8526 = n6224 ^ n3075 ^ 1'b0 ;
  assign n8527 = n3447 ^ n2893 ^ 1'b0 ;
  assign n8528 = n5657 ^ x7 ^ 1'b0 ;
  assign n8529 = n8527 & ~n8528 ;
  assign n8530 = n2633 & ~n4169 ;
  assign n8531 = n1486 & n1954 ;
  assign n8532 = n7932 & n8531 ;
  assign n8533 = n8532 ^ n8459 ^ 1'b0 ;
  assign n8534 = n4024 & n8533 ;
  assign n8538 = n584 | n4225 ;
  assign n8539 = n274 & ~n8538 ;
  assign n8535 = ~n4429 & n7711 ;
  assign n8536 = n364 & n8535 ;
  assign n8537 = n4400 | n8536 ;
  assign n8540 = n8539 ^ n8537 ^ 1'b0 ;
  assign n8541 = n6655 ^ n5264 ^ 1'b0 ;
  assign n8542 = n384 & ~n2848 ;
  assign n8543 = n6392 & n8542 ;
  assign n8544 = n713 | n8112 ;
  assign n8545 = n8544 ^ n1476 ^ 1'b0 ;
  assign n8546 = ~n3640 & n8545 ;
  assign n8547 = n364 & ~n5251 ;
  assign n8548 = n8547 ^ n5844 ^ 1'b0 ;
  assign n8549 = n3806 ^ n1866 ^ 1'b0 ;
  assign n8550 = n7994 ^ n715 ^ 1'b0 ;
  assign n8551 = n2386 & n3926 ;
  assign n8552 = ~n930 & n1656 ;
  assign n8553 = ~n5652 & n8552 ;
  assign n8554 = n1441 | n5903 ;
  assign n8555 = n8554 ^ n2179 ^ 1'b0 ;
  assign n8556 = n3781 & ~n6577 ;
  assign n8557 = ~n2181 & n8556 ;
  assign n8558 = ( n322 & ~n458 ) | ( n322 & n2219 ) | ( ~n458 & n2219 ) ;
  assign n8559 = n8558 ^ n2333 ^ 1'b0 ;
  assign n8560 = n5278 ^ n4024 ^ 1'b0 ;
  assign n8561 = n8560 ^ n5929 ^ 1'b0 ;
  assign n8562 = n500 | n3025 ;
  assign n8563 = n2400 ^ n823 ^ 1'b0 ;
  assign n8564 = n8563 ^ n6306 ^ 1'b0 ;
  assign n8565 = n4812 ^ n2244 ^ 1'b0 ;
  assign n8566 = n6080 | n8565 ;
  assign n8567 = n4559 & ~n8566 ;
  assign n8568 = ~n342 & n495 ;
  assign n8569 = n330 & n8568 ;
  assign n8570 = n8569 ^ n919 ^ 1'b0 ;
  assign n8571 = ~n6072 & n8570 ;
  assign n8572 = n1827 | n5302 ;
  assign n8573 = n8572 ^ n2959 ^ 1'b0 ;
  assign n8574 = n2836 & n5892 ;
  assign n8575 = n4788 | n8574 ;
  assign n8576 = n491 & ~n785 ;
  assign n8577 = ~n1210 & n8576 ;
  assign n8578 = n4342 & ~n8577 ;
  assign n8579 = n7310 & n8578 ;
  assign n8580 = n1304 | n1329 ;
  assign n8581 = n753 & ~n8580 ;
  assign n8582 = ( ~n1001 & n8160 ) | ( ~n1001 & n8581 ) | ( n8160 & n8581 ) ;
  assign n8583 = n1025 & n2136 ;
  assign n8586 = n3408 ^ n444 ^ 1'b0 ;
  assign n8584 = n1447 & ~n3116 ;
  assign n8585 = n4560 | n8584 ;
  assign n8587 = n8586 ^ n8585 ^ 1'b0 ;
  assign n8588 = n1711 | n4116 ;
  assign n8589 = n8588 ^ n4840 ^ 1'b0 ;
  assign n8590 = n577 & ~n4298 ;
  assign n8591 = ~n748 & n8590 ;
  assign n8592 = ~n2176 & n8591 ;
  assign n8593 = n8592 ^ n890 ^ 1'b0 ;
  assign n8594 = n8589 & n8593 ;
  assign n8595 = n1184 & n2166 ;
  assign n8596 = n7388 ^ n4487 ^ 1'b0 ;
  assign n8597 = n4964 & ~n8574 ;
  assign n8598 = n8597 ^ n5793 ^ 1'b0 ;
  assign n8599 = n8598 ^ n1704 ^ 1'b0 ;
  assign n8600 = n1496 & ~n7384 ;
  assign n8601 = n622 & n8600 ;
  assign n8602 = n4257 ^ n2825 ^ 1'b0 ;
  assign n8603 = n1857 & ~n8602 ;
  assign n8604 = n8603 ^ n2130 ^ 1'b0 ;
  assign n8605 = n2572 & n8604 ;
  assign n8606 = ~n5863 & n6785 ;
  assign n8607 = ~n5412 & n8606 ;
  assign n8608 = n2353 & ~n8607 ;
  assign n8609 = n506 & n2636 ;
  assign n8610 = ~n654 & n8062 ;
  assign n8611 = n2426 & n8610 ;
  assign n8614 = n4411 ^ n244 ^ 1'b0 ;
  assign n8612 = n1463 & ~n2014 ;
  assign n8613 = n8612 ^ n4832 ^ 1'b0 ;
  assign n8615 = n8614 ^ n8613 ^ 1'b0 ;
  assign n8616 = n1040 & n8615 ;
  assign n8617 = ~n1814 & n6773 ;
  assign n8618 = n8617 ^ n663 ^ 1'b0 ;
  assign n8619 = ~n3749 & n8618 ;
  assign n8620 = n3744 ^ n284 ^ 1'b0 ;
  assign n8621 = n5251 ^ n3134 ^ 1'b0 ;
  assign n8622 = n5440 & n8621 ;
  assign n8623 = n8622 ^ n2472 ^ 1'b0 ;
  assign n8624 = n3792 ^ n2116 ^ 1'b0 ;
  assign n8625 = ( n727 & n779 ) | ( n727 & ~n1943 ) | ( n779 & ~n1943 ) ;
  assign n8626 = n5953 | n7124 ;
  assign n8627 = n6946 ^ n190 ^ 1'b0 ;
  assign n8628 = n8507 & ~n8574 ;
  assign n8629 = n2645 & ~n4463 ;
  assign n8630 = n7901 ^ n5342 ^ 1'b0 ;
  assign n8631 = n4516 & ~n8630 ;
  assign n8632 = ~n246 & n8631 ;
  assign n8633 = n1304 | n8632 ;
  assign n8634 = n7581 & ~n8633 ;
  assign n8635 = ~n1023 & n1692 ;
  assign n8636 = n8635 ^ n2335 ^ 1'b0 ;
  assign n8637 = x8 & n8636 ;
  assign n8638 = n8637 ^ n1487 ^ 1'b0 ;
  assign n8639 = n1331 & n8638 ;
  assign n8640 = n5134 & n8639 ;
  assign n8641 = n7570 & n8640 ;
  assign n8642 = n7095 | n8641 ;
  assign n8643 = n8634 & ~n8642 ;
  assign n8644 = n1388 & n8583 ;
  assign n8645 = ~n454 & n570 ;
  assign n8646 = ~n1941 & n8645 ;
  assign n8647 = n8646 ^ n1637 ^ 1'b0 ;
  assign n8648 = ~n1159 & n8647 ;
  assign n8649 = n1859 & ~n3976 ;
  assign n8650 = n8649 ^ n8574 ^ 1'b0 ;
  assign n8651 = n121 & ~n8650 ;
  assign n8652 = n8651 ^ n2721 ^ 1'b0 ;
  assign n8653 = n2939 ^ n1359 ^ 1'b0 ;
  assign n8654 = n1463 & ~n5123 ;
  assign n8655 = n8654 ^ n4079 ^ 1'b0 ;
  assign n8656 = n323 & n8655 ;
  assign n8657 = ~n5859 & n8163 ;
  assign n8658 = n2560 | n4169 ;
  assign n8659 = n8658 ^ n5020 ^ 1'b0 ;
  assign n8660 = ( n436 & n4677 ) | ( n436 & n5775 ) | ( n4677 & n5775 ) ;
  assign n8661 = n8660 ^ n273 ^ 1'b0 ;
  assign n8662 = n1975 & ~n8661 ;
  assign n8663 = ~n4924 & n8662 ;
  assign n8664 = n8663 ^ n4037 ^ 1'b0 ;
  assign n8665 = ~n7329 & n8392 ;
  assign n8666 = ~n2316 & n5702 ;
  assign n8667 = n8524 & ~n8666 ;
  assign n8668 = n6125 ^ n851 ^ 1'b0 ;
  assign n8669 = n2541 ^ n2386 ^ 1'b0 ;
  assign n8670 = n4315 | n8294 ;
  assign n8671 = n671 & n7617 ;
  assign n8672 = ~n2252 & n8671 ;
  assign n8673 = n1627 & ~n6236 ;
  assign n8674 = ~n5174 & n8673 ;
  assign n8675 = n1673 ^ n759 ^ 1'b0 ;
  assign n8676 = n2408 & n2652 ;
  assign n8677 = n8676 ^ n6220 ^ 1'b0 ;
  assign n8678 = n8677 ^ n2076 ^ 1'b0 ;
  assign n8679 = n3120 & n8678 ;
  assign n8680 = n8675 & ~n8679 ;
  assign n8681 = n5053 & ~n8680 ;
  assign n8682 = n19 | n1165 ;
  assign n8683 = n1033 | n8682 ;
  assign n8684 = n2813 & n8683 ;
  assign n8685 = n6079 | n6322 ;
  assign n8686 = n8685 ^ n4506 ^ 1'b0 ;
  assign n8687 = ~n4068 & n7734 ;
  assign n8688 = n1671 | n5811 ;
  assign n8689 = ~n148 & n8688 ;
  assign n8690 = n1295 ^ n594 ^ 1'b0 ;
  assign n8691 = ~n3447 & n3535 ;
  assign n8692 = n8690 & n8691 ;
  assign n8700 = n210 | n4979 ;
  assign n8701 = n5537 | n8700 ;
  assign n8693 = n19 | n271 ;
  assign n8694 = n7391 ^ n2883 ^ 1'b0 ;
  assign n8695 = n434 | n2973 ;
  assign n8696 = n428 & ~n8695 ;
  assign n8697 = n8694 & n8696 ;
  assign n8698 = ~n8693 & n8697 ;
  assign n8699 = n4370 & n8698 ;
  assign n8702 = n8701 ^ n8699 ^ 1'b0 ;
  assign n8703 = n8692 | n8702 ;
  assign n8704 = n5691 ^ n4642 ^ 1'b0 ;
  assign n8705 = n983 ^ n483 ^ 1'b0 ;
  assign n8706 = n86 | n1428 ;
  assign n8707 = n8705 & n8706 ;
  assign n8708 = n3734 & n4215 ;
  assign n8709 = n194 & n323 ;
  assign n8710 = n8709 ^ n6162 ^ 1'b0 ;
  assign n8711 = n6439 ^ n1169 ^ 1'b0 ;
  assign n8712 = n287 & n2984 ;
  assign n8713 = n8712 ^ n5193 ^ 1'b0 ;
  assign n8714 = n2881 & n8713 ;
  assign n8715 = n8714 ^ n5920 ^ 1'b0 ;
  assign n8716 = n8715 ^ n8221 ^ 1'b0 ;
  assign n8717 = ~n5454 & n8716 ;
  assign n8718 = n1227 & ~n7193 ;
  assign n8719 = n3089 ^ n2738 ^ 1'b0 ;
  assign n8720 = n450 | n847 ;
  assign n8721 = n6275 & n8720 ;
  assign n8722 = n5716 & n8721 ;
  assign n8723 = ~n4961 & n8722 ;
  assign n8724 = n6248 ^ n1479 ^ 1'b0 ;
  assign n8725 = n6295 & n8724 ;
  assign n8726 = n610 & n8725 ;
  assign n8727 = n3758 ^ n3221 ^ 1'b0 ;
  assign n8728 = n4332 & ~n8727 ;
  assign n8729 = n5986 ^ n3180 ^ 1'b0 ;
  assign n8730 = n472 & n2261 ;
  assign n8731 = n6979 | n8730 ;
  assign n8732 = n5217 & ~n8731 ;
  assign n8733 = ~n602 & n7011 ;
  assign n8734 = ~n6503 & n8733 ;
  assign n8735 = n4830 ^ n185 ^ 1'b0 ;
  assign n8736 = ~n1437 & n8735 ;
  assign n8737 = ~n119 & n4729 ;
  assign n8738 = n8736 & ~n8737 ;
  assign n8739 = n8738 ^ n133 ^ 1'b0 ;
  assign n8744 = n149 & n3638 ;
  assign n8740 = n4125 | n7120 ;
  assign n8741 = ~n876 & n1358 ;
  assign n8742 = n8741 ^ n5024 ^ 1'b0 ;
  assign n8743 = n8740 & n8742 ;
  assign n8745 = n8744 ^ n8743 ^ 1'b0 ;
  assign n8746 = ~n2410 & n4086 ;
  assign n8747 = n5225 & n8746 ;
  assign n8748 = ~n1323 & n6866 ;
  assign n8749 = ~n3398 & n8748 ;
  assign n8750 = n1516 & ~n8749 ;
  assign n8751 = n8750 ^ n4626 ^ 1'b0 ;
  assign n8752 = n557 & ~n5158 ;
  assign n8753 = n8752 ^ n89 ^ 1'b0 ;
  assign n8754 = n3512 & ~n7289 ;
  assign n8755 = ~n2627 & n8754 ;
  assign n8756 = n8753 | n8755 ;
  assign n8757 = n1473 & ~n7310 ;
  assign n8758 = n3338 | n8203 ;
  assign n8759 = n3577 & ~n8758 ;
  assign n8760 = n8759 ^ n1539 ^ 1'b0 ;
  assign n8761 = n417 & ~n694 ;
  assign n8762 = n1038 | n8761 ;
  assign n8763 = n1469 & ~n3354 ;
  assign n8764 = n8762 & n8763 ;
  assign n8765 = n6543 ^ n221 ^ 1'b0 ;
  assign n8766 = n3938 ^ n1628 ^ 1'b0 ;
  assign n8767 = n5455 | n8766 ;
  assign n8768 = n6009 | n8767 ;
  assign n8769 = n7373 ^ n865 ^ 1'b0 ;
  assign n8771 = n4231 & n7810 ;
  assign n8770 = n2546 & n8229 ;
  assign n8772 = n8771 ^ n8770 ^ 1'b0 ;
  assign n8773 = ~n8769 & n8772 ;
  assign n8774 = n8613 ^ n4529 ^ 1'b0 ;
  assign n8775 = ~n880 & n8774 ;
  assign n8776 = n102 & n2191 ;
  assign n8777 = ~n187 & n8776 ;
  assign n8778 = n5702 ^ n5394 ^ 1'b0 ;
  assign n8779 = ~n8777 & n8778 ;
  assign n8780 = n2236 ^ n1443 ^ 1'b0 ;
  assign n8781 = n2912 ^ n1310 ^ 1'b0 ;
  assign n8782 = n507 & n8781 ;
  assign n8783 = n94 & ~n8782 ;
  assign n8784 = n2076 ^ n1764 ^ 1'b0 ;
  assign n8785 = n7686 & ~n8784 ;
  assign n8786 = n1394 & n3298 ;
  assign n8787 = ~n903 & n8786 ;
  assign n8788 = n1418 ^ n1202 ^ 1'b0 ;
  assign n8789 = n86 & ~n1608 ;
  assign n8790 = ~n8788 & n8789 ;
  assign n8791 = n5063 & n8790 ;
  assign n8792 = n8787 & n8791 ;
  assign n8793 = n4236 & n4890 ;
  assign n8794 = n1999 ^ n385 ^ 1'b0 ;
  assign n8795 = n823 & ~n8794 ;
  assign n8796 = n4891 ^ n2477 ^ 1'b0 ;
  assign n8797 = n8795 & n8796 ;
  assign n8798 = n588 | n6100 ;
  assign n8799 = n580 & ~n2348 ;
  assign n8800 = ~n5544 & n8799 ;
  assign n8801 = n7507 ^ n251 ^ 1'b0 ;
  assign n8802 = ~n8800 & n8801 ;
  assign n8803 = n1529 & ~n3166 ;
  assign n8804 = n8296 ^ n2804 ^ 1'b0 ;
  assign n8805 = n3278 & n5617 ;
  assign n8806 = n8805 ^ n5385 ^ 1'b0 ;
  assign n8807 = n1034 | n1501 ;
  assign n8808 = n8807 ^ n273 ^ 1'b0 ;
  assign n8809 = n962 ^ n781 ^ 1'b0 ;
  assign n8810 = n8808 | n8809 ;
  assign n8811 = n8806 | n8810 ;
  assign n8812 = ~n1924 & n2283 ;
  assign n8813 = n1792 ^ n1728 ^ 1'b0 ;
  assign n8814 = n1329 | n4694 ;
  assign n8818 = n1117 | n1389 ;
  assign n8815 = n928 ^ n58 ^ 1'b0 ;
  assign n8816 = n8815 ^ n4756 ^ 1'b0 ;
  assign n8817 = ~n1505 & n8816 ;
  assign n8819 = n8818 ^ n8817 ^ 1'b0 ;
  assign n8820 = ~n1961 & n2087 ;
  assign n8821 = n2370 & ~n5673 ;
  assign n8822 = n4959 & n8821 ;
  assign n8823 = n8822 ^ n4609 ^ 1'b0 ;
  assign n8824 = ~n5201 & n5823 ;
  assign n8825 = n896 ^ n51 ^ 1'b0 ;
  assign n8826 = n2883 | n8825 ;
  assign n8827 = n931 & ~n1922 ;
  assign n8828 = ~n2496 & n8827 ;
  assign n8829 = n5152 & n8828 ;
  assign n8830 = n2873 ^ n158 ^ 1'b0 ;
  assign n8831 = n3477 ^ n2917 ^ 1'b0 ;
  assign n8832 = ~n8830 & n8831 ;
  assign n8833 = n6445 ^ n2432 ^ 1'b0 ;
  assign n8834 = n8833 ^ n5749 ^ n4976 ;
  assign n8835 = n8834 ^ n1165 ^ 1'b0 ;
  assign n8836 = n354 & ~n8835 ;
  assign n8837 = n4406 & n8836 ;
  assign n8838 = n8837 ^ n6254 ^ 1'b0 ;
  assign n8839 = n1314 ^ n493 ^ 1'b0 ;
  assign n8840 = ~n87 & n8839 ;
  assign n8841 = n37 | n8840 ;
  assign n8842 = n261 & n791 ;
  assign n8843 = n6417 | n8842 ;
  assign n8844 = n7972 ^ n1445 ^ 1'b0 ;
  assign n8845 = ~n1337 & n8844 ;
  assign n8846 = n6773 & n7808 ;
  assign n8847 = n46 | n8644 ;
  assign n8848 = n7030 ^ n6089 ^ 1'b0 ;
  assign n8849 = n3861 & ~n6709 ;
  assign n8850 = n8849 ^ n4081 ^ 1'b0 ;
  assign n8851 = n1051 & ~n8850 ;
  assign n8852 = n4264 & ~n4970 ;
  assign n8853 = ~n1431 & n8852 ;
  assign n8854 = n6232 & n7507 ;
  assign n8855 = n7553 | n7690 ;
  assign n8856 = n157 & ~n1193 ;
  assign n8857 = n158 & n8856 ;
  assign n8858 = n6900 ^ n4653 ^ 1'b0 ;
  assign n8859 = n101 & n4040 ;
  assign n8860 = n8859 ^ n4536 ^ 1'b0 ;
  assign n8861 = n690 | n8860 ;
  assign n8862 = n16 | n8861 ;
  assign n8863 = n6827 ^ n1815 ^ 1'b0 ;
  assign n8864 = n174 | n880 ;
  assign n8865 = n6305 | n8864 ;
  assign n8866 = ( n1495 & ~n3624 ) | ( n1495 & n8865 ) | ( ~n3624 & n8865 ) ;
  assign n8867 = n8071 & ~n8250 ;
  assign n8868 = n6485 & n8867 ;
  assign n8869 = ~n3037 & n8868 ;
  assign n8870 = n2817 ^ n384 ^ 1'b0 ;
  assign n8871 = n1879 & n5747 ;
  assign n8872 = n8871 ^ n1346 ^ 1'b0 ;
  assign n8873 = n2795 ^ n1426 ^ 1'b0 ;
  assign n8874 = n324 & ~n8873 ;
  assign n8875 = n339 | n1202 ;
  assign n8876 = n8875 ^ n6458 ^ 1'b0 ;
  assign n8877 = ~n8874 & n8876 ;
  assign n8878 = n257 & n5024 ;
  assign n8879 = n8878 ^ n6286 ^ 1'b0 ;
  assign n8880 = n7254 ^ n914 ^ 1'b0 ;
  assign n8881 = n4445 & n8880 ;
  assign n8882 = ~n1264 & n8881 ;
  assign n8883 = n1058 & n8882 ;
  assign n8884 = n628 & ~n4845 ;
  assign n8885 = ~n2263 & n3068 ;
  assign n8886 = n958 | n2770 ;
  assign n8887 = n8853 & ~n8886 ;
  assign n8888 = ( n4599 & n4613 ) | ( n4599 & ~n5250 ) | ( n4613 & ~n5250 ) ;
  assign n8889 = n8888 ^ n3985 ^ 1'b0 ;
  assign n8890 = n2200 & n3953 ;
  assign n8891 = ~n2817 & n8890 ;
  assign n8892 = n3156 ^ n2689 ^ 1'b0 ;
  assign n8893 = ( n8102 & n8891 ) | ( n8102 & n8892 ) | ( n8891 & n8892 ) ;
  assign n8894 = n356 & ~n687 ;
  assign n8895 = n3473 ^ n309 ^ 1'b0 ;
  assign n8896 = ~n8894 & n8895 ;
  assign n8897 = n1213 | n1987 ;
  assign n8898 = n4851 | n6481 ;
  assign n8899 = n2092 & n3916 ;
  assign n8900 = ~n5179 & n8899 ;
  assign n8901 = n1008 ^ n42 ^ 1'b0 ;
  assign n8902 = n6085 & ~n8901 ;
  assign n8903 = ~n24 & n2136 ;
  assign n8904 = n8903 ^ n5032 ^ n114 ;
  assign n8905 = n2163 | n5982 ;
  assign n8906 = n3158 ^ n310 ^ 1'b0 ;
  assign n8907 = n8210 & ~n8906 ;
  assign n8908 = n8907 ^ n6771 ^ 1'b0 ;
  assign n8909 = n1186 & n4991 ;
  assign n8910 = n8909 ^ n7935 ^ 1'b0 ;
  assign n8911 = n1161 & n6377 ;
  assign n8912 = ~n7511 & n8911 ;
  assign n8913 = n3512 ^ n106 ^ 1'b0 ;
  assign n8914 = n5245 & ~n8913 ;
  assign n8915 = n8912 | n8914 ;
  assign n8916 = n8283 ^ n6966 ^ 1'b0 ;
  assign n8917 = ~n1908 & n8916 ;
  assign n8918 = n690 | n5040 ;
  assign n8919 = n8917 & n8918 ;
  assign n8920 = n2404 & n2513 ;
  assign n8921 = ~n5295 & n8920 ;
  assign n8922 = n5002 ^ n1907 ^ 1'b0 ;
  assign n8923 = n8922 ^ n4253 ^ 1'b0 ;
  assign n8924 = ~n4543 & n5613 ;
  assign n8925 = n8924 ^ n816 ^ 1'b0 ;
  assign n8926 = n3361 ^ n993 ^ 1'b0 ;
  assign n8927 = n2025 & n8926 ;
  assign n8928 = n7868 & ~n8927 ;
  assign n8929 = n938 & n4220 ;
  assign n8930 = n8929 ^ n726 ^ 1'b0 ;
  assign n8931 = n315 & ~n8930 ;
  assign n8932 = n2937 & n8931 ;
  assign n8933 = n4116 ^ n2431 ^ 1'b0 ;
  assign n8934 = n3890 & n6411 ;
  assign n8935 = n8934 ^ n2342 ^ 1'b0 ;
  assign n8936 = n1329 & ~n2305 ;
  assign n8937 = n8936 ^ n759 ^ 1'b0 ;
  assign n8938 = n1638 ^ n1127 ^ n587 ;
  assign n8939 = n573 & n8938 ;
  assign n8940 = n8939 ^ n3797 ^ 1'b0 ;
  assign n8941 = ~n8937 & n8940 ;
  assign n8942 = n4406 ^ n1271 ^ 1'b0 ;
  assign n8943 = n1484 ^ n832 ^ 1'b0 ;
  assign n8944 = n4311 & ~n8943 ;
  assign n8945 = n954 | n5155 ;
  assign n8946 = n387 | n669 ;
  assign n8947 = n283 | n5962 ;
  assign n8948 = n4105 & ~n5889 ;
  assign n8950 = ~n1497 & n4519 ;
  assign n8949 = n175 | n677 ;
  assign n8951 = n8950 ^ n8949 ^ 1'b0 ;
  assign n8953 = n5355 ^ n3663 ^ 1'b0 ;
  assign n8954 = n8953 ^ n1851 ^ n1001 ;
  assign n8955 = n8954 ^ n799 ^ 1'b0 ;
  assign n8956 = n3361 & ~n8955 ;
  assign n8952 = n1659 | n8368 ;
  assign n8957 = n8956 ^ n8952 ^ 1'b0 ;
  assign n8958 = ~n5914 & n7664 ;
  assign n8959 = n8958 ^ n8409 ^ 1'b0 ;
  assign n8960 = ~n2180 & n6966 ;
  assign n8961 = ~n815 & n8960 ;
  assign n8962 = n757 | n8961 ;
  assign n8963 = n8962 ^ n1310 ^ 1'b0 ;
  assign n8964 = ~n7247 & n8963 ;
  assign n8965 = n8964 ^ n2587 ^ 1'b0 ;
  assign n8966 = n1072 & ~n3278 ;
  assign n8967 = n1310 | n8646 ;
  assign n8968 = ~n2665 & n7120 ;
  assign n8969 = ~n8967 & n8968 ;
  assign n8970 = n2490 & ~n8969 ;
  assign n8971 = n161 & n8970 ;
  assign n8972 = ~n1484 & n5210 ;
  assign n8973 = n817 | n1038 ;
  assign n8974 = n2749 ^ n509 ^ 1'b0 ;
  assign n8975 = n3846 & n8974 ;
  assign n8976 = n700 & n8975 ;
  assign n8977 = n2233 & n6331 ;
  assign n8978 = n258 & ~n1270 ;
  assign n8979 = ~n3718 & n8978 ;
  assign n8980 = n2714 & n8979 ;
  assign n8981 = ~n1233 & n6236 ;
  assign n8982 = ~n599 & n8981 ;
  assign n8983 = n38 & n5806 ;
  assign n8984 = n2472 & n8983 ;
  assign n8985 = n4251 & ~n8984 ;
  assign n8986 = ~n8982 & n8985 ;
  assign n8987 = ~n817 & n7713 ;
  assign n8988 = n294 & n618 ;
  assign n8989 = n4081 & n4186 ;
  assign n8990 = n4463 ^ n954 ^ 1'b0 ;
  assign n8991 = n2068 & n3061 ;
  assign n8992 = n8540 ^ n5979 ^ 1'b0 ;
  assign n8993 = n796 & ~n7996 ;
  assign n8994 = n4474 ^ n323 ^ 1'b0 ;
  assign n8995 = n8994 ^ n4378 ^ 1'b0 ;
  assign n8996 = n788 & ~n8552 ;
  assign n8997 = n8996 ^ n2397 ^ 1'b0 ;
  assign n8998 = n3779 & ~n8997 ;
  assign n8999 = ~n2495 & n5706 ;
  assign n9000 = n5148 ^ n4929 ^ 1'b0 ;
  assign n9001 = ~n2811 & n8840 ;
  assign n9002 = n1600 ^ n415 ^ 1'b0 ;
  assign n9003 = n7254 ^ n191 ^ 1'b0 ;
  assign n9004 = n9002 | n9003 ;
  assign n9005 = n4098 | n9004 ;
  assign n9006 = n1372 | n9005 ;
  assign n9007 = ~n9001 & n9006 ;
  assign n9008 = n7935 & n9007 ;
  assign n9009 = ~n1826 & n6127 ;
  assign n9010 = n525 | n1771 ;
  assign n9011 = n1227 | n1714 ;
  assign n9012 = n6897 ^ n5234 ^ 1'b0 ;
  assign n9013 = n2967 ^ n1138 ^ 1'b0 ;
  assign n9014 = n622 | n9013 ;
  assign n9015 = n9014 ^ n1426 ^ 1'b0 ;
  assign n9016 = n229 & n1629 ;
  assign n9017 = n8916 & n9016 ;
  assign n9018 = n1584 & n8823 ;
  assign n9019 = x5 & ~n2730 ;
  assign n9020 = n2043 & n2717 ;
  assign n9021 = n4039 ^ n3049 ^ 1'b0 ;
  assign n9022 = n4629 & n9021 ;
  assign n9023 = ~n2145 & n4952 ;
  assign n9024 = n9022 & ~n9023 ;
  assign n9025 = n666 & ~n7259 ;
  assign n9026 = ~n5639 & n9025 ;
  assign n9027 = n4677 ^ n522 ^ 1'b0 ;
  assign n9028 = ~n853 & n2927 ;
  assign n9029 = n9027 & n9028 ;
  assign n9030 = ~n7910 & n9029 ;
  assign n9031 = n62 | n1410 ;
  assign n9032 = n9031 ^ n1653 ^ 1'b0 ;
  assign n9033 = n1532 & n3290 ;
  assign n9034 = n738 & n9033 ;
  assign n9035 = n9034 ^ n2725 ^ 1'b0 ;
  assign n9036 = n9032 & ~n9035 ;
  assign n9037 = n817 | n1742 ;
  assign n9038 = n5819 & ~n9037 ;
  assign n9039 = n8861 ^ n2924 ^ 1'b0 ;
  assign n9040 = n3348 & ~n4111 ;
  assign n9041 = n9040 ^ n6333 ^ 1'b0 ;
  assign n9042 = n2695 ^ n178 ^ 1'b0 ;
  assign n9043 = ~n141 & n9042 ;
  assign n9044 = n8418 ^ n6167 ^ 1'b0 ;
  assign n9045 = n5849 & ~n9044 ;
  assign n9046 = n3177 & ~n7918 ;
  assign n9047 = n2453 & n6210 ;
  assign n9048 = ~n3786 & n4322 ;
  assign n9049 = n1505 ^ n681 ^ 1'b0 ;
  assign n9050 = n6932 & ~n9049 ;
  assign n9051 = n3081 & n9050 ;
  assign n9052 = n1737 & n4368 ;
  assign n9053 = n1785 ^ x0 ^ 1'b0 ;
  assign n9054 = n9053 ^ n445 ^ 1'b0 ;
  assign n9055 = n5806 & ~n9054 ;
  assign n9056 = n4499 ^ n685 ^ 1'b0 ;
  assign n9057 = n9056 ^ n2773 ^ 1'b0 ;
  assign n9058 = n5453 & n9057 ;
  assign n9059 = ~n3885 & n9058 ;
  assign n9060 = ( n6531 & ~n8843 ) | ( n6531 & n9059 ) | ( ~n8843 & n9059 ) ;
  assign n9061 = n4294 & n8069 ;
  assign n9062 = n3434 ^ n520 ^ 1'b0 ;
  assign n9063 = n7221 ^ n170 ^ 1'b0 ;
  assign n9064 = n1961 & ~n9063 ;
  assign n9065 = n6163 ^ n1106 ^ 1'b0 ;
  assign n9066 = n9065 ^ n226 ^ 1'b0 ;
  assign n9067 = n970 & ~n1329 ;
  assign n9068 = n1931 | n2626 ;
  assign n9069 = n632 | n9068 ;
  assign n9070 = n9069 ^ n6398 ^ 1'b0 ;
  assign n9071 = n89 & n1763 ;
  assign n9072 = n7589 & n9071 ;
  assign n9073 = ~n2268 & n3635 ;
  assign n9074 = n3873 & n9073 ;
  assign n9075 = ( n205 & n2577 ) | ( n205 & ~n9074 ) | ( n2577 & ~n9074 ) ;
  assign n9076 = n9072 | n9075 ;
  assign n9077 = n9076 ^ n945 ^ 1'b0 ;
  assign n9080 = ~n1219 & n2834 ;
  assign n9081 = n9080 ^ n8385 ^ n2059 ;
  assign n9078 = n1714 ^ n252 ^ 1'b0 ;
  assign n9079 = n4728 & ~n9078 ;
  assign n9082 = n9081 ^ n9079 ^ 1'b0 ;
  assign n9083 = n6715 ^ n1707 ^ n1225 ;
  assign n9084 = n376 & n8075 ;
  assign n9085 = n763 & n5254 ;
  assign n9086 = n3866 & ~n7098 ;
  assign n9088 = n1165 | n4942 ;
  assign n9089 = n7483 | n9088 ;
  assign n9090 = n3370 & ~n9089 ;
  assign n9091 = n9090 ^ n1878 ^ 1'b0 ;
  assign n9087 = n1950 & ~n5681 ;
  assign n9092 = n9091 ^ n9087 ^ 1'b0 ;
  assign n9093 = n216 & n787 ;
  assign n9094 = n9093 ^ n5528 ^ 1'b0 ;
  assign n9096 = n7767 ^ n539 ^ 1'b0 ;
  assign n9095 = n908 & ~n7310 ;
  assign n9097 = n9096 ^ n9095 ^ 1'b0 ;
  assign n9098 = n2199 & n9097 ;
  assign n9099 = ~n9094 & n9098 ;
  assign n9101 = n6329 ^ n5085 ^ 1'b0 ;
  assign n9102 = n2170 & ~n9101 ;
  assign n9100 = n8057 ^ n1884 ^ 1'b0 ;
  assign n9103 = n9102 ^ n9100 ^ 1'b0 ;
  assign n9104 = n6170 ^ n1008 ^ 1'b0 ;
  assign n9105 = n4204 ^ n3374 ^ 1'b0 ;
  assign n9106 = n599 | n7866 ;
  assign n9107 = n9106 ^ n233 ^ 1'b0 ;
  assign n9108 = ~n2202 & n3941 ;
  assign n9109 = n1178 & n1845 ;
  assign n9110 = n1133 | n5002 ;
  assign n9111 = n1270 & ~n9110 ;
  assign n9112 = n5760 ^ n5396 ^ 1'b0 ;
  assign n9113 = n9112 ^ n2060 ^ 1'b0 ;
  assign n9114 = n9111 | n9113 ;
  assign n9115 = n342 & ~n9114 ;
  assign n9116 = n9115 ^ n5002 ^ 1'b0 ;
  assign n9117 = ~n6412 & n9116 ;
  assign n9118 = n6062 & n8787 ;
  assign n9119 = n6666 | n9118 ;
  assign n9120 = n1956 ^ n694 ^ 1'b0 ;
  assign n9121 = n9120 ^ n8122 ^ 1'b0 ;
  assign n9122 = n460 | n4650 ;
  assign n9123 = n1783 & ~n9122 ;
  assign n9124 = n9123 ^ n4256 ^ 1'b0 ;
  assign n9125 = n1529 & n3417 ;
  assign n9126 = n9125 ^ n167 ^ 1'b0 ;
  assign n9127 = n1148 | n3015 ;
  assign n9128 = n9127 ^ n1865 ^ 1'b0 ;
  assign n9129 = n4328 ^ n2322 ^ 1'b0 ;
  assign n9130 = n9129 ^ n7353 ^ 1'b0 ;
  assign n9131 = n2155 ^ n977 ^ n390 ;
  assign n9132 = n9131 ^ n2209 ^ 1'b0 ;
  assign n9133 = n1447 & ~n5056 ;
  assign n9134 = n5156 & n9133 ;
  assign n9135 = n4809 | n7661 ;
  assign n9136 = n5980 ^ n484 ^ 1'b0 ;
  assign n9137 = n47 & ~n1276 ;
  assign n9138 = ~n2835 & n9137 ;
  assign n9139 = n9138 ^ n489 ^ 1'b0 ;
  assign n9140 = n9139 ^ n7346 ^ n1748 ;
  assign n9141 = n3377 & ~n3919 ;
  assign n9148 = n3443 & ~n3669 ;
  assign n9142 = n1566 & n3068 ;
  assign n9143 = n2861 & ~n9142 ;
  assign n9144 = n9143 ^ n1191 ^ 1'b0 ;
  assign n9145 = n3526 | n9144 ;
  assign n9146 = n533 & n8575 ;
  assign n9147 = ~n9145 & n9146 ;
  assign n9149 = n9148 ^ n9147 ^ 1'b0 ;
  assign n9150 = n2992 ^ n1097 ^ 1'b0 ;
  assign n9151 = n2615 & n9150 ;
  assign n9152 = n2377 | n6430 ;
  assign n9153 = n7048 & n9152 ;
  assign n9154 = n5355 ^ n750 ^ 1'b0 ;
  assign n9155 = n9154 ^ n741 ^ 1'b0 ;
  assign n9156 = n4575 ^ n4176 ^ 1'b0 ;
  assign n9157 = n4798 & ~n9156 ;
  assign n9158 = n395 | n4889 ;
  assign n9159 = n5160 & ~n9158 ;
  assign n9160 = ~n3843 & n4615 ;
  assign n9161 = n302 & n9160 ;
  assign n9162 = n1533 | n8210 ;
  assign n9163 = n9162 ^ n7034 ^ 1'b0 ;
  assign n9164 = n9163 ^ n5607 ^ n3089 ;
  assign n9165 = n6596 ^ n1088 ^ 1'b0 ;
  assign n9166 = n315 & ~n9165 ;
  assign n9167 = n27 | n977 ;
  assign n9168 = n2865 & ~n9167 ;
  assign n9169 = ~n9166 & n9168 ;
  assign n9170 = n157 & ~n2652 ;
  assign n9171 = n5223 & n7178 ;
  assign n9172 = n1868 & n8239 ;
  assign n9173 = n2799 ^ n489 ^ 1'b0 ;
  assign n9174 = n2245 & ~n9173 ;
  assign n9175 = n113 & ~n6944 ;
  assign n9176 = ~n581 & n9175 ;
  assign n9177 = n6846 ^ n2339 ^ 1'b0 ;
  assign n9178 = n5085 ^ n4812 ^ 1'b0 ;
  assign n9179 = ~n384 & n9178 ;
  assign n9180 = n9179 ^ n205 ^ 1'b0 ;
  assign n9181 = n1146 & ~n2816 ;
  assign n9182 = n7632 & n9181 ;
  assign n9183 = x6 & n367 ;
  assign n9184 = n227 & n9183 ;
  assign n9185 = n9184 ^ n1725 ^ 1'b0 ;
  assign n9186 = n79 & n9185 ;
  assign n9187 = ~n58 & n3144 ;
  assign n9188 = n9187 ^ n8242 ^ n2440 ;
  assign n9189 = ~n3634 & n3960 ;
  assign n9190 = n9189 ^ n2369 ^ 1'b0 ;
  assign n9191 = ~n1766 & n9190 ;
  assign n9192 = n1496 | n3480 ;
  assign n9193 = n5826 ^ n1038 ^ 1'b0 ;
  assign n9194 = n5336 ^ n266 ^ 1'b0 ;
  assign n9196 = n7930 ^ n5223 ^ 1'b0 ;
  assign n9197 = ~n1232 & n9196 ;
  assign n9195 = n5221 ^ n2131 ^ 1'b0 ;
  assign n9198 = n9197 ^ n9195 ^ 1'b0 ;
  assign n9199 = n4119 ^ n2665 ^ 1'b0 ;
  assign n9201 = ( n1103 & n1810 ) | ( n1103 & n4805 ) | ( n1810 & n4805 ) ;
  assign n9200 = n1571 & ~n1705 ;
  assign n9202 = n9201 ^ n9200 ^ 1'b0 ;
  assign n9203 = n5907 & ~n9202 ;
  assign n9204 = n9203 ^ n945 ^ 1'b0 ;
  assign n9206 = n5753 ^ n2060 ^ 1'b0 ;
  assign n9205 = n1982 & ~n8276 ;
  assign n9207 = n9206 ^ n9205 ^ 1'b0 ;
  assign n9208 = n9207 ^ n7055 ^ 1'b0 ;
  assign n9209 = n8888 ^ n2733 ^ 1'b0 ;
  assign n9210 = n5234 & ~n9209 ;
  assign n9211 = n2200 & ~n2377 ;
  assign n9212 = n9211 ^ n6955 ^ 1'b0 ;
  assign n9213 = n3940 & ~n7947 ;
  assign n9214 = ~n2766 & n6393 ;
  assign n9215 = ~n1866 & n9214 ;
  assign n9216 = ~n3991 & n9215 ;
  assign n9217 = ~n1789 & n5397 ;
  assign n9218 = n3342 ^ n874 ^ n268 ;
  assign n9219 = n627 & ~n9218 ;
  assign n9220 = n4052 & ~n9219 ;
  assign n9221 = n4347 ^ n1577 ^ 1'b0 ;
  assign n9222 = n9221 ^ n4365 ^ 1'b0 ;
  assign n9223 = n3345 ^ n1139 ^ 1'b0 ;
  assign n9224 = n6577 | n9104 ;
  assign n9225 = n4392 & ~n9224 ;
  assign n9226 = n3473 & ~n6876 ;
  assign n9227 = n9226 ^ n8277 ^ 1'b0 ;
  assign n9228 = ~n1050 & n9227 ;
  assign n9229 = n2754 ^ x6 ^ 1'b0 ;
  assign n9230 = n9228 | n9229 ;
  assign n9231 = n471 | n1022 ;
  assign n9232 = n414 & n4845 ;
  assign n9233 = ~n9231 & n9232 ;
  assign n9234 = ( ~n1471 & n2572 ) | ( ~n1471 & n6438 ) | ( n2572 & n6438 ) ;
  assign n9235 = ( n271 & n7138 ) | ( n271 & n9234 ) | ( n7138 & n9234 ) ;
  assign n9236 = n4319 & ~n5746 ;
  assign n9237 = n2572 ^ n364 ^ 1'b0 ;
  assign n9238 = n66 & ~n3376 ;
  assign n9239 = n2235 & ~n9238 ;
  assign n9240 = n4390 & n9239 ;
  assign n9241 = n3008 ^ n687 ^ 1'b0 ;
  assign n9242 = n144 & n9241 ;
  assign n9243 = n1790 | n4299 ;
  assign n9244 = n2373 & ~n9243 ;
  assign n9245 = n8495 & n9244 ;
  assign n9246 = ~n997 & n9245 ;
  assign n9247 = n9242 & n9246 ;
  assign n9248 = n5899 & ~n9247 ;
  assign n9249 = n5425 & n9248 ;
  assign n9250 = n3415 & ~n9249 ;
  assign n9251 = n9250 ^ n3585 ^ 1'b0 ;
  assign n9252 = n5842 ^ n1166 ^ 1'b0 ;
  assign n9253 = n2606 & n4440 ;
  assign n9254 = ~n610 & n2934 ;
  assign n9256 = n114 & n865 ;
  assign n9257 = n9256 ^ n3150 ^ 1'b0 ;
  assign n9255 = n1835 & n2004 ;
  assign n9258 = n9257 ^ n9255 ^ 1'b0 ;
  assign n9259 = ~n1979 & n9258 ;
  assign n9260 = n8766 & n9259 ;
  assign n9261 = ~n9254 & n9260 ;
  assign n9262 = n1472 & ~n5133 ;
  assign n9263 = ~n7917 & n9262 ;
  assign n9264 = n2826 ^ n273 ^ 1'b0 ;
  assign n9265 = ~n1688 & n9264 ;
  assign n9266 = n443 & ~n1480 ;
  assign n9267 = ~n1105 & n9266 ;
  assign n9268 = n6250 & ~n9267 ;
  assign n9269 = n4671 ^ n4446 ^ 1'b0 ;
  assign n9270 = n556 | n9269 ;
  assign n9271 = n4034 ^ n671 ^ 1'b0 ;
  assign n9272 = n4897 & ~n9271 ;
  assign n9273 = ~n174 & n1802 ;
  assign n9274 = ~n5210 & n9273 ;
  assign n9275 = n9272 | n9274 ;
  assign n9276 = n9275 ^ n375 ^ 1'b0 ;
  assign n9277 = n2996 | n3320 ;
  assign n9278 = x0 | n3228 ;
  assign n9279 = n9278 ^ n3534 ^ 1'b0 ;
  assign n9280 = n9277 & n9279 ;
  assign n9281 = n5180 ^ n257 ^ 1'b0 ;
  assign n9282 = ~n6121 & n9281 ;
  assign n9283 = n3841 ^ n3592 ^ 1'b0 ;
  assign n9284 = n3922 & n9283 ;
  assign n9285 = n1856 & ~n7380 ;
  assign n9286 = ~n1715 & n9285 ;
  assign n9287 = n1137 & n8685 ;
  assign n9288 = ~n6307 & n6846 ;
  assign n9289 = n3925 & n9288 ;
  assign n9290 = n1430 & n1539 ;
  assign n9291 = ~n1713 & n4418 ;
  assign n9292 = n1252 ^ n114 ^ 1'b0 ;
  assign n9293 = n9291 | n9292 ;
  assign n9294 = n9293 ^ n6182 ^ 1'b0 ;
  assign n9295 = n1505 | n6037 ;
  assign n9296 = ~n594 & n9295 ;
  assign n9297 = n1233 ^ n101 ^ 1'b0 ;
  assign n9298 = n7424 | n9297 ;
  assign n9299 = ~n1549 & n5522 ;
  assign n9301 = n1880 ^ n814 ^ 1'b0 ;
  assign n9300 = n1217 | n6787 ;
  assign n9302 = n9301 ^ n9300 ^ 1'b0 ;
  assign n9303 = n155 & ~n277 ;
  assign n9304 = n1895 & n9303 ;
  assign n9305 = ~n3008 & n5034 ;
  assign n9306 = ~n2166 & n9305 ;
  assign n9307 = n622 | n4606 ;
  assign n9308 = n9307 ^ n8130 ^ 1'b0 ;
  assign n9309 = n9306 | n9308 ;
  assign n9310 = ~n55 & n5467 ;
  assign n9311 = n9310 ^ n3613 ^ 1'b0 ;
  assign n9312 = n406 & n9311 ;
  assign n9313 = n9312 ^ n6488 ^ 1'b0 ;
  assign n9315 = n3128 ^ n931 ^ 1'b0 ;
  assign n9314 = n385 & n5950 ;
  assign n9316 = n9315 ^ n9314 ^ 1'b0 ;
  assign n9317 = n754 | n4004 ;
  assign n9318 = n9317 ^ n687 ^ 1'b0 ;
  assign n9319 = ~n94 & n4961 ;
  assign n9320 = n9319 ^ n498 ^ 1'b0 ;
  assign n9321 = ~n9318 & n9320 ;
  assign n9322 = n5065 & n9321 ;
  assign n9323 = n2872 | n3719 ;
  assign n9324 = n9323 ^ n1036 ^ 1'b0 ;
  assign n9325 = ~n1231 & n9324 ;
  assign n9326 = n1910 & ~n4120 ;
  assign n9327 = n9326 ^ n1899 ^ 1'b0 ;
  assign n9328 = n753 ^ n538 ^ 1'b0 ;
  assign n9329 = n1209 & n9328 ;
  assign n9330 = n9329 ^ n241 ^ 1'b0 ;
  assign n9331 = n2196 & ~n9330 ;
  assign n9332 = n9331 ^ n8832 ^ 1'b0 ;
  assign n9333 = n1565 & n2151 ;
  assign n9334 = ( n158 & n3138 ) | ( n158 & n9333 ) | ( n3138 & n9333 ) ;
  assign n9335 = n587 & n1325 ;
  assign n9337 = n4632 ^ n891 ^ 1'b0 ;
  assign n9344 = n2245 & n4485 ;
  assign n9338 = n697 & ~n1854 ;
  assign n9339 = n6280 ^ n1440 ^ 1'b0 ;
  assign n9340 = n9338 & n9339 ;
  assign n9341 = n5180 & n9340 ;
  assign n9342 = n1384 ^ n657 ^ 1'b0 ;
  assign n9343 = n9341 & ~n9342 ;
  assign n9345 = n9344 ^ n9343 ^ 1'b0 ;
  assign n9346 = n9337 | n9345 ;
  assign n9336 = ~n2254 & n3692 ;
  assign n9347 = n9346 ^ n9336 ^ 1'b0 ;
  assign n9348 = n7443 ^ n2263 ^ 1'b0 ;
  assign n9349 = n3507 | n4086 ;
  assign n9350 = n5752 & ~n9349 ;
  assign n9351 = n178 & ~n462 ;
  assign n9352 = n9351 ^ n15 ^ 1'b0 ;
  assign n9353 = n1096 | n5331 ;
  assign n9354 = n178 & ~n9353 ;
  assign n9355 = ( ~n252 & n9352 ) | ( ~n252 & n9354 ) | ( n9352 & n9354 ) ;
  assign n9356 = n37 & ~n458 ;
  assign n9357 = n748 & n9356 ;
  assign n9358 = n367 | n9357 ;
  assign n9359 = n8552 & ~n9358 ;
  assign n9360 = ~n3377 & n8568 ;
  assign n9361 = n4201 ^ n2268 ^ 1'b0 ;
  assign n9362 = n9361 ^ n1552 ^ 1'b0 ;
  assign n9363 = n3003 & ~n9362 ;
  assign n9364 = n5252 | n6133 ;
  assign n9365 = n372 | n9364 ;
  assign n9366 = n9365 ^ n1499 ^ 1'b0 ;
  assign n9367 = n4385 ^ n1194 ^ 1'b0 ;
  assign n9368 = n9366 | n9367 ;
  assign n9369 = n5626 ^ n4207 ^ 1'b0 ;
  assign n9370 = n7767 & ~n9369 ;
  assign n9371 = n4048 & n7444 ;
  assign n9372 = n9371 ^ n5831 ^ 1'b0 ;
  assign n9373 = n7531 ^ n4123 ^ 1'b0 ;
  assign n9374 = n2243 | n5671 ;
  assign n9376 = n6981 ^ n6713 ^ 1'b0 ;
  assign n9377 = n9376 ^ n6424 ^ 1'b0 ;
  assign n9375 = n538 | n3244 ;
  assign n9378 = n9377 ^ n9375 ^ 1'b0 ;
  assign n9379 = n645 & n9378 ;
  assign n9380 = n3492 ^ n2795 ^ 1'b0 ;
  assign n9381 = n3019 & ~n9380 ;
  assign n9382 = n2659 ^ n158 ^ 1'b0 ;
  assign n9383 = n3408 & ~n9382 ;
  assign n9384 = n1731 & n9383 ;
  assign n9385 = n276 & ~n6466 ;
  assign n9388 = n4961 ^ n2489 ^ 1'b0 ;
  assign n9389 = n2511 & ~n9388 ;
  assign n9390 = ~n109 & n9389 ;
  assign n9386 = n6114 | n7490 ;
  assign n9387 = n4042 | n9386 ;
  assign n9391 = n9390 ^ n9387 ^ 1'b0 ;
  assign n9392 = n3097 & n3741 ;
  assign n9393 = n6102 | n9392 ;
  assign n9394 = n9391 & ~n9393 ;
  assign n9395 = n4609 ^ n327 ^ 1'b0 ;
  assign n9396 = ~n551 & n9395 ;
  assign n9397 = n2166 & ~n9234 ;
  assign n9398 = ~n3882 & n4511 ;
  assign n9399 = n2734 & ~n7913 ;
  assign n9400 = n9399 ^ n1426 ^ 1'b0 ;
  assign n9401 = n5160 | n9400 ;
  assign n9402 = ( n8775 & n9398 ) | ( n8775 & n9401 ) | ( n9398 & n9401 ) ;
  assign n9403 = n938 ^ n343 ^ 1'b0 ;
  assign n9404 = x9 & ~n9403 ;
  assign n9405 = ~n2308 & n9404 ;
  assign n9406 = n1764 & n9405 ;
  assign n9407 = n3141 ^ n2672 ^ 1'b0 ;
  assign n9408 = n7862 & ~n9407 ;
  assign n9409 = n738 & ~n8613 ;
  assign n9410 = n7009 ^ n390 ^ 1'b0 ;
  assign n9411 = n8845 & ~n9410 ;
  assign n9412 = n5359 ^ n288 ^ 1'b0 ;
  assign n9413 = n139 & ~n5622 ;
  assign n9414 = n86 | n5141 ;
  assign n9415 = ~n86 & n5187 ;
  assign n9416 = ~n6029 & n9415 ;
  assign n9417 = n1437 | n6080 ;
  assign n9418 = n9417 ^ n5501 ^ 1'b0 ;
  assign n9419 = n8363 | n9418 ;
  assign n9420 = n4140 | n6060 ;
  assign n9421 = ~n852 & n3803 ;
  assign n9422 = n9421 ^ n710 ^ 1'b0 ;
  assign n9423 = n9422 ^ n5113 ^ 1'b0 ;
  assign n9424 = n2757 & ~n9423 ;
  assign n9425 = n9107 ^ n415 ^ n246 ;
  assign n9426 = ~n3669 & n8005 ;
  assign n9427 = ~n4540 & n9426 ;
  assign n9428 = n1201 & n1235 ;
  assign n9429 = n4256 | n9428 ;
  assign n9430 = n9429 ^ n1945 ^ 1'b0 ;
  assign n9431 = n9427 | n9430 ;
  assign n9432 = n8721 & n9431 ;
  assign n9433 = n1236 & ~n5000 ;
  assign n9434 = ~n4284 & n9433 ;
  assign n9435 = ~n442 & n6181 ;
  assign n9436 = n9435 ^ n7488 ^ 1'b0 ;
  assign n9437 = n5123 | n9436 ;
  assign n9438 = n9437 ^ n4346 ^ 1'b0 ;
  assign n9439 = ~n1227 & n9438 ;
  assign n9440 = ~n1229 & n6127 ;
  assign n9441 = n9440 ^ n1760 ^ 1'b0 ;
  assign n9442 = ~n9439 & n9441 ;
  assign n9443 = ~n259 & n6809 ;
  assign n9444 = n7667 & n9443 ;
  assign n9445 = ~n454 & n5785 ;
  assign n9446 = n6755 & n9445 ;
  assign n9447 = n6514 ^ n426 ^ n175 ;
  assign n9448 = n7701 ^ n359 ^ 1'b0 ;
  assign n9449 = n1345 | n5382 ;
  assign n9450 = n9449 ^ n6121 ^ 1'b0 ;
  assign n9451 = n2969 & n9450 ;
  assign n9452 = n2811 | n8714 ;
  assign n9456 = n42 | n102 ;
  assign n9457 = n102 & ~n9456 ;
  assign n9458 = n183 & ~n9457 ;
  assign n9459 = ~n183 & n9458 ;
  assign n9453 = n1768 & n4063 ;
  assign n9454 = ~n1768 & n9453 ;
  assign n9455 = n587 & n9454 ;
  assign n9460 = n9459 ^ n9455 ^ 1'b0 ;
  assign n9466 = ~n68 & n581 ;
  assign n9467 = n68 & n9466 ;
  assign n9468 = ~n5691 & n9467 ;
  assign n9462 = n788 & n1390 ;
  assign n9463 = ~n1300 & n9462 ;
  assign n9464 = n7814 & ~n9463 ;
  assign n9465 = n9463 & n9464 ;
  assign n9469 = n9468 ^ n9465 ^ 1'b0 ;
  assign n9461 = n2302 | n3037 ;
  assign n9470 = n9469 ^ n9461 ^ 1'b0 ;
  assign n9471 = n9460 & n9470 ;
  assign n9472 = n2961 ^ n472 ^ 1'b0 ;
  assign n9473 = n3997 & n9472 ;
  assign n9474 = n9473 ^ n2083 ^ 1'b0 ;
  assign n9475 = n1375 ^ n593 ^ 1'b0 ;
  assign n9476 = x6 & n9475 ;
  assign n9477 = n1316 & ~n7981 ;
  assign n9478 = ~n9476 & n9477 ;
  assign n9479 = n9474 & ~n9478 ;
  assign n9480 = n5376 ^ n2542 ^ 1'b0 ;
  assign n9481 = n3056 | n9480 ;
  assign n9482 = n9481 ^ n363 ^ 1'b0 ;
  assign n9483 = n6450 & ~n9482 ;
  assign n9484 = n6168 ^ n5528 ^ 1'b0 ;
  assign n9485 = n336 & ~n4493 ;
  assign n9486 = n9485 ^ n3392 ^ 1'b0 ;
  assign n9487 = n4100 & n9486 ;
  assign n9488 = ~n9484 & n9487 ;
  assign n9489 = n9488 ^ n2891 ^ 1'b0 ;
  assign n9490 = n4240 & n9489 ;
  assign n9491 = n5451 ^ n506 ^ 1'b0 ;
  assign n9493 = n3640 ^ n190 ^ 1'b0 ;
  assign n9494 = n1316 & ~n9493 ;
  assign n9492 = n2348 ^ n566 ^ n55 ;
  assign n9495 = n9494 ^ n9492 ^ 1'b0 ;
  assign n9496 = ( n38 & n3219 ) | ( n38 & ~n7185 ) | ( n3219 & ~n7185 ) ;
  assign n9497 = n7247 ^ n662 ^ 1'b0 ;
  assign n9498 = ~n7358 & n9497 ;
  assign n9499 = n2243 ^ n1874 ^ 1'b0 ;
  assign n9500 = n2062 & n9499 ;
  assign n9501 = n9500 ^ n3931 ^ 1'b0 ;
  assign n9502 = n9501 ^ n7791 ^ n3007 ;
  assign n9503 = n2136 ^ n1529 ^ 1'b0 ;
  assign n9504 = n205 & ~n9503 ;
  assign n9505 = n7599 & n9504 ;
  assign n9506 = n9505 ^ n4904 ^ 1'b0 ;
  assign n9507 = n2478 | n6809 ;
  assign n9508 = n5495 ^ n1132 ^ 1'b0 ;
  assign n9509 = n7009 | n9508 ;
  assign n9510 = n9509 ^ n618 ^ 1'b0 ;
  assign n9511 = n7312 ^ n2376 ^ 1'b0 ;
  assign n9512 = n3765 | n9511 ;
  assign n9513 = n1127 & ~n9112 ;
  assign n9514 = n9513 ^ n2370 ^ 1'b0 ;
  assign n9515 = n2513 & ~n6419 ;
  assign n9516 = n6218 & n9515 ;
  assign n9517 = ~n5067 & n8523 ;
  assign n9518 = n9517 ^ n5771 ^ 1'b0 ;
  assign n9519 = n1632 & ~n8725 ;
  assign n9520 = ~n488 & n9519 ;
  assign n9521 = n9193 ^ n2510 ^ 1'b0 ;
  assign n9522 = ~n4551 & n7340 ;
  assign n9523 = ~n3521 & n9522 ;
  assign n9524 = ( ~n879 & n2017 ) | ( ~n879 & n2738 ) | ( n2017 & n2738 ) ;
  assign n9525 = n2572 ^ n252 ^ 1'b0 ;
  assign n9526 = n7336 | n9525 ;
  assign n9527 = n8097 | n9526 ;
  assign n9528 = n107 | n3452 ;
  assign n9529 = n8967 ^ n3325 ^ 1'b0 ;
  assign n9530 = n7952 | n9529 ;
  assign n9531 = n1246 & n2636 ;
  assign n9533 = n470 | n3273 ;
  assign n9534 = n9533 ^ n6295 ^ 1'b0 ;
  assign n9532 = n2509 & n4887 ;
  assign n9535 = n9534 ^ n9532 ^ 1'b0 ;
  assign n9536 = n9531 | n9535 ;
  assign n9537 = n622 ^ n215 ^ 1'b0 ;
  assign n9538 = ~n1637 & n9537 ;
  assign n9539 = n3499 & n9538 ;
  assign n9540 = n135 & ~n7661 ;
  assign n9541 = ~n9539 & n9540 ;
  assign n9542 = n7500 & n9541 ;
  assign n9544 = n5317 & n7457 ;
  assign n9543 = n7545 & n9131 ;
  assign n9545 = n9544 ^ n9543 ^ 1'b0 ;
  assign n9546 = n1449 & ~n2176 ;
  assign n9547 = n8872 ^ n4111 ^ 1'b0 ;
  assign n9548 = n4848 & n9547 ;
  assign n9549 = n3120 & n8088 ;
  assign n9550 = n5913 ^ n1388 ^ 1'b0 ;
  assign n9551 = ~n3273 & n7060 ;
  assign n9552 = ~n2204 & n3601 ;
  assign n9553 = n1974 | n4171 ;
  assign n9554 = n9553 ^ n52 ^ 1'b0 ;
  assign n9555 = n2446 | n5666 ;
  assign n9556 = n9554 | n9555 ;
  assign n9557 = n4367 | n9556 ;
  assign n9558 = n4560 ^ n2501 ^ 1'b0 ;
  assign n9559 = ~n859 & n9558 ;
  assign n9560 = n2497 & ~n2915 ;
  assign n9561 = n9560 ^ n2594 ^ 1'b0 ;
  assign n9562 = n2330 & n4227 ;
  assign n9563 = n139 & ~n1138 ;
  assign n9564 = ~n756 & n9563 ;
  assign n9565 = ~n934 & n4228 ;
  assign n9566 = ~n276 & n6089 ;
  assign n9567 = n414 & n928 ;
  assign n9568 = n9566 & ~n9567 ;
  assign n9569 = ~n9565 & n9568 ;
  assign n9570 = n1718 | n2117 ;
  assign n9571 = n9570 ^ n7860 ^ 1'b0 ;
  assign n9572 = ~n2090 & n4882 ;
  assign n9573 = n958 ^ n50 ^ 1'b0 ;
  assign n9574 = n1458 | n4879 ;
  assign n9575 = n2092 & ~n9574 ;
  assign n9576 = ( n2244 & n2476 ) | ( n2244 & n7353 ) | ( n2476 & n7353 ) ;
  assign n9577 = n434 & n6485 ;
  assign n9578 = n9577 ^ n2493 ^ 1'b0 ;
  assign n9579 = n3929 ^ n1768 ^ 1'b0 ;
  assign n9580 = n322 | n9579 ;
  assign n9581 = n5967 ^ n3051 ^ 1'b0 ;
  assign n9582 = n4249 | n5002 ;
  assign n9583 = n8062 & n9582 ;
  assign n9584 = n4784 ^ n1250 ^ 1'b0 ;
  assign n9585 = n3798 & ~n9584 ;
  assign n9586 = n4830 | n9585 ;
  assign n9587 = n2127 | n2511 ;
  assign n9588 = n9587 ^ n5180 ^ 1'b0 ;
  assign n9589 = n9588 ^ n3156 ^ 1'b0 ;
  assign n9590 = n750 ^ n709 ^ 1'b0 ;
  assign n9591 = n323 & ~n3512 ;
  assign n9592 = n1865 ^ n369 ^ 1'b0 ;
  assign n9593 = n9592 ^ n3204 ^ 1'b0 ;
  assign n9594 = n8910 & n9593 ;
  assign n9595 = n8558 ^ n2136 ^ 1'b0 ;
  assign n9596 = n116 | n2789 ;
  assign n9597 = n825 | n3315 ;
  assign n9598 = n2905 ^ n741 ^ 1'b0 ;
  assign n9599 = n1601 | n9598 ;
  assign n9600 = n3462 | n9599 ;
  assign n9601 = n9600 ^ n9499 ^ 1'b0 ;
  assign n9602 = n7811 | n9601 ;
  assign n9603 = n1130 & ~n3204 ;
  assign n9604 = n9603 ^ n8106 ^ 1'b0 ;
  assign n9605 = n452 | n9604 ;
  assign n9606 = n5443 | n9605 ;
  assign n9607 = ~n2431 & n4739 ;
  assign n9608 = n5200 ^ n3873 ^ n1219 ;
  assign n9609 = n3589 & ~n9608 ;
  assign n9610 = n9607 | n9609 ;
  assign n9611 = ~n1552 & n3539 ;
  assign n9612 = n883 ^ n636 ^ 1'b0 ;
  assign n9613 = n1010 & n9612 ;
  assign n9614 = n7730 ^ n4048 ^ 1'b0 ;
  assign n9615 = n7665 ^ n7483 ^ 1'b0 ;
  assign n9616 = n1502 & ~n9615 ;
  assign n9617 = n6852 & ~n7956 ;
  assign n9618 = n4815 ^ n1401 ^ 1'b0 ;
  assign n9619 = n435 & ~n9618 ;
  assign n9620 = ( n1707 & ~n5752 ) | ( n1707 & n9619 ) | ( ~n5752 & n9619 ) ;
  assign n9621 = n2913 ^ n1193 ^ 1'b0 ;
  assign n9622 = n104 & ~n561 ;
  assign n9623 = ~n9621 & n9622 ;
  assign n9624 = n8411 ^ n3681 ^ 1'b0 ;
  assign n9625 = n3431 & n9624 ;
  assign n9626 = ~n46 & n7666 ;
  assign n9629 = n3581 ^ n1174 ^ 1'b0 ;
  assign n9630 = n6268 ^ n2277 ^ 1'b0 ;
  assign n9631 = n2704 | n9630 ;
  assign n9632 = n9629 & n9631 ;
  assign n9633 = n4570 & n9632 ;
  assign n9627 = ~n2779 & n8241 ;
  assign n9628 = n5422 & ~n9627 ;
  assign n9634 = n9633 ^ n9628 ^ 1'b0 ;
  assign n9635 = ~n764 & n867 ;
  assign n9636 = n5078 | n6581 ;
  assign n9637 = n9636 ^ n3583 ^ 1'b0 ;
  assign n9638 = n9635 & ~n9637 ;
  assign n9639 = n8242 ^ n2022 ^ 1'b0 ;
  assign n9640 = n1372 & ~n9639 ;
  assign n9641 = n9640 ^ n3715 ^ 1'b0 ;
  assign n9642 = n497 & ~n6426 ;
  assign n9643 = n9641 & n9642 ;
  assign n9644 = n4390 ^ n3890 ^ 1'b0 ;
  assign n9645 = ~n357 & n9644 ;
  assign n9646 = ~n3221 & n5769 ;
  assign n9647 = n4403 & ~n8469 ;
  assign n9648 = n1129 ^ n738 ^ 1'b0 ;
  assign n9649 = n5461 & n9648 ;
  assign n9650 = n9649 ^ n1802 ^ 1'b0 ;
  assign n9651 = n527 & ~n9650 ;
  assign n9652 = ~n461 & n883 ;
  assign n9653 = n4241 & n4819 ;
  assign n9654 = n2829 & n9653 ;
  assign n9655 = n9654 ^ n3293 ^ n1026 ;
  assign n9656 = n7285 & n9655 ;
  assign n9657 = n9656 ^ n5380 ^ 1'b0 ;
  assign n9658 = n7046 ^ n3044 ^ 1'b0 ;
  assign n9659 = ~n1575 & n9658 ;
  assign n9660 = n7688 ^ n323 ^ 1'b0 ;
  assign n9661 = n142 | n2078 ;
  assign n9662 = n8613 ^ n3579 ^ n827 ;
  assign n9663 = n4271 ^ n3492 ^ 1'b0 ;
  assign n9664 = n5574 ^ n1388 ^ 1'b0 ;
  assign n9665 = ~n257 & n9664 ;
  assign n9666 = n4966 ^ n4581 ^ 1'b0 ;
  assign n9667 = n86 & ~n9666 ;
  assign n9668 = ~n9665 & n9667 ;
  assign n9669 = n8917 ^ n241 ^ n159 ;
  assign n9670 = n4763 & ~n9669 ;
  assign n9671 = n2417 & n9670 ;
  assign n9672 = n1315 & n9671 ;
  assign n9673 = n6647 ^ n254 ^ 1'b0 ;
  assign n9674 = n6192 ^ n5015 ^ 1'b0 ;
  assign n9675 = ~n146 & n9674 ;
  assign n9676 = n9675 ^ n1716 ^ 1'b0 ;
  assign n9677 = n9673 & n9676 ;
  assign n9679 = n1186 & n6282 ;
  assign n9680 = n6974 & n9679 ;
  assign n9681 = ~n2680 & n4296 ;
  assign n9682 = n9680 & n9681 ;
  assign n9683 = n9682 ^ n5995 ^ 1'b0 ;
  assign n9678 = n271 & ~n1693 ;
  assign n9684 = n9683 ^ n9678 ^ 1'b0 ;
  assign n9686 = ~n2885 & n5332 ;
  assign n9687 = n9686 ^ n1355 ^ 1'b0 ;
  assign n9688 = ~n9118 & n9687 ;
  assign n9685 = n259 | n2611 ;
  assign n9689 = n9688 ^ n9685 ^ 1'b0 ;
  assign n9690 = n4098 | n4904 ;
  assign n9691 = n1044 & ~n9690 ;
  assign n9692 = n246 ^ n177 ^ 1'b0 ;
  assign n9693 = n4593 & n8465 ;
  assign n9694 = ~n3204 & n9693 ;
  assign n9695 = n2734 & n9694 ;
  assign n9696 = n9692 | n9695 ;
  assign n9697 = n4620 ^ n3185 ^ n153 ;
  assign n9698 = n4069 & ~n9697 ;
  assign n9699 = n6023 & n6897 ;
  assign n9700 = ~n5310 & n6023 ;
  assign n9701 = ~n1304 & n9700 ;
  assign n9702 = n9699 & n9701 ;
  assign n9703 = ~n2426 & n7278 ;
  assign n9704 = n3291 & n5194 ;
  assign n9705 = ~n203 & n9704 ;
  assign n9706 = n1203 & ~n4838 ;
  assign n9707 = n131 & n9706 ;
  assign n9708 = n6349 & ~n9707 ;
  assign n9709 = n9708 ^ n3939 ^ 1'b0 ;
  assign n9710 = n321 & ~n1790 ;
  assign n9711 = n9709 | n9710 ;
  assign n9712 = n6189 | n9711 ;
  assign n9713 = n7103 ^ n3939 ^ 1'b0 ;
  assign n9714 = n8269 ^ n2568 ^ n1533 ;
  assign n9715 = n9714 ^ n1385 ^ 1'b0 ;
  assign n9716 = n6360 | n7188 ;
  assign n9717 = n683 & ~n9716 ;
  assign n9718 = n4422 ^ n141 ^ 1'b0 ;
  assign n9721 = n5053 ^ n4439 ^ 1'b0 ;
  assign n9719 = n3837 | n8392 ;
  assign n9720 = ~n6849 & n9719 ;
  assign n9722 = n9721 ^ n9720 ^ 1'b0 ;
  assign n9723 = n5785 ^ n1476 ^ 1'b0 ;
  assign n9724 = ~n7570 & n7593 ;
  assign n9725 = n9724 ^ n2757 ^ 1'b0 ;
  assign n9726 = n9419 ^ n5465 ^ 1'b0 ;
  assign n9727 = ~n684 & n4451 ;
  assign n9728 = ~n357 & n7056 ;
  assign n9729 = n2826 ^ n962 ^ 1'b0 ;
  assign n9730 = n9728 | n9729 ;
  assign n9731 = ~x2 & n7391 ;
  assign n9732 = n9731 ^ n2523 ^ 1'b0 ;
  assign n9733 = ~n9255 & n9732 ;
  assign n9734 = n7550 ^ n6374 ^ 1'b0 ;
  assign n9735 = n9734 ^ n1169 ^ 1'b0 ;
  assign n9736 = ~n4320 & n9735 ;
  assign n9737 = n9727 ^ n7325 ^ 1'b0 ;
  assign n9738 = n1390 ^ n1198 ^ 1'b0 ;
  assign n9739 = n2856 & ~n9738 ;
  assign n9740 = ~n6417 & n9739 ;
  assign n9741 = ~n3101 & n9740 ;
  assign n9742 = n954 ^ n60 ^ 1'b0 ;
  assign n9743 = ~n2846 & n9742 ;
  assign n9744 = n1104 & ~n4619 ;
  assign n9745 = n169 & ~n4619 ;
  assign n9746 = ~n257 & n9745 ;
  assign n9747 = n86 | n359 ;
  assign n9748 = n9747 ^ n2975 ^ 1'b0 ;
  assign n9749 = n1713 & ~n3514 ;
  assign n9750 = ~n9748 & n9749 ;
  assign n9751 = n9750 ^ n400 ^ 1'b0 ;
  assign n9753 = n2577 ^ n598 ^ 1'b0 ;
  assign n9752 = n1081 & ~n6009 ;
  assign n9754 = n9753 ^ n9752 ^ 1'b0 ;
  assign n9755 = n252 | n3626 ;
  assign n9756 = n9755 ^ n1472 ^ 1'b0 ;
  assign n9757 = ~n1226 & n5723 ;
  assign n9758 = n6660 ^ n774 ^ 1'b0 ;
  assign n9759 = n9758 ^ n419 ^ 1'b0 ;
  assign n9760 = ~n5586 & n7195 ;
  assign n9762 = n1917 & n2624 ;
  assign n9763 = n460 & n9762 ;
  assign n9761 = n270 | n5956 ;
  assign n9764 = n9763 ^ n9761 ^ 1'b0 ;
  assign n9765 = n6114 & n6137 ;
  assign n9766 = n1444 & ~n2375 ;
  assign n9767 = ~n1250 & n9766 ;
  assign n9768 = n3171 & n9767 ;
  assign n9769 = n536 ^ n294 ^ 1'b0 ;
  assign n9770 = n9768 & n9769 ;
  assign n9771 = n4906 & n8353 ;
  assign n9775 = n367 ^ x0 ^ 1'b0 ;
  assign n9772 = n3985 & n8832 ;
  assign n9773 = n9772 ^ n8918 ^ 1'b0 ;
  assign n9774 = ~n1469 & n9773 ;
  assign n9776 = n9775 ^ n9774 ^ 1'b0 ;
  assign n9777 = n2551 & ~n5241 ;
  assign n9778 = n2155 & n9777 ;
  assign n9779 = n799 | n3917 ;
  assign n9780 = n9779 ^ n9120 ^ 1'b0 ;
  assign n9781 = n9780 ^ n8163 ^ n1213 ;
  assign n9782 = ~n4700 & n7286 ;
  assign n9783 = ~n7286 & n9782 ;
  assign n9784 = n4057 ^ n16 ^ 1'b0 ;
  assign n9785 = n1117 | n9784 ;
  assign n9786 = n9785 ^ n3709 ^ 1'b0 ;
  assign n9787 = ~n9783 & n9786 ;
  assign n9788 = ~n1608 & n8717 ;
  assign n9789 = n7771 & n9788 ;
  assign n9790 = n117 | n2543 ;
  assign n9791 = n1521 & ~n9790 ;
  assign n9792 = ( n1129 & ~n1360 ) | ( n1129 & n2859 ) | ( ~n1360 & n2859 ) ;
  assign n9793 = ~n403 & n9792 ;
  assign n9794 = ~n1474 & n3651 ;
  assign n9795 = n4129 ^ n3305 ^ 1'b0 ;
  assign n9796 = ~n3514 & n9795 ;
  assign n9797 = n3600 | n7102 ;
  assign n9798 = ~n3276 & n9797 ;
  assign n9799 = n9798 ^ n4223 ^ 1'b0 ;
  assign n9800 = n2849 ^ n1326 ^ 1'b0 ;
  assign n9801 = n9800 ^ n338 ^ 1'b0 ;
  assign n9802 = n3217 & n3430 ;
  assign n9803 = n1320 | n4331 ;
  assign n9804 = n9803 ^ n8720 ^ 1'b0 ;
  assign n9805 = n9804 ^ n9177 ^ 1'b0 ;
  assign n9806 = n3598 ^ n878 ^ 1'b0 ;
  assign n9807 = n1431 & ~n3071 ;
  assign n9808 = n9807 ^ n2406 ^ 1'b0 ;
  assign n9809 = n3694 | n7553 ;
  assign n9810 = n9808 & n9809 ;
  assign n9811 = ( n128 & ~n3775 ) | ( n128 & n5372 ) | ( ~n3775 & n5372 ) ;
  assign n9812 = n85 & ~n9811 ;
  assign n9813 = n4074 & ~n9812 ;
  assign n9814 = n4785 & n9813 ;
  assign n9815 = n3199 ^ n670 ^ 1'b0 ;
  assign n9816 = ~n1769 & n9815 ;
  assign n9817 = n7192 & ~n7239 ;
  assign n9819 = n853 | n1835 ;
  assign n9820 = n2912 ^ n2839 ^ 1'b0 ;
  assign n9821 = n9819 | n9820 ;
  assign n9818 = n2955 & ~n8499 ;
  assign n9822 = n9821 ^ n9818 ^ 1'b0 ;
  assign n9823 = ( ~n2898 & n4697 ) | ( ~n2898 & n8141 ) | ( n4697 & n8141 ) ;
  assign n9824 = n3781 & ~n9823 ;
  assign n9826 = n1130 & ~n5535 ;
  assign n9825 = n3138 | n8169 ;
  assign n9827 = n9826 ^ n9825 ^ 1'b0 ;
  assign n9828 = n907 & n5643 ;
  assign n9829 = n3071 ^ n2281 ^ 1'b0 ;
  assign n9830 = n1961 ^ n257 ^ 1'b0 ;
  assign n9831 = ~n1740 & n9830 ;
  assign n9832 = ~n926 & n9831 ;
  assign n9833 = n5542 & ~n9832 ;
  assign n9834 = ~n1848 & n9833 ;
  assign n9835 = n7368 & n9834 ;
  assign n9836 = n9560 ^ n378 ^ 1'b0 ;
  assign n9837 = n2598 & ~n5621 ;
  assign n9838 = n7355 | n9837 ;
  assign n9839 = n5207 ^ n328 ^ 1'b0 ;
  assign n9840 = n1169 & n9839 ;
  assign n9841 = n8822 & ~n9840 ;
  assign n9842 = n9746 ^ n5383 ^ 1'b0 ;
  assign n9843 = n9211 & n9842 ;
  assign n9844 = n1373 & ~n3632 ;
  assign n9845 = n6209 | n9844 ;
  assign n9847 = n6194 ^ n1609 ^ 1'b0 ;
  assign n9846 = n226 & ~n4037 ;
  assign n9848 = n9847 ^ n9846 ^ 1'b0 ;
  assign n9849 = n1051 & ~n5827 ;
  assign n9850 = n6335 & n9849 ;
  assign n9851 = n7529 ^ n6698 ^ 1'b0 ;
  assign n9852 = n7023 ^ n2273 ^ 1'b0 ;
  assign n9853 = ~n628 & n4819 ;
  assign n9854 = n9853 ^ n3569 ^ 1'b0 ;
  assign n9855 = n3921 & ~n9854 ;
  assign n9856 = ~n6771 & n9045 ;
  assign n9857 = n9856 ^ n1355 ^ 1'b0 ;
  assign n9858 = ~n158 & n3267 ;
  assign n9859 = n8667 ^ n1159 ^ 1'b0 ;
  assign n9860 = n4668 ^ n1369 ^ 1'b0 ;
  assign n9861 = n3202 | n9860 ;
  assign n9862 = n5217 & ~n9861 ;
  assign n9863 = ~n42 & n226 ;
  assign n9864 = ~n226 & n9863 ;
  assign n9865 = n5741 | n9864 ;
  assign n9866 = n5741 & ~n9865 ;
  assign n9867 = n9866 ^ n2282 ^ 1'b0 ;
  assign n9868 = n939 & ~n1418 ;
  assign n9869 = n7894 ^ n165 ^ 1'b0 ;
  assign n9870 = ~n2038 & n9869 ;
  assign n9871 = n366 & n3907 ;
  assign n9872 = n9871 ^ n5146 ^ 1'b0 ;
  assign n9873 = n4703 & n6433 ;
  assign n9874 = n3065 ^ n3005 ^ 1'b0 ;
  assign n9875 = ~n7315 & n9874 ;
  assign n9876 = n1740 & ~n2107 ;
  assign n9877 = n9876 ^ n1880 ^ 1'b0 ;
  assign n9878 = n9877 ^ n1332 ^ 1'b0 ;
  assign n9879 = n9875 & ~n9878 ;
  assign n9880 = ~n5932 & n9879 ;
  assign n9881 = n744 ^ n37 ^ 1'b0 ;
  assign n9882 = n9881 ^ n2510 ^ 1'b0 ;
  assign n9883 = n4123 ^ n3503 ^ 1'b0 ;
  assign n9884 = n4233 ^ n615 ^ 1'b0 ;
  assign n9885 = n8800 ^ n7649 ^ n308 ;
  assign n9886 = n8223 ^ n5926 ^ 1'b0 ;
  assign n9887 = n8433 & n9886 ;
  assign n9888 = ~n9885 & n9887 ;
  assign n9889 = ~n60 & n141 ;
  assign n9890 = ( n4163 & ~n9571 ) | ( n4163 & n9889 ) | ( ~n9571 & n9889 ) ;
  assign n9891 = n1235 & ~n6277 ;
  assign n9892 = n9891 ^ n552 ^ 1'b0 ;
  assign n9893 = n1406 & n7814 ;
  assign n9894 = ~n8453 & n9893 ;
  assign n9895 = n633 | n1165 ;
  assign n9896 = n6163 ^ n4034 ^ 1'b0 ;
  assign n9897 = n1254 & ~n9896 ;
  assign n9898 = n9897 ^ n84 ^ 1'b0 ;
  assign n9899 = n812 & ~n9898 ;
  assign n9900 = n46 | n9527 ;
  assign n9901 = n6827 | n6958 ;
  assign n9902 = n1155 ^ n883 ^ 1'b0 ;
  assign n9903 = n2770 & n9902 ;
  assign n9904 = n9903 ^ n6769 ^ 1'b0 ;
  assign n9905 = ~n5065 & n9904 ;
  assign n9906 = ~n3471 & n6850 ;
  assign n9907 = n2235 & n9341 ;
  assign n9908 = n9907 ^ n4772 ^ 1'b0 ;
  assign n9909 = n9906 & n9908 ;
  assign n9910 = n9909 ^ n8545 ^ 1'b0 ;
  assign n9912 = n154 & ~n1885 ;
  assign n9913 = n35 & n9912 ;
  assign n9911 = n1833 & n6416 ;
  assign n9914 = n9913 ^ n9911 ^ 1'b0 ;
  assign n9915 = n3227 ^ n1584 ^ n76 ;
  assign n9916 = n9915 ^ n16 ^ 1'b0 ;
  assign n9917 = n9914 & n9916 ;
  assign n9918 = n390 | n2722 ;
  assign n9919 = n9918 ^ n8254 ^ 1'b0 ;
  assign n9920 = n2959 & n9919 ;
  assign n9921 = n6062 & n9920 ;
  assign n9922 = ~n9917 & n9921 ;
  assign n9923 = n4697 ^ n2941 ^ 1'b0 ;
  assign n9924 = ~n754 & n4220 ;
  assign n9925 = ~n3290 & n9924 ;
  assign n9926 = n1048 | n5217 ;
  assign n9927 = n9926 ^ n807 ^ 1'b0 ;
  assign n9928 = n9927 ^ n3389 ^ 1'b0 ;
  assign n9929 = n3390 & ~n9928 ;
  assign n9930 = n9925 & n9929 ;
  assign n9931 = n7383 ^ n6397 ^ 1'b0 ;
  assign n9932 = n9775 ^ n5309 ^ 1'b0 ;
  assign n9933 = ~n3613 & n9932 ;
  assign n9934 = ~n339 & n9933 ;
  assign n9935 = n5905 ^ n1790 ^ 1'b0 ;
  assign n9936 = n950 | n4273 ;
  assign n9937 = n9936 ^ n461 ^ 1'b0 ;
  assign n9938 = n4485 ^ n2556 ^ 1'b0 ;
  assign n9939 = ~n9937 & n9938 ;
  assign n9940 = n9939 ^ n6215 ^ n2165 ;
  assign n9941 = n908 | n6335 ;
  assign n9942 = n633 | n5328 ;
  assign n9943 = n203 & n609 ;
  assign n9944 = ~n203 & n9943 ;
  assign n9945 = n527 & ~n9944 ;
  assign n9946 = n89 & n1100 ;
  assign n9947 = ~n1100 & n9946 ;
  assign n9948 = n527 & n1331 ;
  assign n9949 = ~n527 & n9948 ;
  assign n9950 = n2642 & ~n9949 ;
  assign n9951 = ( n9945 & n9947 ) | ( n9945 & n9950 ) | ( n9947 & n9950 ) ;
  assign n9952 = ~n872 & n8165 ;
  assign n9953 = n9952 ^ n1807 ^ 1'b0 ;
  assign n9954 = n577 & ~n9953 ;
  assign n9955 = n760 & ~n9954 ;
  assign n9956 = n5626 & ~n7483 ;
  assign n9957 = n9956 ^ n3699 ^ 1'b0 ;
  assign n9958 = n3304 & ~n5801 ;
  assign n9959 = n9958 ^ n4269 ^ 1'b0 ;
  assign n9960 = n3679 ^ n1129 ^ 1'b0 ;
  assign n9961 = n1316 & ~n9960 ;
  assign n9962 = n1669 & n8622 ;
  assign n9963 = n9962 ^ n6998 ^ 1'b0 ;
  assign n9964 = ~n8572 & n9963 ;
  assign n9965 = n7865 ^ n6536 ^ 1'b0 ;
  assign n9966 = n2519 | n3360 ;
  assign n9967 = n247 & ~n3891 ;
  assign n9968 = n8059 & n9967 ;
  assign n9969 = n9968 ^ n5040 ^ 1'b0 ;
  assign n9970 = n3340 & ~n6487 ;
  assign n9971 = n9970 ^ n6579 ^ 1'b0 ;
  assign n9972 = n1441 & n2995 ;
  assign n9973 = ~n7942 & n9972 ;
  assign n9974 = n2335 ^ n205 ^ 1'b0 ;
  assign n9975 = n2216 & ~n9974 ;
  assign n9976 = ~n5887 & n9975 ;
  assign n9977 = n9976 ^ n2046 ^ 1'b0 ;
  assign n9978 = n5775 & ~n9977 ;
  assign n9979 = ( n1394 & n9973 ) | ( n1394 & n9978 ) | ( n9973 & n9978 ) ;
  assign n9980 = n108 & ~n880 ;
  assign n9981 = ~n144 & n9980 ;
  assign n9982 = n3690 | n7846 ;
  assign n9983 = n6397 & ~n8477 ;
  assign n9984 = ~n1388 & n3498 ;
  assign n9985 = ~n8614 & n9984 ;
  assign n9986 = n5067 ^ n404 ^ 1'b0 ;
  assign n9987 = n8056 & ~n9986 ;
  assign n9988 = n5415 ^ n438 ^ 1'b0 ;
  assign n9989 = ~n5104 & n9734 ;
  assign n9990 = n6168 ^ n3007 ^ 1'b0 ;
  assign n9991 = n1194 & ~n4882 ;
  assign n9992 = ~n5957 & n8347 ;
  assign n9993 = n4790 ^ n62 ^ 1'b0 ;
  assign n9994 = n3826 & n9993 ;
  assign n9995 = n4013 ^ n3599 ^ 1'b0 ;
  assign n9996 = n9994 & ~n9995 ;
  assign n9997 = n6148 ^ n5110 ^ 1'b0 ;
  assign n9998 = n1959 | n9997 ;
  assign n9999 = n8165 ^ n7013 ^ 1'b0 ;
  assign n10000 = n4848 & n8251 ;
  assign n10001 = n290 & n1185 ;
  assign n10002 = ~n2898 & n4991 ;
  assign n10003 = n10002 ^ n113 ^ 1'b0 ;
  assign n10004 = n10001 | n10003 ;
  assign n10005 = n10004 ^ n5447 ^ 1'b0 ;
  assign n10006 = n1254 & ~n9785 ;
  assign n10007 = n10006 ^ n8763 ^ 1'b0 ;
  assign n10008 = n5968 & ~n6417 ;
  assign n10009 = ~n333 & n10008 ;
  assign n10010 = n9860 | n10009 ;
  assign n10011 = n10007 & ~n10010 ;
  assign n10012 = n5363 ^ n2333 ^ n539 ;
  assign n10013 = n10012 ^ n1499 ^ 1'b0 ;
  assign n10014 = n509 | n10013 ;
  assign n10015 = n861 & ~n2270 ;
  assign n10016 = n4492 & n10015 ;
  assign n10017 = n10016 ^ n461 ^ 1'b0 ;
  assign n10018 = n10014 & ~n10017 ;
  assign n10020 = n757 | n905 ;
  assign n10021 = n10020 ^ n2400 ^ n1530 ;
  assign n10019 = n3641 ^ n1233 ^ 1'b0 ;
  assign n10022 = n10021 ^ n10019 ^ 1'b0 ;
  assign n10023 = n8945 ^ n665 ^ 1'b0 ;
  assign n10024 = n10022 & n10023 ;
  assign n10025 = n456 ^ x3 ^ 1'b0 ;
  assign n10026 = n273 & ~n10025 ;
  assign n10027 = n3266 & ~n4044 ;
  assign n10028 = n10027 ^ n1090 ^ 1'b0 ;
  assign n10029 = n3038 & ~n10028 ;
  assign n10030 = n10029 ^ n1162 ^ 1'b0 ;
  assign n10031 = n3545 & n4642 ;
  assign n10032 = n1825 | n5797 ;
  assign n10033 = n3301 ^ n2545 ^ 1'b0 ;
  assign n10034 = ~n1198 & n10033 ;
  assign n10035 = n10034 ^ n4040 ^ 1'b0 ;
  assign n10036 = n10035 ^ n461 ^ 1'b0 ;
  assign n10037 = n2519 & n4264 ;
  assign n10038 = n1870 & n4462 ;
  assign n10039 = ~n10037 & n10038 ;
  assign n10040 = ~n3778 & n10039 ;
  assign n10041 = ~n1758 & n5068 ;
  assign n10042 = n4439 | n6830 ;
  assign n10043 = n1771 & ~n10042 ;
  assign n10044 = n4560 ^ n3027 ^ 1'b0 ;
  assign n10045 = n492 | n6212 ;
  assign n10046 = n3290 | n10045 ;
  assign n10047 = ~n3782 & n5731 ;
  assign n10048 = n2885 ^ n55 ^ 1'b0 ;
  assign n10049 = n4781 ^ n2073 ^ 1'b0 ;
  assign n10050 = n7064 & ~n10049 ;
  assign n10051 = n8350 & n10050 ;
  assign n10052 = n5955 & n10051 ;
  assign n10053 = n4941 ^ n4572 ^ 1'b0 ;
  assign n10054 = n8008 ^ n122 ^ 1'b0 ;
  assign n10055 = n1701 & n10054 ;
  assign n10056 = n2165 & n8086 ;
  assign n10057 = n3047 ^ n998 ^ 1'b0 ;
  assign n10058 = n4313 & ~n10057 ;
  assign n10059 = ( n6456 & n6921 ) | ( n6456 & ~n10058 ) | ( n6921 & ~n10058 ) ;
  assign n10060 = n4708 & ~n9527 ;
  assign n10061 = n8433 ^ n3730 ^ 1'b0 ;
  assign n10062 = n10061 ^ n2269 ^ 1'b0 ;
  assign n10063 = ~n1753 & n10062 ;
  assign n10064 = ~n6595 & n9846 ;
  assign n10065 = n53 | n941 ;
  assign n10066 = n939 & ~n10065 ;
  assign n10067 = n2572 & n6016 ;
  assign n10068 = n3793 & ~n6707 ;
  assign n10069 = n10068 ^ n2294 ^ 1'b0 ;
  assign n10070 = n8075 & ~n10020 ;
  assign n10071 = n10070 ^ n9420 ^ 1'b0 ;
  assign n10072 = n4287 ^ n2261 ^ 1'b0 ;
  assign n10073 = n3477 & ~n10072 ;
  assign n10074 = n10073 ^ n3995 ^ 1'b0 ;
  assign n10075 = n10074 ^ n144 ^ 1'b0 ;
  assign n10076 = n7271 & ~n10075 ;
  assign n10077 = n1360 | n8407 ;
  assign n10078 = ~n1100 & n4569 ;
  assign n10079 = n3300 ^ n2279 ^ 1'b0 ;
  assign n10080 = ( ~n7497 & n8967 ) | ( ~n7497 & n10079 ) | ( n8967 & n10079 ) ;
  assign n10081 = n4441 ^ n1922 ^ 1'b0 ;
  assign n10082 = n9170 ^ n6503 ^ 1'b0 ;
  assign n10083 = n10081 | n10082 ;
  assign n10084 = n3721 | n4001 ;
  assign n10085 = n6709 & n10084 ;
  assign n10086 = n191 | n9601 ;
  assign n10087 = ~n567 & n1372 ;
  assign n10088 = n670 & ~n10087 ;
  assign n10089 = n10088 ^ n7848 ^ 1'b0 ;
  assign n10090 = n5270 & n9137 ;
  assign n10091 = ~n3552 & n10090 ;
  assign n10092 = n10091 ^ n7040 ^ 1'b0 ;
  assign n10094 = n4267 ^ n2619 ^ 1'b0 ;
  assign n10095 = n2571 & n10094 ;
  assign n10093 = ~n954 & n3414 ;
  assign n10096 = n10095 ^ n10093 ^ 1'b0 ;
  assign n10097 = n80 | n5033 ;
  assign n10098 = n10097 ^ n4093 ^ 1'b0 ;
  assign n10099 = n4784 | n10098 ;
  assign n10100 = n7654 ^ n659 ^ 1'b0 ;
  assign n10101 = n3694 | n5112 ;
  assign n10102 = n1918 & ~n10097 ;
  assign n10103 = n7954 & n10102 ;
  assign n10104 = n10103 ^ n1726 ^ 1'b0 ;
  assign n10105 = n3620 ^ n997 ^ 1'b0 ;
  assign n10106 = n10105 ^ n2076 ^ 1'b0 ;
  assign n10107 = n8917 ^ n510 ^ 1'b0 ;
  assign n10108 = n72 & n81 ;
  assign n10109 = ~n81 & n10108 ;
  assign n10110 = ~n841 & n10109 ;
  assign n10111 = n2601 | n10110 ;
  assign n10112 = n10107 | n10111 ;
  assign n10113 = n1677 & n9169 ;
  assign n10114 = n9408 ^ n8566 ^ 1'b0 ;
  assign n10115 = ~n4281 & n10114 ;
  assign n10116 = n4796 ^ n2058 ^ 1'b0 ;
  assign n10117 = n142 | n10116 ;
  assign n10118 = n9281 | n10117 ;
  assign n10119 = n155 & n1946 ;
  assign n10120 = n1157 & ~n4006 ;
  assign n10121 = n5394 & n10120 ;
  assign n10122 = n6229 & n10121 ;
  assign n10123 = n10122 ^ n6456 ^ 1'b0 ;
  assign n10124 = ~n83 & n6063 ;
  assign n10125 = n2567 & n6471 ;
  assign n10126 = n10124 & n10125 ;
  assign n10127 = n7691 ^ n5218 ^ 1'b0 ;
  assign n10128 = ~n7182 & n10127 ;
  assign n10129 = n6407 ^ n6207 ^ 1'b0 ;
  assign n10130 = n7380 | n10129 ;
  assign n10131 = ~n677 & n10130 ;
  assign n10132 = n9242 ^ n2771 ^ 1'b0 ;
  assign n10133 = n1127 & ~n10132 ;
  assign n10134 = ~n2917 & n6873 ;
  assign n10135 = n8132 ^ n79 ^ 1'b0 ;
  assign n10136 = n4348 & ~n10135 ;
  assign n10137 = ~n6862 & n10136 ;
  assign n10138 = n322 & n4742 ;
  assign n10139 = n3874 ^ n364 ^ 1'b0 ;
  assign n10140 = n10138 & ~n10139 ;
  assign n10141 = n3099 ^ n822 ^ 1'b0 ;
  assign n10142 = n1810 & n2658 ;
  assign n10143 = n10141 & n10142 ;
  assign n10144 = n10140 & ~n10143 ;
  assign n10145 = n3382 ^ n1075 ^ 1'b0 ;
  assign n10146 = n10145 ^ n4794 ^ 1'b0 ;
  assign n10147 = n9875 & n10146 ;
  assign n10148 = ~n6730 & n10147 ;
  assign n10149 = n6459 & n10148 ;
  assign n10150 = n121 & n4815 ;
  assign n10151 = n10150 ^ n5234 ^ 1'b0 ;
  assign n10152 = n4488 ^ n2150 ^ 1'b0 ;
  assign n10153 = n3516 & ~n10152 ;
  assign n10154 = n2109 & ~n10153 ;
  assign n10155 = n10154 ^ n3416 ^ 1'b0 ;
  assign n10156 = n9238 ^ n4580 ^ n3585 ;
  assign n10157 = ~n177 & n1768 ;
  assign n10158 = n9372 ^ n2257 ^ 1'b0 ;
  assign n10159 = n2567 & n10158 ;
  assign n10160 = n4342 | n5454 ;
  assign n10161 = n2948 | n10160 ;
  assign n10162 = n1255 & n10161 ;
  assign n10163 = n10162 ^ n148 ^ 1'b0 ;
  assign n10164 = n2910 & n4415 ;
  assign n10165 = n10164 ^ n7779 ^ 1'b0 ;
  assign n10166 = n9973 ^ n8210 ^ 1'b0 ;
  assign n10167 = n10166 ^ n7039 ^ n553 ;
  assign n10168 = n241 & n423 ;
  assign n10169 = n556 ^ n23 ^ 1'b0 ;
  assign n10170 = n8283 & n10169 ;
  assign n10171 = n10170 ^ n7666 ^ 1'b0 ;
  assign n10172 = n654 & n7011 ;
  assign n10173 = n9495 & ~n10172 ;
  assign n10174 = n10173 ^ n4052 ^ 1'b0 ;
  assign n10175 = n1316 & n10174 ;
  assign n10176 = n1048 & ~n2282 ;
  assign n10177 = ~n685 & n10176 ;
  assign n10178 = n7064 & ~n9417 ;
  assign n10179 = n80 | n458 ;
  assign n10180 = n1396 & ~n10179 ;
  assign n10181 = n1205 ^ n1083 ^ 1'b0 ;
  assign n10182 = n4498 & ~n10181 ;
  assign n10183 = n3282 ^ n300 ^ 1'b0 ;
  assign n10184 = n749 & ~n10183 ;
  assign n10185 = n1852 ^ n1285 ^ 1'b0 ;
  assign n10186 = ~n1352 & n10185 ;
  assign n10187 = n10186 ^ n1388 ^ 1'b0 ;
  assign n10188 = n10184 & ~n10187 ;
  assign n10189 = n2180 ^ n883 ^ 1'b0 ;
  assign n10190 = n3203 | n10189 ;
  assign n10191 = n2297 | n9876 ;
  assign n10192 = ~n10190 & n10191 ;
  assign n10193 = n7231 & n10095 ;
  assign n10194 = ( n493 & ~n1999 ) | ( n493 & n2261 ) | ( ~n1999 & n2261 ) ;
  assign n10195 = ~n3483 & n10194 ;
  assign n10196 = n1595 ^ n1511 ^ 1'b0 ;
  assign n10197 = n2463 & n10196 ;
  assign n10198 = n8065 & ~n10197 ;
  assign n10199 = n10198 ^ n3856 ^ 1'b0 ;
  assign n10200 = n6008 & n10199 ;
  assign n10201 = n153 & ~n10072 ;
  assign n10202 = n1070 & n1602 ;
  assign n10204 = n1567 | n6698 ;
  assign n10203 = n7258 ^ n945 ^ 1'b0 ;
  assign n10205 = n10204 ^ n10203 ^ 1'b0 ;
  assign n10206 = n539 | n10205 ;
  assign n10207 = n2665 ^ n1258 ^ 1'b0 ;
  assign n10208 = n46 | n10207 ;
  assign n10209 = n7371 ^ n3143 ^ n2096 ;
  assign n10210 = n7112 & n10209 ;
  assign n10211 = n1084 & ~n5394 ;
  assign n10212 = n10211 ^ n3240 ^ 1'b0 ;
  assign n10213 = n208 & n321 ;
  assign n10214 = n10213 ^ n6102 ^ 1'b0 ;
  assign n10215 = n5103 & ~n10214 ;
  assign n10216 = ( n1041 & n2652 ) | ( n1041 & ~n10215 ) | ( n2652 & ~n10215 ) ;
  assign n10217 = n1354 | n3589 ;
  assign n10218 = n7145 & n10217 ;
  assign n10219 = n10218 ^ n241 ^ 1'b0 ;
  assign n10220 = n10219 ^ n6538 ^ 1'b0 ;
  assign n10221 = n8395 | n10220 ;
  assign n10222 = n6711 & ~n10221 ;
  assign n10223 = ~n9235 & n10222 ;
  assign n10224 = n1934 & n5554 ;
  assign n10225 = n9245 ^ n1546 ^ 1'b0 ;
  assign n10226 = n8112 & ~n10225 ;
  assign n10227 = n1743 | n4644 ;
  assign n10228 = n62 & ~n10227 ;
  assign n10229 = n10228 ^ n2768 ^ 1'b0 ;
  assign n10230 = n3077 ^ n2426 ^ 1'b0 ;
  assign n10231 = n4848 | n10230 ;
  assign n10232 = n2589 & ~n10231 ;
  assign n10233 = n10232 ^ n1138 ^ 1'b0 ;
  assign n10234 = n1445 & ~n4081 ;
  assign n10235 = n9417 | n10234 ;
  assign n10236 = n6084 & ~n10235 ;
  assign n10237 = ~n2120 & n10236 ;
  assign n10238 = n2222 ^ n671 ^ 1'b0 ;
  assign n10239 = ~n10237 & n10238 ;
  assign n10240 = ~n1310 & n10239 ;
  assign n10241 = n10240 ^ n6721 ^ 1'b0 ;
  assign n10245 = n3013 | n4034 ;
  assign n10242 = n2150 ^ n749 ^ 1'b0 ;
  assign n10243 = ~n7614 & n10242 ;
  assign n10244 = ~n876 & n10243 ;
  assign n10246 = n10245 ^ n10244 ^ 1'b0 ;
  assign n10247 = n646 & n1898 ;
  assign n10248 = n7634 ^ n6603 ^ 1'b0 ;
  assign n10249 = n2210 & ~n10248 ;
  assign n10250 = n5380 & n10249 ;
  assign n10251 = n10250 ^ n216 ^ 1'b0 ;
  assign n10252 = ~n294 & n6401 ;
  assign n10253 = ( n713 & n1851 ) | ( n713 & n1937 ) | ( n1851 & n1937 ) ;
  assign n10254 = n2958 ^ n2155 ^ 1'b0 ;
  assign n10255 = n2305 | n10254 ;
  assign n10256 = n5733 ^ n2848 ^ 1'b0 ;
  assign n10257 = n10255 | n10256 ;
  assign n10258 = n4117 ^ n2491 ^ 1'b0 ;
  assign n10259 = ~n10257 & n10258 ;
  assign n10260 = n8395 & n10259 ;
  assign n10261 = n8804 ^ n1622 ^ 1'b0 ;
  assign n10262 = n1063 | n10261 ;
  assign n10263 = n423 & ~n10262 ;
  assign n10264 = ~n7144 & n10263 ;
  assign n10265 = n7683 ^ n615 ^ 1'b0 ;
  assign n10266 = n113 & ~n10265 ;
  assign n10267 = ~n405 & n1656 ;
  assign n10268 = n4000 & n4399 ;
  assign n10269 = n8797 ^ n8410 ^ 1'b0 ;
  assign n10270 = n675 ^ n400 ^ 1'b0 ;
  assign n10271 = n36 & ~n10270 ;
  assign n10272 = ~n995 & n10271 ;
  assign n10273 = ~n3871 & n10272 ;
  assign n10274 = n10273 ^ n2606 ^ n663 ;
  assign n10275 = n7301 & ~n10274 ;
  assign n10276 = n457 & ~n2150 ;
  assign n10277 = ~n4448 & n10276 ;
  assign n10278 = n159 & ~n10277 ;
  assign n10279 = ~n555 & n10278 ;
  assign n10280 = n10275 & n10279 ;
  assign n10281 = n2438 ^ n1465 ^ 1'b0 ;
  assign n10282 = n9307 & ~n10281 ;
  assign n10283 = n278 & ~n5190 ;
  assign n10284 = n10283 ^ n823 ^ 1'b0 ;
  assign n10285 = n1268 & ~n3258 ;
  assign n10286 = ~n5696 & n9585 ;
  assign n10288 = ~n200 & n2049 ;
  assign n10287 = n2295 & ~n4616 ;
  assign n10289 = n10288 ^ n10287 ^ 1'b0 ;
  assign n10290 = n1997 ^ n274 ^ 1'b0 ;
  assign n10291 = n1345 & n10290 ;
  assign n10292 = n7555 | n10291 ;
  assign n10293 = n212 | n906 ;
  assign n10294 = ~n236 & n10293 ;
  assign n10295 = n8560 ^ n128 ^ 1'b0 ;
  assign n10296 = ~n10294 & n10295 ;
  assign n10297 = n3061 | n6571 ;
  assign n10298 = n417 | n10297 ;
  assign n10299 = x3 & n121 ;
  assign n10300 = ~n121 & n10299 ;
  assign n10301 = n27 & n10300 ;
  assign n10302 = n10301 ^ n1802 ^ 1'b0 ;
  assign n10303 = n1606 & ~n2102 ;
  assign n10304 = n4480 & ~n10303 ;
  assign n10305 = n10303 & n10304 ;
  assign n10306 = n10302 & ~n10305 ;
  assign n10307 = n9104 & n10306 ;
  assign n10308 = n3028 ^ n520 ^ 1'b0 ;
  assign n10309 = n8309 & ~n10308 ;
  assign n10310 = n10309 ^ n659 ^ 1'b0 ;
  assign n10311 = n5828 | n7381 ;
  assign n10312 = n8804 | n10311 ;
  assign n10313 = n456 ^ n308 ^ 1'b0 ;
  assign n10314 = ~n393 & n4022 ;
  assign n10315 = n10314 ^ n566 ^ 1'b0 ;
  assign n10316 = n4347 ^ n851 ^ 1'b0 ;
  assign n10317 = n10315 | n10316 ;
  assign n10318 = ~n517 & n10317 ;
  assign n10319 = n3685 & ~n4986 ;
  assign n10320 = ~n6322 & n10319 ;
  assign n10321 = n6704 & n7764 ;
  assign n10322 = n5570 ^ n3154 ^ 1'b0 ;
  assign n10323 = n5234 ^ n2535 ^ 1'b0 ;
  assign n10324 = n5412 & n5420 ;
  assign n10325 = n472 & n10324 ;
  assign n10326 = n1513 | n1632 ;
  assign n10327 = n10326 ^ n5646 ^ 1'b0 ;
  assign n10328 = n10327 ^ n10060 ^ 1'b0 ;
  assign n10329 = n654 | n7872 ;
  assign n10330 = n8276 ^ n6989 ^ 1'b0 ;
  assign n10331 = ~n2409 & n4066 ;
  assign n10332 = n10331 ^ n1957 ^ 1'b0 ;
  assign n10333 = n10332 ^ n7867 ^ 1'b0 ;
  assign n10334 = n9492 ^ n4022 ^ 1'b0 ;
  assign n10335 = n9014 | n10334 ;
  assign n10336 = n1924 & ~n8272 ;
  assign n10337 = ~n1252 & n10336 ;
  assign n10338 = n10337 ^ n4551 ^ 1'b0 ;
  assign n10339 = n1686 & ~n9979 ;
  assign n10340 = n2980 & n4770 ;
  assign n10341 = n2939 | n8329 ;
  assign n10342 = n10340 | n10341 ;
  assign n10343 = n179 | n10342 ;
  assign n10344 = n1020 & n3047 ;
  assign n10345 = n10344 ^ n5837 ^ 1'b0 ;
  assign n10346 = ~n666 & n4585 ;
  assign n10347 = ~n32 & n10346 ;
  assign n10348 = n43 | n10347 ;
  assign n10349 = n3124 ^ n62 ^ 1'b0 ;
  assign n10350 = n1367 & ~n4341 ;
  assign n10351 = n5143 ^ n2104 ^ 1'b0 ;
  assign n10352 = n10350 & ~n10351 ;
  assign n10353 = n302 | n1564 ;
  assign n10354 = n5443 & n10353 ;
  assign n10355 = ~n5080 & n10354 ;
  assign n10356 = n4432 & ~n9897 ;
  assign n10357 = n4595 | n9220 ;
  assign n10358 = n9027 ^ n1733 ^ 1'b0 ;
  assign n10359 = ( ~n1653 & n3742 ) | ( ~n1653 & n5468 ) | ( n3742 & n5468 ) ;
  assign n10360 = ( n8976 & ~n10358 ) | ( n8976 & n10359 ) | ( ~n10358 & n10359 ) ;
  assign n10361 = n5891 ^ n3697 ^ 1'b0 ;
  assign n10362 = n6860 | n7895 ;
  assign n10363 = n6540 & ~n10362 ;
  assign n10364 = ~n5201 & n6938 ;
  assign n10365 = n1957 & n10364 ;
  assign n10366 = ~n4584 & n10365 ;
  assign n10367 = ~n10363 & n10366 ;
  assign n10368 = ~n576 & n9695 ;
  assign n10369 = n10368 ^ n3929 ^ 1'b0 ;
  assign n10370 = ~n5108 & n9237 ;
  assign n10371 = n3817 & ~n8784 ;
  assign n10372 = n5823 & n10371 ;
  assign n10373 = ~x0 & n4916 ;
  assign n10374 = ~n354 & n10373 ;
  assign n10376 = n614 ^ n359 ^ 1'b0 ;
  assign n10377 = n1155 & ~n10376 ;
  assign n10375 = n3125 ^ n1316 ^ 1'b0 ;
  assign n10378 = n10377 ^ n10375 ^ 1'b0 ;
  assign n10379 = ~n2324 & n6133 ;
  assign n10380 = n52 & n1856 ;
  assign n10381 = n10380 ^ n6210 ^ 1'b0 ;
  assign n10382 = n3744 | n10381 ;
  assign n10383 = n653 & ~n2496 ;
  assign n10384 = n532 | n10383 ;
  assign n10385 = n2136 & n3374 ;
  assign n10386 = n8705 & n10385 ;
  assign n10387 = n9752 & n10386 ;
  assign n10388 = n1388 ^ n954 ^ 1'b0 ;
  assign n10389 = n3663 | n10388 ;
  assign n10390 = n10389 ^ n353 ^ 1'b0 ;
  assign n10391 = n799 | n6818 ;
  assign n10392 = n1044 ^ n323 ^ 1'b0 ;
  assign n10393 = n6154 | n10392 ;
  assign n10398 = n6333 ^ n1816 ^ 1'b0 ;
  assign n10394 = ~n4060 & n4746 ;
  assign n10395 = n3068 & ~n5933 ;
  assign n10396 = n10395 ^ n8142 ^ n6506 ;
  assign n10397 = n10394 & ~n10396 ;
  assign n10399 = n10398 ^ n10397 ^ 1'b0 ;
  assign n10400 = n928 & n9381 ;
  assign n10401 = n10400 ^ n461 ^ 1'b0 ;
  assign n10402 = ~n588 & n6254 ;
  assign n10403 = n10402 ^ n6420 ^ 1'b0 ;
  assign n10404 = n8804 & n10403 ;
  assign n10405 = ~n4952 & n10404 ;
  assign n10407 = n1584 | n7221 ;
  assign n10408 = n2261 & ~n10407 ;
  assign n10409 = n10408 ^ n1513 ^ 1'b0 ;
  assign n10406 = n1598 & ~n4475 ;
  assign n10410 = n10409 ^ n10406 ^ 1'b0 ;
  assign n10411 = ~n1538 & n10025 ;
  assign n10412 = n10411 ^ n4337 ^ 1'b0 ;
  assign n10413 = n1990 | n10412 ;
  assign n10414 = n10410 & ~n10413 ;
  assign n10415 = n639 | n4379 ;
  assign n10416 = n4813 ^ n1662 ^ 1'b0 ;
  assign n10417 = n6242 & n10416 ;
  assign n10418 = n10417 ^ n246 ^ 1'b0 ;
  assign n10419 = n10415 & ~n10418 ;
  assign n10420 = n185 | n4791 ;
  assign n10421 = n310 & n2316 ;
  assign n10422 = n1891 & ~n10421 ;
  assign n10423 = n6468 ^ n5152 ^ 1'b0 ;
  assign n10424 = ~n144 & n5617 ;
  assign n10425 = n1362 & ~n4428 ;
  assign n10426 = ( n1608 & ~n4446 ) | ( n1608 & n10425 ) | ( ~n4446 & n10425 ) ;
  assign n10427 = n4449 | n5146 ;
  assign n10428 = n4697 & ~n10427 ;
  assign n10429 = n5068 ^ n1233 ^ 1'b0 ;
  assign n10430 = ( n4493 & n4619 ) | ( n4493 & ~n10429 ) | ( n4619 & ~n10429 ) ;
  assign n10431 = n128 | n2573 ;
  assign n10432 = n6875 | n10431 ;
  assign n10433 = n2297 ^ n1748 ^ 1'b0 ;
  assign n10434 = ~n4031 & n10433 ;
  assign n10435 = n5811 & ~n6129 ;
  assign n10436 = n10435 ^ n2607 ^ 1'b0 ;
  assign n10437 = n5764 & ~n10436 ;
  assign n10438 = ~n294 & n10437 ;
  assign n10439 = n10438 ^ n2289 ^ 1'b0 ;
  assign n10440 = n1497 | n3186 ;
  assign n10441 = n592 & ~n10440 ;
  assign n10442 = n10441 ^ n1937 ^ 1'b0 ;
  assign n10443 = n10442 ^ n10437 ^ n3433 ;
  assign n10444 = n10443 ^ n1379 ^ 1'b0 ;
  assign n10445 = n506 & n748 ;
  assign n10446 = ~n16 & n10445 ;
  assign n10447 = ~n5955 & n10446 ;
  assign n10448 = ~n1881 & n10447 ;
  assign n10449 = n142 & ~n338 ;
  assign n10457 = n2414 ^ n1516 ^ 1'b0 ;
  assign n10450 = n1447 & ~n1631 ;
  assign n10451 = n2194 & n10450 ;
  assign n10452 = n929 ^ n310 ^ 1'b0 ;
  assign n10453 = n4028 | n10452 ;
  assign n10454 = n10451 & ~n10453 ;
  assign n10455 = n2849 & ~n9819 ;
  assign n10456 = n10454 & n10455 ;
  assign n10458 = n10457 ^ n10456 ^ 1'b0 ;
  assign n10459 = n510 & n10458 ;
  assign n10460 = n5542 ^ n1964 ^ 1'b0 ;
  assign n10461 = n281 & n10460 ;
  assign n10462 = n2524 & n10461 ;
  assign n10463 = n5979 & n10462 ;
  assign n10470 = ~n1330 & n3009 ;
  assign n10464 = n2594 | n5263 ;
  assign n10465 = n1081 & ~n2933 ;
  assign n10466 = n10465 ^ n6926 ^ 1'b0 ;
  assign n10467 = ~n10464 & n10466 ;
  assign n10468 = n1928 & n10467 ;
  assign n10469 = ~n8917 & n10468 ;
  assign n10471 = n10470 ^ n10469 ^ 1'b0 ;
  assign n10472 = n10371 & n10471 ;
  assign n10474 = n1235 | n4830 ;
  assign n10475 = n10474 ^ n866 ^ 1'b0 ;
  assign n10473 = ~n9161 & n9563 ;
  assign n10476 = n10475 ^ n10473 ^ 1'b0 ;
  assign n10477 = n3986 | n8392 ;
  assign n10478 = n10477 ^ n9412 ^ 1'b0 ;
  assign n10479 = n10476 | n10478 ;
  assign n10480 = n8279 ^ n3065 ^ 1'b0 ;
  assign n10481 = ~n1318 & n2282 ;
  assign n10482 = n10481 ^ n1933 ^ 1'b0 ;
  assign n10483 = n2022 & ~n7104 ;
  assign n10484 = ~n4329 & n10483 ;
  assign n10485 = n2380 ^ n2216 ^ 1'b0 ;
  assign n10486 = ~n10484 & n10485 ;
  assign n10487 = ~n2017 & n10486 ;
  assign n10488 = n5438 ^ n3693 ^ 1'b0 ;
  assign n10489 = n10392 & n10488 ;
  assign n10490 = n3338 ^ n2059 ^ 1'b0 ;
  assign n10491 = n10235 ^ n5182 ^ 1'b0 ;
  assign n10492 = n1192 & n10491 ;
  assign n10493 = n763 & ~n5123 ;
  assign n10494 = n7431 ^ n192 ^ 1'b0 ;
  assign n10495 = n1174 & n10494 ;
  assign n10496 = n2941 | n10381 ;
  assign n10497 = n10496 ^ n8946 ^ 1'b0 ;
  assign n10498 = n478 | n7853 ;
  assign n10499 = n10497 & ~n10498 ;
  assign n10500 = n9617 ^ n2747 ^ 1'b0 ;
  assign n10501 = ~n1893 & n2523 ;
  assign n10502 = n5362 & n10501 ;
  assign n10503 = n163 ^ n82 ^ 1'b0 ;
  assign n10504 = n227 | n10503 ;
  assign n10505 = n10504 ^ n3399 ^ n2236 ;
  assign n10506 = n10505 ^ n2426 ^ 1'b0 ;
  assign n10507 = n5763 & ~n10506 ;
  assign n10508 = ~n6258 & n8242 ;
  assign n10509 = n666 & n7923 ;
  assign n10510 = n3885 & ~n5134 ;
  assign n10511 = n9763 ^ n4424 ^ 1'b0 ;
  assign n10512 = ( n3886 & ~n10510 ) | ( n3886 & n10511 ) | ( ~n10510 & n10511 ) ;
  assign n10513 = n385 & ~n4315 ;
  assign n10514 = n10513 ^ n10330 ^ 1'b0 ;
  assign n10515 = n840 | n1690 ;
  assign n10516 = n1283 & ~n10515 ;
  assign n10517 = n10516 ^ n5845 ^ 1'b0 ;
  assign n10518 = n16 & ~n3622 ;
  assign n10519 = n10518 ^ n2912 ^ 1'b0 ;
  assign n10521 = n1177 | n2041 ;
  assign n10520 = n10036 ^ n286 ^ 1'b0 ;
  assign n10522 = n10521 ^ n10520 ^ 1'b0 ;
  assign n10523 = ~n769 & n10522 ;
  assign n10524 = n3816 & ~n9251 ;
  assign n10525 = n5574 ^ n56 ^ 1'b0 ;
  assign n10526 = ~n6976 & n10525 ;
  assign n10527 = n10526 ^ n5632 ^ 1'b0 ;
  assign n10528 = n3808 ^ n363 ^ 1'b0 ;
  assign n10529 = n1304 | n10528 ;
  assign n10530 = ( n532 & n10527 ) | ( n532 & n10529 ) | ( n10527 & n10529 ) ;
  assign n10531 = n741 & n10215 ;
  assign n10532 = n8510 ^ n5668 ^ 1'b0 ;
  assign n10533 = n9881 ^ n4116 ^ 1'b0 ;
  assign n10534 = n2969 & n4267 ;
  assign n10535 = n10268 ^ n4774 ^ 1'b0 ;
  assign n10536 = n456 | n6463 ;
  assign n10537 = n1057 & n4048 ;
  assign n10538 = n1052 & ~n3176 ;
  assign n10539 = ~n279 & n9607 ;
  assign n10540 = n4815 & n7596 ;
  assign n10541 = n10540 ^ n748 ^ 1'b0 ;
  assign n10542 = n938 & n1165 ;
  assign n10543 = n10542 ^ n4365 ^ 1'b0 ;
  assign n10544 = n1057 & ~n6866 ;
  assign n10545 = ~n7330 & n10544 ;
  assign n10546 = ~n542 & n10545 ;
  assign n10547 = ~n802 & n5334 ;
  assign n10548 = n433 ^ n55 ^ 1'b0 ;
  assign n10549 = n10548 ^ n3793 ^ 1'b0 ;
  assign n10550 = ~n2254 & n10549 ;
  assign n10551 = n738 & n10550 ;
  assign n10552 = n8664 & n10551 ;
  assign n10553 = n6871 & n10552 ;
  assign n10554 = n1691 ^ n782 ^ 1'b0 ;
  assign n10556 = n7377 ^ n2043 ^ 1'b0 ;
  assign n10557 = n252 | n10556 ;
  assign n10558 = n1425 & ~n10557 ;
  assign n10559 = n10558 ^ n4267 ^ 1'b0 ;
  assign n10555 = ~n2785 & n6896 ;
  assign n10560 = n10559 ^ n10555 ^ 1'b0 ;
  assign n10561 = n259 ^ n139 ^ 1'b0 ;
  assign n10562 = n5207 | n10561 ;
  assign n10563 = n10561 & ~n10562 ;
  assign n10564 = n7808 & ~n10563 ;
  assign n10565 = n10564 ^ n8991 ^ 1'b0 ;
  assign n10566 = n8166 ^ n2939 ^ 1'b0 ;
  assign n10567 = n1057 & n10566 ;
  assign n10568 = n10567 ^ n7424 ^ 1'b0 ;
  assign n10569 = ~n1016 & n10568 ;
  assign n10570 = n1898 & ~n9925 ;
  assign n10571 = n6890 & n10570 ;
  assign n10572 = n9102 & n10571 ;
  assign n10573 = n319 & n3519 ;
  assign n10574 = n10573 ^ n2558 ^ 1'b0 ;
  assign n10575 = n10574 ^ n1770 ^ 1'b0 ;
  assign n10576 = n3338 & ~n3401 ;
  assign n10577 = n811 & ~n5892 ;
  assign n10578 = ~n1975 & n10577 ;
  assign n10579 = n7399 | n10578 ;
  assign n10580 = n2163 ^ n462 ^ 1'b0 ;
  assign n10582 = ~n489 & n1286 ;
  assign n10581 = n9980 ^ n4903 ^ 1'b0 ;
  assign n10583 = n10582 ^ n10581 ^ 1'b0 ;
  assign n10584 = n5158 ^ n527 ^ 1'b0 ;
  assign n10585 = ~n1608 & n1731 ;
  assign n10586 = n10585 ^ n6067 ^ 1'b0 ;
  assign n10587 = n1531 & n2941 ;
  assign n10588 = n4169 & n10587 ;
  assign n10589 = n1430 ^ n456 ^ 1'b0 ;
  assign n10590 = n10588 & ~n10589 ;
  assign n10591 = n497 | n7236 ;
  assign n10592 = n8993 ^ n6755 ^ n3539 ;
  assign n10593 = n8566 ^ n7709 ^ 1'b0 ;
  assign n10596 = n1038 ^ n274 ^ 1'b0 ;
  assign n10595 = ~n3078 & n7064 ;
  assign n10597 = n10596 ^ n10595 ^ 1'b0 ;
  assign n10594 = n259 | n1081 ;
  assign n10598 = n10597 ^ n10594 ^ n2893 ;
  assign n10599 = n4432 & ~n7649 ;
  assign n10600 = n1049 & n8041 ;
  assign n10601 = n10600 ^ n3792 ^ 1'b0 ;
  assign n10602 = n8975 & n10601 ;
  assign n10603 = n10602 ^ n7707 ^ 1'b0 ;
  assign n10604 = n2731 ^ n2432 ^ 1'b0 ;
  assign n10605 = ~n2742 & n3283 ;
  assign n10606 = n8789 ^ n6782 ^ 1'b0 ;
  assign n10607 = n9823 & n10606 ;
  assign n10608 = ~n2752 & n7457 ;
  assign n10609 = n2677 ^ n1768 ^ 1'b0 ;
  assign n10610 = n1826 & n10609 ;
  assign n10611 = ~n1810 & n1825 ;
  assign n10612 = n4770 | n10611 ;
  assign n10613 = ~n387 & n9251 ;
  assign n10614 = n1191 | n5270 ;
  assign n10615 = n10614 ^ n3637 ^ 1'b0 ;
  assign n10616 = n10615 ^ n2164 ^ 1'b0 ;
  assign n10617 = n10613 & ~n10616 ;
  assign n10618 = n119 & n2493 ;
  assign n10619 = n1688 | n10618 ;
  assign n10620 = n954 ^ n382 ^ 1'b0 ;
  assign n10621 = ~n7043 & n10620 ;
  assign n10622 = n10621 ^ n2200 ^ 1'b0 ;
  assign n10623 = n3816 & ~n6541 ;
  assign n10624 = n10622 & n10623 ;
  assign n10625 = n832 & ~n5856 ;
  assign n10626 = n6746 & n10625 ;
  assign n10627 = n8961 & n10626 ;
  assign n10628 = ~n520 & n1316 ;
  assign n10629 = n10628 ^ n1491 ^ 1'b0 ;
  assign n10630 = ~n10627 & n10629 ;
  assign n10631 = n2453 | n7865 ;
  assign n10632 = ~n234 & n1141 ;
  assign n10633 = n258 | n4532 ;
  assign n10634 = n384 & n7289 ;
  assign n10635 = n2876 ^ n1896 ^ 1'b0 ;
  assign n10636 = ~n1482 & n10635 ;
  assign n10637 = n8411 | n10636 ;
  assign n10638 = n616 ^ n372 ^ 1'b0 ;
  assign n10639 = n8465 ^ n1011 ^ 1'b0 ;
  assign n10640 = n279 & n2119 ;
  assign n10641 = n10639 & n10640 ;
  assign n10642 = n10641 ^ n9939 ^ 1'b0 ;
  assign n10643 = n10638 | n10642 ;
  assign n10644 = n5706 & n8552 ;
  assign n10645 = n1304 ^ n713 ^ 1'b0 ;
  assign n10646 = n1986 & n6676 ;
  assign n10647 = n4468 ^ n2885 ^ 1'b0 ;
  assign n10648 = n10647 ^ n4241 ^ n89 ;
  assign n10649 = n448 ^ n85 ^ 1'b0 ;
  assign n10650 = n10649 ^ n596 ^ 1'b0 ;
  assign n10651 = n2543 & n5872 ;
  assign n10652 = n10651 ^ n2733 ^ 1'b0 ;
  assign n10653 = n10650 | n10652 ;
  assign n10654 = n4104 ^ n3940 ^ 1'b0 ;
  assign n10655 = n3025 | n10654 ;
  assign n10656 = n10655 ^ n9289 ^ n4449 ;
  assign n10657 = n6142 ^ n1900 ^ 1'b0 ;
  assign n10658 = n9629 ^ n1048 ^ 1'b0 ;
  assign n10659 = n10658 ^ n9850 ^ 1'b0 ;
  assign n10660 = ~n1724 & n3137 ;
  assign n10661 = n10660 ^ n3449 ^ 1'b0 ;
  assign n10662 = ~n5900 & n6746 ;
  assign n10663 = n2109 ^ x5 ^ 1'b0 ;
  assign n10664 = n10663 ^ n2694 ^ 1'b0 ;
  assign n10665 = n5964 & ~n10664 ;
  assign n10666 = ~n10201 & n10665 ;
  assign n10667 = n208 & n10292 ;
  assign n10668 = n10666 & n10667 ;
  assign n10669 = n310 & n8155 ;
  assign n10670 = ~n7544 & n10669 ;
  assign n10671 = n9478 ^ n4458 ^ 1'b0 ;
  assign n10672 = n3637 & n10671 ;
  assign n10673 = n3512 & n9980 ;
  assign n10674 = n1597 | n10234 ;
  assign n10675 = n8166 ^ n6426 ^ 1'b0 ;
  assign n10677 = ( n928 & n3513 ) | ( n928 & ~n3980 ) | ( n3513 & ~n3980 ) ;
  assign n10676 = ~n5393 & n5635 ;
  assign n10678 = n10677 ^ n10676 ^ 1'b0 ;
  assign n10679 = n3315 | n5686 ;
  assign n10680 = n10679 ^ n4394 ^ 1'b0 ;
  assign n10681 = n10680 ^ n5280 ^ 1'b0 ;
  assign n10682 = ~n10678 & n10681 ;
  assign n10683 = ~n286 & n300 ;
  assign n10684 = n10683 ^ n9387 ^ 1'b0 ;
  assign n10685 = n395 & n10684 ;
  assign n10686 = ( ~n678 & n4581 ) | ( ~n678 & n10685 ) | ( n4581 & n10685 ) ;
  assign n10687 = ~n2483 & n5681 ;
  assign n10688 = n8210 | n10687 ;
  assign n10689 = n10688 ^ n1178 ^ 1'b0 ;
  assign n10690 = n3008 ^ n268 ^ 1'b0 ;
  assign n10691 = n10690 ^ n5469 ^ 1'b0 ;
  assign n10692 = n10691 ^ n3670 ^ 1'b0 ;
  assign n10693 = n1154 | n3293 ;
  assign n10694 = n3293 & ~n10693 ;
  assign n10695 = n534 | n2998 ;
  assign n10696 = n2998 & ~n10695 ;
  assign n10697 = ~n3523 & n8149 ;
  assign n10698 = n3523 & n10697 ;
  assign n10699 = n5393 & ~n10698 ;
  assign n10700 = ~n5393 & n10699 ;
  assign n10701 = ~n929 & n10700 ;
  assign n10702 = n10701 ^ n10509 ^ 1'b0 ;
  assign n10703 = n10696 | n10702 ;
  assign n10704 = n10694 & ~n10703 ;
  assign n10705 = n1904 | n6072 ;
  assign n10706 = n7901 | n10705 ;
  assign n10707 = n2061 | n4361 ;
  assign n10708 = n8216 ^ n3194 ^ 1'b0 ;
  assign n10709 = n10020 ^ n3243 ^ 1'b0 ;
  assign n10710 = x3 & ~n290 ;
  assign n10711 = n290 & n10710 ;
  assign n10712 = n4487 & ~n10711 ;
  assign n10713 = ~n4487 & n10712 ;
  assign n10714 = ~n1191 & n1300 ;
  assign n10715 = n10713 & n10714 ;
  assign n10716 = ~n8321 & n10715 ;
  assign n10717 = n10716 ^ n1423 ^ 1'b0 ;
  assign n10718 = n9626 ^ n779 ^ 1'b0 ;
  assign n10719 = n1304 & ~n7579 ;
  assign n10720 = n1329 ^ n88 ^ 1'b0 ;
  assign n10721 = ~n6740 & n10720 ;
  assign n10722 = n9187 & n10721 ;
  assign n10723 = ~n6237 & n10722 ;
  assign n10724 = n2490 | n3182 ;
  assign n10725 = n10724 ^ n3603 ^ 1'b0 ;
  assign n10726 = n10725 ^ n365 ^ 1'b0 ;
  assign n10727 = n10726 ^ n10447 ^ 1'b0 ;
  assign n10728 = n1597 & n5053 ;
  assign n10729 = n6383 & n6673 ;
  assign n10732 = n4120 | n8784 ;
  assign n10733 = n10732 ^ n1979 ^ 1'b0 ;
  assign n10734 = n2571 & ~n10733 ;
  assign n10735 = ( n2942 & n3774 ) | ( n2942 & ~n10734 ) | ( n3774 & ~n10734 ) ;
  assign n10730 = n10470 ^ n479 ^ 1'b0 ;
  assign n10731 = n5292 & n10730 ;
  assign n10736 = n10735 ^ n10731 ^ 1'b0 ;
  assign n10737 = n3717 & ~n8309 ;
  assign n10738 = ~n3554 & n10737 ;
  assign n10739 = n10738 ^ x0 ^ 1'b0 ;
  assign n10740 = n4152 & n7960 ;
  assign n10741 = n945 | n9707 ;
  assign n10742 = n10032 ^ n2867 ^ 1'b0 ;
  assign n10743 = n2103 & ~n10742 ;
  assign n10744 = n348 & ~n880 ;
  assign n10745 = n10744 ^ n3477 ^ 1'b0 ;
  assign n10746 = n3706 & n10745 ;
  assign n10747 = n1948 | n10746 ;
  assign n10748 = n1676 ^ n19 ^ 1'b0 ;
  assign n10749 = n1080 & ~n10748 ;
  assign n10750 = ~n190 & n10749 ;
  assign n10751 = n10750 ^ n3718 ^ 1'b0 ;
  assign n10752 = n5362 ^ n3839 ^ 1'b0 ;
  assign n10753 = n9244 ^ n4361 ^ n86 ;
  assign n10754 = n10753 ^ n3411 ^ 1'b0 ;
  assign n10755 = n7207 & n10754 ;
  assign n10756 = n3214 ^ n3192 ^ 1'b0 ;
  assign n10757 = n2586 & n10756 ;
  assign n10758 = n10757 ^ n2872 ^ 1'b0 ;
  assign n10760 = ~n212 & n2594 ;
  assign n10759 = n2196 | n9166 ;
  assign n10761 = n10760 ^ n10759 ^ 1'b0 ;
  assign n10762 = n1828 & n9952 ;
  assign n10763 = n938 ^ n813 ^ 1'b0 ;
  assign n10764 = n4399 & n8467 ;
  assign n10765 = ~n6067 & n10764 ;
  assign n10766 = n9443 ^ n3665 ^ 1'b0 ;
  assign n10767 = n5889 ^ n1095 ^ 1'b0 ;
  assign n10768 = n2481 & n5556 ;
  assign n10769 = n204 & n10768 ;
  assign n10770 = n3279 | n8021 ;
  assign n10771 = n7138 ^ n5235 ^ 1'b0 ;
  assign n10772 = ~n7217 & n10771 ;
  assign n10773 = n1976 & ~n6433 ;
  assign n10774 = ~n181 & n10773 ;
  assign n10775 = ~x1 & n4794 ;
  assign n10776 = n10775 ^ n9319 ^ 1'b0 ;
  assign n10777 = n2031 | n4715 ;
  assign n10778 = n9067 & ~n10777 ;
  assign n10779 = n5503 & n9006 ;
  assign n10780 = n10779 ^ n4559 ^ 1'b0 ;
  assign n10781 = n5437 ^ n2348 ^ 1'b0 ;
  assign n10782 = n1023 & ~n4609 ;
  assign n10784 = n3361 | n7374 ;
  assign n10783 = ~n2075 & n5424 ;
  assign n10785 = n10784 ^ n10783 ^ 1'b0 ;
  assign n10786 = n4139 | n4603 ;
  assign n10787 = n4544 | n10786 ;
  assign n10788 = ~n2908 & n10787 ;
  assign n10791 = n700 | n2282 ;
  assign n10789 = n9120 ^ n2759 ^ 1'b0 ;
  assign n10790 = n10789 ^ n4227 ^ 1'b0 ;
  assign n10792 = n10791 ^ n10790 ^ 1'b0 ;
  assign n10793 = n849 & n10792 ;
  assign n10794 = n5111 | n8626 ;
  assign n10795 = n10793 & n10794 ;
  assign n10796 = n1377 & ~n2430 ;
  assign n10797 = n8265 ^ n4809 ^ 1'b0 ;
  assign n10798 = n10797 ^ n1406 ^ 1'b0 ;
  assign n10799 = n3566 & n7747 ;
  assign n10800 = n3335 & n3656 ;
  assign n10801 = n9521 & n10800 ;
  assign n10802 = n290 | n10801 ;
  assign n10803 = n10802 ^ n4033 ^ 1'b0 ;
  assign n10805 = ~n6567 & n7551 ;
  assign n10806 = ( n3542 & n9351 ) | ( n3542 & ~n10805 ) | ( n9351 & ~n10805 ) ;
  assign n10804 = n5963 & n9920 ;
  assign n10807 = n10806 ^ n10804 ^ 1'b0 ;
  assign n10808 = ~n2378 & n7268 ;
  assign n10809 = n906 | n9220 ;
  assign n10810 = ~n1183 & n4519 ;
  assign n10811 = n170 | n10810 ;
  assign n10812 = n8137 & ~n10811 ;
  assign n10813 = n2861 & ~n4807 ;
  assign n10814 = ~n10812 & n10813 ;
  assign n10815 = n6081 ^ n2107 ^ 1'b0 ;
  assign n10816 = n4526 ^ n3550 ^ 1'b0 ;
  assign n10817 = n3575 & n10816 ;
  assign n10818 = ~n10815 & n10817 ;
  assign n10819 = n2101 & ~n5722 ;
  assign n10820 = n4398 ^ n917 ^ 1'b0 ;
  assign n10821 = ~n10819 & n10820 ;
  assign n10822 = ~n865 & n10821 ;
  assign n10823 = ( n1246 & ~n2180 ) | ( n1246 & n7082 ) | ( ~n2180 & n7082 ) ;
  assign n10824 = ~n7021 & n8617 ;
  assign n10825 = n227 & n297 ;
  assign n10826 = n4689 ^ n2109 ^ 1'b0 ;
  assign n10827 = n7341 & n8570 ;
  assign n10828 = n364 | n709 ;
  assign n10829 = n10828 ^ n3340 ^ 1'b0 ;
  assign n10830 = n4761 ^ n3164 ^ 1'b0 ;
  assign n10831 = n3645 ^ n3519 ^ 1'b0 ;
  assign n10832 = ~n8918 & n10831 ;
  assign n10833 = n8632 & n10832 ;
  assign n10834 = n7492 ^ n1488 ^ 1'b0 ;
  assign n10835 = n8488 ^ n7032 ^ 1'b0 ;
  assign n10836 = n4739 | n10835 ;
  assign n10837 = n7011 ^ n3584 ^ 1'b0 ;
  assign n10839 = n4511 & ~n4514 ;
  assign n10840 = n10839 ^ n10377 ^ 1'b0 ;
  assign n10838 = ~n6081 & n6664 ;
  assign n10841 = n10840 ^ n10838 ^ 1'b0 ;
  assign n10842 = n5161 ^ n3053 ^ 1'b0 ;
  assign n10843 = n3477 & ~n10098 ;
  assign n10844 = n10843 ^ n514 ^ 1'b0 ;
  assign n10845 = n10842 | n10844 ;
  assign n10846 = n6207 ^ n4541 ^ 1'b0 ;
  assign n10847 = n613 | n1019 ;
  assign n10848 = n6782 & ~n10847 ;
  assign n10849 = n10846 & n10848 ;
  assign n10850 = n9081 ^ n7661 ^ 1'b0 ;
  assign n10851 = n8125 ^ n4229 ^ 1'b0 ;
  assign n10852 = ~n7429 & n10851 ;
  assign n10853 = n68 & n328 ;
  assign n10855 = ~n3595 & n8523 ;
  assign n10854 = ~n6178 & n6689 ;
  assign n10856 = n10855 ^ n10854 ^ 1'b0 ;
  assign n10858 = n4217 ^ n1430 ^ 1'b0 ;
  assign n10859 = n10858 ^ n3396 ^ n1520 ;
  assign n10857 = ~n670 & n732 ;
  assign n10860 = n10859 ^ n10857 ^ n6039 ;
  assign n10861 = n9846 | n10860 ;
  assign n10862 = n3861 | n4581 ;
  assign n10863 = n10489 & n10862 ;
  assign n10864 = n10861 & n10863 ;
  assign n10865 = n9812 ^ n4625 ^ 1'b0 ;
  assign n10869 = n159 & n2511 ;
  assign n10870 = n5891 & n10869 ;
  assign n10866 = n9159 ^ n5756 ^ 1'b0 ;
  assign n10867 = n1686 & n10866 ;
  assign n10868 = ~n10432 & n10867 ;
  assign n10871 = n10870 ^ n10868 ^ 1'b0 ;
  assign n10872 = n1192 ^ n170 ^ 1'b0 ;
  assign n10873 = n907 | n10872 ;
  assign n10874 = ~n2222 & n10873 ;
  assign n10875 = n4581 ^ n3346 ^ 1'b0 ;
  assign n10876 = n7752 | n10875 ;
  assign n10877 = ( n2920 & ~n4561 ) | ( n2920 & n10876 ) | ( ~n4561 & n10876 ) ;
  assign n10878 = n6136 ^ n5827 ^ 1'b0 ;
  assign n10879 = ~n4172 & n10878 ;
  assign n10880 = n9895 & n10879 ;
  assign n10881 = n5205 ^ n835 ^ 1'b0 ;
  assign n10882 = n815 & ~n1945 ;
  assign n10883 = n602 | n8566 ;
  assign n10884 = n10883 ^ n7277 ^ 1'b0 ;
  assign n10885 = n5116 ^ n1186 ^ 1'b0 ;
  assign n10886 = n6577 & ~n10557 ;
  assign n10887 = n8804 ^ n1774 ^ 1'b0 ;
  assign n10894 = n1598 ^ n713 ^ 1'b0 ;
  assign n10895 = n963 | n10894 ;
  assign n10896 = n1416 | n10895 ;
  assign n10897 = n10896 ^ n2789 ^ 1'b0 ;
  assign n10888 = n7721 & ~n8465 ;
  assign n10889 = n3256 ^ n1034 ^ 1'b0 ;
  assign n10890 = n10889 ^ n423 ^ 1'b0 ;
  assign n10891 = n2880 & n10890 ;
  assign n10892 = ~n9683 & n10891 ;
  assign n10893 = ~n10888 & n10892 ;
  assign n10898 = n10897 ^ n10893 ^ 1'b0 ;
  assign n10899 = ~n10887 & n10898 ;
  assign n10900 = ( n799 & ~n2696 ) | ( n799 & n6121 ) | ( ~n2696 & n6121 ) ;
  assign n10901 = ~n713 & n10900 ;
  assign n10902 = ~n5439 & n10901 ;
  assign n10903 = ~n7597 & n9091 ;
  assign n10904 = n878 & n5294 ;
  assign n10905 = n6279 & n10904 ;
  assign n10906 = n10905 ^ n2472 ^ 1'b0 ;
  assign n10907 = n2551 ^ n2550 ^ 1'b0 ;
  assign n10908 = n3355 & ~n10907 ;
  assign n10909 = n3211 & n10908 ;
  assign n10910 = ~n122 & n3101 ;
  assign n10911 = ~n1090 & n10910 ;
  assign n10912 = ~n3137 & n6095 ;
  assign n10913 = n10911 & n10912 ;
  assign n10914 = n2704 & n3133 ;
  assign n10915 = n4370 ^ n2536 ^ 1'b0 ;
  assign n10916 = n3349 | n10915 ;
  assign n10917 = n715 & n1789 ;
  assign n10918 = n10917 ^ n732 ^ 1'b0 ;
  assign n10919 = n1226 & ~n10918 ;
  assign n10920 = ~n769 & n5254 ;
  assign n10921 = ~n840 & n10920 ;
  assign n10922 = n5273 & n10921 ;
  assign n10923 = n4825 & n10666 ;
  assign n10924 = n10565 ^ n439 ^ 1'b0 ;
  assign n10925 = n102 | n321 ;
  assign n10926 = n7814 ^ n5713 ^ 1'b0 ;
  assign n10927 = ~n2076 & n3022 ;
  assign n10928 = ( ~n2354 & n6735 ) | ( ~n2354 & n9955 ) | ( n6735 & n9955 ) ;
  assign n10929 = n10927 & ~n10928 ;
  assign n10930 = n799 & n10929 ;
  assign n10931 = n4552 | n6156 ;
  assign n10932 = n10931 ^ n630 ^ 1'b0 ;
  assign n10933 = ~n2866 & n10932 ;
  assign n10934 = n6295 & ~n8863 ;
  assign n10935 = n3940 ^ n2101 ^ 1'b0 ;
  assign n10936 = n7087 | n10935 ;
  assign n10937 = n6930 & ~n10936 ;
  assign n10938 = ~n4606 & n10937 ;
  assign n10939 = n5706 ^ n161 ^ 1'b0 ;
  assign n10940 = ~n8827 & n10939 ;
  assign n10941 = n9944 ^ n357 ^ 1'b0 ;
  assign n10942 = n1950 ^ n1096 ^ 1'b0 ;
  assign n10943 = n10942 ^ n2122 ^ 1'b0 ;
  assign n10944 = n10941 | n10943 ;
  assign n10945 = n10941 & ~n10944 ;
  assign n10946 = n5269 ^ n307 ^ n17 ;
  assign n10947 = n10946 ^ n8092 ^ 1'b0 ;
  assign n10948 = n6392 ^ n561 ^ 1'b0 ;
  assign n10949 = n9335 & n10948 ;
  assign n10950 = n10841 & ~n10949 ;
  assign n10951 = n467 ^ n357 ^ 1'b0 ;
  assign n10955 = n9768 ^ n4334 ^ 1'b0 ;
  assign n10956 = ~n2422 & n10955 ;
  assign n10957 = n10956 ^ n1790 ^ 1'b0 ;
  assign n10952 = ~n5223 & n5778 ;
  assign n10953 = n1924 & ~n10952 ;
  assign n10954 = n10953 ^ n794 ^ 1'b0 ;
  assign n10958 = n10957 ^ n10954 ^ 1'b0 ;
  assign n10959 = n2251 & ~n7060 ;
  assign n10960 = ~n497 & n10959 ;
  assign n10961 = n9994 & ~n10960 ;
  assign n10962 = ~n3685 & n10961 ;
  assign n10963 = n4794 | n10962 ;
  assign n10964 = ~n488 & n1750 ;
  assign n10965 = n4860 ^ n1367 ^ 1'b0 ;
  assign n10967 = n5506 ^ n1479 ^ 1'b0 ;
  assign n10966 = n1430 ^ n257 ^ 1'b0 ;
  assign n10968 = n10967 ^ n10966 ^ 1'b0 ;
  assign n10969 = n3341 ^ n784 ^ 1'b0 ;
  assign n10970 = x0 | n10969 ;
  assign n10971 = ~n5343 & n8210 ;
  assign n10973 = n3483 ^ n1112 ^ 1'b0 ;
  assign n10972 = n252 | n1184 ;
  assign n10974 = n10973 ^ n10972 ^ 1'b0 ;
  assign n10975 = n10971 & n10974 ;
  assign n10976 = ~n79 & n4000 ;
  assign n10977 = ( ~n30 & n9212 ) | ( ~n30 & n10976 ) | ( n9212 & n10976 ) ;
  assign n10980 = n2140 | n8276 ;
  assign n10981 = n8412 | n10980 ;
  assign n10982 = n10981 ^ n4088 ^ 1'b0 ;
  assign n10978 = n710 & ~n7596 ;
  assign n10979 = n1026 | n10978 ;
  assign n10983 = n10982 ^ n10979 ^ 1'b0 ;
  assign n10984 = ( n293 & n3648 ) | ( n293 & n10269 ) | ( n3648 & n10269 ) ;
  assign n10985 = n2869 ^ n977 ^ 1'b0 ;
  assign n10990 = n5040 ^ n4564 ^ n659 ;
  assign n10986 = n4453 ^ n1277 ^ 1'b0 ;
  assign n10987 = n133 | n10986 ;
  assign n10988 = ~n5055 & n10987 ;
  assign n10989 = n8763 & ~n10988 ;
  assign n10991 = n10990 ^ n10989 ^ 1'b0 ;
  assign n10992 = n1235 & n3186 ;
  assign n10993 = ~n3033 & n5484 ;
  assign n10994 = ~n4812 & n10993 ;
  assign n10995 = n1473 & ~n10994 ;
  assign n10996 = n4355 ^ n998 ^ 1'b0 ;
  assign n10997 = ~n4907 & n6498 ;
  assign n10998 = n10997 ^ n2295 ^ 1'b0 ;
  assign n10999 = n3106 ^ n167 ^ 1'b0 ;
  assign n11000 = n235 & ~n10999 ;
  assign n11001 = n2367 & n3887 ;
  assign n11002 = n7753 & n11001 ;
  assign n11003 = n2065 & n2352 ;
  assign n11004 = ~n3411 & n11003 ;
  assign n11005 = n6449 & n11004 ;
  assign n11006 = n4180 & ~n6558 ;
  assign n11007 = n11006 ^ n144 ^ 1'b0 ;
  assign n11008 = n2347 & n6406 ;
  assign n11009 = n4777 & ~n7265 ;
  assign n11010 = ~n11008 & n11009 ;
  assign n11011 = n216 | n1003 ;
  assign n11012 = n2494 & ~n11011 ;
  assign n11013 = n3104 & n9808 ;
  assign n11014 = ~n3104 & n11013 ;
  assign n11015 = n6992 & ~n11014 ;
  assign n11016 = n11015 ^ n8701 ^ 1'b0 ;
  assign n11018 = n3896 ^ n2034 ^ 1'b0 ;
  assign n11019 = n11018 ^ n10435 ^ n2819 ;
  assign n11017 = n1453 & ~n4060 ;
  assign n11020 = n11019 ^ n11017 ^ 1'b0 ;
  assign n11021 = n213 & ~n9461 ;
  assign n11022 = n1209 & ~n11021 ;
  assign n11023 = ~n6887 & n11022 ;
  assign n11025 = n172 & n1669 ;
  assign n11024 = ( n685 & ~n2254 ) | ( n685 & n2654 ) | ( ~n2254 & n2654 ) ;
  assign n11026 = n11025 ^ n11024 ^ 1'b0 ;
  assign n11027 = n2356 ^ n1496 ^ 1'b0 ;
  assign n11028 = n4229 ^ n1257 ^ n184 ;
  assign n11029 = ~n5375 & n9179 ;
  assign n11030 = n11029 ^ n816 ^ 1'b0 ;
  assign n11031 = n11028 & ~n11030 ;
  assign n11032 = ~n5193 & n11031 ;
  assign n11033 = n6442 ^ n3188 ^ 1'b0 ;
  assign n11034 = n11033 ^ n406 ^ 1'b0 ;
  assign n11035 = n4722 & ~n11034 ;
  assign n11036 = ( n469 & n4401 ) | ( n469 & ~n6037 ) | ( n4401 & ~n6037 ) ;
  assign n11037 = n7059 & n11036 ;
  assign n11038 = n6745 & ~n9011 ;
  assign n11039 = n11038 ^ n1095 ^ 1'b0 ;
  assign n11040 = ~n1396 & n11039 ;
  assign n11041 = n1619 ^ n1119 ^ 1'b0 ;
  assign n11042 = n8073 & n11041 ;
  assign n11043 = n1431 ^ n1234 ^ 1'b0 ;
  assign n11044 = n6272 & n11043 ;
  assign n11045 = n6133 ^ n2218 ^ 1'b0 ;
  assign n11046 = n17 | n11045 ;
  assign n11047 = n3331 & ~n5964 ;
  assign n11048 = n11046 & n11047 ;
  assign n11049 = ~n11044 & n11048 ;
  assign n11050 = ( ~n3516 & n5242 ) | ( ~n3516 & n11049 ) | ( n5242 & n11049 ) ;
  assign n11051 = ~n5282 & n10064 ;
  assign n11052 = n338 & ~n1048 ;
  assign n11053 = n11052 ^ n1254 ^ 1'b0 ;
  assign n11054 = n1057 & n11053 ;
  assign n11055 = n11054 ^ n7650 ^ 1'b0 ;
  assign n11056 = n4815 & ~n6421 ;
  assign n11062 = n4015 ^ n1759 ^ 1'b0 ;
  assign n11063 = ~n1164 & n11062 ;
  assign n11057 = n458 | n4654 ;
  assign n11058 = n4784 & n10461 ;
  assign n11059 = ~n3415 & n11058 ;
  assign n11060 = n11057 & ~n11059 ;
  assign n11061 = ~n814 & n11060 ;
  assign n11064 = n11063 ^ n11061 ^ 1'b0 ;
  assign n11065 = n4436 & ~n11064 ;
  assign n11066 = ~n231 & n587 ;
  assign n11067 = ~n204 & n11066 ;
  assign n11068 = n6837 | n11067 ;
  assign n11069 = n2496 & ~n11068 ;
  assign n11070 = ~n7110 & n8813 ;
  assign n11071 = n11070 ^ n2607 ^ 1'b0 ;
  assign n11072 = n3787 & ~n4680 ;
  assign n11073 = n11072 ^ n5063 ^ 1'b0 ;
  assign n11074 = ~n11067 & n11073 ;
  assign n11075 = n11074 ^ n7182 ^ 1'b0 ;
  assign n11076 = n6558 | n11075 ;
  assign n11077 = n9667 ^ n1812 ^ 1'b0 ;
  assign n11080 = n3967 ^ n3467 ^ 1'b0 ;
  assign n11078 = n5939 ^ n621 ^ 1'b0 ;
  assign n11079 = n2535 & ~n11078 ;
  assign n11081 = n11080 ^ n11079 ^ 1'b0 ;
  assign n11082 = n2129 & n2436 ;
  assign n11083 = n2959 & n11082 ;
  assign n11084 = n11083 ^ n128 ^ 1'b0 ;
  assign n11085 = ~n3134 & n11084 ;
  assign n11086 = n27 & ~n1348 ;
  assign n11087 = n11086 ^ n252 ^ 1'b0 ;
  assign n11088 = n5904 & n11087 ;
  assign n11089 = n3539 | n9343 ;
  assign n11090 = ( n30 & n4055 ) | ( n30 & n4057 ) | ( n4055 & n4057 ) ;
  assign n11091 = n6268 ^ n1280 ^ 1'b0 ;
  assign n11092 = n8790 & ~n11091 ;
  assign n11093 = n11090 & n11092 ;
  assign n11094 = n2745 & ~n8485 ;
  assign n11095 = n11094 ^ n3532 ^ 1'b0 ;
  assign n11096 = n10981 ^ n2431 ^ n1045 ;
  assign n11097 = n11096 ^ n8245 ^ 1'b0 ;
  assign n11098 = n11095 & n11097 ;
  assign n11099 = ~n2426 & n11098 ;
  assign n11100 = n11099 ^ n4947 ^ 1'b0 ;
  assign n11101 = n1002 ^ n944 ^ 1'b0 ;
  assign n11102 = n4981 ^ n2587 ^ 1'b0 ;
  assign n11103 = n11101 & ~n11102 ;
  assign n11104 = n354 & ~n1490 ;
  assign n11105 = ~n11103 & n11104 ;
  assign n11106 = n11100 | n11105 ;
  assign n11107 = n581 | n4487 ;
  assign n11108 = ~n227 & n9514 ;
  assign n11110 = n8956 ^ n5135 ^ 1'b0 ;
  assign n11111 = ~n4273 & n11110 ;
  assign n11112 = n10636 ^ n2524 ^ 1'b0 ;
  assign n11113 = n11111 & n11112 ;
  assign n11114 = ~n6439 & n11113 ;
  assign n11109 = ~n4796 & n10927 ;
  assign n11115 = n11114 ^ n11109 ^ 1'b0 ;
  assign n11116 = n10985 ^ n9663 ^ 1'b0 ;
  assign n11117 = n748 & ~n3139 ;
  assign n11118 = n2339 ^ n816 ^ 1'b0 ;
  assign n11119 = n2138 | n11118 ;
  assign n11120 = ~n11117 & n11119 ;
  assign n11121 = n11056 ^ n7088 ^ 1'b0 ;
  assign n11122 = n8914 | n11121 ;
  assign n11123 = n3593 | n9118 ;
  assign n11124 = ~n6916 & n10234 ;
  assign n11125 = n666 & n2142 ;
  assign n11126 = n11125 ^ n553 ^ 1'b0 ;
  assign n11127 = n8130 ^ n6999 ^ n3143 ;
  assign n11129 = x0 & ~n514 ;
  assign n11130 = n11129 ^ n520 ^ 1'b0 ;
  assign n11128 = ~n594 & n4193 ;
  assign n11131 = n11130 ^ n11128 ^ 1'b0 ;
  assign n11132 = n1909 | n2611 ;
  assign n11133 = n221 | n4778 ;
  assign n11134 = n3877 | n8886 ;
  assign n11135 = n7149 | n11134 ;
  assign n11136 = n853 & ~n11135 ;
  assign n11137 = n573 & n1640 ;
  assign n11138 = ~n1640 & n11137 ;
  assign n11139 = n775 & ~n11138 ;
  assign n11140 = n11138 & n11139 ;
  assign n11141 = n5162 & n11140 ;
  assign n11142 = n60 | n177 ;
  assign n11143 = n177 & ~n11142 ;
  assign n11144 = n555 & n1008 ;
  assign n11145 = ~n555 & n11144 ;
  assign n11146 = n11143 | n11145 ;
  assign n11147 = n11143 & ~n11146 ;
  assign n11148 = n11147 ^ n7046 ^ 1'b0 ;
  assign n11149 = n279 & ~n1339 ;
  assign n11150 = ~n4814 & n11149 ;
  assign n11151 = n11148 & ~n11150 ;
  assign n11152 = n11141 & n11151 ;
  assign n11153 = ( ~n86 & n441 ) | ( ~n86 & n7445 ) | ( n441 & n7445 ) ;
  assign n11154 = n10177 ^ n931 ^ 1'b0 ;
  assign n11155 = n901 & n11154 ;
  assign n11156 = n2096 & n11155 ;
  assign n11157 = n11156 ^ n8351 ^ 1'b0 ;
  assign n11158 = n4360 ^ n832 ^ 1'b0 ;
  assign n11159 = n6400 ^ n2316 ^ 1'b0 ;
  assign n11160 = n11159 ^ n719 ^ 1'b0 ;
  assign n11163 = ~n2951 & n5713 ;
  assign n11164 = ~n184 & n11163 ;
  assign n11165 = n4070 & ~n11164 ;
  assign n11166 = n721 | n4963 ;
  assign n11167 = n11166 ^ n701 ^ 1'b0 ;
  assign n11168 = n2114 | n11167 ;
  assign n11169 = n6712 ^ n43 ^ 1'b0 ;
  assign n11170 = n11168 | n11169 ;
  assign n11171 = n11165 & ~n11170 ;
  assign n11172 = n11171 ^ n163 ^ 1'b0 ;
  assign n11173 = ~n3561 & n11172 ;
  assign n11174 = n8705 & n11173 ;
  assign n11161 = n6808 & ~n8135 ;
  assign n11162 = n11161 ^ n10080 ^ 1'b0 ;
  assign n11175 = n11174 ^ n11162 ^ n9360 ;
  assign n11176 = ~n5568 & n10968 ;
  assign n11177 = n1229 & n11176 ;
  assign n11178 = n477 ^ x0 ^ 1'b0 ;
  assign n11179 = n2577 & n11178 ;
  assign n11180 = n4295 & n11179 ;
  assign n11181 = n11180 ^ n1090 ^ 1'b0 ;
  assign n11182 = n1888 | n11181 ;
  assign n11183 = n667 | n4453 ;
  assign n11184 = n456 ^ n419 ^ 1'b0 ;
  assign n11185 = n11183 & n11184 ;
  assign n11186 = n11185 ^ n1931 ^ n1469 ;
  assign n11187 = n7126 ^ n1893 ^ 1'b0 ;
  assign n11188 = n11187 ^ n8128 ^ 1'b0 ;
  assign n11189 = n5056 | n10600 ;
  assign n11190 = n7060 & n9094 ;
  assign n11191 = n11190 ^ x2 ^ 1'b0 ;
  assign n11192 = n508 | n8822 ;
  assign n11193 = n11191 & ~n11192 ;
  assign n11196 = n495 & n2130 ;
  assign n11197 = n7710 & n11196 ;
  assign n11194 = n101 & n459 ;
  assign n11195 = ~n5826 & n11194 ;
  assign n11198 = n11197 ^ n11195 ^ 1'b0 ;
  assign n11199 = n7606 & n11198 ;
  assign n11200 = n3692 | n4503 ;
  assign n11201 = n11200 ^ n788 ^ 1'b0 ;
  assign n11202 = ( n3382 & ~n6401 ) | ( n3382 & n11201 ) | ( ~n6401 & n11201 ) ;
  assign n11203 = n11199 & ~n11202 ;
  assign n11204 = n107 & ~n11112 ;
  assign n11205 = ~n3040 & n6090 ;
  assign n11206 = n4139 | n11205 ;
  assign n11207 = n11206 ^ n2272 ^ 1'b0 ;
  assign n11208 = n8566 ^ n1364 ^ 1'b0 ;
  assign n11209 = n10229 | n11208 ;
  assign n11210 = n7045 ^ n6729 ^ 1'b0 ;
  assign n11211 = n7144 ^ n475 ^ 1'b0 ;
  assign n11212 = n1106 & ~n1866 ;
  assign n11213 = n5449 & ~n11212 ;
  assign n11214 = n11212 & n11213 ;
  assign n11215 = n3878 & ~n11214 ;
  assign n11216 = ~n3878 & n11215 ;
  assign n11217 = ~n302 & n704 ;
  assign n11218 = n11217 ^ n252 ^ 1'b0 ;
  assign n11219 = n3487 ^ n3446 ^ n375 ;
  assign n11220 = ~n11218 & n11219 ;
  assign n11221 = n8088 | n11220 ;
  assign n11222 = n11221 ^ n1783 ^ 1'b0 ;
  assign n11223 = n1745 & ~n4842 ;
  assign n11224 = n3311 & n11223 ;
  assign n11225 = n2333 ^ n977 ^ 1'b0 ;
  assign n11226 = n3477 & n11225 ;
  assign n11227 = n1127 | n6843 ;
  assign n11228 = n11227 ^ n7494 ^ 1'b0 ;
  assign n11229 = n5702 & ~n11228 ;
  assign n11230 = n11229 ^ n7290 ^ 1'b0 ;
  assign n11231 = n11230 ^ n8848 ^ 1'b0 ;
  assign n11232 = n11226 & ~n11231 ;
  assign n11233 = n832 & ~n4042 ;
  assign n11234 = n723 | n10618 ;
  assign n11235 = n5409 & ~n11234 ;
  assign n11236 = n11233 & n11235 ;
  assign n11237 = ~n6501 & n11236 ;
  assign n11238 = n2124 | n7726 ;
  assign n11239 = n3787 ^ n3584 ^ 1'b0 ;
  assign n11244 = n6484 ^ n1425 ^ 1'b0 ;
  assign n11240 = n3943 & ~n6558 ;
  assign n11241 = n11240 ^ n4722 ^ 1'b0 ;
  assign n11242 = n4993 | n11241 ;
  assign n11243 = n6308 & n11242 ;
  assign n11245 = n11244 ^ n11243 ^ 1'b0 ;
  assign n11246 = n11245 ^ n4626 ^ 1'b0 ;
  assign n11247 = ~n4537 & n5111 ;
  assign n11248 = n11247 ^ n777 ^ 1'b0 ;
  assign n11249 = n2162 ^ n930 ^ 1'b0 ;
  assign n11250 = n11248 | n11249 ;
  assign n11251 = n7041 & ~n10346 ;
  assign n11252 = ~n3492 & n11251 ;
  assign n11253 = n11252 ^ n8395 ^ 1'b0 ;
  assign n11254 = n4419 & n7678 ;
  assign n11255 = n9105 & ~n11254 ;
  assign n11256 = ~n3679 & n8608 ;
  assign n11257 = n3312 | n9763 ;
  assign n11258 = n3219 | n11257 ;
  assign n11259 = n11258 ^ n2668 ^ n390 ;
  assign n11260 = ~n5752 & n11259 ;
  assign n11261 = n5241 & n11260 ;
  assign n11262 = n2249 ^ n1535 ^ 1'b0 ;
  assign n11263 = n5461 & ~n11262 ;
  assign n11264 = ~n782 & n11263 ;
  assign n11265 = n2883 ^ n1394 ^ 1'b0 ;
  assign n11266 = n457 & n11265 ;
  assign n11267 = n10059 ^ n7424 ^ 1'b0 ;
  assign n11268 = n1263 & ~n9971 ;
  assign n11269 = n89 & ~n1115 ;
  assign n11270 = ( n7977 & ~n10509 ) | ( n7977 & n11269 ) | ( ~n10509 & n11269 ) ;
  assign n11271 = n9492 ^ n1197 ^ 1'b0 ;
  assign n11272 = ~n2819 & n11271 ;
  assign n11273 = n9589 ^ n2733 ^ 1'b0 ;
  assign n11274 = n3579 & ~n11273 ;
  assign n11275 = n6758 ^ n4183 ^ 1'b0 ;
  assign n11276 = n7451 ^ n470 ^ 1'b0 ;
  assign n11277 = n6090 ^ n137 ^ 1'b0 ;
  assign n11278 = n11277 ^ n1081 ^ 1'b0 ;
  assign n11279 = n2835 | n11278 ;
  assign n11280 = n3265 & ~n9535 ;
  assign n11281 = n11280 ^ n3210 ^ 1'b0 ;
  assign n11283 = n30 & n1049 ;
  assign n11282 = ~n1437 & n4441 ;
  assign n11284 = n11283 ^ n11282 ^ 1'b0 ;
  assign n11285 = n1652 | n11284 ;
  assign n11286 = n5653 & ~n11285 ;
  assign n11287 = n3406 & ~n11286 ;
  assign n11288 = ~n2266 & n11287 ;
  assign n11289 = n6349 ^ n1409 ^ x2 ;
  assign n11290 = n1048 & ~n3804 ;
  assign n11291 = n11290 ^ n7444 ^ 1'b0 ;
  assign n11292 = ~n11289 & n11291 ;
  assign n11293 = n11288 & n11292 ;
  assign n11294 = n9394 ^ n163 ^ 1'b0 ;
  assign n11295 = n814 & n1165 ;
  assign n11296 = n10338 ^ n7142 ^ 1'b0 ;
  assign n11297 = n6326 ^ n3180 ^ 1'b0 ;
  assign n11298 = n6463 & n11297 ;
  assign n11299 = n1521 & n11298 ;
  assign n11300 = n2050 & n4884 ;
  assign n11301 = ~n1856 & n11300 ;
  assign n11302 = n9794 ^ n1600 ^ 1'b0 ;
  assign n11303 = ~n5885 & n7108 ;
  assign n11304 = n7201 & n11303 ;
  assign n11305 = n338 & n1539 ;
  assign n11306 = n3559 & n3744 ;
  assign n11307 = n11305 & n11306 ;
  assign n11311 = n3452 & ~n4554 ;
  assign n11310 = n83 & ~n954 ;
  assign n11312 = n11311 ^ n11310 ^ 1'b0 ;
  assign n11313 = n1080 | n11312 ;
  assign n11308 = n2318 ^ x2 ^ 1'b0 ;
  assign n11309 = n6738 & n11308 ;
  assign n11314 = n11313 ^ n11309 ^ 1'b0 ;
  assign n11315 = n5162 & ~n11314 ;
  assign n11316 = n10772 ^ n4677 ^ n3025 ;
  assign n11317 = ( n161 & n2509 ) | ( n161 & ~n2828 ) | ( n2509 & ~n2828 ) ;
  assign n11318 = n1047 | n3080 ;
  assign n11319 = n11318 ^ n5073 ^ 1'b0 ;
  assign n11320 = n2297 | n11319 ;
  assign n11321 = n10084 & ~n11320 ;
  assign n11322 = ~n102 & n1359 ;
  assign n11323 = n9321 & ~n11322 ;
  assign n11324 = ~n2018 & n3803 ;
  assign n11325 = ~n4604 & n11324 ;
  assign n11326 = n1472 & n11325 ;
  assign n11327 = n278 ^ n159 ^ 1'b0 ;
  assign n11328 = ~n445 & n11327 ;
  assign n11329 = n1800 & n11328 ;
  assign n11330 = n7999 ^ n5376 ^ 1'b0 ;
  assign n11333 = n8539 ^ n5749 ^ 1'b0 ;
  assign n11331 = n142 | n532 ;
  assign n11332 = n11331 ^ n6397 ^ 1'b0 ;
  assign n11334 = n11333 ^ n11332 ^ 1'b0 ;
  assign n11335 = n11334 ^ n7787 ^ n294 ;
  assign n11336 = ( n988 & n1496 ) | ( n988 & ~n9441 ) | ( n1496 & ~n9441 ) ;
  assign n11337 = n101 & n501 ;
  assign n11338 = n11336 & n11337 ;
  assign n11339 = n11338 ^ n811 ^ 1'b0 ;
  assign n11340 = n2178 | n11339 ;
  assign n11341 = n10878 ^ n328 ^ 1'b0 ;
  assign n11342 = n10611 | n11341 ;
  assign n11343 = n3009 | n10001 ;
  assign n11344 = ~n2367 & n3603 ;
  assign n11345 = n4647 & n11344 ;
  assign n11346 = n5836 & n11345 ;
  assign n11347 = n665 | n3162 ;
  assign n11348 = n11347 ^ n3998 ^ 1'b0 ;
  assign n11349 = n2386 | n8399 ;
  assign n11350 = n6152 ^ n5525 ^ n5284 ;
  assign n11351 = ( n2460 & n5538 ) | ( n2460 & n11350 ) | ( n5538 & n11350 ) ;
  assign n11352 = n7518 & n8991 ;
  assign n11353 = ~n6746 & n11352 ;
  assign n11354 = n2880 & ~n3586 ;
  assign n11355 = n2771 & n11354 ;
  assign n11356 = n578 & ~n4907 ;
  assign n11357 = n11356 ^ n19 ^ 1'b0 ;
  assign n11358 = n2086 & ~n7331 ;
  assign n11359 = n638 & ~n3844 ;
  assign n11360 = n8415 | n11359 ;
  assign n11361 = ~n5794 & n10691 ;
  assign n11362 = n10576 ^ n1984 ^ 1'b0 ;
  assign n11363 = ~n1545 & n11362 ;
  assign n11364 = n2244 ^ n2075 ^ 1'b0 ;
  assign n11365 = n11364 ^ n653 ^ 1'b0 ;
  assign n11366 = n11365 ^ n8521 ^ 1'b0 ;
  assign n11367 = ~n5650 & n11366 ;
  assign n11368 = n11114 ^ n8220 ^ 1'b0 ;
  assign n11369 = ~n6493 & n9290 ;
  assign n11370 = ~n785 & n4677 ;
  assign n11371 = ~n1431 & n11370 ;
  assign n11372 = n2672 ^ n671 ^ 1'b0 ;
  assign n11373 = n1040 & ~n11372 ;
  assign n11374 = n163 | n11373 ;
  assign n11375 = n7329 ^ n5178 ^ 1'b0 ;
  assign n11376 = ~n3182 & n3785 ;
  assign n11377 = ( n142 & n2899 ) | ( n142 & ~n11376 ) | ( n2899 & ~n11376 ) ;
  assign n11378 = ~n10025 & n11377 ;
  assign n11379 = n6683 | n11378 ;
  assign n11381 = n3276 ^ n1113 ^ 1'b0 ;
  assign n11382 = n1710 & n11381 ;
  assign n11383 = n1800 & n11382 ;
  assign n11384 = n11383 ^ n1734 ^ 1'b0 ;
  assign n11380 = n6846 & ~n7590 ;
  assign n11385 = n11384 ^ n11380 ^ 1'b0 ;
  assign n11386 = n3575 & n5113 ;
  assign n11387 = n2642 & n11386 ;
  assign n11388 = n11387 ^ n9419 ^ n9002 ;
  assign n11389 = ~n9931 & n11388 ;
  assign n11390 = n616 & ~n2059 ;
  assign n11391 = n4904 ^ n273 ^ 1'b0 ;
  assign n11392 = n3176 & n6552 ;
  assign n11393 = n11392 ^ n8254 ^ 1'b0 ;
  assign n11394 = n7208 | n10690 ;
  assign n11395 = n6745 ^ n2983 ^ n522 ;
  assign n11396 = n11395 ^ n3511 ^ 1'b0 ;
  assign n11397 = n3131 & n11396 ;
  assign n11398 = ~n141 & n3796 ;
  assign n11399 = n11398 ^ n532 ^ 1'b0 ;
  assign n11400 = ~n8111 & n11399 ;
  assign n11401 = n10514 ^ n4993 ^ n1137 ;
  assign n11402 = n8998 ^ n8382 ^ 1'b0 ;
  assign n11403 = n4666 ^ n3143 ^ n1958 ;
  assign n11404 = n11403 ^ n5530 ^ 1'b0 ;
  assign n11405 = n7432 & ~n8229 ;
  assign n11406 = ~n1925 & n3600 ;
  assign n11407 = n3366 & n10791 ;
  assign n11408 = n5348 & ~n11407 ;
  assign n11409 = n7647 & n11408 ;
  assign n11410 = n10168 ^ n687 ^ 1'b0 ;
  assign n11411 = n7958 & n8408 ;
  assign n11412 = n695 & n11411 ;
  assign n11413 = n8639 ^ n8161 ^ n7361 ;
  assign n11414 = n470 & ~n7315 ;
  assign n11415 = n1118 & n11414 ;
  assign n11416 = n9096 ^ n690 ^ 1'b0 ;
  assign n11417 = ~n4407 & n11416 ;
  assign n11418 = n2843 | n7380 ;
  assign n11419 = n11417 | n11418 ;
  assign n11420 = n1728 ^ n1673 ^ 1'b0 ;
  assign n11421 = n4511 & ~n11420 ;
  assign n11422 = n11421 ^ n2354 ^ 1'b0 ;
  assign n11423 = n8761 & n11422 ;
  assign n11424 = n10429 ^ n1920 ^ n1164 ;
  assign n11425 = n11424 ^ n1325 ^ 1'b0 ;
  assign n11426 = n4021 & n5650 ;
  assign n11427 = n4479 & ~n7944 ;
  assign n11428 = n11427 ^ n6777 ^ 1'b0 ;
  assign n11429 = n11239 & ~n11428 ;
  assign n11430 = n111 & ~n6725 ;
  assign n11431 = n520 & ~n11430 ;
  assign n11432 = n6445 ^ n159 ^ 1'b0 ;
  assign n11433 = n2880 & ~n11432 ;
  assign n11434 = n11433 ^ n665 ^ 1'b0 ;
  assign n11435 = ~n86 & n276 ;
  assign n11436 = n9022 ^ n2774 ^ 1'b0 ;
  assign n11437 = n4836 | n5739 ;
  assign n11438 = n1601 | n3214 ;
  assign n11439 = n10995 ^ n1974 ^ 1'b0 ;
  assign n11441 = n3717 | n5887 ;
  assign n11442 = n11441 ^ n66 ^ 1'b0 ;
  assign n11440 = n397 & ~n1044 ;
  assign n11443 = n11442 ^ n11440 ^ 1'b0 ;
  assign n11444 = n5704 & ~n11443 ;
  assign n11445 = ~n1835 & n4506 ;
  assign n11446 = n2100 & n11445 ;
  assign n11447 = ~n10685 & n11446 ;
  assign n11448 = n7713 ^ n1274 ^ 1'b0 ;
  assign n11449 = n5922 & ~n8327 ;
  assign n11450 = n9768 ^ n5837 ^ 1'b0 ;
  assign n11451 = n2578 & ~n11450 ;
  assign n11452 = ~n5106 & n11451 ;
  assign n11453 = ~n142 & n2219 ;
  assign n11454 = n3137 & n11453 ;
  assign n11455 = ~n11453 & n11454 ;
  assign n11456 = n2700 & n11455 ;
  assign n11457 = n36 & n11456 ;
  assign n11458 = ~n10575 & n11457 ;
  assign n11459 = ~n444 & n2074 ;
  assign n11460 = ~n387 & n11459 ;
  assign n11461 = n2566 | n11460 ;
  assign n11462 = n1546 & ~n11461 ;
  assign n11463 = n3730 & n10057 ;
  assign n11464 = ( n2822 & n2911 ) | ( n2822 & n11463 ) | ( n2911 & n11463 ) ;
  assign n11465 = n11464 ^ n8370 ^ 1'b0 ;
  assign n11466 = n7046 ^ n55 ^ 1'b0 ;
  assign n11467 = n6933 & ~n11407 ;
  assign n11468 = n11467 ^ n9779 ^ 1'b0 ;
  assign n11469 = n11468 ^ n653 ^ 1'b0 ;
  assign n11470 = n9197 & n11469 ;
  assign n11471 = n11466 & n11470 ;
  assign n11472 = n4879 ^ n4554 ^ 1'b0 ;
  assign n11473 = ~n753 & n5286 ;
  assign n11474 = n11473 ^ n1406 ^ 1'b0 ;
  assign n11475 = ~n3758 & n11474 ;
  assign n11476 = n11475 ^ n7506 ^ 1'b0 ;
  assign n11477 = n11476 ^ n8574 ^ 1'b0 ;
  assign n11478 = n11472 | n11477 ;
  assign n11479 = ~n321 & n677 ;
  assign n11480 = n2414 | n3787 ;
  assign n11481 = n11480 ^ n10427 ^ 1'b0 ;
  assign n11482 = ~n2514 & n10505 ;
  assign n11483 = n11482 ^ n10587 ^ 1'b0 ;
  assign n11484 = n3552 & ~n11483 ;
  assign n11485 = n11484 ^ n1937 ^ 1'b0 ;
  assign n11486 = n3415 & ~n4299 ;
  assign n11487 = n1895 & ~n2426 ;
  assign n11488 = n4034 & n11487 ;
  assign n11489 = n3180 & ~n11049 ;
  assign n11490 = ~n11488 & n11489 ;
  assign n11491 = n11490 ^ n7381 ^ 1'b0 ;
  assign n11492 = n2835 & n7871 ;
  assign n11493 = n4954 ^ n363 ^ 1'b0 ;
  assign n11494 = n1492 & n1734 ;
  assign n11495 = n1213 | n7444 ;
  assign n11496 = n1439 | n11495 ;
  assign n11497 = n1984 & n11496 ;
  assign n11498 = ~n7846 & n11497 ;
  assign n11499 = n11494 | n11498 ;
  assign n11500 = n5501 & ~n6743 ;
  assign n11501 = ~n4507 & n11500 ;
  assign n11502 = n236 & ~n9695 ;
  assign n11503 = n7077 | n11502 ;
  assign n11504 = n7711 ^ n970 ^ 1'b0 ;
  assign n11505 = n4473 | n11504 ;
  assign n11506 = n1880 & ~n11505 ;
  assign n11507 = n7029 ^ n4574 ^ 1'b0 ;
  assign n11508 = n4759 & n11507 ;
  assign n11509 = n1002 & n11508 ;
  assign n11510 = ~n5551 & n11509 ;
  assign n11512 = n3743 & ~n10259 ;
  assign n11511 = n2768 & n4908 ;
  assign n11513 = n11512 ^ n11511 ^ 1'b0 ;
  assign n11514 = n8046 ^ n5914 ^ 1'b0 ;
  assign n11515 = n10053 ^ n7928 ^ 1'b0 ;
  assign n11516 = n3211 | n5152 ;
  assign n11517 = n7261 ^ n862 ^ 1'b0 ;
  assign n11518 = ~n2764 & n11517 ;
  assign n11520 = n1590 | n1851 ;
  assign n11521 = n4369 & n6967 ;
  assign n11522 = ~n288 & n11521 ;
  assign n11523 = ~n11520 & n11522 ;
  assign n11519 = n359 & n614 ;
  assign n11524 = n11523 ^ n11519 ^ 1'b0 ;
  assign n11525 = n1067 & n10674 ;
  assign n11526 = n6910 ^ n2162 ^ 1'b0 ;
  assign n11527 = n6182 | n11526 ;
  assign n11528 = n2085 | n11527 ;
  assign n11529 = n7930 ^ n3507 ^ 1'b0 ;
  assign n11530 = n973 & ~n11529 ;
  assign n11531 = n11530 ^ n4590 ^ 1'b0 ;
  assign n11540 = n76 | n594 ;
  assign n11541 = n5459 & ~n11540 ;
  assign n11532 = n709 & ~n3566 ;
  assign n11533 = n630 | n5513 ;
  assign n11534 = n754 ^ n328 ^ 1'b0 ;
  assign n11535 = n11534 ^ n3238 ^ n1458 ;
  assign n11536 = ~n11533 & n11535 ;
  assign n11537 = ~n4765 & n11536 ;
  assign n11538 = n508 | n11537 ;
  assign n11539 = n11532 & ~n11538 ;
  assign n11542 = n11541 ^ n11539 ^ 1'b0 ;
  assign n11543 = n4838 ^ n2210 ^ 1'b0 ;
  assign n11544 = n9490 & n11464 ;
  assign n11545 = ~n11464 & n11544 ;
  assign n11546 = n1217 & n1287 ;
  assign n11547 = n4482 & ~n7853 ;
  assign n11548 = n11547 ^ n2307 ^ 1'b0 ;
  assign n11549 = n2953 ^ n1601 ^ 1'b0 ;
  assign n11550 = n11549 ^ n3177 ^ 1'b0 ;
  assign n11551 = n8874 | n11550 ;
  assign n11552 = n11551 ^ n6487 ^ 1'b0 ;
  assign n11553 = n9631 ^ n8412 ^ 1'b0 ;
  assign n11554 = ~n4469 & n6739 ;
  assign n11555 = n11553 & ~n11554 ;
  assign n11556 = ~n738 & n2071 ;
  assign n11557 = n11556 ^ n2136 ^ 1'b0 ;
  assign n11558 = n5726 ^ n5015 ^ 1'b0 ;
  assign n11559 = n626 | n11558 ;
  assign n11560 = n11559 ^ n5112 ^ 1'b0 ;
  assign n11561 = n11557 & n11560 ;
  assign n11562 = n8957 ^ n1631 ^ 1'b0 ;
  assign n11563 = n10105 ^ n553 ^ 1'b0 ;
  assign n11564 = n1271 | n2495 ;
  assign n11565 = n6475 & n11564 ;
  assign n11566 = ~n2117 & n11565 ;
  assign n11567 = n7592 & ~n11566 ;
  assign n11568 = n11563 & n11567 ;
  assign n11569 = n2629 ^ n44 ^ 1'b0 ;
  assign n11570 = n11569 ^ n10977 ^ 1'b0 ;
  assign n11577 = n1061 ^ n517 ^ 1'b0 ;
  assign n11578 = n3087 | n11577 ;
  assign n11579 = n11578 ^ n499 ^ 1'b0 ;
  assign n11580 = n11579 ^ n10216 ^ 1'b0 ;
  assign n11581 = ~n6458 & n11580 ;
  assign n11571 = n9035 ^ n1895 ^ 1'b0 ;
  assign n11572 = n5747 & ~n11571 ;
  assign n11574 = ( n1560 & n2261 ) | ( n1560 & n4929 ) | ( n2261 & n4929 ) ;
  assign n11573 = n2562 & ~n6882 ;
  assign n11575 = n11574 ^ n11573 ^ 1'b0 ;
  assign n11576 = n11572 & ~n11575 ;
  assign n11582 = n11581 ^ n11576 ^ 1'b0 ;
  assign n11583 = n4899 & n10285 ;
  assign n11584 = n8147 ^ n2083 ^ 1'b0 ;
  assign n11585 = ~n1538 & n2834 ;
  assign n11586 = n3292 & ~n7091 ;
  assign n11587 = n11585 & n11586 ;
  assign n11588 = n2339 ^ n1031 ^ 1'b0 ;
  assign n11589 = n148 & n227 ;
  assign n11590 = n11589 ^ n5638 ^ 1'b0 ;
  assign n11591 = ~n4084 & n11590 ;
  assign n11592 = n1944 & n5252 ;
  assign n11593 = n9875 & n11200 ;
  assign n11594 = n11593 ^ n817 ^ 1'b0 ;
  assign n11595 = n1061 | n2258 ;
  assign n11596 = n11595 ^ n2083 ^ 1'b0 ;
  assign n11597 = n11594 & n11596 ;
  assign n11598 = n9019 ^ n5708 ^ n4848 ;
  assign n11599 = ~n7624 & n8018 ;
  assign n11600 = ~n11286 & n11599 ;
  assign n11601 = n697 & n11084 ;
  assign n11602 = n11601 ^ n2535 ^ 1'b0 ;
  assign n11603 = n5503 | n8031 ;
  assign n11604 = n9961 ^ n5672 ^ 1'b0 ;
  assign n11608 = n9022 ^ n7642 ^ 1'b0 ;
  assign n11605 = ~n32 & n281 ;
  assign n11606 = ~n2833 & n11605 ;
  assign n11607 = n255 | n11606 ;
  assign n11609 = n11608 ^ n11607 ^ 1'b0 ;
  assign n11610 = n5183 ^ n2412 ^ 1'b0 ;
  assign n11611 = n11609 | n11610 ;
  assign n11612 = n11611 ^ n713 ^ 1'b0 ;
  assign n11613 = n952 ^ n55 ^ 1'b0 ;
  assign n11614 = n11613 ^ n688 ^ 1'b0 ;
  assign n11615 = n1684 | n11614 ;
  assign n11616 = n4491 ^ x1 ^ 1'b0 ;
  assign n11617 = ~n2966 & n11616 ;
  assign n11618 = n11617 ^ n9638 ^ 1'b0 ;
  assign n11619 = n11546 ^ n4304 ^ 1'b0 ;
  assign n11620 = n2953 & ~n4001 ;
  assign n11621 = ~n168 & n11620 ;
  assign n11622 = n11621 ^ n10833 ^ 1'b0 ;
  assign n11623 = n6989 & ~n11622 ;
  assign n11624 = n4198 ^ n1626 ^ 1'b0 ;
  assign n11625 = n2079 & n2403 ;
  assign n11626 = n8808 & n11625 ;
  assign n11627 = n2347 & n10260 ;
  assign n11628 = n10107 ^ n2433 ^ 1'b0 ;
  assign n11629 = ~n6985 & n11628 ;
  assign n11630 = n3545 ^ n1034 ^ 1'b0 ;
  assign n11631 = n939 & ~n11630 ;
  assign n11632 = n580 & n9723 ;
  assign n11633 = ~n11631 & n11632 ;
  assign n11634 = ~n5562 & n11396 ;
  assign n11635 = n8172 ^ n3589 ^ 1'b0 ;
  assign n11636 = ~n432 & n1430 ;
  assign n11637 = n4424 | n11636 ;
  assign n11638 = n2630 & ~n7117 ;
  assign n11641 = n7444 ^ n3735 ^ 1'b0 ;
  assign n11639 = n4127 ^ n412 ^ 1'b0 ;
  assign n11640 = n6781 & ~n11639 ;
  assign n11642 = n11641 ^ n11640 ^ 1'b0 ;
  assign n11643 = n4650 & ~n11642 ;
  assign n11644 = n7545 & ~n11643 ;
  assign n11645 = n2680 ^ n472 ^ 1'b0 ;
  assign n11646 = n957 & ~n11645 ;
  assign n11647 = n3762 ^ n2218 ^ 1'b0 ;
  assign n11648 = n44 & n11647 ;
  assign n11649 = ~n1884 & n6866 ;
  assign n11650 = ~n4815 & n11649 ;
  assign n11651 = n204 ^ n60 ^ 1'b0 ;
  assign n11652 = ~n11650 & n11651 ;
  assign n11653 = ~n11648 & n11652 ;
  assign n11654 = n4445 | n6889 ;
  assign n11655 = n2428 ^ n592 ^ 1'b0 ;
  assign n11656 = ~n2991 & n11655 ;
  assign n11657 = ~n7782 & n8299 ;
  assign n11658 = n11657 ^ n10156 ^ 1'b0 ;
  assign n11659 = n5218 & ~n10545 ;
  assign n11660 = n5427 | n11659 ;
  assign n11661 = n2245 | n9292 ;
  assign n11662 = n11661 ^ n5326 ^ 1'b0 ;
  assign n11663 = n5104 ^ n3150 ^ 1'b0 ;
  assign n11664 = n6303 & ~n11663 ;
  assign n11665 = n11414 ^ n6476 ^ 1'b0 ;
  assign n11666 = ~n255 & n11665 ;
  assign n11667 = ~n10882 & n11666 ;
  assign n11668 = n3925 | n7381 ;
  assign n11669 = ~n10118 & n11668 ;
  assign n11670 = n7608 ^ n4857 ^ 1'b0 ;
  assign n11671 = ~n1308 & n2514 ;
  assign n11672 = n9925 & n11671 ;
  assign n11673 = n11672 ^ n3309 ^ 1'b0 ;
  assign n11674 = n11673 ^ n1394 ^ 1'b0 ;
  assign n11675 = n8281 ^ n1226 ^ 1'b0 ;
  assign n11676 = n3180 & ~n11675 ;
  assign n11677 = n16 & ~n624 ;
  assign n11678 = n11677 ^ n6735 ^ 1'b0 ;
  assign n11679 = n7729 ^ n4446 ^ 1'b0 ;
  assign n11680 = n9032 ^ n5532 ^ 1'b0 ;
  assign n11681 = n3068 ^ n357 ^ 1'b0 ;
  assign n11682 = n11681 ^ n3284 ^ 1'b0 ;
  assign n11683 = n11682 ^ n1095 ^ 1'b0 ;
  assign n11684 = n2205 & ~n11683 ;
  assign n11685 = n417 & ~n7017 ;
  assign n11686 = n11685 ^ n153 ^ 1'b0 ;
  assign n11687 = n3402 | n7374 ;
  assign n11688 = n8558 ^ n7661 ^ 1'b0 ;
  assign n11689 = ~n5507 & n11688 ;
  assign n11690 = n11689 ^ n11261 ^ 1'b0 ;
  assign n11691 = n5646 ^ n519 ^ 1'b0 ;
  assign n11692 = n456 & ~n11691 ;
  assign n11693 = ( ~n3646 & n4136 ) | ( ~n3646 & n4606 ) | ( n4136 & n4606 ) ;
  assign n11694 = n1048 & n6370 ;
  assign n11695 = n495 & n507 ;
  assign n11696 = n11695 ^ n3671 ^ 1'b0 ;
  assign n11697 = ~n385 & n2714 ;
  assign n11698 = n11697 ^ n3338 ^ 1'b0 ;
  assign n11699 = n11698 ^ n4281 ^ 1'b0 ;
  assign n11700 = n4864 | n11699 ;
  assign n11701 = n2664 | n5455 ;
  assign n11702 = n11701 ^ n2373 ^ 1'b0 ;
  assign n11703 = n1810 & n3053 ;
  assign n11704 = n984 & n11703 ;
  assign n11705 = ~n11702 & n11704 ;
  assign n11706 = n8258 & n8412 ;
  assign n11707 = n6230 & n11706 ;
  assign n11708 = n11707 ^ n1771 ^ 1'b0 ;
  assign n11709 = ~n6995 & n11708 ;
  assign n11710 = ~n3199 & n11709 ;
  assign n11711 = n11705 & n11710 ;
  assign n11712 = n7233 ^ n6496 ^ 1'b0 ;
  assign n11713 = n1375 & ~n5308 ;
  assign n11714 = ~n1588 & n11713 ;
  assign n11715 = ~n796 & n4273 ;
  assign n11716 = n5087 | n11715 ;
  assign n11717 = n11716 ^ n4057 ^ 1'b0 ;
  assign n11718 = n2751 & ~n5903 ;
  assign n11719 = n4965 & n6419 ;
  assign n11720 = n11719 ^ n3986 ^ 1'b0 ;
  assign n11721 = n257 & ~n4756 ;
  assign n11722 = n684 & n5033 ;
  assign n11723 = n11722 ^ n11067 ^ 1'b0 ;
  assign n11724 = n989 & ~n3892 ;
  assign n11725 = n2176 ^ n1179 ^ 1'b0 ;
  assign n11726 = ~n11724 & n11725 ;
  assign n11727 = n581 & n1335 ;
  assign n11728 = n11727 ^ n712 ^ 1'b0 ;
  assign n11729 = n11728 ^ n5634 ^ 1'b0 ;
  assign n11730 = n2759 | n3130 ;
  assign n11731 = n1624 & ~n2251 ;
  assign n11732 = ( n7407 & ~n11730 ) | ( n7407 & n11731 ) | ( ~n11730 & n11731 ) ;
  assign n11733 = ~n4533 & n4954 ;
  assign n11734 = n758 | n3509 ;
  assign n11735 = n5796 & ~n6451 ;
  assign n11736 = n8644 ^ n6498 ^ 1'b0 ;
  assign n11737 = n11735 | n11736 ;
  assign n11738 = n5982 | n7973 ;
  assign n11739 = n3971 & ~n10325 ;
  assign n11740 = n11739 ^ n4977 ^ 1'b0 ;
  assign n11741 = ~n3626 & n4112 ;
  assign n11742 = n11741 ^ n4247 ^ 1'b0 ;
  assign n11743 = n3297 & ~n11742 ;
  assign n11744 = ~n839 & n11743 ;
  assign n11745 = n1236 & n11744 ;
  assign n11746 = n11745 ^ n4599 ^ 1'b0 ;
  assign n11747 = n4411 ^ n2479 ^ 1'b0 ;
  assign n11748 = n11746 & n11747 ;
  assign n11749 = n11748 ^ n11597 ^ 1'b0 ;
  assign n11750 = ~n7933 & n11749 ;
  assign n11751 = n3692 | n7278 ;
  assign n11752 = n2599 ^ n1898 ^ 1'b0 ;
  assign n11753 = n11752 ^ n7646 ^ 1'b0 ;
  assign n11754 = n512 & n5963 ;
  assign n11755 = ~n3922 & n11754 ;
  assign n11756 = n6115 ^ n3878 ^ 1'b0 ;
  assign n11757 = n3340 & ~n4660 ;
  assign n11758 = n7936 & n11757 ;
  assign n11759 = n11334 ^ n4492 ^ n4225 ;
  assign n11760 = n11759 ^ n296 ^ 1'b0 ;
  assign n11761 = n7006 ^ n741 ^ 1'b0 ;
  assign n11762 = n984 & n11761 ;
  assign n11763 = n11762 ^ n2951 ^ 1'b0 ;
  assign n11764 = n2235 & n2321 ;
  assign n11765 = n250 & n11764 ;
  assign n11766 = n2573 ^ n1095 ^ 1'b0 ;
  assign n11767 = n5876 & ~n11766 ;
  assign n11768 = n10389 & n11767 ;
  assign n11769 = n2438 & ~n11768 ;
  assign n11770 = n55 & n11769 ;
  assign n11771 = n581 & n4117 ;
  assign n11772 = n5841 | n9939 ;
  assign n11773 = n809 & ~n7949 ;
  assign n11774 = n7450 ^ n688 ^ 1'b0 ;
  assign n11775 = n8381 & n11774 ;
  assign n11776 = ~n642 & n4774 ;
  assign n11777 = n4843 ^ n2948 ^ 1'b0 ;
  assign n11778 = n5554 & n11777 ;
  assign n11779 = n4706 ^ n3856 ^ 1'b0 ;
  assign n11780 = n1287 & n11779 ;
  assign n11781 = n11780 ^ n9925 ^ 1'b0 ;
  assign n11782 = n8760 & ~n11781 ;
  assign n11783 = n4632 | n5821 ;
  assign n11784 = n8422 ^ n1571 ^ n268 ;
  assign n11785 = n8653 | n9397 ;
  assign n11786 = n4846 & ~n11785 ;
  assign n11787 = n2542 & n11786 ;
  assign n11788 = n983 | n3072 ;
  assign n11789 = n983 & ~n11788 ;
  assign n11790 = n2046 & ~n11789 ;
  assign n11791 = ~n2046 & n11790 ;
  assign n11792 = n4799 | n11791 ;
  assign n11793 = ~n3849 & n11792 ;
  assign n11794 = n3849 & n11793 ;
  assign n11795 = n1254 & ~n2939 ;
  assign n11796 = n11795 ^ n4367 ^ 1'b0 ;
  assign n11797 = n8014 ^ n6368 ^ 1'b0 ;
  assign n11798 = n8307 ^ n6845 ^ 1'b0 ;
  assign n11799 = n2613 & ~n3929 ;
  assign n11800 = n8780 & n11799 ;
  assign n11801 = n3929 ^ n395 ^ 1'b0 ;
  assign n11802 = n3861 & n11801 ;
  assign n11803 = n2531 & n11802 ;
  assign n11804 = ~n6469 & n11803 ;
  assign n11805 = n5949 & ~n8479 ;
  assign n11806 = ~n7046 & n11805 ;
  assign n11807 = n7734 & n7755 ;
  assign n11808 = n6567 ^ n28 ^ 1'b0 ;
  assign n11809 = n7383 & n11808 ;
  assign n11810 = n2670 & ~n6818 ;
  assign n11811 = n6818 & n11810 ;
  assign n11812 = ~n7782 & n11811 ;
  assign n11813 = n1632 | n2436 ;
  assign n11814 = n1632 & ~n11813 ;
  assign n11815 = n11814 ^ n5314 ^ 1'b0 ;
  assign n11816 = n11812 & ~n11815 ;
  assign n11817 = n1833 & n11816 ;
  assign n11818 = ~n11816 & n11817 ;
  assign n11819 = n1968 ^ n414 ^ 1'b0 ;
  assign n11820 = n6903 & n11819 ;
  assign n11821 = n10957 | n11820 ;
  assign n11822 = ~n827 & n4072 ;
  assign n11823 = n323 & n11822 ;
  assign n11824 = n7797 & ~n11823 ;
  assign n11825 = n3295 & n5724 ;
  assign n11826 = ~n6921 & n11825 ;
  assign n11827 = n5108 & n6053 ;
  assign n11828 = n169 | n11485 ;
  assign n11829 = n9376 | n11828 ;
  assign n11830 = n7936 | n9925 ;
  assign n11831 = n11830 ^ n937 ^ 1'b0 ;
  assign n11832 = n2216 & ~n11831 ;
  assign n11833 = n11832 ^ n4112 ^ 1'b0 ;
  assign n11834 = n11833 ^ n899 ^ 1'b0 ;
  assign n11835 = n3603 & ~n4845 ;
  assign n11836 = n571 & n11835 ;
  assign n11837 = n6898 & n11836 ;
  assign n11838 = n8455 ^ n1209 ^ 1'b0 ;
  assign n11841 = n506 ^ n283 ^ 1'b0 ;
  assign n11842 = n7007 | n11841 ;
  assign n11839 = n5208 ^ n3338 ^ 1'b0 ;
  assign n11840 = n975 & ~n11839 ;
  assign n11843 = n11842 ^ n11840 ^ 1'b0 ;
  assign n11844 = n6618 & ~n11843 ;
  assign n11846 = n2418 & ~n4256 ;
  assign n11845 = ~n4822 & n5049 ;
  assign n11847 = n11846 ^ n11845 ^ 1'b0 ;
  assign n11848 = n2311 & ~n10644 ;
  assign n11849 = n7140 & n8488 ;
  assign n11850 = n5872 | n11849 ;
  assign n11851 = n4883 ^ n366 ^ 1'b0 ;
  assign n11852 = ~n977 & n10029 ;
  assign n11853 = n6348 ^ x1 ^ 1'b0 ;
  assign n11854 = n7648 | n11853 ;
  assign n11859 = n1712 ^ n144 ^ 1'b0 ;
  assign n11855 = ( ~n493 & n1112 ) | ( ~n493 & n1711 ) | ( n1112 & n1711 ) ;
  assign n11856 = ~n10465 & n11855 ;
  assign n11857 = n11856 ^ n5148 ^ 1'b0 ;
  assign n11858 = ~n5649 & n11857 ;
  assign n11860 = n11859 ^ n11858 ^ 1'b0 ;
  assign n11861 = ~n1637 & n11860 ;
  assign n11862 = n5083 ^ n4968 ^ 1'b0 ;
  assign n11863 = n1932 ^ n1804 ^ 1'b0 ;
  assign n11864 = n1138 | n11863 ;
  assign n11865 = ~n133 & n3663 ;
  assign n11866 = n11865 ^ n690 ^ 1'b0 ;
  assign n11867 = ~n236 & n3418 ;
  assign n11868 = n11867 ^ n2076 ^ 1'b0 ;
  assign n11869 = n744 | n11868 ;
  assign n11871 = n7589 ^ n291 ^ 1'b0 ;
  assign n11872 = n4051 & ~n11871 ;
  assign n11870 = n1307 ^ n246 ^ 1'b0 ;
  assign n11873 = n11872 ^ n11870 ^ 1'b0 ;
  assign n11874 = n6892 | n11873 ;
  assign n11875 = n11777 ^ n10347 ^ 1'b0 ;
  assign n11878 = n144 | n266 ;
  assign n11879 = n144 & ~n11878 ;
  assign n11880 = n6141 | n11879 ;
  assign n11876 = n7553 ^ n929 ^ 1'b0 ;
  assign n11877 = ~n8004 & n11876 ;
  assign n11881 = n11880 ^ n11877 ^ 1'b0 ;
  assign n11882 = n11881 ^ n9428 ^ n656 ;
  assign n11883 = n4860 ^ n4054 ^ 1'b0 ;
  assign n11884 = n11883 ^ n2315 ^ 1'b0 ;
  assign n11885 = n11882 | n11884 ;
  assign n11886 = n7763 & n7814 ;
  assign n11887 = n4959 ^ n3298 ^ 1'b0 ;
  assign n11888 = n939 | n11887 ;
  assign n11889 = n5424 & n7417 ;
  assign n11890 = n8373 & n11889 ;
  assign n11891 = n11888 & n11890 ;
  assign n11892 = n403 | n654 ;
  assign n11893 = n11892 ^ n2086 ^ 1'b0 ;
  assign n11894 = n1673 | n11893 ;
  assign n11895 = n4700 & ~n10936 ;
  assign n11896 = n3219 ^ n2660 ^ 1'b0 ;
  assign n11897 = n6100 | n11896 ;
  assign n11898 = ~n323 & n11897 ;
  assign n11899 = n7461 & ~n11898 ;
  assign n11900 = ~n11895 & n11899 ;
  assign n11901 = ~n5156 & n8234 ;
  assign n11902 = n11901 ^ n850 ^ 1'b0 ;
  assign n11903 = n8629 ^ n1252 ^ 1'b0 ;
  assign n11904 = n11902 & n11903 ;
  assign n11905 = n1011 & ~n9744 ;
  assign n11906 = n9326 | n11905 ;
  assign n11907 = n11904 | n11906 ;
  assign n11908 = n1064 ^ n899 ^ 1'b0 ;
  assign n11909 = n168 & n11908 ;
  assign n11910 = n4319 ^ n3225 ^ 1'b0 ;
  assign n11911 = n2549 & ~n11910 ;
  assign n11912 = ~n3826 & n11911 ;
  assign n11915 = n683 ^ n361 ^ 1'b0 ;
  assign n11913 = ~n231 & n1170 ;
  assign n11914 = ~n2786 & n11913 ;
  assign n11916 = n11915 ^ n11914 ^ 1'b0 ;
  assign n11917 = ~n4473 & n4921 ;
  assign n11918 = ~n4889 & n5124 ;
  assign n11919 = n11918 ^ n8353 ^ 1'b0 ;
  assign n11920 = n1915 & ~n8238 ;
  assign n11921 = n5752 & n10037 ;
  assign n11922 = ~n6339 & n11921 ;
  assign n11923 = n11920 | n11922 ;
  assign n11924 = ~n11919 & n11923 ;
  assign n11925 = ~n10557 & n11924 ;
  assign n11926 = n11925 ^ n8651 ^ 1'b0 ;
  assign n11927 = n246 | n9572 ;
  assign n11928 = n3028 & ~n3162 ;
  assign n11929 = n11928 ^ n6933 ^ 1'b0 ;
  assign n11930 = n6889 ^ n3960 ^ 1'b0 ;
  assign n11931 = n271 & n11930 ;
  assign n11932 = n5394 & n11931 ;
  assign n11933 = n4790 ^ n387 ^ 1'b0 ;
  assign n11934 = ~n6916 & n9608 ;
  assign n11935 = n11934 ^ n4641 ^ 1'b0 ;
  assign n11936 = ~n11933 & n11935 ;
  assign n11937 = ~n11932 & n11936 ;
  assign n11938 = n4504 ^ n670 ^ 1'b0 ;
  assign n11939 = n9255 ^ n4807 ^ 1'b0 ;
  assign n11940 = n4165 | n11939 ;
  assign n11941 = n1887 ^ n1132 ^ 1'b0 ;
  assign n11942 = n11941 ^ n6450 ^ 1'b0 ;
  assign n11943 = ~n11940 & n11942 ;
  assign n11944 = n679 | n3959 ;
  assign n11952 = n727 | n1704 ;
  assign n11947 = ~n4400 & n10033 ;
  assign n11948 = n11947 ^ n168 ^ 1'b0 ;
  assign n11949 = n1106 & ~n11948 ;
  assign n11950 = n11949 ^ n2012 ^ 1'b0 ;
  assign n11951 = n6209 & ~n11950 ;
  assign n11953 = n11952 ^ n11951 ^ 1'b0 ;
  assign n11945 = n945 & n5033 ;
  assign n11946 = n5890 & n11945 ;
  assign n11954 = n11953 ^ n11946 ^ 1'b0 ;
  assign n11955 = ~n536 & n11954 ;
  assign n11956 = n11944 & n11955 ;
  assign n11957 = n9476 ^ n3459 ^ 1'b0 ;
  assign n11958 = n11957 ^ n1664 ^ 1'b0 ;
  assign n11959 = n8019 & ~n11958 ;
  assign n11960 = n7895 | n8472 ;
  assign n11961 = n11960 ^ n587 ^ 1'b0 ;
  assign n11962 = n3178 ^ n1654 ^ 1'b0 ;
  assign n11963 = ~n70 & n11962 ;
  assign n11964 = n88 & n11963 ;
  assign n11965 = n3974 | n11964 ;
  assign n11966 = n10482 ^ n9014 ^ 1'b0 ;
  assign n11967 = n2110 | n11966 ;
  assign n11968 = n3803 ^ n3498 ^ 1'b0 ;
  assign n11969 = ~n4422 & n11968 ;
  assign n11970 = n5123 ^ n3694 ^ 1'b0 ;
  assign n11971 = n7029 ^ n2260 ^ n799 ;
  assign n11972 = n3655 ^ n979 ^ 1'b0 ;
  assign n11973 = n8687 ^ n767 ^ 1'b0 ;
  assign n11974 = n158 | n9306 ;
  assign n11975 = n11974 ^ n903 ^ 1'b0 ;
  assign n11976 = n11975 ^ n11660 ^ 1'b0 ;
  assign n11977 = n52 & ~n11976 ;
  assign n11979 = n7093 ^ n930 ^ 1'b0 ;
  assign n11978 = n4549 & n10444 ;
  assign n11980 = n11979 ^ n11978 ^ 1'b0 ;
  assign n11981 = n6392 & n11712 ;
  assign n11982 = ~n525 & n1112 ;
  assign n11985 = ~n2127 & n2439 ;
  assign n11986 = n11985 ^ n5775 ^ 1'b0 ;
  assign n11987 = n649 | n11986 ;
  assign n11983 = n1425 & ~n2065 ;
  assign n11984 = n11681 & n11983 ;
  assign n11988 = n11987 ^ n11984 ^ 1'b0 ;
  assign n11989 = n10985 ^ n4796 ^ 1'b0 ;
  assign n11990 = n5238 & n11989 ;
  assign n11991 = n630 & n5238 ;
  assign n11992 = ~n5708 & n11991 ;
  assign n11993 = n3960 ^ n1423 ^ 1'b0 ;
  assign n11994 = n3940 | n11993 ;
  assign n11995 = ~n2657 & n5211 ;
  assign n11996 = n204 & ~n2155 ;
  assign n11997 = n11995 & n11996 ;
  assign n11998 = n2732 & ~n11997 ;
  assign n11999 = n2773 ^ n659 ^ 1'b0 ;
  assign n12000 = n2198 & n11999 ;
  assign n12001 = n233 & n12000 ;
  assign n12002 = n12001 ^ n88 ^ 1'b0 ;
  assign n12003 = n9536 ^ n8271 ^ 1'b0 ;
  assign n12004 = n8199 ^ n1940 ^ 1'b0 ;
  assign n12005 = n12003 & ~n12004 ;
  assign n12006 = n1441 & ~n11798 ;
  assign n12007 = n2553 & n4869 ;
  assign n12008 = n11178 & ~n12007 ;
  assign n12009 = n12008 ^ n3558 ^ 1'b0 ;
  assign n12010 = ~n8327 & n12009 ;
  assign n12011 = n191 | n12010 ;
  assign n12012 = n9816 & n12011 ;
  assign n12013 = n12012 ^ n7136 ^ 1'b0 ;
  assign n12014 = n542 | n1005 ;
  assign n12015 = n62 | n257 ;
  assign n12016 = n12015 ^ n75 ^ 1'b0 ;
  assign n12017 = n3742 ^ n528 ^ 1'b0 ;
  assign n12018 = ~n12016 & n12017 ;
  assign n12019 = ~n70 & n12018 ;
  assign n12020 = n5316 & ~n9736 ;
  assign n12021 = n484 | n12020 ;
  assign n12022 = n10203 ^ n3726 ^ 1'b0 ;
  assign n12024 = n5713 ^ n1875 ^ 1'b0 ;
  assign n12025 = n294 & ~n12024 ;
  assign n12023 = ~n1194 & n7548 ;
  assign n12026 = n12025 ^ n12023 ^ 1'b0 ;
  assign n12027 = n7412 ^ n6910 ^ 1'b0 ;
  assign n12028 = ~n6054 & n12027 ;
  assign n12029 = n11057 ^ n9789 ^ n3749 ;
  assign n12030 = n510 & ~n10353 ;
  assign n12031 = n10353 & n12030 ;
  assign n12032 = n12007 | n12031 ;
  assign n12033 = n12007 & ~n12032 ;
  assign n12034 = n9410 ^ n2168 ^ n300 ;
  assign n12035 = n12034 ^ n10180 ^ 1'b0 ;
  assign n12036 = n12035 ^ n8798 ^ 1'b0 ;
  assign n12037 = n1541 | n12036 ;
  assign n12044 = ~n2511 & n9001 ;
  assign n12039 = n1546 & ~n6160 ;
  assign n12038 = n3589 | n4273 ;
  assign n12040 = n12039 ^ n12038 ^ 1'b0 ;
  assign n12041 = ~n345 & n3962 ;
  assign n12042 = n3370 & n12041 ;
  assign n12043 = n12040 | n12042 ;
  assign n12045 = n12044 ^ n12043 ^ 1'b0 ;
  assign n12046 = ~n366 & n3693 ;
  assign n12047 = ~n1185 & n12046 ;
  assign n12048 = n12047 ^ n595 ^ 1'b0 ;
  assign n12049 = n10739 | n12048 ;
  assign n12050 = n3160 & n5447 ;
  assign n12051 = n9705 & n10927 ;
  assign n12052 = n3786 & n11913 ;
  assign n12053 = n3435 & n12052 ;
  assign n12054 = n12053 ^ n3292 ^ 1'b0 ;
  assign n12055 = n3522 ^ n375 ^ 1'b0 ;
  assign n12056 = n4856 | n12055 ;
  assign n12057 = n9831 ^ n3921 ^ n3589 ;
  assign n12058 = n12046 ^ n4807 ^ 1'b0 ;
  assign n12059 = n12057 | n12058 ;
  assign n12060 = ( ~n66 & n1691 ) | ( ~n66 & n7328 ) | ( n1691 & n7328 ) ;
  assign n12061 = n12060 ^ n5449 ^ 1'b0 ;
  assign n12062 = n4292 & ~n12061 ;
  assign n12063 = n6620 ^ n2684 ^ 1'b0 ;
  assign n12064 = n6585 & n12063 ;
  assign n12065 = ( ~n323 & n5267 ) | ( ~n323 & n7534 ) | ( n5267 & n7534 ) ;
  assign n12066 = ~n2136 & n12065 ;
  assign n12067 = n1492 & ~n3492 ;
  assign n12068 = n539 & n3797 ;
  assign n12069 = ~n4822 & n12068 ;
  assign n12070 = n4136 & n12069 ;
  assign n12071 = n1887 | n12070 ;
  assign n12072 = n14 & ~n12071 ;
  assign n12073 = n6691 ^ n2967 ^ 1'b0 ;
  assign n12074 = n2476 & n7894 ;
  assign n12075 = ~n6051 & n12074 ;
  assign n12076 = n208 & n12075 ;
  assign n12077 = n3088 | n4645 ;
  assign n12078 = n12077 ^ n914 ^ 1'b0 ;
  assign n12079 = n290 & n741 ;
  assign n12080 = ~n12078 & n12079 ;
  assign n12081 = n8283 ^ n917 ^ 1'b0 ;
  assign n12082 = n5928 | n12081 ;
  assign n12084 = n6432 & n8360 ;
  assign n12085 = n12084 ^ n7317 ^ 1'b0 ;
  assign n12086 = n2228 & n12085 ;
  assign n12083 = ~n4116 & n6389 ;
  assign n12087 = n12086 ^ n12083 ^ 1'b0 ;
  assign n12090 = n9219 ^ n4314 ^ 1'b0 ;
  assign n12088 = n7024 ^ n2008 ^ 1'b0 ;
  assign n12089 = ~n1159 & n12088 ;
  assign n12091 = n12090 ^ n12089 ^ 1'b0 ;
  assign n12092 = n11433 | n12091 ;
  assign n12093 = ~n2731 & n7624 ;
  assign n12094 = n2059 & n12093 ;
  assign n12095 = n12094 ^ n938 ^ 1'b0 ;
  assign n12096 = n12095 ^ n1379 ^ 1'b0 ;
  assign n12097 = n2584 & ~n12096 ;
  assign n12098 = n8713 & n12097 ;
  assign n12099 = n6128 & n12098 ;
  assign n12100 = n1152 ^ n86 ^ 1'b0 ;
  assign n12101 = n12100 ^ n804 ^ 1'b0 ;
  assign n12102 = n667 & ~n12101 ;
  assign n12103 = n6152 ^ n1645 ^ 1'b0 ;
  assign n12104 = n12102 & n12103 ;
  assign n12105 = n1467 ^ n898 ^ 1'b0 ;
  assign n12106 = n4995 & ~n12105 ;
  assign n12107 = n12106 ^ n1768 ^ 1'b0 ;
  assign n12108 = n12107 ^ n11258 ^ n977 ;
  assign n12109 = n2702 | n8158 ;
  assign n12110 = n367 | n5702 ;
  assign n12111 = n12110 ^ n25 ^ 1'b0 ;
  assign n12112 = n3609 ^ n3320 ^ 1'b0 ;
  assign n12113 = n510 & ~n12112 ;
  assign n12115 = x11 | n4344 ;
  assign n12114 = n7195 ^ n3083 ^ 1'b0 ;
  assign n12116 = n12115 ^ n12114 ^ 1'b0 ;
  assign n12117 = n3781 & n12116 ;
  assign n12118 = ~n12113 & n12117 ;
  assign n12119 = n6510 & n12118 ;
  assign n12120 = n1245 | n12119 ;
  assign n12121 = n1693 & ~n12120 ;
  assign n12122 = n630 & n5397 ;
  assign n12123 = n12122 ^ n1870 ^ 1'b0 ;
  assign n12124 = n5930 | n10346 ;
  assign n12125 = n5347 | n12124 ;
  assign n12130 = x7 & ~n30 ;
  assign n12131 = n30 & n12130 ;
  assign n12132 = x5 & n15 ;
  assign n12133 = n12131 & n12132 ;
  assign n12134 = x5 & ~n12133 ;
  assign n12135 = n12133 & n12134 ;
  assign n12136 = n43 & ~n12135 ;
  assign n12137 = ~n43 & n12136 ;
  assign n12138 = x5 & n101 ;
  assign n12139 = ~n101 & n12138 ;
  assign n12140 = n17 | n12139 ;
  assign n12141 = n12139 & ~n12140 ;
  assign n12142 = n81 & n97 ;
  assign n12143 = n12141 & n12142 ;
  assign n12144 = n96 | n12143 ;
  assign n12145 = n12143 & ~n12144 ;
  assign n12146 = n165 & ~n12145 ;
  assign n12147 = n12137 & n12146 ;
  assign n12148 = n12147 ^ n468 ^ 1'b0 ;
  assign n12149 = n1541 | n7173 ;
  assign n12150 = n4288 & n8840 ;
  assign n12151 = ~n8840 & n12150 ;
  assign n12152 = n12149 & ~n12151 ;
  assign n12153 = ~n12148 & n12152 ;
  assign n12126 = n2933 & ~n10014 ;
  assign n12127 = ~n212 & n12126 ;
  assign n12128 = n212 & n12127 ;
  assign n12129 = ~n7752 & n12128 ;
  assign n12154 = n12153 ^ n12129 ^ 1'b0 ;
  assign n12155 = n12125 & n12154 ;
  assign n12156 = n1765 & n7594 ;
  assign n12157 = n12156 ^ n4078 ^ 1'b0 ;
  assign n12158 = ~n10666 & n12157 ;
  assign n12159 = ~n68 & n12158 ;
  assign n12160 = n3185 & n5930 ;
  assign n12161 = n2762 | n12160 ;
  assign n12162 = n12161 ^ n7632 ^ 1'b0 ;
  assign n12163 = n6296 | n7182 ;
  assign n12164 = n10058 ^ n9231 ^ 1'b0 ;
  assign n12165 = ~n1066 & n12164 ;
  assign n12166 = ~n5673 & n9404 ;
  assign n12167 = n12166 ^ n3089 ^ 1'b0 ;
  assign n12168 = n4040 ^ n1342 ^ 1'b0 ;
  assign n12169 = ~n12167 & n12168 ;
  assign n12170 = n12169 ^ n6463 ^ 1'b0 ;
  assign n12171 = n1186 & n6445 ;
  assign n12172 = n9757 ^ n2509 ^ 1'b0 ;
  assign n12173 = n4804 ^ n1790 ^ 1'b0 ;
  assign n12176 = n503 & n1090 ;
  assign n12177 = n813 & n12176 ;
  assign n12174 = n6097 ^ n5057 ^ 1'b0 ;
  assign n12175 = n5732 | n12174 ;
  assign n12178 = n12177 ^ n12175 ^ 1'b0 ;
  assign n12179 = n2539 & n4320 ;
  assign n12180 = n12179 ^ n1467 ^ 1'b0 ;
  assign n12181 = n4211 ^ n3282 ^ 1'b0 ;
  assign n12182 = ~n7403 & n12181 ;
  assign n12183 = ~n6026 & n12182 ;
  assign n12184 = n12183 ^ n470 ^ 1'b0 ;
  assign n12185 = n6973 | n11266 ;
  assign n12186 = n3917 ^ n3177 ^ 1'b0 ;
  assign n12187 = n5180 ^ n2294 ^ 1'b0 ;
  assign n12188 = n2774 | n10861 ;
  assign n12189 = n963 & n1298 ;
  assign n12190 = n7585 ^ n3100 ^ 1'b0 ;
  assign n12191 = n2686 & ~n12190 ;
  assign n12192 = n12190 & n12191 ;
  assign n12193 = n3603 | n9539 ;
  assign n12194 = n963 | n1023 ;
  assign n12195 = ( n1072 & n12193 ) | ( n1072 & n12194 ) | ( n12193 & n12194 ) ;
  assign n12196 = n5237 ^ n1879 ^ n172 ;
  assign n12197 = n12196 ^ n3067 ^ 1'b0 ;
  assign n12198 = n374 | n12197 ;
  assign n12199 = n1158 & ~n3338 ;
  assign n12200 = n167 & ~n4407 ;
  assign n12201 = ~n11323 & n12200 ;
  assign n12202 = n9959 & n12201 ;
  assign n12203 = n12199 & n12202 ;
  assign n12204 = n1346 ^ n161 ^ 1'b0 ;
  assign n12205 = n4866 & n12204 ;
  assign n12206 = n12205 ^ n4028 ^ 1'b0 ;
  assign n12207 = n5785 ^ n3614 ^ 1'b0 ;
  assign n12208 = n12206 | n12207 ;
  assign n12209 = n12208 ^ n468 ^ 1'b0 ;
  assign n12210 = n2101 & n5625 ;
  assign n12211 = n3407 ^ n1860 ^ 1'b0 ;
  assign n12212 = ~n3138 & n12211 ;
  assign n12213 = ~n361 & n3037 ;
  assign n12214 = n12213 ^ n8922 ^ 1'b0 ;
  assign n12215 = n2887 ^ n976 ^ 1'b0 ;
  assign n12216 = n1134 & n12215 ;
  assign n12217 = n7698 & n12216 ;
  assign n12218 = n12217 ^ x0 ^ 1'b0 ;
  assign n12223 = n8953 ^ n2065 ^ 1'b0 ;
  assign n12219 = n4801 ^ n366 ^ 1'b0 ;
  assign n12220 = n754 & n12219 ;
  assign n12221 = n9585 & n9752 ;
  assign n12222 = ~n12220 & n12221 ;
  assign n12224 = n12223 ^ n12222 ^ 1'b0 ;
  assign n12225 = n11127 ^ n2725 ^ 1'b0 ;
  assign n12226 = n5554 & ~n8515 ;
  assign n12227 = ~n2360 & n12226 ;
  assign n12231 = ~n322 & n8643 ;
  assign n12228 = ~n7380 & n9763 ;
  assign n12229 = n760 | n1139 ;
  assign n12230 = n12228 | n12229 ;
  assign n12232 = n12231 ^ n12230 ^ 1'b0 ;
  assign n12233 = n177 | n1266 ;
  assign n12234 = n3009 | n12233 ;
  assign n12235 = n7541 ^ n70 ^ 1'b0 ;
  assign n12236 = n12234 & n12235 ;
  assign n12237 = ~n5053 & n12236 ;
  assign n12238 = n692 | n4704 ;
  assign n12239 = n4045 & ~n7720 ;
  assign n12240 = n11085 ^ n468 ^ 1'b0 ;
  assign n12241 = n9551 ^ n654 ^ 1'b0 ;
  assign n12242 = n722 | n7865 ;
  assign n12243 = n6120 ^ n2619 ^ 1'b0 ;
  assign n12244 = n4349 | n12243 ;
  assign n12245 = n12244 ^ n4197 ^ 1'b0 ;
  assign n12246 = n1491 & ~n1828 ;
  assign n12247 = n8514 & ~n12246 ;
  assign n12248 = ~n1439 & n12247 ;
  assign n12249 = ~n2784 & n4942 ;
  assign n12250 = ~n4580 & n12249 ;
  assign n12251 = n12250 ^ n423 ^ 1'b0 ;
  assign n12252 = ~n102 & n8838 ;
  assign n12253 = n12252 ^ n7112 ^ 1'b0 ;
  assign n12254 = ~n8737 & n11932 ;
  assign n12255 = ~n4722 & n6655 ;
  assign n12256 = n6003 & ~n7465 ;
  assign n12257 = ~n12255 & n12256 ;
  assign n12258 = n3333 & n7507 ;
  assign n12259 = n700 & n12258 ;
  assign n12260 = n258 | n9799 ;
  assign n12261 = n5330 & ~n12260 ;
  assign n12262 = n114 ^ n68 ^ 1'b0 ;
  assign n12263 = ( n142 & n1456 ) | ( n142 & ~n12262 ) | ( n1456 & ~n12262 ) ;
  assign n12264 = n4825 ^ n2334 ^ 1'b0 ;
  assign n12265 = n2193 & ~n4805 ;
  assign n12266 = n2435 & ~n10981 ;
  assign n12267 = ~n2761 & n11972 ;
  assign n12268 = n12267 ^ n7119 ^ 1'b0 ;
  assign n12269 = n1600 | n5942 ;
  assign n12270 = n892 & ~n1789 ;
  assign n12271 = n12270 ^ n1234 ^ 1'b0 ;
  assign n12272 = n553 | n12271 ;
  assign n12273 = n12272 ^ n10288 ^ n4917 ;
  assign n12274 = n3940 ^ n2477 ^ 1'b0 ;
  assign n12275 = ~n456 & n2142 ;
  assign n12276 = n5439 & n12275 ;
  assign n12277 = n2278 & ~n3798 ;
  assign n12278 = n200 & ~n12277 ;
  assign n12279 = n8804 ^ n1234 ^ 1'b0 ;
  assign n12280 = n12279 ^ n8742 ^ 1'b0 ;
  assign n12281 = n5793 & ~n7333 ;
  assign n12282 = n161 & ~n12281 ;
  assign n12283 = n3965 & n12282 ;
  assign n12284 = n10490 ^ n37 ^ 1'b0 ;
  assign n12285 = n10419 ^ n53 ^ 1'b0 ;
  assign n12286 = n3559 | n12285 ;
  assign n12287 = n7773 ^ n4471 ^ 1'b0 ;
  assign n12288 = ~n364 & n12287 ;
  assign n12289 = ~n1358 & n4742 ;
  assign n12291 = n553 & n1601 ;
  assign n12290 = n782 & n6106 ;
  assign n12292 = n12291 ^ n12290 ^ 1'b0 ;
  assign n12293 = n3968 ^ n743 ^ 1'b0 ;
  assign n12294 = x11 & n12293 ;
  assign n12295 = n12292 & n12294 ;
  assign n12296 = n4778 ^ n741 ^ 1'b0 ;
  assign n12297 = n9695 | n12296 ;
  assign n12298 = n12297 ^ n5894 ^ 1'b0 ;
  assign n12299 = n1730 | n5078 ;
  assign n12300 = n12299 ^ n2148 ^ 1'b0 ;
  assign n12301 = n12300 ^ n10879 ^ 1'b0 ;
  assign n12302 = n7773 & ~n12301 ;
  assign n12303 = n6897 | n7288 ;
  assign n12304 = n4882 & n7948 ;
  assign n12305 = n12304 ^ n205 ^ 1'b0 ;
  assign n12306 = n440 | n12305 ;
  assign n12307 = n1783 ^ n866 ^ 1'b0 ;
  assign n12308 = n2591 | n12307 ;
  assign n12309 = n5083 & ~n6348 ;
  assign n12310 = n12309 ^ n1918 ^ 1'b0 ;
  assign n12311 = n2435 ^ n364 ^ 1'b0 ;
  assign n12312 = n1559 | n12311 ;
  assign n12313 = n7666 ^ n5202 ^ 1'b0 ;
  assign n12314 = ~n1638 & n2060 ;
  assign n12315 = ~n4115 & n12314 ;
  assign n12316 = n4331 & n8790 ;
  assign n12317 = ~n12315 & n12316 ;
  assign n12318 = n5356 & n8921 ;
  assign n12319 = n5275 ^ n164 ^ 1'b0 ;
  assign n12320 = n3642 | n12319 ;
  assign n12323 = n2930 ^ n161 ^ 1'b0 ;
  assign n12324 = n2146 & n12323 ;
  assign n12321 = ~n3554 & n8021 ;
  assign n12322 = ( n5990 & n7083 ) | ( n5990 & ~n12321 ) | ( n7083 & ~n12321 ) ;
  assign n12325 = n12324 ^ n12322 ^ 1'b0 ;
  assign n12326 = n12325 ^ n7579 ^ 1'b0 ;
  assign n12327 = n12320 | n12326 ;
  assign n12328 = ~n4367 & n11125 ;
  assign n12329 = n1476 & ~n4358 ;
  assign n12330 = n2160 & ~n3692 ;
  assign n12331 = n12330 ^ n703 ^ 1'b0 ;
  assign n12332 = n12331 ^ n9978 ^ 1'b0 ;
  assign n12333 = n12329 & n12332 ;
  assign n12334 = n5397 ^ n506 ^ 1'b0 ;
  assign n12335 = ~n1229 & n12334 ;
  assign n12336 = n12335 ^ n10014 ^ 1'b0 ;
  assign n12342 = n908 & n3954 ;
  assign n12343 = n5930 & n12342 ;
  assign n12337 = ~n3080 & n3304 ;
  assign n12338 = n5440 & ~n7081 ;
  assign n12339 = n5701 & n12338 ;
  assign n12340 = n12337 & ~n12339 ;
  assign n12341 = ~n4383 & n12340 ;
  assign n12344 = n12343 ^ n12341 ^ 1'b0 ;
  assign n12345 = n12336 & n12344 ;
  assign n12346 = n988 ^ n432 ^ 1'b0 ;
  assign n12347 = n3141 & ~n12346 ;
  assign n12348 = n4347 & ~n7767 ;
  assign n12349 = n434 & n12348 ;
  assign n12350 = n512 | n8057 ;
  assign n12351 = n9994 ^ n3781 ^ 1'b0 ;
  assign n12352 = n1109 | n10429 ;
  assign n12353 = n12351 & ~n12352 ;
  assign n12354 = n1220 & n4436 ;
  assign n12355 = n75 | n12354 ;
  assign n12356 = n12355 ^ n6107 ^ 1'b0 ;
  assign n12357 = n4927 | n12356 ;
  assign n12358 = ~n1827 & n7907 ;
  assign n12359 = n3732 & n12358 ;
  assign n12360 = n12359 ^ n1158 ^ 1'b0 ;
  assign n12361 = n293 & n4700 ;
  assign n12362 = n4206 | n9337 ;
  assign n12363 = n343 & n12157 ;
  assign n12364 = n5257 ^ n4807 ^ 1'b0 ;
  assign n12365 = n4633 ^ n2395 ^ 1'b0 ;
  assign n12366 = n11846 & n12365 ;
  assign n12367 = n5359 & n5646 ;
  assign n12368 = n12366 & n12367 ;
  assign n12369 = n11711 ^ n3314 ^ 1'b0 ;
  assign n12370 = ~n10644 & n12369 ;
  assign n12371 = n3164 ^ n545 ^ 1'b0 ;
  assign n12372 = n12371 ^ n715 ^ 1'b0 ;
  assign n12373 = n269 & ~n12372 ;
  assign n12374 = n2112 & ~n12373 ;
  assign n12375 = ~n246 & n11673 ;
  assign n12376 = n12375 ^ n2539 ^ 1'b0 ;
  assign n12377 = n448 & n5045 ;
  assign n12378 = n4212 & n12377 ;
  assign n12379 = ~n8948 & n11622 ;
  assign n12380 = n1390 & ~n5070 ;
  assign n12381 = ~n185 & n12380 ;
  assign n12382 = n7486 ^ n239 ^ 1'b0 ;
  assign n12383 = n10676 ^ n7079 ^ 1'b0 ;
  assign n12384 = n3897 & ~n8711 ;
  assign n12385 = ~n5228 & n12384 ;
  assign n12386 = n4339 ^ n832 ^ 1'b0 ;
  assign n12387 = n1077 & n3761 ;
  assign n12388 = ~n461 & n7596 ;
  assign n12389 = n94 | n2549 ;
  assign n12390 = n12389 ^ n805 ^ 1'b0 ;
  assign n12391 = n7258 ^ n4026 ^ 1'b0 ;
  assign n12392 = n489 & n6544 ;
  assign n12393 = n12392 ^ n1219 ^ 1'b0 ;
  assign n12394 = n4790 ^ x9 ^ 1'b0 ;
  assign n12395 = n5359 | n12394 ;
  assign n12396 = n7190 & ~n8312 ;
  assign n12397 = n2535 & ~n10098 ;
  assign n12398 = n12397 ^ n113 ^ 1'b0 ;
  assign n12399 = n1898 & ~n4155 ;
  assign n12400 = n11843 ^ n8819 ^ 1'b0 ;
  assign n12401 = n8341 ^ n1162 ^ 1'b0 ;
  assign n12402 = n79 & n6571 ;
  assign n12403 = n1192 | n12402 ;
  assign n12404 = n12403 ^ n11787 ^ 1'b0 ;
  assign n12405 = n5741 ^ n1768 ^ 1'b0 ;
  assign n12406 = n9058 & ~n12405 ;
  assign n12407 = n519 | n6353 ;
  assign n12408 = n4594 & ~n6065 ;
  assign n12409 = n12407 & n12408 ;
  assign n12410 = n2898 | n5217 ;
  assign n12411 = n12409 & ~n12410 ;
  assign n12412 = ~n3671 & n12184 ;
  assign n12413 = n185 | n7227 ;
  assign n12414 = n12413 ^ n4008 ^ 1'b0 ;
  assign n12415 = n498 ^ n392 ^ 1'b0 ;
  assign n12416 = n12415 ^ n7634 ^ 1'b0 ;
  assign n12417 = n11929 ^ n3097 ^ 1'b0 ;
  assign n12418 = n2770 ^ n2707 ^ 1'b0 ;
  assign n12419 = n12418 ^ n7924 ^ 1'b0 ;
  assign n12420 = n2681 | n8392 ;
  assign n12421 = n2642 | n3894 ;
  assign n12422 = n476 & ~n4749 ;
  assign n12423 = ~n1082 & n12422 ;
  assign n12424 = n12423 ^ n11253 ^ 1'b0 ;
  assign n12425 = n7023 & n11940 ;
  assign n12426 = ~n4827 & n12165 ;
  assign n12427 = n12426 ^ n5326 ^ 1'b0 ;
  assign n12428 = ~n3672 & n6222 ;
  assign n12429 = n6015 | n8001 ;
  assign n12430 = n2560 ^ n2556 ^ 1'b0 ;
  assign n12431 = n2664 | n12430 ;
  assign n12432 = n12431 ^ n3916 ^ 1'b0 ;
  assign n12433 = n12432 ^ n9397 ^ 1'b0 ;
  assign n12434 = n2573 & n3484 ;
  assign n12435 = ~n2046 & n12434 ;
  assign n12436 = n12435 ^ n5232 ^ 1'b0 ;
  assign n12437 = n12237 ^ n7687 ^ 1'b0 ;
  assign n12438 = n532 | n12437 ;
  assign n12439 = ~n1360 & n4765 ;
  assign n12440 = n4088 & n12439 ;
  assign n12441 = n5128 | n12440 ;
  assign n12442 = n1958 ^ n592 ^ 1'b0 ;
  assign n12443 = n119 | n2258 ;
  assign n12444 = n10495 | n12443 ;
  assign n12445 = n7753 ^ n6341 ^ n3247 ;
  assign n12447 = n2611 ^ n2521 ^ 1'b0 ;
  assign n12448 = n2432 & ~n12447 ;
  assign n12449 = n12448 ^ n5286 ^ 1'b0 ;
  assign n12450 = n2762 & n12449 ;
  assign n12446 = ( n3271 & n3636 ) | ( n3271 & ~n7310 ) | ( n3636 & ~n7310 ) ;
  assign n12451 = n12450 ^ n12446 ^ 1'b0 ;
  assign n12452 = n12445 & n12451 ;
  assign n12453 = n3243 ^ n2779 ^ 1'b0 ;
  assign n12454 = n12453 ^ n4916 ^ n1543 ;
  assign n12455 = n92 & n12454 ;
  assign n12456 = n6171 ^ n4763 ^ 1'b0 ;
  assign n12457 = n12455 | n12456 ;
  assign n12458 = n12457 ^ n5704 ^ 1'b0 ;
  assign n12461 = n3738 ^ n2252 ^ 1'b0 ;
  assign n12459 = n1771 ^ n354 ^ 1'b0 ;
  assign n12460 = n9792 | n12459 ;
  assign n12462 = n12461 ^ n12460 ^ 1'b0 ;
  assign n12465 = ~n198 & n963 ;
  assign n12466 = n12465 ^ n9733 ^ 1'b0 ;
  assign n12463 = ~n2344 & n6185 ;
  assign n12464 = ~n1538 & n12463 ;
  assign n12467 = n12466 ^ n12464 ^ 1'b0 ;
  assign n12468 = n10124 ^ n10025 ^ n60 ;
  assign n12469 = n55 & ~n4420 ;
  assign n12470 = ~n12468 & n12469 ;
  assign n12471 = n2813 & ~n6325 ;
  assign n12472 = n9480 & n12471 ;
  assign n12473 = n295 | n3957 ;
  assign n12474 = n12473 ^ n8973 ^ 1'b0 ;
  assign n12475 = ~n12472 & n12474 ;
  assign n12476 = n6185 & ~n6479 ;
  assign n12477 = n12476 ^ n7577 ^ 1'b0 ;
  assign n12478 = n4474 ^ n286 ^ 1'b0 ;
  assign n12479 = n11722 | n12478 ;
  assign n12480 = n3156 ^ n1791 ^ 1'b0 ;
  assign n12481 = ~n12479 & n12480 ;
  assign n12482 = n1552 & n1656 ;
  assign n12483 = n10081 | n12482 ;
  assign n12484 = n9750 | n12483 ;
  assign n12485 = ~n4536 & n10160 ;
  assign n12486 = ~n11481 & n12485 ;
  assign n12487 = ~n3036 & n12486 ;
  assign n12488 = n1110 & ~n6607 ;
  assign n12489 = n12222 ^ n5753 ^ 1'b0 ;
  assign n12490 = n3866 & ~n5269 ;
  assign n12491 = n12490 ^ n6171 ^ 1'b0 ;
  assign n12492 = n7753 | n12491 ;
  assign n12493 = n47 & n12492 ;
  assign n12494 = n12493 ^ n1917 ^ 1'b0 ;
  assign n12495 = n12494 ^ n9186 ^ 1'b0 ;
  assign n12496 = n3594 ^ n1806 ^ 1'b0 ;
  assign n12497 = ~n348 & n12496 ;
  assign n12498 = n965 & ~n5201 ;
  assign n12499 = n12498 ^ n1739 ^ 1'b0 ;
  assign n12500 = n6990 & n12499 ;
  assign n12501 = n1688 ^ n1497 ^ 1'b0 ;
  assign n12502 = n7874 | n12501 ;
  assign n12503 = n2264 & ~n11944 ;
  assign n12504 = n4082 & n7432 ;
  assign n12505 = n5322 & ~n12504 ;
  assign n12506 = n1134 & n5764 ;
  assign n12507 = n12506 ^ n5032 ^ 1'b0 ;
  assign n12508 = n3028 & ~n10098 ;
  assign n12509 = n12508 ^ n3333 ^ 1'b0 ;
  assign n12510 = n9846 ^ n9549 ^ 1'b0 ;
  assign n12511 = n12509 & n12510 ;
  assign n12512 = n9535 | n12511 ;
  assign n12513 = n8341 ^ n6587 ^ n687 ;
  assign n12514 = n1668 & ~n4548 ;
  assign n12515 = n9752 ^ n241 ^ 1'b0 ;
  assign n12516 = n8590 & ~n12515 ;
  assign n12517 = n12514 & n12516 ;
  assign n12518 = n1632 & n2210 ;
  assign n12519 = n1455 ^ n645 ^ 1'b0 ;
  assign n12520 = n12519 ^ n3803 ^ 1'b0 ;
  assign n12521 = n419 & ~n12520 ;
  assign n12525 = n7388 ^ n2689 ^ n1713 ;
  assign n12522 = n9695 ^ n6188 ^ 1'b0 ;
  assign n12523 = ~n1106 & n3940 ;
  assign n12524 = n12522 & ~n12523 ;
  assign n12526 = n12525 ^ n12524 ^ 1'b0 ;
  assign n12527 = n2428 | n2443 ;
  assign n12528 = n3249 ^ n1089 ^ 1'b0 ;
  assign n12529 = n3552 & ~n12528 ;
  assign n12530 = n3449 & ~n12529 ;
  assign n12531 = n8108 | n11870 ;
  assign n12532 = n10902 & ~n12531 ;
  assign n12533 = n9857 | n10384 ;
  assign n12534 = ~n403 & n10954 ;
  assign n12535 = n10479 ^ n5806 ^ 1'b0 ;
  assign n12536 = n9060 | n12535 ;
  assign n12537 = n2942 | n12536 ;
  assign n12538 = ~n576 & n6721 ;
  assign n12539 = ~n4760 & n12538 ;
  assign n12540 = n5085 ^ n354 ^ 1'b0 ;
  assign n12541 = n12540 ^ n9860 ^ 1'b0 ;
  assign n12544 = n1431 & n3451 ;
  assign n12545 = n1672 ^ n121 ^ 1'b0 ;
  assign n12546 = n12544 & ~n12545 ;
  assign n12542 = ~n627 & n4510 ;
  assign n12543 = ~n4334 & n12542 ;
  assign n12547 = n12546 ^ n12543 ^ 1'b0 ;
  assign n12549 = ~n792 & n4589 ;
  assign n12550 = n12549 ^ n1316 ^ 1'b0 ;
  assign n12551 = ~n4018 & n6726 ;
  assign n12552 = n12550 & n12551 ;
  assign n12548 = n1718 | n7380 ;
  assign n12553 = n12552 ^ n12548 ^ 1'b0 ;
  assign n12554 = ~n1824 & n5206 ;
  assign n12555 = n12554 ^ n2342 ^ 1'b0 ;
  assign n12559 = n2027 & ~n3392 ;
  assign n12560 = ~n2611 & n12559 ;
  assign n12561 = n83 & n12560 ;
  assign n12556 = n96 & ~n8363 ;
  assign n12557 = n12556 ^ n1934 ^ 1'b0 ;
  assign n12558 = n4042 & ~n12557 ;
  assign n12562 = n12561 ^ n12558 ^ 1'b0 ;
  assign n12563 = n6725 & ~n7811 ;
  assign n12564 = n3810 & ~n3972 ;
  assign n12565 = n7487 | n9915 ;
  assign n12566 = ~n12564 & n12565 ;
  assign n12567 = n46 & ~n75 ;
  assign n12568 = ~n46 & n12567 ;
  assign n12569 = n253 & n3061 ;
  assign n12570 = ~n3061 & n12569 ;
  assign n12571 = n12570 ^ n191 ^ 1'b0 ;
  assign n12572 = n72 & ~n12571 ;
  assign n12573 = n12568 & n12572 ;
  assign n12574 = n2654 | n12573 ;
  assign n12575 = n12573 & ~n12574 ;
  assign n12576 = ~n6950 & n12575 ;
  assign n12577 = n1129 | n12576 ;
  assign n12578 = n1129 & ~n12577 ;
  assign n12579 = x11 & n107 ;
  assign n12580 = ~x11 & n12579 ;
  assign n12581 = x0 & ~n100 ;
  assign n12582 = ~x0 & n12581 ;
  assign n12583 = x6 & n12582 ;
  assign n12584 = ~n12582 & n12583 ;
  assign n12585 = ~n16 & n12584 ;
  assign n12586 = n34 ^ n14 ^ 1'b0 ;
  assign n12587 = n107 & ~n12586 ;
  assign n12588 = n12587 ^ n55 ^ 1'b0 ;
  assign n12589 = n12585 & ~n12588 ;
  assign n12590 = n36 & n12589 ;
  assign n12591 = n12580 & n12590 ;
  assign n12592 = ~n148 & n456 ;
  assign n12593 = n12591 & n12592 ;
  assign n12594 = n12578 | n12593 ;
  assign n12595 = n12578 & ~n12594 ;
  assign n12596 = n438 & n1716 ;
  assign n12597 = ~n438 & n12596 ;
  assign n12598 = n562 | n12597 ;
  assign n12599 = n562 & ~n12598 ;
  assign n12600 = n12599 ^ n273 ^ 1'b0 ;
  assign n12601 = ~n17 & n37 ;
  assign n12602 = n17 & n12601 ;
  assign n12603 = n55 & ~n12602 ;
  assign n12604 = n12587 & ~n12603 ;
  assign n12605 = ~n12587 & n12604 ;
  assign n12606 = n922 & n12605 ;
  assign n12607 = n7120 & ~n12606 ;
  assign n12608 = n12606 & n12607 ;
  assign n12609 = n25 | n79 ;
  assign n12610 = n25 & ~n12609 ;
  assign n12611 = n848 & ~n12610 ;
  assign n12612 = ~n848 & n12611 ;
  assign n12613 = n678 | n12612 ;
  assign n12614 = n12612 & ~n12613 ;
  assign n12615 = n12608 | n12614 ;
  assign n12616 = n12608 & ~n12615 ;
  assign n12617 = n12600 | n12616 ;
  assign n12618 = n12595 & ~n12617 ;
  assign n12619 = ~n37 & n153 ;
  assign n12620 = ~n153 & n12619 ;
  assign n12621 = n2041 & ~n12620 ;
  assign n12622 = ~n2041 & n12621 ;
  assign n12623 = n8116 & ~n12622 ;
  assign n12624 = n12622 & n12623 ;
  assign n12625 = n1225 | n12624 ;
  assign n12626 = n12618 & ~n12625 ;
  assign n12627 = n4533 ^ n1908 ^ 1'b0 ;
  assign n12628 = n4264 & n12627 ;
  assign n12629 = n7264 & n12628 ;
  assign n12630 = n4285 ^ n257 ^ 1'b0 ;
  assign n12631 = n3088 ^ n1807 ^ 1'b0 ;
  assign n12632 = ~n4706 & n12631 ;
  assign n12635 = n252 | n6979 ;
  assign n12636 = n2639 & ~n12635 ;
  assign n12633 = ( n980 & n1718 ) | ( n980 & n3576 ) | ( n1718 & n3576 ) ;
  assign n12634 = n1718 | n12633 ;
  assign n12637 = n12636 ^ n12634 ^ 1'b0 ;
  assign n12638 = n1304 & n4479 ;
  assign n12639 = n7155 & n12638 ;
  assign n12640 = n513 & n823 ;
  assign n12641 = n12640 ^ n10984 ^ 1'b0 ;
  assign n12642 = n7048 ^ n4790 ^ 1'b0 ;
  assign n12643 = ~n241 & n4805 ;
  assign n12644 = n7697 & n12643 ;
  assign n12645 = ~n37 & n12644 ;
  assign n12646 = n754 | n5053 ;
  assign n12647 = n7096 ^ n4180 ^ 1'b0 ;
  assign n12648 = ~n1306 & n12647 ;
  assign n12649 = n12648 ^ n3503 ^ 1'b0 ;
  assign n12650 = n12646 & n12649 ;
  assign n12651 = ~n12489 & n12650 ;
  assign n12652 = n2130 ^ x8 ^ 1'b0 ;
  assign n12653 = n2506 & n10736 ;
  assign n12654 = n12653 ^ n8056 ^ 1'b0 ;
  assign n12655 = n3991 & ~n12654 ;
  assign n12656 = n4374 ^ n263 ^ 1'b0 ;
  assign n12657 = ~n745 & n2012 ;
  assign n12658 = n278 & n9335 ;
  assign n12659 = n2477 | n12658 ;
  assign n12660 = n5078 | n12659 ;
  assign n12663 = n3135 ^ n3074 ^ 1'b0 ;
  assign n12661 = n689 | n743 ;
  assign n12662 = n11397 | n12661 ;
  assign n12664 = n12663 ^ n12662 ^ 1'b0 ;
  assign n12665 = n1125 & n8392 ;
  assign n12666 = n9607 ^ n3711 ^ 1'b0 ;
  assign n12667 = n6669 ^ n1403 ^ n1254 ;
  assign n12668 = n2607 & ~n8010 ;
  assign n12669 = n12525 & n12668 ;
  assign n12670 = n4756 & ~n12669 ;
  assign n12671 = n12670 ^ n6295 ^ 1'b0 ;
  assign n12672 = n1761 & n6412 ;
  assign n12677 = ~n4266 & n6867 ;
  assign n12673 = n5348 ^ n3537 ^ 1'b0 ;
  assign n12674 = n663 & n12673 ;
  assign n12675 = n12674 ^ n510 ^ 1'b0 ;
  assign n12676 = n1425 & n12675 ;
  assign n12678 = n12677 ^ n12676 ^ 1'b0 ;
  assign n12679 = ~n9641 & n10432 ;
  assign n12680 = n12679 ^ n9060 ^ 1'b0 ;
  assign n12681 = n3875 & ~n4543 ;
  assign n12682 = ~n1476 & n5461 ;
  assign n12683 = ~n8197 & n12682 ;
  assign n12684 = n4053 & n8770 ;
  assign n12685 = ~n1758 & n12684 ;
  assign n12686 = n12685 ^ n10873 ^ 1'b0 ;
  assign n12687 = ~n10079 & n12686 ;
  assign n12688 = n6360 ^ n6040 ^ 1'b0 ;
  assign n12689 = n1886 | n12688 ;
  assign n12690 = n159 & n697 ;
  assign n12691 = n2483 & n11373 ;
  assign n12692 = n7707 & ~n12691 ;
  assign n12693 = n2380 & n4964 ;
  assign n12694 = ~n3807 & n12693 ;
  assign n12695 = n2553 | n9957 ;
  assign n12696 = n12694 & ~n12695 ;
  assign n12697 = n7884 | n9029 ;
  assign n12698 = ~n8120 & n12697 ;
  assign n12699 = n9643 ^ n6472 ^ 1'b0 ;
  assign n12700 = n2898 ^ n785 ^ 1'b0 ;
  assign n12701 = ~n11301 & n12700 ;
  assign n12702 = ~n4024 & n12701 ;
  assign n12703 = n12702 ^ n1492 ^ n250 ;
  assign n12704 = n1929 ^ n634 ^ 1'b0 ;
  assign n12705 = n12042 & n12704 ;
  assign n12707 = ~n1195 & n3882 ;
  assign n12708 = n2260 & n12707 ;
  assign n12709 = n12708 ^ n10636 ^ 1'b0 ;
  assign n12706 = n847 | n3282 ;
  assign n12710 = n12709 ^ n12706 ^ 1'b0 ;
  assign n12711 = n1019 | n9321 ;
  assign n12712 = ~n60 & n2303 ;
  assign n12713 = n12712 ^ n2932 ^ 1'b0 ;
  assign n12714 = ~n9240 & n10313 ;
  assign n12715 = n12277 ^ n4751 ^ 1'b0 ;
  assign n12716 = ~n7656 & n12715 ;
  assign n12717 = n8693 | n12716 ;
  assign n12718 = n2604 & ~n7542 ;
  assign n12719 = ~n10024 & n12718 ;
  assign n12720 = n1737 | n8918 ;
  assign n12721 = n2092 & ~n3127 ;
  assign n12722 = n1822 & ~n12721 ;
  assign n12728 = n7868 ^ n2572 ^ 1'b0 ;
  assign n12729 = ~n567 & n12728 ;
  assign n12730 = n12729 ^ n6346 ^ 1'b0 ;
  assign n12727 = n1348 | n2576 ;
  assign n12731 = n12730 ^ n12727 ^ 1'b0 ;
  assign n12732 = n5270 ^ n1322 ^ 1'b0 ;
  assign n12733 = ~n12731 & n12732 ;
  assign n12734 = ~n1441 & n12733 ;
  assign n12735 = n356 & ~n9581 ;
  assign n12736 = n12734 & n12735 ;
  assign n12723 = n4746 ^ n2481 ^ 1'b0 ;
  assign n12724 = n1577 ^ n1185 ^ 1'b0 ;
  assign n12725 = ~n4267 & n12724 ;
  assign n12726 = n12723 & n12725 ;
  assign n12737 = n12736 ^ n12726 ^ 1'b0 ;
  assign n12738 = n12722 | n12737 ;
  assign n12739 = n1479 ^ n645 ^ 1'b0 ;
  assign n12740 = n2181 & n12739 ;
  assign n12741 = ~n58 & n12740 ;
  assign n12742 = n5686 ^ n4336 ^ 1'b0 ;
  assign n12743 = n5941 & n12742 ;
  assign n12744 = n12743 ^ n7792 ^ 1'b0 ;
  assign n12745 = n12741 & ~n12744 ;
  assign n12746 = n9010 & n12745 ;
  assign n12747 = n94 & n4292 ;
  assign n12748 = ~n4591 & n10659 ;
  assign n12749 = ~n12747 & n12748 ;
  assign n12750 = n4081 ^ n263 ^ 1'b0 ;
  assign n12751 = n6695 | n12750 ;
  assign n12752 = n12751 ^ n2270 ^ 1'b0 ;
  assign n12753 = n3219 ^ n2150 ^ 1'b0 ;
  assign n12754 = ~n9176 & n12753 ;
  assign n12755 = n8644 | n12065 ;
  assign n12756 = n12755 ^ n5857 ^ 1'b0 ;
  assign n12757 = ~n8104 & n11691 ;
  assign n12758 = n3217 & n7112 ;
  assign n12759 = n6065 ^ n3189 ^ 1'b0 ;
  assign n12760 = n10920 & n12759 ;
  assign n12761 = n3138 ^ n1599 ^ 1'b0 ;
  assign n12762 = n954 & ~n1555 ;
  assign n12763 = ~n12761 & n12762 ;
  assign n12765 = n83 | n4061 ;
  assign n12766 = n12765 ^ n1372 ^ 1'b0 ;
  assign n12764 = n958 & n1129 ;
  assign n12767 = n12766 ^ n12764 ^ 1'b0 ;
  assign n12768 = n128 | n12767 ;
  assign n12769 = n10589 | n12768 ;
  assign n12770 = n12769 ^ n4499 ^ 1'b0 ;
  assign n12771 = n3643 ^ n806 ^ 1'b0 ;
  assign n12772 = ~n7798 & n12771 ;
  assign n12773 = n4421 ^ n92 ^ 1'b0 ;
  assign n12774 = ~n299 & n12448 ;
  assign n12775 = n12774 ^ n1407 ^ 1'b0 ;
  assign n12776 = n11542 & n12775 ;
  assign n12777 = n1959 | n4346 ;
  assign n12778 = n159 & n12777 ;
  assign n12779 = n12778 ^ n458 ^ 1'b0 ;
  assign n12780 = n1479 | n8133 ;
  assign n12781 = n12780 ^ n9342 ^ 1'b0 ;
  assign n12782 = n6995 & ~n12781 ;
  assign n12783 = ~n3265 & n12782 ;
  assign n12784 = n12783 ^ n7917 ^ 1'b0 ;
  assign n12785 = ~n3569 & n9217 ;
  assign n12786 = n12777 ^ n12000 ^ 1'b0 ;
  assign n12787 = n10651 & n12786 ;
  assign n12788 = ~n1239 & n1245 ;
  assign n12789 = ~n5964 & n12788 ;
  assign n12790 = n12789 ^ n310 ^ 1'b0 ;
  assign n12791 = n8112 | n12790 ;
  assign n12792 = n133 | n1622 ;
  assign n12793 = n15 | n12792 ;
  assign n12794 = n3643 & n12793 ;
  assign n12795 = ~n6913 & n12794 ;
  assign n12796 = n7265 ^ n148 ^ 1'b0 ;
  assign n12797 = n11696 & n12796 ;
  assign n12798 = n5260 | n6081 ;
  assign n12799 = n2757 & ~n12798 ;
  assign n12800 = ~n3844 & n12799 ;
  assign n12801 = ~n8248 & n10147 ;
  assign n12802 = n12801 ^ n6933 ^ 1'b0 ;
  assign n12803 = n7503 | n12802 ;
  assign n12804 = n540 | n702 ;
  assign n12805 = ~n1936 & n7461 ;
  assign n12806 = ~n2261 & n12805 ;
  assign n12807 = n12804 | n12806 ;
  assign n12808 = n9806 | n10273 ;
  assign n12809 = n3452 & n10472 ;
  assign n12810 = ~n7418 & n12809 ;
  assign n12811 = n149 & n4822 ;
  assign n12824 = n2937 ^ n1965 ^ 1'b0 ;
  assign n12825 = n9459 & ~n12824 ;
  assign n12820 = ~n1117 & n5567 ;
  assign n12821 = ~n5567 & n12820 ;
  assign n12822 = ~n3156 & n12821 ;
  assign n12823 = n12822 ^ n5241 ^ 1'b0 ;
  assign n12826 = n12825 ^ n12823 ^ 1'b0 ;
  assign n12812 = n157 & ~n759 ;
  assign n12813 = n3423 & ~n4407 ;
  assign n12814 = ~n3423 & n12813 ;
  assign n12815 = n12814 ^ n1771 ^ 1'b0 ;
  assign n12816 = n12812 & ~n12815 ;
  assign n12817 = n4842 | n8967 ;
  assign n12818 = n12816 & ~n12817 ;
  assign n12819 = ~n12816 & n12818 ;
  assign n12827 = n12826 ^ n12819 ^ 1'b0 ;
  assign n12828 = ~n86 & n187 ;
  assign n12829 = n86 & n12828 ;
  assign n12830 = n1048 | n2736 ;
  assign n12831 = n2736 & ~n12830 ;
  assign n12832 = n1388 & ~n12831 ;
  assign n12833 = n12829 | n12832 ;
  assign n12834 = n12829 & ~n12833 ;
  assign n12835 = n291 & ~n3116 ;
  assign n12836 = ~n291 & n12835 ;
  assign n12837 = ~n55 & n191 ;
  assign n12838 = ~n191 & n12837 ;
  assign n12839 = n168 & n12838 ;
  assign n12840 = n55 | n12839 ;
  assign n12841 = n12839 & ~n12840 ;
  assign n12842 = n3087 | n12841 ;
  assign n12843 = n3087 & ~n12842 ;
  assign n12844 = ~n12836 & n12843 ;
  assign n12845 = ~n12834 & n12844 ;
  assign n12846 = n12834 & n12845 ;
  assign n12847 = n6230 | n9925 ;
  assign n12848 = n9925 & ~n12847 ;
  assign n12849 = n2707 & ~n12848 ;
  assign n12850 = n12846 & n12849 ;
  assign n12851 = n385 & ~n12850 ;
  assign n12852 = n12827 & n12851 ;
  assign n12853 = n7938 ^ n6230 ^ 1'b0 ;
  assign n12854 = n2176 & n5241 ;
  assign n12855 = n10392 ^ n2912 ^ 1'b0 ;
  assign n12856 = n8156 & ~n12855 ;
  assign n12862 = n609 & ~n6210 ;
  assign n12857 = n4812 ^ n495 ^ 1'b0 ;
  assign n12858 = n3080 | n12857 ;
  assign n12859 = n366 | n12858 ;
  assign n12860 = n12859 ^ n2891 ^ 1'b0 ;
  assign n12861 = n3210 & n12860 ;
  assign n12863 = n12862 ^ n12861 ^ 1'b0 ;
  assign n12864 = n2612 | n12376 ;
  assign n12865 = n12864 ^ n5685 ^ 1'b0 ;
  assign n12866 = n1161 & n6279 ;
  assign n12867 = n12866 ^ n5425 ^ n3431 ;
  assign n12868 = n1320 & ~n12867 ;
  assign n12871 = n11853 ^ n348 ^ 1'b0 ;
  assign n12869 = n3404 & n4761 ;
  assign n12870 = n12869 ^ n5789 ^ 1'b0 ;
  assign n12872 = n12871 ^ n12870 ^ 1'b0 ;
  assign n12873 = n1219 & n12872 ;
  assign n12876 = n5455 ^ n3024 ^ 1'b0 ;
  assign n12877 = ~n2138 & n12876 ;
  assign n12874 = n10639 ^ n721 ^ 1'b0 ;
  assign n12875 = ~n4443 & n12874 ;
  assign n12878 = n12877 ^ n12875 ^ 1'b0 ;
  assign n12879 = n8322 & n12878 ;
  assign n12880 = ~n1632 & n7949 ;
  assign n12881 = n10469 ^ n30 ^ 1'b0 ;
  assign n12882 = n952 ^ n654 ^ 1'b0 ;
  assign n12883 = n3154 & ~n12882 ;
  assign n12884 = n12883 ^ n2932 ^ 1'b0 ;
  assign n12885 = n12884 ^ n1483 ^ 1'b0 ;
  assign n12886 = n3693 | n12885 ;
  assign n12887 = n3240 ^ n653 ^ 1'b0 ;
  assign n12888 = ~n489 & n3655 ;
  assign n12889 = ~n2140 & n10207 ;
  assign n12890 = n12888 & ~n12889 ;
  assign n12891 = ~n6918 & n12890 ;
  assign n12892 = ~n3194 & n12891 ;
  assign n12893 = n1620 & ~n3820 ;
  assign n12894 = n1178 & n8326 ;
  assign n12895 = n12894 ^ n6713 ^ 1'b0 ;
  assign n12896 = n12895 ^ n1172 ^ 1'b0 ;
  assign n12897 = n9344 ^ n2642 ^ 1'b0 ;
  assign n12898 = ~n198 & n12897 ;
  assign n12899 = n7214 | n9832 ;
  assign n12900 = n2432 & n12899 ;
  assign n12901 = ~n12898 & n12900 ;
  assign n12902 = n2027 & n3229 ;
  assign n12903 = n3127 & n4348 ;
  assign n12904 = n12902 & n12903 ;
  assign n12905 = n297 & ~n5823 ;
  assign n12906 = n1441 & n12905 ;
  assign n12907 = n865 & n10652 ;
  assign n12908 = n10481 ^ n7581 ^ 1'b0 ;
  assign n12909 = n338 & n408 ;
  assign n12910 = n86 & n5253 ;
  assign n12911 = n7657 ^ n7344 ^ 1'b0 ;
  assign n12912 = n2843 | n12911 ;
  assign n12913 = n361 & ~n7746 ;
  assign n12914 = n12913 ^ n5788 ^ 1'b0 ;
  assign n12915 = n2013 & ~n12914 ;
  assign n12916 = n12915 ^ n11063 ^ 1'b0 ;
  assign n12917 = n2382 | n11328 ;
  assign n12918 = n9055 ^ n6346 ^ n3841 ;
  assign n12919 = n4216 | n8560 ;
  assign n12920 = n12919 ^ n715 ^ 1'b0 ;
  assign n12921 = n6515 ^ n55 ^ 1'b0 ;
  assign n12922 = n9677 & n12921 ;
  assign n12923 = n12920 & n12922 ;
  assign n12924 = n1722 & n12923 ;
  assign n12925 = n12924 ^ n5023 ^ 1'b0 ;
  assign n12926 = n4548 | n5946 ;
  assign n12927 = n79 & n3988 ;
  assign n12928 = n12295 & n12927 ;
  assign n12929 = ~n497 & n883 ;
  assign n12930 = n16 & n6689 ;
  assign n12931 = n7872 & n12930 ;
  assign n12932 = ~n1893 & n12931 ;
  assign n12933 = n12932 ^ n2060 ^ 1'b0 ;
  assign n12934 = ~n12929 & n12933 ;
  assign n12935 = n10950 ^ n351 ^ 1'b0 ;
  assign n12936 = ~n4844 & n9621 ;
  assign n12937 = n12936 ^ n3643 ^ 1'b0 ;
  assign n12938 = n12937 ^ n12866 ^ 1'b0 ;
  assign n12939 = n4105 & n12938 ;
  assign n12940 = n5647 ^ n4237 ^ n1174 ;
  assign n12941 = n2101 & n7050 ;
  assign n12942 = n1956 & n12941 ;
  assign n12943 = n11897 ^ n3459 ^ 1'b0 ;
  assign n12944 = n10994 | n12943 ;
  assign n12945 = n489 & ~n12740 ;
  assign n12946 = n12944 & n12945 ;
  assign n12947 = n4378 ^ n415 ^ 1'b0 ;
  assign n12948 = n3472 & ~n12947 ;
  assign n12949 = n12948 ^ n2789 ^ 1'b0 ;
  assign n12950 = n7731 | n12949 ;
  assign n12952 = n2932 ^ n1222 ^ 1'b0 ;
  assign n12953 = n12952 ^ n3567 ^ 1'b0 ;
  assign n12954 = n5234 | n12953 ;
  assign n12951 = n700 & n8479 ;
  assign n12955 = n12954 ^ n12951 ^ n1479 ;
  assign n12957 = n6286 ^ n3402 ^ 1'b0 ;
  assign n12958 = n4024 | n12957 ;
  assign n12956 = n616 & n1381 ;
  assign n12959 = n12958 ^ n12956 ^ 1'b0 ;
  assign n12960 = n7942 & n12959 ;
  assign n12961 = n6933 & n12960 ;
  assign n12962 = ~n1033 & n6450 ;
  assign n12963 = n2844 & ~n12962 ;
  assign n12964 = n12215 ^ n2761 ^ n2055 ;
  assign n12965 = n9393 ^ n2967 ^ 1'b0 ;
  assign n12966 = n1956 | n12965 ;
  assign n12967 = n10719 ^ n9655 ^ n4246 ;
  assign n12968 = n2623 ^ n1695 ^ 1'b0 ;
  assign n12969 = n12968 ^ n11831 ^ 1'b0 ;
  assign n12971 = n364 | n2339 ;
  assign n12970 = n2131 | n10438 ;
  assign n12972 = n12971 ^ n12970 ^ 1'b0 ;
  assign n12973 = n8759 ^ n1550 ^ 1'b0 ;
  assign n12974 = n3807 & n12973 ;
  assign n12975 = n1300 & n12034 ;
  assign n12976 = ~n532 & n12975 ;
  assign n12977 = n10132 | n11265 ;
  assign n12978 = n2850 & ~n3931 ;
  assign n12979 = n627 & ~n3064 ;
  assign n12980 = n10878 | n12979 ;
  assign n12981 = n4856 & n5440 ;
  assign n12982 = n3602 | n8331 ;
  assign n12983 = ( n513 & n7673 ) | ( n513 & n12982 ) | ( n7673 & n12982 ) ;
  assign n12984 = n12983 ^ n4406 ^ 1'b0 ;
  assign n12985 = ~n6944 & n11707 ;
  assign n12986 = n7863 ^ n4889 ^ 1'b0 ;
  assign n12987 = n549 & n10657 ;
  assign n12988 = n5917 ^ n1388 ^ 1'b0 ;
  assign n12989 = ~n2303 & n12988 ;
  assign n12990 = n3542 ^ n497 ^ 1'b0 ;
  assign n12991 = n8167 | n12990 ;
  assign n12992 = n11513 ^ n1020 ^ 1'b0 ;
  assign n12993 = n4812 & ~n6320 ;
  assign n12994 = n729 & ~n9429 ;
  assign n12995 = n12993 & n12994 ;
  assign n12996 = n10107 & n12995 ;
  assign n12997 = n7416 ^ n3885 ^ 1'b0 ;
  assign n12998 = n12996 & ~n12997 ;
  assign n12999 = n382 & ~n649 ;
  assign n13000 = n6923 ^ n5270 ^ 1'b0 ;
  assign n13001 = n4640 ^ n3899 ^ 1'b0 ;
  assign n13002 = n872 | n6885 ;
  assign n13003 = n12057 | n13002 ;
  assign n13004 = n13001 & n13003 ;
  assign n13005 = ~n13001 & n13004 ;
  assign n13008 = n144 | n6060 ;
  assign n13006 = n673 | n2814 ;
  assign n13007 = n13006 ^ n722 ^ 1'b0 ;
  assign n13009 = n13008 ^ n13007 ^ 1'b0 ;
  assign n13010 = n4436 ^ n1029 ^ 1'b0 ;
  assign n13011 = ( ~n364 & n2162 ) | ( ~n364 & n3223 ) | ( n2162 & n3223 ) ;
  assign n13012 = n1815 & n5128 ;
  assign n13013 = n1710 & n13012 ;
  assign n13014 = n1768 & n3406 ;
  assign n13015 = ~n7803 & n13014 ;
  assign n13016 = n9055 & n13015 ;
  assign n13017 = n11117 ^ n1849 ^ 1'b0 ;
  assign n13018 = n1316 & ~n13017 ;
  assign n13019 = n6974 & n13018 ;
  assign n13020 = n149 | n7066 ;
  assign n13021 = n13020 ^ n1174 ^ 1'b0 ;
  assign n13022 = n4365 | n4990 ;
  assign n13023 = n5971 ^ n1344 ^ 1'b0 ;
  assign n13024 = n8291 ^ n800 ^ 1'b0 ;
  assign n13025 = ~n12976 & n13024 ;
  assign n13026 = n1602 ^ n495 ^ 1'b0 ;
  assign n13027 = n13026 ^ n5890 ^ 1'b0 ;
  assign n13028 = n1898 & ~n10154 ;
  assign n13029 = n8107 ^ n3193 ^ 1'b0 ;
  assign n13031 = n2083 & n8075 ;
  assign n13030 = n273 & ~n5161 ;
  assign n13032 = n13031 ^ n13030 ^ 1'b0 ;
  assign n13033 = n2967 & n5261 ;
  assign n13034 = n13033 ^ n6234 ^ 1'b0 ;
  assign n13035 = n13034 ^ n10098 ^ n850 ;
  assign n13036 = n7544 ^ n3929 ^ 1'b0 ;
  assign n13037 = n2933 & ~n13036 ;
  assign n13039 = n6253 ^ n461 ^ 1'b0 ;
  assign n13038 = n4037 & ~n11334 ;
  assign n13040 = n13039 ^ n13038 ^ 1'b0 ;
  assign n13041 = n1933 & n8764 ;
  assign n13042 = ~n7955 & n13041 ;
  assign n13043 = n10198 ^ n2214 ^ 1'b0 ;
  assign n13044 = n3788 & ~n6575 ;
  assign n13045 = n5458 & n13044 ;
  assign n13046 = ~n1370 & n13045 ;
  assign n13047 = n5041 & ~n13046 ;
  assign n13048 = n13047 ^ n4434 ^ 1'b0 ;
  assign n13049 = n4274 & n5348 ;
  assign n13050 = n2370 & ~n13049 ;
  assign n13051 = ~n9486 & n13050 ;
  assign n13052 = n1627 & ~n7707 ;
  assign n13053 = n3353 & ~n6769 ;
  assign n13054 = n13053 ^ n11570 ^ 1'b0 ;
  assign n13055 = n6349 ^ n1650 ^ 1'b0 ;
  assign n13056 = n8497 ^ n1060 ^ 1'b0 ;
  assign n13057 = n13055 & n13056 ;
  assign n13058 = n5659 & n13057 ;
  assign n13059 = n10464 | n13058 ;
  assign n13060 = n8611 & ~n13059 ;
  assign n13061 = n12114 ^ n5856 ^ 1'b0 ;
  assign n13062 = n2925 & ~n13061 ;
  assign n13063 = n13060 & n13062 ;
  assign n13064 = n13063 ^ n5529 ^ 1'b0 ;
  assign n13065 = n3469 & n9631 ;
  assign n13066 = ~n3803 & n13065 ;
  assign n13067 = n11105 ^ n3214 ^ 1'b0 ;
  assign n13068 = n3939 ^ n3753 ^ 1'b0 ;
  assign n13069 = n3643 ^ n1011 ^ 1'b0 ;
  assign n13070 = n13068 | n13069 ;
  assign n13071 = n13070 ^ n3025 ^ 1'b0 ;
  assign n13072 = n898 | n2446 ;
  assign n13073 = n9102 & n11197 ;
  assign n13074 = n814 & n2061 ;
  assign n13075 = ~n7067 & n13074 ;
  assign n13076 = n9793 & n13075 ;
  assign n13077 = n3604 | n5363 ;
  assign n13078 = n8399 & ~n13077 ;
  assign n13079 = n6660 & n13078 ;
  assign n13080 = n6995 ^ n520 ^ 1'b0 ;
  assign n13081 = n2519 | n4930 ;
  assign n13082 = n1078 & ~n13081 ;
  assign n13083 = n13082 ^ n3141 ^ n937 ;
  assign n13084 = n878 & ~n7922 ;
  assign n13085 = n13084 ^ n3074 ^ 1'b0 ;
  assign n13086 = ~n11409 & n13085 ;
  assign n13087 = ~n1375 & n2311 ;
  assign n13088 = n13087 ^ n11254 ^ 1'b0 ;
  assign n13089 = n13088 ^ n9705 ^ 1'b0 ;
  assign n13090 = n3803 ^ n128 ^ 1'b0 ;
  assign n13091 = n12989 & ~n13090 ;
  assign n13092 = n1443 ^ n1329 ^ 1'b0 ;
  assign n13093 = n13092 ^ n7008 ^ 1'b0 ;
  assign n13094 = ~n2987 & n7439 ;
  assign n13095 = n13094 ^ n2186 ^ 1'b0 ;
  assign n13096 = n3584 ^ n88 ^ 1'b0 ;
  assign n13097 = n12875 ^ n7272 ^ 1'b0 ;
  assign n13098 = ( n3516 & ~n4972 ) | ( n3516 & n9255 ) | ( ~n4972 & n9255 ) ;
  assign n13099 = n10819 & n13098 ;
  assign n13100 = n1133 & n13099 ;
  assign n13101 = n13097 & n13100 ;
  assign n13102 = n13101 ^ n6024 ^ 1'b0 ;
  assign n13103 = n13096 | n13102 ;
  assign n13104 = n13103 ^ n7771 ^ 1'b0 ;
  assign n13105 = n3748 ^ n3405 ^ 1'b0 ;
  assign n13106 = ~n3522 & n13105 ;
  assign n13107 = n5326 ^ n5286 ^ 1'b0 ;
  assign n13108 = n1537 & ~n13107 ;
  assign n13109 = ~n8130 & n13108 ;
  assign n13110 = n2254 | n5369 ;
  assign n13111 = n4016 & n9997 ;
  assign n13112 = n5415 ^ n14 ^ 1'b0 ;
  assign n13113 = ~n599 & n13112 ;
  assign n13114 = ~n2312 & n5971 ;
  assign n13115 = n9213 & ~n13114 ;
  assign n13116 = n4497 & n13115 ;
  assign n13117 = n12968 ^ n7508 ^ 1'b0 ;
  assign n13118 = n3717 | n13117 ;
  assign n13119 = n4899 | n5255 ;
  assign n13120 = n1357 & ~n13119 ;
  assign n13121 = n135 & ~n7669 ;
  assign n13122 = n6780 & ~n13121 ;
  assign n13123 = ~n9770 & n13122 ;
  assign n13124 = n13123 ^ n12242 ^ 1'b0 ;
  assign n13125 = n79 & ~n13124 ;
  assign n13126 = n1095 ^ n815 ^ 1'b0 ;
  assign n13127 = ~n510 & n3793 ;
  assign n13128 = ~n188 & n13127 ;
  assign n13129 = n7091 | n9691 ;
  assign n13130 = n13129 ^ n5436 ^ 1'b0 ;
  assign n13131 = n709 | n8079 ;
  assign n13132 = n8545 & n13131 ;
  assign n13133 = n1184 | n4835 ;
  assign n13134 = n13133 ^ n9058 ^ 1'b0 ;
  assign n13135 = n9100 ^ n300 ^ 1'b0 ;
  assign n13136 = n5677 | n13135 ;
  assign n13137 = n13136 ^ n3993 ^ 1'b0 ;
  assign n13138 = n13134 & ~n13137 ;
  assign n13139 = n13132 & n13138 ;
  assign n13140 = n3095 & ~n9019 ;
  assign n13141 = n36 & n749 ;
  assign n13142 = ~n749 & n13141 ;
  assign n13143 = n703 & ~n13142 ;
  assign n13144 = ~n703 & n13143 ;
  assign n13145 = n1398 | n13144 ;
  assign n13146 = n1398 & ~n13145 ;
  assign n13147 = n1687 & n13146 ;
  assign n13148 = ~n5415 & n13147 ;
  assign n13149 = n13148 ^ n4659 ^ 1'b0 ;
  assign n13150 = n3990 ^ n1543 ^ 1'b0 ;
  assign n13151 = n13150 ^ n325 ^ 1'b0 ;
  assign n13152 = n68 | n7182 ;
  assign n13153 = n8330 | n13152 ;
  assign n13154 = n3546 & n5970 ;
  assign n13155 = n1898 | n13154 ;
  assign n13156 = n13073 ^ n10942 ^ 1'b0 ;
  assign n13157 = n11935 ^ n10925 ^ 1'b0 ;
  assign n13158 = n736 & n13157 ;
  assign n13159 = n13158 ^ n2842 ^ 1'b0 ;
  assign n13160 = ~n11637 & n13159 ;
  assign n13161 = n9045 & n13160 ;
  assign n13162 = ~n13160 & n13161 ;
  assign n13163 = n8759 ^ n2101 ^ n178 ;
  assign n13164 = n13163 ^ n3037 ^ 1'b0 ;
  assign n13167 = ~n1207 & n3126 ;
  assign n13165 = n3941 ^ n1349 ^ 1'b0 ;
  assign n13166 = n4283 & ~n13165 ;
  assign n13168 = n13167 ^ n13166 ^ 1'b0 ;
  assign n13169 = n5863 ^ n1929 ^ n1330 ;
  assign n13170 = n13169 ^ n5963 ^ 1'b0 ;
  assign n13171 = n11332 & n11587 ;
  assign n13172 = n8299 | n10421 ;
  assign n13173 = ( n6434 & n7355 ) | ( n6434 & ~n13172 ) | ( n7355 & ~n13172 ) ;
  assign n13174 = n10664 ^ n1315 ^ 1'b0 ;
  assign n13175 = n4848 & n11064 ;
  assign n13176 = n13175 ^ n963 ^ 1'b0 ;
  assign n13177 = n236 | n13176 ;
  assign n13178 = n8053 | n10392 ;
  assign n13179 = n2529 | n13178 ;
  assign n13180 = n2150 | n5701 ;
  assign n13181 = n13180 ^ n4898 ^ 1'b0 ;
  assign n13182 = n941 | n7380 ;
  assign n13183 = n724 & ~n13182 ;
  assign n13184 = ~n2453 & n13183 ;
  assign n13185 = n1431 ^ n1227 ^ n1019 ;
  assign n13186 = ~n11417 & n13185 ;
  assign n13187 = n5421 & ~n5551 ;
  assign n13188 = n13186 & n13187 ;
  assign n13189 = n80 & ~n1476 ;
  assign n13190 = n8411 & n13189 ;
  assign n13191 = n13190 ^ n5447 ^ 1'b0 ;
  assign n13193 = ~n4336 & n8527 ;
  assign n13192 = n1399 & n12173 ;
  assign n13194 = n13193 ^ n13192 ^ 1'b0 ;
  assign n13195 = ( n2537 & n5217 ) | ( n2537 & ~n9542 ) | ( n5217 & ~n9542 ) ;
  assign n13196 = n5254 & n11430 ;
  assign n13198 = n37 | n3464 ;
  assign n13199 = n2096 & ~n13198 ;
  assign n13197 = n2547 & ~n4085 ;
  assign n13200 = n13199 ^ n13197 ^ 1'b0 ;
  assign n13201 = n9212 & n13200 ;
  assign n13202 = n581 & ~n1772 ;
  assign n13203 = n13202 ^ n5694 ^ 1'b0 ;
  assign n13204 = n4312 & ~n13203 ;
  assign n13205 = n5859 ^ n2963 ^ 1'b0 ;
  assign n13206 = n1225 | n13205 ;
  assign n13207 = ~n9627 & n13206 ;
  assign n13208 = n995 & n13207 ;
  assign n13209 = n7261 & ~n13208 ;
  assign n13210 = n80 | n3735 ;
  assign n13211 = n3735 & ~n13210 ;
  assign n13212 = n3690 | n13211 ;
  assign n13213 = n13211 & ~n13212 ;
  assign n13214 = n2311 | n13213 ;
  assign n13215 = n2311 & ~n13214 ;
  assign n13216 = n13215 ^ n11274 ^ 1'b0 ;
  assign n13217 = n5551 | n13216 ;
  assign n13218 = n865 & ~n8737 ;
  assign n13219 = ~n4556 & n13218 ;
  assign n13220 = n3988 ^ n2082 ^ 1'b0 ;
  assign n13221 = n5586 ^ n614 ^ 1'b0 ;
  assign n13222 = n13220 & ~n13221 ;
  assign n13223 = n11150 & n13222 ;
  assign n13226 = n50 & n310 ;
  assign n13227 = ~n310 & n13226 ;
  assign n13228 = n1467 & ~n13227 ;
  assign n13229 = n13227 & n13228 ;
  assign n13230 = n616 | n13229 ;
  assign n13231 = n616 & ~n13230 ;
  assign n13232 = n1852 & ~n2131 ;
  assign n13233 = n13231 & n13232 ;
  assign n13224 = ~n1323 & n1731 ;
  assign n13225 = n1323 & n13224 ;
  assign n13234 = n13233 ^ n13225 ^ 1'b0 ;
  assign n13235 = n6950 & ~n7299 ;
  assign n13236 = n1627 & n4899 ;
  assign n13237 = n13236 ^ n3479 ^ 1'b0 ;
  assign n13238 = n13237 ^ n5002 ^ 1'b0 ;
  assign n13239 = n13235 | n13238 ;
  assign n13240 = n13235 & ~n13239 ;
  assign n13241 = n13234 & n13240 ;
  assign n13242 = n2395 & n4336 ;
  assign n13243 = n13242 ^ n4440 ^ 1'b0 ;
  assign n13244 = n5178 & n13243 ;
  assign n13245 = n3264 & n13244 ;
  assign n13246 = n556 | n13245 ;
  assign n13247 = n168 & ~n5885 ;
  assign n13248 = n13247 ^ n3080 ^ 1'b0 ;
  assign n13249 = ~n5554 & n13248 ;
  assign n13250 = n13246 & n13249 ;
  assign n13251 = n6095 ^ n4299 ^ 1'b0 ;
  assign n13252 = n11840 | n13251 ;
  assign n13253 = ~n10241 & n13252 ;
  assign n13254 = n3193 ^ n434 ^ 1'b0 ;
  assign n13255 = n161 & ~n13254 ;
  assign n13256 = n8234 & ~n13255 ;
  assign n13257 = n13256 ^ n3171 ^ 1'b0 ;
  assign n13258 = n1885 | n13257 ;
  assign n13259 = n675 & ~n13258 ;
  assign n13260 = ~n2163 & n13259 ;
  assign n13261 = n5953 & ~n13260 ;
  assign n13262 = n2733 & ~n6388 ;
  assign n13263 = n13262 ^ n4269 ^ 1'b0 ;
  assign n13264 = n11694 ^ n9153 ^ 1'b0 ;
  assign n13265 = n10736 & n13264 ;
  assign n13266 = ~n662 & n6541 ;
  assign n13267 = n8199 & n9086 ;
  assign n13268 = n13267 ^ n4434 ^ 1'b0 ;
  assign n13269 = n5316 & n7056 ;
  assign n13270 = ~n3939 & n13269 ;
  assign n13271 = n3484 ^ n3407 ^ 1'b0 ;
  assign n13272 = ~n7476 & n13271 ;
  assign n13273 = n13272 ^ n12259 ^ 1'b0 ;
  assign n13274 = n5603 & ~n13273 ;
  assign n13275 = n754 & n13274 ;
  assign n13278 = n6300 ^ n5179 ^ 1'b0 ;
  assign n13276 = ~n1505 & n5096 ;
  assign n13277 = n13276 ^ n3009 ^ 1'b0 ;
  assign n13279 = n13278 ^ n13277 ^ 1'b0 ;
  assign n13280 = ~n5856 & n6945 ;
  assign n13281 = n13280 ^ n4689 ^ 1'b0 ;
  assign n13282 = n279 & n13281 ;
  assign n13283 = ~n9026 & n11744 ;
  assign n13284 = n2654 & n6434 ;
  assign n13285 = n3693 & ~n13284 ;
  assign n13287 = n2014 | n2455 ;
  assign n13288 = n1359 | n13287 ;
  assign n13289 = n1887 & ~n13288 ;
  assign n13286 = n2828 ^ n2759 ^ 1'b0 ;
  assign n13290 = n13289 ^ n13286 ^ 1'b0 ;
  assign n13291 = n2200 & n13290 ;
  assign n13292 = n7395 ^ n1582 ^ 1'b0 ;
  assign n13293 = n578 ^ n532 ^ 1'b0 ;
  assign n13294 = n5180 ^ n3567 ^ 1'b0 ;
  assign n13295 = n13293 & n13294 ;
  assign n13296 = n1178 | n8900 ;
  assign n13297 = n13296 ^ n8982 ^ 1'b0 ;
  assign n13298 = n13297 ^ n7408 ^ 1'b0 ;
  assign n13299 = n2076 | n5528 ;
  assign n13300 = ~n4216 & n6300 ;
  assign n13301 = n13300 ^ n4899 ^ 1'b0 ;
  assign n13302 = ~n190 & n1547 ;
  assign n13303 = ~n940 & n13302 ;
  assign n13304 = n1087 & ~n13303 ;
  assign n13305 = n2549 & n7399 ;
  assign n13306 = n13305 ^ n8946 ^ 1'b0 ;
  assign n13307 = ~n567 & n5915 ;
  assign n13308 = n13307 ^ n6916 ^ 1'b0 ;
  assign n13309 = n385 | n13308 ;
  assign n13310 = n6880 & n13309 ;
  assign n13311 = n6773 & n9000 ;
  assign n13312 = n2560 & n13311 ;
  assign n13319 = n4169 & ~n7647 ;
  assign n13320 = ~n4169 & n13319 ;
  assign n13313 = ~n324 & n552 ;
  assign n13314 = ~n552 & n13313 ;
  assign n13315 = ~n481 & n13314 ;
  assign n13316 = ~n3940 & n13315 ;
  assign n13317 = n13316 ^ n68 ^ 1'b0 ;
  assign n13318 = ~n9099 & n13317 ;
  assign n13321 = n13320 ^ n13318 ^ 1'b0 ;
  assign n13322 = n13321 ^ n82 ^ 1'b0 ;
  assign n13323 = x2 | n4125 ;
  assign n13324 = n13323 ^ n4737 ^ 1'b0 ;
  assign n13325 = n406 & ~n1739 ;
  assign n13326 = n13325 ^ n5328 ^ 1'b0 ;
  assign n13327 = n7767 & n13326 ;
  assign n13328 = n13324 & n13327 ;
  assign n13329 = n2582 & n13328 ;
  assign n13330 = n6128 & n7376 ;
  assign n13331 = ~n13329 & n13330 ;
  assign n13332 = n13331 ^ n7040 ^ 1'b0 ;
  assign n13333 = ~n280 & n1920 ;
  assign n13334 = n13333 ^ n2604 ^ 1'b0 ;
  assign n13335 = n9221 ^ n1716 ^ 1'b0 ;
  assign n13336 = n2222 | n13335 ;
  assign n13337 = n3440 & ~n6060 ;
  assign n13338 = ~n754 & n3583 ;
  assign n13339 = n6534 & n13338 ;
  assign n13340 = ~n10760 & n13339 ;
  assign n13341 = n27 | n5566 ;
  assign n13342 = n1001 | n12213 ;
  assign n13343 = n13342 ^ n114 ^ 1'b0 ;
  assign n13344 = n13343 ^ n519 ^ 1'b0 ;
  assign n13345 = n432 | n8814 ;
  assign n13346 = n13345 ^ n1566 ^ 1'b0 ;
  assign n13347 = n79 | n4543 ;
  assign n13348 = n7244 | n13347 ;
  assign n13349 = n7827 ^ n6039 ^ 1'b0 ;
  assign n13350 = n3584 & n13349 ;
  assign n13351 = n13350 ^ n3068 ^ 1'b0 ;
  assign n13352 = n7408 | n13351 ;
  assign n13353 = n2623 & n6194 ;
  assign n13354 = n13353 ^ n958 ^ 1'b0 ;
  assign n13355 = n4523 & ~n5571 ;
  assign n13356 = ~n9091 & n13355 ;
  assign n13357 = n6631 & ~n8792 ;
  assign n13358 = n1458 & ~n13357 ;
  assign n13359 = n10668 ^ n68 ^ 1'b0 ;
  assign n13360 = ~n908 & n5428 ;
  assign n13361 = n13360 ^ n3483 ^ 1'b0 ;
  assign n13362 = n6247 & ~n13361 ;
  assign n13363 = n12062 ^ n3173 ^ 1'b0 ;
  assign n13364 = n310 | n5228 ;
  assign n13365 = n491 & n3741 ;
  assign n13366 = ~n13364 & n13365 ;
  assign n13367 = ~n1229 & n5551 ;
  assign n13368 = n12180 ^ n3001 ^ 1'b0 ;
  assign n13369 = n2092 & n13368 ;
  assign n13370 = n3820 & n9149 ;
  assign n13371 = n13370 ^ n7862 ^ 1'b0 ;
  assign n13372 = n9810 ^ n3806 ^ 1'b0 ;
  assign n13373 = n10303 ^ n9666 ^ 1'b0 ;
  assign n13374 = n8972 & ~n13373 ;
  assign n13375 = n13374 ^ n9164 ^ 1'b0 ;
  assign n13376 = n203 & ~n1644 ;
  assign n13377 = n13376 ^ n12984 ^ 1'b0 ;
  assign n13378 = ( ~n540 & n4653 ) | ( ~n540 & n8130 ) | ( n4653 & n8130 ) ;
  assign n13379 = n13364 ^ n2166 ^ 1'b0 ;
  assign n13380 = n327 ^ n252 ^ 1'b0 ;
  assign n13381 = ~n5568 & n6953 ;
  assign n13382 = n13381 ^ n6981 ^ n1499 ;
  assign n13383 = n9428 ^ n2222 ^ 1'b0 ;
  assign n13384 = n3093 & n13383 ;
  assign n13385 = ~n11311 & n13384 ;
  assign n13386 = n7277 & n13385 ;
  assign n13387 = n3211 | n10656 ;
  assign n13388 = n2849 & ~n11301 ;
  assign n13389 = ~n6089 & n6822 ;
  assign n13390 = n616 | n5004 ;
  assign n13391 = n4485 ^ n2100 ^ 1'b0 ;
  assign n13392 = n2076 ^ n1668 ^ 1'b0 ;
  assign n13393 = n1642 & ~n13392 ;
  assign n13394 = n13393 ^ n9194 ^ 1'b0 ;
  assign n13395 = n13391 & n13394 ;
  assign n13396 = n2984 ^ n1212 ^ n410 ;
  assign n13397 = n13396 ^ n323 ^ 1'b0 ;
  assign n13398 = n6037 ^ n3183 ^ 1'b0 ;
  assign n13399 = ~n55 & n5562 ;
  assign n13400 = ~n5562 & n13399 ;
  assign n13401 = ~n9578 & n10805 ;
  assign n13402 = n9578 & n13401 ;
  assign n13403 = n13400 | n13402 ;
  assign n13404 = n13400 & ~n13403 ;
  assign n13407 = n12046 ^ n3998 ^ 1'b0 ;
  assign n13405 = ( n2376 & n2714 ) | ( n2376 & n7155 ) | ( n2714 & n7155 ) ;
  assign n13406 = ~n7106 & n13405 ;
  assign n13408 = n13407 ^ n13406 ^ 1'b0 ;
  assign n13409 = n9794 ^ n246 ^ 1'b0 ;
  assign n13410 = n13409 ^ n7849 ^ 1'b0 ;
  assign n13411 = n13408 & ~n13410 ;
  assign n13412 = n2501 ^ n2385 ^ 1'b0 ;
  assign n13413 = n3866 & ~n9791 ;
  assign n13414 = n13412 & n13413 ;
  assign n13421 = n6262 & ~n7087 ;
  assign n13422 = n13421 ^ n6700 ^ 1'b0 ;
  assign n13415 = n807 | n2469 ;
  assign n13416 = n1965 & ~n13415 ;
  assign n13417 = n228 & n3144 ;
  assign n13418 = n34 | n13417 ;
  assign n13419 = n741 & ~n13418 ;
  assign n13420 = n13416 & ~n13419 ;
  assign n13423 = n13422 ^ n13420 ^ 1'b0 ;
  assign n13424 = n628 & n13423 ;
  assign n13425 = n12310 ^ n6090 ^ 1'b0 ;
  assign n13426 = n8868 & ~n13425 ;
  assign n13427 = ~n8923 & n13426 ;
  assign n13428 = n5127 & ~n5170 ;
  assign n13429 = n13428 ^ n9691 ^ 1'b0 ;
  assign n13430 = n9900 & ~n13429 ;
  assign n13431 = n4241 ^ n1184 ^ 1'b0 ;
  assign n13432 = n2236 | n13431 ;
  assign n13433 = n13432 ^ n3007 ^ 1'b0 ;
  assign n13434 = ~n5207 & n13433 ;
  assign n13437 = n1438 & ~n2494 ;
  assign n13435 = n1285 | n7043 ;
  assign n13436 = n4203 & ~n13435 ;
  assign n13438 = n13437 ^ n13436 ^ 1'b0 ;
  assign n13439 = n308 & ~n364 ;
  assign n13440 = n9061 ^ n5979 ^ 1'b0 ;
  assign n13441 = n2608 ^ n382 ^ 1'b0 ;
  assign n13442 = ~n3583 & n13441 ;
  assign n13443 = ~n3431 & n13442 ;
  assign n13444 = n3185 & n10255 ;
  assign n13445 = ~n847 & n3360 ;
  assign n13446 = n13445 ^ n2919 ^ 1'b0 ;
  assign n13447 = n6857 & ~n13446 ;
  assign n13448 = ~n3326 & n13274 ;
  assign n13449 = n4660 & n13448 ;
  assign n13450 = n4708 ^ n2260 ^ 1'b0 ;
  assign n13451 = n3459 & n5094 ;
  assign n13452 = ~n689 & n5846 ;
  assign n13453 = n13452 ^ n573 ^ 1'b0 ;
  assign n13454 = n9020 & ~n13453 ;
  assign n13455 = n13451 & n13454 ;
  assign n13458 = n9227 ^ n4189 ^ 1'b0 ;
  assign n13459 = n4757 & n13458 ;
  assign n13460 = ~n4294 & n13459 ;
  assign n13461 = n13460 ^ n233 ^ 1'b0 ;
  assign n13456 = n1927 & ~n6192 ;
  assign n13457 = n10475 & n13456 ;
  assign n13462 = n13461 ^ n13457 ^ 1'b0 ;
  assign n13463 = n5849 ^ n28 ^ 1'b0 ;
  assign n13464 = n1255 & n4720 ;
  assign n13465 = ~n1255 & n13464 ;
  assign n13466 = n13463 | n13465 ;
  assign n13467 = n3426 | n13466 ;
  assign n13470 = ~n3780 & n4434 ;
  assign n13471 = n13470 ^ n6094 ^ 1'b0 ;
  assign n13468 = ~n158 & n3096 ;
  assign n13469 = n4241 & n13468 ;
  assign n13472 = n13471 ^ n13469 ^ 1'b0 ;
  assign n13473 = ~n4846 & n13472 ;
  assign n13474 = n5551 & ~n7981 ;
  assign n13475 = ~n4121 & n4155 ;
  assign n13476 = n13475 ^ n11588 ^ 1'b0 ;
  assign n13477 = n4044 | n8950 ;
  assign n13478 = n13477 ^ n12046 ^ 1'b0 ;
  assign n13479 = n19 & ~n10966 ;
  assign n13480 = ~n7476 & n13479 ;
  assign n13481 = ~n3637 & n6753 ;
  assign n13482 = n274 | n11046 ;
  assign n13483 = n11895 ^ n501 ^ 1'b0 ;
  assign n13484 = n5503 | n8221 ;
  assign n13485 = n13483 | n13484 ;
  assign n13486 = n6219 ^ n3036 ^ 1'b0 ;
  assign n13487 = n3603 & n13486 ;
  assign n13488 = n13487 ^ n10481 ^ 1'b0 ;
  assign n13489 = n1915 ^ n452 ^ 1'b0 ;
  assign n13490 = n5452 & n13489 ;
  assign n13491 = n2346 & n13490 ;
  assign n13492 = n7737 & n13491 ;
  assign n13493 = n1519 & n3263 ;
  assign n13494 = n13493 ^ n4700 ^ 1'b0 ;
  assign n13495 = n148 | n592 ;
  assign n13496 = n592 & ~n13495 ;
  assign n13497 = n3890 & ~n13496 ;
  assign n13498 = ~n3890 & n13497 ;
  assign n13499 = n2586 & ~n2941 ;
  assign n13500 = ~n2586 & n13499 ;
  assign n13501 = n2732 & ~n2861 ;
  assign n13502 = ~n484 & n13501 ;
  assign n13503 = ~n1323 & n13502 ;
  assign n13504 = n13500 & n13503 ;
  assign n13505 = n766 & n13504 ;
  assign n13506 = n557 & n7830 ;
  assign n13507 = n294 | n1573 ;
  assign n13508 = n1573 & ~n13507 ;
  assign n13509 = ~n35 & n46 ;
  assign n13510 = n35 & n13509 ;
  assign n13511 = n50 & n13510 ;
  assign n13512 = n291 & n13511 ;
  assign n13513 = ~n291 & n13512 ;
  assign n13514 = n830 & n13513 ;
  assign n13515 = n13514 ^ n158 ^ 1'b0 ;
  assign n13516 = ( ~n13506 & n13508 ) | ( ~n13506 & n13515 ) | ( n13508 & n13515 ) ;
  assign n13517 = n13505 & ~n13516 ;
  assign n13518 = n13498 & n13517 ;
  assign n13519 = ~n3017 & n3931 ;
  assign n13520 = n6763 & n10942 ;
  assign n13521 = n13519 & n13520 ;
  assign n13522 = n5261 | n10025 ;
  assign n13523 = n13522 ^ n6992 ^ 1'b0 ;
  assign n13524 = n4183 & ~n13523 ;
  assign n13525 = ~n10012 & n13524 ;
  assign n13526 = n7707 & ~n13525 ;
  assign n13527 = ~n542 & n2244 ;
  assign n13528 = n5393 ^ n4575 ^ 1'b0 ;
  assign n13529 = n5612 | n6133 ;
  assign n13530 = n13529 ^ n763 ^ 1'b0 ;
  assign n13531 = n653 & ~n12354 ;
  assign n13532 = n1026 & ~n4267 ;
  assign n13533 = n5359 & n6343 ;
  assign n13534 = n13533 ^ n3402 ^ 1'b0 ;
  assign n13535 = n6260 | n13534 ;
  assign n13536 = n13309 & ~n13535 ;
  assign n13537 = n8309 ^ n2124 ^ 1'b0 ;
  assign n13538 = n5758 & ~n7289 ;
  assign n13539 = n13537 & ~n13538 ;
  assign n13540 = n12908 & n13539 ;
  assign n13543 = n9131 ^ n1802 ^ 1'b0 ;
  assign n13541 = n1546 & ~n10389 ;
  assign n13542 = ~n4941 & n13541 ;
  assign n13544 = n13543 ^ n13542 ^ 1'b0 ;
  assign n13546 = n4249 ^ n3467 ^ 1'b0 ;
  assign n13545 = n141 | n8272 ;
  assign n13547 = n13546 ^ n13545 ^ 1'b0 ;
  assign n13548 = x0 & n3013 ;
  assign n13549 = n13548 ^ n2236 ^ 1'b0 ;
  assign n13550 = ~n2754 & n13549 ;
  assign n13551 = n12301 & n13550 ;
  assign n13552 = n356 & n6464 ;
  assign n13553 = n13552 ^ n4081 ^ 1'b0 ;
  assign n13554 = n13553 ^ n6995 ^ x0 ;
  assign n13555 = n3229 & ~n3622 ;
  assign n13556 = n6474 | n6878 ;
  assign n13557 = n13556 ^ n6923 ^ 1'b0 ;
  assign n13558 = n2469 | n13557 ;
  assign n13559 = n2576 & ~n13558 ;
  assign n13560 = n3886 & ~n9121 ;
  assign n13561 = n13559 & n13560 ;
  assign n13562 = n2085 & ~n7597 ;
  assign n13563 = n2222 | n9437 ;
  assign n13564 = n13563 ^ n12290 ^ n7784 ;
  assign n13565 = n1015 | n13564 ;
  assign n13566 = n13562 | n13565 ;
  assign n13567 = n3292 ^ n3116 ^ 1'b0 ;
  assign n13568 = n7391 & ~n13567 ;
  assign n13569 = n13568 ^ n2721 ^ 1'b0 ;
  assign n13570 = ~n5364 & n13286 ;
  assign n13571 = n3775 & n13570 ;
  assign n13572 = n11040 | n12541 ;
  assign n13573 = n1961 & ~n4533 ;
  assign n13574 = n1937 ^ n683 ^ 1'b0 ;
  assign n13575 = n7926 | n13574 ;
  assign n13576 = n13573 | n13575 ;
  assign n13577 = n8747 ^ n1010 ^ 1'b0 ;
  assign n13578 = n1591 & n4104 ;
  assign n13579 = ~n17 & n6865 ;
  assign n13580 = n1276 & n13579 ;
  assign n13581 = n13580 ^ n6377 ^ 1'b0 ;
  assign n13583 = n734 & ~n1946 ;
  assign n13582 = ~n4407 & n4972 ;
  assign n13584 = n13583 ^ n13582 ^ 1'b0 ;
  assign n13585 = n1455 ^ n469 ^ 1'b0 ;
  assign n13586 = n9405 ^ n3882 ^ 1'b0 ;
  assign n13587 = n9272 ^ n1810 ^ 1'b0 ;
  assign n13588 = n1166 & n13587 ;
  assign n13589 = ~n11758 & n13588 ;
  assign n13590 = n1766 & n13589 ;
  assign n13591 = n10309 ^ n2992 ^ 1'b0 ;
  assign n13592 = n378 | n13591 ;
  assign n13593 = n364 | n5659 ;
  assign n13594 = n13592 & ~n13593 ;
  assign n13595 = n737 | n11638 ;
  assign n13596 = n6653 ^ n3118 ^ 1'b0 ;
  assign n13597 = n1879 & n4419 ;
  assign n13598 = n1860 | n12407 ;
  assign n13599 = n13598 ^ n1956 ^ 1'b0 ;
  assign n13600 = n3166 & n9136 ;
  assign n13601 = n532 | n2187 ;
  assign n13605 = n7330 ^ n4878 ^ 1'b0 ;
  assign n13606 = n8349 | n13605 ;
  assign n13602 = n9187 ^ n34 ^ 1'b0 ;
  assign n13603 = n2129 & n13602 ;
  assign n13604 = n2537 & n13603 ;
  assign n13607 = n13606 ^ n13604 ^ 1'b0 ;
  assign n13608 = n892 | n7669 ;
  assign n13609 = ~n1829 & n1929 ;
  assign n13610 = n13608 & n13609 ;
  assign n13611 = n13610 ^ n3369 ^ 1'b0 ;
  assign n13612 = n636 ^ n17 ^ 1'b0 ;
  assign n13613 = n13612 ^ n8183 ^ 1'b0 ;
  assign n13614 = ( n4815 & n5760 ) | ( n4815 & ~n12263 ) | ( n5760 & ~n12263 ) ;
  assign n13615 = n10265 ^ n5714 ^ 1'b0 ;
  assign n13616 = n12706 ^ n6700 ^ 1'b0 ;
  assign n13617 = ~n7310 & n13616 ;
  assign n13618 = ~n1129 & n5749 ;
  assign n13619 = n4355 & ~n7054 ;
  assign n13620 = ~n9538 & n12761 ;
  assign n13621 = n7294 ^ n3853 ^ n2547 ;
  assign n13622 = n4407 | n5043 ;
  assign n13623 = n1080 | n7103 ;
  assign n13624 = n9292 | n13623 ;
  assign n13625 = n7777 & ~n7936 ;
  assign n13626 = n5545 & n13625 ;
  assign n13627 = n4037 & n9939 ;
  assign n13628 = n5196 ^ n4606 ^ 1'b0 ;
  assign n13629 = n8514 ^ n3269 ^ 1'b0 ;
  assign n13630 = n13629 ^ n12721 ^ 1'b0 ;
  assign n13631 = n13628 | n13630 ;
  assign n13632 = n13631 ^ n9520 ^ 1'b0 ;
  assign n13633 = ~n7258 & n13632 ;
  assign n13634 = n1645 & n8574 ;
  assign n13635 = ~n690 & n4668 ;
  assign n13636 = n415 & n958 ;
  assign n13637 = n13636 ^ n6540 ^ 1'b0 ;
  assign n13638 = n1645 & n4448 ;
  assign n13639 = n13638 ^ n9986 ^ 1'b0 ;
  assign n13640 = n3297 & n12169 ;
  assign n13641 = n109 & n13640 ;
  assign n13642 = n2266 & ~n9792 ;
  assign n13643 = n2661 & n13642 ;
  assign n13644 = n13643 ^ n86 ^ 1'b0 ;
  assign n13645 = n187 & ~n8876 ;
  assign n13646 = ~n6498 & n13645 ;
  assign n13647 = n561 & ~n5821 ;
  assign n13648 = n13356 & n13647 ;
  assign n13649 = n1155 & n1872 ;
  assign n13650 = n13649 ^ n12765 ^ 1'b0 ;
  assign n13652 = n3570 ^ n2483 ^ 1'b0 ;
  assign n13651 = n8106 | n9074 ;
  assign n13653 = n13652 ^ n13651 ^ 1'b0 ;
  assign n13654 = n11486 & ~n13653 ;
  assign n13655 = n1575 | n2233 ;
  assign n13656 = n86 & ~n13655 ;
  assign n13657 = n6102 & n8024 ;
  assign n13658 = n489 & n596 ;
  assign n13659 = n1010 & n7523 ;
  assign n13660 = n13659 ^ n7735 ^ 1'b0 ;
  assign n13661 = ~n7803 & n13660 ;
  assign n13662 = n8783 ^ n4939 ^ 1'b0 ;
  assign n13663 = ~n13661 & n13662 ;
  assign n13664 = ~n142 & n2910 ;
  assign n13665 = n8575 & n13664 ;
  assign n13666 = ~n3509 & n9789 ;
  assign n13667 = n13666 ^ n6046 ^ 1'b0 ;
  assign n13668 = n2617 | n8994 ;
  assign n13669 = n13668 ^ n4121 ^ 1'b0 ;
  assign n13670 = n13669 ^ n6620 ^ 1'b0 ;
  assign n13671 = n4300 | n8022 ;
  assign n13672 = ~n11266 & n13671 ;
  assign n13673 = n13672 ^ n5575 ^ 1'b0 ;
  assign n13674 = n190 | n4131 ;
  assign n13675 = n12350 & ~n13674 ;
  assign n13676 = n13675 ^ n3676 ^ 1'b0 ;
  assign n13677 = n507 & n3589 ;
  assign n13678 = n9102 & n13677 ;
  assign n13679 = n4872 ^ n2604 ^ 1'b0 ;
  assign n13680 = ~n6972 & n13679 ;
  assign n13681 = ~n13678 & n13680 ;
  assign n13682 = n483 | n1671 ;
  assign n13683 = n13682 ^ n1227 ^ 1'b0 ;
  assign n13684 = n5056 ^ n4698 ^ 1'b0 ;
  assign n13685 = n10384 & ~n13684 ;
  assign n13686 = n6418 & n9019 ;
  assign n13687 = ~n1530 & n4487 ;
  assign n13688 = n4207 & ~n4733 ;
  assign n13689 = n8488 ^ n3719 ^ 1'b0 ;
  assign n13690 = n12742 ^ n2799 ^ 1'b0 ;
  assign n13691 = n963 ^ n915 ^ 1'b0 ;
  assign n13692 = n8602 & n13691 ;
  assign n13693 = n13692 ^ n5089 ^ 1'b0 ;
  assign n13694 = n1820 & n13693 ;
  assign n13695 = n4315 & n9996 ;
  assign n13696 = n13695 ^ n7619 ^ 1'b0 ;
  assign n13697 = n5805 | n11136 ;
  assign n13698 = n10664 & ~n13697 ;
  assign n13699 = ~n3887 & n4480 ;
  assign n13700 = x11 & ~n745 ;
  assign n13701 = n3049 ^ n364 ^ 1'b0 ;
  assign n13702 = n13700 & n13701 ;
  assign n13704 = n4540 ^ n1052 ^ 1'b0 ;
  assign n13705 = n328 | n13704 ;
  assign n13703 = n1929 | n7336 ;
  assign n13706 = n13705 ^ n13703 ^ 1'b0 ;
  assign n13707 = n13706 ^ n5716 ^ 1'b0 ;
  assign n13708 = n7189 ^ n5725 ^ 1'b0 ;
  assign n13709 = n9692 ^ n2542 ^ 1'b0 ;
  assign n13710 = n13709 ^ n6190 ^ 1'b0 ;
  assign n13711 = n2238 ^ n1307 ^ 1'b0 ;
  assign n13713 = n6349 ^ n986 ^ 1'b0 ;
  assign n13712 = n724 & n1519 ;
  assign n13714 = n13713 ^ n13712 ^ 1'b0 ;
  assign n13715 = n1205 | n2252 ;
  assign n13716 = n10606 & ~n13715 ;
  assign n13717 = n252 | n13716 ;
  assign n13718 = n6607 ^ n2221 ^ 1'b0 ;
  assign n13719 = n13717 & n13718 ;
  assign n13720 = n11553 ^ n8134 ^ 1'b0 ;
  assign n13721 = n4051 & ~n12200 ;
  assign n13722 = n4137 ^ n159 ^ 1'b0 ;
  assign n13723 = n3037 | n13722 ;
  assign n13724 = n5714 & ~n8130 ;
  assign n13725 = n13724 ^ n1281 ^ 1'b0 ;
  assign n13726 = n13723 | n13725 ;
  assign n13727 = n3312 | n7597 ;
  assign n13728 = n13727 ^ n280 ^ 1'b0 ;
  assign n13729 = n13728 ^ n7214 ^ n618 ;
  assign n13730 = n1373 ^ n1246 ^ 1'b0 ;
  assign n13731 = n198 | n6156 ;
  assign n13732 = n2915 | n13731 ;
  assign n13733 = n13730 & n13732 ;
  assign n13734 = n13733 ^ n982 ^ 1'b0 ;
  assign n13735 = n10922 | n13734 ;
  assign n13736 = n3779 ^ n2790 ^ 1'b0 ;
  assign n13737 = n13736 ^ n3843 ^ 1'b0 ;
  assign n13738 = n9718 ^ x10 ^ 1'b0 ;
  assign n13739 = n7045 & ~n9753 ;
  assign n13740 = n13739 ^ n257 ^ 1'b0 ;
  assign n13741 = n12496 & n13740 ;
  assign n13742 = n7597 | n12991 ;
  assign n13743 = n7088 ^ n111 ^ 1'b0 ;
  assign n13744 = n13743 ^ n2303 ^ 1'b0 ;
  assign n13745 = n4227 & n13744 ;
  assign n13746 = n5557 & ~n5568 ;
  assign n13747 = ~n2157 & n13746 ;
  assign n13748 = ~n2577 & n3737 ;
  assign n13749 = n5208 & ~n13748 ;
  assign n13750 = n366 & ~n985 ;
  assign n13751 = n7994 & ~n13750 ;
  assign n13752 = n89 & ~n204 ;
  assign n13753 = n5090 & ~n13752 ;
  assign n13754 = n116 | n12110 ;
  assign n13755 = n3988 | n13754 ;
  assign n13756 = n3186 & n8637 ;
  assign n13757 = n2064 | n13756 ;
  assign n13758 = ~n2440 & n13757 ;
  assign n13759 = n5083 | n6028 ;
  assign n13760 = n4096 | n9619 ;
  assign n13761 = n5241 & ~n9014 ;
  assign n13762 = ~n1974 & n5144 ;
  assign n13763 = n1810 ^ x11 ^ 1'b0 ;
  assign n13764 = n4513 | n13763 ;
  assign n13765 = n60 | n10172 ;
  assign n13766 = n4460 & ~n13765 ;
  assign n13767 = n210 | n13766 ;
  assign n13768 = n13764 & ~n13767 ;
  assign n13769 = n581 & n4186 ;
  assign n13770 = n1693 | n13769 ;
  assign n13771 = n13768 & ~n13770 ;
  assign n13772 = n1655 ^ n456 ^ 1'b0 ;
  assign n13773 = n5708 | n8056 ;
  assign n13774 = n3133 ^ n787 ^ 1'b0 ;
  assign n13775 = n284 & ~n13774 ;
  assign n13776 = n13775 ^ n2430 ^ 1'b0 ;
  assign n13777 = n10922 ^ n5610 ^ n1860 ;
  assign n13782 = n170 ^ n102 ^ 1'b0 ;
  assign n13778 = ~n7539 & n12025 ;
  assign n13779 = n984 & n1469 ;
  assign n13780 = n13779 ^ n10001 ^ 1'b0 ;
  assign n13781 = n13778 & n13780 ;
  assign n13783 = n13782 ^ n13781 ^ 1'b0 ;
  assign n13784 = ~n2717 & n13783 ;
  assign n13785 = n2676 | n10386 ;
  assign n13786 = n2176 & ~n13785 ;
  assign n13787 = n605 | n13786 ;
  assign n13788 = n13787 ^ n585 ^ 1'b0 ;
  assign n13789 = n13788 ^ n6250 ^ 1'b0 ;
  assign n13790 = ~n2090 & n13789 ;
  assign n13791 = n3888 & n13790 ;
  assign n13792 = n274 & ~n4927 ;
  assign n13793 = ~n6595 & n8925 ;
  assign n13794 = n6780 & ~n9898 ;
  assign n13795 = n1518 & n1920 ;
  assign n13796 = ~n6072 & n13795 ;
  assign n13797 = n13794 & n13796 ;
  assign n13798 = n4355 & ~n6887 ;
  assign n13799 = n13797 | n13798 ;
  assign n13800 = n2843 ^ n2460 ^ 1'b0 ;
  assign n13801 = n4249 & ~n13800 ;
  assign n13802 = n9384 ^ n19 ^ 1'b0 ;
  assign n13803 = n12097 & ~n13802 ;
  assign n13804 = n7726 ^ n3927 ^ 1'b0 ;
  assign n13805 = n6194 & ~n13804 ;
  assign n13806 = n6320 ^ n273 ^ 1'b0 ;
  assign n13807 = n13806 ^ n10651 ^ 1'b0 ;
  assign n13808 = n10718 & n13807 ;
  assign n13809 = ~n1759 & n11476 ;
  assign n13810 = n13809 ^ n891 ^ 1'b0 ;
  assign n13811 = n2774 | n3514 ;
  assign n13812 = n5613 & n8126 ;
  assign n13813 = ~n296 & n13812 ;
  assign n13814 = n1900 & ~n13813 ;
  assign n13815 = n13814 ^ n6166 ^ 1'b0 ;
  assign n13816 = ~n58 & n220 ;
  assign n13817 = n2065 | n13816 ;
  assign n13818 = ~n5067 & n7289 ;
  assign n13819 = n13818 ^ n6289 ^ 1'b0 ;
  assign n13820 = n294 ^ n30 ^ 1'b0 ;
  assign n13821 = n3707 & ~n7639 ;
  assign n13822 = n1959 | n11098 ;
  assign n13823 = n13822 ^ n713 ^ 1'b0 ;
  assign n13824 = ~n4533 & n13823 ;
  assign n13825 = n2633 ^ n1058 ^ 1'b0 ;
  assign n13826 = ~n4023 & n13825 ;
  assign n13827 = n13826 ^ n4915 ^ 1'b0 ;
  assign n13828 = n1740 & ~n9925 ;
  assign n13829 = n3868 ^ n1079 ^ 1'b0 ;
  assign n13830 = n6323 | n12125 ;
  assign n13831 = n13830 ^ n98 ^ 1'b0 ;
  assign n13832 = n9104 ^ n3791 ^ 1'b0 ;
  assign n13833 = n3389 & n4869 ;
  assign n13834 = n13833 ^ n2305 ^ 1'b0 ;
  assign n13835 = ~n13563 & n13834 ;
  assign n13836 = ~n11003 & n13835 ;
  assign n13837 = n6933 ^ n308 ^ 1'b0 ;
  assign n13838 = ~n12913 & n13837 ;
  assign n13839 = n2573 ^ n236 ^ 1'b0 ;
  assign n13840 = n1660 ^ n1529 ^ 1'b0 ;
  assign n13841 = n13839 & ~n13840 ;
  assign n13842 = n551 ^ n378 ^ 1'b0 ;
  assign n13843 = ~n1851 & n13620 ;
  assign n13844 = n310 | n10327 ;
  assign n13845 = n11745 ^ n6248 ^ 1'b0 ;
  assign n13846 = ~n747 & n802 ;
  assign n13847 = n1655 ^ n1473 ^ 1'b0 ;
  assign n13848 = n6991 & ~n13847 ;
  assign n13849 = n3701 | n4537 ;
  assign n13850 = n13849 ^ n2484 ^ 1'b0 ;
  assign n13851 = n2997 & n13850 ;
  assign n13852 = ~n4550 & n7678 ;
  assign n13853 = n1987 ^ n129 ^ 1'b0 ;
  assign n13854 = ~n336 & n874 ;
  assign n13855 = n2400 & ~n9819 ;
  assign n13856 = n236 & n1712 ;
  assign n13857 = n13856 ^ n6721 ^ 1'b0 ;
  assign n13858 = n13857 ^ n11843 ^ 1'b0 ;
  assign n13859 = ~n13855 & n13858 ;
  assign n13860 = n5977 ^ n5241 ^ 1'b0 ;
  assign n13861 = ~n363 & n13860 ;
  assign n13862 = n13861 ^ n2083 ^ 1'b0 ;
  assign n13863 = n3014 & ~n13862 ;
  assign n13864 = n11281 & n13863 ;
  assign n13865 = n2564 | n6062 ;
  assign n13866 = n335 & n8718 ;
  assign n13867 = n13866 ^ n520 ^ 1'b0 ;
  assign n13868 = n9977 ^ n2885 ^ 1'b0 ;
  assign n13869 = n13868 ^ n2183 ^ 1'b0 ;
  assign n13870 = n13869 ^ n2941 ^ 1'b0 ;
  assign n13871 = n142 | n6028 ;
  assign n13872 = n3524 | n13871 ;
  assign n13873 = n2476 & n13872 ;
  assign n13874 = ~n5772 & n13873 ;
  assign n13875 = n643 | n13874 ;
  assign n13876 = n10086 ^ n2462 ^ 1'b0 ;
  assign n13877 = n11606 ^ n777 ^ 1'b0 ;
  assign n13878 = n8672 & ~n13877 ;
  assign n13879 = n2773 & ~n4865 ;
  assign n13880 = n4653 & ~n7056 ;
  assign n13881 = ~n4653 & n13880 ;
  assign n13882 = n4270 & ~n13881 ;
  assign n13883 = n197 & n769 ;
  assign n13884 = n5369 ^ n3665 ^ 1'b0 ;
  assign n13885 = n2300 ^ n1774 ^ 1'b0 ;
  assign n13886 = n113 & ~n12765 ;
  assign n13887 = n1344 & ~n13886 ;
  assign n13888 = n5743 | n8098 ;
  assign n13889 = n5743 ^ n5313 ^ 1'b0 ;
  assign n13890 = n9327 & n13889 ;
  assign n13891 = n7106 | n9649 ;
  assign n13892 = n10771 & n13891 ;
  assign n13893 = n5802 & ~n11239 ;
  assign n13894 = n2414 | n8579 ;
  assign n13895 = n3743 | n13894 ;
  assign n13896 = n1447 | n3812 ;
  assign n13897 = n215 | n1324 ;
  assign n13898 = n690 & ~n13897 ;
  assign n13899 = n4090 & ~n13898 ;
  assign n13900 = n13899 ^ n2049 ^ 1'b0 ;
  assign n13901 = n3180 | n9857 ;
  assign n13902 = n339 & n10436 ;
  assign n13903 = ~n7263 & n13902 ;
  assign n13904 = ( ~n2187 & n6133 ) | ( ~n2187 & n13816 ) | ( n6133 & n13816 ) ;
  assign n13905 = n10356 ^ n962 ^ 1'b0 ;
  assign n13906 = ~n216 & n13905 ;
  assign n13907 = n13606 ^ n3527 ^ 1'b0 ;
  assign n13908 = n5856 ^ n3570 ^ 1'b0 ;
  assign n13909 = n13908 ^ n12483 ^ 1'b0 ;
  assign n13910 = n13909 ^ n9895 ^ 1'b0 ;
  assign n13911 = n3406 | n13910 ;
  assign n13912 = n1562 | n11485 ;
  assign n13913 = n1833 & ~n13912 ;
  assign n13914 = n3095 | n9416 ;
  assign n13915 = n2377 & ~n13914 ;
  assign n13916 = n1476 & ~n12402 ;
  assign n13917 = n9036 & n13916 ;
  assign n13918 = n2272 | n13917 ;
  assign n13920 = n9370 ^ n5237 ^ 1'b0 ;
  assign n13919 = n4740 & n5862 ;
  assign n13921 = n13920 ^ n13919 ^ 1'b0 ;
  assign n13922 = n2041 & ~n5310 ;
  assign n13923 = ~n7439 & n13922 ;
  assign n13924 = n7714 | n10370 ;
  assign n13925 = ~n501 & n1543 ;
  assign n13926 = n101 & ~n7817 ;
  assign n13927 = n3901 & n13926 ;
  assign n13928 = n13927 ^ n169 ^ 1'b0 ;
  assign n13929 = ~n2880 & n13928 ;
  assign n13930 = ~n183 & n1329 ;
  assign n13931 = n10753 ^ n9215 ^ 1'b0 ;
  assign n13934 = n2533 & n3680 ;
  assign n13932 = n5891 & n7696 ;
  assign n13933 = n13932 ^ n4607 ^ 1'b0 ;
  assign n13935 = n13934 ^ n13933 ^ 1'b0 ;
  assign n13936 = n8464 ^ n8056 ^ 1'b0 ;
  assign n13937 = ~n13935 & n13936 ;
  assign n13938 = n813 | n2297 ;
  assign n13939 = n13938 ^ n3141 ^ 1'b0 ;
  assign n13940 = n10837 ^ n5470 ^ 1'b0 ;
  assign n13941 = n1257 | n13940 ;
  assign n13942 = ~x0 & n1017 ;
  assign n13943 = n13942 ^ n6238 ^ 1'b0 ;
  assign n13944 = n13943 ^ n339 ^ 1'b0 ;
  assign n13945 = ~n6368 & n13944 ;
  assign n13946 = n7116 ^ n321 ^ 1'b0 ;
  assign n13947 = n6269 | n12779 ;
  assign n13948 = n608 & ~n1935 ;
  assign n13949 = n7690 & n13948 ;
  assign n13950 = n1349 | n13766 ;
  assign n13951 = n13949 | n13950 ;
  assign n13952 = n5833 ^ n3687 ^ 1'b0 ;
  assign n13953 = n5169 ^ n340 ^ 1'b0 ;
  assign n13954 = n342 & ~n1895 ;
  assign n13955 = n9029 ^ n6403 ^ 1'b0 ;
  assign n13956 = n2244 | n13955 ;
  assign n13957 = n6447 | n13956 ;
  assign n13959 = n2159 & n7112 ;
  assign n13960 = ~n5089 & n13959 ;
  assign n13958 = n2900 & ~n5741 ;
  assign n13961 = n13960 ^ n13958 ^ 1'b0 ;
  assign n13962 = n1104 & ~n13961 ;
  assign n13963 = n6519 ^ n2144 ^ 1'b0 ;
  assign n13964 = n4869 ^ n1545 ^ 1'b0 ;
  assign n13967 = ~n3719 & n5263 ;
  assign n13968 = n13967 ^ x5 ^ 1'b0 ;
  assign n13965 = n1039 | n6586 ;
  assign n13966 = n13965 ^ n1865 ^ 1'b0 ;
  assign n13969 = n13968 ^ n13966 ^ 1'b0 ;
  assign n13970 = n8829 & ~n13969 ;
  assign n13971 = n11360 ^ n5649 ^ 1'b0 ;
  assign n13972 = n7786 & ~n7845 ;
  assign n13973 = n6389 | n13972 ;
  assign n13974 = n3095 ^ n1027 ^ 1'b0 ;
  assign n13975 = n1904 & n13974 ;
  assign n13976 = ~n2433 & n13975 ;
  assign n13977 = n142 & ~n594 ;
  assign n13978 = ~n5428 & n13977 ;
  assign n13979 = n13976 & n13978 ;
  assign n13980 = n3704 & n9151 ;
  assign n13981 = n13980 ^ n2929 ^ 1'b0 ;
  assign n13982 = n13981 ^ n3868 ^ 1'b0 ;
  assign n13983 = n5610 & ~n13982 ;
  assign n13984 = n3947 | n13983 ;
  assign n13985 = n769 & n5208 ;
  assign n13986 = ( n7909 & ~n7968 ) | ( n7909 & n13985 ) | ( ~n7968 & n13985 ) ;
  assign n13987 = n2362 ^ n1559 ^ 1'b0 ;
  assign n13988 = n11872 & n13987 ;
  assign n13989 = n2584 & n13988 ;
  assign n13990 = n13989 ^ n9208 ^ 1'b0 ;
  assign n13991 = n6475 ^ n1992 ^ 1'b0 ;
  assign n13992 = ~n12310 & n13991 ;
  assign n13993 = n13992 ^ n7301 ^ 1'b0 ;
  assign n13994 = n4485 & ~n13993 ;
  assign n13995 = n9304 ^ n2449 ^ 1'b0 ;
  assign n13996 = ~n310 & n13995 ;
  assign n13997 = n13996 ^ n4003 ^ 1'b0 ;
  assign n13998 = n13997 ^ n12241 ^ 1'b0 ;
  assign n13999 = n11192 & n13998 ;
  assign n14001 = n2074 & n4251 ;
  assign n14000 = n2556 & n3761 ;
  assign n14002 = n14001 ^ n14000 ^ 1'b0 ;
  assign n14003 = n14002 ^ n8156 ^ n2311 ;
  assign n14004 = n9161 ^ n4935 ^ 1'b0 ;
  assign n14005 = ~n13324 & n14004 ;
  assign n14006 = ~n3034 & n8775 ;
  assign n14007 = n904 & ~n14006 ;
  assign n14029 = n193 & ~n2426 ;
  assign n14030 = n2426 & n14029 ;
  assign n14031 = ~n5542 & n14030 ;
  assign n14032 = ~n4072 & n14031 ;
  assign n14033 = n14032 ^ n553 ^ 1'b0 ;
  assign n14008 = n5106 & ~n6933 ;
  assign n14009 = n6933 & n14008 ;
  assign n14010 = n9053 & ~n14009 ;
  assign n14011 = n122 & ~n7829 ;
  assign n14012 = ~n122 & n14011 ;
  assign n14013 = n810 & n2441 ;
  assign n14014 = n14012 & n14013 ;
  assign n14015 = n17 & ~n179 ;
  assign n14016 = n48 | n404 ;
  assign n14017 = n404 & ~n14016 ;
  assign n14018 = n14015 | n14017 ;
  assign n14019 = n14015 & ~n14018 ;
  assign n14020 = ~x8 & n2236 ;
  assign n14021 = n14019 & n14020 ;
  assign n14022 = n2348 & ~n14021 ;
  assign n14023 = n86 & ~n1688 ;
  assign n14024 = ~n86 & n14023 ;
  assign n14025 = n14022 | n14024 ;
  assign n14026 = n14014 & ~n14025 ;
  assign n14027 = n14010 & ~n14026 ;
  assign n14028 = ~n14010 & n14027 ;
  assign n14034 = n14033 ^ n14028 ^ 1'b0 ;
  assign n14035 = n2637 & n14034 ;
  assign n14036 = n11678 ^ n2151 ^ 1'b0 ;
  assign n14043 = n9682 ^ n1002 ^ 1'b0 ;
  assign n14044 = n12078 | n14043 ;
  assign n14038 = n1599 & n4090 ;
  assign n14039 = ~n2879 & n14038 ;
  assign n14040 = n1790 & n14039 ;
  assign n14041 = n14040 ^ n9340 ^ 1'b0 ;
  assign n14042 = n7696 & ~n14041 ;
  assign n14037 = n144 ^ n122 ^ 1'b0 ;
  assign n14045 = n14044 ^ n14042 ^ n14037 ;
  assign n14046 = ~n740 & n7442 ;
  assign n14047 = n14046 ^ n11870 ^ 1'b0 ;
  assign n14048 = n3693 ^ n628 ^ 1'b0 ;
  assign n14049 = ~n1118 & n14048 ;
  assign n14050 = n14047 & n14049 ;
  assign n14051 = n107 | n10882 ;
  assign n14052 = n14051 ^ n1581 ^ 1'b0 ;
  assign n14053 = n5322 & ~n7034 ;
  assign n14054 = n9409 ^ n107 ^ 1'b0 ;
  assign n14055 = ~n1015 & n14054 ;
  assign n14056 = n9808 & ~n11036 ;
  assign n14057 = n1854 & ~n11324 ;
  assign n14058 = n9026 ^ n2254 ^ 1'b0 ;
  assign n14059 = ~n12525 & n14058 ;
  assign n14060 = n14059 ^ n2624 ^ 1'b0 ;
  assign n14061 = n10924 ^ n4981 ^ 1'b0 ;
  assign n14062 = ~n14060 & n14061 ;
  assign n14063 = n11389 ^ n2599 ^ 1'b0 ;
  assign n14064 = n9764 ^ n6644 ^ 1'b0 ;
  assign n14065 = n9074 ^ n5355 ^ 1'b0 ;
  assign n14066 = n5800 | n14065 ;
  assign n14067 = n9696 | n14066 ;
  assign n14068 = n343 | n11671 ;
  assign n14069 = n13710 ^ n10194 ^ 1'b0 ;
  assign n14070 = n2676 ^ n814 ^ 1'b0 ;
  assign n14071 = n1622 | n14070 ;
  assign n14072 = n6297 & n6876 ;
  assign n14073 = n472 & ~n7741 ;
  assign n14074 = n8278 | n11025 ;
  assign n14075 = n406 | n4299 ;
  assign n14076 = n7090 | n14075 ;
  assign n14077 = n9492 & ~n14076 ;
  assign n14078 = ~n12175 & n14077 ;
  assign n14079 = n2222 & n5532 ;
  assign n14080 = n9767 & n14079 ;
  assign n14081 = n6376 & n14080 ;
  assign n14082 = n14081 ^ n1652 ^ 1'b0 ;
  assign n14083 = n8998 | n11967 ;
  assign n14084 = n14083 ^ n1691 ^ 1'b0 ;
  assign n14085 = n6618 ^ n760 ^ 1'b0 ;
  assign n14086 = n5825 ^ n128 ^ 1'b0 ;
  assign n14087 = n14085 | n14086 ;
  assign n14088 = n14087 ^ n3366 ^ 1'b0 ;
  assign n14089 = n8891 ^ n1508 ^ 1'b0 ;
  assign n14090 = n8329 & n12304 ;
  assign n14091 = n14089 & n14090 ;
  assign n14092 = n56 & n83 ;
  assign n14093 = n12180 ^ n9210 ^ 1'b0 ;
  assign n14094 = n1073 | n1804 ;
  assign n14095 = ~n1825 & n14094 ;
  assign n14096 = n13073 ^ n9175 ^ 1'b0 ;
  assign n14097 = n11703 ^ n2032 ^ 1'b0 ;
  assign n14098 = ~n8276 & n14097 ;
  assign n14099 = n2551 & n9461 ;
  assign n14100 = n8352 & n14099 ;
  assign n14101 = n14100 ^ n1342 ^ 1'b0 ;
  assign n14102 = n14098 & ~n14101 ;
  assign n14105 = ~x0 & n4646 ;
  assign n14103 = n1112 & ~n8488 ;
  assign n14104 = n8320 & n14103 ;
  assign n14106 = n14105 ^ n14104 ^ 1'b0 ;
  assign n14107 = n3559 | n4959 ;
  assign n14108 = n14106 & ~n14107 ;
  assign n14109 = ~n2275 & n2504 ;
  assign n14110 = n6935 & n14109 ;
  assign n14111 = n14110 ^ n2745 ^ 1'b0 ;
  assign n14112 = n14111 ^ n1959 ^ 1'b0 ;
  assign n14113 = n6200 ^ n4626 ^ 1'b0 ;
  assign n14114 = n1732 | n14113 ;
  assign n14115 = n1121 & n14114 ;
  assign n14116 = n1186 & ~n12060 ;
  assign n14117 = n14116 ^ n4538 ^ 1'b0 ;
  assign n14118 = n3014 & ~n14117 ;
  assign n14119 = n2533 & n9918 ;
  assign n14120 = n14118 & n14119 ;
  assign n14124 = n4379 | n5663 ;
  assign n14125 = n14124 ^ n8988 ^ 1'b0 ;
  assign n14121 = ~n3855 & n5256 ;
  assign n14122 = n14121 ^ n3023 ^ 1'b0 ;
  assign n14123 = n5126 & n14122 ;
  assign n14126 = n14125 ^ n14123 ^ n4529 ;
  assign n14127 = n2531 & ~n4855 ;
  assign n14128 = n6571 ^ n1710 ^ 1'b0 ;
  assign n14129 = n14127 & ~n14128 ;
  assign n14130 = n2929 ^ n501 ^ 1'b0 ;
  assign n14131 = ~n229 & n14130 ;
  assign n14132 = n9275 & ~n14131 ;
  assign n14133 = n14132 ^ n2480 ^ 1'b0 ;
  assign n14134 = n7034 ^ n878 ^ 1'b0 ;
  assign n14135 = n5162 & n14134 ;
  assign n14137 = ~n3134 & n3706 ;
  assign n14138 = ~n1810 & n14137 ;
  assign n14139 = n14138 ^ n2159 ^ 1'b0 ;
  assign n14140 = n5121 | n14139 ;
  assign n14136 = n5882 & n11915 ;
  assign n14141 = n14140 ^ n14136 ^ 1'b0 ;
  assign n14142 = n4004 & ~n6307 ;
  assign n14143 = n14142 ^ n12654 ^ 1'b0 ;
  assign n14144 = ~n7870 & n11192 ;
  assign n14145 = n85 | n3116 ;
  assign n14146 = n4842 & ~n14145 ;
  assign n14147 = n4853 & ~n14146 ;
  assign n14148 = n5501 ^ n2501 ^ 1'b0 ;
  assign n14149 = n4618 & n13001 ;
  assign n14150 = ~n1927 & n9304 ;
  assign n14151 = n14150 ^ n6590 ^ 1'b0 ;
  assign n14152 = n14151 ^ n6212 ^ 1'b0 ;
  assign n14153 = n10435 ^ n10259 ^ 1'b0 ;
  assign n14154 = n7214 ^ n6220 ^ 1'b0 ;
  assign n14155 = ~n55 & n14154 ;
  assign n14156 = ~n10963 & n12967 ;
  assign n14157 = ~n14155 & n14156 ;
  assign n14158 = n12633 ^ n2676 ^ 1'b0 ;
  assign n14159 = n12902 ^ n7483 ^ 1'b0 ;
  assign n14160 = ~n8641 & n12529 ;
  assign n14161 = n6405 ^ n6186 ^ 1'b0 ;
  assign n14162 = n713 & n14161 ;
  assign n14163 = n359 & n2261 ;
  assign n14164 = ~n6855 & n14163 ;
  assign n14165 = n6348 & ~n14164 ;
  assign n14166 = n988 & n2021 ;
  assign n14167 = n8121 ^ n7968 ^ 1'b0 ;
  assign n14168 = n1192 & ~n14167 ;
  assign n14169 = n2178 | n14168 ;
  assign n14170 = n8966 ^ n2450 ^ 1'b0 ;
  assign n14174 = n5853 & n6349 ;
  assign n14175 = n14174 ^ n2523 ^ 1'b0 ;
  assign n14171 = n6160 ^ n727 ^ 1'b0 ;
  assign n14172 = n1081 & ~n14171 ;
  assign n14173 = ~n5369 & n14172 ;
  assign n14176 = n14175 ^ n14173 ^ 1'b0 ;
  assign n14177 = ~n3063 & n14176 ;
  assign n14178 = n7319 ^ n1019 ^ 1'b0 ;
  assign n14179 = n6421 & ~n14178 ;
  assign n14180 = n6184 ^ n625 ^ 1'b0 ;
  assign n14181 = n14179 & n14180 ;
  assign n14182 = n4976 & n14181 ;
  assign n14183 = ~n2948 & n10829 ;
  assign n14184 = n14183 ^ n12213 ^ 1'b0 ;
  assign n14186 = n551 & n1060 ;
  assign n14185 = ~n2314 & n4760 ;
  assign n14187 = n14186 ^ n14185 ^ 1'b0 ;
  assign n14188 = n2725 | n4163 ;
  assign n14189 = n14188 ^ n14171 ^ 1'b0 ;
  assign n14190 = n13935 & ~n14189 ;
  assign n14191 = n2747 ^ n1814 ^ 1'b0 ;
  assign n14192 = n8523 & n14191 ;
  assign n14193 = n862 & n11067 ;
  assign n14194 = ~n9966 & n14193 ;
  assign n14199 = ~n2059 & n3653 ;
  assign n14200 = ~n3279 & n14199 ;
  assign n14195 = n462 | n5425 ;
  assign n14196 = n14195 ^ n1159 ^ 1'b0 ;
  assign n14197 = n4671 | n14196 ;
  assign n14198 = n5495 & ~n14197 ;
  assign n14201 = n14200 ^ n14198 ^ 1'b0 ;
  assign n14202 = n800 & ~n14201 ;
  assign n14203 = n11898 ^ n3529 ^ 1'b0 ;
  assign n14204 = n14203 ^ n12281 ^ n2578 ;
  assign n14205 = n767 | n5444 ;
  assign n14206 = n14205 ^ n3916 ^ 1'b0 ;
  assign n14207 = n14206 ^ n246 ^ 1'b0 ;
  assign n14208 = n8441 | n11289 ;
  assign n14209 = ~n5431 & n9114 ;
  assign n14210 = n1687 & n9571 ;
  assign n14211 = ~n847 & n6188 ;
  assign n14212 = ~n3814 & n14211 ;
  assign n14213 = n14212 ^ n4927 ^ 1'b0 ;
  assign n14214 = ~n14086 & n14213 ;
  assign n14215 = ~n185 & n14214 ;
  assign n14216 = n8973 ^ n5041 ^ 1'b0 ;
  assign n14217 = ~n10429 & n14216 ;
  assign n14218 = n113 & ~n5455 ;
  assign n14219 = n11233 ^ n2551 ^ 1'b0 ;
  assign n14220 = n14219 ^ x2 ^ 1'b0 ;
  assign n14221 = n6476 & ~n14220 ;
  assign n14222 = n234 | n2604 ;
  assign n14223 = n13541 & ~n14222 ;
  assign n14224 = ~n14221 & n14223 ;
  assign n14225 = n520 | n1835 ;
  assign n14226 = n14225 ^ n2351 ^ 1'b0 ;
  assign n14227 = ~n1743 & n14226 ;
  assign n14228 = n7904 & n14227 ;
  assign n14229 = ~n6755 & n8407 ;
  assign n14230 = n12223 ^ n7654 ^ 1'b0 ;
  assign n14231 = n4078 | n14230 ;
  assign n14232 = n2348 & n2929 ;
  assign n14233 = n10050 & ~n14232 ;
  assign n14234 = n4227 | n9122 ;
  assign n14235 = ~n11948 & n14234 ;
  assign n14236 = ( n3868 & ~n5808 ) | ( n3868 & n13874 ) | ( ~n5808 & n13874 ) ;
  assign n14237 = n1194 & n1879 ;
  assign n14238 = ~n14236 & n14237 ;
  assign n14239 = n3125 & ~n14238 ;
  assign n14240 = n14239 ^ n3567 ^ 1'b0 ;
  assign n14241 = n3262 & ~n13870 ;
  assign n14242 = n624 ^ n191 ^ 1'b0 ;
  assign n14243 = n5110 & n14242 ;
  assign n14244 = n6889 & n11778 ;
  assign n14245 = n14244 ^ n5013 ^ 1'b0 ;
  assign n14246 = ~n7464 & n8461 ;
  assign n14247 = ~n3229 & n12468 ;
  assign n14248 = ~n13220 & n14247 ;
  assign n14249 = n8969 ^ n6102 ^ 1'b0 ;
  assign n14250 = n8861 | n11950 ;
  assign n14251 = n443 | n14250 ;
  assign n14252 = n8946 ^ n4920 ^ 1'b0 ;
  assign n14253 = n5844 & ~n14252 ;
  assign n14254 = n259 & n14179 ;
  assign n14255 = ~n5280 & n14254 ;
  assign n14256 = n3493 & n9572 ;
  assign n14257 = n2517 ^ n2456 ^ 1'b0 ;
  assign n14258 = n7096 & ~n14257 ;
  assign n14259 = n14258 ^ n2619 ^ 1'b0 ;
  assign n14260 = n3845 | n4093 ;
  assign n14261 = n6090 & ~n11105 ;
  assign n14262 = ~n4712 & n9210 ;
  assign n14263 = n8054 ^ n1893 ^ 1'b0 ;
  assign n14264 = n4700 | n14263 ;
  assign n14265 = n11195 ^ n506 ^ 1'b0 ;
  assign n14266 = n5726 ^ n4774 ^ 1'b0 ;
  assign n14267 = n14265 & ~n14266 ;
  assign n14268 = n12717 & n14267 ;
  assign n14269 = n2721 | n9122 ;
  assign n14270 = n8419 ^ n7497 ^ n6209 ;
  assign n14271 = n4256 ^ n1070 ^ n536 ;
  assign n14272 = n1174 & n5161 ;
  assign n14273 = n12761 & ~n14272 ;
  assign n14274 = ~n14271 & n14273 ;
  assign n14275 = n9327 ^ n1912 ^ 1'b0 ;
  assign n14276 = n5562 & n7572 ;
  assign n14277 = n14276 ^ n7144 ^ 1'b0 ;
  assign n14278 = n12223 ^ n4121 ^ n471 ;
  assign n14279 = ~n2933 & n3226 ;
  assign n14295 = ~n357 & n405 ;
  assign n14296 = n38 & n336 ;
  assign n14297 = ~n38 & n14296 ;
  assign n14298 = n14295 & ~n14297 ;
  assign n14299 = ~n12310 & n14298 ;
  assign n14300 = ~n56 & n14299 ;
  assign n14280 = ~n192 & n287 ;
  assign n14281 = ~n287 & n14280 ;
  assign n14282 = n2022 & n14281 ;
  assign n14283 = ~n2022 & n14282 ;
  assign n14284 = n1230 & n14283 ;
  assign n14285 = n269 & ~n307 ;
  assign n14286 = ~n269 & n14285 ;
  assign n14287 = n195 & n14286 ;
  assign n14288 = n4683 | n14287 ;
  assign n14289 = n14287 & ~n14288 ;
  assign n14290 = n14284 & ~n14289 ;
  assign n14291 = ~n14284 & n14290 ;
  assign n14292 = n250 & ~n10917 ;
  assign n14293 = ~n250 & n14292 ;
  assign n14294 = n14291 | n14293 ;
  assign n14301 = n14300 ^ n14294 ^ 1'b0 ;
  assign n14302 = n7706 ^ n7147 ^ 1'b0 ;
  assign n14303 = ~n7926 & n14302 ;
  assign n14304 = n5010 & n14303 ;
  assign n14305 = n2659 ^ n1314 ^ 1'b0 ;
  assign n14306 = n2448 ^ n1225 ^ 1'b0 ;
  assign n14307 = n14306 ^ n246 ^ 1'b0 ;
  assign n14308 = n11826 ^ n958 ^ 1'b0 ;
  assign n14309 = ~n14307 & n14308 ;
  assign n14310 = n163 & ~n2131 ;
  assign n14311 = n471 & n7924 ;
  assign n14312 = n14311 ^ n907 ^ 1'b0 ;
  assign n14313 = n12645 ^ n8525 ^ 1'b0 ;
  assign n14314 = n13029 ^ n113 ^ 1'b0 ;
  assign n14315 = n850 | n14314 ;
  assign n14316 = n2432 ^ n1804 ^ 1'b0 ;
  assign n14317 = n5983 | n14316 ;
  assign n14318 = n6238 ^ n1884 ^ 1'b0 ;
  assign n14319 = n2228 & n14318 ;
  assign n14320 = ~n9750 & n14319 ;
  assign n14321 = n3709 & n14320 ;
  assign n14322 = n174 | n14321 ;
  assign n14323 = n14317 | n14322 ;
  assign n14324 = n5416 ^ n3771 ^ n1506 ;
  assign n14325 = n14324 ^ n5626 ^ 1'b0 ;
  assign n14326 = n2661 | n2953 ;
  assign n14327 = n6210 ^ n3706 ^ 1'b0 ;
  assign n14328 = ~n12167 & n14327 ;
  assign n14329 = n14326 & n14328 ;
  assign n14330 = n812 & n1537 ;
  assign n14331 = n14330 ^ n5467 ^ 1'b0 ;
  assign n14332 = n330 & n13493 ;
  assign n14333 = n4322 & n14332 ;
  assign n14338 = n1226 & n3183 ;
  assign n14339 = ~n4206 & n14338 ;
  assign n14334 = n4407 & ~n6028 ;
  assign n14335 = ~n1865 & n5046 ;
  assign n14336 = n14334 & n14335 ;
  assign n14337 = n7077 & ~n14336 ;
  assign n14340 = n14339 ^ n14337 ^ 1'b0 ;
  assign n14341 = ~n14333 & n14340 ;
  assign n14342 = n14341 ^ n1039 ^ 1'b0 ;
  assign n14343 = n14331 | n14342 ;
  assign n14344 = ~n2460 & n3290 ;
  assign n14345 = n2846 | n14344 ;
  assign n14346 = n14345 ^ n12747 ^ 1'b0 ;
  assign n14347 = n382 | n8373 ;
  assign n14348 = n3203 | n14347 ;
  assign n14349 = n1152 & ~n8532 ;
  assign n14350 = n7056 ^ n3344 ^ 1'b0 ;
  assign n14351 = ( n205 & n412 ) | ( n205 & n13733 ) | ( n412 & n13733 ) ;
  assign n14352 = n10790 & ~n14351 ;
  assign n14353 = n281 & n14352 ;
  assign n14354 = n14353 ^ n11948 ^ 1'b0 ;
  assign n14355 = ~n8349 & n14354 ;
  assign n14356 = n11738 | n12284 ;
  assign n14357 = n4700 & ~n8448 ;
  assign n14358 = n1329 & n14357 ;
  assign n14359 = n11843 ^ n4432 ^ 1'b0 ;
  assign n14360 = n6690 | n14359 ;
  assign n14364 = x8 & n581 ;
  assign n14365 = ~x8 & n14364 ;
  assign n14366 = n14365 ^ n2509 ^ 1'b0 ;
  assign n14361 = n441 | n5369 ;
  assign n14362 = n5369 & ~n14361 ;
  assign n14363 = n12912 | n14362 ;
  assign n14367 = n14366 ^ n14363 ^ 1'b0 ;
  assign n14368 = n7449 ^ n1771 ^ 1'b0 ;
  assign n14369 = n3487 & ~n14368 ;
  assign n14370 = n2321 | n10479 ;
  assign n14371 = n7924 & n10652 ;
  assign n14372 = ~n1129 & n11680 ;
  assign n14379 = ~n1562 & n4525 ;
  assign n14380 = n14379 ^ n104 ^ 1'b0 ;
  assign n14381 = n1577 & ~n5366 ;
  assign n14382 = n14381 ^ n5520 ^ 1'b0 ;
  assign n14383 = n14380 | n14382 ;
  assign n14373 = n632 & n7401 ;
  assign n14374 = n14373 ^ n3836 ^ 1'b0 ;
  assign n14375 = ~n3896 & n14374 ;
  assign n14376 = n690 & n14375 ;
  assign n14377 = n14376 ^ n116 ^ 1'b0 ;
  assign n14378 = n1143 | n14377 ;
  assign n14384 = n14383 ^ n14378 ^ 1'b0 ;
  assign n14385 = ~x5 & n14384 ;
  assign n14386 = n10736 & n13312 ;
  assign n14387 = ~n200 & n2134 ;
  assign n14388 = n986 ^ n60 ^ 1'b0 ;
  assign n14389 = ~n820 & n14388 ;
  assign n14390 = n14389 ^ n8523 ^ 1'b0 ;
  assign n14391 = n14387 & ~n14390 ;
  assign n14392 = ~x1 & n2420 ;
  assign n14393 = n5401 | n5826 ;
  assign n14394 = n12435 ^ n6170 ^ 1'b0 ;
  assign n14395 = n905 | n10583 ;
  assign n14396 = n2813 | n7124 ;
  assign n14397 = n8582 & n10327 ;
  assign n14398 = n14120 ^ n5538 ^ 1'b0 ;
  assign n14399 = n8993 & n9499 ;
  assign n14400 = ~n11525 & n14399 ;
  assign n14401 = n7582 & n12408 ;
  assign n14402 = n848 & ~n2637 ;
  assign n14403 = n14402 ^ n378 ^ 1'b0 ;
  assign n14404 = n7523 & ~n14403 ;
  assign n14409 = n1127 & ~n4346 ;
  assign n14405 = n1372 | n8226 ;
  assign n14406 = n5456 & n9009 ;
  assign n14407 = n14405 & n14406 ;
  assign n14408 = n14407 ^ n11970 ^ 1'b0 ;
  assign n14410 = n14409 ^ n14408 ^ 1'b0 ;
  assign n14411 = n1849 & n5741 ;
  assign n14412 = n1789 & ~n14411 ;
  assign n14413 = n14412 ^ n9793 ^ n9422 ;
  assign n14414 = n3178 & n14413 ;
  assign n14415 = n1195 & ~n3542 ;
  assign n14417 = n1688 | n6687 ;
  assign n14416 = n3068 & ~n9695 ;
  assign n14418 = n14417 ^ n14416 ^ n11516 ;
  assign n14419 = n14088 ^ n6740 ^ 1'b0 ;
  assign n14420 = ~n2752 & n14419 ;
  assign n14421 = n7060 ^ n3664 ^ 1'b0 ;
  assign n14422 = n3309 | n14421 ;
  assign n14423 = n14309 & n14422 ;
  assign n14424 = n2487 | n8665 ;
  assign n14425 = n10915 ^ n10046 ^ 1'b0 ;
  assign n14426 = ~n469 & n7111 ;
  assign n14427 = n14426 ^ n6644 ^ 1'b0 ;
  assign n14433 = n6349 & ~n10105 ;
  assign n14428 = n5024 ^ n3459 ^ 1'b0 ;
  assign n14429 = ~n940 & n14428 ;
  assign n14430 = ~n8306 & n8403 ;
  assign n14431 = n14430 ^ n5334 ^ 1'b0 ;
  assign n14432 = n14429 & n14431 ;
  assign n14434 = n14433 ^ n14432 ^ 1'b0 ;
  assign n14435 = n10058 & n14434 ;
  assign n14436 = n12222 ^ n19 ^ 1'b0 ;
  assign n14437 = n1348 & ~n1613 ;
  assign n14438 = n14437 ^ n3532 ^ 1'b0 ;
  assign n14439 = n14438 ^ n3928 ^ 1'b0 ;
  assign n14440 = n14439 ^ n1984 ^ 1'b0 ;
  assign n14441 = n7136 ^ n2684 ^ 1'b0 ;
  assign n14442 = n13344 & n14441 ;
  assign n14443 = ~n14440 & n14442 ;
  assign n14444 = n3341 ^ n3068 ^ 1'b0 ;
  assign n14445 = n14444 ^ n7043 ^ 1'b0 ;
  assign n14446 = n6200 ^ n3490 ^ 1'b0 ;
  assign n14447 = n297 & n14446 ;
  assign n14448 = n14447 ^ n13260 ^ 1'b0 ;
  assign n14449 = n12181 ^ n203 ^ 1'b0 ;
  assign n14450 = n1263 & n4013 ;
  assign n14451 = n3389 ^ n3264 ^ 1'b0 ;
  assign n14452 = n7208 | n14451 ;
  assign n14453 = n2476 & ~n3395 ;
  assign n14454 = n14452 & n14453 ;
  assign n14455 = ~n14450 & n14454 ;
  assign n14456 = n14449 & n14455 ;
  assign n14457 = n14456 ^ n13252 ^ 1'b0 ;
  assign n14458 = n12993 | n14400 ;
  assign n14461 = n1597 | n5197 ;
  assign n14462 = n243 & ~n14461 ;
  assign n14459 = ~n520 & n9086 ;
  assign n14460 = ~n9934 & n14459 ;
  assign n14463 = n14462 ^ n14460 ^ n1975 ;
  assign n14464 = n12663 ^ n758 ^ 1'b0 ;
  assign n14465 = n4275 & ~n5169 ;
  assign n14466 = n14464 & n14465 ;
  assign n14467 = n5099 & ~n14466 ;
  assign n14468 = n14467 ^ n5894 ^ 1'b0 ;
  assign n14469 = n11728 & n14468 ;
  assign n14470 = n13206 ^ n1756 ^ 1'b0 ;
  assign n14471 = n7487 & ~n8819 ;
  assign n14472 = n5302 ^ n263 ^ 1'b0 ;
  assign n14473 = ~n328 & n14472 ;
  assign n14474 = n1250 & ~n8135 ;
  assign n14475 = n4404 ^ n627 ^ 1'b0 ;
  assign n14476 = n3335 & n14475 ;
  assign n14477 = n8398 ^ n4979 ^ 1'b0 ;
  assign n14478 = ~n4182 & n14477 ;
  assign n14479 = ~n133 & n2626 ;
  assign n14480 = n4838 ^ n2239 ^ 1'b0 ;
  assign n14481 = n4077 & n14480 ;
  assign n14482 = n14479 | n14481 ;
  assign n14483 = ( n1444 & n6244 ) | ( n1444 & ~n14482 ) | ( n6244 & ~n14482 ) ;
  assign n14484 = n2776 & ~n6463 ;
  assign n14485 = n6296 & ~n14484 ;
  assign n14486 = ~n6296 & n14485 ;
  assign n14487 = n133 | n5570 ;
  assign n14488 = n9211 | n14487 ;
  assign n14489 = n6246 ^ n3985 ^ 1'b0 ;
  assign n14490 = n3745 & ~n14489 ;
  assign n14491 = ~n6137 & n12868 ;
  assign n14492 = n3053 & ~n12431 ;
  assign n14493 = n3735 ^ n1469 ^ 1'b0 ;
  assign n14494 = ~n8203 & n14493 ;
  assign n14495 = n4426 & n14494 ;
  assign n14496 = n2569 & ~n4976 ;
  assign n14497 = n82 & ~n1165 ;
  assign n14498 = n14497 ^ n10486 ^ 1'b0 ;
  assign n14499 = n1934 & ~n2155 ;
  assign n14500 = n10641 & n14499 ;
  assign n14501 = n14500 ^ n12416 ^ 1'b0 ;
  assign n14502 = n2391 & ~n14501 ;
  assign n14503 = n1794 | n3767 ;
  assign n14504 = n1794 & ~n14503 ;
  assign n14505 = ~n3506 & n5258 ;
  assign n14506 = n14504 & n14505 ;
  assign n14507 = n2971 & n6880 ;
  assign n14508 = ~n6880 & n14507 ;
  assign n14509 = n13930 | n14508 ;
  assign n14510 = ~n1058 & n4853 ;
  assign n14511 = n14509 | n14510 ;
  assign n14512 = n14506 & ~n14511 ;
  assign n14513 = n123 | n5814 ;
  assign n14514 = n4774 & ~n9291 ;
  assign n14515 = ~n101 & n14514 ;
  assign n14516 = ( ~n2263 & n10390 ) | ( ~n2263 & n14515 ) | ( n10390 & n14515 ) ;
  assign n14517 = n6679 | n14516 ;
  assign n14519 = n7424 | n13017 ;
  assign n14518 = n812 & ~n3220 ;
  assign n14520 = n14519 ^ n14518 ^ 1'b0 ;
  assign n14521 = n9572 ^ n2489 ^ 1'b0 ;
  assign n14522 = n13389 & n14521 ;
  assign n14523 = ~n10798 & n14522 ;
  assign n14524 = n336 & n9655 ;
  assign n14525 = ~n1112 & n14524 ;
  assign n14526 = ~n2896 & n14525 ;
  assign n14527 = n7388 | n11224 ;
  assign n14528 = n14526 & ~n14527 ;
  assign n14529 = n8999 ^ n154 ^ 1'b0 ;
  assign n14530 = n1002 | n3423 ;
  assign n14531 = n14529 | n14530 ;
  assign n14532 = n8411 | n12385 ;
  assign n14533 = n4904 | n8233 ;
  assign n14534 = n14533 ^ n6748 ^ 1'b0 ;
  assign n14535 = n14534 ^ n7082 ^ 1'b0 ;
  assign n14536 = ( n520 & n1252 ) | ( n520 & n6008 ) | ( n1252 & n6008 ) ;
  assign n14537 = n11234 ^ n726 ^ 1'b0 ;
  assign n14538 = n7153 | n14537 ;
  assign n14539 = n2166 | n14538 ;
  assign n14540 = n612 & n4498 ;
  assign n14541 = n14540 ^ n1152 ^ 1'b0 ;
  assign n14542 = n86 & ~n1188 ;
  assign n14543 = n14542 ^ n299 ^ 1'b0 ;
  assign n14544 = n14543 ^ n4942 ^ 1'b0 ;
  assign n14545 = n2140 | n8004 ;
  assign n14546 = n14544 | n14545 ;
  assign n14547 = n9696 & n14546 ;
  assign n14548 = n3137 | n5265 ;
  assign n14549 = n14548 ^ n2933 ^ 1'b0 ;
  assign n14550 = n4180 ^ n353 ^ 1'b0 ;
  assign n14551 = ~n4966 & n14550 ;
  assign n14552 = n14551 ^ n9877 ^ 1'b0 ;
  assign n14553 = n4055 ^ n3764 ^ 1'b0 ;
  assign n14554 = ~n6071 & n14553 ;
  assign n14555 = n4523 & n7644 ;
  assign n14556 = ~n9890 & n14555 ;
  assign n14557 = ( n181 & ~n4570 ) | ( n181 & n7589 ) | ( ~n4570 & n7589 ) ;
  assign n14558 = n556 ^ n512 ^ 1'b0 ;
  assign n14559 = n14558 ^ n8439 ^ 1'b0 ;
  assign n14560 = n1587 & n11359 ;
  assign n14561 = n7455 ^ n281 ^ 1'b0 ;
  assign n14562 = n7483 ^ n575 ^ 1'b0 ;
  assign n14563 = ~n158 & n14562 ;
  assign n14564 = n5805 ^ n1096 ^ 1'b0 ;
  assign n14565 = n7696 ^ n2148 ^ 1'b0 ;
  assign n14566 = n6481 | n14565 ;
  assign n14567 = n336 & ~n14566 ;
  assign n14568 = n14567 ^ n12673 ^ 1'b0 ;
  assign n14569 = ~n709 & n12804 ;
  assign n14570 = ~n14551 & n14569 ;
  assign n14571 = n1110 & ~n4926 ;
  assign n14572 = n14571 ^ n5056 ^ n2939 ;
  assign n14573 = n12186 | n14572 ;
  assign n14574 = n185 & n3293 ;
  assign n14575 = n4341 & ~n5415 ;
  assign n14576 = n5415 & n14575 ;
  assign n14577 = n520 & ~n14576 ;
  assign n14578 = n4142 | n14577 ;
  assign n14579 = n14577 & ~n14578 ;
  assign n14580 = n10655 | n10943 ;
  assign n14581 = n10655 & ~n14580 ;
  assign n14582 = n14579 | n14581 ;
  assign n14583 = n14579 & ~n14582 ;
  assign n14584 = n6160 | n14583 ;
  assign n14585 = n14584 ^ n8739 ^ 1'b0 ;
  assign n14586 = n5666 | n14585 ;
  assign n14587 = ~n847 & n9284 ;
  assign n14588 = ~n163 & n1968 ;
  assign n14589 = n1529 & ~n9357 ;
  assign n14590 = n14589 ^ n1765 ^ 1'b0 ;
  assign n14591 = n14590 ^ n12075 ^ 1'b0 ;
  assign n14592 = ~n5913 & n6181 ;
  assign n14593 = n14592 ^ n7487 ^ 1'b0 ;
  assign n14594 = n13118 ^ n5317 ^ 1'b0 ;
  assign n14595 = ~n6187 & n14594 ;
  assign n14596 = n2542 | n6060 ;
  assign n14597 = n1756 & n14596 ;
  assign n14598 = ~n14596 & n14597 ;
  assign n14599 = n9482 ^ n5532 ^ 1'b0 ;
  assign n14600 = ~n14598 & n14599 ;
  assign n14601 = n6154 & ~n9049 ;
  assign n14602 = n14601 ^ n2109 ^ 1'b0 ;
  assign n14603 = n241 | n581 ;
  assign n14604 = n5778 | n5903 ;
  assign n14605 = n14604 ^ n1966 ^ 1'b0 ;
  assign n14606 = n5621 ^ n624 ^ n286 ;
  assign n14607 = ~n14605 & n14606 ;
  assign n14611 = n2011 | n7338 ;
  assign n14608 = n2107 ^ n1822 ^ 1'b0 ;
  assign n14609 = n14608 ^ n5193 ^ 1'b0 ;
  assign n14610 = n4584 & ~n14609 ;
  assign n14612 = n14611 ^ n14610 ^ 1'b0 ;
  assign n14613 = n2654 | n12193 ;
  assign n14614 = n2388 | n14613 ;
  assign n14615 = n14614 ^ n7216 ^ 1'b0 ;
  assign n14616 = ~n1991 & n14615 ;
  assign n14617 = n79 & n8307 ;
  assign n14618 = ~n935 & n1297 ;
  assign n14619 = n14617 | n14618 ;
  assign n14620 = n2491 | n13757 ;
  assign n14621 = n1166 & n7917 ;
  assign n14622 = n14621 ^ n325 ^ 1'b0 ;
  assign n14623 = n14622 ^ n6345 ^ 1'b0 ;
  assign n14624 = n1416 | n14623 ;
  assign n14625 = n11346 ^ n1684 ^ 1'b0 ;
  assign n14626 = n1260 & n5452 ;
  assign n14627 = ~n528 & n562 ;
  assign n14628 = ~n562 & n14627 ;
  assign n14629 = ~x3 & n14628 ;
  assign n14630 = n8071 & n14629 ;
  assign n14631 = n14626 & n14630 ;
  assign n14632 = n566 | n10561 ;
  assign n14633 = n566 & ~n14632 ;
  assign n14634 = n4076 & ~n14633 ;
  assign n14635 = n14633 & n14634 ;
  assign n14636 = n14631 | n14635 ;
  assign n14637 = n14631 & ~n14636 ;
  assign n14638 = n2790 & ~n14637 ;
  assign n14639 = ~n11019 & n14638 ;
  assign n14640 = ~n814 & n6439 ;
  assign n14641 = n2432 & n14640 ;
  assign n14642 = n14641 ^ n2079 ^ 1'b0 ;
  assign n14643 = n391 | n5797 ;
  assign n14644 = n14643 ^ n817 ^ 1'b0 ;
  assign n14645 = n2727 & n12948 ;
  assign n14646 = n5873 & ~n7551 ;
  assign n14648 = ~n4893 & n8652 ;
  assign n14647 = n7203 ^ n7107 ^ 1'b0 ;
  assign n14649 = n14648 ^ n14647 ^ 1'b0 ;
  assign n14650 = n12978 & n13208 ;
  assign n14651 = n5756 & n12242 ;
  assign n14652 = n618 | n10107 ;
  assign n14653 = n14652 ^ n4374 ^ 1'b0 ;
  assign n14654 = n12659 ^ n2067 ^ 1'b0 ;
  assign n14655 = n1929 | n6242 ;
  assign n14656 = n541 | n14655 ;
  assign n14657 = n14656 ^ n7683 ^ 1'b0 ;
  assign n14658 = n2074 & n5700 ;
  assign n14659 = ~n1332 & n14658 ;
  assign n14660 = ~n14131 & n14659 ;
  assign n14661 = n3533 | n13058 ;
  assign n14662 = n14661 ^ n161 ^ 1'b0 ;
  assign n14663 = n6871 | n7650 ;
  assign n14664 = n14663 ^ n11659 ^ 1'b0 ;
  assign n14665 = n9925 ^ n109 ^ 1'b0 ;
  assign n14666 = n64 & n1847 ;
  assign n14667 = n14666 ^ n3088 ^ 1'b0 ;
  assign n14668 = n6156 ^ n4779 ^ 1'b0 ;
  assign n14669 = n1125 & ~n14668 ;
  assign n14670 = n6816 ^ n3624 ^ 1'b0 ;
  assign n14671 = n14670 ^ n11528 ^ 1'b0 ;
  assign n14672 = n14669 & ~n14671 ;
  assign n14673 = n5819 | n13968 ;
  assign n14674 = n8505 & ~n14673 ;
  assign n14675 = ~n2752 & n9961 ;
  assign n14676 = n8357 ^ n456 ^ 1'b0 ;
  assign n14677 = n5858 | n6853 ;
  assign n14679 = n4872 & n5744 ;
  assign n14680 = ~n5642 & n14679 ;
  assign n14678 = ~n942 & n1362 ;
  assign n14681 = n14680 ^ n14678 ^ 1'b0 ;
  assign n14682 = n14681 ^ n7249 ^ 1'b0 ;
  assign n14683 = n2455 | n4870 ;
  assign n14684 = n13792 & ~n14683 ;
  assign n14685 = n6400 ^ n628 ^ 1'b0 ;
  assign n14686 = ~n3287 & n14685 ;
  assign n14687 = ~n8286 & n14686 ;
  assign n14688 = n14687 ^ n4403 ^ 1'b0 ;
  assign n14689 = ~x3 & n3917 ;
  assign n14690 = ~n1644 & n1834 ;
  assign n14691 = n14689 & ~n14690 ;
  assign n14692 = ~n1866 & n14691 ;
  assign n14693 = n186 & n5053 ;
  assign n14694 = n14693 ^ n6907 ^ 1'b0 ;
  assign n14695 = n14694 ^ n8358 ^ 1'b0 ;
  assign n14696 = n3394 & n14695 ;
  assign n14697 = n6325 ^ n2348 ^ 1'b0 ;
  assign n14698 = ~n5481 & n14697 ;
  assign n14699 = ~n14696 & n14698 ;
  assign n14701 = n3333 & n13693 ;
  assign n14700 = n11192 & n14664 ;
  assign n14702 = n14701 ^ n14700 ^ 1'b0 ;
  assign n14703 = n1505 ^ n89 ^ 1'b0 ;
  assign n14704 = n5154 & n14703 ;
  assign n14705 = n5666 | n14704 ;
  assign n14706 = n14705 ^ n295 ^ 1'b0 ;
  assign n14707 = n3464 | n14706 ;
  assign n14708 = n12673 & ~n14707 ;
  assign n14709 = n13285 ^ n2730 ^ 1'b0 ;
  assign n14710 = n3219 ^ n1708 ^ 1'b0 ;
  assign n14712 = n4227 ^ n2298 ^ 1'b0 ;
  assign n14711 = n1396 | n4060 ;
  assign n14713 = n14712 ^ n14711 ^ 1'b0 ;
  assign n14714 = n14713 ^ n2348 ^ 1'b0 ;
  assign n14715 = n14714 ^ n2125 ^ 1'b0 ;
  assign n14718 = n13453 ^ n286 ^ 1'b0 ;
  assign n14719 = n4965 & n14718 ;
  assign n14717 = ( n3329 & n4961 ) | ( n3329 & n9274 ) | ( n4961 & n9274 ) ;
  assign n14716 = ~n3584 & n4469 ;
  assign n14720 = n14719 ^ n14717 ^ n14716 ;
  assign n14721 = n906 | n9659 ;
  assign n14722 = n1922 | n9849 ;
  assign n14723 = n3497 & ~n14722 ;
  assign n14724 = n5447 | n14723 ;
  assign n14725 = n9539 ^ n1480 ^ 1'b0 ;
  assign n14726 = n4369 ^ n860 ^ 1'b0 ;
  assign n14727 = n2526 & n14726 ;
  assign n14728 = n9391 ^ n570 ^ 1'b0 ;
  assign n14729 = ~n3990 & n14728 ;
  assign n14730 = n14729 ^ n5387 ^ 1'b0 ;
  assign n14731 = n1742 & ~n5545 ;
  assign n14732 = ~n5095 & n14731 ;
  assign n14733 = n10663 ^ n8761 ^ 1'b0 ;
  assign n14734 = n7475 ^ n284 ^ 1'b0 ;
  assign n14735 = n14734 ^ n6691 ^ 1'b0 ;
  assign n14736 = n5462 | n5831 ;
  assign n14740 = n11833 ^ n2747 ^ 1'b0 ;
  assign n14737 = ( ~n263 & n726 ) | ( ~n263 & n1050 ) | ( n726 & n1050 ) ;
  assign n14738 = n5663 ^ n1260 ^ 1'b0 ;
  assign n14739 = n14737 | n14738 ;
  assign n14741 = n14740 ^ n14739 ^ 1'b0 ;
  assign n14742 = ~n2704 & n3171 ;
  assign n14743 = n14742 ^ n7394 ^ 1'b0 ;
  assign n14744 = ~n1165 & n14743 ;
  assign n14745 = n3398 & ~n5880 ;
  assign n14746 = n10920 ^ n5121 ^ 1'b0 ;
  assign n14747 = ~n5292 & n7023 ;
  assign n14748 = n14746 & ~n14747 ;
  assign n14749 = ~n4365 & n5364 ;
  assign n14750 = n14749 ^ n6235 ^ 1'b0 ;
  assign n14751 = n958 & ~n7450 ;
  assign n14752 = n14751 ^ n4367 ^ 1'b0 ;
  assign n14753 = n14750 | n14752 ;
  assign n14754 = n14753 ^ n11775 ^ 1'b0 ;
  assign n14755 = n5070 | n14754 ;
  assign n14756 = n14755 ^ n286 ^ 1'b0 ;
  assign n14757 = n1368 & ~n14756 ;
  assign n14758 = ~n2038 & n2302 ;
  assign n14759 = n14758 ^ n7630 ^ 1'b0 ;
  assign n14760 = n9692 ^ x0 ^ 1'b0 ;
  assign n14761 = n14759 & ~n14760 ;
  assign n14762 = n14761 ^ n1926 ^ 1'b0 ;
  assign n14763 = n7988 ^ n622 ^ 1'b0 ;
  assign n14764 = ~n14762 & n14763 ;
  assign n14765 = ~n1895 & n9750 ;
  assign n14766 = ~n2532 & n12561 ;
  assign n14767 = n1880 & ~n13803 ;
  assign n14768 = n4875 & n6349 ;
  assign n14769 = n1701 & ~n10546 ;
  assign n14770 = ~n6265 & n14769 ;
  assign n14771 = n6383 & n7625 ;
  assign n14772 = n813 & ~n6894 ;
  assign n14773 = n3378 | n5459 ;
  assign n14774 = n5362 & ~n14773 ;
  assign n14775 = n7148 & ~n14774 ;
  assign n14776 = n14775 ^ n3503 ^ 1'b0 ;
  assign n14777 = ~n86 & n14776 ;
  assign n14778 = n7999 ^ n1388 ^ 1'b0 ;
  assign n14779 = n796 | n14778 ;
  assign n14780 = n2947 & ~n5780 ;
  assign n14781 = n823 & ~n14780 ;
  assign n14782 = n14781 ^ n11407 ^ 1'b0 ;
  assign n14783 = n9340 ^ n7265 ^ 1'b0 ;
  assign n14784 = n2790 | n14783 ;
  assign n14785 = n14784 ^ n318 ^ 1'b0 ;
  assign n14786 = n14785 ^ n522 ^ 1'b0 ;
  assign n14787 = n763 & n2538 ;
  assign n14788 = n14787 ^ n1049 ^ 1'b0 ;
  assign n14789 = n2883 & n5144 ;
  assign n14790 = ~n378 & n5620 ;
  assign n14791 = n1774 & ~n14790 ;
  assign n14792 = ~n4965 & n14791 ;
  assign n14793 = n14792 ^ n9010 ^ 1'b0 ;
  assign n14795 = n330 | n439 ;
  assign n14796 = n48 & ~n14795 ;
  assign n14797 = n8714 & ~n14796 ;
  assign n14794 = n7435 | n7882 ;
  assign n14798 = n14797 ^ n14794 ^ 1'b0 ;
  assign n14799 = n4075 & ~n12395 ;
  assign n14800 = n14799 ^ n1205 ^ 1'b0 ;
  assign n14801 = n2263 ^ n46 ^ 1'b0 ;
  assign n14802 = n1817 | n14801 ;
  assign n14803 = n14802 ^ n13446 ^ 1'b0 ;
  assign n14804 = n7383 & n13610 ;
  assign n14805 = n5378 | n10293 ;
  assign n14809 = n11881 ^ n1864 ^ 1'b0 ;
  assign n14806 = n23 | n3957 ;
  assign n14807 = ( ~n6436 & n6763 ) | ( ~n6436 & n14806 ) | ( n6763 & n14806 ) ;
  assign n14808 = n14807 ^ n2565 ^ 1'b0 ;
  assign n14810 = n14809 ^ n14808 ^ 1'b0 ;
  assign n14811 = n14805 & n14810 ;
  assign n14812 = n2136 & n8972 ;
  assign n14813 = n3139 | n4597 ;
  assign n14814 = ~n924 & n3574 ;
  assign n14815 = n14814 ^ n506 ^ 1'b0 ;
  assign n14816 = n7051 ^ n1178 ^ 1'b0 ;
  assign n14817 = n14815 & ~n14816 ;
  assign n14818 = n4060 ^ n3226 ^ 1'b0 ;
  assign n14819 = n3423 | n14818 ;
  assign n14820 = n13384 ^ n497 ^ 1'b0 ;
  assign n14821 = n352 | n14820 ;
  assign n14822 = n14819 | n14821 ;
  assign n14823 = n2270 ^ n1693 ^ 1'b0 ;
  assign n14824 = n1736 & n14823 ;
  assign n14825 = n10926 & n14824 ;
  assign n14826 = n3297 & ~n3968 ;
  assign n14827 = n14721 ^ n5221 ^ 1'b0 ;
  assign n14828 = ~n7227 & n14827 ;
  assign n14829 = n2420 | n6876 ;
  assign n14830 = n14829 ^ n7051 ^ 1'b0 ;
  assign n14831 = n4949 & ~n14830 ;
  assign n14832 = n14831 ^ n14131 ^ 1'b0 ;
  assign n14833 = n10905 ^ n37 ^ 1'b0 ;
  assign n14834 = n1280 & n14833 ;
  assign n14835 = ~n315 & n5297 ;
  assign n14836 = n14835 ^ n3570 ^ 1'b0 ;
  assign n14838 = n3221 ^ n3099 ^ 1'b0 ;
  assign n14837 = n3030 | n6117 ;
  assign n14839 = n14838 ^ n14837 ^ 1'b0 ;
  assign n14840 = ~n2436 & n8614 ;
  assign n14841 = ~n847 & n926 ;
  assign n14842 = n7433 & n14686 ;
  assign n14843 = n859 & n14842 ;
  assign n14844 = n14841 & n14843 ;
  assign n14845 = n5522 & n5704 ;
  assign n14848 = n2209 & ~n5071 ;
  assign n14846 = ~n594 & n3620 ;
  assign n14847 = n4551 & n14846 ;
  assign n14849 = n14848 ^ n14847 ^ 1'b0 ;
  assign n14850 = ~n713 & n14849 ;
  assign n14851 = n1255 & n10841 ;
  assign n14852 = n14851 ^ n2278 ^ 1'b0 ;
  assign n14853 = ~n102 & n3665 ;
  assign n14854 = n14853 ^ n6633 ^ 1'b0 ;
  assign n14857 = n239 | n2212 ;
  assign n14858 = n239 & ~n14857 ;
  assign n14855 = n5761 & n6916 ;
  assign n14856 = ~n5761 & n14855 ;
  assign n14859 = n14858 ^ n14856 ^ 1'b0 ;
  assign n14860 = n14854 & n14859 ;
  assign n14861 = n68 | n1673 ;
  assign n14862 = n9164 & n14861 ;
  assign n14863 = n7894 ^ n1314 ^ 1'b0 ;
  assign n14864 = n11586 & ~n14863 ;
  assign n14865 = n14864 ^ n3516 ^ 1'b0 ;
  assign n14866 = n6331 & ~n14865 ;
  assign n14867 = n12688 & n14866 ;
  assign n14868 = n1435 & n13816 ;
  assign n14869 = n14868 ^ n6743 ^ 1'b0 ;
  assign n14870 = ~n5891 & n8873 ;
  assign n14871 = n14870 ^ n2865 ^ 1'b0 ;
  assign n14872 = n5982 | n14871 ;
  assign n14873 = n13837 ^ n2704 ^ 1'b0 ;
  assign n14874 = n14872 | n14873 ;
  assign n14875 = n14869 & ~n14874 ;
  assign n14876 = ~n6822 & n14875 ;
  assign n14877 = n678 & ~n2885 ;
  assign n14878 = n10097 ^ n6887 ^ 1'b0 ;
  assign n14879 = ~n14877 & n14878 ;
  assign n14880 = ~n1637 & n14879 ;
  assign n14881 = ~n1100 & n14880 ;
  assign n14882 = n1268 & n11539 ;
  assign n14884 = n7221 ^ n5884 ^ 1'b0 ;
  assign n14883 = n4174 | n8500 ;
  assign n14885 = n14884 ^ n14883 ^ 1'b0 ;
  assign n14887 = ~n4371 & n5323 ;
  assign n14886 = ( ~n119 & n3821 ) | ( ~n119 & n4322 ) | ( n3821 & n4322 ) ;
  assign n14888 = n14887 ^ n14886 ^ 1'b0 ;
  assign n14889 = n14885 & ~n14888 ;
  assign n14890 = n14889 ^ n4969 ^ 1'b0 ;
  assign n14891 = n9748 & n14890 ;
  assign n14892 = n328 & n1573 ;
  assign n14893 = ~n2064 & n3466 ;
  assign n14894 = n3181 | n14893 ;
  assign n14895 = n14892 | n14894 ;
  assign n14896 = n14895 ^ n84 ^ 1'b0 ;
  assign n14897 = n10223 | n10403 ;
  assign n14898 = n9887 & ~n13768 ;
  assign n14899 = ~n512 & n14898 ;
  assign n14900 = n2062 & ~n2727 ;
  assign n14901 = n14900 ^ n2817 ^ 1'b0 ;
  assign n14902 = n10812 & n13185 ;
  assign n14903 = ~n233 & n7751 ;
  assign n14904 = n14903 ^ n6275 ^ 1'b0 ;
  assign n14905 = ( n10431 & n14902 ) | ( n10431 & n14904 ) | ( n14902 & n14904 ) ;
  assign n14906 = n2917 & ~n14462 ;
  assign n14907 = n2367 | n5833 ;
  assign n14908 = ~n3522 & n10861 ;
  assign n14909 = n5884 ^ n3564 ^ 1'b0 ;
  assign n14910 = n351 | n14909 ;
  assign n14911 = n2618 & ~n14910 ;
  assign n14912 = ~n11645 & n14911 ;
  assign n14913 = n6401 & ~n14912 ;
  assign n14914 = n14908 & n14913 ;
  assign n14915 = n5065 | n6689 ;
  assign n14919 = n4247 ^ n2667 ^ 1'b0 ;
  assign n14920 = ~n6633 & n14919 ;
  assign n14921 = ~n4131 & n4340 ;
  assign n14922 = ~n14920 & n14921 ;
  assign n14916 = n2983 ^ n1900 ^ 1'b0 ;
  assign n14917 = n862 & n14916 ;
  assign n14918 = n14917 ^ n338 ^ 1'b0 ;
  assign n14923 = n14922 ^ n14918 ^ 1'b0 ;
  assign n14924 = n14915 | n14923 ;
  assign n14925 = n6846 ^ n5152 ^ 1'b0 ;
  assign n14926 = ~n622 & n14925 ;
  assign n14927 = n14926 ^ n8278 ^ 1'b0 ;
  assign n14928 = n10598 | n14927 ;
  assign n14929 = n14928 ^ n8056 ^ 1'b0 ;
  assign n14930 = n7497 & ~n7796 ;
  assign n14931 = n8552 ^ n408 ^ 1'b0 ;
  assign n14932 = ~n4850 & n14931 ;
  assign n14933 = n555 & n14932 ;
  assign n14934 = ~n6385 & n14933 ;
  assign n14935 = n14080 & n14934 ;
  assign n14936 = n1691 & ~n5505 ;
  assign n14937 = n14935 & ~n14936 ;
  assign n14940 = n3456 ^ n271 ^ 1'b0 ;
  assign n14941 = n281 & n14940 ;
  assign n14938 = ~n10014 & n14863 ;
  assign n14939 = n1078 | n14938 ;
  assign n14942 = n14941 ^ n14939 ^ 1'b0 ;
  assign n14943 = n412 | n7442 ;
  assign n14944 = ~n6387 & n13171 ;
  assign n14945 = ~n4564 & n6953 ;
  assign n14946 = ~n4548 & n10733 ;
  assign n14947 = n14946 ^ n5434 ^ 1'b0 ;
  assign n14948 = n5248 | n12680 ;
  assign n14949 = n1267 ^ n1117 ^ 1'b0 ;
  assign n14950 = ~n10117 & n14949 ;
  assign n14951 = n14950 ^ n6629 ^ 1'b0 ;
  assign n14953 = n888 ^ n492 ^ 1'b0 ;
  assign n14954 = n14953 ^ n4671 ^ n475 ;
  assign n14952 = ~n7479 & n12313 ;
  assign n14955 = n14954 ^ n14952 ^ 1'b0 ;
  assign n14956 = n14955 ^ n10865 ^ 1'b0 ;
  assign n14957 = n10459 & ~n14956 ;
  assign n14958 = n246 & n5686 ;
  assign n14959 = n1982 ^ n1467 ^ 1'b0 ;
  assign n14960 = n863 & n14959 ;
  assign n14961 = n922 & n14960 ;
  assign n14962 = n717 & n14961 ;
  assign n14963 = n14958 & n14962 ;
  assign n14964 = ~n2556 & n10512 ;
  assign n14965 = n8523 & n14964 ;
  assign n14966 = n5541 & n14965 ;
  assign n14967 = n1974 & n7920 ;
  assign n14968 = n128 & ~n4677 ;
  assign n14969 = ~n5681 & n14968 ;
  assign n14970 = n14969 ^ n3176 ^ 1'b0 ;
  assign n14971 = n5259 & n14970 ;
  assign n14972 = ~n1061 & n2204 ;
  assign n14973 = n292 & n14972 ;
  assign n14974 = n1597 | n14973 ;
  assign n14975 = n14974 ^ n12095 ^ 1'b0 ;
  assign n14976 = n14975 ^ n3483 ^ 1'b0 ;
  assign n14977 = n5258 ^ n2893 ^ 1'b0 ;
  assign n14978 = ~n3649 & n14977 ;
  assign n14979 = ~n3993 & n9287 ;
  assign n14980 = n14979 ^ n16 ^ 1'b0 ;
  assign n14981 = n4041 ^ n3976 ^ 1'b0 ;
  assign n14982 = n10055 & n14981 ;
  assign n14983 = ~n1742 & n4577 ;
  assign n14984 = n2979 | n6894 ;
  assign n14985 = ~n4700 & n14984 ;
  assign n14986 = n14985 ^ n2441 ^ 1'b0 ;
  assign n14987 = n2710 & n3684 ;
  assign n14988 = ~n1069 & n8508 ;
  assign n14989 = n1627 & n3552 ;
  assign n14990 = n14989 ^ n12185 ^ 1'b0 ;
  assign n14991 = x0 | n68 ;
  assign n14992 = n14991 ^ n14458 ^ 1'b0 ;
  assign n14993 = n4409 ^ n3651 ^ 1'b0 ;
  assign n14994 = n1929 & ~n14993 ;
  assign n14995 = ~n6981 & n14994 ;
  assign n14996 = n357 & n14995 ;
  assign n14997 = ~n1804 & n14996 ;
  assign n14998 = n139 & n14997 ;
  assign n14999 = n1913 | n10303 ;
  assign n15000 = n1802 | n14999 ;
  assign n15001 = n1966 & ~n2771 ;
  assign n15002 = ~n15000 & n15001 ;
  assign n15003 = n6245 & ~n9754 ;
  assign n15004 = n15003 ^ n726 ^ 1'b0 ;
  assign n15005 = n8517 ^ n371 ^ 1'b0 ;
  assign n15006 = n3851 ^ n380 ^ 1'b0 ;
  assign n15007 = n4764 & n15006 ;
  assign n15008 = ~n6685 & n15007 ;
  assign n15009 = ~n2984 & n15008 ;
  assign n15010 = n6922 & ~n15009 ;
  assign n15011 = n2443 | n14712 ;
  assign n15012 = n2598 | n15011 ;
  assign n15013 = ~n769 & n12539 ;
  assign n15014 = n2840 & n3897 ;
  assign n15015 = n5673 ^ n627 ^ 1'b0 ;
  assign n15016 = n15015 ^ n116 ^ 1'b0 ;
  assign n15017 = n6965 ^ n6453 ^ 1'b0 ;
  assign n15018 = ~n12299 & n15017 ;
  assign n15019 = n11997 ^ n5763 ^ 1'b0 ;
  assign n15020 = n15018 & ~n15019 ;
  assign n15021 = n685 | n11460 ;
  assign n15022 = n613 & n3857 ;
  assign n15023 = n8402 & n15022 ;
  assign n15024 = n10785 | n15023 ;
  assign n15025 = n4567 | n15024 ;
  assign n15026 = n2316 | n5021 ;
  assign n15027 = n3477 & ~n9654 ;
  assign n15028 = n15027 ^ n2031 ^ 1'b0 ;
  assign n15029 = n369 & ~n15028 ;
  assign n15030 = n1831 & n5452 ;
  assign n15031 = n13444 ^ n982 ^ 1'b0 ;
  assign n15032 = n15030 & ~n15031 ;
  assign n15033 = n8630 ^ n6102 ^ 1'b0 ;
  assign n15034 = ~n1167 & n13258 ;
  assign n15035 = n1760 | n2025 ;
  assign n15036 = ~n8969 & n15035 ;
  assign n15037 = ~n3801 & n15036 ;
  assign n15038 = n5161 & ~n15037 ;
  assign n15039 = n15038 ^ n4274 ^ 1'b0 ;
  assign n15040 = n15034 | n15039 ;
  assign n15041 = n2789 ^ n1048 ^ 1'b0 ;
  assign n15042 = n5041 | n5067 ;
  assign n15043 = n15041 | n15042 ;
  assign n15044 = n212 | n14690 ;
  assign n15045 = n4074 | n15044 ;
  assign n15046 = x2 | n692 ;
  assign n15047 = n960 | n15046 ;
  assign n15048 = n15047 ^ n5128 ^ 1'b0 ;
  assign n15053 = n9554 ^ n7794 ^ 1'b0 ;
  assign n15054 = n11827 | n15053 ;
  assign n15049 = n7187 ^ n6655 ^ 1'b0 ;
  assign n15050 = n2303 & n15049 ;
  assign n15051 = n3770 | n15050 ;
  assign n15052 = n15051 ^ n7710 ^ 1'b0 ;
  assign n15055 = n15054 ^ n15052 ^ 1'b0 ;
  assign n15056 = ~n3690 & n15055 ;
  assign n15057 = n7995 & ~n8685 ;
  assign n15058 = ~n1258 & n13915 ;
  assign n15059 = ~n58 & n6665 ;
  assign n15060 = n15059 ^ n9895 ^ 1'b0 ;
  assign n15061 = n13189 & ~n15060 ;
  assign n15062 = n15061 ^ n2618 ^ 1'b0 ;
  assign n15063 = n2308 & n8351 ;
  assign n15065 = ~n7194 & n12804 ;
  assign n15066 = n340 | n15065 ;
  assign n15064 = n10137 ^ n2246 ^ 1'b0 ;
  assign n15067 = n15066 ^ n15064 ^ 1'b0 ;
  assign n15068 = n14351 ^ n1601 ^ 1'b0 ;
  assign n15069 = n6880 ^ n928 ^ 1'b0 ;
  assign n15070 = n15069 ^ n1220 ^ 1'b0 ;
  assign n15071 = n532 | n15070 ;
  assign n15072 = ~n2148 & n7528 ;
  assign n15073 = n8885 ^ n4412 ^ 1'b0 ;
  assign n15074 = n15072 & ~n15073 ;
  assign n15075 = n15074 ^ n1704 ^ 1'b0 ;
  assign n15076 = n4965 | n9599 ;
  assign n15077 = n4347 & ~n15076 ;
  assign n15078 = n1822 & n11340 ;
  assign n15080 = ~n146 & n7439 ;
  assign n15081 = n5897 & ~n15080 ;
  assign n15079 = n3943 & n10544 ;
  assign n15082 = n15081 ^ n15079 ^ 1'b0 ;
  assign n15083 = n5739 ^ n1087 ^ 1'b0 ;
  assign n15084 = ~n9255 & n15083 ;
  assign n15085 = ~n1445 & n15084 ;
  assign n15086 = ~n15082 & n15085 ;
  assign n15090 = n102 & ~n310 ;
  assign n15091 = n15090 ^ n5889 ^ 1'b0 ;
  assign n15087 = n1936 | n2273 ;
  assign n15088 = n15087 ^ n8283 ^ 1'b0 ;
  assign n15089 = n6906 | n15088 ;
  assign n15092 = n15091 ^ n15089 ^ 1'b0 ;
  assign n15093 = n15092 ^ n4586 ^ n4121 ;
  assign n15094 = n290 & n11809 ;
  assign n15095 = n8271 & n15094 ;
  assign n15096 = n274 & ~n13599 ;
  assign n15097 = n3511 ^ n719 ^ 1'b0 ;
  assign n15098 = n1695 & ~n2068 ;
  assign n15099 = ~n10077 & n15098 ;
  assign n15100 = ~n12445 & n15099 ;
  assign n15101 = n4772 | n15100 ;
  assign n15102 = n9208 ^ n2856 ^ 1'b0 ;
  assign n15103 = n2506 & ~n15102 ;
  assign n15104 = n10784 & n15103 ;
  assign n15105 = ~n6438 & n15104 ;
  assign n15106 = n192 & ~n441 ;
  assign n15107 = n15106 ^ n520 ^ 1'b0 ;
  assign n15108 = ~n11606 & n15107 ;
  assign n15109 = n1523 | n14822 ;
  assign n15110 = n1010 & n2408 ;
  assign n15111 = n15110 ^ n5973 ^ 1'b0 ;
  assign n15112 = n310 | n5516 ;
  assign n15113 = ~n6886 & n15112 ;
  assign n15114 = ~n15111 & n15113 ;
  assign n15115 = n6152 & ~n12488 ;
  assign n15116 = n7116 ^ n5543 ^ 1'b0 ;
  assign n15117 = ( n1246 & ~n6433 ) | ( n1246 & n7771 ) | ( ~n6433 & n7771 ) ;
  assign n15118 = n13931 ^ n9461 ^ 1'b0 ;
  assign n15119 = ( ~n1020 & n15117 ) | ( ~n1020 & n15118 ) | ( n15117 & n15118 ) ;
  assign n15120 = n3260 & n14007 ;
  assign n15121 = n12721 & n15120 ;
  assign n15122 = n4365 | n14520 ;
  assign n15123 = n2779 & n3037 ;
  assign n15124 = ~n2705 & n15123 ;
  assign n15125 = n11916 | n15124 ;
  assign n15126 = n15125 ^ n1516 ^ 1'b0 ;
  assign n15127 = n7732 & ~n8634 ;
  assign n15128 = n6761 & n15127 ;
  assign n15129 = n4439 | n6253 ;
  assign n15130 = n15129 ^ n4933 ^ 1'b0 ;
  assign n15131 = ~n8596 & n15130 ;
  assign n15132 = n15131 ^ n14213 ^ 1'b0 ;
  assign n15133 = n7326 | n11584 ;
  assign n15134 = n5792 & ~n15133 ;
  assign n15135 = n2418 & n9797 ;
  assign n15136 = n958 ^ n310 ^ 1'b0 ;
  assign n15137 = n15136 ^ n10208 ^ 1'b0 ;
  assign n15138 = n613 & ~n1086 ;
  assign n15139 = n5800 & n15138 ;
  assign n15140 = n5031 & n9267 ;
  assign n15141 = n15140 ^ n10390 ^ 1'b0 ;
  assign n15142 = n13794 | n15141 ;
  assign n15143 = n2450 & ~n15142 ;
  assign n15144 = n15143 ^ n6875 ^ 1'b0 ;
  assign n15145 = n6995 ^ n3074 ^ 1'b0 ;
  assign n15146 = n12432 & n15145 ;
  assign n15147 = n11795 ^ n4968 ^ 1'b0 ;
  assign n15148 = n9292 & n15147 ;
  assign n15149 = n5196 ^ n2097 ^ 1'b0 ;
  assign n15150 = n2116 | n15149 ;
  assign n15151 = ~n15148 & n15150 ;
  assign n15152 = n501 | n9574 ;
  assign n15153 = n8373 ^ n591 ^ 1'b0 ;
  assign n15154 = n294 & ~n15153 ;
  assign n15155 = n715 & n10448 ;
  assign n15156 = n15155 ^ n3311 ^ 1'b0 ;
  assign n15157 = n3065 ^ n1106 ^ 1'b0 ;
  assign n15158 = n12929 ^ n2040 ^ 1'b0 ;
  assign n15159 = n4327 & ~n15158 ;
  assign n15160 = ~n833 & n908 ;
  assign n15161 = ~n15159 & n15160 ;
  assign n15162 = x10 & n4751 ;
  assign n15163 = ~n5326 & n11715 ;
  assign n15165 = ~n4726 & n11521 ;
  assign n15164 = n9645 & n13817 ;
  assign n15166 = n15165 ^ n15164 ^ 1'b0 ;
  assign n15167 = n9698 ^ n308 ^ 1'b0 ;
  assign n15168 = n5013 & ~n15167 ;
  assign n15169 = n13015 ^ n1178 ^ 1'b0 ;
  assign n15170 = n2851 ^ n592 ^ 1'b0 ;
  assign n15171 = ~n9218 & n15170 ;
  assign n15172 = n14321 & n15171 ;
  assign n15173 = n1637 | n2144 ;
  assign n15174 = n2172 & ~n15173 ;
  assign n15175 = n15174 ^ n5424 ^ n5248 ;
  assign n15176 = ~n2020 & n5657 ;
  assign n15177 = n5218 | n15176 ;
  assign n15180 = ~n613 & n3037 ;
  assign n15178 = n10794 ^ n6681 ^ 1'b0 ;
  assign n15179 = n9053 & ~n15178 ;
  assign n15181 = n15180 ^ n15179 ^ 1'b0 ;
  assign n15182 = n495 & ~n11722 ;
  assign n15183 = n15182 ^ n832 ^ 1'b0 ;
  assign n15184 = n4356 & ~n15183 ;
  assign n15185 = n15184 ^ n7596 ^ 1'b0 ;
  assign n15186 = n12472 ^ n4076 ^ 1'b0 ;
  assign n15187 = n2388 & ~n15186 ;
  assign n15188 = n3559 | n15187 ;
  assign n15189 = n1710 | n15188 ;
  assign n15190 = ~n882 & n2130 ;
  assign n15191 = n615 & n15190 ;
  assign n15192 = ~n495 & n15131 ;
  assign n15193 = n684 & n5021 ;
  assign n15194 = ( ~n962 & n2580 ) | ( ~n962 & n5523 ) | ( n2580 & n5523 ) ;
  assign n15195 = n1414 & n2714 ;
  assign n15196 = n15195 ^ n12339 ^ 1'b0 ;
  assign n15198 = n685 & ~n690 ;
  assign n15197 = n5495 & ~n14605 ;
  assign n15199 = n15198 ^ n15197 ^ 1'b0 ;
  assign n15200 = n8226 ^ n4600 ^ 1'b0 ;
  assign n15201 = n3939 ^ n2879 ^ 1'b0 ;
  assign n15202 = n4537 ^ n594 ^ 1'b0 ;
  assign n15203 = ~n15201 & n15202 ;
  assign n15204 = n15200 & n15203 ;
  assign n15205 = n15204 ^ n6458 ^ 1'b0 ;
  assign n15206 = n7074 & ~n8874 ;
  assign n15207 = n15206 ^ n10771 ^ 1'b0 ;
  assign n15208 = n4426 & n9043 ;
  assign n15209 = ~n3805 & n5189 ;
  assign n15210 = n5067 & n15209 ;
  assign n15211 = n2347 & ~n15210 ;
  assign n15212 = n15211 ^ n14037 ^ 1'b0 ;
  assign n15213 = n10634 ^ n6575 ^ 1'b0 ;
  assign n15214 = n7118 | n15213 ;
  assign n15215 = n13591 ^ n5499 ^ 1'b0 ;
  assign n15216 = ~n2517 & n15215 ;
  assign n15217 = ~n8389 & n15216 ;
  assign n15218 = n15217 ^ n7850 ^ 1'b0 ;
  assign n15219 = ~n2568 & n6852 ;
  assign n15220 = ~n8723 & n15219 ;
  assign n15221 = n773 & n15220 ;
  assign n15222 = n15045 | n15221 ;
  assign n15223 = n8994 | n14975 ;
  assign n15224 = n2853 & ~n10255 ;
  assign n15225 = n596 | n3988 ;
  assign n15226 = n15225 ^ n9811 ^ 1'b0 ;
  assign n15227 = n15226 ^ n9526 ^ 1'b0 ;
  assign n15228 = ~n3629 & n9504 ;
  assign n15229 = n15227 & n15228 ;
  assign n15230 = ~n4330 & n9059 ;
  assign n15231 = n15230 ^ n5297 ^ 1'b0 ;
  assign n15232 = n5956 | n10707 ;
  assign n15233 = n4453 ^ n454 ^ 1'b0 ;
  assign n15234 = n7420 ^ n4212 ^ 1'b0 ;
  assign n15235 = n1205 | n15234 ;
  assign n15236 = ~n1324 & n2377 ;
  assign n15237 = n15236 ^ n1474 ^ 1'b0 ;
  assign n15238 = ( n1668 & n15235 ) | ( n1668 & ~n15237 ) | ( n15235 & ~n15237 ) ;
  assign n15239 = n9611 & n15238 ;
  assign n15240 = ~n10508 & n15239 ;
  assign n15241 = n1565 & ~n5625 ;
  assign n15242 = n7516 & n10914 ;
  assign n15243 = n15242 ^ n6191 ^ 1'b0 ;
  assign n15244 = ~n857 & n15243 ;
  assign n15245 = n8513 | n12295 ;
  assign n15246 = n2460 | n8672 ;
  assign n15247 = n9244 ^ n321 ^ 1'b0 ;
  assign n15248 = n2289 & n15247 ;
  assign n15249 = n15248 ^ n6332 ^ 1'b0 ;
  assign n15250 = ( ~n476 & n512 ) | ( ~n476 & n547 ) | ( n512 & n547 ) ;
  assign n15251 = n9029 | n15250 ;
  assign n15252 = n1447 | n15251 ;
  assign n15253 = ~n2129 & n2562 ;
  assign n15254 = n7896 & ~n15253 ;
  assign n15255 = n15254 ^ n596 ^ 1'b0 ;
  assign n15256 = n15255 ^ n11859 ^ 1'b0 ;
  assign n15257 = n7928 | n13186 ;
  assign n15258 = n7323 & ~n15257 ;
  assign n15259 = n1432 ^ n817 ^ 1'b0 ;
  assign n15260 = n15259 ^ n1901 ^ 1'b0 ;
  assign n15261 = n12025 & ~n15260 ;
  assign n15262 = n4115 | n6927 ;
  assign n15263 = n1933 | n6704 ;
  assign n15264 = n6982 & n9124 ;
  assign n15265 = n1810 & ~n15264 ;
  assign n15266 = n8401 ^ n2352 ^ 1'b0 ;
  assign n15267 = n2361 & n6644 ;
  assign n15268 = n5080 & n11761 ;
  assign n15269 = ~n11355 & n15268 ;
  assign n15270 = n8549 | n15269 ;
  assign n15271 = n15267 | n15270 ;
  assign n15272 = n13710 & ~n13743 ;
  assign n15273 = n15272 ^ n13088 ^ 1'b0 ;
  assign n15274 = n7390 & ~n9805 ;
  assign n15275 = n4171 & ~n4241 ;
  assign n15276 = n15275 ^ n3674 ^ 1'b0 ;
  assign n15277 = n966 & n4961 ;
  assign n15278 = n372 & n15277 ;
  assign n15279 = n3617 ^ n963 ^ 1'b0 ;
  assign n15280 = ~n11096 & n15279 ;
  assign n15281 = n15280 ^ n11039 ^ 1'b0 ;
  assign n15282 = n1007 & ~n14525 ;
  assign n15283 = n4976 & n15282 ;
  assign n15284 = n2542 & n15283 ;
  assign n15285 = n294 | n6067 ;
  assign n15286 = n13829 ^ n2097 ^ 1'b0 ;
  assign n15287 = ~n385 & n15286 ;
  assign n15288 = n2142 ^ n1816 ^ 1'b0 ;
  assign n15289 = n7319 & n15288 ;
  assign n15290 = n11167 & n13338 ;
  assign n15291 = n15290 ^ n5914 ^ 1'b0 ;
  assign n15292 = ~n8139 & n9985 ;
  assign n15293 = n10786 ^ n1181 ^ 1'b0 ;
  assign n15294 = n15293 ^ n8054 ^ 1'b0 ;
  assign n15295 = ~n52 & n10734 ;
  assign n15296 = ~n6871 & n15295 ;
  assign n15297 = ~n8435 & n15296 ;
  assign n15298 = n15232 ^ n6444 ^ 1'b0 ;
  assign n15299 = n10551 ^ n2162 ^ 1'b0 ;
  assign n15300 = n13196 ^ n1031 ^ 1'b0 ;
  assign n15301 = n6587 ^ n4791 ^ 1'b0 ;
  assign n15302 = n7523 & n15301 ;
  assign n15303 = n3398 ^ n2930 ^ 1'b0 ;
  assign n15304 = n1774 & n15303 ;
  assign n15305 = n1243 & n7865 ;
  assign n15306 = n15305 ^ n7596 ^ 1'b0 ;
  assign n15307 = n695 | n15306 ;
  assign n15308 = ~n227 & n3089 ;
  assign n15309 = n1488 | n2933 ;
  assign n15310 = n2157 & ~n2979 ;
  assign n15311 = n1714 | n6709 ;
  assign n15312 = n4700 & ~n15311 ;
  assign n15315 = n549 & n14932 ;
  assign n15316 = n15315 ^ n2014 ^ 1'b0 ;
  assign n15314 = n5668 & ~n11180 ;
  assign n15317 = n15316 ^ n15314 ^ 1'b0 ;
  assign n15313 = n1772 ^ n1398 ^ 1'b0 ;
  assign n15318 = n15317 ^ n15313 ^ 1'b0 ;
  assign n15319 = n1263 & ~n8723 ;
  assign n15323 = ~n2478 & n11855 ;
  assign n15324 = ~n8414 & n15323 ;
  assign n15321 = ( n489 & ~n498 ) | ( n489 & n957 ) | ( ~n498 & n957 ) ;
  assign n15320 = n12162 | n12190 ;
  assign n15322 = n15321 ^ n15320 ^ 1'b0 ;
  assign n15325 = n15324 ^ n15322 ^ 1'b0 ;
  assign n15326 = ~n2288 & n8666 ;
  assign n15327 = n2261 & ~n7780 ;
  assign n15328 = n11242 & n15327 ;
  assign n15329 = n13806 ^ n8331 ^ 1'b0 ;
  assign n15330 = n6887 & ~n15154 ;
  assign n15331 = n13175 ^ n2462 ^ 1'b0 ;
  assign n15332 = n13954 & ~n15331 ;
  assign n15333 = n8662 & ~n11288 ;
  assign n15358 = n3187 & ~n14790 ;
  assign n15359 = n14790 & n15358 ;
  assign n15360 = n15359 ^ n5465 ^ 1'b0 ;
  assign n15334 = n2496 | n7420 ;
  assign n15335 = ~n14080 & n15334 ;
  assign n15336 = n15335 ^ n10035 ^ 1'b0 ;
  assign n15337 = ~n9966 & n15336 ;
  assign n15338 = n9966 & n15337 ;
  assign n15339 = n601 | n5739 ;
  assign n15340 = n601 & ~n15339 ;
  assign n15341 = ~n35 & n512 ;
  assign n15342 = ~n512 & n15341 ;
  assign n15343 = n15340 & n15342 ;
  assign n15344 = n1183 & n15343 ;
  assign n15345 = n744 | n15344 ;
  assign n15346 = n15344 & ~n15345 ;
  assign n15347 = n170 & ~n2582 ;
  assign n15348 = n6793 & n15347 ;
  assign n15349 = n423 & ~n15348 ;
  assign n15350 = ~n423 & n15349 ;
  assign n15351 = n15346 | n15350 ;
  assign n15352 = n15346 & ~n15351 ;
  assign n15353 = n8581 | n15352 ;
  assign n15354 = n8581 & ~n15353 ;
  assign n15355 = n7033 & ~n15354 ;
  assign n15356 = ~n7033 & n15355 ;
  assign n15357 = n15338 | n15356 ;
  assign n15361 = n15360 ^ n15357 ^ 1'b0 ;
  assign n15362 = n1143 & n12239 ;
  assign n15363 = n10439 & ~n14264 ;
  assign n15364 = n15363 ^ n10976 ^ 1'b0 ;
  assign n15365 = n12541 ^ n11382 ^ 1'b0 ;
  assign n15366 = n4000 | n15365 ;
  assign n15367 = n939 | n1293 ;
  assign n15368 = n15367 ^ n13111 ^ 1'b0 ;
  assign n15369 = ~n2914 & n3601 ;
  assign n15370 = n15369 ^ n2176 ^ 1'b0 ;
  assign n15371 = n15370 ^ n12373 ^ 1'b0 ;
  assign n15372 = ~n15368 & n15371 ;
  assign n15373 = x1 | n2771 ;
  assign n15374 = x1 & ~n15373 ;
  assign n15375 = n1227 | n15374 ;
  assign n15376 = n1227 & ~n15375 ;
  assign n15377 = ( n3049 & ~n3329 ) | ( n3049 & n3753 ) | ( ~n3329 & n3753 ) ;
  assign n15378 = n15376 & n15377 ;
  assign n15379 = ( n6265 & n13183 ) | ( n6265 & n15378 ) | ( n13183 & n15378 ) ;
  assign n15380 = n14961 ^ n10584 ^ n5716 ;
  assign n15381 = n1388 & ~n2648 ;
  assign n15382 = n5560 ^ n1412 ^ 1'b0 ;
  assign n15383 = n2780 & n15382 ;
  assign n15384 = ~n2947 & n15383 ;
  assign n15385 = ~n3653 & n15384 ;
  assign n15386 = n2112 & ~n4850 ;
  assign n15387 = n4850 & n15386 ;
  assign n15388 = n105 & ~n9949 ;
  assign n15389 = ~n105 & n15388 ;
  assign n15390 = n3783 ^ n1181 ^ 1'b0 ;
  assign n15391 = n15389 & ~n15390 ;
  assign n15392 = n15387 | n15391 ;
  assign n15393 = n10191 | n15392 ;
  assign n15394 = n15392 & ~n15393 ;
  assign n15395 = n705 ^ n321 ^ 1'b0 ;
  assign n15396 = n2307 | n15395 ;
  assign n15397 = n15396 ^ n1959 ^ 1'b0 ;
  assign n15398 = n15397 ^ n13208 ^ 1'b0 ;
  assign n15399 = ~n6050 & n9154 ;
  assign n15400 = n86 | n13895 ;
  assign n15401 = n15084 ^ n4114 ^ 1'b0 ;
  assign n15402 = ~n10995 & n15401 ;
  assign n15403 = n3103 & ~n15402 ;
  assign n15404 = n4700 & n11296 ;
  assign n15405 = ( ~n1061 & n3120 ) | ( ~n1061 & n3286 ) | ( n3120 & n3286 ) ;
  assign n15406 = n15405 ^ n2432 ^ 1'b0 ;
  assign n15407 = n11313 ^ n5733 ^ 1'b0 ;
  assign n15408 = n151 & ~n3003 ;
  assign n15409 = n13755 & n15408 ;
  assign n15410 = n1898 & ~n11941 ;
  assign n15411 = n15012 ^ n6973 ^ 1'b0 ;
  assign n15412 = ~n11574 & n12540 ;
  assign n15413 = n561 & n1157 ;
  assign n15414 = n7863 & n15413 ;
  assign n15415 = ~n3063 & n10644 ;
  assign n15416 = n11269 ^ n4898 ^ 1'b0 ;
  assign n15417 = n15416 ^ n3240 ^ 1'b0 ;
  assign n15418 = n3941 & ~n15417 ;
  assign n15419 = n149 | n11829 ;
  assign n15420 = n10874 ^ n10396 ^ 1'b0 ;
  assign n15421 = n9474 | n15420 ;
  assign n15422 = ~n951 & n15421 ;
  assign n15423 = n6315 ^ n3485 ^ 1'b0 ;
  assign n15424 = ~n15422 & n15423 ;
  assign n15425 = n3907 ^ n616 ^ 1'b0 ;
  assign n15426 = n2568 | n15425 ;
  assign n15427 = n5551 | n11973 ;
  assign n15428 = n12766 ^ n4532 ^ 1'b0 ;
  assign n15429 = n1695 & n15428 ;
  assign n15430 = n4256 & n15429 ;
  assign n15431 = n364 & n737 ;
  assign n15432 = n1917 & n3514 ;
  assign n15433 = ~n15431 & n15432 ;
  assign n15434 = n7381 | n12324 ;
  assign n15435 = n9890 & ~n14040 ;
  assign n15436 = n3459 | n10273 ;
  assign n15437 = n11272 | n15436 ;
  assign n15439 = n614 & ~n4483 ;
  assign n15438 = n10166 ^ n1588 ^ 1'b0 ;
  assign n15440 = n15439 ^ n15438 ^ 1'b0 ;
  assign n15441 = n1822 | n15440 ;
  assign n15442 = n700 & ~n9571 ;
  assign n15443 = n15442 ^ n5569 ^ 1'b0 ;
  assign n15444 = n15443 ^ n2291 ^ 1'b0 ;
  assign n15445 = n4439 ^ n1559 ^ 1'b0 ;
  assign n15446 = n15445 ^ n13206 ^ 1'b0 ;
  assign n15447 = n10031 & n15446 ;
  assign n15448 = ~n2925 & n15447 ;
  assign n15449 = n2591 | n3527 ;
  assign n15450 = n15449 ^ n7981 ^ 1'b0 ;
  assign n15451 = n15450 ^ n7427 ^ n1987 ;
  assign n15452 = n4202 & n4872 ;
  assign n15453 = n15452 ^ n1737 ^ 1'b0 ;
  assign n15454 = n7523 & ~n15453 ;
  assign n15455 = n10309 & ~n11764 ;
  assign n15456 = n14978 ^ n3335 ^ 1'b0 ;
  assign n15457 = n8760 ^ n2261 ^ 1'b0 ;
  assign n15458 = n15129 ^ n4279 ^ 1'b0 ;
  assign n15459 = n268 & n1833 ;
  assign n15460 = n6361 | n7374 ;
  assign n15461 = n6361 & ~n15460 ;
  assign n15462 = n5470 | n10624 ;
  assign n15463 = n15462 ^ n10793 ^ 1'b0 ;
  assign n15464 = n6558 ^ n1903 ^ 1'b0 ;
  assign n15465 = n9697 | n15464 ;
  assign n15466 = ~x3 & n5144 ;
  assign n15467 = n5942 & n15466 ;
  assign n15468 = ~n5978 & n11375 ;
  assign n15469 = n11777 ^ n2546 ^ 1'b0 ;
  assign n15470 = n323 | n2842 ;
  assign n15471 = n2311 & n3093 ;
  assign n15472 = n15471 ^ n482 ^ 1'b0 ;
  assign n15473 = n723 & ~n15472 ;
  assign n15474 = ~n3993 & n15473 ;
  assign n15475 = n15470 & n15474 ;
  assign n15476 = n15475 ^ n6440 ^ 1'b0 ;
  assign n15477 = n2953 & n8869 ;
  assign n15478 = n13898 & n15477 ;
  assign n15479 = n13844 ^ n10274 ^ 1'b0 ;
  assign n15480 = n70 | n1810 ;
  assign n15481 = n10756 ^ n8897 ^ 1'b0 ;
  assign n15482 = n9767 ^ n5016 ^ 1'b0 ;
  assign n15483 = n15482 ^ n3262 ^ 1'b0 ;
  assign n15484 = n7487 ^ n1426 ^ 1'b0 ;
  assign n15485 = n4511 ^ n1992 ^ 1'b0 ;
  assign n15486 = n624 & n15485 ;
  assign n15487 = n81 & n15486 ;
  assign n15488 = n15487 ^ n14323 ^ 1'b0 ;
  assign n15489 = n11025 & n13359 ;
  assign n15490 = n11295 & n15489 ;
  assign n15491 = n3523 | n8198 ;
  assign n15492 = n15491 ^ n5837 ^ 1'b0 ;
  assign n15493 = ~n9261 & n15492 ;
  assign n15494 = n7609 ^ n6420 ^ 1'b0 ;
  assign n15495 = n274 | n15494 ;
  assign n15496 = n11322 ^ n1110 ^ 1'b0 ;
  assign n15497 = n1929 & ~n15496 ;
  assign n15498 = n10992 ^ n619 ^ 1'b0 ;
  assign n15499 = n9992 & ~n15498 ;
  assign n15505 = n2256 ^ n791 ^ 1'b0 ;
  assign n15506 = n12504 | n15505 ;
  assign n15501 = ~n3263 & n5172 ;
  assign n15502 = n15501 ^ n2826 ^ 1'b0 ;
  assign n15500 = n475 & n3345 ;
  assign n15503 = n15502 ^ n15500 ^ 1'b0 ;
  assign n15504 = n1414 & n15503 ;
  assign n15507 = n15506 ^ n15504 ^ 1'b0 ;
  assign n15508 = n227 | n5299 ;
  assign n15509 = n594 & ~n15508 ;
  assign n15510 = n4322 | n4972 ;
  assign n15511 = n9001 & ~n15510 ;
  assign n15512 = n15509 & ~n15511 ;
  assign n15513 = n6763 ^ n619 ^ 1'b0 ;
  assign n15514 = ~n5887 & n15513 ;
  assign n15515 = n4054 | n7325 ;
  assign n15516 = n2367 & n15515 ;
  assign n15517 = n15066 ^ n2535 ^ 1'b0 ;
  assign n15518 = n15516 | n15517 ;
  assign n15519 = n4052 & n12678 ;
  assign n15520 = n3887 | n8690 ;
  assign n15521 = ~n1763 & n8409 ;
  assign n15522 = n852 | n3064 ;
  assign n15523 = n3152 & ~n15522 ;
  assign n15524 = ~n15521 & n15523 ;
  assign n15525 = n10383 | n15524 ;
  assign n15526 = ~n1473 & n5234 ;
  assign n15527 = n2351 & n5580 ;
  assign n15528 = n15527 ^ n36 ^ 1'b0 ;
  assign n15529 = n15526 | n15528 ;
  assign n15530 = n7978 ^ n1430 ^ 1'b0 ;
  assign n15531 = ~n12512 & n15530 ;
  assign n15532 = n14874 & n15531 ;
  assign n15533 = ~n5140 & n15532 ;
  assign n15534 = n4664 ^ n958 ^ 1'b0 ;
  assign n15535 = n13108 ^ n3864 ^ 1'b0 ;
  assign n15536 = n10228 | n15535 ;
  assign n15537 = n10327 & ~n15536 ;
  assign n15538 = ~n79 & n6667 ;
  assign n15539 = ~n8082 & n15538 ;
  assign n15540 = n15537 | n15539 ;
  assign n15541 = n15540 ^ n4039 ^ 1'b0 ;
  assign n15542 = n501 ^ n335 ^ 1'b0 ;
  assign n15543 = ~n1039 & n5059 ;
  assign n15544 = n2495 & ~n4606 ;
  assign n15545 = n2752 | n15544 ;
  assign n15546 = n15539 & ~n15545 ;
  assign n15547 = n509 & ~n3808 ;
  assign n15548 = n622 ^ n246 ^ 1'b0 ;
  assign n15549 = n10153 & n15548 ;
  assign n15550 = n5679 & n15549 ;
  assign n15551 = n8784 & n15550 ;
  assign n15552 = n15547 | n15551 ;
  assign n15553 = ~n6935 & n11417 ;
  assign n15554 = ~n1072 & n15553 ;
  assign n15555 = n15554 ^ n1924 ^ 1'b0 ;
  assign n15556 = n616 | n7609 ;
  assign n15557 = n4883 & ~n15556 ;
  assign n15558 = n616 & n11226 ;
  assign n15559 = n2377 | n15558 ;
  assign n15560 = n3464 & ~n7679 ;
  assign n15561 = n2733 & n4302 ;
  assign n15562 = n1688 | n4990 ;
  assign n15563 = n1688 & ~n15562 ;
  assign n15564 = n1174 & n4440 ;
  assign n15565 = ~n4440 & n15564 ;
  assign n15566 = n1707 | n15565 ;
  assign n15567 = n15563 | n15566 ;
  assign n15568 = n15561 & ~n15567 ;
  assign n15569 = ~n15561 & n15568 ;
  assign n15570 = n8057 ^ n6885 ^ 1'b0 ;
  assign n15571 = n15570 ^ x7 ^ 1'b0 ;
  assign n15572 = n15431 & n15571 ;
  assign n15573 = n200 | n10861 ;
  assign n15574 = n13853 | n15573 ;
  assign n15576 = n9819 ^ n254 ^ 1'b0 ;
  assign n15575 = n2613 & ~n10448 ;
  assign n15577 = n15576 ^ n15575 ^ n4832 ;
  assign n15578 = ~n6090 & n10862 ;
  assign n15579 = n4463 & n15578 ;
  assign n15580 = n3449 ^ n1874 ^ n1095 ;
  assign n15581 = n6245 & ~n7330 ;
  assign n15582 = ~n15580 & n15581 ;
  assign n15583 = ~n3227 & n15582 ;
  assign n15584 = n5208 & ~n6096 ;
  assign n15585 = n38 & n15584 ;
  assign n15586 = n10055 ^ n497 ^ 1'b0 ;
  assign n15587 = n3817 & ~n15586 ;
  assign n15588 = n15585 & n15587 ;
  assign n15589 = n1039 | n11447 ;
  assign n15590 = n12682 | n15589 ;
  assign n15591 = ~n4710 & n15590 ;
  assign n15592 = n8278 ^ n6665 ^ 1'b0 ;
  assign n15593 = n5551 & ~n15592 ;
  assign n15594 = ~n3464 & n15593 ;
  assign n15595 = ~n12249 & n15594 ;
  assign n15596 = n3701 ^ n94 ^ 1'b0 ;
  assign n15597 = n15596 ^ n8106 ^ 1'b0 ;
  assign n15598 = n3354 ^ n1426 ^ 1'b0 ;
  assign n15599 = ~n7943 & n15598 ;
  assign n15600 = n15599 ^ n488 ^ 1'b0 ;
  assign n15601 = ~n338 & n4191 ;
  assign n15602 = n9218 & n15601 ;
  assign n15603 = n3228 | n15602 ;
  assign n15604 = n15603 ^ n612 ^ 1'b0 ;
  assign n15605 = n1747 | n15604 ;
  assign n15606 = n2348 | n5891 ;
  assign n15607 = n2517 | n2753 ;
  assign n15608 = n302 | n460 ;
  assign n15609 = n15608 ^ n14493 ^ 1'b0 ;
  assign n15610 = n15609 ^ n11723 ^ 1'b0 ;
  assign n15611 = n15607 | n15610 ;
  assign n15612 = n4805 ^ n4031 ^ 1'b0 ;
  assign n15613 = n7545 & n15612 ;
  assign n15614 = n4913 & ~n15613 ;
  assign n15615 = n4936 | n7466 ;
  assign n15616 = ~n1162 & n8836 ;
  assign n15617 = n15616 ^ n6306 ^ 1'b0 ;
  assign n15618 = ~n8830 & n15617 ;
  assign n15619 = n798 ^ n273 ^ 1'b0 ;
  assign n15620 = n212 | n15619 ;
  assign n15621 = n15620 ^ n62 ^ 1'b0 ;
  assign n15622 = n15621 ^ n188 ^ 1'b0 ;
  assign n15623 = n7504 | n15622 ;
  assign n15624 = n12382 ^ n5122 ^ 1'b0 ;
  assign n15625 = n5802 & n14253 ;
  assign n15626 = n11937 ^ n9796 ^ n3196 ;
  assign n15627 = n4261 & ~n7981 ;
  assign n15628 = n671 & n749 ;
  assign n15629 = n929 & n15628 ;
  assign n15630 = n7399 & ~n15629 ;
  assign n15631 = n15630 ^ n9732 ^ 1'b0 ;
  assign n15632 = n4618 ^ n2647 ^ 1'b0 ;
  assign n15633 = n15632 ^ n1766 ^ 1'b0 ;
  assign n15634 = n5217 ^ n1552 ^ 1'b0 ;
  assign n15635 = ~n11626 & n15634 ;
  assign n15636 = n4607 | n15132 ;
  assign n15637 = n15636 ^ n7516 ^ 1'b0 ;
  assign n15638 = n7355 | n11197 ;
  assign n15639 = ~n3969 & n15638 ;
  assign n15640 = n484 | n5702 ;
  assign n15641 = n3858 & ~n15640 ;
  assign n15642 = n15641 ^ n3280 ^ 1'b0 ;
  assign n15643 = n542 & ~n15255 ;
  assign n15644 = n119 & ~n15643 ;
  assign n15645 = n10982 ^ n8910 ^ 1'b0 ;
  assign n15646 = n8461 & n15645 ;
  assign n15647 = n8584 ^ n5273 ^ 1'b0 ;
  assign n15648 = n15646 & n15647 ;
  assign n15649 = ~n833 & n8128 ;
  assign n15650 = ~n375 & n2059 ;
  assign n15651 = n15650 ^ n12709 ^ n5730 ;
  assign n15652 = n15651 ^ n6220 ^ 1'b0 ;
  assign n15653 = n15652 ^ n5813 ^ 1'b0 ;
  assign n15654 = n5232 & ~n15653 ;
  assign n15655 = ~n10180 & n15654 ;
  assign n15656 = n417 & n7535 ;
  assign n15657 = n1410 & n15656 ;
  assign n15658 = x2 | n6963 ;
  assign n15659 = n15658 ^ n9204 ^ 1'b0 ;
  assign n15660 = n3221 & ~n4269 ;
  assign n15661 = n15660 ^ n3253 ^ 1'b0 ;
  assign n15662 = n3738 | n15661 ;
  assign n15663 = n15662 ^ n4622 ^ 1'b0 ;
  assign n15664 = n2193 | n15663 ;
  assign n15665 = n6498 ^ n4241 ^ 1'b0 ;
  assign n15666 = n366 & n15665 ;
  assign n15667 = n15666 ^ n1821 ^ 1'b0 ;
  assign n15668 = n7608 ^ n4590 ^ 1'b0 ;
  assign n15669 = n15667 | n15668 ;
  assign n15670 = n15669 ^ n11195 ^ 1'b0 ;
  assign n15671 = n11998 ^ n690 ^ 1'b0 ;
  assign n15672 = ~n6449 & n13042 ;
  assign n15674 = n3859 ^ n1165 ^ 1'b0 ;
  assign n15673 = n2945 & n6085 ;
  assign n15675 = n15674 ^ n15673 ^ 1'b0 ;
  assign n15676 = n2289 & n10855 ;
  assign n15677 = n3100 | n5643 ;
  assign n15678 = n8977 & ~n11611 ;
  assign n15679 = n9952 & n15390 ;
  assign n15680 = n15679 ^ n12325 ^ 1'b0 ;
  assign n15681 = n7848 & n8488 ;
  assign n15682 = n15681 ^ n6473 ^ 1'b0 ;
  assign n15683 = n9388 & n10991 ;
  assign n15684 = n2122 | n14457 ;
  assign n15685 = n9760 ^ n7322 ^ 1'b0 ;
  assign n15686 = ~n970 & n15685 ;
  assign n15687 = n6782 & ~n10194 ;
  assign n15688 = n10685 & n15687 ;
  assign n15689 = ~n2269 & n4549 ;
  assign n15690 = ~n963 & n1887 ;
  assign n15691 = n3643 & ~n15232 ;
  assign n15692 = n5559 & ~n6963 ;
  assign n15693 = n3431 | n5354 ;
  assign n15694 = ~n15692 & n15693 ;
  assign n15695 = n2127 | n4591 ;
  assign n15696 = n15695 ^ n968 ^ 1'b0 ;
  assign n15697 = ~n4600 & n5443 ;
  assign n15698 = n7856 ^ n7707 ^ 1'b0 ;
  assign n15699 = n1109 | n15698 ;
  assign n15700 = ~n5041 & n15699 ;
  assign n15701 = n14953 | n15700 ;
  assign n15702 = n2307 & ~n5568 ;
  assign n15703 = n15702 ^ n6070 ^ 1'b0 ;
  assign n15704 = ~n5128 & n15703 ;
  assign n15705 = n15704 ^ n15180 ^ 1'b0 ;
  assign n15706 = n10650 ^ n7497 ^ n1444 ;
  assign n15707 = n2328 & n13901 ;
  assign n15708 = n8295 ^ n3300 ^ 1'b0 ;
  assign n15709 = n2804 & n15708 ;
  assign n15710 = n524 & ~n4033 ;
  assign n15711 = ~n9504 & n15710 ;
  assign n15712 = n15711 ^ n7511 ^ 1'b0 ;
  assign n15713 = n10584 ^ n1856 ^ 1'b0 ;
  assign n15714 = ~n8189 & n8251 ;
  assign n15715 = n5060 & n6617 ;
  assign n15716 = n10976 ^ n3040 ^ 1'b0 ;
  assign n15717 = n3666 & ~n15716 ;
  assign n15718 = n1674 & n15717 ;
  assign n15719 = ~n472 & n15718 ;
  assign n15720 = n9417 & n15719 ;
  assign n15721 = ~n9318 & n9338 ;
  assign n15722 = n15013 ^ n5412 ^ 1'b0 ;
  assign n15723 = n3127 | n15722 ;
  assign n15724 = n8750 | n15516 ;
  assign n15726 = ~n64 & n7831 ;
  assign n15727 = n64 & n15726 ;
  assign n15728 = n153 & n581 ;
  assign n15729 = n15727 & n15728 ;
  assign n15730 = n749 & n15729 ;
  assign n15731 = n15730 ^ n354 ^ 1'b0 ;
  assign n15732 = n5475 | n13506 ;
  assign n15733 = n5475 & ~n15732 ;
  assign n15734 = n3059 & ~n15733 ;
  assign n15735 = ~n3059 & n15734 ;
  assign n15736 = n15731 & n15735 ;
  assign n15725 = n3849 | n5239 ;
  assign n15737 = n15736 ^ n15725 ^ 1'b0 ;
  assign n15744 = n995 | n2136 ;
  assign n15745 = n10181 | n15744 ;
  assign n15738 = n459 | n2978 ;
  assign n15739 = n12836 & ~n15738 ;
  assign n15740 = n5606 | n15739 ;
  assign n15741 = n5845 ^ n1043 ^ 1'b0 ;
  assign n15742 = n1891 & ~n15741 ;
  assign n15743 = ~n15740 & n15742 ;
  assign n15746 = n15745 ^ n15743 ^ 1'b0 ;
  assign n15747 = ( n3648 & n15737 ) | ( n3648 & n15746 ) | ( n15737 & n15746 ) ;
  assign n15748 = ~n694 & n1903 ;
  assign n15749 = n3321 & n15748 ;
  assign n15750 = n1699 & n7590 ;
  assign n15758 = n2538 ^ n737 ^ 1'b0 ;
  assign n15759 = n6857 & n15758 ;
  assign n15751 = n5241 & n7655 ;
  assign n15752 = n10772 & n15751 ;
  assign n15753 = n7611 ^ n7458 ^ 1'b0 ;
  assign n15754 = n2360 & n15753 ;
  assign n15755 = n3725 & n15754 ;
  assign n15756 = n15752 & n15755 ;
  assign n15757 = n10066 | n15756 ;
  assign n15760 = n15759 ^ n15757 ^ 1'b0 ;
  assign n15761 = n2977 ^ n622 ^ 1'b0 ;
  assign n15762 = n68 | n3264 ;
  assign n15763 = n15316 | n15762 ;
  assign n15764 = n1325 & n15763 ;
  assign n15765 = n10076 & n15764 ;
  assign n15766 = n15765 ^ n8318 ^ 1'b0 ;
  assign n15767 = ~n3037 & n4700 ;
  assign n15768 = n15767 ^ n1883 ^ 1'b0 ;
  assign n15769 = n958 & ~n11403 ;
  assign n15770 = n3311 | n7251 ;
  assign n15771 = n15770 ^ n1827 ^ 1'b0 ;
  assign n15772 = n15771 ^ n5696 ^ 1'b0 ;
  assign n15773 = n15769 & n15772 ;
  assign n15777 = n1263 & n1350 ;
  assign n15778 = n5313 | n15777 ;
  assign n15774 = n901 | n3967 ;
  assign n15775 = n15774 ^ n11745 ^ 1'b0 ;
  assign n15776 = n5344 & ~n15775 ;
  assign n15779 = n15778 ^ n15776 ^ 1'b0 ;
  assign n15780 = n13719 & ~n15779 ;
  assign n15781 = n15780 ^ n196 ^ 1'b0 ;
  assign n15782 = n3186 ^ n310 ^ 1'b0 ;
  assign n15783 = ~n66 & n1887 ;
  assign n15784 = n684 & n15783 ;
  assign n15785 = n7272 | n10534 ;
  assign n15786 = ~n2915 & n15785 ;
  assign n15787 = n503 & ~n1928 ;
  assign n15788 = n11842 ^ n4473 ^ 1'b0 ;
  assign n15789 = n6238 ^ n4976 ^ 1'b0 ;
  assign n15790 = ~n15788 & n15789 ;
  assign n15791 = n254 & n1304 ;
  assign n15792 = n1460 & ~n3640 ;
  assign n15793 = n15792 ^ n3130 ^ 1'b0 ;
  assign n15794 = n15791 | n15793 ;
  assign n15795 = n15794 ^ n12788 ^ 1'b0 ;
  assign n15796 = n15790 & ~n15795 ;
  assign n15797 = n15787 & n15796 ;
  assign n15798 = n11827 ^ n3053 ^ 1'b0 ;
  assign n15799 = ~n4816 & n15798 ;
  assign n15800 = n2526 & n10968 ;
  assign n15801 = n15800 ^ n9688 ^ 1'b0 ;
  assign n15802 = n2124 ^ n741 ^ 1'b0 ;
  assign n15803 = n10180 ^ n6434 ^ 1'b0 ;
  assign n15804 = n13419 | n15803 ;
  assign n15806 = n9056 ^ n4314 ^ 1'b0 ;
  assign n15807 = n15806 ^ n7047 ^ 1'b0 ;
  assign n15808 = ~n3633 & n15807 ;
  assign n15809 = ~n3346 & n6914 ;
  assign n15810 = ~n15808 & n15809 ;
  assign n15805 = n6819 & n8112 ;
  assign n15811 = n15810 ^ n15805 ^ 1'b0 ;
  assign n15812 = n7580 ^ n6644 ^ 1'b0 ;
  assign n15813 = n1668 & ~n14246 ;
  assign n15814 = n15813 ^ n615 ^ 1'b0 ;
  assign n15815 = n11263 & n15814 ;
  assign n15816 = ~n512 & n15815 ;
  assign n15817 = n14863 ^ n1674 ^ 1'b0 ;
  assign n15818 = n8470 | n15817 ;
  assign n15819 = n270 & n2866 ;
  assign n15820 = ~n11323 & n15819 ;
  assign n15821 = n10359 & ~n12877 ;
  assign n15822 = n15820 & ~n15821 ;
  assign n15823 = n2762 ^ n653 ^ 1'b0 ;
  assign n15826 = n627 & ~n1598 ;
  assign n15828 = n2693 ^ n274 ^ 1'b0 ;
  assign n15829 = n3075 & n15828 ;
  assign n15830 = n1469 ^ n688 ^ 1'b0 ;
  assign n15831 = n2584 & ~n15830 ;
  assign n15832 = n15829 & ~n15831 ;
  assign n15827 = n5967 & n9175 ;
  assign n15833 = n15832 ^ n15827 ^ 1'b0 ;
  assign n15834 = ( ~n6087 & n15826 ) | ( ~n6087 & n15833 ) | ( n15826 & n15833 ) ;
  assign n15824 = n636 & n832 ;
  assign n15825 = n15205 & ~n15824 ;
  assign n15835 = n15834 ^ n15825 ^ 1'b0 ;
  assign n15836 = n378 | n3631 ;
  assign n15837 = n15836 ^ n15316 ^ 1'b0 ;
  assign n15838 = n5256 | n15837 ;
  assign n15839 = n2458 | n3333 ;
  assign n15840 = n8404 | n15839 ;
  assign n15841 = n14712 ^ n6461 ^ 1'b0 ;
  assign n15842 = n14554 & n15841 ;
  assign n15843 = n5372 & n11963 ;
  assign n15844 = ~n844 & n15843 ;
  assign n15845 = n4809 ^ n4357 ^ 1'b0 ;
  assign n15846 = n9242 & ~n15845 ;
  assign n15847 = n15846 ^ n9554 ^ n9428 ;
  assign n15848 = ~n7609 & n11671 ;
  assign n15849 = ~n510 & n15848 ;
  assign n15850 = n30 & ~n15849 ;
  assign n15851 = n15850 ^ n8041 ^ 1'b0 ;
  assign n15854 = n348 & n6463 ;
  assign n15852 = n2142 & n5877 ;
  assign n15853 = n15852 ^ n133 ^ 1'b0 ;
  assign n15855 = n15854 ^ n15853 ^ 1'b0 ;
  assign n15856 = n7046 & ~n15855 ;
  assign n15857 = ~n4865 & n15856 ;
  assign n15858 = n1917 & ~n4004 ;
  assign n15859 = ~n6552 & n15858 ;
  assign n15860 = n12560 | n15859 ;
  assign n15861 = n2717 | n15860 ;
  assign n15862 = n15861 ^ n2397 ^ 1'b0 ;
  assign n15863 = ~n7386 & n13153 ;
  assign n15864 = n10995 ^ n3642 ^ 1'b0 ;
  assign n15865 = n1311 & n14068 ;
  assign n15866 = n3672 & n15865 ;
  assign n15867 = n15866 ^ n3595 ^ 1'b0 ;
  assign n15869 = n15576 ^ n5457 ^ 1'b0 ;
  assign n15868 = n1363 & ~n12817 ;
  assign n15870 = n15869 ^ n15868 ^ 1'b0 ;
  assign n15871 = n15870 ^ n8966 ^ 1'b0 ;
  assign n15872 = n9645 & ~n14202 ;
  assign n15873 = n1947 & n11036 ;
  assign n15874 = n15873 ^ n2545 ^ 1'b0 ;
  assign n15875 = ~n5338 & n15874 ;
  assign n15876 = n4746 | n6533 ;
  assign n15877 = ~n891 & n15876 ;
  assign n15878 = n15877 ^ n6339 ^ 1'b0 ;
  assign n15879 = ( n2187 & ~n2487 ) | ( n2187 & n4185 ) | ( ~n2487 & n4185 ) ;
  assign n15880 = n1988 & ~n15879 ;
  assign n15881 = ~n1988 & n15880 ;
  assign n15882 = n12284 | n15881 ;
  assign n15883 = n10687 ^ n6418 ^ 1'b0 ;
  assign n15884 = ~n3864 & n4840 ;
  assign n15885 = n3864 & n15884 ;
  assign n15886 = n2010 | n3613 ;
  assign n15887 = n15885 & ~n15886 ;
  assign n15888 = ~n15883 & n15887 ;
  assign n15889 = ~n9960 & n15888 ;
  assign n15890 = n15882 & n15889 ;
  assign n15891 = n4367 & ~n14712 ;
  assign n15892 = n15891 ^ n369 ^ 1'b0 ;
  assign n15893 = ~n3193 & n15892 ;
  assign n15894 = n8810 & n15893 ;
  assign n15895 = n3423 & n10083 ;
  assign n15896 = n2560 ^ n1714 ^ 1'b0 ;
  assign n15897 = n7683 & n15896 ;
  assign n15898 = n274 | n1170 ;
  assign n15899 = n2719 & ~n15898 ;
  assign n15900 = n4686 & n15899 ;
  assign n15901 = n15900 ^ n2907 ^ 1'b0 ;
  assign n15902 = n15901 ^ n101 ^ 1'b0 ;
  assign n15903 = n782 & ~n8946 ;
  assign n15904 = ( n489 & ~n2547 ) | ( n489 & n15903 ) | ( ~n2547 & n15903 ) ;
  assign n15905 = n2227 & n15259 ;
  assign n15906 = n4449 | n10644 ;
  assign n15907 = n809 & n9198 ;
  assign n15908 = n15906 & n15907 ;
  assign n15909 = n15908 ^ n7445 ^ 1'b0 ;
  assign n15912 = n1411 & n2221 ;
  assign n15910 = ~n1237 & n2917 ;
  assign n15911 = n158 | n15910 ;
  assign n15913 = n15912 ^ n15911 ^ n11269 ;
  assign n15914 = n13713 ^ n3014 ^ 1'b0 ;
  assign n15915 = n9668 | n15914 ;
  assign n15916 = n4221 & n6916 ;
  assign n15917 = n15916 ^ n1648 ^ 1'b0 ;
  assign n15918 = ~n15915 & n15917 ;
  assign n15919 = n128 | n729 ;
  assign n15920 = n3088 & ~n15919 ;
  assign n15921 = n553 & n6999 ;
  assign n15922 = n7377 ^ n2939 ^ 1'b0 ;
  assign n15923 = ~n15921 & n15922 ;
  assign n15924 = ~n3759 & n15923 ;
  assign n15925 = n5382 & n15924 ;
  assign n15926 = n13654 ^ n3424 ^ 1'b0 ;
  assign n15927 = n11413 ^ n8581 ^ 1'b0 ;
  assign n15928 = n1207 & n15927 ;
  assign n15929 = n14975 ^ n536 ^ 1'b0 ;
  assign n15930 = n15321 | n15929 ;
  assign n15931 = n2142 ^ n1715 ^ 1'b0 ;
  assign n15932 = ~n200 & n15931 ;
  assign n15933 = n15229 & n15862 ;
  assign n15934 = n17 & ~n1407 ;
  assign n15935 = ~n17 & n15934 ;
  assign n15938 = n34 & n387 ;
  assign n15939 = ~n387 & n15938 ;
  assign n15936 = n28 & ~n2469 ;
  assign n15937 = ~n28 & n15936 ;
  assign n15940 = n15939 ^ n15937 ^ 1'b0 ;
  assign n15941 = n15935 & n15940 ;
  assign n15942 = n8309 ^ n5364 ^ 1'b0 ;
  assign n15943 = n5714 & ~n15942 ;
  assign n15944 = n15941 & n15943 ;
  assign n15945 = ~n15941 & n15944 ;
  assign n15946 = ~n158 & n5404 ;
  assign n15947 = n158 & n15946 ;
  assign n15948 = n15945 & ~n15947 ;
  assign n15950 = n2448 & ~n12817 ;
  assign n15951 = ~n5286 & n15950 ;
  assign n15949 = ~n3674 & n10743 ;
  assign n15952 = n15951 ^ n15949 ^ 1'b0 ;
  assign n15953 = n4748 & n14776 ;
  assign n15954 = n15953 ^ n11123 ^ 1'b0 ;
  assign n15955 = n5894 & ~n12080 ;
  assign n15956 = ~n8697 & n15955 ;
  assign n15957 = n11040 & ~n15956 ;
  assign n15958 = ~n15954 & n15957 ;
  assign n15959 = n2028 & ~n8254 ;
  assign n15960 = n2785 & n4416 ;
  assign n15961 = n200 & ~n11840 ;
  assign n15962 = ~n4396 & n15961 ;
  assign n15963 = n15962 ^ n9629 ^ 1'b0 ;
  assign n15964 = n6080 ^ n1346 ^ 1'b0 ;
  assign n15965 = n5710 & ~n15964 ;
  assign n15966 = n6579 & ~n10544 ;
  assign n15968 = ~n880 & n5349 ;
  assign n15969 = ~n5349 & n15968 ;
  assign n15970 = ~n3030 & n4036 ;
  assign n15971 = n15969 & n15970 ;
  assign n15972 = n418 | n15971 ;
  assign n15973 = n418 & ~n15972 ;
  assign n15974 = ~n10475 & n15973 ;
  assign n15967 = n3586 | n13711 ;
  assign n15975 = n15974 ^ n15967 ^ 1'b0 ;
  assign n15976 = ~n9270 & n15975 ;
  assign n15977 = n15976 ^ n14879 ^ 1'b0 ;
  assign n15978 = n324 & ~n11742 ;
  assign n15979 = n387 & n1530 ;
  assign n15980 = n3068 ^ n2599 ^ 1'b0 ;
  assign n15981 = n6406 & ~n15980 ;
  assign n15982 = n5530 & ~n6479 ;
  assign n15983 = ~n15981 & n15982 ;
  assign n15984 = n15983 ^ n2165 ^ 1'b0 ;
  assign n15985 = ~n3901 & n15984 ;
  assign n15986 = n1874 & n3476 ;
  assign n15987 = n15986 ^ n2236 ^ 1'b0 ;
  assign n15988 = n13854 ^ n443 ^ 1'b0 ;
  assign n15989 = n3793 & ~n15988 ;
  assign n15990 = n15989 ^ n7734 ^ 1'b0 ;
  assign n15991 = n15987 & n15990 ;
  assign n15992 = n3878 | n9763 ;
  assign n15993 = n11673 ^ n11471 ^ 1'b0 ;
  assign n15994 = n1893 & ~n15993 ;
  assign n15995 = n553 | n1103 ;
  assign n15996 = n553 & ~n15995 ;
  assign n15997 = n1254 & n15996 ;
  assign n15998 = n1359 & n15997 ;
  assign n15999 = ~n15997 & n15998 ;
  assign n16000 = ~n1162 & n2397 ;
  assign n16001 = n1162 & n16000 ;
  assign n16002 = n16001 ^ n12304 ^ 1'b0 ;
  assign n16003 = n16002 ^ n2474 ^ 1'b0 ;
  assign n16004 = ~n15999 & n16003 ;
  assign n16005 = n7868 ^ n4379 ^ 1'b0 ;
  assign n16006 = n2848 | n16005 ;
  assign n16007 = n12873 & n16006 ;
  assign n16008 = ~n6244 & n14768 ;
  assign n16009 = n16008 ^ n7114 ^ 1'b0 ;
  assign n16010 = n3034 & ~n14258 ;
  assign n16014 = n5534 ^ n553 ^ 1'b0 ;
  assign n16015 = n2785 | n16014 ;
  assign n16011 = n1157 & ~n3038 ;
  assign n16012 = n5043 & ~n16011 ;
  assign n16013 = n16012 ^ n3892 ^ 1'b0 ;
  assign n16016 = n16015 ^ n16013 ^ 1'b0 ;
  assign n16017 = n3774 | n16016 ;
  assign n16018 = n1017 & n16017 ;
  assign n16019 = n1218 & n6897 ;
  assign n16020 = n16019 ^ n9116 ^ 1'b0 ;
  assign n16021 = ~n1098 & n16020 ;
  assign n16022 = n16021 ^ n177 ^ 1'b0 ;
  assign n16023 = ~n1572 & n3803 ;
  assign n16024 = ~n3784 & n16023 ;
  assign n16025 = n7770 & ~n10521 ;
  assign n16026 = n16025 ^ n4480 ^ 1'b0 ;
  assign n16027 = n13949 & n16026 ;
  assign n16028 = n3637 & ~n14484 ;
  assign n16029 = n16028 ^ n7489 ^ 1'b0 ;
  assign n16030 = n14181 & n15210 ;
  assign n16031 = ~n328 & n8290 ;
  assign n16032 = n7451 ^ n7395 ^ n5418 ;
  assign n16033 = n5897 | n7322 ;
  assign n16034 = n16033 ^ n1329 ^ 1'b0 ;
  assign n16035 = n14863 | n16034 ;
  assign n16036 = ~n4907 & n12547 ;
  assign n16037 = n1326 & n2839 ;
  assign n16038 = ~n1924 & n16037 ;
  assign n16039 = n16038 ^ n3088 ^ 1'b0 ;
  assign n16040 = n16039 ^ n5924 ^ 1'b0 ;
  assign n16041 = n13327 ^ n5806 ^ 1'b0 ;
  assign n16042 = ~n3849 & n16041 ;
  assign n16043 = n258 ^ n205 ^ 1'b0 ;
  assign n16044 = n9435 ^ n2270 ^ 1'b0 ;
  assign n16045 = n12225 & ~n16044 ;
  assign n16046 = ~n16043 & n16045 ;
  assign n16047 = n6730 | n10600 ;
  assign n16048 = n785 & ~n5603 ;
  assign n16049 = n1370 & n16048 ;
  assign n16050 = n588 | n16049 ;
  assign n16051 = n5389 | n6031 ;
  assign n16052 = n3940 & ~n16051 ;
  assign n16053 = n16052 ^ n8685 ^ 1'b0 ;
  assign n16054 = n5936 & ~n16053 ;
  assign n16055 = n10399 | n13357 ;
  assign n16056 = ~n566 & n13964 ;
  assign n16057 = n16056 ^ n3637 ^ 1'b0 ;
  assign n16058 = ~n1124 & n9194 ;
  assign n16059 = n284 | n481 ;
  assign n16060 = n6485 & ~n16059 ;
  assign n16061 = n11806 | n16060 ;
  assign n16062 = n55 & ~n16061 ;
  assign n16063 = n542 & ~n740 ;
  assign n16064 = ~n700 & n16063 ;
  assign n16065 = n1810 & ~n13468 ;
  assign n16066 = n16065 ^ n2633 ^ 1'b0 ;
  assign n16067 = n1390 & n10849 ;
  assign n16068 = n6011 & n11373 ;
  assign n16069 = n3116 & n16068 ;
  assign n16070 = n2880 & n12742 ;
  assign n16071 = n16070 ^ n7981 ^ 1'b0 ;
  assign n16072 = n8620 | n16071 ;
  assign n16073 = n9189 & ~n16072 ;
  assign n16074 = n5113 | n6615 ;
  assign n16075 = n86 & n1613 ;
  assign n16076 = n4977 & n16075 ;
  assign n16077 = ~n5425 & n15770 ;
  assign n16078 = n16077 ^ n3827 ^ 1'b0 ;
  assign n16079 = n1571 ^ n613 ^ 1'b0 ;
  assign n16080 = ~n8290 & n8442 ;
  assign n16081 = n16079 & n16080 ;
  assign n16082 = n16078 | n16081 ;
  assign n16083 = n6194 ^ n1406 ^ 1'b0 ;
  assign n16084 = n8763 & ~n16083 ;
  assign n16085 = n382 | n10728 ;
  assign n16086 = n16085 ^ n2382 ^ 1'b0 ;
  assign n16088 = n58 & ~n1235 ;
  assign n16087 = n1673 & ~n5754 ;
  assign n16089 = n16088 ^ n16087 ^ 1'b0 ;
  assign n16090 = n16086 | n16089 ;
  assign n16091 = n599 ^ n363 ^ 1'b0 ;
  assign n16092 = n229 & n16091 ;
  assign n16093 = ~n1528 & n3239 ;
  assign n16094 = n16093 ^ n8517 ^ n1225 ;
  assign n16095 = n3333 & n16094 ;
  assign n16096 = n5033 & n12193 ;
  assign n16097 = n16096 ^ n2672 ^ 1'b0 ;
  assign n16098 = n13120 & ~n16097 ;
  assign n16099 = n2542 & n6253 ;
  assign n16100 = n3267 & ~n7283 ;
  assign n16101 = n16100 ^ n15580 ^ n75 ;
  assign n16102 = n3311 | n12817 ;
  assign n16103 = n13265 ^ n4332 ^ 1'b0 ;
  assign n16104 = n724 & ~n16103 ;
  assign n16105 = n2003 & ~n8186 ;
  assign n16106 = n16105 ^ n8654 ^ 1'b0 ;
  assign n16107 = ~n13610 & n16106 ;
  assign n16108 = n4326 | n6553 ;
  assign n16109 = n16108 ^ n382 ^ 1'b0 ;
  assign n16110 = n1061 & ~n16109 ;
  assign n16111 = n3820 & n7231 ;
  assign n16112 = n1141 & ~n16111 ;
  assign n16113 = n16112 ^ n6270 ^ 1'b0 ;
  assign n16114 = n3878 & n7624 ;
  assign n16115 = n8732 & n16114 ;
  assign n16116 = n16113 | n16115 ;
  assign n16117 = n16116 ^ n12042 ^ 1'b0 ;
  assign n16118 = n624 | n13220 ;
  assign n16119 = n2082 & ~n9261 ;
  assign n16120 = n14147 ^ n2789 ^ 1'b0 ;
  assign n16121 = n6770 & ~n9447 ;
  assign n16122 = n16120 & n16121 ;
  assign n16123 = n1658 ^ n1304 ^ 1'b0 ;
  assign n16124 = n7110 | n16123 ;
  assign n16125 = n997 | n16124 ;
  assign n16126 = n8680 | n16125 ;
  assign n16127 = ~n8739 & n11872 ;
  assign n16128 = n3472 & n14608 ;
  assign n16129 = n2858 ^ n131 ^ 1'b0 ;
  assign n16130 = n16128 & n16129 ;
  assign n16131 = n284 & n5094 ;
  assign n16132 = n5256 & n16131 ;
  assign n16133 = n12639 ^ n3452 ^ 1'b0 ;
  assign n16134 = ~n11604 & n13842 ;
  assign n16135 = n5364 & n16134 ;
  assign n16136 = ~n7408 & n14339 ;
  assign n16137 = n16136 ^ n11346 ^ 1'b0 ;
  assign n16138 = n9351 ^ n4683 ^ 1'b0 ;
  assign n16139 = ~n1087 & n1719 ;
  assign n16140 = n16139 ^ n741 ^ 1'b0 ;
  assign n16141 = n16138 & ~n16140 ;
  assign n16142 = ~n1447 & n9223 ;
  assign n16143 = n16142 ^ n3059 ^ 1'b0 ;
  assign n16144 = n7450 & n15066 ;
  assign n16145 = n16144 ^ n5418 ^ 1'b0 ;
  assign n16146 = n12118 ^ n8963 ^ 1'b0 ;
  assign n16147 = n497 | n2542 ;
  assign n16148 = n6374 & ~n11334 ;
  assign n16149 = n16148 ^ n3857 ^ 1'b0 ;
  assign n16150 = n13585 & n16149 ;
  assign n16151 = ~n2681 & n3559 ;
  assign n16152 = n1633 & ~n10207 ;
  assign n16153 = n16152 ^ n3585 ^ 1'b0 ;
  assign n16154 = n16153 ^ n1811 ^ 1'b0 ;
  assign n16155 = n1412 & n16154 ;
  assign n16156 = ~n47 & n6333 ;
  assign n16157 = n837 & n5549 ;
  assign n16158 = n1293 & n3431 ;
  assign n16159 = n12659 ^ n2347 ^ 1'b0 ;
  assign n16160 = n16158 & n16159 ;
  assign n16161 = n2864 | n7825 ;
  assign n16162 = n7617 & n16161 ;
  assign n16163 = n2403 ^ n1283 ^ 1'b0 ;
  assign n16164 = n2633 | n10375 ;
  assign n16165 = n13795 ^ n798 ^ 1'b0 ;
  assign n16166 = n16165 ^ n1133 ^ 1'b0 ;
  assign n16167 = n14265 ^ n1845 ^ 1'b0 ;
  assign n16168 = n3569 | n14550 ;
  assign n16170 = n1380 ^ x0 ^ 1'b0 ;
  assign n16169 = ~n458 & n7140 ;
  assign n16171 = n16170 ^ n16169 ^ 1'b0 ;
  assign n16172 = n2101 & n16171 ;
  assign n16173 = n16172 ^ n12242 ^ 1'b0 ;
  assign n16175 = n3502 ^ n1663 ^ 1'b0 ;
  assign n16174 = n12458 ^ n10053 ^ 1'b0 ;
  assign n16176 = n16175 ^ n16174 ^ n5010 ;
  assign n16177 = n2313 | n12523 ;
  assign n16178 = n3063 | n16177 ;
  assign n16179 = n8739 & n12219 ;
  assign n16180 = ~n16178 & n16179 ;
  assign n16181 = ~n1263 & n4763 ;
  assign n16182 = n16181 ^ n2873 ^ 1'b0 ;
  assign n16183 = n12470 ^ n6416 ^ 1'b0 ;
  assign n16184 = n13777 | n16183 ;
  assign n16185 = n14920 ^ n1684 ^ 1'b0 ;
  assign n16186 = ( n2554 & n7490 ) | ( n2554 & n12723 ) | ( n7490 & n12723 ) ;
  assign n16187 = ~n2173 & n16186 ;
  assign n16188 = ~n12348 & n16187 ;
  assign n16189 = n859 & ~n4420 ;
  assign n16190 = n16189 ^ n1791 ^ 1'b0 ;
  assign n16191 = n2356 ^ n2326 ^ 1'b0 ;
  assign n16192 = n1224 & n16191 ;
  assign n16193 = n16192 ^ n1266 ^ 1'b0 ;
  assign n16194 = n9161 | n16193 ;
  assign n16195 = n8715 ^ n1329 ^ 1'b0 ;
  assign n16196 = ~n5194 & n16195 ;
  assign n16197 = n1565 & n13544 ;
  assign n16198 = n6433 & n16197 ;
  assign n16199 = n9556 ^ n9435 ^ 1'b0 ;
  assign n16200 = ~n364 & n16199 ;
  assign n16201 = ~n8253 & n16200 ;
  assign n16202 = n1704 & n16201 ;
  assign n16203 = n6547 ^ n724 ^ 1'b0 ;
  assign n16204 = n2595 & ~n3334 ;
  assign n16205 = n3334 & n16204 ;
  assign n16206 = n16205 ^ n4157 ^ 1'b0 ;
  assign n16207 = n3088 | n15192 ;
  assign n16208 = n8220 ^ n6017 ^ 1'b0 ;
  assign n16209 = n1384 & n16208 ;
  assign n16210 = n16209 ^ n4186 ^ 1'b0 ;
  assign n16211 = n818 & n16210 ;
  assign n16212 = n5534 | n9074 ;
  assign n16213 = n16212 ^ n15426 ^ 1'b0 ;
  assign n16214 = n731 & n16213 ;
  assign n16215 = n16214 ^ n11186 ^ 1'b0 ;
  assign n16216 = n13753 | n16215 ;
  assign n16217 = n8822 ^ n6450 ^ 1'b0 ;
  assign n16218 = n16217 ^ n849 ^ 1'b0 ;
  assign n16219 = n6835 ^ n3477 ^ 1'b0 ;
  assign n16220 = n14052 ^ n748 ^ 1'b0 ;
  assign n16221 = n8081 & ~n16220 ;
  assign n16222 = n1777 ^ n104 ^ 1'b0 ;
  assign n16223 = n283 & ~n16222 ;
  assign n16224 = n11187 & n16223 ;
  assign n16225 = ~n6871 & n10789 ;
  assign n16226 = ~n4466 & n16225 ;
  assign n16227 = n16226 ^ n1056 ^ 1'b0 ;
  assign n16228 = n2386 | n16227 ;
  assign n16229 = ~n2834 & n14444 ;
  assign n16230 = n16229 ^ n70 ^ 1'b0 ;
  assign n16231 = n16230 ^ n1728 ^ 1'b0 ;
  assign n16232 = n190 | n5253 ;
  assign n16233 = n5253 & ~n16232 ;
  assign n16234 = n16233 ^ n7265 ^ 1'b0 ;
  assign n16235 = n2261 & n16234 ;
  assign n16236 = n4181 ^ n167 ^ 1'b0 ;
  assign n16237 = n2779 ^ n2240 ^ 1'b0 ;
  assign n16238 = n7732 & n11846 ;
  assign n16239 = n16238 ^ n7947 ^ 1'b0 ;
  assign n16240 = n16239 ^ n14904 ^ 1'b0 ;
  assign n16241 = n7193 & ~n11466 ;
  assign n16242 = n16241 ^ n11136 ^ 1'b0 ;
  assign n16243 = ~n2073 & n7489 ;
  assign n16244 = n207 & n12737 ;
  assign n16245 = n1947 & n16244 ;
  assign n16246 = n16245 ^ n8460 ^ 1'b0 ;
  assign n16247 = n2491 & n4549 ;
  assign n16248 = n2068 & ~n6492 ;
  assign n16249 = ~n9745 & n16248 ;
  assign n16250 = n4774 & ~n9499 ;
  assign n16251 = ~n7263 & n12052 ;
  assign n16252 = ~n5661 & n16251 ;
  assign n16253 = ~n16250 & n16252 ;
  assign n16254 = n10788 ^ n7227 ^ 1'b0 ;
  assign n16255 = n4237 & n16254 ;
  assign n16256 = n6870 ^ n5905 ^ 1'b0 ;
  assign n16257 = n1968 & ~n16256 ;
  assign n16258 = n15368 ^ n3539 ^ 1'b0 ;
  assign n16259 = n12225 & ~n16258 ;
  assign n16260 = n13126 ^ n9108 ^ 1'b0 ;
  assign n16261 = n12234 ^ n11578 ^ 1'b0 ;
  assign n16262 = n14822 ^ n382 ^ 1'b0 ;
  assign n16263 = n4326 & n10282 ;
  assign n16264 = n11822 ^ n4446 ^ 1'b0 ;
  assign n16265 = n14093 ^ n10381 ^ 1'b0 ;
  assign n16266 = n7056 & ~n16265 ;
  assign n16267 = n8141 & n14194 ;
  assign n16268 = n1341 & n16105 ;
  assign n16269 = ~n16267 & n16268 ;
  assign n16270 = n5962 ^ n2229 ^ 1'b0 ;
  assign n16271 = n11735 ^ n6809 ^ n6071 ;
  assign n16272 = ~n16270 & n16271 ;
  assign n16273 = n592 | n11574 ;
  assign n16274 = n4819 ^ n4379 ^ 1'b0 ;
  assign n16275 = n16274 ^ n695 ^ 1'b0 ;
  assign n16276 = n4448 ^ n3931 ^ 1'b0 ;
  assign n16277 = n16276 ^ n4965 ^ 1'b0 ;
  assign n16278 = ~n9744 & n16277 ;
  assign n16279 = n16278 ^ n6186 ^ 1'b0 ;
  assign n16280 = ( n1227 & n2027 ) | ( n1227 & n5342 ) | ( n2027 & n5342 ) ;
  assign n16281 = n12357 & ~n16280 ;
  assign n16283 = n4964 ^ n643 ^ 1'b0 ;
  assign n16282 = ~n96 & n1821 ;
  assign n16284 = n16283 ^ n16282 ^ 1'b0 ;
  assign n16285 = n16284 ^ n13952 ^ 1'b0 ;
  assign n16286 = ~n5983 & n16285 ;
  assign n16287 = n8450 | n11127 ;
  assign n16288 = n16287 ^ n2071 ^ 1'b0 ;
  assign n16289 = n16288 ^ n7507 ^ n7480 ;
  assign n16290 = n1713 & n10271 ;
  assign n16291 = n16290 ^ n4644 ^ 1'b0 ;
  assign n16292 = n16291 ^ n10153 ^ 1'b0 ;
  assign n16293 = n11604 ^ n1020 ^ 1'b0 ;
  assign n16294 = n364 & n16293 ;
  assign n16295 = n9368 ^ n938 ^ 1'b0 ;
  assign n16296 = ~n3803 & n5024 ;
  assign n16297 = ~n10514 & n16296 ;
  assign n16298 = n1775 & n16297 ;
  assign n16299 = n14968 & n16298 ;
  assign n16300 = n16299 ^ n9727 ^ 1'b0 ;
  assign n16301 = n7377 & n9839 ;
  assign n16302 = n3171 ^ n1705 ^ 1'b0 ;
  assign n16303 = n1831 & n4842 ;
  assign n16304 = n6438 & ~n16303 ;
  assign n16305 = n16302 & n16304 ;
  assign n16306 = n16305 ^ n694 ^ 1'b0 ;
  assign n16307 = n2294 | n16306 ;
  assign n16308 = n8667 | n16307 ;
  assign n16309 = n250 & n1421 ;
  assign n16311 = n11888 ^ n2951 ^ 1'b0 ;
  assign n16310 = n2902 ^ n2367 ^ 1'b0 ;
  assign n16312 = n16311 ^ n16310 ^ 1'b0 ;
  assign n16313 = ~n7404 & n16312 ;
  assign n16314 = ~n4544 & n6099 ;
  assign n16315 = n16314 ^ n2046 ^ 1'b0 ;
  assign n16316 = ~n683 & n8472 ;
  assign n16317 = ~n1802 & n16316 ;
  assign n16318 = n2010 & ~n16317 ;
  assign n16319 = n16318 ^ n13424 ^ 1'b0 ;
  assign n16320 = n1095 & ~n16319 ;
  assign n16321 = n1491 ^ n157 ^ 1'b0 ;
  assign n16322 = n287 & ~n5056 ;
  assign n16323 = n1995 ^ n363 ^ 1'b0 ;
  assign n16324 = n16322 & n16323 ;
  assign n16325 = n8810 & n15796 ;
  assign n16326 = n2021 & ~n9326 ;
  assign n16327 = n4412 & n16326 ;
  assign n16328 = ~n4412 & n16327 ;
  assign n16329 = n1348 & ~n9299 ;
  assign n16330 = ~n872 & n16329 ;
  assign n16331 = n2163 & ~n8041 ;
  assign n16332 = ~n15050 & n16331 ;
  assign n16333 = ~n4449 & n16332 ;
  assign n16334 = ~n2043 & n10470 ;
  assign n16335 = ~n2362 & n9231 ;
  assign n16336 = ~n3211 & n3642 ;
  assign n16337 = n4878 & ~n6363 ;
  assign n16338 = n653 & n16337 ;
  assign n16339 = n1707 ^ n907 ^ 1'b0 ;
  assign n16340 = n7676 | n13501 ;
  assign n16341 = n2805 & n5373 ;
  assign n16342 = ~n4688 & n16341 ;
  assign n16343 = ~n6758 & n16342 ;
  assign n16344 = n8486 ^ n4501 ^ 1'b0 ;
  assign n16345 = n10887 ^ n4247 ^ 1'b0 ;
  assign n16346 = ( n10121 & n16344 ) | ( n10121 & n16345 ) | ( n16344 & n16345 ) ;
  assign n16347 = n14179 ^ n3244 ^ 1'b0 ;
  assign n16348 = n414 & n1763 ;
  assign n16349 = n8769 & n16348 ;
  assign n16350 = n7589 ^ n5225 ^ 1'b0 ;
  assign n16351 = ~n16349 & n16350 ;
  assign n16352 = n3745 ^ n2486 ^ 1'b0 ;
  assign n16353 = n10946 & ~n16352 ;
  assign n16354 = n7472 & n13326 ;
  assign n16355 = ~n7223 & n8320 ;
  assign n16356 = n1598 ^ n395 ^ 1'b0 ;
  assign n16357 = n16356 ^ n3071 ^ 1'b0 ;
  assign n16358 = n294 & n13961 ;
  assign n16359 = n13439 & ~n16358 ;
  assign n16360 = ~n1772 & n4840 ;
  assign n16361 = n10104 & n15961 ;
  assign n16362 = n6170 & n16361 ;
  assign n16363 = n1323 & n9808 ;
  assign n16364 = n10044 ^ n501 ^ 1'b0 ;
  assign n16365 = n16363 & ~n16364 ;
  assign n16366 = ~n1829 & n12709 ;
  assign n16367 = n16366 ^ n14441 ^ 1'b0 ;
  assign n16368 = n14194 | n16367 ;
  assign n16369 = n4645 ^ n3890 ^ 1'b0 ;
  assign n16370 = n9252 | n16369 ;
  assign n16371 = n4503 & ~n12126 ;
  assign n16372 = ~n216 & n4668 ;
  assign n16373 = n16372 ^ n1112 ^ 1'b0 ;
  assign n16374 = n15521 ^ n10536 ^ 1'b0 ;
  assign n16375 = n16373 | n16374 ;
  assign n16376 = n6329 & ~n14819 ;
  assign n16377 = n16376 ^ n12258 ^ 1'b0 ;
  assign n16378 = n11556 ^ n322 ^ 1'b0 ;
  assign n16379 = n16378 ^ n1455 ^ 1'b0 ;
  assign n16380 = ~n3193 & n16379 ;
  assign n16381 = ~n13048 & n16380 ;
  assign n16382 = n11763 ^ n9252 ^ 1'b0 ;
  assign n16383 = n16382 ^ n15426 ^ 1'b0 ;
  assign n16384 = n2776 & n16383 ;
  assign n16385 = n641 & n4996 ;
  assign n16386 = n1491 & n16385 ;
  assign n16387 = n629 & n10057 ;
  assign n16388 = n9638 & n16387 ;
  assign n16389 = n16386 & n16388 ;
  assign n16390 = n9422 ^ n3248 ^ 1'b0 ;
  assign n16391 = ~n7119 & n16390 ;
  assign n16392 = ~n4747 & n16391 ;
  assign n16393 = ~n448 & n16392 ;
  assign n16394 = ~n1906 & n2004 ;
  assign n16395 = n16394 ^ n867 ^ 1'b0 ;
  assign n16396 = ~n3947 & n16395 ;
  assign n16397 = n16393 & n16396 ;
  assign n16398 = n5716 & ~n6933 ;
  assign n16399 = n321 & ~n3707 ;
  assign n16400 = n6363 & n16399 ;
  assign n16401 = n622 | n8165 ;
  assign n16402 = ~n1066 & n16401 ;
  assign n16403 = n16143 | n16402 ;
  assign n16404 = n9461 & n11771 ;
  assign n16405 = n1961 & n12057 ;
  assign n16406 = n16405 ^ n11876 ^ 1'b0 ;
  assign n16407 = n13453 ^ n6400 ^ 1'b0 ;
  assign n16408 = n16407 ^ n274 ^ 1'b0 ;
  assign n16409 = n64 | n16408 ;
  assign n16410 = ( n4857 & ~n4969 ) | ( n4857 & n6331 ) | ( ~n4969 & n6331 ) ;
  assign n16411 = n16410 ^ n9561 ^ n101 ;
  assign n16412 = n6780 ^ n2687 ^ 1'b0 ;
  assign n16413 = n484 & n2929 ;
  assign n16414 = n16267 ^ n6924 ^ 1'b0 ;
  assign n16415 = n16413 | n16414 ;
  assign n16416 = n2249 & ~n7495 ;
  assign n16417 = n16416 ^ n2075 ^ 1'b0 ;
  assign n16418 = n468 & n5389 ;
  assign n16419 = n14225 ^ n1155 ^ 1'b0 ;
  assign n16420 = n16418 | n16419 ;
  assign n16421 = n2542 ^ n1924 ^ 1'b0 ;
  assign n16422 = n1089 & ~n1800 ;
  assign n16423 = n16422 ^ n14836 ^ 1'b0 ;
  assign n16424 = n2611 & n2914 ;
  assign n16425 = n12952 ^ n11496 ^ 1'b0 ;
  assign n16426 = ~n13006 & n16425 ;
  assign n16427 = n16426 ^ n9954 ^ n5686 ;
  assign n16428 = n357 | n3099 ;
  assign n16429 = n12674 ^ n3390 ^ 1'b0 ;
  assign n16430 = n390 | n1441 ;
  assign n16431 = n1506 & ~n16430 ;
  assign n16432 = n12363 & ~n16431 ;
  assign n16433 = n16432 ^ n6682 ^ 1'b0 ;
  assign n16437 = n25 & n11931 ;
  assign n16438 = n16437 ^ n3206 ^ 1'b0 ;
  assign n16439 = n6887 & n16438 ;
  assign n16440 = n16439 ^ n13556 ^ 1'b0 ;
  assign n16441 = n16440 ^ n874 ^ 1'b0 ;
  assign n16434 = n2882 | n6407 ;
  assign n16435 = n9401 & ~n16434 ;
  assign n16436 = n460 | n16435 ;
  assign n16442 = n16441 ^ n16436 ^ 1'b0 ;
  assign n16447 = n7656 ^ n3245 ^ 1'b0 ;
  assign n16448 = n175 | n16447 ;
  assign n16449 = n7431 ^ n3744 ^ n1895 ;
  assign n16450 = n83 & n2728 ;
  assign n16451 = n799 | n16450 ;
  assign n16452 = n16449 | n16451 ;
  assign n16453 = n16452 ^ n3646 ^ 1'b0 ;
  assign n16454 = n16448 | n16453 ;
  assign n16443 = n11019 ^ n919 ^ 1'b0 ;
  assign n16444 = n16443 ^ n7264 ^ 1'b0 ;
  assign n16445 = n9829 ^ n6079 ^ 1'b0 ;
  assign n16446 = n16444 & n16445 ;
  assign n16455 = n16454 ^ n16446 ^ 1'b0 ;
  assign n16456 = n1070 & ~n7909 ;
  assign n16457 = n16456 ^ n850 ^ 1'b0 ;
  assign n16458 = ( n6809 & n7660 ) | ( n6809 & n16457 ) | ( n7660 & n16457 ) ;
  assign n16459 = n5264 ^ n4326 ^ 1'b0 ;
  assign n16460 = n5554 ^ n1471 ^ 1'b0 ;
  assign n16461 = n2431 & ~n7301 ;
  assign n16462 = n233 | n12454 ;
  assign n16463 = n6464 ^ n938 ^ 1'b0 ;
  assign n16465 = ~n2771 & n9913 ;
  assign n16464 = n1089 & ~n2072 ;
  assign n16466 = n16465 ^ n16464 ^ 1'b0 ;
  assign n16467 = n16463 | n16466 ;
  assign n16468 = ( n1087 & n11360 ) | ( n1087 & n16467 ) | ( n11360 & n16467 ) ;
  assign n16469 = n11559 ^ n2371 ^ 1'b0 ;
  assign n16470 = ~n7646 & n9422 ;
  assign n16471 = ~n4864 & n4869 ;
  assign n16472 = n16471 ^ n4474 ^ 1'b0 ;
  assign n16473 = n13837 & ~n15482 ;
  assign n16474 = n13087 ^ n729 ^ 1'b0 ;
  assign n16475 = n16474 ^ n16101 ^ 1'b0 ;
  assign n16477 = ~n239 & n3758 ;
  assign n16476 = n415 & ~n3154 ;
  assign n16478 = n16477 ^ n16476 ^ 1'b0 ;
  assign n16480 = n3221 ^ n47 ^ 1'b0 ;
  assign n16479 = n2209 ^ n415 ^ 1'b0 ;
  assign n16481 = n16480 ^ n16479 ^ 1'b0 ;
  assign n16482 = n4782 & n16481 ;
  assign n16483 = n1165 & n3247 ;
  assign n16484 = n16483 ^ n3348 ^ 1'b0 ;
  assign n16485 = n9588 & n16484 ;
  assign n16486 = n8957 ^ n5727 ^ 1'b0 ;
  assign n16487 = n4436 ^ n3418 ^ 1'b0 ;
  assign n16488 = n14046 & n16126 ;
  assign n16489 = n1159 & n16488 ;
  assign n16490 = n7688 ^ n1825 ^ 1'b0 ;
  assign n16491 = n4734 ^ n3727 ^ 1'b0 ;
  assign n16492 = ~n3593 & n16491 ;
  assign n16493 = n1209 & n2239 ;
  assign n16494 = ~n2239 & n16493 ;
  assign n16495 = n2606 & ~n16494 ;
  assign n16496 = n16494 & n16495 ;
  assign n16497 = n16053 | n16496 ;
  assign n16498 = ~n6023 & n12363 ;
  assign n16499 = n16498 ^ n5444 ^ 1'b0 ;
  assign n16500 = n16497 | n16499 ;
  assign n16501 = n4077 | n14772 ;
  assign n16502 = n66 & n5338 ;
  assign n16503 = n952 | n1705 ;
  assign n16504 = n4752 & ~n16503 ;
  assign n16505 = n190 & n16504 ;
  assign n16506 = ~n1539 & n6732 ;
  assign n16507 = ~n6034 & n15485 ;
  assign n16508 = n3447 | n16507 ;
  assign n16509 = n2682 | n16508 ;
  assign n16510 = n16509 ^ n8863 ^ n470 ;
  assign n16511 = n16510 ^ n8763 ^ 1'b0 ;
  assign n16512 = n1915 & ~n11616 ;
  assign n16513 = n458 & ~n12550 ;
  assign n16514 = n8214 & n16513 ;
  assign n16515 = n16011 & n16514 ;
  assign n16516 = n16152 ^ n4169 ^ 1'b0 ;
  assign n16517 = ~n3226 & n3722 ;
  assign n16518 = n11012 & n16517 ;
  assign n16519 = n13979 ^ n823 ^ 1'b0 ;
  assign n16520 = n8984 | n9597 ;
  assign n16521 = n16520 ^ n5502 ^ 1'b0 ;
  assign n16522 = n3176 & ~n5302 ;
  assign n16523 = n16522 ^ n10265 ^ 1'b0 ;
  assign n16524 = ~n2577 & n16523 ;
  assign n16525 = n16521 & n16524 ;
  assign n16526 = n3532 & n4615 ;
  assign n16527 = ~n9284 & n16526 ;
  assign n16528 = n310 & ~n16527 ;
  assign n16529 = n6109 | n16528 ;
  assign n16530 = ~n1811 & n8036 ;
  assign n16531 = ~n6438 & n16530 ;
  assign n16532 = n16531 ^ n3356 ^ 1'b0 ;
  assign n16533 = n10973 ^ n1349 ^ 1'b0 ;
  assign n16534 = n16532 & ~n16533 ;
  assign n16535 = n16534 ^ n4548 ^ 1'b0 ;
  assign n16538 = n10859 ^ n1105 ^ 1'b0 ;
  assign n16536 = ~n328 & n703 ;
  assign n16537 = n6973 & n16536 ;
  assign n16539 = n16538 ^ n16537 ^ 1'b0 ;
  assign n16540 = n4153 & n14887 ;
  assign n16541 = ~n11698 & n16540 ;
  assign n16542 = n1349 | n4449 ;
  assign n16543 = n7126 & ~n16542 ;
  assign n16544 = n9077 | n12689 ;
  assign n16548 = ~n1744 & n14439 ;
  assign n16546 = n7481 & n7586 ;
  assign n16547 = n3861 & ~n16546 ;
  assign n16549 = n16548 ^ n16547 ^ 1'b0 ;
  assign n16545 = n4482 | n11204 ;
  assign n16550 = n16549 ^ n16545 ^ 1'b0 ;
  assign n16551 = ~n1794 & n1937 ;
  assign n16552 = n16551 ^ n12171 ^ 1'b0 ;
  assign n16553 = n4548 ^ n2397 ^ 1'b0 ;
  assign n16554 = n7194 | n16553 ;
  assign n16555 = n1467 & ~n2311 ;
  assign n16556 = ~n8149 & n16555 ;
  assign n16557 = n8027 ^ n30 ^ 1'b0 ;
  assign n16558 = n6188 & n16557 ;
  assign n16559 = n7753 | n11835 ;
  assign n16560 = n2951 | n16559 ;
  assign n16561 = n16560 ^ n2558 ^ 1'b0 ;
  assign n16562 = ~n13437 & n14195 ;
  assign n16563 = n16562 ^ n598 ^ 1'b0 ;
  assign n16564 = n5065 | n16563 ;
  assign n16565 = ~n7129 & n16564 ;
  assign n16566 = n2032 & n10261 ;
  assign n16567 = n1588 | n11578 ;
  assign n16568 = n16567 ^ n294 ^ 1'b0 ;
  assign n16569 = n1745 & ~n2943 ;
  assign n16570 = n16569 ^ n15210 ^ 1'b0 ;
  assign n16571 = n14611 & n16570 ;
  assign n16572 = n16571 ^ n1699 ^ n321 ;
  assign n16573 = n616 ^ n469 ^ 1'b0 ;
  assign n16574 = n10064 & ~n16573 ;
  assign n16575 = n16574 ^ n257 ^ 1'b0 ;
  assign n16576 = ~n1027 & n2973 ;
  assign n16577 = n16576 ^ n9673 ^ 1'b0 ;
  assign n16578 = n1414 & ~n16577 ;
  assign n16579 = n16578 ^ n8971 ^ 1'b0 ;
  assign n16580 = n5990 & ~n10943 ;
  assign n16581 = n2021 & ~n4085 ;
  assign n16582 = n16581 ^ n7290 ^ 1'b0 ;
  assign n16583 = n4155 & ~n13116 ;
  assign n16584 = n16583 ^ n12059 ^ 1'b0 ;
  assign n16585 = n549 & ~n1865 ;
  assign n16586 = ~n1835 & n5714 ;
  assign n16587 = n468 | n8261 ;
  assign n16588 = n6272 & ~n16587 ;
  assign n16589 = n3489 ^ n1833 ^ 1'b0 ;
  assign n16590 = n3044 & n16589 ;
  assign n16591 = n16590 ^ n8499 ^ 1'b0 ;
  assign n16592 = n15255 ^ n694 ^ 1'b0 ;
  assign n16593 = n7580 & n16592 ;
  assign n16594 = n14669 & ~n16593 ;
  assign n16595 = n1096 ^ n635 ^ 1'b0 ;
  assign n16596 = ~n16594 & n16595 ;
  assign n16600 = n1818 ^ n656 ^ 1'b0 ;
  assign n16601 = n3373 | n16600 ;
  assign n16602 = n3320 & ~n16601 ;
  assign n16603 = n7988 & n16602 ;
  assign n16597 = n2566 & ~n5663 ;
  assign n16598 = n3206 & n16597 ;
  assign n16599 = n539 | n16598 ;
  assign n16604 = n16603 ^ n16599 ^ 1'b0 ;
  assign n16605 = n16604 ^ n10879 ^ 1'b0 ;
  assign n16606 = ~n1370 & n16605 ;
  assign n16607 = n2556 & ~n3369 ;
  assign n16608 = n7151 & n16607 ;
  assign n16609 = n1349 & n16608 ;
  assign n16610 = n2110 | n16609 ;
  assign n16611 = n2681 ^ n158 ^ 1'b0 ;
  assign n16612 = n13008 ^ n950 ^ n891 ;
  assign n16613 = n12269 ^ n5930 ^ 1'b0 ;
  assign n16614 = n6731 & n10759 ;
  assign n16615 = n16614 ^ n4527 ^ 1'b0 ;
  assign n16616 = n6746 & n14394 ;
  assign n16617 = n789 & n16616 ;
  assign n16618 = ~n1933 & n2701 ;
  assign n16619 = n16618 ^ n2092 ^ 1'b0 ;
  assign n16620 = n759 | n16619 ;
  assign n16621 = n16620 ^ n1064 ^ 1'b0 ;
  assign n16622 = n2269 | n10014 ;
  assign n16623 = n3249 | n16622 ;
  assign n16624 = n5547 ^ n988 ^ 1'b0 ;
  assign n16625 = n4976 | n16624 ;
  assign n16626 = n3452 & ~n16625 ;
  assign n16627 = ~n16623 & n16626 ;
  assign n16628 = n1502 & ~n1800 ;
  assign n16629 = n16628 ^ n2155 ^ 1'b0 ;
  assign n16630 = n16629 ^ n4176 ^ 1'b0 ;
  assign n16631 = n8830 & ~n13706 ;
  assign n16632 = ~n5551 & n5817 ;
  assign n16633 = n348 | n1447 ;
  assign n16634 = ( n595 & n2682 ) | ( n595 & ~n9349 ) | ( n2682 & ~n9349 ) ;
  assign n16635 = n16421 ^ n7383 ^ n128 ;
  assign n16636 = n314 & n2514 ;
  assign n16637 = n8813 & ~n16636 ;
  assign n16638 = n16637 ^ n1026 ^ 1'b0 ;
  assign n16639 = ~n638 & n8309 ;
  assign n16640 = n8318 ^ n4112 ^ 1'b0 ;
  assign n16641 = n9211 & n10181 ;
  assign n16642 = n7269 ^ n3514 ^ 1'b0 ;
  assign n16643 = n6250 & ~n16642 ;
  assign n16644 = ~n7253 & n16643 ;
  assign n16645 = n16644 ^ n7596 ^ 1'b0 ;
  assign n16646 = n12039 & ~n16645 ;
  assign n16647 = n4315 ^ n782 ^ 1'b0 ;
  assign n16648 = n16647 ^ n3796 ^ 1'b0 ;
  assign n16649 = n4893 ^ n2736 ^ 1'b0 ;
  assign n16650 = ~n3484 & n16649 ;
  assign n16652 = n553 & ~n8891 ;
  assign n16651 = n6348 ^ n2440 ^ 1'b0 ;
  assign n16653 = n16652 ^ n16651 ^ 1'b0 ;
  assign n16654 = n16653 ^ n4568 ^ 1'b0 ;
  assign n16655 = n16654 ^ n137 ^ 1'b0 ;
  assign n16656 = n469 ^ n28 ^ 1'b0 ;
  assign n16657 = n512 | n16656 ;
  assign n16658 = n5525 & n12194 ;
  assign n16659 = n16657 & n16658 ;
  assign n16660 = n3663 & ~n4787 ;
  assign n16661 = n7268 & ~n16660 ;
  assign n16662 = ~n4315 & n9523 ;
  assign n16663 = n16662 ^ n2154 ^ 1'b0 ;
  assign n16664 = n14622 & ~n14680 ;
  assign n16665 = ~n14622 & n16664 ;
  assign n16666 = n16665 ^ n2136 ^ 1'b0 ;
  assign n16667 = n1720 ^ n178 ^ 1'b0 ;
  assign n16668 = n767 & ~n16667 ;
  assign n16669 = ~n9424 & n16668 ;
  assign n16670 = n16669 ^ n10322 ^ 1'b0 ;
  assign n16671 = n787 & n1839 ;
  assign n16672 = n566 | n16671 ;
  assign n16673 = n3594 & ~n4513 ;
  assign n16674 = ~n9902 & n16673 ;
  assign n16675 = ( n9234 & ~n11065 ) | ( n9234 & n14928 ) | ( ~n11065 & n14928 ) ;
  assign n16676 = n1339 & n1968 ;
  assign n16677 = n16676 ^ n8277 ^ 1'b0 ;
  assign n16678 = n2994 & ~n16677 ;
  assign n16679 = n1878 & ~n16678 ;
  assign n16680 = n16679 ^ n9263 ^ 1'b0 ;
  assign n16681 = ( n1360 & n5301 ) | ( n1360 & ~n5314 ) | ( n5301 & ~n5314 ) ;
  assign n16682 = n16681 ^ n2542 ^ 1'b0 ;
  assign n16683 = ~n1739 & n13855 ;
  assign n16684 = n7671 & ~n16683 ;
  assign n16686 = ~n3095 & n12673 ;
  assign n16685 = n6348 & n15483 ;
  assign n16687 = n16686 ^ n16685 ^ 1'b0 ;
  assign n16688 = n5280 ^ n2235 ^ 1'b0 ;
  assign n16689 = ~n11504 & n16688 ;
  assign n16690 = n1083 & n6573 ;
  assign n16691 = n16690 ^ n2141 ^ 1'b0 ;
  assign n16692 = n6185 & n16691 ;
  assign n16693 = n7327 & n16692 ;
  assign n16694 = n16693 ^ n12265 ^ 1'b0 ;
  assign n16695 = n15 | n16694 ;
  assign n16696 = n3526 & n7245 ;
  assign n16697 = ~n6579 & n16696 ;
  assign n16698 = n5332 ^ n1323 ^ 1'b0 ;
  assign n16699 = n16697 | n16698 ;
  assign n16700 = ~n4025 & n14863 ;
  assign n16702 = n4045 & n6421 ;
  assign n16703 = ~n1358 & n16702 ;
  assign n16701 = n15200 ^ n13461 ^ 1'b0 ;
  assign n16704 = n16703 ^ n16701 ^ n1915 ;
  assign n16705 = n2029 & ~n16704 ;
  assign n16706 = n2999 | n5868 ;
  assign n16707 = ~n10105 & n16706 ;
  assign n16708 = n16707 ^ n1105 ^ 1'b0 ;
  assign n16709 = n10836 ^ n8363 ^ 1'b0 ;
  assign n16710 = ~n16126 & n16709 ;
  assign n16711 = n12353 ^ n5427 ^ 1'b0 ;
  assign n16712 = ~n3151 & n16711 ;
  assign n16713 = n15537 ^ n1017 ^ n234 ;
  assign n16714 = n919 & n10909 ;
  assign n16715 = n16714 ^ n4889 ^ 1'b0 ;
  assign n16716 = n15093 | n16715 ;
  assign n16717 = n1794 & ~n8536 ;
  assign n16718 = n5205 ^ n1165 ^ 1'b0 ;
  assign n16719 = n16717 & ~n16718 ;
  assign n16720 = n16719 ^ n2369 ^ 1'b0 ;
  assign n16721 = n6622 & ~n16720 ;
  assign n16722 = n1080 ^ n227 ^ 1'b0 ;
  assign n16723 = n10962 ^ n8216 ^ 1'b0 ;
  assign n16724 = n16722 | n16723 ;
  assign n16725 = n9930 | n16724 ;
  assign n16726 = x9 | n16725 ;
  assign n16727 = n4125 ^ n1320 ^ 1'b0 ;
  assign n16728 = n2796 & n16727 ;
  assign n16729 = ~n852 & n16728 ;
  assign n16730 = n1372 ^ n376 ^ 1'b0 ;
  assign n16731 = n4591 ^ n30 ^ 1'b0 ;
  assign n16732 = n2814 | n16731 ;
  assign n16733 = n16732 ^ n13852 ^ 1'b0 ;
  assign n16734 = ~n11714 & n16733 ;
  assign n16735 = ~n16730 & n16734 ;
  assign n16736 = n3438 | n4419 ;
  assign n16737 = n7678 & ~n12523 ;
  assign n16738 = n16737 ^ n6735 ^ 1'b0 ;
  assign n16739 = ~n14331 & n16738 ;
  assign n16740 = n1355 & n15479 ;
  assign n16741 = n8314 | n15231 ;
  assign n16742 = n2847 ^ n2352 ^ 1'b0 ;
  assign n16743 = ~n14910 & n15783 ;
  assign n16744 = ~n16742 & n16743 ;
  assign n16745 = n1934 ^ n715 ^ 1'b0 ;
  assign n16746 = n1245 | n16745 ;
  assign n16747 = n11630 | n16746 ;
  assign n16748 = n16747 ^ n7288 ^ 1'b0 ;
  assign n16750 = n731 ^ n274 ^ 1'b0 ;
  assign n16749 = n2479 & ~n7696 ;
  assign n16751 = n16750 ^ n16749 ^ 1'b0 ;
  assign n16752 = n78 & ~n16751 ;
  assign n16753 = n16752 ^ n6060 ^ 1'b0 ;
  assign n16754 = n1173 & ~n16753 ;
  assign n16755 = n9811 ^ n7693 ^ n6462 ;
  assign n16756 = n16755 ^ n11205 ^ 1'b0 ;
  assign n16757 = n6011 & n16756 ;
  assign n16758 = n16313 ^ n1307 ^ 1'b0 ;
  assign n16759 = ~n804 & n5776 ;
  assign n16760 = ~n14601 & n16759 ;
  assign n16763 = n8286 & ~n10255 ;
  assign n16764 = n16763 ^ n632 ^ 1'b0 ;
  assign n16761 = n561 | n1581 ;
  assign n16762 = n16761 ^ n1817 ^ 1'b0 ;
  assign n16765 = n16764 ^ n16762 ^ 1'b0 ;
  assign n16766 = n3624 | n7737 ;
  assign n16767 = n13820 | n16766 ;
  assign n16768 = n13099 ^ n6318 ^ 1'b0 ;
  assign n16769 = ~n12168 & n16768 ;
  assign n16773 = ~n4169 & n9952 ;
  assign n16770 = ~n43 & n333 ;
  assign n16771 = ~n4753 & n16770 ;
  assign n16772 = ~n419 & n16771 ;
  assign n16774 = n16773 ^ n16772 ^ 1'b0 ;
  assign n16775 = n6545 & n15853 ;
  assign n16777 = n5205 & n7616 ;
  assign n16778 = n4400 ^ n2567 ^ 1'b0 ;
  assign n16779 = n16777 & ~n16778 ;
  assign n16776 = n4867 & ~n10644 ;
  assign n16780 = n16779 ^ n16776 ^ 1'b0 ;
  assign n16781 = ~n5780 & n10931 ;
  assign n16782 = n16781 ^ n8030 ^ 1'b0 ;
  assign n16783 = ~n15546 & n16782 ;
  assign n16784 = n16783 ^ n4422 ^ 1'b0 ;
  assign n16785 = n323 | n5621 ;
  assign n16786 = n16785 ^ n281 ^ 1'b0 ;
  assign n16787 = n16786 ^ n12252 ^ 1'b0 ;
  assign n16788 = n11479 ^ n419 ^ 1'b0 ;
  assign n16789 = n11609 | n16788 ;
  assign n16790 = n16789 ^ n208 ^ 1'b0 ;
  assign n16791 = n1168 ^ x0 ^ 1'b0 ;
  assign n16792 = n4179 ^ n535 ^ 1'b0 ;
  assign n16793 = n3211 & n16792 ;
  assign n16794 = n5626 & n16793 ;
  assign n16795 = n1165 | n3354 ;
  assign n16796 = n16795 ^ n2558 ^ 1'b0 ;
  assign n16797 = n5031 | n9291 ;
  assign n16798 = n5128 | n16797 ;
  assign n16799 = n16798 ^ n12964 ^ 1'b0 ;
  assign n16801 = ~n2391 & n8183 ;
  assign n16802 = ~n483 & n8117 ;
  assign n16803 = n16801 & n16802 ;
  assign n16800 = ~n8760 & n14334 ;
  assign n16804 = n16803 ^ n16800 ^ n4189 ;
  assign n16805 = n188 | n3423 ;
  assign n16806 = n535 & ~n5955 ;
  assign n16807 = n16806 ^ n9197 ^ 1'b0 ;
  assign n16808 = n3891 ^ n553 ^ 1'b0 ;
  assign n16809 = n16808 ^ n1645 ^ 1'b0 ;
  assign n16810 = n4220 & ~n16809 ;
  assign n16811 = ~n16807 & n16810 ;
  assign n16812 = ~n16805 & n16811 ;
  assign n16813 = n908 & n1880 ;
  assign n16814 = n13324 ^ n11239 ^ 1'b0 ;
  assign n16815 = n12511 & ~n16814 ;
  assign n16816 = n16813 & n16815 ;
  assign n16817 = n581 | n7930 ;
  assign n16818 = n7545 | n16817 ;
  assign n16819 = n11908 ^ n10584 ^ n3120 ;
  assign n16820 = n10879 ^ n4508 ^ n3057 ;
  assign n16821 = n3154 & n16820 ;
  assign n16822 = n8827 ^ n2119 ^ n84 ;
  assign n16823 = n2799 & n16822 ;
  assign n16824 = n16823 ^ n1571 ^ 1'b0 ;
  assign n16825 = n3980 | n10035 ;
  assign n16830 = n1273 | n2618 ;
  assign n16826 = n4328 & n4336 ;
  assign n16827 = n16826 ^ n10936 ^ n1994 ;
  assign n16828 = n5514 | n16827 ;
  assign n16829 = ~n16126 & n16828 ;
  assign n16831 = n16830 ^ n16829 ^ 1'b0 ;
  assign n16832 = n13578 ^ n3123 ^ 1'b0 ;
  assign n16833 = n1645 & ~n10923 ;
  assign n16834 = n4221 | n7289 ;
  assign n16835 = ~n4733 & n16834 ;
  assign n16836 = n11646 ^ n9852 ^ 1'b0 ;
  assign n16837 = n16835 & n16836 ;
  assign n16838 = n1722 & n8165 ;
  assign n16839 = n5075 | n16838 ;
  assign n16840 = n227 & ~n16839 ;
  assign n16841 = n630 & ~n16840 ;
  assign n16842 = ~n216 & n16841 ;
  assign n16843 = n3019 | n16842 ;
  assign n16844 = ~n4577 & n6194 ;
  assign n16845 = n7371 & n16844 ;
  assign n16846 = n1777 & ~n5284 ;
  assign n16847 = n16846 ^ n6722 ^ 1'b0 ;
  assign n16848 = ~n6761 & n13532 ;
  assign n16849 = ~n5413 & n16848 ;
  assign n16850 = n16849 ^ n11155 ^ n602 ;
  assign n16851 = n491 | n914 ;
  assign n16852 = n4169 & n14376 ;
  assign n16853 = n2339 | n14370 ;
  assign n16854 = n1331 | n5863 ;
  assign n16855 = n1271 | n16854 ;
  assign n16856 = ~n12027 & n16855 ;
  assign n16857 = n5148 & n16856 ;
  assign n16858 = n16857 ^ n10691 ^ 1'b0 ;
  assign n16859 = n436 | n1348 ;
  assign n16860 = n16859 ^ n14481 ^ 1'b0 ;
  assign n16861 = n616 | n9342 ;
  assign n16862 = n16860 | n16861 ;
  assign n16863 = ~n307 & n16862 ;
  assign n16864 = n307 & n16863 ;
  assign n16865 = n6021 & n16864 ;
  assign n16866 = ~n3149 & n9486 ;
  assign n16867 = n3149 & n16866 ;
  assign n16868 = n5040 | n15042 ;
  assign n16869 = n15042 & ~n16868 ;
  assign n16870 = n16867 & ~n16869 ;
  assign n16871 = n12979 & n16870 ;
  assign n16872 = n5826 & ~n16871 ;
  assign n16873 = ~n5826 & n16872 ;
  assign n16874 = ~n1162 & n2856 ;
  assign n16875 = ~n2856 & n16874 ;
  assign n16876 = n16873 | n16875 ;
  assign n16877 = n16873 & ~n16876 ;
  assign n16878 = n1146 & ~n16877 ;
  assign n16879 = ~n1146 & n16878 ;
  assign n16880 = n16865 | n16879 ;
  assign n16881 = n16865 & ~n16880 ;
  assign n16882 = n487 & ~n1707 ;
  assign n16883 = n12716 & n16882 ;
  assign n16884 = n16883 ^ n2817 ^ 1'b0 ;
  assign n16885 = n1416 | n2937 ;
  assign n16886 = ~n167 & n495 ;
  assign n16887 = ~n495 & n16886 ;
  assign n16888 = n125 | n16887 ;
  assign n16889 = n125 & ~n16888 ;
  assign n16890 = n16889 ^ n713 ^ 1'b0 ;
  assign n16891 = n16890 ^ n1933 ^ 1'b0 ;
  assign n16892 = n1061 | n16891 ;
  assign n16893 = n6538 & ~n16892 ;
  assign n16894 = n16893 ^ n4560 ^ 1'b0 ;
  assign n16895 = n16885 | n16894 ;
  assign n16897 = n8789 ^ n1368 ^ 1'b0 ;
  assign n16898 = ~n7254 & n16897 ;
  assign n16896 = ~n52 & n185 ;
  assign n16899 = n16898 ^ n16896 ^ 1'b0 ;
  assign n16900 = n16895 | n16899 ;
  assign n16901 = n6646 & ~n8181 ;
  assign n16902 = n16901 ^ n3320 ^ 1'b0 ;
  assign n16903 = n3739 & n16902 ;
  assign n16904 = n104 | n13546 ;
  assign n16905 = n16904 ^ n2923 ^ 1'b0 ;
  assign n16906 = n3033 | n11178 ;
  assign n16907 = n5361 & ~n5409 ;
  assign n16908 = n16906 & n16907 ;
  assign n16909 = n83 & ~n7862 ;
  assign n16910 = n2012 & n10751 ;
  assign n16911 = n16910 ^ n632 ^ 1'b0 ;
  assign n16912 = n16911 ^ n1831 ^ 1'b0 ;
  assign n16913 = n3604 & n16912 ;
  assign n16914 = n1851 ^ n570 ^ 1'b0 ;
  assign n16915 = n14990 ^ n12883 ^ 1'b0 ;
  assign n16916 = n16452 & n16915 ;
  assign n16917 = ~n2819 & n5040 ;
  assign n16918 = n10893 & n16917 ;
  assign n16919 = n3334 | n5542 ;
  assign n16920 = n3311 | n5161 ;
  assign n16921 = n16920 ^ n2150 ^ 1'b0 ;
  assign n16922 = n16921 ^ n4127 ^ 1'b0 ;
  assign n16923 = n649 | n15537 ;
  assign n16924 = n1100 | n1339 ;
  assign n16925 = n16923 | n16924 ;
  assign n16926 = ~n3100 & n6602 ;
  assign n16927 = n12929 | n13366 ;
  assign n16928 = n16926 & ~n16927 ;
  assign n16929 = n3254 & ~n7011 ;
  assign n16930 = n10583 & n16929 ;
  assign n16931 = n4743 ^ n2917 ^ 1'b0 ;
  assign n16932 = n232 & ~n16931 ;
  assign n16934 = ~n483 & n2284 ;
  assign n16935 = ~n2284 & n16934 ;
  assign n16936 = n16935 ^ n7416 ^ 1'b0 ;
  assign n16933 = n7523 & ~n9815 ;
  assign n16937 = n16936 ^ n16933 ^ 1'b0 ;
  assign n16938 = n7344 & n16937 ;
  assign n16939 = n14865 ^ n8081 ^ 1'b0 ;
  assign n16940 = n638 & n16939 ;
  assign n16941 = ~n11588 & n15783 ;
  assign n16942 = n16941 ^ n7425 ^ 1'b0 ;
  assign n16943 = n7685 & n7954 ;
  assign n16944 = n16943 ^ n7646 ^ 1'b0 ;
  assign n16945 = n15652 | n16944 ;
  assign n16946 = n6150 & ~n15509 ;
  assign n16947 = n2512 & ~n7454 ;
  assign n16948 = n8845 ^ n7038 ^ 1'b0 ;
  assign n16949 = n6897 & ~n16948 ;
  assign n16950 = n16949 ^ n5261 ^ 1'b0 ;
  assign n16951 = n16947 & n16950 ;
  assign n16952 = n2289 & ~n16951 ;
  assign n16953 = n4916 ^ n390 ^ 1'b0 ;
  assign n16954 = n7604 & n16953 ;
  assign n16955 = ~n2301 & n16954 ;
  assign n16956 = n9714 & n16955 ;
  assign n16957 = n10130 | n16956 ;
  assign n16958 = n1148 & ~n16957 ;
  assign n16959 = n941 | n16958 ;
  assign n16960 = n16959 ^ n3033 ^ 1'b0 ;
  assign n16961 = n4404 | n6076 ;
  assign n16962 = n16961 ^ n9729 ^ 1'b0 ;
  assign n16963 = n7179 & n16962 ;
  assign n16964 = n10340 ^ n475 ^ 1'b0 ;
  assign n16965 = ~n10303 & n16964 ;
  assign n16966 = n2273 & ~n14161 ;
  assign n16967 = n3980 & ~n8632 ;
  assign n16968 = n636 ^ n268 ^ 1'b0 ;
  assign n16969 = n6008 & ~n16968 ;
  assign n16970 = n1303 | n16969 ;
  assign n16971 = n16970 ^ n1137 ^ 1'b0 ;
  assign n16972 = n1668 & ~n10303 ;
  assign n16973 = n6762 & n16972 ;
  assign n16974 = ~n38 & n16973 ;
  assign n16975 = n1082 ^ n178 ^ 1'b0 ;
  assign n16976 = n190 & ~n16627 ;
  assign n16977 = n16975 & n16976 ;
  assign n16978 = n8864 ^ n2733 ^ 1'b0 ;
  assign n16979 = n434 & ~n16978 ;
  assign n16980 = ~n274 & n15255 ;
  assign n16981 = n16979 & n16980 ;
  assign n16982 = n15203 | n16981 ;
  assign n16986 = n489 ^ n294 ^ 1'b0 ;
  assign n16987 = n5752 & ~n16986 ;
  assign n16988 = n3609 & n16987 ;
  assign n16983 = n48 | n15439 ;
  assign n16984 = n16983 ^ n6885 ^ 1'b0 ;
  assign n16985 = n198 | n16984 ;
  assign n16989 = n16988 ^ n16985 ^ 1'b0 ;
  assign n16990 = n4193 ^ n2870 ^ 1'b0 ;
  assign n16991 = ~n3423 & n6642 ;
  assign n16992 = n2205 & n16991 ;
  assign n16993 = ~n16990 & n16992 ;
  assign n16997 = n5488 & ~n10190 ;
  assign n16998 = n1268 & n4416 ;
  assign n16999 = n16997 & n16998 ;
  assign n17000 = ~n3227 & n9831 ;
  assign n17001 = n17000 ^ n15640 ^ 1'b0 ;
  assign n17002 = ( n2403 & n16999 ) | ( n2403 & n17001 ) | ( n16999 & n17001 ) ;
  assign n16994 = n444 | n7608 ;
  assign n16995 = n4085 | n16994 ;
  assign n16996 = ~n2623 & n16995 ;
  assign n17003 = n17002 ^ n16996 ^ n5826 ;
  assign n17004 = n17003 ^ n8410 ^ n1798 ;
  assign n17005 = n17004 ^ n4155 ^ 1'b0 ;
  assign n17006 = n1620 | n17005 ;
  assign n17007 = ~n621 & n5502 ;
  assign n17008 = ~n1733 & n2556 ;
  assign n17009 = n17007 | n17008 ;
  assign n17010 = n6762 & ~n13017 ;
  assign n17011 = ~n8714 & n17010 ;
  assign n17012 = n17009 & n17011 ;
  assign n17013 = ~n410 & n17012 ;
  assign n17015 = n12704 ^ n4059 ^ 1'b0 ;
  assign n17016 = n10624 & ~n17015 ;
  assign n17014 = ~n891 & n10942 ;
  assign n17017 = n17016 ^ n17014 ^ 1'b0 ;
  assign n17018 = n9860 ^ n1880 ^ n194 ;
  assign n17019 = n3933 & ~n13892 ;
  assign n17020 = n800 & n2137 ;
  assign n17021 = n12039 | n17020 ;
  assign n17022 = n17021 ^ n7506 ^ 1'b0 ;
  assign n17023 = n4403 & n10195 ;
  assign n17024 = n17023 ^ n5789 ^ 1'b0 ;
  assign n17025 = n17022 & ~n17024 ;
  assign n17026 = n7574 ^ n6449 ^ 1'b0 ;
  assign n17031 = n8767 ^ n6730 ^ 1'b0 ;
  assign n17027 = n5284 ^ n4611 ^ 1'b0 ;
  assign n17028 = n2589 ^ n1201 ^ 1'b0 ;
  assign n17029 = ~n460 & n17028 ;
  assign n17030 = ~n17027 & n17029 ;
  assign n17032 = n17031 ^ n17030 ^ 1'b0 ;
  assign n17033 = n2839 & ~n17032 ;
  assign n17035 = n10664 ^ n122 ^ 1'b0 ;
  assign n17036 = ~n8167 & n17035 ;
  assign n17034 = ~n5842 & n10367 ;
  assign n17037 = n17036 ^ n17034 ^ 1'b0 ;
  assign n17038 = n7403 ^ n3221 ^ 1'b0 ;
  assign n17039 = n17038 ^ n1399 ^ 1'b0 ;
  assign n17040 = n10682 & ~n17039 ;
  assign n17041 = ~n741 & n15047 ;
  assign n17042 = ~n351 & n17041 ;
  assign n17043 = n4919 ^ n414 ^ 1'b0 ;
  assign n17044 = n17042 | n17043 ;
  assign n17045 = n7980 ^ n4937 ^ 1'b0 ;
  assign n17046 = n17045 ^ n10050 ^ 1'b0 ;
  assign n17047 = ~n17044 & n17046 ;
  assign n17048 = n17047 ^ n5389 ^ 1'b0 ;
  assign n17051 = n1918 | n7406 ;
  assign n17052 = n86 & ~n17051 ;
  assign n17049 = n327 & n922 ;
  assign n17050 = ~n6017 & n17049 ;
  assign n17053 = n17052 ^ n17050 ^ 1'b0 ;
  assign n17054 = n5205 ^ n3036 ^ 1'b0 ;
  assign n17055 = n2639 | n17054 ;
  assign n17056 = n11985 ^ n8639 ^ 1'b0 ;
  assign n17057 = n567 ^ n148 ^ 1'b0 ;
  assign n17058 = ( n37 & ~n10377 ) | ( n37 & n17057 ) | ( ~n10377 & n17057 ) ;
  assign n17059 = n4296 & ~n17058 ;
  assign n17060 = n2611 ^ n253 ^ 1'b0 ;
  assign n17061 = n4679 | n8084 ;
  assign n17062 = n7431 | n15707 ;
  assign n17063 = n17061 | n17062 ;
  assign n17064 = n3540 | n14044 ;
  assign n17065 = n14869 & n16993 ;
  assign n17066 = ( n2424 & n3356 ) | ( n2424 & ~n9736 ) | ( n3356 & ~n9736 ) ;
  assign n17067 = n817 | n3435 ;
  assign n17068 = ~n7116 & n17067 ;
  assign n17069 = ~n2495 & n7590 ;
  assign n17070 = n11421 | n15241 ;
  assign n17071 = n12078 & n12376 ;
  assign n17072 = n7056 ^ n760 ^ 1'b0 ;
  assign n17073 = ~n1904 & n17072 ;
  assign n17074 = n28 | n3080 ;
  assign n17075 = n1766 | n8067 ;
  assign n17081 = n73 & n433 ;
  assign n17082 = n375 & n17081 ;
  assign n17083 = n17082 ^ n671 ^ 1'b0 ;
  assign n17076 = n419 | n2924 ;
  assign n17077 = n419 & ~n17076 ;
  assign n17078 = n5308 ^ n2364 ^ 1'b0 ;
  assign n17079 = n17077 & n17078 ;
  assign n17080 = ~n5661 & n17079 ;
  assign n17084 = n17083 ^ n17080 ^ 1'b0 ;
  assign n17085 = n17084 ^ n1406 ^ 1'b0 ;
  assign n17086 = n3640 | n16750 ;
  assign n17087 = ~n4421 & n4584 ;
  assign n17088 = n17087 ^ n13801 ^ 1'b0 ;
  assign n17089 = n11263 ^ n2977 ^ 1'b0 ;
  assign n17090 = n6229 ^ n175 ^ 1'b0 ;
  assign n17091 = n17090 ^ n14897 ^ 1'b0 ;
  assign n17092 = ~n6065 & n17091 ;
  assign n17093 = n13155 ^ n10651 ^ 1'b0 ;
  assign n17094 = n3670 ^ n2161 ^ 1'b0 ;
  assign n17095 = n3433 | n6753 ;
  assign n17096 = n17095 ^ n15775 ^ 1'b0 ;
  assign n17097 = n14462 & n16931 ;
  assign n17098 = n17096 & ~n17097 ;
  assign n17099 = n1385 & ~n2903 ;
  assign n17100 = n17099 ^ n83 ^ 1'b0 ;
  assign n17101 = n17100 ^ n9649 ^ 1'b0 ;
  assign n17102 = n679 & n3907 ;
  assign n17103 = ~n10677 & n17102 ;
  assign n17104 = n4893 & n8341 ;
  assign n17105 = n17104 ^ n2112 ^ 1'b0 ;
  assign n17106 = ~n11002 & n17105 ;
  assign n17107 = n5130 ^ n3064 ^ 1'b0 ;
  assign n17108 = n446 | n17107 ;
  assign n17109 = n542 & n4560 ;
  assign n17110 = n17109 ^ n9592 ^ n8617 ;
  assign n17111 = n13203 ^ n2362 ^ 1'b0 ;
  assign n17112 = n7609 & ~n11611 ;
  assign n17113 = n6323 ^ n454 ^ 1'b0 ;
  assign n17114 = n804 & ~n1151 ;
  assign n17115 = n8586 & ~n17114 ;
  assign n17116 = n6098 ^ n2260 ^ 1'b0 ;
  assign n17117 = n627 & n17116 ;
  assign n17118 = n11071 & n17117 ;
  assign n17119 = n1707 & ~n17118 ;
  assign n17120 = n328 & n2953 ;
  assign n17121 = n17120 ^ n5283 ^ n4939 ;
  assign n17122 = n6704 & ~n17121 ;
  assign n17123 = n5428 | n9957 ;
  assign n17124 = n17122 & ~n17123 ;
  assign n17125 = ~n16251 & n17124 ;
  assign n17127 = n957 & ~n10928 ;
  assign n17126 = n13983 ^ n8409 ^ 1'b0 ;
  assign n17128 = n17127 ^ n17126 ^ 1'b0 ;
  assign n17129 = n9646 ^ n8000 ^ 1'b0 ;
  assign n17130 = n5465 | n17129 ;
  assign n17131 = n15987 & n16949 ;
  assign n17132 = n17131 ^ n9954 ^ 1'b0 ;
  assign n17133 = n4483 & n5370 ;
  assign n17134 = n17133 ^ n517 ^ 1'b0 ;
  assign n17135 = ~n17003 & n17134 ;
  assign n17136 = n17135 ^ n15605 ^ 1'b0 ;
  assign n17137 = n6954 | n17136 ;
  assign n17138 = n8445 & n11378 ;
  assign n17139 = n7750 ^ n1668 ^ 1'b0 ;
  assign n17140 = n17138 & ~n17139 ;
  assign n17141 = ~n894 & n3415 ;
  assign n17142 = ~n8674 & n8832 ;
  assign n17143 = ( n13437 & n17141 ) | ( n13437 & n17142 ) | ( n17141 & n17142 ) ;
  assign n17144 = ~n901 & n4966 ;
  assign n17145 = n5538 & n17144 ;
  assign n17146 = n17145 ^ n15103 ^ 1'b0 ;
  assign n17147 = n2408 & ~n9161 ;
  assign n17148 = n17147 ^ n11283 ^ 1'b0 ;
  assign n17149 = n3371 & n9839 ;
  assign n17150 = n17149 ^ n12462 ^ 1'b0 ;
  assign n17151 = n16108 ^ n14044 ^ 1'b0 ;
  assign n17152 = n749 & ~n3876 ;
  assign n17153 = n17152 ^ n11479 ^ 1'b0 ;
  assign n17154 = n2078 | n3929 ;
  assign n17155 = n1246 ^ n75 ^ 1'b0 ;
  assign n17156 = n17154 & ~n17155 ;
  assign n17157 = ~n11095 & n17156 ;
  assign n17158 = n4270 ^ n1067 ^ 1'b0 ;
  assign n17159 = n8502 & ~n17158 ;
  assign n17160 = n4647 & ~n13203 ;
  assign n17161 = n17160 ^ n5484 ^ 1'b0 ;
  assign n17162 = n16057 ^ n3333 ^ 1'b0 ;
  assign n17163 = ~n677 & n17162 ;
  assign n17164 = n4770 ^ n4189 ^ 1'b0 ;
  assign n17165 = n15607 | n17164 ;
  assign n17166 = n1474 | n11288 ;
  assign n17167 = ~n3309 & n4029 ;
  assign n17168 = n5071 & n6700 ;
  assign n17169 = n17168 ^ n3653 ^ 1'b0 ;
  assign n17170 = n17169 ^ n3229 ^ 1'b0 ;
  assign n17171 = n6477 & ~n13887 ;
  assign n17176 = n1350 ^ n363 ^ 1'b0 ;
  assign n17177 = n3574 ^ n107 ^ 1'b0 ;
  assign n17178 = ~n17176 & n17177 ;
  assign n17174 = n2812 | n10255 ;
  assign n17173 = n3832 | n9476 ;
  assign n17175 = n17174 ^ n17173 ^ 1'b0 ;
  assign n17179 = n17178 ^ n17175 ^ 1'b0 ;
  assign n17180 = n4482 & n17179 ;
  assign n17172 = n2595 & ~n9184 ;
  assign n17181 = n17180 ^ n17172 ^ 1'b0 ;
  assign n17182 = n8075 & n17181 ;
  assign n17183 = n9641 ^ n390 ^ 1'b0 ;
  assign n17184 = n3969 ^ n3287 ^ 1'b0 ;
  assign n17185 = x0 | n17184 ;
  assign n17186 = n4088 | n7203 ;
  assign n17189 = n7104 ^ n3804 ^ 1'b0 ;
  assign n17190 = n375 | n17189 ;
  assign n17188 = n2501 | n3156 ;
  assign n17191 = n17190 ^ n17188 ^ 1'b0 ;
  assign n17187 = n7737 & ~n12902 ;
  assign n17192 = n17191 ^ n17187 ^ 1'b0 ;
  assign n17193 = n17192 ^ n4799 ^ 1'b0 ;
  assign n17194 = n11631 ^ n6476 ^ 1'b0 ;
  assign n17195 = n930 & n15093 ;
  assign n17196 = n17194 & n17195 ;
  assign n17197 = n13972 ^ n3037 ^ 1'b0 ;
  assign n17198 = n2612 & n17197 ;
  assign n17199 = n3359 & n17198 ;
  assign n17200 = n1891 & n17199 ;
  assign n17201 = n11933 & n17200 ;
  assign n17202 = n5903 & ~n12048 ;
  assign n17203 = n3665 & ~n9691 ;
  assign n17204 = n6125 & ~n13067 ;
  assign n17205 = ~n17203 & n17204 ;
  assign n17206 = ~n3303 & n5420 ;
  assign n17207 = n17206 ^ n4748 ^ 1'b0 ;
  assign n17208 = n17207 ^ n10858 ^ n8965 ;
  assign n17209 = n13416 | n17208 ;
  assign n17210 = n328 ^ n261 ^ 1'b0 ;
  assign n17212 = ~n19 & n1252 ;
  assign n17213 = ~n1252 & n17212 ;
  assign n17214 = ~n2023 & n17213 ;
  assign n17215 = n17214 ^ n3718 ^ 1'b0 ;
  assign n17211 = n11069 ^ n6109 ^ 1'b0 ;
  assign n17216 = n17215 ^ n17211 ^ 1'b0 ;
  assign n17217 = n1326 & ~n8013 ;
  assign n17218 = n17217 ^ n1396 ^ 1'b0 ;
  assign n17219 = n340 | n5996 ;
  assign n17220 = n810 | n17219 ;
  assign n17221 = n7856 | n15515 ;
  assign n17222 = n17221 ^ n16236 ^ 1'b0 ;
  assign n17223 = n12971 & n17222 ;
  assign n17224 = n427 & ~n5830 ;
  assign n17225 = n17224 ^ n6237 ^ 1'b0 ;
  assign n17226 = n4263 & ~n17225 ;
  assign n17227 = n4181 & n5776 ;
  assign n17228 = n5134 ^ n4649 ^ 1'b0 ;
  assign n17229 = n5942 ^ x11 ^ 1'b0 ;
  assign n17230 = n7975 & ~n17229 ;
  assign n17231 = n182 & n3242 ;
  assign n17232 = n17231 ^ n12892 ^ 1'b0 ;
  assign n17233 = n2909 & n17232 ;
  assign n17234 = n15983 ^ n1300 ^ 1'b0 ;
  assign n17235 = n4765 & ~n17234 ;
  assign n17236 = n929 & ~n3387 ;
  assign n17237 = n9531 | n17236 ;
  assign n17238 = n8864 & ~n17237 ;
  assign n17239 = n17235 & n17238 ;
  assign n17240 = n694 & ~n17239 ;
  assign n17241 = n17240 ^ n11355 ^ 1'b0 ;
  assign n17242 = n6458 ^ n2431 ^ 1'b0 ;
  assign n17243 = n1263 | n17242 ;
  assign n17244 = n1445 | n2714 ;
  assign n17245 = n763 & ~n17244 ;
  assign n17246 = n2681 & n2911 ;
  assign n17247 = n17246 ^ n414 ^ 1'b0 ;
  assign n17248 = n107 & n417 ;
  assign n17249 = n581 & ~n17248 ;
  assign n17250 = n1704 | n12479 ;
  assign n17251 = n17250 ^ n7824 ^ 1'b0 ;
  assign n17252 = n1537 & n17251 ;
  assign n17253 = n1080 & ~n17252 ;
  assign n17254 = ~n12381 & n17253 ;
  assign n17255 = n17254 ^ n1108 ^ 1'b0 ;
  assign n17256 = n8602 & ~n17255 ;
  assign n17257 = n1462 & ~n15279 ;
  assign n17258 = n17257 ^ n3032 ^ 1'b0 ;
  assign n17259 = ( n68 & ~n184 ) | ( n68 & n14080 ) | ( ~n184 & n14080 ) ;
  assign n17260 = n17259 ^ n8507 ^ 1'b0 ;
  assign n17261 = n1458 | n15201 ;
  assign n17262 = n4883 ^ n692 ^ 1'b0 ;
  assign n17263 = n5234 & n17262 ;
  assign n17264 = n10798 & n17263 ;
  assign n17265 = n2236 & n6627 ;
  assign n17266 = n10271 ^ n6706 ^ 1'b0 ;
  assign n17267 = n340 | n14618 ;
  assign n17268 = n311 | n17267 ;
  assign n17269 = n14470 ^ n8868 ^ 1'b0 ;
  assign n17275 = n343 | n15050 ;
  assign n17276 = n17275 ^ n2027 ^ 1'b0 ;
  assign n17270 = n2778 & ~n4737 ;
  assign n17271 = n1474 & n17270 ;
  assign n17272 = n6128 & n17271 ;
  assign n17273 = n7102 & ~n17272 ;
  assign n17274 = n17273 ^ n12274 ^ 1'b0 ;
  assign n17277 = n17276 ^ n17274 ^ 1'b0 ;
  assign n17278 = n6048 ^ n2495 ^ 1'b0 ;
  assign n17279 = n533 & ~n17278 ;
  assign n17280 = n16079 ^ n4750 ^ 1'b0 ;
  assign n17281 = n6739 & ~n17280 ;
  assign n17282 = n4116 ^ n121 ^ 1'b0 ;
  assign n17283 = n6873 & n17282 ;
  assign n17284 = n17281 | n17283 ;
  assign n17285 = n12657 ^ n2020 ^ n1600 ;
  assign n17286 = n7876 ^ n4090 ^ 1'b0 ;
  assign n17287 = n3761 & n4990 ;
  assign n17288 = n17287 ^ n2104 ^ 1'b0 ;
  assign n17289 = n5775 | n6277 ;
  assign n17290 = n17289 ^ n8973 ^ 1'b0 ;
  assign n17291 = n812 & ~n2509 ;
  assign n17292 = n7244 ^ n862 ^ 1'b0 ;
  assign n17293 = n17291 & n17292 ;
  assign n17294 = n40 & ~n1968 ;
  assign n17295 = n17294 ^ n6256 ^ 1'b0 ;
  assign n17296 = n4904 & ~n13087 ;
  assign n17297 = ~n3940 & n17296 ;
  assign n17298 = n15901 & ~n17297 ;
  assign n17299 = n17298 ^ n7319 ^ 1'b0 ;
  assign n17300 = n3208 & ~n4745 ;
  assign n17301 = n191 & n8639 ;
  assign n17302 = n13110 ^ n8530 ^ 1'b0 ;
  assign n17303 = n9275 & n12279 ;
  assign n17304 = n17303 ^ n4899 ^ 1'b0 ;
  assign n17305 = n12706 & ~n17304 ;
  assign n17306 = ( n8986 & n10366 ) | ( n8986 & n11924 ) | ( n10366 & n11924 ) ;
  assign n17307 = n495 & ~n11119 ;
  assign n17308 = n17307 ^ n1933 ^ 1'b0 ;
  assign n17309 = ~n4606 & n10636 ;
  assign n17310 = n17309 ^ n1961 ^ 1'b0 ;
  assign n17311 = ~n13114 & n17310 ;
  assign n17312 = n10025 & n17311 ;
  assign n17313 = n17312 ^ n4084 ^ 1'b0 ;
  assign n17315 = n4273 & ~n5737 ;
  assign n17314 = ~n153 & n2939 ;
  assign n17316 = n17315 ^ n17314 ^ 1'b0 ;
  assign n17317 = n2138 | n8116 ;
  assign n17318 = n2619 & ~n15194 ;
  assign n17319 = n17318 ^ n6188 ^ 1'b0 ;
  assign n17321 = n144 | n614 ;
  assign n17322 = n13330 & n17321 ;
  assign n17323 = n17322 ^ n4075 ^ 1'b0 ;
  assign n17320 = ~n6849 & n9583 ;
  assign n17324 = n17323 ^ n17320 ^ 1'b0 ;
  assign n17325 = ~n5812 & n17324 ;
  assign n17326 = n2679 & ~n5343 ;
  assign n17327 = n9832 & n17326 ;
  assign n17328 = n2495 & n17327 ;
  assign n17329 = n271 & n5818 ;
  assign n17330 = n4983 & n8405 ;
  assign n17331 = n2908 | n17330 ;
  assign n17332 = n17330 & ~n17331 ;
  assign n17333 = n13670 | n17332 ;
  assign n17334 = n7241 & ~n17333 ;
  assign n17335 = ~n11585 & n15806 ;
  assign n17336 = ~n15293 & n17335 ;
  assign n17341 = n2486 ^ n159 ^ 1'b0 ;
  assign n17337 = n4550 | n10557 ;
  assign n17338 = ~n286 & n4328 ;
  assign n17339 = n17338 ^ n5530 ^ 1'b0 ;
  assign n17340 = n17337 | n17339 ;
  assign n17342 = n17341 ^ n17340 ^ 1'b0 ;
  assign n17343 = n1873 & n17342 ;
  assign n17344 = n17343 ^ n15695 ^ 1'b0 ;
  assign n17345 = n17336 | n17344 ;
  assign n17346 = n17345 ^ n14662 ^ 1'b0 ;
  assign n17347 = n5452 & ~n12658 ;
  assign n17348 = n11155 & n17347 ;
  assign n17349 = n338 & n1308 ;
  assign n17350 = n17349 ^ n3424 ^ 1'b0 ;
  assign n17351 = n17350 ^ n10761 ^ 1'b0 ;
  assign n17352 = n5721 & n5771 ;
  assign n17353 = ~n5096 & n17352 ;
  assign n17354 = ~n310 & n9372 ;
  assign n17355 = n16346 | n17354 ;
  assign n17356 = n8172 & ~n17355 ;
  assign n17357 = n3074 & ~n4996 ;
  assign n17358 = n17357 ^ n810 ^ 1'b0 ;
  assign n17359 = ~n2458 & n2942 ;
  assign n17360 = ~n8014 & n17359 ;
  assign n17361 = n715 & ~n7245 ;
  assign n17362 = ~n11707 & n17361 ;
  assign n17363 = n6160 & n17362 ;
  assign n17364 = n4574 ^ n250 ^ 1'b0 ;
  assign n17365 = ~n15434 & n17364 ;
  assign n17366 = n10797 & n11124 ;
  assign n17369 = n14694 ^ n5729 ^ n279 ;
  assign n17367 = ~n7439 & n9914 ;
  assign n17368 = ~n7367 & n17367 ;
  assign n17370 = n17369 ^ n17368 ^ 1'b0 ;
  assign n17371 = n4432 | n16445 ;
  assign n17372 = n3693 ^ n2012 ^ 1'b0 ;
  assign n17373 = n2155 | n7236 ;
  assign n17374 = n17373 ^ n5996 ^ 1'b0 ;
  assign n17375 = n10664 ^ n9422 ^ 1'b0 ;
  assign n17376 = ~n1619 & n17375 ;
  assign n17377 = n2200 & n2700 ;
  assign n17378 = ~n2700 & n17377 ;
  assign n17379 = n17378 ^ n11931 ^ 1'b0 ;
  assign n17380 = n17376 & ~n17379 ;
  assign n17381 = n17374 & n17380 ;
  assign n17382 = n86 ^ n55 ^ 1'b0 ;
  assign n17383 = n8639 | n17382 ;
  assign n17384 = n1966 | n17383 ;
  assign n17385 = n17384 ^ n11379 ^ 1'b0 ;
  assign n17386 = n11863 & n17385 ;
  assign n17387 = n10178 ^ n243 ^ 1'b0 ;
  assign n17388 = ~n7669 & n17387 ;
  assign n17389 = n2156 | n5005 ;
  assign n17390 = n5761 ^ n2949 ^ n1622 ;
  assign n17391 = n17390 ^ n6464 ^ 1'b0 ;
  assign n17392 = ~n8414 & n17391 ;
  assign n17393 = n6602 & n13297 ;
  assign n17394 = n7933 & n17393 ;
  assign n17395 = ~n4660 & n6159 ;
  assign n17396 = n15067 ^ n1113 ^ 1'b0 ;
  assign n17397 = n1469 | n12242 ;
  assign n17398 = n17396 | n17397 ;
  assign n17403 = n43 & n12587 ;
  assign n17404 = ~n36 & n17403 ;
  assign n17405 = n690 | n1573 ;
  assign n17406 = n1573 & ~n17405 ;
  assign n17407 = ~n381 & n15727 ;
  assign n17408 = ~n243 & n249 ;
  assign n17409 = n243 & n17408 ;
  assign n17410 = n17407 & ~n17409 ;
  assign n17411 = n17406 & n17410 ;
  assign n17412 = ~n12831 & n17411 ;
  assign n17413 = n2397 & ~n17412 ;
  assign n17414 = ~n2397 & n17413 ;
  assign n17415 = n81 & n170 ;
  assign n17416 = ~n170 & n17415 ;
  assign n17417 = n17416 ^ n83 ^ 1'b0 ;
  assign n17418 = n21 & n40 ;
  assign n17419 = ~n40 & n17418 ;
  assign n17420 = n88 & ~n17419 ;
  assign n17421 = ~n88 & n17420 ;
  assign n17422 = n1173 & n17421 ;
  assign n17423 = n178 & n17422 ;
  assign n17424 = n17417 & n17423 ;
  assign n17425 = n1315 & n17424 ;
  assign n17426 = n17414 | n17425 ;
  assign n17427 = n17404 & ~n17426 ;
  assign n17399 = n338 & n1381 ;
  assign n17400 = ~n338 & n17399 ;
  assign n17401 = n107 & n17400 ;
  assign n17402 = n15066 | n17401 ;
  assign n17428 = n17427 ^ n17402 ^ 1'b0 ;
  assign n17429 = ~n6797 & n12205 ;
  assign n17430 = n17429 ^ n8602 ^ 1'b0 ;
  assign n17431 = ~n17428 & n17430 ;
  assign n17432 = n15781 ^ n11982 ^ 1'b0 ;
  assign n17435 = n227 & ~n11566 ;
  assign n17436 = n17435 ^ n363 ^ 1'b0 ;
  assign n17434 = n3845 & n12562 ;
  assign n17437 = n17436 ^ n17434 ^ 1'b0 ;
  assign n17433 = n8283 | n9697 ;
  assign n17438 = n17437 ^ n17433 ^ 1'b0 ;
  assign n17439 = n310 | n6266 ;
  assign n17440 = ~x8 & n17439 ;
  assign n17441 = n1246 & n17440 ;
  assign n17442 = n10963 ^ n1309 ^ 1'b0 ;
  assign n17443 = n892 & n17442 ;
  assign n17444 = ~n3576 & n17443 ;
  assign n17445 = ~n3010 & n7126 ;
  assign n17446 = n542 & n7120 ;
  assign n17447 = n17446 ^ n11735 ^ 1'b0 ;
  assign n17448 = n2136 & n9325 ;
  assign n17449 = n747 | n17448 ;
  assign n17450 = n9534 ^ n2302 ^ 1'b0 ;
  assign n17451 = n6817 & ~n17450 ;
  assign n17452 = ~n14976 & n17451 ;
  assign n17459 = n8860 ^ n3263 ^ 1'b0 ;
  assign n17460 = n616 | n17459 ;
  assign n17453 = n270 | n551 ;
  assign n17454 = n270 & ~n17453 ;
  assign n17455 = ~n119 & n178 ;
  assign n17456 = n17454 & n17455 ;
  assign n17457 = n4840 & n12002 ;
  assign n17458 = n17456 | n17457 ;
  assign n17461 = n17460 ^ n17458 ^ 1'b0 ;
  assign n17462 = n7821 ^ n4432 ^ 1'b0 ;
  assign n17463 = n861 | n5067 ;
  assign n17464 = n258 & ~n17463 ;
  assign n17465 = n10377 ^ n7195 ^ 1'b0 ;
  assign n17466 = n5995 & ~n8290 ;
  assign n17467 = n3874 & n17466 ;
  assign n17468 = n17467 ^ n14182 ^ 1'b0 ;
  assign n17469 = n7988 ^ n4917 ^ 1'b0 ;
  assign n17470 = n13579 ^ n227 ^ 1'b0 ;
  assign n17471 = n3533 | n17470 ;
  assign n17472 = n17471 ^ n3206 ^ 1'b0 ;
  assign n17473 = n1081 & n17472 ;
  assign n17474 = n17473 ^ n6468 ^ 1'b0 ;
  assign n17475 = n1309 | n16653 ;
  assign n17476 = n2059 & n10567 ;
  assign n17477 = n17476 ^ n8862 ^ 1'b0 ;
  assign n17478 = ~n17317 & n17477 ;
  assign n17479 = x6 & n2467 ;
  assign n17480 = n223 & n2159 ;
  assign n17481 = n17479 & n17480 ;
  assign n17482 = n14539 ^ n2450 ^ 1'b0 ;
  assign n17483 = n5313 ^ n183 ^ 1'b0 ;
  assign n17484 = n17483 ^ n1877 ^ 1'b0 ;
  assign n17485 = n7747 & n11972 ;
  assign n17486 = n698 & n17485 ;
  assign n17487 = ( n1467 & ~n7459 ) | ( n1467 & n10275 ) | ( ~n7459 & n10275 ) ;
  assign n17488 = n11618 ^ n8598 ^ 1'b0 ;
  assign n17489 = n2661 | n12749 ;
  assign n17490 = n15117 & ~n17489 ;
  assign n17491 = n567 | n13892 ;
  assign n17492 = n17491 ^ n10360 ^ 1'b0 ;
  assign n17493 = n456 & ~n17492 ;
  assign n17494 = n6730 | n9036 ;
  assign n17495 = n5255 & ~n17494 ;
  assign n17497 = n3940 | n6230 ;
  assign n17496 = n46 & n11525 ;
  assign n17498 = n17497 ^ n17496 ^ 1'b0 ;
  assign n17499 = ~n2747 & n2828 ;
  assign n17500 = n17499 ^ n14544 ^ 1'b0 ;
  assign n17501 = n17500 ^ n11696 ^ 1'b0 ;
  assign n17502 = n7392 & n17501 ;
  assign n17503 = n17502 ^ n10658 ^ 1'b0 ;
  assign n17504 = ~n8921 & n17503 ;
  assign n17505 = n461 & ~n1095 ;
  assign n17506 = n17505 ^ n1759 ^ 1'b0 ;
  assign n17507 = n5237 | n11678 ;
  assign n17508 = n8523 & n17507 ;
  assign n17509 = ~n7419 & n17508 ;
  assign n17510 = n1224 & ~n2844 ;
  assign n17511 = n2844 & n17510 ;
  assign n17512 = n15867 | n17511 ;
  assign n17513 = n14213 & ~n17512 ;
  assign n17514 = ~n14213 & n17513 ;
  assign n17515 = n6636 | n12422 ;
  assign n17516 = n17515 ^ x5 ^ 1'b0 ;
  assign n17517 = ~n2872 & n6443 ;
  assign n17521 = n11645 ^ n9410 ^ 1'b0 ;
  assign n17522 = n11820 & ~n17521 ;
  assign n17523 = n17522 ^ n10627 ^ n10345 ;
  assign n17518 = n5796 & n5799 ;
  assign n17519 = n4823 & n17518 ;
  assign n17520 = n14759 & ~n17519 ;
  assign n17524 = n17523 ^ n17520 ^ 1'b0 ;
  assign n17525 = n4081 ^ n975 ^ 1'b0 ;
  assign n17526 = n17525 ^ n1008 ^ 1'b0 ;
  assign n17527 = n17526 ^ n12457 ^ 1'b0 ;
  assign n17528 = n11806 | n17527 ;
  assign n17529 = n957 & ~n3162 ;
  assign n17530 = ~n3627 & n17529 ;
  assign n17531 = n1386 ^ n277 ^ 1'b0 ;
  assign n17532 = n17531 ^ n6919 ^ 1'b0 ;
  assign n17533 = n3579 & n17532 ;
  assign n17534 = n4406 | n13068 ;
  assign n17537 = n327 & n1491 ;
  assign n17535 = n942 & n11057 ;
  assign n17536 = ~n8261 & n17535 ;
  assign n17538 = n17537 ^ n17536 ^ 1'b0 ;
  assign n17539 = n1143 & ~n7388 ;
  assign n17540 = n17539 ^ n8756 ^ 1'b0 ;
  assign n17541 = n5396 & n17540 ;
  assign n17544 = ~n963 & n7120 ;
  assign n17545 = n17544 ^ n4488 ^ 1'b0 ;
  assign n17546 = ~n9739 & n17545 ;
  assign n17542 = n1130 & n12167 ;
  assign n17543 = n8234 & ~n17542 ;
  assign n17547 = n17546 ^ n17543 ^ 1'b0 ;
  assign n17548 = ~n4031 & n12488 ;
  assign n17549 = n14323 & ~n17341 ;
  assign n17550 = n1901 | n14863 ;
  assign n17551 = ( n882 & n7995 ) | ( n882 & n11360 ) | ( n7995 & n11360 ) ;
  assign n17552 = n4037 | n9240 ;
  assign n17553 = n17552 ^ n10878 ^ 1'b0 ;
  assign n17554 = n86 & n6960 ;
  assign n17555 = n1775 & n17554 ;
  assign n17556 = n17555 ^ n17007 ^ 1'b0 ;
  assign n17557 = ( ~n4819 & n8823 ) | ( ~n4819 & n17556 ) | ( n8823 & n17556 ) ;
  assign n17558 = n495 & n7261 ;
  assign n17559 = n7503 ^ n727 ^ 1'b0 ;
  assign n17560 = n148 & ~n17559 ;
  assign n17561 = n17560 ^ n777 ^ 1'b0 ;
  assign n17562 = n2012 ^ n384 ^ 1'b0 ;
  assign n17563 = ~n418 & n17562 ;
  assign n17564 = n395 & n17563 ;
  assign n17565 = n1347 & ~n10374 ;
  assign n17566 = n1060 & ~n2902 ;
  assign n17567 = ~n5102 & n17566 ;
  assign n17568 = n2948 & n11088 ;
  assign n17569 = n928 & n3166 ;
  assign n17570 = n17569 ^ n8333 ^ n1726 ;
  assign n17571 = ~n14734 & n17570 ;
  assign n17572 = n1733 & ~n7866 ;
  assign n17573 = n17572 ^ n16509 ^ 1'b0 ;
  assign n17574 = ( n3301 & n8505 ) | ( n3301 & ~n9655 ) | ( n8505 & ~n9655 ) ;
  assign n17575 = ~n131 & n299 ;
  assign n17576 = n131 & n17575 ;
  assign n17577 = n142 & ~n17576 ;
  assign n17578 = n7552 & n17577 ;
  assign n17579 = ~n17577 & n17578 ;
  assign n17580 = n622 & ~n8181 ;
  assign n17581 = n7237 & n17580 ;
  assign n17582 = n7338 | n17581 ;
  assign n17583 = n17582 ^ n16643 ^ 1'b0 ;
  assign n17584 = n17583 ^ n9199 ^ n1910 ;
  assign n17585 = n11641 ^ n8197 ^ 1'b0 ;
  assign n17586 = n9245 & ~n17585 ;
  assign n17587 = ~n216 & n14143 ;
  assign n17588 = n17587 ^ n6322 ^ 1'b0 ;
  assign n17589 = ~n1283 & n13007 ;
  assign n17590 = n6834 | n13870 ;
  assign n17591 = n2163 | n17590 ;
  assign n17592 = n6647 ^ n2422 ^ 1'b0 ;
  assign n17593 = n8370 & n9541 ;
  assign n17594 = n1672 & n17593 ;
  assign n17595 = n340 & ~n17594 ;
  assign n17596 = n3598 & n17595 ;
  assign n17597 = ~n8333 & n15631 ;
  assign n17598 = n17597 ^ n6226 ^ 1'b0 ;
  assign n17599 = n13391 ^ n7853 ^ 1'b0 ;
  assign n17600 = ~n9039 & n12760 ;
  assign n17601 = n3267 & n5811 ;
  assign n17602 = n2515 & ~n6562 ;
  assign n17603 = ~n7001 & n17602 ;
  assign n17604 = n14185 & ~n17603 ;
  assign n17605 = n17604 ^ n9884 ^ 1'b0 ;
  assign n17606 = n5084 ^ n3121 ^ 1'b0 ;
  assign n17607 = n1479 & n17606 ;
  assign n17608 = n13572 & ~n17607 ;
  assign n17609 = n1652 ^ n690 ^ 1'b0 ;
  assign n17610 = n129 & n17609 ;
  assign n17611 = n12980 & ~n15194 ;
  assign n17612 = n17611 ^ n2982 ^ 1'b0 ;
  assign n17613 = ~n1806 & n4406 ;
  assign n17614 = n12889 | n16246 ;
  assign n17615 = n55 & ~n17614 ;
  assign n17616 = n16572 ^ n10996 ^ 1'b0 ;
  assign n17617 = n17616 ^ n12362 ^ 1'b0 ;
  assign n17618 = n3927 ^ n1564 ^ 1'b0 ;
  assign n17619 = n11178 ^ n8426 ^ 1'b0 ;
  assign n17620 = n17618 | n17619 ;
  assign n17621 = n677 & ~n9060 ;
  assign n17622 = n618 & ~n7845 ;
  assign n17623 = ~n4540 & n17622 ;
  assign n17624 = n17623 ^ n5359 ^ 1'b0 ;
  assign n17625 = n10002 & n16566 ;
  assign n17626 = ~n6742 & n9501 ;
  assign n17627 = n17626 ^ n4460 ^ 1'b0 ;
  assign n17628 = n17627 ^ n12046 ^ 1'b0 ;
  assign n17630 = n1748 ^ n86 ^ 1'b0 ;
  assign n17629 = n255 | n1348 ;
  assign n17631 = n17630 ^ n17629 ^ 1'b0 ;
  assign n17632 = n7409 & ~n17631 ;
  assign n17633 = n17632 ^ n9225 ^ 1'b0 ;
  assign n17634 = n14210 & ~n17633 ;
  assign n17635 = n2687 & ~n3803 ;
  assign n17636 = n17635 ^ n15723 ^ 1'b0 ;
  assign n17637 = ~n1790 & n2879 ;
  assign n17638 = n7471 | n17637 ;
  assign n17639 = ~n1186 & n7599 ;
  assign n17640 = n1779 & ~n9751 ;
  assign n17641 = n5884 ^ n5758 ^ 1'b0 ;
  assign n17642 = ~n5084 & n17641 ;
  assign n17643 = n1699 ^ n1556 ^ 1'b0 ;
  assign n17649 = n4547 ^ n4381 ^ 1'b0 ;
  assign n17644 = n180 | n5310 ;
  assign n17645 = n159 & ~n17644 ;
  assign n17646 = n9233 | n17645 ;
  assign n17647 = n17646 ^ n12725 ^ 1'b0 ;
  assign n17648 = ~n8916 & n17647 ;
  assign n17650 = n17649 ^ n17648 ^ 1'b0 ;
  assign n17651 = n6539 ^ n4517 ^ 1'b0 ;
  assign n17652 = n4820 & ~n10084 ;
  assign n17653 = n3920 & n11367 ;
  assign n17654 = n3346 ^ n627 ^ 1'b0 ;
  assign n17655 = n5232 & ~n17654 ;
  assign n17656 = n9428 ^ n5255 ^ 1'b0 ;
  assign n17657 = n17656 ^ n6887 ^ 1'b0 ;
  assign n17658 = n2873 & ~n5444 ;
  assign n17659 = n5444 & n17658 ;
  assign n17660 = ~n1026 & n8056 ;
  assign n17661 = ~n8056 & n17660 ;
  assign n17662 = n7464 & ~n17661 ;
  assign n17663 = n17661 & n17662 ;
  assign n17664 = n17663 ^ n489 ^ 1'b0 ;
  assign n17665 = n17659 | n17664 ;
  assign n17667 = n3969 ^ n3721 ^ 1'b0 ;
  assign n17668 = n17667 ^ n5872 ^ 1'b0 ;
  assign n17666 = n4890 & n10816 ;
  assign n17669 = n17668 ^ n17666 ^ 1'b0 ;
  assign n17670 = n2784 ^ n1673 ^ 1'b0 ;
  assign n17671 = n5083 ^ n1506 ^ 1'b0 ;
  assign n17672 = n10990 ^ n2377 ^ 1'b0 ;
  assign n17673 = ~n3481 & n17672 ;
  assign n17674 = ~n12656 & n17673 ;
  assign n17675 = n1286 | n8382 ;
  assign n17676 = n7140 & n12890 ;
  assign n17677 = ~n3748 & n17676 ;
  assign n17678 = n17677 ^ n1785 ^ 1'b0 ;
  assign n17679 = n295 ^ n16 ^ 1'b0 ;
  assign n17680 = n6849 & n17679 ;
  assign n17681 = ~n1115 & n9693 ;
  assign n17682 = n9172 & n17681 ;
  assign n17683 = n14772 ^ n5347 ^ n2117 ;
  assign n17685 = n7221 & ~n7726 ;
  assign n17684 = n9582 ^ n5547 ^ 1'b0 ;
  assign n17686 = n17685 ^ n17684 ^ 1'b0 ;
  assign n17687 = ~n17683 & n17686 ;
  assign n17688 = n12628 ^ n736 ^ 1'b0 ;
  assign n17689 = ~n16296 & n17197 ;
  assign n17690 = n1940 & n17689 ;
  assign n17691 = n7439 & n17690 ;
  assign n17692 = n2738 | n13237 ;
  assign n17694 = n1655 ^ n1652 ^ 1'b0 ;
  assign n17693 = ~n5217 & n11382 ;
  assign n17695 = n17694 ^ n17693 ^ 1'b0 ;
  assign n17699 = n1130 & n4042 ;
  assign n17700 = ~n2825 & n17699 ;
  assign n17696 = x6 & ~n5060 ;
  assign n17697 = ~n5959 & n17696 ;
  assign n17698 = n17044 | n17697 ;
  assign n17701 = n17700 ^ n17698 ^ 1'b0 ;
  assign n17702 = n11735 | n12021 ;
  assign n17703 = ~n5853 & n6762 ;
  assign n17704 = ~n13168 & n15831 ;
  assign n17708 = n254 ^ n177 ^ 1'b0 ;
  assign n17709 = n2261 & ~n17708 ;
  assign n17710 = n17709 ^ n14324 ^ 1'b0 ;
  assign n17705 = n1743 & n10213 ;
  assign n17706 = n14185 & ~n17705 ;
  assign n17707 = n17706 ^ n3511 ^ 1'b0 ;
  assign n17711 = n17710 ^ n17707 ^ 1'b0 ;
  assign n17712 = n12895 ^ n3653 ^ 1'b0 ;
  assign n17713 = n3135 & ~n17712 ;
  assign n17714 = n2017 & n4595 ;
  assign n17715 = n8957 & n15718 ;
  assign n17716 = ~n17714 & n17715 ;
  assign n17717 = n16663 & ~n17716 ;
  assign n17718 = n185 & ~n1898 ;
  assign n17719 = n17718 ^ n2460 ^ 1'b0 ;
  assign n17723 = ~n3193 & n4311 ;
  assign n17724 = n17723 ^ n1036 ^ 1'b0 ;
  assign n17725 = n5809 & n17724 ;
  assign n17720 = n4662 & n7120 ;
  assign n17721 = n4618 & n17720 ;
  assign n17722 = n10475 & ~n17721 ;
  assign n17726 = n17725 ^ n17722 ^ 1'b0 ;
  assign n17727 = n17726 ^ n2964 ^ 1'b0 ;
  assign n17728 = n17719 & ~n17727 ;
  assign n17732 = n3097 & ~n6755 ;
  assign n17733 = n17732 ^ n5776 ^ 1'b0 ;
  assign n17729 = n3180 | n7501 ;
  assign n17730 = n17729 ^ n628 ^ 1'b0 ;
  assign n17731 = n5867 & n17730 ;
  assign n17734 = n17733 ^ n17731 ^ n16835 ;
  assign n17735 = n708 | n2157 ;
  assign n17736 = n17735 ^ n616 ^ 1'b0 ;
  assign n17737 = ~n5481 & n8858 ;
  assign n17738 = ~n1523 & n17737 ;
  assign n17739 = ( ~n12325 & n12954 ) | ( ~n12325 & n17738 ) | ( n12954 & n17738 ) ;
  assign n17740 = ~n461 & n17739 ;
  assign n17741 = n1202 | n1396 ;
  assign n17742 = n17740 & ~n17741 ;
  assign n17743 = n2574 | n8437 ;
  assign n17744 = n195 & ~n17743 ;
  assign n17745 = n9132 ^ n2316 ^ 1'b0 ;
  assign n17746 = ~n11245 & n17745 ;
  assign n17747 = ~n5831 & n5884 ;
  assign n17748 = n640 & n17747 ;
  assign n17753 = n4961 | n4998 ;
  assign n17749 = n98 | n5055 ;
  assign n17750 = n4025 & n17749 ;
  assign n17751 = n17750 ^ n6125 ^ 1'b0 ;
  assign n17752 = n340 & n17751 ;
  assign n17754 = n17753 ^ n17752 ^ 1'b0 ;
  assign n17755 = n5161 ^ n313 ^ 1'b0 ;
  assign n17756 = ( n3007 & n5025 ) | ( n3007 & n17755 ) | ( n5025 & n17755 ) ;
  assign n17757 = n17756 ^ n13949 ^ 1'b0 ;
  assign n17758 = n11645 | n17757 ;
  assign n17759 = n5059 & n15943 ;
  assign n17760 = n13275 ^ n8825 ^ 1'b0 ;
  assign n17761 = n10059 ^ n7355 ^ 1'b0 ;
  assign n17762 = n6055 ^ n3179 ^ 1'b0 ;
  assign n17763 = n1790 | n5588 ;
  assign n17764 = n17763 ^ n1227 ^ 1'b0 ;
  assign n17765 = n3017 ^ n2155 ^ 1'b0 ;
  assign n17766 = n4694 & n13983 ;
  assign n17769 = n8745 & ~n14611 ;
  assign n17770 = n17769 ^ n7934 ^ 1'b0 ;
  assign n17767 = n14425 ^ n3498 ^ 1'b0 ;
  assign n17768 = n5267 | n17767 ;
  assign n17771 = n17770 ^ n17768 ^ 1'b0 ;
  assign n17772 = n1429 & n7659 ;
  assign n17773 = n442 | n1044 ;
  assign n17774 = n17773 ^ n83 ^ 1'b0 ;
  assign n17775 = n105 & n17774 ;
  assign n17776 = n17775 ^ n779 ^ 1'b0 ;
  assign n17777 = n17776 ^ n1149 ^ 1'b0 ;
  assign n17778 = n4815 | n17777 ;
  assign n17779 = n17778 ^ n11020 ^ 1'b0 ;
  assign n17780 = n17637 & n17669 ;
  assign n17781 = n17233 ^ n863 ^ 1'b0 ;
  assign n17782 = n11593 & ~n12386 ;
  assign n17783 = ~n16209 & n17782 ;
  assign n17784 = ~n42 & n7917 ;
  assign n17785 = ~n7199 & n17784 ;
  assign n17786 = n17785 ^ n8597 ^ 1'b0 ;
  assign n17787 = ~n12477 & n17786 ;
  assign n17788 = ~n3156 & n17787 ;
  assign n17789 = ~n624 & n17788 ;
  assign n17790 = n17783 & ~n17789 ;
  assign n17791 = n17479 ^ n13961 ^ 1'b0 ;
  assign n17792 = n798 & n7980 ;
  assign n17793 = ~n2246 & n17792 ;
  assign n17794 = ( n16639 & ~n17791 ) | ( n16639 & n17793 ) | ( ~n17791 & n17793 ) ;
  assign n17795 = n4460 ^ n2032 ^ 1'b0 ;
  assign n17796 = n17795 ^ n7734 ^ 1'b0 ;
  assign n17799 = n4098 ^ n781 ^ 1'b0 ;
  assign n17797 = n2542 & n5623 ;
  assign n17798 = n17797 ^ n2932 ^ 1'b0 ;
  assign n17800 = n17799 ^ n17798 ^ n300 ;
  assign n17801 = ~n6636 & n11787 ;
  assign n17802 = n17801 ^ n6512 ^ 1'b0 ;
  assign n17803 = n5080 & n8014 ;
  assign n17804 = n15532 & n17803 ;
  assign n17805 = n4231 & ~n10067 ;
  assign n17806 = ~n627 & n17805 ;
  assign n17807 = ~n2912 & n9897 ;
  assign n17808 = ~n4241 & n16971 ;
  assign n17809 = ~n530 & n17808 ;
  assign n17810 = n9376 & ~n15144 ;
  assign n17811 = ~n5467 & n17810 ;
  assign n17812 = n16897 | n17811 ;
  assign n17813 = n3959 ^ n3894 ^ 1'b0 ;
  assign n17815 = n3796 & ~n5468 ;
  assign n17814 = n6608 & n12877 ;
  assign n17816 = n17815 ^ n17814 ^ 1'b0 ;
  assign n17817 = ~n14224 & n17717 ;
  assign n17818 = n963 | n2681 ;
  assign n17819 = n1533 & ~n5394 ;
  assign n17820 = n17819 ^ n1143 ^ 1'b0 ;
  assign n17821 = n17820 ^ n12980 ^ n3437 ;
  assign n17822 = n4274 | n7599 ;
  assign n17823 = ~n273 & n804 ;
  assign n17824 = n17823 ^ n8072 ^ 1'b0 ;
  assign n17825 = ~n17822 & n17824 ;
  assign n17826 = n2120 & n17825 ;
  assign n17827 = n17826 ^ n3088 ^ 1'b0 ;
  assign n17828 = n10853 ^ n294 ^ 1'b0 ;
  assign n17829 = n11857 | n17828 ;
  assign n17830 = n17829 ^ n6476 ^ 1'b0 ;
  assign n17831 = n4120 | n14537 ;
  assign n17832 = n4516 & ~n17831 ;
  assign n17833 = ~n17830 & n17832 ;
  assign n17834 = n2721 ^ n713 ^ 1'b0 ;
  assign n17835 = n556 | n17834 ;
  assign n17836 = n11253 ^ n9792 ^ n5025 ;
  assign n17837 = n16276 & n17836 ;
  assign n17838 = n4625 ^ n536 ^ 1'b0 ;
  assign n17839 = n13437 ^ n7368 ^ 1'b0 ;
  assign n17840 = n8726 & n8867 ;
  assign n17841 = n6266 & n17840 ;
  assign n17842 = n4510 & n10215 ;
  assign n17843 = n12320 & n17842 ;
  assign n17844 = n5393 & ~n17843 ;
  assign n17845 = n3369 | n4136 ;
  assign n17846 = n17845 ^ n7425 ^ 1'b0 ;
  assign n17847 = n2426 ^ n891 ^ 1'b0 ;
  assign n17848 = ~n465 & n17847 ;
  assign n17849 = n1743 | n17848 ;
  assign n17850 = n5895 & ~n17849 ;
  assign n17851 = n17850 ^ n3803 ^ 1'b0 ;
  assign n17852 = n11037 & ~n17851 ;
  assign n17853 = ~n2065 & n17852 ;
  assign n17854 = n1541 & n7109 ;
  assign n17855 = n4491 | n17125 ;
  assign n17856 = n14432 & ~n17855 ;
  assign n17857 = n10789 ^ n6136 ^ 1'b0 ;
  assign n17858 = n3684 ^ n622 ^ 1'b0 ;
  assign n17859 = n5437 | n17858 ;
  assign n17860 = n6908 ^ n1547 ^ 1'b0 ;
  assign n17861 = n17860 ^ n5419 ^ 1'b0 ;
  assign n17862 = n17861 ^ n5559 ^ n4509 ;
  assign n17863 = n4180 & n17862 ;
  assign n17864 = n17863 ^ n11434 ^ 1'b0 ;
  assign n17865 = n193 & n11382 ;
  assign n17866 = n37 & n17865 ;
  assign n17867 = ( n37 & n1300 ) | ( n37 & n13930 ) | ( n1300 & n13930 ) ;
  assign n17868 = n3344 ^ n616 ^ 1'b0 ;
  assign n17869 = n4140 & n4585 ;
  assign n17870 = n5979 & n17869 ;
  assign n17871 = n16548 & n17870 ;
  assign n17872 = n812 & n1826 ;
  assign n17873 = n628 & n11421 ;
  assign n17874 = ~n17872 & n17873 ;
  assign n17875 = ~n17871 & n17874 ;
  assign n17876 = n2049 | n2784 ;
  assign n17877 = n17876 ^ n8630 ^ 1'b0 ;
  assign n17878 = ~n4379 & n16225 ;
  assign n17879 = n17878 ^ n17667 ^ 1'b0 ;
  assign n17880 = n1226 & n1543 ;
  assign n17881 = ~n17879 & n17880 ;
  assign n17882 = n3589 | n9792 ;
  assign n17883 = n12210 | n17882 ;
  assign n17884 = n17883 ^ n9292 ^ 1'b0 ;
  assign n17885 = n10682 | n11234 ;
  assign n17886 = n14272 ^ n12723 ^ n6515 ;
  assign n17887 = n241 & n17886 ;
  assign n17888 = n9344 ^ n7870 ^ n432 ;
  assign n17889 = n850 | n17888 ;
  assign n17890 = n15674 & n17889 ;
  assign n17891 = ( n820 & n2577 ) | ( n820 & n7905 ) | ( n2577 & n7905 ) ;
  assign n17892 = n6602 & ~n17891 ;
  assign n17893 = n7744 & n17892 ;
  assign n17894 = n2535 & n17893 ;
  assign n17895 = n17894 ^ n2869 ^ 1'b0 ;
  assign n17896 = ~n1158 & n14404 ;
  assign n17897 = ~n1060 & n5752 ;
  assign n17898 = n17236 ^ n6695 ^ 1'b0 ;
  assign n17899 = n3646 | n17898 ;
  assign n17900 = n14372 ^ n977 ^ 1'b0 ;
  assign n17901 = n1571 | n7424 ;
  assign n17902 = n5061 ^ n1748 ^ 1'b0 ;
  assign n17903 = n290 | n17902 ;
  assign n17904 = n2313 | n7607 ;
  assign n17905 = n8684 & ~n17904 ;
  assign n17906 = n17903 | n17905 ;
  assign n17907 = n13584 | n17906 ;
  assign n17910 = n1106 & ~n10634 ;
  assign n17908 = n980 & n1836 ;
  assign n17909 = n17908 ^ n1582 ^ 1'b0 ;
  assign n17911 = n17910 ^ n17909 ^ 1'b0 ;
  assign n17912 = n14747 ^ n643 ^ 1'b0 ;
  assign n17913 = ( n25 & ~n5180 ) | ( n25 & n8115 ) | ( ~n5180 & n8115 ) ;
  assign n17914 = ( n956 & n5335 ) | ( n956 & ~n5343 ) | ( n5335 & ~n5343 ) ;
  assign n17915 = ~n7731 & n17914 ;
  assign n17916 = n17915 ^ n2779 ^ 1'b0 ;
  assign n17917 = n17916 ^ n16814 ^ 1'b0 ;
  assign n17918 = ~n17913 & n17917 ;
  assign n17919 = n7780 ^ n2320 ^ 1'b0 ;
  assign n17920 = n47 & n17919 ;
  assign n17921 = n17920 ^ n4916 ^ 1'b0 ;
  assign n17922 = n133 | n1790 ;
  assign n17923 = n17921 & ~n17922 ;
  assign n17924 = n7328 & ~n14274 ;
  assign n17925 = n17924 ^ n12934 ^ 1'b0 ;
  assign n17926 = ~n17923 & n17925 ;
  assign n17927 = n2435 & n13730 ;
  assign n17928 = ~n6080 & n13252 ;
  assign n17929 = ~n17927 & n17928 ;
  assign n17930 = n1148 | n17929 ;
  assign n17931 = n11159 & ~n17930 ;
  assign n17932 = n367 | n2220 ;
  assign n17933 = n17932 ^ n5394 ^ 1'b0 ;
  assign n17934 = ~n11187 & n17933 ;
  assign n17935 = n3295 ^ n2068 ^ 1'b0 ;
  assign n17936 = n17935 ^ n748 ^ 1'b0 ;
  assign n17937 = n8031 ^ n2817 ^ 1'b0 ;
  assign n17938 = n17937 ^ n14003 ^ 1'b0 ;
  assign n17939 = n6051 & ~n17938 ;
  assign n17940 = n4848 & n9108 ;
  assign n17941 = ~n3270 & n13120 ;
  assign n17942 = n17941 ^ n11950 ^ 1'b0 ;
  assign n17943 = n13781 ^ n12542 ^ 1'b0 ;
  assign n17944 = n14168 ^ n321 ^ 1'b0 ;
  assign n17945 = n9111 | n17944 ;
  assign n17946 = n17945 ^ n17580 ^ 1'b0 ;
  assign n17947 = n8210 ^ n675 ^ 1'b0 ;
  assign n17948 = n8410 ^ n8269 ^ 1'b0 ;
  assign n17949 = n1064 & n17948 ;
  assign n17950 = ~n1619 & n17949 ;
  assign n17951 = n14200 | n17950 ;
  assign n17952 = n336 | n3801 ;
  assign n17953 = n743 | n17952 ;
  assign n17954 = n14382 ^ n190 ^ 1'b0 ;
  assign n17955 = n8868 & ~n17954 ;
  assign n17956 = ~n9986 & n17955 ;
  assign n17957 = ~n158 & n15146 ;
  assign n17958 = n4593 | n14114 ;
  assign n17959 = n17958 ^ n3722 ^ 1'b0 ;
  assign n17960 = n1080 & ~n4339 ;
  assign n17961 = ~n1745 & n17960 ;
  assign n17962 = n2642 & ~n17961 ;
  assign n17963 = n17962 ^ n11164 ^ 1'b0 ;
  assign n17964 = n8505 & n17134 ;
  assign n17965 = n17598 ^ n5462 ^ 1'b0 ;
  assign n17968 = n235 & n5735 ;
  assign n17969 = n17968 ^ n11012 ^ 1'b0 ;
  assign n17970 = n17969 ^ n754 ^ 1'b0 ;
  assign n17971 = n573 | n17970 ;
  assign n17966 = n1895 | n11083 ;
  assign n17967 = n8969 & ~n17966 ;
  assign n17972 = n17971 ^ n17967 ^ 1'b0 ;
  assign n17973 = n4277 ^ n3389 ^ 1'b0 ;
  assign n17974 = n17972 & n17973 ;
  assign n17975 = n15902 ^ n15469 ^ 1'b0 ;
  assign n17976 = n281 & ~n17975 ;
  assign n17984 = n89 | n7561 ;
  assign n17985 = n89 & ~n17984 ;
  assign n17977 = ~n1608 & n2804 ;
  assign n17978 = ~n2804 & n17977 ;
  assign n17979 = n9454 | n17978 ;
  assign n17980 = n9454 & ~n17979 ;
  assign n17981 = n2958 & ~n5749 ;
  assign n17982 = n17980 & n17981 ;
  assign n17983 = ~n2163 & n17982 ;
  assign n17986 = n17985 ^ n17983 ^ 1'b0 ;
  assign n17987 = n2236 & ~n14141 ;
  assign n17988 = n1125 & ~n2720 ;
  assign n17989 = n10532 & ~n17988 ;
  assign n17990 = n5800 & ~n7072 ;
  assign n17991 = n17990 ^ n2307 ^ 1'b0 ;
  assign n17992 = n15675 & n17991 ;
  assign n17993 = n813 ^ n748 ^ 1'b0 ;
  assign n17994 = ~n1516 & n7263 ;
  assign n17995 = n17994 ^ n4740 ^ 1'b0 ;
  assign n17996 = n17854 & n17995 ;
  assign n17997 = n15544 ^ n14782 ^ 1'b0 ;
  assign n17998 = n17997 ^ n14068 ^ n83 ;
  assign n17999 = n1844 ^ n1679 ^ 1'b0 ;
  assign n18000 = n17999 ^ n9371 ^ 1'b0 ;
  assign n18001 = n18000 ^ n2028 ^ 1'b0 ;
  assign n18002 = ~n5909 & n8457 ;
  assign n18003 = n9352 | n18002 ;
  assign n18004 = n13070 ^ n2601 ^ 1'b0 ;
  assign n18005 = n17477 ^ n3761 ^ 1'b0 ;
  assign n18006 = n6965 & n14168 ;
  assign n18007 = n10684 & n18006 ;
  assign n18008 = n9118 ^ n750 ^ 1'b0 ;
  assign n18009 = n18007 | n18008 ;
  assign n18010 = n315 & n18009 ;
  assign n18011 = n6258 ^ n616 ^ 1'b0 ;
  assign n18012 = n18011 ^ n7624 ^ 1'b0 ;
  assign n18013 = n9855 & n18012 ;
  assign n18016 = n7192 ^ n3741 ^ 1'b0 ;
  assign n18017 = n570 & n11053 ;
  assign n18018 = ~n18016 & n18017 ;
  assign n18014 = n9834 ^ n246 ^ 1'b0 ;
  assign n18015 = ~n13720 & n18014 ;
  assign n18019 = n18018 ^ n18015 ^ 1'b0 ;
  assign n18020 = n12974 ^ n1254 ^ 1'b0 ;
  assign n18021 = n4409 | n18020 ;
  assign n18022 = ( n1671 & n2927 ) | ( n1671 & n17561 ) | ( n2927 & n17561 ) ;
  assign n18023 = n2969 & ~n18022 ;
  assign n18024 = n14138 & n18023 ;
  assign n18025 = n11469 ^ n489 ^ 1'b0 ;
  assign n18026 = ~n3839 & n7710 ;
  assign n18027 = n7702 & ~n18026 ;
  assign n18028 = n18027 ^ n1266 ^ 1'b0 ;
  assign n18029 = n8874 ^ n6263 ^ 1'b0 ;
  assign n18030 = n18029 ^ n16534 ^ 1'b0 ;
  assign n18031 = n3693 & n3928 ;
  assign n18032 = n13857 ^ n223 ^ 1'b0 ;
  assign n18033 = n10100 & n14393 ;
  assign n18034 = n12877 ^ n7634 ^ 1'b0 ;
  assign n18035 = n6427 ^ n4261 ^ n3382 ;
  assign n18036 = n10186 & n18035 ;
  assign n18037 = n18036 ^ n938 ^ 1'b0 ;
  assign n18038 = ~n1170 & n6633 ;
  assign n18039 = n18037 & n18038 ;
  assign n18040 = n9478 | n17700 ;
  assign n18041 = n12300 & ~n18040 ;
  assign n18042 = n18041 ^ n8504 ^ 1'b0 ;
  assign n18043 = n939 & n18042 ;
  assign n18044 = n1252 & n4120 ;
  assign n18045 = n3696 & n18044 ;
  assign n18046 = n14464 ^ n9311 ^ 1'b0 ;
  assign n18047 = ( ~n7685 & n7866 ) | ( ~n7685 & n18046 ) | ( n7866 & n18046 ) ;
  assign n18048 = ~n4054 & n4913 ;
  assign n18049 = n18048 ^ n1533 ^ 1'b0 ;
  assign n18050 = n13435 ^ n7114 ^ 1'b0 ;
  assign n18051 = n12252 | n18050 ;
  assign n18052 = n5713 ^ n673 ^ 1'b0 ;
  assign n18053 = n18052 ^ n5751 ^ 1'b0 ;
  assign n18054 = ~n9849 & n18053 ;
  assign n18055 = n18054 ^ n3579 ^ 1'b0 ;
  assign n18056 = n1702 & n3282 ;
  assign n18057 = n18056 ^ n9377 ^ 1'b0 ;
  assign n18058 = n879 & ~n18057 ;
  assign n18059 = n18058 ^ n13321 ^ 1'b0 ;
  assign n18060 = n9837 | n18059 ;
  assign n18061 = ( n5128 & n7541 ) | ( n5128 & n18060 ) | ( n7541 & n18060 ) ;
  assign n18062 = n257 | n16416 ;
  assign n18063 = n1693 ^ n404 ^ 1'b0 ;
  assign n18064 = ~n556 & n18063 ;
  assign n18065 = n241 & n18064 ;
  assign n18066 = n5507 | n18065 ;
  assign n18067 = n2326 & ~n18066 ;
  assign n18068 = n18067 ^ n2432 ^ 1'b0 ;
  assign n18069 = n9623 | n18068 ;
  assign n18070 = n404 | n8086 ;
  assign n18071 = n5814 & ~n18070 ;
  assign n18072 = n1564 & n18071 ;
  assign n18073 = n931 ^ n114 ^ 1'b0 ;
  assign n18074 = ~n12098 & n13790 ;
  assign n18075 = n198 | n954 ;
  assign n18076 = n954 & ~n18075 ;
  assign n18077 = ~n4025 & n18076 ;
  assign n18078 = n609 | n18077 ;
  assign n18079 = n609 & ~n18078 ;
  assign n18080 = n1863 | n18079 ;
  assign n18081 = n18079 & ~n18080 ;
  assign n18082 = ~n3442 & n8282 ;
  assign n18083 = n6417 ^ n4934 ^ 1'b0 ;
  assign n18084 = n3527 | n15879 ;
  assign n18085 = n5366 & n6330 ;
  assign n18086 = n18085 ^ n191 ^ 1'b0 ;
  assign n18087 = n12255 ^ n9043 ^ 1'b0 ;
  assign n18088 = n1067 & ~n1722 ;
  assign n18089 = n9697 & n12868 ;
  assign n18090 = ~n10635 & n18089 ;
  assign n18091 = x6 & n6043 ;
  assign n18092 = n18091 ^ n212 ^ 1'b0 ;
  assign n18093 = n14226 & n18092 ;
  assign n18094 = n839 & n8649 ;
  assign n18095 = n18094 ^ n2818 ^ 1'b0 ;
  assign n18096 = n977 & ~n18095 ;
  assign n18097 = n15139 & ~n18096 ;
  assign n18098 = n2778 & n4076 ;
  assign n18099 = ~n6162 & n18098 ;
  assign n18100 = n18099 ^ n1118 ^ 1'b0 ;
  assign n18101 = n6682 & ~n13121 ;
  assign n18102 = n18101 ^ n2331 ^ 1'b0 ;
  assign n18103 = n18102 ^ n726 ^ 1'b0 ;
  assign n18105 = n7433 ^ n122 ^ 1'b0 ;
  assign n18106 = n1686 & n18105 ;
  assign n18104 = ~n1522 & n8898 ;
  assign n18107 = n18106 ^ n18104 ^ 1'b0 ;
  assign n18108 = n1342 & ~n10212 ;
  assign n18109 = n18108 ^ n15034 ^ 1'b0 ;
  assign n18110 = n2467 ^ n169 ^ 1'b0 ;
  assign n18111 = n17092 ^ n14408 ^ 1'b0 ;
  assign n18112 = n3074 | n18111 ;
  assign n18113 = ~n866 & n10452 ;
  assign n18114 = n11521 & n18113 ;
  assign n18115 = n439 & n596 ;
  assign n18116 = n588 | n18115 ;
  assign n18117 = n13447 & ~n16762 ;
  assign n18118 = n18117 ^ n2585 ^ 1'b0 ;
  assign n18119 = n6487 & n13691 ;
  assign n18120 = n18119 ^ n2930 ^ 1'b0 ;
  assign n18121 = ~n1447 & n18120 ;
  assign n18122 = n4419 & ~n18121 ;
  assign n18123 = n6174 & n18122 ;
  assign n18124 = n5070 ^ n1898 ^ 1'b0 ;
  assign n18125 = n2361 ^ n1663 ^ 1'b0 ;
  assign n18126 = ~n4095 & n18125 ;
  assign n18127 = ~n18124 & n18126 ;
  assign n18128 = n10217 ^ n294 ^ 1'b0 ;
  assign n18129 = ~n6385 & n8992 ;
  assign n18130 = n18129 ^ n5050 ^ 1'b0 ;
  assign n18131 = n6677 | n14203 ;
  assign n18132 = n18131 ^ n14924 ^ 1'b0 ;
  assign n18133 = n2185 & n14806 ;
  assign n18134 = ~n14928 & n18133 ;
  assign n18135 = ~n11298 & n18134 ;
  assign n18136 = n18135 ^ n11586 ^ 1'b0 ;
  assign n18137 = n5264 ^ n73 ^ 1'b0 ;
  assign n18138 = ~n46 & n18137 ;
  assign n18139 = n9794 ^ n2426 ^ 1'b0 ;
  assign n18140 = n619 & n5237 ;
  assign n18141 = n1910 & ~n18140 ;
  assign n18142 = n18141 ^ n13028 ^ 1'b0 ;
  assign n18143 = n671 & ~n9968 ;
  assign n18144 = n9326 & n18143 ;
  assign n18145 = n7428 ^ n3995 ^ 1'b0 ;
  assign n18146 = n10026 | n10074 ;
  assign n18147 = n18146 ^ n1281 ^ 1'b0 ;
  assign n18148 = n495 | n4628 ;
  assign n18149 = n1886 | n18148 ;
  assign n18150 = n11542 | n18149 ;
  assign n18151 = n6250 & ~n12082 ;
  assign n18152 = n302 & n18151 ;
  assign n18153 = n8747 & ~n16746 ;
  assign n18154 = n151 & n18153 ;
  assign n18155 = n4487 & n6490 ;
  assign n18156 = ~n519 & n18155 ;
  assign n18158 = ~n7450 & n10938 ;
  assign n18157 = n4321 & ~n10978 ;
  assign n18159 = n18158 ^ n18157 ^ 1'b0 ;
  assign n18160 = n40 & ~n66 ;
  assign n18161 = n66 & n18160 ;
  assign n18162 = n279 | n989 ;
  assign n18163 = n989 & ~n18162 ;
  assign n18164 = n2364 & ~n18163 ;
  assign n18165 = ~n2364 & n18164 ;
  assign n18166 = n1431 & n18165 ;
  assign n18167 = n414 & n18166 ;
  assign n18168 = ~n1179 & n18167 ;
  assign n18169 = n18168 ^ n6333 ^ 1'b0 ;
  assign n18170 = n18161 | n18169 ;
  assign n18171 = n1569 | n8994 ;
  assign n18172 = n3406 & ~n18171 ;
  assign n18173 = n18172 ^ n4549 ^ 1'b0 ;
  assign n18174 = n1155 & ~n15060 ;
  assign n18175 = n5471 | n12457 ;
  assign n18176 = n1060 & n16043 ;
  assign n18177 = n5749 | n11111 ;
  assign n18178 = n17502 & ~n18177 ;
  assign n18179 = n8660 ^ n6512 ^ n5673 ;
  assign n18180 = n7469 & ~n13160 ;
  assign n18181 = n18180 ^ n17156 ^ 1'b0 ;
  assign n18182 = n4550 ^ n540 ^ 1'b0 ;
  assign n18183 = ~n11333 & n18182 ;
  assign n18184 = n3584 & n18183 ;
  assign n18185 = n18184 ^ n14984 ^ 1'b0 ;
  assign n18186 = n7494 ^ n4436 ^ 1'b0 ;
  assign n18187 = n18186 ^ n2824 ^ 1'b0 ;
  assign n18188 = n18187 ^ n1947 ^ 1'b0 ;
  assign n18189 = n3957 & n14797 ;
  assign n18190 = n719 | n5040 ;
  assign n18191 = ~n86 & n1355 ;
  assign n18192 = n311 | n18191 ;
  assign n18193 = ~n310 & n12859 ;
  assign n18194 = n5977 ^ n161 ^ 1'b0 ;
  assign n18195 = ~n68 & n18194 ;
  assign n18196 = n929 & ~n8365 ;
  assign n18197 = n18196 ^ n2168 ^ 1'b0 ;
  assign n18198 = n18195 & n18197 ;
  assign n18199 = n18198 ^ n5953 ^ 1'b0 ;
  assign n18200 = n18199 ^ n455 ^ 1'b0 ;
  assign n18201 = n1469 ^ n227 ^ 1'b0 ;
  assign n18202 = ~n2853 & n12454 ;
  assign n18203 = ~n4013 & n18202 ;
  assign n18204 = ~n1339 & n6441 ;
  assign n18205 = n18204 ^ n5319 ^ 1'b0 ;
  assign n18206 = n9493 ^ n3122 ^ 1'b0 ;
  assign n18207 = ~n79 & n18206 ;
  assign n18208 = n1854 ^ n820 ^ 1'b0 ;
  assign n18209 = n6011 & n18208 ;
  assign n18210 = n18207 & n18209 ;
  assign n18211 = n18210 ^ n9307 ^ 1'b0 ;
  assign n18212 = n8789 ^ n6104 ^ 1'b0 ;
  assign n18213 = ~n3791 & n11777 ;
  assign n18215 = n478 | n17776 ;
  assign n18216 = n6079 | n18215 ;
  assign n18217 = n18216 ^ n6016 ^ 1'b0 ;
  assign n18214 = n6629 | n15862 ;
  assign n18218 = n18217 ^ n18214 ^ 1'b0 ;
  assign n18219 = n197 & n11254 ;
  assign n18224 = n6617 ^ n2418 ^ 1'b0 ;
  assign n18220 = n4949 & ~n6339 ;
  assign n18221 = ~n3040 & n18220 ;
  assign n18222 = n8117 & n18221 ;
  assign n18223 = ~n12114 & n18222 ;
  assign n18225 = n18224 ^ n18223 ^ 1'b0 ;
  assign n18226 = n8262 & ~n18225 ;
  assign n18227 = n5612 | n10241 ;
  assign n18228 = n10156 ^ n2618 ^ n1227 ;
  assign n18229 = n991 & n13172 ;
  assign n18230 = n17115 ^ n15985 ^ 1'b0 ;
  assign n18231 = n18229 & ~n18230 ;
  assign n18232 = n13594 ^ n11063 ^ 1'b0 ;
  assign n18233 = n16100 & ~n18232 ;
  assign n18235 = n2936 ^ n2181 ^ 1'b0 ;
  assign n18236 = n16931 & ~n18235 ;
  assign n18234 = n8971 & ~n14134 ;
  assign n18237 = n18236 ^ n18234 ^ 1'b0 ;
  assign n18238 = n9166 & n11373 ;
  assign n18239 = n18238 ^ n832 ^ 1'b0 ;
  assign n18240 = n8318 ^ n172 ^ 1'b0 ;
  assign n18241 = n10509 | n18240 ;
  assign n18242 = n2644 ^ n216 ^ 1'b0 ;
  assign n18243 = n3939 | n13409 ;
  assign n18244 = n15244 ^ n13119 ^ 1'b0 ;
  assign n18245 = n18244 ^ n461 ^ 1'b0 ;
  assign n18246 = n18243 & n18245 ;
  assign n18247 = ~n11025 & n18246 ;
  assign n18248 = n726 & ~n6645 ;
  assign n18249 = n6133 & n6655 ;
  assign n18250 = ~n4183 & n18249 ;
  assign n18251 = n532 & n2085 ;
  assign n18252 = n18251 ^ n1193 ^ 1'b0 ;
  assign n18253 = n1937 & n18252 ;
  assign n18254 = n7449 & n18253 ;
  assign n18255 = n9233 & n18254 ;
  assign n18256 = n6579 ^ n3134 ^ 1'b0 ;
  assign n18257 = n2311 & n6061 ;
  assign n18258 = ~n18256 & n18257 ;
  assign n18259 = n11295 & ~n13170 ;
  assign n18260 = n5890 & ~n13753 ;
  assign n18261 = n18260 ^ n1704 ^ 1'b0 ;
  assign n18262 = n2662 & n15067 ;
  assign n18263 = n717 & n6618 ;
  assign n18264 = ~n9219 & n18263 ;
  assign n18265 = n18264 ^ n16568 ^ 1'b0 ;
  assign n18266 = n6878 | n18265 ;
  assign n18267 = ( n393 & n3855 ) | ( n393 & n17013 ) | ( n3855 & n17013 ) ;
  assign n18268 = n664 | n1194 ;
  assign n18269 = n129 & n12862 ;
  assign n18270 = n18269 ^ n3764 ^ 1'b0 ;
  assign n18271 = n5566 ^ n2618 ^ 1'b0 ;
  assign n18272 = ~n2539 & n14918 ;
  assign n18273 = n107 | n17952 ;
  assign n18274 = n18273 ^ n364 ^ 1'b0 ;
  assign n18275 = n297 & ~n621 ;
  assign n18276 = ~n18274 & n18275 ;
  assign n18277 = ~n4374 & n5324 ;
  assign n18280 = n3584 ^ n3146 ^ 1'b0 ;
  assign n18281 = n2103 ^ n1739 ^ 1'b0 ;
  assign n18282 = n1337 | n18281 ;
  assign n18283 = n6399 ^ n1384 ^ 1'b0 ;
  assign n18284 = ~n1170 & n18283 ;
  assign n18285 = ~n18282 & n18284 ;
  assign n18286 = n18280 & n18285 ;
  assign n18278 = n2007 & n14409 ;
  assign n18279 = n17157 & ~n18278 ;
  assign n18287 = n18286 ^ n18279 ^ 1'b0 ;
  assign n18288 = n18277 & n18287 ;
  assign n18289 = n10751 ^ n7460 ^ 1'b0 ;
  assign n18290 = n16601 ^ n15602 ^ 1'b0 ;
  assign n18291 = n6139 & ~n18290 ;
  assign n18292 = n18291 ^ n15770 ^ 1'b0 ;
  assign n18293 = n4690 & n13528 ;
  assign n18294 = ~n1051 & n5150 ;
  assign n18295 = n6244 | n7340 ;
  assign n18296 = n2880 ^ n2183 ^ 1'b0 ;
  assign n18297 = n18295 & ~n18296 ;
  assign n18298 = ~n4734 & n6131 ;
  assign n18299 = n16153 | n18298 ;
  assign n18300 = n4122 ^ n94 ^ 1'b0 ;
  assign n18301 = n6356 ^ n2549 ^ 1'b0 ;
  assign n18302 = ~n13455 & n18301 ;
  assign n18303 = n10982 ^ n7329 ^ 1'b0 ;
  assign n18304 = ~n1452 & n11425 ;
  assign n18305 = n8668 ^ n7409 ^ 1'b0 ;
  assign n18306 = n9072 ^ n1235 ^ 1'b0 ;
  assign n18307 = n18306 ^ n15720 ^ 1'b0 ;
  assign n18308 = n9398 ^ n4377 ^ 1'b0 ;
  assign n18309 = n717 & n15775 ;
  assign n18310 = n18308 & n18309 ;
  assign n18311 = n6174 & n10184 ;
  assign n18312 = n5445 & ~n5815 ;
  assign n18315 = n5025 | n10080 ;
  assign n18313 = n11174 ^ n3072 ^ 1'b0 ;
  assign n18314 = ~n11797 & n18313 ;
  assign n18316 = n18315 ^ n18314 ^ n139 ;
  assign n18317 = n9954 & ~n12366 ;
  assign n18318 = n18317 ^ n6150 ^ 1'b0 ;
  assign n18319 = n246 | n18318 ;
  assign n18320 = ~n1229 & n3669 ;
  assign n18321 = n43 & n3034 ;
  assign n18322 = n18321 ^ n8692 ^ 1'b0 ;
  assign n18323 = n7981 ^ n6281 ^ 1'b0 ;
  assign n18324 = ~n1284 & n18323 ;
  assign n18325 = ~n6274 & n13238 ;
  assign n18326 = ~n1109 & n5996 ;
  assign n18327 = n18326 ^ n16719 ^ 1'b0 ;
  assign n18328 = ~n745 & n18327 ;
  assign n18329 = n16577 | n18317 ;
  assign n18330 = n18329 ^ n4329 ^ 1'b0 ;
  assign n18331 = n1165 & ~n3793 ;
  assign n18332 = ~n8974 & n18331 ;
  assign n18333 = n8288 & ~n15853 ;
  assign n18334 = n5288 & ~n18333 ;
  assign n18335 = n4424 | n7288 ;
  assign n18336 = n10251 & ~n18335 ;
  assign n18337 = n17308 ^ n10662 ^ n1144 ;
  assign n18338 = n8967 ^ n4181 ^ 1'b0 ;
  assign n18339 = n2899 & ~n18338 ;
  assign n18340 = ~n8212 & n18339 ;
  assign n18341 = ~n252 & n5284 ;
  assign n18342 = n18341 ^ n2870 ^ 1'b0 ;
  assign n18343 = n1637 | n18342 ;
  assign n18344 = n6534 | n18343 ;
  assign n18345 = ~n743 & n3655 ;
  assign n18346 = ~n1292 & n18345 ;
  assign n18347 = ~n1169 & n5894 ;
  assign n18348 = n18347 ^ n6939 ^ 1'b0 ;
  assign n18349 = n4749 ^ n2270 ^ 1'b0 ;
  assign n18350 = n18349 ^ n2941 ^ 1'b0 ;
  assign n18351 = n2549 | n3682 ;
  assign n18352 = n1529 & n18351 ;
  assign n18353 = n555 & ~n1218 ;
  assign n18354 = n18353 ^ n1686 ^ 1'b0 ;
  assign n18355 = n17537 & ~n18354 ;
  assign n18356 = n14165 | n18355 ;
  assign n18357 = ( n6933 & n18352 ) | ( n6933 & ~n18356 ) | ( n18352 & ~n18356 ) ;
  assign n18358 = ~n1785 & n4121 ;
  assign n18359 = n1418 | n5428 ;
  assign n18360 = n13961 ^ n12954 ^ 1'b0 ;
  assign n18361 = ~n5055 & n18360 ;
  assign n18362 = n6558 ^ n4650 ^ 1'b0 ;
  assign n18363 = ~n7181 & n18362 ;
  assign n18365 = ~n64 & n5556 ;
  assign n18364 = n3848 & ~n17605 ;
  assign n18366 = n18365 ^ n18364 ^ 1'b0 ;
  assign n18367 = n1827 ^ n1406 ^ 1'b0 ;
  assign n18368 = n3598 | n5655 ;
  assign n18369 = n18368 ^ n3384 ^ 1'b0 ;
  assign n18370 = n18369 ^ n2194 ^ n2072 ;
  assign n18371 = ~n1840 & n18370 ;
  assign n18372 = n18367 & n18371 ;
  assign n18373 = n18372 ^ n3273 ^ 1'b0 ;
  assign n18374 = ~n6536 & n18373 ;
  assign n18375 = ~n2106 & n18374 ;
  assign n18376 = n257 & ~n9158 ;
  assign n18377 = n18376 ^ n94 ^ 1'b0 ;
  assign n18378 = n16424 & n18377 ;
  assign n18379 = ~n9023 & n11968 ;
  assign n18380 = n2699 & n18379 ;
  assign n18381 = n9166 ^ n1613 ^ 1'b0 ;
  assign n18382 = ~n9534 & n16792 ;
  assign n18383 = n2440 ^ n1912 ^ 1'b0 ;
  assign n18384 = n69 & n2193 ;
  assign n18385 = ~n18383 & n18384 ;
  assign n18387 = n13308 ^ n10831 ^ 1'b0 ;
  assign n18386 = ~n2036 & n3321 ;
  assign n18388 = n18387 ^ n18386 ^ 1'b0 ;
  assign n18389 = n8102 ^ n3946 ^ 1'b0 ;
  assign n18390 = n784 & n18389 ;
  assign n18391 = n6971 | n18390 ;
  assign n18392 = n2001 & n4703 ;
  assign n18393 = n2532 | n3749 ;
  assign n18394 = n17656 | n18393 ;
  assign n18395 = n7093 | n17141 ;
  assign n18396 = n2983 & ~n18395 ;
  assign n18397 = n7469 & ~n18396 ;
  assign n18398 = ~n18394 & n18397 ;
  assign n18399 = n17594 ^ n16833 ^ 1'b0 ;
  assign n18400 = n3514 & ~n18399 ;
  assign n18401 = ~n4966 & n8513 ;
  assign n18402 = n18401 ^ n133 ^ 1'b0 ;
  assign n18403 = n6871 & n17160 ;
  assign n18404 = n11225 ^ n7104 ^ 1'b0 ;
  assign n18405 = n4261 & ~n18404 ;
  assign n18406 = n10743 & ~n18405 ;
  assign n18407 = ( n2932 & n18403 ) | ( n2932 & n18406 ) | ( n18403 & n18406 ) ;
  assign n18408 = n3512 & n8749 ;
  assign n18409 = ~n1515 & n16835 ;
  assign n18410 = n18409 ^ n9375 ^ 1'b0 ;
  assign n18411 = n9544 ^ n87 ^ 1'b0 ;
  assign n18412 = n8488 & ~n18411 ;
  assign n18413 = n18410 & n18412 ;
  assign n18414 = n18413 ^ n9319 ^ 1'b0 ;
  assign n18415 = n13801 ^ n8081 ^ 1'b0 ;
  assign n18416 = ~n941 & n7870 ;
  assign n18417 = n2059 & n18416 ;
  assign n18418 = ~n4322 & n18417 ;
  assign n18419 = n18418 ^ n6874 ^ n4780 ;
  assign n18420 = n12649 | n18419 ;
  assign n18421 = n532 | n18420 ;
  assign n18422 = n18421 ^ n5223 ^ 1'b0 ;
  assign n18423 = n6596 | n6786 ;
  assign n18424 = n172 & n5451 ;
  assign n18425 = ~n2260 & n3743 ;
  assign n18426 = n18424 & n18425 ;
  assign n18427 = n18426 ^ n16820 ^ 1'b0 ;
  assign n18428 = n4169 & ~n18427 ;
  assign n18429 = n6368 ^ n3802 ^ 1'b0 ;
  assign n18430 = n1310 & n18429 ;
  assign n18431 = ~n704 & n18430 ;
  assign n18432 = ~n18428 & n18431 ;
  assign n18433 = n1652 & n13298 ;
  assign n18434 = n10141 ^ n2575 ^ 1'b0 ;
  assign n18438 = n7825 ^ n116 ^ 1'b0 ;
  assign n18439 = n18438 ^ n8574 ^ 1'b0 ;
  assign n18435 = n7328 & ~n10107 ;
  assign n18436 = n18435 ^ n14500 ^ 1'b0 ;
  assign n18437 = n2027 | n18436 ;
  assign n18440 = n18439 ^ n18437 ^ 1'b0 ;
  assign n18441 = ~n11934 & n18440 ;
  assign n18442 = ~n18440 & n18441 ;
  assign n18443 = n18442 ^ n3112 ^ 1'b0 ;
  assign n18444 = n18434 & ~n18443 ;
  assign n18445 = ~n18434 & n18444 ;
  assign n18446 = n8628 & ~n9292 ;
  assign n18447 = n876 | n15582 ;
  assign n18448 = n11024 & ~n18447 ;
  assign n18449 = n13295 ^ n8064 ^ 1'b0 ;
  assign n18450 = n37 | n3598 ;
  assign n18451 = ~n18449 & n18450 ;
  assign n18452 = n6401 & ~n7736 ;
  assign n18453 = n18452 ^ n3692 ^ 1'b0 ;
  assign n18454 = n18453 ^ n11555 ^ 1'b0 ;
  assign n18455 = n3374 & ~n18454 ;
  assign n18456 = n12440 & ~n18455 ;
  assign n18461 = ~n495 & n3479 ;
  assign n18462 = n8448 & n18461 ;
  assign n18457 = n6590 & ~n8201 ;
  assign n18458 = n18457 ^ n123 ^ 1'b0 ;
  assign n18459 = n10678 | n18458 ;
  assign n18460 = n11242 | n18459 ;
  assign n18463 = n18462 ^ n18460 ^ 1'b0 ;
  assign n18464 = n51 & n18463 ;
  assign n18465 = ~n7216 & n8377 ;
  assign n18466 = n18465 ^ n9833 ^ 1'b0 ;
  assign n18467 = n570 & ~n18466 ;
  assign n18468 = n18467 ^ n15820 ^ 1'b0 ;
  assign n18469 = ~n1298 & n3352 ;
  assign n18470 = n8239 ^ n7019 ^ 1'b0 ;
  assign n18471 = n8381 & ~n18470 ;
  assign n18472 = ~n2017 & n18471 ;
  assign n18473 = n9898 ^ n6937 ^ 1'b0 ;
  assign n18474 = n5073 & ~n9507 ;
  assign n18475 = n2769 ^ n1425 ^ 1'b0 ;
  assign n18476 = ~n9051 & n18475 ;
  assign n18477 = n3408 & ~n7504 ;
  assign n18478 = n8765 & n18477 ;
  assign n18479 = n2235 & ~n18478 ;
  assign n18480 = n13750 & n18479 ;
  assign n18481 = n4228 ^ n2110 ^ 1'b0 ;
  assign n18482 = n18481 ^ n4748 ^ 1'b0 ;
  assign n18483 = n764 & n18482 ;
  assign n18484 = n3027 & ~n6176 ;
  assign n18485 = n4300 ^ n164 ^ 1'b0 ;
  assign n18486 = ~n6187 & n18485 ;
  assign n18487 = n18486 ^ n633 ^ 1'b0 ;
  assign n18488 = n5554 & n12679 ;
  assign n18489 = n5707 & n7955 ;
  assign n18490 = ~n1045 & n18489 ;
  assign n18491 = n11721 | n16310 ;
  assign n18492 = n18490 & ~n18491 ;
  assign n18493 = n6210 ^ n628 ^ 1'b0 ;
  assign n18494 = n622 & n18493 ;
  assign n18495 = n10942 & n18494 ;
  assign n18496 = n9257 & n18495 ;
  assign n18497 = n5560 ^ n5551 ^ 1'b0 ;
  assign n18498 = ~x0 & n147 ;
  assign n18499 = n2294 & ~n18498 ;
  assign n18500 = ~n2294 & n18499 ;
  assign n18501 = n18500 ^ n4827 ^ 1'b0 ;
  assign n18502 = n12167 | n18501 ;
  assign n18503 = n18497 & ~n18502 ;
  assign n18504 = ( n114 & n2726 ) | ( n114 & n13610 ) | ( n2726 & n13610 ) ;
  assign n18505 = n18504 ^ n10908 ^ n561 ;
  assign n18506 = n2512 | n6320 ;
  assign n18507 = n2489 ^ n25 ^ 1'b0 ;
  assign n18508 = n18507 ^ n713 ^ 1'b0 ;
  assign n18509 = ~n10828 & n14098 ;
  assign n18510 = n519 & n3083 ;
  assign n18511 = n18510 ^ n828 ^ 1'b0 ;
  assign n18512 = ~n6360 & n8649 ;
  assign n18513 = n18512 ^ n11780 ^ 1'b0 ;
  assign n18514 = n13108 & ~n18513 ;
  assign n18515 = n18514 ^ n7185 ^ 1'b0 ;
  assign n18516 = n2797 & ~n6385 ;
  assign n18517 = ~n2848 & n18516 ;
  assign n18518 = n14696 & n18517 ;
  assign n18519 = n9959 & ~n14007 ;
  assign n18520 = n182 & ~n5269 ;
  assign n18521 = n8705 ^ n1619 ^ 1'b0 ;
  assign n18522 = n7297 ^ n3263 ^ 1'b0 ;
  assign n18523 = n1533 | n15247 ;
  assign n18524 = ~n1539 & n18523 ;
  assign n18525 = n18524 ^ n5551 ^ 1'b0 ;
  assign n18526 = n18525 ^ n3694 ^ 1'b0 ;
  assign n18529 = n532 | n1804 ;
  assign n18530 = n18529 ^ n4043 ^ 1'b0 ;
  assign n18527 = n5735 & n8365 ;
  assign n18528 = n18527 ^ n12090 ^ 1'b0 ;
  assign n18531 = n18530 ^ n18528 ^ 1'b0 ;
  assign n18532 = n1560 | n18531 ;
  assign n18533 = n18532 ^ n12404 ^ 1'b0 ;
  assign n18534 = n10746 ^ n5774 ^ n2072 ;
  assign n18535 = ~n348 & n18534 ;
  assign n18536 = n7981 & n18535 ;
  assign n18537 = n6258 & n12948 ;
  assign n18543 = n4263 | n6244 ;
  assign n18544 = n785 | n18543 ;
  assign n18539 = n1048 & ~n1864 ;
  assign n18540 = n18539 ^ n3251 ^ 1'b0 ;
  assign n18541 = n18540 ^ n1441 ^ n372 ;
  assign n18542 = n18541 ^ n6067 ^ 1'b0 ;
  assign n18538 = ~n712 & n15117 ;
  assign n18545 = n18544 ^ n18542 ^ n18538 ;
  assign n18546 = n7210 ^ n4185 ^ 1'b0 ;
  assign n18547 = ~n2117 & n18546 ;
  assign n18548 = n18547 ^ n1194 ^ 1'b0 ;
  assign n18549 = n863 & n3493 ;
  assign n18550 = n18549 ^ n2732 ^ 1'b0 ;
  assign n18551 = n1888 | n18550 ;
  assign n18552 = n18551 ^ n3007 ^ 1'b0 ;
  assign n18553 = n18552 ^ n8070 ^ 1'b0 ;
  assign n18554 = n14737 | n18553 ;
  assign n18555 = n6890 ^ x1 ^ 1'b0 ;
  assign n18556 = n15629 ^ n5891 ^ 1'b0 ;
  assign n18557 = n4453 | n11313 ;
  assign n18558 = ( n4510 & n5713 ) | ( n4510 & n18557 ) | ( n5713 & n18557 ) ;
  assign n18559 = n11324 ^ n4463 ^ 1'b0 ;
  assign n18560 = n18558 | n18559 ;
  assign n18561 = n9714 ^ n8114 ^ 1'b0 ;
  assign n18562 = ~n8351 & n18561 ;
  assign n18563 = n13732 & ~n16792 ;
  assign n18564 = n5868 & n17889 ;
  assign n18565 = ~n2502 & n10959 ;
  assign n18566 = n18565 ^ n12177 ^ 1'b0 ;
  assign n18567 = n4688 & n18566 ;
  assign n18568 = n4292 & n18567 ;
  assign n18569 = ~n1088 & n3988 ;
  assign n18570 = n13174 ^ n5568 ^ 1'b0 ;
  assign n18571 = n6345 ^ n3635 ^ 1'b0 ;
  assign n18572 = n18570 & ~n18571 ;
  assign n18573 = n218 & ~n1491 ;
  assign n18574 = n18573 ^ n3306 ^ 1'b0 ;
  assign n18575 = n15799 ^ n8910 ^ 1'b0 ;
  assign n18579 = n2655 & ~n6884 ;
  assign n18576 = ~n2465 & n7670 ;
  assign n18577 = n18576 ^ n4573 ^ 1'b0 ;
  assign n18578 = n18577 ^ n14910 ^ 1'b0 ;
  assign n18580 = n18579 ^ n18578 ^ 1'b0 ;
  assign n18581 = n17218 ^ n7365 ^ 1'b0 ;
  assign n18582 = n1671 & ~n7688 ;
  assign n18583 = ~n133 & n3509 ;
  assign n18584 = n12655 ^ n8644 ^ 1'b0 ;
  assign n18585 = n628 & ~n18584 ;
  assign n18586 = n6519 | n7128 ;
  assign n18587 = n8587 | n18586 ;
  assign n18588 = n7093 & n18587 ;
  assign n18589 = ~n1366 & n1693 ;
  assign n18590 = ~n1137 & n12797 ;
  assign n18591 = n384 & ~n666 ;
  assign n18592 = n9090 | n18591 ;
  assign n18593 = n15718 & n18592 ;
  assign n18594 = n4660 & n13857 ;
  assign n18595 = n18594 ^ n1707 ^ 1'b0 ;
  assign n18596 = n18595 ^ n6162 ^ 1'b0 ;
  assign n18597 = ~n512 & n11316 ;
  assign n18598 = ~n7311 & n18597 ;
  assign n18599 = n2225 & ~n18598 ;
  assign n18600 = ~n18596 & n18599 ;
  assign n18601 = n15866 ^ n1887 ^ 1'b0 ;
  assign n18602 = n13971 & ~n14905 ;
  assign n18603 = n18602 ^ n10368 ^ 1'b0 ;
  assign n18604 = n8885 | n9986 ;
  assign n18605 = n1662 | n18604 ;
  assign n18606 = n7265 | n8226 ;
  assign n18607 = n11409 & ~n18606 ;
  assign n18608 = n11119 ^ n8065 ^ 1'b0 ;
  assign n18612 = n270 & ~n9992 ;
  assign n18613 = ~n10285 & n18612 ;
  assign n18609 = n8651 ^ n5041 ^ 1'b0 ;
  assign n18610 = n3990 & ~n18609 ;
  assign n18611 = ~n17109 & n18610 ;
  assign n18614 = n18613 ^ n18611 ^ 1'b0 ;
  assign n18616 = n1547 & ~n2073 ;
  assign n18617 = n2073 & n18616 ;
  assign n18615 = n2738 | n7007 ;
  assign n18618 = n18617 ^ n18615 ^ 1'b0 ;
  assign n18619 = ~n2509 & n5825 ;
  assign n18620 = n11283 ^ n5551 ^ 1'b0 ;
  assign n18621 = n2537 & ~n18620 ;
  assign n18622 = n8082 & ~n18621 ;
  assign n18623 = n4057 & ~n4918 ;
  assign n18624 = n4532 ^ n3599 ^ 1'b0 ;
  assign n18625 = n18624 ^ n12046 ^ 1'b0 ;
  assign n18626 = n18625 ^ n13800 ^ n3559 ;
  assign n18627 = n3376 & ~n6916 ;
  assign n18628 = n18627 ^ n4927 ^ 1'b0 ;
  assign n18629 = n293 & ~n18628 ;
  assign n18630 = n3380 & ~n4453 ;
  assign n18631 = ~n2349 & n18630 ;
  assign n18632 = n18631 ^ n627 ^ 1'b0 ;
  assign n18633 = ~n3591 & n7715 ;
  assign n18634 = n18633 ^ n6653 ^ 1'b0 ;
  assign n18635 = n14089 ^ n8629 ^ 1'b0 ;
  assign n18636 = n102 | n9383 ;
  assign n18637 = n7457 & n8018 ;
  assign n18638 = n10235 ^ n1367 ^ 1'b0 ;
  assign n18639 = n11963 & ~n18504 ;
  assign n18640 = n18639 ^ n10874 ^ 1'b0 ;
  assign n18641 = n8768 & ~n18640 ;
  assign n18642 = n10239 ^ n6025 ^ 1'b0 ;
  assign n18643 = n2059 & ~n7476 ;
  assign n18644 = n9577 & n11561 ;
  assign n18645 = n18644 ^ n2515 ^ 1'b0 ;
  assign n18646 = n18645 ^ n13065 ^ 1'b0 ;
  assign n18647 = n1466 & n6106 ;
  assign n18648 = n8005 & n18647 ;
  assign n18649 = n7026 & n13656 ;
  assign n18650 = n18649 ^ n12438 ^ 1'b0 ;
  assign n18651 = n3311 & n17463 ;
  assign n18652 = n2038 & ~n8519 ;
  assign n18653 = n1968 & ~n18652 ;
  assign n18654 = ~n7489 & n18653 ;
  assign n18658 = n354 & n581 ;
  assign n18659 = n18658 ^ n3141 ^ 1'b0 ;
  assign n18660 = n2964 & ~n18659 ;
  assign n18655 = ~n1310 & n13408 ;
  assign n18656 = n5835 | n18655 ;
  assign n18657 = n16678 & ~n18656 ;
  assign n18661 = n18660 ^ n18657 ^ 1'b0 ;
  assign n18662 = n2567 & ~n18661 ;
  assign n18663 = n16356 ^ n12903 ^ 1'b0 ;
  assign n18664 = n18663 ^ n18097 ^ 1'b0 ;
  assign n18665 = ~n7947 & n16712 ;
  assign n18666 = n18665 ^ n15269 ^ 1'b0 ;
  assign n18674 = ~n2395 & n2882 ;
  assign n18675 = n17412 & n18674 ;
  assign n18676 = n149 & n635 ;
  assign n18677 = ~n149 & n18676 ;
  assign n18678 = n412 & ~n18677 ;
  assign n18679 = n18677 & n18678 ;
  assign n18680 = n292 & n18679 ;
  assign n18681 = n83 & n18680 ;
  assign n18682 = n3911 | n18681 ;
  assign n18683 = n18675 & ~n18682 ;
  assign n18684 = n73 & n121 ;
  assign n18685 = ~n121 & n18684 ;
  assign n18686 = n16 & ~n80 ;
  assign n18687 = n18685 & n18686 ;
  assign n18688 = n12829 | n18687 ;
  assign n18689 = n12829 & ~n18688 ;
  assign n18690 = n294 & ~n18689 ;
  assign n18691 = n18689 & n18690 ;
  assign n18692 = ~n266 & n18691 ;
  assign n18696 = ~n60 & n4902 ;
  assign n18697 = n60 & n18696 ;
  assign n18693 = n538 | n576 ;
  assign n18694 = n538 & ~n18693 ;
  assign n18695 = n6753 | n18694 ;
  assign n18698 = n18697 ^ n18695 ^ 1'b0 ;
  assign n18699 = n18698 ^ n2629 ^ 1'b0 ;
  assign n18700 = n18692 & n18699 ;
  assign n18701 = n1426 & ~n5362 ;
  assign n18702 = ~n1426 & n18701 ;
  assign n18703 = n18702 ^ n43 ^ 1'b0 ;
  assign n18704 = n18703 ^ n2403 ^ 1'b0 ;
  assign n18705 = n18700 & n18704 ;
  assign n18706 = ~n18683 & n18705 ;
  assign n18707 = ~n547 & n6575 ;
  assign n18708 = n18706 & n18707 ;
  assign n18667 = x2 & ~n180 ;
  assign n18668 = n180 & n18667 ;
  assign n18669 = n481 | n18668 ;
  assign n18670 = n481 & ~n18669 ;
  assign n18671 = n361 & n18670 ;
  assign n18672 = ~n4909 & n18671 ;
  assign n18673 = n4909 & n18672 ;
  assign n18709 = n18708 ^ n18673 ^ 1'b0 ;
  assign n18710 = ~n2005 & n18709 ;
  assign n18711 = n5418 ^ x6 ^ 1'b0 ;
  assign n18712 = ( ~n527 & n4602 ) | ( ~n527 & n18711 ) | ( n4602 & n18711 ) ;
  assign n18713 = ~n216 & n5301 ;
  assign n18714 = n18713 ^ n11429 ^ 1'b0 ;
  assign n18715 = n2450 & ~n4820 ;
  assign n18716 = n18714 & n18715 ;
  assign n18717 = n963 & ~n13766 ;
  assign n18718 = ~n8674 & n12232 ;
  assign n18719 = n18718 ^ n12436 ^ 1'b0 ;
  assign n18720 = n6133 & ~n10879 ;
  assign n18721 = n5528 ^ n3292 ^ 1'b0 ;
  assign n18722 = n18721 ^ n18290 ^ 1'b0 ;
  assign n18723 = n3960 | n6661 ;
  assign n18724 = n1323 | n18723 ;
  assign n18725 = n18724 ^ n12400 ^ 1'b0 ;
  assign n18726 = ~n2362 & n4254 ;
  assign n18727 = n18725 & n18726 ;
  assign n18728 = n3713 ^ n3037 ^ 1'b0 ;
  assign n18729 = ~n6376 & n18728 ;
  assign n18730 = ~n8201 & n18729 ;
  assign n18731 = n8819 & n18730 ;
  assign n18732 = n6636 | n18731 ;
  assign n18733 = n18732 ^ n8829 ^ 1'b0 ;
  assign n18734 = n841 | n4041 ;
  assign n18735 = n15042 ^ n3360 ^ 1'b0 ;
  assign n18736 = ~n18734 & n18735 ;
  assign n18737 = n18736 ^ n4983 ^ 1'b0 ;
  assign n18738 = n1475 & n18737 ;
  assign n18739 = n1203 & ~n9905 ;
  assign n18740 = n16044 ^ n1556 ^ 1'b0 ;
  assign n18741 = ~n11490 & n14551 ;
  assign n18748 = n7980 & n10751 ;
  assign n18742 = n552 & ~n2222 ;
  assign n18743 = n18742 ^ n16440 ^ 1'b0 ;
  assign n18744 = ~n6251 & n18743 ;
  assign n18745 = n18744 ^ n1192 ^ 1'b0 ;
  assign n18746 = ~n4541 & n18745 ;
  assign n18747 = ~n3449 & n18746 ;
  assign n18749 = n18748 ^ n18747 ^ 1'b0 ;
  assign n18750 = n7884 | n17190 ;
  assign n18751 = n18750 ^ n499 ^ 1'b0 ;
  assign n18752 = n3561 & ~n5126 ;
  assign n18753 = n18752 ^ n2733 ^ 1'b0 ;
  assign n18754 = n17507 ^ n5326 ^ 1'b0 ;
  assign n18755 = n4482 & ~n18754 ;
  assign n18756 = n11803 ^ n7497 ^ n4782 ;
  assign n18757 = n495 & ~n5639 ;
  assign n18758 = ~n5317 & n18757 ;
  assign n18759 = n13435 & n18758 ;
  assign n18760 = ~n3270 & n4549 ;
  assign n18761 = n18760 ^ n2446 ^ 1'b0 ;
  assign n18762 = n18570 & n18761 ;
  assign n18763 = n3493 & ~n12220 ;
  assign n18764 = n7130 ^ n880 ^ 1'b0 ;
  assign n18765 = n3019 & ~n18764 ;
  assign n18766 = ~n11056 & n18765 ;
  assign n18767 = n14800 ^ n8271 ^ 1'b0 ;
  assign n18768 = n5506 & n5688 ;
  assign n18769 = ~n1748 & n18768 ;
  assign n18770 = n5733 ^ n3659 ^ 1'b0 ;
  assign n18771 = n18769 | n18770 ;
  assign n18772 = n2728 ^ n520 ^ 1'b0 ;
  assign n18773 = n10032 & ~n18772 ;
  assign n18774 = n18773 ^ n15129 ^ 1'b0 ;
  assign n18775 = ~n18771 & n18774 ;
  assign n18776 = n18775 ^ n9657 ^ 1'b0 ;
  assign n18777 = n18776 ^ n5180 ^ 1'b0 ;
  assign n18778 = n8689 ^ n5302 ^ 1'b0 ;
  assign n18780 = n159 & n4595 ;
  assign n18781 = ~n3452 & n6291 ;
  assign n18782 = ~n18780 & n18781 ;
  assign n18779 = ~n2792 & n7908 ;
  assign n18783 = n18782 ^ n18779 ^ 1'b0 ;
  assign n18784 = ~n4227 & n5986 ;
  assign n18785 = ~n3844 & n18784 ;
  assign n18786 = n3414 & n5244 ;
  assign n18788 = n951 | n1798 ;
  assign n18787 = ~n6322 & n11278 ;
  assign n18789 = n18788 ^ n18787 ^ 1'b0 ;
  assign n18790 = n4015 ^ n2975 ^ 1'b0 ;
  assign n18791 = ~n3373 & n16731 ;
  assign n18792 = n439 | n13828 ;
  assign n18793 = n1162 | n12351 ;
  assign n18794 = ~n2649 & n6981 ;
  assign n18795 = n12207 & n18794 ;
  assign n18796 = ~n4495 & n7675 ;
  assign n18797 = ~n472 & n18796 ;
  assign n18798 = n18797 ^ n4803 ^ 1'b0 ;
  assign n18799 = n3226 & ~n6878 ;
  assign n18800 = n18799 ^ n2767 ^ 1'b0 ;
  assign n18801 = n7862 | n14852 ;
  assign n18802 = n16424 | n18801 ;
  assign n18803 = n16202 ^ n11742 ^ n4875 ;
  assign n18804 = n10221 ^ n5363 ^ 1'b0 ;
  assign n18805 = x9 | n5310 ;
  assign n18806 = n1455 & ~n16755 ;
  assign n18807 = n18806 ^ n9146 ^ 1'b0 ;
  assign n18808 = ( n1441 & n18305 ) | ( n1441 & n18807 ) | ( n18305 & n18807 ) ;
  assign n18809 = n16969 ^ n10751 ^ n9114 ;
  assign n18810 = n13061 ^ n1134 ^ 1'b0 ;
  assign n18811 = n3074 & ~n18810 ;
  assign n18812 = n8792 ^ n332 ^ 1'b0 ;
  assign n18813 = n18811 & ~n18812 ;
  assign n18814 = n18813 ^ n11334 ^ 1'b0 ;
  assign n18815 = n809 & ~n15129 ;
  assign n18816 = ~n5910 & n18815 ;
  assign n18817 = n18816 ^ n9978 ^ 1'b0 ;
  assign n18818 = ~n11462 & n18817 ;
  assign n18821 = n6260 ^ n2577 ^ 1'b0 ;
  assign n18819 = n4327 & ~n10787 ;
  assign n18820 = ~n12488 & n18819 ;
  assign n18822 = n18821 ^ n18820 ^ 1'b0 ;
  assign n18823 = n1615 & n13532 ;
  assign n18824 = n7675 & n18823 ;
  assign n18825 = n974 | n4361 ;
  assign n18826 = n18825 ^ n5182 ^ 1'b0 ;
  assign n18827 = n5853 ^ n1467 ^ 1'b0 ;
  assign n18828 = n8411 & ~n18827 ;
  assign n18829 = n18516 & n18828 ;
  assign n18830 = n18826 & n18829 ;
  assign n18831 = n3567 | n17169 ;
  assign n18832 = ~n18830 & n18831 ;
  assign n18833 = n18370 ^ n2105 ^ 1'b0 ;
  assign n18835 = n14877 ^ n10124 ^ 1'b0 ;
  assign n18834 = n9910 & ~n18113 ;
  assign n18836 = n18835 ^ n18834 ^ 1'b0 ;
  assign n18837 = n5501 & ~n18836 ;
  assign n18838 = n5973 & n18837 ;
  assign n18839 = n2497 & n14622 ;
  assign n18840 = ~n1840 & n18839 ;
  assign n18841 = n18840 ^ n1533 ^ 1'b0 ;
  assign n18842 = ~n2371 & n15238 ;
  assign n18843 = n4241 & ~n6094 ;
  assign n18846 = n1314 ^ n87 ^ 1'b0 ;
  assign n18847 = n12040 | n18846 ;
  assign n18844 = n11120 & ~n11865 ;
  assign n18845 = n18844 ^ n13585 ^ 1'b0 ;
  assign n18848 = n18847 ^ n18845 ^ 1'b0 ;
  assign n18849 = n2107 & ~n10378 ;
  assign n18850 = n18849 ^ n5148 ^ 1'b0 ;
  assign n18851 = ( n5237 & n6469 ) | ( n5237 & ~n11645 ) | ( n6469 & ~n11645 ) ;
  assign n18852 = ~n283 & n2613 ;
  assign n18853 = n13806 ^ n10180 ^ 1'b0 ;
  assign n18854 = n18853 ^ n15703 ^ 1'b0 ;
  assign n18855 = n634 & n18854 ;
  assign n18857 = n10525 ^ n6954 ^ 1'b0 ;
  assign n18858 = n17337 & n18857 ;
  assign n18856 = n269 & ~n11705 ;
  assign n18859 = n18858 ^ n18856 ^ n9035 ;
  assign n18860 = n10537 ^ n3992 ^ 1'b0 ;
  assign n18861 = n11622 | n18860 ;
  assign n18862 = n2712 & n18861 ;
  assign n18863 = n10523 ^ n6272 ^ 1'b0 ;
  assign n18865 = n18099 ^ n15089 ^ n218 ;
  assign n18864 = n1668 & ~n15604 ;
  assign n18866 = n18865 ^ n18864 ^ 1'b0 ;
  assign n18867 = ( n14819 & n18376 ) | ( n14819 & ~n18592 ) | ( n18376 & ~n18592 ) ;
  assign n18868 = n475 | n11233 ;
  assign n18869 = n3260 & ~n7236 ;
  assign n18870 = n18869 ^ n11491 ^ 1'b0 ;
  assign n18871 = n18870 ^ n2477 ^ 1'b0 ;
  assign n18872 = n2065 & ~n13067 ;
  assign n18873 = n18872 ^ n690 ^ 1'b0 ;
  assign n18874 = n1842 & ~n17723 ;
  assign n18876 = ~n8277 & n16656 ;
  assign n18875 = n3423 & n9599 ;
  assign n18877 = n18876 ^ n18875 ^ 1'b0 ;
  assign n18878 = n18874 & n18877 ;
  assign n18879 = n177 | n14422 ;
  assign n18880 = n18878 | n18879 ;
  assign n18881 = n6159 & ~n8838 ;
  assign n18882 = n18881 ^ n10190 ^ 1'b0 ;
  assign n18883 = n12225 & n18882 ;
  assign n18884 = n2439 & n3452 ;
  assign n18885 = n10184 ^ n7497 ^ 1'b0 ;
  assign n18886 = n8279 ^ n7095 ^ n1441 ;
  assign n18887 = n5304 | n18886 ;
  assign n18888 = n8406 & ~n18887 ;
  assign n18889 = n12898 ^ n5463 ^ 1'b0 ;
  assign n18890 = ~n4990 & n18889 ;
  assign n18891 = ~n10359 & n18890 ;
  assign n18892 = n1010 & ~n14476 ;
  assign n18893 = ~n113 & n10829 ;
  assign n18894 = n13974 | n14240 ;
  assign n18895 = n1995 ^ n633 ^ 1'b0 ;
  assign n18896 = ~n16175 & n18895 ;
  assign n18897 = n3827 | n7880 ;
  assign n18898 = n18897 ^ n1945 ^ 1'b0 ;
  assign n18899 = n18896 & ~n18898 ;
  assign n18900 = n517 & n628 ;
  assign n18901 = n254 & n1165 ;
  assign n18902 = ~n1165 & n18901 ;
  assign n18903 = n18900 & n18902 ;
  assign n18904 = n2739 & ~n18903 ;
  assign n18905 = n18903 & n18904 ;
  assign n18906 = n18905 ^ n2484 ^ 1'b0 ;
  assign n18907 = n16262 & n18906 ;
  assign n18908 = ~n18906 & n18907 ;
  assign n18909 = ~n1906 & n4314 ;
  assign n18910 = n191 | n18909 ;
  assign n18911 = n3887 | n12299 ;
  assign n18912 = n18911 ^ n2120 ^ 1'b0 ;
  assign n18913 = ~n2696 & n8253 ;
  assign n18914 = ~n18912 & n18913 ;
  assign n18915 = n2541 & n18914 ;
  assign n18916 = n6776 ^ n3546 ^ 1'b0 ;
  assign n18917 = ~n3732 & n18916 ;
  assign n18918 = n18917 ^ n7954 ^ 1'b0 ;
  assign n18919 = n2424 & n5947 ;
  assign n18920 = ~n158 & n2964 ;
  assign n18921 = n18920 ^ n4357 ^ 1'b0 ;
  assign n18922 = n4197 | n6769 ;
  assign n18923 = n18922 ^ n2155 ^ 1'b0 ;
  assign n18924 = n18923 ^ n11861 ^ 1'b0 ;
  assign n18925 = ~n18921 & n18924 ;
  assign n18926 = n5507 | n7668 ;
  assign n18927 = n10470 & ~n18926 ;
  assign n18928 = n935 | n3355 ;
  assign n18929 = n18928 ^ n142 ^ 1'b0 ;
  assign n18930 = ~n18927 & n18929 ;
  assign n18931 = n161 & n613 ;
  assign n18932 = ~n666 & n18931 ;
  assign n18933 = n2023 | n18932 ;
  assign n18934 = n18933 ^ n11707 ^ 1'b0 ;
  assign n18935 = n15509 | n18934 ;
  assign n18936 = n5401 | n13016 ;
  assign n18937 = n10692 ^ n3552 ^ 1'b0 ;
  assign n18938 = n6718 ^ n1052 ^ 1'b0 ;
  assign n18939 = ~n139 & n18938 ;
  assign n18940 = n7930 ^ n2165 ^ 1'b0 ;
  assign n18941 = n18769 ^ n861 ^ 1'b0 ;
  assign n18942 = n18940 & ~n18941 ;
  assign n18943 = n2097 | n3407 ;
  assign n18944 = n18943 ^ n3084 ^ 1'b0 ;
  assign n18945 = ( n6194 & n18942 ) | ( n6194 & n18944 ) | ( n18942 & n18944 ) ;
  assign n18946 = n7669 & n18945 ;
  assign n18947 = n6919 & n18946 ;
  assign n18948 = n1226 ^ n43 ^ 1'b0 ;
  assign n18949 = ~n4918 & n18948 ;
  assign n18950 = ( n2406 & ~n2900 ) | ( n2406 & n18949 ) | ( ~n2900 & n18949 ) ;
  assign n18951 = n17802 | n18950 ;
  assign n18952 = n257 & n14179 ;
  assign n18953 = n18952 ^ n4368 ^ 1'b0 ;
  assign n18954 = n105 & ~n18953 ;
  assign n18955 = n18954 ^ n46 ^ 1'b0 ;
  assign n18956 = n14870 ^ n8973 ^ 1'b0 ;
  assign n18957 = n18956 ^ n16680 ^ 1'b0 ;
  assign n18958 = ~n18955 & n18957 ;
  assign n18959 = n17320 ^ n10930 ^ 1'b0 ;
  assign n18960 = n16803 | n18959 ;
  assign n18963 = n2964 & ~n9424 ;
  assign n18961 = n3946 ^ n2360 ^ n1991 ;
  assign n18962 = n18961 ^ n3356 ^ 1'b0 ;
  assign n18964 = n18963 ^ n18962 ^ 1'b0 ;
  assign n18965 = n8392 | n18964 ;
  assign n18966 = n5506 ^ n2661 ^ 1'b0 ;
  assign n18967 = n7717 & n18966 ;
  assign n18968 = n18967 ^ n1426 ^ 1'b0 ;
  assign n18969 = n10021 ^ n8956 ^ 1'b0 ;
  assign n18970 = n86 | n18969 ;
  assign n18971 = n18970 ^ n12291 ^ 1'b0 ;
  assign n18972 = n15015 ^ n910 ^ 1'b0 ;
  assign n18973 = n1597 | n18972 ;
  assign n18974 = n18120 ^ n1358 ^ 1'b0 ;
  assign n18975 = n13038 & ~n18974 ;
  assign n18976 = n18975 ^ n7641 ^ 1'b0 ;
  assign n18977 = n3873 ^ n2331 ^ 1'b0 ;
  assign n18978 = ~n732 & n9227 ;
  assign n18979 = n18978 ^ n3264 ^ 1'b0 ;
  assign n18980 = n588 & n8751 ;
  assign n18981 = n18980 ^ n6427 ^ 1'b0 ;
  assign n18982 = n6385 | n18981 ;
  assign n18983 = n18982 ^ n13612 ^ 1'b0 ;
  assign n18987 = n602 | n1782 ;
  assign n18988 = n1782 & ~n18987 ;
  assign n18989 = n18988 ^ n18876 ^ 1'b0 ;
  assign n18984 = ~n1392 & n10635 ;
  assign n18985 = ~n10635 & n18984 ;
  assign n18986 = n11261 & ~n18985 ;
  assign n18990 = n18989 ^ n18986 ^ 1'b0 ;
  assign n18995 = n890 ^ n323 ^ 1'b0 ;
  assign n18991 = n4358 & n7892 ;
  assign n18992 = n615 | n13015 ;
  assign n18993 = n18991 | n18992 ;
  assign n18994 = n333 & n18993 ;
  assign n18996 = n18995 ^ n18994 ^ 1'b0 ;
  assign n18997 = n6081 ^ n1388 ^ 1'b0 ;
  assign n18998 = n9666 ^ n5774 ^ 1'b0 ;
  assign n18999 = n247 & n18998 ;
  assign n19000 = n8601 & n18999 ;
  assign n19001 = n7585 & n13899 ;
  assign n19002 = n11709 & n19001 ;
  assign n19003 = n12857 | n19002 ;
  assign n19004 = n1726 ^ n741 ^ 1'b0 ;
  assign n19005 = ~n252 & n19004 ;
  assign n19006 = n833 | n6385 ;
  assign n19007 = n17471 & ~n19006 ;
  assign n19008 = ~n11842 & n15033 ;
  assign n19009 = n7555 | n19008 ;
  assign n19010 = n3939 & ~n8173 ;
  assign n19011 = n9292 ^ n2865 ^ 1'b0 ;
  assign n19012 = n11413 ^ n1342 ^ 1'b0 ;
  assign n19013 = n3567 ^ n2461 ^ 1'b0 ;
  assign n19014 = n19013 ^ n748 ^ 1'b0 ;
  assign n19015 = n8114 & ~n19014 ;
  assign n19016 = n3535 | n17068 ;
  assign n19017 = ~n11002 & n14992 ;
  assign n19018 = n2618 & n19017 ;
  assign n19019 = ~n2618 & n19018 ;
  assign n19020 = ( n114 & ~n3576 ) | ( n114 & n9292 ) | ( ~n3576 & n9292 ) ;
  assign n19021 = n19020 ^ n17700 ^ 1'b0 ;
  assign n19022 = n5251 | n19021 ;
  assign n19023 = n6174 ^ n2882 ^ n290 ;
  assign n19024 = ~n19022 & n19023 ;
  assign n19025 = n9983 ^ n2519 ^ 1'b0 ;
  assign n19026 = n18778 ^ n2314 ^ 1'b0 ;
  assign n19033 = n10470 ^ n1555 ^ 1'b0 ;
  assign n19030 = ~n10421 & n16931 ;
  assign n19031 = n19030 ^ n11682 ^ 1'b0 ;
  assign n19027 = n18798 ^ n4917 ^ 1'b0 ;
  assign n19028 = n938 & n19027 ;
  assign n19029 = ~n4349 & n19028 ;
  assign n19032 = n19031 ^ n19029 ^ 1'b0 ;
  assign n19034 = n19033 ^ n19032 ^ 1'b0 ;
  assign n19038 = n4823 ^ n2635 ^ 1'b0 ;
  assign n19035 = n2201 ^ n645 ^ 1'b0 ;
  assign n19036 = n1360 | n19035 ;
  assign n19037 = ~n6378 & n19036 ;
  assign n19039 = n19038 ^ n19037 ^ 1'b0 ;
  assign n19040 = ~n2751 & n2874 ;
  assign n19041 = n5014 & n7051 ;
  assign n19042 = n3507 ^ n1933 ^ 1'b0 ;
  assign n19043 = n19042 ^ n17196 ^ 1'b0 ;
  assign n19044 = n5267 & ~n19043 ;
  assign n19047 = n9096 & n16158 ;
  assign n19045 = n3137 ^ n2984 ^ 1'b0 ;
  assign n19046 = n975 & n19045 ;
  assign n19048 = n19047 ^ n19046 ^ 1'b0 ;
  assign n19049 = ( n2122 & n11061 ) | ( n2122 & ~n19048 ) | ( n11061 & ~n19048 ) ;
  assign n19050 = n19049 ^ n1345 ^ 1'b0 ;
  assign n19051 = ~n19 & n13813 ;
  assign n19052 = n19051 ^ n11080 ^ 1'b0 ;
  assign n19053 = n281 & n19052 ;
  assign n19054 = n205 & ~n741 ;
  assign n19055 = n19054 ^ n12222 ^ 1'b0 ;
  assign n19057 = n5314 ^ n3120 ^ 1'b0 ;
  assign n19058 = n9131 & n19057 ;
  assign n19056 = n14062 & ~n17603 ;
  assign n19059 = n19058 ^ n19056 ^ 1'b0 ;
  assign n19060 = n19055 & ~n19059 ;
  assign n19063 = ~n2577 & n4746 ;
  assign n19064 = n2217 & n19063 ;
  assign n19061 = ~n5892 & n14102 ;
  assign n19062 = n19061 ^ n16289 ^ 1'b0 ;
  assign n19065 = n19064 ^ n19062 ^ 1'b0 ;
  assign n19066 = n19060 & n19065 ;
  assign n19067 = n3514 & n16691 ;
  assign n19068 = ~n9775 & n19067 ;
  assign n19069 = ~n2790 & n19068 ;
  assign n19070 = n3959 & ~n10873 ;
  assign n19071 = n9306 | n19070 ;
  assign n19072 = n3437 | n19071 ;
  assign n19073 = n5681 & n19072 ;
  assign n19074 = n19073 ^ n17618 ^ 1'b0 ;
  assign n19075 = n2604 & ~n19074 ;
  assign n19076 = n375 | n2233 ;
  assign n19077 = n19076 ^ n16646 ^ 1'b0 ;
  assign n19078 = n2980 & ~n13430 ;
  assign n19079 = n520 & n19078 ;
  assign n19080 = n7497 & n19079 ;
  assign n19081 = ~n4618 & n17707 ;
  assign n19082 = n3423 ^ n1023 ^ 1'b0 ;
  assign n19083 = n364 & ~n679 ;
  assign n19084 = n5957 ^ n1827 ^ 1'b0 ;
  assign n19085 = n749 & ~n19084 ;
  assign n19086 = n19085 ^ n535 ^ 1'b0 ;
  assign n19087 = n19083 & n19086 ;
  assign n19088 = ~n2005 & n11502 ;
  assign n19089 = n6562 | n19088 ;
  assign n19090 = n6562 & ~n19089 ;
  assign n19091 = n10012 ^ n3971 ^ 1'b0 ;
  assign n19092 = n16552 & n16753 ;
  assign n19093 = n9811 ^ n1831 ^ 1'b0 ;
  assign n19094 = n9785 | n19093 ;
  assign n19095 = ~n3767 & n19094 ;
  assign n19096 = n180 ^ n149 ^ 1'b0 ;
  assign n19097 = n3327 ^ n1584 ^ 1'b0 ;
  assign n19103 = n5756 & ~n11338 ;
  assign n19104 = n12073 & n19103 ;
  assign n19100 = n2252 & n2604 ;
  assign n19101 = n5890 & n19100 ;
  assign n19098 = ~n5016 & n9307 ;
  assign n19099 = n19098 ^ n1127 ^ 1'b0 ;
  assign n19102 = n19101 ^ n19099 ^ n12982 ;
  assign n19105 = n19104 ^ n19102 ^ n10911 ;
  assign n19106 = n12299 ^ n3287 ^ 1'b0 ;
  assign n19107 = n2566 & ~n3304 ;
  assign n19108 = ~n19106 & n19107 ;
  assign n19109 = n19108 ^ n10245 ^ 1'b0 ;
  assign n19110 = n16577 | n17356 ;
  assign n19111 = n6897 ^ n2011 ^ 1'b0 ;
  assign n19112 = n1369 ^ n208 ^ 1'b0 ;
  assign n19113 = n8108 & ~n19112 ;
  assign n19114 = n7108 & n10728 ;
  assign n19115 = n19114 ^ n18975 ^ n5030 ;
  assign n19116 = n16977 ^ n3826 ^ 1'b0 ;
  assign n19117 = n5434 | n9166 ;
  assign n19118 = n19117 ^ n271 ^ 1'b0 ;
  assign n19119 = n2927 & n19118 ;
  assign n19120 = n19119 ^ n423 ^ 1'b0 ;
  assign n19121 = ~n294 & n13660 ;
  assign n19122 = n7419 ^ n4210 ^ 1'b0 ;
  assign n19123 = n1835 | n6440 ;
  assign n19124 = n19123 ^ n907 ^ 1'b0 ;
  assign n19125 = n2104 & n4586 ;
  assign n19126 = n19125 ^ n4033 ^ 1'b0 ;
  assign n19127 = n3985 | n4939 ;
  assign n19128 = n1506 | n3855 ;
  assign n19129 = n4867 ^ n375 ^ 1'b0 ;
  assign n19130 = ~n2454 & n19129 ;
  assign n19131 = n8108 & n19130 ;
  assign n19132 = n19128 | n19131 ;
  assign n19133 = n9210 | n19132 ;
  assign n19134 = n19133 ^ n13966 ^ 1'b0 ;
  assign n19135 = ~n19127 & n19134 ;
  assign n19136 = ~n3539 & n7642 ;
  assign n19137 = n1432 ^ n116 ^ 1'b0 ;
  assign n19138 = ~n3939 & n5613 ;
  assign n19139 = n19138 ^ n15330 ^ 1'b0 ;
  assign n19140 = n4133 & ~n19139 ;
  assign n19141 = n5862 & n10024 ;
  assign n19142 = n5202 & ~n16770 ;
  assign n19143 = n4873 ^ n284 ^ 1'b0 ;
  assign n19144 = ~n8276 & n9022 ;
  assign n19145 = n17266 ^ n3101 ^ 1'b0 ;
  assign n19146 = n19144 & ~n19145 ;
  assign n19147 = ~n5697 & n8504 ;
  assign n19148 = n19147 ^ n3091 ^ 1'b0 ;
  assign n19149 = n14448 & n19148 ;
  assign n19150 = n3753 & n5041 ;
  assign n19151 = n748 & ~n2784 ;
  assign n19152 = n11168 ^ n343 ^ 1'b0 ;
  assign n19153 = n12922 & ~n19152 ;
  assign n19154 = n12961 & n19153 ;
  assign n19155 = n1951 & n19154 ;
  assign n19156 = n13027 ^ n2710 ^ 1'b0 ;
  assign n19157 = ~n2075 & n2106 ;
  assign n19158 = n19157 ^ n1441 ^ 1'b0 ;
  assign n19159 = n6571 | n14848 ;
  assign n19160 = n18508 | n19159 ;
  assign n19161 = n11931 ^ n4623 ^ 1'b0 ;
  assign n19162 = n8620 | n10958 ;
  assign n19163 = n19162 ^ n3577 ^ 1'b0 ;
  assign n19164 = n17383 ^ n10658 ^ 1'b0 ;
  assign n19165 = n19163 & ~n19164 ;
  assign n19166 = n2047 & ~n7263 ;
  assign n19167 = n15288 | n19166 ;
  assign n19168 = n4654 ^ n2987 ^ 1'b0 ;
  assign n19169 = n2460 & n19168 ;
  assign n19170 = ~n461 & n9191 ;
  assign n19171 = n1974 & n19170 ;
  assign n19172 = n18595 | n19171 ;
  assign n19173 = n14059 ^ n3580 ^ 1'b0 ;
  assign n19174 = n553 & n7205 ;
  assign n19175 = n19174 ^ n1359 ^ 1'b0 ;
  assign n19176 = n19175 ^ n14094 ^ 1'b0 ;
  assign n19177 = n8863 ^ n97 ^ 1'b0 ;
  assign n19178 = n677 & n19177 ;
  assign n19179 = n3522 & n19178 ;
  assign n19180 = n19176 | n19179 ;
  assign n19181 = n19180 ^ n7071 ^ 1'b0 ;
  assign n19182 = n19181 ^ n4075 ^ 1'b0 ;
  assign n19183 = n5011 | n14400 ;
  assign n19184 = ( n191 & n1463 ) | ( n191 & ~n3550 ) | ( n1463 & ~n3550 ) ;
  assign n19185 = n14822 & ~n19184 ;
  assign n19186 = n216 | n235 ;
  assign n19187 = n216 | n1671 ;
  assign n19188 = n2955 | n4070 ;
  assign n19189 = n1463 & ~n10618 ;
  assign n19190 = ~n19188 & n19189 ;
  assign n19191 = n4728 & ~n19190 ;
  assign n19192 = n13532 & n19191 ;
  assign n19193 = n15081 & ~n19192 ;
  assign n19195 = n2105 | n9561 ;
  assign n19196 = n19195 ^ n4475 ^ 1'b0 ;
  assign n19194 = n435 & n7668 ;
  assign n19197 = n19196 ^ n19194 ^ 1'b0 ;
  assign n19198 = n9431 ^ n119 ^ 1'b0 ;
  assign n19199 = ~n1720 & n14608 ;
  assign n19200 = n120 & n19199 ;
  assign n19201 = n6230 | n19200 ;
  assign n19202 = n8764 & ~n19201 ;
  assign n19203 = n19202 ^ n702 ^ 1'b0 ;
  assign n19204 = ~n19198 & n19203 ;
  assign n19205 = n10544 & n15543 ;
  assign n19206 = n10971 ^ n6005 ^ 1'b0 ;
  assign n19207 = ~n5502 & n19206 ;
  assign n19209 = n8013 ^ n2542 ^ 1'b0 ;
  assign n19210 = n258 & ~n19209 ;
  assign n19208 = ~n9567 & n11494 ;
  assign n19211 = n19210 ^ n19208 ^ 1'b0 ;
  assign n19212 = n19211 ^ n3851 ^ n2252 ;
  assign n19213 = n5905 & ~n19212 ;
  assign n19214 = n9491 ^ n7301 ^ 1'b0 ;
  assign n19215 = n4864 | n19214 ;
  assign n19216 = n9279 & n18379 ;
  assign n19217 = n19216 ^ n10239 ^ 1'b0 ;
  assign n19218 = n2086 ^ n934 ^ 1'b0 ;
  assign n19219 = ~n3216 & n19218 ;
  assign n19220 = ~n965 & n14684 ;
  assign n19221 = n965 & n19220 ;
  assign n19222 = n73 & ~n19221 ;
  assign n19223 = n19222 ^ n2072 ^ 1'b0 ;
  assign n19224 = n2238 & n10216 ;
  assign n19225 = n3280 ^ n3249 ^ 1'b0 ;
  assign n19226 = n13206 ^ n1304 ^ 1'b0 ;
  assign n19227 = n19225 | n19226 ;
  assign n19228 = n19227 ^ n9750 ^ 1'b0 ;
  assign n19229 = n3042 | n6876 ;
  assign n19230 = n13150 ^ n11597 ^ 1'b0 ;
  assign n19231 = n19229 & n19230 ;
  assign n19232 = n2655 & ~n7657 ;
  assign n19233 = n19232 ^ n14181 ^ 1'b0 ;
  assign n19234 = n9649 ^ n4575 ^ 1'b0 ;
  assign n19235 = n18729 ^ n3221 ^ 1'b0 ;
  assign n19236 = ~n6156 & n19235 ;
  assign n19237 = n5260 & ~n10544 ;
  assign n19238 = n12455 ^ n10676 ^ 1'b0 ;
  assign n19239 = ( n2067 & n13747 ) | ( n2067 & ~n19238 ) | ( n13747 & ~n19238 ) ;
  assign n19240 = n1179 & n19239 ;
  assign n19242 = n10636 ^ n5799 ^ 1'b0 ;
  assign n19241 = ~n4495 & n7130 ;
  assign n19243 = n19242 ^ n19241 ^ 1'b0 ;
  assign n19244 = n14884 ^ n2360 ^ 1'b0 ;
  assign n19245 = ~n8915 & n19244 ;
  assign n19246 = n12049 | n19120 ;
  assign n19248 = n5024 & ~n9155 ;
  assign n19247 = n5698 & ~n9550 ;
  assign n19249 = n19248 ^ n19247 ^ 1'b0 ;
  assign n19250 = n963 | n5394 ;
  assign n19251 = n6150 & ~n8286 ;
  assign n19252 = n19250 & n19251 ;
  assign n19253 = n19252 ^ n9294 ^ 1'b0 ;
  assign n19254 = n19253 ^ n8834 ^ n328 ;
  assign n19255 = n14765 | n19254 ;
  assign n19256 = ~n6023 & n8104 ;
  assign n19257 = n19256 ^ n17920 ^ 1'b0 ;
  assign n19258 = n4322 | n19257 ;
  assign n19259 = n1080 & n10676 ;
  assign n19260 = ~n1531 & n19259 ;
  assign n19261 = n927 & n7857 ;
  assign n19262 = n281 & n2482 ;
  assign n19263 = n19262 ^ n2566 ^ 1'b0 ;
  assign n19264 = ~n495 & n19263 ;
  assign n19265 = n14608 ^ n12664 ^ 1'b0 ;
  assign n19266 = n13128 | n19265 ;
  assign n19267 = n832 & n4036 ;
  assign n19268 = ~n4036 & n19267 ;
  assign n19269 = n4684 & n19268 ;
  assign n19273 = n1085 & n1207 ;
  assign n19274 = ~n1085 & n19273 ;
  assign n19270 = ~n7435 & n9592 ;
  assign n19271 = n7435 & n19270 ;
  assign n19272 = n1026 | n19271 ;
  assign n19275 = n19274 ^ n19272 ^ 1'b0 ;
  assign n19276 = n15711 | n19275 ;
  assign n19277 = n378 & ~n664 ;
  assign n19278 = ~n378 & n19277 ;
  assign n19279 = n121 & ~n19278 ;
  assign n19280 = ~n121 & n19279 ;
  assign n19281 = n13035 ^ n5625 ^ 1'b0 ;
  assign n19282 = n19280 & n19281 ;
  assign n19283 = n8081 & n19282 ;
  assign n19284 = n19276 & n19283 ;
  assign n19285 = n19269 & ~n19284 ;
  assign n19286 = ~n404 & n17421 ;
  assign n19287 = n404 & n19286 ;
  assign n19288 = n19287 ^ n2961 ^ 1'b0 ;
  assign n19289 = n846 | n19288 ;
  assign n19290 = n19289 ^ n1660 ^ 1'b0 ;
  assign n19291 = n19290 ^ n18039 ^ 1'b0 ;
  assign n19292 = ~n19285 & n19291 ;
  assign n19293 = ~n18798 & n18886 ;
  assign n19294 = n4804 ^ n2420 ^ 1'b0 ;
  assign n19295 = n1149 & ~n19294 ;
  assign n19296 = n4349 & n19295 ;
  assign n19297 = n1227 & n4214 ;
  assign n19298 = n19297 ^ n4972 ^ 1'b0 ;
  assign n19299 = n19298 ^ n2270 ^ 1'b0 ;
  assign n19302 = n8099 ^ n4970 ^ 1'b0 ;
  assign n19303 = n15765 & n19302 ;
  assign n19304 = n1860 & n19303 ;
  assign n19305 = n704 | n19304 ;
  assign n19306 = n292 | n19305 ;
  assign n19300 = ~n405 & n13529 ;
  assign n19301 = n19300 ^ n8869 ^ 1'b0 ;
  assign n19307 = n19306 ^ n19301 ^ 1'b0 ;
  assign n19308 = n6589 & n8771 ;
  assign n19309 = ~n2921 & n19308 ;
  assign n19310 = n2558 & ~n19309 ;
  assign n19311 = n19310 ^ n15145 ^ 1'b0 ;
  assign n19312 = n19311 ^ n3098 ^ 1'b0 ;
  assign n19313 = ~n3869 & n6464 ;
  assign n19314 = n19313 ^ n1252 ^ 1'b0 ;
  assign n19315 = n1431 | n19314 ;
  assign n19316 = n5156 | n19315 ;
  assign n19317 = n6890 & ~n17531 ;
  assign n19318 = n19317 ^ n3355 ^ 1'b0 ;
  assign n19319 = n1072 | n14423 ;
  assign n19320 = n4889 ^ n1329 ^ 1'b0 ;
  assign n19321 = n5747 & n19320 ;
  assign n19322 = n5709 & n19321 ;
  assign n19323 = n19322 ^ n6365 ^ 1'b0 ;
  assign n19324 = n19323 ^ n16443 ^ 1'b0 ;
  assign n19325 = n931 & ~n19324 ;
  assign n19326 = n11460 ^ n917 ^ 1'b0 ;
  assign n19327 = n2364 & n19326 ;
  assign n19328 = n2680 & ~n19327 ;
  assign n19329 = n624 ^ n163 ^ 1'b0 ;
  assign n19330 = n3459 ^ n354 ^ 1'b0 ;
  assign n19331 = ~n5805 & n9629 ;
  assign n19332 = n19331 ^ n11656 ^ 1'b0 ;
  assign n19334 = n1148 | n3911 ;
  assign n19335 = n3911 & ~n19334 ;
  assign n19336 = n246 | n19335 ;
  assign n19337 = n246 & ~n19336 ;
  assign n19338 = n8552 | n19337 ;
  assign n19339 = n19337 & ~n19338 ;
  assign n19340 = n2007 & n19339 ;
  assign n19341 = n7410 | n19340 ;
  assign n19333 = n12223 ^ n6349 ^ 1'b0 ;
  assign n19342 = n19341 ^ n19333 ^ 1'b0 ;
  assign n19343 = ~n8609 & n19342 ;
  assign n19344 = n4357 & n19343 ;
  assign n19345 = n19344 ^ n15151 ^ 1'b0 ;
  assign n19347 = n4741 ^ n1169 ^ 1'b0 ;
  assign n19348 = ( n11586 & n18007 ) | ( n11586 & ~n19347 ) | ( n18007 & ~n19347 ) ;
  assign n19346 = n2573 & ~n7283 ;
  assign n19349 = n19348 ^ n19346 ^ 1'b0 ;
  assign n19350 = n6539 & n19349 ;
  assign n19351 = n3449 & n3862 ;
  assign n19352 = n18268 | n19351 ;
  assign n19353 = n17859 & ~n19352 ;
  assign n19354 = n234 & n19353 ;
  assign n19355 = n4314 ^ n4297 ^ 1'b0 ;
  assign n19356 = n5144 & ~n19355 ;
  assign n19357 = n5525 ^ n4037 ^ 1'b0 ;
  assign n19358 = n19356 & n19357 ;
  assign n19359 = ~n2295 & n19358 ;
  assign n19360 = n2726 ^ n1662 ^ 1'b0 ;
  assign n19361 = ~n3007 & n19360 ;
  assign n19362 = n1130 ^ n608 ^ 1'b0 ;
  assign n19363 = n13237 | n19362 ;
  assign n19364 = n19363 ^ n8495 ^ 1'b0 ;
  assign n19365 = n19364 ^ n2864 ^ 1'b0 ;
  assign n19366 = n11360 ^ n4531 ^ 1'b0 ;
  assign n19367 = n14321 | n19366 ;
  assign n19368 = n19367 ^ n13588 ^ 1'b0 ;
  assign n19369 = n4924 | n19368 ;
  assign n19370 = ~n3750 & n11033 ;
  assign n19371 = ( n321 & n5566 ) | ( n321 & n9889 ) | ( n5566 & n9889 ) ;
  assign n19372 = ~n14838 & n19371 ;
  assign n19373 = n8470 ^ n1929 ^ 1'b0 ;
  assign n19374 = n11272 & n19373 ;
  assign n19375 = n1433 ^ n1226 ^ 1'b0 ;
  assign n19376 = n17052 | n19375 ;
  assign n19377 = n5322 | n19376 ;
  assign n19378 = ~n4589 & n19377 ;
  assign n19379 = n1854 | n2036 ;
  assign n19380 = n19379 ^ n3739 ^ 1'b0 ;
  assign n19381 = n9506 & n19380 ;
  assign n19382 = n19381 ^ n3027 ^ 1'b0 ;
  assign n19383 = n8785 ^ n233 ^ 1'b0 ;
  assign n19384 = n7330 & ~n19383 ;
  assign n19385 = n19384 ^ n4840 ^ 1'b0 ;
  assign n19386 = n19382 | n19385 ;
  assign n19387 = n19386 ^ n3177 ^ 1'b0 ;
  assign n19388 = n4728 & ~n10158 ;
  assign n19389 = n12119 & ~n19388 ;
  assign n19390 = n3868 & n8657 ;
  assign n19391 = n295 | n19390 ;
  assign n19392 = n1730 & ~n4853 ;
  assign n19393 = n478 | n604 ;
  assign n19394 = n19393 ^ n495 ^ 1'b0 ;
  assign n19395 = n2193 & ~n2472 ;
  assign n19396 = n2472 & n19395 ;
  assign n19397 = n10025 | n19396 ;
  assign n19398 = n19396 & ~n19397 ;
  assign n19399 = n17119 & ~n18916 ;
  assign n19400 = n16906 ^ n16570 ^ n15933 ;
  assign n19401 = n11889 ^ n8082 ^ 1'b0 ;
  assign n19402 = ~n1982 & n15905 ;
  assign n19403 = n4063 & ~n17151 ;
  assign n19404 = n7136 ^ n83 ^ 1'b0 ;
  assign n19405 = n2456 & n6090 ;
  assign n19406 = n19405 ^ n817 ^ 1'b0 ;
  assign n19407 = ~n382 & n3335 ;
  assign n19408 = n19407 ^ n4505 ^ 1'b0 ;
  assign n19409 = n2179 & n7634 ;
  assign n19410 = ~n19408 & n19409 ;
  assign n19411 = n19410 ^ n5362 ^ 1'b0 ;
  assign n19412 = n2733 & n8907 ;
  assign n19413 = ~n40 & n19412 ;
  assign n19414 = n3329 | n19413 ;
  assign n19415 = n850 | n5185 ;
  assign n19416 = n1917 | n13258 ;
  assign n19417 = n18552 ^ n1271 ^ 1'b0 ;
  assign n19418 = n4455 | n5535 ;
  assign n19419 = n19418 ^ n4418 ^ 1'b0 ;
  assign n19420 = n1388 & ~n2437 ;
  assign n19421 = n10208 & n19420 ;
  assign n19422 = n12385 ^ n8893 ^ n764 ;
  assign n19423 = n19422 ^ n5603 ^ 1'b0 ;
  assign n19424 = n4055 | n19423 ;
  assign n19425 = n540 | n19424 ;
  assign n19426 = ~n1011 & n6160 ;
  assign n19427 = n19426 ^ n6571 ^ 1'b0 ;
  assign n19428 = ~n671 & n15219 ;
  assign n19429 = n13583 & n19428 ;
  assign n19430 = n450 & ~n4544 ;
  assign n19431 = n3049 & ~n10996 ;
  assign n19435 = ~n1660 & n1891 ;
  assign n19436 = n19435 ^ n3871 ^ 1'b0 ;
  assign n19432 = n8322 ^ n1472 ^ 1'b0 ;
  assign n19433 = ~n3293 & n19432 ;
  assign n19434 = n5952 & n19433 ;
  assign n19437 = n19436 ^ n19434 ^ 1'b0 ;
  assign n19438 = n310 & ~n3566 ;
  assign n19439 = n7384 | n7421 ;
  assign n19440 = n5657 | n11435 ;
  assign n19441 = n12688 & ~n19440 ;
  assign n19442 = n443 & n13253 ;
  assign n19443 = n3373 & n19442 ;
  assign n19444 = ( n183 & n2551 ) | ( n183 & n16501 ) | ( n2551 & n16501 ) ;
  assign n19445 = n2931 | n12519 ;
  assign n19446 = n1113 | n3112 ;
  assign n19447 = n6277 & ~n6327 ;
  assign n19448 = ~n2732 & n19447 ;
  assign n19449 = n19448 ^ n12048 ^ 1'b0 ;
  assign n19450 = n3219 & n19449 ;
  assign n19451 = ~n19446 & n19450 ;
  assign n19452 = n19451 ^ n1961 ^ 1'b0 ;
  assign n19453 = ~n4015 & n19452 ;
  assign n19454 = n458 | n13094 ;
  assign n19455 = n19454 ^ n5326 ^ 1'b0 ;
  assign n19456 = n157 & ~n19455 ;
  assign n19457 = n19456 ^ n16557 ^ 1'b0 ;
  assign n19458 = n8660 ^ n2566 ^ 1'b0 ;
  assign n19459 = n66 & ~n19458 ;
  assign n19460 = n19459 ^ n4906 ^ 1'b0 ;
  assign n19461 = n13966 & n19460 ;
  assign n19462 = ~n11041 & n19461 ;
  assign n19463 = n727 & n19462 ;
  assign n19464 = n16671 ^ n4923 ^ 1'b0 ;
  assign n19465 = n19464 ^ n9789 ^ 1'b0 ;
  assign n19466 = n205 | n19465 ;
  assign n19467 = n446 | n853 ;
  assign n19468 = n853 & ~n19467 ;
  assign n19469 = n388 & n1747 ;
  assign n19470 = n7594 & n19469 ;
  assign n19471 = ~n19469 & n19470 ;
  assign n19472 = ~n19468 & n19471 ;
  assign n19473 = n2254 | n19472 ;
  assign n19474 = n19472 & ~n19473 ;
  assign n19475 = n7604 ^ n2998 ^ n1355 ;
  assign n19476 = n7729 | n9625 ;
  assign n19477 = ~n2719 & n11802 ;
  assign n19478 = n19476 & n19477 ;
  assign n19479 = n8441 | n19478 ;
  assign n19480 = n861 & ~n16219 ;
  assign n19481 = n1668 & n5716 ;
  assign n19482 = n19481 ^ n3068 ^ 1'b0 ;
  assign n19483 = ~n7570 & n7697 ;
  assign n19484 = n19482 & n19483 ;
  assign n19485 = n905 ^ n501 ^ 1'b0 ;
  assign n19486 = n19485 ^ n149 ^ 1'b0 ;
  assign n19487 = n19486 ^ n432 ^ 1'b0 ;
  assign n19488 = n5331 | n19487 ;
  assign n19490 = ~n7312 & n12871 ;
  assign n19489 = n8279 & ~n8518 ;
  assign n19491 = n19490 ^ n19489 ^ 1'b0 ;
  assign n19492 = n18579 & n19491 ;
  assign n19493 = n1061 & ~n4075 ;
  assign n19496 = n6365 & ~n6942 ;
  assign n19497 = n19496 ^ n9184 ^ 1'b0 ;
  assign n19494 = n3584 & n7137 ;
  assign n19495 = n19494 ^ n4891 ^ 1'b0 ;
  assign n19498 = n19497 ^ n19495 ^ 1'b0 ;
  assign n19499 = n7661 ^ n3928 ^ 1'b0 ;
  assign n19500 = n1110 & ~n8696 ;
  assign n19501 = ~n13634 & n19500 ;
  assign n19502 = n19501 ^ n13586 ^ 1'b0 ;
  assign n19503 = n7849 ^ n1879 ^ 1'b0 ;
  assign n19508 = ~n7812 & n12875 ;
  assign n19505 = n1274 | n11111 ;
  assign n19504 = n148 & n6453 ;
  assign n19506 = n19505 ^ n19504 ^ 1'b0 ;
  assign n19507 = n5125 & n19506 ;
  assign n19509 = n19508 ^ n19507 ^ 1'b0 ;
  assign n19510 = n3219 | n14204 ;
  assign n19511 = n19510 ^ n5252 ^ 1'b0 ;
  assign n19512 = n10414 ^ n8223 ^ 1'b0 ;
  assign n19513 = n8422 & ~n14425 ;
  assign n19514 = n19513 ^ n17535 ^ 1'b0 ;
  assign n19515 = n1419 | n10303 ;
  assign n19516 = n2773 | n19515 ;
  assign n19517 = n7279 & n8326 ;
  assign n19518 = n19517 ^ n13079 ^ 1'b0 ;
  assign n19519 = n6880 ^ n3542 ^ 1'b0 ;
  assign n19520 = n4643 & n14226 ;
  assign n19521 = n19520 ^ n10201 ^ 1'b0 ;
  assign n19522 = ~n5685 & n11619 ;
  assign n19523 = n14806 ^ n1090 ^ 1'b0 ;
  assign n19524 = ~n2136 & n19523 ;
  assign n19526 = n17777 ^ n13026 ^ 1'b0 ;
  assign n19527 = ~n4267 & n19526 ;
  assign n19525 = n512 & n10064 ;
  assign n19528 = n19527 ^ n19525 ^ 1'b0 ;
  assign n19529 = n2303 | n19528 ;
  assign n19530 = n19403 | n19529 ;
  assign n19531 = n665 | n14537 ;
  assign n19532 = n7988 & ~n19531 ;
  assign n19533 = n408 & n12709 ;
  assign n19534 = n167 & n19533 ;
  assign n19535 = n1632 & n2633 ;
  assign n19536 = n8437 ^ n2659 ^ 1'b0 ;
  assign n19537 = n2101 & ~n19536 ;
  assign n19538 = n8614 ^ n3078 ^ 1'b0 ;
  assign n19539 = n10784 & n19538 ;
  assign n19540 = n8639 | n9346 ;
  assign n19541 = n10368 ^ n4361 ^ 1'b0 ;
  assign n19542 = n148 | n19541 ;
  assign n19543 = n70 | n274 ;
  assign n19544 = n1025 & ~n19543 ;
  assign n19545 = n19544 ^ n1642 ^ 1'b0 ;
  assign n19546 = n3196 & ~n19545 ;
  assign n19547 = n1057 & ~n19546 ;
  assign n19548 = n19547 ^ n3816 ^ 1'b0 ;
  assign n19549 = n19542 | n19548 ;
  assign n19550 = n2754 ^ n1354 ^ 1'b0 ;
  assign n19551 = n7183 | n11666 ;
  assign n19552 = n19551 ^ n1438 ^ 1'b0 ;
  assign n19553 = n15062 & ~n19552 ;
  assign n19554 = n512 & n7846 ;
  assign n19555 = n11965 ^ n1425 ^ 1'b0 ;
  assign n19556 = n1668 & n9723 ;
  assign n19557 = n2082 & n19556 ;
  assign n19558 = n18453 ^ n3359 ^ 1'b0 ;
  assign n19559 = n12317 & ~n19558 ;
  assign n19560 = n19559 ^ n642 ^ 1'b0 ;
  assign n19561 = n4373 ^ n254 ^ 1'b0 ;
  assign n19562 = n1592 ^ n622 ^ 1'b0 ;
  assign n19563 = n19562 ^ n16782 ^ 1'b0 ;
  assign n19564 = n7564 | n10520 ;
  assign n19565 = n1284 & n19564 ;
  assign n19566 = n6432 & ~n19565 ;
  assign n19567 = n19566 ^ n8461 ^ 1'b0 ;
  assign n19568 = ~n55 & n2151 ;
  assign n19569 = ~n4545 & n19568 ;
  assign n19570 = n19569 ^ n19055 ^ 1'b0 ;
  assign n19571 = n3405 | n13748 ;
  assign n19572 = n17697 & ~n19571 ;
  assign n19573 = n19572 ^ n14155 ^ n9244 ;
  assign n19574 = ~n769 & n7221 ;
  assign n19575 = n908 & ~n2014 ;
  assign n19576 = n15553 ^ n1523 ^ 1'b0 ;
  assign n19577 = n3483 ^ n497 ^ 1'b0 ;
  assign n19578 = ~n9780 & n19577 ;
  assign n19579 = n144 | n18735 ;
  assign n19580 = n799 & n1254 ;
  assign n19581 = n19580 ^ n14967 ^ 1'b0 ;
  assign n19582 = n497 | n1822 ;
  assign n19583 = n19582 ^ n403 ^ 1'b0 ;
  assign n19584 = n7729 & ~n19583 ;
  assign n19585 = n19584 ^ n2752 ^ 1'b0 ;
  assign n19586 = ~n4870 & n5551 ;
  assign n19587 = ~n2316 & n13696 ;
  assign n19588 = ~n14586 & n19587 ;
  assign n19589 = n5252 & ~n7383 ;
  assign n19590 = n227 & ~n19589 ;
  assign n19591 = n19544 & n19590 ;
  assign n19592 = ~n19588 & n19591 ;
  assign n19593 = n8757 | n11541 ;
  assign n19594 = n8067 & ~n19593 ;
  assign n19595 = n9594 ^ n1887 ^ n129 ;
  assign n19596 = n5124 & ~n12058 ;
  assign n19597 = n19596 ^ n6046 ^ n4903 ;
  assign n19598 = n756 & ~n8830 ;
  assign n19599 = n19598 ^ n15219 ^ 1'b0 ;
  assign n19600 = n2136 & ~n19599 ;
  assign n19601 = n19597 & ~n19600 ;
  assign n19602 = n19601 ^ n13908 ^ 1'b0 ;
  assign n19604 = n1139 ^ n55 ^ 1'b0 ;
  assign n19605 = n6933 & ~n19604 ;
  assign n19606 = ~n1050 & n19605 ;
  assign n19603 = n653 & n6439 ;
  assign n19607 = n19606 ^ n19603 ^ 1'b0 ;
  assign n19608 = n274 & ~n19607 ;
  assign n19609 = n2961 ^ n1217 ^ n348 ;
  assign n19610 = n568 & n10876 ;
  assign n19611 = n19610 ^ n8298 ^ 1'b0 ;
  assign n19612 = n19611 ^ n5350 ^ 1'b0 ;
  assign n19613 = n2298 & ~n13720 ;
  assign n19614 = ~n12388 & n19613 ;
  assign n19615 = n12462 | n13523 ;
  assign n19617 = n7652 ^ n1883 ^ 1'b0 ;
  assign n19616 = n5629 & ~n12207 ;
  assign n19618 = n19617 ^ n19616 ^ 1'b0 ;
  assign n19619 = n13843 ^ n628 ^ 1'b0 ;
  assign n19620 = n19618 | n19619 ;
  assign n19621 = n19620 ^ n12879 ^ 1'b0 ;
  assign n19622 = ~n3300 & n6331 ;
  assign n19623 = n1437 | n2116 ;
  assign n19624 = n607 | n19623 ;
  assign n19625 = n9091 ^ n3053 ^ 1'b0 ;
  assign n19626 = n19625 ^ n5326 ^ n609 ;
  assign n19627 = n13960 | n19088 ;
  assign n19628 = n10437 | n12777 ;
  assign n19629 = n8617 & n12453 ;
  assign n19630 = n2554 & n19629 ;
  assign n19631 = n12178 ^ n11827 ^ 1'b0 ;
  assign n19632 = ~n1929 & n17836 ;
  assign n19633 = ~n2661 & n16701 ;
  assign n19634 = n5862 & ~n17700 ;
  assign n19635 = n19633 & n19634 ;
  assign n19636 = n5270 | n10191 ;
  assign n19637 = n14472 | n19636 ;
  assign n19638 = n10154 ^ n290 ^ 1'b0 ;
  assign n19639 = n527 & ~n3285 ;
  assign n19640 = ~n5321 & n19639 ;
  assign n19641 = ~n5131 & n19640 ;
  assign n19642 = n19638 & n19641 ;
  assign n19643 = n666 ^ n153 ^ 1'b0 ;
  assign n19644 = n6709 & ~n19643 ;
  assign n19645 = ~n1061 & n19644 ;
  assign n19646 = n19645 ^ n25 ^ 1'b0 ;
  assign n19647 = n19646 ^ n977 ^ 1'b0 ;
  assign n19648 = n19642 & n19647 ;
  assign n19649 = n6577 ^ n328 ^ 1'b0 ;
  assign n19650 = n18002 ^ n1541 ^ n104 ;
  assign n19651 = n9195 ^ n2906 ^ 1'b0 ;
  assign n19652 = n812 & n13408 ;
  assign n19653 = n3068 & n19652 ;
  assign n19654 = n13028 & ~n19296 ;
  assign n19655 = n8291 & n10224 ;
  assign n19656 = n5851 ^ n164 ^ 1'b0 ;
  assign n19657 = n19656 ^ n6060 ^ 1'b0 ;
  assign n19658 = n7190 & n19657 ;
  assign n19659 = n16701 ^ n13248 ^ 1'b0 ;
  assign n19660 = n4740 & ~n10906 ;
  assign n19661 = n7032 ^ n467 ^ 1'b0 ;
  assign n19662 = n19661 ^ n2862 ^ 1'b0 ;
  assign n19663 = n19660 & n19662 ;
  assign n19664 = ~n382 & n6332 ;
  assign n19665 = n5136 ^ n434 ^ 1'b0 ;
  assign n19666 = ~n60 & n19665 ;
  assign n19667 = n12537 | n13101 ;
  assign n19668 = n8280 ^ n2978 ^ 1'b0 ;
  assign n19669 = n4603 & n18880 ;
  assign n19670 = n12409 & n19669 ;
  assign n19671 = n6234 ^ n2995 ^ 1'b0 ;
  assign n19672 = n4846 ^ n2768 ^ 1'b0 ;
  assign n19673 = n1390 & n15397 ;
  assign n19674 = n19672 | n19673 ;
  assign n19675 = n12804 ^ n10293 ^ 1'b0 ;
  assign n19676 = n4884 & n6887 ;
  assign n19677 = ~n4884 & n19676 ;
  assign n19678 = n6334 | n19677 ;
  assign n19679 = n19678 ^ n7259 ^ 1'b0 ;
  assign n19680 = ~n6398 & n19679 ;
  assign n19681 = n726 & n5156 ;
  assign n19682 = n8908 & ~n12512 ;
  assign n19683 = n19682 ^ n10064 ^ 1'b0 ;
  assign n19684 = n12657 & n15656 ;
  assign n19685 = ~n16152 & n19684 ;
  assign n19686 = n364 & n8526 ;
  assign n19687 = n2977 ^ n1831 ^ 1'b0 ;
  assign n19688 = n16742 ^ n5133 ^ n433 ;
  assign n19689 = n19687 | n19688 ;
  assign n19690 = n159 & n19689 ;
  assign n19691 = ( n1529 & n4117 ) | ( n1529 & ~n19690 ) | ( n4117 & ~n19690 ) ;
  assign n19692 = n7130 ^ n3483 ^ 1'b0 ;
  assign n19693 = n19691 & ~n19692 ;
  assign n19694 = n2144 & n7777 ;
  assign n19695 = n19694 ^ n843 ^ 1'b0 ;
  assign n19696 = n9927 ^ n6417 ^ 1'b0 ;
  assign n19697 = n233 | n525 ;
  assign n19698 = n19697 ^ n17811 ^ 1'b0 ;
  assign n19699 = n713 | n5376 ;
  assign n19700 = n12213 & ~n19699 ;
  assign n19701 = ~n15439 & n19700 ;
  assign n19702 = n19701 ^ n721 ^ 1'b0 ;
  assign n19703 = n17031 ^ n6768 ^ 1'b0 ;
  assign n19704 = n13048 | n19703 ;
  assign n19705 = n1606 & n2762 ;
  assign n19706 = n1399 & ~n6788 ;
  assign n19707 = n2969 & n8654 ;
  assign n19708 = n19707 ^ n2414 ^ 1'b0 ;
  assign n19709 = n19708 ^ n2005 ^ 1'b0 ;
  assign n19710 = ~n5727 & n14001 ;
  assign n19711 = n19710 ^ n9027 ^ 1'b0 ;
  assign n19712 = ~n712 & n11330 ;
  assign n19713 = ~n2414 & n12007 ;
  assign n19714 = n19713 ^ n12089 ^ 1'b0 ;
  assign n19715 = ( ~n6187 & n8529 ) | ( ~n6187 & n8810 ) | ( n8529 & n8810 ) ;
  assign n19716 = n945 & ~n958 ;
  assign n19717 = n19716 ^ n894 ^ 1'b0 ;
  assign n19718 = n11311 ^ n7380 ^ 1'b0 ;
  assign n19719 = n19717 | n19718 ;
  assign n19720 = n5927 & ~n19719 ;
  assign n19721 = n3493 ^ n128 ^ 1'b0 ;
  assign n19722 = n4880 | n19721 ;
  assign n19723 = n19722 ^ n1532 ^ 1'b0 ;
  assign n19724 = n19723 ^ n8064 ^ 1'b0 ;
  assign n19725 = n55 | n6222 ;
  assign n19726 = n1283 & ~n19725 ;
  assign n19727 = ~n5900 & n19726 ;
  assign n19728 = n19727 ^ n9670 ^ 1'b0 ;
  assign n19729 = n16236 & ~n19728 ;
  assign n19730 = n14423 & n19729 ;
  assign n19731 = n86 & n13872 ;
  assign n19732 = ~n2880 & n19731 ;
  assign n19733 = n4247 & n19314 ;
  assign n19734 = n11579 ^ n7646 ^ 1'b0 ;
  assign n19735 = n2497 ^ n1668 ^ 1'b0 ;
  assign n19736 = n7188 | n11957 ;
  assign n19737 = n19735 & ~n19736 ;
  assign n19738 = n1747 & ~n19737 ;
  assign n19739 = ~n1848 & n19738 ;
  assign n19740 = n5338 | n18490 ;
  assign n19741 = ~n1020 & n4952 ;
  assign n19742 = ~n3793 & n19741 ;
  assign n19743 = n1274 ^ n1198 ^ 1'b0 ;
  assign n19744 = n75 | n7059 ;
  assign n19745 = ~n4351 & n19744 ;
  assign n19746 = n16074 | n19745 ;
  assign n19747 = n12065 & ~n19746 ;
  assign n19748 = n19747 ^ n43 ^ 1'b0 ;
  assign n19749 = n7464 & n17122 ;
  assign n19750 = ~n1732 & n15770 ;
  assign n19751 = n9750 & n19750 ;
  assign n19752 = n3939 & n19751 ;
  assign n19753 = n17156 ^ n3566 ^ 1'b0 ;
  assign n19754 = ~n832 & n6868 ;
  assign n19755 = n8827 ^ n1447 ^ 1'b0 ;
  assign n19756 = n7685 ^ n2220 ^ 1'b0 ;
  assign n19757 = n5377 & ~n7812 ;
  assign n19758 = n456 | n10618 ;
  assign n19759 = ~n5799 & n19758 ;
  assign n19760 = n19757 | n19759 ;
  assign n19761 = ~n3290 & n17568 ;
  assign n19762 = ~n155 & n10041 ;
  assign n19763 = n19762 ^ n3139 ^ 1'b0 ;
  assign n19764 = n11064 ^ n3285 ^ 1'b0 ;
  assign n19765 = n9765 & ~n19764 ;
  assign n19766 = n9998 & n10379 ;
  assign n19767 = n19766 ^ n5090 ^ 1'b0 ;
  assign n19768 = n4750 & n10996 ;
  assign n19769 = ~n17199 & n19768 ;
  assign n19770 = ~n2349 & n5551 ;
  assign n19771 = n1406 & n19770 ;
  assign n19772 = n1095 & ~n4856 ;
  assign n19773 = n3280 & ~n19772 ;
  assign n19775 = n998 | n6830 ;
  assign n19774 = ~n7500 & n9376 ;
  assign n19776 = n19775 ^ n19774 ^ 1'b0 ;
  assign n19777 = n19776 ^ n13619 ^ 1'b0 ;
  assign n19778 = n7487 | n19777 ;
  assign n19779 = n9385 ^ n6131 ^ 1'b0 ;
  assign n19780 = ~n2546 & n19779 ;
  assign n19781 = n18488 & n19780 ;
  assign n19782 = n5727 & n10425 ;
  assign n19783 = n19782 ^ n5286 ^ 1'b0 ;
  assign n19784 = n520 & ~n10536 ;
  assign n19785 = n10261 ^ n7301 ^ 1'b0 ;
  assign n19786 = n1716 | n19785 ;
  assign n19787 = n1096 & ~n7185 ;
  assign n19788 = ~n2915 & n19787 ;
  assign n19789 = ~n1144 & n2549 ;
  assign n19790 = n17537 ^ n2634 ^ 1'b0 ;
  assign n19791 = n5495 & ~n19790 ;
  assign n19792 = n19791 ^ n4387 ^ 1'b0 ;
  assign n19793 = ~n19789 & n19792 ;
  assign n19794 = ~n649 & n19793 ;
  assign n19795 = n8548 & ~n19794 ;
  assign n19796 = n17597 & n19795 ;
  assign n19797 = n169 & n3065 ;
  assign n19798 = ~n14495 & n19797 ;
  assign n19799 = n19798 ^ n5118 ^ 1'b0 ;
  assign n19800 = n19799 ^ n16244 ^ 1'b0 ;
  assign n19801 = n1100 & n19800 ;
  assign n19802 = n5316 & ~n6878 ;
  assign n19803 = n19802 ^ n3915 ^ 1'b0 ;
  assign n19804 = n19803 ^ n9216 ^ 1'b0 ;
  assign n19805 = n8918 | n13729 ;
  assign n19806 = n15465 | n19805 ;
  assign n19807 = n7399 & n11910 ;
  assign n19808 = n10548 | n19807 ;
  assign n19809 = n68 | n296 ;
  assign n19810 = n296 & ~n19809 ;
  assign n19811 = ~n7609 & n19810 ;
  assign n19812 = n3256 & n19811 ;
  assign n19813 = n9434 ^ n1959 ^ 1'b0 ;
  assign n19814 = ~n19812 & n19813 ;
  assign n19815 = n19812 & n19814 ;
  assign n19816 = n19815 ^ n17308 ^ 1'b0 ;
  assign n19817 = n666 & n13023 ;
  assign n19818 = n484 & n19817 ;
  assign n19819 = n10421 & n10424 ;
  assign n19820 = n6764 ^ n2680 ^ 1'b0 ;
  assign n19824 = n60 | n613 ;
  assign n19825 = n11200 | n19824 ;
  assign n19826 = n19825 ^ n4509 ^ 1'b0 ;
  assign n19821 = n532 | n637 ;
  assign n19822 = n532 & ~n19821 ;
  assign n19823 = n3752 & ~n19822 ;
  assign n19827 = n19826 ^ n19823 ^ 1'b0 ;
  assign n19828 = ( n3939 & n12335 ) | ( n3939 & n19673 ) | ( n12335 & n19673 ) ;
  assign n19829 = n18227 ^ n1172 ^ 1'b0 ;
  assign n19830 = n13856 ^ n624 ^ 1'b0 ;
  assign n19831 = n2969 & n8883 ;
  assign n19832 = n19831 ^ n6041 ^ 1'b0 ;
  assign n19833 = n1388 | n9596 ;
  assign n19834 = n4169 | n19833 ;
  assign n19835 = n8590 ^ n1227 ^ 1'b0 ;
  assign n19836 = n5968 & n19835 ;
  assign n19837 = n17603 ^ n812 ^ 1'b0 ;
  assign n19838 = n2425 & n7706 ;
  assign n19839 = n16808 & ~n19838 ;
  assign n19840 = n17050 & n19839 ;
  assign n19841 = n7782 ^ n1141 ^ 1'b0 ;
  assign n19842 = ( n2375 & n3519 ) | ( n2375 & ~n19841 ) | ( n3519 & ~n19841 ) ;
  assign n19843 = ~n6076 & n19842 ;
  assign n19844 = n6618 ^ n701 ^ 1'b0 ;
  assign n19845 = n1309 & ~n19844 ;
  assign n19846 = n19843 & ~n19845 ;
  assign n19847 = n4879 & n19846 ;
  assign n19848 = n5950 ^ n4594 ^ n615 ;
  assign n19849 = n19848 ^ n14386 ^ 1'b0 ;
  assign n19850 = n5146 & ~n19849 ;
  assign n19851 = n1810 & n15025 ;
  assign n19852 = n19083 ^ n638 ^ 1'b0 ;
  assign n19853 = ~n1851 & n11559 ;
  assign n19854 = n258 & n448 ;
  assign n19855 = n11670 & n19854 ;
  assign n19856 = n19855 ^ n16193 ^ 1'b0 ;
  assign n19857 = n19856 ^ n9062 ^ n7872 ;
  assign n19858 = ~n158 & n9758 ;
  assign n19859 = n19858 ^ n14182 ^ 1'b0 ;
  assign n19860 = n626 ^ n595 ^ 1'b0 ;
  assign n19861 = n8439 & ~n19860 ;
  assign n19862 = n19861 ^ n11518 ^ 1'b0 ;
  assign n19863 = n19862 ^ n794 ^ 1'b0 ;
  assign n19864 = n19859 & n19863 ;
  assign n19865 = n17653 ^ n3181 ^ 1'b0 ;
  assign n19866 = n2103 & n2186 ;
  assign n19867 = ~n12258 & n19866 ;
  assign n19868 = n7674 & ~n19867 ;
  assign n19869 = n2566 | n13928 ;
  assign n19875 = n6967 ^ n2538 ^ 1'b0 ;
  assign n19874 = n873 | n5854 ;
  assign n19876 = n19875 ^ n19874 ^ 1'b0 ;
  assign n19870 = n2352 & n6647 ;
  assign n19871 = n9606 ^ n4560 ^ 1'b0 ;
  assign n19872 = ~n19870 & n19871 ;
  assign n19873 = ~n18731 & n19872 ;
  assign n19877 = n19876 ^ n19873 ^ 1'b0 ;
  assign n19878 = n5245 & n19708 ;
  assign n19879 = n19878 ^ n11643 ^ 1'b0 ;
  assign n19880 = n14376 ^ n4436 ^ 1'b0 ;
  assign n19881 = n14085 & ~n19880 ;
  assign n19882 = n2103 & ~n14233 ;
  assign n19891 = n2553 & n4734 ;
  assign n19892 = n19891 ^ n6432 ^ 1'b0 ;
  assign n19893 = n9402 & n19892 ;
  assign n19883 = n7665 & n11200 ;
  assign n19884 = n19883 ^ n2519 ^ 1'b0 ;
  assign n19886 = n2185 & ~n11568 ;
  assign n19885 = n768 | n9930 ;
  assign n19887 = n19886 ^ n19885 ^ 1'b0 ;
  assign n19888 = ~n12661 & n19887 ;
  assign n19889 = n3293 & n19888 ;
  assign n19890 = n19884 & ~n19889 ;
  assign n19894 = n19893 ^ n19890 ^ 1'b0 ;
  assign n19895 = ~n1804 & n1845 ;
  assign n19896 = n19895 ^ n4938 ^ 1'b0 ;
  assign n19897 = n10180 | n19896 ;
  assign n19898 = n163 & n16663 ;
  assign n19899 = n19898 ^ n4684 ^ 1'b0 ;
  assign n19900 = n4547 & n6683 ;
  assign n19901 = n19364 ^ n5366 ^ 1'b0 ;
  assign n19902 = n3137 & ~n19901 ;
  assign n19903 = ~n2549 & n14123 ;
  assign n19904 = n19903 ^ n17248 ^ 1'b0 ;
  assign n19905 = ~n687 & n1106 ;
  assign n19906 = n1705 | n11685 ;
  assign n19907 = n2439 ^ n1186 ^ 1'b0 ;
  assign n19908 = n1276 & ~n19907 ;
  assign n19909 = n8584 | n19908 ;
  assign n19910 = n4748 | n19909 ;
  assign n19911 = ~n1453 & n5953 ;
  assign n19912 = n3526 ^ n2161 ^ 1'b0 ;
  assign n19913 = ~n534 & n19912 ;
  assign n19914 = ~n13096 & n18069 ;
  assign n19915 = n2786 | n9252 ;
  assign n19916 = n161 & n4247 ;
  assign n19917 = ~n4247 & n19916 ;
  assign n19918 = n40 & ~n19917 ;
  assign n19919 = ~n40 & n19918 ;
  assign n19920 = n14466 ^ n6609 ^ 1'b0 ;
  assign n19921 = n11520 & ~n19920 ;
  assign n19922 = n15983 | n19921 ;
  assign n19923 = n19919 | n19922 ;
  assign n19924 = n19919 & ~n19923 ;
  assign n19925 = n70 | n867 ;
  assign n19926 = n70 & ~n19925 ;
  assign n19927 = n1645 & n19926 ;
  assign n19928 = ~n1318 & n19927 ;
  assign n19929 = ~n487 & n19928 ;
  assign n19930 = n19929 ^ n8723 ^ 1'b0 ;
  assign n19931 = n7394 & ~n19930 ;
  assign n19932 = n19924 & n19931 ;
  assign n19933 = n1366 | n2640 ;
  assign n19934 = n13831 ^ n985 ^ 1'b0 ;
  assign n19935 = ( ~n702 & n2448 ) | ( ~n702 & n12971 ) | ( n2448 & n12971 ) ;
  assign n19936 = ~n19934 & n19935 ;
  assign n19937 = ~n4504 & n19936 ;
  assign n19938 = n14779 ^ n7955 ^ 1'b0 ;
  assign n19939 = ~n7704 & n19938 ;
  assign n19940 = ( n6006 & n8916 ) | ( n6006 & ~n19939 ) | ( n8916 & ~n19939 ) ;
  assign n19941 = n940 | n1447 ;
  assign n19942 = n15915 ^ n5696 ^ 1'b0 ;
  assign n19943 = n2883 & ~n19942 ;
  assign n19944 = n15621 ^ n14569 ^ 1'b0 ;
  assign n19945 = n19944 ^ n10981 ^ 1'b0 ;
  assign n19946 = n9019 & n16108 ;
  assign n19947 = n19946 ^ n3749 ^ 1'b0 ;
  assign n19948 = n16981 | n19947 ;
  assign n19949 = n8903 | n19948 ;
  assign n19950 = n9338 | n19949 ;
  assign n19951 = n1019 & n6079 ;
  assign n19952 = n9121 & n19951 ;
  assign n19953 = n19952 ^ n542 ^ 1'b0 ;
  assign n19954 = n19950 & n19953 ;
  assign n19955 = n8056 | n15775 ;
  assign n19956 = n19955 ^ n310 ^ 1'b0 ;
  assign n19957 = n17341 ^ n1133 ^ 1'b0 ;
  assign n19958 = n1412 & n19957 ;
  assign n19959 = n11845 & ~n19958 ;
  assign n19960 = n19959 ^ n5609 ^ 1'b0 ;
  assign n19961 = ~n8734 & n19960 ;
  assign n19962 = ~n12525 & n19961 ;
  assign n19963 = n19962 ^ n8819 ^ 1'b0 ;
  assign n19964 = n8325 ^ n3443 ^ 1'b0 ;
  assign n19965 = n19963 & ~n19964 ;
  assign n19966 = ~n11748 & n19965 ;
  assign n19967 = n10824 | n17531 ;
  assign n19968 = n16819 | n19967 ;
  assign n19969 = n3789 ^ n2448 ^ 1'b0 ;
  assign n19970 = n4689 | n19969 ;
  assign n19971 = ~n2288 & n7369 ;
  assign n19972 = n12563 & n19971 ;
  assign n19973 = n4018 & n19972 ;
  assign n19974 = ~n2627 & n4469 ;
  assign n19975 = n1812 | n3756 ;
  assign n19976 = n19975 ^ n13700 ^ 1'b0 ;
  assign n19977 = n2670 & n19976 ;
  assign n19978 = n19977 ^ n8398 ^ 1'b0 ;
  assign n19979 = n423 & n1668 ;
  assign n19980 = ~n19978 & n19979 ;
  assign n19981 = n13643 ^ n378 ^ 1'b0 ;
  assign n19982 = n19981 ^ n8928 ^ 1'b0 ;
  assign n19983 = ~n19980 & n19982 ;
  assign n19984 = n8037 & n19983 ;
  assign n19985 = n19984 ^ n8242 ^ 1'b0 ;
  assign n19986 = n3993 ^ n715 ^ 1'b0 ;
  assign n19987 = n12361 ^ n9401 ^ 1'b0 ;
  assign n19988 = n6361 | n19987 ;
  assign n19989 = n5032 | n5235 ;
  assign n19990 = n3678 & ~n19989 ;
  assign n19991 = ~n310 & n3481 ;
  assign n19992 = n5340 ^ n3960 ^ 1'b0 ;
  assign n19993 = ~n19991 & n19992 ;
  assign n19994 = n19993 ^ n14674 ^ 1'b0 ;
  assign n19995 = n2155 | n19994 ;
  assign n19996 = n19995 ^ n2082 ^ 1'b0 ;
  assign n19997 = n1082 | n6431 ;
  assign n19998 = n19997 ^ n8784 ^ 1'b0 ;
  assign n19999 = n3307 & n19998 ;
  assign n20000 = n7667 | n19999 ;
  assign n20002 = ~n4879 & n12390 ;
  assign n20003 = n20002 ^ n1165 ^ 1'b0 ;
  assign n20004 = n15987 & n20003 ;
  assign n20005 = n20004 ^ n3501 ^ 1'b0 ;
  assign n20001 = n1447 & n5826 ;
  assign n20006 = n20005 ^ n20001 ^ n14221 ;
  assign n20007 = n2668 & ~n4790 ;
  assign n20008 = ~n3459 & n14768 ;
  assign n20009 = n20007 & n20008 ;
  assign n20010 = n20009 ^ n4166 ^ 1'b0 ;
  assign n20011 = n7288 & ~n17138 ;
  assign n20012 = n11323 ^ n5060 ^ 1'b0 ;
  assign n20013 = n5355 & ~n11405 ;
  assign n20016 = n7283 | n10086 ;
  assign n20014 = ~n3533 & n5364 ;
  assign n20015 = n14960 & ~n20014 ;
  assign n20017 = n20016 ^ n20015 ^ 1'b0 ;
  assign n20018 = n6284 ^ n294 ^ 1'b0 ;
  assign n20019 = n20018 ^ n15915 ^ n8828 ;
  assign n20020 = n11089 | n19014 ;
  assign n20021 = n20020 ^ n799 ^ 1'b0 ;
  assign n20022 = n9004 & n20021 ;
  assign n20023 = n804 & n8272 ;
  assign n20024 = n14254 ^ n8820 ^ 1'b0 ;
  assign n20025 = n20023 | n20024 ;
  assign n20026 = n20025 ^ n2067 ^ 1'b0 ;
  assign n20027 = n3929 & n20026 ;
  assign n20028 = ~n15473 & n20027 ;
  assign n20029 = n17804 ^ n13137 ^ 1'b0 ;
  assign n20030 = n4356 ^ n492 ^ 1'b0 ;
  assign n20031 = ~n594 & n20030 ;
  assign n20032 = n541 | n1560 ;
  assign n20033 = n20032 ^ n1377 ^ 1'b0 ;
  assign n20035 = ~n8140 & n11569 ;
  assign n20034 = ~n1673 & n7815 ;
  assign n20036 = n20035 ^ n20034 ^ 1'b0 ;
  assign n20037 = n4992 ^ n866 ^ 1'b0 ;
  assign n20038 = n16091 ^ n4273 ^ 1'b0 ;
  assign n20039 = ~n15232 & n20038 ;
  assign n20040 = n557 & ~n12382 ;
  assign n20041 = n257 | n11355 ;
  assign n20042 = n19879 & ~n20041 ;
  assign n20043 = n950 ^ n532 ^ n461 ;
  assign n20044 = ~n1794 & n20043 ;
  assign n20045 = n793 | n20044 ;
  assign n20046 = n7749 ^ n351 ^ 1'b0 ;
  assign n20047 = n2312 & ~n8432 ;
  assign n20048 = ~n5294 & n19317 ;
  assign n20049 = n10840 ^ n8230 ^ 1'b0 ;
  assign n20050 = n3028 & n20049 ;
  assign n20052 = n9106 ^ n7311 ^ 1'b0 ;
  assign n20051 = n8316 ^ n3081 ^ n663 ;
  assign n20053 = n20052 ^ n20051 ^ 1'b0 ;
  assign n20054 = n11533 ^ n7435 ^ 1'b0 ;
  assign n20055 = ~n3382 & n7759 ;
  assign n20057 = n18912 ^ n6272 ^ 1'b0 ;
  assign n20058 = n5716 & n20057 ;
  assign n20056 = ~n3649 & n4924 ;
  assign n20059 = n20058 ^ n20056 ^ 1'b0 ;
  assign n20060 = n622 & n6950 ;
  assign n20061 = n17834 ^ n820 ^ 1'b0 ;
  assign n20062 = n1231 & ~n13286 ;
  assign n20063 = ~n1165 & n6011 ;
  assign n20064 = n1165 & n20063 ;
  assign n20065 = n2542 & ~n17272 ;
  assign n20066 = n17272 & n20065 ;
  assign n20067 = n20064 & ~n20066 ;
  assign n20068 = n501 | n20067 ;
  assign n20069 = n20062 & ~n20068 ;
  assign n20070 = n366 & ~n2849 ;
  assign n20071 = n11359 & ~n20070 ;
  assign n20072 = n5534 ^ n2348 ^ 1'b0 ;
  assign n20073 = ~n8404 & n20072 ;
  assign n20074 = n6235 ^ n4028 ^ 1'b0 ;
  assign n20075 = n5116 | n20074 ;
  assign n20076 = n20075 ^ n1260 ^ 1'b0 ;
  assign n20077 = n20073 & n20076 ;
  assign n20078 = n20077 ^ n8081 ^ 1'b0 ;
  assign n20079 = n1390 & ~n6610 ;
  assign n20080 = n9768 & n20079 ;
  assign n20081 = ~n4396 & n20080 ;
  assign n20082 = n9682 ^ n5038 ^ 1'b0 ;
  assign n20083 = n3604 & n15336 ;
  assign n20084 = ~n15336 & n20083 ;
  assign n20085 = n1209 & ~n12395 ;
  assign n20086 = ~n7391 & n20085 ;
  assign n20087 = n13700 ^ n2403 ^ 1'b0 ;
  assign n20088 = n3492 & ~n8192 ;
  assign n20089 = ~n20087 & n20088 ;
  assign n20090 = n14418 ^ n6316 ^ 1'b0 ;
  assign n20091 = ~n1283 & n20090 ;
  assign n20092 = n5059 | n5252 ;
  assign n20093 = n2640 & ~n9531 ;
  assign n20094 = n3940 & n20093 ;
  assign n20095 = n20094 ^ n3579 ^ 1'b0 ;
  assign n20096 = n10676 & n20095 ;
  assign n20097 = n6955 ^ n5700 ^ 1'b0 ;
  assign n20098 = ~n3916 & n20097 ;
  assign n20099 = n3936 ^ n2822 ^ 1'b0 ;
  assign n20100 = ( n2719 & n10937 ) | ( n2719 & n15775 ) | ( n10937 & n15775 ) ;
  assign n20101 = n9531 | n18106 ;
  assign n20102 = n11105 ^ n8586 ^ 1'b0 ;
  assign n20103 = n1476 & ~n5891 ;
  assign n20104 = n10575 & ~n12222 ;
  assign n20105 = n3998 & n8935 ;
  assign n20106 = n20105 ^ n799 ^ 1'b0 ;
  assign n20107 = n20104 & ~n20106 ;
  assign n20109 = n1716 & n5561 ;
  assign n20110 = n6966 & n20109 ;
  assign n20111 = n20110 ^ n6240 ^ 1'b0 ;
  assign n20108 = n11323 ^ n3602 ^ n532 ;
  assign n20112 = n20111 ^ n20108 ^ 1'b0 ;
  assign n20113 = n13733 & ~n15426 ;
  assign n20114 = ~n14590 & n20113 ;
  assign n20115 = n20114 ^ n14557 ^ 1'b0 ;
  assign n20116 = ~n789 & n15334 ;
  assign n20117 = n4844 ^ n4171 ^ 1'b0 ;
  assign n20118 = n20116 & n20117 ;
  assign n20119 = n8910 ^ n1083 ^ 1'b0 ;
  assign n20120 = n18405 ^ n16058 ^ 1'b0 ;
  assign n20121 = n11636 | n20120 ;
  assign n20122 = n20121 ^ n18632 ^ 1'b0 ;
  assign n20123 = n608 & ~n1704 ;
  assign n20124 = n5179 & ~n20123 ;
  assign n20125 = ~n5805 & n20124 ;
  assign n20126 = n20125 ^ n14422 ^ 1'b0 ;
  assign n20127 = n4267 ^ n1423 ^ 1'b0 ;
  assign n20128 = n5569 & n20127 ;
  assign n20129 = n20128 ^ n11865 ^ 1'b0 ;
  assign n20130 = ~n2977 & n6330 ;
  assign n20131 = ~n5043 & n10041 ;
  assign n20132 = n20131 ^ n20107 ^ 1'b0 ;
  assign n20133 = ~n15711 & n17603 ;
  assign n20134 = n13988 ^ n9661 ^ 1'b0 ;
  assign n20135 = n8042 ^ n5343 ^ 1'b0 ;
  assign n20136 = ~n1388 & n3228 ;
  assign n20137 = n2011 | n18357 ;
  assign n20138 = n20137 ^ n6661 ^ 1'b0 ;
  assign n20139 = n4976 & ~n15368 ;
  assign n20140 = n3449 | n8006 ;
  assign n20141 = n20140 ^ n3765 ^ 1'b0 ;
  assign n20142 = n20141 ^ n18156 ^ n15029 ;
  assign n20143 = n14046 ^ n9614 ^ 1'b0 ;
  assign n20144 = ~n13308 & n15811 ;
  assign n20145 = n20144 ^ n11783 ^ 1'b0 ;
  assign n20146 = ~n6349 & n13074 ;
  assign n20147 = ~n3670 & n20146 ;
  assign n20148 = ~n12854 & n20147 ;
  assign n20149 = n11556 ^ n1642 ^ 1'b0 ;
  assign n20150 = n7848 & ~n20149 ;
  assign n20151 = n20150 ^ n7975 ^ 1'b0 ;
  assign n20180 = ~n604 & n1280 ;
  assign n20181 = n604 & n20180 ;
  assign n20182 = n4640 & ~n20181 ;
  assign n20152 = ~n117 & n443 ;
  assign n20153 = ~n443 & n20152 ;
  assign n20154 = n789 | n20153 ;
  assign n20155 = n789 & ~n20154 ;
  assign n20156 = n135 & ~n481 ;
  assign n20157 = n20155 & n20156 ;
  assign n20158 = n1609 & n20157 ;
  assign n20159 = ~n130 & n183 ;
  assign n20160 = ~n183 & n20159 ;
  assign n20161 = ~n7829 & n20160 ;
  assign n20162 = ~n380 & n20161 ;
  assign n20163 = ~n278 & n20162 ;
  assign n20164 = n34 & ~n60 ;
  assign n20165 = ~n34 & n20164 ;
  assign n20166 = n369 & n20165 ;
  assign n20167 = n492 & ~n20166 ;
  assign n20168 = n1105 & n13142 ;
  assign n20169 = n20167 | n20168 ;
  assign n20170 = n20163 & ~n20169 ;
  assign n20171 = n20158 | n20170 ;
  assign n20172 = n20158 & ~n20171 ;
  assign n20173 = ~n6306 & n20172 ;
  assign n20174 = n5673 & n20173 ;
  assign n20175 = n3592 & n12866 ;
  assign n20176 = ~n6073 & n20175 ;
  assign n20177 = ~n20175 & n20176 ;
  assign n20178 = n20174 & ~n20177 ;
  assign n20179 = n20178 ^ n18016 ^ 1'b0 ;
  assign n20183 = n20182 ^ n20179 ^ 1'b0 ;
  assign n20184 = ~n20151 & n20183 ;
  assign n20185 = n1425 ^ n102 ^ 1'b0 ;
  assign n20186 = n269 & ~n20185 ;
  assign n20187 = n20186 ^ n19719 ^ 1'b0 ;
  assign n20188 = n18226 & n18339 ;
  assign n20189 = n20188 ^ n9335 ^ 1'b0 ;
  assign n20190 = n16425 ^ n8366 ^ 1'b0 ;
  assign n20191 = n18587 & n19293 ;
  assign n20192 = n7454 | n15329 ;
  assign n20193 = n4815 ^ n1291 ^ 1'b0 ;
  assign n20194 = n6689 & n20193 ;
  assign n20195 = n15231 ^ n5090 ^ 1'b0 ;
  assign n20196 = n9999 ^ n4304 ^ 1'b0 ;
  assign n20197 = n6139 | n20196 ;
  assign n20198 = n4754 | n20197 ;
  assign n20199 = n7225 ^ n258 ^ 1'b0 ;
  assign n20200 = n20199 ^ n17390 ^ 1'b0 ;
  assign n20201 = n3803 & n20200 ;
  assign n20202 = n20201 ^ n1479 ^ 1'b0 ;
  assign n20203 = ~n5201 & n20202 ;
  assign n20204 = ~n9335 & n9978 ;
  assign n20205 = n498 | n2491 ;
  assign n20206 = ~n7639 & n9055 ;
  assign n20207 = ~n5457 & n20206 ;
  assign n20208 = n713 | n20207 ;
  assign n20209 = x3 & ~n6531 ;
  assign n20210 = n20209 ^ n13364 ^ 1'b0 ;
  assign n20212 = n984 & ~n5328 ;
  assign n20213 = ~n15183 & n20212 ;
  assign n20211 = n8457 & ~n10915 ;
  assign n20214 = n20213 ^ n20211 ^ 1'b0 ;
  assign n20215 = n7722 & n14387 ;
  assign n20216 = ~n1025 & n7355 ;
  assign n20217 = ( n4603 & n5373 ) | ( n4603 & ~n20216 ) | ( n5373 & ~n20216 ) ;
  assign n20218 = ~n4074 & n20217 ;
  assign n20219 = n20218 ^ n690 ^ 1'b0 ;
  assign n20220 = ~n20215 & n20219 ;
  assign n20221 = ~n3636 & n20220 ;
  assign n20222 = n2670 | n5771 ;
  assign n20223 = n3857 ^ n332 ^ 1'b0 ;
  assign n20224 = n1425 & n20223 ;
  assign n20225 = n14588 & n20224 ;
  assign n20226 = ~n2449 & n20181 ;
  assign n20227 = n350 & n14125 ;
  assign n20228 = ~n14125 & n20227 ;
  assign n20229 = n20226 & ~n20228 ;
  assign n20230 = ~n20226 & n20229 ;
  assign n20231 = n9197 | n18521 ;
  assign n20232 = n6148 | n20231 ;
  assign n20233 = n2842 & n17007 ;
  assign n20234 = n989 & n3965 ;
  assign n20235 = n20234 ^ n5372 ^ n2075 ;
  assign n20236 = n19332 ^ n15408 ^ 1'b0 ;
  assign n20237 = n4632 & ~n20236 ;
  assign n20238 = n19 | n5462 ;
  assign n20239 = n2043 ^ n53 ^ 1'b0 ;
  assign n20240 = n20239 ^ n2849 ^ 1'b0 ;
  assign n20241 = n1008 | n20240 ;
  assign n20242 = n8373 | n20241 ;
  assign n20243 = n7922 & n14048 ;
  assign n20244 = n16575 ^ n2148 ^ 1'b0 ;
  assign n20245 = x9 & ~n387 ;
  assign n20246 = n1036 & ~n7657 ;
  assign n20247 = n7988 | n14886 ;
  assign n20248 = n2657 | n20247 ;
  assign n20249 = n13976 ^ n6896 ^ 1'b0 ;
  assign n20250 = n6136 ^ n4780 ^ 1'b0 ;
  assign n20251 = n8777 | n20250 ;
  assign n20252 = n327 | n20251 ;
  assign n20253 = n17950 ^ n3103 ^ 1'b0 ;
  assign n20254 = n541 & n7814 ;
  assign n20255 = n1426 & n1619 ;
  assign n20256 = n3682 ^ n767 ^ 1'b0 ;
  assign n20257 = n9170 | n20256 ;
  assign n20258 = n5355 | n20257 ;
  assign n20259 = n3778 & n7427 ;
  assign n20260 = n4068 ^ n1063 ^ 1'b0 ;
  assign n20261 = n3637 & n20260 ;
  assign n20262 = ~n9364 & n20261 ;
  assign n20263 = n20259 & n20262 ;
  assign n20264 = n4165 ^ n274 ^ 1'b0 ;
  assign n20265 = n17300 ^ n146 ^ 1'b0 ;
  assign n20266 = n20264 & ~n20265 ;
  assign n20267 = n6080 & n6565 ;
  assign n20268 = n52 & n290 ;
  assign n20269 = n20268 ^ n5370 ^ 1'b0 ;
  assign n20270 = n221 | n15334 ;
  assign n20271 = n20270 ^ n4563 ^ 1'b0 ;
  assign n20272 = n20269 | n20271 ;
  assign n20273 = n7157 ^ n3103 ^ 1'b0 ;
  assign n20274 = n16243 & n20273 ;
  assign n20275 = n8946 | n20274 ;
  assign n20276 = n4133 & ~n5535 ;
  assign n20277 = ~n1109 & n5619 ;
  assign n20278 = ( ~n1880 & n6242 ) | ( ~n1880 & n20277 ) | ( n6242 & n20277 ) ;
  assign n20279 = n5283 ^ n2449 ^ 1'b0 ;
  assign n20280 = n12862 & n20279 ;
  assign n20281 = ~n2911 & n3833 ;
  assign n20282 = n8707 ^ n2510 ^ 1'b0 ;
  assign n20283 = n5076 & n20282 ;
  assign n20284 = n1026 ^ n715 ^ 1'b0 ;
  assign n20285 = n3133 | n17547 ;
  assign n20286 = n536 & ~n20285 ;
  assign n20287 = ~n3978 & n4279 ;
  assign n20288 = n17820 ^ n412 ^ 1'b0 ;
  assign n20289 = n20288 ^ n5326 ^ 1'b0 ;
  assign n20290 = n15602 ^ n4358 ^ 1'b0 ;
  assign n20291 = n10118 & n10169 ;
  assign n20292 = n1995 & n8104 ;
  assign n20293 = n15210 | n16126 ;
  assign n20294 = n9175 | n20293 ;
  assign n20295 = n20294 ^ n2943 ^ 1'b0 ;
  assign n20296 = n13126 | n20295 ;
  assign n20297 = n8115 ^ n2333 ^ 1'b0 ;
  assign n20298 = ~n17050 & n20297 ;
  assign n20299 = ( n10870 & n13163 ) | ( n10870 & n20298 ) | ( n13163 & n20298 ) ;
  assign n20300 = ~n12656 & n20299 ;
  assign n20301 = n20300 ^ n14443 ^ 1'b0 ;
  assign n20302 = n14396 ^ n2819 ^ 1'b0 ;
  assign n20303 = n4029 | n20302 ;
  assign n20304 = ~n13544 & n14455 ;
  assign n20305 = n4549 & n6296 ;
  assign n20306 = ~n6296 & n20305 ;
  assign n20307 = n9539 & ~n20306 ;
  assign n20308 = n16276 ^ n10261 ^ 1'b0 ;
  assign n20309 = n20307 & n20308 ;
  assign n20310 = n16476 ^ n1191 ^ 1'b0 ;
  assign n20311 = n6371 & n11783 ;
  assign n20312 = n10172 ^ n468 ^ 1'b0 ;
  assign n20313 = n498 & ~n872 ;
  assign n20314 = ~n1560 & n1693 ;
  assign n20315 = ( n1685 & n20313 ) | ( n1685 & ~n20314 ) | ( n20313 & ~n20314 ) ;
  assign n20316 = ( n736 & ~n8628 ) | ( n736 & n9191 ) | ( ~n8628 & n9191 ) ;
  assign n20317 = ~n532 & n20316 ;
  assign n20318 = n14452 & ~n16029 ;
  assign n20319 = n3219 & ~n15607 ;
  assign n20320 = n20318 & n20319 ;
  assign n20321 = n5083 & ~n15811 ;
  assign n20322 = n19327 ^ n2582 ^ 1'b0 ;
  assign n20323 = n14438 & n15673 ;
  assign n20324 = ( n16222 & n20322 ) | ( n16222 & n20323 ) | ( n20322 & n20323 ) ;
  assign n20325 = n1163 & ~n12639 ;
  assign n20326 = n14064 ^ n13196 ^ 1'b0 ;
  assign n20327 = n4915 | n20326 ;
  assign n20328 = n20327 ^ n5170 ^ 1'b0 ;
  assign n20329 = n8450 ^ n3999 ^ 1'b0 ;
  assign n20330 = ~n4277 & n7855 ;
  assign n20331 = ~n500 & n20330 ;
  assign n20332 = n11724 & n20331 ;
  assign n20333 = n20329 & ~n20332 ;
  assign n20334 = n641 & n11350 ;
  assign n20335 = n653 & ~n11384 ;
  assign n20336 = ~n235 & n20335 ;
  assign n20337 = n14991 & ~n20336 ;
  assign n20338 = ~n7717 & n20337 ;
  assign n20339 = n12887 | n20338 ;
  assign n20340 = n1271 & n9994 ;
  assign n20341 = n20340 ^ n19958 ^ 1'b0 ;
  assign n20342 = ~n4373 & n20341 ;
  assign n20343 = n6089 ^ n3696 ^ 1'b0 ;
  assign n20344 = n11096 | n20343 ;
  assign n20345 = n20344 ^ n1359 ^ n1226 ;
  assign n20346 = n19627 ^ n2542 ^ 1'b0 ;
  assign n20347 = n20345 & ~n20346 ;
  assign n20348 = n340 | n15909 ;
  assign n20349 = n4640 | n9242 ;
  assign n20350 = n6843 | n20349 ;
  assign n20351 = n20348 & ~n20350 ;
  assign n20352 = n15703 ^ n8819 ^ 1'b0 ;
  assign n20353 = n3292 & ~n20352 ;
  assign n20354 = n3210 & ~n12502 ;
  assign n20355 = n2905 ^ n481 ^ 1'b0 ;
  assign n20356 = ~n1867 & n20355 ;
  assign n20357 = n20296 ^ n4054 ^ 1'b0 ;
  assign n20358 = n2440 & n10167 ;
  assign n20359 = n20358 ^ n2120 ^ 1'b0 ;
  assign n20360 = ~n9657 & n20036 ;
  assign n20361 = ( n2531 & ~n4435 ) | ( n2531 & n12902 ) | ( ~n4435 & n12902 ) ;
  assign n20362 = n633 | n7138 ;
  assign n20363 = n2550 | n20362 ;
  assign n20364 = n7234 & ~n17442 ;
  assign n20365 = n20364 ^ n690 ^ 1'b0 ;
  assign n20366 = n1394 & n5211 ;
  assign n20367 = ~n5211 & n20366 ;
  assign n20368 = n6830 | n20367 ;
  assign n20369 = n6830 & ~n20368 ;
  assign n20370 = n15149 & ~n20369 ;
  assign n20371 = n20370 ^ n9064 ^ 1'b0 ;
  assign n20372 = n20371 ^ n19961 ^ n4687 ;
  assign n20373 = n3853 & ~n6785 ;
  assign n20374 = n8571 & ~n20373 ;
  assign n20375 = ~n678 & n4677 ;
  assign n20376 = n20375 ^ n2410 ^ 1'b0 ;
  assign n20377 = ~n1098 & n20376 ;
  assign n20378 = n9906 ^ n5826 ^ 1'b0 ;
  assign n20379 = n20377 & ~n20378 ;
  assign n20380 = ( n4801 & n6306 ) | ( n4801 & n6594 ) | ( n6306 & n6594 ) ;
  assign n20381 = n5795 & ~n20380 ;
  assign n20382 = n20381 ^ n6055 ^ 1'b0 ;
  assign n20383 = n20382 ^ n11322 ^ 1'b0 ;
  assign n20384 = n9839 & n11698 ;
  assign n20385 = n8988 & ~n20384 ;
  assign n20386 = n20385 ^ n19747 ^ 1'b0 ;
  assign n20387 = n6964 & n8770 ;
  assign n20388 = n582 & ~n7142 ;
  assign n20389 = ~n9484 & n20388 ;
  assign n20390 = n18009 ^ n8309 ^ 1'b0 ;
  assign n20391 = ~n8459 & n20390 ;
  assign n20392 = n5819 ^ n80 ^ 1'b0 ;
  assign n20393 = n5164 ^ n5125 ^ 1'b0 ;
  assign n20394 = n2951 | n20393 ;
  assign n20395 = n2511 ^ n908 ^ 1'b0 ;
  assign n20396 = ~n190 & n20395 ;
  assign n20397 = n20396 ^ n3346 ^ 1'b0 ;
  assign n20398 = n3037 & n11696 ;
  assign n20399 = n20398 ^ n2661 ^ 1'b0 ;
  assign n20400 = n15276 & ~n20399 ;
  assign n20401 = n1922 & ~n10670 ;
  assign n20402 = n3713 & n11405 ;
  assign n20405 = n924 ^ n565 ^ 1'b0 ;
  assign n20406 = n3479 & n20405 ;
  assign n20403 = n14174 ^ n325 ^ 1'b0 ;
  assign n20404 = n4754 & ~n20403 ;
  assign n20407 = n20406 ^ n20404 ^ n15509 ;
  assign n20408 = n9592 & n20407 ;
  assign n20409 = n20408 ^ n10635 ^ n2141 ;
  assign n20410 = n6464 & n20409 ;
  assign n20411 = n1631 & n20410 ;
  assign n20412 = n16384 ^ n4563 ^ 1'b0 ;
  assign n20413 = n13352 | n16877 ;
  assign n20414 = n16877 & ~n20413 ;
  assign n20415 = n415 | n9756 ;
  assign n20416 = n20415 ^ n12066 ^ 1'b0 ;
  assign n20417 = n2987 & n14955 ;
  assign n20418 = n2541 | n3791 ;
  assign n20419 = n12225 | n20418 ;
  assign n20420 = n3567 | n14254 ;
  assign n20421 = n5161 | n9623 ;
  assign n20422 = n20421 ^ n14922 ^ n6683 ;
  assign n20423 = n5682 ^ n5583 ^ 1'b0 ;
  assign n20424 = n15967 ^ n1929 ^ 1'b0 ;
  assign n20425 = n14978 & ~n20424 ;
  assign n20426 = ~n1109 & n10107 ;
  assign n20427 = ~n6875 & n20426 ;
  assign n20428 = ~n10430 & n18852 ;
  assign n20429 = n19505 ^ n2566 ^ 1'b0 ;
  assign n20430 = ~n1790 & n20429 ;
  assign n20431 = n1880 & n15869 ;
  assign n20432 = ( n1310 & n3559 ) | ( n1310 & n20431 ) | ( n3559 & n20431 ) ;
  assign n20433 = n1344 & n11185 ;
  assign n20434 = n20433 ^ n20289 ^ 1'b0 ;
  assign n20435 = n7935 & ~n17009 ;
  assign n20436 = ~n4223 & n20435 ;
  assign n20437 = n1898 ^ n1704 ^ 1'b0 ;
  assign n20438 = n20437 ^ n5227 ^ 1'b0 ;
  assign n20439 = n1602 & ~n20438 ;
  assign n20440 = n11756 & ~n15604 ;
  assign n20441 = n20440 ^ n11593 ^ 1'b0 ;
  assign n20442 = n14120 & n14491 ;
  assign n20443 = n20442 ^ n1491 ^ 1'b0 ;
  assign n20444 = n7249 | n9281 ;
  assign n20445 = n1237 & ~n20444 ;
  assign n20446 = n15291 & n20445 ;
  assign n20447 = ~n1219 & n20446 ;
  assign n20448 = n7698 | n9394 ;
  assign n20449 = n20448 ^ n11827 ^ 1'b0 ;
  assign n20450 = n10725 | n12390 ;
  assign n20451 = n20450 ^ n356 ^ 1'b0 ;
  assign n20452 = n7732 & ~n8950 ;
  assign n20453 = n20452 ^ n4964 ^ 1'b0 ;
  assign n20454 = ~n9397 & n20453 ;
  assign n20455 = n931 & n3744 ;
  assign n20456 = n20455 ^ n7520 ^ 1'b0 ;
  assign n20457 = n9764 | n20456 ;
  assign n20458 = n20457 ^ n6758 ^ 1'b0 ;
  assign n20459 = n5317 | n20458 ;
  assign n20460 = n20459 ^ n16286 ^ 1'b0 ;
  assign n20461 = n17229 | n20460 ;
  assign n20462 = n461 | n662 ;
  assign n20463 = n20462 ^ n825 ^ 1'b0 ;
  assign n20464 = n3007 | n4935 ;
  assign n20465 = n1339 & ~n20464 ;
  assign n20466 = n20465 ^ n19149 ^ 1'b0 ;
  assign n20467 = n20463 & ~n20466 ;
  assign n20468 = n1958 ^ n1571 ^ 1'b0 ;
  assign n20469 = n12694 ^ n2786 ^ 1'b0 ;
  assign n20470 = n16070 ^ n9673 ^ 1'b0 ;
  assign n20471 = n3226 & ~n5885 ;
  assign n20472 = n20471 ^ n8614 ^ 1'b0 ;
  assign n20473 = n9828 ^ n5241 ^ 1'b0 ;
  assign n20474 = n13857 ^ n2580 ^ 1'b0 ;
  assign n20475 = n2547 & ~n7008 ;
  assign n20476 = n20475 ^ n9923 ^ 1'b0 ;
  assign n20477 = ~n3080 & n13362 ;
  assign n20478 = n20477 ^ n1432 ^ 1'b0 ;
  assign n20479 = n5827 | n13558 ;
  assign n20480 = n9881 & ~n20479 ;
  assign n20481 = n3784 & ~n20480 ;
  assign n20482 = n5995 & n20481 ;
  assign n20483 = n8764 & n13857 ;
  assign n20484 = n2452 & n7111 ;
  assign n20485 = ~n17486 & n20484 ;
  assign n20486 = n1829 & n20485 ;
  assign n20487 = n1545 | n8568 ;
  assign n20488 = ~n3856 & n20487 ;
  assign n20489 = n322 & n10188 ;
  assign n20490 = ~n5193 & n20489 ;
  assign n20491 = n5910 & ~n8489 ;
  assign n20492 = ~n1172 & n20491 ;
  assign n20493 = ( n16603 & ~n17843 ) | ( n16603 & n20492 ) | ( ~n17843 & n20492 ) ;
  assign n20495 = n1227 | n2400 ;
  assign n20494 = n14339 | n19831 ;
  assign n20496 = n20495 ^ n20494 ^ 1'b0 ;
  assign n20497 = n6043 | n13781 ;
  assign n20498 = ~n3939 & n10343 ;
  assign n20499 = n12115 & n20498 ;
  assign n20500 = n20499 ^ n5707 ^ 1'b0 ;
  assign n20501 = n20497 | n20500 ;
  assign n20502 = n8730 ^ n2173 ^ 1'b0 ;
  assign n20503 = n13554 & n20502 ;
  assign n20504 = n11039 & ~n16680 ;
  assign n20505 = n3015 & n11453 ;
  assign n20506 = n2840 & ~n5155 ;
  assign n20507 = ( n6942 & n8105 ) | ( n6942 & ~n15900 ) | ( n8105 & ~n15900 ) ;
  assign n20508 = n20506 | n20507 ;
  assign n20509 = n185 & n20508 ;
  assign n20510 = n20505 & n20509 ;
  assign n20511 = n7896 ^ n4181 ^ 1'b0 ;
  assign n20512 = ~n4274 & n9357 ;
  assign n20513 = n3924 & n5775 ;
  assign n20514 = n4123 & ~n4650 ;
  assign n20515 = ( n11650 & ~n15131 ) | ( n11650 & n15893 ) | ( ~n15131 & n15893 ) ;
  assign n20516 = ~n2485 & n10846 ;
  assign n20517 = n5549 ^ n5263 ^ n5083 ;
  assign n20518 = n105 & ~n2785 ;
  assign n20519 = n20518 ^ n14845 ^ 1'b0 ;
  assign n20520 = ~n20517 & n20519 ;
  assign n20521 = n15204 ^ n5002 ^ n1106 ;
  assign n20522 = n1199 | n17479 ;
  assign n20523 = n1186 & ~n9493 ;
  assign n20524 = x3 & ~n1177 ;
  assign n20525 = n20524 ^ n1759 ^ 1'b0 ;
  assign n20526 = n20525 ^ n5225 ^ 1'b0 ;
  assign n20527 = ~n14730 & n20526 ;
  assign n20528 = ~n3990 & n7116 ;
  assign n20529 = n8360 ^ n268 ^ 1'b0 ;
  assign n20530 = n4626 ^ n3074 ^ 1'b0 ;
  assign n20531 = n20529 & ~n20530 ;
  assign n20532 = n1944 & n20531 ;
  assign n20533 = n20532 ^ n5780 ^ 1'b0 ;
  assign n20534 = n16527 ^ n2945 ^ 1'b0 ;
  assign n20535 = n104 & n20534 ;
  assign n20536 = ~n10521 & n20535 ;
  assign n20537 = ~n20535 & n20536 ;
  assign n20538 = n9768 & ~n20537 ;
  assign n20539 = n8206 & n20538 ;
  assign n20540 = x7 | n8486 ;
  assign n20541 = n20540 ^ n12269 ^ 1'b0 ;
  assign n20542 = n10084 ^ n1385 ^ 1'b0 ;
  assign n20543 = n1888 & n12205 ;
  assign n20544 = n20543 ^ n3715 ^ 1'b0 ;
  assign n20545 = n20542 & ~n20544 ;
  assign n20546 = n20545 ^ n8107 ^ 1'b0 ;
  assign n20547 = n11235 | n20546 ;
  assign n20548 = n6867 ^ n1043 ^ 1'b0 ;
  assign n20549 = n19175 | n20548 ;
  assign n20550 = n2534 | n2610 ;
  assign n20551 = n20550 ^ n10897 ^ 1'b0 ;
  assign n20552 = n4969 | n9495 ;
  assign n20553 = n15549 ^ n3877 ^ 1'b0 ;
  assign n20554 = n4819 & n10007 ;
  assign n20555 = n20554 ^ n6402 ^ 1'b0 ;
  assign n20556 = n20555 ^ n4986 ^ 1'b0 ;
  assign n20557 = n20556 ^ n1718 ^ 1'b0 ;
  assign n20558 = n8541 & ~n20557 ;
  assign n20559 = n10739 ^ n8828 ^ 1'b0 ;
  assign n20560 = n14132 | n20559 ;
  assign n20561 = n20560 ^ n18624 ^ 1'b0 ;
  assign n20566 = n7075 | n13422 ;
  assign n20562 = n540 & ~n6290 ;
  assign n20563 = n2936 | n20562 ;
  assign n20564 = ~n15221 & n20563 ;
  assign n20565 = ~n6039 & n20564 ;
  assign n20567 = n20566 ^ n20565 ^ 1'b0 ;
  assign n20568 = n12680 ^ n5643 ^ 1'b0 ;
  assign n20569 = ~n12175 & n20568 ;
  assign n20570 = n10718 ^ n8148 ^ n4274 ;
  assign n20571 = n12699 | n16981 ;
  assign n20572 = n20570 & ~n20571 ;
  assign n20573 = n3315 & n11178 ;
  assign n20574 = n527 & ~n20573 ;
  assign n20575 = n20574 ^ n1322 ^ 1'b0 ;
  assign n20576 = n6093 & ~n8842 ;
  assign n20578 = n7061 ^ n2608 ^ 1'b0 ;
  assign n20577 = ~n10344 & n15777 ;
  assign n20579 = n20578 ^ n20577 ^ 1'b0 ;
  assign n20580 = n3032 | n20579 ;
  assign n20581 = n1765 & ~n20580 ;
  assign n20582 = n5643 & ~n5774 ;
  assign n20583 = n5984 & n10033 ;
  assign n20584 = ~n1537 & n20583 ;
  assign n20585 = n8153 | n20584 ;
  assign n20586 = n3997 & n7288 ;
  assign n20587 = ~n8363 & n16013 ;
  assign n20588 = n12378 & n20587 ;
  assign n20589 = n6198 | n17713 ;
  assign n20590 = n10591 | n17791 ;
  assign n20591 = n20590 ^ n19038 ^ 1'b0 ;
  assign n20592 = n13628 | n20105 ;
  assign n20593 = n15748 | n20592 ;
  assign n20594 = n1963 ^ n408 ^ 1'b0 ;
  assign n20595 = ~n8987 & n16506 ;
  assign n20596 = n607 | n1842 ;
  assign n20597 = n20596 ^ n3742 ^ 1'b0 ;
  assign n20600 = n212 | n1396 ;
  assign n20601 = n14737 & ~n20600 ;
  assign n20598 = n11476 & ~n15725 ;
  assign n20599 = ~n7368 & n20598 ;
  assign n20602 = n20601 ^ n20599 ^ 1'b0 ;
  assign n20603 = n19542 | n20602 ;
  assign n20604 = n2209 & ~n20603 ;
  assign n20605 = ~n9687 & n15050 ;
  assign n20606 = n986 ^ n767 ^ 1'b0 ;
  assign n20607 = ~n2894 & n20606 ;
  assign n20608 = n4728 ^ n4537 ^ 1'b0 ;
  assign n20609 = n9229 ^ n573 ^ 1'b0 ;
  assign n20610 = n15319 | n20609 ;
  assign n20611 = ~n20608 & n20610 ;
  assign n20612 = n1520 & ~n16138 ;
  assign n20613 = ~n5775 & n10870 ;
  assign n20614 = n20613 ^ n1444 ^ 1'b0 ;
  assign n20615 = n15626 & n15929 ;
  assign n20616 = n16862 & n20615 ;
  assign n20617 = n1637 & ~n7497 ;
  assign n20618 = ~n20616 & n20617 ;
  assign n20619 = n10940 | n17044 ;
  assign n20620 = n20619 ^ n2303 ^ 1'b0 ;
  assign n20625 = n1310 & ~n16137 ;
  assign n20621 = ~n991 & n2059 ;
  assign n20622 = ~n266 & n20621 ;
  assign n20623 = n20622 ^ n2535 ^ 1'b0 ;
  assign n20624 = ~n2140 & n20623 ;
  assign n20626 = n20625 ^ n20624 ^ 1'b0 ;
  assign n20627 = n8773 & n11795 ;
  assign n20628 = n18026 & n20627 ;
  assign n20629 = n1283 & ~n2745 ;
  assign n20630 = n14713 & ~n20629 ;
  assign n20631 = n20630 ^ n2681 ^ 1'b0 ;
  assign n20635 = n7261 ^ n458 ^ 1'b0 ;
  assign n20636 = n503 & n20635 ;
  assign n20632 = n15310 & ~n17165 ;
  assign n20633 = ~n18622 & n20632 ;
  assign n20634 = n3645 & ~n20633 ;
  assign n20637 = n20636 ^ n20634 ^ 1'b0 ;
  assign n20638 = n13877 ^ n847 ^ 1'b0 ;
  assign n20639 = n1154 | n13885 ;
  assign n20640 = n20638 & ~n20639 ;
  assign n20641 = n4031 | n11714 ;
  assign n20642 = n10169 ^ n7604 ^ 1'b0 ;
  assign n20643 = n6498 & n20642 ;
  assign n20644 = n17924 & ~n20643 ;
  assign n20645 = n2751 | n7673 ;
  assign n20646 = ~n9324 & n10977 ;
  assign n20647 = n20646 ^ n9889 ^ 1'b0 ;
  assign n20648 = n20647 ^ n7718 ^ n865 ;
  assign n20649 = n3493 ^ n3374 ^ 1'b0 ;
  assign n20650 = n2549 & ~n12402 ;
  assign n20651 = n10315 ^ n6320 ^ 1'b0 ;
  assign n20652 = n3114 & n20651 ;
  assign n20653 = ~n8236 & n20652 ;
  assign n20654 = n20650 & n20653 ;
  assign n20655 = n20654 ^ n7681 ^ 1'b0 ;
  assign n20656 = n7938 | n20655 ;
  assign n20657 = n1133 & ~n6436 ;
  assign n20658 = ~n11365 & n20657 ;
  assign n20659 = ~n9175 & n20658 ;
  assign n20661 = n3429 ^ n949 ^ 1'b0 ;
  assign n20662 = n2564 | n20661 ;
  assign n20663 = n20662 ^ n2011 ^ 1'b0 ;
  assign n20660 = ~n6942 & n12297 ;
  assign n20664 = n20663 ^ n20660 ^ 1'b0 ;
  assign n20665 = n7495 ^ n5005 ^ 1'b0 ;
  assign n20666 = ( n1174 & n8843 ) | ( n1174 & n20665 ) | ( n8843 & n20665 ) ;
  assign n20667 = n956 & n10879 ;
  assign n20668 = n10546 ^ n5934 ^ 1'b0 ;
  assign n20669 = ~n20667 & n20668 ;
  assign n20670 = ~n16362 & n17342 ;
  assign n20671 = ~n13691 & n17303 ;
  assign n20672 = n20671 ^ n10559 ^ 1'b0 ;
  assign n20673 = n4756 & ~n7140 ;
  assign n20674 = n15042 & n20673 ;
  assign n20675 = n722 & n11703 ;
  assign n20676 = ~n4034 & n20675 ;
  assign n20677 = n56 & ~n5292 ;
  assign n20678 = n3546 & ~n19364 ;
  assign n20679 = n20678 ^ n11465 ^ 1'b0 ;
  assign n20680 = n9082 ^ n4919 ^ 1'b0 ;
  assign n20681 = n20679 | n20680 ;
  assign n20682 = n3046 ^ n2059 ^ 1'b0 ;
  assign n20683 = n20128 & ~n20682 ;
  assign n20684 = n20683 ^ n4984 ^ 1'b0 ;
  assign n20685 = n261 & n7392 ;
  assign n20686 = ( n3221 & n9963 ) | ( n3221 & ~n20685 ) | ( n9963 & ~n20685 ) ;
  assign n20687 = n2642 & ~n16655 ;
  assign n20688 = n20687 ^ n15896 ^ 1'b0 ;
  assign n20689 = n10414 ^ n1822 ^ 1'b0 ;
  assign n20690 = n15090 & ~n20689 ;
  assign n20691 = n719 | n7740 ;
  assign n20692 = n20691 ^ n15032 ^ 1'b0 ;
  assign n20693 = n1034 ^ n281 ^ 1'b0 ;
  assign n20694 = n4349 & ~n12913 ;
  assign n20695 = n16443 & n20694 ;
  assign n20696 = n17174 ^ n4256 ^ 1'b0 ;
  assign n20697 = n20695 & ~n20696 ;
  assign n20698 = n20697 ^ n1908 ^ 1'b0 ;
  assign n20699 = n20698 ^ n4514 ^ 1'b0 ;
  assign n20700 = ~n462 & n20699 ;
  assign n20701 = n19 | n60 ;
  assign n20702 = n18163 & ~n20701 ;
  assign n20703 = n20702 ^ n4574 ^ 1'b0 ;
  assign n20704 = ( n1875 & n6078 ) | ( n1875 & n20703 ) | ( n6078 & n20703 ) ;
  assign n20705 = ~n5979 & n20704 ;
  assign n20706 = ~n817 & n20705 ;
  assign n20707 = n367 | n20706 ;
  assign n20708 = n20707 ^ n3479 ^ 1'b0 ;
  assign n20709 = n6955 & n18103 ;
  assign n20710 = ~n767 & n13009 ;
  assign n20711 = n1289 | n4406 ;
  assign n20712 = ~n4732 & n5785 ;
  assign n20713 = ~n9410 & n20712 ;
  assign n20714 = n20713 ^ n19770 ^ 1'b0 ;
  assign n20715 = n20711 & n20714 ;
  assign n20716 = n9212 ^ n960 ^ 1'b0 ;
  assign n20717 = n6378 | n14886 ;
  assign n20718 = n8508 & ~n20717 ;
  assign n20719 = n5256 & ~n6244 ;
  assign n20720 = n13006 & ~n20719 ;
  assign n20721 = n20720 ^ n12649 ^ 1'b0 ;
  assign n20722 = n12859 & n20456 ;
  assign n20723 = n2883 & n20722 ;
  assign n20724 = ~n2594 & n14165 ;
  assign n20725 = ~n20723 & n20724 ;
  assign n20726 = n745 | n20601 ;
  assign n20727 = n20726 ^ n1462 ^ 1'b0 ;
  assign n20728 = n20727 ^ n15661 ^ n10691 ;
  assign n20729 = n20728 ^ n5533 ^ 1'b0 ;
  assign n20730 = n5713 | n16318 ;
  assign n20731 = ~n15843 & n20730 ;
  assign n20732 = n17884 ^ n11111 ^ 1'b0 ;
  assign n20733 = n2078 & ~n20732 ;
  assign n20734 = n236 & ~n6145 ;
  assign n20735 = n20734 ^ n10967 ^ 1'b0 ;
  assign n20736 = n5769 ^ n821 ^ 1'b0 ;
  assign n20737 = n302 & ~n10269 ;
  assign n20738 = ~n20736 & n20737 ;
  assign n20739 = n16375 | n16525 ;
  assign n20740 = n20739 ^ n20696 ^ 1'b0 ;
  assign n20741 = n20740 ^ n16221 ^ 1'b0 ;
  assign n20742 = n20738 | n20741 ;
  assign n20743 = n15528 | n19796 ;
  assign n20744 = n367 & ~n20743 ;
  assign n20745 = ( n144 & ~n2209 ) | ( n144 & n5537 ) | ( ~n2209 & n5537 ) ;
  assign n20746 = n83 & ~n6831 ;
  assign n20747 = n9193 & n20746 ;
  assign n20748 = n20747 ^ n3871 ^ 1'b0 ;
  assign n20749 = n800 & n20748 ;
  assign n20750 = n425 & ~n20749 ;
  assign n20751 = ~n1177 & n20750 ;
  assign n20752 = n11403 & n18953 ;
  assign n20753 = n18719 | n20752 ;
  assign n20754 = n3826 & n15814 ;
  assign n20755 = n15390 ^ n11164 ^ 1'b0 ;
  assign n20756 = n10101 ^ n1132 ^ 1'b0 ;
  assign n20757 = n11115 & n20756 ;
  assign n20758 = ~n231 & n20757 ;
  assign n20759 = n17528 ^ n8429 ^ 1'b0 ;
  assign n20760 = ~n20758 & n20759 ;
  assign n20761 = ( ~n4899 & n5070 ) | ( ~n4899 & n5588 ) | ( n5070 & n5588 ) ;
  assign n20762 = ~n3632 & n20761 ;
  assign n20763 = n20762 ^ n18634 ^ 1'b0 ;
  assign n20764 = n18308 ^ n10025 ^ 1'b0 ;
  assign n20765 = ~n18478 & n20764 ;
  assign n20766 = n3423 & n20765 ;
  assign n20767 = n6664 & n14232 ;
  assign n20768 = n17030 ^ n15064 ^ 1'b0 ;
  assign n20769 = n284 | n8415 ;
  assign n20770 = n20769 ^ n11468 ^ 1'b0 ;
  assign n20771 = n4869 & ~n20770 ;
  assign n20772 = n2016 ^ x5 ^ 1'b0 ;
  assign n20773 = n187 & ~n16347 ;
  assign n20774 = n20773 ^ n4977 ^ 1'b0 ;
  assign n20775 = n15900 & n20774 ;
  assign n20776 = n18811 ^ n6087 ^ 1'b0 ;
  assign n20777 = n14316 | n20776 ;
  assign n20778 = n19651 ^ n11929 ^ 1'b0 ;
  assign n20779 = n12397 & n13831 ;
  assign n20780 = n14534 ^ n2027 ^ 1'b0 ;
  assign n20781 = n19099 ^ n2978 ^ 1'b0 ;
  assign n20782 = n3552 & n10650 ;
  assign n20783 = ~n10360 & n16409 ;
  assign n20784 = n775 & ~n1472 ;
  assign n20785 = n20784 ^ n8714 ^ 1'b0 ;
  assign n20786 = n5048 & n20785 ;
  assign n20787 = n20786 ^ n15288 ^ 1'b0 ;
  assign n20788 = n4749 | n20787 ;
  assign n20789 = n663 & n9490 ;
  assign n20790 = n16572 ^ n9368 ^ 1'b0 ;
  assign n20791 = ~n7326 & n9081 ;
  assign n20792 = n20791 ^ n330 ^ 1'b0 ;
  assign n20793 = n4618 & n5099 ;
  assign n20794 = n20793 ^ n934 ^ 1'b0 ;
  assign n20795 = n3183 & n20794 ;
  assign n20800 = n984 & n2072 ;
  assign n20801 = n4048 & n20800 ;
  assign n20802 = n20801 ^ n142 ^ 1'b0 ;
  assign n20803 = n2657 & n20802 ;
  assign n20804 = ~n3489 & n20803 ;
  assign n20805 = n20804 ^ n15596 ^ 1'b0 ;
  assign n20796 = n840 & ~n11174 ;
  assign n20797 = n1867 | n20796 ;
  assign n20798 = n1523 & ~n20797 ;
  assign n20799 = n20480 | n20798 ;
  assign n20806 = n20805 ^ n20799 ^ 1'b0 ;
  assign n20807 = n20795 | n20806 ;
  assign n20808 = n4878 & ~n8175 ;
  assign n20809 = n3616 | n20808 ;
  assign n20810 = n1994 & n2433 ;
  assign n20811 = ~n1982 & n20810 ;
  assign n20812 = n9075 & ~n20811 ;
  assign n20813 = n19870 & ~n20812 ;
  assign n20814 = ~n1388 & n3178 ;
  assign n20815 = n1884 | n2885 ;
  assign n20816 = n20815 ^ n12098 ^ 1'b0 ;
  assign n20817 = ~n9491 & n20816 ;
  assign n20818 = ~n16585 & n20817 ;
  assign n20819 = ~n37 & n1649 ;
  assign n20820 = ( n3635 & ~n10988 ) | ( n3635 & n11678 ) | ( ~n10988 & n11678 ) ;
  assign n20821 = n1831 & ~n10203 ;
  assign n20822 = n20821 ^ n5625 ^ 1'b0 ;
  assign n20823 = n3227 | n14911 ;
  assign n20824 = n2866 & ~n11613 ;
  assign n20825 = n10437 & ~n20824 ;
  assign n20826 = ~n20823 & n20825 ;
  assign n20830 = n5739 ^ n5737 ^ n3929 ;
  assign n20831 = n20830 ^ n9523 ^ 1'b0 ;
  assign n20832 = n12302 | n20831 ;
  assign n20827 = n4662 ^ n3885 ^ 1'b0 ;
  assign n20828 = n2900 & n20827 ;
  assign n20829 = ~n198 & n20828 ;
  assign n20833 = n20832 ^ n20829 ^ 1'b0 ;
  assign n20834 = n2382 | n14734 ;
  assign n20835 = n20834 ^ n3431 ^ 1'b0 ;
  assign n20836 = ~n3131 & n6608 ;
  assign n20837 = n20836 ^ n405 ^ 1'b0 ;
  assign n20838 = ( n466 & n6580 ) | ( n466 & ~n20837 ) | ( n6580 & ~n20837 ) ;
  assign n20839 = n20838 ^ n8411 ^ n592 ;
  assign n20840 = n20839 ^ n3200 ^ 1'b0 ;
  assign n20841 = n20835 | n20840 ;
  assign n20842 = n963 | n1522 ;
  assign n20843 = n12716 & n20842 ;
  assign n20844 = n833 & n20843 ;
  assign n20845 = n20844 ^ n20728 ^ 1'b0 ;
  assign n20846 = n3512 & n20845 ;
  assign n20847 = n8599 ^ n5443 ^ 1'b0 ;
  assign n20848 = n12937 & ~n20847 ;
  assign n20849 = n6626 ^ n666 ^ 1'b0 ;
  assign n20850 = n7994 & n8450 ;
  assign n20851 = n304 | n17576 ;
  assign n20852 = n304 & ~n20851 ;
  assign n20853 = n191 | n20852 ;
  assign n20854 = n20852 & ~n20853 ;
  assign n20855 = n89 & ~n20854 ;
  assign n20856 = ~n89 & n20855 ;
  assign n20857 = n109 & n283 ;
  assign n20858 = n14015 & n20857 ;
  assign n20859 = n20856 | n20858 ;
  assign n20860 = n20856 & ~n20859 ;
  assign n20867 = n471 | n2928 ;
  assign n20868 = n471 & ~n20867 ;
  assign n20869 = n6392 & ~n20868 ;
  assign n20861 = n17 & n101 ;
  assign n20862 = ~n101 & n20861 ;
  assign n20863 = n1236 & n20862 ;
  assign n20864 = n3627 & n20863 ;
  assign n20865 = n9307 & ~n20864 ;
  assign n20866 = ~n9307 & n20865 ;
  assign n20870 = n20869 ^ n20866 ^ 1'b0 ;
  assign n20871 = ~n20860 & n20870 ;
  assign n20872 = n11209 | n18312 ;
  assign n20873 = n11259 ^ n7492 ^ 1'b0 ;
  assign n20874 = n7143 & n16897 ;
  assign n20875 = ~n107 & n20874 ;
  assign n20876 = x8 & n19 ;
  assign n20877 = n141 | n20876 ;
  assign n20878 = n12602 & ~n20877 ;
  assign n20879 = n487 & ~n20878 ;
  assign n20880 = n20878 & n20879 ;
  assign n20881 = n142 | n20880 ;
  assign n20882 = n20880 & ~n20881 ;
  assign n20883 = n3837 | n20882 ;
  assign n20884 = n20882 & ~n20883 ;
  assign n20885 = n5864 & ~n20884 ;
  assign n20886 = ~n14463 & n20885 ;
  assign n20887 = n20886 ^ n15458 ^ 1'b0 ;
  assign n20888 = n4211 ^ n1132 ^ 1'b0 ;
  assign n20889 = n19807 & ~n20888 ;
  assign n20890 = n20889 ^ n4485 ^ 1'b0 ;
  assign n20891 = n13832 & ~n20890 ;
  assign n20892 = n20887 & n20891 ;
  assign n20895 = n7564 | n17673 ;
  assign n20896 = n367 & n13417 ;
  assign n20897 = n20896 ^ n3001 ^ 1'b0 ;
  assign n20898 = ~n17944 & n20897 ;
  assign n20899 = ~n20895 & n20898 ;
  assign n20893 = n16171 ^ n6014 ^ 1'b0 ;
  assign n20894 = n3096 & ~n20893 ;
  assign n20900 = n20899 ^ n20894 ^ n9542 ;
  assign n20901 = n15470 ^ n3921 ^ 1'b0 ;
  assign n20902 = n7424 & ~n20901 ;
  assign n20903 = n20902 ^ n817 ^ 1'b0 ;
  assign n20904 = n20903 ^ n11981 ^ 1'b0 ;
  assign n20905 = n310 & ~n8577 ;
  assign n20906 = n8577 & n20905 ;
  assign n20907 = n11141 | n20906 ;
  assign n20908 = n20906 & ~n20907 ;
  assign n20909 = n30 | n66 ;
  assign n20910 = n30 & ~n20909 ;
  assign n20911 = n55 | n164 ;
  assign n20912 = n164 & ~n20911 ;
  assign n20913 = n20910 | n20912 ;
  assign n20914 = n20910 & ~n20913 ;
  assign n20916 = n98 & ~n117 ;
  assign n20917 = n117 & n20916 ;
  assign n20918 = n20917 ^ x3 ^ 1'b0 ;
  assign n20915 = ~n336 & n15727 ;
  assign n20919 = n20918 ^ n20915 ^ 1'b0 ;
  assign n20920 = n661 | n20919 ;
  assign n20921 = n20914 & ~n20920 ;
  assign n20922 = n14015 | n20921 ;
  assign n20923 = n14015 & ~n20922 ;
  assign n20924 = n12193 & ~n20923 ;
  assign n20925 = ~n12193 & n20924 ;
  assign n20926 = x9 & ~n228 ;
  assign n20927 = ~x9 & n20926 ;
  assign n20928 = n937 | n20927 ;
  assign n20929 = n20927 & ~n20928 ;
  assign n20930 = n107 & ~n146 ;
  assign n20931 = ~n107 & n20930 ;
  assign n20932 = n556 & ~n20931 ;
  assign n20933 = n149 & ~n20932 ;
  assign n20934 = n20929 & n20933 ;
  assign n20935 = n46 & ~n687 ;
  assign n20936 = n687 & n20935 ;
  assign n20937 = n20936 ^ n694 ^ 1'b0 ;
  assign n20938 = n20934 | n20937 ;
  assign n20939 = n20925 | n20938 ;
  assign n20940 = n20925 & ~n20939 ;
  assign n20941 = n20908 | n20940 ;
  assign n20942 = n20941 ^ n20499 ^ 1'b0 ;
  assign n20943 = ~n13242 & n13629 ;
  assign n20944 = ~n5376 & n6524 ;
  assign n20945 = n6718 & n20944 ;
  assign n20946 = n227 | n15656 ;
  assign n20947 = n18201 ^ n17492 ^ 1'b0 ;
  assign n20948 = n6078 | n6611 ;
  assign n20949 = ~n5821 & n9719 ;
  assign n20950 = n6269 & n20949 ;
  assign n20951 = n461 & n20950 ;
  assign n20952 = n11821 ^ n9934 ^ n3349 ;
  assign n20953 = ~n8022 & n20952 ;
  assign n20954 = n20953 ^ n4042 ^ 1'b0 ;
  assign n20955 = n567 & n17229 ;
  assign n20956 = n3724 & n8409 ;
  assign n20957 = n4155 ^ n2049 ^ 1'b0 ;
  assign n20958 = n14478 ^ x1 ^ 1'b0 ;
  assign n20959 = n4439 | n20958 ;
  assign n20960 = ~n14706 & n19013 ;
  assign n20961 = n20960 ^ n15915 ^ 1'b0 ;
  assign n20962 = n17546 ^ n9880 ^ 1'b0 ;
  assign n20963 = n2696 & n17264 ;
  assign n20964 = n20963 ^ n19050 ^ 1'b0 ;
  assign n20966 = n3374 & ~n3640 ;
  assign n20967 = ~n2650 & n20966 ;
  assign n20965 = n8948 & n10171 ;
  assign n20968 = n20967 ^ n20965 ^ n20323 ;
  assign n20969 = n14081 ^ n9092 ^ 1'b0 ;
  assign n20970 = n3270 & ~n13769 ;
  assign n20971 = n1914 & n6316 ;
  assign n20972 = n1237 | n20971 ;
  assign n20973 = n1825 & n10862 ;
  assign n20974 = n14303 & n20973 ;
  assign n20975 = n1705 | n8244 ;
  assign n20976 = n20975 ^ n4647 ^ 1'b0 ;
  assign n20977 = ~n9145 & n13225 ;
  assign n20978 = n20977 ^ n3632 ^ 1'b0 ;
  assign n20987 = n1019 & ~n5038 ;
  assign n20983 = ~n432 & n477 ;
  assign n20984 = n432 & n20983 ;
  assign n20985 = ~n1851 & n20984 ;
  assign n20979 = n2478 | n4885 ;
  assign n20980 = n4885 & ~n20979 ;
  assign n20981 = n5831 | n19363 ;
  assign n20982 = n20980 & ~n20981 ;
  assign n20986 = n20985 ^ n20982 ^ 1'b0 ;
  assign n20988 = n20987 ^ n20986 ^ 1'b0 ;
  assign n20989 = n20978 | n20988 ;
  assign n20990 = ~n7188 & n20948 ;
  assign n20991 = n14311 ^ n1325 ^ 1'b0 ;
  assign n20992 = n20506 | n20991 ;
  assign n20993 = n9750 ^ n9581 ^ 1'b0 ;
  assign n20994 = n19302 & n20993 ;
  assign n20995 = n6361 ^ n4161 ^ 1'b0 ;
  assign n20996 = n20994 & n20995 ;
  assign n20997 = n1310 | n9341 ;
  assign n20998 = n20997 ^ n7767 ^ 1'b0 ;
  assign n20999 = n534 | n5583 ;
  assign n21000 = n3627 ^ n2774 ^ 1'b0 ;
  assign n21001 = ~n231 & n21000 ;
  assign n21002 = n395 & ~n964 ;
  assign n21003 = n2817 ^ n107 ^ 1'b0 ;
  assign n21004 = n21002 & ~n21003 ;
  assign n21005 = n364 & n21004 ;
  assign n21006 = n1891 ^ n1810 ^ 1'b0 ;
  assign n21007 = ~n444 & n21006 ;
  assign n21008 = n21007 ^ n2252 ^ 1'b0 ;
  assign n21009 = n15045 ^ n5828 ^ 1'b0 ;
  assign n21010 = n15093 & ~n21009 ;
  assign n21011 = ( n4308 & ~n6915 ) | ( n4308 & n21010 ) | ( ~n6915 & n21010 ) ;
  assign n21012 = ~n13661 & n18175 ;
  assign n21013 = n21012 ^ n55 ^ 1'b0 ;
  assign n21014 = ~n5076 & n21013 ;
  assign n21015 = ~n5808 & n19713 ;
  assign n21016 = n9695 ^ n6188 ^ n4020 ;
  assign n21017 = n10867 & n21016 ;
  assign n21018 = ~n1958 & n2537 ;
  assign n21019 = n21018 ^ n4843 ^ 1'b0 ;
  assign n21020 = n799 ^ n715 ^ 1'b0 ;
  assign n21021 = ~n11768 & n21020 ;
  assign n21022 = n3873 ^ n1530 ^ 1'b0 ;
  assign n21023 = n8453 & ~n21022 ;
  assign n21024 = n21023 ^ n18058 ^ 1'b0 ;
  assign n21025 = ~n16527 & n21024 ;
  assign n21026 = n2352 | n11483 ;
  assign n21027 = n14751 | n21026 ;
  assign n21028 = ~n3183 & n21027 ;
  assign n21029 = ~n4600 & n21028 ;
  assign n21030 = ~n6660 & n10219 ;
  assign n21031 = n21030 ^ n35 ^ 1'b0 ;
  assign n21032 = n715 & ~n21031 ;
  assign n21033 = n21032 ^ n430 ^ 1'b0 ;
  assign n21034 = n10983 ^ n7984 ^ 1'b0 ;
  assign n21035 = n5261 & n21034 ;
  assign n21036 = n21035 ^ n6055 ^ 1'b0 ;
  assign n21037 = ~n14200 & n21036 ;
  assign n21038 = n4221 & n20323 ;
  assign n21039 = n21038 ^ n1382 ^ 1'b0 ;
  assign n21040 = ~n11159 & n12530 ;
  assign n21041 = ~n13080 & n21040 ;
  assign n21042 = n3498 & ~n5326 ;
  assign n21043 = ~n1731 & n9994 ;
  assign n21044 = n2305 | n20142 ;
  assign n21045 = n21044 ^ n1947 ^ 1'b0 ;
  assign n21047 = n2064 & n10194 ;
  assign n21046 = n9032 & n10538 ;
  assign n21048 = n21047 ^ n21046 ^ 1'b0 ;
  assign n21049 = ~n8411 & n21048 ;
  assign n21050 = n10195 | n18383 ;
  assign n21051 = ~n10156 & n21050 ;
  assign n21052 = n8070 ^ n315 ^ 1'b0 ;
  assign n21053 = n254 & ~n21052 ;
  assign n21054 = n19 & n2380 ;
  assign n21055 = ~n21053 & n21054 ;
  assign n21056 = ~n4560 & n10940 ;
  assign n21057 = n8904 & n12014 ;
  assign n21058 = n119 | n2681 ;
  assign n21059 = n878 & ~n21058 ;
  assign n21060 = n21059 ^ n15756 ^ 1'b0 ;
  assign n21061 = n4590 & n21060 ;
  assign n21062 = n16643 ^ n2154 ^ 1'b0 ;
  assign n21063 = n55 & n1598 ;
  assign n21064 = ~n8617 & n18106 ;
  assign n21065 = n2937 & n21064 ;
  assign n21066 = ~n6477 & n21065 ;
  assign n21067 = n21066 ^ n258 ^ 1'b0 ;
  assign n21068 = n1375 & ~n21067 ;
  assign n21069 = n1878 ^ n646 ^ 1'b0 ;
  assign n21071 = n30 | n246 ;
  assign n21072 = n785 & ~n21071 ;
  assign n21073 = n1027 | n1763 ;
  assign n21074 = n21072 & ~n21073 ;
  assign n21070 = ~n17281 & n21049 ;
  assign n21075 = n21074 ^ n21070 ^ 1'b0 ;
  assign n21076 = n1704 & ~n18497 ;
  assign n21077 = n2705 & n6809 ;
  assign n21078 = n2353 & n21077 ;
  assign n21079 = n13169 | n18828 ;
  assign n21080 = n9336 | n21079 ;
  assign n21081 = n21078 | n21080 ;
  assign n21082 = n1670 & n7498 ;
  assign n21083 = n832 | n21082 ;
  assign n21084 = ~n17750 & n21083 ;
  assign n21085 = ~n159 & n193 ;
  assign n21086 = n21085 ^ n9287 ^ 1'b0 ;
  assign n21087 = n18956 ^ n3010 ^ 1'b0 ;
  assign n21088 = n2135 & ~n18592 ;
  assign n21089 = ~n304 & n6476 ;
  assign n21090 = n21089 ^ n16320 ^ 1'b0 ;
  assign n21091 = n6619 ^ n236 ^ 1'b0 ;
  assign n21092 = ~n3995 & n4063 ;
  assign n21093 = n6810 & n21092 ;
  assign n21094 = n21093 ^ n5452 ^ 1'b0 ;
  assign n21095 = n506 & ~n13939 ;
  assign n21096 = n21094 & n21095 ;
  assign n21097 = n3437 & n11658 ;
  assign n21098 = ~n3364 & n21097 ;
  assign n21105 = n9994 & ~n11384 ;
  assign n21106 = ~n2574 & n21105 ;
  assign n21107 = n7607 | n21106 ;
  assign n21108 = n942 | n21107 ;
  assign n21099 = ~n6194 & n7960 ;
  assign n21100 = n21099 ^ n6711 ^ 1'b0 ;
  assign n21101 = n8033 | n14226 ;
  assign n21102 = ~n1217 & n21101 ;
  assign n21103 = n3646 & n21102 ;
  assign n21104 = n21100 | n21103 ;
  assign n21109 = n21108 ^ n21104 ^ 1'b0 ;
  assign n21111 = n2720 & n8062 ;
  assign n21110 = ~n6586 & n14192 ;
  assign n21112 = n21111 ^ n21110 ^ 1'b0 ;
  assign n21113 = n8922 ^ n5283 ^ 1'b0 ;
  assign n21114 = n7996 ^ n5063 ^ 1'b0 ;
  assign n21115 = n16058 ^ n566 ^ 1'b0 ;
  assign n21116 = n5245 & n21115 ;
  assign n21117 = n1666 & n3411 ;
  assign n21118 = n594 | n21117 ;
  assign n21119 = n21118 ^ n764 ^ 1'b0 ;
  assign n21120 = n157 & n21119 ;
  assign n21121 = n21120 ^ n1067 ^ 1'b0 ;
  assign n21122 = ~n86 & n6732 ;
  assign n21123 = n21122 ^ n19886 ^ 1'b0 ;
  assign n21124 = n16423 ^ n2435 ^ 1'b0 ;
  assign n21125 = n4115 & n9914 ;
  assign n21126 = n3940 & n21125 ;
  assign n21127 = n2023 & n13359 ;
  assign n21128 = n21127 ^ n3449 ^ 1'b0 ;
  assign n21129 = n4199 & ~n21128 ;
  assign n21130 = ~n3859 & n7810 ;
  assign n21131 = n1902 & ~n13836 ;
  assign n21132 = n13875 & ~n21131 ;
  assign n21133 = n5808 | n10751 ;
  assign n21134 = n21133 ^ n15397 ^ 1'b0 ;
  assign n21135 = n1252 & ~n10588 ;
  assign n21136 = n21135 ^ n3243 ^ 1'b0 ;
  assign n21137 = ( n1849 & n14932 ) | ( n1849 & n21136 ) | ( n14932 & n21136 ) ;
  assign n21138 = ( n2376 & n21134 ) | ( n2376 & n21137 ) | ( n21134 & n21137 ) ;
  assign n21139 = n10223 & n12509 ;
  assign n21140 = n2524 ^ n197 ^ 1'b0 ;
  assign n21141 = n21140 ^ n18305 ^ 1'b0 ;
  assign n21142 = n16977 ^ n3175 ^ 1'b0 ;
  assign n21143 = n13869 | n21142 ;
  assign n21144 = n1388 & ~n12708 ;
  assign n21145 = n19901 ^ n384 ^ 1'b0 ;
  assign n21146 = ~n4655 & n6026 ;
  assign n21147 = n3969 & n4740 ;
  assign n21148 = n7360 & n21147 ;
  assign n21149 = n10282 & ~n13250 ;
  assign n21150 = n4117 & ~n8111 ;
  assign n21151 = n11433 ^ n9316 ^ n1183 ;
  assign n21152 = n21150 & ~n21151 ;
  assign n21153 = n21152 ^ n5256 ^ 1'b0 ;
  assign n21154 = n15122 ^ n1884 ^ 1'b0 ;
  assign n21155 = n4078 | n21154 ;
  assign n21156 = n6021 | n21155 ;
  assign n21157 = n6353 | n19119 ;
  assign n21158 = n3032 | n5164 ;
  assign n21159 = ~n55 & n14824 ;
  assign n21160 = n21159 ^ n14596 ^ 1'b0 ;
  assign n21161 = n21158 & ~n21160 ;
  assign n21162 = n21157 & n21161 ;
  assign n21166 = ~n4874 & n12450 ;
  assign n21167 = ~n8037 & n21166 ;
  assign n21163 = n1031 ^ n461 ^ 1'b0 ;
  assign n21164 = n7683 & ~n21163 ;
  assign n21165 = n11760 & n21164 ;
  assign n21168 = n21167 ^ n21165 ^ 1'b0 ;
  assign n21169 = n7148 | n21168 ;
  assign n21170 = n11631 ^ n1007 ^ 1'b0 ;
  assign n21171 = n11965 ^ n6907 ^ 1'b0 ;
  assign n21172 = ~n3406 & n21171 ;
  assign n21173 = ~n7714 & n21172 ;
  assign n21174 = n2209 | n2687 ;
  assign n21175 = ~n2733 & n20553 ;
  assign n21176 = n4024 & ~n5694 ;
  assign n21177 = n5694 & n21176 ;
  assign n21179 = n3681 & n20409 ;
  assign n21180 = ~n3681 & n21179 ;
  assign n21178 = n804 & ~n15210 ;
  assign n21181 = n21180 ^ n21178 ^ 1'b0 ;
  assign n21182 = ~n21177 & n21181 ;
  assign n21183 = n21177 & n21182 ;
  assign n21184 = n339 & n1194 ;
  assign n21185 = ~n1194 & n21184 ;
  assign n21186 = n20615 | n21185 ;
  assign n21187 = n20615 & ~n21186 ;
  assign n21188 = n21183 | n21187 ;
  assign n21189 = n342 | n21188 ;
  assign n21190 = n3611 | n18120 ;
  assign n21191 = n21190 ^ n7417 ^ 1'b0 ;
  assign n21192 = ~n3663 & n15673 ;
  assign n21193 = n21192 ^ n520 ^ 1'b0 ;
  assign n21194 = n21191 & ~n21193 ;
  assign n21195 = n21194 ^ n11150 ^ 1'b0 ;
  assign n21196 = n6687 ^ n527 ^ 1'b0 ;
  assign n21197 = n1306 | n18634 ;
  assign n21198 = n21197 ^ n11074 ^ 1'b0 ;
  assign n21199 = n7622 & n11041 ;
  assign n21200 = n466 & ~n21199 ;
  assign n21201 = ~n8648 & n21200 ;
  assign n21202 = n3586 & ~n18579 ;
  assign n21203 = ~n1777 & n6332 ;
  assign n21204 = n51 & ~n13786 ;
  assign n21205 = n7249 | n21204 ;
  assign n21206 = n21203 | n21205 ;
  assign n21207 = n359 & ~n21206 ;
  assign n21208 = n3368 & ~n9330 ;
  assign n21209 = n3180 & ~n5842 ;
  assign n21210 = n20828 ^ n14464 ^ 1'b0 ;
  assign n21211 = n17342 & ~n21210 ;
  assign n21212 = n1095 & ~n12100 ;
  assign n21213 = n21212 ^ n8195 ^ 1'b0 ;
  assign n21214 = n13028 & n21213 ;
  assign n21215 = ~n6710 & n21214 ;
  assign n21216 = n21215 ^ n14662 ^ 1'b0 ;
  assign n21217 = n14996 ^ n9055 ^ 1'b0 ;
  assign n21218 = ~n6519 & n14540 ;
  assign n21219 = n21217 & n21218 ;
  assign n21220 = ( ~n1526 & n3803 ) | ( ~n1526 & n21219 ) | ( n3803 & n21219 ) ;
  assign n21221 = n4087 ^ n977 ^ 1'b0 ;
  assign n21222 = n21221 ^ n16822 ^ 1'b0 ;
  assign n21223 = n11557 ^ n759 ^ 1'b0 ;
  assign n21224 = ~n5934 & n16708 ;
  assign n21225 = n8225 & ~n9038 ;
  assign n21226 = n19450 ^ n16190 ^ 1'b0 ;
  assign n21227 = n21225 | n21226 ;
  assign n21228 = n6953 & ~n15674 ;
  assign n21229 = n21228 ^ n12544 ^ 1'b0 ;
  assign n21230 = n21229 ^ n19406 ^ 1'b0 ;
  assign n21231 = n1851 & ~n21230 ;
  assign n21232 = n13110 ^ n8910 ^ 1'b0 ;
  assign n21233 = n8050 ^ n330 ^ 1'b0 ;
  assign n21234 = n3580 | n21233 ;
  assign n21237 = n15 | n2642 ;
  assign n21236 = n3899 | n9821 ;
  assign n21238 = n21237 ^ n21236 ^ 1'b0 ;
  assign n21239 = n21238 ^ n448 ^ 1'b0 ;
  assign n21235 = n2286 & n10761 ;
  assign n21240 = n21239 ^ n21235 ^ 1'b0 ;
  assign n21241 = n21240 ^ n9038 ^ 1'b0 ;
  assign n21242 = n9039 & n11533 ;
  assign n21243 = ~n6493 & n7599 ;
  assign n21244 = n1098 | n9364 ;
  assign n21245 = ~n2120 & n11003 ;
  assign n21246 = n4590 ^ n3485 ^ 1'b0 ;
  assign n21247 = n9195 | n21246 ;
  assign n21248 = n21247 ^ n19607 ^ 1'b0 ;
  assign n21249 = ~n1595 & n3014 ;
  assign n21250 = n837 & n21249 ;
  assign n21251 = n18229 ^ n1872 ^ 1'b0 ;
  assign n21252 = ~n14850 & n21251 ;
  assign n21253 = ~n1270 & n4898 ;
  assign n21254 = n18950 | n21253 ;
  assign n21255 = n1505 & ~n17649 ;
  assign n21256 = n14751 ^ n2050 ^ 1'b0 ;
  assign n21257 = ~n200 & n21256 ;
  assign n21258 = n16820 & ~n21257 ;
  assign n21270 = ~n604 & n996 ;
  assign n21271 = n604 & n21270 ;
  assign n21269 = n7539 ^ n4655 ^ 1'b0 ;
  assign n21259 = ~n177 & n809 ;
  assign n21260 = n177 & n21259 ;
  assign n21261 = n21260 ^ n6349 ^ 1'b0 ;
  assign n21262 = n257 | n1239 ;
  assign n21263 = n1239 & ~n21262 ;
  assign n21264 = ~n1295 & n21263 ;
  assign n21265 = n266 & n21264 ;
  assign n21266 = n21265 ^ x0 ^ 1'b0 ;
  assign n21267 = ~n215 & n21266 ;
  assign n21268 = n21261 & n21267 ;
  assign n21272 = n21271 ^ n21269 ^ n21268 ;
  assign n21273 = n8073 ^ n1065 ^ 1'b0 ;
  assign n21274 = n646 ^ n43 ^ 1'b0 ;
  assign n21275 = n5495 & ~n21274 ;
  assign n21276 = n2354 | n3036 ;
  assign n21277 = n21276 ^ n11768 ^ 1'b0 ;
  assign n21278 = n21275 & n21277 ;
  assign n21279 = n2549 & n21278 ;
  assign n21280 = n21279 ^ n1571 ^ 1'b0 ;
  assign n21281 = n177 & n11164 ;
  assign n21282 = n20099 ^ n3739 ^ 1'b0 ;
  assign n21283 = n497 & n21282 ;
  assign n21284 = n9242 & n13250 ;
  assign n21285 = ~n7265 & n14435 ;
  assign n21286 = ~n748 & n21285 ;
  assign n21287 = n1856 & ~n3219 ;
  assign n21288 = ~n10417 & n21287 ;
  assign n21289 = n19095 ^ n12359 ^ 1'b0 ;
  assign n21290 = ~n3931 & n8628 ;
  assign n21291 = n12898 ^ n495 ^ 1'b0 ;
  assign n21292 = n8755 & n21291 ;
  assign n21293 = n15269 ^ n12168 ^ 1'b0 ;
  assign n21294 = n3841 & n21293 ;
  assign n21295 = n11692 & ~n21294 ;
  assign n21296 = ~n6335 & n21295 ;
  assign n21297 = n21296 ^ n7821 ^ 1'b0 ;
  assign n21298 = n4623 & n21297 ;
  assign n21299 = n5796 & ~n11258 ;
  assign n21300 = n566 | n21299 ;
  assign n21317 = n1166 & n1529 ;
  assign n21318 = ~n1166 & n21317 ;
  assign n21301 = n11829 & ~n11866 ;
  assign n21302 = ~n14177 & n21301 ;
  assign n21307 = n7229 & ~n13320 ;
  assign n21308 = n390 & n3097 ;
  assign n21309 = ~n390 & n21308 ;
  assign n21310 = ~n1100 & n4326 ;
  assign n21311 = n21309 & n21310 ;
  assign n21312 = ~n1090 & n21311 ;
  assign n21313 = n21307 & n21312 ;
  assign n21314 = n8208 & n21313 ;
  assign n21303 = n5312 ^ n4390 ^ 1'b0 ;
  assign n21304 = n194 & n7720 ;
  assign n21305 = ~n21303 & n21304 ;
  assign n21306 = n21305 ^ n2227 ^ 1'b0 ;
  assign n21315 = n21314 ^ n21306 ^ 1'b0 ;
  assign n21316 = ~n21302 & n21315 ;
  assign n21319 = n21318 ^ n21316 ^ 1'b0 ;
  assign n21320 = n2869 | n21319 ;
  assign n21321 = n9086 ^ n4657 ^ 1'b0 ;
  assign n21322 = n21321 ^ n21050 ^ 1'b0 ;
  assign n21323 = n101 & n300 ;
  assign n21324 = n21323 ^ n3329 ^ 1'b0 ;
  assign n21325 = n21324 ^ n11895 ^ n9592 ;
  assign n21326 = n6272 & ~n21325 ;
  assign n21327 = n21326 ^ n8263 ^ 1'b0 ;
  assign n21328 = ~n13119 & n21327 ;
  assign n21329 = n1640 & n2017 ;
  assign n21330 = n3005 | n12227 ;
  assign n21331 = n21330 ^ n18308 ^ n3127 ;
  assign n21332 = n9209 & n13459 ;
  assign n21333 = n21332 ^ n1193 ^ 1'b0 ;
  assign n21334 = n19626 ^ n7694 ^ 1'b0 ;
  assign n21335 = n21333 & ~n21334 ;
  assign n21336 = n3352 ^ n1597 ^ 1'b0 ;
  assign n21337 = n761 & ~n21336 ;
  assign n21338 = ( n4245 & n6011 ) | ( n4245 & ~n21337 ) | ( n6011 & ~n21337 ) ;
  assign n21339 = n1838 ^ n1143 ^ 1'b0 ;
  assign n21340 = ~n47 & n21339 ;
  assign n21341 = n21340 ^ n18057 ^ 1'b0 ;
  assign n21342 = n21338 & ~n21341 ;
  assign n21343 = n6907 ^ n4929 ^ 1'b0 ;
  assign n21344 = n11319 & ~n21343 ;
  assign n21345 = n21344 ^ n16231 ^ 1'b0 ;
  assign n21346 = n21345 ^ n18199 ^ n3219 ;
  assign n21348 = n12028 ^ n1227 ^ 1'b0 ;
  assign n21349 = n2824 | n21348 ;
  assign n21347 = n8047 | n8512 ;
  assign n21350 = n21349 ^ n21347 ^ 1'b0 ;
  assign n21353 = n830 & n3125 ;
  assign n21351 = n1672 ^ n1622 ^ 1'b0 ;
  assign n21352 = n491 & n21351 ;
  assign n21354 = n21353 ^ n21352 ^ 1'b0 ;
  assign n21355 = ~n16450 & n21354 ;
  assign n21357 = n497 & n1207 ;
  assign n21356 = n5260 | n12855 ;
  assign n21358 = n21357 ^ n21356 ^ n6981 ;
  assign n21359 = ~n6060 & n10572 ;
  assign n21360 = ( n11891 & ~n13255 ) | ( n11891 & n18046 ) | ( ~n13255 & n18046 ) ;
  assign n21361 = n4552 | n21360 ;
  assign n21362 = n2721 & ~n2779 ;
  assign n21365 = n9778 & ~n9827 ;
  assign n21363 = n9211 ^ n6496 ^ n3767 ;
  assign n21364 = n13106 & ~n21363 ;
  assign n21366 = n21365 ^ n21364 ^ 1'b0 ;
  assign n21367 = ~n15035 & n18133 ;
  assign n21368 = ~n17250 & n21367 ;
  assign n21369 = n8466 ^ n6135 ^ 1'b0 ;
  assign n21370 = ~n10318 & n21369 ;
  assign n21371 = ~n8932 & n10743 ;
  assign n21372 = n16138 ^ n8288 ^ 1'b0 ;
  assign n21373 = n12669 ^ n6711 ^ 1'b0 ;
  assign n21374 = n21373 ^ n15688 ^ 1'b0 ;
  assign n21375 = n4392 & n21374 ;
  assign n21376 = n213 | n20240 ;
  assign n21377 = n21376 ^ n10105 ^ 1'b0 ;
  assign n21378 = n8764 | n21377 ;
  assign n21379 = ~n3040 & n21014 ;
  assign n21380 = n21379 ^ n11824 ^ 1'b0 ;
  assign n21381 = n2921 & n15792 ;
  assign n21382 = ~n20554 & n21381 ;
  assign n21383 = n532 & n18858 ;
  assign n21384 = n21383 ^ n5842 ^ 1'b0 ;
  assign n21385 = ~n7217 & n8836 ;
  assign n21386 = n16338 ^ n7967 ^ 1'b0 ;
  assign n21387 = n20516 & ~n21386 ;
  assign n21388 = n2495 & n6051 ;
  assign n21389 = n21388 ^ n6067 ^ 1'b0 ;
  assign n21390 = n962 & ~n21389 ;
  assign n21391 = n13256 & n21390 ;
  assign n21392 = n4000 ^ n1499 ^ 1'b0 ;
  assign n21393 = n4228 & ~n21392 ;
  assign n21394 = n21393 ^ n1325 ^ 1'b0 ;
  assign n21395 = n21394 ^ n12306 ^ 1'b0 ;
  assign n21396 = n5543 | n21395 ;
  assign n21397 = n257 & ~n21396 ;
  assign n21398 = ~n5241 & n5525 ;
  assign n21399 = n21398 ^ n142 ^ 1'b0 ;
  assign n21400 = n19550 ^ n5386 ^ 1'b0 ;
  assign n21401 = n21399 & ~n21400 ;
  assign n21402 = n11021 & ~n12315 ;
  assign n21403 = n5761 ^ n509 ^ 1'b0 ;
  assign n21404 = n883 & n21403 ;
  assign n21405 = n21404 ^ n12455 ^ 1'b0 ;
  assign n21406 = n19117 ^ n13522 ^ 1'b0 ;
  assign n21407 = ~n10099 & n21406 ;
  assign n21408 = n21407 ^ n8010 ^ 1'b0 ;
  assign n21409 = n20676 & n21408 ;
  assign n21410 = n1760 | n12518 ;
  assign n21411 = n3567 & ~n4416 ;
  assign n21412 = n2316 & ~n21411 ;
  assign n21413 = n17364 ^ n9509 ^ n4976 ;
  assign n21414 = n10588 & n21413 ;
  assign n21415 = n6588 & n12511 ;
  assign n21416 = ~n6588 & n21415 ;
  assign n21417 = n3365 & ~n11967 ;
  assign n21418 = ~n839 & n21417 ;
  assign n21419 = n7529 ^ n97 ^ 1'b0 ;
  assign n21420 = n236 | n21419 ;
  assign n21421 = n21420 ^ n2092 ^ 1'b0 ;
  assign n21422 = n6242 & ~n7605 ;
  assign n21423 = ( ~n2204 & n21421 ) | ( ~n2204 & n21422 ) | ( n21421 & n21422 ) ;
  assign n21424 = ~n12391 & n21423 ;
  assign n21425 = n2987 | n3156 ;
  assign n21426 = n21425 ^ n3794 ^ 1'b0 ;
  assign n21427 = n259 | n2424 ;
  assign n21428 = n3771 ^ n2252 ^ 1'b0 ;
  assign n21429 = ~n3434 & n21428 ;
  assign n21430 = n10982 & n21429 ;
  assign n21431 = n1385 & ~n21430 ;
  assign n21432 = n9829 & n21431 ;
  assign n21433 = n4093 & ~n12948 ;
  assign n21434 = n21433 ^ n12645 ^ 1'b0 ;
  assign n21435 = n191 | n21434 ;
  assign n21436 = n1329 ^ n169 ^ 1'b0 ;
  assign n21437 = ~n4763 & n21436 ;
  assign n21438 = n66 & ~n169 ;
  assign n21439 = n169 & n21438 ;
  assign n21440 = ~n20663 & n21439 ;
  assign n21441 = n2102 & ~n21440 ;
  assign n21442 = ~n2102 & n21441 ;
  assign n21443 = n9326 | n10337 ;
  assign n21444 = n21443 ^ n2817 ^ 1'b0 ;
  assign n21445 = ~n21442 & n21444 ;
  assign n21446 = n21442 & n21445 ;
  assign n21447 = n3793 ^ n37 ^ 1'b0 ;
  assign n21448 = n8271 ^ n7475 ^ 1'b0 ;
  assign n21449 = n12242 & ~n21448 ;
  assign n21450 = n2038 & n5222 ;
  assign n21451 = ~n1054 & n9737 ;
  assign n21452 = ~n3183 & n21451 ;
  assign n21453 = ~n55 & n6933 ;
  assign n21454 = n11008 & ~n20890 ;
  assign n21455 = n21453 & n21454 ;
  assign n21456 = n9858 ^ n2987 ^ 1'b0 ;
  assign n21457 = n7444 & ~n21456 ;
  assign n21458 = ~n4684 & n6373 ;
  assign n21459 = n21458 ^ n3075 ^ 1'b0 ;
  assign n21460 = n1526 | n21459 ;
  assign n21464 = n419 & n9301 ;
  assign n21465 = n21464 ^ n2260 ^ 1'b0 ;
  assign n21466 = n2303 & n21465 ;
  assign n21461 = n2295 & ~n13743 ;
  assign n21462 = ~n16663 & n21461 ;
  assign n21463 = n1730 & ~n21462 ;
  assign n21467 = n21466 ^ n21463 ^ 1'b0 ;
  assign n21468 = n318 | n1572 ;
  assign n21469 = n13646 ^ n1608 ^ 1'b0 ;
  assign n21470 = n11158 & n21469 ;
  assign n21471 = n1471 ^ n917 ^ 1'b0 ;
  assign n21472 = n2948 & n21471 ;
  assign n21473 = ~n927 & n5461 ;
  assign n21474 = n21472 & n21473 ;
  assign n21475 = ~n3767 & n21474 ;
  assign n21476 = n21475 ^ n10507 ^ 1'b0 ;
  assign n21477 = ~n21470 & n21476 ;
  assign n21478 = ~n1308 & n18590 ;
  assign n21479 = n21478 ^ n236 ^ 1'b0 ;
  assign n21480 = n2939 | n15707 ;
  assign n21481 = n1608 | n5826 ;
  assign n21482 = ~n9206 & n21481 ;
  assign n21483 = n13795 ^ n4522 ^ 1'b0 ;
  assign n21484 = ~n6847 & n21483 ;
  assign n21485 = n6196 ^ n475 ^ 1'b0 ;
  assign n21486 = n10537 | n20086 ;
  assign n21487 = n21486 ^ n6910 ^ 1'b0 ;
  assign n21488 = n7506 ^ n4574 ^ 1'b0 ;
  assign n21489 = ~n6538 & n21488 ;
  assign n21490 = n21489 ^ n7665 ^ 1'b0 ;
  assign n21491 = ~n3202 & n21490 ;
  assign n21492 = n6453 & n17180 ;
  assign n21493 = n21492 ^ n11308 ^ 1'b0 ;
  assign n21494 = n9709 ^ n5823 ^ 1'b0 ;
  assign n21495 = n647 & ~n21494 ;
  assign n21496 = n21495 ^ n9163 ^ 1'b0 ;
  assign n21497 = ~n14146 & n21496 ;
  assign n21498 = n21493 & n21497 ;
  assign n21499 = n21498 ^ n13741 ^ 1'b0 ;
  assign n21500 = ~n14225 & n21499 ;
  assign n21501 = n6897 & n12416 ;
  assign n21502 = n21501 ^ n1704 ^ 1'b0 ;
  assign n21503 = n14200 ^ n14165 ^ 1'b0 ;
  assign n21504 = n4965 | n21503 ;
  assign n21505 = n3408 ^ n2203 ^ n2176 ;
  assign n21506 = n2235 & n20401 ;
  assign n21507 = n271 & ~n17542 ;
  assign n21508 = n9595 & ~n17495 ;
  assign n21509 = ~n2582 & n2606 ;
  assign n21510 = n11635 & n21509 ;
  assign n21511 = ~n16750 & n21510 ;
  assign n21512 = n2637 & ~n6228 ;
  assign n21513 = n1173 & ~n15041 ;
  assign n21514 = n4895 & ~n10913 ;
  assign n21515 = n21514 ^ n14715 ^ 1'b0 ;
  assign n21516 = ~n10333 & n21515 ;
  assign n21517 = n21516 ^ n14573 ^ 1'b0 ;
  assign n21518 = n15495 & ~n15559 ;
  assign n21519 = n21518 ^ n5131 ^ 1'b0 ;
  assign n21520 = n7572 ^ n1342 ^ 1'b0 ;
  assign n21521 = n3362 & ~n21520 ;
  assign n21522 = n3742 & ~n21521 ;
  assign n21523 = n1207 ^ n1025 ^ 1'b0 ;
  assign n21524 = n11471 | n21523 ;
  assign n21525 = ~n2917 & n16745 ;
  assign n21526 = n1029 | n4159 ;
  assign n21527 = ~n1355 & n13652 ;
  assign n21528 = n17721 | n19426 ;
  assign n21529 = n21528 ^ n382 ^ 1'b0 ;
  assign n21530 = n14645 ^ n2279 ^ 1'b0 ;
  assign n21531 = ~n21529 & n21530 ;
  assign n21532 = ~n4746 & n13839 ;
  assign n21533 = n9449 & n20736 ;
  assign n21534 = ~n19978 & n21533 ;
  assign n21535 = ( n4326 & n21532 ) | ( n4326 & n21534 ) | ( n21532 & n21534 ) ;
  assign n21536 = n3825 & ~n7325 ;
  assign n21537 = n21536 ^ n17104 ^ 1'b0 ;
  assign n21538 = n21535 | n21537 ;
  assign n21539 = n1874 & n4749 ;
  assign n21540 = n13928 & n21539 ;
  assign n21541 = n6466 & ~n17339 ;
  assign n21542 = ~n21540 & n21541 ;
  assign n21543 = n1143 & ~n16504 ;
  assign n21544 = n9189 & ~n10976 ;
  assign n21545 = n3180 & n21078 ;
  assign n21546 = n15759 ^ n3121 ^ 1'b0 ;
  assign n21547 = n4991 | n9971 ;
  assign n21548 = n11248 ^ n770 ^ 1'b0 ;
  assign n21549 = n21548 ^ n363 ^ 1'b0 ;
  assign n21550 = ~n15426 & n21549 ;
  assign n21551 = n21550 ^ n4613 ^ 1'b0 ;
  assign n21552 = n6269 & ~n21551 ;
  assign n21553 = n19546 ^ n6669 ^ 1'b0 ;
  assign n21554 = n21552 & n21553 ;
  assign n21555 = n6410 ^ n481 ^ 1'b0 ;
  assign n21556 = n6721 & ~n21555 ;
  assign n21557 = n5889 | n6142 ;
  assign n21558 = n15318 ^ n1087 ^ 1'b0 ;
  assign n21559 = n7442 | n21558 ;
  assign n21560 = n21559 ^ n5115 ^ 1'b0 ;
  assign n21561 = n102 | n11309 ;
  assign n21562 = ~n5782 & n8828 ;
  assign n21563 = n1458 & ~n4123 ;
  assign n21564 = n21563 ^ n232 ^ 1'b0 ;
  assign n21565 = n2071 & ~n6880 ;
  assign n21566 = n13151 & n21565 ;
  assign n21567 = n21564 & n21566 ;
  assign n21568 = n9986 & n12903 ;
  assign n21569 = ~n12257 & n12280 ;
  assign n21570 = n364 | n17187 ;
  assign n21571 = n340 & ~n21570 ;
  assign n21572 = n10443 | n21571 ;
  assign n21573 = n11202 & n21572 ;
  assign n21574 = n21573 ^ n14704 ^ 1'b0 ;
  assign n21575 = n2162 & n3443 ;
  assign n21576 = ~n2162 & n21575 ;
  assign n21577 = n1655 & ~n21576 ;
  assign n21578 = ~n1655 & n21577 ;
  assign n21579 = n2220 | n21578 ;
  assign n21580 = n3477 & n13408 ;
  assign n21581 = n17531 & n21580 ;
  assign n21582 = n21581 ^ n8053 ^ 1'b0 ;
  assign n21583 = n21579 & n21582 ;
  assign n21584 = n7192 | n13422 ;
  assign n21585 = ~n7330 & n19993 ;
  assign n21586 = n21585 ^ n4228 ^ 1'b0 ;
  assign n21587 = n21586 ^ n335 ^ 1'b0 ;
  assign n21588 = n9823 & n21587 ;
  assign n21589 = n21584 & n21588 ;
  assign n21590 = n5802 & n7867 ;
  assign n21591 = ~n11624 & n15150 ;
  assign n21592 = n9852 ^ n2432 ^ 1'b0 ;
  assign n21593 = ~n1782 & n21592 ;
  assign n21594 = n21593 ^ n15041 ^ n5722 ;
  assign n21595 = n9039 ^ n7390 ^ 1'b0 ;
  assign n21596 = n9847 | n21595 ;
  assign n21597 = n998 & ~n6577 ;
  assign n21598 = ~n2403 & n21597 ;
  assign n21599 = n21598 ^ n7056 ^ 1'b0 ;
  assign n21600 = n21599 ^ n14181 ^ 1'b0 ;
  assign n21601 = n1194 & ~n21600 ;
  assign n21602 = ~n15801 & n21601 ;
  assign n21603 = n21596 & n21602 ;
  assign n21604 = n13376 ^ n52 ^ 1'b0 ;
  assign n21605 = n6537 & n21604 ;
  assign n21606 = n12453 ^ n4942 ^ 1'b0 ;
  assign n21607 = n7266 | n21606 ;
  assign n21608 = n2088 & n2885 ;
  assign n21609 = ( ~n3451 & n21372 ) | ( ~n3451 & n21608 ) | ( n21372 & n21608 ) ;
  assign n21610 = n11266 & n17390 ;
  assign n21611 = n395 & ~n2904 ;
  assign n21612 = n13408 ^ n653 ^ 1'b0 ;
  assign n21613 = n13572 ^ n4872 ^ 1'b0 ;
  assign n21614 = n5205 | n5698 ;
  assign n21615 = n21614 ^ n8158 ^ 1'b0 ;
  assign n21616 = n4559 ^ n1233 ^ 1'b0 ;
  assign n21617 = n21616 ^ n553 ^ 1'b0 ;
  assign n21618 = n13635 & ~n21617 ;
  assign n21619 = n21615 & ~n21618 ;
  assign n21620 = n1248 & n10489 ;
  assign n21621 = ~n4976 & n21620 ;
  assign n21622 = n6864 & ~n21621 ;
  assign n21623 = n817 & ~n12089 ;
  assign n21624 = n21623 ^ n2594 ^ 1'b0 ;
  assign n21625 = ~n3459 & n21624 ;
  assign n21626 = n5183 ^ n2282 ^ 1'b0 ;
  assign n21627 = n3575 & ~n21626 ;
  assign n21628 = n21627 ^ n18186 ^ 1'b0 ;
  assign n21629 = n19559 ^ n1304 ^ 1'b0 ;
  assign n21630 = n6850 & n16216 ;
  assign n21631 = n21630 ^ n10707 ^ 1'b0 ;
  assign n21632 = n1887 & n2774 ;
  assign n21633 = n4332 | n18091 ;
  assign n21634 = n21633 ^ n3211 ^ 1'b0 ;
  assign n21635 = n14044 & ~n21634 ;
  assign n21636 = n10765 ^ n8046 ^ n2665 ;
  assign n21637 = n9315 & ~n9794 ;
  assign n21638 = n1219 & n21637 ;
  assign n21639 = ~n6087 & n7322 ;
  assign n21640 = n16808 & n21639 ;
  assign n21641 = n1604 & ~n14454 ;
  assign n21642 = ~n5076 & n16431 ;
  assign n21643 = ( ~n1368 & n1441 ) | ( ~n1368 & n5899 ) | ( n1441 & n5899 ) ;
  assign n21644 = n21643 ^ n5115 ^ 1'b0 ;
  assign n21645 = ~n2004 & n17572 ;
  assign n21646 = n8202 & n21645 ;
  assign n21647 = n21646 ^ n8795 ^ 1'b0 ;
  assign n21648 = n2996 | n10273 ;
  assign n21649 = n21648 ^ n18932 ^ 1'b0 ;
  assign n21650 = n9554 ^ n3901 ^ 1'b0 ;
  assign n21651 = n1388 ^ n798 ^ 1'b0 ;
  assign n21652 = n19801 & ~n21651 ;
  assign n21653 = ~n13023 & n21652 ;
  assign n21654 = ~n4191 & n9833 ;
  assign n21655 = n13903 ^ n9366 ^ 1'b0 ;
  assign n21656 = n2752 | n19293 ;
  assign n21657 = n5135 ^ n5076 ^ 1'b0 ;
  assign n21658 = n6730 & n14422 ;
  assign n21659 = n1945 & ~n10582 ;
  assign n21660 = n21659 ^ n3413 ^ 1'b0 ;
  assign n21661 = n1007 & n13320 ;
  assign n21662 = n12223 & n21661 ;
  assign n21663 = n272 | n9390 ;
  assign n21664 = n175 | n21663 ;
  assign n21665 = n21663 & ~n21664 ;
  assign n21666 = n21665 ^ n11526 ^ 1'b0 ;
  assign n21667 = n21662 & n21666 ;
  assign n21668 = n9062 ^ n2209 ^ 1'b0 ;
  assign n21669 = n19830 & n21668 ;
  assign n21671 = n6370 & n12236 ;
  assign n21670 = ~n12016 & n15711 ;
  assign n21672 = n21671 ^ n21670 ^ 1'b0 ;
  assign n21673 = n14549 & ~n21455 ;
  assign n21674 = ~n223 & n21673 ;
  assign n21675 = n13861 | n19721 ;
  assign n21676 = ~n19796 & n21675 ;
  assign n21677 = n21676 ^ n2951 ^ 1'b0 ;
  assign n21678 = n243 & ~n8510 ;
  assign n21679 = ~n236 & n2757 ;
  assign n21680 = n21678 & n21679 ;
  assign n21681 = ~n8935 & n10282 ;
  assign n21682 = ~n58 & n12881 ;
  assign n21683 = n21682 ^ n83 ^ 1'b0 ;
  assign n21684 = n538 | n3221 ;
  assign n21685 = n10355 ^ n10246 ^ 1'b0 ;
  assign n21686 = n9287 & ~n10443 ;
  assign n21711 = ~n627 & n4220 ;
  assign n21712 = n20819 ^ n13135 ^ 1'b0 ;
  assign n21713 = n21711 | n21712 ;
  assign n21703 = n151 | n236 ;
  assign n21704 = n236 & ~n21703 ;
  assign n21705 = n46 & n21704 ;
  assign n21706 = ~n991 & n21705 ;
  assign n21707 = n21706 ^ n1992 ^ 1'b0 ;
  assign n21687 = n183 & ~n357 ;
  assign n21688 = n357 & n21687 ;
  assign n21689 = x4 & ~n21688 ;
  assign n21690 = ~x4 & n21689 ;
  assign n21691 = n15729 & ~n21690 ;
  assign n21692 = n376 | n1115 ;
  assign n21693 = n21691 & ~n21692 ;
  assign n21694 = n21693 ^ n11355 ^ 1'b0 ;
  assign n21695 = n1465 | n4563 ;
  assign n21696 = n4563 & ~n21695 ;
  assign n21697 = n900 | n8245 ;
  assign n21698 = n8245 & ~n21697 ;
  assign n21699 = n21696 | n21698 ;
  assign n21700 = n21696 & ~n21699 ;
  assign n21701 = n21700 ^ n9835 ^ 1'b0 ;
  assign n21702 = n21694 & ~n21701 ;
  assign n21708 = n21707 ^ n21702 ^ 1'b0 ;
  assign n21709 = n4077 & n21708 ;
  assign n21710 = n2774 | n21709 ;
  assign n21714 = n21713 ^ n21710 ^ 1'b0 ;
  assign n21715 = n7943 ^ n3464 ^ 1'b0 ;
  assign n21716 = n16592 & ~n21715 ;
  assign n21717 = n21716 ^ n6552 ^ 1'b0 ;
  assign n21718 = n21717 ^ n15631 ^ 1'b0 ;
  assign n21719 = n16930 ^ n6529 ^ 1'b0 ;
  assign n21720 = n5158 & ~n17789 ;
  assign n21721 = ~n1460 & n4972 ;
  assign n21722 = n10442 ^ n1961 ^ 1'b0 ;
  assign n21723 = n2378 | n21722 ;
  assign n21724 = n21723 ^ n7442 ^ 1'b0 ;
  assign n21725 = n14541 ^ n6631 ^ 1'b0 ;
  assign n21726 = n12887 ^ n1472 ^ 1'b0 ;
  assign n21727 = n21725 & n21726 ;
  assign n21728 = n20010 ^ x3 ^ 1'b0 ;
  assign n21729 = n6115 ^ n2723 ^ 1'b0 ;
  assign n21730 = n1470 & n15144 ;
  assign n21731 = n4171 ^ n292 ^ 1'b0 ;
  assign n21732 = n5785 & ~n8946 ;
  assign n21733 = n21732 ^ n7179 ^ 1'b0 ;
  assign n21734 = n18579 & ~n18842 ;
  assign n21735 = n7901 & ~n16827 ;
  assign n21736 = n8230 | n10441 ;
  assign n21737 = ~n20694 & n21736 ;
  assign n21738 = n508 & n1498 ;
  assign n21739 = n10018 & n12366 ;
  assign n21740 = n21738 & n21739 ;
  assign n21741 = n21212 & n21740 ;
  assign n21742 = n9033 & n21741 ;
  assign n21743 = n7435 | n7924 ;
  assign n21744 = n3732 | n4694 ;
  assign n21745 = n20763 ^ n20270 ^ 1'b0 ;
  assign n21746 = ~n21744 & n21745 ;
  assign n21747 = n4337 ^ n654 ^ 1'b0 ;
  assign n21748 = n10661 & ~n21747 ;
  assign n21749 = n16124 | n21748 ;
  assign n21750 = n21749 ^ n13579 ^ 1'b0 ;
  assign n21751 = n1304 & ~n21750 ;
  assign n21752 = n6439 ^ n3484 ^ 1'b0 ;
  assign n21753 = n21752 ^ n15866 ^ 1'b0 ;
  assign n21754 = n7973 & ~n8031 ;
  assign n21755 = n1263 | n6753 ;
  assign n21756 = n21755 ^ n322 ^ 1'b0 ;
  assign n21757 = n10364 ^ n4963 ^ 1'b0 ;
  assign n21758 = n364 & n2046 ;
  assign n21759 = n21758 ^ n3074 ^ 1'b0 ;
  assign n21760 = n20723 & ~n21759 ;
  assign n21761 = n21760 ^ n7185 ^ 1'b0 ;
  assign n21762 = n18326 & n21761 ;
  assign n21763 = n359 & ~n11629 ;
  assign n21764 = n21763 ^ n5885 ^ 1'b0 ;
  assign n21765 = n21764 ^ n8109 ^ 1'b0 ;
  assign n21766 = n6209 ^ n5788 ^ 1'b0 ;
  assign n21767 = n21766 ^ n17100 ^ n11364 ;
  assign n21768 = n1655 & ~n21767 ;
  assign n21769 = ~n6866 & n21768 ;
  assign n21770 = ~n546 & n2644 ;
  assign n21771 = n21770 ^ n3061 ^ 1'b0 ;
  assign n21772 = n2341 & n13947 ;
  assign n21773 = n21771 | n21772 ;
  assign n21774 = n1714 & n10078 ;
  assign n21775 = n21774 ^ n1310 ^ 1'b0 ;
  assign n21776 = n21775 ^ n1118 ^ 1'b0 ;
  assign n21777 = n11178 & ~n21776 ;
  assign n21778 = n21773 | n21777 ;
  assign n21779 = n4832 | n10998 ;
  assign n21780 = n21779 ^ n14948 ^ 1'b0 ;
  assign n21781 = ~n6571 & n21780 ;
  assign n21782 = n7610 & ~n9422 ;
  assign n21783 = n21209 & n21782 ;
  assign n21784 = n3306 ^ n1748 ^ 1'b0 ;
  assign n21785 = n20650 & ~n21784 ;
  assign n21786 = n13797 ^ n13246 ^ 1'b0 ;
  assign n21787 = ~n8226 & n21786 ;
  assign n21788 = ~n1273 & n6667 ;
  assign n21789 = n21788 ^ n535 ^ 1'b0 ;
  assign n21790 = n6552 & ~n21789 ;
  assign n21791 = n5501 & ~n21790 ;
  assign n21792 = n934 & n5083 ;
  assign n21793 = n21792 ^ n11338 ^ 1'b0 ;
  assign n21794 = ~n5128 & n7377 ;
  assign n21795 = n7045 ^ n4864 ^ 1'b0 ;
  assign n21796 = ~n2855 & n21795 ;
  assign n21797 = n14385 | n21796 ;
  assign n21798 = n21794 & ~n21797 ;
  assign n21799 = n9758 & ~n12661 ;
  assign n21800 = ~n627 & n8220 ;
  assign n21801 = n15687 ^ n9152 ^ 1'b0 ;
  assign n21802 = ~n11578 & n21801 ;
  assign n21803 = n21802 ^ n12690 ^ 1'b0 ;
  assign n21804 = n6244 | n21803 ;
  assign n21805 = ( ~n3718 & n5164 ) | ( ~n3718 & n11158 ) | ( n5164 & n11158 ) ;
  assign n21806 = n4468 | n11106 ;
  assign n21807 = n18329 ^ n8990 ^ 1'b0 ;
  assign n21808 = n1452 & ~n10446 ;
  assign n21809 = n11672 ^ n1702 ^ 1'b0 ;
  assign n21810 = n10449 & ~n15244 ;
  assign n21811 = ( n512 & ~n8782 ) | ( n512 & n21810 ) | ( ~n8782 & n21810 ) ;
  assign n21812 = n21811 ^ n1283 ^ 1'b0 ;
  assign n21817 = ~n963 & n1057 ;
  assign n21818 = n393 & n21817 ;
  assign n21819 = n13956 ^ n1549 ^ 1'b0 ;
  assign n21820 = ~n21818 & n21819 ;
  assign n21821 = ~n4332 & n21820 ;
  assign n21822 = n3037 & n21821 ;
  assign n21815 = ~n3539 & n7670 ;
  assign n21813 = n2310 & ~n2740 ;
  assign n21814 = n539 & n21813 ;
  assign n21816 = n21815 ^ n21814 ^ n14043 ;
  assign n21823 = n21822 ^ n21816 ^ 1'b0 ;
  assign n21824 = n6585 & ~n14544 ;
  assign n21825 = n3588 ^ n857 ^ 1'b0 ;
  assign n21826 = n1802 & ~n21825 ;
  assign n21827 = n21824 & n21826 ;
  assign n21828 = n7780 & ~n21827 ;
  assign n21829 = n21828 ^ n13073 ^ 1'b0 ;
  assign n21830 = n191 | n10992 ;
  assign n21831 = n21830 ^ n1388 ^ 1'b0 ;
  assign n21832 = ~n6398 & n10459 ;
  assign n21833 = ~n5204 & n21832 ;
  assign n21834 = ~n133 & n20788 ;
  assign n21835 = n14235 ^ n2157 ^ 1'b0 ;
  assign n21836 = n133 | n21835 ;
  assign n21837 = n10100 & ~n21836 ;
  assign n21838 = n68 | n19014 ;
  assign n21839 = n21838 ^ n11520 ^ 1'b0 ;
  assign n21840 = n21839 ^ n9569 ^ 1'b0 ;
  assign n21841 = n3292 & n21840 ;
  assign n21842 = n2252 & ~n7185 ;
  assign n21843 = ~n13278 & n21842 ;
  assign n21844 = n13382 & ~n21843 ;
  assign n21846 = ~n5778 & n9577 ;
  assign n21847 = ~n5282 & n21846 ;
  assign n21848 = n9194 & ~n21847 ;
  assign n21845 = ~n1497 & n4019 ;
  assign n21849 = n21848 ^ n21845 ^ 1'b0 ;
  assign n21850 = ~n5196 & n21849 ;
  assign n21851 = n16679 ^ n10444 ^ 1'b0 ;
  assign n21852 = n2604 & ~n21851 ;
  assign n21856 = n6481 & ~n11803 ;
  assign n21853 = n823 ^ n384 ^ 1'b0 ;
  assign n21854 = n18201 & ~n21853 ;
  assign n21855 = n7582 & n21854 ;
  assign n21857 = n21856 ^ n21855 ^ 1'b0 ;
  assign n21858 = n21852 | n21857 ;
  assign n21859 = n10787 ^ n9284 ^ 1'b0 ;
  assign n21862 = n6376 & ~n17229 ;
  assign n21863 = n5068 | n21862 ;
  assign n21860 = ~n690 & n5412 ;
  assign n21861 = n1414 & n21860 ;
  assign n21864 = n21863 ^ n21861 ^ 1'b0 ;
  assign n21865 = n1086 | n18694 ;
  assign n21866 = n9851 & ~n21865 ;
  assign n21867 = n11357 | n14556 ;
  assign n21868 = n5293 & ~n21867 ;
  assign n21869 = ~n8825 & n9140 ;
  assign n21870 = n10009 & n21869 ;
  assign n21871 = n800 & ~n19600 ;
  assign n21872 = n21871 ^ n7079 ^ 1'b0 ;
  assign n21873 = n21326 ^ n7350 ^ 1'b0 ;
  assign n21874 = n5169 & ~n21873 ;
  assign n21875 = n14647 ^ n9979 ^ 1'b0 ;
  assign n21876 = n20111 & n21875 ;
  assign n21877 = n2577 & ~n2733 ;
  assign n21878 = n12688 ^ n2394 ^ 1'b0 ;
  assign n21879 = n16170 & n21878 ;
  assign n21880 = n14067 | n21879 ;
  assign n21881 = n361 & n2001 ;
  assign n21882 = ~n14236 & n21881 ;
  assign n21884 = n567 & ~n3452 ;
  assign n21883 = n10392 ^ n5953 ^ 1'b0 ;
  assign n21885 = n21884 ^ n21883 ^ 1'b0 ;
  assign n21886 = ~n11690 & n21885 ;
  assign n21887 = n2955 & n4197 ;
  assign n21888 = ~n3395 & n21887 ;
  assign n21889 = n751 & ~n17295 ;
  assign n21890 = n21889 ^ n11934 ^ 1'b0 ;
  assign n21891 = n532 | n11549 ;
  assign n21892 = n21891 ^ n18909 ^ 1'b0 ;
  assign n21893 = n323 | n12133 ;
  assign n21894 = n12133 | n21893 ;
  assign n21895 = n12133 & ~n21894 ;
  assign n21896 = n43 & n12139 ;
  assign n21897 = n109 & n12580 ;
  assign n21898 = n21896 | n21897 ;
  assign n21899 = n21896 & ~n21898 ;
  assign n21900 = n21899 ^ n100 ^ 1'b0 ;
  assign n21901 = n21895 | n21900 ;
  assign n21902 = n21895 & ~n21901 ;
  assign n21903 = x6 & n56 ;
  assign n21904 = n12135 & n21903 ;
  assign n21905 = n69 | n21904 ;
  assign n21906 = n101 ^ n36 ^ 1'b0 ;
  assign n21907 = n36 & n21906 ;
  assign n21908 = n34 & ~n100 ;
  assign n21909 = ~n34 & n21908 ;
  assign n21910 = n20876 | n21909 ;
  assign n21911 = n20876 & ~n21910 ;
  assign n21912 = n12580 | n21911 ;
  assign n21913 = n12580 & ~n21912 ;
  assign n21914 = n21907 | n21913 ;
  assign n21915 = n21905 | n21914 ;
  assign n21916 = n21902 & ~n21915 ;
  assign n21917 = n198 | n467 ;
  assign n21918 = n21916 & ~n21917 ;
  assign n21919 = n6196 | n10407 ;
  assign n21920 = n10407 & ~n21919 ;
  assign n21921 = ~n870 & n4203 ;
  assign n21922 = ~n4203 & n21921 ;
  assign n21923 = n2874 & n21922 ;
  assign n21924 = ~n21920 & n21923 ;
  assign n21925 = n1841 & n15346 ;
  assign n21926 = ~n177 & n21925 ;
  assign n21927 = n4737 & n21926 ;
  assign n21928 = n2235 & n21927 ;
  assign n21929 = ~n3773 & n21928 ;
  assign n21930 = n3221 & n21929 ;
  assign n21931 = n21924 & ~n21930 ;
  assign n21932 = ~n21924 & n21931 ;
  assign n21933 = n21918 | n21932 ;
  assign n21934 = n21918 & ~n21933 ;
  assign n21935 = n21263 | n21934 ;
  assign n21936 = n14551 & ~n21935 ;
  assign n21937 = n6843 & ~n16170 ;
  assign n21938 = n6523 | n21937 ;
  assign n21939 = n1550 & n6282 ;
  assign n21940 = n21939 ^ n3047 ^ 1'b0 ;
  assign n21941 = n18869 & n21940 ;
  assign n21942 = n142 & ~n2577 ;
  assign n21943 = n1838 & ~n2575 ;
  assign n21944 = n8994 & ~n21943 ;
  assign n21945 = n6999 & ~n8892 ;
  assign n21946 = n10463 ^ n1388 ^ 1'b0 ;
  assign n21947 = n6995 & n21946 ;
  assign n21948 = n14066 ^ n9177 ^ 1'b0 ;
  assign n21949 = ~n17741 & n18286 ;
  assign n21950 = n21948 & n21949 ;
  assign n21951 = n9398 & n12446 ;
  assign n21952 = n21299 & n21951 ;
  assign n21953 = ~n12411 & n13096 ;
  assign n21954 = n11664 & ~n21953 ;
  assign n21955 = n21954 ^ n2001 ^ 1'b0 ;
  assign n21956 = n3786 | n16098 ;
  assign n21957 = n17969 ^ n3466 ^ 1'b0 ;
  assign n21958 = n14158 & n21957 ;
  assign n21959 = n3818 & ~n8571 ;
  assign n21960 = n9340 & n21959 ;
  assign n21962 = n4399 ^ n4327 ^ 1'b0 ;
  assign n21961 = n2497 & n9758 ;
  assign n21963 = n21962 ^ n21961 ^ n15879 ;
  assign n21964 = ~n4281 & n8416 ;
  assign n21965 = n21964 ^ n1388 ^ 1'b0 ;
  assign n21966 = n4824 & ~n16332 ;
  assign n21967 = n1130 & n13694 ;
  assign n21968 = ~n8900 & n21967 ;
  assign n21969 = n21968 ^ n20903 ^ 1'b0 ;
  assign n21970 = n2816 ^ n1873 ^ 1'b0 ;
  assign n21971 = ~n2843 & n21970 ;
  assign n21972 = ~n1440 & n21971 ;
  assign n21973 = n21972 ^ n3036 ^ 1'b0 ;
  assign n21974 = ~n13188 & n16217 ;
  assign n21975 = n12953 & n21974 ;
  assign n21976 = n13608 ^ n2513 ^ 1'b0 ;
  assign n21977 = ~n6207 & n6222 ;
  assign n21978 = n18133 & ~n21977 ;
  assign n21979 = n5391 & n20698 ;
  assign n21980 = n6525 & n7090 ;
  assign n21981 = n21980 ^ n2668 ^ 1'b0 ;
  assign n21982 = n2991 & ~n21970 ;
  assign n21983 = n1660 & ~n21982 ;
  assign n21984 = ~n402 & n21983 ;
  assign n21985 = n12639 ^ n5286 ^ 1'b0 ;
  assign n21986 = n43 | n21985 ;
  assign n21987 = n3750 & n5694 ;
  assign n21988 = n19611 | n20059 ;
  assign n21989 = n4426 ^ n1765 ^ 1'b0 ;
  assign n21990 = n21989 ^ n4969 ^ 1'b0 ;
  assign n21991 = n9606 & ~n15201 ;
  assign n21992 = ~x3 & n21991 ;
  assign n21993 = n254 | n2414 ;
  assign n21994 = n21993 ^ n13792 ^ n10291 ;
  assign n21995 = n2911 | n21994 ;
  assign n21996 = n21995 ^ n16479 ^ 1'b0 ;
  assign n21997 = ~n2277 & n12777 ;
  assign n21999 = n12495 | n17253 ;
  assign n21998 = ~n3433 & n4855 ;
  assign n22000 = n21999 ^ n21998 ^ 1'b0 ;
  assign n22001 = n154 & ~n163 ;
  assign n22002 = n163 & n22001 ;
  assign n22003 = n182 & n22002 ;
  assign n22004 = n1407 | n22003 ;
  assign n22005 = n22003 & ~n22004 ;
  assign n22006 = n16 & n121 ;
  assign n22007 = ~n121 & n22006 ;
  assign n22008 = n22007 ^ n7829 ^ 1'b0 ;
  assign n22009 = n22005 | n22008 ;
  assign n22010 = n22005 & ~n22009 ;
  assign n22011 = n1011 | n1039 ;
  assign n22012 = n22010 & ~n22011 ;
  assign n22013 = n255 | n20157 ;
  assign n22014 = n255 & ~n22013 ;
  assign n22015 = n88 & ~n22014 ;
  assign n22016 = ~n88 & n22015 ;
  assign n22017 = n4535 & ~n13682 ;
  assign n22018 = n13682 & n22017 ;
  assign n22019 = n22016 & ~n22018 ;
  assign n22020 = n1820 & n22019 ;
  assign n22021 = n22012 & n22020 ;
  assign n22022 = n6421 & ~n22021 ;
  assign n22023 = n16001 & n22022 ;
  assign n22024 = ~n2709 & n3526 ;
  assign n22025 = ~n3526 & n22024 ;
  assign n22026 = ~n410 & n22025 ;
  assign n22027 = n22023 | n22026 ;
  assign n22028 = n22023 & ~n22027 ;
  assign n22029 = ~n371 & n7005 ;
  assign n22030 = n12371 ^ n5264 ^ 1'b0 ;
  assign n22031 = n5625 & n22030 ;
  assign n22032 = n12453 ^ n461 ^ 1'b0 ;
  assign n22033 = n6959 & n22032 ;
  assign n22034 = n339 | n17189 ;
  assign n22035 = n8857 | n19789 ;
  assign n22036 = n6915 & ~n22035 ;
  assign n22037 = n3894 | n22036 ;
  assign n22038 = ~n5735 & n10991 ;
  assign n22039 = n1053 | n5943 ;
  assign n22040 = n12407 ^ n5254 ^ 1'b0 ;
  assign n22041 = n22039 & ~n22040 ;
  assign n22042 = n9959 ^ n1693 ^ 1'b0 ;
  assign n22043 = ~n9691 & n18622 ;
  assign n22044 = ~n1368 & n22043 ;
  assign n22045 = n278 & ~n782 ;
  assign n22046 = n1235 ^ n105 ^ 1'b0 ;
  assign n22047 = n3663 & n16050 ;
  assign n22048 = n4674 | n21475 ;
  assign n22049 = n3007 | n7051 ;
  assign n22050 = n9495 & n21586 ;
  assign n22051 = n102 & ~n21299 ;
  assign n22052 = n22051 ^ n10208 ^ 1'b0 ;
  assign n22053 = n6281 ^ n4550 ^ 1'b0 ;
  assign n22054 = n9472 & ~n11957 ;
  assign n22055 = n22054 ^ n6405 ^ 1'b0 ;
  assign n22056 = n22055 ^ n7792 ^ 1'b0 ;
  assign n22057 = ~n7713 & n22056 ;
  assign n22058 = n20101 & n22057 ;
  assign n22059 = n16362 & n22058 ;
  assign n22060 = n22059 ^ n11946 ^ 1'b0 ;
  assign n22061 = ~n3133 & n22060 ;
  assign n22062 = n13708 ^ n545 ^ 1'b0 ;
  assign n22063 = ~n8497 & n22062 ;
  assign n22064 = n15040 ^ n1243 ^ 1'b0 ;
  assign n22065 = n440 & ~n22064 ;
  assign n22066 = n2410 | n12272 ;
  assign n22067 = n14235 ^ n7909 ^ 1'b0 ;
  assign n22068 = n957 & n22067 ;
  assign n22071 = n2371 & ~n2828 ;
  assign n22072 = n22071 ^ n1995 ^ 1'b0 ;
  assign n22069 = n4295 ^ n3476 ^ 1'b0 ;
  assign n22070 = n107 | n22069 ;
  assign n22073 = n22072 ^ n22070 ^ 1'b0 ;
  assign n22074 = n15100 | n22073 ;
  assign n22075 = n10122 ^ n4222 ^ 1'b0 ;
  assign n22076 = ~n14784 & n22075 ;
  assign n22077 = n3402 & n22076 ;
  assign n22078 = n22077 ^ n9881 ^ 1'b0 ;
  assign n22079 = n3431 | n9588 ;
  assign n22080 = n3422 | n21808 ;
  assign n22081 = n354 & n17967 ;
  assign n22083 = n14885 ^ n8415 ^ 1'b0 ;
  assign n22082 = ~n7741 & n12968 ;
  assign n22084 = n22083 ^ n22082 ^ 1'b0 ;
  assign n22085 = n5348 ^ n3539 ^ 1'b0 ;
  assign n22086 = n22085 ^ n13735 ^ n3509 ;
  assign n22087 = n375 ^ n227 ^ 1'b0 ;
  assign n22088 = n3220 | n22087 ;
  assign n22089 = n22088 ^ n15015 ^ n7722 ;
  assign n22090 = n22089 ^ n10947 ^ 1'b0 ;
  assign n22091 = n13011 | n22090 ;
  assign n22092 = n13094 | n22091 ;
  assign n22093 = n7401 ^ n1467 ^ 1'b0 ;
  assign n22094 = n11803 & n22093 ;
  assign n22097 = ~n5338 & n9563 ;
  assign n22095 = n338 & n3472 ;
  assign n22096 = n14515 & n22095 ;
  assign n22098 = n22097 ^ n22096 ^ 1'b0 ;
  assign n22099 = ~n3797 & n12804 ;
  assign n22100 = n2751 & n22099 ;
  assign n22101 = ( n3861 & n11689 ) | ( n3861 & n22100 ) | ( n11689 & n22100 ) ;
  assign n22102 = ( ~n3452 & n4895 ) | ( ~n3452 & n9408 ) | ( n4895 & n9408 ) ;
  assign n22103 = n18289 | n22102 ;
  assign n22104 = n19083 ^ n17955 ^ 1'b0 ;
  assign n22105 = n19020 ^ n12541 ^ 1'b0 ;
  assign n22106 = ~n7430 & n22105 ;
  assign n22109 = n1526 | n3928 ;
  assign n22110 = n7615 & ~n22109 ;
  assign n22107 = n1588 & n3844 ;
  assign n22108 = n18125 & n22107 ;
  assign n22111 = n22110 ^ n22108 ^ 1'b0 ;
  assign n22112 = ~n4271 & n16742 ;
  assign n22113 = n11827 | n12470 ;
  assign n22114 = n11904 | n22113 ;
  assign n22115 = n141 & ~n17903 ;
  assign n22116 = n9018 & ~n19758 ;
  assign n22117 = n9409 & n22116 ;
  assign n22118 = n7301 ^ n6449 ^ 1'b0 ;
  assign n22119 = n178 | n767 ;
  assign n22120 = ~n8210 & n22119 ;
  assign n22121 = ~n6278 & n22120 ;
  assign n22122 = n18217 & n22121 ;
  assign n22123 = n405 | n20432 ;
  assign n22124 = n22123 ^ n15441 ^ 1'b0 ;
  assign n22125 = n13909 ^ n8622 ^ 1'b0 ;
  assign n22126 = n14186 | n22125 ;
  assign n22127 = n2007 & n16545 ;
  assign n22128 = n11940 & n22127 ;
  assign n22129 = ~n16190 & n22128 ;
  assign n22130 = n3965 ^ n2017 ^ 1'b0 ;
  assign n22131 = n14991 ^ n1345 ^ 1'b0 ;
  assign n22132 = n4214 ^ n924 ^ 1'b0 ;
  assign n22133 = n15448 | n22132 ;
  assign n22134 = n1016 & n18216 ;
  assign n22135 = n17899 & n22134 ;
  assign n22136 = ~n4025 & n7148 ;
  assign n22137 = n22136 ^ n979 ^ 1'b0 ;
  assign n22138 = n22137 ^ n8886 ^ 1'b0 ;
  assign n22139 = ~n22135 & n22138 ;
  assign n22140 = n20077 & n22139 ;
  assign n22141 = n7491 ^ n340 ^ 1'b0 ;
  assign n22142 = n2159 & ~n8769 ;
  assign n22143 = ~n338 & n22142 ;
  assign n22144 = n4306 & ~n5463 ;
  assign n22145 = n12280 & n19713 ;
  assign n22146 = n3774 & ~n4899 ;
  assign n22147 = n22146 ^ n20623 ^ 1'b0 ;
  assign n22148 = x3 & ~n10441 ;
  assign n22149 = n296 & n22148 ;
  assign n22150 = n22149 ^ n18610 ^ 1'b0 ;
  assign n22151 = n621 | n1866 ;
  assign n22152 = n22151 ^ n2334 ^ 1'b0 ;
  assign n22153 = n4400 | n4787 ;
  assign n22154 = n4455 & ~n22153 ;
  assign n22155 = n22152 & ~n22154 ;
  assign n22156 = n22155 ^ n17738 ^ 1'b0 ;
  assign n22157 = n2842 | n5053 ;
  assign n22158 = n17176 | n22157 ;
  assign n22159 = n22158 ^ n12509 ^ 1'b0 ;
  assign n22160 = n17349 ^ n6865 ^ 1'b0 ;
  assign n22161 = n12982 ^ n5749 ^ 1'b0 ;
  assign n22162 = n16853 ^ n13329 ^ 1'b0 ;
  assign n22163 = n22161 | n22162 ;
  assign n22164 = n5626 & ~n14430 ;
  assign n22165 = n622 & n6868 ;
  assign n22166 = ~n4618 & n22165 ;
  assign n22167 = n9925 | n12702 ;
  assign n22168 = n8333 | n22167 ;
  assign n22169 = n1552 & n22168 ;
  assign n22170 = ~n11946 & n19629 ;
  assign n22171 = n4169 & ~n6370 ;
  assign n22172 = n22171 ^ n2825 ^ 1'b0 ;
  assign n22173 = n17016 & ~n22172 ;
  assign n22174 = n791 & ~n995 ;
  assign n22175 = n22174 ^ n1149 ^ 1'b0 ;
  assign n22176 = n22175 ^ n6043 ^ 1'b0 ;
  assign n22177 = n6278 | n22176 ;
  assign n22178 = n6137 ^ n1771 ^ 1'b0 ;
  assign n22179 = n4437 | n22178 ;
  assign n22180 = ~n6412 & n14172 ;
  assign n22181 = n13449 | n22180 ;
  assign n22182 = n14378 ^ n4921 ^ 1'b0 ;
  assign n22183 = n13693 ^ n817 ^ 1'b0 ;
  assign n22185 = ~n2412 & n3144 ;
  assign n22184 = n6644 ^ n4838 ^ 1'b0 ;
  assign n22186 = n22185 ^ n22184 ^ 1'b0 ;
  assign n22187 = n17621 & n22186 ;
  assign n22188 = n14450 ^ n3940 ^ 1'b0 ;
  assign n22189 = n22188 ^ n15834 ^ 1'b0 ;
  assign n22190 = n14080 | n22189 ;
  assign n22191 = n5927 | n22190 ;
  assign n22192 = n14727 ^ n6424 ^ 1'b0 ;
  assign n22193 = n12429 ^ n10442 ^ 1'b0 ;
  assign n22194 = n5583 ^ n1478 ^ 1'b0 ;
  assign n22195 = n16097 & n22194 ;
  assign n22196 = n4155 & ~n8389 ;
  assign n22197 = ( ~n1495 & n14235 ) | ( ~n1495 & n22196 ) | ( n14235 & n22196 ) ;
  assign n22198 = ( n8825 & ~n22195 ) | ( n8825 & n22197 ) | ( ~n22195 & n22197 ) ;
  assign n22200 = n12407 ^ n12315 ^ 1'b0 ;
  assign n22199 = n6303 & n12888 ;
  assign n22201 = n22200 ^ n22199 ^ 1'b0 ;
  assign n22202 = n22201 ^ n1879 ^ 1'b0 ;
  assign n22203 = ~n21607 & n22202 ;
  assign n22204 = n2440 | n6960 ;
  assign n22205 = n22204 ^ n7456 ^ 1'b0 ;
  assign n22206 = ~n5011 & n21610 ;
  assign n22207 = n1997 & n16738 ;
  assign n22208 = n20104 ^ n5284 ^ 1'b0 ;
  assign n22209 = n1165 & n3947 ;
  assign n22210 = n16687 ^ n1770 ^ 1'b0 ;
  assign n22211 = ~n2222 & n8489 ;
  assign n22212 = n4708 & ~n6586 ;
  assign n22213 = n5239 & n22212 ;
  assign n22214 = n3407 & n22213 ;
  assign n22215 = n22214 ^ n19783 ^ 1'b0 ;
  assign n22216 = n22215 ^ n3574 ^ 1'b0 ;
  assign n22217 = n13759 ^ n4161 ^ 1'b0 ;
  assign n22218 = n664 | n19476 ;
  assign n22219 = ( ~n3635 & n8842 ) | ( ~n3635 & n10439 ) | ( n8842 & n10439 ) ;
  assign n22220 = n18636 ^ n2108 ^ 1'b0 ;
  assign n22221 = ~n8387 & n22220 ;
  assign n22222 = n4525 & n6689 ;
  assign n22223 = n22222 ^ n9541 ^ 1'b0 ;
  assign n22224 = ~n2998 & n16572 ;
  assign n22225 = n7927 & n22224 ;
  assign n22226 = n22225 ^ n11178 ^ 1'b0 ;
  assign n22227 = ( ~n773 & n22223 ) | ( ~n773 & n22226 ) | ( n22223 & n22226 ) ;
  assign n22228 = n5219 ^ n615 ^ 1'b0 ;
  assign n22229 = n1676 & n22228 ;
  assign n22230 = ~n1914 & n1968 ;
  assign n22231 = n1490 & ~n2469 ;
  assign n22232 = n13839 & n22231 ;
  assign n22233 = n22230 & n22232 ;
  assign n22234 = n22233 ^ n3263 ^ 1'b0 ;
  assign n22235 = ~n4835 & n22234 ;
  assign n22236 = n22235 ^ n9992 ^ 1'b0 ;
  assign n22237 = ~n3855 & n6074 ;
  assign n22239 = ~n4766 & n6078 ;
  assign n22238 = ~n2904 & n3100 ;
  assign n22240 = n22239 ^ n22238 ^ 1'b0 ;
  assign n22241 = n4550 | n15163 ;
  assign n22242 = ~n1165 & n22241 ;
  assign n22243 = n2562 | n18973 ;
  assign n22244 = n22243 ^ n5319 ^ 1'b0 ;
  assign n22245 = ~n910 & n22244 ;
  assign n22246 = n616 | n22245 ;
  assign n22247 = n4697 | n17851 ;
  assign n22248 = n5691 & n22247 ;
  assign n22249 = n22248 ^ n8966 ^ 1'b0 ;
  assign n22250 = n1463 & n4722 ;
  assign n22251 = n16474 & n22250 ;
  assign n22252 = n7500 ^ n1918 ^ 1'b0 ;
  assign n22253 = n4374 & n16580 ;
  assign n22254 = n8596 & n21777 ;
  assign n22255 = n17445 ^ n842 ^ 1'b0 ;
  assign n22256 = n22255 ^ n6017 ^ 1'b0 ;
  assign n22257 = n6647 & ~n20801 ;
  assign n22258 = ~n8937 & n11433 ;
  assign n22259 = n22258 ^ n12223 ^ 1'b0 ;
  assign n22260 = n11036 ^ n5238 ^ 1'b0 ;
  assign n22261 = n2252 & n22260 ;
  assign n22262 = n13196 & n22261 ;
  assign n22263 = n22259 & n22262 ;
  assign n22264 = n489 & ~n18052 ;
  assign n22265 = n6040 & n22264 ;
  assign n22266 = n16572 & ~n22265 ;
  assign n22267 = n22266 ^ n13455 ^ 1'b0 ;
  assign n22268 = n3466 & ~n10067 ;
  assign n22269 = ~n7304 & n22268 ;
  assign n22270 = n5722 & ~n22269 ;
  assign n22271 = ~n6270 & n18828 ;
  assign n22272 = n9667 & n14805 ;
  assign n22273 = n22272 ^ n1213 ^ 1'b0 ;
  assign n22274 = n3471 & n22273 ;
  assign n22275 = ~n3567 & n4961 ;
  assign n22276 = n5167 & n22275 ;
  assign n22277 = n8508 ^ n894 ^ 1'b0 ;
  assign n22278 = n22276 | n22277 ;
  assign n22279 = n15203 ^ n1556 ^ 1'b0 ;
  assign n22280 = n17580 ^ n8992 ^ 1'b0 ;
  assign n22281 = n22280 ^ n15319 ^ n2578 ;
  assign n22282 = n4320 ^ n3221 ^ 1'b0 ;
  assign n22283 = n22282 ^ n3061 ^ 1'b0 ;
  assign n22284 = ~n12053 & n22283 ;
  assign n22285 = ~n15065 & n22284 ;
  assign n22286 = n22285 ^ n10511 ^ 1'b0 ;
  assign n22287 = n17530 & n22286 ;
  assign n22288 = n13278 ^ n3338 ^ n1090 ;
  assign n22289 = ~n13519 & n15252 ;
  assign n22290 = n12237 & n22289 ;
  assign n22291 = n2109 & ~n6610 ;
  assign n22292 = ~n6619 & n22291 ;
  assign n22293 = n22292 ^ n7611 ^ 1'b0 ;
  assign n22294 = ~n55 & n2112 ;
  assign n22295 = n2680 ^ n928 ^ 1'b0 ;
  assign n22296 = ~n5685 & n6471 ;
  assign n22297 = n22296 ^ n16138 ^ 1'b0 ;
  assign n22298 = n19971 & ~n22297 ;
  assign n22299 = n22298 ^ n232 ^ 1'b0 ;
  assign n22300 = ~n4400 & n13261 ;
  assign n22301 = ( ~n3408 & n9986 ) | ( ~n3408 & n14813 ) | ( n9986 & n14813 ) ;
  assign n22302 = n21978 ^ n11053 ^ 1'b0 ;
  assign n22303 = n19790 | n22302 ;
  assign n22304 = n4604 & n18029 ;
  assign n22305 = ~n5335 & n22304 ;
  assign n22306 = n302 & ~n22305 ;
  assign n22307 = n22306 ^ n4482 ^ 1'b0 ;
  assign n22308 = n4513 | n22193 ;
  assign n22309 = n12363 & ~n13693 ;
  assign n22310 = n940 & ~n983 ;
  assign n22311 = n7904 & n22310 ;
  assign n22312 = n11504 & n21839 ;
  assign n22313 = n1739 & ~n14910 ;
  assign n22314 = n2934 & ~n6222 ;
  assign n22315 = n10658 ^ n4968 ^ 1'b0 ;
  assign n22316 = n1683 | n22315 ;
  assign n22317 = n3254 & n17276 ;
  assign n22318 = ~n206 & n549 ;
  assign n22319 = n206 & n22318 ;
  assign n22320 = n627 & ~n22319 ;
  assign n22321 = n2310 & ~n8067 ;
  assign n22322 = n8067 & n22321 ;
  assign n22323 = n22320 & ~n22322 ;
  assign n22324 = ~n22320 & n22323 ;
  assign n22325 = n15930 ^ n6716 ^ 1'b0 ;
  assign n22326 = ~n22324 & n22325 ;
  assign n22327 = n1992 & n22326 ;
  assign n22328 = ~n22326 & n22327 ;
  assign n22329 = n7799 ^ n582 ^ 1'b0 ;
  assign n22330 = ~n1000 & n22329 ;
  assign n22331 = ~n5713 & n22330 ;
  assign n22332 = n12855 & n14850 ;
  assign n22333 = ~n3303 & n4039 ;
  assign n22334 = ~n22332 & n22333 ;
  assign n22335 = n2955 | n14051 ;
  assign n22336 = n22335 ^ n19773 ^ 1'b0 ;
  assign n22337 = n19408 & n22336 ;
  assign n22338 = n5281 & n10431 ;
  assign n22339 = n14696 & ~n22338 ;
  assign n22340 = n2203 | n2547 ;
  assign n22341 = n4565 ^ n2463 ^ 1'b0 ;
  assign n22342 = n4157 & n22341 ;
  assign n22343 = n216 | n4508 ;
  assign n22344 = n22343 ^ n7367 ^ 1'b0 ;
  assign n22345 = n2426 ^ n587 ^ 1'b0 ;
  assign n22346 = n22344 & n22345 ;
  assign n22347 = n9375 ^ n1815 ^ 1'b0 ;
  assign n22348 = n6479 | n22347 ;
  assign n22349 = ~n318 & n22348 ;
  assign n22350 = n3430 | n16065 ;
  assign n22351 = n5400 & ~n22350 ;
  assign n22352 = ~n11089 & n11228 ;
  assign n22353 = n22352 ^ n19025 ^ 1'b0 ;
  assign n22354 = ~n9062 & n22353 ;
  assign n22355 = n22354 ^ n19528 ^ 1'b0 ;
  assign n22356 = n22355 ^ n9963 ^ 1'b0 ;
  assign n22357 = ~n22351 & n22356 ;
  assign n22358 = n17527 ^ n9823 ^ 1'b0 ;
  assign n22359 = n6936 & n22358 ;
  assign n22360 = ~n4171 & n22359 ;
  assign n22361 = n10430 ^ n475 ^ 1'b0 ;
  assign n22362 = n16225 & n22361 ;
  assign n22363 = n5891 | n8945 ;
  assign n22364 = n10523 ^ n5040 ^ 1'b0 ;
  assign n22365 = ~n22363 & n22364 ;
  assign n22366 = n12485 & n18721 ;
  assign n22367 = n375 & n22366 ;
  assign n22368 = n18513 ^ n16758 ^ 1'b0 ;
  assign n22369 = n186 & ~n22368 ;
  assign n22370 = n22369 ^ n19371 ^ 1'b0 ;
  assign n22371 = n7331 & ~n10636 ;
  assign n22372 = n8488 & ~n18759 ;
  assign n22373 = n22371 & n22372 ;
  assign n22374 = n832 ^ n684 ^ 1'b0 ;
  assign n22375 = n22374 ^ n2627 ^ 1'b0 ;
  assign n22376 = n376 | n5359 ;
  assign n22377 = n22375 | n22376 ;
  assign n22378 = n1587 & ~n21973 ;
  assign n22379 = n5865 & ~n12058 ;
  assign n22380 = n12424 | n13729 ;
  assign n22381 = n22380 ^ n11556 ^ 1'b0 ;
  assign n22382 = n9090 | n21711 ;
  assign n22383 = n22381 | n22382 ;
  assign n22384 = ~n1426 & n21031 ;
  assign n22385 = n2611 & n10436 ;
  assign n22386 = n3498 & ~n20075 ;
  assign n22387 = n205 | n2463 ;
  assign n22388 = n20288 ^ n12926 ^ n2472 ;
  assign n22389 = n11192 & ~n22388 ;
  assign n22390 = n22389 ^ n9074 ^ 1'b0 ;
  assign n22391 = n880 | n13997 ;
  assign n22392 = n10395 ^ n6266 ^ 1'b0 ;
  assign n22397 = n13715 ^ n2978 ^ n2441 ;
  assign n22393 = n7687 & n13660 ;
  assign n22394 = n7634 & n22393 ;
  assign n22395 = ~n2448 & n22394 ;
  assign n22396 = ~n7406 & n22395 ;
  assign n22398 = n22397 ^ n22396 ^ 1'b0 ;
  assign n22399 = n460 | n7851 ;
  assign n22400 = n22399 ^ n6730 ^ 1'b0 ;
  assign n22401 = n545 & ~n22400 ;
  assign n22402 = n15468 & n22401 ;
  assign n22403 = n22402 ^ n17508 ^ 1'b0 ;
  assign n22404 = n3669 ^ n2773 ^ 1'b0 ;
  assign n22405 = n770 & ~n19000 ;
  assign n22410 = ~n265 & n767 ;
  assign n22406 = n12877 ^ n10142 ^ 1'b0 ;
  assign n22407 = n13422 | n22406 ;
  assign n22408 = n13422 & ~n22407 ;
  assign n22409 = n2624 & ~n22408 ;
  assign n22411 = n22410 ^ n22409 ^ 1'b0 ;
  assign n22413 = n802 | n7678 ;
  assign n22414 = n22413 ^ n7769 ^ 1'b0 ;
  assign n22412 = n1838 & ~n6016 ;
  assign n22415 = n22414 ^ n22412 ^ 1'b0 ;
  assign n22416 = n412 & ~n17326 ;
  assign n22417 = ~n498 & n8265 ;
  assign n22418 = n22417 ^ n11765 ^ 1'b0 ;
  assign n22419 = n9911 & ~n13715 ;
  assign n22420 = n2324 | n6412 ;
  assign n22421 = ~n684 & n2183 ;
  assign n22422 = n17903 & n22421 ;
  assign n22423 = n6946 ^ n3604 ^ 1'b0 ;
  assign n22424 = ~n2851 & n22423 ;
  assign n22425 = n10292 & n22424 ;
  assign n22426 = n5065 ^ n2121 ^ 1'b0 ;
  assign n22427 = n19020 & n22426 ;
  assign n22428 = n2925 & ~n8137 ;
  assign n22429 = n22428 ^ n3679 ^ 1'b0 ;
  assign n22430 = n6571 ^ n4195 ^ 1'b0 ;
  assign n22431 = n7160 & n22430 ;
  assign n22432 = n1250 ^ n495 ^ 1'b0 ;
  assign n22433 = n22432 ^ n19414 ^ 1'b0 ;
  assign n22434 = n487 & ~n8221 ;
  assign n22435 = n4407 ^ n3065 ^ 1'b0 ;
  assign n22436 = ~n10386 & n22435 ;
  assign n22437 = ~n3972 & n22436 ;
  assign n22438 = n22437 ^ n17525 ^ 1'b0 ;
  assign n22439 = n15467 ^ n4222 ^ 1'b0 ;
  assign n22440 = n7792 ^ n7383 ^ 1'b0 ;
  assign n22441 = n4312 | n22440 ;
  assign n22442 = ~n1254 & n22441 ;
  assign n22444 = n688 & ~n1097 ;
  assign n22443 = n14125 & ~n17339 ;
  assign n22445 = n22444 ^ n22443 ^ 1'b0 ;
  assign n22448 = n6983 | n7754 ;
  assign n22449 = n7465 | n22448 ;
  assign n22450 = n22449 ^ n6986 ^ 1'b0 ;
  assign n22446 = ~n1794 & n2572 ;
  assign n22447 = n7506 & n22446 ;
  assign n22451 = n22450 ^ n22447 ^ 1'b0 ;
  assign n22452 = n7797 ^ n495 ^ 1'b0 ;
  assign n22453 = n8352 | n8823 ;
  assign n22454 = n2819 & n22453 ;
  assign n22455 = n22454 ^ n18187 ^ 1'b0 ;
  assign n22456 = n2082 & n2648 ;
  assign n22457 = n22456 ^ n9357 ^ 1'b0 ;
  assign n22458 = n4567 & ~n10984 ;
  assign n22459 = ~n22457 & n22458 ;
  assign n22460 = n22459 ^ n21420 ^ 1'b0 ;
  assign n22461 = n6862 & ~n7608 ;
  assign n22462 = n22461 ^ n10476 ^ n2162 ;
  assign n22463 = n21885 | n22462 ;
  assign n22464 = n17590 ^ n13777 ^ 1'b0 ;
  assign n22465 = n3423 & ~n22464 ;
  assign n22466 = n627 & n8656 ;
  assign n22467 = n1584 | n11533 ;
  assign n22468 = n1584 & ~n22467 ;
  assign n22469 = n157 & ~n22468 ;
  assign n22470 = n22468 & n22469 ;
  assign n22471 = n294 & ~n10097 ;
  assign n22472 = n19575 & n19701 ;
  assign n22473 = n8812 & n22472 ;
  assign n22474 = n367 & n22473 ;
  assign n22475 = n2784 | n7148 ;
  assign n22476 = n16 & ~n233 ;
  assign n22477 = n122 | n2955 ;
  assign n22478 = n22477 ^ n679 ^ 1'b0 ;
  assign n22479 = n4219 | n22478 ;
  assign n22480 = n1677 & ~n22479 ;
  assign n22481 = ~n164 & n10728 ;
  assign n22482 = ~n2990 & n22481 ;
  assign n22483 = n10364 ^ n2991 ^ 1'b0 ;
  assign n22484 = n4155 & ~n10650 ;
  assign n22485 = n22484 ^ n4976 ^ 1'b0 ;
  assign n22486 = n7429 | n12806 ;
  assign n22487 = n22485 & ~n22486 ;
  assign n22488 = n5978 ^ n5469 ^ 1'b0 ;
  assign n22489 = ~n22487 & n22488 ;
  assign n22490 = n7596 & ~n17567 ;
  assign n22491 = ~n14474 & n22490 ;
  assign n22492 = n20316 ^ n10374 ^ 1'b0 ;
  assign n22493 = n12728 ^ n2885 ^ 1'b0 ;
  assign n22494 = n22493 ^ n1337 ^ 1'b0 ;
  assign n22495 = n11241 & ~n21136 ;
  assign n22496 = n3197 ^ n207 ^ 1'b0 ;
  assign n22497 = n22496 ^ n15052 ^ 1'b0 ;
  assign n22498 = ~n131 & n4913 ;
  assign n22499 = n8052 | n10451 ;
  assign n22500 = n3180 & n12236 ;
  assign n22501 = ~n722 & n22500 ;
  assign n22502 = ~n22499 & n22501 ;
  assign n22503 = n7388 ^ n340 ^ 1'b0 ;
  assign n22504 = n8251 & ~n20264 ;
  assign n22506 = n17776 ^ n9476 ^ n1324 ;
  assign n22505 = n8276 | n18292 ;
  assign n22507 = n22506 ^ n22505 ^ 1'b0 ;
  assign n22508 = n7497 & n10282 ;
  assign n22509 = n17255 ^ n16346 ^ 1'b0 ;
  assign n22521 = n123 & ~n1499 ;
  assign n22522 = ~n123 & n22521 ;
  assign n22523 = n1588 & ~n7269 ;
  assign n22524 = n22522 & n22523 ;
  assign n22510 = n1701 & n7894 ;
  assign n22511 = ~n7894 & n22510 ;
  assign n22512 = n22511 ^ n1203 ^ 1'b0 ;
  assign n22513 = ~n133 & n14295 ;
  assign n22514 = n300 & n22513 ;
  assign n22515 = n22512 & n22514 ;
  assign n22516 = ~n22512 & n22515 ;
  assign n22517 = ~n636 & n22516 ;
  assign n22518 = n318 | n12742 ;
  assign n22519 = n12742 & ~n22518 ;
  assign n22520 = n22517 | n22519 ;
  assign n22525 = n22524 ^ n22520 ^ 1'b0 ;
  assign n22526 = n88 & n19976 ;
  assign n22527 = ~n21007 & n22526 ;
  assign n22528 = n6224 & n8679 ;
  assign n22529 = n22527 & n22528 ;
  assign n22530 = n3529 & n3746 ;
  assign n22531 = ~n1370 & n7380 ;
  assign n22532 = ( ~n1292 & n15966 ) | ( ~n1292 & n22531 ) | ( n15966 & n22531 ) ;
  assign n22533 = n15524 ^ n1860 ^ 1'b0 ;
  assign n22534 = ~n8162 & n22533 ;
  assign n22535 = n7378 ^ n3985 ^ 1'b0 ;
  assign n22536 = ~n844 & n8672 ;
  assign n22537 = n15434 & ~n22536 ;
  assign n22538 = n22535 | n22537 ;
  assign n22539 = ~n1020 & n1260 ;
  assign n22540 = ~n5327 & n6609 ;
  assign n22541 = n14961 & ~n16821 ;
  assign n22542 = n7490 & n22541 ;
  assign n22543 = n2003 & n7892 ;
  assign n22544 = n1688 & ~n22543 ;
  assign n22545 = n9135 & n14165 ;
  assign n22546 = n940 & n6218 ;
  assign n22547 = ~n5273 & n22546 ;
  assign n22548 = n22547 ^ n22175 ^ 1'b0 ;
  assign n22549 = n8967 ^ n323 ^ 1'b0 ;
  assign n22550 = n13588 & n22549 ;
  assign n22551 = n19544 & n22550 ;
  assign n22552 = n10322 | n22462 ;
  assign n22553 = n22551 & ~n22552 ;
  assign n22560 = n977 & n1958 ;
  assign n22561 = n799 & n22560 ;
  assign n22554 = n917 & n1139 ;
  assign n22555 = n2303 & n12862 ;
  assign n22556 = n18769 & n22555 ;
  assign n22557 = n11355 | n22556 ;
  assign n22558 = n22554 | n22557 ;
  assign n22559 = n22558 ^ n15145 ^ 1'b0 ;
  assign n22562 = n22561 ^ n22559 ^ 1'b0 ;
  assign n22563 = n22553 | n22562 ;
  assign n22564 = n9227 & ~n9965 ;
  assign n22565 = n4460 | n13312 ;
  assign n22566 = n4642 | n5702 ;
  assign n22567 = ~n1782 & n14142 ;
  assign n22568 = n9846 & n22567 ;
  assign n22569 = n6217 ^ n2142 ^ 1'b0 ;
  assign n22570 = n13870 ^ n4155 ^ 1'b0 ;
  assign n22571 = n2155 & ~n3431 ;
  assign n22572 = n186 & ~n19175 ;
  assign n22573 = n22571 & n22572 ;
  assign n22574 = n2992 & n21375 ;
  assign n22575 = n22574 ^ n501 ^ 1'b0 ;
  assign n22576 = n6682 ^ n2099 ^ 1'b0 ;
  assign n22577 = n20713 ^ n3449 ^ 1'b0 ;
  assign n22578 = ~n13094 & n22577 ;
  assign n22579 = ( n88 & n3533 ) | ( n88 & ~n22578 ) | ( n3533 & ~n22578 ) ;
  assign n22580 = n425 & n9222 ;
  assign n22583 = n58 & ~n13108 ;
  assign n22581 = n5776 ^ n5574 ^ 1'b0 ;
  assign n22582 = n2874 & n22581 ;
  assign n22584 = n22583 ^ n22582 ^ 1'b0 ;
  assign n22585 = n12007 ^ n3106 ^ 1'b0 ;
  assign n22586 = n161 | n22585 ;
  assign n22587 = n22586 ^ n3653 ^ 1'b0 ;
  assign n22588 = n592 | n22587 ;
  assign n22589 = n19169 & n20055 ;
  assign n22590 = n22589 ^ n3007 ^ 1'b0 ;
  assign n22591 = n21101 ^ n2980 ^ 1'b0 ;
  assign n22592 = n1798 & ~n11239 ;
  assign n22593 = n3839 ^ n117 ^ 1'b0 ;
  assign n22594 = n13199 | n22593 ;
  assign n22595 = n7508 | n22594 ;
  assign n22596 = n8053 ^ n2924 ^ 1'b0 ;
  assign n22597 = ~n12082 & n22596 ;
  assign n22598 = n1679 & n22597 ;
  assign n22599 = n13170 & n22598 ;
  assign n22600 = n18579 & n22599 ;
  assign n22601 = n2506 ^ n758 ^ 1'b0 ;
  assign n22602 = n6493 ^ n5297 ^ 1'b0 ;
  assign n22603 = n22601 | n22602 ;
  assign n22604 = n22603 ^ n1704 ^ 1'b0 ;
  assign n22605 = ~n3371 & n7130 ;
  assign n22606 = n22605 ^ n2317 ^ 1'b0 ;
  assign n22607 = ~n7500 & n22606 ;
  assign n22608 = n22607 ^ n128 ^ 1'b0 ;
  assign n22609 = ~n6406 & n7624 ;
  assign n22610 = ~n4716 & n5955 ;
  assign n22611 = ~n13238 & n22610 ;
  assign n22612 = ~n22609 & n22611 ;
  assign n22613 = n20974 ^ n135 ^ 1'b0 ;
  assign n22614 = n1947 | n2225 ;
  assign n22615 = n4531 | n13455 ;
  assign n22616 = n9062 & ~n13548 ;
  assign n22617 = n883 & n19420 ;
  assign n22618 = n1480 & n22617 ;
  assign n22619 = n556 & ~n22618 ;
  assign n22620 = n12441 ^ n2377 ^ 1'b0 ;
  assign n22621 = n19618 | n22620 ;
  assign n22622 = ~n2136 & n22621 ;
  assign n22623 = n2244 | n5977 ;
  assign n22624 = n22623 ^ n1895 ^ n378 ;
  assign n22625 = n18484 ^ n2486 ^ 1'b0 ;
  assign n22627 = n12272 & ~n13483 ;
  assign n22626 = ~n4424 & n8656 ;
  assign n22628 = n22627 ^ n22626 ^ 1'b0 ;
  assign n22632 = n404 & ~n3069 ;
  assign n22629 = n5899 ^ n364 ^ 1'b0 ;
  assign n22630 = ~n644 & n22629 ;
  assign n22631 = n22630 ^ n4765 ^ 1'b0 ;
  assign n22633 = n22632 ^ n22631 ^ n19390 ;
  assign n22634 = n10107 & ~n18523 ;
  assign n22635 = ~n4873 & n20762 ;
  assign n22639 = n2768 ^ n556 ^ 1'b0 ;
  assign n22640 = n229 & ~n22639 ;
  assign n22636 = n9588 & ~n11612 ;
  assign n22637 = ~n5154 & n22636 ;
  assign n22638 = n22637 ^ n1714 ^ 1'b0 ;
  assign n22641 = n22640 ^ n22638 ^ 1'b0 ;
  assign n22642 = n1198 | n5749 ;
  assign n22643 = n13720 | n22642 ;
  assign n22644 = n9666 & n22643 ;
  assign n22645 = n1497 | n2978 ;
  assign n22646 = n3821 & ~n22645 ;
  assign n22648 = n13220 ^ n4732 ^ 1'b0 ;
  assign n22649 = n5183 & ~n22648 ;
  assign n22647 = n8128 & ~n12702 ;
  assign n22650 = n22649 ^ n22647 ^ 1'b0 ;
  assign n22651 = n1117 | n9247 ;
  assign n22652 = n11201 | n22651 ;
  assign n22653 = ( n6224 & n8891 ) | ( n6224 & n10076 ) | ( n8891 & n10076 ) ;
  assign n22654 = ~n10634 & n22653 ;
  assign n22656 = n5950 ^ n388 ^ 1'b0 ;
  assign n22657 = n2639 | n22656 ;
  assign n22655 = n6471 & n8409 ;
  assign n22658 = n22657 ^ n22655 ^ 1'b0 ;
  assign n22659 = n6822 & ~n15748 ;
  assign n22660 = n8863 | n14786 ;
  assign n22661 = n22660 ^ n1817 ^ n578 ;
  assign n22662 = n2200 & n9242 ;
  assign n22663 = ~n11451 & n22662 ;
  assign n22664 = n1285 & ~n6040 ;
  assign n22665 = ~n1684 & n22664 ;
  assign n22666 = ( n1246 & n22663 ) | ( n1246 & n22665 ) | ( n22663 & n22665 ) ;
  assign n22667 = n7944 & ~n22666 ;
  assign n22668 = n22667 ^ n3540 ^ 1'b0 ;
  assign n22669 = ~n14370 & n17733 ;
  assign n22670 = ~n22163 & n22669 ;
  assign n22671 = n11624 ^ n1961 ^ 1'b0 ;
  assign n22672 = n11260 ^ n10835 ^ n1345 ;
  assign n22673 = n21411 ^ n3885 ^ 1'b0 ;
  assign n22674 = ~n17038 & n22673 ;
  assign n22675 = n21999 ^ n10983 ^ 1'b0 ;
  assign n22676 = n9291 | n22675 ;
  assign n22677 = n2819 ^ n1789 ^ 1'b0 ;
  assign n22678 = n17050 ^ n3121 ^ 1'b0 ;
  assign n22679 = n3783 | n22678 ;
  assign n22680 = n22679 ^ n2546 ^ 1'b0 ;
  assign n22681 = ~n139 & n22680 ;
  assign n22682 = n4559 ^ n1235 ^ 1'b0 ;
  assign n22683 = n9010 & n22682 ;
  assign n22684 = n2288 | n12853 ;
  assign n22685 = n22684 ^ n7668 ^ 1'b0 ;
  assign n22686 = n2536 & n6157 ;
  assign n22687 = n1349 | n4533 ;
  assign n22688 = n2936 & n22687 ;
  assign n22689 = n7512 | n11948 ;
  assign n22690 = ~n3156 & n3423 ;
  assign n22691 = n22690 ^ n7526 ^ 1'b0 ;
  assign n22692 = ~n8766 & n22163 ;
  assign n22693 = n364 | n6962 ;
  assign n22694 = n9592 & ~n13082 ;
  assign n22695 = ~n22693 & n22694 ;
  assign n22696 = n22695 ^ n1926 ^ 1'b0 ;
  assign n22697 = n9596 ^ n9211 ^ n133 ;
  assign n22698 = n22697 ^ n20806 ^ n5424 ;
  assign n22699 = n1934 & ~n20495 ;
  assign n22700 = ~n3454 & n22699 ;
  assign n22701 = ~n538 & n2773 ;
  assign n22702 = n22701 ^ n13652 ^ 1'b0 ;
  assign n22703 = ~n22700 & n22702 ;
  assign n22704 = n22703 ^ n6277 ^ 1'b0 ;
  assign n22705 = n3465 | n20841 ;
  assign n22706 = n21635 ^ n14916 ^ 1'b0 ;
  assign n22707 = n4062 | n19935 ;
  assign n22708 = n22707 ^ n16693 ^ 1'b0 ;
  assign n22709 = ~n1497 & n6107 ;
  assign n22710 = n15576 | n22709 ;
  assign n22711 = n16658 & ~n22710 ;
  assign n22712 = n22711 ^ n1826 ^ 1'b0 ;
  assign n22713 = n15201 ^ n82 ^ 1'b0 ;
  assign n22714 = n547 & n22713 ;
  assign n22715 = n3717 & ~n4927 ;
  assign n22716 = n18363 & n22715 ;
  assign n22717 = n6645 & n22716 ;
  assign n22718 = n6682 & n9108 ;
  assign n22719 = ~n7579 & n22718 ;
  assign n22720 = n5827 & ~n8674 ;
  assign n22721 = n2585 ^ n701 ^ 1'b0 ;
  assign n22722 = n22721 ^ n11478 ^ 1'b0 ;
  assign n22724 = n3837 | n9578 ;
  assign n22725 = n22724 ^ n14647 ^ 1'b0 ;
  assign n22723 = n3744 & n10791 ;
  assign n22726 = n22725 ^ n22723 ^ 1'b0 ;
  assign n22727 = n3771 ^ n928 ^ 1'b0 ;
  assign n22728 = ~n14652 & n22727 ;
  assign n22729 = n5070 | n18508 ;
  assign n22730 = n9877 | n22729 ;
  assign n22731 = n4753 ^ n2726 ^ 1'b0 ;
  assign n22732 = n5205 ^ n2531 ^ 1'b0 ;
  assign n22733 = n22732 ^ n9088 ^ 1'b0 ;
  assign n22734 = n17843 ^ n14539 ^ 1'b0 ;
  assign n22735 = n22414 | n22734 ;
  assign n22736 = n15368 | n18923 ;
  assign n22737 = n3262 ^ n2569 ^ 1'b0 ;
  assign n22738 = n7464 ^ n3506 ^ 1'b0 ;
  assign n22739 = n9520 | n22738 ;
  assign n22740 = ~n21475 & n22739 ;
  assign n22741 = n6560 & n9911 ;
  assign n22742 = ~n9033 & n22741 ;
  assign n22743 = ~n837 & n11973 ;
  assign n22744 = n22743 ^ n8263 ^ 1'b0 ;
  assign n22745 = ~n22742 & n22744 ;
  assign n22746 = n22745 ^ n11764 ^ 1'b0 ;
  assign n22747 = ~n2677 & n9180 ;
  assign n22748 = n22747 ^ n22459 ^ n5194 ;
  assign n22749 = n7589 | n9881 ;
  assign n22750 = n3845 | n21221 ;
  assign n22751 = n8596 & ~n22750 ;
  assign n22752 = n7578 ^ n6098 ^ 1'b0 ;
  assign n22753 = n1431 & ~n22752 ;
  assign n22754 = n8354 & ~n16733 ;
  assign n22755 = n663 & n18795 ;
  assign n22756 = ( n2876 & ~n9803 ) | ( n2876 & n22755 ) | ( ~n9803 & n22755 ) ;
  assign n22757 = n8971 ^ n1165 ^ 1'b0 ;
  assign n22758 = n2155 | n22757 ;
  assign n22759 = n22758 ^ n3692 ^ 1'b0 ;
  assign n22761 = n3346 & n9023 ;
  assign n22762 = ~n12073 & n22761 ;
  assign n22763 = n13554 & ~n22762 ;
  assign n22764 = n11248 & n22763 ;
  assign n22760 = n3946 | n9155 ;
  assign n22765 = n22764 ^ n22760 ^ 1'b0 ;
  assign n22766 = n6646 & n7290 ;
  assign n22767 = n6019 & n22766 ;
  assign n22768 = n16307 ^ n3037 ^ n440 ;
  assign n22769 = n2096 & ~n9899 ;
  assign n22770 = n22769 ^ n13620 ^ 1'b0 ;
  assign n22771 = ~n2961 & n10465 ;
  assign n22772 = n22771 ^ n3509 ^ 1'b0 ;
  assign n22774 = n2467 & ~n5299 ;
  assign n22773 = n10974 & ~n11444 ;
  assign n22775 = n22774 ^ n22773 ^ 1'b0 ;
  assign n22776 = n5225 & ~n16507 ;
  assign n22777 = n12441 | n22776 ;
  assign n22778 = ~n7694 & n22777 ;
  assign n22779 = n19700 & n22778 ;
  assign n22780 = n16952 ^ n10504 ^ 1'b0 ;
  assign n22781 = n10064 & n14941 ;
  assign n22782 = n16411 & n16849 ;
  assign n22783 = n2165 & n18563 ;
  assign n22784 = n4866 & n22783 ;
  assign n22785 = n22784 ^ n1748 ^ 1'b0 ;
  assign n22786 = n13660 & ~n18782 ;
  assign n22787 = n10446 & n22786 ;
  assign n22788 = n4741 & n14478 ;
  assign n22789 = n1302 & n22788 ;
  assign n22790 = n17723 ^ n4062 ^ 1'b0 ;
  assign n22791 = n6365 & ~n8688 ;
  assign n22792 = n22790 & n22791 ;
  assign n22793 = n613 | n6740 ;
  assign n22794 = n22793 ^ n9927 ^ 1'b0 ;
  assign n22795 = n22794 ^ n8755 ^ 1'b0 ;
  assign n22796 = n3664 | n16519 ;
  assign n22797 = n22796 ^ n4318 ^ 1'b0 ;
  assign n22798 = ~n7269 & n9159 ;
  assign n22799 = ~n558 & n18387 ;
  assign n22800 = n8183 & n22799 ;
  assign n22801 = n3138 & ~n22800 ;
  assign n22802 = n22801 ^ n12643 ^ 1'b0 ;
  assign n22803 = n22802 ^ n18039 ^ 1'b0 ;
  assign n22804 = n22798 & n22803 ;
  assign n22805 = n2948 & n17795 ;
  assign n22806 = n22805 ^ n13864 ^ 1'b0 ;
  assign n22807 = n15115 & n15659 ;
  assign n22808 = ~n1226 & n15760 ;
  assign n22809 = n22808 ^ n13948 ^ 1'b0 ;
  assign n22810 = n10674 | n11212 ;
  assign n22811 = n3376 | n22810 ;
  assign n22812 = n3670 ^ n200 ^ 1'b0 ;
  assign n22813 = n3101 & n14490 ;
  assign n22814 = ~n22812 & n22813 ;
  assign n22815 = n3459 ^ n2399 ^ 1'b0 ;
  assign n22816 = ~n22814 & n22815 ;
  assign n22817 = n22816 ^ n719 ^ 1'b0 ;
  assign n22818 = n216 & ~n8446 ;
  assign n22819 = n22818 ^ n15087 ^ 1'b0 ;
  assign n22820 = n22819 ^ n19785 ^ n8656 ;
  assign n22821 = n792 | n22820 ;
  assign n22822 = n17621 | n22821 ;
  assign n22823 = ~n6502 & n22822 ;
  assign n22824 = n10159 & n22325 ;
  assign n22825 = n15561 ^ n1415 ^ 1'b0 ;
  assign n22826 = n22824 & n22825 ;
  assign n22827 = n22826 ^ n9697 ^ 1'b0 ;
  assign n22828 = n5625 & ~n22827 ;
  assign n22829 = n10457 ^ n8365 ^ 1'b0 ;
  assign n22830 = ~n1396 & n10395 ;
  assign n22831 = ~n11586 & n22830 ;
  assign n22832 = n2594 & ~n18789 ;
  assign n22833 = n6315 & ~n18882 ;
  assign n22834 = n21081 ^ n10101 ^ 1'b0 ;
  assign n22835 = n22833 & ~n22834 ;
  assign n22836 = n3042 & ~n10905 ;
  assign n22837 = ~n7666 & n7736 ;
  assign n22838 = ~n406 & n1406 ;
  assign n22839 = n2789 ^ n2635 ^ 1'b0 ;
  assign n22840 = n635 & ~n22839 ;
  assign n22841 = n9086 ^ n758 ^ 1'b0 ;
  assign n22842 = n1817 | n22841 ;
  assign n22843 = n17451 | n22842 ;
  assign n22844 = ~n21423 & n22843 ;
  assign n22845 = n22840 & n22844 ;
  assign n22846 = n4875 ^ n4392 ^ 1'b0 ;
  assign n22847 = n6738 | n22846 ;
  assign n22848 = n22847 ^ n3626 ^ 1'b0 ;
  assign n22849 = n4304 & n22848 ;
  assign n22850 = n4126 ^ n3188 ^ 1'b0 ;
  assign n22851 = n14683 ^ n964 ^ 1'b0 ;
  assign n22852 = n11377 ^ n8620 ^ 1'b0 ;
  assign n22853 = n8763 & n22852 ;
  assign n22854 = n251 & ~n6126 ;
  assign n22855 = ~n18379 & n22854 ;
  assign n22856 = ( n4495 & n11000 ) | ( n4495 & ~n20585 ) | ( n11000 & ~n20585 ) ;
  assign n22857 = n13461 ^ n12441 ^ 1'b0 ;
  assign n22858 = n339 & ~n5749 ;
  assign n22859 = n1179 & n22858 ;
  assign n22860 = n5210 & n5348 ;
  assign n22861 = n443 & ~n22860 ;
  assign n22862 = x0 & ~n19 ;
  assign n22863 = ~n433 & n22862 ;
  assign n22864 = n8198 | n22863 ;
  assign n22865 = n2294 | n18025 ;
  assign n22866 = ~n7400 & n17948 ;
  assign n22867 = n14333 & n22866 ;
  assign n22868 = n22867 ^ n9898 ^ 1'b0 ;
  assign n22869 = n17947 | n22868 ;
  assign n22870 = n1344 | n22869 ;
  assign n22871 = n3882 & n11077 ;
  assign n22872 = n22871 ^ n9873 ^ 1'b0 ;
  assign n22873 = n2584 ^ n542 ^ 1'b0 ;
  assign n22874 = n3988 & ~n13480 ;
  assign n22875 = n461 | n5194 ;
  assign n22876 = n22875 ^ n4756 ^ 1'b0 ;
  assign n22877 = n8613 ^ n1184 ^ 1'b0 ;
  assign n22878 = ~n22876 & n22877 ;
  assign n22879 = n769 | n13242 ;
  assign n22880 = n5850 & ~n22543 ;
  assign n22881 = ~n7201 & n11709 ;
  assign n22882 = n22880 & n22881 ;
  assign n22883 = ~n294 & n1750 ;
  assign n22884 = ~n6008 & n22883 ;
  assign n22885 = n22884 ^ n14742 ^ 1'b0 ;
  assign n22886 = n167 & n11556 ;
  assign n22887 = n3741 & ~n22886 ;
  assign n22888 = n10047 & n12469 ;
  assign n22889 = n19691 ^ n5465 ^ n2377 ;
  assign n22890 = n10390 ^ n1390 ^ 1'b0 ;
  assign n22891 = ~n1396 & n3369 ;
  assign n22892 = n22890 & n22891 ;
  assign n22893 = n12393 ^ n6416 ^ 1'b0 ;
  assign n22894 = n19978 ^ n10328 ^ 1'b0 ;
  assign n22895 = n1838 & ~n22894 ;
  assign n22896 = ~n5505 & n22895 ;
  assign n22897 = n22896 ^ n21836 ^ 1'b0 ;
  assign n22898 = n9091 & ~n22897 ;
  assign n22899 = n187 | n8415 ;
  assign n22900 = n22899 ^ n12784 ^ 1'b0 ;
  assign n22901 = n3321 & ~n22900 ;
  assign n22902 = n960 & n20578 ;
  assign n22903 = ~n20483 & n22902 ;
  assign n22907 = n200 & n7053 ;
  assign n22906 = n13253 & ~n15124 ;
  assign n22908 = n22907 ^ n22906 ^ 1'b0 ;
  assign n22904 = n10052 & n10797 ;
  assign n22905 = n7649 & ~n22904 ;
  assign n22909 = n22908 ^ n22905 ^ 1'b0 ;
  assign n22910 = ~n9837 & n19165 ;
  assign n22911 = n22910 ^ n6442 ^ 1'b0 ;
  assign n22912 = n7879 | n10004 ;
  assign n22913 = n4293 ^ n1787 ^ 1'b0 ;
  assign n22914 = n1763 & n22913 ;
  assign n22915 = n7383 | n14470 ;
  assign n22916 = n4626 ^ n1175 ^ 1'b0 ;
  assign n22917 = n7652 ^ n1715 ^ 1'b0 ;
  assign n22918 = n8246 | n22917 ;
  assign n22919 = n22918 ^ n7159 ^ 1'b0 ;
  assign n22920 = n14861 ^ n12423 ^ 1'b0 ;
  assign n22921 = ~n6442 & n15606 ;
  assign n22922 = n22921 ^ n3803 ^ 1'b0 ;
  assign n22923 = n9227 ^ n6849 ^ 1'b0 ;
  assign n22924 = n5639 & ~n22923 ;
  assign n22925 = n22924 ^ n13343 ^ 1'b0 ;
  assign n22926 = n2849 & n22925 ;
  assign n22927 = ~n2607 & n19843 ;
  assign n22928 = ~n458 & n12700 ;
  assign n22929 = ~n22927 & n22928 ;
  assign n22930 = n16360 & n22929 ;
  assign n22931 = n13155 & ~n19990 ;
  assign n22932 = n7827 & n22931 ;
  assign n22934 = n806 & ~n8525 ;
  assign n22935 = n2626 | n6028 ;
  assign n22936 = n22934 | n22935 ;
  assign n22933 = n726 & ~n7338 ;
  assign n22937 = n22936 ^ n22933 ^ 1'b0 ;
  assign n22938 = n3135 ^ n2012 ^ 1'b0 ;
  assign n22939 = x2 & ~n22938 ;
  assign n22940 = ~n9737 & n22939 ;
  assign n22941 = ~n21072 & n22940 ;
  assign n22942 = ~n3980 & n11178 ;
  assign n22943 = n22942 ^ n929 ^ 1'b0 ;
  assign n22944 = n22941 | n22943 ;
  assign n22945 = n15307 & ~n22944 ;
  assign n22946 = n10788 ^ n6562 ^ 1'b0 ;
  assign n22947 = n21126 ^ n17169 ^ 1'b0 ;
  assign n22948 = n88 & ~n20403 ;
  assign n22949 = ~n18131 & n22948 ;
  assign n22950 = n11910 ^ n7112 ^ n1486 ;
  assign n22951 = n2571 & n22950 ;
  assign n22952 = ~n423 & n22951 ;
  assign n22953 = n34 | n22952 ;
  assign n22954 = n22949 & ~n22953 ;
  assign n22955 = n13856 & n15717 ;
  assign n22956 = n2633 | n3931 ;
  assign n22957 = ~n2991 & n5971 ;
  assign n22958 = n22957 ^ n432 ^ 1'b0 ;
  assign n22959 = n710 & n10798 ;
  assign n22960 = ~n1701 & n22959 ;
  assign n22961 = n21635 ^ n15264 ^ 1'b0 ;
  assign n22962 = n5331 | n8419 ;
  assign n22963 = n22962 ^ n8825 ^ 1'b0 ;
  assign n22964 = n9561 | n15434 ;
  assign n22965 = n22964 ^ n14779 ^ 1'b0 ;
  assign n22966 = n958 ^ n297 ^ 1'b0 ;
  assign n22967 = n5524 & ~n22966 ;
  assign n22968 = n22343 ^ n6334 ^ 1'b0 ;
  assign n22969 = n1004 & n22968 ;
  assign n22970 = n22271 ^ n6210 ^ 1'b0 ;
  assign n22971 = ~n6940 & n22970 ;
  assign n22972 = n22971 ^ n11298 ^ 1'b0 ;
  assign n22975 = n940 & n8582 ;
  assign n22976 = n22975 ^ n4799 ^ 1'b0 ;
  assign n22973 = n22907 ^ n3793 ^ 1'b0 ;
  assign n22974 = ~n3589 & n22973 ;
  assign n22977 = n22976 ^ n22974 ^ 1'b0 ;
  assign n22978 = n4853 | n22977 ;
  assign n22979 = n22978 ^ n12632 ^ 1'b0 ;
  assign n22980 = n1396 | n16315 ;
  assign n22981 = n9447 & ~n22980 ;
  assign n22982 = n22981 ^ n4084 ^ 1'b0 ;
  assign n22983 = n22979 & n22982 ;
  assign n22984 = n12803 & n17867 ;
  assign n22985 = n814 & ~n9692 ;
  assign n22986 = ~n10107 & n22985 ;
  assign n22987 = n1169 | n22986 ;
  assign n22988 = n12231 & n22987 ;
  assign n22989 = ~n4525 & n21735 ;
  assign n22990 = n1431 & ~n10876 ;
  assign n22991 = n1080 | n22990 ;
  assign n22992 = n22991 ^ n962 ^ 1'b0 ;
  assign n22993 = n6540 & n22992 ;
  assign n22994 = ~n11471 & n22993 ;
  assign n22995 = n22994 ^ n128 ^ 1'b0 ;
  assign n22996 = n2318 | n10105 ;
  assign n22997 = n12073 & ~n22996 ;
  assign n22998 = n22997 ^ n20492 ^ 1'b0 ;
  assign n22999 = n5406 ^ n2985 ^ 1'b0 ;
  assign n23000 = n22999 ^ n708 ^ 1'b0 ;
  assign n23001 = ~n159 & n22248 ;
  assign n23002 = n8460 ^ n4686 ^ 1'b0 ;
  assign n23003 = n11403 & ~n23002 ;
  assign n23004 = n19837 & n23003 ;
  assign n23005 = ~n22681 & n23004 ;
  assign n23006 = n3223 | n13022 ;
  assign n23007 = ~n468 & n12000 ;
  assign n23008 = ~n3663 & n4781 ;
  assign n23009 = n11265 & n23008 ;
  assign n23010 = n16295 & n23009 ;
  assign n23011 = n11972 & n20508 ;
  assign n23012 = n1441 & n23011 ;
  assign n23013 = n17249 & n20027 ;
  assign n23014 = n23012 | n23013 ;
  assign n23015 = n388 & ~n3808 ;
  assign n23016 = n23015 ^ n16661 ^ 1'b0 ;
  assign n23017 = n4355 ^ n296 ^ 1'b0 ;
  assign n23018 = n13727 ^ n1167 ^ 1'b0 ;
  assign n23019 = n23017 & n23018 ;
  assign n23020 = n17519 & n23019 ;
  assign n23021 = n16697 | n17282 ;
  assign n23022 = ~n2294 & n4575 ;
  assign n23023 = n23022 ^ n10760 ^ 1'b0 ;
  assign n23024 = n9889 | n23023 ;
  assign n23025 = n20254 | n23024 ;
  assign n23026 = n2194 | n8787 ;
  assign n23027 = n23026 ^ n11804 ^ 1'b0 ;
  assign n23028 = n8627 ^ n5575 ^ 1'b0 ;
  assign n23029 = n15862 ^ n7497 ^ 1'b0 ;
  assign n23030 = ~n960 & n8897 ;
  assign n23031 = n9719 ^ n156 ^ 1'b0 ;
  assign n23032 = n622 & n23031 ;
  assign n23033 = ~n1690 & n4872 ;
  assign n23034 = ~n23032 & n23033 ;
  assign n23035 = n6194 ^ n2759 ^ 1'b0 ;
  assign n23036 = ~n758 & n4117 ;
  assign n23037 = n9360 & n19720 ;
  assign n23038 = ~n477 & n3178 ;
  assign n23039 = n8653 | n15244 ;
  assign n23040 = n7783 ^ n7217 ^ 1'b0 ;
  assign n23041 = n23039 | n23040 ;
  assign n23043 = n1626 & n4166 ;
  assign n23044 = n7780 & ~n14537 ;
  assign n23045 = ~n23043 & n23044 ;
  assign n23042 = n96 | n15792 ;
  assign n23046 = n23045 ^ n23042 ^ 1'b0 ;
  assign n23047 = n6880 | n9788 ;
  assign n23048 = n21509 ^ n10060 ^ n665 ;
  assign n23049 = n6876 & ~n23048 ;
  assign n23050 = n15966 ^ n7706 ^ 1'b0 ;
  assign n23051 = n12501 | n23050 ;
  assign n23052 = n23051 ^ n10119 ^ 1'b0 ;
  assign n23053 = n108 | n493 ;
  assign n23054 = n23053 ^ n553 ^ 1'b0 ;
  assign n23055 = n19000 & n23054 ;
  assign n23056 = n2248 & ~n16906 ;
  assign n23057 = n23056 ^ n1845 ^ 1'b0 ;
  assign n23058 = ~n14316 & n23057 ;
  assign n23059 = n22057 ^ n5903 ^ 1'b0 ;
  assign n23060 = n483 | n14457 ;
  assign n23061 = n23060 ^ x0 ^ 1'b0 ;
  assign n23062 = n142 | n23061 ;
  assign n23063 = n273 & ~n2924 ;
  assign n23064 = n23063 ^ n16384 ^ 1'b0 ;
  assign n23065 = n89 & ~n23064 ;
  assign n23066 = n2689 | n21836 ;
  assign n23067 = n7491 & n19017 ;
  assign n23068 = ~n1638 & n23067 ;
  assign n23069 = ~n14682 & n21763 ;
  assign n23070 = ~n418 & n17802 ;
  assign n23071 = ~n6432 & n23070 ;
  assign n23072 = n2738 ^ n1260 ^ 1'b0 ;
  assign n23073 = n1922 ^ n203 ^ 1'b0 ;
  assign n23074 = ~n8326 & n23073 ;
  assign n23075 = n10816 & ~n18403 ;
  assign n23076 = n23075 ^ n1995 ^ 1'b0 ;
  assign n23077 = n23076 ^ n3493 ^ 1'b0 ;
  assign n23078 = n3542 & ~n12371 ;
  assign n23079 = n23078 ^ n3707 ^ 1'b0 ;
  assign n23080 = n16507 | n23079 ;
  assign n23081 = n4770 | n9412 ;
  assign n23082 = n18052 ^ n3631 ^ 1'b0 ;
  assign n23083 = ~n5443 & n23082 ;
  assign n23084 = n4840 & n15090 ;
  assign n23085 = n5041 & n23084 ;
  assign n23086 = n23083 & ~n23085 ;
  assign n23087 = ~n1964 & n13255 ;
  assign n23088 = n23087 ^ n10083 ^ 1'b0 ;
  assign n23089 = n11516 ^ n5397 ^ 1'b0 ;
  assign n23090 = n23089 ^ n6907 ^ 1'b0 ;
  assign n23091 = n23088 & ~n23090 ;
  assign n23092 = n19058 ^ n14572 ^ 1'b0 ;
  assign n23093 = n7480 | n23092 ;
  assign n23094 = ~n1219 & n5725 ;
  assign n23095 = n23094 ^ n13094 ^ 1'b0 ;
  assign n23096 = n14179 & n14911 ;
  assign n23097 = n2581 ^ n255 ^ 1'b0 ;
  assign n23098 = n17282 & n23097 ;
  assign n23099 = n3152 & ~n23098 ;
  assign n23100 = n23099 ^ n15700 ^ 1'b0 ;
  assign n23101 = n12044 | n23100 ;
  assign n23102 = n23096 & ~n23101 ;
  assign n23103 = ~n532 & n23102 ;
  assign n23104 = n273 | n3837 ;
  assign n23105 = n13178 | n23104 ;
  assign n23106 = ~n4643 & n5256 ;
  assign n23107 = ~n8630 & n23106 ;
  assign n23108 = n20967 & n23107 ;
  assign n23109 = n23105 & n23108 ;
  assign n23110 = n8497 ^ n101 ^ 1'b0 ;
  assign n23111 = ~n12928 & n23110 ;
  assign n23112 = n5076 ^ n2577 ^ 1'b0 ;
  assign n23113 = n148 & n23112 ;
  assign n23114 = n1036 | n1152 ;
  assign n23115 = n2301 | n17044 ;
  assign n23116 = n23114 & ~n23115 ;
  assign n23117 = n3974 & ~n16212 ;
  assign n23118 = n3068 ^ n2615 ^ n366 ;
  assign n23119 = n9689 & ~n11775 ;
  assign n23120 = n823 & n7949 ;
  assign n23121 = n23120 ^ n17844 ^ 1'b0 ;
  assign n23123 = ~n1096 & n1293 ;
  assign n23124 = ~n1293 & n23123 ;
  assign n23125 = n6620 & ~n23124 ;
  assign n23126 = n608 | n12570 ;
  assign n23130 = ~n1622 & n2391 ;
  assign n23131 = ~n2391 & n23130 ;
  assign n23132 = ~n3270 & n9201 ;
  assign n23133 = n23131 & n23132 ;
  assign n23127 = ~n2260 & n6579 ;
  assign n23128 = n2260 & n23127 ;
  assign n23129 = ~n5376 & n23128 ;
  assign n23134 = n23133 ^ n23129 ^ 1'b0 ;
  assign n23135 = n23126 | n23134 ;
  assign n23136 = n23125 | n23135 ;
  assign n23122 = n265 & ~n3221 ;
  assign n23137 = n23136 ^ n23122 ^ 1'b0 ;
  assign n23138 = n302 | n2898 ;
  assign n23139 = n4918 & ~n23138 ;
  assign n23140 = ~n5033 & n21722 ;
  assign n23141 = n12206 & n16382 ;
  assign n23142 = ~n23140 & n23141 ;
  assign n23143 = n23139 | n23142 ;
  assign n23144 = n2240 ^ n1349 ^ 1'b0 ;
  assign n23145 = n9492 & ~n23144 ;
  assign n23146 = n5570 ^ n2484 ^ 1'b0 ;
  assign n23147 = n1655 & ~n9253 ;
  assign n23148 = n14218 ^ n450 ^ 1'b0 ;
  assign n23149 = n813 & ~n14706 ;
  assign n23150 = ~n22917 & n23149 ;
  assign n23151 = ~n3084 & n18519 ;
  assign n23152 = ~n23150 & n23151 ;
  assign n23153 = n6019 ^ n4034 ^ 1'b0 ;
  assign n23154 = ( n18125 & n21752 ) | ( n18125 & n23153 ) | ( n21752 & n23153 ) ;
  assign n23155 = ~n5156 & n23154 ;
  assign n23156 = ~n14690 & n23155 ;
  assign n23157 = n13851 & ~n19482 ;
  assign n23158 = n23157 ^ n10071 ^ 1'b0 ;
  assign n23159 = n6730 & n23158 ;
  assign n23160 = n11326 ^ n553 ^ 1'b0 ;
  assign n23161 = n6194 & n22214 ;
  assign n23162 = n673 & n23161 ;
  assign n23163 = n17250 & n23162 ;
  assign n23164 = ( ~n1880 & n14161 ) | ( ~n1880 & n14515 ) | ( n14161 & n14515 ) ;
  assign n23166 = n20472 ^ n8971 ^ 1'b0 ;
  assign n23165 = n1385 & n5179 ;
  assign n23167 = n23166 ^ n23165 ^ 1'b0 ;
  assign n23168 = n4237 & ~n15849 ;
  assign n23169 = n23168 ^ n2448 ^ 1'b0 ;
  assign n23170 = n2491 ^ n997 ^ 1'b0 ;
  assign n23171 = ~n23169 & n23170 ;
  assign n23172 = n23171 ^ n14824 ^ 1'b0 ;
  assign n23173 = n6316 & ~n23172 ;
  assign n23174 = n23167 & n23173 ;
  assign n23175 = n13470 & ~n15034 ;
  assign n23176 = n9340 & ~n13617 ;
  assign n23177 = ( n5894 & ~n17207 ) | ( n5894 & n22847 ) | ( ~n17207 & n22847 ) ;
  assign n23178 = n5700 & ~n23177 ;
  assign n23179 = n9253 ^ n581 ^ 1'b0 ;
  assign n23180 = n7626 | n21567 ;
  assign n23181 = n17815 & ~n23180 ;
  assign n23182 = n13299 ^ n10990 ^ 1'b0 ;
  assign n23183 = ~n5575 & n20682 ;
  assign n23184 = ~n4179 & n9569 ;
  assign n23185 = n5771 | n23184 ;
  assign n23186 = n23185 ^ n8097 ^ 1'b0 ;
  assign n23187 = ~n17519 & n23186 ;
  assign n23188 = n23187 ^ n18406 ^ 1'b0 ;
  assign n23189 = n20146 & ~n20850 ;
  assign n23190 = n23189 ^ n21029 ^ 1'b0 ;
  assign n23191 = n6269 & ~n15923 ;
  assign n23192 = n5525 & ~n7265 ;
  assign n23193 = ~n4334 & n23192 ;
  assign n23194 = n23193 ^ n19250 ^ 1'b0 ;
  assign n23195 = n391 & ~n7322 ;
  assign n23196 = ~n5652 & n5719 ;
  assign n23197 = n23196 ^ n8666 ^ 1'b0 ;
  assign n23198 = n3446 | n5731 ;
  assign n23199 = n14306 ^ n6923 ^ 1'b0 ;
  assign n23200 = n23198 & n23199 ;
  assign n23201 = n17190 ^ n1458 ^ 1'b0 ;
  assign n23202 = n20997 & n23201 ;
  assign n23203 = n278 & ~n4332 ;
  assign n23204 = n14731 & ~n17319 ;
  assign n23205 = ~n2946 & n23204 ;
  assign n23206 = n5557 & ~n12863 ;
  assign n23207 = n5513 ^ n3413 ^ 1'b0 ;
  assign n23208 = n23207 ^ n15925 ^ 1'b0 ;
  assign n23209 = n19367 | n23208 ;
  assign n23210 = n23209 ^ n8375 ^ n5891 ;
  assign n23211 = n4217 & ~n11021 ;
  assign n23212 = ~n6655 & n23211 ;
  assign n23213 = n21683 & n23212 ;
  assign n23214 = n15770 ^ n7806 ^ 1'b0 ;
  assign n23215 = ~n576 & n23214 ;
  assign n23216 = ~n294 & n10777 ;
  assign n23217 = n19845 | n23216 ;
  assign n23218 = n23217 ^ n634 ^ 1'b0 ;
  assign n23221 = ~n1387 & n13752 ;
  assign n23222 = n2003 & n23221 ;
  assign n23219 = n3074 & ~n15310 ;
  assign n23220 = n10262 | n23219 ;
  assign n23223 = n23222 ^ n23220 ^ 1'b0 ;
  assign n23224 = n3089 & ~n23223 ;
  assign n23225 = n8917 ^ n3231 ^ 1'b0 ;
  assign n23226 = n23225 ^ n6161 ^ 1'b0 ;
  assign n23227 = n23226 ^ n6866 ^ n6001 ;
  assign n23228 = n6305 & ~n12007 ;
  assign n23229 = n23228 ^ n5941 ^ 1'b0 ;
  assign n23230 = ~n8769 & n23229 ;
  assign n23231 = n2943 & ~n4522 ;
  assign n23232 = ~n10618 & n23231 ;
  assign n23233 = n2618 | n4499 ;
  assign n23234 = n23233 ^ n3638 ^ 1'b0 ;
  assign n23235 = n6028 ^ n1431 ^ 1'b0 ;
  assign n23236 = n19403 & n23235 ;
  assign n23241 = n7612 & ~n22371 ;
  assign n23242 = n23241 ^ n16752 ^ 1'b0 ;
  assign n23243 = n18514 | n23242 ;
  assign n23237 = ( n1768 & ~n3437 ) | ( n1768 & n16814 ) | ( ~n3437 & n16814 ) ;
  assign n23238 = n9826 ^ n8107 ^ 1'b0 ;
  assign n23239 = ~n20819 & n23238 ;
  assign n23240 = ~n23237 & n23239 ;
  assign n23244 = n23243 ^ n23240 ^ 1'b0 ;
  assign n23245 = x1 & ~n2991 ;
  assign n23246 = n2148 & n23245 ;
  assign n23247 = ( n2043 & n8173 ) | ( n2043 & ~n23246 ) | ( n8173 & ~n23246 ) ;
  assign n23248 = ~n1492 & n8974 ;
  assign n23249 = n15602 & n23248 ;
  assign n23250 = n23249 ^ n142 ^ 1'b0 ;
  assign n23251 = n23247 & ~n23250 ;
  assign n23252 = n16144 & n23251 ;
  assign n23253 = n17517 ^ n3267 ^ n1768 ;
  assign n23254 = n23253 ^ n10347 ^ 1'b0 ;
  assign n23255 = n184 & n1463 ;
  assign n23256 = n9718 & n23255 ;
  assign n23257 = n7353 ^ n1560 ^ 1'b0 ;
  assign n23258 = n23256 | n23257 ;
  assign n23259 = n23258 ^ n16636 ^ 1'b0 ;
  assign n23260 = n12867 | n18853 ;
  assign n23261 = n16510 & ~n23260 ;
  assign n23262 = n5205 ^ n2751 ^ 1'b0 ;
  assign n23263 = n8519 ^ n1318 ^ 1'b0 ;
  assign n23264 = n23262 | n23263 ;
  assign n23265 = n23264 ^ n3394 ^ 1'b0 ;
  assign n23266 = n23261 | n23265 ;
  assign n23267 = ~n2318 & n8854 ;
  assign n23268 = ~n9192 & n23267 ;
  assign n23269 = n21219 & n23268 ;
  assign n23270 = n415 & ~n23269 ;
  assign n23271 = n23270 ^ n18977 ^ 1'b0 ;
  assign n23272 = n715 | n6488 ;
  assign n23273 = n23272 ^ n3392 ^ 1'b0 ;
  assign n23274 = n8319 ^ n4419 ^ 1'b0 ;
  assign n23275 = n177 | n18282 ;
  assign n23276 = n5554 | n23275 ;
  assign n23277 = n23274 & n23276 ;
  assign n23278 = n630 & ~n9333 ;
  assign n23279 = ( n3219 & ~n16184 ) | ( n3219 & n19954 ) | ( ~n16184 & n19954 ) ;
  assign n23280 = n23279 ^ n3919 ^ n962 ;
  assign n23282 = n4850 & n5428 ;
  assign n23281 = n9636 & n13918 ;
  assign n23283 = n23282 ^ n23281 ^ 1'b0 ;
  assign n23284 = n1918 ^ n1688 ^ 1'b0 ;
  assign n23285 = n4799 & n23284 ;
  assign n23286 = n2044 | n2494 ;
  assign n23287 = n23285 | n23286 ;
  assign n23288 = n5053 ^ n2339 ^ 1'b0 ;
  assign n23289 = n4924 & n5402 ;
  assign n23290 = ~n13992 & n23289 ;
  assign n23291 = ~n23288 & n23290 ;
  assign n23292 = n18477 & n23291 ;
  assign n23293 = ~n23287 & n23292 ;
  assign n23295 = ( ~n9379 & n11229 ) | ( ~n9379 & n11631 ) | ( n11229 & n11631 ) ;
  assign n23294 = ~n17946 & n20284 ;
  assign n23296 = n23295 ^ n23294 ^ 1'b0 ;
  assign n23297 = n8257 & ~n16827 ;
  assign n23299 = n1739 | n2485 ;
  assign n23300 = n23299 ^ n6197 ^ n149 ;
  assign n23301 = ~n190 & n6418 ;
  assign n23302 = ~n23300 & n23301 ;
  assign n23303 = n1701 ^ n16 ^ 1'b0 ;
  assign n23304 = ~n23302 & n23303 ;
  assign n23305 = n23304 ^ n753 ^ 1'b0 ;
  assign n23306 = n8081 & ~n23305 ;
  assign n23298 = n6725 & ~n10533 ;
  assign n23307 = n23306 ^ n23298 ^ 1'b0 ;
  assign n23308 = n23307 ^ n14341 ^ 1'b0 ;
  assign n23309 = n5802 & ~n23308 ;
  assign n23310 = n9141 & ~n13411 ;
  assign n23311 = n1950 | n2273 ;
  assign n23312 = n23311 ^ n532 ^ 1'b0 ;
  assign n23313 = n15650 & n23312 ;
  assign n23314 = n12889 | n14440 ;
  assign n23316 = n8362 | n14930 ;
  assign n23315 = n325 | n11239 ;
  assign n23317 = n23316 ^ n23315 ^ 1'b0 ;
  assign n23318 = n4241 & n6079 ;
  assign n23319 = n23318 ^ n1098 ^ 1'b0 ;
  assign n23320 = n2810 & n13384 ;
  assign n23321 = n7114 ^ n6628 ^ 1'b0 ;
  assign n23322 = n23321 ^ n5922 ^ 1'b0 ;
  assign n23323 = n23322 ^ n11080 ^ 1'b0 ;
  assign n23324 = n23320 & ~n23323 ;
  assign n23325 = n23319 & ~n23324 ;
  assign n23326 = n10794 ^ n4840 ^ 1'b0 ;
  assign n23327 = n23326 ^ n17169 ^ n10242 ;
  assign n23328 = n53 | n12079 ;
  assign n23329 = n22602 | n23328 ;
  assign n23330 = n23329 ^ n3368 ^ 1'b0 ;
  assign n23331 = ~n13132 & n23330 ;
  assign n23332 = ~n7956 & n23331 ;
  assign n23336 = ~n241 & n1663 ;
  assign n23337 = n23336 ^ n3929 ^ 1'b0 ;
  assign n23333 = n388 & n541 ;
  assign n23334 = n23333 ^ n4936 ^ 1'b0 ;
  assign n23335 = n5561 | n23334 ;
  assign n23338 = n23337 ^ n23335 ^ 1'b0 ;
  assign n23339 = n323 & ~n5713 ;
  assign n23340 = n23339 ^ n830 ^ 1'b0 ;
  assign n23341 = n12095 & ~n23340 ;
  assign n23342 = n20254 ^ n2324 ^ 1'b0 ;
  assign n23343 = n128 | n21986 ;
  assign n23344 = n11564 | n21561 ;
  assign n23345 = n23344 ^ n2870 ^ 1'b0 ;
  assign n23346 = n3256 | n6280 ;
  assign n23347 = n5956 ^ n592 ^ 1'b0 ;
  assign n23348 = n2173 & n2910 ;
  assign n23349 = n23348 ^ n4480 ^ 1'b0 ;
  assign n23350 = n23347 | n23349 ;
  assign n23351 = n52 & n4714 ;
  assign n23352 = ~n744 & n5030 ;
  assign n23353 = n8116 ^ n7605 ^ 1'b0 ;
  assign n23354 = n1174 & n16759 ;
  assign n23355 = n7512 | n19096 ;
  assign n23356 = n228 | n8860 ;
  assign n23357 = n7231 | n9302 ;
  assign n23358 = n23357 ^ n8624 ^ 1'b0 ;
  assign n23359 = n581 | n1112 ;
  assign n23360 = n581 & ~n23359 ;
  assign n23361 = ~n6321 & n23360 ;
  assign n23362 = n12895 & n23361 ;
  assign n23366 = n297 & n860 ;
  assign n23367 = ~n860 & n23366 ;
  assign n23363 = n3479 & ~n4992 ;
  assign n23364 = n4992 & n23363 ;
  assign n23365 = n5538 | n23364 ;
  assign n23368 = n23367 ^ n23365 ^ 1'b0 ;
  assign n23369 = n23368 ^ n19009 ^ 1'b0 ;
  assign n23370 = n23362 & n23369 ;
  assign n23371 = n709 & ~n23370 ;
  assign n23372 = n177 & n14112 ;
  assign n23373 = n23372 ^ n15108 ^ 1'b0 ;
  assign n23374 = n5187 | n21029 ;
  assign n23375 = n5083 & ~n23374 ;
  assign n23376 = n7107 ^ n3946 ^ 1'b0 ;
  assign n23377 = n16559 & n23376 ;
  assign n23378 = n9588 ^ n1235 ^ 1'b0 ;
  assign n23379 = n16652 & n23378 ;
  assign n23380 = n23379 ^ n1255 ^ 1'b0 ;
  assign n23381 = n9149 ^ n3765 ^ 1'b0 ;
  assign n23382 = n15021 & ~n23275 ;
  assign n23383 = ~n15137 & n23382 ;
  assign n23384 = n23381 & n23383 ;
  assign n23385 = n14713 | n23384 ;
  assign n23386 = n12289 & ~n23020 ;
  assign n23387 = n8418 ^ n128 ^ 1'b0 ;
  assign n23388 = n8562 | n23387 ;
  assign n23389 = n4749 ^ n2833 ^ 1'b0 ;
  assign n23390 = n20023 & n23389 ;
  assign n23391 = ~n8347 & n23199 ;
  assign n23392 = n23390 & n23391 ;
  assign n23398 = n6281 & n14513 ;
  assign n23393 = n4381 | n23144 ;
  assign n23394 = n23393 ^ n18205 ^ 1'b0 ;
  assign n23395 = n3115 ^ n851 ^ 1'b0 ;
  assign n23396 = n23394 | n23395 ;
  assign n23397 = n23396 ^ n15707 ^ 1'b0 ;
  assign n23399 = n23398 ^ n23397 ^ 1'b0 ;
  assign n23400 = n18390 ^ n339 ^ 1'b0 ;
  assign n23401 = n1372 ^ n423 ^ 1'b0 ;
  assign n23402 = n5660 | n23401 ;
  assign n23404 = n3434 ^ n161 ^ 1'b0 ;
  assign n23405 = ~n938 & n23404 ;
  assign n23406 = n4446 & n23405 ;
  assign n23407 = n23406 ^ n4666 ^ 1'b0 ;
  assign n23403 = ~n5317 & n19765 ;
  assign n23408 = n23407 ^ n23403 ^ 1'b0 ;
  assign n23409 = n3718 ^ n2408 ^ 1'b0 ;
  assign n23410 = n6552 & n23409 ;
  assign n23411 = ~n6419 & n11656 ;
  assign n23412 = ~n14055 & n23411 ;
  assign n23413 = n23412 ^ n4332 ^ 1'b0 ;
  assign n23414 = n3559 & n23413 ;
  assign n23415 = n6025 ^ n4037 ^ 1'b0 ;
  assign n23416 = n23414 & n23415 ;
  assign n23417 = ~n5527 & n6441 ;
  assign n23418 = n23417 ^ n17796 ^ 1'b0 ;
  assign n23419 = n2542 & n18798 ;
  assign n23420 = ~n678 & n16913 ;
  assign n23421 = n23420 ^ n6197 ^ 1'b0 ;
  assign n23422 = n273 & ~n419 ;
  assign n23423 = n419 & n23422 ;
  assign n23424 = n23423 ^ n158 ^ 1'b0 ;
  assign n23425 = n8337 | n23424 ;
  assign n23426 = n79 & n7171 ;
  assign n23427 = ~n273 & n23426 ;
  assign n23428 = ~n157 & n23427 ;
  assign n23429 = n2011 | n23428 ;
  assign n23430 = n2011 & ~n23429 ;
  assign n23431 = n6745 & ~n13496 ;
  assign n23432 = n13496 & n23431 ;
  assign n23433 = n23430 & ~n23432 ;
  assign n23434 = n23425 | n23433 ;
  assign n23435 = n23425 & ~n23434 ;
  assign n23436 = n16499 & ~n18472 ;
  assign n23437 = n23435 & n23436 ;
  assign n23438 = n1893 & ~n16940 ;
  assign n23439 = n6025 | n7647 ;
  assign n23440 = n2494 | n23439 ;
  assign n23441 = n10086 ^ n8972 ^ 1'b0 ;
  assign n23442 = ~n23440 & n23441 ;
  assign n23443 = n23442 ^ n3744 ^ 1'b0 ;
  assign n23444 = n23438 & ~n23443 ;
  assign n23445 = n5811 & n18995 ;
  assign n23446 = n23445 ^ n3990 ^ 1'b0 ;
  assign n23447 = ~n3793 & n15126 ;
  assign n23448 = ~n169 & n1125 ;
  assign n23449 = n983 & n23448 ;
  assign n23450 = n8097 | n23449 ;
  assign n23451 = n3447 ^ n2273 ^ n1198 ;
  assign n23452 = ~n15986 & n19495 ;
  assign n23453 = n3049 & n23452 ;
  assign n23454 = ~n23451 & n23453 ;
  assign n23455 = n2007 ^ n378 ^ 1'b0 ;
  assign n23456 = n12689 & ~n13299 ;
  assign n23457 = n18494 | n19721 ;
  assign n23458 = n23457 ^ n3524 ^ 1'b0 ;
  assign n23459 = ~n23456 & n23458 ;
  assign n23460 = n592 | n5914 ;
  assign n23461 = n23460 ^ x5 ^ 1'b0 ;
  assign n23462 = n14699 ^ n1537 ^ 1'b0 ;
  assign n23463 = n16284 & ~n23462 ;
  assign n23464 = n82 | n5513 ;
  assign n23465 = n258 & n21300 ;
  assign n23466 = ~n19148 & n23465 ;
  assign n23467 = ~n130 & n4349 ;
  assign n23468 = ~n8092 & n23467 ;
  assign n23469 = n6295 & n15429 ;
  assign n23470 = n23469 ^ n10519 ^ 1'b0 ;
  assign n23471 = n23470 ^ n14235 ^ 1'b0 ;
  assign n23472 = n2038 | n23471 ;
  assign n23473 = ~n5891 & n19761 ;
  assign n23474 = n18562 & n23473 ;
  assign n23475 = n5227 & n23474 ;
  assign n23476 = n5193 & ~n19544 ;
  assign n23477 = n169 & n23476 ;
  assign n23478 = n17683 ^ n1927 ^ 1'b0 ;
  assign n23479 = n2969 & n5275 ;
  assign n23480 = n322 | n23479 ;
  assign n23481 = n20541 | n21994 ;
  assign n23482 = n11266 & ~n23481 ;
  assign n23483 = n4033 ^ n1959 ^ 1'b0 ;
  assign n23485 = n8510 & n10383 ;
  assign n23484 = n2348 ^ n1015 ^ 1'b0 ;
  assign n23486 = n23485 ^ n23484 ^ 1'b0 ;
  assign n23487 = n23486 ^ n5253 ^ 1'b0 ;
  assign n23488 = ~n23483 & n23487 ;
  assign n23489 = ~n15023 & n22640 ;
  assign n23490 = n23489 ^ n22496 ^ 1'b0 ;
  assign n23491 = ( n7855 & n17599 ) | ( n7855 & n22987 ) | ( n17599 & n22987 ) ;
  assign n23492 = n6946 ^ n113 ^ 1'b0 ;
  assign n23493 = ~n15229 & n23492 ;
  assign n23496 = n1900 & n2594 ;
  assign n23494 = n11820 | n19583 ;
  assign n23495 = n23494 ^ n6766 ^ 1'b0 ;
  assign n23497 = n23496 ^ n23495 ^ 1'b0 ;
  assign n23498 = n17860 & n23497 ;
  assign n23499 = n6611 ^ n356 ^ 1'b0 ;
  assign n23500 = n400 | n23499 ;
  assign n23501 = ( n3801 & n12046 ) | ( n3801 & n16759 ) | ( n12046 & n16759 ) ;
  assign n23502 = n23500 | n23501 ;
  assign n23503 = n210 | n410 ;
  assign n23504 = n122 & ~n23503 ;
  assign n23505 = ( n18896 & n19212 ) | ( n18896 & ~n23504 ) | ( n19212 & ~n23504 ) ;
  assign n23507 = ~n1073 & n2418 ;
  assign n23508 = ~n23320 & n23507 ;
  assign n23506 = n734 ^ n436 ^ 1'b0 ;
  assign n23509 = n23508 ^ n23506 ^ 1'b0 ;
  assign n23510 = n23505 & n23509 ;
  assign n23511 = n907 | n21229 ;
  assign n23512 = n23511 ^ n7994 ^ 1'b0 ;
  assign n23513 = n5950 | n14678 ;
  assign n23514 = n23513 ^ n973 ^ 1'b0 ;
  assign n23515 = n4473 & ~n6033 ;
  assign n23516 = n9236 ^ n6656 ^ 1'b0 ;
  assign n23517 = n2714 & ~n21717 ;
  assign n23518 = ~n3223 & n5025 ;
  assign n23519 = n23518 ^ n23247 ^ 1'b0 ;
  assign n23520 = n4904 & n12060 ;
  assign n23521 = n23520 ^ n13573 ^ 1'b0 ;
  assign n23522 = n8266 & n12689 ;
  assign n23523 = ~n662 & n10052 ;
  assign n23524 = n398 & n23523 ;
  assign n23525 = ~n857 & n23524 ;
  assign n23526 = n10317 ^ x9 ^ 1'b0 ;
  assign n23527 = n4616 | n23526 ;
  assign n23528 = n23527 ^ n128 ^ 1'b0 ;
  assign n23529 = ~n954 & n14218 ;
  assign n23530 = n4574 & n23529 ;
  assign n23531 = ~n5749 & n13827 ;
  assign n23532 = n23531 ^ n7032 ^ 1'b0 ;
  assign n23533 = n8568 & ~n23532 ;
  assign n23534 = n5584 & n6061 ;
  assign n23535 = n23534 ^ n3983 ^ 1'b0 ;
  assign n23536 = n5956 & ~n23535 ;
  assign n23537 = n932 | n2291 ;
  assign n23538 = n11963 | n23537 ;
  assign n23539 = n800 & ~n23538 ;
  assign n23540 = n2303 ^ n1637 ^ 1'b0 ;
  assign n23541 = n8479 | n9111 ;
  assign n23542 = n10262 & ~n23541 ;
  assign n23543 = ~n15864 & n22674 ;
  assign n23544 = n10338 ^ n339 ^ 1'b0 ;
  assign n23545 = n2238 & ~n3030 ;
  assign n23546 = ~n1852 & n23545 ;
  assign n23547 = n23546 ^ n11272 ^ 1'b0 ;
  assign n23548 = n23544 & n23547 ;
  assign n23549 = n3724 ^ n1465 ^ 1'b0 ;
  assign n23550 = n4812 & n23549 ;
  assign n23551 = n23550 ^ n2141 ^ 1'b0 ;
  assign n23552 = n6862 | n9441 ;
  assign n23553 = n5419 | n23552 ;
  assign n23554 = ~n2843 & n9213 ;
  assign n23555 = n23554 ^ n23379 ^ 1'b0 ;
  assign n23556 = n11618 | n15655 ;
  assign n23557 = n12457 & ~n23556 ;
  assign n23558 = n6546 & ~n23557 ;
  assign n23559 = n415 | n15173 ;
  assign n23560 = n23559 ^ n984 ^ 1'b0 ;
  assign n23561 = n11412 ^ n8688 ^ 1'b0 ;
  assign n23562 = ~n599 & n23561 ;
  assign n23563 = n12482 ^ n6558 ^ 1'b0 ;
  assign n23564 = ~n7657 & n23563 ;
  assign n23565 = n23564 ^ n10216 ^ 1'b0 ;
  assign n23566 = n23562 & n23565 ;
  assign n23567 = ~n1352 & n8939 ;
  assign n23568 = ~n2199 & n13364 ;
  assign n23569 = n13709 ^ n8827 ^ 1'b0 ;
  assign n23570 = n23569 ^ n13981 ^ n9004 ;
  assign n23571 = n9364 | n23570 ;
  assign n23576 = n10926 ^ n1600 ^ 1'b0 ;
  assign n23572 = n8258 & ~n11487 ;
  assign n23573 = n10966 & n23572 ;
  assign n23574 = n23038 ^ n236 ^ 1'b0 ;
  assign n23575 = ~n23573 & n23574 ;
  assign n23577 = n23576 ^ n23575 ^ n8149 ;
  assign n23578 = n1154 | n5629 ;
  assign n23579 = n23578 ^ n4996 ^ 1'b0 ;
  assign n23580 = n19688 ^ n4646 ^ n232 ;
  assign n23581 = n884 & ~n1416 ;
  assign n23582 = n23581 ^ n3348 ^ 1'b0 ;
  assign n23583 = ~n23580 & n23582 ;
  assign n23584 = n532 ^ n80 ^ 1'b0 ;
  assign n23585 = n1008 | n23584 ;
  assign n23586 = n4114 | n23585 ;
  assign n23587 = n6330 | n23586 ;
  assign n23588 = n23587 ^ n23583 ^ 1'b0 ;
  assign n23589 = n23583 | n23588 ;
  assign n23590 = n6011 & n23589 ;
  assign n23591 = n23590 ^ n12407 ^ 1'b0 ;
  assign n23592 = n962 ^ n142 ^ 1'b0 ;
  assign n23593 = n23592 ^ n9281 ^ 1'b0 ;
  assign n23594 = n12094 | n23593 ;
  assign n23595 = n16659 & ~n23594 ;
  assign n23596 = ( ~n3634 & n18137 ) | ( ~n3634 & n23595 ) | ( n18137 & n23595 ) ;
  assign n23597 = n23596 ^ n7227 ^ n3593 ;
  assign n23598 = n7424 | n23401 ;
  assign n23599 = n7700 | n23598 ;
  assign n23600 = ~n11360 & n23599 ;
  assign n23601 = n8823 ^ n2572 ^ 1'b0 ;
  assign n23602 = n2942 & n10507 ;
  assign n23603 = n23602 ^ n7181 ^ 1'b0 ;
  assign n23604 = n23601 & ~n23603 ;
  assign n23605 = ( n1529 & n8053 ) | ( n1529 & ~n16660 ) | ( n8053 & ~n16660 ) ;
  assign n23606 = n23605 ^ n2535 ^ 1'b0 ;
  assign n23607 = x4 & n23606 ;
  assign n23610 = ~n9322 & n15159 ;
  assign n23611 = n332 & n23610 ;
  assign n23608 = n1814 & ~n6230 ;
  assign n23609 = ~n4449 & n23608 ;
  assign n23612 = n23611 ^ n23609 ^ 1'b0 ;
  assign n23613 = n8291 ^ n294 ^ 1'b0 ;
  assign n23614 = ~n23612 & n23613 ;
  assign n23616 = n16983 ^ n954 ^ 1'b0 ;
  assign n23615 = n4446 & ~n10660 ;
  assign n23617 = n23616 ^ n23615 ^ 1'b0 ;
  assign n23618 = n1673 | n23195 ;
  assign n23619 = n22371 ^ n6178 ^ 1'b0 ;
  assign n23620 = n12777 & ~n23619 ;
  assign n23621 = ~n10543 & n23620 ;
  assign n23622 = n23621 ^ n1579 ^ 1'b0 ;
  assign n23623 = n1960 & n2351 ;
  assign n23624 = ~n4818 & n23623 ;
  assign n23625 = n18029 ^ n15931 ^ 1'b0 ;
  assign n23626 = n6647 & ~n23625 ;
  assign n23627 = ~n23624 & n23626 ;
  assign n23628 = n23627 ^ n10886 ^ 1'b0 ;
  assign n23629 = ( n3003 & ~n10429 ) | ( n3003 & n11508 ) | ( ~n10429 & n11508 ) ;
  assign n23630 = n12381 ^ n3990 ^ 1'b0 ;
  assign n23631 = n15009 | n23630 ;
  assign n23632 = n11768 ^ n5632 ^ 1'b0 ;
  assign n23633 = n4840 | n23632 ;
  assign n23634 = n5771 | n23633 ;
  assign n23635 = n14114 | n23634 ;
  assign n23636 = n5024 & ~n8109 ;
  assign n23637 = n23636 ^ n18522 ^ 1'b0 ;
  assign n23638 = n958 & n10852 ;
  assign n23639 = n23638 ^ n7135 ^ 1'b0 ;
  assign n23640 = ~n3663 & n9723 ;
  assign n23641 = n23640 ^ n4757 ^ 1'b0 ;
  assign n23642 = n8850 ^ n2020 ^ 1'b0 ;
  assign n23643 = n958 & ~n17845 ;
  assign n23644 = ~n23642 & n23643 ;
  assign n23645 = n23641 & ~n23644 ;
  assign n23646 = n13821 ^ n12898 ^ 1'b0 ;
  assign n23647 = ~n5135 & n23646 ;
  assign n23648 = ~n3782 & n15987 ;
  assign n23649 = ~n21785 & n23648 ;
  assign n23650 = n13108 ^ n7690 ^ 1'b0 ;
  assign n23651 = n281 & ~n1026 ;
  assign n23652 = n963 & n23651 ;
  assign n23653 = n23652 ^ n12968 ^ 1'b0 ;
  assign n23654 = n7316 | n10511 ;
  assign n23655 = n10428 & n23654 ;
  assign n23656 = n1520 & ~n3116 ;
  assign n23657 = ~n1520 & n23656 ;
  assign n23658 = n15727 & ~n23657 ;
  assign n23661 = ~n308 & n659 ;
  assign n23662 = n308 & n23661 ;
  assign n23659 = ~n55 & n484 ;
  assign n23660 = n55 & n23659 ;
  assign n23663 = n23662 ^ n23660 ^ 1'b0 ;
  assign n23664 = n23658 & n23663 ;
  assign n23665 = n1441 & n23664 ;
  assign n23666 = ~n963 & n23665 ;
  assign n23667 = n23666 ^ n367 ^ 1'b0 ;
  assign n23668 = n1766 | n3743 ;
  assign n23669 = n1766 & ~n23668 ;
  assign n23670 = n596 & ~n8279 ;
  assign n23671 = n23669 & n23670 ;
  assign n23672 = ~n4947 & n23671 ;
  assign n23673 = n23672 ^ n5792 ^ 1'b0 ;
  assign n23674 = n23667 | n23673 ;
  assign n23675 = n12441 & n16906 ;
  assign n23676 = n23675 ^ n13462 ^ 1'b0 ;
  assign n23677 = n4856 ^ n1315 ^ 1'b0 ;
  assign n23678 = n23677 ^ n6922 ^ 1'b0 ;
  assign n23679 = n20787 & ~n23678 ;
  assign n23680 = n1956 | n17668 ;
  assign n23681 = n2582 & ~n23680 ;
  assign n23682 = n81 & ~n9718 ;
  assign n23683 = n23681 & n23682 ;
  assign n23684 = n7900 ^ n249 ^ 1'b0 ;
  assign n23685 = ( n94 & n1637 ) | ( n94 & n3598 ) | ( n1637 & n3598 ) ;
  assign n23686 = n23684 | n23685 ;
  assign n23687 = n5467 ^ n246 ^ 1'b0 ;
  assign n23688 = n330 & n18191 ;
  assign n23689 = n23688 ^ n13798 ^ 1'b0 ;
  assign n23690 = n14152 & ~n23689 ;
  assign n23691 = ( n6246 & ~n21586 ) | ( n6246 & n23690 ) | ( ~n21586 & n23690 ) ;
  assign n23692 = n18643 & n21624 ;
  assign n23693 = n596 & ~n2546 ;
  assign n23694 = n23693 ^ n15312 ^ 1'b0 ;
  assign n23695 = n19490 ^ n533 ^ 1'b0 ;
  assign n23696 = ~n9009 & n18021 ;
  assign n23697 = n3634 & ~n3710 ;
  assign n23698 = n14142 | n23697 ;
  assign n23699 = n4998 & n23698 ;
  assign n23700 = n2189 & n11322 ;
  assign n23701 = n565 | n6894 ;
  assign n23702 = n12225 | n23701 ;
  assign n23705 = n1477 & n3572 ;
  assign n23706 = n2217 & n23705 ;
  assign n23703 = n16302 & ~n21398 ;
  assign n23704 = n2074 & n23703 ;
  assign n23707 = n23706 ^ n23704 ^ 1'b0 ;
  assign n23708 = n6758 | n11532 ;
  assign n23709 = n11532 & ~n23708 ;
  assign n23710 = ~n6428 & n23709 ;
  assign n23711 = n512 & ~n748 ;
  assign n23712 = n23711 ^ n853 ^ 1'b0 ;
  assign n23715 = n1477 & n1790 ;
  assign n23716 = ~n1302 & n23715 ;
  assign n23717 = n782 | n23716 ;
  assign n23718 = n178 | n23717 ;
  assign n23719 = ~n1714 & n12453 ;
  assign n23720 = ~n23718 & n23719 ;
  assign n23721 = n23720 ^ n555 ^ 1'b0 ;
  assign n23713 = ~n128 & n1683 ;
  assign n23714 = n2932 | n23713 ;
  assign n23722 = n23721 ^ n23714 ^ 1'b0 ;
  assign n23723 = ~n23712 & n23722 ;
  assign n23724 = n23723 ^ n18847 ^ 1'b0 ;
  assign n23725 = n8415 ^ n5041 ^ 1'b0 ;
  assign n23726 = n20322 & n23725 ;
  assign n23727 = n2168 & ~n17246 ;
  assign n23728 = n23727 ^ n21199 ^ n2951 ;
  assign n23729 = n13538 | n13748 ;
  assign n23730 = n10973 ^ n9137 ^ 1'b0 ;
  assign n23731 = n7006 | n7676 ;
  assign n23732 = n6602 | n23731 ;
  assign n23733 = ~n4724 & n13487 ;
  assign n23734 = n23733 ^ n13056 ^ 1'b0 ;
  assign n23735 = n23734 ^ n4294 ^ 1'b0 ;
  assign n23736 = ~n23732 & n23735 ;
  assign n23737 = n5075 | n5856 ;
  assign n23738 = n18099 | n23737 ;
  assign n23739 = n23738 ^ n252 ^ 1'b0 ;
  assign n23740 = n23739 ^ n2836 ^ 1'b0 ;
  assign n23741 = n9592 & n13607 ;
  assign n23742 = n1246 & ~n4273 ;
  assign n23743 = ( n4897 & n18807 ) | ( n4897 & n20010 ) | ( n18807 & n20010 ) ;
  assign n23744 = ~n14844 & n23743 ;
  assign n23745 = n6587 & n23744 ;
  assign n23746 = ~n2848 & n7038 ;
  assign n23747 = ~n812 & n23746 ;
  assign n23748 = ~n2665 & n23747 ;
  assign n23749 = ~n14159 & n23748 ;
  assign n23750 = n16294 ^ n8377 ^ n5617 ;
  assign n23751 = n19760 & n23750 ;
  assign n23752 = n1851 | n14174 ;
  assign n23753 = ~n14106 & n15124 ;
  assign n23754 = n23753 ^ n3685 ^ 1'b0 ;
  assign n23755 = n14824 & n15866 ;
  assign n23756 = ~n11848 & n18266 ;
  assign n23757 = n19948 & n23756 ;
  assign n23758 = n3368 & ~n23246 ;
  assign n23759 = n8590 ^ n2662 ^ 1'b0 ;
  assign n23760 = n3475 & n23759 ;
  assign n23761 = ~n8427 & n23760 ;
  assign n23764 = n15725 ^ n4836 ^ 1'b0 ;
  assign n23762 = n241 & ~n15108 ;
  assign n23763 = ~n2117 & n23762 ;
  assign n23765 = n23764 ^ n23763 ^ 1'b0 ;
  assign n23766 = n10030 & n11981 ;
  assign n23767 = n1704 & n23766 ;
  assign n23768 = n23767 ^ n11436 ^ 1'b0 ;
  assign n23769 = n14550 ^ n5416 ^ 1'b0 ;
  assign n23770 = n156 & n7114 ;
  assign n23771 = n23770 ^ n5758 ^ 1'b0 ;
  assign n23772 = n5186 ^ n996 ^ 1'b0 ;
  assign n23773 = ~n758 & n23772 ;
  assign n23774 = n23771 | n23773 ;
  assign n23775 = n205 & n8767 ;
  assign n23776 = n23775 ^ n15060 ^ 1'b0 ;
  assign n23777 = n19744 | n23776 ;
  assign n23778 = n23777 ^ n5856 ^ 1'b0 ;
  assign n23779 = ~n6129 & n14326 ;
  assign n23780 = ~n1155 & n23779 ;
  assign n23781 = n23780 ^ n7006 ^ 1'b0 ;
  assign n23782 = n14075 ^ n2260 ^ 1'b0 ;
  assign n23783 = n4353 & n23782 ;
  assign n23784 = n2209 & n23783 ;
  assign n23785 = n20128 & ~n23784 ;
  assign n23786 = n19518 ^ n1245 ^ 1'b0 ;
  assign n23787 = n5439 & n22487 ;
  assign n23788 = n23787 ^ n6901 ^ 1'b0 ;
  assign n23789 = n19641 ^ n4750 ^ 1'b0 ;
  assign n23790 = n15485 & ~n23789 ;
  assign n23791 = n4283 & n13627 ;
  assign n23792 = ~n1100 & n23791 ;
  assign n23793 = n9635 & ~n10001 ;
  assign n23794 = ~n3175 & n23793 ;
  assign n23795 = n23794 ^ n366 ^ 1'b0 ;
  assign n23796 = ~n3352 & n6719 ;
  assign n23797 = n23795 & ~n23796 ;
  assign n23801 = n638 & ~n5423 ;
  assign n23802 = ~n4862 & n23801 ;
  assign n23800 = n292 | n1802 ;
  assign n23803 = n23802 ^ n23800 ^ 1'b0 ;
  assign n23798 = n7063 & n22843 ;
  assign n23799 = n23798 ^ n6458 ^ 1'b0 ;
  assign n23804 = n23803 ^ n23799 ^ 1'b0 ;
  assign n23805 = n11493 ^ n3078 ^ 1'b0 ;
  assign n23806 = n5278 | n23805 ;
  assign n23807 = n23806 ^ n11514 ^ 1'b0 ;
  assign n23808 = n9472 & ~n13142 ;
  assign n23809 = ~n9472 & n23808 ;
  assign n23810 = n582 & n23809 ;
  assign n23811 = n907 & n23810 ;
  assign n23812 = ~n22175 & n23811 ;
  assign n23813 = n22175 & n23812 ;
  assign n23814 = n13956 ^ n9434 ^ 1'b0 ;
  assign n23815 = ( ~n2022 & n7285 ) | ( ~n2022 & n8685 ) | ( n7285 & n8685 ) ;
  assign n23816 = n13091 ^ n3318 ^ n1052 ;
  assign n23817 = n18811 & n23816 ;
  assign n23818 = n246 | n8130 ;
  assign n23819 = n799 | n23818 ;
  assign n23820 = n1326 & n3589 ;
  assign n23821 = ~n1370 & n23820 ;
  assign n23822 = n23819 | n23821 ;
  assign n23823 = n2176 & ~n5981 ;
  assign n23824 = ~n258 & n23823 ;
  assign n23825 = n7824 | n23824 ;
  assign n23826 = n2380 | n23825 ;
  assign n23827 = n2549 ^ n1644 ^ 1'b0 ;
  assign n23828 = n310 & n23827 ;
  assign n23829 = n7619 ^ n1653 ^ 1'b0 ;
  assign n23830 = n10499 | n15674 ;
  assign n23831 = n23829 & ~n23830 ;
  assign n23832 = ~n14337 & n20420 ;
  assign n23833 = n23832 ^ n12341 ^ 1'b0 ;
  assign n23834 = ~n2964 & n7033 ;
  assign n23835 = ~n16136 & n23834 ;
  assign n23836 = n5760 & n6225 ;
  assign n23837 = n23836 ^ n9292 ^ 1'b0 ;
  assign n23838 = n23837 ^ n3187 ^ n2011 ;
  assign n23839 = n10858 | n16745 ;
  assign n23840 = n7126 ^ n2068 ^ 1'b0 ;
  assign n23841 = n12738 & ~n23840 ;
  assign n23842 = n2797 & ~n14955 ;
  assign n23843 = n4830 | n7870 ;
  assign n23844 = n2087 ^ n1029 ^ 1'b0 ;
  assign n23845 = n23843 | n23844 ;
  assign n23846 = n23845 ^ n5187 ^ 1'b0 ;
  assign n23847 = n7673 ^ n6904 ^ 1'b0 ;
  assign n23848 = n148 | n9834 ;
  assign n23849 = n23848 ^ n13892 ^ 1'b0 ;
  assign n23850 = n13462 ^ n5005 ^ 1'b0 ;
  assign n23851 = ~n3890 & n23850 ;
  assign n23852 = n14422 & n23496 ;
  assign n23853 = n9998 & ~n19653 ;
  assign n23854 = n23853 ^ n6226 ^ 1'b0 ;
  assign n23855 = n1960 & n8614 ;
  assign n23856 = n23855 ^ n17845 ^ n79 ;
  assign n23857 = n7466 | n23856 ;
  assign n23858 = n1642 & ~n17125 ;
  assign n23859 = n23858 ^ n3146 ^ 1'b0 ;
  assign n23860 = ~n1058 & n7153 ;
  assign n23861 = n7029 & n18807 ;
  assign n23862 = n892 & ~n5223 ;
  assign n23863 = n12552 | n23862 ;
  assign n23864 = n3392 & n9053 ;
  assign n23865 = n4049 & n13913 ;
  assign n23866 = n3101 & n3567 ;
  assign n23867 = ~n23865 & n23866 ;
  assign n23868 = n3240 & n23239 ;
  assign n23869 = n5295 & n18592 ;
  assign n23870 = n6989 & n15495 ;
  assign n23871 = ( ~n8139 & n17189 ) | ( ~n8139 & n21423 ) | ( n17189 & n21423 ) ;
  assign n23873 = n10488 ^ n6519 ^ 1'b0 ;
  assign n23874 = n6476 & ~n23873 ;
  assign n23872 = n5980 ^ n1022 ^ 1'b0 ;
  assign n23875 = n23874 ^ n23872 ^ 1'b0 ;
  assign n23876 = n23875 ^ n695 ^ 1'b0 ;
  assign n23877 = n960 | n1528 ;
  assign n23878 = n23877 ^ n3928 ^ 1'b0 ;
  assign n23881 = n2286 & ~n11882 ;
  assign n23879 = n378 & ~n9613 ;
  assign n23880 = n2477 | n23879 ;
  assign n23882 = n23881 ^ n23880 ^ 1'b0 ;
  assign n23883 = n22874 & n23882 ;
  assign n23884 = n23883 ^ n19950 ^ 1'b0 ;
  assign n23885 = n1081 & ~n14164 ;
  assign n23886 = n23885 ^ n8219 ^ 1'b0 ;
  assign n23887 = ~n7483 & n13058 ;
  assign n23888 = ( ~n16621 & n23382 ) | ( ~n16621 & n23887 ) | ( n23382 & n23887 ) ;
  assign n23889 = n8703 ^ n616 ^ 1'b0 ;
  assign n23890 = n23889 ^ n17830 ^ 1'b0 ;
  assign n23891 = n11377 ^ n4506 ^ n3951 ;
  assign n23892 = n83 | n9041 ;
  assign n23893 = ~n3158 & n9116 ;
  assign n23894 = n11365 & n23893 ;
  assign n23895 = n2672 | n23894 ;
  assign n23896 = n2704 | n23895 ;
  assign n23897 = n11764 | n19484 ;
  assign n23898 = n23896 | n23897 ;
  assign n23899 = n16842 ^ n322 ^ 1'b0 ;
  assign n23900 = ~n6764 & n23899 ;
  assign n23901 = n23900 ^ n5516 ^ 1'b0 ;
  assign n23902 = ~n212 & n4129 ;
  assign n23903 = n16 & ~n5343 ;
  assign n23904 = n23902 & n23903 ;
  assign n23905 = n722 | n12438 ;
  assign n23906 = n15271 ^ n395 ^ 1'b0 ;
  assign n23907 = n1236 & ~n23906 ;
  assign n23908 = ~n498 & n3457 ;
  assign n23909 = ~n9441 & n23908 ;
  assign n23910 = n2138 & ~n2242 ;
  assign n23911 = n23910 ^ n20277 ^ 1'b0 ;
  assign n23912 = n13359 & n23911 ;
  assign n23913 = n23909 & n23912 ;
  assign n23914 = n16708 ^ n6421 ^ 1'b0 ;
  assign n23915 = n23913 | n23914 ;
  assign n23916 = ~n15711 & n16321 ;
  assign n23917 = n23916 ^ n2453 ^ 1'b0 ;
  assign n23918 = n12168 ^ n3227 ^ 1'b0 ;
  assign n23919 = n23917 & n23918 ;
  assign n23922 = n16477 ^ n9049 ^ n7542 ;
  assign n23920 = n294 & n2333 ;
  assign n23921 = n13931 & ~n23920 ;
  assign n23923 = n23922 ^ n23921 ^ 1'b0 ;
  assign n23924 = n3069 & ~n23923 ;
  assign n23925 = n5828 | n13806 ;
  assign n23926 = n18191 | n23925 ;
  assign n23927 = n17483 & ~n23926 ;
  assign n23928 = n3664 | n10203 ;
  assign n23929 = n12463 | n23928 ;
  assign n23930 = n5623 | n8886 ;
  assign n23931 = n9507 ^ n7799 ^ 1'b0 ;
  assign n23932 = n6995 ^ n3368 ^ 1'b0 ;
  assign n23933 = ~n3892 & n23932 ;
  assign n23934 = n23933 ^ n4363 ^ 1'b0 ;
  assign n23935 = n20967 | n23934 ;
  assign n23936 = n17432 ^ n9567 ^ 1'b0 ;
  assign n23937 = n2476 & n23936 ;
  assign n23938 = n20415 ^ n20231 ^ 1'b0 ;
  assign n23939 = n23937 & n23938 ;
  assign n23940 = n16344 & n18144 ;
  assign n23941 = n23940 ^ n5884 ^ 1'b0 ;
  assign n23942 = n15677 ^ n6870 ^ 1'b0 ;
  assign n23943 = n3339 ^ n2650 ^ 1'b0 ;
  assign n23944 = n13800 & n23943 ;
  assign n23945 = n2618 ^ n687 ^ 1'b0 ;
  assign n23946 = n20478 & n23945 ;
  assign n23947 = ~n935 & n16029 ;
  assign n23948 = ( n252 & n1414 ) | ( n252 & ~n2862 ) | ( n1414 & ~n2862 ) ;
  assign n23949 = n23948 ^ n12973 ^ n2911 ;
  assign n23950 = n2282 | n23949 ;
  assign n23951 = ~n4657 & n14727 ;
  assign n23952 = n23951 ^ n8130 ^ 1'b0 ;
  assign n23953 = n2819 & n7918 ;
  assign n23954 = n23953 ^ n6476 ^ 1'b0 ;
  assign n23955 = n18557 ^ n17630 ^ 1'b0 ;
  assign n23956 = n11845 ^ n3758 ^ 1'b0 ;
  assign n23957 = n20278 ^ n3311 ^ 1'b0 ;
  assign n23959 = ~n200 & n392 ;
  assign n23960 = ~n392 & n23959 ;
  assign n23961 = n3077 | n23960 ;
  assign n23958 = ~n1953 & n3784 ;
  assign n23962 = n23961 ^ n23958 ^ 1'b0 ;
  assign n23963 = n23962 ^ n5202 ^ 1'b0 ;
  assign n23964 = n19599 & n23963 ;
  assign n23965 = ~n1637 & n6232 ;
  assign n23966 = n21963 & n23965 ;
  assign n23967 = n23966 ^ n18596 ^ 1'b0 ;
  assign n23968 = ~n1426 & n19561 ;
  assign n23969 = n5915 & ~n12903 ;
  assign n23970 = n9639 | n23969 ;
  assign n23971 = n1483 & n3926 ;
  assign n23972 = n23971 ^ n7418 ^ 1'b0 ;
  assign n23973 = n6900 & n23972 ;
  assign n23977 = n3156 & n3546 ;
  assign n23975 = n3027 ^ n156 ^ 1'b0 ;
  assign n23974 = n13293 & n15686 ;
  assign n23976 = n23975 ^ n23974 ^ 1'b0 ;
  assign n23978 = n23977 ^ n23976 ^ n310 ;
  assign n23979 = n11330 ^ n10132 ^ 1'b0 ;
  assign n23980 = n23979 ^ n3452 ^ 1'b0 ;
  assign n23982 = n3101 | n9880 ;
  assign n23983 = n9435 ^ n901 ^ 1'b0 ;
  assign n23984 = n23982 | n23983 ;
  assign n23981 = n6419 ^ n1608 ^ 1'b0 ;
  assign n23985 = n23984 ^ n23981 ^ 1'b0 ;
  assign n23987 = n3193 | n7438 ;
  assign n23988 = n2549 & ~n14893 ;
  assign n23989 = n23987 & n23988 ;
  assign n23986 = n9952 & n17364 ;
  assign n23990 = n23989 ^ n23986 ^ 1'b0 ;
  assign n23991 = n133 | n11220 ;
  assign n23992 = n23991 ^ n2264 ^ 1'b0 ;
  assign n23993 = ~n10973 & n23992 ;
  assign n23994 = n4231 ^ n938 ^ 1'b0 ;
  assign n23995 = n12163 ^ n8797 ^ 1'b0 ;
  assign n23996 = n2572 & n23995 ;
  assign n23997 = n1316 & n1415 ;
  assign n23998 = ~n450 & n23997 ;
  assign n23999 = n19039 ^ n2418 ^ 1'b0 ;
  assign n24000 = n2813 & n4334 ;
  assign n24001 = n19311 & ~n24000 ;
  assign n24002 = n24001 ^ n15916 ^ 1'b0 ;
  assign n24003 = ~n21254 & n24002 ;
  assign n24005 = n1518 & ~n10178 ;
  assign n24006 = ~n7447 & n24005 ;
  assign n24004 = n5691 | n12014 ;
  assign n24007 = n24006 ^ n24004 ^ n8497 ;
  assign n24008 = n18172 ^ n11863 ^ 1'b0 ;
  assign n24009 = n20683 ^ n495 ^ 1'b0 ;
  assign n24010 = n10053 & n12993 ;
  assign n24011 = n323 & ~n11778 ;
  assign n24012 = n2811 & ~n9326 ;
  assign n24013 = n6664 & n24012 ;
  assign n24014 = n3526 & ~n24013 ;
  assign n24015 = n24014 ^ n14422 ^ 1'b0 ;
  assign n24016 = n1785 ^ n804 ^ 1'b0 ;
  assign n24017 = ~n7093 & n24016 ;
  assign n24018 = n24017 ^ n22278 ^ 1'b0 ;
  assign n24019 = n13782 & n17953 ;
  assign n24020 = n12078 ^ n2223 ^ 1'b0 ;
  assign n24021 = n8405 & ~n22387 ;
  assign n24022 = n17959 & n24021 ;
  assign n24023 = n17272 ^ n4577 ^ 1'b0 ;
  assign n24024 = n13920 ^ n12448 ^ 1'b0 ;
  assign n24025 = n18403 ^ n11758 ^ 1'b0 ;
  assign n24026 = n22535 & n24025 ;
  assign n24027 = n7487 & n13450 ;
  assign n24028 = n10664 ^ n2484 ^ 1'b0 ;
  assign n24029 = n8034 & ~n24028 ;
  assign n24031 = ~n6595 & n12692 ;
  assign n24032 = n24031 ^ n16803 ^ 1'b0 ;
  assign n24030 = ~n10873 & n15512 ;
  assign n24033 = n24032 ^ n24030 ^ 1'b0 ;
  assign n24034 = n8897 ^ n8477 ^ 1'b0 ;
  assign n24035 = n23384 | n24034 ;
  assign n24036 = n1598 & ~n2449 ;
  assign n24037 = ~n3744 & n18832 ;
  assign n24038 = ~n24036 & n24037 ;
  assign n24039 = n857 | n9368 ;
  assign n24040 = n24039 ^ n6923 ^ 1'b0 ;
  assign n24041 = n1364 & ~n1662 ;
  assign n24042 = n2929 & n24041 ;
  assign n24043 = n24042 ^ n1877 ^ 1'b0 ;
  assign n24044 = n24040 & ~n24043 ;
  assign n24045 = n3941 & ~n7460 ;
  assign n24046 = n22924 ^ n6417 ^ 1'b0 ;
  assign n24047 = ~n18061 & n24046 ;
  assign n24048 = n24047 ^ n3135 ^ 1'b0 ;
  assign n24049 = n24045 | n24048 ;
  assign n24050 = ~n7674 & n23696 ;
  assign n24051 = n24050 ^ n4629 ^ 1'b0 ;
  assign n24052 = n21064 ^ n6407 ^ 1'b0 ;
  assign n24053 = n17323 ^ n1155 ^ n567 ;
  assign n24054 = n14185 ^ n8755 ^ 1'b0 ;
  assign n24055 = n24053 & n24054 ;
  assign n24056 = n2686 & n19138 ;
  assign n24057 = ~n624 & n24056 ;
  assign n24058 = n8630 ^ n2322 ^ 1'b0 ;
  assign n24059 = n15631 ^ n7155 ^ 1'b0 ;
  assign n24060 = n1368 ^ n907 ^ 1'b0 ;
  assign n24061 = n24060 ^ n977 ^ 1'b0 ;
  assign n24062 = n19689 ^ n12436 ^ 1'b0 ;
  assign n24063 = n24062 ^ n113 ^ 1'b0 ;
  assign n24065 = n2472 & n5152 ;
  assign n24064 = ~n10777 & n18977 ;
  assign n24066 = n24065 ^ n24064 ^ 1'b0 ;
  assign n24067 = n21969 ^ n10261 ^ 1'b0 ;
  assign n24068 = n5048 & n21085 ;
  assign n24069 = n24068 ^ n5564 ^ 1'b0 ;
  assign n24070 = ( n901 & n8253 ) | ( n901 & n24069 ) | ( n8253 & n24069 ) ;
  assign n24071 = ~n2784 & n6944 ;
  assign n24072 = n24071 ^ n229 ^ 1'b0 ;
  assign n24073 = ~n24070 & n24072 ;
  assign n24074 = n2109 & n4629 ;
  assign n24075 = n4297 & n9918 ;
  assign n24076 = n17581 & n24075 ;
  assign n24077 = x6 | n5143 ;
  assign n24082 = ~n1323 & n3007 ;
  assign n24081 = n7812 & ~n15421 ;
  assign n24083 = n24082 ^ n24081 ^ 1'b0 ;
  assign n24078 = n4097 & n11324 ;
  assign n24079 = n24078 ^ n7254 ^ 1'b0 ;
  assign n24080 = n19804 | n24079 ;
  assign n24084 = n24083 ^ n24080 ^ 1'b0 ;
  assign n24085 = n2107 & n2910 ;
  assign n24086 = n24085 ^ n9434 ^ 1'b0 ;
  assign n24087 = n14933 ^ n3318 ^ 1'b0 ;
  assign n24088 = n1458 & ~n24087 ;
  assign n24089 = n12935 ^ n10347 ^ n3950 ;
  assign n24090 = n24088 | n24089 ;
  assign n24091 = ~n11319 & n19584 ;
  assign n24092 = ~n2216 & n8990 ;
  assign n24093 = n3477 & n17765 ;
  assign n24094 = n24093 ^ n489 ^ 1'b0 ;
  assign n24095 = n4171 | n8705 ;
  assign n24096 = n24095 ^ n9971 ^ 1'b0 ;
  assign n24097 = n10847 ^ n3452 ^ 1'b0 ;
  assign n24098 = n2916 | n24097 ;
  assign n24099 = n24096 & ~n24098 ;
  assign n24100 = n1206 | n4698 ;
  assign n24101 = n21647 & ~n24100 ;
  assign n24102 = n19617 ^ n10389 ^ n2281 ;
  assign n24103 = n24102 ^ n469 ^ 1'b0 ;
  assign n24104 = ~n1868 & n2921 ;
  assign n24105 = ~n1464 & n2371 ;
  assign n24106 = ~n1877 & n24105 ;
  assign n24107 = n1655 & n24106 ;
  assign n24108 = n24107 ^ n576 ^ 1'b0 ;
  assign n24109 = ~n4018 & n15676 ;
  assign n24110 = ~n2848 & n23209 ;
  assign n24111 = ~n6206 & n7968 ;
  assign n24112 = n24111 ^ n2757 ^ 1'b0 ;
  assign n24113 = n3690 | n4439 ;
  assign n24114 = n24112 | n24113 ;
  assign n24115 = n24114 ^ n979 ^ 1'b0 ;
  assign n24116 = ~n339 & n24115 ;
  assign n24117 = n10827 & n16967 ;
  assign n24118 = ~n24116 & n24117 ;
  assign n24119 = n382 | n2380 ;
  assign n24120 = n2851 ^ n2644 ^ 1'b0 ;
  assign n24121 = n8730 | n24120 ;
  assign n24122 = n7495 | n24121 ;
  assign n24123 = n2949 & n24122 ;
  assign n24124 = ~n19296 & n22085 ;
  assign n24125 = n7735 & n12099 ;
  assign n24126 = n3841 ^ n883 ^ 1'b0 ;
  assign n24127 = ~n1164 & n24126 ;
  assign n24128 = ~n2959 & n24127 ;
  assign n24129 = n11859 | n15624 ;
  assign n24130 = n1531 | n24129 ;
  assign n24131 = n24130 ^ n10769 ^ 1'b0 ;
  assign n24132 = ~n1999 & n24131 ;
  assign n24133 = n8231 ^ n7936 ^ 1'b0 ;
  assign n24134 = n3137 & n3539 ;
  assign n24135 = n1385 | n24134 ;
  assign n24136 = n1248 | n7673 ;
  assign n24137 = n6541 & ~n24136 ;
  assign n24138 = n14395 ^ n6281 ^ 1'b0 ;
  assign n24139 = n1531 & ~n15490 ;
  assign n24140 = n16202 ^ n1867 ^ 1'b0 ;
  assign n24141 = n5625 & ~n24140 ;
  assign n24142 = n1231 | n22259 ;
  assign n24143 = n2933 & ~n6327 ;
  assign n24144 = n22609 ^ n7054 ^ 1'b0 ;
  assign n24145 = n24143 & n24144 ;
  assign n24147 = n194 & n330 ;
  assign n24148 = n24147 ^ n8990 ^ 1'b0 ;
  assign n24146 = n2107 | n4054 ;
  assign n24149 = n24148 ^ n24146 ^ n3642 ;
  assign n24150 = n24149 ^ n3586 ^ 1'b0 ;
  assign n24151 = n19563 & n24150 ;
  assign n24152 = n14483 | n21999 ;
  assign n24153 = ~n1117 & n1660 ;
  assign n24154 = n24153 ^ n2412 ^ 1'b0 ;
  assign n24155 = ~n20577 & n24154 ;
  assign n24156 = n24155 ^ n475 ^ 1'b0 ;
  assign n24157 = n14731 & n24156 ;
  assign n24158 = n5873 & n24157 ;
  assign n24159 = n323 & n2850 ;
  assign n24160 = ~n12680 & n24159 ;
  assign n24161 = n13197 & n24160 ;
  assign n24162 = n5911 & n15792 ;
  assign n24163 = n4516 & n8750 ;
  assign n24164 = ~n7250 & n24163 ;
  assign n24165 = ~n9346 & n24164 ;
  assign n24166 = n469 | n24165 ;
  assign n24167 = n24166 ^ n4584 ^ 1'b0 ;
  assign n24168 = n15963 ^ n14072 ^ 1'b0 ;
  assign n24169 = n9823 & n24168 ;
  assign n24170 = n21509 & ~n22471 ;
  assign n24171 = n21412 & n24170 ;
  assign n24172 = n848 & n1053 ;
  assign n24173 = n1944 & ~n4295 ;
  assign n24174 = n24173 ^ n1957 ^ 1'b0 ;
  assign n24175 = ~n24172 & n24174 ;
  assign n24176 = n1258 | n2869 ;
  assign n24177 = n8760 | n24176 ;
  assign n24178 = n3032 ^ n497 ^ 1'b0 ;
  assign n24179 = n3037 & n24178 ;
  assign n24180 = n24179 ^ n6345 ^ 1'b0 ;
  assign n24181 = n22669 & ~n24180 ;
  assign n24182 = n2064 & n16905 ;
  assign n24183 = ~n5507 & n24182 ;
  assign n24184 = n1025 ^ n367 ^ 1'b0 ;
  assign n24185 = n6250 & ~n24184 ;
  assign n24186 = n14241 ^ n8442 ^ 1'b0 ;
  assign n24187 = n4793 & n8705 ;
  assign n24188 = ~n8705 & n24187 ;
  assign n24189 = n2925 & n5186 ;
  assign n24190 = ~n2925 & n24189 ;
  assign n24191 = n2862 & n24190 ;
  assign n24192 = ~n15931 & n24191 ;
  assign n24193 = n2885 & n24192 ;
  assign n24194 = n24193 ^ n4784 ^ 1'b0 ;
  assign n24195 = n24188 | n24194 ;
  assign n24196 = n3218 & ~n9291 ;
  assign n24197 = n9447 & n24196 ;
  assign n24198 = ~n15532 & n24197 ;
  assign n24199 = ( n4645 & n9566 ) | ( n4645 & ~n18550 ) | ( n9566 & ~n18550 ) ;
  assign n24200 = n24199 ^ n3063 ^ 1'b0 ;
  assign n24201 = n15773 & n24200 ;
  assign n24202 = ~n21479 & n24201 ;
  assign n24203 = n15602 ^ n3651 ^ 1'b0 ;
  assign n24204 = n12804 & ~n24203 ;
  assign n24205 = n10749 & n24204 ;
  assign n24206 = n24205 ^ n20875 ^ 1'b0 ;
  assign n24207 = n97 & n5626 ;
  assign n24208 = n9381 ^ n255 ^ 1'b0 ;
  assign n24209 = n4466 | n24208 ;
  assign n24210 = n294 & n11379 ;
  assign n24211 = ~n6085 & n24210 ;
  assign n24212 = n5780 & n8881 ;
  assign n24213 = n5358 & ~n11904 ;
  assign n24214 = n19358 ^ n14834 ^ 1'b0 ;
  assign n24215 = n19263 ^ n1138 ^ 1'b0 ;
  assign n24216 = n7455 & n24215 ;
  assign n24217 = ( n6647 & n24214 ) | ( n6647 & n24216 ) | ( n24214 & n24216 ) ;
  assign n24218 = n21597 ^ n10288 ^ 1'b0 ;
  assign n24219 = n2278 | n14386 ;
  assign n24220 = n24219 ^ n13277 ^ 1'b0 ;
  assign n24221 = n1608 | n8503 ;
  assign n24222 = n6709 & ~n24221 ;
  assign n24223 = ( n7512 & n18091 ) | ( n7512 & ~n21298 ) | ( n18091 & ~n21298 ) ;
  assign n24224 = n9739 ^ n8110 ^ 1'b0 ;
  assign n24225 = ~n10818 & n24224 ;
  assign n24226 = ~n9791 & n14714 ;
  assign n24227 = n6876 & n24226 ;
  assign n24228 = n10741 ^ n5554 ^ 1'b0 ;
  assign n24229 = n24228 ^ n16625 ^ n15674 ;
  assign n24230 = ~n3845 & n9566 ;
  assign n24231 = n24230 ^ n6376 ^ 1'b0 ;
  assign n24232 = n5645 ^ n4937 ^ 1'b0 ;
  assign n24233 = n6296 & n23872 ;
  assign n24234 = n23455 ^ n3278 ^ 1'b0 ;
  assign n24235 = ~n15414 & n24234 ;
  assign n24236 = n3775 ^ n2145 ^ 1'b0 ;
  assign n24237 = n24236 ^ n5428 ^ 1'b0 ;
  assign n24238 = ~n7192 & n24237 ;
  assign n24239 = n16379 ^ n10982 ^ 1'b0 ;
  assign n24240 = n24239 ^ n19131 ^ n19129 ;
  assign n24241 = ~n1778 & n10837 ;
  assign n24242 = n24241 ^ n12687 ^ 1'b0 ;
  assign n24243 = n5410 ^ n1964 ^ 1'b0 ;
  assign n24244 = n68 & n24243 ;
  assign n24245 = n24244 ^ n5067 ^ 1'b0 ;
  assign n24246 = n11275 | n24245 ;
  assign n24247 = n24246 ^ n1048 ^ 1'b0 ;
  assign n24248 = n615 | n9065 ;
  assign n24249 = n24247 & ~n24248 ;
  assign n24250 = n3380 | n24249 ;
  assign n24251 = n24250 ^ n4794 ^ 1'b0 ;
  assign n24252 = n4812 & n10161 ;
  assign n24253 = ( n113 & ~n14708 ) | ( n113 & n18436 ) | ( ~n14708 & n18436 ) ;
  assign n24254 = n8466 & ~n24253 ;
  assign n24255 = n2101 & ~n3563 ;
  assign n24256 = n6102 ^ n97 ^ 1'b0 ;
  assign n24257 = n24256 ^ n10842 ^ 1'b0 ;
  assign n24258 = ~n13869 & n24257 ;
  assign n24259 = n24258 ^ n12242 ^ 1'b0 ;
  assign n24260 = ~n5793 & n6569 ;
  assign n24261 = n19580 ^ n5205 ^ 1'b0 ;
  assign n24262 = ~n17589 & n24261 ;
  assign n24263 = n24262 ^ n15866 ^ 1'b0 ;
  assign n24264 = n24260 & n24263 ;
  assign n24265 = ~n13887 & n24264 ;
  assign n24268 = n8061 & n20175 ;
  assign n24269 = n1526 & n24268 ;
  assign n24266 = n20713 ^ n6653 ^ 1'b0 ;
  assign n24267 = n8192 | n24266 ;
  assign n24270 = n24269 ^ n24267 ^ n15569 ;
  assign n24271 = n3483 & ~n3771 ;
  assign n24272 = n215 | n1205 ;
  assign n24273 = n23449 | n24272 ;
  assign n24274 = n16916 & ~n24273 ;
  assign n24275 = n24271 & n24274 ;
  assign n24276 = n6493 | n15786 ;
  assign n24277 = n950 | n24276 ;
  assign n24278 = n17227 | n23242 ;
  assign n24279 = n922 | n24278 ;
  assign n24286 = n3940 ^ n1219 ^ 1'b0 ;
  assign n24287 = n4550 & n24286 ;
  assign n24280 = n3535 ^ n1210 ^ 1'b0 ;
  assign n24281 = ~n4137 & n24280 ;
  assign n24282 = n229 & n24281 ;
  assign n24283 = n19583 & n24282 ;
  assign n24284 = ~n5463 & n7967 ;
  assign n24285 = ~n24283 & n24284 ;
  assign n24288 = n24287 ^ n24285 ^ 1'b0 ;
  assign n24289 = n20121 ^ n443 ^ 1'b0 ;
  assign n24290 = n8128 & ~n24289 ;
  assign n24291 = n740 & n24290 ;
  assign n24292 = n653 | n12284 ;
  assign n24293 = n24292 ^ n1198 ^ 1'b0 ;
  assign n24294 = n19264 ^ n5250 ^ 1'b0 ;
  assign n24295 = ~n16039 & n24294 ;
  assign n24296 = ~n12928 & n24295 ;
  assign n24297 = n24296 ^ n6388 ^ 1'b0 ;
  assign n24298 = n13086 ^ n1790 ^ 1'b0 ;
  assign n24299 = n15204 & n24298 ;
  assign n24300 = n1602 | n4700 ;
  assign n24301 = n19202 & ~n19332 ;
  assign n24302 = n24301 ^ n14561 ^ 1'b0 ;
  assign n24303 = n812 & ~n1940 ;
  assign n24304 = n988 | n21010 ;
  assign n24305 = n24303 | n24304 ;
  assign n24306 = ~n177 & n7476 ;
  assign n24307 = n24306 ^ n13901 ^ 1'b0 ;
  assign n24308 = ~n10513 & n22875 ;
  assign n24309 = n24308 ^ n3037 ^ 1'b0 ;
  assign n24310 = n14158 & ~n24309 ;
  assign n24311 = n6814 | n21456 ;
  assign n24312 = n24310 | n24311 ;
  assign n24313 = ~n6080 & n19013 ;
  assign n24314 = ~n13648 & n24313 ;
  assign n24315 = n24314 ^ n3321 ^ 1'b0 ;
  assign n24316 = n17238 ^ n963 ^ 1'b0 ;
  assign n24317 = n8718 & ~n24316 ;
  assign n24318 = n6150 & n24317 ;
  assign n24319 = ~n4451 & n24075 ;
  assign n24320 = n24319 ^ n20322 ^ 1'b0 ;
  assign n24321 = n1058 | n8021 ;
  assign n24322 = n24321 ^ n633 ^ 1'b0 ;
  assign n24323 = n24322 ^ n9577 ^ 1'b0 ;
  assign n24324 = ~n10113 & n24323 ;
  assign n24325 = n662 | n24089 ;
  assign n24326 = ~n302 & n11277 ;
  assign n24327 = n8295 | n24326 ;
  assign n24328 = n24327 ^ n77 ^ 1'b0 ;
  assign n24329 = n3718 & ~n7548 ;
  assign n24330 = ~n82 & n3794 ;
  assign n24331 = n13385 & ~n24330 ;
  assign n24332 = ~n12757 & n24331 ;
  assign n24333 = n10191 | n13556 ;
  assign n24334 = n158 | n10735 ;
  assign n24335 = n2764 & ~n24334 ;
  assign n24337 = ~n1438 & n22597 ;
  assign n24338 = n23286 & n24337 ;
  assign n24336 = n3141 & n4482 ;
  assign n24339 = n24338 ^ n24336 ^ 1'b0 ;
  assign n24340 = n10030 ^ n8033 ^ n97 ;
  assign n24341 = n11343 | n13432 ;
  assign n24342 = n155 & n4227 ;
  assign n24343 = n24342 ^ n4320 ^ 1'b0 ;
  assign n24344 = n6475 & ~n6833 ;
  assign n24345 = ~n24343 & n24344 ;
  assign n24346 = n2303 & n24345 ;
  assign n24347 = ~n1591 & n20011 ;
  assign n24348 = n532 | n5250 ;
  assign n24349 = n24348 ^ n12997 ^ 1'b0 ;
  assign n24350 = n24349 ^ n20220 ^ 1'b0 ;
  assign n24351 = n24350 ^ n12171 ^ 1'b0 ;
  assign n24352 = n15910 ^ n1315 ^ 1'b0 ;
  assign n24353 = n3269 ^ n1198 ^ 1'b0 ;
  assign n24354 = n2279 & ~n4385 ;
  assign n24355 = ( n2316 & n24353 ) | ( n2316 & ~n24354 ) | ( n24353 & ~n24354 ) ;
  assign n24356 = ~n1491 & n2910 ;
  assign n24357 = n9029 | n15627 ;
  assign n24358 = n15905 & ~n24357 ;
  assign n24359 = n24356 & ~n24358 ;
  assign n24360 = n24359 ^ n2027 ^ 1'b0 ;
  assign n24361 = n142 | n17367 ;
  assign n24362 = n638 & ~n8135 ;
  assign n24363 = n24362 ^ n8410 ^ 1'b0 ;
  assign n24364 = ~n1961 & n2945 ;
  assign n24365 = n24363 & n24364 ;
  assign n24366 = n3485 | n20313 ;
  assign n24367 = n24366 ^ n2922 ^ 1'b0 ;
  assign n24368 = ~n4580 & n23274 ;
  assign n24369 = n4493 ^ n535 ^ 1'b0 ;
  assign n24370 = n5861 & ~n24369 ;
  assign n24371 = n3127 | n19377 ;
  assign n24372 = n3061 & ~n5806 ;
  assign n24373 = n321 & n758 ;
  assign n24376 = n17439 ^ n3827 ^ 1'b0 ;
  assign n24377 = n5187 | n24376 ;
  assign n24374 = n458 | n9019 ;
  assign n24375 = n24374 ^ n800 ^ 1'b0 ;
  assign n24378 = n24377 ^ n24375 ^ 1'b0 ;
  assign n24379 = n15304 & ~n19772 ;
  assign n24380 = n24379 ^ n10584 ^ 1'b0 ;
  assign n24381 = n5710 & n19826 ;
  assign n24382 = n24380 | n24381 ;
  assign n24383 = n1157 ^ n512 ^ 1'b0 ;
  assign n24384 = n1953 & ~n24383 ;
  assign n24385 = n1469 & n5590 ;
  assign n24386 = ~n10358 & n24385 ;
  assign n24389 = n20599 ^ n6539 ^ 1'b0 ;
  assign n24387 = ~n2320 & n2565 ;
  assign n24388 = n11351 | n24387 ;
  assign n24390 = n24389 ^ n24388 ^ 1'b0 ;
  assign n24391 = n11551 ^ n847 ^ 1'b0 ;
  assign n24392 = n3385 ^ n1645 ^ 1'b0 ;
  assign n24393 = n13588 & ~n24392 ;
  assign n24394 = n16675 ^ n397 ^ 1'b0 ;
  assign n24395 = n4332 & ~n20807 ;
  assign n24396 = ~n24394 & n24395 ;
  assign n24397 = ~n12411 & n21123 ;
  assign n24398 = ( n6095 & n6426 ) | ( n6095 & ~n23583 ) | ( n6426 & ~n23583 ) ;
  assign n24399 = n20694 ^ n2751 ^ 1'b0 ;
  assign n24400 = n4552 & ~n8226 ;
  assign n24401 = n9581 | n24400 ;
  assign n24402 = n2545 | n3674 ;
  assign n24403 = n5468 | n24402 ;
  assign n24404 = n24403 ^ n5904 ^ 1'b0 ;
  assign n24405 = ~n10168 & n24404 ;
  assign n24406 = ~n3765 & n15367 ;
  assign n24407 = n24406 ^ n2097 ^ 1'b0 ;
  assign n24408 = ~n10625 & n23911 ;
  assign n24409 = n23377 ^ n1816 ^ 1'b0 ;
  assign n24410 = n21773 | n24409 ;
  assign n24411 = n198 | n11302 ;
  assign n24412 = n9077 | n24411 ;
  assign n24413 = ( n10534 & n15045 ) | ( n10534 & n24412 ) | ( n15045 & n24412 ) ;
  assign n24414 = n1142 & n10707 ;
  assign n24415 = n24414 ^ n1934 ^ 1'b0 ;
  assign n24416 = ~n715 & n23197 ;
  assign n24417 = n6758 ^ n44 ^ 1'b0 ;
  assign n24418 = n24416 & ~n24417 ;
  assign n24419 = n7195 & n19933 ;
  assign n24420 = n24419 ^ n16311 ^ n5639 ;
  assign n24421 = ~n4098 & n24420 ;
  assign n24422 = n24421 ^ n3483 ^ n1852 ;
  assign n24423 = n24418 & ~n24422 ;
  assign n24424 = ~n7399 & n24423 ;
  assign n24425 = n1081 & ~n13608 ;
  assign n24426 = ~n4307 & n24425 ;
  assign n24427 = n24426 ^ n7670 ^ 1'b0 ;
  assign n24428 = ( n1855 & ~n7909 ) | ( n1855 & n18555 ) | ( ~n7909 & n18555 ) ;
  assign n24429 = n19364 ^ n78 ^ 1'b0 ;
  assign n24430 = ~n24428 & n24429 ;
  assign n24431 = n24430 ^ n1318 ^ 1'b0 ;
  assign n24432 = n7958 ^ n6589 ^ n880 ;
  assign n24433 = n12692 & ~n24432 ;
  assign n24434 = n5950 & ~n6154 ;
  assign n24435 = n24434 ^ n817 ^ 1'b0 ;
  assign n24436 = n24435 ^ n8195 ^ 1'b0 ;
  assign n24437 = n24433 & ~n24436 ;
  assign n24438 = n4904 ^ n1185 ^ 1'b0 ;
  assign n24439 = n2799 & n24438 ;
  assign n24440 = n10383 & n24439 ;
  assign n24441 = n14321 & n24440 ;
  assign n24442 = n19198 ^ n6948 ^ 1'b0 ;
  assign n24443 = n2218 & n3243 ;
  assign n24444 = n24443 ^ n21993 ^ 1'b0 ;
  assign n24445 = ~n24442 & n24444 ;
  assign n24446 = n17637 ^ n3137 ^ 1'b0 ;
  assign n24447 = n1304 & ~n24446 ;
  assign n24448 = ~n1856 & n24447 ;
  assign n24449 = ~n4387 & n14077 ;
  assign n24450 = ~n653 & n17774 ;
  assign n24451 = n9840 & n24450 ;
  assign n24452 = n24451 ^ n8869 ^ 1'b0 ;
  assign n24454 = n281 | n1396 ;
  assign n24453 = n11272 & ~n19751 ;
  assign n24455 = n24454 ^ n24453 ^ 1'b0 ;
  assign n24456 = n3099 & ~n15824 ;
  assign n24457 = n1824 & n24456 ;
  assign n24458 = n23626 | n24457 ;
  assign n24459 = n23681 ^ n2949 ^ 1'b0 ;
  assign n24460 = n24164 | n24459 ;
  assign n24461 = n3233 | n13763 ;
  assign n24462 = n3141 | n24461 ;
  assign n24463 = n5520 & n24462 ;
  assign n24464 = n24463 ^ n15613 ^ 1'b0 ;
  assign n24465 = n23079 | n24464 ;
  assign n24466 = n11542 | n11766 ;
  assign n24467 = n448 & n16654 ;
  assign n24468 = ~n24466 & n24467 ;
  assign n24469 = n24468 ^ n10058 ^ 1'b0 ;
  assign n24470 = n24469 ^ n5922 ^ 1'b0 ;
  assign n24471 = n3557 & n12057 ;
  assign n24472 = n13768 & n24471 ;
  assign n24473 = n24470 & ~n24472 ;
  assign n24474 = n3827 & ~n24473 ;
  assign n24475 = n24474 ^ n21212 ^ 1'b0 ;
  assign n24476 = n12318 ^ n1010 ^ 1'b0 ;
  assign n24477 = n14936 | n24476 ;
  assign n24478 = n8896 ^ n2767 ^ 1'b0 ;
  assign n24479 = n828 & n7827 ;
  assign n24480 = n4814 ^ n2382 ^ 1'b0 ;
  assign n24481 = n8377 & ~n24480 ;
  assign n24482 = n593 & ~n24481 ;
  assign n24483 = n2137 | n4784 ;
  assign n24486 = n19003 & n19420 ;
  assign n24487 = n24486 ^ n5564 ^ 1'b0 ;
  assign n24484 = n8500 ^ n2963 ^ 1'b0 ;
  assign n24485 = n4927 & ~n24484 ;
  assign n24488 = n24487 ^ n24485 ^ 1'b0 ;
  assign n24490 = n7449 ^ n7247 ^ 1'b0 ;
  assign n24489 = n252 | n7438 ;
  assign n24491 = n24490 ^ n24489 ^ 1'b0 ;
  assign n24492 = n3295 & ~n4726 ;
  assign n24493 = n6230 ^ n2927 ^ 1'b0 ;
  assign n24494 = n17631 & ~n24493 ;
  assign n24495 = n14066 ^ n9327 ^ 1'b0 ;
  assign n24496 = n19482 | n24495 ;
  assign n24497 = ~n1858 & n7179 ;
  assign n24498 = ( n835 & ~n5194 ) | ( n835 & n24497 ) | ( ~n5194 & n24497 ) ;
  assign n24499 = n2700 & ~n14344 ;
  assign n24500 = n24499 ^ n4902 ^ 1'b0 ;
  assign n24501 = n9988 & ~n24500 ;
  assign n24502 = n30 & n8072 ;
  assign n24503 = n3561 ^ n649 ^ 1'b0 ;
  assign n24504 = n13743 | n14355 ;
  assign n24505 = n3845 & n24504 ;
  assign n24506 = n22611 & n24505 ;
  assign n24507 = n18191 & ~n20738 ;
  assign n24509 = n8305 | n10028 ;
  assign n24510 = n4580 & ~n24509 ;
  assign n24508 = n6929 | n14906 ;
  assign n24511 = n24510 ^ n24508 ^ 1'b0 ;
  assign n24512 = ~n10774 & n20109 ;
  assign n24513 = n3504 | n15866 ;
  assign n24514 = n4194 & ~n24513 ;
  assign n24515 = n24512 & ~n24514 ;
  assign n24516 = n1763 & ~n2136 ;
  assign n24517 = n446 | n9488 ;
  assign n24518 = n24517 ^ n11067 ^ 1'b0 ;
  assign n24519 = n8242 & ~n24518 ;
  assign n24520 = n13407 & n24519 ;
  assign n24521 = n21360 | n23940 ;
  assign n24522 = n9901 | n24521 ;
  assign n24523 = ~n9536 & n20301 ;
  assign n24524 = ~n16157 & n24523 ;
  assign n24525 = ~n2080 & n5034 ;
  assign n24526 = ~n7391 & n24525 ;
  assign n24527 = n17507 ^ n11371 ^ 1'b0 ;
  assign n24528 = n24526 | n24527 ;
  assign n24529 = n1144 | n8969 ;
  assign n24530 = n24529 ^ n4404 ^ 1'b0 ;
  assign n24531 = n9662 & n16090 ;
  assign n24532 = n24531 ^ n4620 ^ 1'b0 ;
  assign n24533 = n2060 & n11175 ;
  assign n24534 = ~n4450 & n9409 ;
  assign n24535 = ~n2022 & n22453 ;
  assign n24536 = n19504 ^ n11309 ^ 1'b0 ;
  assign n24537 = ~n4495 & n12249 ;
  assign n24538 = n24537 ^ n14808 ^ 1'b0 ;
  assign n24539 = n1318 & ~n5283 ;
  assign n24540 = n1350 & ~n19383 ;
  assign n24541 = ~n532 & n24540 ;
  assign n24542 = ~n318 & n2388 ;
  assign n24543 = n7403 | n24542 ;
  assign n24544 = n24543 ^ n8790 ^ 1'b0 ;
  assign n24545 = n24544 ^ n11866 ^ 1'b0 ;
  assign n24546 = n24545 ^ n22099 ^ n233 ;
  assign n24547 = n15663 ^ n274 ^ 1'b0 ;
  assign n24548 = n24547 ^ n4156 ^ 1'b0 ;
  assign n24549 = n21719 ^ n2967 ^ 1'b0 ;
  assign n24550 = n21028 & ~n24549 ;
  assign n24551 = n2465 & n5999 ;
  assign n24552 = n20313 ^ n1401 ^ 1'b0 ;
  assign n24553 = ~n6168 & n24552 ;
  assign n24554 = n5825 & n24553 ;
  assign n24555 = n24554 ^ n16637 ^ 1'b0 ;
  assign n24556 = n40 & n9969 ;
  assign n24557 = n7440 & n24556 ;
  assign n24558 = n24557 ^ n467 ^ 1'b0 ;
  assign n24559 = ~n15631 & n24558 ;
  assign n24560 = n10279 | n14608 ;
  assign n24561 = n19880 ^ n151 ^ 1'b0 ;
  assign n24562 = n18803 ^ n11061 ^ 1'b0 ;
  assign n24563 = n1318 ^ n419 ^ 1'b0 ;
  assign n24564 = n19154 ^ x6 ^ 1'b0 ;
  assign n24565 = n24563 | n24564 ;
  assign n24566 = n24565 ^ n2829 ^ n583 ;
  assign n24567 = n14062 ^ n1209 ^ 1'b0 ;
  assign n24568 = n8763 & n23209 ;
  assign n24569 = n5110 ^ n4763 ^ 1'b0 ;
  assign n24570 = n18099 & ~n24569 ;
  assign n24571 = n5836 | n12368 ;
  assign n24572 = n7605 ^ n6544 ^ 1'b0 ;
  assign n24573 = n5245 & ~n24572 ;
  assign n24574 = n8106 ^ n653 ^ 1'b0 ;
  assign n24575 = ~n7283 & n24574 ;
  assign n24576 = n24573 & n24575 ;
  assign n24577 = n10486 | n18579 ;
  assign n24578 = n3334 & n24577 ;
  assign n24579 = n9335 | n24578 ;
  assign n24580 = ~n541 & n12681 ;
  assign n24581 = n24580 ^ n19250 ^ 1'b0 ;
  assign n24582 = n24581 ^ n21324 ^ 1'b0 ;
  assign n24583 = n169 | n19210 ;
  assign n24584 = n2459 & n24583 ;
  assign n24585 = ~n4818 & n21938 ;
  assign n24586 = n24585 ^ n9776 ^ 1'b0 ;
  assign n24587 = n2670 & ~n16828 ;
  assign n24588 = n21749 ^ n17479 ^ 1'b0 ;
  assign n24589 = n24375 & n24588 ;
  assign n24590 = ~n1513 & n3318 ;
  assign n24591 = n12482 & ~n24590 ;
  assign n24592 = n12509 & ~n24591 ;
  assign n24593 = n22355 & ~n24592 ;
  assign n24594 = n2560 | n4740 ;
  assign n24595 = n24594 ^ n18284 ^ 1'b0 ;
  assign n24596 = ( n19 & n1770 ) | ( n19 & ~n24595 ) | ( n1770 & ~n24595 ) ;
  assign n24597 = n2849 | n2998 ;
  assign n24598 = n24597 ^ n184 ^ 1'b0 ;
  assign n24599 = n6262 & ~n24598 ;
  assign n24600 = n2263 & ~n21296 ;
  assign n24601 = n5995 & ~n15370 ;
  assign n24602 = ~n13623 & n24601 ;
  assign n24604 = n5621 ^ n1026 ^ 1'b0 ;
  assign n24605 = n24604 ^ n19478 ^ 1'b0 ;
  assign n24606 = n10635 & ~n24605 ;
  assign n24603 = ~n5465 & n19158 ;
  assign n24607 = n24606 ^ n24603 ^ 1'b0 ;
  assign n24608 = n24607 ^ n7572 ^ 1'b0 ;
  assign n24609 = n7411 & ~n14146 ;
  assign n24610 = n22205 & ~n24609 ;
  assign n24611 = n24610 ^ n2566 ^ 1'b0 ;
  assign n24612 = n24611 ^ n18053 ^ 1'b0 ;
  assign n24613 = n535 & n15691 ;
  assign n24614 = n958 | n7138 ;
  assign n24615 = n24614 ^ n1036 ^ 1'b0 ;
  assign n24616 = n10079 | n24615 ;
  assign n24617 = n24616 ^ n9326 ^ 1'b0 ;
  assign n24618 = n24617 ^ n8472 ^ 1'b0 ;
  assign n24619 = n13682 & ~n17118 ;
  assign n24620 = ~n12887 & n19495 ;
  assign n24621 = n11478 ^ n6723 ^ 1'b0 ;
  assign n24622 = n7241 | n24621 ;
  assign n24623 = ~n2761 & n24622 ;
  assign n24624 = n13532 | n24623 ;
  assign n24625 = n9131 & ~n9727 ;
  assign n24626 = n22621 & n24625 ;
  assign n24627 = n15668 ^ n4754 ^ 1'b0 ;
  assign n24628 = n627 & n23282 ;
  assign n24629 = n13450 & ~n24628 ;
  assign n24630 = ~n192 & n12529 ;
  assign n24631 = n24630 ^ n16812 ^ 1'b0 ;
  assign n24632 = n1907 | n13419 ;
  assign n24633 = n348 | n24632 ;
  assign n24634 = n24633 ^ n4852 ^ 1'b0 ;
  assign n24635 = n12725 & ~n24634 ;
  assign n24636 = n2657 & n24635 ;
  assign n24637 = n690 & n24636 ;
  assign n24638 = ~n3346 & n3650 ;
  assign n24639 = n24637 | n24638 ;
  assign n24640 = n24639 ^ n8485 ^ 1'b0 ;
  assign n24641 = n4784 | n24640 ;
  assign n24642 = n2517 | n10423 ;
  assign n24643 = n419 & ~n6275 ;
  assign n24644 = n9107 & n19632 ;
  assign n24645 = n24644 ^ n4274 ^ 1'b0 ;
  assign n24646 = ~n11645 & n14681 ;
  assign n24647 = n24646 ^ n21384 ^ 1'b0 ;
  assign n24648 = n137 & ~n10303 ;
  assign n24649 = ~n348 & n24648 ;
  assign n24650 = ~n954 & n7908 ;
  assign n24651 = ~n342 & n24650 ;
  assign n24652 = n13407 | n24651 ;
  assign n24653 = ~n16385 & n24652 ;
  assign n24654 = n24649 & n24653 ;
  assign n24655 = n5793 | n13563 ;
  assign n24656 = n13874 | n24655 ;
  assign n24657 = n1017 & ~n22715 ;
  assign n24658 = n60 | n20555 ;
  assign n24659 = n24658 ^ n9006 ^ 1'b0 ;
  assign n24660 = ( n178 & ~n755 ) | ( n178 & n15679 ) | ( ~n755 & n15679 ) ;
  assign n24661 = n8370 & n15901 ;
  assign n24662 = ~n10881 & n24661 ;
  assign n24663 = n12425 ^ n9514 ^ 1'b0 ;
  assign n24664 = n10352 & n24663 ;
  assign n24665 = n4247 ^ n2538 ^ 1'b0 ;
  assign n24666 = ~n1418 & n5897 ;
  assign n24667 = n3929 ^ n2792 ^ 1'b0 ;
  assign n24668 = n4694 | n24667 ;
  assign n24669 = n227 & ~n24668 ;
  assign n24670 = n1458 & ~n24669 ;
  assign n24671 = n24670 ^ n8263 ^ 1'b0 ;
  assign n24672 = n4788 & ~n24671 ;
  assign n24673 = n8908 & n24672 ;
  assign n24674 = n24666 & n24673 ;
  assign n24675 = n5968 ^ n2834 ^ 1'b0 ;
  assign n24676 = ~n10925 & n24675 ;
  assign n24677 = n15395 & n24676 ;
  assign n24678 = n13393 & ~n24677 ;
  assign n24679 = ~n5643 & n11953 ;
  assign n24680 = ~n7472 & n17203 ;
  assign n24681 = n21586 ^ n8587 ^ 1'b0 ;
  assign n24682 = n2566 | n24681 ;
  assign n24683 = n7063 | n10255 ;
  assign n24684 = n24683 ^ n9342 ^ 1'b0 ;
  assign n24685 = n24684 ^ n4697 ^ n434 ;
  assign n24686 = ~n1421 & n15700 ;
  assign n24687 = n24686 ^ n7350 ^ 1'b0 ;
  assign n24688 = ~n21157 & n24687 ;
  assign n24689 = n24542 & n24688 ;
  assign n24690 = n5550 & ~n24689 ;
  assign n24691 = n1865 ^ n308 ^ 1'b0 ;
  assign n24692 = ~n18039 & n24691 ;
  assign n24693 = n19663 ^ n2476 ^ 1'b0 ;
  assign n24694 = n9925 | n24693 ;
  assign n24695 = n3267 & n17531 ;
  assign n24696 = n5660 | n24695 ;
  assign n24697 = n24696 ^ n12411 ^ 1'b0 ;
  assign n24698 = n51 & n727 ;
  assign n24699 = ~n17958 & n24698 ;
  assign n24700 = ~n7284 & n24699 ;
  assign n24701 = n23513 & n24700 ;
  assign n24702 = n16842 ^ n3260 ^ 1'b0 ;
  assign n24703 = n16750 | n19455 ;
  assign n24704 = n12879 | n24703 ;
  assign n24705 = n6567 | n13619 ;
  assign n24706 = ~n174 & n4582 ;
  assign n24707 = ~n7608 & n24706 ;
  assign n24708 = n4163 & n18013 ;
  assign n24709 = ~n12290 & n14667 ;
  assign n24710 = n24708 & n24709 ;
  assign n24711 = n21594 ^ n8662 ^ 1'b0 ;
  assign n24712 = n7681 ^ n5574 ^ 1'b0 ;
  assign n24713 = n7555 | n24712 ;
  assign n24714 = n5858 & n12000 ;
  assign n24715 = n24713 | n24714 ;
  assign n24716 = n6617 | n9072 ;
  assign n24717 = ( n3820 & n15098 ) | ( n3820 & ~n24716 ) | ( n15098 & ~n24716 ) ;
  assign n24718 = n23735 ^ n8788 ^ 1'b0 ;
  assign n24719 = n4097 & n24718 ;
  assign n24720 = n581 & n16347 ;
  assign n24721 = ~n3430 & n24720 ;
  assign n24722 = x5 | n338 ;
  assign n24723 = n246 & n24722 ;
  assign n24724 = n24723 ^ n8976 ^ 1'b0 ;
  assign n24725 = ~n14395 & n14789 ;
  assign n24726 = ~n8128 & n24725 ;
  assign n24727 = n24724 | n24726 ;
  assign n24728 = n8285 ^ n7676 ^ 1'b0 ;
  assign n24729 = n5227 | n24728 ;
  assign n24730 = n2477 & n6150 ;
  assign n24731 = n24730 ^ n1418 ^ 1'b0 ;
  assign n24732 = ~n21545 & n24731 ;
  assign n24733 = n20076 ^ n4129 ^ n2964 ;
  assign n24734 = n3769 & n6019 ;
  assign n24735 = ~n3769 & n24734 ;
  assign n24736 = x8 & ~n6799 ;
  assign n24737 = ~x8 & n24736 ;
  assign n24738 = n17421 | n24737 ;
  assign n24739 = n12585 & ~n24738 ;
  assign n24740 = n111 & ~n17421 ;
  assign n24741 = n17421 & n24740 ;
  assign n24742 = n24739 & ~n24741 ;
  assign n24743 = n74 | n94 ;
  assign n24744 = n74 & ~n24743 ;
  assign n24745 = n89 & ~n24744 ;
  assign n24746 = n24744 & n24745 ;
  assign n24747 = n122 & ~n24746 ;
  assign n24748 = ~n122 & n24747 ;
  assign n24749 = n9457 | n24748 ;
  assign n24750 = n24742 & ~n24749 ;
  assign n24751 = ~n24742 & n24750 ;
  assign n24752 = n15485 & ~n24751 ;
  assign n24753 = ~n15485 & n24752 ;
  assign n24754 = n24753 ^ n20719 ^ 1'b0 ;
  assign n24755 = ~n24735 & n24754 ;
  assign n24756 = n2267 | n4320 ;
  assign n24757 = n24756 ^ n5333 ^ 1'b0 ;
  assign n24759 = n21814 ^ n8220 ^ 1'b0 ;
  assign n24758 = n8529 & ~n10203 ;
  assign n24760 = n24759 ^ n24758 ^ 1'b0 ;
  assign n24761 = ~n14376 & n20951 ;
  assign n24762 = ~n8762 & n24761 ;
  assign n24763 = n24762 ^ n5131 ^ 1'b0 ;
  assign n24764 = ~n5205 & n24763 ;
  assign n24765 = ~n865 & n8090 ;
  assign n24766 = n15528 ^ n246 ^ 1'b0 ;
  assign n24767 = n16834 & ~n24766 ;
  assign n24768 = n24767 ^ n15012 ^ 1'b0 ;
  assign n24769 = n4574 ^ n678 ^ 1'b0 ;
  assign n24770 = n24769 ^ n7309 ^ 1'b0 ;
  assign n24771 = n9120 ^ n2694 ^ 1'b0 ;
  assign n24772 = n6720 | n12118 ;
  assign n24773 = n7244 | n24772 ;
  assign n24774 = n10490 & n24773 ;
  assign n24775 = ~n24771 & n24774 ;
  assign n24776 = n5451 ^ n83 ^ 1'b0 ;
  assign n24777 = n24776 ^ n7553 ^ 1'b0 ;
  assign n24778 = n532 & n7586 ;
  assign n24779 = n19490 & n24778 ;
  assign n24780 = n14943 | n24779 ;
  assign n24781 = n226 & n8646 ;
  assign n24782 = n553 & ~n16755 ;
  assign n24783 = n11114 & n24782 ;
  assign n24784 = n6487 | n12309 ;
  assign n24785 = n14564 | n24784 ;
  assign n24786 = n24784 & ~n24785 ;
  assign n24795 = ~n922 & n9864 ;
  assign n24796 = ~n498 & n18692 ;
  assign n24797 = ~n5830 & n24796 ;
  assign n24798 = ~n24795 & n24797 ;
  assign n24799 = n5350 & ~n24798 ;
  assign n24800 = n24798 & n24799 ;
  assign n24801 = ~n290 & n2376 ;
  assign n24802 = n290 & n24801 ;
  assign n24803 = n7528 ^ n4629 ^ 1'b0 ;
  assign n24804 = ~n24802 & n24803 ;
  assign n24805 = n24802 & n24804 ;
  assign n24806 = n24805 ^ n6887 ^ 1'b0 ;
  assign n24807 = n24800 & n24806 ;
  assign n24808 = ~n390 & n1064 ;
  assign n24809 = ~n1064 & n24808 ;
  assign n24810 = n633 & n24809 ;
  assign n24811 = n2983 & ~n24810 ;
  assign n24812 = n24807 | n24811 ;
  assign n24813 = n24807 & ~n24812 ;
  assign n24790 = n964 | n1020 ;
  assign n24791 = n964 & ~n24790 ;
  assign n24792 = n3774 | n24791 ;
  assign n24793 = n3774 & ~n24792 ;
  assign n24787 = ~n158 & n417 ;
  assign n24788 = n14 & n24787 ;
  assign n24789 = n17638 & ~n24788 ;
  assign n24794 = n24793 ^ n24789 ^ 1'b0 ;
  assign n24814 = n24813 ^ n24794 ^ 1'b0 ;
  assign n24815 = n24786 | n24814 ;
  assign n24823 = n21421 ^ n6073 ^ 1'b0 ;
  assign n24824 = n24823 ^ n1426 ^ n156 ;
  assign n24825 = ( n2076 & n3118 ) | ( n2076 & ~n24824 ) | ( n3118 & ~n24824 ) ;
  assign n24820 = n3669 ^ n2233 ^ 1'b0 ;
  assign n24821 = n24820 ^ n24244 ^ 1'b0 ;
  assign n24816 = n9094 ^ n2972 ^ 1'b0 ;
  assign n24817 = n3742 | n6645 ;
  assign n24818 = n24817 ^ n5206 ^ 1'b0 ;
  assign n24819 = ~n24816 & n24818 ;
  assign n24822 = n24821 ^ n24819 ^ 1'b0 ;
  assign n24826 = n24825 ^ n24822 ^ 1'b0 ;
  assign n24827 = n2822 & ~n24826 ;
  assign n24828 = n4111 | n8041 ;
  assign n24829 = n24828 ^ n9461 ^ 1'b0 ;
  assign n24830 = ( n9254 & ~n15591 ) | ( n9254 & n24829 ) | ( ~n15591 & n24829 ) ;
  assign n24831 = n16792 ^ n3527 ^ 1'b0 ;
  assign n24832 = ~n19091 & n19150 ;
  assign n24833 = n22307 & n24832 ;
  assign n24834 = n14987 & n16440 ;
  assign n24835 = n24834 ^ n2601 ^ 1'b0 ;
  assign n24838 = n6176 ^ n5399 ^ 1'b0 ;
  assign n24836 = ~n12175 & n17825 ;
  assign n24837 = n24836 ^ n8107 ^ 1'b0 ;
  assign n24839 = n24838 ^ n24837 ^ 1'b0 ;
  assign n24840 = n1388 | n3027 ;
  assign n24841 = n24840 ^ n9898 ^ 1'b0 ;
  assign n24842 = n22952 & ~n24841 ;
  assign n24843 = ~n1787 & n24842 ;
  assign n24844 = n2431 & ~n24843 ;
  assign n24845 = ~n21338 & n24844 ;
  assign n24846 = n14125 & ~n20415 ;
  assign n24847 = n15470 & n24846 ;
  assign n24848 = n15840 ^ n236 ^ 1'b0 ;
  assign n24849 = n24847 | n24848 ;
  assign n24850 = n24849 ^ n16777 ^ 1'b0 ;
  assign n24851 = n22840 ^ n2853 ^ 1'b0 ;
  assign n24852 = ~n9092 & n24851 ;
  assign n24853 = n2913 & n23566 ;
  assign n24854 = n10531 & n14142 ;
  assign n24855 = n8327 & n10107 ;
  assign n24856 = ~n24854 & n24855 ;
  assign n24857 = n10347 ^ n726 ^ 1'b0 ;
  assign n24858 = ~n20667 & n24857 ;
  assign n24859 = ~n12488 & n24858 ;
  assign n24860 = ~n10149 & n24859 ;
  assign n24861 = n24513 ^ n10990 ^ 1'b0 ;
  assign n24862 = n17854 & n24861 ;
  assign n24863 = n10273 ^ n3608 ^ 1'b0 ;
  assign n24864 = ~n119 & n24863 ;
  assign n24865 = n1449 | n5179 ;
  assign n24866 = n7532 | n22638 ;
  assign n24867 = n5144 | n24866 ;
  assign n24868 = n934 ^ n300 ^ 1'b0 ;
  assign n24869 = n24868 ^ n17976 ^ 1'b0 ;
  assign n24870 = n5377 | n21448 ;
  assign n24871 = n24870 ^ n11129 ^ 1'b0 ;
  assign n24872 = n21826 ^ n1325 ^ 1'b0 ;
  assign n24873 = n24871 & ~n24872 ;
  assign n24874 = n2577 | n14699 ;
  assign n24875 = n34 & n5892 ;
  assign n24876 = ~n2478 & n24875 ;
  assign n24877 = n2478 & n24876 ;
  assign n24878 = ( ~n20549 & n21568 ) | ( ~n20549 & n24877 ) | ( n21568 & n24877 ) ;
  assign n24879 = n16606 ^ n14854 ^ 1'b0 ;
  assign n24880 = n4931 & ~n24879 ;
  assign n24881 = n3597 & n11763 ;
  assign n24882 = n10303 & n24881 ;
  assign n24883 = n11913 ^ n1789 ^ 1'b0 ;
  assign n24884 = ~n10177 & n24883 ;
  assign n24885 = n270 & n24884 ;
  assign n24886 = n20501 ^ n5764 ^ 1'b0 ;
  assign n24888 = n1406 ^ n903 ^ n367 ;
  assign n24887 = n1818 & n17142 ;
  assign n24889 = n24888 ^ n24887 ^ 1'b0 ;
  assign n24890 = ~n3021 & n15145 ;
  assign n24891 = n22254 & ~n24890 ;
  assign n24892 = ~n4559 & n13844 ;
  assign n24893 = n24892 ^ n8916 ^ 1'b0 ;
  assign n24894 = n278 & n24893 ;
  assign n24895 = n24894 ^ n2233 ^ 1'b0 ;
  assign n24896 = n5544 & ~n8777 ;
  assign n24897 = n24896 ^ n23989 ^ 1'b0 ;
  assign n24898 = n8699 ^ n2059 ^ 1'b0 ;
  assign n24899 = n688 | n24898 ;
  assign n24900 = n21999 | n24899 ;
  assign n24901 = ~n1501 & n24261 ;
  assign n24902 = n24901 ^ n5394 ^ 1'b0 ;
  assign n24903 = n2631 & n15112 ;
  assign n24904 = n5612 ^ n4927 ^ 1'b0 ;
  assign n24905 = ~n16326 & n24904 ;
  assign n24906 = n24905 ^ n16564 ^ 1'b0 ;
  assign n24907 = n15544 ^ n9626 ^ n4332 ;
  assign n24908 = ~n24906 & n24907 ;
  assign n24909 = n18953 ^ n2449 ^ 1'b0 ;
  assign n24910 = n24909 ^ n5871 ^ 1'b0 ;
  assign n24911 = n2790 | n24910 ;
  assign n24912 = n6784 ^ n4531 ^ 1'b0 ;
  assign n24913 = n18334 & n24912 ;
  assign n24914 = n24913 ^ n7472 ^ 1'b0 ;
  assign n24915 = n17781 ^ n17194 ^ 1'b0 ;
  assign n24916 = n1958 & n24915 ;
  assign n24917 = n24916 ^ n6552 ^ 1'b0 ;
  assign n24918 = n10728 ^ n2982 ^ 1'b0 ;
  assign n24919 = n2148 | n24918 ;
  assign n24920 = n24919 ^ n4875 ^ 1'b0 ;
  assign n24921 = n11944 ^ n5823 ^ 1'b0 ;
  assign n24922 = n3579 | n11995 ;
  assign n24923 = n24921 | n24922 ;
  assign n24924 = n24923 ^ n24215 ^ 1'b0 ;
  assign n24925 = n378 & n24924 ;
  assign n24926 = n6023 ^ n3156 ^ n1159 ;
  assign n24927 = ( ~n9913 & n24925 ) | ( ~n9913 & n24926 ) | ( n24925 & n24926 ) ;
  assign n24928 = n10858 & ~n14450 ;
  assign n24929 = n1027 ^ n737 ^ 1'b0 ;
  assign n24930 = n24928 & ~n24929 ;
  assign n24931 = n24930 ^ n5161 ^ 1'b0 ;
  assign n24932 = n14970 & n22897 ;
  assign n24933 = n220 & ~n14086 ;
  assign n24934 = ~n9088 & n10398 ;
  assign n24935 = n3451 & n24934 ;
  assign n24936 = n1179 & n6265 ;
  assign n24937 = n4690 | n24936 ;
  assign n24938 = n32 & n24937 ;
  assign n24939 = n6712 & n24490 ;
  assign n24941 = n906 | n1130 ;
  assign n24942 = n906 & ~n24941 ;
  assign n24943 = ~n13096 & n24942 ;
  assign n24944 = ~n4061 & n14297 ;
  assign n24945 = n1137 | n1318 ;
  assign n24946 = n1137 & ~n24945 ;
  assign n24947 = n24944 | n24946 ;
  assign n24948 = n24944 & ~n24947 ;
  assign n24949 = n24948 ^ n19144 ^ 1'b0 ;
  assign n24950 = ~n24943 & n24949 ;
  assign n24951 = n24950 ^ n1445 ^ 1'b0 ;
  assign n24940 = n1129 & n8842 ;
  assign n24952 = n24951 ^ n24940 ^ 1'b0 ;
  assign n24953 = n1452 | n5835 ;
  assign n24954 = n235 & ~n4853 ;
  assign n24955 = x5 | n21072 ;
  assign n24956 = n24955 ^ n191 ^ 1'b0 ;
  assign n24957 = n1354 & n4604 ;
  assign n24958 = n21124 ^ n1254 ^ 1'b0 ;
  assign n24959 = n10762 & n13830 ;
  assign n24960 = n177 & n6970 ;
  assign n24961 = n24960 ^ n3269 ^ 1'b0 ;
  assign n24962 = n18219 ^ n11387 ^ 1'b0 ;
  assign n24963 = n16313 ^ n6817 ^ 1'b0 ;
  assign n24964 = n636 | n4572 ;
  assign n24965 = n16275 & ~n24964 ;
  assign n24966 = n2266 & n8551 ;
  assign n24967 = n512 & n24966 ;
  assign n24968 = n962 & n6932 ;
  assign n24969 = ~n24483 & n24968 ;
  assign n24970 = n3219 | n4191 ;
  assign n24971 = n5764 | n24970 ;
  assign n24972 = n1760 & ~n24971 ;
  assign n24973 = n9539 & ~n20365 ;
  assign n24974 = n24973 ^ n18785 ^ 1'b0 ;
  assign n24975 = n13055 & ~n24974 ;
  assign n24980 = n1777 ^ n395 ^ 1'b0 ;
  assign n24976 = n70 & ~n2171 ;
  assign n24977 = n24976 ^ n2572 ^ 1'b0 ;
  assign n24978 = n17937 ^ n2655 ^ 1'b0 ;
  assign n24979 = ~n24977 & n24978 ;
  assign n24981 = n24980 ^ n24979 ^ 1'b0 ;
  assign n24982 = n740 | n6236 ;
  assign n24983 = ~n364 & n880 ;
  assign n24984 = ~n1650 & n24983 ;
  assign n24985 = n24984 ^ n1982 ^ 1'b0 ;
  assign n24986 = n24985 ^ n5538 ^ 1'b0 ;
  assign n24987 = ~n6732 & n24986 ;
  assign n24988 = n8393 & ~n21978 ;
  assign n24989 = n14936 ^ n6364 ^ 1'b0 ;
  assign n24990 = n15198 ^ n2608 ^ 1'b0 ;
  assign n24991 = n2185 & ~n24990 ;
  assign n24992 = n10977 & n24991 ;
  assign n24993 = ~n1932 & n24992 ;
  assign n24994 = n16506 | n24993 ;
  assign n24996 = n207 & ~n2536 ;
  assign n24995 = ~n273 & n1598 ;
  assign n24997 = n24996 ^ n24995 ^ n6247 ;
  assign n24998 = n2910 | n15516 ;
  assign n24999 = n5493 ^ n4623 ^ 1'b0 ;
  assign n25000 = ~n5730 & n24999 ;
  assign n25001 = n754 | n23954 ;
  assign n25002 = n23096 ^ n15092 ^ 1'b0 ;
  assign n25003 = ~n553 & n25002 ;
  assign n25004 = ~n1842 & n5956 ;
  assign n25005 = n22114 ^ n20735 ^ 1'b0 ;
  assign n25006 = n7185 ^ n497 ^ 1'b0 ;
  assign n25007 = n6589 & n25006 ;
  assign n25008 = ~n4266 & n25007 ;
  assign n25009 = n7731 & ~n25008 ;
  assign n25010 = n12477 ^ n156 ^ 1'b0 ;
  assign n25011 = n20022 ^ n19981 ^ 1'b0 ;
  assign n25012 = n25010 & n25011 ;
  assign n25013 = n325 & n2278 ;
  assign n25014 = n22461 ^ n1227 ^ 1'b0 ;
  assign n25015 = n16990 | n25014 ;
  assign n25016 = n12242 ^ n1630 ^ 1'b0 ;
  assign n25017 = ~n1172 & n25016 ;
  assign n25018 = n3346 ^ n133 ^ 1'b0 ;
  assign n25019 = n7064 & ~n24386 ;
  assign n25020 = n25019 ^ n9627 ^ 1'b0 ;
  assign n25021 = ~n10288 & n11829 ;
  assign n25022 = ~n7130 & n25021 ;
  assign n25023 = n1010 & n25022 ;
  assign n25024 = ~n2300 & n2695 ;
  assign n25025 = n25024 ^ n3271 ^ 1'b0 ;
  assign n25026 = n10739 | n25025 ;
  assign n25027 = n1449 | n3300 ;
  assign n25028 = n37 & n25027 ;
  assign n25029 = n2064 ^ n567 ^ 1'b0 ;
  assign n25030 = n1073 & n10055 ;
  assign n25031 = n25030 ^ n1254 ^ n968 ;
  assign n25032 = n25029 | n25031 ;
  assign n25033 = n25032 ^ n7134 ^ 1'b0 ;
  assign n25034 = ~n5835 & n14579 ;
  assign n25035 = n25034 ^ n2414 ^ 1'b0 ;
  assign n25036 = n25035 ^ n2078 ^ 1'b0 ;
  assign n25037 = n1226 & ~n3437 ;
  assign n25038 = ~n6249 & n17268 ;
  assign n25039 = n17293 ^ n11433 ^ 1'b0 ;
  assign n25040 = n18302 & ~n19227 ;
  assign n25041 = n19227 & n25040 ;
  assign n25042 = n11858 | n14466 ;
  assign n25043 = n25042 ^ n12523 ^ 1'b0 ;
  assign n25044 = ~n20338 & n21639 ;
  assign n25045 = n25043 & n25044 ;
  assign n25046 = n5192 & n10137 ;
  assign n25047 = n2637 & n25046 ;
  assign n25048 = n21807 ^ n14970 ^ 1'b0 ;
  assign n25049 = n475 & ~n2864 ;
  assign n25050 = ~n8107 & n12242 ;
  assign n25051 = ~n25049 & n25050 ;
  assign n25052 = ( n5635 & ~n9885 ) | ( n5635 & n13299 ) | ( ~n9885 & n13299 ) ;
  assign n25053 = n11833 & ~n25052 ;
  assign n25054 = n17021 ^ n6487 ^ 1'b0 ;
  assign n25055 = n15052 & n25054 ;
  assign n25056 = n9059 ^ n3526 ^ 1'b0 ;
  assign n25057 = n25 | n25056 ;
  assign n25058 = n25057 ^ n8192 ^ 1'b0 ;
  assign n25059 = n7544 | n14226 ;
  assign n25060 = n5873 ^ n4791 ^ 1'b0 ;
  assign n25061 = n10590 & ~n16219 ;
  assign n25062 = n5978 ^ n5239 ^ 1'b0 ;
  assign n25063 = n17196 | n25062 ;
  assign n25064 = n15652 | n17330 ;
  assign n25065 = n25064 ^ n15859 ^ 1'b0 ;
  assign n25066 = n2759 | n22527 ;
  assign n25067 = n7764 | n10588 ;
  assign n25068 = n25067 ^ n6194 ^ 1'b0 ;
  assign n25069 = n5832 | n6720 ;
  assign n25070 = n2967 & ~n10774 ;
  assign n25071 = n25070 ^ n3983 ^ 1'b0 ;
  assign n25072 = n25069 & ~n25071 ;
  assign n25073 = n1822 & n20971 ;
  assign n25074 = ~n1169 & n4186 ;
  assign n25075 = n25074 ^ n11917 ^ 1'b0 ;
  assign n25076 = n19404 ^ n3687 ^ 1'b0 ;
  assign n25077 = n16822 ^ n4377 ^ 1'b0 ;
  assign n25078 = ~n15866 & n25077 ;
  assign n25079 = n8399 & n25078 ;
  assign n25080 = n18302 & n20095 ;
  assign n25081 = n25080 ^ n20625 ^ 1'b0 ;
  assign n25082 = n163 & n20408 ;
  assign n25083 = n8601 & n25082 ;
  assign n25084 = n24007 ^ n5880 ^ 1'b0 ;
  assign n25085 = n15216 & ~n25084 ;
  assign n25086 = n7273 ^ n1368 ^ 1'b0 ;
  assign n25087 = n12867 ^ n6702 ^ 1'b0 ;
  assign n25088 = n25086 & ~n25087 ;
  assign n25089 = n5586 & n11535 ;
  assign n25090 = n4708 & n12345 ;
  assign n25091 = n25090 ^ n3121 ^ 1'b0 ;
  assign n25092 = n25091 ^ n13891 ^ 1'b0 ;
  assign n25093 = n1664 & ~n7488 ;
  assign n25094 = n23169 & n25093 ;
  assign n25095 = n7391 & ~n25094 ;
  assign n25096 = n25095 ^ n12657 ^ 1'b0 ;
  assign n25097 = ~n6178 & n25096 ;
  assign n25098 = ~n1714 & n25097 ;
  assign n25099 = n25098 ^ n5264 ^ 1'b0 ;
  assign n25100 = n16040 ^ n12263 ^ 1'b0 ;
  assign n25101 = ~n520 & n1040 ;
  assign n25102 = ~n5760 & n25101 ;
  assign n25103 = n25102 ^ n4626 ^ 1'b0 ;
  assign n25104 = n3976 & ~n25103 ;
  assign n25105 = n412 & ~n25104 ;
  assign n25106 = n24236 ^ n13764 ^ 1'b0 ;
  assign n25107 = n2110 ^ n1631 ^ 1'b0 ;
  assign n25108 = n4331 | n25107 ;
  assign n25109 = n25108 ^ n8242 ^ 1'b0 ;
  assign n25110 = n1081 | n25109 ;
  assign n25111 = n25110 ^ n11592 ^ n7080 ;
  assign n25112 = n10477 ^ n4195 ^ 1'b0 ;
  assign n25113 = n25112 ^ n21872 ^ 1'b0 ;
  assign n25114 = n327 | n1966 ;
  assign n25115 = n5205 | n25114 ;
  assign n25116 = n25114 & ~n25115 ;
  assign n25117 = ~n7185 & n16013 ;
  assign n25118 = n25117 ^ n1329 ^ 1'b0 ;
  assign n25119 = n24356 & ~n25118 ;
  assign n25120 = n4000 & n25119 ;
  assign n25121 = n3580 & ~n3931 ;
  assign n25122 = n1070 & n25121 ;
  assign n25123 = n25122 ^ n1904 ^ 1'b0 ;
  assign n25124 = n1954 ^ n226 ^ 1'b0 ;
  assign n25125 = n178 & n25124 ;
  assign n25126 = n25125 ^ n23461 ^ 1'b0 ;
  assign n25127 = n25123 | n25126 ;
  assign n25128 = n11446 | n21389 ;
  assign n25129 = n25128 ^ n9447 ^ 1'b0 ;
  assign n25130 = n25129 ^ n7535 ^ 1'b0 ;
  assign n25131 = n8939 & n21376 ;
  assign n25132 = n5204 & n9154 ;
  assign n25133 = n2848 & n25132 ;
  assign n25134 = n827 & ~n25133 ;
  assign n25136 = n8022 | n13043 ;
  assign n25135 = n3469 | n18264 ;
  assign n25137 = n25136 ^ n25135 ^ 1'b0 ;
  assign n25138 = n6873 & ~n25137 ;
  assign n25139 = n17313 ^ n3370 ^ 1'b0 ;
  assign n25143 = n4936 ^ n2288 ^ 1'b0 ;
  assign n25140 = n4537 | n7448 ;
  assign n25141 = n14452 & ~n25140 ;
  assign n25142 = ~n3873 & n25141 ;
  assign n25144 = n25143 ^ n25142 ^ 1'b0 ;
  assign n25145 = n1966 & ~n3980 ;
  assign n25146 = ~n9234 & n25145 ;
  assign n25147 = n4780 & n6179 ;
  assign n25148 = n12898 ^ n4899 ^ 1'b0 ;
  assign n25149 = n12511 ^ n1474 ^ 1'b0 ;
  assign n25150 = n22365 & ~n25149 ;
  assign n25151 = n11826 | n25150 ;
  assign n25152 = ~n375 & n4535 ;
  assign n25153 = n7066 & n25152 ;
  assign n25154 = n25153 ^ n23269 ^ 1'b0 ;
  assign n25155 = n2975 & ~n12982 ;
  assign n25156 = ~n290 & n13614 ;
  assign n25157 = ~n22329 & n25156 ;
  assign n25158 = ~n2864 & n4769 ;
  assign n25159 = ~n713 & n25158 ;
  assign n25160 = n98 & ~n25159 ;
  assign n25161 = ~n1645 & n25160 ;
  assign n25162 = ~n9255 & n21276 ;
  assign n25163 = n25162 ^ n8151 ^ 1'b0 ;
  assign n25164 = n17545 ^ n37 ^ 1'b0 ;
  assign n25169 = n10837 & ~n19301 ;
  assign n25165 = n17016 ^ n8467 ^ 1'b0 ;
  assign n25166 = n22451 | n25165 ;
  assign n25167 = n14242 | n25166 ;
  assign n25168 = n20365 & n25167 ;
  assign n25170 = n25169 ^ n25168 ^ 1'b0 ;
  assign n25171 = n7391 ^ n4929 ^ 1'b0 ;
  assign n25172 = n6184 & ~n25171 ;
  assign n25173 = ~n3569 & n18594 ;
  assign n25174 = n1686 & n12951 ;
  assign n25175 = ~n25173 & n25174 ;
  assign n25176 = n14394 & ~n25175 ;
  assign n25177 = n22535 & n25176 ;
  assign n25179 = n2458 & n2644 ;
  assign n25178 = n299 & n731 ;
  assign n25180 = n25179 ^ n25178 ^ 1'b0 ;
  assign n25181 = n233 & ~n16444 ;
  assign n25185 = n2183 & ~n3586 ;
  assign n25186 = ~n17117 & n25185 ;
  assign n25182 = n20662 ^ x5 ^ 1'b0 ;
  assign n25183 = n20185 | n25182 ;
  assign n25184 = n8362 | n25183 ;
  assign n25187 = n25186 ^ n25184 ^ 1'b0 ;
  assign n25188 = n7710 | n25187 ;
  assign n25189 = n5520 & n9142 ;
  assign n25190 = n25189 ^ n19380 ^ 1'b0 ;
  assign n25191 = n6089 ^ n1763 ^ 1'b0 ;
  assign n25192 = n489 & n25191 ;
  assign n25193 = n3075 & ~n13121 ;
  assign n25194 = n25193 ^ n5354 ^ 1'b0 ;
  assign n25195 = n25192 | n25194 ;
  assign n25196 = n4176 & n10891 ;
  assign n25197 = n1730 | n2742 ;
  assign n25198 = n25197 ^ n158 ^ 1'b0 ;
  assign n25199 = n2191 & n25198 ;
  assign n25200 = n4543 ^ n252 ^ 1'b0 ;
  assign n25201 = n921 & n25200 ;
  assign n25202 = ~n11283 & n25201 ;
  assign n25203 = n938 & ~n5063 ;
  assign n25204 = n25203 ^ n22102 ^ 1'b0 ;
  assign n25205 = n288 & n25204 ;
  assign n25206 = n6713 & n25205 ;
  assign n25207 = n25202 & n25206 ;
  assign n25208 = n7675 & ~n9763 ;
  assign n25209 = ~n330 & n25208 ;
  assign n25211 = n3311 & n6603 ;
  assign n25210 = n788 & n2809 ;
  assign n25212 = n25211 ^ n25210 ^ 1'b0 ;
  assign n25213 = n25212 ^ n888 ^ 1'b0 ;
  assign n25214 = n477 & ~n25213 ;
  assign n25215 = n25214 ^ n2553 ^ n1390 ;
  assign n25216 = ~n6658 & n17652 ;
  assign n25217 = n951 ^ n241 ^ 1'b0 ;
  assign n25218 = ~n164 & n694 ;
  assign n25219 = n4406 & ~n25218 ;
  assign n25220 = n5111 & n25219 ;
  assign n25221 = n14961 & n21085 ;
  assign n25222 = n8539 & n25221 ;
  assign n25223 = n5218 | n10279 ;
  assign n25224 = n24516 & ~n25223 ;
  assign n25225 = ~n24116 & n25224 ;
  assign n25226 = n2036 ^ n346 ^ 1'b0 ;
  assign n25227 = n5978 | n25226 ;
  assign n25228 = n6817 & ~n25227 ;
  assign n25229 = ~n14046 & n25228 ;
  assign n25230 = n8928 ^ n4749 ^ 1'b0 ;
  assign n25231 = n15233 & n21164 ;
  assign n25232 = n25230 & n25231 ;
  assign n25233 = n8134 | n25232 ;
  assign n25234 = n1802 ^ n898 ^ 1'b0 ;
  assign n25235 = ~n5355 & n15522 ;
  assign n25236 = n7812 ^ n3511 ^ 1'b0 ;
  assign n25237 = n2964 & n15455 ;
  assign n25238 = n4451 ^ n616 ^ 1'b0 ;
  assign n25239 = n19076 & n25238 ;
  assign n25240 = n24 & ~n15060 ;
  assign n25241 = n25240 ^ n13854 ^ 1'b0 ;
  assign n25242 = ~n4121 & n10447 ;
  assign n25243 = n3552 | n13574 ;
  assign n25244 = n25243 ^ n10774 ^ n7805 ;
  assign n25245 = n330 & ~n3877 ;
  assign n25246 = n25245 ^ n6361 ^ 1'b0 ;
  assign n25247 = ~n10925 & n25246 ;
  assign n25248 = n6764 & n12442 ;
  assign n25249 = ~n11868 & n25248 ;
  assign n25250 = n24606 ^ n1379 ^ 1'b0 ;
  assign n25251 = ~n5691 & n25250 ;
  assign n25252 = n25251 ^ n7904 ^ 1'b0 ;
  assign n25254 = n4076 & n10651 ;
  assign n25255 = n25254 ^ n23819 ^ 1'b0 ;
  assign n25253 = n763 & n20280 ;
  assign n25256 = n25255 ^ n25253 ^ 1'b0 ;
  assign n25257 = n10100 | n20415 ;
  assign n25258 = n23619 & ~n25257 ;
  assign n25259 = n9498 & ~n19224 ;
  assign n25260 = ~n364 & n25259 ;
  assign n25261 = n19460 & ~n25260 ;
  assign n25262 = n25258 & n25261 ;
  assign n25263 = n101 | n25262 ;
  assign n25264 = n17876 ^ n9062 ^ n768 ;
  assign n25265 = n436 | n25264 ;
  assign n25266 = n25265 ^ n23864 ^ 1'b0 ;
  assign n25267 = n22159 & ~n25266 ;
  assign n25268 = n14226 ^ n2751 ^ 1'b0 ;
  assign n25269 = ~n234 & n25268 ;
  assign n25270 = n7384 ^ n324 ^ 1'b0 ;
  assign n25271 = n14936 | n25270 ;
  assign n25272 = n6463 & n6669 ;
  assign n25273 = n1152 & n4024 ;
  assign n25274 = n25273 ^ n5583 ^ 1'b0 ;
  assign n25275 = n17211 & n22329 ;
  assign n25276 = ~n25274 & n25275 ;
  assign n25277 = n3352 | n25276 ;
  assign n25278 = n719 & ~n19562 ;
  assign n25279 = n25278 ^ n6487 ^ 1'b0 ;
  assign n25280 = ( n11462 & n17182 ) | ( n11462 & ~n25279 ) | ( n17182 & ~n25279 ) ;
  assign n25281 = ~n9065 & n19725 ;
  assign n25282 = ~n13869 & n25281 ;
  assign n25283 = n25282 ^ n4150 ^ 1'b0 ;
  assign n25284 = ~n144 & n2034 ;
  assign n25285 = n25284 ^ n3851 ^ 1'b0 ;
  assign n25286 = n3300 & ~n17812 ;
  assign n25287 = n6172 & n25286 ;
  assign n25288 = n4400 & n15192 ;
  assign n25289 = n9130 & n13964 ;
  assign n25290 = n3346 & ~n15870 ;
  assign n25291 = n19485 ^ n5856 ^ 1'b0 ;
  assign n25292 = n24096 ^ n281 ^ 1'b0 ;
  assign n25293 = n25291 & n25292 ;
  assign n25295 = n11061 ^ n3007 ^ 1'b0 ;
  assign n25296 = n3434 | n25295 ;
  assign n25294 = n5030 & ~n17169 ;
  assign n25297 = n25296 ^ n25294 ^ 1'b0 ;
  assign n25298 = n7528 ^ n4667 ^ 1'b0 ;
  assign n25299 = n6876 & n7263 ;
  assign n25300 = n25299 ^ n16589 ^ 1'b0 ;
  assign n25301 = ~n3793 & n13820 ;
  assign n25302 = n25301 ^ n11376 ^ 1'b0 ;
  assign n25303 = n1083 & ~n18627 ;
  assign n25304 = n2460 & ~n13171 ;
  assign n25305 = ~n1438 & n14531 ;
  assign n25306 = n1541 & n4949 ;
  assign n25307 = n23689 & n25306 ;
  assign n25308 = n25305 & ~n25307 ;
  assign n25309 = n25308 ^ n769 ^ 1'b0 ;
  assign n25310 = ~n9903 & n25309 ;
  assign n25311 = n802 | n22230 ;
  assign n25312 = n25311 ^ n9435 ^ 1'b0 ;
  assign n25313 = ~n43 & n25312 ;
  assign n25314 = n2064 & n25313 ;
  assign n25315 = n8523 & n23451 ;
  assign n25316 = n1216 & ~n8183 ;
  assign n25317 = n3210 & ~n9366 ;
  assign n25318 = n25317 ^ n3707 ^ 1'b0 ;
  assign n25319 = n2910 | n3935 ;
  assign n25320 = n25319 ^ n3371 ^ 1'b0 ;
  assign n25321 = n10662 ^ n8503 ^ 1'b0 ;
  assign n25322 = n1473 | n3502 ;
  assign n25323 = n25322 ^ n21510 ^ 1'b0 ;
  assign n25324 = n19672 & ~n25323 ;
  assign n25325 = n2236 & n25324 ;
  assign n25326 = n415 | n9639 ;
  assign n25327 = n18492 & n25326 ;
  assign n25328 = n24725 ^ n17931 ^ 1'b0 ;
  assign n25329 = n5160 | n25328 ;
  assign n25330 = n11021 ^ n5555 ^ 1'b0 ;
  assign n25331 = n4180 & ~n9476 ;
  assign n25332 = n14848 & n25331 ;
  assign n25333 = ~n3564 & n25332 ;
  assign n25335 = n20511 & n20805 ;
  assign n25334 = n17530 & ~n17685 ;
  assign n25336 = n25335 ^ n25334 ^ 1'b0 ;
  assign n25337 = ~n754 & n2386 ;
  assign n25338 = n3583 & ~n25337 ;
  assign n25339 = n1961 & n10785 ;
  assign n25340 = ~n2092 & n25339 ;
  assign n25341 = n3718 & n15166 ;
  assign n25342 = n5466 ^ n4791 ^ 1'b0 ;
  assign n25343 = ~n23952 & n25342 ;
  assign n25344 = n4677 & n9195 ;
  assign n25345 = n7225 & n12683 ;
  assign n25346 = ~n10046 & n25345 ;
  assign n25348 = n9234 & ~n10673 ;
  assign n25347 = n8466 | n10392 ;
  assign n25349 = n25348 ^ n25347 ^ 1'b0 ;
  assign n25350 = n622 & ~n12507 ;
  assign n25351 = ~n8049 & n13970 ;
  assign n25352 = n25351 ^ n17252 ^ 1'b0 ;
  assign n25353 = ~n3523 & n9645 ;
  assign n25354 = n25353 ^ n3396 ^ 1'b0 ;
  assign n25355 = n8995 ^ n7498 ^ 1'b0 ;
  assign n25356 = n3992 & ~n25355 ;
  assign n25357 = n18317 ^ n2087 ^ 1'b0 ;
  assign n25358 = n5836 | n25357 ;
  assign n25359 = n25358 ^ n22950 ^ 1'b0 ;
  assign n25360 = n25356 & ~n25359 ;
  assign n25361 = n553 & n9910 ;
  assign n25362 = n309 & n25361 ;
  assign n25363 = n25362 ^ n5054 ^ 1'b0 ;
  assign n25364 = n921 & ~n25363 ;
  assign n25365 = n3646 | n15866 ;
  assign n25366 = n1622 & ~n25365 ;
  assign n25367 = n15785 & ~n25366 ;
  assign n25368 = n25367 ^ n2964 ^ 1'b0 ;
  assign n25369 = n11465 & ~n16677 ;
  assign n25370 = n25369 ^ n1772 ^ 1'b0 ;
  assign n25371 = n18458 | n25370 ;
  assign n25372 = n1480 & ~n25371 ;
  assign n25373 = n25372 ^ n1668 ^ 1'b0 ;
  assign n25374 = n653 & n13411 ;
  assign n25375 = n25374 ^ n38 ^ 1'b0 ;
  assign n25376 = n8414 & ~n25375 ;
  assign n25377 = n15981 ^ n6541 ^ 1'b0 ;
  assign n25378 = n3185 & ~n15292 ;
  assign n25379 = n11681 ^ n2619 ^ 1'b0 ;
  assign n25380 = n765 & n11694 ;
  assign n25387 = n6655 | n9302 ;
  assign n25382 = ~n9088 & n20652 ;
  assign n25383 = n25382 ^ n14701 ^ 1'b0 ;
  assign n25384 = n279 & n25383 ;
  assign n25385 = n25384 ^ n3025 ^ n2497 ;
  assign n25386 = ~n12362 & n25385 ;
  assign n25388 = n25387 ^ n25386 ^ 1'b0 ;
  assign n25389 = n25388 ^ n364 ^ 1'b0 ;
  assign n25381 = n4318 & n18433 ;
  assign n25390 = n25389 ^ n25381 ^ 1'b0 ;
  assign n25397 = n294 & ~n5471 ;
  assign n25394 = n2655 | n6303 ;
  assign n25391 = ~n11756 & n18650 ;
  assign n25392 = ~n1814 & n25391 ;
  assign n25393 = n21450 | n25392 ;
  assign n25395 = n25394 ^ n25393 ^ 1'b0 ;
  assign n25396 = n3138 & n25395 ;
  assign n25398 = n25397 ^ n25396 ^ 1'b0 ;
  assign n25399 = n983 | n7108 ;
  assign n25401 = n460 & ~n14790 ;
  assign n25402 = ~n14703 & n25401 ;
  assign n25400 = n310 & n5709 ;
  assign n25403 = n25402 ^ n25400 ^ 1'b0 ;
  assign n25404 = ~n116 & n23684 ;
  assign n25405 = ~n7798 & n13798 ;
  assign n25406 = n25405 ^ n11087 ^ 1'b0 ;
  assign n25407 = n8065 ^ n6764 ^ n4662 ;
  assign n25408 = ( n7225 & ~n11552 ) | ( n7225 & n25407 ) | ( ~n11552 & n25407 ) ;
  assign n25409 = ~n25406 & n25408 ;
  assign n25411 = ~n3303 & n8370 ;
  assign n25412 = n18861 & n25411 ;
  assign n25410 = n7217 ^ n5303 ^ n3557 ;
  assign n25413 = n25412 ^ n25410 ^ 1'b0 ;
  assign n25414 = n3386 ^ n55 ^ 1'b0 ;
  assign n25415 = ~n23814 & n24149 ;
  assign n25416 = n8552 ^ n6810 ^ 1'b0 ;
  assign n25417 = n16459 | n25416 ;
  assign n25418 = n25417 ^ n19910 ^ 1'b0 ;
  assign n25419 = n23972 & n25418 ;
  assign n25420 = n11745 ^ n6577 ^ n4531 ;
  assign n25421 = n25420 ^ n10029 ^ 1'b0 ;
  assign n25422 = n2322 ^ n1396 ^ 1'b0 ;
  assign n25423 = ~n12385 & n25422 ;
  assign n25424 = ~n2183 & n25423 ;
  assign n25425 = ~n4929 & n5844 ;
  assign n25426 = n25425 ^ n22110 ^ 1'b0 ;
  assign n25427 = n14712 ^ n3899 ^ 1'b0 ;
  assign n25428 = n22614 ^ n9359 ^ 1'b0 ;
  assign n25429 = ~n17238 & n25428 ;
  assign n25430 = n5205 ^ n4759 ^ 1'b0 ;
  assign n25431 = n8765 | n25430 ;
  assign n25432 = n1966 | n5857 ;
  assign n25433 = ~n1812 & n11658 ;
  assign n25434 = n18782 & n25433 ;
  assign n25435 = n19747 ^ n11035 ^ 1'b0 ;
  assign n25436 = n15485 & ~n25435 ;
  assign n25437 = n8224 & ~n13913 ;
  assign n25438 = n4422 & n25437 ;
  assign n25439 = n2032 & n8705 ;
  assign n25440 = ~n23039 & n25439 ;
  assign n25441 = ~n20652 & n25440 ;
  assign n25445 = n4439 ^ n1335 ^ 1'b0 ;
  assign n25446 = n5261 & ~n25445 ;
  assign n25442 = n4586 | n13583 ;
  assign n25443 = n25442 ^ n14172 ^ 1'b0 ;
  assign n25444 = ( n3684 & n9357 ) | ( n3684 & n25443 ) | ( n9357 & n25443 ) ;
  assign n25447 = n25446 ^ n25444 ^ 1'b0 ;
  assign n25448 = n18818 ^ n17439 ^ 1'b0 ;
  assign n25449 = n6903 & ~n11471 ;
  assign n25450 = n22234 & n25449 ;
  assign n25451 = ~n146 & n19358 ;
  assign n25452 = ~n16660 & n25451 ;
  assign n25453 = n3841 ^ n1311 ^ 1'b0 ;
  assign n25454 = n22423 ^ n21085 ^ 1'b0 ;
  assign n25455 = n382 | n16264 ;
  assign n25456 = n2956 | n6716 ;
  assign n25457 = n25456 ^ n5048 ^ 1'b0 ;
  assign n25458 = n25457 ^ n25337 ^ 1'b0 ;
  assign n25459 = n5716 & n10107 ;
  assign n25460 = ~n128 & n25459 ;
  assign n25461 = n1392 | n25460 ;
  assign n25462 = n15196 | n25461 ;
  assign n25464 = n5771 ^ n5201 ^ 1'b0 ;
  assign n25463 = n2624 & ~n17750 ;
  assign n25465 = n25464 ^ n25463 ^ 1'b0 ;
  assign n25466 = n9620 ^ n2176 ^ 1'b0 ;
  assign n25467 = ~n3122 & n25466 ;
  assign n25468 = ~n4098 & n23484 ;
  assign n25469 = ~n25467 & n25468 ;
  assign n25470 = n11539 ^ n2281 ^ 1'b0 ;
  assign n25471 = n19161 ^ n10589 ^ 1'b0 ;
  assign n25472 = n8366 ^ n7888 ^ 1'b0 ;
  assign n25473 = n25472 ^ n293 ^ 1'b0 ;
  assign n25474 = n512 & ~n4392 ;
  assign n25475 = ~n25473 & n25474 ;
  assign n25476 = n25473 & n25475 ;
  assign n25477 = n697 & ~n25476 ;
  assign n25478 = n25476 & n25477 ;
  assign n25479 = n4053 & n16344 ;
  assign n25480 = ~n14306 & n25479 ;
  assign n25481 = n3749 ^ n1695 ^ 1'b0 ;
  assign n25482 = n25481 ^ n5643 ^ 1'b0 ;
  assign n25483 = n9275 & ~n25482 ;
  assign n25484 = n9247 | n13906 ;
  assign n25485 = n11897 | n18156 ;
  assign n25486 = n25485 ^ n5455 ^ 1'b0 ;
  assign n25487 = n688 ^ n228 ^ 1'b0 ;
  assign n25488 = n10477 & ~n25487 ;
  assign n25489 = n20263 ^ n13896 ^ 1'b0 ;
  assign n25490 = n23098 ^ n7360 ^ 1'b0 ;
  assign n25491 = ~n81 & n15154 ;
  assign n25492 = n25491 ^ n20399 ^ 1'b0 ;
  assign n25493 = n10430 & ~n25492 ;
  assign n25494 = ~n4574 & n10632 ;
  assign n25495 = n18652 ^ n284 ^ 1'b0 ;
  assign n25496 = n25337 & n25495 ;
  assign n25497 = n25496 ^ n16052 ^ 1'b0 ;
  assign n25498 = ~n6172 & n6191 ;
  assign n25499 = n764 & n25498 ;
  assign n25501 = n321 & n5452 ;
  assign n25500 = n1766 | n22432 ;
  assign n25502 = n25501 ^ n25500 ^ 1'b0 ;
  assign n25503 = n15276 & n23354 ;
  assign n25504 = n5386 | n14713 ;
  assign n25505 = n4746 | n25504 ;
  assign n25506 = ~n328 & n25505 ;
  assign n25507 = ~n9255 & n25506 ;
  assign n25508 = n5827 ^ n2951 ^ 1'b0 ;
  assign n25509 = ~n119 & n25508 ;
  assign n25510 = n6375 & ~n6749 ;
  assign n25511 = n25510 ^ n5206 ^ 1'b0 ;
  assign n25513 = n11711 ^ n8389 ^ 1'b0 ;
  assign n25512 = n1098 & n3915 ;
  assign n25514 = n25513 ^ n25512 ^ 1'b0 ;
  assign n25515 = n1447 & ~n8958 ;
  assign n25516 = n23197 ^ n5630 ^ 1'b0 ;
  assign n25517 = n25515 | n25516 ;
  assign n25518 = ~n7233 & n19178 ;
  assign n25519 = ~n1763 & n25518 ;
  assign n25520 = n2092 & ~n6823 ;
  assign n25521 = n25520 ^ n13063 ^ 1'b0 ;
  assign n25522 = n17235 ^ n11042 ^ 1'b0 ;
  assign n25523 = ~n6487 & n25522 ;
  assign n25532 = n776 & n4045 ;
  assign n25533 = n3204 & n25532 ;
  assign n25534 = n83 | n3346 ;
  assign n25535 = n6711 | n25534 ;
  assign n25536 = ~n6521 & n25535 ;
  assign n25537 = n25533 & n25536 ;
  assign n25538 = n25537 ^ n13470 ^ 1'b0 ;
  assign n25526 = n2642 & n3187 ;
  assign n25527 = n908 | n25526 ;
  assign n25528 = n3757 | n5495 ;
  assign n25529 = n25527 | n25528 ;
  assign n25524 = n130 & ~n5691 ;
  assign n25525 = ~n11641 & n25524 ;
  assign n25530 = n25529 ^ n25525 ^ 1'b0 ;
  assign n25531 = n22044 | n25530 ;
  assign n25539 = n25538 ^ n25531 ^ 1'b0 ;
  assign n25540 = n291 & ~n15210 ;
  assign n25541 = n14258 ^ n7237 ^ 1'b0 ;
  assign n25542 = n6055 ^ n1179 ^ 1'b0 ;
  assign n25543 = n8170 ^ n666 ^ 1'b0 ;
  assign n25544 = n280 | n1001 ;
  assign n25545 = n25544 ^ n23871 ^ 1'b0 ;
  assign n25546 = n11067 | n20197 ;
  assign n25547 = n25546 ^ n815 ^ 1'b0 ;
  assign n25548 = ~n16313 & n25547 ;
  assign n25549 = n14046 & ~n24544 ;
  assign n25550 = n787 & n6617 ;
  assign n25551 = n8572 & n25550 ;
  assign n25552 = n25551 ^ n8614 ^ 1'b0 ;
  assign n25553 = ~n10670 & n14143 ;
  assign n25554 = n19327 ^ n12388 ^ n4740 ;
  assign n25555 = n25553 & ~n25554 ;
  assign n25556 = n15173 ^ n2672 ^ 1'b0 ;
  assign n25557 = n9486 & n25556 ;
  assign n25558 = n5613 & n12089 ;
  assign n25559 = n52 & n4334 ;
  assign n25560 = n8319 & n25559 ;
  assign n25561 = n25560 ^ n330 ^ 1'b0 ;
  assign n25562 = n9152 & n25561 ;
  assign n25563 = n24231 ^ n1179 ^ 1'b0 ;
  assign n25564 = n3171 ^ n1193 ^ 1'b0 ;
  assign n25565 = n25564 ^ n7271 ^ 1'b0 ;
  assign n25566 = ~n243 & n25565 ;
  assign n25567 = n25566 ^ n22669 ^ n2964 ;
  assign n25568 = n9126 & ~n25567 ;
  assign n25569 = n3472 & ~n9048 ;
  assign n25570 = n25569 ^ n9201 ^ 1'b0 ;
  assign n25571 = n6971 | n7056 ;
  assign n25572 = n1254 | n25571 ;
  assign n25573 = n4788 & ~n5794 ;
  assign n25574 = n25573 ^ n3616 ^ 1'b0 ;
  assign n25575 = n25574 ^ n20807 ^ 1'b0 ;
  assign n25576 = ( n958 & n8750 ) | ( n958 & ~n21117 ) | ( n8750 & ~n21117 ) ;
  assign n25577 = n25576 ^ n7888 ^ 1'b0 ;
  assign n25578 = n3269 & ~n17882 ;
  assign n25579 = ~n330 & n25578 ;
  assign n25580 = n5793 | n17183 ;
  assign n25581 = n1011 | n4483 ;
  assign n25582 = n2937 ^ n2047 ^ n1355 ;
  assign n25583 = n9601 & ~n25582 ;
  assign n25584 = n25583 ^ n25055 ^ 1'b0 ;
  assign n25585 = ~n9377 & n25584 ;
  assign n25586 = n20339 ^ n18271 ^ 1'b0 ;
  assign n25587 = ~n19068 & n25586 ;
  assign n25588 = n2267 | n18624 ;
  assign n25589 = n25588 ^ n1283 ^ 1'b0 ;
  assign n25590 = n9096 ^ n3743 ^ 1'b0 ;
  assign n25591 = n8258 & n25590 ;
  assign n25592 = n9447 | n25591 ;
  assign n25593 = ~n950 & n22130 ;
  assign n25594 = n4203 & n7009 ;
  assign n25596 = n79 & ~n24172 ;
  assign n25595 = n7455 & ~n12412 ;
  assign n25597 = n25596 ^ n25595 ^ 1'b0 ;
  assign n25598 = n19383 ^ n6933 ^ 1'b0 ;
  assign n25599 = n23496 ^ n9789 ^ 1'b0 ;
  assign n25600 = ~n11487 & n25599 ;
  assign n25601 = ~n12795 & n25281 ;
  assign n25602 = n2626 & n25601 ;
  assign n25603 = n18970 ^ n1842 ^ 1'b0 ;
  assign n25604 = n17483 & n25603 ;
  assign n25605 = ~n423 & n25604 ;
  assign n25606 = n10924 | n22282 ;
  assign n25607 = n3329 & n13186 ;
  assign n25610 = n16418 ^ n2320 ^ 1'b0 ;
  assign n25608 = n2148 & n14310 ;
  assign n25609 = ~n21521 & n25608 ;
  assign n25611 = n25610 ^ n25609 ^ n16041 ;
  assign n25612 = n452 & ~n25611 ;
  assign n25613 = n8050 & ~n9551 ;
  assign n25614 = n5522 & n25613 ;
  assign n25615 = n14369 ^ n5245 ^ 1'b0 ;
  assign n25616 = n25614 & ~n25615 ;
  assign n25617 = n6272 ^ n4361 ^ 1'b0 ;
  assign n25618 = n520 | n9747 ;
  assign n25619 = n1933 | n25618 ;
  assign n25620 = n25291 ^ n18812 ^ 1'b0 ;
  assign n25621 = n4258 & n9284 ;
  assign n25622 = n8319 & n25621 ;
  assign n25623 = ~n7439 & n10971 ;
  assign n25624 = n25622 & n25623 ;
  assign n25625 = n11968 ^ n741 ^ 1'b0 ;
  assign n25626 = n5466 ^ n2364 ^ 1'b0 ;
  assign n25627 = n14194 ^ n9514 ^ 1'b0 ;
  assign n25628 = n975 & ~n25627 ;
  assign n25629 = n294 & n6907 ;
  assign n25630 = n25629 ^ n7698 ^ 1'b0 ;
  assign n25631 = ~n14400 & n25630 ;
  assign n25632 = ~n17752 & n25631 ;
  assign n25633 = n2948 | n6609 ;
  assign n25634 = ( n1963 & n19364 ) | ( n1963 & ~n25633 ) | ( n19364 & ~n25633 ) ;
  assign n25635 = n25634 ^ n12412 ^ 1'b0 ;
  assign n25636 = n2767 | n5545 ;
  assign n25637 = n51 & n8294 ;
  assign n25638 = n25637 ^ n2172 ^ 1'b0 ;
  assign n25639 = n10288 ^ n9578 ^ 1'b0 ;
  assign n25640 = n8401 & n25639 ;
  assign n25641 = n7227 ^ n2812 ^ 1'b0 ;
  assign n25642 = n17525 & n25641 ;
  assign n25643 = n21140 ^ n2817 ^ 1'b0 ;
  assign n25644 = n19048 & ~n25643 ;
  assign n25645 = n545 & ~n11570 ;
  assign n25646 = n5406 | n11922 ;
  assign n25647 = n16265 | n25646 ;
  assign n25648 = n17621 ^ n3684 ^ 1'b0 ;
  assign n25649 = n5823 & ~n25648 ;
  assign n25650 = n16813 ^ n7034 ^ 1'b0 ;
  assign n25651 = n25649 & n25650 ;
  assign n25652 = n2145 & ~n5155 ;
  assign n25653 = n5590 & n21884 ;
  assign n25654 = n25653 ^ n5135 ^ 1'b0 ;
  assign n25655 = n25652 | n25654 ;
  assign n25656 = n4087 & ~n25655 ;
  assign n25657 = n2289 & ~n19099 ;
  assign n25658 = ~n609 & n15321 ;
  assign n25659 = ~n83 & n1684 ;
  assign n25660 = n3312 | n4098 ;
  assign n25661 = n25659 & n25660 ;
  assign n25662 = n2486 & ~n12958 ;
  assign n25663 = n25662 ^ n23780 ^ 1'b0 ;
  assign n25664 = n3748 | n13334 ;
  assign n25665 = n25663 | n25664 ;
  assign n25666 = n4748 ^ n3017 ^ 1'b0 ;
  assign n25667 = n10288 & ~n16342 ;
  assign n25668 = n5880 & ~n25667 ;
  assign n25669 = n3746 & n9102 ;
  assign n25670 = n1743 & n25669 ;
  assign n25671 = ( n4927 & n17834 ) | ( n4927 & ~n25670 ) | ( n17834 & ~n25670 ) ;
  assign n25672 = ~n3542 & n10099 ;
  assign n25673 = ~n876 & n25672 ;
  assign n25674 = n5700 ^ n1003 ^ 1'b0 ;
  assign n25675 = n2546 & n25674 ;
  assign n25676 = n25675 ^ n6045 ^ 1'b0 ;
  assign n25677 = n3217 & n3552 ;
  assign n25678 = n25677 ^ n6468 ^ 1'b0 ;
  assign n25679 = n15438 & ~n15627 ;
  assign n25680 = n8930 ^ n8876 ^ 1'b0 ;
  assign n25681 = n616 & ~n1796 ;
  assign n25682 = ~n15672 & n25681 ;
  assign n25683 = ~n2813 & n15146 ;
  assign n25684 = ~n533 & n6763 ;
  assign n25685 = n25684 ^ n7483 ^ 1'b0 ;
  assign n25686 = n4785 & ~n12242 ;
  assign n25688 = n7080 & ~n11742 ;
  assign n25689 = n25688 ^ n6277 ^ 1'b0 ;
  assign n25687 = ~n4165 & n10909 ;
  assign n25690 = n25689 ^ n25687 ^ 1'b0 ;
  assign n25691 = n23062 ^ n4377 ^ 1'b0 ;
  assign n25693 = ~n954 & n15961 ;
  assign n25692 = n3061 & n20830 ;
  assign n25694 = n25693 ^ n25692 ^ 1'b0 ;
  assign n25695 = n2933 | n25694 ;
  assign n25696 = n16387 ^ n4033 ^ 1'b0 ;
  assign n25697 = ~n7439 & n25696 ;
  assign n25698 = n142 | n25697 ;
  assign n25699 = ~n16681 & n18521 ;
  assign n25700 = n1708 ^ n776 ^ 1'b0 ;
  assign n25701 = ~n22531 & n25700 ;
  assign n25702 = n25701 ^ n11590 ^ 1'b0 ;
  assign n25703 = n616 | n25702 ;
  assign n25704 = n798 & n9857 ;
  assign n25705 = n25704 ^ n21369 ^ 1'b0 ;
  assign n25706 = n1019 & ~n25705 ;
  assign n25707 = n25706 ^ n23753 ^ 1'b0 ;
  assign n25708 = n3566 ^ n984 ^ 1'b0 ;
  assign n25709 = ~n10171 & n20248 ;
  assign n25710 = n6643 & ~n12857 ;
  assign n25711 = ~n484 & n25710 ;
  assign n25712 = n2799 & ~n12669 ;
  assign n25713 = n25712 ^ n4311 ^ 1'b0 ;
  assign n25714 = n24449 ^ n2751 ^ 1'b0 ;
  assign n25715 = n25713 | n25714 ;
  assign n25716 = n2136 | n7646 ;
  assign n25717 = n24356 & ~n25716 ;
  assign n25718 = n4412 & n22867 ;
  assign n25719 = n3359 & ~n7612 ;
  assign n25720 = n8399 & ~n10009 ;
  assign n25721 = n8042 & n25720 ;
  assign n25722 = n2551 | n8203 ;
  assign n25723 = n20546 ^ n9722 ^ 1'b0 ;
  assign n25724 = ~n25722 & n25723 ;
  assign n25725 = n12064 ^ n4732 ^ 1'b0 ;
  assign n25726 = n3903 ^ n757 ^ 1'b0 ;
  assign n25727 = n18646 | n25726 ;
  assign n25728 = n25727 ^ n15821 ^ 1'b0 ;
  assign n25729 = n10926 | n25728 ;
  assign n25730 = n4891 & ~n8995 ;
  assign n25731 = n7061 & n22122 ;
  assign n25732 = n1152 & ~n24977 ;
  assign n25733 = n24977 & n25732 ;
  assign n25734 = n6245 ^ n4389 ^ 1'b0 ;
  assign n25735 = n1902 | n2626 ;
  assign n25736 = n2626 & ~n25735 ;
  assign n25737 = n1690 | n25736 ;
  assign n25738 = ( n18095 & n25734 ) | ( n18095 & n25737 ) | ( n25734 & n25737 ) ;
  assign n25739 = n25738 ^ n11438 ^ 1'b0 ;
  assign n25740 = ~n25733 & n25739 ;
  assign n25741 = ~n556 & n5842 ;
  assign n25742 = n24726 & n25741 ;
  assign n25743 = n9507 | n20676 ;
  assign n25744 = n25743 ^ n2236 ^ 1'b0 ;
  assign n25745 = n19066 ^ n18663 ^ 1'b0 ;
  assign n25746 = n3957 ^ n157 ^ 1'b0 ;
  assign n25747 = n25746 ^ n18382 ^ n10277 ;
  assign n25748 = ~n9983 & n20652 ;
  assign n25749 = n5033 & n25748 ;
  assign n25750 = n11842 & ~n25749 ;
  assign n25751 = n6903 ^ x2 ^ 1'b0 ;
  assign n25752 = n7483 | n25751 ;
  assign n25753 = n8104 & ~n25752 ;
  assign n25754 = n4915 | n6698 ;
  assign n25755 = ~n14901 & n17892 ;
  assign n25756 = n13550 ^ n1020 ^ 1'b0 ;
  assign n25757 = n23743 & n25756 ;
  assign n25758 = ~n6552 & n24040 ;
  assign n25759 = ( n169 & n1364 ) | ( n169 & n9914 ) | ( n1364 & n9914 ) ;
  assign n25760 = ~n2828 & n4122 ;
  assign n25761 = n2025 & n22815 ;
  assign n25762 = n5613 & ~n18388 ;
  assign n25763 = n25762 ^ n20095 ^ 1'b0 ;
  assign n25764 = n278 | n25763 ;
  assign n25765 = ~n11204 & n25764 ;
  assign n25766 = n25765 ^ n10602 ^ 1'b0 ;
  assign n25767 = n25766 ^ n18329 ^ n2987 ;
  assign n25768 = ( n235 & n9718 ) | ( n235 & n25767 ) | ( n9718 & n25767 ) ;
  assign n25769 = n2361 & ~n11426 ;
  assign n25770 = n11175 ^ n1593 ^ 1'b0 ;
  assign n25771 = n393 & n25770 ;
  assign n25775 = ~n7303 & n15429 ;
  assign n25776 = n25775 ^ n3015 ^ 1'b0 ;
  assign n25772 = n20060 | n21091 ;
  assign n25773 = n25772 ^ n8756 ^ 1'b0 ;
  assign n25774 = ~n2917 & n25773 ;
  assign n25777 = n25776 ^ n25774 ^ 1'b0 ;
  assign n25779 = n9913 ^ n2911 ^ 1'b0 ;
  assign n25780 = n6414 | n25779 ;
  assign n25781 = n16283 | n25780 ;
  assign n25782 = n25781 ^ n5321 ^ 1'b0 ;
  assign n25778 = n2112 & ~n11164 ;
  assign n25783 = n25782 ^ n25778 ^ 1'b0 ;
  assign n25784 = n25783 ^ n3793 ^ 1'b0 ;
  assign n25785 = n1502 & n8648 ;
  assign n25786 = n10422 ^ n8629 ^ 1'b0 ;
  assign n25787 = n13793 | n23225 ;
  assign n25788 = n12095 ^ n4044 ^ 1'b0 ;
  assign n25789 = n21395 | n24633 ;
  assign n25790 = n2767 & ~n25789 ;
  assign n25791 = n25788 | n25790 ;
  assign n25792 = n25791 ^ n21353 ^ 1'b0 ;
  assign n25793 = n3138 & ~n5698 ;
  assign n25794 = n15 & ~n25793 ;
  assign n25795 = n51 & n1368 ;
  assign n25796 = ~n7103 & n10510 ;
  assign n25797 = n17617 ^ n940 ^ 1'b0 ;
  assign n25798 = n25796 & ~n25797 ;
  assign n25799 = n2879 & ~n3138 ;
  assign n25800 = n9975 ^ n962 ^ n609 ;
  assign n25801 = n25800 ^ n7458 ^ 1'b0 ;
  assign n25802 = n5615 & n10141 ;
  assign n25803 = ~n2747 & n25802 ;
  assign n25804 = ~n1249 & n25803 ;
  assign n25805 = n2295 & n25804 ;
  assign n25806 = n20757 ^ n4677 ^ 1'b0 ;
  assign n25807 = n6265 ^ n3367 ^ 1'b0 ;
  assign n25808 = n2142 & ~n25807 ;
  assign n25809 = n10547 & n25808 ;
  assign n25810 = ~n2680 & n5806 ;
  assign n25811 = n4239 & ~n4563 ;
  assign n25812 = n25811 ^ n3939 ^ 1'b0 ;
  assign n25813 = n25812 ^ n3877 ^ 1'b0 ;
  assign n25814 = n13913 | n25813 ;
  assign n25815 = n5010 ^ n1798 ^ 1'b0 ;
  assign n25816 = n8488 ^ n280 ^ 1'b0 ;
  assign n25817 = n15509 ^ n1437 ^ 1'b0 ;
  assign n25818 = n3621 & n25817 ;
  assign n25819 = ~n3931 & n14593 ;
  assign n25820 = n615 & n998 ;
  assign n25821 = n25820 ^ n17207 ^ 1'b0 ;
  assign n25822 = n22864 | n25821 ;
  assign n25823 = n2060 | n12339 ;
  assign n25824 = n25823 ^ n18735 ^ 1'b0 ;
  assign n25825 = n25824 ^ n10223 ^ 1'b0 ;
  assign n25826 = n434 | n3744 ;
  assign n25827 = n1118 & ~n11404 ;
  assign n25828 = n25827 ^ n25037 ^ 1'b0 ;
  assign n25829 = n24291 & n25828 ;
  assign n25830 = ~n13960 & n25829 ;
  assign n25831 = n8064 | n11355 ;
  assign n25832 = ~n17913 & n25831 ;
  assign n25833 = n2179 | n3354 ;
  assign n25834 = n25833 ^ n16212 ^ 1'b0 ;
  assign n25835 = n16313 & n22554 ;
  assign n25836 = n2912 & n25835 ;
  assign n25837 = n8199 & n14706 ;
  assign n25838 = n13111 & n14537 ;
  assign n25839 = n25838 ^ n7221 ^ n863 ;
  assign n25840 = n5013 & ~n25839 ;
  assign n25841 = n25840 ^ n14780 ^ 1'b0 ;
  assign n25842 = ~n10053 & n19688 ;
  assign n25843 = n25842 ^ n22502 ^ 1'b0 ;
  assign n25844 = n348 & n1786 ;
  assign n25845 = ~n348 & n25844 ;
  assign n25846 = n19518 & ~n25845 ;
  assign n25847 = ~n19518 & n25846 ;
  assign n25848 = n5754 ^ n273 ^ 1'b0 ;
  assign n25849 = ~n25847 & n25848 ;
  assign n25850 = ~n23 & n2436 ;
  assign n25851 = n7214 ^ n1124 ^ 1'b0 ;
  assign n25852 = n27 & ~n25851 ;
  assign n25853 = ~n12408 & n25852 ;
  assign n25854 = n25850 & ~n25853 ;
  assign n25855 = n25854 ^ n6764 ^ 1'b0 ;
  assign n25856 = n4346 ^ n3557 ^ 1'b0 ;
  assign n25857 = ( n2014 & ~n8827 ) | ( n2014 & n23684 ) | ( ~n8827 & n23684 ) ;
  assign n25858 = n3032 & ~n25857 ;
  assign n25859 = ~n20452 & n25858 ;
  assign n25860 = n11521 ^ n1219 ^ 1'b0 ;
  assign n25861 = n25746 | n25860 ;
  assign n25862 = n7346 & ~n10260 ;
  assign n25863 = ~n14121 & n25862 ;
  assign n25864 = n104 & n13165 ;
  assign n25865 = n16140 ^ n3921 ^ 1'b0 ;
  assign n25866 = ~n169 & n6240 ;
  assign n25867 = n25866 ^ n2830 ^ 1'b0 ;
  assign n25868 = n2766 & ~n3589 ;
  assign n25869 = n25868 ^ n395 ^ 1'b0 ;
  assign n25870 = n11968 & n16595 ;
  assign n25871 = ~n1704 & n25870 ;
  assign n25872 = ( ~n11827 & n25869 ) | ( ~n11827 & n25871 ) | ( n25869 & n25871 ) ;
  assign n25873 = n5083 & ~n8864 ;
  assign n25874 = n8144 & ~n11724 ;
  assign n25875 = n3146 | n25874 ;
  assign n25876 = n19475 ^ n4112 ^ 1'b0 ;
  assign n25877 = n1022 & n6062 ;
  assign n25878 = ~n9284 & n25877 ;
  assign n25879 = n11375 & ~n25878 ;
  assign n25880 = ~n2312 & n25879 ;
  assign n25881 = n11615 | n25880 ;
  assign n25882 = n25881 ^ n3034 ^ 1'b0 ;
  assign n25883 = ~n469 & n1577 ;
  assign n25884 = n25883 ^ n2403 ^ 1'b0 ;
  assign n25885 = n6316 ^ n1277 ^ 1'b0 ;
  assign n25886 = n3099 & ~n6198 ;
  assign n25887 = n25885 & n25886 ;
  assign n25888 = n11891 | n25887 ;
  assign n25889 = n14059 & n25888 ;
  assign n25890 = n25884 & n25889 ;
  assign n25892 = n6557 & n6867 ;
  assign n25893 = n25892 ^ n1602 ^ 1'b0 ;
  assign n25891 = n509 & ~n15582 ;
  assign n25894 = n25893 ^ n25891 ^ 1'b0 ;
  assign n25895 = ~n8067 & n23076 ;
  assign n25896 = n7773 & n25895 ;
  assign n25897 = n2086 ^ n512 ^ 1'b0 ;
  assign n25898 = n20446 & n25897 ;
  assign n25899 = n6084 & n7217 ;
  assign n25900 = n4373 ^ n378 ^ 1'b0 ;
  assign n25901 = n159 & ~n12429 ;
  assign n25902 = n19893 ^ n6242 ^ 1'b0 ;
  assign n25903 = n9006 & ~n25902 ;
  assign n25904 = n8547 ^ n7369 ^ 1'b0 ;
  assign n25905 = ( ~n592 & n2851 ) | ( ~n592 & n25904 ) | ( n2851 & n25904 ) ;
  assign n25906 = n7479 ^ n5245 ^ 1'b0 ;
  assign n25907 = n1248 & ~n25906 ;
  assign n25908 = n25907 ^ n14803 ^ 1'b0 ;
  assign n25909 = ~n4578 & n20408 ;
  assign n25910 = n23577 | n25909 ;
  assign n25911 = n932 | n3412 ;
  assign n25912 = n607 | n25911 ;
  assign n25913 = n25912 ^ n23762 ^ 1'b0 ;
  assign n25914 = ~n79 & n2700 ;
  assign n25915 = ~n2700 & n25914 ;
  assign n25916 = n461 & ~n25915 ;
  assign n25917 = ~n461 & n25916 ;
  assign n25918 = n6228 | n25917 ;
  assign n25919 = n3340 & ~n25918 ;
  assign n25920 = n3797 & n5568 ;
  assign n25921 = n1385 & n25920 ;
  assign n25922 = n8933 & n19705 ;
  assign n25923 = ~n7483 & n7699 ;
  assign n25924 = n8562 & ~n11245 ;
  assign n25925 = x5 & n6849 ;
  assign n25926 = n25925 ^ n6008 ^ 1'b0 ;
  assign n25927 = n25926 ^ n8170 ^ 1'b0 ;
  assign n25928 = n9855 | n16448 ;
  assign n25929 = n7271 & n25928 ;
  assign n25930 = n25929 ^ n236 ^ 1'b0 ;
  assign n25931 = n19642 & ~n25930 ;
  assign n25932 = ~n3507 & n25931 ;
  assign n25933 = n20510 & n25932 ;
  assign n25934 = n2424 & ~n6784 ;
  assign n25935 = n24045 & n25934 ;
  assign n25936 = n2514 | n5562 ;
  assign n25937 = ~n7110 & n25936 ;
  assign n25938 = ~n19762 & n25937 ;
  assign n25939 = ~n709 & n6090 ;
  assign n25941 = n16703 ^ n2070 ^ 1'b0 ;
  assign n25940 = n4339 & ~n11284 ;
  assign n25942 = n25941 ^ n25940 ^ 1'b0 ;
  assign n25943 = n3580 ^ n2604 ^ 1'b0 ;
  assign n25944 = n25943 ^ n13706 ^ 1'b0 ;
  assign n25945 = n10509 ^ n2785 ^ 1'b0 ;
  assign n25946 = ~n22700 & n25945 ;
  assign n25947 = n15986 ^ n11943 ^ 1'b0 ;
  assign n25948 = n6097 & n8987 ;
  assign n25949 = ~n13338 & n20101 ;
  assign n25954 = n16759 & n21229 ;
  assign n25955 = ~n2494 & n25954 ;
  assign n25951 = n3457 ^ n1431 ^ 1'b0 ;
  assign n25950 = n3757 | n15210 ;
  assign n25952 = n25951 ^ n25950 ^ 1'b0 ;
  assign n25953 = ~n16750 & n25952 ;
  assign n25956 = n25955 ^ n25953 ^ 1'b0 ;
  assign n25957 = n12123 & ~n21778 ;
  assign n25958 = n337 & ~n11965 ;
  assign n25959 = ~n6051 & n8365 ;
  assign n25960 = n8070 ^ n1829 ^ 1'b0 ;
  assign n25961 = n18857 ^ n1025 ^ n55 ;
  assign n25962 = n1883 & ~n20998 ;
  assign n25963 = n11520 ^ n3514 ^ 1'b0 ;
  assign n25964 = n3346 & ~n9639 ;
  assign n25965 = n11332 & n25964 ;
  assign n25966 = n5590 | n25965 ;
  assign n25967 = n22037 & ~n25966 ;
  assign n25968 = n5683 & ~n24347 ;
  assign n25969 = n21245 ^ n8617 ^ 1'b0 ;
  assign n25970 = n7753 | n16081 ;
  assign n25971 = n18430 ^ n13272 ^ 1'b0 ;
  assign n25972 = n13076 & n24664 ;
  assign n25973 = n3680 & n22092 ;
  assign n25974 = n25973 ^ n12000 ^ 1'b0 ;
  assign n25975 = n25974 ^ n12875 ^ 1'b0 ;
  assign n25976 = n6445 & ~n8053 ;
  assign n25977 = n17 | n19051 ;
  assign n25978 = n25977 ^ n21860 ^ 1'b0 ;
  assign n25979 = n7472 & ~n19538 ;
  assign n25980 = ~n25978 & n25979 ;
  assign n25981 = n216 | n25980 ;
  assign n25982 = n25981 ^ n9197 ^ 1'b0 ;
  assign n25983 = ~n476 & n18392 ;
  assign n25984 = n8311 ^ n1645 ^ 1'b0 ;
  assign n25985 = n2923 & ~n20025 ;
  assign n25986 = n2028 & n11088 ;
  assign n25987 = n2199 & ~n2933 ;
  assign n25988 = n1423 & ~n25987 ;
  assign n25989 = n8329 & ~n19837 ;
  assign n25990 = n6758 ^ n278 ^ 1'b0 ;
  assign n25991 = n25990 ^ n19198 ^ 1'b0 ;
  assign n25992 = n3326 | n25991 ;
  assign n25993 = n15673 ^ n713 ^ 1'b0 ;
  assign n25994 = n16777 ^ n13244 ^ 1'b0 ;
  assign n25995 = n2780 & n25994 ;
  assign n25996 = n12169 & ~n25995 ;
  assign n25997 = n8887 ^ n6715 ^ 1'b0 ;
  assign n25998 = n1112 & ~n14498 ;
  assign n25999 = n2362 | n25998 ;
  assign n26000 = n25997 & ~n25999 ;
  assign n26001 = n13806 ^ n1673 ^ 1'b0 ;
  assign n26002 = n11581 & n26001 ;
  assign n26003 = ~n23506 & n26002 ;
  assign n26004 = n22583 | n26003 ;
  assign n26005 = n26004 ^ n10223 ^ 1'b0 ;
  assign n26006 = n7641 & n19491 ;
  assign n26009 = n1794 & n6955 ;
  assign n26007 = n11177 ^ n5458 ^ 1'b0 ;
  assign n26008 = n26007 ^ n4911 ^ n2497 ;
  assign n26010 = n26009 ^ n26008 ^ 1'b0 ;
  assign n26011 = n1280 & n26010 ;
  assign n26012 = n14771 ^ n13614 ^ n6168 ;
  assign n26013 = n22312 | n26012 ;
  assign n26014 = n8939 ^ n1325 ^ 1'b0 ;
  assign n26015 = n1268 & n18253 ;
  assign n26016 = n16485 ^ n5255 ^ 1'b0 ;
  assign n26017 = n8208 ^ n995 ^ 1'b0 ;
  assign n26019 = n24383 ^ n5826 ^ 1'b0 ;
  assign n26020 = n9145 | n26019 ;
  assign n26018 = n18517 & n23451 ;
  assign n26021 = n26020 ^ n26018 ^ 1'b0 ;
  assign n26022 = n26017 & n26021 ;
  assign n26023 = n1765 & n20954 ;
  assign n26024 = n1235 & n6364 ;
  assign n26025 = n26024 ^ n17573 ^ 1'b0 ;
  assign n26026 = ~n1229 & n18019 ;
  assign n26027 = n26026 ^ n19776 ^ 1'b0 ;
  assign n26028 = n23683 ^ n14850 ^ 1'b0 ;
  assign n26029 = n6867 & n21002 ;
  assign n26030 = ~n1624 & n26029 ;
  assign n26031 = n13841 ^ n9432 ^ 1'b0 ;
  assign n26032 = n7091 | n26031 ;
  assign n26033 = ~n5193 & n21793 ;
  assign n26034 = n26033 ^ n17119 ^ 1'b0 ;
  assign n26035 = ~n3237 & n10019 ;
  assign n26036 = n14233 ^ n12017 ^ 1'b0 ;
  assign n26037 = n15908 ^ n2547 ^ 1'b0 ;
  assign n26038 = n804 & n25419 ;
  assign n26039 = n26038 ^ n15604 ^ 1'b0 ;
  assign n26040 = n5854 ^ n5071 ^ 1'b0 ;
  assign n26041 = n506 | n26040 ;
  assign n26042 = n4815 & ~n26041 ;
  assign n26043 = ~n11447 & n26042 ;
  assign n26044 = n5313 | n11667 ;
  assign n26045 = n26044 ^ n17683 ^ 1'b0 ;
  assign n26046 = n21657 | n26045 ;
  assign n26047 = n20449 ^ n1550 ^ 1'b0 ;
  assign n26048 = ~n22666 & n26047 ;
  assign n26049 = n14571 & ~n26048 ;
  assign n26050 = x11 & n1707 ;
  assign n26051 = n14943 ^ n8008 ^ 1'b0 ;
  assign n26052 = n1673 & n26051 ;
  assign n26053 = n6536 & ~n12217 ;
  assign n26054 = n26053 ^ n15077 ^ 1'b0 ;
  assign n26055 = n4714 & n5231 ;
  assign n26056 = ~n9239 & n26055 ;
  assign n26057 = n18940 ^ n3173 ^ 1'b0 ;
  assign n26058 = n24857 & n26057 ;
  assign n26059 = ( n791 & n12101 ) | ( n791 & ~n12955 ) | ( n12101 & ~n12955 ) ;
  assign n26060 = n14458 & n26059 ;
  assign n26061 = ~n86 & n26060 ;
  assign n26062 = n2569 & ~n26061 ;
  assign n26063 = n11089 ^ n6544 ^ 1'b0 ;
  assign n26064 = ~n4563 & n6719 ;
  assign n26065 = n26064 ^ n2898 ^ 1'b0 ;
  assign n26066 = ~n8635 & n10569 ;
  assign n26067 = n26066 ^ n8959 ^ 1'b0 ;
  assign n26068 = n356 & ~n1097 ;
  assign n26069 = n26068 ^ n3093 ^ 1'b0 ;
  assign n26070 = n1591 & ~n26069 ;
  assign n26071 = ~n1591 & n26070 ;
  assign n26072 = n19743 & ~n26071 ;
  assign n26073 = ~n11582 & n26072 ;
  assign n26074 = n11582 & n26073 ;
  assign n26075 = n21818 ^ n4497 ^ 1'b0 ;
  assign n26076 = ~n3162 & n19795 ;
  assign n26077 = n3249 & n11378 ;
  assign n26078 = n26077 ^ n252 ^ 1'b0 ;
  assign n26079 = n20716 & n26078 ;
  assign n26081 = ~n3846 & n24350 ;
  assign n26080 = n11681 & n12772 ;
  assign n26082 = n26081 ^ n26080 ^ 1'b0 ;
  assign n26083 = n26082 ^ n14335 ^ 1'b0 ;
  assign n26084 = n17196 ^ n8891 ^ 1'b0 ;
  assign n26085 = n2615 & n26014 ;
  assign n26086 = ~n26014 & n26085 ;
  assign n26087 = n10370 | n13797 ;
  assign n26088 = ~n4214 & n6339 ;
  assign n26091 = n1474 & n3785 ;
  assign n26092 = ~n1474 & n26091 ;
  assign n26093 = ~n3767 & n26092 ;
  assign n26089 = n9566 ^ n2263 ^ 1'b0 ;
  assign n26090 = n7548 & ~n26089 ;
  assign n26094 = n26093 ^ n26090 ^ 1'b0 ;
  assign n26095 = n26088 & ~n26094 ;
  assign n26096 = n11085 & n26095 ;
  assign n26097 = n13646 ^ n5979 ^ 1'b0 ;
  assign n26098 = n627 | n3189 ;
  assign n26099 = n26097 | n26098 ;
  assign n26100 = n2542 & n3668 ;
  assign n26101 = n6096 | n19117 ;
  assign n26102 = ~n26100 & n26101 ;
  assign n26103 = n8330 | n26102 ;
  assign n26104 = n4640 & n22282 ;
  assign n26105 = ~n12879 & n26104 ;
  assign n26106 = ~n6058 & n13343 ;
  assign n26107 = n26105 & n26106 ;
  assign n26108 = n4508 ^ n3489 ^ 1'b0 ;
  assign n26109 = n1326 & n23557 ;
  assign n26110 = n10882 ^ n10417 ^ 1'b0 ;
  assign n26111 = n26110 ^ n1212 ^ 1'b0 ;
  assign n26112 = n15931 ^ n7944 ^ 1'b0 ;
  assign n26113 = ~n22858 & n26112 ;
  assign n26114 = ~n6271 & n26113 ;
  assign n26115 = n26111 | n26114 ;
  assign n26116 = n2961 & n26115 ;
  assign n26117 = n22450 ^ n14681 ^ 1'b0 ;
  assign n26118 = n15790 & n26117 ;
  assign n26119 = n14834 ^ n547 ^ 1'b0 ;
  assign n26120 = n16789 | n26119 ;
  assign n26121 = n17483 & ~n26120 ;
  assign n26122 = n26121 ^ n16669 ^ 1'b0 ;
  assign n26123 = ~n10465 & n12724 ;
  assign n26124 = n26123 ^ n3100 ^ 1'b0 ;
  assign n26125 = n1588 & n8948 ;
  assign n26126 = n26125 ^ n20301 ^ 1'b0 ;
  assign n26127 = ( ~n364 & n8958 ) | ( ~n364 & n10536 ) | ( n8958 & n10536 ) ;
  assign n26128 = n328 | n5507 ;
  assign n26129 = n16407 | n26128 ;
  assign n26130 = n26129 ^ n1201 ^ 1'b0 ;
  assign n26131 = n23114 ^ n8810 ^ 1'b0 ;
  assign n26132 = n22083 ^ n19544 ^ 1'b0 ;
  assign n26133 = n671 | n23780 ;
  assign n26134 = n4616 & ~n26133 ;
  assign n26135 = n7410 | n26134 ;
  assign n26136 = n26135 ^ n12632 ^ 1'b0 ;
  assign n26137 = ~n19184 & n24985 ;
  assign n26138 = n5890 & n26137 ;
  assign n26139 = ~n26136 & n26138 ;
  assign n26140 = n7981 | n26139 ;
  assign n26141 = n119 & ~n26140 ;
  assign n26142 = n8064 ^ n36 ^ 1'b0 ;
  assign n26143 = ~x11 & n18049 ;
  assign n26144 = n20694 ^ n18485 ^ n5939 ;
  assign n26145 = n10662 ^ n133 ^ 1'b0 ;
  assign n26146 = n547 & n26145 ;
  assign n26147 = ~n768 & n26146 ;
  assign n26148 = n4879 | n13993 ;
  assign n26150 = n2875 ^ n1748 ^ 1'b0 ;
  assign n26151 = n12366 & n26150 ;
  assign n26152 = n26151 ^ n1354 ^ 1'b0 ;
  assign n26149 = ~n1401 & n21572 ;
  assign n26153 = n26152 ^ n26149 ^ 1'b0 ;
  assign n26154 = n16324 ^ n4088 ^ 1'b0 ;
  assign n26155 = ~n11837 & n26154 ;
  assign n26156 = ~n924 & n26155 ;
  assign n26157 = n18152 & n26156 ;
  assign n26158 = n7048 | n26157 ;
  assign n26159 = n26158 ^ n14742 ^ 1'b0 ;
  assign n26160 = ~n3446 & n4525 ;
  assign n26161 = ~n741 & n26160 ;
  assign n26165 = n3550 & n6303 ;
  assign n26166 = ~n3550 & n26165 ;
  assign n26162 = ~n7048 & n10197 ;
  assign n26163 = n7048 & n26162 ;
  assign n26164 = n4322 & ~n26163 ;
  assign n26167 = n26166 ^ n26164 ^ 1'b0 ;
  assign n26168 = ~n26161 & n26167 ;
  assign n26169 = n2621 & n4181 ;
  assign n26170 = n2822 & n24939 ;
  assign n26171 = ~n2822 & n26170 ;
  assign n26172 = n2556 & ~n4037 ;
  assign n26173 = n26172 ^ n288 ^ 1'b0 ;
  assign n26174 = n22441 ^ n3219 ^ 1'b0 ;
  assign n26175 = n12280 ^ n3265 ^ 1'b0 ;
  assign n26176 = n12341 | n26175 ;
  assign n26177 = n26174 & ~n26176 ;
  assign n26178 = n21597 & ~n26177 ;
  assign n26179 = n26173 & n26178 ;
  assign n26180 = n6552 ^ n3663 ^ 1'b0 ;
  assign n26181 = n188 & ~n1078 ;
  assign n26182 = n3974 & n26181 ;
  assign n26183 = ~n18968 & n26182 ;
  assign n26184 = n13490 & ~n25922 ;
  assign n26185 = n1880 & n8088 ;
  assign n26186 = n86 & n832 ;
  assign n26187 = ( n3214 & n23786 ) | ( n3214 & ~n24938 ) | ( n23786 & ~n24938 ) ;
  assign n26188 = n17181 ^ n2073 ^ 1'b0 ;
  assign n26189 = n19756 ^ n10076 ^ 1'b0 ;
  assign n26190 = n24633 ^ n17737 ^ 1'b0 ;
  assign n26191 = n16981 | n17617 ;
  assign n26192 = n19837 | n26191 ;
  assign n26193 = n11072 ^ n8548 ^ 1'b0 ;
  assign n26194 = n26192 & ~n26193 ;
  assign n26195 = n24271 ^ n3793 ^ n901 ;
  assign n26196 = n9461 ^ n2932 ^ 1'b0 ;
  assign n26197 = n3957 | n10578 ;
  assign n26198 = n8161 ^ n3189 ^ 1'b0 ;
  assign n26199 = n12379 ^ n7430 ^ 1'b0 ;
  assign n26200 = n26198 | n26199 ;
  assign n26201 = n7111 | n22230 ;
  assign n26205 = ~n2356 & n13389 ;
  assign n26202 = n3656 & n4870 ;
  assign n26203 = n26202 ^ n4900 ^ n1986 ;
  assign n26204 = n10829 & ~n26203 ;
  assign n26206 = n26205 ^ n26204 ^ 1'b0 ;
  assign n26208 = n3063 & ~n3758 ;
  assign n26207 = n8059 ^ n594 ^ 1'b0 ;
  assign n26209 = n26208 ^ n26207 ^ n22461 ;
  assign n26210 = ~n12322 & n18523 ;
  assign n26211 = n776 & ~n16751 ;
  assign n26212 = n2001 & n4746 ;
  assign n26213 = ~n8464 & n26212 ;
  assign n26214 = n332 & n26213 ;
  assign n26215 = n5939 & n7920 ;
  assign n26223 = n5613 & n17325 ;
  assign n26224 = n21136 & n26223 ;
  assign n26218 = n252 | n1739 ;
  assign n26217 = n966 & n1330 ;
  assign n26219 = n26218 ^ n26217 ^ 1'b0 ;
  assign n26220 = n12423 & ~n26219 ;
  assign n26216 = n9449 & ~n15605 ;
  assign n26221 = n26220 ^ n26216 ^ 1'b0 ;
  assign n26222 = n2822 & ~n26221 ;
  assign n26225 = n26224 ^ n26222 ^ 1'b0 ;
  assign n26226 = n20375 ^ n13984 ^ 1'b0 ;
  assign n26227 = n1668 & n26226 ;
  assign n26228 = n4247 & n9273 ;
  assign n26229 = ~n1054 & n4855 ;
  assign n26230 = n26229 ^ n1300 ^ 1'b0 ;
  assign n26231 = n13275 | n26230 ;
  assign n26232 = n18511 ^ n10607 ^ 1'b0 ;
  assign n26233 = n7524 & ~n26232 ;
  assign n26234 = n6991 & n10266 ;
  assign n26235 = n13801 ^ n7180 ^ 1'b0 ;
  assign n26236 = n16462 & ~n26235 ;
  assign n26237 = n18041 & n26236 ;
  assign n26238 = x8 & n15087 ;
  assign n26239 = n6828 & n26238 ;
  assign n26240 = n23172 ^ n6045 ^ 1'b0 ;
  assign n26241 = n26240 ^ n5626 ^ 1'b0 ;
  assign n26242 = n3420 & n26241 ;
  assign n26243 = n5724 & ~n8730 ;
  assign n26244 = n26243 ^ n9344 ^ 1'b0 ;
  assign n26245 = n26244 ^ n15434 ^ 1'b0 ;
  assign n26246 = n10444 | n26245 ;
  assign n26247 = n3150 & n26246 ;
  assign n26248 = n1740 | n8093 ;
  assign n26249 = n846 & ~n26248 ;
  assign n26250 = ~n4392 & n20535 ;
  assign n26251 = n26249 & n26250 ;
  assign n26252 = ~n4811 & n10794 ;
  assign n26253 = ~n10794 & n26252 ;
  assign n26254 = n16217 ^ n3791 ^ 1'b0 ;
  assign n26255 = n26253 | n26254 ;
  assign n26256 = n8946 ^ n302 ^ 1'b0 ;
  assign n26257 = n5776 | n21614 ;
  assign n26258 = n10007 ^ n7191 ^ 1'b0 ;
  assign n26259 = n10548 & ~n26258 ;
  assign n26260 = n15069 ^ n9478 ^ 1'b0 ;
  assign n26261 = n12888 & n26260 ;
  assign n26262 = n26261 ^ n385 ^ 1'b0 ;
  assign n26263 = ~n1974 & n18014 ;
  assign n26264 = n26263 ^ n2463 ^ 1'b0 ;
  assign n26265 = n2680 | n26264 ;
  assign n26266 = n27 & n205 ;
  assign n26267 = ~n27 & n26266 ;
  assign n26268 = n11219 & n26267 ;
  assign n26269 = n8617 | n15080 ;
  assign n26270 = n15080 & ~n26269 ;
  assign n26271 = n26270 ^ n15052 ^ 1'b0 ;
  assign n26272 = n21744 | n26271 ;
  assign n26273 = n26272 ^ n17268 ^ 1'b0 ;
  assign n26274 = n26273 ^ n7746 ^ 1'b0 ;
  assign n26275 = n26268 & n26274 ;
  assign n26276 = n23847 & n26275 ;
  assign n26277 = ~n26275 & n26276 ;
  assign n26278 = n20089 ^ n8389 ^ 1'b0 ;
  assign n26279 = n3480 ^ n715 ^ 1'b0 ;
  assign n26280 = n5845 & ~n26279 ;
  assign n26281 = n17580 & n26280 ;
  assign n26283 = n1487 & n1515 ;
  assign n26282 = n2254 & n5295 ;
  assign n26284 = n26283 ^ n26282 ^ 1'b0 ;
  assign n26289 = n8320 | n13913 ;
  assign n26287 = ~n5429 & n10081 ;
  assign n26285 = n5361 & ~n8764 ;
  assign n26286 = n8183 & n26285 ;
  assign n26288 = n26287 ^ n26286 ^ 1'b0 ;
  assign n26290 = n26289 ^ n26288 ^ n20175 ;
  assign n26291 = ~n3349 & n12110 ;
  assign n26292 = n15490 ^ n6664 ^ 1'b0 ;
  assign n26293 = ~n9925 & n26292 ;
  assign n26294 = n791 | n5626 ;
  assign n26295 = n5270 | n26294 ;
  assign n26296 = n24244 & ~n26295 ;
  assign n26297 = n17684 ^ n1246 ^ 1'b0 ;
  assign n26298 = n4965 & n7746 ;
  assign n26299 = n26297 & n26298 ;
  assign n26300 = n700 & n12879 ;
  assign n26301 = ~n18979 & n26300 ;
  assign n26302 = ~n13114 & n19028 ;
  assign n26303 = n23262 & n26302 ;
  assign n26306 = n20270 ^ n1089 ^ 1'b0 ;
  assign n26307 = n7580 & ~n26306 ;
  assign n26304 = n4473 ^ n2733 ^ 1'b0 ;
  assign n26305 = n3267 & n26304 ;
  assign n26308 = n26307 ^ n26305 ^ 1'b0 ;
  assign n26309 = ~n26303 & n26308 ;
  assign n26310 = n1175 & n25943 ;
  assign n26311 = n1772 & n3803 ;
  assign n26312 = n5205 ^ n2371 ^ 1'b0 ;
  assign n26313 = n26311 & ~n26312 ;
  assign n26314 = n10143 & ~n26313 ;
  assign n26315 = n13534 ^ n552 ^ 1'b0 ;
  assign n26316 = n16203 ^ n12926 ^ 1'b0 ;
  assign n26317 = n8918 ^ n1945 ^ 1'b0 ;
  assign n26318 = n11943 & ~n26317 ;
  assign n26319 = ~n8246 & n16160 ;
  assign n26320 = n26319 ^ n1909 ^ 1'b0 ;
  assign n26321 = n4963 & n20238 ;
  assign n26322 = n119 & n26321 ;
  assign n26323 = n9090 | n9251 ;
  assign n26324 = ( n3946 & n9911 ) | ( n3946 & n18466 ) | ( n9911 & n18466 ) ;
  assign n26325 = n9272 ^ n19 ^ 1'b0 ;
  assign n26326 = ( n7737 & n11374 ) | ( n7737 & ~n26325 ) | ( n11374 & ~n26325 ) ;
  assign n26327 = n13473 ^ n4590 ^ 1'b0 ;
  assign n26328 = n18587 ^ n3836 ^ 1'b0 ;
  assign n26329 = n8639 & ~n26328 ;
  assign n26330 = ~n3890 & n16728 ;
  assign n26331 = n3592 & n8145 ;
  assign n26332 = n2990 & n26331 ;
  assign n26333 = n26332 ^ n17845 ^ n4475 ;
  assign n26334 = n18414 ^ n3481 ^ 1'b0 ;
  assign n26335 = n5229 & n26334 ;
  assign n26336 = ( n1476 & ~n1979 ) | ( n1476 & n21614 ) | ( ~n1979 & n21614 ) ;
  assign n26337 = n11355 & n26336 ;
  assign n26338 = ~n13341 & n14929 ;
  assign n26339 = ~n3138 & n26338 ;
  assign n26340 = n247 | n747 ;
  assign n26341 = n21854 & ~n26340 ;
  assign n26342 = n26341 ^ n13996 ^ 1'b0 ;
  assign n26343 = n1931 & n3888 ;
  assign n26344 = n17976 ^ n9066 ^ 1'b0 ;
  assign n26345 = n26343 & n26344 ;
  assign n26346 = n3701 ^ n2135 ^ 1'b0 ;
  assign n26347 = n26346 ^ n1631 ^ 1'b0 ;
  assign n26348 = n10330 ^ n9228 ^ 1'b0 ;
  assign n26349 = ~n20336 & n26348 ;
  assign n26350 = n2704 & n10273 ;
  assign n26351 = n6981 ^ n6897 ^ 1'b0 ;
  assign n26352 = n26351 ^ n2939 ^ 1'b0 ;
  assign n26353 = ~n5260 & n26352 ;
  assign n26354 = n4400 | n26353 ;
  assign n26355 = n1052 & ~n14798 ;
  assign n26356 = n26354 & n26355 ;
  assign n26357 = n1688 ^ n844 ^ 1'b0 ;
  assign n26358 = n1140 & n26357 ;
  assign n26359 = n278 & n26358 ;
  assign n26360 = n26359 ^ n23320 ^ n12207 ;
  assign n26361 = n10470 ^ n4387 ^ 1'b0 ;
  assign n26362 = ~n8061 & n26361 ;
  assign n26363 = n26362 ^ n5582 ^ 1'b0 ;
  assign n26364 = n26363 ^ n636 ^ 1'b0 ;
  assign n26365 = n1795 & n26364 ;
  assign n26366 = ~n19 & n25384 ;
  assign n26367 = ~n8004 & n26366 ;
  assign n26368 = n11968 & n24454 ;
  assign n26369 = n13028 & ~n26368 ;
  assign n26370 = n26369 ^ n7319 ^ 1'b0 ;
  assign n26371 = n13679 & ~n25190 ;
  assign n26372 = n6407 & n26371 ;
  assign n26373 = n10480 ^ n8520 ^ 1'b0 ;
  assign n26374 = n3676 & n8500 ;
  assign n26375 = n26373 & ~n26374 ;
  assign n26376 = ~n310 & n17522 ;
  assign n26377 = n15142 ^ n5252 ^ 1'b0 ;
  assign n26378 = n178 | n20745 ;
  assign n26379 = n26378 ^ n9447 ^ 1'b0 ;
  assign n26380 = ~n1506 & n7662 ;
  assign n26381 = n20549 ^ n19416 ^ 1'b0 ;
  assign n26382 = n18221 ^ n14303 ^ 1'b0 ;
  assign n26383 = n6444 & n26382 ;
  assign n26384 = ~n951 & n3744 ;
  assign n26385 = n26384 ^ n3324 ^ 1'b0 ;
  assign n26386 = n26383 & ~n26385 ;
  assign n26387 = n26386 ^ n5802 ^ 1'b0 ;
  assign n26388 = n215 | n1437 ;
  assign n26389 = n9001 | n26388 ;
  assign n26390 = n402 | n26389 ;
  assign n26391 = n1418 | n6165 ;
  assign n26392 = n1264 | n25481 ;
  assign n26393 = ~n3311 & n4036 ;
  assign n26394 = ~n18252 & n26393 ;
  assign n26395 = n7564 | n24498 ;
  assign n26396 = n11907 & n12924 ;
  assign n26397 = n6135 & ~n26396 ;
  assign n26398 = n4163 & n26397 ;
  assign n26399 = n24102 | n26398 ;
  assign n26400 = n3663 | n3674 ;
  assign n26401 = n6421 | n26400 ;
  assign n26402 = n26401 ^ n9696 ^ n8616 ;
  assign n26403 = n4436 ^ x11 ^ 1'b0 ;
  assign n26404 = n3461 & ~n4055 ;
  assign n26405 = n26404 ^ n765 ^ 1'b0 ;
  assign n26406 = n12683 & ~n26405 ;
  assign n26407 = ~n26403 & n26406 ;
  assign n26408 = n23048 ^ n2808 ^ 1'b0 ;
  assign n26409 = n1115 | n13123 ;
  assign n26410 = n26408 | n26409 ;
  assign n26411 = n26410 ^ n3634 ^ 1'b0 ;
  assign n26412 = n1584 | n26411 ;
  assign n26413 = n26412 ^ n5837 ^ 1'b0 ;
  assign n26414 = n24284 ^ n2728 ^ 1'b0 ;
  assign n26418 = n7384 ^ n890 ^ 1'b0 ;
  assign n26415 = n6248 & n16906 ;
  assign n26416 = ~n7650 & n14481 ;
  assign n26417 = n26415 & n26416 ;
  assign n26419 = n26418 ^ n26417 ^ 1'b0 ;
  assign n26420 = n26414 | n26419 ;
  assign n26421 = n5386 & ~n9447 ;
  assign n26422 = ~n616 & n2899 ;
  assign n26423 = ~n3150 & n26422 ;
  assign n26424 = n9914 ^ n1491 ^ 1'b0 ;
  assign n26425 = n11535 & ~n26424 ;
  assign n26426 = ~n832 & n26425 ;
  assign n26427 = n12472 ^ n7253 ^ 1'b0 ;
  assign n26428 = n20347 & n26427 ;
  assign n26429 = ~n2294 & n3110 ;
  assign n26430 = n259 ^ n148 ^ 1'b0 ;
  assign n26431 = ~n26429 & n26430 ;
  assign n26432 = n16307 | n26431 ;
  assign n26433 = n10861 & ~n26432 ;
  assign n26434 = n26433 ^ n8480 ^ 1'b0 ;
  assign n26445 = n2843 ^ n2322 ^ 1'b0 ;
  assign n26435 = n10846 ^ n6198 ^ 1'b0 ;
  assign n26436 = n18043 ^ n9222 ^ 1'b0 ;
  assign n26437 = ~n9375 & n26436 ;
  assign n26438 = ~n820 & n14682 ;
  assign n26439 = n26438 ^ n16909 ^ 1'b0 ;
  assign n26440 = n26439 ^ n22108 ^ 1'b0 ;
  assign n26441 = n15791 | n26440 ;
  assign n26442 = n16821 | n26441 ;
  assign n26443 = n26437 | n26442 ;
  assign n26444 = ~n26435 & n26443 ;
  assign n26446 = n26445 ^ n26444 ^ 1'b0 ;
  assign n26447 = n8660 | n22777 ;
  assign n26448 = n18598 ^ n18461 ^ n12101 ;
  assign n26449 = n2196 & ~n4263 ;
  assign n26450 = n19922 & n26449 ;
  assign n26451 = ~n1525 & n5325 ;
  assign n26452 = ~n4303 & n26451 ;
  assign n26459 = n3329 & ~n19410 ;
  assign n26460 = n26459 ^ n1345 ^ 1'b0 ;
  assign n26456 = n1184 | n3451 ;
  assign n26457 = n26456 ^ n919 ^ 1'b0 ;
  assign n26453 = n1659 ^ n294 ^ 1'b0 ;
  assign n26454 = n24769 ^ n14941 ^ 1'b0 ;
  assign n26455 = n26453 | n26454 ;
  assign n26458 = n26457 ^ n26455 ^ 1'b0 ;
  assign n26461 = n26460 ^ n26458 ^ 1'b0 ;
  assign n26462 = n26461 ^ n14528 ^ 1'b0 ;
  assign n26463 = n13529 ^ n9039 ^ n7472 ;
  assign n26464 = n26463 ^ n2278 ^ 1'b0 ;
  assign n26465 = n3456 ^ n3344 ^ 1'b0 ;
  assign n26466 = n1957 & ~n26465 ;
  assign n26467 = n10451 ^ n6090 ^ 1'b0 ;
  assign n26468 = n24856 ^ n23781 ^ 1'b0 ;
  assign n26469 = n3699 & n14203 ;
  assign n26470 = n19158 & n20401 ;
  assign n26471 = n26470 ^ n17861 ^ 1'b0 ;
  assign n26472 = ~n8800 & n15047 ;
  assign n26473 = n26472 ^ n23246 ^ 1'b0 ;
  assign n26474 = ~n2879 & n23569 ;
  assign n26475 = n15631 & ~n20527 ;
  assign n26476 = n5498 ^ n1480 ^ 1'b0 ;
  assign n26477 = n17272 | n26476 ;
  assign n26478 = n18484 & ~n26477 ;
  assign n26479 = n55 | n9402 ;
  assign n26480 = n17885 & ~n18286 ;
  assign n26481 = n3396 & n26480 ;
  assign n26482 = x0 | n26481 ;
  assign n26483 = n10787 & ~n26482 ;
  assign n26484 = n15435 & ~n17361 ;
  assign n26485 = n16643 & n24885 ;
  assign n26486 = n26484 & n26485 ;
  assign n26487 = n1887 & n8587 ;
  assign n26488 = ~n23781 & n26487 ;
  assign n26489 = n22352 ^ n7193 ^ 1'b0 ;
  assign n26490 = ~n6870 & n18935 ;
  assign n26491 = n26490 ^ n15539 ^ 1'b0 ;
  assign n26492 = n1179 & n26491 ;
  assign n26493 = n26492 ^ n21059 ^ n297 ;
  assign n26494 = n6822 ^ n191 ^ 1'b0 ;
  assign n26495 = n26494 ^ n10734 ^ 1'b0 ;
  assign n26496 = n16993 ^ n6242 ^ 1'b0 ;
  assign n26497 = n26495 & ~n26496 ;
  assign n26498 = n5752 & ~n10908 ;
  assign n26499 = n12349 & n26498 ;
  assign n26500 = n25818 | n26499 ;
  assign n26501 = ~n3663 & n15862 ;
  assign n26502 = n2095 | n26501 ;
  assign n26503 = x11 & ~n3067 ;
  assign n26504 = n1891 & n26503 ;
  assign n26505 = n26504 ^ n23440 ^ n17695 ;
  assign n26506 = n15814 ^ n2205 ^ 1'b0 ;
  assign n26507 = ~n18067 & n26506 ;
  assign n26508 = n685 | n17349 ;
  assign n26509 = n26508 ^ n12974 ^ 1'b0 ;
  assign n26510 = n34 & n26509 ;
  assign n26511 = n636 | n4346 ;
  assign n26512 = n26511 ^ n19600 ^ 1'b0 ;
  assign n26513 = ~n11167 & n19521 ;
  assign n26514 = n4586 & n5527 ;
  assign n26515 = n26514 ^ n6580 ^ 1'b0 ;
  assign n26516 = n26515 ^ n9614 ^ 1'b0 ;
  assign n26517 = n13588 & ~n24019 ;
  assign n26518 = n26517 ^ n18031 ^ 1'b0 ;
  assign n26519 = ~n2148 & n3186 ;
  assign n26520 = n1533 & ~n18589 ;
  assign n26521 = n3389 & ~n5429 ;
  assign n26522 = n26521 ^ n4974 ^ 1'b0 ;
  assign n26523 = ( n914 & n24770 ) | ( n914 & n26522 ) | ( n24770 & n26522 ) ;
  assign n26524 = n5241 & ~n6552 ;
  assign n26525 = ~n25154 & n26524 ;
  assign n26526 = n1878 | n4485 ;
  assign n26527 = n3899 | n18663 ;
  assign n26528 = n26527 ^ n11845 ^ 1'b0 ;
  assign n26529 = n6481 ^ n4396 ^ 1'b0 ;
  assign n26530 = n19881 ^ n14907 ^ 1'b0 ;
  assign n26531 = n20578 ^ n11935 ^ n8512 ;
  assign n26532 = n13781 ^ n11157 ^ 1'b0 ;
  assign n26533 = n6104 & ~n21647 ;
  assign n26534 = n26533 ^ n6539 ^ 1'b0 ;
  assign n26535 = ~n2730 & n3338 ;
  assign n26536 = n26535 ^ n1450 ^ 1'b0 ;
  assign n26537 = n4320 & n26536 ;
  assign n26538 = n26537 ^ n281 ^ 1'b0 ;
  assign n26539 = n7694 | n10786 ;
  assign n26540 = n7694 & ~n26539 ;
  assign n26541 = n1572 & ~n26540 ;
  assign n26542 = n26541 ^ n7902 ^ 1'b0 ;
  assign n26543 = n16298 | n26542 ;
  assign n26544 = n196 & ~n294 ;
  assign n26545 = n294 & n26544 ;
  assign n26546 = ~n2414 & n26545 ;
  assign n26547 = ~n10592 & n11239 ;
  assign n26548 = n26546 | n26547 ;
  assign n26549 = n26543 & ~n26548 ;
  assign n26550 = n3896 & n19158 ;
  assign n26551 = n12199 ^ n5068 ^ 1'b0 ;
  assign n26552 = n16 | n13055 ;
  assign n26553 = ~n13326 & n26552 ;
  assign n26554 = n15495 & n26553 ;
  assign n26555 = n8543 & n22507 ;
  assign n26556 = n161 & n17409 ;
  assign n26557 = ~n471 & n26556 ;
  assign n26558 = n471 & n26557 ;
  assign n26559 = n4203 & n14626 ;
  assign n26560 = n939 & ~n10655 ;
  assign n26561 = n26559 & n26560 ;
  assign n26562 = n5952 & ~n26561 ;
  assign n26563 = ~n26558 & n26562 ;
  assign n26564 = n26558 & n26563 ;
  assign n26565 = n1895 | n11377 ;
  assign n26566 = n25108 ^ n1734 ^ n757 ;
  assign n26567 = ~n7008 & n26566 ;
  assign n26568 = n2263 | n17891 ;
  assign n26569 = n1686 & n14759 ;
  assign n26570 = n2194 & n26569 ;
  assign n26571 = n84 & n26570 ;
  assign n26572 = ~n6134 & n11531 ;
  assign n26573 = n25878 ^ n1711 ^ 1'b0 ;
  assign n26574 = n11724 ^ n7450 ^ 1'b0 ;
  assign n26575 = n3624 | n5812 ;
  assign n26576 = n26575 ^ n637 ^ 1'b0 ;
  assign n26577 = n9335 & n26576 ;
  assign n26578 = n1523 ^ n1366 ^ 1'b0 ;
  assign n26579 = n21557 | n26578 ;
  assign n26580 = n26577 | n26579 ;
  assign n26581 = ( n1957 & n11464 ) | ( n1957 & n13088 ) | ( n11464 & n13088 ) ;
  assign n26582 = n10475 & ~n26581 ;
  assign n26583 = ~n26580 & n26582 ;
  assign n26584 = n7717 & ~n8720 ;
  assign n26586 = n1567 & ~n6285 ;
  assign n26585 = n6383 & n19420 ;
  assign n26587 = n26586 ^ n26585 ^ 1'b0 ;
  assign n26588 = n26587 ^ n12660 ^ 1'b0 ;
  assign n26589 = n26584 | n26588 ;
  assign n26590 = n708 | n12982 ;
  assign n26591 = n2280 | n26590 ;
  assign n26592 = n13261 ^ n610 ^ 1'b0 ;
  assign n26593 = ~n666 & n26592 ;
  assign n26594 = n26591 & ~n26593 ;
  assign n26595 = ( n760 & n7792 ) | ( n760 & ~n17178 ) | ( n7792 & ~n17178 ) ;
  assign n26596 = n26595 ^ n25622 ^ 1'b0 ;
  assign n26597 = n6009 ^ n163 ^ 1'b0 ;
  assign n26598 = n10835 ^ n2893 ^ 1'b0 ;
  assign n26599 = n82 | n10383 ;
  assign n26600 = n1693 & n26599 ;
  assign n26601 = n769 | n26600 ;
  assign n26602 = n26598 & ~n26601 ;
  assign n26606 = ~n616 & n3818 ;
  assign n26607 = n545 & n26606 ;
  assign n26603 = n942 & n11796 ;
  assign n26604 = n26603 ^ n22059 ^ 1'b0 ;
  assign n26605 = n12798 & n26604 ;
  assign n26608 = n26607 ^ n26605 ^ 1'b0 ;
  assign n26609 = ~n13855 & n26608 ;
  assign n26610 = n3552 & ~n12674 ;
  assign n26611 = n12013 & n26610 ;
  assign n26612 = n26611 ^ n1315 ^ 1'b0 ;
  assign n26613 = n3589 & ~n11328 ;
  assign n26614 = n6608 | n26613 ;
  assign n26615 = n6463 & ~n15718 ;
  assign n26616 = n25810 ^ n11153 ^ 1'b0 ;
  assign n26617 = n15198 & n19058 ;
  assign n26618 = ~n14231 & n26617 ;
  assign n26619 = n17998 | n23394 ;
  assign n26620 = n9655 | n26619 ;
  assign n26621 = n10780 & n26620 ;
  assign n26622 = ~n1692 & n25526 ;
  assign n26623 = ~n15450 & n26622 ;
  assign n26624 = n6249 & n26623 ;
  assign n26625 = n15576 ^ n4757 ^ n2509 ;
  assign n26626 = n1699 & ~n8450 ;
  assign n26627 = n1950 & ~n20641 ;
  assign n26628 = n26627 ^ n233 ^ 1'b0 ;
  assign n26629 = n20495 ^ n336 ^ 1'b0 ;
  assign n26630 = n14737 | n26629 ;
  assign n26631 = n11943 | n26611 ;
  assign n26632 = ( n2694 & ~n26630 ) | ( n2694 & n26631 ) | ( ~n26630 & n26631 ) ;
  assign n26635 = n2432 ^ n1482 ^ 1'b0 ;
  assign n26633 = n13687 ^ n12324 ^ 1'b0 ;
  assign n26634 = n2270 | n26633 ;
  assign n26636 = n26635 ^ n26634 ^ 1'b0 ;
  assign n26637 = n8988 & n12913 ;
  assign n26638 = n2472 & ~n2894 ;
  assign n26639 = n17613 ^ n15915 ^ 1'b0 ;
  assign n26640 = n1175 & n1872 ;
  assign n26641 = ~n5686 & n10914 ;
  assign n26642 = n26641 ^ n1744 ^ 1'b0 ;
  assign n26643 = n9151 & n17252 ;
  assign n26644 = n19438 ^ n1010 ^ 1'b0 ;
  assign n26645 = n6543 & n26644 ;
  assign n26646 = n8523 & ~n13690 ;
  assign n26647 = n9088 ^ n4533 ^ 1'b0 ;
  assign n26648 = n26646 & n26647 ;
  assign n26649 = n15478 ^ n14884 ^ 1'b0 ;
  assign n26650 = n13183 | n26649 ;
  assign n26651 = n685 & ~n24512 ;
  assign n26652 = n26651 ^ n10482 ^ n3560 ;
  assign n26654 = n8412 | n20108 ;
  assign n26655 = n26654 ^ n6903 ^ 1'b0 ;
  assign n26656 = n10192 & ~n26655 ;
  assign n26657 = n26656 ^ n9897 ^ 1'b0 ;
  assign n26658 = n1385 & n26657 ;
  assign n26653 = n1207 & ~n2452 ;
  assign n26659 = n26658 ^ n26653 ^ 1'b0 ;
  assign n26660 = n18035 ^ n15163 ^ 1'b0 ;
  assign n26661 = n9420 & ~n26660 ;
  assign n26662 = ~n19211 & n26661 ;
  assign n26663 = n26662 ^ n11761 ^ 1'b0 ;
  assign n26664 = n7520 | n13094 ;
  assign n26665 = n5283 & ~n26664 ;
  assign n26666 = n507 & n26665 ;
  assign n26667 = n5326 | n7096 ;
  assign n26668 = ~n19527 & n26667 ;
  assign n26669 = n5996 | n22590 ;
  assign n26670 = n1718 & ~n26669 ;
  assign n26671 = n9043 ^ n1460 ^ 1'b0 ;
  assign n26672 = n17772 & n26671 ;
  assign n26673 = n24665 ^ n3037 ^ 1'b0 ;
  assign n26674 = ~n23234 & n24141 ;
  assign n26675 = ~n8850 & n26674 ;
  assign n26677 = n703 & ~n21855 ;
  assign n26676 = n8360 | n15606 ;
  assign n26678 = n26677 ^ n26676 ^ 1'b0 ;
  assign n26680 = n3527 | n10973 ;
  assign n26679 = n8429 & ~n25519 ;
  assign n26681 = n26680 ^ n26679 ^ 1'b0 ;
  assign n26682 = n1851 & ~n12053 ;
  assign n26683 = n26682 ^ n15515 ^ 1'b0 ;
  assign n26684 = n8510 | n24828 ;
  assign n26685 = n3355 | n26684 ;
  assign n26686 = n1218 & n2078 ;
  assign n26687 = ~n1218 & n26686 ;
  assign n26688 = n55 | n26687 ;
  assign n26689 = n55 & ~n26688 ;
  assign n26690 = n489 & n5597 ;
  assign n26691 = ~n489 & n26690 ;
  assign n26692 = n10973 | n26691 ;
  assign n26693 = n1166 & ~n26692 ;
  assign n26694 = n26689 & n26693 ;
  assign n26695 = n15971 ^ n8093 ^ 1'b0 ;
  assign n26696 = n338 & n20854 ;
  assign n26697 = ~n20702 & n26696 ;
  assign n26698 = n2433 & n26697 ;
  assign n26699 = n26695 | n26698 ;
  assign n26700 = n26695 & ~n26699 ;
  assign n26701 = n4306 & ~n14683 ;
  assign n26702 = ~n4306 & n26701 ;
  assign n26703 = n2315 | n26702 ;
  assign n26704 = n2315 & ~n26703 ;
  assign n26705 = n26700 | n26704 ;
  assign n26706 = n26694 & ~n26705 ;
  assign n26707 = n13109 ^ n828 ^ n737 ;
  assign n26708 = ~n1880 & n12079 ;
  assign n26709 = n26708 ^ n10751 ^ 1'b0 ;
  assign n26710 = ( n2112 & n9672 ) | ( n2112 & ~n26709 ) | ( n9672 & ~n26709 ) ;
  assign n26711 = n17118 ^ n5832 ^ 1'b0 ;
  assign n26712 = n7654 | n26711 ;
  assign n26713 = n6001 ^ n839 ^ 1'b0 ;
  assign n26714 = n26713 ^ n4929 ^ 1'b0 ;
  assign n26715 = n2420 | n9785 ;
  assign n26716 = n220 & n26715 ;
  assign n26717 = n26716 ^ n15484 ^ 1'b0 ;
  assign n26718 = n19934 | n26717 ;
  assign n26719 = n1575 | n9796 ;
  assign n26720 = n14808 & n26719 ;
  assign n26721 = n1138 ^ n187 ^ 1'b0 ;
  assign n26722 = n5309 & ~n26721 ;
  assign n26723 = n6143 & n26722 ;
  assign n26724 = ~n3305 & n26723 ;
  assign n26725 = n5002 & ~n26724 ;
  assign n26726 = n18367 | n26185 ;
  assign n26728 = n3645 & ~n7330 ;
  assign n26727 = ~n5637 & n17315 ;
  assign n26729 = n26728 ^ n26727 ^ 1'b0 ;
  assign n26730 = n83 & n2414 ;
  assign n26731 = ~n19830 & n26730 ;
  assign n26732 = n15931 & ~n19392 ;
  assign n26733 = n19129 ^ n142 ^ 1'b0 ;
  assign n26735 = n66 & n8412 ;
  assign n26736 = n2724 | n26735 ;
  assign n26734 = n10876 & ~n18280 ;
  assign n26737 = n26736 ^ n26734 ^ 1'b0 ;
  assign n26738 = n26737 ^ n799 ^ 1'b0 ;
  assign n26739 = n6864 & n12220 ;
  assign n26740 = n1505 | n9108 ;
  assign n26741 = n1645 & ~n14440 ;
  assign n26742 = ~n541 & n6338 ;
  assign n26743 = n2842 & n10407 ;
  assign n26744 = n5908 & n26743 ;
  assign n26745 = n26744 ^ n7003 ^ 1'b0 ;
  assign n26746 = n16826 & n22814 ;
  assign n26747 = n26746 ^ n1857 ^ 1'b0 ;
  assign n26748 = n7892 ^ n1655 ^ 1'b0 ;
  assign n26749 = n25274 & ~n26748 ;
  assign n26750 = n26749 ^ n12040 ^ 1'b0 ;
  assign n26751 = ~n7996 & n17607 ;
  assign n26752 = n26751 ^ n1274 ^ 1'b0 ;
  assign n26753 = n19998 ^ n6661 ^ 1'b0 ;
  assign n26754 = n26752 & n26753 ;
  assign n26755 = ~n7266 & n10420 ;
  assign n26756 = ~n2408 & n26755 ;
  assign n26757 = ~n5378 & n26756 ;
  assign n26758 = n26757 ^ n5775 ^ 1'b0 ;
  assign n26759 = n5280 & ~n6224 ;
  assign n26760 = n26759 ^ n6772 ^ 1'b0 ;
  assign n26761 = n26760 ^ n7144 ^ 1'b0 ;
  assign n26762 = n11003 & ~n26761 ;
  assign n26763 = n549 & ~n3037 ;
  assign n26764 = ~n4171 & n26763 ;
  assign n26765 = ~n26762 & n26764 ;
  assign n26766 = n4483 & n10057 ;
  assign n26767 = n10547 & n26766 ;
  assign n26768 = n5330 & ~n14085 ;
  assign n26769 = n26768 ^ n9166 ^ 1'b0 ;
  assign n26770 = n8275 | n26769 ;
  assign n26771 = n121 & ~n151 ;
  assign n26772 = n423 | n1347 ;
  assign n26773 = n26772 ^ n13125 ^ n12562 ;
  assign n26774 = ~n84 & n26773 ;
  assign n26775 = ~n26771 & n26774 ;
  assign n26776 = ~n11992 & n15224 ;
  assign n26777 = n15626 | n23167 ;
  assign n26778 = n26777 ^ n5789 ^ 1'b0 ;
  assign n26779 = n9862 ^ n847 ^ 1'b0 ;
  assign n26780 = n19533 & n26779 ;
  assign n26781 = n26780 ^ n1396 ^ 1'b0 ;
  assign n26782 = n26781 ^ n24637 ^ n10673 ;
  assign n26783 = n25501 ^ n6477 ^ 1'b0 ;
  assign n26784 = n10186 & n26783 ;
  assign n26785 = ~n8648 & n26784 ;
  assign n26786 = n20652 & ~n26785 ;
  assign n26787 = n1112 & n23207 ;
  assign n26788 = ~n11042 & n12952 ;
  assign n26789 = n7096 & n26788 ;
  assign n26790 = ~n2060 & n26789 ;
  assign n26791 = n7227 ^ n6951 ^ 1'b0 ;
  assign n26792 = n233 & n292 ;
  assign n26793 = n13171 ^ n4109 ^ 1'b0 ;
  assign n26794 = n11566 & n26793 ;
  assign n26795 = n2898 | n26794 ;
  assign n26800 = n3993 ^ n2220 ^ n533 ;
  assign n26796 = n1868 ^ n747 ^ 1'b0 ;
  assign n26797 = n26796 ^ n4347 ^ 1'b0 ;
  assign n26798 = n2075 & n26797 ;
  assign n26799 = n26798 ^ n15557 ^ 1'b0 ;
  assign n26801 = n26800 ^ n26799 ^ 1'b0 ;
  assign n26802 = ~n325 & n26801 ;
  assign n26803 = n26802 ^ n12457 ^ 1'b0 ;
  assign n26804 = n3951 & ~n23887 ;
  assign n26822 = n3721 & n7357 ;
  assign n26823 = ~n7357 & n26822 ;
  assign n26824 = n5972 | n26823 ;
  assign n26805 = n255 | n403 ;
  assign n26806 = n7829 & ~n26805 ;
  assign n26807 = n1975 & n26806 ;
  assign n26808 = n26807 ^ n782 ^ 1'b0 ;
  assign n26809 = n412 & n466 ;
  assign n26810 = ~n466 & n26809 ;
  assign n26811 = n1412 & ~n26810 ;
  assign n26812 = n609 & ~n821 ;
  assign n26813 = ~n609 & n26812 ;
  assign n26814 = ~n24802 & n26813 ;
  assign n26815 = ~n1284 & n26814 ;
  assign n26816 = ~n26811 & n26815 ;
  assign n26817 = n4061 & n26816 ;
  assign n26818 = n3150 & n26817 ;
  assign n26819 = n15231 | n26818 ;
  assign n26820 = n26818 & ~n26819 ;
  assign n26821 = n26808 & ~n26820 ;
  assign n26825 = n26824 ^ n26821 ^ 1'b0 ;
  assign n26826 = n624 | n4590 ;
  assign n26827 = n9760 ^ n5912 ^ 1'b0 ;
  assign n26828 = ~n6361 & n19550 ;
  assign n26829 = n26828 ^ n19630 ^ 1'b0 ;
  assign n26830 = n5097 & ~n18097 ;
  assign n26831 = n16972 ^ n5118 ^ 1'b0 ;
  assign n26832 = n10121 | n26831 ;
  assign n26833 = n26832 ^ n2932 ^ 1'b0 ;
  assign n26834 = n2150 & ~n13266 ;
  assign n26835 = n26834 ^ n6417 ^ n290 ;
  assign n26836 = n43 & ~n6046 ;
  assign n26837 = n23057 ^ n553 ^ 1'b0 ;
  assign n26838 = n1854 | n18925 ;
  assign n26839 = n423 & n7419 ;
  assign n26840 = n26839 ^ n2693 ^ 1'b0 ;
  assign n26841 = n11740 & ~n26840 ;
  assign n26842 = n26841 ^ n612 ^ 1'b0 ;
  assign n26843 = n1795 | n17176 ;
  assign n26844 = n18778 ^ n9758 ^ n7135 ;
  assign n26845 = ~n26843 & n26844 ;
  assign n26846 = n7965 | n12913 ;
  assign n26847 = n26846 ^ n34 ^ 1'b0 ;
  assign n26848 = n4864 ^ n3107 ^ 1'b0 ;
  assign n26849 = n22867 | n26848 ;
  assign n26850 = n10158 & ~n20014 ;
  assign n26851 = n8384 & n26850 ;
  assign n26852 = n21791 ^ n1310 ^ 1'b0 ;
  assign n26853 = n15065 ^ n8942 ^ 1'b0 ;
  assign n26854 = ~n75 & n7661 ;
  assign n26855 = ( n3645 & ~n24824 ) | ( n3645 & n26854 ) | ( ~n24824 & n26854 ) ;
  assign n26856 = n26855 ^ n759 ^ 1'b0 ;
  assign n26857 = n20505 ^ n9208 ^ 1'b0 ;
  assign n26858 = n4756 & ~n8878 ;
  assign n26859 = ~n7714 & n19302 ;
  assign n26860 = n5917 | n15725 ;
  assign n26861 = n9541 | n26860 ;
  assign n26862 = n26861 ^ n17791 ^ 1'b0 ;
  assign n26863 = n6194 | n20505 ;
  assign n26864 = n18131 ^ n14206 ^ 1'b0 ;
  assign n26865 = n6534 & ~n26864 ;
  assign n26866 = n26865 ^ n8067 ^ 1'b0 ;
  assign n26867 = n433 & n3986 ;
  assign n26868 = ~n433 & n26867 ;
  assign n26869 = n32 | n26868 ;
  assign n26870 = n32 & ~n26869 ;
  assign n26871 = n13231 | n26870 ;
  assign n26872 = n13231 & ~n26871 ;
  assign n26873 = ~n6906 & n16855 ;
  assign n26874 = ~n16855 & n26873 ;
  assign n26875 = n26872 | n26874 ;
  assign n26876 = n26866 | n26875 ;
  assign n26877 = n5002 | n17592 ;
  assign n26878 = n17063 ^ n9778 ^ 1'b0 ;
  assign n26879 = n94 & ~n26878 ;
  assign n26880 = ~n11888 & n15426 ;
  assign n26881 = n26880 ^ n940 ^ 1'b0 ;
  assign n26882 = ( n278 & ~n2593 ) | ( n278 & n10625 ) | ( ~n2593 & n10625 ) ;
  assign n26883 = n4288 & ~n12641 ;
  assign n26884 = ~n12987 & n13471 ;
  assign n26885 = n26884 ^ n5802 ^ 1'b0 ;
  assign n26886 = n10990 ^ n836 ^ 1'b0 ;
  assign n26887 = n9152 ^ n5350 ^ 1'b0 ;
  assign n26888 = n5733 & n26887 ;
  assign n26889 = n26888 ^ n24491 ^ 1'b0 ;
  assign n26893 = ~n9514 & n13588 ;
  assign n26890 = n3255 ^ n1686 ^ 1'b0 ;
  assign n26891 = ~n14573 & n26890 ;
  assign n26892 = ~n18748 & n26891 ;
  assign n26894 = n26893 ^ n26892 ^ 1'b0 ;
  assign n26895 = n7285 & n26894 ;
  assign n26896 = n9235 ^ n8683 ^ 1'b0 ;
  assign n26897 = ( n2437 & n16677 ) | ( n2437 & ~n26896 ) | ( n16677 & ~n26896 ) ;
  assign n26898 = n13425 & n14768 ;
  assign n26899 = n26898 ^ n22970 ^ 1'b0 ;
  assign n26900 = n11207 & n26681 ;
  assign n26901 = n13778 ^ n5336 ^ 1'b0 ;
  assign n26902 = n21194 & ~n22265 ;
  assign n26903 = n461 | n8562 ;
  assign n26904 = n17229 & ~n26903 ;
  assign n26905 = ~n1283 & n1309 ;
  assign n26906 = n21772 & ~n24333 ;
  assign n26907 = n26906 ^ n13769 ^ 1'b0 ;
  assign n26908 = n11079 ^ n5370 ^ 1'b0 ;
  assign n26909 = n1865 | n26908 ;
  assign n26910 = n7802 ^ n2943 ^ 1'b0 ;
  assign n26911 = ~n26909 & n26910 ;
  assign n26912 = n26911 ^ n12072 ^ 1'b0 ;
  assign n26913 = n5202 | n6912 ;
  assign n26914 = n26913 ^ n8392 ^ 1'b0 ;
  assign n26915 = n3687 & ~n26914 ;
  assign n26918 = ~n1113 & n14046 ;
  assign n26919 = ~n14046 & n26918 ;
  assign n26916 = n14398 ^ n7483 ^ 1'b0 ;
  assign n26917 = ~n19388 & n26916 ;
  assign n26920 = n26919 ^ n26917 ^ n7264 ;
  assign n26921 = n5412 & n18826 ;
  assign n26922 = n26921 ^ n782 ^ 1'b0 ;
  assign n26923 = n26922 ^ n23843 ^ 1'b0 ;
  assign n26924 = n7780 ^ n2403 ^ 1'b0 ;
  assign n26925 = n26924 ^ n9776 ^ 1'b0 ;
  assign n26926 = n26923 & n26925 ;
  assign n26927 = n9892 ^ n2983 ^ 1'b0 ;
  assign n26928 = n484 | n26927 ;
  assign n26929 = ~n6599 & n14614 ;
  assign n26930 = n6752 & n26929 ;
  assign n26931 = n11849 | n26930 ;
  assign n26932 = n26928 & ~n26931 ;
  assign n26933 = n1026 & ~n10578 ;
  assign n26934 = n8967 | n26933 ;
  assign n26935 = n26934 ^ n1676 ^ 1'b0 ;
  assign n26936 = n8036 & ~n26935 ;
  assign n26937 = n508 | n1777 ;
  assign n26938 = n7147 & ~n26937 ;
  assign n26939 = n26938 ^ n55 ^ 1'b0 ;
  assign n26940 = ( n649 & n7649 ) | ( n649 & ~n21525 ) | ( n7649 & ~n21525 ) ;
  assign n26941 = n26940 ^ n5820 ^ 1'b0 ;
  assign n26942 = n26939 & ~n26941 ;
  assign n26943 = n3899 | n6519 ;
  assign n26944 = n26943 ^ n2001 ^ 1'b0 ;
  assign n26945 = n12944 | n21627 ;
  assign n26946 = n11189 ^ n8963 ^ 1'b0 ;
  assign n26947 = ~n11501 & n16303 ;
  assign n26948 = n26947 ^ n9397 ^ 1'b0 ;
  assign n26949 = ~n14219 & n19575 ;
  assign n26950 = ~n20078 & n26949 ;
  assign n26951 = ~n200 & n8711 ;
  assign n26952 = ~n14694 & n26951 ;
  assign n26953 = n8233 & n26952 ;
  assign n26954 = n1281 & ~n9463 ;
  assign n26955 = n14 & n26954 ;
  assign n26956 = ( n4700 & n15165 ) | ( n4700 & n26955 ) | ( n15165 & n26955 ) ;
  assign n26957 = ~n1968 & n26956 ;
  assign n26958 = n25746 ^ n10061 ^ 1'b0 ;
  assign n26959 = n25154 ^ n22958 ^ 1'b0 ;
  assign n26960 = n24083 ^ n3437 ^ 1'b0 ;
  assign n26961 = n11448 | n26960 ;
  assign n26962 = n3098 | n26605 ;
  assign n26963 = n26962 ^ n26827 ^ 1'b0 ;
  assign n26968 = n942 & n22721 ;
  assign n26969 = n26968 ^ n1511 ^ 1'b0 ;
  assign n26964 = n4131 | n14877 ;
  assign n26965 = n6336 ^ n1003 ^ 1'b0 ;
  assign n26966 = n26964 & ~n26965 ;
  assign n26967 = n3947 & n26966 ;
  assign n26970 = n26969 ^ n26967 ^ 1'b0 ;
  assign n26971 = n7214 | n17999 ;
  assign n26972 = n4236 ^ n2805 ^ 1'b0 ;
  assign n26973 = n7674 & ~n26972 ;
  assign n26974 = n26973 ^ n4774 ^ 1'b0 ;
  assign n26975 = n26971 & ~n26974 ;
  assign n26976 = n268 & ~n16808 ;
  assign n26977 = n6090 & ~n15117 ;
  assign n26978 = n26977 ^ n3151 ^ 1'b0 ;
  assign n26979 = n20495 & ~n26978 ;
  assign n26980 = n3256 & ~n13841 ;
  assign n26981 = n12236 & n21306 ;
  assign n26982 = n3189 | n26981 ;
  assign n26983 = n12958 ^ n11523 ^ 1'b0 ;
  assign n26984 = n258 | n22981 ;
  assign n26985 = ~n3072 & n5453 ;
  assign n26986 = n26985 ^ n532 ^ 1'b0 ;
  assign n26987 = n252 & ~n26986 ;
  assign n26988 = n7625 & n26987 ;
  assign n26989 = n1033 & n25095 ;
  assign n26990 = n1975 & n21103 ;
  assign n26991 = ~n2209 & n4121 ;
  assign n26992 = ~n2904 & n20927 ;
  assign n26993 = n10340 & n26992 ;
  assign n26994 = n2010 & n26993 ;
  assign n26995 = n5106 & ~n26994 ;
  assign n26996 = n26994 & n26995 ;
  assign n26997 = n13363 & ~n26996 ;
  assign n26998 = n24147 & n26997 ;
  assign n26999 = n26998 ^ n22256 ^ 1'b0 ;
  assign n27000 = n79 | n2820 ;
  assign n27001 = n1184 | n2818 ;
  assign n27002 = n6250 & n27001 ;
  assign n27003 = ( n619 & ~n4115 ) | ( n619 & n27002 ) | ( ~n4115 & n27002 ) ;
  assign n27004 = n27000 & ~n27003 ;
  assign n27005 = n27004 ^ n5543 ^ 1'b0 ;
  assign n27006 = n10534 | n19033 ;
  assign n27007 = n2072 ^ n596 ^ 1'b0 ;
  assign n27008 = n16143 ^ n3658 ^ 1'b0 ;
  assign n27009 = n4927 | n27008 ;
  assign n27010 = n24696 ^ n12411 ^ n9566 ;
  assign n27011 = n7064 ^ n3859 ^ 1'b0 ;
  assign n27012 = n27011 ^ n19527 ^ 1'b0 ;
  assign n27013 = n27012 ^ n5827 ^ 1'b0 ;
  assign n27014 = ~n1366 & n13155 ;
  assign n27015 = n27014 ^ n15050 ^ 1'b0 ;
  assign n27016 = ~n15177 & n17135 ;
  assign n27017 = n19625 ^ n175 ^ 1'b0 ;
  assign n27018 = n10519 & ~n27017 ;
  assign n27019 = n3850 | n17603 ;
  assign n27020 = n13554 | n27019 ;
  assign n27021 = n21479 & n27020 ;
  assign n27022 = n27021 ^ n12673 ^ 1'b0 ;
  assign n27023 = n12757 & ~n17959 ;
  assign n27024 = n1613 & ~n3711 ;
  assign n27025 = ~n27023 & n27024 ;
  assign n27028 = n6348 ^ n2889 ^ 1'b0 ;
  assign n27029 = ~n5140 & n27028 ;
  assign n27030 = n27029 ^ n1392 ^ 1'b0 ;
  assign n27026 = ~n397 & n20244 ;
  assign n27027 = ~n534 & n27026 ;
  assign n27031 = n27030 ^ n27027 ^ 1'b0 ;
  assign n27032 = n9287 & ~n12902 ;
  assign n27033 = n27032 ^ n16462 ^ 1'b0 ;
  assign n27034 = n4273 & ~n27033 ;
  assign n27035 = n7529 | n8238 ;
  assign n27036 = n5065 & ~n27035 ;
  assign n27037 = n6671 | n27036 ;
  assign n27055 = n1469 & ~n2136 ;
  assign n27056 = n2136 & n27055 ;
  assign n27057 = n4996 | n27056 ;
  assign n27058 = n27057 ^ n9465 ^ 1'b0 ;
  assign n27038 = n1203 & ~n4734 ;
  assign n27039 = n4734 & n27038 ;
  assign n27040 = n278 | n27039 ;
  assign n27041 = n278 & ~n27040 ;
  assign n27042 = n5413 & n27041 ;
  assign n27043 = n22747 & n27042 ;
  assign n27044 = n1314 & n27043 ;
  assign n27048 = n508 | n1165 ;
  assign n27049 = n508 & ~n27048 ;
  assign n27050 = n4036 & ~n27049 ;
  assign n27051 = n27049 & n27050 ;
  assign n27045 = n1693 | n1935 ;
  assign n27046 = n1693 & ~n27045 ;
  assign n27047 = n27046 ^ n24513 ^ 1'b0 ;
  assign n27052 = n27051 ^ n27047 ^ 1'b0 ;
  assign n27053 = ~n27044 & n27052 ;
  assign n27054 = n9512 & n27053 ;
  assign n27059 = n27058 ^ n27054 ^ 1'b0 ;
  assign n27060 = n5846 ^ n4275 ^ 1'b0 ;
  assign n27061 = ~n364 & n27060 ;
  assign n27062 = n3209 & n3239 ;
  assign n27063 = n27062 ^ n2828 ^ 1'b0 ;
  assign n27064 = n1688 & ~n27063 ;
  assign n27065 = n27064 ^ n18107 ^ 1'b0 ;
  assign n27066 = n1693 & ~n7007 ;
  assign n27067 = n6251 & n27066 ;
  assign n27068 = n14771 ^ n6168 ^ 1'b0 ;
  assign n27069 = n27068 ^ n1372 ^ 1'b0 ;
  assign n27070 = n8067 | n27069 ;
  assign n27071 = n27067 | n27070 ;
  assign n27072 = n1564 & ~n2495 ;
  assign n27073 = n5794 & n27072 ;
  assign n27074 = ~n22161 & n27073 ;
  assign n27075 = ~n17361 & n27074 ;
  assign n27076 = n14975 ^ n2470 ^ 1'b0 ;
  assign n27077 = n18621 & n21082 ;
  assign n27078 = n7413 ^ n86 ^ 1'b0 ;
  assign n27079 = x6 & n1355 ;
  assign n27080 = n27079 ^ n12731 ^ 1'b0 ;
  assign n27081 = n27080 ^ n3074 ^ 1'b0 ;
  assign n27082 = n17221 ^ n8654 ^ 1'b0 ;
  assign n27083 = n25051 ^ n12206 ^ n814 ;
  assign n27084 = n4407 | n4766 ;
  assign n27085 = n27084 ^ n26986 ^ 1'b0 ;
  assign n27086 = n4680 & ~n27085 ;
  assign n27087 = n12732 ^ n6901 ^ 1'b0 ;
  assign n27088 = n4772 & ~n27087 ;
  assign n27089 = n24544 ^ n1631 ^ 1'b0 ;
  assign n27090 = ~n8054 & n11845 ;
  assign n27091 = n27090 ^ n10461 ^ 1'b0 ;
  assign n27092 = n23702 ^ n4943 ^ 1'b0 ;
  assign n27093 = ~n16190 & n21987 ;
  assign n27094 = n784 & n13629 ;
  assign n27095 = n754 ^ n322 ^ 1'b0 ;
  assign n27096 = n8107 & n10680 ;
  assign n27097 = n19876 ^ n4575 ^ 1'b0 ;
  assign n27098 = ~n27096 & n27097 ;
  assign n27099 = n27098 ^ n19902 ^ 1'b0 ;
  assign n27100 = n10004 | n27099 ;
  assign n27101 = n5567 & n23601 ;
  assign n27102 = n27100 & n27101 ;
  assign n27103 = n13362 | n13727 ;
  assign n27104 = n1699 & ~n25025 ;
  assign n27105 = n27104 ^ n8158 ^ 1'b0 ;
  assign n27106 = n16985 ^ n3726 ^ 1'b0 ;
  assign n27107 = ~n12366 & n24669 ;
  assign n27108 = n6165 | n27107 ;
  assign n27109 = n1135 | n4546 ;
  assign n27110 = n323 & n22279 ;
  assign n27111 = n2774 | n10313 ;
  assign n27112 = n784 | n27111 ;
  assign n27113 = ~n8387 & n27112 ;
  assign n27114 = ~n1924 & n27113 ;
  assign n27115 = n8977 ^ n1117 ^ 1'b0 ;
  assign n27116 = n5953 & n27115 ;
  assign n27117 = n7096 & ~n27116 ;
  assign n27118 = n573 | n10067 ;
  assign n27119 = n8630 & ~n27118 ;
  assign n27120 = n24611 | n27119 ;
  assign n27121 = n9810 | n10414 ;
  assign n27122 = n27121 ^ n15859 ^ 1'b0 ;
  assign n27123 = ( n7304 & n20058 ) | ( n7304 & n27122 ) | ( n20058 & n27122 ) ;
  assign n27124 = ~n3297 & n11040 ;
  assign n27125 = n24222 | n27124 ;
  assign n27126 = n1588 | n27125 ;
  assign n27127 = ~n330 & n16964 ;
  assign n27128 = n27127 ^ n10823 ^ 1'b0 ;
  assign n27129 = n6667 ^ n3720 ^ n1878 ;
  assign n27130 = n257 & n10025 ;
  assign n27131 = n1421 & n27130 ;
  assign n27132 = n27131 ^ n14144 ^ 1'b0 ;
  assign n27133 = n18716 & ~n27132 ;
  assign n27134 = n24585 & n27133 ;
  assign n27135 = n27134 ^ n22974 ^ 1'b0 ;
  assign n27136 = ~n5147 & n23328 ;
  assign n27137 = ~n7388 & n14432 ;
  assign n27138 = n27137 ^ n22474 ^ 1'b0 ;
  assign n27139 = n6449 & n22979 ;
  assign n27140 = n3997 & n14675 ;
  assign n27141 = n17948 ^ n10429 ^ 1'b0 ;
  assign n27142 = n2075 & ~n27141 ;
  assign n27143 = n27142 ^ n1235 ^ 1'b0 ;
  assign n27144 = n16082 | n27143 ;
  assign n27145 = ~n6595 & n18587 ;
  assign n27146 = n3535 & ~n13534 ;
  assign n27147 = n5461 ^ n1090 ^ 1'b0 ;
  assign n27148 = ~n382 & n27147 ;
  assign n27151 = ( n2183 & n5288 ) | ( n2183 & n12472 ) | ( n5288 & n12472 ) ;
  assign n27149 = n12877 ^ n1939 ^ 1'b0 ;
  assign n27150 = n23783 & n27149 ;
  assign n27152 = n27151 ^ n27150 ^ 1'b0 ;
  assign n27153 = ( n17537 & ~n27148 ) | ( n17537 & n27152 ) | ( ~n27148 & n27152 ) ;
  assign n27154 = n13154 ^ n419 ^ 1'b0 ;
  assign n27155 = n23767 | n27154 ;
  assign n27156 = n1081 | n27155 ;
  assign n27161 = n22076 ^ n7104 ^ 1'b0 ;
  assign n27162 = n6277 & ~n27161 ;
  assign n27157 = n4105 & ~n4236 ;
  assign n27158 = n27157 ^ n3015 ^ 1'b0 ;
  assign n27159 = n7271 & n16160 ;
  assign n27160 = ~n27158 & n27159 ;
  assign n27163 = n27162 ^ n27160 ^ 1'b0 ;
  assign n27164 = n218 | n27163 ;
  assign n27165 = n1668 & n3417 ;
  assign n27166 = n22853 ^ n7697 ^ 1'b0 ;
  assign n27167 = ~n27165 & n27166 ;
  assign n27168 = ~n1425 & n9319 ;
  assign n27169 = n1026 & ~n2377 ;
  assign n27170 = n3589 | n27169 ;
  assign n27171 = n25243 ^ n4660 ^ 1'b0 ;
  assign n27172 = ~n18330 & n18510 ;
  assign n27173 = n17001 & ~n18192 ;
  assign n27174 = ~n8037 & n13992 ;
  assign n27175 = n6959 & n27174 ;
  assign n27176 = n3131 | n23982 ;
  assign n27177 = n14469 | n27176 ;
  assign n27178 = n13777 ^ n12269 ^ 1'b0 ;
  assign n27179 = n2217 | n2912 ;
  assign n27180 = n2912 & ~n27179 ;
  assign n27181 = n2311 & ~n27180 ;
  assign n27182 = n27180 & n27181 ;
  assign n27183 = n8594 & n11895 ;
  assign n27184 = n7736 & n27183 ;
  assign n27185 = n4874 | n27184 ;
  assign n27186 = n27182 & ~n27185 ;
  assign n27187 = n22343 ^ n18275 ^ 1'b0 ;
  assign n27188 = n12027 ^ n6933 ^ 1'b0 ;
  assign n27189 = ~n471 & n10736 ;
  assign n27190 = n27189 ^ n11453 ^ 1'b0 ;
  assign n27191 = n8681 & ~n27190 ;
  assign n27192 = n27191 ^ n2283 ^ 1'b0 ;
  assign n27193 = n66 | n25179 ;
  assign n27198 = n478 ^ n354 ^ 1'b0 ;
  assign n27197 = n2248 & ~n2485 ;
  assign n27199 = n27198 ^ n27197 ^ 1'b0 ;
  assign n27194 = n4400 & ~n6082 ;
  assign n27195 = n7088 | n27194 ;
  assign n27196 = n27194 & ~n27195 ;
  assign n27200 = n27199 ^ n27196 ^ n10705 ;
  assign n27201 = n653 & ~n7119 ;
  assign n27202 = ~n117 & n27201 ;
  assign n27203 = n27202 ^ n20752 ^ 1'b0 ;
  assign n27205 = ~n713 & n8534 ;
  assign n27206 = n27205 ^ n11682 ^ 1'b0 ;
  assign n27204 = n12072 | n14204 ;
  assign n27207 = n27206 ^ n27204 ^ 1'b0 ;
  assign n27208 = n4809 & ~n22230 ;
  assign n27209 = n4970 & ~n27208 ;
  assign n27210 = n17339 | n18921 ;
  assign n27211 = n17326 | n27210 ;
  assign n27212 = n2031 | n27211 ;
  assign n27213 = n19889 ^ n3597 ^ 1'b0 ;
  assign n27214 = ~n17 & n154 ;
  assign n27215 = n27214 ^ n514 ^ 1'b0 ;
  assign n27216 = ~n23894 & n27215 ;
  assign n27217 = n27216 ^ n16910 ^ 1'b0 ;
  assign n27218 = n3095 | n18290 ;
  assign n27219 = n3749 & ~n27218 ;
  assign n27220 = n8679 | n11343 ;
  assign n27221 = n12972 & n27220 ;
  assign n27222 = n27221 ^ n1848 ^ 1'b0 ;
  assign n27223 = ~n27219 & n27222 ;
  assign n27224 = n27223 ^ n6359 ^ 1'b0 ;
  assign n27225 = n7514 | n12982 ;
  assign n27226 = n507 | n27225 ;
  assign n27227 = ~n20999 & n26843 ;
  assign n27228 = n12240 ^ x0 ^ 1'b0 ;
  assign n27229 = n5927 & ~n27228 ;
  assign n27230 = ~n27227 & n27229 ;
  assign n27231 = n3882 & ~n15405 ;
  assign n27232 = ~n13446 & n27231 ;
  assign n27233 = n539 | n27232 ;
  assign n27234 = ~n2472 & n27233 ;
  assign n27235 = n10097 & ~n27234 ;
  assign n27236 = n7265 | n20103 ;
  assign n27237 = n14804 | n19963 ;
  assign n27238 = ~n7071 & n27237 ;
  assign n27239 = ~n7425 & n27238 ;
  assign n27240 = n8685 & n27239 ;
  assign n27241 = n4882 ^ n322 ^ 1'b0 ;
  assign n27242 = ~n2792 & n27241 ;
  assign n27243 = n24477 ^ n3643 ^ 1'b0 ;
  assign n27244 = n2004 | n27243 ;
  assign n27246 = n9197 & ~n27219 ;
  assign n27245 = n3100 & ~n24919 ;
  assign n27247 = n27246 ^ n27245 ^ 1'b0 ;
  assign n27248 = n23746 ^ n4655 ^ 1'b0 ;
  assign n27249 = n27247 & n27248 ;
  assign n27250 = n55 & ~n236 ;
  assign n27251 = n27250 ^ n6753 ^ 1'b0 ;
  assign n27252 = n14089 ^ n6376 ^ 1'b0 ;
  assign n27253 = ~n15469 & n24672 ;
  assign n27254 = n27253 ^ n1226 ^ 1'b0 ;
  assign n27255 = ~n27252 & n27254 ;
  assign n27256 = n2593 | n15336 ;
  assign n27257 = n2361 & ~n14198 ;
  assign n27258 = n16729 & n17691 ;
  assign n27259 = n27258 ^ n14006 ^ 1'b0 ;
  assign n27260 = n5733 | n13258 ;
  assign n27261 = n4551 | n11626 ;
  assign n27262 = n27261 ^ n930 ^ 1'b0 ;
  assign n27263 = n736 & n11970 ;
  assign n27264 = n27263 ^ n3327 ^ 1'b0 ;
  assign n27265 = n27264 ^ n2644 ^ 1'b0 ;
  assign n27266 = n27262 & n27265 ;
  assign n27267 = n982 & n15263 ;
  assign n27268 = n4061 & n27267 ;
  assign n27269 = n17127 ^ n318 ^ 1'b0 ;
  assign n27270 = ~n27268 & n27269 ;
  assign n27271 = n2032 & n10655 ;
  assign n27272 = n507 | n10344 ;
  assign n27273 = n6530 ^ n3447 ^ 1'b0 ;
  assign n27274 = ( ~n7731 & n14440 ) | ( ~n7731 & n27273 ) | ( n14440 & n27273 ) ;
  assign n27275 = n27274 ^ n22899 ^ 1'b0 ;
  assign n27276 = n6329 & ~n27275 ;
  assign n27277 = n6301 & n27276 ;
  assign n27278 = n18316 ^ n10554 ^ 1'b0 ;
  assign n27279 = x8 & n17207 ;
  assign n27280 = n7395 & ~n7582 ;
  assign n27281 = ~n18566 & n27280 ;
  assign n27282 = ~n1790 & n9815 ;
  assign n27283 = n27282 ^ n339 ^ 1'b0 ;
  assign n27284 = n3532 & n27283 ;
  assign n27285 = n5812 ^ n5322 ^ 1'b0 ;
  assign n27286 = n1560 | n27285 ;
  assign n27287 = n27284 & n27286 ;
  assign n27288 = n8842 & n8885 ;
  assign n27289 = n5947 ^ n1350 ^ 1'b0 ;
  assign n27290 = n24127 & ~n27289 ;
  assign n27291 = ~n4760 & n27290 ;
  assign n27292 = n3262 ^ n241 ^ 1'b0 ;
  assign n27293 = n27291 | n27292 ;
  assign n27294 = n1300 | n27293 ;
  assign n27295 = ~n12028 & n27294 ;
  assign n27296 = ~n13074 & n27295 ;
  assign n27297 = n11427 ^ n86 ^ 1'b0 ;
  assign n27298 = n10447 & ~n22556 ;
  assign n27299 = n5356 | n15176 ;
  assign n27300 = n27299 ^ n14170 ^ 1'b0 ;
  assign n27301 = n817 | n2261 ;
  assign n27302 = n914 | n22088 ;
  assign n27303 = n9872 ^ n659 ^ 1'b0 ;
  assign n27304 = n15438 & n27303 ;
  assign n27305 = ( n159 & n15227 ) | ( n159 & ~n27304 ) | ( n15227 & ~n27304 ) ;
  assign n27306 = ( n12201 & ~n13428 ) | ( n12201 & n27305 ) | ( ~n13428 & n27305 ) ;
  assign n27307 = n2919 ^ n2874 ^ 1'b0 ;
  assign n27308 = n2455 | n27307 ;
  assign n27309 = n5943 | n26972 ;
  assign n27310 = n27308 & ~n27309 ;
  assign n27311 = n19641 ^ n3851 ^ 1'b0 ;
  assign n27312 = ~n14147 & n17284 ;
  assign n27313 = n9751 & n27312 ;
  assign n27314 = n7792 & n12993 ;
  assign n27315 = n5529 ^ n4590 ^ 1'b0 ;
  assign n27316 = n2194 & ~n10105 ;
  assign n27317 = n8392 ^ n4327 ^ 1'b0 ;
  assign n27318 = n16318 | n27317 ;
  assign n27319 = n11508 & ~n26680 ;
  assign n27320 = ~n26959 & n27319 ;
  assign n27321 = ~n5241 & n21740 ;
  assign n27322 = n27321 ^ n13377 ^ 1'b0 ;
  assign n27323 = n22287 & ~n27322 ;
  assign n27324 = n3941 ^ n1008 ^ 1'b0 ;
  assign n27325 = n4273 & ~n27324 ;
  assign n27326 = n1246 ^ n135 ^ 1'b0 ;
  assign n27327 = n8769 | n10815 ;
  assign n27328 = n16100 & n21614 ;
  assign n27329 = ~n1100 & n12366 ;
  assign n27330 = n6244 & n22947 ;
  assign n27332 = n8156 ^ n4357 ^ 1'b0 ;
  assign n27331 = n5258 & n20566 ;
  assign n27333 = n27332 ^ n27331 ^ 1'b0 ;
  assign n27334 = n7093 & ~n16803 ;
  assign n27335 = n11379 ^ n2814 ^ 1'b0 ;
  assign n27336 = n1235 ^ n765 ^ 1'b0 ;
  assign n27337 = n8637 & n27336 ;
  assign n27338 = ~n27335 & n27337 ;
  assign n27339 = n27338 ^ n9564 ^ 1'b0 ;
  assign n27340 = n1772 | n7664 ;
  assign n27341 = n770 & ~n8628 ;
  assign n27342 = n2930 & n27341 ;
  assign n27343 = x9 & n9649 ;
  assign n27344 = n11874 & n27343 ;
  assign n27345 = n24770 ^ n3516 ^ 1'b0 ;
  assign n27346 = ~n14423 & n27345 ;
  assign n27347 = n27346 ^ n8219 ^ 1'b0 ;
  assign n27348 = n1292 & n4132 ;
  assign n27349 = ~n8541 & n27348 ;
  assign n27350 = n4893 | n27349 ;
  assign n27351 = n4400 & ~n15103 ;
  assign n27352 = ~n11401 & n27351 ;
  assign n27353 = n18471 ^ n8950 ^ 1'b0 ;
  assign n27354 = n724 & ~n25406 ;
  assign n27355 = ~n3211 & n24353 ;
  assign n27356 = ( n4639 & n12046 ) | ( n4639 & n13015 ) | ( n12046 & n13015 ) ;
  assign n27357 = n13058 ^ n328 ^ 1'b0 ;
  assign n27358 = ~n5265 & n8197 ;
  assign n27359 = ~n26982 & n27358 ;
  assign n27360 = n1979 & ~n12865 ;
  assign n27361 = ~n6643 & n27360 ;
  assign n27362 = n68 | n2956 ;
  assign n27363 = ( ~n594 & n10527 ) | ( ~n594 & n17944 ) | ( n10527 & n17944 ) ;
  assign n27364 = n719 & n27363 ;
  assign n27365 = n27364 ^ n2657 ^ 1'b0 ;
  assign n27366 = n27362 | n27365 ;
  assign n27367 = n7397 ^ n770 ^ 1'b0 ;
  assign n27368 = n27367 ^ n7704 ^ 1'b0 ;
  assign n27369 = ~n6387 & n7013 ;
  assign n27370 = ~n24310 & n27369 ;
  assign n27371 = ~n883 & n6097 ;
  assign n27372 = n27371 ^ n2921 ^ 1'b0 ;
  assign n27373 = n22227 ^ n13337 ^ 1'b0 ;
  assign n27374 = ~n21363 & n27373 ;
  assign n27375 = n8056 ^ n7615 ^ 1'b0 ;
  assign n27377 = n16990 ^ n938 ^ 1'b0 ;
  assign n27378 = n985 & ~n2948 ;
  assign n27379 = ~n27377 & n27378 ;
  assign n27380 = n27379 ^ n13747 ^ 1'b0 ;
  assign n27381 = n11415 & n27380 ;
  assign n27376 = n1041 | n11360 ;
  assign n27382 = n27381 ^ n27376 ^ 1'b0 ;
  assign n27383 = n15769 ^ n3292 ^ 1'b0 ;
  assign n27384 = ~n8803 & n27383 ;
  assign n27385 = n18187 & ~n27384 ;
  assign n27386 = n827 & n20104 ;
  assign n27387 = n3405 ^ n2862 ^ 1'b0 ;
  assign n27388 = n4332 & ~n27387 ;
  assign n27389 = ~n13585 & n18121 ;
  assign n27390 = n11384 & ~n12297 ;
  assign n27391 = n27390 ^ n9659 ^ 1'b0 ;
  assign n27392 = n6061 & ~n20652 ;
  assign n27393 = n27391 | n27392 ;
  assign n27394 = ~n10850 & n18326 ;
  assign n27395 = n23992 & ~n27394 ;
  assign n27396 = n15027 ^ n8107 ^ n3049 ;
  assign n27397 = ~n17667 & n27396 ;
  assign n27398 = n27397 ^ n10644 ^ 1'b0 ;
  assign n27399 = n16311 & ~n27398 ;
  assign n27400 = n20615 ^ n291 ^ 1'b0 ;
  assign n27401 = n2261 & ~n6442 ;
  assign n27402 = n27401 ^ n27011 ^ 1'b0 ;
  assign n27403 = n27400 & ~n27402 ;
  assign n27404 = n2849 & ~n22914 ;
  assign n27405 = n27404 ^ n10083 ^ 1'b0 ;
  assign n27406 = n270 | n1868 ;
  assign n27407 = n4279 & n25263 ;
  assign n27408 = ~n702 & n10096 ;
  assign n27409 = ~n3277 & n27408 ;
  assign n27410 = n17935 & n27409 ;
  assign n27411 = n16979 & n17921 ;
  assign n27412 = n19117 ^ n246 ^ 1'b0 ;
  assign n27413 = n1626 ^ n104 ^ 1'b0 ;
  assign n27414 = n4807 | n21303 ;
  assign n27415 = n25431 ^ n24619 ^ 1'b0 ;
  assign n27416 = ~n27414 & n27415 ;
  assign n27417 = n24308 ^ n9145 ^ 1'b0 ;
  assign n27418 = n5303 | n27417 ;
  assign n27419 = n12409 & ~n27418 ;
  assign n27420 = n16913 & n24350 ;
  assign n27421 = ~n23479 & n27420 ;
  assign n27422 = n9768 & ~n27421 ;
  assign n27423 = n9043 & n11272 ;
  assign n27424 = ~n14739 & n27423 ;
  assign n27425 = n27424 ^ n5918 ^ 1'b0 ;
  assign n27426 = n12514 ^ n6154 ^ 1'b0 ;
  assign n27427 = n1856 & ~n5394 ;
  assign n27428 = ~n2639 & n15642 ;
  assign n27429 = ~n27427 & n27428 ;
  assign n27430 = ~n2124 & n3655 ;
  assign n27431 = ~n23279 & n27430 ;
  assign n27435 = n457 ^ n342 ^ 1'b0 ;
  assign n27436 = n6114 ^ n1673 ^ 1'b0 ;
  assign n27437 = n27435 | n27436 ;
  assign n27433 = n4361 & ~n5393 ;
  assign n27432 = n2418 & ~n15933 ;
  assign n27434 = n27433 ^ n27432 ^ 1'b0 ;
  assign n27438 = n27437 ^ n27434 ^ 1'b0 ;
  assign n27439 = ~n22762 & n27438 ;
  assign n27440 = n27431 | n27439 ;
  assign n27441 = n255 | n951 ;
  assign n27442 = ~n13707 & n27441 ;
  assign n27443 = n27442 ^ n6631 ^ 1'b0 ;
  assign n27444 = n7060 & n20218 ;
  assign n27445 = n27444 ^ n5903 ^ 1'b0 ;
  assign n27446 = n628 & ~n27445 ;
  assign n27447 = n26108 ^ n1844 ^ 1'b0 ;
  assign n27448 = n24713 | n27447 ;
  assign n27449 = n27446 | n27448 ;
  assign n27450 = n27112 ^ n24874 ^ 1'b0 ;
  assign n27451 = n7185 & ~n27450 ;
  assign n27452 = n5412 ^ n4158 ^ 1'b0 ;
  assign n27453 = n4936 & n7039 ;
  assign n27454 = ~n7783 & n27453 ;
  assign n27455 = n27454 ^ n4964 ^ 1'b0 ;
  assign n27456 = ~n15879 & n27455 ;
  assign n27457 = ~n2517 & n25125 ;
  assign n27458 = ~n7709 & n27457 ;
  assign n27459 = ~n9273 & n27458 ;
  assign n27460 = n27459 ^ n7943 ^ 1'b0 ;
  assign n27461 = ~n15117 & n27460 ;
  assign n27462 = n27461 ^ n9614 ^ 1'b0 ;
  assign n27463 = n20097 & n27462 ;
  assign n27464 = n9574 | n15954 ;
  assign n27465 = n3099 & ~n18095 ;
  assign n27466 = n27464 & n27465 ;
  assign n27467 = n14254 & ~n22966 ;
  assign n27468 = ~n9931 & n27467 ;
  assign n27469 = n10940 & ~n16081 ;
  assign n27470 = n8269 & ~n15931 ;
  assign n27471 = ~n3012 & n27470 ;
  assign n27472 = n27471 ^ n642 ^ 1'b0 ;
  assign n27473 = n5655 ^ n2930 ^ 1'b0 ;
  assign n27474 = ~n7431 & n27473 ;
  assign n27475 = n5510 & ~n8341 ;
  assign n27476 = n27475 ^ n9635 ^ 1'b0 ;
  assign n27477 = n27476 ^ n1350 ^ 1'b0 ;
  assign n27478 = n27474 & ~n27477 ;
  assign n27479 = n9846 ^ n212 ^ 1'b0 ;
  assign n27480 = n9209 & n16030 ;
  assign n27481 = n10982 & n27480 ;
  assign n27482 = n68 | n17180 ;
  assign n27483 = n7875 & n27482 ;
  assign n27484 = n213 & ~n27483 ;
  assign n27485 = x3 | n17703 ;
  assign n27486 = n26020 & ~n27485 ;
  assign n27487 = n22100 & ~n27486 ;
  assign n27488 = n27487 ^ n7943 ^ 1'b0 ;
  assign n27489 = n4311 | n18532 ;
  assign n27490 = n1934 & n8115 ;
  assign n27491 = n325 & n27490 ;
  assign n27492 = ~n15766 & n27491 ;
  assign n27493 = n27492 ^ n14165 ^ 1'b0 ;
  assign n27494 = n23336 | n27493 ;
  assign n27495 = n1019 ^ n82 ^ 1'b0 ;
  assign n27496 = n24569 & ~n27495 ;
  assign n27497 = n13529 & n27496 ;
  assign n27498 = n18839 ^ n8071 ^ 1'b0 ;
  assign n27499 = n25489 & ~n27498 ;
  assign n27500 = n62 | n3216 ;
  assign n27501 = n27500 ^ n9850 ^ 1'b0 ;
  assign n27502 = n13803 ^ n4321 ^ 1'b0 ;
  assign n27503 = n27502 ^ n26493 ^ 1'b0 ;
  assign n27504 = n15336 & n17191 ;
  assign n27505 = n2315 | n16981 ;
  assign n27506 = n7775 & ~n27288 ;
  assign n27507 = ~n19144 & n27506 ;
  assign n27508 = n11374 & ~n15055 ;
  assign n27509 = n343 & n2513 ;
  assign n27510 = n10475 & n14392 ;
  assign n27511 = ~n9155 & n11317 ;
  assign n27512 = n8632 & n27511 ;
  assign n27513 = n861 & ~n6224 ;
  assign n27514 = n8011 & n27513 ;
  assign n27515 = n27514 ^ n6068 ^ 1'b0 ;
  assign n27516 = ~n27512 & n27515 ;
  assign n27517 = ( n27509 & n27510 ) | ( n27509 & n27516 ) | ( n27510 & n27516 ) ;
  assign n27518 = ~n458 & n11535 ;
  assign n27519 = n1217 ^ n231 ^ 1'b0 ;
  assign n27520 = n5501 & ~n27519 ;
  assign n27521 = n20276 & n27520 ;
  assign n27522 = n23500 & n27521 ;
  assign n27523 = n27522 ^ n19922 ^ 1'b0 ;
  assign n27524 = n10818 & n10837 ;
  assign n27525 = n335 & n3178 ;
  assign n27526 = n4533 ^ n2637 ^ 1'b0 ;
  assign n27527 = n27525 & ~n27526 ;
  assign n27528 = n1712 & ~n2268 ;
  assign n27529 = n7231 ^ n3485 ^ 1'b0 ;
  assign n27530 = ~n9507 & n27529 ;
  assign n27531 = n11160 ^ n9634 ^ 1'b0 ;
  assign n27532 = n10358 & n27531 ;
  assign n27533 = n9593 & ~n23536 ;
  assign n27534 = n27533 ^ n18150 ^ 1'b0 ;
  assign n27535 = n2774 | n4485 ;
  assign n27536 = ~n8810 & n9335 ;
  assign n27537 = n27536 ^ n18494 ^ 1'b0 ;
  assign n27538 = n5758 | n27537 ;
  assign n27539 = n27535 & ~n27538 ;
  assign n27540 = n1193 | n11039 ;
  assign n27541 = n27540 ^ n10500 ^ n1774 ;
  assign n27542 = n4914 | n21346 ;
  assign n27543 = n1630 ^ n1040 ^ 1'b0 ;
  assign n27544 = ~n122 & n27543 ;
  assign n27545 = n7427 | n12292 ;
  assign n27546 = n4794 & ~n27545 ;
  assign n27547 = ~n21155 & n22159 ;
  assign n27548 = ~n557 & n27547 ;
  assign n27549 = n9492 ^ n5503 ^ 1'b0 ;
  assign n27550 = n1687 ^ n1260 ^ 1'b0 ;
  assign n27551 = n2484 & n27550 ;
  assign n27552 = n27551 ^ n3476 ^ 1'b0 ;
  assign n27553 = ~n8360 & n27552 ;
  assign n27554 = n27553 ^ n14712 ^ 1'b0 ;
  assign n27555 = ( n36 & n724 ) | ( n36 & n6904 ) | ( n724 & n6904 ) ;
  assign n27556 = n16799 ^ n5336 ^ 1'b0 ;
  assign n27557 = ~n1909 & n20113 ;
  assign n27558 = n23439 ^ n5206 ^ 1'b0 ;
  assign n27559 = ~n21816 & n27558 ;
  assign n27560 = n18052 ^ n13073 ^ 1'b0 ;
  assign n27561 = n27559 & n27560 ;
  assign n27562 = n22905 ^ n20490 ^ 1'b0 ;
  assign n27563 = n4582 ^ n4060 ^ 1'b0 ;
  assign n27564 = n27011 | n27563 ;
  assign n27565 = n7263 ^ n2513 ^ n1879 ;
  assign n27566 = n27564 | n27565 ;
  assign n27567 = n27566 ^ n5232 ^ 1'b0 ;
  assign n27568 = n709 & ~n1267 ;
  assign n27569 = n14306 | n27568 ;
  assign n27570 = n27569 ^ n19887 ^ 1'b0 ;
  assign n27571 = n9852 & n27570 ;
  assign n27572 = n15873 & n27571 ;
  assign n27573 = n23472 & ~n27572 ;
  assign n27574 = n21548 ^ n722 ^ 1'b0 ;
  assign n27575 = n27574 ^ n758 ^ 1'b0 ;
  assign n27576 = ~n11061 & n14102 ;
  assign n27577 = ~n19976 & n27576 ;
  assign n27578 = n5278 & ~n9359 ;
  assign n27579 = n11731 & n14803 ;
  assign n27580 = n1109 | n15368 ;
  assign n27581 = n27580 ^ n2167 ^ 1'b0 ;
  assign n27582 = ~n4899 & n22999 ;
  assign n27583 = n2093 | n27582 ;
  assign n27585 = n16305 ^ n11528 ^ n954 ;
  assign n27584 = ~n741 & n21111 ;
  assign n27586 = n27585 ^ n27584 ^ 1'b0 ;
  assign n27588 = n4850 ^ n3697 ^ n3053 ;
  assign n27589 = ~n6028 & n27588 ;
  assign n27590 = ~n3506 & n27589 ;
  assign n27591 = n15707 & n27590 ;
  assign n27587 = ~n1898 & n3685 ;
  assign n27592 = n27591 ^ n27587 ^ 1'b0 ;
  assign n27593 = ~n685 & n7954 ;
  assign n27594 = n310 & n27593 ;
  assign n27595 = n17303 ^ n10480 ^ 1'b0 ;
  assign n27596 = n4115 | n27595 ;
  assign n27597 = n20795 ^ n11690 ^ 1'b0 ;
  assign n27598 = n105 & n9588 ;
  assign n27599 = n24006 & n27598 ;
  assign n27600 = n7581 | n22610 ;
  assign n27601 = n10766 & ~n14228 ;
  assign n27602 = ~n3487 & n27601 ;
  assign n27603 = n27602 ^ n25630 ^ 1'b0 ;
  assign n27604 = n1737 | n19790 ;
  assign n27605 = ~n6306 & n27604 ;
  assign n27606 = n27605 ^ n18059 ^ n4491 ;
  assign n27607 = n20130 & n27606 ;
  assign n27608 = n3423 & n27607 ;
  assign n27609 = n23783 ^ n2254 ^ 1'b0 ;
  assign n27610 = n7865 & ~n15050 ;
  assign n27611 = n16966 & ~n27610 ;
  assign n27612 = ~n804 & n27611 ;
  assign n27613 = ~n101 & n9707 ;
  assign n27614 = n813 | n27613 ;
  assign n27615 = n4549 | n13519 ;
  assign n27616 = n10756 & ~n27615 ;
  assign n27617 = ~n12641 & n27616 ;
  assign n27618 = n16472 ^ n8915 ^ 1'b0 ;
  assign n27619 = n10753 ^ n6070 ^ 1'b0 ;
  assign n27620 = ~n10968 & n27619 ;
  assign n27621 = ( n1845 & ~n6971 ) | ( n1845 & n27620 ) | ( ~n6971 & n27620 ) ;
  assign n27622 = n16158 ^ n419 ^ 1'b0 ;
  assign n27623 = n16124 | n27622 ;
  assign n27624 = n11338 & ~n27623 ;
  assign n27625 = n25661 & n27624 ;
  assign n27626 = ~n27621 & n27625 ;
  assign n27627 = n294 & ~n5756 ;
  assign n27628 = n27627 ^ n12269 ^ 1'b0 ;
  assign n27629 = n5421 ^ n2909 ^ 1'b0 ;
  assign n27630 = ( n4883 & ~n11064 ) | ( n4883 & n27629 ) | ( ~n11064 & n27629 ) ;
  assign n27631 = n5623 & n14534 ;
  assign n27632 = n27631 ^ n7825 ^ 1'b0 ;
  assign n27633 = n27630 & n27632 ;
  assign n27634 = ~n307 & n2491 ;
  assign n27635 = n27634 ^ n6272 ^ 1'b0 ;
  assign n27636 = n27635 ^ n22166 ^ 1'b0 ;
  assign n27637 = ~n23045 & n27636 ;
  assign n27638 = n24043 ^ n19681 ^ 1'b0 ;
  assign n27639 = n5370 & n7814 ;
  assign n27640 = n27639 ^ n12556 ^ 1'b0 ;
  assign n27641 = n865 & ~n27640 ;
  assign n27642 = n27641 ^ n6645 ^ 1'b0 ;
  assign n27643 = n17104 ^ n3382 ^ 1'b0 ;
  assign n27644 = n10822 ^ n5085 ^ 1'b0 ;
  assign n27645 = ~n3645 & n13709 ;
  assign n27646 = n27645 ^ n11745 ^ 1'b0 ;
  assign n27647 = n16786 ^ n4897 ^ 1'b0 ;
  assign n27648 = ~n2813 & n27647 ;
  assign n27649 = n17694 & n27648 ;
  assign n27650 = ~n745 & n27649 ;
  assign n27651 = ~n25850 & n27650 ;
  assign n27652 = n12210 ^ n9548 ^ 1'b0 ;
  assign n27653 = n13876 | n18058 ;
  assign n27654 = n2714 & ~n13064 ;
  assign n27655 = n18925 ^ n4852 ^ 1'b0 ;
  assign n27656 = n3442 | n27655 ;
  assign n27657 = n10031 & ~n15760 ;
  assign n27658 = n1050 | n4733 ;
  assign n27659 = n21764 & ~n27658 ;
  assign n27660 = n4851 | n8705 ;
  assign n27661 = n27660 ^ n16910 ^ 1'b0 ;
  assign n27662 = n19486 ^ n2288 ^ 1'b0 ;
  assign n27663 = n4245 & ~n27662 ;
  assign n27664 = n656 | n1015 ;
  assign n27665 = n27664 ^ n20828 ^ 1'b0 ;
  assign n27666 = n24816 & n27665 ;
  assign n27667 = n8730 & ~n19049 ;
  assign n27668 = ~n254 & n27667 ;
  assign n27669 = ( n27663 & n27666 ) | ( n27663 & ~n27668 ) | ( n27666 & ~n27668 ) ;
  assign n27670 = n5295 | n15605 ;
  assign n27671 = n14037 & n14321 ;
  assign n27672 = n27670 & ~n27671 ;
  assign n27673 = n27672 ^ n27302 ^ 1'b0 ;
  assign n27674 = n12740 & n16523 ;
  assign n27675 = n27674 ^ n1812 ^ 1'b0 ;
  assign n27676 = ~n14046 & n17750 ;
  assign n27677 = n26842 ^ n3773 ^ 1'b0 ;
  assign n27678 = n27676 & n27677 ;
  assign n27679 = n25505 | n27206 ;
  assign n27680 = n403 | n5205 ;
  assign n27681 = n27680 ^ n1198 ^ 1'b0 ;
  assign n27682 = n27681 ^ n15103 ^ 1'b0 ;
  assign n27683 = n27679 | n27682 ;
  assign n27684 = ~n11586 & n11936 ;
  assign n27685 = n879 | n18372 ;
  assign n27686 = n12014 ^ n9039 ^ 1'b0 ;
  assign n27687 = n12020 & n25684 ;
  assign n27688 = n27687 ^ n11656 ^ 1'b0 ;
  assign n27689 = n15718 & n27688 ;
  assign n27690 = n177 | n17484 ;
  assign n27691 = n3382 & ~n21394 ;
  assign n27692 = n4482 | n4842 ;
  assign n27693 = n3646 | n27692 ;
  assign n27694 = n4211 & ~n8652 ;
  assign n27695 = n15931 ^ n270 ^ 1'b0 ;
  assign n27696 = n14943 & n27695 ;
  assign n27697 = n828 & ~n1225 ;
  assign n27698 = n27697 ^ n14086 ^ 1'b0 ;
  assign n27699 = n24238 ^ n18514 ^ 1'b0 ;
  assign n27700 = n10861 ^ n489 ^ 1'b0 ;
  assign n27701 = n965 | n1041 ;
  assign n27702 = n6842 | n27701 ;
  assign n27703 = ~n21778 & n27702 ;
  assign n27704 = ~n3692 & n11294 ;
  assign n27705 = n3692 & n27704 ;
  assign n27706 = n27705 ^ n9242 ^ 1'b0 ;
  assign n27707 = n10141 ^ n806 ^ 1'b0 ;
  assign n27708 = ~n5284 & n27707 ;
  assign n27711 = n9344 ^ n2942 ^ 1'b0 ;
  assign n27712 = n25674 & n27711 ;
  assign n27709 = n3139 | n10759 ;
  assign n27710 = n8648 & n27709 ;
  assign n27713 = n27712 ^ n27710 ^ 1'b0 ;
  assign n27714 = n27713 ^ n5413 ^ 1'b0 ;
  assign n27715 = n323 | n27714 ;
  assign n27716 = n5304 & ~n27715 ;
  assign n27717 = n19962 ^ n6907 ^ 1'b0 ;
  assign n27718 = ~x2 & n27717 ;
  assign n27719 = ~n2924 & n11298 ;
  assign n27720 = ~n11298 & n27719 ;
  assign n27722 = n8965 ^ n2145 ^ 1'b0 ;
  assign n27721 = n2005 & n3413 ;
  assign n27723 = n27722 ^ n27721 ^ 1'b0 ;
  assign n27724 = n18123 ^ n13921 ^ 1'b0 ;
  assign n27725 = n5718 & n27724 ;
  assign n27727 = ~n1768 & n2040 ;
  assign n27728 = n18252 | n27727 ;
  assign n27726 = n17317 & n26458 ;
  assign n27729 = n27728 ^ n27726 ^ 1'b0 ;
  assign n27730 = n16501 ^ n4317 ^ 1'b0 ;
  assign n27731 = n27729 & ~n27730 ;
  assign n27732 = ~n23889 & n27731 ;
  assign n27733 = n6892 ^ n6721 ^ 1'b0 ;
  assign n27734 = ~n38 & n27733 ;
  assign n27735 = n14077 & ~n22598 ;
  assign n27736 = n21078 ^ n2415 ^ 1'b0 ;
  assign n27737 = n21764 ^ n3687 ^ 1'b0 ;
  assign n27738 = n3467 | n27737 ;
  assign n27739 = n27736 | n27738 ;
  assign n27740 = n23184 ^ n14395 ^ 1'b0 ;
  assign n27741 = n27740 ^ n14973 ^ 1'b0 ;
  assign n27742 = n13623 ^ n5663 ^ 1'b0 ;
  assign n27743 = ~n7043 & n27742 ;
  assign n27744 = ~n16040 & n23743 ;
  assign n27745 = n27744 ^ n13017 ^ 1'b0 ;
  assign n27746 = n21023 ^ n9151 ^ 1'b0 ;
  assign n27747 = ~n2875 & n27746 ;
  assign n27748 = n13732 & ~n27747 ;
  assign n27749 = n19799 & n27748 ;
  assign n27750 = n907 & ~n3776 ;
  assign n27751 = n12223 ^ n6784 ^ 1'b0 ;
  assign n27752 = n27750 | n27751 ;
  assign n27753 = n21354 & ~n26509 ;
  assign n27755 = n16745 ^ n13806 ^ n3443 ;
  assign n27754 = n5905 | n7056 ;
  assign n27756 = n27755 ^ n27754 ^ 1'b0 ;
  assign n27757 = n5063 | n16838 ;
  assign n27758 = n22493 | n27757 ;
  assign n27759 = n23226 & ~n27758 ;
  assign n27760 = n4546 & ~n20844 ;
  assign n27761 = ~n27759 & n27760 ;
  assign n27762 = n4078 & n26220 ;
  assign n27763 = n16906 & n25563 ;
  assign n27764 = n27763 ^ n14987 ^ 1'b0 ;
  assign n27765 = n10255 ^ n5650 ^ 1'b0 ;
  assign n27766 = ~n4998 & n27765 ;
  assign n27767 = n27766 ^ n13550 ^ 1'b0 ;
  assign n27768 = ~n16207 & n17135 ;
  assign n27769 = n27768 ^ n22225 ^ 1'b0 ;
  assign n27770 = n2278 | n6365 ;
  assign n27771 = n4246 & n27770 ;
  assign n27772 = n21339 ^ n3653 ^ 1'b0 ;
  assign n27773 = n18000 ^ n12953 ^ n1638 ;
  assign n27774 = n7546 & ~n15873 ;
  assign n27775 = n8049 & n8502 ;
  assign n27776 = n27775 ^ n9592 ^ 1'b0 ;
  assign n27777 = n5206 ^ n1118 ^ 1'b0 ;
  assign n27778 = n3520 ^ n614 ^ 1'b0 ;
  assign n27779 = n27778 ^ n12002 ^ 1'b0 ;
  assign n27780 = n5860 | n27779 ;
  assign n27781 = n3718 ^ n1901 ^ 1'b0 ;
  assign n27782 = n1602 & ~n27781 ;
  assign n27783 = n3101 & n4198 ;
  assign n27784 = n1106 | n8239 ;
  assign n27785 = n26065 & ~n27784 ;
  assign n27787 = ~n1158 & n9699 ;
  assign n27786 = n5917 & n10078 ;
  assign n27788 = n27787 ^ n27786 ^ 1'b0 ;
  assign n27789 = n11260 ^ n5885 ^ 1'b0 ;
  assign n27790 = n20472 | n27789 ;
  assign n27791 = n27790 ^ n2292 ^ 1'b0 ;
  assign n27792 = n1423 & ~n14151 ;
  assign n27793 = n7875 & ~n21966 ;
  assign n27794 = n16576 ^ n279 ^ 1'b0 ;
  assign n27795 = n25159 | n27794 ;
  assign n27796 = n13759 ^ n9502 ^ 1'b0 ;
  assign n27797 = n9069 ^ n632 ^ 1'b0 ;
  assign n27798 = ~n4351 & n27797 ;
  assign n27799 = n5241 & n27798 ;
  assign n27800 = n1135 | n3845 ;
  assign n27801 = n1662 & ~n6224 ;
  assign n27802 = n5385 & n27801 ;
  assign n27803 = n12208 & ~n19854 ;
  assign n27804 = ~n12444 & n27803 ;
  assign n27805 = n27802 & ~n27804 ;
  assign n27806 = n3706 | n14186 ;
  assign n27807 = n25181 | n27806 ;
  assign n27808 = ~n7646 & n7681 ;
  assign n27809 = n27807 & n27808 ;
  assign n27810 = n7429 ^ n3337 ^ 1'b0 ;
  assign n27811 = n5397 & n20077 ;
  assign n27812 = n27811 ^ n13626 ^ 1'b0 ;
  assign n27813 = n22423 ^ n4673 ^ 1'b0 ;
  assign n27814 = n3823 | n15788 ;
  assign n27815 = n15185 ^ n246 ^ 1'b0 ;
  assign n27816 = n3853 ^ n158 ^ 1'b0 ;
  assign n27817 = n27816 ^ n11245 ^ 1'b0 ;
  assign n27818 = n19948 ^ n11827 ^ 1'b0 ;
  assign n27819 = n14120 ^ n5854 ^ 1'b0 ;
  assign n27820 = ~n10370 & n27819 ;
  assign n27821 = n1933 | n6335 ;
  assign n27822 = n27821 ^ n13656 ^ 1'b0 ;
  assign n27823 = n27822 ^ n2430 ^ 1'b0 ;
  assign n27824 = ~n7964 & n27823 ;
  assign n27825 = n5844 & ~n9707 ;
  assign n27826 = n27825 ^ n26367 ^ 1'b0 ;
  assign n27827 = n3210 ^ n1347 ^ 1'b0 ;
  assign n27828 = n27827 ^ n9299 ^ 1'b0 ;
  assign n27829 = n6687 ^ n1331 ^ 1'b0 ;
  assign n27830 = n9977 ^ n1199 ^ 1'b0 ;
  assign n27831 = n178 | n7467 ;
  assign n27832 = n4122 & n27831 ;
  assign n27833 = n357 & n27832 ;
  assign n27834 = n13706 ^ n1533 ^ 1'b0 ;
  assign n27835 = ~n15873 & n27834 ;
  assign n27836 = n8932 & n21325 ;
  assign n27837 = ~n27835 & n27836 ;
  assign n27838 = n3539 | n27837 ;
  assign n27839 = n6706 | n27838 ;
  assign n27840 = n13242 & n14701 ;
  assign n27841 = ~n14953 & n18515 ;
  assign n27842 = n3370 & n27841 ;
  assign n27844 = n470 ^ n15 ^ 1'b0 ;
  assign n27843 = n12966 | n14736 ;
  assign n27845 = n27844 ^ n27843 ^ 1'b0 ;
  assign n27846 = n26374 ^ n24010 ^ 1'b0 ;
  assign n27847 = n12966 | n17337 ;
  assign n27848 = n27847 ^ n13884 ^ 1'b0 ;
  assign n27849 = n5752 & n13928 ;
  assign n27850 = n4769 & ~n16570 ;
  assign n27851 = n11787 & n13671 ;
  assign n27852 = n4572 & n27851 ;
  assign n27853 = n13490 ^ n12237 ^ n3180 ;
  assign n27854 = ~n12207 & n16057 ;
  assign n27855 = ~n469 & n27854 ;
  assign n27856 = ~n153 & n12972 ;
  assign n27857 = n24667 ^ n15626 ^ 1'b0 ;
  assign n27858 = n15473 & n20664 ;
  assign n27859 = n27858 ^ n10288 ^ 1'b0 ;
  assign n27860 = n10156 & ~n21178 ;
  assign n27861 = n26909 ^ n23154 ^ n16029 ;
  assign n27862 = n3774 | n27861 ;
  assign n27863 = n158 | n3931 ;
  assign n27864 = n27863 ^ n832 ^ 1'b0 ;
  assign n27865 = ~n3418 & n27864 ;
  assign n27866 = n5497 & n27865 ;
  assign n27867 = ( n2825 & n3561 ) | ( n2825 & n9212 ) | ( n3561 & n9212 ) ;
  assign n27868 = ~n8081 & n12993 ;
  assign n27869 = ~n27867 & n27868 ;
  assign n27870 = n3741 & ~n27869 ;
  assign n27871 = ~n274 & n27870 ;
  assign n27872 = n8110 & n8686 ;
  assign n27873 = n2220 & n23677 ;
  assign n27874 = n27872 & n27873 ;
  assign n27875 = n13847 ^ n13665 ^ 1'b0 ;
  assign n27876 = n8620 ^ n3801 ^ 1'b0 ;
  assign n27877 = n27876 ^ n5812 ^ 1'b0 ;
  assign n27878 = n5317 & n24857 ;
  assign n27879 = n2294 & n19708 ;
  assign n27880 = ~n14854 & n27879 ;
  assign n27881 = n11931 & ~n22535 ;
  assign n27882 = n6728 & n22613 ;
  assign n27883 = ~n20325 & n27882 ;
  assign n27884 = n8408 ^ n2848 ^ 1'b0 ;
  assign n27885 = n8107 ^ n2173 ^ 1'b0 ;
  assign n27886 = n27885 ^ n4883 ^ 1'b0 ;
  assign n27887 = n5368 & ~n27886 ;
  assign n27888 = ~n2659 & n26511 ;
  assign n27889 = n7217 | n27888 ;
  assign n27890 = n27887 | n27889 ;
  assign n27891 = n1909 | n14532 ;
  assign n27892 = n872 | n15792 ;
  assign n27893 = ~n3616 & n27892 ;
  assign n27894 = n9544 ^ n1208 ^ 1'b0 ;
  assign n27895 = n4044 | n25651 ;
  assign n27896 = n14394 ^ n12920 ^ 1'b0 ;
  assign n27897 = ~n24378 & n27896 ;
  assign n27898 = ~n5719 & n7683 ;
  assign n27899 = n1036 | n4965 ;
  assign n27900 = n141 & ~n5317 ;
  assign n27901 = ( n18558 & n27899 ) | ( n18558 & n27900 ) | ( n27899 & n27900 ) ;
  assign n27902 = n27901 ^ n68 ^ 1'b0 ;
  assign n27903 = n5155 | n27902 ;
  assign n27904 = n4297 & ~n27903 ;
  assign n27905 = n1496 | n25926 ;
  assign n27906 = n27905 ^ n3346 ^ 1'b0 ;
  assign n27907 = n15633 ^ n13644 ^ 1'b0 ;
  assign n27908 = n2909 & ~n17374 ;
  assign n27909 = ~n17929 & n27908 ;
  assign n27910 = n27909 ^ n9707 ^ 1'b0 ;
  assign n27911 = n18968 ^ n977 ^ 1'b0 ;
  assign n27912 = n1401 | n6341 ;
  assign n27913 = n6341 & ~n27912 ;
  assign n27914 = n27787 ^ n24730 ^ 1'b0 ;
  assign n27915 = ~n5819 & n27914 ;
  assign n27916 = n22218 ^ n1048 ^ 1'b0 ;
  assign n27917 = n25102 ^ n2920 ^ 1'b0 ;
  assign n27918 = ~n330 & n27917 ;
  assign n27919 = n14519 & n27918 ;
  assign n27920 = n27370 ^ n7112 ^ 1'b0 ;
  assign n27923 = n2155 ^ n1851 ^ 1'b0 ;
  assign n27921 = n25588 ^ n12645 ^ 1'b0 ;
  assign n27922 = n15913 | n27921 ;
  assign n27924 = n27923 ^ n27922 ^ 1'b0 ;
  assign n27925 = ~n119 & n7140 ;
  assign n27926 = n12308 & n27925 ;
  assign n27927 = n11405 | n14609 ;
  assign n27928 = n27927 ^ n10887 ^ 1'b0 ;
  assign n27929 = n19358 & ~n27928 ;
  assign n27930 = n4526 & n27929 ;
  assign n27931 = n1793 & ~n18942 ;
  assign n27932 = n10658 & n27931 ;
  assign n27933 = n23747 ^ n632 ^ 1'b0 ;
  assign n27934 = n27933 ^ n3435 ^ 1'b0 ;
  assign n27935 = n21158 & n27934 ;
  assign n27936 = n27935 ^ n6887 ^ 1'b0 ;
  assign n27937 = n15271 ^ n6165 ^ 1'b0 ;
  assign n27938 = n898 | n4419 ;
  assign n27939 = n818 & n1841 ;
  assign n27940 = n23276 & n26667 ;
  assign n27941 = n16339 ^ n12175 ^ 1'b0 ;
  assign n27942 = n5205 & n7540 ;
  assign n27943 = n2275 ^ n627 ^ 1'b0 ;
  assign n27944 = n27943 ^ n5192 ^ 1'b0 ;
  assign n27945 = n2843 & n27944 ;
  assign n27946 = n13532 ^ n4700 ^ 1'b0 ;
  assign n27947 = n7007 | n27946 ;
  assign n27948 = n2150 & n18212 ;
  assign n27949 = n27947 & n27948 ;
  assign n27950 = ( ~n8634 & n10590 ) | ( ~n8634 & n15161 ) | ( n10590 & n15161 ) ;
  assign n27951 = n17866 ^ n1134 ^ 1'b0 ;
  assign n27952 = n820 | n27951 ;
  assign n27953 = n6074 ^ n4864 ^ 1'b0 ;
  assign n27954 = n17719 & ~n27953 ;
  assign n27955 = n6334 | n10395 ;
  assign n27956 = ~n18636 & n21322 ;
  assign n27957 = n20005 ^ n3880 ^ 1'b0 ;
  assign n27958 = n26495 & n27957 ;
  assign n27959 = ~n5034 & n12366 ;
  assign n27960 = n334 & n9134 ;
  assign n27961 = n24413 & n27960 ;
  assign n27962 = ~n27066 & n27961 ;
  assign n27963 = n3144 & n11641 ;
  assign n27964 = n18652 & n27963 ;
  assign n27965 = n549 & ~n27964 ;
  assign n27968 = n5890 | n27670 ;
  assign n27966 = n6540 ^ n1920 ^ 1'b0 ;
  assign n27967 = n19403 & ~n27966 ;
  assign n27969 = n27968 ^ n27967 ^ 1'b0 ;
  assign n27970 = n5471 & ~n27969 ;
  assign n27971 = ~n21005 & n27970 ;
  assign n27973 = n83 & ~n11944 ;
  assign n27972 = n3081 & ~n15695 ;
  assign n27974 = n27973 ^ n27972 ^ n23992 ;
  assign n27975 = n2478 | n8646 ;
  assign n27976 = n27975 ^ n26946 ^ 1'b0 ;
  assign n27977 = n13549 & n20347 ;
  assign n27978 = ~n865 & n27977 ;
  assign n27979 = n11155 ^ n6139 ^ n2572 ;
  assign n27980 = n15438 & n27979 ;
  assign n27981 = n27980 ^ n5176 ^ 1'b0 ;
  assign n27982 = n2796 & n14435 ;
  assign n27983 = ~n24573 & n27982 ;
  assign n27984 = n21643 & ~n27306 ;
  assign n27985 = n27983 | n27984 ;
  assign n27986 = n1151 & n7799 ;
  assign n27987 = n907 | n14566 ;
  assign n27988 = n2301 & ~n27987 ;
  assign n27989 = n1089 & ~n4830 ;
  assign n27990 = n8499 | n27989 ;
  assign n27991 = n12982 ^ n55 ^ 1'b0 ;
  assign n27992 = n10909 & n22639 ;
  assign n27994 = ~n1003 & n2107 ;
  assign n27995 = ~n2509 & n27994 ;
  assign n27993 = n5939 | n8686 ;
  assign n27996 = n27995 ^ n27993 ^ 1'b0 ;
  assign n27997 = ~n1559 & n27996 ;
  assign n27998 = n13470 & n13685 ;
  assign n27999 = n27998 ^ x7 ^ 1'b0 ;
  assign n28000 = ( ~n15295 & n26964 ) | ( ~n15295 & n27999 ) | ( n26964 & n27999 ) ;
  assign n28001 = n16557 ^ n6094 ^ 1'b0 ;
  assign n28002 = n14792 ^ n3343 ^ 1'b0 ;
  assign n28003 = n11399 ^ n5516 ^ 1'b0 ;
  assign n28004 = n23099 | n28003 ;
  assign n28005 = n2724 & ~n4883 ;
  assign n28006 = n28005 ^ n7978 ^ 1'b0 ;
  assign n28007 = n3277 | n28006 ;
  assign n28008 = ~n7236 & n28007 ;
  assign n28009 = n24169 ^ n22485 ^ 1'b0 ;
  assign n28010 = n6530 & n11745 ;
  assign n28011 = n10987 & n28010 ;
  assign n28012 = n8115 & ~n24249 ;
  assign n28013 = n28012 ^ n9414 ^ 1'b0 ;
  assign n28014 = n18195 ^ n12099 ^ 1'b0 ;
  assign n28015 = n3180 & n28014 ;
  assign n28016 = n25371 ^ n9069 ^ 1'b0 ;
  assign n28017 = n257 & n2700 ;
  assign n28018 = ~n2700 & n28017 ;
  assign n28019 = n1212 | n28018 ;
  assign n28020 = n28018 & ~n28019 ;
  assign n28021 = n18076 | n28020 ;
  assign n28022 = n28020 & ~n28021 ;
  assign n28023 = n28022 ^ n2100 ^ 1'b0 ;
  assign n28024 = n3452 & ~n23638 ;
  assign n28025 = ~n28023 & n28024 ;
  assign n28026 = n5607 | n17920 ;
  assign n28027 = n1763 | n28026 ;
  assign n28028 = n28027 ^ n12455 ^ 1'b0 ;
  assign n28029 = n28028 ^ n22254 ^ 1'b0 ;
  assign n28030 = ~n6287 & n18067 ;
  assign n28031 = n15034 ^ n1178 ^ 1'b0 ;
  assign n28032 = ~n28030 & n28031 ;
  assign n28033 = n25529 ^ n14683 ^ 1'b0 ;
  assign n28034 = n17948 & ~n28033 ;
  assign n28035 = n10504 ^ n8147 ^ 1'b0 ;
  assign n28036 = ~n10431 & n25227 ;
  assign n28037 = n28036 ^ n17323 ^ 1'b0 ;
  assign n28038 = ~n23531 & n28037 ;
  assign n28039 = n12674 ^ n3571 ^ 1'b0 ;
  assign n28040 = n28038 & ~n28039 ;
  assign n28041 = n10855 ^ n7430 ^ 1'b0 ;
  assign n28042 = n28041 ^ n17092 ^ 1'b0 ;
  assign n28043 = n13706 & n28042 ;
  assign n28044 = n894 & n1505 ;
  assign n28045 = ( n3774 & n4469 ) | ( n3774 & ~n9751 ) | ( n4469 & ~n9751 ) ;
  assign n28046 = n7983 | n10366 ;
  assign n28047 = n4686 & n18932 ;
  assign n28048 = n28047 ^ n2517 ^ 1'b0 ;
  assign n28049 = ~n5586 & n16421 ;
  assign n28050 = n709 & n4934 ;
  assign n28051 = n12007 & n28050 ;
  assign n28052 = n28051 ^ n16791 ^ 1'b0 ;
  assign n28053 = n2733 & n16853 ;
  assign n28054 = n2212 ^ n1600 ^ 1'b0 ;
  assign n28055 = n11630 | n28054 ;
  assign n28056 = n14874 | n28055 ;
  assign n28057 = n28056 ^ n15910 ^ 1'b0 ;
  assign n28058 = ~n22278 & n26351 ;
  assign n28059 = n25995 ^ n4689 ^ n592 ;
  assign n28060 = n10657 | n11837 ;
  assign n28061 = n19419 | n28060 ;
  assign n28062 = ~n300 & n13405 ;
  assign n28063 = n7383 & n28062 ;
  assign n28064 = n28063 ^ n17008 ^ 1'b0 ;
  assign n28065 = n14955 ^ n8914 ^ 1'b0 ;
  assign n28066 = n3566 ^ n457 ^ 1'b0 ;
  assign n28067 = n18317 | n28066 ;
  assign n28068 = n24628 ^ n15192 ^ 1'b0 ;
  assign n28069 = n19904 ^ n18150 ^ 1'b0 ;
  assign n28070 = n84 | n13425 ;
  assign n28071 = n19253 & ~n23392 ;
  assign n28072 = n28071 ^ n3857 ^ 1'b0 ;
  assign n28073 = n8833 ^ n7608 ^ 1'b0 ;
  assign n28074 = n1235 & n12348 ;
  assign n28075 = n28073 & n28074 ;
  assign n28076 = n28075 ^ n10727 ^ 1'b0 ;
  assign n28077 = n1017 & ~n28076 ;
  assign n28078 = n27463 ^ n9971 ^ 1'b0 ;
  assign n28079 = n5981 & ~n9794 ;
  assign n28080 = n28079 ^ n24060 ^ 1'b0 ;
  assign n28081 = n13186 | n28080 ;
  assign n28082 = n11239 | n13435 ;
  assign n28083 = n14845 & ~n15777 ;
  assign n28084 = ~n10536 & n28083 ;
  assign n28085 = n2017 & n4329 ;
  assign n28086 = n3264 & ~n7194 ;
  assign n28087 = n446 & n16641 ;
  assign n28088 = ~n15150 & n21884 ;
  assign n28089 = n28088 ^ n22122 ^ 1'b0 ;
  assign n28090 = n25853 | n28089 ;
  assign n28091 = n10266 | n28090 ;
  assign n28092 = n3717 & ~n28091 ;
  assign n28093 = ~n5663 & n12683 ;
  assign n28094 = ~n16469 & n21751 ;
  assign n28095 = n8067 & n28094 ;
  assign n28096 = n5032 & n8149 ;
  assign n28097 = n15319 & n28096 ;
  assign n28098 = n7923 ^ n769 ^ 1'b0 ;
  assign n28099 = n28098 ^ n9966 ^ 1'b0 ;
  assign n28100 = n6421 & ~n14385 ;
  assign n28101 = n9163 & n28100 ;
  assign n28102 = n12239 ^ n3279 ^ 1'b0 ;
  assign n28103 = ~n6080 & n8090 ;
  assign n28104 = n18116 ^ n16533 ^ 1'b0 ;
  assign n28105 = n12860 & ~n28104 ;
  assign n28106 = n8994 | n22255 ;
  assign n28107 = ~n11501 & n12242 ;
  assign n28108 = n7134 ^ n5533 ^ 1'b0 ;
  assign n28109 = n1585 & ~n28108 ;
  assign n28110 = n28109 ^ n19020 ^ 1'b0 ;
  assign n28111 = n8226 ^ n6833 ^ n2796 ;
  assign n28112 = n11046 & ~n12027 ;
  assign n28113 = n28112 ^ n23222 ^ 1'b0 ;
  assign n28114 = n7701 ^ n3597 ^ 1'b0 ;
  assign n28115 = ( n1081 & ~n5772 ) | ( n1081 & n8306 ) | ( ~n5772 & n8306 ) ;
  assign n28116 = n28115 ^ n1684 ^ 1'b0 ;
  assign n28117 = ~n2117 & n28116 ;
  assign n28118 = ~n28114 & n28117 ;
  assign n28119 = ~n8352 & n28118 ;
  assign n28120 = ~n310 & n1250 ;
  assign n28121 = ~n28119 & n28120 ;
  assign n28122 = n55 & ~n16763 ;
  assign n28123 = n28122 ^ n1052 ^ 1'b0 ;
  assign n28124 = ( n28113 & ~n28121 ) | ( n28113 & n28123 ) | ( ~n28121 & n28123 ) ;
  assign n28125 = n11126 & ~n11526 ;
  assign n28126 = n14197 & n28125 ;
  assign n28127 = n14790 ^ n1825 ^ 1'b0 ;
  assign n28128 = n28127 ^ n8710 ^ 1'b0 ;
  assign n28129 = n13051 | n16065 ;
  assign n28130 = n1645 | n28129 ;
  assign n28131 = n1033 & ~n19785 ;
  assign n28132 = n28131 ^ n1478 ^ 1'b0 ;
  assign n28133 = n6713 & ~n28132 ;
  assign n28134 = ~n28130 & n28133 ;
  assign n28136 = n11433 ^ n715 ^ 1'b0 ;
  assign n28137 = ~n3056 & n28136 ;
  assign n28135 = ~n5590 & n24664 ;
  assign n28138 = n28137 ^ n28135 ^ 1'b0 ;
  assign n28139 = n14908 | n19891 ;
  assign n28140 = n17010 & n28139 ;
  assign n28141 = n28140 ^ n3827 ^ 1'b0 ;
  assign n28142 = n4070 | n8086 ;
  assign n28143 = n2736 | n28142 ;
  assign n28144 = n556 & ~n28143 ;
  assign n28145 = n1768 & ~n7338 ;
  assign n28146 = ( n14662 & n22197 ) | ( n14662 & n24699 ) | ( n22197 & n24699 ) ;
  assign n28147 = ~n13077 & n28146 ;
  assign n28148 = n28147 ^ n5501 ^ 1'b0 ;
  assign n28149 = ~n2751 & n15657 ;
  assign n28150 = n1770 & n3360 ;
  assign n28151 = n28150 ^ n24675 ^ 1'b0 ;
  assign n28152 = ~n2680 & n9831 ;
  assign n28154 = ~n1023 & n10661 ;
  assign n28153 = ~n671 & n872 ;
  assign n28155 = n28154 ^ n28153 ^ 1'b0 ;
  assign n28156 = n4508 ^ n1110 ^ 1'b0 ;
  assign n28157 = ( n19479 & n27406 ) | ( n19479 & n28156 ) | ( n27406 & n28156 ) ;
  assign n28158 = n8408 & ~n16082 ;
  assign n28159 = n25519 & n28158 ;
  assign n28160 = n3398 & n9697 ;
  assign n28161 = n116 & ~n24415 ;
  assign n28162 = n28161 ^ n17457 ^ 1'b0 ;
  assign n28163 = n28160 | n28162 ;
  assign n28164 = n4127 ^ n1227 ^ 1'b0 ;
  assign n28165 = n119 | n28164 ;
  assign n28166 = n28165 ^ n1705 ^ 1'b0 ;
  assign n28167 = ~n3064 & n3684 ;
  assign n28168 = ~n9585 & n28167 ;
  assign n28169 = ~n8749 & n18923 ;
  assign n28170 = n4902 | n12186 ;
  assign n28171 = n15336 & n28170 ;
  assign n28172 = n1537 & n4485 ;
  assign n28173 = ~n3694 & n15465 ;
  assign n28174 = n8586 & n9595 ;
  assign n28175 = ~n6323 & n28174 ;
  assign n28176 = ~n12360 & n28175 ;
  assign n28177 = n764 | n23973 ;
  assign n28178 = n2973 ^ n175 ^ 1'b0 ;
  assign n28179 = n24645 ^ n21735 ^ 1'b0 ;
  assign n28180 = n2017 & ~n22228 ;
  assign n28181 = n28180 ^ n14534 ^ 1'b0 ;
  assign n28182 = ~n21449 & n28181 ;
  assign n28183 = n2652 & ~n4981 ;
  assign n28184 = ~n10247 & n11379 ;
  assign n28185 = n13419 ^ n10195 ^ 1'b0 ;
  assign n28186 = n17163 & ~n28185 ;
  assign n28187 = n13077 ^ n7105 ^ 1'b0 ;
  assign n28188 = n5860 | n28187 ;
  assign n28189 = n17670 & n22036 ;
  assign n28190 = n3339 & n28189 ;
  assign n28191 = n3378 | n25118 ;
  assign n28192 = n1194 | n28191 ;
  assign n28193 = n2565 ^ n2245 ^ 1'b0 ;
  assign n28194 = n1105 | n28193 ;
  assign n28195 = n14569 | n28194 ;
  assign n28196 = n7641 & ~n8856 ;
  assign n28197 = n28195 & n28196 ;
  assign n28198 = n164 & n2870 ;
  assign n28199 = ~n149 & n2439 ;
  assign n28200 = ~n2439 & n28199 ;
  assign n28201 = n11691 & ~n28200 ;
  assign n28202 = ~n547 & n28201 ;
  assign n28203 = n547 & n28202 ;
  assign n28204 = n24598 ^ n11201 ^ 1'b0 ;
  assign n28205 = n10447 & ~n28204 ;
  assign n28206 = n5046 ^ n21 ^ 1'b0 ;
  assign n28207 = n272 & n18477 ;
  assign n28208 = n28206 & n28207 ;
  assign n28210 = n3144 & n6969 ;
  assign n28209 = n2384 & ~n8446 ;
  assign n28211 = n28210 ^ n28209 ^ 1'b0 ;
  assign n28213 = n3580 & n8948 ;
  assign n28214 = n12498 | n28213 ;
  assign n28215 = n2331 | n28214 ;
  assign n28212 = n6414 | n9137 ;
  assign n28216 = n28215 ^ n28212 ^ 1'b0 ;
  assign n28217 = n6863 | n28216 ;
  assign n28218 = n26146 ^ n6588 ^ 1'b0 ;
  assign n28219 = n6636 | n28218 ;
  assign n28220 = n2027 & ~n28219 ;
  assign n28221 = n14353 ^ n6772 ^ 1'b0 ;
  assign n28222 = ( ~n68 & n3744 ) | ( ~n68 & n4817 ) | ( n3744 & n4817 ) ;
  assign n28223 = n12200 ^ n371 ^ 1'b0 ;
  assign n28224 = n8991 & ~n28223 ;
  assign n28225 = n17297 ^ n15748 ^ 1'b0 ;
  assign n28226 = n446 | n20123 ;
  assign n28227 = n1175 | n21545 ;
  assign n28228 = n1065 & n10280 ;
  assign n28229 = n6126 | n11608 ;
  assign n28230 = n28229 ^ n2185 ^ 1'b0 ;
  assign n28231 = n2995 & n3931 ;
  assign n28232 = ~n9159 & n16288 ;
  assign n28233 = n28232 ^ n4256 ^ 1'b0 ;
  assign n28234 = n28233 ^ n10213 ^ 1'b0 ;
  assign n28235 = n13422 ^ n9682 ^ 1'b0 ;
  assign n28236 = n591 | n28235 ;
  assign n28237 = n23721 | n28236 ;
  assign n28238 = n11125 ^ n5580 ^ 1'b0 ;
  assign n28239 = n3871 & n28238 ;
  assign n28240 = n10673 & ~n28239 ;
  assign n28241 = n1860 | n10005 ;
  assign n28242 = n23972 ^ n19540 ^ n19104 ;
  assign n28243 = n6919 & ~n13068 ;
  assign n28245 = ~n4606 & n5890 ;
  assign n28246 = n28245 ^ n10535 ^ 1'b0 ;
  assign n28244 = n7217 & ~n21843 ;
  assign n28247 = n28246 ^ n28244 ^ 1'b0 ;
  assign n28248 = n21321 ^ n1047 ^ 1'b0 ;
  assign n28249 = n4522 & n28248 ;
  assign n28250 = n3614 & n28249 ;
  assign n28251 = ~n236 & n13660 ;
  assign n28252 = n18007 ^ n7679 ^ 1'b0 ;
  assign n28253 = ~n28251 & n28252 ;
  assign n28254 = ~n440 & n23689 ;
  assign n28255 = ~n616 & n28254 ;
  assign n28256 = n2187 & ~n19804 ;
  assign n28257 = n22746 ^ n709 ^ 1'b0 ;
  assign n28258 = n25342 ^ n21377 ^ n9871 ;
  assign n28259 = ~n1690 & n14054 ;
  assign n28260 = ~n1430 & n10561 ;
  assign n28261 = n28260 ^ n17861 ^ 1'b0 ;
  assign n28262 = n28259 & n28261 ;
  assign n28263 = n1366 | n27483 ;
  assign n28264 = n23057 | n28263 ;
  assign n28265 = n6610 ^ n3924 ^ 1'b0 ;
  assign n28266 = n6729 ^ n4361 ^ 1'b0 ;
  assign n28267 = n28265 & ~n28266 ;
  assign n28268 = n9592 ^ n7754 ^ n4706 ;
  assign n28269 = n28268 ^ n7187 ^ 1'b0 ;
  assign n28270 = ~n1283 & n18731 ;
  assign n28271 = n5501 ^ n1048 ^ 1'b0 ;
  assign n28272 = n15157 ^ n7523 ^ 1'b0 ;
  assign n28273 = n15687 & ~n22649 ;
  assign n28274 = n5002 & ~n28273 ;
  assign n28275 = n4077 ^ n1132 ^ 1'b0 ;
  assign n28276 = n24628 ^ n22850 ^ 1'b0 ;
  assign n28277 = ~n8321 & n9542 ;
  assign n28278 = n28276 & n28277 ;
  assign n28279 = ~n15698 & n21077 ;
  assign n28280 = n28279 ^ n949 ^ 1'b0 ;
  assign n28281 = n9631 ^ n3344 ^ 1'b0 ;
  assign n28282 = ~n912 & n28281 ;
  assign n28283 = n3660 & n28282 ;
  assign n28284 = n4687 & ~n28283 ;
  assign n28285 = n25419 ^ n25085 ^ 1'b0 ;
  assign n28287 = ~n5454 & n10255 ;
  assign n28286 = n5452 & n8613 ;
  assign n28288 = n28287 ^ n28286 ^ 1'b0 ;
  assign n28289 = ( ~n832 & n7412 ) | ( ~n832 & n15699 ) | ( n7412 & n15699 ) ;
  assign n28290 = n11672 & ~n17094 ;
  assign n28291 = n22265 & n28290 ;
  assign n28292 = n11590 ^ n8692 ^ 1'b0 ;
  assign n28293 = n1961 & n28292 ;
  assign n28294 = ~n1449 & n2321 ;
  assign n28295 = n23848 & n28294 ;
  assign n28296 = n23948 & n28295 ;
  assign n28297 = n1168 | n28296 ;
  assign n28298 = ~n556 & n4372 ;
  assign n28299 = ~n15902 & n28298 ;
  assign n28300 = n10728 & ~n28299 ;
  assign n28301 = n28300 ^ n15766 ^ 1'b0 ;
  assign n28302 = ~n4976 & n28301 ;
  assign n28303 = n7497 | n14771 ;
  assign n28304 = n1790 & ~n28303 ;
  assign n28305 = ~n149 & n9032 ;
  assign n28306 = ~n4203 & n28305 ;
  assign n28308 = n280 & ~n23252 ;
  assign n28309 = n556 & ~n28308 ;
  assign n28307 = n11603 & ~n14780 ;
  assign n28310 = n28309 ^ n28307 ^ 1'b0 ;
  assign n28311 = n25302 ^ n13338 ^ 1'b0 ;
  assign n28312 = n5451 ^ n3021 ^ 1'b0 ;
  assign n28313 = n3537 & ~n4505 ;
  assign n28314 = ~n7588 & n28313 ;
  assign n28315 = n7433 ^ n3613 ^ 1'b0 ;
  assign n28316 = n1444 & ~n13960 ;
  assign n28317 = n4891 & n28316 ;
  assign n28318 = n28315 & ~n28317 ;
  assign n28319 = n16007 ^ n12291 ^ 1'b0 ;
  assign n28320 = n11024 | n28319 ;
  assign n28321 = ~n5857 & n19564 ;
  assign n28323 = n3141 & ~n3598 ;
  assign n28324 = n9715 & n28323 ;
  assign n28322 = n9979 & ~n14690 ;
  assign n28325 = n28324 ^ n28322 ^ n5697 ;
  assign n28326 = n207 & n6234 ;
  assign n28327 = ~n24297 & n28326 ;
  assign n28328 = n28327 ^ n18953 ^ 1'b0 ;
  assign n28329 = n14409 & n28328 ;
  assign n28330 = ~n129 & n4440 ;
  assign n28331 = n12266 & ~n28330 ;
  assign n28332 = ( n6752 & ~n23771 ) | ( n6752 & n28331 ) | ( ~n23771 & n28331 ) ;
  assign n28333 = n11419 ^ n5327 ^ 1'b0 ;
  assign n28334 = n19725 | n28333 ;
  assign n28335 = n25349 | n28334 ;
  assign n28336 = n3177 & ~n13781 ;
  assign n28337 = ~n22168 & n28336 ;
  assign n28338 = n28215 ^ n9132 ^ 1'b0 ;
  assign n28339 = n11659 & ~n28338 ;
  assign n28340 = n12308 & ~n22223 ;
  assign n28341 = ~n8811 & n28340 ;
  assign n28342 = n5846 & ~n18217 ;
  assign n28343 = n28342 ^ n4817 ^ 1'b0 ;
  assign n28344 = n8980 ^ n6751 ^ 1'b0 ;
  assign n28345 = ~n28343 & n28344 ;
  assign n28346 = ~n28341 & n28345 ;
  assign n28347 = ~n9607 & n28346 ;
  assign n28356 = n2733 | n6134 ;
  assign n28357 = n28356 ^ n2221 ^ 1'b0 ;
  assign n28348 = n2482 & n26304 ;
  assign n28349 = ~n6037 & n12272 ;
  assign n28350 = n28349 ^ n3793 ^ 1'b0 ;
  assign n28351 = n28348 | n28350 ;
  assign n28352 = n28351 ^ n12512 ^ 1'b0 ;
  assign n28353 = n9928 ^ n5860 ^ 1'b0 ;
  assign n28354 = n28352 | n28353 ;
  assign n28355 = n16041 | n28354 ;
  assign n28358 = n28357 ^ n28355 ^ 1'b0 ;
  assign n28359 = n1802 ^ n246 ^ 1'b0 ;
  assign n28360 = n10833 ^ n1922 ^ 1'b0 ;
  assign n28361 = n18505 & ~n28360 ;
  assign n28362 = ~n7868 & n22247 ;
  assign n28363 = ~n810 & n3966 ;
  assign n28364 = n14324 | n28363 ;
  assign n28365 = n13525 ^ n274 ^ 1'b0 ;
  assign n28366 = n3519 | n8644 ;
  assign n28367 = n28365 | n28366 ;
  assign n28368 = n21244 | n27718 ;
  assign n28369 = n18190 ^ n185 ^ 1'b0 ;
  assign n28370 = n14967 ^ n7887 ^ n294 ;
  assign n28371 = n9870 & ~n28370 ;
  assign n28372 = ~n13364 & n28371 ;
  assign n28373 = n28372 ^ n18096 ^ 1'b0 ;
  assign n28374 = n15775 ^ n5890 ^ 1'b0 ;
  assign n28375 = n3064 & n15287 ;
  assign n28376 = n17360 | n28375 ;
  assign n28377 = n9192 & n28376 ;
  assign n28378 = n11224 ^ n1705 ^ 1'b0 ;
  assign n28379 = n2603 & ~n12887 ;
  assign n28380 = n467 & ~n28379 ;
  assign n28381 = n21764 ^ n10733 ^ 1'b0 ;
  assign n28382 = n14262 & ~n28381 ;
  assign n28383 = x9 & ~n8984 ;
  assign n28384 = n10115 & n21033 ;
  assign n28385 = n3559 & n28384 ;
  assign n28386 = n9449 & n27412 ;
  assign n28387 = n17012 & n28386 ;
  assign n28388 = n14203 ^ n233 ^ 1'b0 ;
  assign n28389 = n1592 & ~n12300 ;
  assign n28390 = ~n1469 & n28389 ;
  assign n28391 = n13551 ^ n6664 ^ 1'b0 ;
  assign n28392 = n28390 & n28391 ;
  assign n28393 = n428 | n28392 ;
  assign n28394 = n5850 | n7071 ;
  assign n28395 = n28394 ^ n17581 ^ 1'b0 ;
  assign n28396 = n1990 & n20004 ;
  assign n28397 = ( n9871 & ~n13556 ) | ( n9871 & n19299 ) | ( ~n13556 & n19299 ) ;
  assign n28398 = n726 & ~n6090 ;
  assign n28399 = n604 | n11116 ;
  assign n28400 = n8527 ^ n4312 ^ 1'b0 ;
  assign n28401 = n28400 ^ n12123 ^ 1'b0 ;
  assign n28402 = ~n3663 & n28401 ;
  assign n28403 = n10046 & ~n28402 ;
  assign n28404 = n28399 & n28403 ;
  assign n28405 = n8515 & n16193 ;
  assign n28406 = ~n10684 & n10995 ;
  assign n28407 = n28406 ^ n6090 ^ 1'b0 ;
  assign n28408 = n21625 ^ n4258 ^ 1'b0 ;
  assign n28409 = ~n12777 & n28408 ;
  assign n28410 = ( n479 & n5858 ) | ( n479 & n6656 ) | ( n5858 & n6656 ) ;
  assign n28411 = n28410 ^ n12169 ^ 1'b0 ;
  assign n28412 = n22193 & n28411 ;
  assign n28413 = ~n1637 & n28412 ;
  assign n28414 = n13977 ^ n233 ^ 1'b0 ;
  assign n28415 = n11323 & n28414 ;
  assign n28416 = n12466 ^ n390 ^ 1'b0 ;
  assign n28417 = ~n10059 & n15098 ;
  assign n28418 = n28417 ^ n3356 ^ 1'b0 ;
  assign n28419 = ~n3931 & n28418 ;
  assign n28420 = n1394 | n2843 ;
  assign n28421 = n19351 ^ n1318 ^ 1'b0 ;
  assign n28422 = n12188 ^ n11820 ^ 1'b0 ;
  assign n28423 = n3270 & ~n9286 ;
  assign n28424 = n9739 & ~n16308 ;
  assign n28425 = n18401 ^ n227 ^ 1'b0 ;
  assign n28426 = n9596 & ~n28425 ;
  assign n28427 = n28426 ^ n3237 ^ 1'b0 ;
  assign n28428 = n3143 & ~n28427 ;
  assign n28429 = n3154 | n23780 ;
  assign n28430 = n2025 & ~n4817 ;
  assign n28431 = n11272 & ~n24081 ;
  assign n28432 = n28430 & n28431 ;
  assign n28433 = ( n1060 & n22485 ) | ( n1060 & n28432 ) | ( n22485 & n28432 ) ;
  assign n28435 = n10394 ^ n37 ^ 1'b0 ;
  assign n28436 = n9195 & n28435 ;
  assign n28437 = n4250 & ~n20415 ;
  assign n28438 = ~n28436 & n28437 ;
  assign n28434 = n9721 | n20807 ;
  assign n28439 = n28438 ^ n28434 ^ 1'b0 ;
  assign n28440 = n2263 & ~n28439 ;
  assign n28441 = n28440 ^ n25741 ^ 1'b0 ;
  assign n28442 = ~n7338 & n18268 ;
  assign n28443 = n2179 | n28442 ;
  assign n28444 = n11209 | n27683 ;
  assign n28445 = n6094 & n16478 ;
  assign n28477 = n1463 & ~n4538 ;
  assign n28478 = n4538 & n28477 ;
  assign n28479 = n6361 | n28478 ;
  assign n28480 = n2041 & n4283 ;
  assign n28481 = ~n4283 & n28480 ;
  assign n28482 = n10790 & n28481 ;
  assign n28483 = n28479 | n28482 ;
  assign n28484 = n28479 & ~n28483 ;
  assign n28473 = n756 & n1626 ;
  assign n28474 = ~n1626 & n28473 ;
  assign n28475 = ~n6916 & n28474 ;
  assign n28476 = ~n17721 & n28475 ;
  assign n28485 = n28484 ^ n28476 ^ 1'b0 ;
  assign n28446 = n10018 ^ n6944 ^ 1'b0 ;
  assign n28447 = n6439 & n23960 ;
  assign n28448 = ~n277 & n28447 ;
  assign n28449 = n28448 ^ n5252 ^ 1'b0 ;
  assign n28450 = n1475 & n1997 ;
  assign n28451 = ~n1997 & n28450 ;
  assign n28452 = n1482 & ~n6876 ;
  assign n28453 = n28451 & n28452 ;
  assign n28454 = ~n2603 & n28453 ;
  assign n28455 = ~n139 & n220 ;
  assign n28456 = ~n220 & n28455 ;
  assign n28457 = n273 & n28456 ;
  assign n28458 = n232 & n28457 ;
  assign n28459 = n590 & n28458 ;
  assign n28460 = ~n75 & n28459 ;
  assign n28461 = n28460 ^ n7839 ^ 1'b0 ;
  assign n28462 = ~n133 & n21896 ;
  assign n28463 = ~n20858 & n28462 ;
  assign n28464 = n265 & ~n18498 ;
  assign n28465 = n18498 & n28464 ;
  assign n28466 = n28465 ^ n1135 ^ 1'b0 ;
  assign n28467 = n28463 & n28466 ;
  assign n28468 = ~n28461 & n28467 ;
  assign n28469 = n28454 & n28468 ;
  assign n28470 = n28449 | n28469 ;
  assign n28471 = n28446 & ~n28470 ;
  assign n28472 = n1588 | n28471 ;
  assign n28486 = n28485 ^ n28472 ^ 1'b0 ;
  assign n28487 = n19674 | n27444 ;
  assign n28488 = n25607 | n28487 ;
  assign n28489 = n6249 | n28488 ;
  assign n28490 = n8385 | n8705 ;
  assign n28491 = ~n15192 & n28490 ;
  assign n28492 = ~n4591 & n28491 ;
  assign n28493 = n23334 ^ n17946 ^ 1'b0 ;
  assign n28494 = n4687 & ~n7358 ;
  assign n28495 = n28494 ^ n9899 ^ 1'b0 ;
  assign n28496 = n13613 | n22107 ;
  assign n28497 = ~n79 & n3504 ;
  assign n28498 = ( n622 & ~n5065 ) | ( n622 & n28497 ) | ( ~n5065 & n28497 ) ;
  assign n28499 = n17861 ^ n5968 ^ 1'b0 ;
  assign n28500 = n6039 & n20540 ;
  assign n28501 = n28500 ^ n6911 ^ 1'b0 ;
  assign n28502 = n3699 & n4622 ;
  assign n28503 = n28502 ^ n2819 ^ 1'b0 ;
  assign n28504 = ~n8278 & n28503 ;
  assign n28505 = n8018 & n28504 ;
  assign n28506 = ~n8018 & n28505 ;
  assign n28507 = ( n4611 & n16612 ) | ( n4611 & n28506 ) | ( n16612 & n28506 ) ;
  assign n28508 = n24973 ^ n1323 ^ 1'b0 ;
  assign n28509 = n15151 & ~n28508 ;
  assign n28510 = n1783 & ~n17854 ;
  assign n28511 = n28510 ^ n14646 ^ 1'b0 ;
  assign n28512 = ~n2618 & n28511 ;
  assign n28513 = n28512 ^ n104 ^ 1'b0 ;
  assign n28516 = n323 & n928 ;
  assign n28517 = ~n928 & n28516 ;
  assign n28514 = ~n1499 & n8088 ;
  assign n28515 = n1499 & n28514 ;
  assign n28518 = n28517 ^ n28515 ^ 1'b0 ;
  assign n28519 = ~n1225 & n28518 ;
  assign n28520 = n3888 & n28519 ;
  assign n28521 = n12679 & n28520 ;
  assign n28522 = n22744 ^ n13379 ^ 1'b0 ;
  assign n28523 = n16336 ^ n9141 ^ 1'b0 ;
  assign n28524 = n10464 | n28523 ;
  assign n28525 = n2107 & n5718 ;
  assign n28526 = ~n9391 & n27335 ;
  assign n28527 = n28526 ^ n13308 ^ 1'b0 ;
  assign n28528 = n28525 & ~n28527 ;
  assign n28529 = n4740 & ~n28528 ;
  assign n28530 = n24393 ^ n532 ^ 1'b0 ;
  assign n28531 = ~n15246 & n28530 ;
  assign n28532 = ~n654 & n5165 ;
  assign n28533 = ~n6818 & n28532 ;
  assign n28534 = n25904 ^ n1310 ^ 1'b0 ;
  assign n28535 = n28533 & n28534 ;
  assign n28536 = n1555 | n25130 ;
  assign n28537 = n5202 | n17674 ;
  assign n28538 = n13759 & n16545 ;
  assign n28539 = n28538 ^ n22856 ^ 1'b0 ;
  assign n28540 = n28537 | n28539 ;
  assign n28541 = n23508 ^ n9209 ^ 1'b0 ;
  assign n28542 = n9667 & n27431 ;
  assign n28543 = n4196 & ~n10403 ;
  assign n28544 = n28543 ^ n1959 ^ 1'b0 ;
  assign n28545 = n3340 & ~n28544 ;
  assign n28546 = n814 & ~n28545 ;
  assign n28547 = n880 & n2130 ;
  assign n28548 = ~n21394 & n28547 ;
  assign n28549 = n11338 & ~n15790 ;
  assign n28550 = n3412 | n4817 ;
  assign n28551 = n28550 ^ n22234 ^ 1'b0 ;
  assign n28552 = n24179 & ~n28551 ;
  assign n28553 = n23154 ^ n2705 ^ 1'b0 ;
  assign n28554 = n27753 & ~n28553 ;
  assign n28555 = n28554 ^ n2578 ^ 1'b0 ;
  assign n28556 = n11776 ^ n776 ^ 1'b0 ;
  assign n28557 = n2165 & n4358 ;
  assign n28558 = n17119 & n28557 ;
  assign n28559 = ~n28556 & n28558 ;
  assign n28560 = ~n4990 & n9751 ;
  assign n28561 = n28560 ^ n20118 ^ 1'b0 ;
  assign n28562 = n14920 ^ n2404 ^ 1'b0 ;
  assign n28563 = n23472 ^ n2680 ^ 1'b0 ;
  assign n28564 = n8416 & n9371 ;
  assign n28565 = ~n16748 & n20474 ;
  assign n28566 = n1527 & n20931 ;
  assign n28567 = x6 & n186 ;
  assign n28568 = ~x6 & n28567 ;
  assign n28569 = n28568 ^ n1475 ^ 1'b0 ;
  assign n28570 = n28566 & ~n28569 ;
  assign n28574 = n732 & n3921 ;
  assign n28575 = ~n732 & n28574 ;
  assign n28576 = n6837 | n28575 ;
  assign n28577 = n28575 & ~n28576 ;
  assign n28571 = n1419 | n7898 ;
  assign n28572 = n7898 & ~n28571 ;
  assign n28573 = n28572 ^ n7714 ^ 1'b0 ;
  assign n28578 = n28577 ^ n28573 ^ 1'b0 ;
  assign n28579 = n6793 & ~n28578 ;
  assign n28580 = n2034 & n28579 ;
  assign n28581 = ~n28570 & n28580 ;
  assign n28582 = n23896 & ~n28581 ;
  assign n28583 = n28582 ^ n21296 ^ 1'b0 ;
  assign n28584 = ~n372 & n15121 ;
  assign n28585 = n4075 & ~n28584 ;
  assign n28586 = ~n5119 & n28585 ;
  assign n28587 = n12560 & n15472 ;
  assign n28595 = ~n159 & n1506 ;
  assign n28596 = n159 & n28595 ;
  assign n28588 = n1588 | n4970 ;
  assign n28589 = n4970 & ~n28588 ;
  assign n28590 = n28589 ^ n1961 ^ 1'b0 ;
  assign n28591 = ~n1008 & n3583 ;
  assign n28592 = n1008 & n28591 ;
  assign n28593 = n6148 & ~n28592 ;
  assign n28594 = n28590 & n28593 ;
  assign n28597 = n28596 ^ n28594 ^ 1'b0 ;
  assign n28598 = n28597 ^ n3423 ^ 1'b0 ;
  assign n28599 = n9739 ^ n9540 ^ 1'b0 ;
  assign n28600 = n24097 & n28599 ;
  assign n28601 = n7920 & n9593 ;
  assign n28602 = n28600 & n28601 ;
  assign n28603 = n4604 ^ n3371 ^ 1'b0 ;
  assign n28604 = n17649 | n28603 ;
  assign n28605 = n2967 & n28604 ;
  assign n28606 = n2509 & ~n8162 ;
  assign n28607 = n20525 & n28606 ;
  assign n28608 = n11443 & ~n28607 ;
  assign n28609 = n28608 ^ n2943 ^ 1'b0 ;
  assign n28610 = n8207 & n16038 ;
  assign n28611 = n14953 & n28610 ;
  assign n28612 = n8918 ^ n2140 ^ 1'b0 ;
  assign n28613 = ~n6474 & n28612 ;
  assign n28614 = n28613 ^ n2732 ^ 1'b0 ;
  assign n28615 = ~n18156 & n23759 ;
  assign n28616 = n9922 & n28615 ;
  assign n28617 = ~n5994 & n24154 ;
  assign n28618 = ~n22853 & n25527 ;
  assign n28619 = n28618 ^ n3462 ^ 1'b0 ;
  assign n28620 = n5802 & ~n12291 ;
  assign n28621 = ~n20276 & n28620 ;
  assign n28622 = n4123 | n14841 ;
  assign n28623 = n28622 ^ n9601 ^ 1'b0 ;
  assign n28624 = n23314 & ~n28623 ;
  assign n28625 = n6596 ^ n4155 ^ 1'b0 ;
  assign n28626 = n16803 ^ n13983 ^ 1'b0 ;
  assign n28627 = n2606 & n8276 ;
  assign n28628 = ~n16443 & n28627 ;
  assign n28629 = n2668 & ~n3803 ;
  assign n28630 = n10785 & n28629 ;
  assign n28631 = ~n12749 & n24094 ;
  assign n28632 = n28631 ^ n12269 ^ 1'b0 ;
  assign n28633 = n28632 ^ n19316 ^ n7217 ;
  assign n28634 = ~n2842 & n14690 ;
  assign n28635 = n6536 ^ n1096 ^ 1'b0 ;
  assign n28636 = n2647 & n16243 ;
  assign n28637 = n28636 ^ n4684 ^ 1'b0 ;
  assign n28638 = n1390 & ~n6515 ;
  assign n28639 = n15576 | n24713 ;
  assign n28640 = n28638 & ~n28639 ;
  assign n28641 = n962 & n23739 ;
  assign n28642 = ( n236 & ~n3820 ) | ( n236 & n18546 ) | ( ~n3820 & n18546 ) ;
  assign n28643 = n922 & n19789 ;
  assign n28644 = n28643 ^ n12643 ^ 1'b0 ;
  assign n28645 = n24907 & n28644 ;
  assign n28646 = n8128 ^ n1385 ^ 1'b0 ;
  assign n28647 = n6154 & n10352 ;
  assign n28648 = n7311 | n14376 ;
  assign n28649 = n10658 ^ n1165 ^ 1'b0 ;
  assign n28650 = ~n1631 & n6923 ;
  assign n28651 = n12495 | n28650 ;
  assign n28652 = n4419 & n6713 ;
  assign n28653 = n28652 ^ n8624 ^ 1'b0 ;
  assign n28654 = n28653 ^ n5621 ^ 1'b0 ;
  assign n28655 = n7144 & n24959 ;
  assign n28656 = n28655 ^ n14872 ^ 1'b0 ;
  assign n28657 = n6700 ^ n1433 ^ 1'b0 ;
  assign n28658 = n28657 ^ n20399 ^ 1'b0 ;
  assign n28659 = n1414 & ~n18324 ;
  assign n28660 = ( n2947 & n2974 ) | ( n2947 & n28659 ) | ( n2974 & n28659 ) ;
  assign n28661 = n15596 ^ n3559 ^ 1'b0 ;
  assign n28662 = n4358 & n12887 ;
  assign n28663 = n6225 & n7751 ;
  assign n28664 = n13431 & n28663 ;
  assign n28665 = n14739 ^ n6263 ^ 1'b0 ;
  assign n28666 = n28664 | n28665 ;
  assign n28667 = n8256 & ~n28666 ;
  assign n28668 = ~n28662 & n28667 ;
  assign n28669 = n10959 ^ n10031 ^ 1'b0 ;
  assign n28670 = n321 & n9910 ;
  assign n28671 = n1834 & n5232 ;
  assign n28672 = n1179 & n13356 ;
  assign n28674 = n1105 & ~n11731 ;
  assign n28673 = ~n567 & n22424 ;
  assign n28675 = n28674 ^ n28673 ^ 1'b0 ;
  assign n28676 = n12117 & ~n28675 ;
  assign n28677 = ~n1958 & n13164 ;
  assign n28678 = n28676 & n28677 ;
  assign n28679 = n22494 ^ n4972 ^ 1'b0 ;
  assign n28680 = n6911 | n28679 ;
  assign n28681 = n13874 ^ n1235 ^ 1'b0 ;
  assign n28682 = n1677 & n28681 ;
  assign n28683 = n2316 ^ n1793 ^ n1041 ;
  assign n28684 = ~n1831 & n28683 ;
  assign n28685 = ~n19150 & n22669 ;
  assign n28686 = n23950 ^ n18035 ^ 1'b0 ;
  assign n28687 = n16817 | n28686 ;
  assign n28688 = n18302 ^ n14657 ^ 1'b0 ;
  assign n28689 = n23732 & n28688 ;
  assign n28692 = ~n9267 & n13985 ;
  assign n28693 = ~n19516 & n28692 ;
  assign n28690 = n19868 ^ n12655 ^ 1'b0 ;
  assign n28691 = n27840 & ~n28690 ;
  assign n28694 = n28693 ^ n28691 ^ 1'b0 ;
  assign n28695 = n14466 ^ n599 ^ 1'b0 ;
  assign n28697 = ~n11091 & n12856 ;
  assign n28696 = n24900 & ~n26202 ;
  assign n28698 = n28697 ^ n28696 ^ 1'b0 ;
  assign n28699 = n993 & ~n2052 ;
  assign n28700 = n2052 & n28699 ;
  assign n28701 = n562 & n28700 ;
  assign n28702 = n194 & n618 ;
  assign n28703 = ~n194 & n28702 ;
  assign n28704 = n6581 & ~n28703 ;
  assign n28705 = n28701 & n28704 ;
  assign n28706 = ~n1322 & n24606 ;
  assign n28707 = n28705 & n28706 ;
  assign n28712 = n942 ^ n622 ^ 1'b0 ;
  assign n28713 = ~n8764 & n28712 ;
  assign n28714 = ~n28712 & n28713 ;
  assign n28708 = n1233 & ~n9459 ;
  assign n28709 = n3461 ^ n715 ^ 1'b0 ;
  assign n28710 = ~n7554 & n28709 ;
  assign n28711 = ~n28708 & n28710 ;
  assign n28715 = n28714 ^ n28711 ^ 1'b0 ;
  assign n28716 = ~n28707 & n28715 ;
  assign n28717 = n28716 ^ n21856 ^ 1'b0 ;
  assign n28718 = n20700 & n24654 ;
  assign n28719 = ~n1166 & n10298 ;
  assign n28720 = n25785 ^ n19347 ^ 1'b0 ;
  assign n28721 = n1613 & ~n22474 ;
  assign n28722 = n26486 ^ n18197 ^ 1'b0 ;
  assign n28723 = ~n13449 & n21035 ;
  assign n28724 = n28723 ^ n11827 ^ 1'b0 ;
  assign n28725 = n4307 & ~n28724 ;
  assign n28726 = ~n2991 & n23113 ;
  assign n28727 = ~n16136 & n28726 ;
  assign n28728 = n17203 ^ n4088 ^ 1'b0 ;
  assign n28729 = n7511 ^ n5885 ^ 1'b0 ;
  assign n28730 = n743 & ~n2163 ;
  assign n28731 = n28729 | n28730 ;
  assign n28733 = n5860 & n12293 ;
  assign n28734 = n19619 & n28733 ;
  assign n28732 = ( ~n3008 & n8988 ) | ( ~n3008 & n16161 ) | ( n8988 & n16161 ) ;
  assign n28735 = n28734 ^ n28732 ^ n9272 ;
  assign n28736 = ~n12507 & n24720 ;
  assign n28737 = n28736 ^ n10234 ^ 1'b0 ;
  assign n28738 = n22426 ^ n17678 ^ 1'b0 ;
  assign n28739 = ~n6192 & n28738 ;
  assign n28740 = n4264 & ~n14876 ;
  assign n28741 = ~n292 & n6331 ;
  assign n28742 = n20513 ^ n14443 ^ 1'b0 ;
  assign n28745 = n7481 | n13108 ;
  assign n28743 = n190 | n2556 ;
  assign n28744 = n28743 ^ n12387 ^ 1'b0 ;
  assign n28746 = n28745 ^ n28744 ^ 1'b0 ;
  assign n28747 = ~n28742 & n28746 ;
  assign n28748 = ~n26518 & n28747 ;
  assign n28749 = ( n5582 & n22897 ) | ( n5582 & ~n28748 ) | ( n22897 & ~n28748 ) ;
  assign n28750 = n19575 ^ n3663 ^ 1'b0 ;
  assign n28751 = n3928 | n28750 ;
  assign n28752 = n15200 ^ n7870 ^ 1'b0 ;
  assign n28753 = ~n1590 & n18308 ;
  assign n28754 = n4710 | n25756 ;
  assign n28755 = ( ~n9536 & n15810 ) | ( ~n9536 & n24803 ) | ( n15810 & n24803 ) ;
  assign n28756 = n4652 & ~n8402 ;
  assign n28757 = n6775 & n28756 ;
  assign n28758 = n8249 ^ n1739 ^ 1'b0 ;
  assign n28759 = ~n28757 & n28758 ;
  assign n28761 = n30 | n1431 ;
  assign n28762 = n1848 | n28761 ;
  assign n28763 = n25416 & n28762 ;
  assign n28764 = n28763 ^ n9808 ^ 1'b0 ;
  assign n28760 = ~n4334 & n11696 ;
  assign n28765 = n28764 ^ n28760 ^ 1'b0 ;
  assign n28766 = n335 & n28627 ;
  assign n28767 = n7767 & n28766 ;
  assign n28768 = n2848 | n28767 ;
  assign n28769 = n5323 & ~n28768 ;
  assign n28770 = n13974 & n19914 ;
  assign n28771 = n28770 ^ n22657 ^ 1'b0 ;
  assign n28772 = n6580 & ~n25208 ;
  assign n28773 = n28772 ^ n25407 ^ 1'b0 ;
  assign n28774 = n10678 ^ n330 ^ 1'b0 ;
  assign n28775 = n10815 & ~n28774 ;
  assign n28776 = ~n4604 & n5180 ;
  assign n28777 = n28775 & ~n28776 ;
  assign n28778 = n7943 | n14443 ;
  assign n28779 = n4392 | n28778 ;
  assign n28780 = n28779 ^ n2205 ^ 1'b0 ;
  assign n28781 = n6492 | n21778 ;
  assign n28782 = n28781 ^ n27757 ^ 1'b0 ;
  assign n28783 = ~n27635 & n28782 ;
  assign n28784 = n3115 | n4848 ;
  assign n28785 = n23145 | n28784 ;
  assign n28790 = n148 | n483 ;
  assign n28791 = n483 & ~n28790 ;
  assign n28792 = n697 & n861 ;
  assign n28793 = ~n697 & n28792 ;
  assign n28794 = n9864 ^ n1659 ^ 1'b0 ;
  assign n28795 = n28793 | n28794 ;
  assign n28796 = n28791 & ~n28795 ;
  assign n28797 = n774 & n28796 ;
  assign n28798 = n9455 & ~n28797 ;
  assign n28786 = n966 & n7681 ;
  assign n28787 = ~n966 & n28786 ;
  assign n28788 = ~n17246 & n28787 ;
  assign n28789 = n28788 ^ n11024 ^ 1'b0 ;
  assign n28799 = n28798 ^ n28789 ^ 1'b0 ;
  assign n28800 = n24334 | n28799 ;
  assign n28801 = n22188 ^ n18355 ^ 1'b0 ;
  assign n28802 = ~n28800 & n28801 ;
  assign n28803 = n873 | n2612 ;
  assign n28804 = n28803 ^ n3561 ^ 1'b0 ;
  assign n28805 = n4120 | n28804 ;
  assign n28806 = n28805 ^ n10627 ^ 1'b0 ;
  assign n28807 = n13389 & n14127 ;
  assign n28808 = n28807 ^ n3321 ^ 1'b0 ;
  assign n28809 = n7112 & ~n28287 ;
  assign n28810 = n11549 & n28809 ;
  assign n28811 = n11573 ^ n4088 ^ 1'b0 ;
  assign n28812 = ~n7427 & n12329 ;
  assign n28813 = n28812 ^ n7144 ^ 1'b0 ;
  assign n28814 = n14228 ^ n8692 ^ 1'b0 ;
  assign n28815 = n23449 & n28804 ;
  assign n28816 = n28815 ^ n679 ^ 1'b0 ;
  assign n28817 = ( n11203 & n28439 ) | ( n11203 & ~n28816 ) | ( n28439 & ~n28816 ) ;
  assign n28818 = n3764 & ~n23256 ;
  assign n28819 = n12651 & n28818 ;
  assign n28820 = n17218 & n28819 ;
  assign n28821 = n28251 & n28820 ;
  assign n28822 = n4246 & ~n12710 ;
  assign n28823 = ~n1479 & n28822 ;
  assign n28824 = n25940 & n28823 ;
  assign n28825 = n1676 & ~n17944 ;
  assign n28826 = n28825 ^ n599 ^ 1'b0 ;
  assign n28827 = ~n16525 & n28826 ;
  assign n28828 = n28827 ^ n754 ^ 1'b0 ;
  assign n28829 = ~n36 & n1854 ;
  assign n28830 = n28829 ^ n14884 ^ 1'b0 ;
  assign n28831 = n28323 | n28830 ;
  assign n28832 = n11164 & ~n28831 ;
  assign n28833 = n1884 & ~n17756 ;
  assign n28834 = n28833 ^ n10194 ^ 1'b0 ;
  assign n28835 = n7572 & ~n28834 ;
  assign n28836 = n20472 ^ n10509 ^ 1'b0 ;
  assign n28837 = ~n11766 & n28836 ;
  assign n28838 = n28837 ^ n10415 ^ 1'b0 ;
  assign n28839 = n20793 ^ n5929 ^ 1'b0 ;
  assign n28840 = n6933 & ~n10721 ;
  assign n28841 = ~n9756 & n28840 ;
  assign n28842 = n28841 ^ n883 ^ 1'b0 ;
  assign n28843 = ~n4363 & n11311 ;
  assign n28844 = n3407 | n27085 ;
  assign n28845 = n25943 ^ n15147 ^ 1'b0 ;
  assign n28846 = n129 & n28845 ;
  assign n28847 = ~n1428 & n23389 ;
  assign n28848 = n28847 ^ n14670 ^ 1'b0 ;
  assign n28849 = n895 | n28848 ;
  assign n28850 = ~n4683 & n13757 ;
  assign n28851 = n10180 | n18921 ;
  assign n28852 = n28850 | n28851 ;
  assign n28853 = n13086 | n26286 ;
  assign n28854 = n28853 ^ n7368 ^ 1'b0 ;
  assign n28855 = n28854 ^ n9143 ^ 1'b0 ;
  assign n28856 = n26146 & n28855 ;
  assign n28857 = n13992 ^ n3778 ^ 1'b0 ;
  assign n28858 = ~n3938 & n28857 ;
  assign n28859 = n4233 & n28227 ;
  assign n28860 = n28859 ^ n3262 ^ 1'b0 ;
  assign n28861 = n15625 ^ n12217 ^ 1'b0 ;
  assign n28862 = n19033 & ~n28861 ;
  assign n28863 = n7503 & n28862 ;
  assign n28864 = ( n141 & ~n3398 ) | ( n141 & n9207 ) | ( ~n3398 & n9207 ) ;
  assign n28865 = n26295 & n28864 ;
  assign n28866 = n12379 & n17176 ;
  assign n28867 = n28866 ^ n16840 ^ 1'b0 ;
  assign n28868 = n27935 ^ n3735 ^ 1'b0 ;
  assign n28869 = n28867 & ~n28868 ;
  assign n28870 = n15009 ^ n2239 ^ 1'b0 ;
  assign n28871 = ~n2450 & n22393 ;
  assign n28872 = n28871 ^ n17448 ^ 1'b0 ;
  assign n28873 = n8148 & ~n25543 ;
  assign n28874 = ~n4726 & n28873 ;
  assign n28875 = n1141 & n3322 ;
  assign n28876 = ~n7622 & n15244 ;
  assign n28877 = n28876 ^ n17383 ^ 1'b0 ;
  assign n28878 = n22374 ^ n2116 ^ 1'b0 ;
  assign n28879 = n19229 & ~n20596 ;
  assign n28880 = n24418 ^ n17584 ^ 1'b0 ;
  assign n28881 = ~n458 & n28880 ;
  assign n28882 = n28881 ^ n10126 ^ 1'b0 ;
  assign n28883 = n28879 | n28882 ;
  assign n28884 = n15307 | n28883 ;
  assign n28885 = n28884 ^ n5566 ^ 1'b0 ;
  assign n28886 = n10217 ^ n8091 ^ 1'b0 ;
  assign n28887 = n28886 ^ n9364 ^ 1'b0 ;
  assign n28888 = ~n1480 & n1937 ;
  assign n28889 = n5011 & n28888 ;
  assign n28890 = n28889 ^ n6168 ^ 1'b0 ;
  assign n28891 = n5709 ^ n1946 ^ 1'b0 ;
  assign n28893 = n6999 ^ n2311 ^ 1'b0 ;
  assign n28894 = n2618 & ~n28893 ;
  assign n28892 = n4320 | n9957 ;
  assign n28895 = n28894 ^ n28892 ^ 1'b0 ;
  assign n28896 = n24559 & ~n28895 ;
  assign n28897 = n1817 | n25133 ;
  assign n28898 = ~n3939 & n9934 ;
  assign n28899 = n28898 ^ n18772 ^ 1'b0 ;
  assign n28900 = n8570 & ~n24611 ;
  assign n28901 = n5697 & n9542 ;
  assign n28902 = n542 & ~n9406 ;
  assign n28903 = n28121 ^ n18348 ^ 1'b0 ;
  assign n28904 = n18305 & n28903 ;
  assign n28905 = n11334 | n13083 ;
  assign n28906 = ~n6376 & n7960 ;
  assign n28907 = ~n13923 & n28906 ;
  assign n28908 = n28907 ^ n4419 ^ 1'b0 ;
  assign n28909 = n748 | n7495 ;
  assign n28910 = n1349 | n26796 ;
  assign n28911 = n28910 ^ n22737 ^ 1'b0 ;
  assign n28912 = n11039 & ~n16786 ;
  assign n28913 = n14184 ^ n3735 ^ 1'b0 ;
  assign n28914 = n10934 | n28623 ;
  assign n28915 = n7026 & ~n9779 ;
  assign n28916 = n28915 ^ n6498 ^ 1'b0 ;
  assign n28917 = n4934 & n28916 ;
  assign n28918 = n1019 ^ n1016 ^ 1'b0 ;
  assign n28919 = ~n4580 & n28918 ;
  assign n28920 = ~n16091 & n28919 ;
  assign n28921 = ~n28917 & n28920 ;
  assign n28922 = n7282 & ~n17020 ;
  assign n28923 = n630 & ~n28922 ;
  assign n28924 = ~n1108 & n28923 ;
  assign n28925 = n8290 | n26120 ;
  assign n28926 = n15117 & ~n28925 ;
  assign n28927 = n988 | n9461 ;
  assign n28928 = n7082 | n28927 ;
  assign n28929 = n542 | n14665 ;
  assign n28930 = n9162 & ~n16625 ;
  assign n28932 = n7449 & n16120 ;
  assign n28933 = n28932 ^ n11159 ^ 1'b0 ;
  assign n28931 = n13939 | n20505 ;
  assign n28934 = n28933 ^ n28931 ^ 1'b0 ;
  assign n28935 = n3219 & n28306 ;
  assign n28936 = n28935 ^ n12546 ^ 1'b0 ;
  assign n28937 = n6503 & ~n12553 ;
  assign n28938 = n28936 & n28937 ;
  assign n28939 = n10274 ^ n3074 ^ 1'b0 ;
  assign n28940 = n2547 | n28208 ;
  assign n28941 = ~n2787 & n23032 ;
  assign n28942 = n28941 ^ n20563 ^ 1'b0 ;
  assign n28943 = n3826 ^ n924 ^ 1'b0 ;
  assign n28944 = n2785 | n28943 ;
  assign n28945 = ~n12184 & n28944 ;
  assign n28946 = n1087 & ~n2463 ;
  assign n28947 = n28946 ^ n2964 ^ 1'b0 ;
  assign n28948 = n14495 ^ n2138 ^ 1'b0 ;
  assign n28949 = n469 & ~n28948 ;
  assign n28950 = n28949 ^ n9654 ^ 1'b0 ;
  assign n28951 = n7149 ^ n25 ^ 1'b0 ;
  assign n28952 = ~n5182 & n16504 ;
  assign n28953 = n498 & ~n7118 ;
  assign n28954 = ~n23325 & n28953 ;
  assign n28955 = n16506 | n28954 ;
  assign n28956 = n25526 ^ n16585 ^ 1'b0 ;
  assign n28957 = n28956 ^ n13963 ^ 1'b0 ;
  assign n28958 = ~n3732 & n28957 ;
  assign n28959 = n2722 & ~n7462 ;
  assign n28960 = n1832 & ~n6281 ;
  assign n28961 = n21815 ^ n2817 ^ n882 ;
  assign n28962 = n294 & ~n1718 ;
  assign n28965 = n11494 ^ n3744 ^ 1'b0 ;
  assign n28963 = n562 ^ n339 ^ 1'b0 ;
  assign n28964 = n278 & ~n28963 ;
  assign n28966 = n28965 ^ n28964 ^ n7160 ;
  assign n28967 = n28966 ^ n11044 ^ 1'b0 ;
  assign n28968 = n16764 ^ n4300 ^ 1'b0 ;
  assign n28969 = n28968 ^ n1233 ^ 1'b0 ;
  assign n28970 = ~n16193 & n17638 ;
  assign n28971 = n28970 ^ n741 ^ 1'b0 ;
  assign n28972 = n4904 ^ n3524 ^ 1'b0 ;
  assign n28973 = n28972 ^ n1258 ^ 1'b0 ;
  assign n28974 = n12300 & ~n28973 ;
  assign n28975 = n2542 ^ n2148 ^ 1'b0 ;
  assign n28976 = n28975 ^ n11298 ^ n5376 ;
  assign n28977 = ~n578 & n14986 ;
  assign n28978 = n13781 & n28977 ;
  assign n28979 = n594 & n1572 ;
  assign n28980 = n5138 ^ n833 ^ 1'b0 ;
  assign n28981 = ~n28979 & n28980 ;
  assign n28982 = n9837 & n12873 ;
  assign n28983 = n28982 ^ n9593 ^ 1'b0 ;
  assign n28984 = n28983 ^ n15649 ^ 1'b0 ;
  assign n28985 = n257 | n15457 ;
  assign n28986 = n28985 ^ n4191 ^ 1'b0 ;
  assign n28987 = n11463 & ~n11680 ;
  assign n28988 = ~n3007 & n28987 ;
  assign n28989 = n104 & ~n28988 ;
  assign n28990 = ~n4749 & n28989 ;
  assign n28991 = n11076 ^ n1878 ^ 1'b0 ;
  assign n28992 = ~n7503 & n28991 ;
  assign n28993 = n25709 & ~n28992 ;
  assign n28994 = n14616 ^ n7234 ^ 1'b0 ;
  assign n28995 = n1479 & n28994 ;
  assign n28996 = n28995 ^ n1406 ^ 1'b0 ;
  assign n28997 = n509 & n28996 ;
  assign n28998 = n653 | n2924 ;
  assign n28999 = ~n11753 & n28998 ;
  assign n29000 = n22665 ^ n1125 ^ 1'b0 ;
  assign n29001 = n9741 | n29000 ;
  assign n29002 = n848 | n29001 ;
  assign n29003 = n3666 | n27861 ;
  assign n29004 = n8079 & n8705 ;
  assign n29005 = ~n6287 & n29004 ;
  assign n29007 = ( n9159 & ~n10137 ) | ( n9159 & n28133 ) | ( ~n10137 & n28133 ) ;
  assign n29006 = ~n2401 & n3548 ;
  assign n29008 = n29007 ^ n29006 ^ 1'b0 ;
  assign n29009 = n29008 ^ n13590 ^ 1'b0 ;
  assign n29010 = n2524 | n8725 ;
  assign n29011 = n1323 | n20148 ;
  assign n29012 = n20275 ^ n6019 ^ 1'b0 ;
  assign n29013 = ~n27228 & n29012 ;
  assign n29014 = ~n5083 & n7879 ;
  assign n29015 = n8148 ^ n6421 ^ 1'b0 ;
  assign n29017 = n10409 ^ n3735 ^ n1895 ;
  assign n29016 = n2660 | n20472 ;
  assign n29018 = n29017 ^ n29016 ^ 1'b0 ;
  assign n29019 = n29018 ^ n22907 ^ 1'b0 ;
  assign n29020 = n29019 ^ n24356 ^ 1'b0 ;
  assign n29021 = n6082 & n14055 ;
  assign n29022 = n29021 ^ n2430 ^ 1'b0 ;
  assign n29023 = n52 | n29022 ;
  assign n29024 = n29020 | n29023 ;
  assign n29025 = n1838 & n4314 ;
  assign n29026 = n24651 & n29025 ;
  assign n29027 = n1529 & ~n12702 ;
  assign n29028 = n8517 & n29027 ;
  assign n29029 = n29028 ^ n5010 ^ 1'b0 ;
  assign n29030 = n29029 ^ n15932 ^ 1'b0 ;
  assign n29031 = n6432 & ~n29030 ;
  assign n29032 = n10718 & ~n16090 ;
  assign n29033 = n630 | n1947 ;
  assign n29034 = n827 | n28296 ;
  assign n29035 = n16773 | n29034 ;
  assign n29036 = n29033 | n29035 ;
  assign n29037 = n22481 ^ n4668 ^ 1'b0 ;
  assign n29038 = n13994 ^ n13063 ^ 1'b0 ;
  assign n29039 = ~n13088 & n29038 ;
  assign n29040 = n16491 | n20659 ;
  assign n29041 = n29039 | n29040 ;
  assign n29042 = n27570 ^ n11797 ^ 1'b0 ;
  assign n29043 = n9220 & ~n29042 ;
  assign n29044 = n2667 ^ n1810 ^ 1'b0 ;
  assign n29045 = n252 & n29044 ;
  assign n29046 = ~n7348 & n17857 ;
  assign n29047 = n10635 & n29046 ;
  assign n29048 = n29047 ^ n20774 ^ 1'b0 ;
  assign n29049 = ~n10298 & n28970 ;
  assign n29050 = n15892 ^ n3663 ^ 1'b0 ;
  assign n29051 = n7130 & n29050 ;
  assign n29052 = n29051 ^ n3812 ^ 1'b0 ;
  assign n29053 = n2268 | n4264 ;
  assign n29054 = n28335 ^ n13878 ^ 1'b0 ;
  assign n29055 = n25721 ^ n903 ^ 1'b0 ;
  assign n29056 = n20472 ^ n7665 ^ 1'b0 ;
  assign n29057 = n14225 ^ n1112 ^ 1'b0 ;
  assign n29058 = n29057 ^ n8589 ^ 1'b0 ;
  assign n29059 = n4640 & ~n29058 ;
  assign n29060 = ~n29056 & n29059 ;
  assign n29061 = n10194 ^ n4874 ^ 1'b0 ;
  assign n29062 = n25063 & ~n29061 ;
  assign n29063 = n29060 & n29062 ;
  assign n29064 = ~n55 & n4917 ;
  assign n29065 = n5603 ^ n1473 ^ 1'b0 ;
  assign n29066 = n390 & ~n29065 ;
  assign n29067 = n29066 ^ n6595 ^ 1'b0 ;
  assign n29068 = n5992 ^ n2842 ^ 1'b0 ;
  assign n29069 = n23848 ^ n10651 ^ 1'b0 ;
  assign n29070 = n29068 & n29069 ;
  assign n29073 = n5018 & n10195 ;
  assign n29074 = n29073 ^ n8219 ^ 1'b0 ;
  assign n29071 = n5012 | n13046 ;
  assign n29072 = n20284 & n29071 ;
  assign n29075 = n29074 ^ n29072 ^ 1'b0 ;
  assign n29076 = n8502 & ~n9039 ;
  assign n29077 = n29076 ^ n7475 ^ 1'b0 ;
  assign n29078 = ~n6365 & n29077 ;
  assign n29079 = n29078 ^ n1263 ^ 1'b0 ;
  assign n29080 = n24045 ^ n11630 ^ 1'b0 ;
  assign n29081 = ~n21367 & n29080 ;
  assign n29082 = n562 & n9492 ;
  assign n29083 = n5823 & n29082 ;
  assign n29084 = n17961 ^ n17479 ^ 1'b0 ;
  assign n29085 = n13198 ^ n288 ^ 1'b0 ;
  assign n29086 = n489 | n4696 ;
  assign n29087 = n6651 | n7056 ;
  assign n29088 = n2734 | n12515 ;
  assign n29089 = n29088 ^ n15422 ^ 1'b0 ;
  assign n29090 = ~n382 & n7286 ;
  assign n29091 = n29090 ^ n2194 ^ 1'b0 ;
  assign n29092 = ~n14528 & n29091 ;
  assign n29093 = ~n19437 & n29092 ;
  assign n29094 = n29093 ^ n18186 ^ 1'b0 ;
  assign n29095 = n26575 & n28366 ;
  assign n29096 = n10721 ^ n2335 ^ 1'b0 ;
  assign n29097 = n6244 | n29096 ;
  assign n29098 = n29097 ^ n364 ^ 1'b0 ;
  assign n29099 = n26591 & ~n29098 ;
  assign n29100 = n9739 ^ n2571 ^ 1'b0 ;
  assign n29101 = n861 ^ n483 ^ 1'b0 ;
  assign n29102 = n7594 & ~n19559 ;
  assign n29103 = n6921 ^ n671 ^ 1'b0 ;
  assign n29104 = n12489 | n13420 ;
  assign n29105 = ~n29103 & n29104 ;
  assign n29106 = n1250 & n12732 ;
  assign n29107 = ~n16126 & n29106 ;
  assign n29108 = ~n10632 & n23997 ;
  assign n29109 = n29107 | n29108 ;
  assign n29110 = n8262 | n26213 ;
  assign n29111 = n984 & n3620 ;
  assign n29112 = ~n22700 & n29111 ;
  assign n29113 = n29112 ^ n4401 ^ 1'b0 ;
  assign n29114 = n12368 & ~n13160 ;
  assign n29115 = n29114 ^ n153 ^ 1'b0 ;
  assign n29116 = ~n568 & n22257 ;
  assign n29117 = n1950 & ~n4840 ;
  assign n29118 = n29117 ^ n6333 ^ 1'b0 ;
  assign n29119 = n21023 & ~n29118 ;
  assign n29120 = n23171 ^ n10784 ^ n278 ;
  assign n29121 = n1711 | n18016 ;
  assign n29122 = n16086 & ~n29121 ;
  assign n29123 = n6162 & ~n9332 ;
  assign n29124 = n10637 & ~n14998 ;
  assign n29125 = n4361 ^ n722 ^ 1'b0 ;
  assign n29126 = n29125 ^ n24841 ^ 1'b0 ;
  assign n29127 = n13855 ^ n10286 ^ n4641 ;
  assign n29128 = ~n12470 & n29127 ;
  assign n29129 = n29128 ^ n10815 ^ 1'b0 ;
  assign n29130 = n29129 ^ n5065 ^ 1'b0 ;
  assign n29131 = n6371 & n7792 ;
  assign n29132 = n10647 & n29131 ;
  assign n29133 = n12123 & ~n29132 ;
  assign n29135 = ~n246 & n2674 ;
  assign n29134 = ~n10136 & n17997 ;
  assign n29136 = n29135 ^ n29134 ^ 1'b0 ;
  assign n29137 = n16658 ^ n5871 ^ 1'b0 ;
  assign n29138 = ~n13564 & n29137 ;
  assign n29139 = n14185 & n29138 ;
  assign n29140 = n6141 ^ n5193 ^ 1'b0 ;
  assign n29141 = n7952 ^ n2569 ^ 1'b0 ;
  assign n29142 = n4196 & ~n29141 ;
  assign n29143 = n8389 & ~n12817 ;
  assign n29144 = n4063 & n14236 ;
  assign n29145 = n4482 & n29144 ;
  assign n29146 = n29145 ^ n25267 ^ 1'b0 ;
  assign n29147 = n20506 ^ n7124 ^ 1'b0 ;
  assign n29148 = n917 & ~n29147 ;
  assign n29149 = ( n6870 & n17361 ) | ( n6870 & n29148 ) | ( n17361 & n29148 ) ;
  assign n29150 = n2769 & ~n15271 ;
  assign n29151 = n1246 & ~n1710 ;
  assign n29152 = n5283 | n15605 ;
  assign n29153 = n7227 ^ n5943 ^ 1'b0 ;
  assign n29154 = n378 & n29153 ;
  assign n29155 = n23796 ^ n2130 ^ 1'b0 ;
  assign n29156 = n5905 & n14645 ;
  assign n29157 = n29155 & n29156 ;
  assign n29158 = n23594 ^ n297 ^ 1'b0 ;
  assign n29159 = ~n3915 & n9197 ;
  assign n29160 = n29159 ^ n13875 ^ 1'b0 ;
  assign n29161 = n11588 | n29160 ;
  assign n29162 = n9883 | n29161 ;
  assign n29163 = n29162 ^ n1958 ^ 1'b0 ;
  assign n29164 = n7540 & n29163 ;
  assign n29165 = n8409 & ~n27162 ;
  assign n29166 = ~n6876 & n11434 ;
  assign n29167 = n3369 | n29166 ;
  assign n29168 = n29167 ^ n6565 ^ 1'b0 ;
  assign n29169 = n297 & n29168 ;
  assign n29170 = n7732 ^ n5031 ^ 1'b0 ;
  assign n29171 = ~n5887 & n29170 ;
  assign n29172 = ~n2893 & n6284 ;
  assign n29173 = n24473 | n29172 ;
  assign n29174 = n16070 ^ n5103 ^ 1'b0 ;
  assign n29175 = n1245 | n29174 ;
  assign n29176 = n364 | n5347 ;
  assign n29177 = n6884 & n8654 ;
  assign n29178 = n29177 ^ n7730 ^ 1'b0 ;
  assign n29179 = n25766 | n29178 ;
  assign n29180 = ~n12310 & n16719 ;
  assign n29181 = n29180 ^ n9814 ^ 1'b0 ;
  assign n29182 = n22282 & n29181 ;
  assign n29183 = n9512 ^ n8662 ^ 1'b0 ;
  assign n29184 = n128 & ~n29183 ;
  assign n29185 = ~n1054 & n29184 ;
  assign n29186 = n29185 ^ n20557 ^ 1'b0 ;
  assign n29187 = ~n15395 & n29186 ;
  assign n29188 = n4350 & ~n13083 ;
  assign n29189 = n29188 ^ n5839 ^ 1'b0 ;
  assign n29190 = n10357 & n29189 ;
  assign n29191 = n29190 ^ n17647 ^ 1'b0 ;
  assign n29192 = ~n12310 & n29191 ;
  assign n29197 = n6414 ^ n3542 ^ 1'b0 ;
  assign n29194 = n318 | n20102 ;
  assign n29195 = n24698 | n29194 ;
  assign n29193 = ~n14606 & n21406 ;
  assign n29196 = n29195 ^ n29193 ^ 1'b0 ;
  assign n29198 = n29197 ^ n29196 ^ n13164 ;
  assign n29199 = n2714 ^ n1844 ^ 1'b0 ;
  assign n29202 = n22554 ^ n9124 ^ 1'b0 ;
  assign n29200 = n27869 ^ n22108 ^ 1'b0 ;
  assign n29201 = ~n2328 & n29200 ;
  assign n29203 = n29202 ^ n29201 ^ 1'b0 ;
  assign n29204 = n5527 & ~n7501 ;
  assign n29206 = n7459 ^ n3431 ^ 1'b0 ;
  assign n29205 = n6722 & n12416 ;
  assign n29207 = n29206 ^ n29205 ^ 1'b0 ;
  assign n29208 = n29207 ^ n24360 ^ 1'b0 ;
  assign n29209 = n21999 ^ n15045 ^ n10936 ;
  assign n29210 = ~n19210 & n21764 ;
  assign n29211 = n481 | n19710 ;
  assign n29212 = ~n26655 & n29211 ;
  assign n29215 = n1645 & n5053 ;
  assign n29216 = n11677 & n29215 ;
  assign n29213 = n15087 ^ n2060 ^ 1'b0 ;
  assign n29214 = n823 & n29213 ;
  assign n29217 = n29216 ^ n29214 ^ 1'b0 ;
  assign n29218 = n15377 & ~n29217 ;
  assign n29219 = n1565 & n29218 ;
  assign n29220 = ~n3781 & n15785 ;
  assign n29221 = n29220 ^ n21244 ^ n3061 ;
  assign n29222 = n2595 & ~n15542 ;
  assign n29223 = n19674 & n28512 ;
  assign n29224 = ~n384 & n29223 ;
  assign n29225 = n2842 & n3245 ;
  assign n29226 = n29225 ^ n4270 ^ 1'b0 ;
  assign n29227 = n29226 ^ n24041 ^ n20238 ;
  assign n29228 = ~n17255 & n29227 ;
  assign n29229 = n25159 & ~n26575 ;
  assign n29230 = n13933 ^ n12743 ^ 1'b0 ;
  assign n29231 = n7386 | n29230 ;
  assign n29232 = n29231 ^ n9309 ^ 1'b0 ;
  assign n29233 = ~n782 & n28968 ;
  assign n29234 = n2662 & ~n27973 ;
  assign n29235 = n2606 & n12215 ;
  assign n29236 = ~n25557 & n29235 ;
  assign n29237 = n10590 ^ n524 ^ 1'b0 ;
  assign n29238 = ~n512 & n2542 ;
  assign n29239 = n29238 ^ n1913 ^ 1'b0 ;
  assign n29240 = n1419 & n29239 ;
  assign n29241 = n18466 ^ n16712 ^ 1'b0 ;
  assign n29242 = n6150 ^ n2476 ^ n2029 ;
  assign n29243 = ~n4108 & n17259 ;
  assign n29244 = n29242 | n29243 ;
  assign n29245 = n29241 | n29244 ;
  assign n29246 = n3197 ^ n1368 ^ 1'b0 ;
  assign n29247 = n4319 & n13741 ;
  assign n29248 = n24185 ^ n20487 ^ 1'b0 ;
  assign n29249 = ~n29247 & n29248 ;
  assign n29250 = n4521 ^ n3134 ^ 1'b0 ;
  assign n29251 = n1191 & ~n28968 ;
  assign n29252 = n20097 & n22967 ;
  assign n29253 = n29252 ^ n16226 ^ 1'b0 ;
  assign n29254 = n10500 & n29253 ;
  assign n29255 = n815 & ~n29254 ;
  assign n29256 = n29255 ^ n5143 ^ 1'b0 ;
  assign n29257 = n3353 | n6136 ;
  assign n29258 = n23485 ^ n8763 ^ 1'b0 ;
  assign n29259 = ~n24097 & n29258 ;
  assign n29260 = n21384 ^ n4915 ^ 1'b0 ;
  assign n29261 = n11042 & n29260 ;
  assign n29262 = n19911 ^ n6163 ^ 1'b0 ;
  assign n29263 = ~n1687 & n29262 ;
  assign n29264 = n29263 ^ n7734 ^ 1'b0 ;
  assign n29265 = n3366 | n9697 ;
  assign n29266 = n6282 ^ n141 ^ 1'b0 ;
  assign n29267 = n7051 & ~n29266 ;
  assign n29268 = ~n395 & n5586 ;
  assign n29269 = n21427 ^ n1192 ^ 1'b0 ;
  assign n29270 = n15451 & n29269 ;
  assign n29271 = n20105 & n29270 ;
  assign n29272 = n2900 ^ n989 ^ 1'b0 ;
  assign n29273 = n3292 ^ n2134 ^ 1'b0 ;
  assign n29274 = n29272 & ~n29273 ;
  assign n29275 = n832 ^ n760 ^ 1'b0 ;
  assign n29276 = n23783 & ~n29275 ;
  assign n29277 = n29274 & n29276 ;
  assign n29278 = n3260 ^ n2813 ^ 1'b0 ;
  assign n29279 = n22949 ^ n17127 ^ 1'b0 ;
  assign n29280 = n20795 & ~n29279 ;
  assign n29281 = n29280 ^ n28670 ^ 1'b0 ;
  assign n29282 = ~n3616 & n8840 ;
  assign n29283 = ~n19042 & n29282 ;
  assign n29284 = ~n129 & n29283 ;
  assign n29285 = n12180 & ~n20332 ;
  assign n29286 = n12237 & n29285 ;
  assign n29287 = n3611 & n11376 ;
  assign n29288 = n1747 & ~n7406 ;
  assign n29289 = n22479 ^ n19363 ^ 1'b0 ;
  assign n29290 = n15159 ^ n1112 ^ 1'b0 ;
  assign n29291 = n11412 & n23235 ;
  assign n29292 = n12313 ^ n4367 ^ 1'b0 ;
  assign n29293 = n10292 & ~n29292 ;
  assign n29294 = ~n5033 & n29293 ;
  assign n29295 = n615 & ~n2825 ;
  assign n29296 = n29294 & n29295 ;
  assign n29297 = n839 & ~n9880 ;
  assign n29298 = n21195 & ~n29297 ;
  assign n29299 = n29296 & n29298 ;
  assign n29300 = ~n1521 & n14337 ;
  assign n29302 = n3784 & ~n4533 ;
  assign n29301 = n11174 | n17452 ;
  assign n29303 = n29302 ^ n29301 ^ 1'b0 ;
  assign n29306 = n675 & ~n5330 ;
  assign n29307 = ~n9548 & n29306 ;
  assign n29308 = n29307 ^ n14865 ^ 1'b0 ;
  assign n29309 = ~n10765 & n29308 ;
  assign n29310 = n29309 ^ n378 ^ 1'b0 ;
  assign n29304 = n14571 ^ n8587 ^ 1'b0 ;
  assign n29305 = ~n2835 & n29304 ;
  assign n29311 = n29310 ^ n29305 ^ 1'b0 ;
  assign n29312 = n9108 & n29311 ;
  assign n29313 = n1769 & n29312 ;
  assign n29314 = ~n458 & n584 ;
  assign n29315 = ~n584 & n29314 ;
  assign n29316 = n9162 | n29315 ;
  assign n29317 = n29315 & ~n29316 ;
  assign n29318 = ~n5428 & n9843 ;
  assign n29319 = n29318 ^ n19565 ^ 1'b0 ;
  assign n29320 = n14265 & ~n19404 ;
  assign n29321 = n13501 & n29320 ;
  assign n29322 = n13801 | n24465 ;
  assign n29323 = n29322 ^ n25878 ^ 1'b0 ;
  assign n29324 = n2558 ^ n513 ^ 1'b0 ;
  assign n29325 = ~n15528 & n29324 ;
  assign n29326 = n4640 & ~n29325 ;
  assign n29327 = n108 | n148 ;
  assign n29328 = n148 & ~n29327 ;
  assign n29329 = ~n19 & n14281 ;
  assign n29330 = n1105 & ~n17409 ;
  assign n29331 = ~n29329 & n29330 ;
  assign n29332 = n29328 & ~n29331 ;
  assign n29333 = n29332 ^ n1827 ^ 1'b0 ;
  assign n29334 = n3433 ^ n2254 ^ 1'b0 ;
  assign n29335 = ~n29333 & n29334 ;
  assign n29336 = n29335 ^ n6062 ^ 1'b0 ;
  assign n29337 = n29326 & n29336 ;
  assign n29338 = n12458 ^ n9240 ^ 1'b0 ;
  assign n29339 = n7596 ^ n3104 ^ 1'b0 ;
  assign n29340 = n29338 & n29339 ;
  assign n29341 = n22447 ^ n5254 ^ n2767 ;
  assign n29343 = n6488 ^ n6464 ^ 1'b0 ;
  assign n29344 = n8365 & n29343 ;
  assign n29342 = n16528 ^ n1877 ^ 1'b0 ;
  assign n29345 = n29344 ^ n29342 ^ 1'b0 ;
  assign n29346 = n24366 ^ n16090 ^ 1'b0 ;
  assign n29347 = n29345 & n29346 ;
  assign n29348 = n6509 ^ n1531 ^ 1'b0 ;
  assign n29349 = n5957 ^ n3007 ^ 1'b0 ;
  assign n29350 = n6250 & ~n14730 ;
  assign n29351 = n3595 ^ n732 ^ 1'b0 ;
  assign n29352 = n29350 & ~n29351 ;
  assign n29353 = n1741 ^ n963 ^ 1'b0 ;
  assign n29354 = ~n2842 & n29353 ;
  assign n29355 = n4401 ^ n2474 ^ 1'b0 ;
  assign n29356 = ~n669 & n29355 ;
  assign n29358 = n5221 & n11761 ;
  assign n29357 = n2853 & n4966 ;
  assign n29359 = n29358 ^ n29357 ^ n5128 ;
  assign n29360 = n104 & ~n29359 ;
  assign n29361 = ~n28979 & n29360 ;
  assign n29362 = n3367 & n29361 ;
  assign n29363 = n310 & n28194 ;
  assign n29364 = ~n3395 & n29363 ;
  assign n29365 = n12866 & n29364 ;
  assign n29366 = n8128 ^ n8106 ^ 1'b0 ;
  assign n29367 = n29366 ^ n2415 ^ 1'b0 ;
  assign n29368 = ~n7822 & n29367 ;
  assign n29372 = n9419 | n12118 ;
  assign n29373 = ( ~n3338 & n6436 ) | ( ~n3338 & n29372 ) | ( n6436 & n29372 ) ;
  assign n29369 = n2090 & ~n6529 ;
  assign n29370 = n29369 ^ n9015 ^ 1'b0 ;
  assign n29371 = n23103 | n29370 ;
  assign n29374 = n29373 ^ n29371 ^ 1'b0 ;
  assign n29375 = n21426 ^ n16321 ^ 1'b0 ;
  assign n29376 = n4214 | n20054 ;
  assign n29377 = ~n5535 & n19144 ;
  assign n29378 = n15547 & ~n29066 ;
  assign n29379 = ~n18471 & n29378 ;
  assign n29380 = n12363 | n29379 ;
  assign n29381 = n4748 ^ n3887 ^ 1'b0 ;
  assign n29382 = n4939 ^ n246 ^ 1'b0 ;
  assign n29383 = n2991 | n29382 ;
  assign n29384 = n931 & n29383 ;
  assign n29385 = n5439 ^ n4203 ^ 1'b0 ;
  assign n29386 = n5284 | n29385 ;
  assign n29387 = n6901 | n10957 ;
  assign n29388 = n14571 | n29387 ;
  assign n29389 = n29388 ^ n7360 ^ 1'b0 ;
  assign n29390 = n8946 & ~n29389 ;
  assign n29391 = n7915 ^ n7180 ^ 1'b0 ;
  assign n29392 = n5990 & ~n29391 ;
  assign n29393 = n8056 ^ n6424 ^ 1'b0 ;
  assign n29394 = n27606 & ~n29393 ;
  assign n29395 = n5713 ^ n1105 ^ 1'b0 ;
  assign n29396 = n281 & ~n29395 ;
  assign n29397 = n29396 ^ n1106 ^ 1'b0 ;
  assign n29398 = n751 & n1335 ;
  assign n29399 = ~n751 & n29398 ;
  assign n29400 = n374 | n29399 ;
  assign n29401 = n374 & ~n29400 ;
  assign n29402 = n957 & ~n2680 ;
  assign n29403 = ~n957 & n29402 ;
  assign n29404 = n278 & ~n29403 ;
  assign n29405 = n29401 & n29404 ;
  assign n29406 = ~n141 & n2415 ;
  assign n29407 = n29405 & n29406 ;
  assign n29408 = n3444 | n29407 ;
  assign n29409 = n29407 & ~n29408 ;
  assign n29410 = ~n29397 & n29409 ;
  assign n29411 = ~x2 & n7450 ;
  assign n29412 = ~n7450 & n29411 ;
  assign n29413 = n12299 | n29412 ;
  assign n29414 = n12299 & ~n29413 ;
  assign n29415 = n17528 & ~n29414 ;
  assign n29416 = ~n29410 & n29415 ;
  assign n29418 = n11585 & n14171 ;
  assign n29417 = x6 & ~n17247 ;
  assign n29419 = n29418 ^ n29417 ^ 1'b0 ;
  assign n29420 = ~n24599 & n29419 ;
  assign n29421 = n18114 ^ n14766 ^ 1'b0 ;
  assign n29422 = n16250 & n21810 ;
  assign n29423 = ~n6885 & n29422 ;
  assign n29424 = n29423 ^ n9858 ^ 1'b0 ;
  assign n29425 = n1900 | n29424 ;
  assign n29426 = n16838 | n27302 ;
  assign n29427 = ~n9845 & n15872 ;
  assign n29428 = n29427 ^ n11309 ^ 1'b0 ;
  assign n29429 = n10833 & ~n13420 ;
  assign n29431 = n3405 | n16060 ;
  assign n29432 = n10228 & ~n29431 ;
  assign n29433 = n12316 & ~n29432 ;
  assign n29434 = ~n456 & n29433 ;
  assign n29435 = n12883 & n29434 ;
  assign n29430 = n4051 & ~n4421 ;
  assign n29436 = n29435 ^ n29430 ^ 1'b0 ;
  assign n29437 = n7935 & n23159 ;
  assign n29438 = n973 & ~n23590 ;
  assign n29439 = n3211 ^ n1027 ^ n294 ;
  assign n29440 = n24383 & ~n29439 ;
  assign n29441 = n1840 ^ n856 ^ n442 ;
  assign n29442 = n25551 ^ n3354 ^ 1'b0 ;
  assign n29443 = n11802 & n29442 ;
  assign n29444 = ( n12680 & ~n21617 ) | ( n12680 & n29443 ) | ( ~n21617 & n29443 ) ;
  assign n29445 = n257 & ~n15923 ;
  assign n29446 = n6291 ^ n4233 ^ 1'b0 ;
  assign n29447 = ~n68 & n29446 ;
  assign n29448 = n7467 & n13720 ;
  assign n29449 = n15185 | n29448 ;
  assign n29450 = n2409 | n29449 ;
  assign n29451 = n15137 ^ n279 ^ 1'b0 ;
  assign n29452 = n8703 | n17526 ;
  assign n29453 = ( n10394 & n12123 ) | ( n10394 & n14125 ) | ( n12123 & n14125 ) ;
  assign n29454 = n10794 & ~n17172 ;
  assign n29455 = n3014 ^ n1697 ^ 1'b0 ;
  assign n29456 = ~n21953 & n29455 ;
  assign n29457 = n8145 & ~n11537 ;
  assign n29458 = n27508 & ~n29457 ;
  assign n29459 = n29457 & n29458 ;
  assign n29460 = n22461 ^ n10685 ^ 1'b0 ;
  assign n29461 = n3729 & ~n21100 ;
  assign n29462 = n29461 ^ n26342 ^ 1'b0 ;
  assign n29463 = ~n17882 & n29462 ;
  assign n29464 = n19356 ^ n15555 ^ 1'b0 ;
  assign n29465 = n7704 & ~n29464 ;
  assign n29466 = n4586 & n5345 ;
  assign n29467 = n113 & ~n29466 ;
  assign n29468 = ~n2512 & n29467 ;
  assign n29469 = n29465 | n29468 ;
  assign n29470 = n27174 ^ n20055 ^ n11975 ;
  assign n29471 = n867 & ~n25177 ;
  assign n29472 = n13456 ^ n7424 ^ 1'b0 ;
  assign n29473 = n9120 & n12738 ;
  assign n29474 = ~n899 & n29473 ;
  assign n29475 = ~n302 & n2121 ;
  assign n29476 = n19045 & n29475 ;
  assign n29477 = ~n2860 & n6217 ;
  assign n29478 = ~n29476 & n29477 ;
  assign n29479 = n15759 & ~n16407 ;
  assign n29480 = ~n14824 & n29479 ;
  assign n29481 = ( n10158 & ~n27334 ) | ( n10158 & n29480 ) | ( ~n27334 & n29480 ) ;
  assign n29482 = n10266 & n23691 ;
  assign n29483 = n11865 & n29482 ;
  assign n29484 = n16753 & n28745 ;
  assign n29485 = n7970 & ~n9966 ;
  assign n29486 = ~n17941 & n29485 ;
  assign n29487 = n1347 | n12982 ;
  assign n29488 = n29486 & ~n29487 ;
  assign n29489 = n2129 | n3598 ;
  assign n29490 = n11712 ^ n2572 ^ 1'b0 ;
  assign n29491 = n29489 | n29490 ;
  assign n29492 = n12255 ^ n1674 ^ 1'b0 ;
  assign n29493 = ~n3527 & n25633 ;
  assign n29494 = ~n29492 & n29493 ;
  assign n29495 = ~n19152 & n29494 ;
  assign n29496 = n14091 ^ n2129 ^ 1'b0 ;
  assign n29497 = n18339 & ~n29496 ;
  assign n29498 = n1693 ^ n294 ^ 1'b0 ;
  assign n29499 = n14941 & n29498 ;
  assign n29500 = ~n12299 & n29499 ;
  assign n29501 = n29500 ^ n14225 ^ 1'b0 ;
  assign n29502 = n8959 & n24628 ;
  assign n29503 = n5923 & n29502 ;
  assign n29504 = n13389 ^ n2092 ^ 1'b0 ;
  assign n29505 = n24983 & n29504 ;
  assign n29506 = n29505 ^ n20839 ^ 1'b0 ;
  assign n29507 = n6333 ^ n2933 ^ 1'b0 ;
  assign n29508 = n6737 | n10965 ;
  assign n29509 = n13327 & ~n29508 ;
  assign n29510 = n29509 ^ n10386 ^ 1'b0 ;
  assign n29511 = n10197 ^ n2358 ^ 1'b0 ;
  assign n29512 = n12185 | n29511 ;
  assign n29513 = ~n2812 & n14218 ;
  assign n29514 = ~n9680 & n23872 ;
  assign n29515 = ~n1023 & n1492 ;
  assign n29516 = n6514 | n29515 ;
  assign n29517 = n29516 ^ n1091 ^ 1'b0 ;
  assign n29518 = n384 & n5825 ;
  assign n29519 = n1286 & n14535 ;
  assign n29520 = n29018 & n29519 ;
  assign n29521 = n2431 & ~n10510 ;
  assign n29522 = n5419 & n29521 ;
  assign n29523 = ~n767 & n3648 ;
  assign n29524 = ~n743 & n29523 ;
  assign n29525 = n5428 & ~n8317 ;
  assign n29526 = ~n1608 & n18919 ;
  assign n29527 = n1541 | n18121 ;
  assign n29528 = n17187 & ~n29527 ;
  assign n29529 = ~n1349 & n10942 ;
  assign n29530 = n29429 & n29529 ;
  assign n29531 = n12723 ^ n2494 ^ 1'b0 ;
  assign n29532 = n6889 & ~n29531 ;
  assign n29533 = n18181 & ~n22872 ;
  assign n29534 = n792 | n16099 ;
  assign n29535 = n29534 ^ n17347 ^ 1'b0 ;
  assign n29536 = n10002 ^ n1081 ^ 1'b0 ;
  assign n29537 = n9142 ^ n5913 ^ 1'b0 ;
  assign n29538 = n26571 ^ n5923 ^ 1'b0 ;
  assign n29539 = n13917 | n29538 ;
  assign n29540 = n10539 ^ n5820 ^ 1'b0 ;
  assign n29541 = x3 | n29540 ;
  assign n29542 = n29541 ^ n6055 ^ 1'b0 ;
  assign n29543 = ~n4770 & n29542 ;
  assign n29544 = n2577 | n6084 ;
  assign n29545 = n23684 ^ n5445 ^ n3512 ;
  assign n29546 = n2354 & ~n20480 ;
  assign n29547 = n12309 ^ n2130 ^ 1'b0 ;
  assign n29548 = n1904 & n29547 ;
  assign n29549 = n29548 ^ n11506 ^ 1'b0 ;
  assign n29550 = n12084 | n29549 ;
  assign n29551 = n3707 & ~n29550 ;
  assign n29552 = n29551 ^ n484 ^ 1'b0 ;
  assign n29553 = n4586 | n8549 ;
  assign n29554 = n16445 & n29553 ;
  assign n29556 = ~n2888 & n9764 ;
  assign n29557 = n16090 & ~n29556 ;
  assign n29555 = n3969 & n6085 ;
  assign n29558 = n29557 ^ n29555 ^ 1'b0 ;
  assign n29559 = ~n1508 & n5398 ;
  assign n29560 = n29559 ^ n8392 ^ 1'b0 ;
  assign n29564 = ~n142 & n2514 ;
  assign n29565 = ( n8865 & n12870 ) | ( n8865 & n29564 ) | ( n12870 & n29564 ) ;
  assign n29566 = n11922 & n29565 ;
  assign n29561 = n336 | n8013 ;
  assign n29562 = n29561 ^ n9975 ^ 1'b0 ;
  assign n29563 = n29562 ^ n3636 ^ 1'b0 ;
  assign n29567 = n29566 ^ n29563 ^ 1'b0 ;
  assign n29568 = ~n37 & n1048 ;
  assign n29569 = n29568 ^ n8822 ^ 1'b0 ;
  assign n29570 = n22375 | n22863 ;
  assign n29571 = n26593 & ~n29570 ;
  assign n29572 = ~n29569 & n29571 ;
  assign n29573 = n2773 & n4992 ;
  assign n29574 = n258 & ~n11897 ;
  assign n29575 = n29573 & n29574 ;
  assign n29576 = n27080 ^ n1956 ^ 1'b0 ;
  assign n29577 = n6889 & n27670 ;
  assign n29578 = n29577 ^ n11076 ^ 1'b0 ;
  assign n29579 = n13027 ^ n1373 ^ 1'b0 ;
  assign n29581 = n3769 ^ n2268 ^ 1'b0 ;
  assign n29582 = n14089 | n29581 ;
  assign n29580 = n3514 ^ n448 ^ 1'b0 ;
  assign n29583 = n29582 ^ n29580 ^ 1'b0 ;
  assign n29584 = n11474 & n29583 ;
  assign n29585 = n24667 ^ n3484 ^ 1'b0 ;
  assign n29586 = n29585 ^ n22089 ^ 1'b0 ;
  assign n29587 = n29584 & n29586 ;
  assign n29588 = ~n25513 & n29587 ;
  assign n29589 = n29588 ^ n28335 ^ 1'b0 ;
  assign n29590 = n18280 ^ n4312 ^ 1'b0 ;
  assign n29591 = ( n9635 & ~n21389 ) | ( n9635 & n26103 ) | ( ~n21389 & n26103 ) ;
  assign n29592 = ~n200 & n6174 ;
  assign n29593 = n16391 & n29592 ;
  assign n29594 = n17341 ^ x0 ^ 1'b0 ;
  assign n29595 = n1183 | n29594 ;
  assign n29596 = n12798 ^ n7179 ^ 1'b0 ;
  assign n29597 = n29596 ^ n27075 ^ 1'b0 ;
  assign n29598 = n4029 | n24454 ;
  assign n29599 = n22616 | n29598 ;
  assign n29600 = n21880 ^ n507 ^ 1'b0 ;
  assign n29601 = n11513 & n18207 ;
  assign n29602 = n29601 ^ n215 ^ 1'b0 ;
  assign n29603 = n10928 & n13694 ;
  assign n29604 = n6385 & ~n21343 ;
  assign n29605 = ~n23862 & n29604 ;
  assign n29606 = n22872 | n29605 ;
  assign n29607 = n21355 | n29606 ;
  assign n29608 = n12463 ^ n6341 ^ n233 ;
  assign n29609 = n6502 ^ n4482 ^ 1'b0 ;
  assign n29610 = n27299 ^ n20788 ^ 1'b0 ;
  assign n29611 = n24784 | n29610 ;
  assign n29612 = n10527 ^ n322 ^ 1'b0 ;
  assign n29613 = n20039 ^ n9210 ^ n6280 ;
  assign n29615 = n10919 & ~n16143 ;
  assign n29616 = ~n817 & n29615 ;
  assign n29614 = n7802 & n24818 ;
  assign n29617 = n29616 ^ n29614 ^ 1'b0 ;
  assign n29618 = n21823 ^ n10072 ^ 1'b0 ;
  assign n29619 = n323 & ~n1326 ;
  assign n29620 = n29618 | n29619 ;
  assign n29621 = n12995 ^ n4965 ^ 1'b0 ;
  assign n29622 = n19316 ^ n18107 ^ 1'b0 ;
  assign n29623 = n29583 ^ n46 ^ 1'b0 ;
  assign n29624 = n13396 | n29623 ;
  assign n29625 = n4626 & ~n15782 ;
  assign n29626 = ~n20748 & n29625 ;
  assign n29627 = n22747 ^ n1588 ^ 1'b0 ;
  assign n29628 = n24606 & n29627 ;
  assign n29629 = n11309 & n29628 ;
  assign n29630 = n439 | n16749 ;
  assign n29631 = n29630 ^ n16284 ^ 1'b0 ;
  assign n29632 = n9721 ^ n9357 ^ 1'b0 ;
  assign n29633 = n22735 ^ n1255 ^ 1'b0 ;
  assign n29634 = n6492 ^ n726 ^ 1'b0 ;
  assign n29635 = n17707 & n29634 ;
  assign n29637 = n1724 | n5256 ;
  assign n29638 = n16178 | n29637 ;
  assign n29639 = n29638 ^ n2883 ^ 1'b0 ;
  assign n29636 = n17086 | n22966 ;
  assign n29640 = n29639 ^ n29636 ^ 1'b0 ;
  assign n29641 = n26249 ^ n19490 ^ 1'b0 ;
  assign n29642 = n29640 & ~n29641 ;
  assign n29643 = n37 & n29080 ;
  assign n29644 = n979 | n2514 ;
  assign n29645 = n29644 ^ n2532 ^ 1'b0 ;
  assign n29647 = n3637 & ~n12527 ;
  assign n29648 = n7657 | n29647 ;
  assign n29646 = n1034 & ~n7605 ;
  assign n29649 = n29648 ^ n29646 ^ 1'b0 ;
  assign n29650 = n20244 ^ n3586 ^ 1'b0 ;
  assign n29651 = n663 | n13169 ;
  assign n29652 = n29651 ^ n10476 ^ 1'b0 ;
  assign n29653 = n5410 & ~n29652 ;
  assign n29654 = n6780 & ~n29653 ;
  assign n29655 = n29654 ^ n28098 ^ 1'b0 ;
  assign n29656 = n4053 & n4836 ;
  assign n29657 = ~n27870 & n29656 ;
  assign n29659 = n6552 & n12642 ;
  assign n29660 = n13049 ^ n9952 ^ n3049 ;
  assign n29661 = ~n29659 & n29660 ;
  assign n29658 = n2800 & n3882 ;
  assign n29662 = n29661 ^ n29658 ^ 1'b0 ;
  assign n29663 = n29569 ^ n23246 ^ n18099 ;
  assign n29664 = n2313 & n19653 ;
  assign n29665 = n3624 & n10810 ;
  assign n29666 = n10213 ^ n7144 ^ 1'b0 ;
  assign n29667 = ~n26460 & n29666 ;
  assign n29668 = n24516 ^ n17851 ^ 1'b0 ;
  assign n29669 = ~n16954 & n21597 ;
  assign n29670 = ~n653 & n29669 ;
  assign n29671 = ~n3972 & n23083 ;
  assign n29672 = n1480 & n8939 ;
  assign n29673 = n5905 | n22689 ;
  assign n29674 = n9227 & ~n9360 ;
  assign n29675 = n18874 ^ n14544 ^ 1'b0 ;
  assign n29676 = n726 & ~n29675 ;
  assign n29677 = ~n6906 & n29676 ;
  assign n29678 = n29677 ^ n4748 ^ 1'b0 ;
  assign n29679 = n24361 & n28352 ;
  assign n29680 = n5229 & ~n21055 ;
  assign n29681 = ~n18106 & n29680 ;
  assign n29682 = n1115 | n21136 ;
  assign n29683 = n29682 ^ n3411 ^ 1'b0 ;
  assign n29684 = n1662 & ~n29683 ;
  assign n29685 = ~n8472 & n11069 ;
  assign n29686 = n6045 & n29685 ;
  assign n29687 = ~n29684 & n29686 ;
  assign n29688 = n5227 | n29687 ;
  assign n29689 = n457 & ~n5295 ;
  assign n29690 = n5621 | n8326 ;
  assign n29691 = n20848 | n27466 ;
  assign n29692 = n29691 ^ n28818 ^ 1'b0 ;
  assign n29693 = n5169 & ~n7288 ;
  assign n29697 = n3068 | n4322 ;
  assign n29694 = n13732 ^ n8064 ^ 1'b0 ;
  assign n29695 = n29694 ^ n310 ^ 1'b0 ;
  assign n29696 = ~n17436 & n29695 ;
  assign n29698 = n29697 ^ n29696 ^ 1'b0 ;
  assign n29699 = n22737 ^ n3965 ^ 1'b0 ;
  assign n29700 = ( ~n7789 & n19690 ) | ( ~n7789 & n22501 ) | ( n19690 & n22501 ) ;
  assign n29701 = n2872 & ~n9424 ;
  assign n29702 = n29701 ^ n8523 ^ 1'b0 ;
  assign n29703 = n9009 ^ n7805 ^ 1'b0 ;
  assign n29704 = n28725 ^ n15981 ^ 1'b0 ;
  assign n29705 = ~n29703 & n29704 ;
  assign n29706 = ~n687 & n23655 ;
  assign n29707 = n29706 ^ n15334 ^ 1'b0 ;
  assign n29708 = n6711 & ~n9267 ;
  assign n29709 = n29708 ^ n10132 ^ 1'b0 ;
  assign n29710 = n17464 & ~n29709 ;
  assign n29711 = n21106 ^ n11730 ^ n8543 ;
  assign n29712 = n29711 ^ n7265 ^ n2196 ;
  assign n29713 = n13425 ^ n3050 ^ 1'b0 ;
  assign n29714 = n880 | n29713 ;
  assign n29715 = n104 & ~n1361 ;
  assign n29716 = n4290 | n7350 ;
  assign n29717 = n13205 | n29716 ;
  assign n29718 = n20647 ^ n1178 ^ 1'b0 ;
  assign n29719 = n29717 & ~n29718 ;
  assign n29720 = ~n2462 & n29719 ;
  assign n29721 = n29720 ^ n12997 ^ 1'b0 ;
  assign n29722 = n7011 & n14181 ;
  assign n29723 = n26069 | n29722 ;
  assign n29724 = n276 & ~n8282 ;
  assign n29725 = n11241 | n12443 ;
  assign n29726 = n29725 ^ n5928 ^ 1'b0 ;
  assign n29727 = n5308 & n11057 ;
  assign n29728 = n6315 & n29727 ;
  assign n29729 = n29728 ^ n8192 ^ 1'b0 ;
  assign n29730 = n461 | n29729 ;
  assign n29731 = n29726 | n29730 ;
  assign n29738 = ~n2942 & n7104 ;
  assign n29732 = n14840 ^ n3083 ^ 1'b0 ;
  assign n29733 = n15711 | n29732 ;
  assign n29734 = n3244 & ~n24262 ;
  assign n29735 = n24262 & n29734 ;
  assign n29736 = n29735 ^ n25057 ^ 1'b0 ;
  assign n29737 = ~n29733 & n29736 ;
  assign n29739 = n29738 ^ n29737 ^ n2624 ;
  assign n29740 = n24281 ^ n12039 ^ 1'b0 ;
  assign n29741 = n29740 ^ n1225 ^ 1'b0 ;
  assign n29742 = n22549 ^ n2878 ^ 1'b0 ;
  assign n29743 = n29742 ^ n19668 ^ 1'b0 ;
  assign n29744 = n25010 & n29743 ;
  assign n29745 = n1530 & n15012 ;
  assign n29746 = n29745 ^ n6885 ^ 1'b0 ;
  assign n29747 = n29746 ^ n15916 ^ 1'b0 ;
  assign n29748 = n1865 | n6703 ;
  assign n29749 = n12982 | n29541 ;
  assign n29750 = n29749 ^ n8489 ^ 1'b0 ;
  assign n29751 = n5018 & n29750 ;
  assign n29752 = ~n2567 & n3361 ;
  assign n29753 = ( n2235 & n17882 ) | ( n2235 & n29752 ) | ( n17882 & n29752 ) ;
  assign n29755 = n13876 ^ n5310 ^ 1'b0 ;
  assign n29754 = n3804 & ~n13301 ;
  assign n29756 = n29755 ^ n29754 ^ 1'b0 ;
  assign n29757 = n1263 & ~n1608 ;
  assign n29758 = n21742 ^ n11025 ^ 1'b0 ;
  assign n29759 = n29757 & n29758 ;
  assign n29760 = n27995 ^ n14647 ^ 1'b0 ;
  assign n29761 = n4254 ^ n1654 ^ 1'b0 ;
  assign n29762 = n13098 & n29761 ;
  assign n29763 = n10366 & ~n29762 ;
  assign n29764 = ~n1274 & n17674 ;
  assign n29766 = n2263 ^ n553 ^ 1'b0 ;
  assign n29767 = n29766 ^ n1986 ^ 1'b0 ;
  assign n29765 = ~n6141 & n10621 ;
  assign n29768 = n29767 ^ n29765 ^ 1'b0 ;
  assign n29769 = n290 & n1412 ;
  assign n29770 = ~n4485 & n29769 ;
  assign n29771 = ( ~n8883 & n18110 ) | ( ~n8883 & n29770 ) | ( n18110 & n29770 ) ;
  assign n29772 = n29771 ^ n15783 ^ 1'b0 ;
  assign n29773 = n1286 | n12049 ;
  assign n29774 = n2007 & ~n29773 ;
  assign n29775 = ~n26332 & n29774 ;
  assign n29776 = n29775 ^ n16604 ^ 1'b0 ;
  assign n29777 = ~n8198 & n26566 ;
  assign n29778 = n9675 | n18196 ;
  assign n29779 = n28230 ^ n4179 ^ 1'b0 ;
  assign n29780 = ~n4139 & n29779 ;
  assign n29781 = ~n19591 & n29780 ;
  assign n29782 = n29781 ^ n21539 ^ 1'b0 ;
  assign n29783 = ~n3355 & n9739 ;
  assign n29784 = n2920 & ~n23519 ;
  assign n29785 = n29784 ^ n6981 ^ 1'b0 ;
  assign n29786 = n3947 & ~n29785 ;
  assign n29787 = n17770 & ~n24262 ;
  assign n29788 = n29787 ^ n15561 ^ 1'b0 ;
  assign n29789 = n4349 ^ n1619 ^ 1'b0 ;
  assign n29790 = ~n9647 & n29789 ;
  assign n29791 = n15012 ^ n510 ^ 1'b0 ;
  assign n29792 = n1649 & ~n6170 ;
  assign n29793 = n6170 & n29792 ;
  assign n29794 = n29793 ^ n4088 ^ 1'b0 ;
  assign n29795 = ~n26825 & n29794 ;
  assign n29796 = n2410 & ~n7933 ;
  assign n29797 = n3178 & n6099 ;
  assign n29798 = n2792 | n29797 ;
  assign n29799 = n2156 & n17451 ;
  assign n29800 = n1920 | n29799 ;
  assign n29801 = n10632 & n29800 ;
  assign n29802 = ~n29798 & n29801 ;
  assign n29803 = n3580 & ~n10201 ;
  assign n29804 = n29803 ^ n1562 ^ 1'b0 ;
  assign n29805 = ~n3878 & n13612 ;
  assign n29806 = ( n3186 & ~n14821 ) | ( n3186 & n22610 ) | ( ~n14821 & n22610 ) ;
  assign n29807 = n10976 | n22940 ;
  assign n29808 = n7805 & ~n29807 ;
  assign n29809 = n8059 | n21043 ;
  assign n29810 = n7594 | n29809 ;
  assign n29811 = n614 ^ n322 ^ 1'b0 ;
  assign n29812 = ( ~n7454 & n12052 ) | ( ~n7454 & n29811 ) | ( n12052 & n29811 ) ;
  assign n29813 = n3001 ^ n390 ^ 1'b0 ;
  assign n29814 = n15618 & n29813 ;
  assign n29815 = ~n2689 & n29814 ;
  assign n29816 = n29812 | n29815 ;
  assign n29817 = n12472 | n27971 ;
  assign n29818 = n29816 | n29817 ;
  assign n29819 = n20269 ^ n1926 ^ 1'b0 ;
  assign n29820 = n47 & n8283 ;
  assign n29821 = ~n239 & n25450 ;
  assign n29822 = ~n912 & n4560 ;
  assign n29823 = ~n11861 & n29822 ;
  assign n29824 = n5208 & n5963 ;
  assign n29825 = n29824 ^ n4404 ^ 1'b0 ;
  assign n29826 = n4774 & ~n29825 ;
  assign n29827 = n29823 & n29826 ;
  assign n29828 = n8282 ^ n6607 ^ 1'b0 ;
  assign n29829 = n28587 ^ n6378 ^ 1'b0 ;
  assign n29830 = n28866 ^ n5950 ^ 1'b0 ;
  assign n29831 = n8851 ^ n2352 ^ 1'b0 ;
  assign n29832 = ~n3648 & n10285 ;
  assign n29833 = n6923 ^ n3209 ^ 1'b0 ;
  assign n29834 = ~n2896 & n4185 ;
  assign n29835 = ~n1940 & n29834 ;
  assign n29836 = ( n4400 & n15595 ) | ( n4400 & ~n29835 ) | ( n15595 & ~n29835 ) ;
  assign n29837 = ~n23525 & n29836 ;
  assign n29838 = n23525 & n29837 ;
  assign n29839 = ( n300 & ~n2784 ) | ( n300 & n24343 ) | ( ~n2784 & n24343 ) ;
  assign n29840 = n26866 & ~n29839 ;
  assign n29841 = n17323 ^ n6620 ^ 1'b0 ;
  assign n29842 = n16691 ^ n12721 ^ 1'b0 ;
  assign n29843 = n3032 | n29842 ;
  assign n29844 = n16634 & ~n29843 ;
  assign n29845 = n20597 ^ n14986 ^ 1'b0 ;
  assign n29846 = n12649 ^ n10025 ^ 1'b0 ;
  assign n29847 = ~n185 & n4934 ;
  assign n29848 = ~n2399 & n5076 ;
  assign n29849 = n3866 | n8711 ;
  assign n29850 = ( ~n72 & n1825 ) | ( ~n72 & n29849 ) | ( n1825 & n29849 ) ;
  assign n29851 = n17831 ^ n11975 ^ 1'b0 ;
  assign n29852 = n119 | n29851 ;
  assign n29853 = n13800 & ~n29852 ;
  assign n29854 = n404 | n19725 ;
  assign n29855 = n3104 & ~n29854 ;
  assign n29856 = n29855 ^ n15742 ^ 1'b0 ;
  assign n29857 = n28134 ^ n9516 ^ 1'b0 ;
  assign n29858 = n29856 & n29857 ;
  assign n29859 = n506 & n2574 ;
  assign n29860 = n29859 ^ n2736 ^ 1'b0 ;
  assign n29861 = n14462 | n29860 ;
  assign n29862 = n29861 ^ n6512 ^ 1'b0 ;
  assign n29863 = n863 & n29862 ;
  assign n29864 = n784 & n29863 ;
  assign n29865 = n29864 ^ n25129 ^ 1'b0 ;
  assign n29866 = n20888 ^ n3078 ^ 1'b0 ;
  assign n29867 = n29865 & n29866 ;
  assign n29868 = n26128 & n29867 ;
  assign n29869 = ~n2075 & n8637 ;
  assign n29870 = n29869 ^ n6713 ^ 1'b0 ;
  assign n29871 = n7488 | n29870 ;
  assign n29872 = n29871 ^ n114 ^ 1'b0 ;
  assign n29873 = n29872 ^ n12170 ^ 1'b0 ;
  assign n29874 = n11542 & ~n18654 ;
  assign n29875 = n29874 ^ n2945 ^ 1'b0 ;
  assign n29876 = n1396 | n3988 ;
  assign n29877 = n22332 | n29876 ;
  assign n29878 = n12740 ^ n3176 ^ 1'b0 ;
  assign n29879 = n7520 | n28781 ;
  assign n29880 = n29878 & ~n29879 ;
  assign n29881 = n8019 | n16981 ;
  assign n29882 = n2674 | n29881 ;
  assign n29883 = n29882 ^ n21101 ^ 1'b0 ;
  assign n29884 = ~n8402 & n28253 ;
  assign n29885 = n14665 & n29884 ;
  assign n29886 = n14204 | n16203 ;
  assign n29887 = n29886 ^ n10167 ^ 1'b0 ;
  assign n29888 = ~n17750 & n18026 ;
  assign n29889 = n44 & n123 ;
  assign n29890 = ~n123 & n29889 ;
  assign n29891 = ~n227 & n29890 ;
  assign n29892 = ~n1499 & n29891 ;
  assign n29893 = ~n442 & n29892 ;
  assign n29894 = ~n4091 & n29893 ;
  assign n29895 = n9930 | n29894 ;
  assign n29896 = n29894 & ~n29895 ;
  assign n29897 = n22789 | n29896 ;
  assign n29898 = n22096 & ~n29897 ;
  assign n29899 = n3335 & ~n6436 ;
  assign n29900 = n23486 | n29899 ;
  assign n29901 = n29900 ^ n15579 ^ 1'b0 ;
  assign n29902 = n10252 & n28146 ;
  assign n29903 = n161 & ~n16518 ;
  assign n29904 = n2566 ^ n1872 ^ 1'b0 ;
  assign n29905 = ~n2107 & n29904 ;
  assign n29906 = n2982 & n29905 ;
  assign n29907 = n29906 ^ n25346 ^ 1'b0 ;
  assign n29908 = n10282 ^ n4344 ^ 1'b0 ;
  assign n29909 = n13768 | n29908 ;
  assign n29910 = n7915 & n14714 ;
  assign n29911 = n29910 ^ n28650 ^ 1'b0 ;
  assign n29912 = n14689 & ~n28804 ;
  assign n29913 = ~n21411 & n29912 ;
  assign n29914 = n15312 ^ n5797 ^ 1'b0 ;
  assign n29915 = n24820 ^ n475 ^ 1'b0 ;
  assign n29916 = n20566 & n29915 ;
  assign n29917 = n18451 ^ n1431 ^ 1'b0 ;
  assign n29918 = ~n5952 & n29917 ;
  assign n29919 = n10078 & ~n21938 ;
  assign n29920 = n5616 & ~n15325 ;
  assign n29921 = n29920 ^ n12962 ^ 1'b0 ;
  assign n29922 = ~n1217 & n27831 ;
  assign n29923 = n29922 ^ n5201 ^ 1'b0 ;
  assign n29924 = n19300 | n21868 ;
  assign n29925 = ~n19466 & n29924 ;
  assign n29926 = n10644 & n19743 ;
  assign n29927 = n9892 & ~n29926 ;
  assign n29928 = n24906 ^ n14190 ^ 1'b0 ;
  assign n29929 = n10635 & ~n15785 ;
  assign n29930 = ~n16209 & n22898 ;
  assign n29931 = ~n7430 & n7508 ;
  assign n29932 = n13087 & n29931 ;
  assign n29933 = n10992 | n15591 ;
  assign n29934 = n11085 ^ n715 ^ 1'b0 ;
  assign n29935 = ~n16189 & n29934 ;
  assign n29936 = ~n2914 & n8825 ;
  assign n29937 = n13326 & n29936 ;
  assign n29938 = n2571 & ~n12683 ;
  assign n29939 = n29938 ^ n7323 ^ 1'b0 ;
  assign n29940 = ~n818 & n1713 ;
  assign n29941 = n29940 ^ n13574 ^ 1'b0 ;
  assign n29942 = n10741 & ~n29941 ;
  assign n29945 = n15544 | n17483 ;
  assign n29943 = n365 & ~n4856 ;
  assign n29944 = n11640 & n29943 ;
  assign n29946 = n29945 ^ n29944 ^ 1'b0 ;
  assign n29947 = n15799 & ~n19870 ;
  assign n29948 = n29946 & n29947 ;
  assign n29949 = n14272 | n26956 ;
  assign n29950 = n8234 ^ n227 ^ 1'b0 ;
  assign n29951 = n1095 & ~n29950 ;
  assign n29952 = n4297 ^ n273 ^ 1'b0 ;
  assign n29953 = n25326 & ~n29952 ;
  assign n29954 = n29953 ^ n10965 ^ 1'b0 ;
  assign n29955 = n5835 | n29954 ;
  assign n29956 = n14678 ^ n1987 ^ 1'b0 ;
  assign n29957 = n22504 & n24852 ;
  assign n29958 = ~n3567 & n8396 ;
  assign n29959 = n22768 & n29958 ;
  assign n29960 = n2618 | n5583 ;
  assign n29961 = n4256 & ~n29960 ;
  assign n29962 = n1024 & ~n26435 ;
  assign n29963 = ~n27844 & n29962 ;
  assign n29964 = n29963 ^ n12438 ^ 1'b0 ;
  assign n29965 = ~n18440 & n29964 ;
  assign n29966 = n15468 ^ n1505 ^ 1'b0 ;
  assign n29967 = n12991 | n29966 ;
  assign n29968 = ~n55 & n20890 ;
  assign n29969 = ~n5347 & n29968 ;
  assign n29970 = ~n23894 & n29969 ;
  assign n29971 = n3033 & n29970 ;
  assign n29973 = n16534 ^ n5049 ^ 1'b0 ;
  assign n29972 = n415 & ~n1758 ;
  assign n29974 = n29973 ^ n29972 ^ 1'b0 ;
  assign n29975 = n6107 | n29974 ;
  assign n29976 = n5447 & ~n26609 ;
  assign n29977 = n75 & ~n528 ;
  assign n29978 = n7969 & n7999 ;
  assign n29979 = ~n16800 & n29978 ;
  assign n29980 = n3283 & n4334 ;
  assign n29981 = n27302 ^ n4549 ^ 1'b0 ;
  assign n29982 = n8552 ^ n5551 ^ 1'b0 ;
  assign n29983 = n29296 ^ n3598 ^ 1'b0 ;
  assign n29984 = n22739 ^ n3202 ^ 1'b0 ;
  assign n29985 = n2001 & n29984 ;
  assign n29986 = n6649 & ~n29985 ;
  assign n29987 = n13865 ^ n8084 ^ 1'b0 ;
  assign n29988 = n4654 & ~n29987 ;
  assign n29989 = ~n24147 & n29988 ;
  assign n29990 = n3369 ^ n2500 ^ 1'b0 ;
  assign n29991 = n2888 | n29990 ;
  assign n29992 = n8915 ^ n743 ^ 1'b0 ;
  assign n29993 = n15225 & n29992 ;
  assign n29994 = n24349 & n29993 ;
  assign n29995 = n25764 & ~n29994 ;
  assign n29996 = n5711 ^ n954 ^ 1'b0 ;
  assign n29997 = n23299 & ~n29996 ;
  assign n29998 = n8323 ^ n7459 ^ 1'b0 ;
  assign n29999 = n22399 & ~n29998 ;
  assign n30000 = n23772 ^ n7590 ^ 1'b0 ;
  assign n30001 = n5128 | n27351 ;
  assign n30002 = n23759 ^ n3692 ^ 1'b0 ;
  assign n30003 = n15367 & ~n30002 ;
  assign n30004 = n30003 ^ n14689 ^ 1'b0 ;
  assign n30005 = n3743 | n23581 ;
  assign n30006 = n7742 | n11546 ;
  assign n30007 = n30005 & ~n30006 ;
  assign n30008 = n3423 & ~n28760 ;
  assign n30009 = n30008 ^ n3664 ^ 1'b0 ;
  assign n30010 = n7667 & n13603 ;
  assign n30011 = n30010 ^ n1940 ^ 1'b0 ;
  assign n30012 = n30011 ^ n6553 ^ 1'b0 ;
  assign n30013 = ~n10902 & n30012 ;
  assign n30014 = n6258 | n17815 ;
  assign n30015 = n11395 ^ n5801 ^ n3816 ;
  assign n30016 = n7508 & ~n30015 ;
  assign n30017 = n27366 ^ n13852 ^ 1'b0 ;
  assign n30018 = n30016 & ~n30017 ;
  assign n30019 = n2129 & n17678 ;
  assign n30020 = n27917 & n30019 ;
  assign n30021 = n5183 & n7859 ;
  assign n30022 = ~n12298 & n30021 ;
  assign n30023 = n3939 & ~n5241 ;
  assign n30024 = n7786 | n17337 ;
  assign n30025 = n3567 & ~n30024 ;
  assign n30026 = n210 | n30025 ;
  assign n30027 = n1165 | n30026 ;
  assign n30028 = n1213 | n6365 ;
  assign n30029 = n888 | n1219 ;
  assign n30030 = n888 & ~n30029 ;
  assign n30031 = ~n567 & n30030 ;
  assign n30032 = ~n917 & n955 ;
  assign n30033 = n917 & n30032 ;
  assign n30034 = ~n2201 & n30033 ;
  assign n30035 = ~n4311 & n30034 ;
  assign n30036 = n30031 & n30035 ;
  assign n30037 = n5865 & ~n14877 ;
  assign n30038 = ( n2531 & n30036 ) | ( n2531 & ~n30037 ) | ( n30036 & ~n30037 ) ;
  assign n30039 = n2538 & ~n30038 ;
  assign n30040 = n2291 & ~n30039 ;
  assign n30041 = n30028 & n30040 ;
  assign n30042 = ~n614 & n1748 ;
  assign n30043 = n8756 | n10861 ;
  assign n30044 = n6543 & n16373 ;
  assign n30045 = n614 & n30044 ;
  assign n30048 = ~n2311 & n15225 ;
  assign n30046 = n810 & n1394 ;
  assign n30047 = ~n2495 & n30046 ;
  assign n30049 = n30048 ^ n30047 ^ 1'b0 ;
  assign n30050 = n9326 | n16703 ;
  assign n30051 = n30050 ^ n689 ^ 1'b0 ;
  assign n30052 = n7497 & ~n22371 ;
  assign n30053 = n26203 ^ n17328 ^ 1'b0 ;
  assign n30054 = n16656 & n30053 ;
  assign n30055 = n327 & n2260 ;
  assign n30056 = n10391 ^ n499 ^ 1'b0 ;
  assign n30057 = x0 & n30056 ;
  assign n30058 = n7495 & n27151 ;
  assign n30059 = n5646 ^ n300 ^ 1'b0 ;
  assign n30060 = n30059 ^ n5273 ^ 1'b0 ;
  assign n30061 = n30060 ^ n6940 ^ 1'b0 ;
  assign n30062 = ( n2959 & n5637 ) | ( n2959 & n30061 ) | ( n5637 & n30061 ) ;
  assign n30063 = n30058 | n30062 ;
  assign n30064 = n21539 ^ n4954 ^ 1'b0 ;
  assign n30065 = n7596 & ~n30064 ;
  assign n30066 = ~n5701 & n29653 ;
  assign n30067 = n23072 ^ n4399 ^ 1'b0 ;
  assign n30068 = n9188 ^ n284 ^ 1'b0 ;
  assign n30069 = n24041 & n30068 ;
  assign n30070 = n30069 ^ n5043 ^ 1'b0 ;
  assign n30071 = n3887 & n30070 ;
  assign n30072 = n7057 | n7736 ;
  assign n30073 = n30072 ^ n15512 ^ 1'b0 ;
  assign n30074 = ~n7217 & n16556 ;
  assign n30075 = n18308 ^ n16303 ^ 1'b0 ;
  assign n30076 = n24598 ^ n13322 ^ n6578 ;
  assign n30083 = n17927 ^ n1165 ^ 1'b0 ;
  assign n30084 = n26772 | n30083 ;
  assign n30085 = n30084 ^ n1979 ^ 1'b0 ;
  assign n30078 = n9452 & n10582 ;
  assign n30079 = n8195 & ~n30078 ;
  assign n30080 = n18530 & n30079 ;
  assign n30077 = n229 & n1254 ;
  assign n30081 = n30080 ^ n30077 ^ n5845 ;
  assign n30082 = n7239 & ~n30081 ;
  assign n30086 = n30085 ^ n30082 ^ 1'b0 ;
  assign n30087 = n6762 & ~n9523 ;
  assign n30088 = ~n10134 & n30087 ;
  assign n30089 = n30088 ^ n27426 ^ 1'b0 ;
  assign n30090 = n9641 ^ n7706 ^ 1'b0 ;
  assign n30091 = n23981 ^ n5825 ^ 1'b0 ;
  assign n30092 = ~n27502 & n30091 ;
  assign n30093 = n3632 ^ n351 ^ 1'b0 ;
  assign n30094 = n2289 & ~n30093 ;
  assign n30095 = n30094 ^ n5726 ^ 1'b0 ;
  assign n30096 = n3271 ^ n2973 ^ 1'b0 ;
  assign n30097 = n30096 ^ n13172 ^ 1'b0 ;
  assign n30098 = ~n16329 & n30097 ;
  assign n30099 = n19735 | n30098 ;
  assign n30100 = n229 | n1102 ;
  assign n30101 = n30100 ^ n12963 ^ 1'b0 ;
  assign n30102 = n4485 & ~n30101 ;
  assign n30103 = ~n246 & n13949 ;
  assign n30104 = n6816 & n30103 ;
  assign n30105 = n6620 & n30104 ;
  assign n30106 = ~n20638 & n30105 ;
  assign n30107 = n30106 ^ n10831 ^ 1'b0 ;
  assign n30108 = n3892 | n25169 ;
  assign n30109 = n4157 | n5118 ;
  assign n30110 = n30109 ^ n30 ^ 1'b0 ;
  assign n30111 = n287 & n1685 ;
  assign n30112 = ~n4793 & n30111 ;
  assign n30113 = n30112 ^ n6610 ^ 1'b0 ;
  assign n30115 = ~n10687 & n11042 ;
  assign n30116 = n30115 ^ n9461 ^ 1'b0 ;
  assign n30114 = n1785 | n24010 ;
  assign n30117 = n30116 ^ n30114 ^ 1'b0 ;
  assign n30118 = n1739 & ~n16072 ;
  assign n30119 = n24553 ^ n16738 ^ 1'b0 ;
  assign n30120 = n1066 & n1384 ;
  assign n30121 = ( n47 & ~n24955 ) | ( n47 & n30120 ) | ( ~n24955 & n30120 ) ;
  assign n30122 = n11302 ^ n6048 ^ 1'b0 ;
  assign n30123 = n26763 & ~n30122 ;
  assign n30124 = n20662 ^ n4569 ^ 1'b0 ;
  assign n30125 = n30123 & ~n30124 ;
  assign n30126 = n19349 & n25217 ;
  assign n30127 = n20459 & n30126 ;
  assign n30128 = n4840 & ~n22615 ;
  assign n30129 = ~n4403 & n30128 ;
  assign n30130 = n2767 & n5623 ;
  assign n30131 = n6109 ^ n670 ^ 1'b0 ;
  assign n30132 = n4927 | n5778 ;
  assign n30133 = n6442 & ~n30132 ;
  assign n30134 = n1471 | n30133 ;
  assign n30135 = n6476 | n14252 ;
  assign n30136 = n3624 | n3951 ;
  assign n30137 = n9574 & ~n30136 ;
  assign n30138 = n337 | n30137 ;
  assign n30139 = n25030 | n30138 ;
  assign n30140 = ~n21630 & n28821 ;
  assign n30141 = n257 & ~n26525 ;
  assign n30142 = n1054 & n30141 ;
  assign n30143 = n195 & ~n21741 ;
  assign n30144 = n14771 & n30143 ;
  assign n30145 = n1431 & n13908 ;
  assign n30146 = n4312 & n30145 ;
  assign n30147 = n30146 ^ n268 ^ 1'b0 ;
  assign n30148 = n703 & ~n30147 ;
  assign n30149 = n18453 & n30148 ;
  assign n30150 = n30149 ^ n10900 ^ 1'b0 ;
  assign n30151 = n26373 ^ n19876 ^ 1'b0 ;
  assign n30152 = n11074 & n30151 ;
  assign n30153 = n10429 ^ n1501 ^ 1'b0 ;
  assign n30154 = n3797 & n30153 ;
  assign n30155 = n15148 & n16425 ;
  assign n30156 = n84 & ~n30155 ;
  assign n30157 = n896 & n30156 ;
  assign n30158 = ~n114 & n30157 ;
  assign n30159 = n4105 ^ n1668 ^ 1'b0 ;
  assign n30160 = n11083 ^ n8967 ^ 1'b0 ;
  assign n30161 = n9210 & n30160 ;
  assign n30162 = ~n468 & n30161 ;
  assign n30163 = n7358 | n19561 ;
  assign n30164 = n11253 | n21464 ;
  assign n30165 = n30163 | n30164 ;
  assign n30173 = ~n86 & n3063 ;
  assign n30174 = n86 & n30173 ;
  assign n30175 = n1886 | n3091 ;
  assign n30176 = n30174 & ~n30175 ;
  assign n30177 = n7188 | n30176 ;
  assign n30178 = n30176 & ~n30177 ;
  assign n30179 = n508 | n1304 ;
  assign n30180 = n1304 & ~n30179 ;
  assign n30181 = n30180 ^ n2302 ^ 1'b0 ;
  assign n30182 = n30178 | n30181 ;
  assign n30183 = n30178 & ~n30182 ;
  assign n30166 = n598 & ~n2070 ;
  assign n30167 = ~n598 & n30166 ;
  assign n30168 = n3110 & ~n30167 ;
  assign n30169 = ~n3110 & n30168 ;
  assign n30170 = n367 & ~n1705 ;
  assign n30171 = ~n367 & n30170 ;
  assign n30172 = n30169 & ~n30171 ;
  assign n30184 = n30183 ^ n30172 ^ 1'b0 ;
  assign n30185 = n748 & n2067 ;
  assign n30186 = ~n748 & n30185 ;
  assign n30187 = n11579 & n30186 ;
  assign n30188 = n21607 | n30187 ;
  assign n30189 = n30184 | n30188 ;
  assign n30190 = n20612 ^ n4514 ^ 1'b0 ;
  assign n30191 = n21057 ^ n14195 ^ 1'b0 ;
  assign n30192 = n1937 & n30191 ;
  assign n30193 = n250 & ~n11211 ;
  assign n30194 = n18955 & n30193 ;
  assign n30195 = n4051 & ~n10279 ;
  assign n30196 = n6474 & n30195 ;
  assign n30197 = n227 & n30196 ;
  assign n30198 = n18052 ^ n3679 ^ n2695 ;
  assign n30199 = n2249 | n5549 ;
  assign n30201 = n1608 | n8034 ;
  assign n30200 = n1990 & n13926 ;
  assign n30202 = n30201 ^ n30200 ^ 1'b0 ;
  assign n30203 = n148 | n12157 ;
  assign n30204 = n30203 ^ n9832 ^ 1'b0 ;
  assign n30205 = n7590 | n7853 ;
  assign n30206 = n5010 ^ n1672 ^ 1'b0 ;
  assign n30207 = n30206 ^ n26950 ^ 1'b0 ;
  assign n30208 = n2005 & ~n30207 ;
  assign n30209 = n9265 | n11939 ;
  assign n30210 = n364 & n512 ;
  assign n30211 = ~n3267 & n30210 ;
  assign n30212 = n30211 ^ n17266 ^ 1'b0 ;
  assign n30213 = n3776 | n26424 ;
  assign n30214 = n1241 | n30213 ;
  assign n30215 = n2373 & ~n3709 ;
  assign n30216 = ~n9188 & n30215 ;
  assign n30217 = n5606 ^ n1690 ^ 1'b0 ;
  assign n30218 = ~n30216 & n30217 ;
  assign n30219 = n19184 ^ n7019 ^ 1'b0 ;
  assign n30220 = n14447 & ~n15327 ;
  assign n30221 = n23197 ^ n10495 ^ 1'b0 ;
  assign n30222 = n25674 & n30221 ;
  assign n30224 = n12647 ^ n10651 ^ 1'b0 ;
  assign n30223 = ~n391 & n23602 ;
  assign n30225 = n30224 ^ n30223 ^ 1'b0 ;
  assign n30226 = ( n1948 & ~n10121 ) | ( n1948 & n30225 ) | ( ~n10121 & n30225 ) ;
  assign n30227 = n13453 ^ n8648 ^ n1810 ;
  assign n30228 = n16358 ^ n16035 ^ 1'b0 ;
  assign n30229 = n128 & n30228 ;
  assign n30230 = n310 | n12063 ;
  assign n30231 = n30230 ^ n9486 ^ 1'b0 ;
  assign n30232 = n945 | n4664 ;
  assign n30233 = n22721 ^ n19475 ^ 1'b0 ;
  assign n30234 = n8307 & n10422 ;
  assign n30235 = n30234 ^ n25008 ^ 1'b0 ;
  assign n30236 = n19364 | n30235 ;
  assign n30237 = n3620 | n30236 ;
  assign n30238 = n10493 & ~n12884 ;
  assign n30239 = n30238 ^ n27668 ^ 1'b0 ;
  assign n30240 = n3604 & ~n4751 ;
  assign n30241 = n6594 & n30240 ;
  assign n30242 = n8521 & n30241 ;
  assign n30243 = n1565 | n30242 ;
  assign n30244 = n814 & n26566 ;
  assign n30245 = n30244 ^ n14242 ^ 1'b0 ;
  assign n30246 = ( n2104 & n9275 ) | ( n2104 & n30245 ) | ( n9275 & n30245 ) ;
  assign n30247 = ~n1902 & n5124 ;
  assign n30248 = n8864 & n30247 ;
  assign n30249 = n30248 ^ n7038 ^ 1'b0 ;
  assign n30250 = n7650 | n30249 ;
  assign n30251 = ~n688 & n7043 ;
  assign n30252 = n3046 | n10332 ;
  assign n30253 = n30252 ^ n227 ^ 1'b0 ;
  assign n30254 = n12564 & ~n30253 ;
  assign n30255 = ~n8296 & n30254 ;
  assign n30256 = ~n30251 & n30255 ;
  assign n30257 = n22858 ^ n577 ^ 1'b0 ;
  assign n30258 = n28504 ^ n10052 ^ 1'b0 ;
  assign n30259 = n15 | n19387 ;
  assign n30260 = n2331 & ~n17016 ;
  assign n30261 = n27666 ^ n18121 ^ 1'b0 ;
  assign n30262 = n10500 & ~n16921 ;
  assign n30263 = n11125 ^ n3537 ^ 1'b0 ;
  assign n30264 = n62 & n30263 ;
  assign n30265 = n8889 & n10390 ;
  assign n30266 = n14441 & n30265 ;
  assign n30267 = ~n13220 & n30266 ;
  assign n30268 = n21531 ^ n726 ^ 1'b0 ;
  assign n30269 = n30268 ^ n15136 ^ n547 ;
  assign n30270 = n22228 ^ n10435 ^ 1'b0 ;
  assign n30271 = n15135 & n26457 ;
  assign n30272 = n23523 ^ n22099 ^ 1'b0 ;
  assign n30273 = n30271 | n30272 ;
  assign n30274 = ~n4683 & n13032 ;
  assign n30275 = ~n30273 & n30274 ;
  assign n30276 = ~n15448 & n20100 ;
  assign n30277 = n15242 & n22634 ;
  assign n30278 = n30277 ^ n5675 ^ 1'b0 ;
  assign n30281 = n16513 & n18525 ;
  assign n30282 = n6709 & n30281 ;
  assign n30279 = n10055 & ~n11212 ;
  assign n30280 = n30279 ^ n8347 ^ 1'b0 ;
  assign n30283 = n30282 ^ n30280 ^ 1'b0 ;
  assign n30284 = n325 | n12237 ;
  assign n30286 = n21617 ^ n15429 ^ 1'b0 ;
  assign n30285 = ~n6307 & n27588 ;
  assign n30287 = n30286 ^ n30285 ^ 1'b0 ;
  assign n30288 = n11523 | n15711 ;
  assign n30289 = n7697 | n30288 ;
  assign n30290 = n26147 & n30289 ;
  assign n30291 = ~n21729 & n30290 ;
  assign n30292 = n7807 & n19829 ;
  assign n30293 = ~n9280 & n24708 ;
  assign n30294 = n10115 & n17347 ;
  assign n30295 = n3941 & ~n17031 ;
  assign n30296 = n30294 & n30295 ;
  assign n30297 = n7221 ^ n2574 ^ 1'b0 ;
  assign n30298 = n4121 | n30297 ;
  assign n30299 = n6179 & ~n30298 ;
  assign n30300 = ~n12542 & n30299 ;
  assign n30301 = n17630 ^ n1854 ^ 1'b0 ;
  assign n30302 = n10122 ^ n2560 ^ 1'b0 ;
  assign n30303 = n1081 & ~n30302 ;
  assign n30304 = ( ~n520 & n3109 ) | ( ~n520 & n23753 ) | ( n3109 & n23753 ) ;
  assign n30305 = n5884 ^ n90 ^ 1'b0 ;
  assign n30306 = n30305 ^ n14534 ^ 1'b0 ;
  assign n30307 = ~n10118 & n30306 ;
  assign n30308 = n524 & n30307 ;
  assign n30309 = ~n15321 & n30308 ;
  assign n30310 = n10454 | n18550 ;
  assign n30311 = n23496 | n30310 ;
  assign n30312 = n5607 & n6986 ;
  assign n30313 = n25786 | n30312 ;
  assign n30314 = n19691 | n30313 ;
  assign n30315 = n18086 & ~n30116 ;
  assign n30316 = ~n30314 & n30315 ;
  assign n30317 = ~n1015 & n3570 ;
  assign n30318 = ~n23697 & n30317 ;
  assign n30319 = n13121 & n30318 ;
  assign n30320 = n30319 ^ n12297 ^ n5189 ;
  assign n30321 = n19096 ^ n6012 ^ 1'b0 ;
  assign n30322 = n20099 ^ n19859 ^ 1'b0 ;
  assign n30323 = n38 & n1662 ;
  assign n30324 = ~n1662 & n30323 ;
  assign n30325 = n901 & ~n30324 ;
  assign n30326 = ~n2366 & n7383 ;
  assign n30327 = ~n7383 & n30326 ;
  assign n30328 = n2449 & ~n30327 ;
  assign n30329 = ~n18640 & n30328 ;
  assign n30330 = n30325 & n30329 ;
  assign n30331 = n25356 ^ n6322 ^ 1'b0 ;
  assign n30332 = ~n7419 & n30331 ;
  assign n30333 = n15903 & n30332 ;
  assign n30334 = n608 & ~n8177 ;
  assign n30335 = n3418 ^ n2034 ^ 1'b0 ;
  assign n30350 = x7 & n107 ;
  assign n30351 = ~n107 & n30350 ;
  assign n30352 = n30351 ^ n310 ^ 1'b0 ;
  assign n30353 = n114 & n21911 ;
  assign n30354 = n30352 & ~n30353 ;
  assign n30355 = ~n30352 & n30354 ;
  assign n30356 = n90 | n12141 ;
  assign n30357 = n90 & ~n30356 ;
  assign n30358 = n80 | n30357 ;
  assign n30359 = n80 & ~n30358 ;
  assign n30360 = ~n12580 & n12589 ;
  assign n30361 = n56 & ~n30360 ;
  assign n30362 = ~n56 & n30361 ;
  assign n30363 = n15727 | n30362 ;
  assign n30364 = n30362 & ~n30363 ;
  assign n30365 = n14015 | n30364 ;
  assign n30366 = n30364 & ~n30365 ;
  assign n30367 = n30359 | n30366 ;
  assign n30368 = n30355 & ~n30367 ;
  assign n30369 = n35 & ~n12583 ;
  assign n30370 = n30353 | n30369 ;
  assign n30371 = n30369 & ~n30370 ;
  assign n30372 = n19 | n30351 ;
  assign n30373 = n19 & ~n30372 ;
  assign n30374 = n55 | n255 ;
  assign n30375 = n55 & ~n30374 ;
  assign n30376 = n30373 | n30375 ;
  assign n30377 = n30371 & ~n30376 ;
  assign n30378 = n30368 | n30377 ;
  assign n30379 = n30368 & ~n30378 ;
  assign n30337 = n188 & ~n1479 ;
  assign n30338 = n1479 & n30337 ;
  assign n30339 = n86 & n30338 ;
  assign n30340 = n997 | n30339 ;
  assign n30341 = n30339 & ~n30340 ;
  assign n30342 = x3 | n1202 ;
  assign n30343 = n1202 & ~n30342 ;
  assign n30344 = n32 | n499 ;
  assign n30345 = n30343 & ~n30344 ;
  assign n30346 = n102 & ~n30345 ;
  assign n30347 = n30341 & n30346 ;
  assign n30348 = ~n3717 & n30347 ;
  assign n30349 = n6224 | n30348 ;
  assign n30380 = n30379 ^ n30349 ^ 1'b0 ;
  assign n30381 = ~n491 & n18692 ;
  assign n30386 = n198 | n28791 ;
  assign n30387 = n198 & ~n30386 ;
  assign n30382 = n821 | n3894 ;
  assign n30383 = n3894 & ~n30382 ;
  assign n30384 = n1394 & ~n30383 ;
  assign n30385 = n30383 & n30384 ;
  assign n30388 = n30387 ^ n30385 ^ 1'b0 ;
  assign n30389 = n30381 & n30388 ;
  assign n30390 = ~n5112 & n30389 ;
  assign n30391 = n2178 & n30390 ;
  assign n30392 = n252 & n800 ;
  assign n30393 = ~n800 & n30392 ;
  assign n30394 = ~n698 & n903 ;
  assign n30395 = n698 & n30394 ;
  assign n30396 = n292 & ~n30395 ;
  assign n30397 = ~n292 & n30396 ;
  assign n30398 = n1560 | n30397 ;
  assign n30399 = n30393 & ~n30398 ;
  assign n30400 = n622 & ~n30399 ;
  assign n30401 = ~n622 & n30400 ;
  assign n30402 = n30401 ^ n2542 ^ 1'b0 ;
  assign n30403 = ~n30391 & n30402 ;
  assign n30404 = n30391 & n30403 ;
  assign n30405 = n2090 | n30404 ;
  assign n30406 = n2090 & ~n30405 ;
  assign n30407 = n5574 | n30406 ;
  assign n30408 = n30380 & ~n30407 ;
  assign n30336 = ~n1602 & n23852 ;
  assign n30409 = n30408 ^ n30336 ^ 1'b0 ;
  assign n30410 = n133 | n16647 ;
  assign n30411 = ~n16784 & n30410 ;
  assign n30412 = n12547 ^ n6251 ^ 1'b0 ;
  assign n30413 = n1113 & n6046 ;
  assign n30414 = n30413 ^ n2303 ^ 1'b0 ;
  assign n30415 = ~n139 & n4126 ;
  assign n30416 = n20323 | n30415 ;
  assign n30417 = n7497 & n7503 ;
  assign n30418 = n15426 ^ n8362 ^ 1'b0 ;
  assign n30419 = n30417 & n30418 ;
  assign n30420 = ~n9362 & n14648 ;
  assign n30421 = n30420 ^ n2843 ^ 1'b0 ;
  assign n30422 = ~n1885 & n20492 ;
  assign n30423 = n30421 & n30422 ;
  assign n30424 = n5573 | n15458 ;
  assign n30425 = n20030 & ~n21721 ;
  assign n30426 = n10767 & n30425 ;
  assign n30427 = n30426 ^ n14466 ^ 1'b0 ;
  assign n30428 = n2332 & n18107 ;
  assign n30429 = n30427 & n30428 ;
  assign n30430 = n14881 | n30429 ;
  assign n30431 = n5218 & n14469 ;
  assign n30432 = n15015 & n23299 ;
  assign n30433 = n23681 ^ n6997 ^ 1'b0 ;
  assign n30434 = n30433 ^ n4019 ^ n3394 ;
  assign n30435 = n5928 & n30434 ;
  assign n30436 = n7051 & n13501 ;
  assign n30437 = n7627 | n26061 ;
  assign n30438 = ~n3742 & n30437 ;
  assign n30440 = n12741 ^ n1036 ^ 1'b0 ;
  assign n30441 = n323 & ~n30440 ;
  assign n30442 = n9197 | n10180 ;
  assign n30443 = n1368 & ~n30442 ;
  assign n30444 = ~n30441 & n30443 ;
  assign n30439 = ~n5747 & n13554 ;
  assign n30445 = n30444 ^ n30439 ^ 1'b0 ;
  assign n30446 = n30445 ^ n9364 ^ 1'b0 ;
  assign n30447 = n7737 & ~n15288 ;
  assign n30448 = ~n12976 & n30447 ;
  assign n30449 = n29742 ^ n5285 ^ 1'b0 ;
  assign n30450 = n30092 ^ n8870 ^ 1'b0 ;
  assign n30451 = n8247 ^ n5938 ^ 1'b0 ;
  assign n30452 = n9890 & n30451 ;
  assign n30453 = ~n3367 & n11193 ;
  assign n30454 = n30453 ^ n22267 ^ 1'b0 ;
  assign n30455 = n30452 & ~n30454 ;
  assign n30456 = n17812 ^ n917 ^ 1'b0 ;
  assign n30457 = n4197 & n5533 ;
  assign n30458 = ~n30456 & n30457 ;
  assign n30459 = n30458 ^ n5713 ^ n3793 ;
  assign n30460 = n13810 | n30459 ;
  assign n30461 = ( n2917 & n8219 ) | ( n2917 & ~n9806 ) | ( n8219 & ~n9806 ) ;
  assign n30462 = n5428 ^ n2463 ^ 1'b0 ;
  assign n30463 = n30462 ^ n16255 ^ 1'b0 ;
  assign n30464 = n30461 | n30463 ;
  assign n30465 = ~n10426 & n27670 ;
  assign n30466 = n30465 ^ n5567 ^ 1'b0 ;
  assign n30467 = n3131 | n25499 ;
  assign n30468 = n25990 | n30467 ;
  assign n30469 = ~n4237 & n7237 ;
  assign n30470 = ~n1188 & n15126 ;
  assign n30471 = ~n929 & n30470 ;
  assign n30472 = ~n2799 & n4115 ;
  assign n30473 = n30085 ^ n10190 ^ 1'b0 ;
  assign n30474 = n11047 ^ n4872 ^ 1'b0 ;
  assign n30475 = ~n12996 & n30474 ;
  assign n30480 = n27802 ^ n19895 ^ 1'b0 ;
  assign n30476 = n560 & n1572 ;
  assign n30477 = ~n18721 & n30476 ;
  assign n30478 = n5461 | n30477 ;
  assign n30479 = ~n2497 & n30478 ;
  assign n30481 = n30480 ^ n30479 ^ 1'b0 ;
  assign n30482 = ~n7355 & n10122 ;
  assign n30483 = n30482 ^ n9322 ^ 1'b0 ;
  assign n30484 = n23956 & n26431 ;
  assign n30485 = n30484 ^ n27527 ^ 1'b0 ;
  assign n30486 = n1909 | n9357 ;
  assign n30487 = n1771 | n30486 ;
  assign n30488 = ~n7056 & n30487 ;
  assign n30489 = n47 & n27555 ;
  assign n30490 = ~n13926 & n30489 ;
  assign n30491 = n5237 & ~n19789 ;
  assign n30492 = n21495 & ~n27063 ;
  assign n30493 = n16020 | n30492 ;
  assign n30494 = n16302 ^ n5806 ^ 1'b0 ;
  assign n30495 = n11586 & ~n30494 ;
  assign n30496 = n30495 ^ n3007 ^ 1'b0 ;
  assign n30497 = n8527 & ~n25782 ;
  assign n30498 = n30497 ^ n5538 ^ n3877 ;
  assign n30499 = n25075 ^ n8264 ^ 1'b0 ;
  assign n30500 = n7667 | n26586 ;
  assign n30501 = n18977 & ~n30500 ;
  assign n30502 = n5928 & n30501 ;
  assign n30503 = n83 & ~n6392 ;
  assign n30504 = n30503 ^ n2850 ^ 1'b0 ;
  assign n30505 = n16607 & ~n30504 ;
  assign n30506 = ~n5610 & n30505 ;
  assign n30507 = ~n30502 & n30506 ;
  assign n30508 = ( n4919 & ~n8396 ) | ( n4919 & n11977 ) | ( ~n8396 & n11977 ) ;
  assign n30509 = n4109 | n27246 ;
  assign n30510 = n1961 & ~n30509 ;
  assign n30511 = n18186 & ~n23842 ;
  assign n30512 = n30511 ^ n10203 ^ 1'b0 ;
  assign n30513 = n30512 ^ n7301 ^ 1'b0 ;
  assign n30514 = ~n30510 & n30513 ;
  assign n30515 = n13121 ^ n3452 ^ 1'b0 ;
  assign n30516 = n19299 & ~n30515 ;
  assign n30517 = n22312 ^ n2661 ^ 1'b0 ;
  assign n30518 = n8470 | n14544 ;
  assign n30519 = n15469 & ~n30518 ;
  assign n30520 = n30519 ^ n12193 ^ 1'b0 ;
  assign n30521 = n2906 & n30520 ;
  assign n30522 = n7728 & n30521 ;
  assign n30523 = n5063 ^ n4561 ^ 1'b0 ;
  assign n30524 = ~n8764 & n30523 ;
  assign n30525 = n15680 ^ n6301 ^ 1'b0 ;
  assign n30526 = n30524 & ~n30525 ;
  assign n30527 = n662 | n2178 ;
  assign n30528 = n30527 ^ n817 ^ 1'b0 ;
  assign n30529 = n11498 & n30528 ;
  assign n30530 = n2733 & n30529 ;
  assign n30531 = ~n565 & n2686 ;
  assign n30532 = n30531 ^ n5956 ^ 1'b0 ;
  assign n30533 = n30532 ^ n6001 ^ 1'b0 ;
  assign n30534 = ~n1113 & n30533 ;
  assign n30535 = n30534 ^ n12271 ^ 1'b0 ;
  assign n30536 = n501 | n3869 ;
  assign n30537 = n7789 | n8793 ;
  assign n30538 = n30537 ^ n16598 ^ n3408 ;
  assign n30539 = n1217 | n6596 ;
  assign n30540 = ~n4646 & n19012 ;
  assign n30541 = n1227 | n12257 ;
  assign n30542 = ~n10253 & n30541 ;
  assign n30543 = n20819 ^ n17197 ^ 1'b0 ;
  assign n30544 = ~n599 & n5590 ;
  assign n30545 = n5652 & n26489 ;
  assign n30546 = n2929 & n13417 ;
  assign n30547 = n27353 | n30546 ;
  assign n30548 = ~n7667 & n7857 ;
  assign n30549 = n1804 | n30548 ;
  assign n30550 = n8121 ^ x3 ^ 1'b0 ;
  assign n30551 = ~n30549 & n30550 ;
  assign n30552 = n24185 & ~n30551 ;
  assign n30553 = n1817 | n30552 ;
  assign n30554 = n9134 & ~n30553 ;
  assign n30555 = ~n15210 & n25954 ;
  assign n30556 = n22832 & n30555 ;
  assign n30557 = n11260 & n30556 ;
  assign n30558 = ~n670 & n23057 ;
  assign n30559 = n30558 ^ n25782 ^ n3237 ;
  assign n30560 = n4712 ^ n144 ^ 1'b0 ;
  assign n30561 = ~n6474 & n11414 ;
  assign n30562 = n27610 & n30561 ;
  assign n30563 = n23553 & ~n30562 ;
  assign n30564 = ~n7523 & n30563 ;
  assign n30565 = n12500 ^ n5423 ^ 1'b0 ;
  assign n30566 = n10743 & n30565 ;
  assign n30567 = ~n3176 & n30566 ;
  assign n30568 = n156 & n715 ;
  assign n30569 = n1124 & ~n3967 ;
  assign n30570 = n3967 & n30569 ;
  assign n30571 = ~n6307 & n30570 ;
  assign n30572 = n17176 & n30571 ;
  assign n30585 = ~n17 & n1052 ;
  assign n30586 = n17 & n30585 ;
  assign n30587 = ~n17082 & n30586 ;
  assign n30573 = n423 & n3729 ;
  assign n30574 = ~n423 & n30573 ;
  assign n30575 = ~n159 & n30574 ;
  assign n30576 = n30575 ^ n1933 ^ 1'b0 ;
  assign n30577 = n263 & n1152 ;
  assign n30578 = ~n263 & n30577 ;
  assign n30579 = ~n1672 & n30578 ;
  assign n30580 = ~n321 & n1519 ;
  assign n30581 = n30579 & n30580 ;
  assign n30582 = n4202 & ~n30581 ;
  assign n30583 = ~n4202 & n30582 ;
  assign n30584 = n30576 & ~n30583 ;
  assign n30588 = n30587 ^ n30584 ^ 1'b0 ;
  assign n30589 = n8904 | n30588 ;
  assign n30590 = n30572 | n30589 ;
  assign n30591 = n21119 ^ n1102 ^ 1'b0 ;
  assign n30592 = n11159 & ~n30591 ;
  assign n30593 = n2260 & ~n10451 ;
  assign n30594 = n6492 & n30593 ;
  assign n30595 = n21082 & n30594 ;
  assign n30596 = n8937 | n29585 ;
  assign n30597 = n4700 ^ n231 ^ 1'b0 ;
  assign n30598 = ~n6538 & n30597 ;
  assign n30599 = n9937 | n14411 ;
  assign n30600 = n4236 & ~n30599 ;
  assign n30601 = n8280 & ~n30600 ;
  assign n30602 = n7753 & n30601 ;
  assign n30603 = n1541 | n4419 ;
  assign n30604 = n817 & ~n30603 ;
  assign n30605 = n14561 | n18402 ;
  assign n30606 = n235 | n30605 ;
  assign n30607 = n30606 ^ n10019 ^ 1'b0 ;
  assign n30608 = n11178 & ~n14561 ;
  assign n30609 = n30608 ^ n18711 ^ 1'b0 ;
  assign n30610 = n25060 & ~n30609 ;
  assign n30611 = n27405 ^ n24986 ^ 1'b0 ;
  assign n30612 = n3800 & n30611 ;
  assign n30613 = n16519 ^ n5380 ^ 1'b0 ;
  assign n30614 = n16983 ^ n9980 ^ 1'b0 ;
  assign n30615 = n30613 & n30614 ;
  assign n30616 = n8186 | n8959 ;
  assign n30617 = n30616 ^ n12252 ^ n2511 ;
  assign n30618 = n14083 ^ n4803 ^ 1'b0 ;
  assign n30619 = n2436 & n30618 ;
  assign n30620 = ~n5269 & n10232 ;
  assign n30621 = n11596 ^ n1415 ^ 1'b0 ;
  assign n30622 = n12982 | n30621 ;
  assign n30623 = n15915 | n30622 ;
  assign n30624 = n2155 & n5128 ;
  assign n30625 = n5146 & n5332 ;
  assign n30626 = n17156 ^ n16065 ^ 1'b0 ;
  assign n30627 = n17078 & ~n30626 ;
  assign n30628 = n2162 & ~n30627 ;
  assign n30629 = n3042 | n6536 ;
  assign n30630 = ~n12284 & n30629 ;
  assign n30631 = n14164 & n30630 ;
  assign n30632 = n1947 & ~n2786 ;
  assign n30633 = n30632 ^ n1867 ^ 1'b0 ;
  assign n30634 = n26385 ^ n8764 ^ 1'b0 ;
  assign n30635 = n17283 | n30634 ;
  assign n30636 = n102 & n24756 ;
  assign n30637 = n14618 & n30636 ;
  assign n30638 = n28826 ^ n3698 ^ 1'b0 ;
  assign n30639 = n26403 & ~n30638 ;
  assign n30640 = ~n12734 & n30639 ;
  assign n30641 = ~n14356 & n30640 ;
  assign n30642 = n7524 ^ n6663 ^ 1'b0 ;
  assign n30643 = n3412 | n4899 ;
  assign n30644 = ~n962 & n11731 ;
  assign n30645 = n15475 & n30644 ;
  assign n30646 = n30645 ^ n22131 ^ 1'b0 ;
  assign n30647 = ~n20263 & n21146 ;
  assign n30648 = n19298 & n30647 ;
  assign n30649 = ~n10561 & n30648 ;
  assign n30650 = n25315 ^ n14138 ^ 1'b0 ;
  assign n30651 = n17014 ^ n62 ^ 1'b0 ;
  assign n30652 = ~n10504 & n30651 ;
  assign n30653 = n16 & n15552 ;
  assign n30654 = n4245 & ~n10751 ;
  assign n30655 = ~n3032 & n30654 ;
  assign n30656 = n30655 ^ n16363 ^ 1'b0 ;
  assign n30658 = n6897 & n16283 ;
  assign n30657 = n1473 | n2694 ;
  assign n30659 = n30658 ^ n30657 ^ 1'b0 ;
  assign n30662 = n5685 | n25460 ;
  assign n30660 = n16088 & n26262 ;
  assign n30661 = ~n439 & n30660 ;
  assign n30663 = n30662 ^ n30661 ^ 1'b0 ;
  assign n30664 = n8396 ^ n1716 ^ 1'b0 ;
  assign n30665 = n30664 ^ n3369 ^ 1'b0 ;
  assign n30667 = n901 & ~n1409 ;
  assign n30668 = n4549 ^ n1768 ^ 1'b0 ;
  assign n30669 = ~n30667 & n30668 ;
  assign n30670 = ~n5185 & n30669 ;
  assign n30671 = n30670 ^ n15782 ^ 1'b0 ;
  assign n30666 = n3642 | n15493 ;
  assign n30672 = n30671 ^ n30666 ^ 1'b0 ;
  assign n30673 = n26776 ^ n3265 ^ 1'b0 ;
  assign n30674 = n9661 & ~n22299 ;
  assign n30675 = n30674 ^ n30528 ^ 1'b0 ;
  assign n30676 = n8034 ^ n5917 ^ 1'b0 ;
  assign n30677 = n16170 | n30676 ;
  assign n30678 = n4400 & n8833 ;
  assign n30679 = ( n2627 & ~n30677 ) | ( n2627 & n30678 ) | ( ~n30677 & n30678 ) ;
  assign n30680 = ~n231 & n5685 ;
  assign n30681 = n8412 | n13263 ;
  assign n30682 = n30681 ^ n2883 ^ 1'b0 ;
  assign n30683 = n13678 ^ n397 ^ 1'b0 ;
  assign n30684 = n6777 | n30683 ;
  assign n30685 = n1902 | n27933 ;
  assign n30686 = n14995 & ~n30685 ;
  assign n30687 = n30686 ^ n20676 ^ n5794 ;
  assign n30688 = n4559 | n6016 ;
  assign n30689 = n30687 & ~n30688 ;
  assign n30690 = n21848 & n25700 ;
  assign n30691 = n30690 ^ n2378 ^ 1'b0 ;
  assign n30692 = n5241 | n20758 ;
  assign n30693 = n2205 | n30692 ;
  assign n30694 = n30693 ^ n15441 ^ 1'b0 ;
  assign n30695 = n18735 ^ n3857 ^ 1'b0 ;
  assign n30696 = n5011 & ~n30695 ;
  assign n30697 = n13687 ^ n1608 ^ n374 ;
  assign n30698 = n30696 & ~n30697 ;
  assign n30699 = ~n1130 & n16714 ;
  assign n30700 = n213 | n7038 ;
  assign n30701 = n30700 ^ n10586 ^ 1'b0 ;
  assign n30702 = n15468 & ~n30701 ;
  assign n30703 = n13277 & n30702 ;
  assign n30704 = n6408 & ~n30703 ;
  assign n30705 = n30704 ^ n8416 ^ 1'b0 ;
  assign n30706 = n310 | n23288 ;
  assign n30707 = n15814 & ~n18824 ;
  assign n30708 = n30706 & n30707 ;
  assign n30709 = n29109 | n30708 ;
  assign n30710 = n30709 ^ n599 ^ 1'b0 ;
  assign n30711 = n1560 | n19554 ;
  assign n30712 = n30711 ^ n6944 ^ 1'b0 ;
  assign n30713 = n942 & n30712 ;
  assign n30714 = n5685 & ~n12016 ;
  assign n30715 = n24449 ^ n14706 ^ 1'b0 ;
  assign n30716 = n10429 | n17502 ;
  assign n30717 = n12777 ^ n12400 ^ n419 ;
  assign n30718 = n1501 & n15292 ;
  assign n30719 = n23152 ^ n23001 ^ 1'b0 ;
  assign n30720 = n18276 | n30719 ;
  assign n30721 = n2200 | n23734 ;
  assign n30722 = n30721 ^ n16582 ^ 1'b0 ;
  assign n30723 = n22185 ^ n12418 ^ 1'b0 ;
  assign n30724 = ~n16360 & n22215 ;
  assign n30725 = ~n3177 & n10153 ;
  assign n30732 = n5253 | n13263 ;
  assign n30733 = n13263 & ~n30732 ;
  assign n30726 = n4869 & n19927 ;
  assign n30727 = n11722 & ~n30726 ;
  assign n30728 = n21311 & ~n30727 ;
  assign n30729 = n2311 & n30728 ;
  assign n30730 = n30729 ^ n10060 ^ 1'b0 ;
  assign n30731 = n25808 & n30730 ;
  assign n30734 = n30733 ^ n30731 ^ 1'b0 ;
  assign n30735 = n323 & ~n1458 ;
  assign n30736 = n6152 & ~n30735 ;
  assign n30737 = n17872 & ~n24097 ;
  assign n30738 = n30737 ^ n12866 ^ 1'b0 ;
  assign n30739 = n12517 ^ n3347 ^ 1'b0 ;
  assign n30740 = n7040 | n18315 ;
  assign n30741 = ( n18144 & ~n22130 ) | ( n18144 & n24057 ) | ( ~n22130 & n24057 ) ;
  assign n30742 = n5640 | n13682 ;
  assign n30743 = n30742 ^ n26388 ^ 1'b0 ;
  assign n30744 = ~n15883 & n28335 ;
  assign n30745 = n17969 | n26007 ;
  assign n30746 = ( n7596 & n10571 ) | ( n7596 & n17475 ) | ( n10571 & n17475 ) ;
  assign n30747 = n17854 ^ n495 ^ 1'b0 ;
  assign n30748 = n11895 & ~n30747 ;
  assign n30749 = n16416 | n24511 ;
  assign n30750 = n3040 | n5684 ;
  assign n30751 = n154 & n30750 ;
  assign n30752 = ~n14701 & n30751 ;
  assign n30753 = n3459 & ~n12730 ;
  assign n30754 = n30753 ^ n2730 ^ 1'b0 ;
  assign n30755 = n2433 & ~n30754 ;
  assign n30756 = n18033 ^ n12211 ^ 1'b0 ;
  assign n30757 = n11531 ^ n3600 ^ 1'b0 ;
  assign n30758 = n12976 ^ n5187 ^ 1'b0 ;
  assign n30759 = n8680 & ~n14686 ;
  assign n30760 = n14556 & ~n19226 ;
  assign n30761 = n2294 & ~n15147 ;
  assign n30762 = n22070 ^ n7531 ^ 1'b0 ;
  assign n30763 = n30761 | n30762 ;
  assign n30764 = n5286 & n14422 ;
  assign n30765 = ~n10124 & n30764 ;
  assign n30766 = n1547 & n24890 ;
  assign n30767 = n12810 & n30766 ;
  assign n30768 = n1795 & n3068 ;
  assign n30769 = n8326 ^ n2924 ^ 1'b0 ;
  assign n30770 = n16513 & n30769 ;
  assign n30771 = n30770 ^ n23038 ^ 1'b0 ;
  assign n30772 = n7550 | n11827 ;
  assign n30773 = n4400 & ~n30772 ;
  assign n30774 = ~n17612 & n25267 ;
  assign n30775 = n30774 ^ n3459 ^ 1'b0 ;
  assign n30776 = ~n11466 & n19437 ;
  assign n30777 = ~n2022 & n13847 ;
  assign n30778 = n6295 ^ n520 ^ 1'b0 ;
  assign n30779 = n11740 ^ n7915 ^ 1'b0 ;
  assign n30780 = ~n10429 & n30779 ;
  assign n30781 = ~n8734 & n30780 ;
  assign n30782 = n11027 ^ n290 ^ 1'b0 ;
  assign n30783 = n258 & n22876 ;
  assign n30784 = ~n395 & n18430 ;
  assign n30785 = ~n30783 & n30784 ;
  assign n30786 = n21411 | n30785 ;
  assign n30787 = n2168 | n3380 ;
  assign n30788 = n4419 ^ n3933 ^ 1'b0 ;
  assign n30789 = n9697 ^ n6919 ^ 1'b0 ;
  assign n30790 = ~n1602 & n5683 ;
  assign n30791 = n2435 ^ n137 ^ 1'b0 ;
  assign n30792 = n915 | n26786 ;
  assign n30793 = n4092 & n25069 ;
  assign n30794 = n9131 ^ n5196 ^ 1'b0 ;
  assign n30795 = ~n13748 & n30794 ;
  assign n30796 = n20224 | n30795 ;
  assign n30797 = n5056 | n30796 ;
  assign n30798 = n30797 ^ n8862 ^ 1'b0 ;
  assign n30799 = n3211 & n30798 ;
  assign n30800 = n25948 & ~n26061 ;
  assign n30801 = n5562 & n11656 ;
  assign n30802 = ~n2150 & n2506 ;
  assign n30803 = ~n9119 & n9131 ;
  assign n30804 = n43 & n30803 ;
  assign n30805 = n2136 & n8933 ;
  assign n30806 = n13887 | n30805 ;
  assign n30807 = ( n2005 & ~n3138 ) | ( n2005 & n7288 ) | ( ~n3138 & n7288 ) ;
  assign n30808 = n654 & ~n3423 ;
  assign n30809 = n14789 & n29741 ;
  assign n30810 = ~n22215 & n30809 ;
  assign n30811 = n27854 ^ n27240 ^ 1'b0 ;
  assign n30812 = n13099 & ~n30811 ;
  assign n30813 = ~n5161 & n29836 ;
  assign n30814 = n30813 ^ n16102 ^ 1'b0 ;
  assign n30815 = n581 | n11615 ;
  assign n30816 = n7652 & ~n30815 ;
  assign n30817 = n6755 | n23546 ;
  assign n30818 = n30817 ^ n13874 ^ 1'b0 ;
  assign n30819 = n9384 & n30818 ;
  assign n30820 = n7448 & n7468 ;
  assign n30821 = n4748 & ~n13089 ;
  assign n30822 = n30821 ^ n28274 ^ 1'b0 ;
  assign n30823 = n3807 | n16677 ;
  assign n30824 = n14739 ^ n10076 ^ 1'b0 ;
  assign n30825 = n16315 | n16748 ;
  assign n30826 = n30825 ^ n4552 ^ 1'b0 ;
  assign n30827 = ~n4853 & n21045 ;
  assign n30828 = n6165 ^ n6037 ^ 1'b0 ;
  assign n30829 = ~n7596 & n30828 ;
  assign n30830 = n12547 ^ n6385 ^ 1'b0 ;
  assign n30831 = ~n23057 & n30830 ;
  assign n30832 = ~n4314 & n5882 ;
  assign n30833 = n25493 | n30832 ;
  assign n30834 = n2939 | n30833 ;
  assign n30835 = ~n932 & n10384 ;
  assign n30836 = n30835 ^ n1666 ^ 1'b0 ;
  assign n30837 = n4483 & n30836 ;
  assign n30838 = n30837 ^ n7381 ^ 1'b0 ;
  assign n30839 = n6454 ^ n2388 ^ 1'b0 ;
  assign n30840 = ( ~n4373 & n8500 ) | ( ~n4373 & n30839 ) | ( n8500 & n30839 ) ;
  assign n30841 = n14043 ^ n7936 ^ 1'b0 ;
  assign n30842 = n5290 & ~n12440 ;
  assign n30843 = n22744 ^ n567 ^ 1'b0 ;
  assign n30844 = n30842 | n30843 ;
  assign n30845 = n14235 ^ n12105 ^ 1'b0 ;
  assign n30846 = ~n9427 & n30845 ;
  assign n30847 = n28817 & n30846 ;
  assign n30848 = n19875 ^ n13348 ^ 1'b0 ;
  assign n30849 = n4194 & ~n22231 ;
  assign n30850 = n24722 & ~n30849 ;
  assign n30851 = n30850 ^ n23700 ^ 1'b0 ;
  assign n30852 = ~n19933 & n30851 ;
  assign n30853 = n4878 & n30532 ;
  assign n30854 = ~n3071 & n30853 ;
  assign n30855 = n10976 ^ n552 ^ 1'b0 ;
  assign n30856 = n286 & ~n30855 ;
  assign n30857 = n30856 ^ n16310 ^ 1'b0 ;
  assign n30858 = n30854 & ~n30857 ;
  assign n30859 = n8818 | n13079 ;
  assign n30860 = ~n390 & n3828 ;
  assign n30863 = n17275 ^ n6773 ^ 1'b0 ;
  assign n30864 = n18624 ^ n14954 ^ 1'b0 ;
  assign n30865 = ~n30863 & n30864 ;
  assign n30861 = n5801 ^ n3816 ^ 1'b0 ;
  assign n30862 = n26462 | n30861 ;
  assign n30866 = n30865 ^ n30862 ^ 1'b0 ;
  assign n30867 = n4660 & ~n9335 ;
  assign n30868 = n20288 & ~n29466 ;
  assign n30869 = ~n24079 & n25952 ;
  assign n30870 = n9697 & ~n25926 ;
  assign n30871 = n25047 ^ n12119 ^ 1'b0 ;
  assign n30872 = ~n158 & n13298 ;
  assign n30873 = n21157 ^ n9307 ^ n3164 ;
  assign n30874 = n17519 ^ n12265 ^ 1'b0 ;
  assign n30875 = n29066 | n30874 ;
  assign n30876 = n7388 ^ n4250 ^ 1'b0 ;
  assign n30877 = n30875 & ~n30876 ;
  assign n30878 = n17684 & n27872 ;
  assign n30879 = x6 & n10393 ;
  assign n30880 = n30879 ^ n6073 ^ 1'b0 ;
  assign n30881 = ~n2324 & n30880 ;
  assign n30882 = ~n30878 & n30881 ;
  assign n30883 = n8623 & ~n30882 ;
  assign n30884 = n2591 & n30883 ;
  assign n30885 = n30884 ^ n12998 ^ 1'b0 ;
  assign n30886 = ~n3773 & n5707 ;
  assign n30887 = ~n13915 & n30886 ;
  assign n30888 = ~n10790 & n30887 ;
  assign n30889 = n30888 ^ n7193 ^ 1'b0 ;
  assign n30890 = n9247 | n16305 ;
  assign n30891 = ~n1638 & n30890 ;
  assign n30892 = n30891 ^ n27486 ^ 1'b0 ;
  assign n30893 = n4156 | n9482 ;
  assign n30894 = n11806 ^ n7801 ^ 1'b0 ;
  assign n30895 = ( n931 & ~n2790 ) | ( n931 & n30894 ) | ( ~n2790 & n30894 ) ;
  assign n30896 = n1927 & n15054 ;
  assign n30897 = ~n3939 & n30896 ;
  assign n30898 = n2199 | n17935 ;
  assign n30899 = ~n5178 & n30898 ;
  assign n30900 = n7145 & n30899 ;
  assign n30901 = n30900 ^ n4883 ^ 1'b0 ;
  assign n30902 = n11673 & ~n16777 ;
  assign n30903 = n30902 ^ n380 ^ 1'b0 ;
  assign n30904 = ~n7422 & n24933 ;
  assign n30905 = n7422 & n30904 ;
  assign n30906 = n944 & ~n30905 ;
  assign n30907 = n11764 & n30906 ;
  assign n30908 = ~n21291 & n29724 ;
  assign n30909 = n23558 ^ n10398 ^ 1'b0 ;
  assign n30910 = ~n28838 & n30909 ;
  assign n30911 = n4860 & n5201 ;
  assign n30912 = n12387 & n30911 ;
  assign n30913 = n4250 | n12444 ;
  assign n30914 = n158 & ~n2538 ;
  assign n30915 = ~n4069 & n30914 ;
  assign n30916 = ~n8804 & n30915 ;
  assign n30917 = ~n1814 & n4112 ;
  assign n30918 = n30917 ^ n294 ^ 1'b0 ;
  assign n30919 = n30916 | n30918 ;
  assign n30920 = n30913 | n30919 ;
  assign n30921 = n10559 ^ n4850 ^ 1'b0 ;
  assign n30922 = n5180 | n30921 ;
  assign n30923 = n3788 & ~n10937 ;
  assign n30924 = n30922 & n30923 ;
  assign n30925 = n1048 & n30924 ;
  assign n30926 = n16651 | n30925 ;
  assign n30927 = n15910 & n30926 ;
  assign n30928 = n25808 ^ n4954 ^ 1'b0 ;
  assign n30929 = n3744 & ~n30928 ;
  assign n30930 = n25464 & n30929 ;
  assign n30931 = n11044 | n15322 ;
  assign n30932 = n30931 ^ n26336 ^ 1'b0 ;
  assign n30933 = n23594 ^ n364 ^ 1'b0 ;
  assign n30934 = n348 & ~n30933 ;
  assign n30935 = n30934 ^ n23865 ^ 1'b0 ;
  assign n30936 = n5957 ^ n4650 ^ 1'b0 ;
  assign n30937 = n27370 ^ n14432 ^ 1'b0 ;
  assign n30938 = n30936 & n30937 ;
  assign n30939 = n3837 | n17253 ;
  assign n30940 = n2034 & ~n9757 ;
  assign n30941 = n3663 & n30940 ;
  assign n30942 = n30941 ^ n5542 ^ 1'b0 ;
  assign n30943 = ~n14566 & n23508 ;
  assign n30945 = n6745 ^ n1865 ^ 1'b0 ;
  assign n30944 = n20395 & ~n27771 ;
  assign n30946 = n30945 ^ n30944 ^ 1'b0 ;
  assign n30947 = ~n5575 & n6082 ;
  assign n30948 = ~n24469 & n30947 ;
  assign n30949 = ~n2061 & n5288 ;
  assign n30950 = n1254 & n10740 ;
  assign n30951 = n30950 ^ n10581 ^ 1'b0 ;
  assign n30952 = n6045 ^ n5560 ^ n5551 ;
  assign n30953 = n10936 & ~n30952 ;
  assign n30954 = ~n2853 & n30953 ;
  assign n30955 = n11726 & n24273 ;
  assign n30956 = n30955 ^ n6085 ^ 1'b0 ;
  assign n30957 = n310 & ~n8389 ;
  assign n30958 = n30956 & n30957 ;
  assign n30959 = n28165 ^ n21404 ^ 1'b0 ;
  assign n30960 = n10242 | n28102 ;
  assign n30961 = n3366 & n16136 ;
  assign n30962 = n2883 ^ n653 ^ 1'b0 ;
  assign n30963 = n3108 & n11296 ;
  assign n30964 = ~n14432 & n30963 ;
  assign n30965 = n30962 | n30964 ;
  assign n30966 = n292 & n24852 ;
  assign n30967 = ~n11551 & n20484 ;
  assign n30968 = n5936 & n30967 ;
  assign n30969 = n23678 ^ n14427 ^ 1'b0 ;
  assign n30970 = n30968 & ~n30969 ;
  assign n30971 = n2627 | n3594 ;
  assign n30972 = n5033 ^ n1619 ^ 1'b0 ;
  assign n30973 = n1385 & ~n21642 ;
  assign n30974 = n10224 & ~n27240 ;
  assign n30975 = ~n6748 & n30974 ;
  assign n30976 = n9429 & n19843 ;
  assign n30977 = n2303 & ~n14339 ;
  assign n30978 = n928 & ~n13090 ;
  assign n30979 = n5726 & ~n30978 ;
  assign n30980 = n16358 ^ n62 ^ 1'b0 ;
  assign n30981 = n11931 & ~n13693 ;
  assign n30982 = ~n9901 & n30981 ;
  assign n30983 = ~n2324 & n30982 ;
  assign n30984 = ~n390 & n15293 ;
  assign n30985 = n30984 ^ n11588 ^ 1'b0 ;
  assign n30987 = n11755 ^ n8674 ^ 1'b0 ;
  assign n30986 = ~n4286 & n28131 ;
  assign n30988 = n30987 ^ n30986 ^ 1'b0 ;
  assign n30989 = n16675 | n30988 ;
  assign n30990 = n30985 | n30989 ;
  assign n30991 = n4029 ^ n1655 ^ 1'b0 ;
  assign n30992 = ( ~n12298 & n12799 ) | ( ~n12298 & n30991 ) | ( n12799 & n30991 ) ;
  assign n30993 = n17942 & n30992 ;
  assign n30994 = n6106 & n13760 ;
  assign n30995 = n4061 | n30994 ;
  assign n30996 = n8904 ^ n7951 ^ 1'b0 ;
  assign n30997 = ~n882 & n17787 ;
  assign n30998 = ~n729 & n30997 ;
  assign n31004 = n632 & ~n670 ;
  assign n30999 = n603 & n5707 ;
  assign n31000 = n30999 ^ n7646 ^ 1'b0 ;
  assign n31001 = ~n1309 & n31000 ;
  assign n31002 = n31001 ^ n9051 ^ 1'b0 ;
  assign n31003 = n13040 & n31002 ;
  assign n31005 = n31004 ^ n31003 ^ 1'b0 ;
  assign n31006 = n21784 ^ n4774 ^ n1300 ;
  assign n31007 = n22819 ^ n4036 ^ 1'b0 ;
  assign n31008 = n30240 ^ n10438 ^ 1'b0 ;
  assign n31009 = n31007 & ~n31008 ;
  assign n31010 = n3579 & n31009 ;
  assign n31011 = ~n2378 & n19332 ;
  assign n31012 = ~n2762 & n31011 ;
  assign n31013 = n2102 & n5971 ;
  assign n31014 = ~n21433 & n31013 ;
  assign n31015 = n3643 & ~n31014 ;
  assign n31016 = ~n11673 & n31015 ;
  assign n31017 = n11187 ^ n2029 ^ 1'b0 ;
  assign n31018 = n562 & n4568 ;
  assign n31019 = n13098 ^ n582 ^ 1'b0 ;
  assign n31020 = ~n6429 & n31019 ;
  assign n31021 = n31020 ^ n8251 ^ 1'b0 ;
  assign n31022 = ~n3586 & n22325 ;
  assign n31023 = n18148 ^ n10607 ^ 1'b0 ;
  assign n31024 = n20364 & ~n31023 ;
  assign n31025 = n31024 ^ n21145 ^ 1'b0 ;
  assign n31026 = n29511 ^ n6989 ^ n5542 ;
  assign n31027 = n15492 & n18028 ;
  assign n31028 = n28116 ^ n19110 ^ 1'b0 ;
  assign n31029 = n22485 & ~n31028 ;
  assign n31030 = n754 | n2076 ;
  assign n31031 = n23396 | n25289 ;
  assign n31032 = n31031 ^ n30945 ^ 1'b0 ;
  assign n31033 = n227 | n1635 ;
  assign n31034 = n31033 ^ n8860 ^ 1'b0 ;
  assign n31035 = n955 ^ n279 ^ 1'b0 ;
  assign n31036 = n14393 ^ n1112 ^ 1'b0 ;
  assign n31037 = ~n24366 & n31036 ;
  assign n31038 = n31037 ^ n5725 ^ 1'b0 ;
  assign n31039 = n2431 & n31038 ;
  assign n31041 = n2655 ^ n2092 ^ 1'b0 ;
  assign n31040 = ~n1337 & n3799 ;
  assign n31042 = n31041 ^ n31040 ^ 1'b0 ;
  assign n31043 = n11980 | n25670 ;
  assign n31044 = n86 | n9627 ;
  assign n31045 = n22908 ^ n15717 ^ 1'b0 ;
  assign n31046 = n31045 ^ n13820 ^ 1'b0 ;
  assign n31047 = n4419 & ~n7480 ;
  assign n31048 = n567 & n31047 ;
  assign n31049 = n20214 & n20529 ;
  assign n31050 = ~n3186 & n3794 ;
  assign n31051 = n31050 ^ n2689 ^ 1'b0 ;
  assign n31052 = n5724 & n31051 ;
  assign n31053 = n31052 ^ n3287 ^ 1'b0 ;
  assign n31054 = ~n3359 & n29863 ;
  assign n31055 = n31054 ^ n26746 ^ 1'b0 ;
  assign n31056 = n26890 & n28055 ;
  assign n31057 = n31056 ^ n25865 ^ 1'b0 ;
  assign n31058 = n3583 & ~n31057 ;
  assign n31059 = n16882 ^ n470 ^ 1'b0 ;
  assign n31060 = n4662 & ~n31059 ;
  assign n31061 = n31060 ^ n2460 ^ 1'b0 ;
  assign n31062 = n31061 ^ n4319 ^ 1'b0 ;
  assign n31063 = n9399 | n31062 ;
  assign n31064 = n9603 & n18655 ;
  assign n31065 = n1001 & n13974 ;
  assign n31066 = ~n30 & n17872 ;
  assign n31067 = n9596 | n22579 ;
  assign n31068 = n1439 | n3735 ;
  assign n31069 = n3338 & n31068 ;
  assign n31070 = ~n24404 & n31069 ;
  assign n31071 = n4865 | n31070 ;
  assign n31072 = n11438 & ~n20839 ;
  assign n31073 = n6933 & n29953 ;
  assign n31074 = n4695 & n11053 ;
  assign n31075 = n12223 & n21116 ;
  assign n31076 = n20322 ^ n6166 ^ 1'b0 ;
  assign n31077 = n27844 & ~n28744 ;
  assign n31078 = ~n1197 & n5634 ;
  assign n31079 = n17849 & n31078 ;
  assign n31080 = n616 & ~n31079 ;
  assign n31081 = n31080 ^ n2165 ^ 1'b0 ;
  assign n31082 = ~n3138 & n13782 ;
  assign n31083 = n31081 & n31082 ;
  assign n31084 = n10415 & n22032 ;
  assign n31085 = n31084 ^ n10175 ^ 1'b0 ;
  assign n31086 = n31085 ^ n29079 ^ 1'b0 ;
  assign n31087 = n1560 & ~n2617 ;
  assign n31088 = n31087 ^ n4246 ^ 1'b0 ;
  assign n31089 = ~n3743 & n6822 ;
  assign n31090 = n31089 ^ n18152 ^ 1'b0 ;
  assign n31091 = ~n4815 & n12280 ;
  assign n31092 = n51 & n19789 ;
  assign n31093 = ~n4671 & n10175 ;
  assign n31094 = n12308 | n20263 ;
  assign n31095 = n6281 | n28353 ;
  assign n31096 = n4510 | n11447 ;
  assign n31097 = n10946 & n23357 ;
  assign n31098 = n5484 & ~n31097 ;
  assign n31099 = n16906 ^ n6170 ^ 1'b0 ;
  assign n31100 = n28837 & n31099 ;
  assign n31101 = n5721 & ~n27260 ;
  assign n31102 = n1920 & n27686 ;
  assign n31103 = ~n31101 & n31102 ;
  assign n31104 = n20967 ^ n5625 ^ n3718 ;
  assign n31105 = ~n1067 & n17974 ;
  assign n31106 = n5877 ^ n2604 ^ 1'b0 ;
  assign n31107 = n23506 | n31106 ;
  assign n31108 = n12010 & n18440 ;
  assign n31109 = ( ~n5263 & n31107 ) | ( ~n5263 & n31108 ) | ( n31107 & n31108 ) ;
  assign n31110 = n553 & ~n2873 ;
  assign n31111 = n16758 & n31110 ;
  assign n31112 = n31111 ^ n105 ^ 1'b0 ;
  assign n31113 = n9134 & n31112 ;
  assign n31114 = n7632 ^ n3492 ^ 1'b0 ;
  assign n31115 = n8747 | n31114 ;
  assign n31116 = n19789 & ~n31115 ;
  assign n31117 = ~n2199 & n8619 ;
  assign n31118 = ~n4288 & n28712 ;
  assign n31119 = n14935 | n28806 ;
  assign n31120 = n31118 | n31119 ;
  assign n31121 = n20299 ^ n1003 ^ 1'b0 ;
  assign n31122 = n3928 & ~n31121 ;
  assign n31123 = n31122 ^ n11513 ^ 1'b0 ;
  assign n31124 = ( n4547 & ~n16401 ) | ( n4547 & n20728 ) | ( ~n16401 & n20728 ) ;
  assign n31125 = n2067 & n22857 ;
  assign n31126 = n4281 & n31125 ;
  assign n31127 = n7355 & n11872 ;
  assign n31128 = n8231 ^ n840 ^ 1'b0 ;
  assign n31129 = ~n1744 & n17233 ;
  assign n31130 = n31128 & n31129 ;
  assign n31131 = n31130 ^ n5939 ^ 1'b0 ;
  assign n31132 = n158 & ~n1320 ;
  assign n31133 = n4815 & n31132 ;
  assign n31134 = n6538 & n31133 ;
  assign n31135 = n8856 & ~n13736 ;
  assign n31136 = n6357 & n17645 ;
  assign n31137 = n19687 ^ n1103 ^ 1'b0 ;
  assign n31138 = ~n31136 & n31137 ;
  assign n31139 = n19922 & ~n20517 ;
  assign n31140 = n11483 ^ n1106 ^ 1'b0 ;
  assign n31141 = ~n461 & n31140 ;
  assign n31142 = ~n31139 & n31141 ;
  assign n31143 = n12669 & n31142 ;
  assign n31144 = n30289 ^ n12242 ^ n2973 ;
  assign n31145 = ~n9994 & n19789 ;
  assign n31146 = n24186 & n31145 ;
  assign n31147 = ~n560 & n31146 ;
  assign n31148 = n31147 ^ n11210 ^ 1'b0 ;
  assign n31149 = ~n1652 & n31148 ;
  assign n31150 = ~n18106 & n19055 ;
  assign n31151 = n29103 ^ n6666 ^ n1025 ;
  assign n31153 = n1406 | n17537 ;
  assign n31154 = n31153 ^ n5095 ^ 1'b0 ;
  assign n31152 = n19327 ^ n15048 ^ 1'b0 ;
  assign n31155 = n31154 ^ n31152 ^ 1'b0 ;
  assign n31156 = n785 | n13777 ;
  assign n31157 = n31156 ^ n3154 ^ 1'b0 ;
  assign n31158 = n3980 | n16485 ;
  assign n31159 = n14903 ^ n10676 ^ n4584 ;
  assign n31160 = ~n5663 & n13660 ;
  assign n31161 = ~n31159 & n31160 ;
  assign n31162 = n22373 ^ n19437 ^ 1'b0 ;
  assign n31163 = n7452 & n31162 ;
  assign n31164 = n31163 ^ n1876 ^ 1'b0 ;
  assign n31165 = n1050 & ~n3339 ;
  assign n31166 = n424 ^ n423 ^ n246 ;
  assign n31167 = n31166 ^ n3493 ^ 1'b0 ;
  assign n31168 = n15287 | n17045 ;
  assign n31169 = n31167 & ~n31168 ;
  assign n31170 = n3346 ^ n476 ^ 1'b0 ;
  assign n31171 = n7090 | n31170 ;
  assign n31172 = n11186 | n31171 ;
  assign n31173 = n31172 ^ n19175 ^ 1'b0 ;
  assign n31174 = n21126 ^ n2964 ^ 1'b0 ;
  assign n31175 = n31173 | n31174 ;
  assign n31176 = n7134 & n12967 ;
  assign n31177 = n2439 & ~n2973 ;
  assign n31178 = n465 | n18481 ;
  assign n31179 = n31178 ^ n1833 ^ 1'b0 ;
  assign n31180 = n8002 ^ n5073 ^ 1'b0 ;
  assign n31181 = n1157 ^ n585 ^ 1'b0 ;
  assign n31182 = n31181 ^ n8199 ^ 1'b0 ;
  assign n31183 = n23310 ^ n78 ^ 1'b0 ;
  assign n31184 = n477 | n26484 ;
  assign n31185 = n15074 | n31184 ;
  assign n31186 = n10535 | n15319 ;
  assign n31187 = n10092 & ~n21350 ;
  assign n31188 = ~n3524 & n31187 ;
  assign n31189 = ~n13678 & n21988 ;
  assign n31190 = ~n3697 & n31189 ;
  assign n31191 = n15038 ^ n10534 ^ 1'b0 ;
  assign n31192 = n4291 & ~n22502 ;
  assign n31193 = n31192 ^ n24510 ^ 1'b0 ;
  assign n31194 = n2967 ^ n809 ^ 1'b0 ;
  assign n31195 = ~n5831 & n31194 ;
  assign n31196 = n891 | n24404 ;
  assign n31197 = n4510 & ~n31196 ;
  assign n31198 = n31197 ^ n6673 ^ 1'b0 ;
  assign n31199 = n17714 & n18873 ;
  assign n31200 = n31199 ^ n9536 ^ 1'b0 ;
  assign n31201 = ~n2789 & n3131 ;
  assign n31202 = n20715 & n31201 ;
  assign n31203 = n1555 | n27292 ;
  assign n31204 = n836 & n2316 ;
  assign n31205 = n16164 | n31204 ;
  assign n31206 = n14315 ^ n1081 ^ 1'b0 ;
  assign n31207 = n2554 & ~n31206 ;
  assign n31208 = ~n21013 & n29268 ;
  assign n31209 = n16808 ^ n2553 ^ 1'b0 ;
  assign n31210 = n31209 ^ n28392 ^ 1'b0 ;
  assign n31215 = n2753 & ~n8105 ;
  assign n31211 = n8088 ^ n6558 ^ 1'b0 ;
  assign n31212 = n17889 & ~n31211 ;
  assign n31213 = n5382 & n31212 ;
  assign n31214 = n1821 & ~n31213 ;
  assign n31216 = n31215 ^ n31214 ^ 1'b0 ;
  assign n31217 = n16923 & n22055 ;
  assign n31218 = ( ~n142 & n5102 ) | ( ~n142 & n6091 ) | ( n5102 & n6091 ) ;
  assign n31219 = n6932 ^ n2397 ^ 1'b0 ;
  assign n31220 = n31218 | n31219 ;
  assign n31221 = ( n1139 & ~n14731 ) | ( n1139 & n19002 ) | ( ~n14731 & n19002 ) ;
  assign n31222 = n6222 & n31221 ;
  assign n31223 = n31222 ^ n23624 ^ n318 ;
  assign n31224 = ~n10813 & n18053 ;
  assign n31225 = n13604 ^ n9498 ^ 1'b0 ;
  assign n31226 = n13183 & ~n31225 ;
  assign n31227 = n17886 ^ n4133 ^ 1'b0 ;
  assign n31230 = n24502 & n29882 ;
  assign n31228 = n4987 ^ n281 ^ 1'b0 ;
  assign n31229 = n19095 | n31228 ;
  assign n31231 = n31230 ^ n31229 ^ 1'b0 ;
  assign n31232 = ~n5696 & n10113 ;
  assign n31237 = n8156 ^ n3442 ^ 1'b0 ;
  assign n31234 = n9589 | n18428 ;
  assign n31235 = n31234 ^ n627 ^ 1'b0 ;
  assign n31233 = n2154 & ~n15794 ;
  assign n31236 = n31235 ^ n31233 ^ n17756 ;
  assign n31238 = n31237 ^ n31236 ^ 1'b0 ;
  assign n31239 = n2578 & ~n4824 ;
  assign n31240 = n9139 & n31239 ;
  assign n31241 = n1606 ^ n128 ^ 1'b0 ;
  assign n31242 = n2773 & ~n31241 ;
  assign n31243 = n17315 & ~n31242 ;
  assign n31244 = n22165 | n31243 ;
  assign n31245 = n8106 | n31244 ;
  assign n31246 = ~n2260 & n12550 ;
  assign n31247 = n30009 ^ n15367 ^ 1'b0 ;
  assign n31248 = n11359 | n13093 ;
  assign n31250 = n2589 | n3037 ;
  assign n31251 = n3037 & ~n31250 ;
  assign n31249 = n599 & ~n3378 ;
  assign n31252 = n31251 ^ n31249 ^ 1'b0 ;
  assign n31253 = n2017 & n31252 ;
  assign n31254 = n1227 & ~n31253 ;
  assign n31255 = n5529 & ~n31254 ;
  assign n31256 = n652 | n13856 ;
  assign n31257 = n24999 | n31256 ;
  assign n31258 = n4311 & ~n27965 ;
  assign n31259 = n3387 & n4505 ;
  assign n31260 = n7019 ^ n667 ^ 1'b0 ;
  assign n31261 = n6315 & ~n31260 ;
  assign n31262 = ~n21961 & n31261 ;
  assign n31263 = ~n12063 & n21520 ;
  assign n31264 = n31263 ^ n9583 ^ 1'b0 ;
  assign n31265 = n31264 ^ n594 ^ 1'b0 ;
  assign n31266 = n7810 & ~n31265 ;
  assign n31267 = n86 & ~n27629 ;
  assign n31268 = n3817 ^ n1103 ^ 1'b0 ;
  assign n31269 = n205 & n29863 ;
  assign n31270 = n31269 ^ n10261 ^ 1'b0 ;
  assign n31272 = n10033 ^ n697 ^ 1'b0 ;
  assign n31271 = n9179 & ~n9273 ;
  assign n31273 = n31272 ^ n31271 ^ 1'b0 ;
  assign n31274 = n10923 | n31273 ;
  assign n31275 = n22282 | n31274 ;
  assign n31276 = ~n1867 & n31275 ;
  assign n31277 = n31276 ^ n7767 ^ 1'b0 ;
  assign n31278 = ~n16122 & n16445 ;
  assign n31279 = n8829 & ~n31278 ;
  assign n31280 = n4396 | n6951 ;
  assign n31281 = n31280 ^ n865 ^ 1'b0 ;
  assign n31282 = n16505 | n26634 ;
  assign n31283 = n20951 ^ n1366 ^ n1197 ;
  assign n31284 = n19527 | n20013 ;
  assign n31285 = ~n8121 & n17827 ;
  assign n31286 = n31285 ^ n16753 ^ 1'b0 ;
  assign n31287 = ~n9239 & n9435 ;
  assign n31288 = n12961 ^ n10625 ^ 1'b0 ;
  assign n31289 = n31287 & ~n31288 ;
  assign n31290 = n10831 ^ n837 ^ 1'b0 ;
  assign n31291 = ~n20527 & n31290 ;
  assign n31292 = ~n4253 & n5345 ;
  assign n31293 = n31292 ^ n10541 ^ n9408 ;
  assign n31294 = n1441 & ~n31293 ;
  assign n31295 = n31294 ^ n14830 ^ 1'b0 ;
  assign n31296 = n17238 ^ n114 ^ 1'b0 ;
  assign n31297 = ( n11462 & ~n22335 ) | ( n11462 & n31296 ) | ( ~n22335 & n31296 ) ;
  assign n31298 = n9623 | n21005 ;
  assign n31299 = n18746 ^ n10950 ^ 1'b0 ;
  assign n31300 = n1441 ^ n866 ^ 1'b0 ;
  assign n31301 = n288 & n31300 ;
  assign n31302 = n2509 | n8281 ;
  assign n31303 = n1396 & n18778 ;
  assign n31304 = ( n31301 & n31302 ) | ( n31301 & ~n31303 ) | ( n31302 & ~n31303 ) ;
  assign n31305 = n18300 ^ n16800 ^ 1'b0 ;
  assign n31306 = n12373 & ~n31305 ;
  assign n31307 = n7289 ^ n3804 ^ 1'b0 ;
  assign n31308 = n29986 & ~n31307 ;
  assign n31309 = n31308 ^ n24582 ^ 1'b0 ;
  assign n31310 = n6758 ^ n5749 ^ 1'b0 ;
  assign n31311 = ~n17519 & n31310 ;
  assign n31312 = n7927 & n31311 ;
  assign n31313 = n9439 | n31312 ;
  assign n31314 = n1851 | n16309 ;
  assign n31315 = n31314 ^ n3370 ^ 1'b0 ;
  assign n31316 = n4415 & ~n9221 ;
  assign n31317 = ~x0 & n1425 ;
  assign n31318 = n31317 ^ n9588 ^ 1'b0 ;
  assign n31319 = n1763 & ~n4176 ;
  assign n31320 = n31318 & n31319 ;
  assign n31321 = n31320 ^ n2624 ^ 1'b0 ;
  assign n31322 = n31321 ^ n1329 ^ 1'b0 ;
  assign n31323 = n4666 ^ n114 ^ 1'b0 ;
  assign n31324 = n14452 | n31323 ;
  assign n31325 = n9223 & ~n30978 ;
  assign n31326 = n8472 ^ n6098 ^ n1048 ;
  assign n31327 = ~n207 & n14865 ;
  assign n31328 = n28083 | n31327 ;
  assign n31329 = n31328 ^ n18966 ^ 1'b0 ;
  assign n31330 = n832 & n6536 ;
  assign n31331 = n3779 & ~n15419 ;
  assign n31332 = n31331 ^ n10882 ^ 1'b0 ;
  assign n31333 = n3844 & n7981 ;
  assign n31334 = n31333 ^ n6927 ^ 1'b0 ;
  assign n31335 = n19970 ^ n137 ^ 1'b0 ;
  assign n31336 = n20951 | n31335 ;
  assign n31337 = n1777 & n4334 ;
  assign n31338 = n31337 ^ n4801 ^ 1'b0 ;
  assign n31339 = n13569 | n31338 ;
  assign n31340 = n4060 & n8362 ;
  assign n31341 = n4057 | n4263 ;
  assign n31342 = n8360 | n31341 ;
  assign n31343 = n31340 | n31342 ;
  assign n31344 = n1178 & n7983 ;
  assign n31345 = n348 & ~n6531 ;
  assign n31346 = ~n3732 & n17021 ;
  assign n31347 = n4580 | n10246 ;
  assign n31348 = n4652 | n31347 ;
  assign n31349 = n23274 ^ n758 ^ 1'b0 ;
  assign n31350 = n2072 & ~n16996 ;
  assign n31351 = n23942 | n30798 ;
  assign n31352 = ~n5978 & n9667 ;
  assign n31353 = n1505 & ~n15821 ;
  assign n31354 = n25751 ^ n2260 ^ 1'b0 ;
  assign n31357 = n7277 & n27424 ;
  assign n31358 = n6054 & n31357 ;
  assign n31355 = n24046 ^ n1795 ^ 1'b0 ;
  assign n31356 = n10033 & n31355 ;
  assign n31359 = n31358 ^ n31356 ^ 1'b0 ;
  assign n31360 = n11733 ^ n4048 ^ 1'b0 ;
  assign n31361 = ~n2304 & n31360 ;
  assign n31362 = n9791 ^ n8014 ^ 1'b0 ;
  assign n31363 = n31362 ^ n11493 ^ 1'b0 ;
  assign n31364 = n31361 & n31363 ;
  assign n31365 = n4918 ^ n3452 ^ 1'b0 ;
  assign n31366 = ~n259 & n31365 ;
  assign n31367 = n594 & n27412 ;
  assign n31368 = n31367 ^ n3718 ^ 1'b0 ;
  assign n31369 = n18899 ^ n1697 ^ 1'b0 ;
  assign n31370 = n5559 | n17815 ;
  assign n31371 = n28732 & ~n31370 ;
  assign n31372 = n1202 & ~n2945 ;
  assign n31373 = n23621 ^ n6846 ^ 1'b0 ;
  assign n31374 = ~n12495 & n13954 ;
  assign n31375 = n31374 ^ n2258 ^ 1'b0 ;
  assign n31376 = ~n3732 & n31375 ;
  assign n31377 = n31376 ^ n28535 ^ 1'b0 ;
  assign n31378 = n6333 | n31377 ;
  assign n31379 = n25990 ^ n5445 ^ 1'b0 ;
  assign n31380 = ~n6484 & n14160 ;
  assign n31381 = n18528 & n31380 ;
  assign n31382 = n2001 & ~n15678 ;
  assign n31383 = n3061 | n4636 ;
  assign n31384 = n31383 ^ n2318 ^ 1'b0 ;
  assign n31385 = n17025 ^ n713 ^ 1'b0 ;
  assign n31386 = n5140 | n31385 ;
  assign n31387 = n2904 ^ n279 ^ 1'b0 ;
  assign n31388 = ~n20269 & n31387 ;
  assign n31389 = ~n5445 & n13449 ;
  assign n31390 = n1681 & n13890 ;
  assign n31391 = ~n1681 & n31390 ;
  assign n31396 = ~n556 & n1834 ;
  assign n31397 = n556 & n31396 ;
  assign n31398 = n1785 | n2260 ;
  assign n31399 = n2260 & ~n31398 ;
  assign n31400 = n31397 & ~n31399 ;
  assign n31392 = n4440 & n5826 ;
  assign n31393 = ~n4440 & n31392 ;
  assign n31394 = n15879 ^ n5367 ^ 1'b0 ;
  assign n31395 = n31393 | n31394 ;
  assign n31401 = n31400 ^ n31395 ^ 1'b0 ;
  assign n31402 = n31391 | n31401 ;
  assign n31403 = n10676 ^ n820 ^ 1'b0 ;
  assign n31404 = ~n16029 & n31403 ;
  assign n31405 = n12019 ^ n832 ^ 1'b0 ;
  assign n31406 = ~n7654 & n18746 ;
  assign n31408 = n13442 ^ n1429 ^ 1'b0 ;
  assign n31409 = n306 & ~n31408 ;
  assign n31407 = n7569 | n8711 ;
  assign n31410 = n31409 ^ n31407 ^ 1'b0 ;
  assign n31411 = n278 | n19862 ;
  assign n31412 = n6091 & ~n31411 ;
  assign n31413 = n13196 & ~n31412 ;
  assign n31414 = n31413 ^ n15054 ^ 1'b0 ;
  assign n31415 = n10816 & n14472 ;
  assign n31416 = n21552 & ~n21994 ;
  assign n31417 = n3693 & n31416 ;
  assign n31418 = n2339 & ~n4680 ;
  assign n31419 = n20796 & ~n31418 ;
  assign n31420 = n13943 ^ n389 ^ 1'b0 ;
  assign n31422 = n8172 | n9197 ;
  assign n31423 = n412 | n31422 ;
  assign n31421 = n12184 ^ n8939 ^ 1'b0 ;
  assign n31424 = n31423 ^ n31421 ^ n12053 ;
  assign n31425 = n22886 ^ n3900 ^ 1'b0 ;
  assign n31426 = n31425 ^ n12502 ^ n12205 ;
  assign n31427 = n7805 | n31426 ;
  assign n31428 = n12918 ^ n962 ^ 1'b0 ;
  assign n31429 = ~n10976 & n31428 ;
  assign n31430 = n16158 & ~n28324 ;
  assign n31431 = n12193 ^ n2063 ^ 1'b0 ;
  assign n31432 = n412 & n5495 ;
  assign n31433 = n3649 ^ n1934 ^ 1'b0 ;
  assign n31434 = ( n1355 & ~n21616 ) | ( n1355 & n31433 ) | ( ~n21616 & n31433 ) ;
  assign n31435 = n31434 ^ n23183 ^ 1'b0 ;
  assign n31436 = n31432 & ~n31435 ;
  assign n31437 = n2380 | n6417 ;
  assign n31438 = n24256 | n31437 ;
  assign n31439 = n22583 ^ n6911 ^ 1'b0 ;
  assign n31440 = n25291 & n31439 ;
  assign n31441 = n6950 | n31440 ;
  assign n31442 = ~n17263 & n22721 ;
  assign n31443 = n31442 ^ n4004 ^ 1'b0 ;
  assign n31444 = n835 | n4565 ;
  assign n31445 = n6810 & n31444 ;
  assign n31446 = n31445 ^ n4217 ^ 1'b0 ;
  assign n31447 = n13650 | n31446 ;
  assign n31448 = n27414 & ~n31447 ;
  assign n31449 = n24722 ^ n23198 ^ 1'b0 ;
  assign n31450 = ~n340 & n15902 ;
  assign n31451 = n2547 & ~n31450 ;
  assign n31452 = n26083 ^ n2792 ^ 1'b0 ;
  assign n31453 = ~n10878 & n22693 ;
  assign n31454 = n9206 ^ n7612 ^ n44 ;
  assign n31455 = n7669 & ~n31454 ;
  assign n31456 = n2664 & n14054 ;
  assign n31457 = n857 & ~n2766 ;
  assign n31458 = n16706 & ~n31457 ;
  assign n31459 = n31458 ^ n6011 ^ 1'b0 ;
  assign n31460 = n6945 | n31459 ;
  assign n31461 = n2500 & ~n29466 ;
  assign n31462 = n16645 ^ n12777 ^ 1'b0 ;
  assign n31463 = ~n14316 & n31462 ;
  assign n31464 = n6558 ^ n364 ^ 1'b0 ;
  assign n31465 = n2662 ^ n1854 ^ 1'b0 ;
  assign n31466 = ~n25352 & n31465 ;
  assign n31467 = ~n12388 & n31466 ;
  assign n31468 = n6611 ^ n2485 ^ 1'b0 ;
  assign n31469 = n809 | n10282 ;
  assign n31470 = ~n628 & n6166 ;
  assign n31471 = n31470 ^ n24439 ^ 1'b0 ;
  assign n31472 = ~n1368 & n31471 ;
  assign n31473 = n19759 | n31472 ;
  assign n31475 = ~n7706 & n8718 ;
  assign n31474 = n2633 | n2769 ;
  assign n31476 = n31475 ^ n31474 ^ 1'b0 ;
  assign n31477 = n6729 & ~n31476 ;
  assign n31478 = n17508 ^ n10476 ^ 1'b0 ;
  assign n31479 = n7943 | n31478 ;
  assign n31480 = n233 & ~n16269 ;
  assign n31481 = n30924 & n31480 ;
  assign n31482 = ~n15553 & n25267 ;
  assign n31483 = n8689 | n12316 ;
  assign n31484 = n2410 ^ n253 ^ 1'b0 ;
  assign n31485 = n7806 & ~n7821 ;
  assign n31486 = n31484 & n31485 ;
  assign n31487 = n10621 ^ n4374 ^ 1'b0 ;
  assign n31488 = n9443 & n31487 ;
  assign n31489 = ~n13070 & n22120 ;
  assign n31490 = n31489 ^ n4640 ^ 1'b0 ;
  assign n31491 = n31488 | n31490 ;
  assign n31492 = ( n1309 & n1896 ) | ( n1309 & n2941 ) | ( n1896 & n2941 ) ;
  assign n31493 = n7401 & ~n31492 ;
  assign n31494 = n31493 ^ n9060 ^ 1'b0 ;
  assign n31495 = n4649 & n31494 ;
  assign n31496 = n11539 ^ n5517 ^ 1'b0 ;
  assign n31497 = n719 | n2440 ;
  assign n31498 = n50 & n19113 ;
  assign n31499 = n5609 & n6618 ;
  assign n31500 = n323 & n10367 ;
  assign n31501 = ~n9180 & n31500 ;
  assign n31502 = n673 & n31501 ;
  assign n31503 = n14235 ^ n9263 ^ 1'b0 ;
  assign n31504 = n4763 & n31503 ;
  assign n31505 = n5094 | n31504 ;
  assign n31506 = n512 & n6957 ;
  assign n31507 = n9599 & n31506 ;
  assign n31508 = ~n19535 & n31507 ;
  assign n31509 = ~n1138 & n11904 ;
  assign n31510 = n3738 & n9014 ;
  assign n31511 = n1444 | n4407 ;
  assign n31512 = n6622 & n22494 ;
  assign n31513 = n25125 ^ n12951 ^ 1'b0 ;
  assign n31514 = n4015 ^ n2978 ^ 1'b0 ;
  assign n31515 = n31513 | n31514 ;
  assign n31516 = n31515 ^ n10589 ^ 1'b0 ;
  assign n31517 = n6278 & n31516 ;
  assign n31518 = n3028 ^ n566 ^ 1'b0 ;
  assign n31519 = ~n4439 & n14884 ;
  assign n31520 = x1 & n22096 ;
  assign n31521 = ~n4893 & n31520 ;
  assign n31522 = ~n9666 & n31521 ;
  assign n31523 = n12118 ^ n4976 ^ 1'b0 ;
  assign n31524 = n11105 & n23030 ;
  assign n31525 = n7476 | n12412 ;
  assign n31526 = n31524 & ~n31525 ;
  assign n31527 = n14601 ^ n2585 ^ 1'b0 ;
  assign n31528 = n31527 ^ n16779 ^ 1'b0 ;
  assign n31529 = ( n5155 & ~n10117 ) | ( n5155 & n15012 ) | ( ~n10117 & n15012 ) ;
  assign n31530 = n25131 ^ n970 ^ 1'b0 ;
  assign n31531 = n847 | n31530 ;
  assign n31532 = n8271 & ~n31531 ;
  assign n31533 = n475 | n2553 ;
  assign n31534 = n31533 ^ n4473 ^ 1'b0 ;
  assign n31535 = n2141 | n30059 ;
  assign n31536 = n31535 ^ n5304 ^ 1'b0 ;
  assign n31537 = n31534 & n31536 ;
  assign n31538 = n9242 & ~n10427 ;
  assign n31539 = ~n31537 & n31538 ;
  assign n31540 = n15623 ^ n3803 ^ 1'b0 ;
  assign n31541 = ~n901 & n17026 ;
  assign n31542 = n1516 & ~n31541 ;
  assign n31543 = n9817 ^ n5856 ^ 1'b0 ;
  assign n31544 = n6849 & n16995 ;
  assign n31545 = n31544 ^ n7907 ^ 1'b0 ;
  assign n31546 = n4196 | n20847 ;
  assign n31547 = n17867 & ~n31546 ;
  assign n31548 = n31547 ^ n30529 ^ 1'b0 ;
  assign n31549 = n16940 ^ n14225 ^ 1'b0 ;
  assign n31550 = n31548 & n31549 ;
  assign n31551 = n4373 ^ n3451 ^ n1602 ;
  assign n31552 = n4660 | n19959 ;
  assign n31553 = n31552 ^ n9659 ^ 1'b0 ;
  assign n31554 = n31553 ^ n10333 ^ 1'b0 ;
  assign n31555 = n27587 | n31554 ;
  assign n31556 = n3225 | n25315 ;
  assign n31557 = ~n3434 & n31556 ;
  assign n31558 = n2136 | n28270 ;
  assign n31559 = n7231 ^ n2595 ^ 1'b0 ;
  assign n31560 = n18326 & ~n31559 ;
  assign n31561 = ~n4879 & n18542 ;
  assign n31562 = n31561 ^ n10644 ^ 1'b0 ;
  assign n31563 = n10423 ^ n1460 ^ 1'b0 ;
  assign n31564 = ~n3845 & n11716 ;
  assign n31565 = n77 | n31564 ;
  assign n31566 = n31565 ^ n17094 ^ 1'b0 ;
  assign n31567 = ~n31563 & n31566 ;
  assign n31568 = n3120 & ~n12477 ;
  assign n31571 = n2436 ^ n1872 ^ 1'b0 ;
  assign n31570 = n2068 & ~n5187 ;
  assign n31572 = n31571 ^ n31570 ^ 1'b0 ;
  assign n31569 = n25634 ^ n23043 ^ 1'b0 ;
  assign n31573 = n31572 ^ n31569 ^ 1'b0 ;
  assign n31574 = n18606 ^ n16025 ^ 1'b0 ;
  assign n31575 = n31574 ^ n26088 ^ 1'b0 ;
  assign n31576 = ~n7704 & n31575 ;
  assign n31577 = n30459 ^ n9364 ^ 1'b0 ;
  assign n31578 = ~n13352 & n17146 ;
  assign n31579 = n14193 & n31578 ;
  assign n31600 = n11232 & n18949 ;
  assign n31601 = ~n11232 & n31600 ;
  assign n31580 = ~n378 & n1064 ;
  assign n31581 = n378 & n31580 ;
  assign n31582 = ~n20160 & n30362 ;
  assign n31583 = n24744 ^ n715 ^ 1'b0 ;
  assign n31584 = n31582 & ~n31583 ;
  assign n31585 = n468 | n17404 ;
  assign n31586 = n31584 & ~n31585 ;
  assign n31587 = n31581 & n31586 ;
  assign n31588 = n227 | n403 ;
  assign n31589 = n227 & ~n31588 ;
  assign n31590 = n31589 ^ n862 ^ 1'b0 ;
  assign n31591 = ~n158 & n238 ;
  assign n31592 = ~n238 & n31591 ;
  assign n31593 = n1744 & ~n31592 ;
  assign n31594 = ~n1744 & n31593 ;
  assign n31595 = n31590 & ~n31594 ;
  assign n31596 = ~n31590 & n31595 ;
  assign n31597 = n3100 & ~n31596 ;
  assign n31598 = ~n3100 & n31597 ;
  assign n31599 = n31587 | n31598 ;
  assign n31602 = n31601 ^ n31599 ^ 1'b0 ;
  assign n31603 = n31602 ^ n23559 ^ n21277 ;
  assign n31604 = n25262 ^ n10255 ^ 1'b0 ;
  assign n31605 = ( n4867 & ~n7217 ) | ( n4867 & n16548 ) | ( ~n7217 & n16548 ) ;
  assign n31606 = n18624 & ~n31605 ;
  assign n31607 = ~n27606 & n31606 ;
  assign n31608 = n16660 ^ n227 ^ 1'b0 ;
  assign n31609 = n28154 & n31608 ;
  assign n31610 = n14727 & ~n17683 ;
  assign n31611 = n7188 & n31610 ;
  assign n31612 = n4642 & ~n31611 ;
  assign n31613 = n542 & ~n19579 ;
  assign n31614 = n31613 ^ n24615 ^ 1'b0 ;
  assign n31615 = n27976 ^ n1650 ^ 1'b0 ;
  assign n31616 = ~n3127 & n31615 ;
  assign n31617 = n5498 | n13727 ;
  assign n31618 = n21373 & ~n31617 ;
  assign n31619 = n13150 & n31618 ;
  assign n31620 = ~n4396 & n19715 ;
  assign n31621 = n26435 & n31620 ;
  assign n31622 = n21604 ^ n7954 ^ 1'b0 ;
  assign n31623 = n31621 | n31622 ;
  assign n31624 = n11235 | n27464 ;
  assign n31625 = n3446 | n3452 ;
  assign n31626 = n31624 & ~n31625 ;
  assign n31627 = n12777 | n15299 ;
  assign n31628 = n2260 | n5827 ;
  assign n31629 = n4034 & n11608 ;
  assign n31630 = ~n3221 & n31629 ;
  assign n31631 = n30844 ^ n22940 ^ 1'b0 ;
  assign n31632 = n31630 & n31631 ;
  assign n31633 = n258 & n4787 ;
  assign n31634 = n4211 & ~n4660 ;
  assign n31635 = n31634 ^ n1372 ^ 1'b0 ;
  assign n31636 = n26727 & n31635 ;
  assign n31637 = n4784 | n31636 ;
  assign n31638 = n1559 | n31637 ;
  assign n31639 = n15605 ^ n13398 ^ 1'b0 ;
  assign n31640 = n11111 & n13357 ;
  assign n31641 = n15614 ^ n6246 ^ 1'b0 ;
  assign n31642 = n19015 ^ n2686 ^ 1'b0 ;
  assign n31643 = n2403 & ~n31642 ;
  assign n31644 = n18538 & ~n31643 ;
  assign n31646 = n16653 ^ n1388 ^ 1'b0 ;
  assign n31647 = n619 & ~n31646 ;
  assign n31645 = n8219 & ~n12291 ;
  assign n31648 = n31647 ^ n31645 ^ 1'b0 ;
  assign n31649 = ~n7915 & n10315 ;
  assign n31650 = n5813 & ~n31649 ;
  assign n31651 = n31650 ^ n849 ^ 1'b0 ;
  assign n31652 = n29941 ^ n374 ^ 1'b0 ;
  assign n31653 = n715 & n4228 ;
  assign n31654 = n10337 ^ n8559 ^ 1'b0 ;
  assign n31655 = ~n16459 & n31654 ;
  assign n31656 = n5677 | n9654 ;
  assign n31657 = n31655 & ~n31656 ;
  assign n31658 = n31657 ^ n29237 ^ 1'b0 ;
  assign n31659 = n8818 & n31658 ;
  assign n31660 = n8994 | n11797 ;
  assign n31661 = n16251 | n31660 ;
  assign n31662 = ~n3368 & n31661 ;
  assign n31663 = n12457 ^ n4367 ^ 1'b0 ;
  assign n31667 = n5024 ^ n1005 ^ 1'b0 ;
  assign n31668 = ~n3408 & n31667 ;
  assign n31664 = n5218 & n29272 ;
  assign n31665 = n31664 ^ n26110 ^ 1'b0 ;
  assign n31666 = n6196 | n31665 ;
  assign n31669 = n31668 ^ n31666 ^ 1'b0 ;
  assign n31670 = n2373 & n23014 ;
  assign n31671 = n10553 | n31670 ;
  assign n31672 = n235 & n21379 ;
  assign n31673 = n17247 & n31672 ;
  assign n31674 = n7311 & n17122 ;
  assign n31675 = n3509 | n12714 ;
  assign n31676 = n31675 ^ n25966 ^ 1'b0 ;
  assign n31677 = ~n10708 & n29563 ;
  assign n31679 = n30048 ^ n638 ^ 1'b0 ;
  assign n31678 = n1060 | n12512 ;
  assign n31680 = n31679 ^ n31678 ^ 1'b0 ;
  assign n31681 = n3333 & n6191 ;
  assign n31682 = ~n13085 & n31681 ;
  assign n31683 = ~n5076 & n24024 ;
  assign n31684 = ( n5796 & n5867 ) | ( n5796 & n11254 ) | ( n5867 & n11254 ) ;
  assign n31685 = n25 | n6322 ;
  assign n31686 = n31684 & ~n31685 ;
  assign n31687 = n31686 ^ n12252 ^ 1'b0 ;
  assign n31689 = ~n8611 & n17506 ;
  assign n31690 = n30462 & n31689 ;
  assign n31688 = n2228 & n20662 ;
  assign n31691 = n31690 ^ n31688 ^ 1'b0 ;
  assign n31692 = n16322 | n25780 ;
  assign n31693 = n3557 & n19364 ;
  assign n31694 = n3896 ^ n1325 ^ 1'b0 ;
  assign n31695 = ~n31693 & n31694 ;
  assign n31696 = n25000 & ~n31695 ;
  assign n31697 = n11115 & ~n13592 ;
  assign n31698 = n31697 ^ n7203 ^ 1'b0 ;
  assign n31699 = n25094 & ~n31698 ;
  assign n31700 = n13954 & ~n31699 ;
  assign n31701 = n200 | n10705 ;
  assign n31702 = ~n715 & n31701 ;
  assign n31703 = n715 | n12689 ;
  assign n31704 = n18091 ^ n738 ^ 1'b0 ;
  assign n31705 = n21737 & ~n31184 ;
  assign n31706 = n6849 ^ n5551 ^ 1'b0 ;
  assign n31707 = n31706 ^ n23377 ^ 1'b0 ;
  assign n31708 = n18214 & n31707 ;
  assign n31709 = n879 & n12747 ;
  assign n31710 = n6249 & n23145 ;
  assign n31711 = n31710 ^ n25868 ^ 1'b0 ;
  assign n31712 = n18525 ^ n5280 ^ 1'b0 ;
  assign n31713 = n6414 ^ n354 ^ 1'b0 ;
  assign n31715 = n11064 ^ n9114 ^ 1'b0 ;
  assign n31714 = ~n4885 & n27227 ;
  assign n31716 = n31715 ^ n31714 ^ 1'b0 ;
  assign n31717 = ~n2723 & n12741 ;
  assign n31718 = ( ~n14438 & n24097 ) | ( ~n14438 & n29216 ) | ( n24097 & n29216 ) ;
  assign n31719 = n2814 | n14566 ;
  assign n31720 = n31719 ^ n1668 ^ 1'b0 ;
  assign n31721 = n2686 ^ n34 ^ 1'b0 ;
  assign n31722 = n31720 & ~n31721 ;
  assign n31723 = n15614 | n31722 ;
  assign n31724 = n25053 ^ n18173 ^ 1'b0 ;
  assign n31725 = n30863 | n31724 ;
  assign n31726 = n31725 ^ n20797 ^ 1'b0 ;
  assign n31727 = ~n5666 & n8990 ;
  assign n31728 = n23155 & n31727 ;
  assign n31729 = ~n17564 & n31728 ;
  assign n31730 = n17546 & n31729 ;
  assign n31731 = n11218 & n24077 ;
  assign n31732 = n31731 ^ n24279 ^ 1'b0 ;
  assign n31733 = n9841 ^ n2358 ^ 1'b0 ;
  assign n31734 = n2733 & n31733 ;
  assign n31735 = n5979 ^ n2751 ^ 1'b0 ;
  assign n31736 = n7307 & n31735 ;
  assign n31737 = n6618 & n31736 ;
  assign n31738 = n621 & n16660 ;
  assign n31739 = ~n19799 & n31738 ;
  assign n31740 = n23038 ^ n18004 ^ 1'b0 ;
  assign n31741 = ~n18975 & n19868 ;
  assign n31742 = n12225 & n31741 ;
  assign n31743 = n19475 | n27928 ;
  assign n31744 = n31743 ^ n12396 ^ 1'b0 ;
  assign n31745 = n10927 & ~n31744 ;
  assign n31746 = n13586 ^ n9304 ^ 1'b0 ;
  assign n31747 = n5540 ^ n3050 ^ 1'b0 ;
  assign n31748 = n2414 ^ n1233 ^ n726 ;
  assign n31749 = n22527 ^ n6543 ^ 1'b0 ;
  assign n31750 = n532 | n13948 ;
  assign n31751 = n8122 | n9009 ;
  assign n31752 = n31750 & ~n31751 ;
  assign n31753 = n6510 & ~n31752 ;
  assign n31754 = n8715 | n23843 ;
  assign n31755 = n31754 ^ n3880 ^ 1'b0 ;
  assign n31757 = n9199 ^ n602 ^ 1'b0 ;
  assign n31758 = n7311 & n31757 ;
  assign n31756 = n2337 & n22145 ;
  assign n31759 = n31758 ^ n31756 ^ 1'b0 ;
  assign n31760 = n16521 ^ n10719 ^ 1'b0 ;
  assign n31761 = n773 & n14949 ;
  assign n31762 = n13113 ^ n4807 ^ 1'b0 ;
  assign n31763 = n4193 & n31762 ;
  assign n31764 = n20875 | n31763 ;
  assign n31765 = n6927 & ~n30807 ;
  assign n31766 = n21959 & n31765 ;
  assign n31767 = n5397 | n31766 ;
  assign n31768 = n21735 | n31767 ;
  assign n31769 = n7288 & ~n25456 ;
  assign n31770 = n8583 & n31769 ;
  assign n31771 = n8813 ^ n8767 ^ 1'b0 ;
  assign n31772 = n4045 & ~n31771 ;
  assign n31773 = ~n2099 & n19390 ;
  assign n31774 = n10984 & ~n26405 ;
  assign n31777 = n774 & ~n2400 ;
  assign n31778 = n31777 ^ n14258 ^ 1'b0 ;
  assign n31779 = ( ~n782 & n1740 ) | ( ~n782 & n31778 ) | ( n1740 & n31778 ) ;
  assign n31780 = ~n345 & n6067 ;
  assign n31781 = ~n31779 & n31780 ;
  assign n31775 = n5914 & n9381 ;
  assign n31776 = n6746 & n31775 ;
  assign n31782 = n31781 ^ n31776 ^ 1'b0 ;
  assign n31783 = ~n21124 & n25990 ;
  assign n31784 = n16504 & n31783 ;
  assign n31785 = n19941 & n31784 ;
  assign n31786 = n2078 & n23171 ;
  assign n31787 = n1693 & n31786 ;
  assign n31788 = n31787 ^ n4404 ^ 1'b0 ;
  assign n31789 = n958 & n18097 ;
  assign n31790 = n26362 ^ n13883 ^ 1'b0 ;
  assign n31791 = ~n6944 & n14355 ;
  assign n31792 = ~n31790 & n31791 ;
  assign n31793 = n2680 | n18372 ;
  assign n31794 = n483 & ~n7088 ;
  assign n31795 = ( n18096 & n29290 ) | ( n18096 & ~n31794 ) | ( n29290 & ~n31794 ) ;
  assign n31796 = n31793 & ~n31795 ;
  assign n31797 = ~n1110 & n18826 ;
  assign n31798 = n3793 ^ n183 ^ 1'b0 ;
  assign n31799 = ~n4264 & n9137 ;
  assign n31800 = n31799 ^ n2780 ^ 1'b0 ;
  assign n31801 = n3827 & n4274 ;
  assign n31802 = n2982 | n14865 ;
  assign n31803 = n31801 & n31802 ;
  assign n31804 = n31800 & ~n31803 ;
  assign n31805 = n4703 & n22546 ;
  assign n31806 = n1602 & ~n22193 ;
  assign n31807 = n3277 & n16251 ;
  assign n31808 = ( n12724 & n24165 ) | ( n12724 & n29448 ) | ( n24165 & n29448 ) ;
  assign n31809 = n1473 | n19304 ;
  assign n31810 = n9736 | n31809 ;
  assign n31811 = n627 & n31810 ;
  assign n31812 = n31811 ^ n6284 ^ 1'b0 ;
  assign n31813 = ~n17999 & n31812 ;
  assign n31815 = n10599 & ~n22504 ;
  assign n31816 = n29586 & n31815 ;
  assign n31817 = n31816 ^ n1112 ^ 1'b0 ;
  assign n31814 = n213 | n7353 ;
  assign n31818 = n31817 ^ n31814 ^ 1'b0 ;
  assign n31820 = ~n1472 & n1769 ;
  assign n31819 = ~n227 & n2331 ;
  assign n31821 = n31820 ^ n31819 ^ 1'b0 ;
  assign n31822 = n21078 & n28753 ;
  assign n31823 = n10607 & ~n13997 ;
  assign n31824 = ~n12232 & n31823 ;
  assign n31825 = n31824 ^ n27128 ^ 1'b0 ;
  assign n31826 = n20252 & n31825 ;
  assign n31827 = n16926 | n22719 ;
  assign n31828 = n31826 | n31827 ;
  assign n31829 = n2260 | n7500 ;
  assign n31830 = n8156 ^ n5269 ^ 1'b0 ;
  assign n31831 = n29366 ^ n4623 ^ 1'b0 ;
  assign n31832 = ~n25131 & n31831 ;
  assign n31833 = n1463 & n16359 ;
  assign n31834 = n31833 ^ n5293 ^ 1'b0 ;
  assign n31835 = n21771 ^ n13911 ^ 1'b0 ;
  assign n31836 = ~n5101 & n31835 ;
  assign n31837 = ~n1038 & n4949 ;
  assign n31838 = ~n1256 & n31837 ;
  assign n31839 = n12310 | n21597 ;
  assign n31840 = n517 & n1791 ;
  assign n31841 = n14926 ^ n8767 ^ 1'b0 ;
  assign n31842 = ~n148 & n31841 ;
  assign n31843 = n593 & ~n16010 ;
  assign n31844 = n31843 ^ n22533 ^ 1'b0 ;
  assign n31845 = n28051 ^ n1303 ^ 1'b0 ;
  assign n31846 = ~n13590 & n31845 ;
  assign n31847 = n25569 ^ n4788 ^ 1'b0 ;
  assign n31848 = n29239 & n31847 ;
  assign n31849 = n16199 & n19550 ;
  assign n31850 = n31849 ^ n24924 ^ n1229 ;
  assign n31851 = n31436 ^ n13949 ^ 1'b0 ;
  assign n31852 = ~n16053 & n31851 ;
  assign n31853 = n12677 & ~n27861 ;
  assign n31854 = n1815 & n6655 ;
  assign n31855 = n31854 ^ n20517 ^ 1'b0 ;
  assign n31856 = n10347 & n19196 ;
  assign n31857 = n31856 ^ n3194 ^ 1'b0 ;
  assign n31858 = ~n18120 & n31857 ;
  assign n31859 = n31858 ^ n4429 ^ 1'b0 ;
  assign n31860 = n10535 ^ n2547 ^ 1'b0 ;
  assign n31861 = ~n512 & n14676 ;
  assign n31862 = n31861 ^ n619 ^ 1'b0 ;
  assign n31863 = n2027 & ~n31862 ;
  assign n31864 = n83 & n151 ;
  assign n31865 = n83 & ~n31864 ;
  assign n31866 = ~n279 & n2883 ;
  assign n31867 = n279 & n31866 ;
  assign n31868 = n1851 & ~n31867 ;
  assign n31869 = ~n96 & n359 ;
  assign n31870 = ~n359 & n31869 ;
  assign n31871 = ~n669 & n823 ;
  assign n31872 = n31870 & n31871 ;
  assign n31873 = ~n2100 & n31872 ;
  assign n31874 = n3718 & n31873 ;
  assign n31875 = n31868 & ~n31874 ;
  assign n31876 = n31865 & n31875 ;
  assign n31877 = n31876 ^ n30971 ^ 1'b0 ;
  assign n31878 = n20508 | n28908 ;
  assign n31879 = n675 & n21990 ;
  assign n31881 = n1213 ^ n159 ^ 1'b0 ;
  assign n31882 = n2578 & n31881 ;
  assign n31883 = n18387 & n31882 ;
  assign n31884 = n26203 & n31883 ;
  assign n31880 = n2850 & n31181 ;
  assign n31885 = n31884 ^ n31880 ^ 1'b0 ;
  assign n31886 = ~n29491 & n30046 ;
  assign n31887 = n1339 & n31886 ;
  assign n31888 = n13244 ^ n715 ^ 1'b0 ;
  assign n31889 = ~n4025 & n8277 ;
  assign n31890 = ~n3985 & n25734 ;
  assign n31891 = n31889 & n31890 ;
  assign n31892 = n9937 & ~n10705 ;
  assign n31893 = n10322 & n31892 ;
  assign n31894 = n16771 ^ n14218 ^ n4449 ;
  assign n31895 = ~n30433 & n31894 ;
  assign n31896 = ~n16209 & n31895 ;
  assign n31897 = n6887 & n11677 ;
  assign n31898 = n31897 ^ n22657 ^ 1'b0 ;
  assign n31899 = n467 & ~n11069 ;
  assign n31900 = n22357 | n31899 ;
  assign n31901 = ~n2938 & n6524 ;
  assign n31902 = ~n26886 & n31901 ;
  assign n31903 = n27822 & n31902 ;
  assign n31904 = n8088 ^ n4526 ^ 1'b0 ;
  assign n31905 = ~n30 & n31904 ;
  assign n31906 = n8665 ^ n6397 ^ 1'b0 ;
  assign n31907 = n1447 | n31906 ;
  assign n31908 = n28011 | n30746 ;
  assign n31909 = n17939 & n28906 ;
  assign n31910 = n31909 ^ n11851 ^ 1'b0 ;
  assign n31911 = n4167 ^ n3965 ^ 1'b0 ;
  assign n31912 = ~n1361 & n31911 ;
  assign n31913 = n31912 ^ n9104 ^ 1'b0 ;
  assign n31914 = n9617 & n11409 ;
  assign n31915 = n16975 ^ n8049 ^ 1'b0 ;
  assign n31916 = ~n3025 & n31915 ;
  assign n31917 = n3475 & n31916 ;
  assign n31918 = n21848 ^ n12561 ^ 1'b0 ;
  assign n31919 = n23581 & ~n31918 ;
  assign n31920 = n7913 ^ n3394 ^ 1'b0 ;
  assign n31921 = n736 | n24553 ;
  assign n31922 = n13459 ^ n1684 ^ 1'b0 ;
  assign n31923 = n16898 & n31922 ;
  assign n31924 = n27479 & n31923 ;
  assign n31925 = ~n25472 & n31924 ;
  assign n31926 = n12692 & ~n20211 ;
  assign n31927 = n31926 ^ n29239 ^ 1'b0 ;
  assign n31928 = ~n6653 & n8416 ;
  assign n31929 = ~n3270 & n31928 ;
  assign n31930 = n3211 & n31929 ;
  assign n31932 = n13242 & n24445 ;
  assign n31933 = n31932 ^ n7943 ^ 1'b0 ;
  assign n31931 = n4560 | n24701 ;
  assign n31934 = n31933 ^ n31931 ^ 1'b0 ;
  assign n31935 = n28917 ^ n4126 ^ 1'b0 ;
  assign n31936 = n13794 | n31935 ;
  assign n31937 = n2067 & ~n29853 ;
  assign n31938 = n31937 ^ n16176 ^ 1'b0 ;
  assign n31939 = ~n1148 & n7717 ;
  assign n31940 = n1460 & ~n4112 ;
  assign n31941 = n23629 | n31940 ;
  assign n31942 = n1859 & ~n2040 ;
  assign n31943 = n18229 ^ n13583 ^ 1'b0 ;
  assign n31944 = n9107 ^ n4108 ^ 1'b0 ;
  assign n31945 = n2041 & ~n3429 ;
  assign n31946 = ~n3915 & n31945 ;
  assign n31947 = n4394 ^ n3279 ^ 1'b0 ;
  assign n31948 = n31946 & n31947 ;
  assign n31949 = n31948 ^ n82 ^ 1'b0 ;
  assign n31950 = n31944 | n31949 ;
  assign n31951 = n14219 ^ n7908 ^ 1'b0 ;
  assign n31952 = ~n10374 & n31951 ;
  assign n31953 = n879 | n4091 ;
  assign n31954 = n2431 | n3636 ;
  assign n31955 = n31954 ^ n9277 ^ 1'b0 ;
  assign n31956 = n4495 | n9652 ;
  assign n31957 = n7288 & ~n31956 ;
  assign n31958 = n31957 ^ n5979 ^ 1'b0 ;
  assign n31959 = n12185 | n16137 ;
  assign n31960 = n17046 | n31959 ;
  assign n31961 = ~n7077 & n31960 ;
  assign n31962 = ~n9359 & n13759 ;
  assign n31964 = n6015 | n6399 ;
  assign n31965 = n31964 ^ n6475 ^ 1'b0 ;
  assign n31963 = n14676 & n19347 ;
  assign n31966 = n31965 ^ n31963 ^ 1'b0 ;
  assign n31967 = n3022 & n31541 ;
  assign n31968 = n21269 & n31967 ;
  assign n31969 = n5607 & n11516 ;
  assign n31970 = n1360 | n4968 ;
  assign n31971 = n31970 ^ n785 ^ 1'b0 ;
  assign n31972 = n27215 ^ n20638 ^ 1'b0 ;
  assign n31973 = n7040 & n31972 ;
  assign n31974 = n31973 ^ n31060 ^ 1'b0 ;
  assign n31975 = n31971 & n31974 ;
  assign n31976 = ~n3128 & n5424 ;
  assign n31977 = n1249 & n31976 ;
  assign n31978 = n1286 | n31977 ;
  assign n31979 = ~n10370 & n23276 ;
  assign n31980 = ~x0 & n31979 ;
  assign n31981 = n24973 ^ n10442 ^ 1'b0 ;
  assign n31982 = n3770 ^ n895 ^ 1'b0 ;
  assign n31983 = n30155 ^ n16940 ^ 1'b0 ;
  assign n31984 = ~n8185 & n31983 ;
  assign n31985 = n9927 | n30735 ;
  assign n31986 = n21729 ^ n13419 ^ 1'b0 ;
  assign n31987 = n3120 ^ x0 ^ 1'b0 ;
  assign n31988 = n2741 & n31987 ;
  assign n31989 = n8574 ^ n2916 ^ 1'b0 ;
  assign n31990 = n254 & n31989 ;
  assign n31991 = n31988 & ~n31990 ;
  assign n31993 = n3732 | n5011 ;
  assign n31994 = n31993 ^ n30 ^ 1'b0 ;
  assign n31992 = ~n5215 & n25569 ;
  assign n31995 = n31994 ^ n31992 ^ 1'b0 ;
  assign n31996 = n31995 ^ n3843 ^ 1'b0 ;
  assign n31997 = n3467 ^ n3449 ^ 1'b0 ;
  assign n31998 = ~n2302 & n31997 ;
  assign n31999 = n2893 & ~n17493 ;
  assign n32000 = ( n4495 & ~n31998 ) | ( n4495 & n31999 ) | ( ~n31998 & n31999 ) ;
  assign n32001 = n5465 | n7006 ;
  assign n32002 = ~n16262 & n19724 ;
  assign n32003 = ~n9757 & n26604 ;
  assign n32004 = ~n31124 & n31492 ;
  assign n32005 = n7754 & n32004 ;
  assign n32006 = n7871 ^ n4784 ^ 1'b0 ;
  assign n32007 = ~n8347 & n32006 ;
  assign n32008 = n32007 ^ n20329 ^ 1'b0 ;
  assign n32009 = ~n241 & n14798 ;
  assign n32011 = n15639 & n31444 ;
  assign n32010 = n6527 | n13238 ;
  assign n32012 = n32011 ^ n32010 ^ 1'b0 ;
  assign n32013 = n30146 ^ n21638 ^ 1'b0 ;
  assign n32014 = n677 & n32013 ;
  assign n32015 = ~n384 & n10234 ;
  assign n32017 = ~n461 & n1831 ;
  assign n32018 = n32017 ^ n2180 ^ 1'b0 ;
  assign n32019 = n18011 & ~n32018 ;
  assign n32016 = ~n1674 & n2160 ;
  assign n32020 = n32019 ^ n32016 ^ 1'b0 ;
  assign n32021 = n8935 ^ n5501 ^ 1'b0 ;
  assign n32022 = n32020 | n32021 ;
  assign n32023 = n12366 & ~n27501 ;
  assign n32024 = n32023 ^ n3767 ^ 1'b0 ;
  assign n32025 = ~n1368 & n18412 ;
  assign n32026 = ~n13481 & n17134 ;
  assign n32027 = n32026 ^ n3997 ^ 1'b0 ;
  assign n32028 = ~n1789 & n32027 ;
  assign n32029 = n3042 & ~n5158 ;
  assign n32030 = ( n666 & ~n4079 ) | ( n666 & n13682 ) | ( ~n4079 & n13682 ) ;
  assign n32031 = n32030 ^ n14863 ^ n253 ;
  assign n32032 = ~n32029 & n32031 ;
  assign n32033 = ~n10298 & n32032 ;
  assign n32034 = ~n5455 & n32033 ;
  assign n32035 = n32034 ^ n2076 ^ 1'b0 ;
  assign n32036 = n11263 & ~n32035 ;
  assign n32037 = n22195 & ~n32036 ;
  assign n32039 = n14213 & n20021 ;
  assign n32040 = n7379 | n8609 ;
  assign n32041 = n32039 | n32040 ;
  assign n32038 = n5685 | n24536 ;
  assign n32042 = n32041 ^ n32038 ^ 1'b0 ;
  assign n32043 = n8466 & ~n15034 ;
  assign n32044 = n5040 ^ n4700 ^ 1'b0 ;
  assign n32045 = n4626 & ~n5835 ;
  assign n32046 = n32044 & n32045 ;
  assign n32047 = n27264 ^ n3095 ^ 1'b0 ;
  assign n32048 = n5187 ^ n4890 ^ 1'b0 ;
  assign n32049 = ~n13729 & n21808 ;
  assign n32050 = n32049 ^ n29719 ^ 1'b0 ;
  assign n32051 = n13849 ^ n2762 ^ 1'b0 ;
  assign n32052 = n26923 & n32051 ;
  assign n32053 = ~n2865 & n23438 ;
  assign n32054 = ( n30693 & n32052 ) | ( n30693 & ~n32053 ) | ( n32052 & ~n32053 ) ;
  assign n32055 = ~n12854 & n24890 ;
  assign n32056 = n9692 ^ n5310 ^ 1'b0 ;
  assign n32057 = n7640 | n18843 ;
  assign n32058 = n292 & n3660 ;
  assign n32059 = ( n684 & n18423 ) | ( n684 & n31235 ) | ( n18423 & n31235 ) ;
  assign n32060 = ~n3303 & n7578 ;
  assign n32061 = ~n9094 & n32060 ;
  assign n32062 = ~n11939 & n32061 ;
  assign n32063 = n6810 & ~n31428 ;
  assign n32064 = n22880 ^ n11220 ^ 1'b0 ;
  assign n32065 = n1033 | n14543 ;
  assign n32066 = ~n2312 & n19568 ;
  assign n32067 = n10419 | n32066 ;
  assign n32068 = n3131 & ~n23774 ;
  assign n32069 = ~n3131 & n32068 ;
  assign n32070 = n18010 ^ n11433 ^ 1'b0 ;
  assign n32071 = ~n7728 & n24306 ;
  assign n32072 = ~n32070 & n32071 ;
  assign n32073 = n23238 & ~n27501 ;
  assign n32074 = n32073 ^ n1086 ^ 1'b0 ;
  assign n32075 = n32074 ^ n10482 ^ 1'b0 ;
  assign n32076 = n23051 | n26726 ;
  assign n32077 = n17750 & ~n32076 ;
  assign n32079 = n8403 & ~n24389 ;
  assign n32078 = ~n27870 & n31470 ;
  assign n32080 = n32079 ^ n32078 ^ 1'b0 ;
  assign n32081 = n14701 ^ n3150 ^ 1'b0 ;
  assign n32082 = n8863 & n32081 ;
  assign n32083 = n32082 ^ n10246 ^ n3339 ;
  assign n32084 = n31019 ^ n624 ^ 1'b0 ;
  assign n32085 = n425 & ~n11752 ;
  assign n32086 = ( ~n142 & n483 ) | ( ~n142 & n32085 ) | ( n483 & n32085 ) ;
  assign n32087 = n1219 & ~n32086 ;
  assign n32088 = n32087 ^ n1043 ^ 1'b0 ;
  assign n32089 = n1811 & n26595 ;
  assign n32090 = n28532 ^ n16979 ^ 1'b0 ;
  assign n32091 = ~n345 & n11167 ;
  assign n32092 = ( n408 & n32090 ) | ( n408 & ~n32091 ) | ( n32090 & ~n32091 ) ;
  assign n32093 = ~n32089 & n32092 ;
  assign n32094 = n32093 ^ n1613 ^ 1'b0 ;
  assign n32095 = n3745 & ~n32094 ;
  assign n32096 = n3378 & n5877 ;
  assign n32097 = n32096 ^ n2332 ^ 1'b0 ;
  assign n32098 = n2619 & ~n32097 ;
  assign n32099 = n27435 ^ n339 ^ 1'b0 ;
  assign n32100 = n3426 & n18923 ;
  assign n32101 = ~n13576 & n32100 ;
  assign n32102 = n27996 & ~n32101 ;
  assign n32103 = n19527 ^ n6689 ^ 1'b0 ;
  assign n32104 = n32103 ^ n232 ^ 1'b0 ;
  assign n32105 = n2278 | n8081 ;
  assign n32106 = n26991 ^ n9925 ^ 1'b0 ;
  assign n32107 = n231 & n6291 ;
  assign n32108 = ~n24626 & n32107 ;
  assign n32109 = n3581 & ~n17763 ;
  assign n32110 = n4267 & n12103 ;
  assign n32111 = n17517 & ~n25513 ;
  assign n32112 = n637 & ~n13197 ;
  assign n32113 = n6403 & ~n32112 ;
  assign n32114 = n32113 ^ n6265 ^ 1'b0 ;
  assign n32115 = n28810 & ~n32114 ;
  assign n32116 = n32115 ^ n13085 ^ 1'b0 ;
  assign n32117 = n89 & n6331 ;
  assign n32118 = n32117 ^ n2337 ^ 1'b0 ;
  assign n32119 = n8186 ^ n6287 ^ 1'b0 ;
  assign n32120 = ~n32118 & n32119 ;
  assign n32121 = n1431 & ~n9074 ;
  assign n32122 = n32121 ^ n1412 ^ 1'b0 ;
  assign n32123 = n927 & ~n12734 ;
  assign n32124 = n25197 ^ n4446 ^ 1'b0 ;
  assign n32125 = ~n32123 & n32124 ;
  assign n32126 = n2225 | n31014 ;
  assign n32127 = n11831 | n13126 ;
  assign n32128 = n32126 & ~n32127 ;
  assign n32129 = n5551 | n18342 ;
  assign n32130 = n1358 & n16654 ;
  assign n32131 = n4109 & n32130 ;
  assign n32132 = n12236 | n14249 ;
  assign n32133 = ~n13678 & n20694 ;
  assign n32134 = n22279 & n32133 ;
  assign n32135 = n32134 ^ n25305 ^ 1'b0 ;
  assign n32136 = ~n10845 & n32135 ;
  assign n32137 = n12561 | n18219 ;
  assign n32138 = ( n17794 & n27620 ) | ( n17794 & n29046 ) | ( n27620 & n29046 ) ;
  assign n32139 = n32138 ^ n18492 ^ 1'b0 ;
  assign n32140 = ~n4919 & n32139 ;
  assign n32141 = ~n883 & n26966 ;
  assign n32142 = n32141 ^ n12095 ^ 1'b0 ;
  assign n32143 = n15333 ^ n102 ^ 1'b0 ;
  assign n32144 = ( n11263 & n15609 ) | ( n11263 & n32143 ) | ( n15609 & n32143 ) ;
  assign n32145 = n32144 ^ n20051 ^ n1538 ;
  assign n32146 = n32145 ^ n27437 ^ 1'b0 ;
  assign n32147 = n22426 ^ n142 ^ 1'b0 ;
  assign n32148 = ~n10787 & n13083 ;
  assign n32149 = ~n17668 & n32148 ;
  assign n32150 = n729 & n6412 ;
  assign n32151 = n823 & n32150 ;
  assign n32152 = n23438 & n32151 ;
  assign n32153 = n32152 ^ n56 ^ 1'b0 ;
  assign n32154 = n2948 & ~n12194 ;
  assign n32155 = n32154 ^ n18534 ^ 1'b0 ;
  assign n32156 = ~n32153 & n32155 ;
  assign n32157 = n27679 ^ n15454 ^ 1'b0 ;
  assign n32158 = n18921 | n32157 ;
  assign n32159 = n15047 & n23926 ;
  assign n32160 = n19829 ^ n5968 ^ 1'b0 ;
  assign n32161 = n8191 & n25104 ;
  assign n32162 = n32161 ^ n9672 ^ 1'b0 ;
  assign n32163 = n23059 ^ n14889 ^ 1'b0 ;
  assign n32164 = n4796 & ~n8515 ;
  assign n32165 = n23 & ~n2155 ;
  assign n32166 = ~n7516 & n32165 ;
  assign n32167 = ~n32164 & n32166 ;
  assign n32168 = n7147 | n32167 ;
  assign n32169 = n32168 ^ n10067 ^ 1'b0 ;
  assign n32173 = n3786 ^ n1670 ^ 1'b0 ;
  assign n32171 = n2096 & ~n16548 ;
  assign n32170 = n15237 | n15325 ;
  assign n32172 = n32171 ^ n32170 ^ 1'b0 ;
  assign n32174 = n32173 ^ n32172 ^ 1'b0 ;
  assign n32175 = ~n9119 & n9992 ;
  assign n32176 = n3182 & n32175 ;
  assign n32177 = n32176 ^ n3793 ^ 1'b0 ;
  assign n32178 = ~n11478 & n21453 ;
  assign n32179 = n3269 & ~n28058 ;
  assign n32180 = ~n23001 & n32179 ;
  assign n32181 = n1929 | n32180 ;
  assign n32182 = n10930 ^ n1431 ^ 1'b0 ;
  assign n32183 = n20059 | n32182 ;
  assign n32184 = n19426 ^ n11298 ^ 1'b0 ;
  assign n32185 = ~n11893 & n17063 ;
  assign n32186 = n13422 & ~n17616 ;
  assign n32187 = ~n3007 & n3219 ;
  assign n32188 = n10621 | n24058 ;
  assign n32189 = n13131 ^ n12561 ^ 1'b0 ;
  assign n32190 = n23321 & n32189 ;
  assign n32191 = n2842 & n26181 ;
  assign n32192 = n32191 ^ n6538 ^ 1'b0 ;
  assign n32193 = n7599 ^ n6187 ^ n5363 ;
  assign n32194 = n4348 & ~n32193 ;
  assign n32195 = n86 & n205 ;
  assign n32196 = ( ~n1119 & n32194 ) | ( ~n1119 & n32195 ) | ( n32194 & n32195 ) ;
  assign n32197 = n21818 ^ n334 ^ 1'b0 ;
  assign n32198 = n3282 & ~n32197 ;
  assign n32199 = n1984 & ~n12214 ;
  assign n32200 = ~n191 & n32199 ;
  assign n32201 = ( n16803 & n32198 ) | ( n16803 & ~n32200 ) | ( n32198 & ~n32200 ) ;
  assign n32202 = n7221 & n8430 ;
  assign n32203 = n32202 ^ n18856 ^ 1'b0 ;
  assign n32204 = n32201 & ~n32203 ;
  assign n32205 = n3297 & n13385 ;
  assign n32206 = n32205 ^ n25716 ^ 1'b0 ;
  assign n32207 = n10069 & n15415 ;
  assign n32208 = ~n18874 & n32207 ;
  assign n32209 = n12967 & ~n32208 ;
  assign n32210 = ~n1458 & n32209 ;
  assign n32211 = n5322 ^ n3418 ^ 1'b0 ;
  assign n32212 = n78 & n32211 ;
  assign n32213 = n10543 ^ n86 ^ 1'b0 ;
  assign n32214 = ~n1707 & n14694 ;
  assign n32215 = ~n661 & n23907 ;
  assign n32216 = ~n1158 & n32215 ;
  assign n32217 = ~n11400 & n30229 ;
  assign n32218 = n2117 | n2909 ;
  assign n32219 = n32218 ^ n17891 ^ 1'b0 ;
  assign n32220 = ~n8563 & n12219 ;
  assign n32221 = n32219 & n32220 ;
  assign n32222 = n213 & n666 ;
  assign n32223 = ~n213 & n32222 ;
  assign n32224 = n1501 | n32223 ;
  assign n32225 = n1501 & ~n32224 ;
  assign n32226 = n29407 | n32225 ;
  assign n32227 = n29407 & ~n32226 ;
  assign n32228 = ~n294 & n32227 ;
  assign n32229 = n5046 | n32228 ;
  assign n32230 = n43 & n28589 ;
  assign n32231 = n32230 ^ n1034 ^ 1'b0 ;
  assign n32232 = ~n4253 & n32231 ;
  assign n32233 = ~n32229 & n32232 ;
  assign n32234 = n5006 & ~n11106 ;
  assign n32235 = n5534 ^ n618 ^ 1'b0 ;
  assign n32236 = n32234 & ~n32235 ;
  assign n32237 = n20048 & n32236 ;
  assign n32238 = n32237 ^ n29027 ^ 1'b0 ;
  assign n32239 = n9149 & ~n14269 ;
  assign n32240 = ~n7875 & n32239 ;
  assign n32241 = n24156 & ~n27169 ;
  assign n32242 = n32240 & n32241 ;
  assign n32243 = n13791 & ~n32242 ;
  assign n32244 = n16645 ^ n2988 ^ 1'b0 ;
  assign n32245 = ~n5507 & n32244 ;
  assign n32246 = n4495 ^ n1710 ^ 1'b0 ;
  assign n32247 = n4009 & ~n32246 ;
  assign n32248 = n32247 ^ n32086 ^ 1'b0 ;
  assign n32249 = ~n15754 & n18235 ;
  assign n32250 = n13128 | n29572 ;
  assign n32251 = n6809 & ~n32250 ;
  assign n32252 = n9744 & n16339 ;
  assign n32254 = n14211 & n25010 ;
  assign n32255 = ~n14234 & n32254 ;
  assign n32253 = n6897 & n22086 ;
  assign n32256 = n32255 ^ n32253 ^ 1'b0 ;
  assign n32257 = ~n1456 & n11487 ;
  assign n32258 = n32150 ^ n22204 ^ 1'b0 ;
  assign n32259 = n1354 & ~n30964 ;
  assign n32260 = n246 ^ n38 ^ 1'b0 ;
  assign n32261 = n18614 ^ n9362 ^ 1'b0 ;
  assign n32262 = ~n1946 & n18275 ;
  assign n32263 = n32262 ^ n10638 ^ 1'b0 ;
  assign n32264 = n10899 ^ n9977 ^ 1'b0 ;
  assign n32267 = n777 & ~n2116 ;
  assign n32268 = ~n777 & n32267 ;
  assign n32269 = n495 & n32268 ;
  assign n32270 = n2567 & ~n32269 ;
  assign n32271 = n32270 ^ n18697 ^ 1'b0 ;
  assign n32265 = ~n1515 & n11680 ;
  assign n32266 = n1515 & n32265 ;
  assign n32272 = n32271 ^ n32266 ^ 1'b0 ;
  assign n32273 = n32272 ^ n26687 ^ 1'b0 ;
  assign n32274 = ~n28438 & n32273 ;
  assign n32275 = n7973 ^ n34 ^ 1'b0 ;
  assign n32276 = n32275 ^ n4326 ^ 1'b0 ;
  assign n32277 = n32276 ^ n10228 ^ 1'b0 ;
  assign n32278 = n4424 | n7981 ;
  assign n32279 = n32278 ^ n8253 ^ 1'b0 ;
  assign n32280 = n3929 | n6025 ;
  assign n32281 = n32280 ^ n2773 ^ 1'b0 ;
  assign n32282 = ~n2567 & n32281 ;
  assign n32283 = n32282 ^ n2117 ^ 1'b0 ;
  assign n32284 = ~n21526 & n32283 ;
  assign n32285 = ~n32279 & n32284 ;
  assign n32286 = n27747 ^ n3223 ^ 1'b0 ;
  assign n32287 = n2017 & n24773 ;
  assign n32288 = n32287 ^ n9154 ^ 1'b0 ;
  assign n32289 = n9988 | n32288 ;
  assign n32290 = n14159 ^ n1315 ^ 1'b0 ;
  assign n32291 = n13591 | n32290 ;
  assign n32292 = n14240 ^ n7487 ^ 1'b0 ;
  assign n32293 = n6246 & ~n32292 ;
  assign n32294 = n1989 & n18004 ;
  assign n32295 = ~n8392 & n27272 ;
  assign n32296 = n32295 ^ n21752 ^ 1'b0 ;
  assign n32297 = n20596 ^ n12781 ^ 1'b0 ;
  assign n32298 = ~n8654 & n10022 ;
  assign n32299 = n19390 & ~n32298 ;
  assign n32300 = n25113 & ~n32299 ;
  assign n32301 = n32297 & n32300 ;
  assign n32302 = n5385 ^ n2571 ^ 1'b0 ;
  assign n32303 = ~n29985 & n32302 ;
  assign n32306 = n15906 ^ n5130 ^ 1'b0 ;
  assign n32304 = n11376 ^ n6131 ^ 1'b0 ;
  assign n32305 = n1325 | n32304 ;
  assign n32307 = n32306 ^ n32305 ^ n25154 ;
  assign n32308 = n30750 & ~n32307 ;
  assign n32310 = n2269 & ~n8245 ;
  assign n32311 = n20934 & n32310 ;
  assign n32312 = n7357 & ~n32311 ;
  assign n32313 = ~n7357 & n32312 ;
  assign n32314 = ~n446 & n32313 ;
  assign n32309 = n139 & ~n31492 ;
  assign n32315 = n32314 ^ n32309 ^ n23583 ;
  assign n32316 = n5758 & n25444 ;
  assign n32317 = ( n4422 & ~n22941 ) | ( n4422 & n31213 ) | ( ~n22941 & n31213 ) ;
  assign n32318 = n22261 | n32317 ;
  assign n32319 = n16102 ^ n13583 ^ 1'b0 ;
  assign n32320 = n32318 & n32319 ;
  assign n32321 = n3027 & ~n7641 ;
  assign n32322 = n32321 ^ n7895 ^ n3567 ;
  assign n32323 = n5444 & ~n17652 ;
  assign n32324 = n3810 & n32323 ;
  assign n32325 = n9925 & n32324 ;
  assign n32326 = n17527 ^ n9577 ^ n1637 ;
  assign n32327 = n22840 ^ n5471 ^ 1'b0 ;
  assign n32328 = n3415 & ~n30682 ;
  assign n32329 = n32328 ^ n8463 ^ 1'b0 ;
  assign n32330 = n31459 ^ n14549 ^ 1'b0 ;
  assign n32331 = n814 & n8197 ;
  assign n32332 = n372 & ~n16311 ;
  assign n32333 = n17096 ^ n13435 ^ 1'b0 ;
  assign n32334 = n4931 ^ n4538 ^ 1'b0 ;
  assign n32335 = n15183 ^ n968 ^ 1'b0 ;
  assign n32336 = n32335 ^ n1790 ^ 1'b0 ;
  assign n32337 = n32336 ^ n24442 ^ 1'b0 ;
  assign n32338 = ~n4174 & n19580 ;
  assign n32339 = n32338 ^ n14815 ^ 1'b0 ;
  assign n32340 = n24025 | n32339 ;
  assign n32341 = n10265 | n11833 ;
  assign n32342 = n28283 & ~n32341 ;
  assign n32343 = ~n13707 & n16808 ;
  assign n32344 = n12354 ^ n11696 ^ 1'b0 ;
  assign n32345 = n11919 | n28365 ;
  assign n32346 = n6784 ^ n6277 ^ n3138 ;
  assign n32347 = n500 | n32346 ;
  assign n32348 = n14043 & ~n32347 ;
  assign n32349 = n3428 & ~n7667 ;
  assign n32350 = n252 & n9920 ;
  assign n32351 = ( n23197 & n32349 ) | ( n23197 & n32350 ) | ( n32349 & n32350 ) ;
  assign n32352 = n9398 & n17279 ;
  assign n32353 = ~n26208 & n32352 ;
  assign n32354 = n20145 ^ n5308 ^ 1'b0 ;
  assign n32355 = n3406 | n8530 ;
  assign n32356 = n11494 & n21793 ;
  assign n32357 = ~n497 & n6006 ;
  assign n32358 = n25102 ^ n5261 ^ 1'b0 ;
  assign n32359 = n32357 & ~n32358 ;
  assign n32360 = n2391 ^ n158 ^ 1'b0 ;
  assign n32361 = ( ~n8450 & n32359 ) | ( ~n8450 & n32360 ) | ( n32359 & n32360 ) ;
  assign n32362 = ~n21890 & n32361 ;
  assign n32363 = n9399 & n32362 ;
  assign n32364 = n10651 & ~n10818 ;
  assign n32365 = n32364 ^ n19249 ^ 1'b0 ;
  assign n32366 = n1886 & n7040 ;
  assign n32367 = n17178 & ~n32366 ;
  assign n32368 = n13870 ^ n11838 ^ 1'b0 ;
  assign n32369 = ~n25764 & n32368 ;
  assign n32370 = n3103 | n28400 ;
  assign n32371 = n32370 ^ n27427 ^ 1'b0 ;
  assign n32372 = n2511 | n2684 ;
  assign n32373 = n19910 & ~n21656 ;
  assign n32374 = n32373 ^ n10617 ^ 1'b0 ;
  assign n32375 = n361 & n31087 ;
  assign n32376 = n32375 ^ n27590 ^ 1'b0 ;
  assign n32377 = n12865 ^ n10296 ^ 1'b0 ;
  assign n32378 = n14716 & ~n32377 ;
  assign n32379 = n3680 & ~n6739 ;
  assign n32380 = n32378 & n32379 ;
  assign n32381 = ~n1178 & n32380 ;
  assign n32382 = n27656 ^ n24837 ^ n7117 ;
  assign n32383 = ~n1065 & n24868 ;
  assign n32384 = ~n158 & n7294 ;
  assign n32385 = n28734 ^ n1608 ^ 1'b0 ;
  assign n32386 = n849 & ~n12214 ;
  assign n32387 = n32386 ^ n22076 ^ 1'b0 ;
  assign n32389 = n8321 ^ n1760 ^ 1'b0 ;
  assign n32388 = n2878 | n11003 ;
  assign n32390 = n32389 ^ n32388 ^ 1'b0 ;
  assign n32391 = n13751 & ~n32390 ;
  assign n32392 = n13434 & ~n19022 ;
  assign n32393 = n32392 ^ n9915 ^ 1'b0 ;
  assign n32394 = ~n20672 & n31837 ;
  assign n32395 = ~n30317 & n32394 ;
  assign n32396 = n32395 ^ n30537 ^ n8561 ;
  assign n32397 = n478 | n17456 ;
  assign n32398 = n478 & ~n32397 ;
  assign n32399 = n32398 ^ n1688 ^ 1'b0 ;
  assign n32400 = n20456 & ~n32399 ;
  assign n32401 = ~n20456 & n32400 ;
  assign n32402 = n685 | n8570 ;
  assign n32403 = n459 & n5264 ;
  assign n32404 = n2294 & n10635 ;
  assign n32405 = n227 & n32404 ;
  assign n32406 = n323 & n10030 ;
  assign n32407 = n32405 & n32406 ;
  assign n32409 = n1316 | n1416 ;
  assign n32408 = n1105 & n15126 ;
  assign n32410 = n32409 ^ n32408 ^ 1'b0 ;
  assign n32411 = n32410 ^ n14120 ^ 1'b0 ;
  assign n32412 = ~n13997 & n32411 ;
  assign n32413 = n8624 & n32412 ;
  assign n32414 = n10461 & ~n17884 ;
  assign n32415 = n30956 ^ n843 ^ 1'b0 ;
  assign n32416 = n18899 & n32415 ;
  assign n32417 = n1222 & n32416 ;
  assign n32418 = n32417 ^ n6420 ^ 1'b0 ;
  assign n32419 = n28549 ^ n3928 ^ 1'b0 ;
  assign n32420 = n7522 | n9521 ;
  assign n32421 = n13628 & ~n32420 ;
  assign n32422 = n32421 ^ n17466 ^ n10215 ;
  assign n32423 = n13087 | n32070 ;
  assign n32424 = ~n556 & n25356 ;
  assign n32425 = n32424 ^ n9291 ^ 1'b0 ;
  assign n32426 = ~n7179 & n21884 ;
  assign n32427 = n32426 ^ n12205 ^ 1'b0 ;
  assign n32428 = n3729 & n32427 ;
  assign n32429 = n2681 ^ n1227 ^ 1'b0 ;
  assign n32430 = n16474 ^ n4227 ^ n1988 ;
  assign n32431 = ( n891 & ~n32429 ) | ( n891 & n32430 ) | ( ~n32429 & n32430 ) ;
  assign n32432 = n13118 & ~n21103 ;
  assign n32433 = n9033 & n11153 ;
  assign n32434 = ( n4165 & ~n9619 ) | ( n4165 & n11691 ) | ( ~n9619 & n11691 ) ;
  assign n32435 = n20375 | n32434 ;
  assign n32436 = n165 | n32435 ;
  assign n32437 = ~n21811 & n32436 ;
  assign n32438 = n4936 ^ n3452 ^ 1'b0 ;
  assign n32439 = n7615 | n32438 ;
  assign n32440 = n10797 & n20549 ;
  assign n32441 = n32440 ^ n4668 ^ 1'b0 ;
  assign n32442 = n3931 & ~n8457 ;
  assign n32443 = n32442 ^ n29850 ^ 1'b0 ;
  assign n32444 = n18798 & n32443 ;
  assign n32445 = n12324 | n19609 ;
  assign n32446 = ~n10962 & n12273 ;
  assign n32447 = n1674 & n32446 ;
  assign n32448 = n32447 ^ n2295 ^ 1'b0 ;
  assign n32449 = n31348 & n31916 ;
  assign n32450 = ~n10806 & n17010 ;
  assign n32451 = n32450 ^ n23381 ^ n4292 ;
  assign n32452 = n32451 ^ n32361 ^ 1'b0 ;
  assign n32453 = n21860 & n32452 ;
  assign n32454 = ~n12382 & n20997 ;
  assign n32455 = n32454 ^ n11722 ^ 1'b0 ;
  assign n32456 = n1960 & n16830 ;
  assign n32457 = n1003 | n9211 ;
  assign n32458 = n32457 ^ n17030 ^ 1'b0 ;
  assign n32459 = ~n32456 & n32458 ;
  assign n32460 = n12165 ^ n1912 ^ 1'b0 ;
  assign n32461 = n3103 | n32460 ;
  assign n32462 = n6477 ^ n3337 ^ 1'b0 ;
  assign n32463 = n16230 | n32462 ;
  assign n32464 = n313 & ~n7153 ;
  assign n32465 = ~n32463 & n32464 ;
  assign n32466 = n32465 ^ n6384 ^ 1'b0 ;
  assign n32467 = ( n3078 & ~n7943 ) | ( n3078 & n8562 ) | ( ~n7943 & n8562 ) ;
  assign n32468 = n15867 & ~n32467 ;
  assign n32469 = n177 | n27166 ;
  assign n32470 = n489 & ~n9422 ;
  assign n32471 = ~n11674 & n32470 ;
  assign n32472 = n1768 | n32471 ;
  assign n32473 = ~n18530 & n32472 ;
  assign n32474 = n32360 ^ n785 ^ 1'b0 ;
  assign n32475 = ~n5570 & n25397 ;
  assign n32476 = n32475 ^ n12222 ^ 1'b0 ;
  assign n32477 = n2984 & n3049 ;
  assign n32478 = n5684 ^ n2191 ^ 1'b0 ;
  assign n32479 = n32477 & ~n32478 ;
  assign n32480 = n4462 & n6926 ;
  assign n32481 = n13478 ^ n729 ^ 1'b0 ;
  assign n32482 = n11855 ^ n7681 ^ 1'b0 ;
  assign n32483 = ~n6461 & n32482 ;
  assign n32484 = n32481 & n32483 ;
  assign n32485 = n4191 & n24582 ;
  assign n32486 = ~n2100 & n18778 ;
  assign n32487 = ~n16294 & n32486 ;
  assign n32488 = n6230 & ~n32487 ;
  assign n32489 = n28331 ^ n15400 ^ 1'b0 ;
  assign n32490 = n24669 | n30069 ;
  assign n32491 = n14241 & n32490 ;
  assign n32492 = ~n3162 & n32491 ;
  assign n32493 = n26264 ^ n17475 ^ 1'b0 ;
  assign n32494 = n32493 ^ n16910 ^ n52 ;
  assign n32495 = n32492 | n32494 ;
  assign n32496 = n7754 ^ n7430 ^ 1'b0 ;
  assign n32497 = n4003 & n32496 ;
  assign n32498 = n32497 ^ n3363 ^ 1'b0 ;
  assign n32499 = ~n500 & n11968 ;
  assign n32500 = n32498 & n32499 ;
  assign n32501 = ~n6376 & n27491 ;
  assign n32502 = n22422 | n32501 ;
  assign n32503 = n32502 ^ n21496 ^ 1'b0 ;
  assign n32505 = n1004 & ~n14238 ;
  assign n32504 = n284 & n22387 ;
  assign n32506 = n32505 ^ n32504 ^ 1'b0 ;
  assign n32507 = ~n4668 & n21988 ;
  assign n32508 = n77 & n29056 ;
  assign n32509 = n16621 ^ n5359 ^ 1'b0 ;
  assign n32510 = ~n17623 & n32509 ;
  assign n32511 = n24083 ^ n2235 ^ 1'b0 ;
  assign n32513 = n3997 & ~n4519 ;
  assign n32514 = n32513 ^ n2200 ^ 1'b0 ;
  assign n32515 = n28137 | n32514 ;
  assign n32512 = n415 & ~n1552 ;
  assign n32516 = n32515 ^ n32512 ^ 1'b0 ;
  assign n32517 = n10392 & ~n19020 ;
  assign n32518 = ~n6942 & n16196 ;
  assign n32519 = n11821 & n32518 ;
  assign n32520 = n14539 & ~n17621 ;
  assign n32521 = n32520 ^ n5180 ^ 1'b0 ;
  assign n32522 = n9758 & ~n32521 ;
  assign n32523 = n11401 & ~n17831 ;
  assign n32524 = n1865 & ~n3483 ;
  assign n32525 = n8253 & ~n32524 ;
  assign n32526 = n21651 ^ n9625 ^ 1'b0 ;
  assign n32527 = n5336 | n32526 ;
  assign n32528 = ~n11933 & n13588 ;
  assign n32529 = n16782 & n29140 ;
  assign n32530 = n5345 | n8827 ;
  assign n32531 = n3053 | n6539 ;
  assign n32532 = n4533 | n22107 ;
  assign n32533 = n32531 | n32532 ;
  assign n32534 = n27302 & n32533 ;
  assign n32535 = n5758 & ~n18433 ;
  assign n32536 = ~n7503 & n32535 ;
  assign n32537 = n24888 ^ n14272 ^ 1'b0 ;
  assign n32538 = n32148 ^ n3396 ^ 1'b0 ;
  assign n32539 = n2202 | n14089 ;
  assign n32540 = ~n5419 & n13206 ;
  assign n32541 = ~n32539 & n32540 ;
  assign n32542 = n4437 & ~n32541 ;
  assign n32543 = n190 ^ n169 ^ 1'b0 ;
  assign n32544 = n1965 ^ n905 ^ 1'b0 ;
  assign n32545 = ~n32543 & n32544 ;
  assign n32546 = n3820 & n32545 ;
  assign n32547 = n2509 & n25684 ;
  assign n32548 = n32547 ^ n12697 ^ 1'b0 ;
  assign n32549 = n626 | n12092 ;
  assign n32550 = n32549 ^ n1874 ^ 1'b0 ;
  assign n32551 = ~n621 & n17561 ;
  assign n32552 = n32551 ^ n10881 ^ 1'b0 ;
  assign n32553 = n32552 ^ n2545 ^ n542 ;
  assign n32554 = n14269 ^ n12265 ^ 1'b0 ;
  assign n32555 = n12457 | n32554 ;
  assign n32556 = ~n4657 & n13930 ;
  assign n32557 = n32556 ^ n26854 ^ 1'b0 ;
  assign n32558 = n1825 & n8302 ;
  assign n32559 = n17497 & n32558 ;
  assign n32560 = n3850 ^ n3056 ^ 1'b0 ;
  assign n32561 = n4155 & n32560 ;
  assign n32562 = ( n1404 & ~n6855 ) | ( n1404 & n32561 ) | ( ~n6855 & n32561 ) ;
  assign n32563 = n6210 & n14433 ;
  assign n32564 = ~n4217 & n32563 ;
  assign n32565 = n2266 & ~n2664 ;
  assign n32566 = n32565 ^ n1878 ^ 1'b0 ;
  assign n32567 = ~n3211 & n32361 ;
  assign n32568 = n32567 ^ n5161 ^ 1'b0 ;
  assign n32569 = ~n2490 & n10572 ;
  assign n32570 = ~n31433 & n32569 ;
  assign n32572 = n297 & n14088 ;
  assign n32571 = ~n3467 & n21375 ;
  assign n32573 = n32572 ^ n32571 ^ 1'b0 ;
  assign n32574 = n4580 & n28848 ;
  assign n32575 = n32574 ^ n2198 ^ 1'b0 ;
  assign n32576 = n7327 | n28356 ;
  assign n32577 = n32576 ^ n6488 ^ 1'b0 ;
  assign n32578 = n16728 ^ n1098 ^ 1'b0 ;
  assign n32579 = ~n68 & n5180 ;
  assign n32580 = ~n32578 & n32579 ;
  assign n32581 = n16338 ^ n3668 ^ 1'b0 ;
  assign n32582 = n19455 ^ n9019 ^ n3394 ;
  assign n32583 = n9195 ^ n2436 ^ 1'b0 ;
  assign n32584 = n4674 & ~n6712 ;
  assign n32585 = n22180 & n27308 ;
  assign n32586 = ~n468 & n21394 ;
  assign n32587 = ~n181 & n32586 ;
  assign n32588 = n3074 ^ n2790 ^ 1'b0 ;
  assign n32589 = ~n32587 & n32588 ;
  assign n32590 = n21340 & n32589 ;
  assign n32591 = ~n29703 & n30410 ;
  assign n32592 = n11436 & n29882 ;
  assign n32593 = n6154 | n27748 ;
  assign n32594 = n32593 ^ n7998 ^ 1'b0 ;
  assign n32595 = ~n27876 & n29916 ;
  assign n32596 = n3966 ^ n1183 ^ 1'b0 ;
  assign n32597 = ( n7717 & ~n8167 ) | ( n7717 & n32596 ) | ( ~n8167 & n32596 ) ;
  assign n32598 = n3348 | n5801 ;
  assign n32599 = n27366 & ~n27473 ;
  assign n32600 = n7140 ^ n5164 ^ 1'b0 ;
  assign n32601 = ~n13967 & n32600 ;
  assign n32602 = ~n13198 & n32601 ;
  assign n32603 = n16820 & n32602 ;
  assign n32604 = n4478 | n32603 ;
  assign n32605 = n6889 & n23317 ;
  assign n32606 = n32605 ^ n1213 ^ 1'b0 ;
  assign n32607 = n3850 ^ n3443 ^ 1'b0 ;
  assign n32608 = n3526 | n32607 ;
  assign n32609 = n14986 & ~n20618 ;
  assign n32610 = n7241 & n14325 ;
  assign n32611 = ~n24784 & n29144 ;
  assign n32612 = n32611 ^ n6714 ^ 1'b0 ;
  assign n32613 = ~n1933 & n8318 ;
  assign n32614 = n323 | n5128 ;
  assign n32615 = n3221 & ~n32614 ;
  assign n32616 = n31690 ^ n12993 ^ 1'b0 ;
  assign n32617 = n32616 ^ n1406 ^ 1'b0 ;
  assign n32618 = n7120 & ~n32617 ;
  assign n32619 = ~n940 & n25657 ;
  assign n32620 = n10124 | n30080 ;
  assign n32621 = n32620 ^ n628 ^ 1'b0 ;
  assign n32622 = n29152 | n31618 ;
  assign n32623 = n22817 ^ n15725 ^ 1'b0 ;
  assign n32624 = ~n32622 & n32623 ;
  assign n32631 = n7216 ^ n2499 ^ 1'b0 ;
  assign n32632 = n32405 | n32631 ;
  assign n32625 = n9306 | n12730 ;
  assign n32626 = n32625 ^ n6506 ^ 1'b0 ;
  assign n32627 = ~n10998 & n15334 ;
  assign n32628 = n32627 ^ n2059 ^ 1'b0 ;
  assign n32629 = n11108 | n32628 ;
  assign n32630 = n32626 & ~n32629 ;
  assign n32633 = n32632 ^ n32630 ^ 1'b0 ;
  assign n32634 = n20000 | n32633 ;
  assign n32635 = ( n986 & ~n4018 ) | ( n986 & n9623 ) | ( ~n4018 & n9623 ) ;
  assign n32636 = n26105 ^ n20512 ^ 1'b0 ;
  assign n32637 = ~n32635 & n32636 ;
  assign n32638 = n4784 & n4991 ;
  assign n32639 = n32638 ^ n20494 ^ 1'b0 ;
  assign n32640 = n6019 & n24657 ;
  assign n32641 = n26081 ^ n18839 ^ 1'b0 ;
  assign n32642 = n5583 & n11594 ;
  assign n32643 = n24335 ^ n13726 ^ 1'b0 ;
  assign n32644 = ~x3 & n10658 ;
  assign n32645 = n8042 ^ n2012 ^ 1'b0 ;
  assign n32646 = n32644 | n32645 ;
  assign n32647 = n8946 | n17221 ;
  assign n32648 = n32647 ^ n83 ^ 1'b0 ;
  assign n32649 = n2076 | n10527 ;
  assign n32650 = n32649 ^ n479 ^ 1'b0 ;
  assign n32651 = n14110 & n32650 ;
  assign n32652 = n6569 & ~n12924 ;
  assign n32653 = ~n21257 & n32652 ;
  assign n32658 = n8785 | n13822 ;
  assign n32659 = n2279 | n32658 ;
  assign n32654 = n9117 ^ n2696 ^ 1'b0 ;
  assign n32655 = n832 | n4891 ;
  assign n32656 = n32654 & ~n32655 ;
  assign n32657 = n24827 & ~n32656 ;
  assign n32660 = n32659 ^ n32657 ^ 1'b0 ;
  assign n32661 = n2150 ^ n741 ^ 1'b0 ;
  assign n32662 = n4098 | n32661 ;
  assign n32663 = n14813 | n16069 ;
  assign n32664 = n2314 | n7407 ;
  assign n32665 = n32664 ^ n10280 ^ 1'b0 ;
  assign n32667 = n16351 ^ n13913 ^ 1'b0 ;
  assign n32668 = n20610 | n32667 ;
  assign n32666 = ~n3939 & n25572 ;
  assign n32669 = n32668 ^ n32666 ^ 1'b0 ;
  assign n32671 = n27737 | n30506 ;
  assign n32672 = n7227 & ~n32671 ;
  assign n32670 = ~n15788 & n27920 ;
  assign n32673 = n32672 ^ n32670 ^ 1'b0 ;
  assign n32674 = n3398 & n18780 ;
  assign n32675 = n2044 ^ n671 ^ 1'b0 ;
  assign n32676 = n32674 & n32675 ;
  assign n32677 = n175 | n19094 ;
  assign n32678 = n6027 | n32677 ;
  assign n32679 = n21004 ^ n17923 ^ 1'b0 ;
  assign n32680 = n21373 ^ n7920 ^ 1'b0 ;
  assign n32681 = n25444 & ~n32680 ;
  assign n32682 = n32681 ^ n43 ^ 1'b0 ;
  assign n32683 = n1246 & n12776 ;
  assign n32684 = n11246 & ~n13726 ;
  assign n32685 = n23979 ^ n13487 ^ 1'b0 ;
  assign n32686 = n421 & ~n6549 ;
  assign n32687 = n32686 ^ n27827 ^ 1'b0 ;
  assign n32688 = ~n8448 & n9839 ;
  assign n32689 = ~n17113 & n25562 ;
  assign n32690 = ~n15225 & n18930 ;
  assign n32691 = ~n855 & n3928 ;
  assign n32692 = n6721 & n32691 ;
  assign n32693 = ~n13114 & n26489 ;
  assign n32694 = ~n6229 & n32693 ;
  assign n32695 = n3110 | n19293 ;
  assign n32696 = n3748 | n7033 ;
  assign n32697 = n32696 ^ n31446 ^ n820 ;
  assign n32698 = n27933 ^ n13238 ^ 1'b0 ;
  assign n32699 = n1435 & n32698 ;
  assign n32700 = n10583 & ~n12734 ;
  assign n32701 = n1585 & ~n32700 ;
  assign n32702 = n9212 & n32701 ;
  assign n32703 = n32702 ^ n17029 ^ 1'b0 ;
  assign n32704 = n10047 ^ n7625 ^ 1'b0 ;
  assign n32705 = n12717 ^ n2679 ^ 1'b0 ;
  assign n32706 = n11008 & ~n32705 ;
  assign n32707 = n7263 & n32706 ;
  assign n32708 = n11685 ^ n5254 ^ 1'b0 ;
  assign n32709 = n200 | n16400 ;
  assign n32710 = n24072 & ~n32709 ;
  assign n32711 = n1947 & ~n32710 ;
  assign n32712 = n869 & ~n11024 ;
  assign n32713 = n32712 ^ n13098 ^ 1'b0 ;
  assign n32714 = n2438 & n7866 ;
  assign n32715 = n719 & n4203 ;
  assign n32716 = n13634 | n23309 ;
  assign n32717 = n10092 ^ n4058 ^ 1'b0 ;
  assign n32718 = n1152 & n21956 ;
  assign n32719 = n32718 ^ n16007 ^ 1'b0 ;
  assign n32720 = n32719 ^ n4133 ^ 1'b0 ;
  assign n32721 = n7327 & n15172 ;
  assign n32722 = n31162 & n32721 ;
  assign n32723 = n9134 & n32722 ;
  assign n32724 = n227 & ~n14822 ;
  assign n32725 = n8686 | n23581 ;
  assign n32726 = n5099 & ~n13592 ;
  assign n32727 = n13098 ^ n2497 ^ 1'b0 ;
  assign n32728 = n10531 & n32727 ;
  assign n32729 = ~n1208 & n4607 ;
  assign n32730 = n9977 | n32729 ;
  assign n32731 = n31171 & ~n32730 ;
  assign n32732 = n6194 & ~n20612 ;
  assign n32733 = n32732 ^ n25526 ^ 1'b0 ;
  assign n32734 = n3741 ^ n272 ^ 1'b0 ;
  assign n32735 = n32734 ^ n21546 ^ 1'b0 ;
  assign n32736 = n2872 | n32735 ;
  assign n32748 = n787 & n2397 ;
  assign n32749 = n26697 & n32748 ;
  assign n32750 = n442 | n474 ;
  assign n32751 = n32749 & ~n32750 ;
  assign n32752 = ~n1082 & n32751 ;
  assign n32753 = ~n1183 & n2624 ;
  assign n32754 = n1183 & n32753 ;
  assign n32755 = n3633 | n32754 ;
  assign n32756 = n32752 & ~n32755 ;
  assign n32737 = n1267 & ~n13314 ;
  assign n32738 = ~n1267 & n32737 ;
  assign n32739 = n2623 & ~n27281 ;
  assign n32740 = n27281 & n32739 ;
  assign n32741 = n32738 | n32740 ;
  assign n32742 = n32738 & ~n32741 ;
  assign n32743 = x8 & n2331 ;
  assign n32744 = ~n2331 & n32743 ;
  assign n32745 = n8687 & ~n32744 ;
  assign n32746 = n32744 & n32745 ;
  assign n32747 = n32742 | n32746 ;
  assign n32757 = n32756 ^ n32747 ^ 1'b0 ;
  assign n32758 = n2980 & n32757 ;
  assign n32759 = n2757 & ~n16213 ;
  assign n32760 = n1380 & n5259 ;
  assign n32761 = n32760 ^ n34 ^ 1'b0 ;
  assign n32762 = n10581 ^ n2964 ^ 1'b0 ;
  assign n32763 = n3194 & n32762 ;
  assign n32764 = n5297 & ~n30109 ;
  assign n32765 = n32764 ^ n2070 ^ 1'b0 ;
  assign n32766 = n26227 ^ n10957 ^ 1'b0 ;
  assign n32767 = n32765 & ~n32766 ;
  assign n32768 = ~n8690 & n11578 ;
  assign n32769 = n20535 ^ n6698 ^ 1'b0 ;
  assign n32770 = n6198 | n18191 ;
  assign n32771 = n32770 ^ n14742 ^ n3859 ;
  assign n32772 = n9789 & n32771 ;
  assign n32773 = n26124 ^ n25289 ^ 1'b0 ;
  assign n32774 = n27835 & n32773 ;
  assign n32775 = n8236 | n24667 ;
  assign n32776 = n26041 & ~n32775 ;
  assign n32777 = n852 | n26385 ;
  assign n32778 = n7770 & ~n32777 ;
  assign n32779 = n32778 ^ n4613 ^ 1'b0 ;
  assign n32780 = ~n21599 & n32779 ;
  assign n32781 = n1649 | n25806 ;
  assign n32782 = ~n4668 & n32781 ;
  assign n32783 = n5736 & n10078 ;
  assign n32784 = n23295 ^ n8236 ^ 1'b0 ;
  assign n32785 = n5011 & ~n16216 ;
  assign n32786 = ~n2391 & n32785 ;
  assign n32787 = n6728 ^ n3378 ^ 1'b0 ;
  assign n32788 = n2128 & ~n6964 ;
  assign n32789 = n21982 | n32788 ;
  assign n32790 = n32789 ^ n3085 ^ 1'b0 ;
  assign n32791 = ~n8959 & n28866 ;
  assign n32792 = ~x3 & n32791 ;
  assign n32793 = n15237 ^ n2969 ^ 1'b0 ;
  assign n32794 = n2270 | n32793 ;
  assign n32795 = n32794 ^ n3484 ^ 1'b0 ;
  assign n32796 = n16243 ^ n4543 ^ 1'b0 ;
  assign n32797 = n4378 & ~n32796 ;
  assign n32798 = n3224 & n4600 ;
  assign n32799 = ~n32797 & n32798 ;
  assign n32800 = n4640 & ~n13886 ;
  assign n32801 = n144 | n1001 ;
  assign n32802 = n7069 ^ n839 ^ 1'b0 ;
  assign n32803 = n7110 & n32802 ;
  assign n32804 = ~n3559 & n32803 ;
  assign n32805 = n878 & ~n17330 ;
  assign n32806 = n32805 ^ n10534 ^ 1'b0 ;
  assign n32807 = n3139 ^ n1685 ^ 1'b0 ;
  assign n32808 = n14586 | n32807 ;
  assign n32811 = n1975 & ~n19064 ;
  assign n32810 = n1048 & n29214 ;
  assign n32812 = n32811 ^ n32810 ^ 1'b0 ;
  assign n32809 = ~n8482 & n21333 ;
  assign n32813 = n32812 ^ n32809 ^ 1'b0 ;
  assign n32814 = n19854 ^ n2012 ^ n1263 ;
  assign n32815 = n6325 & n32814 ;
  assign n32816 = ~n461 & n18566 ;
  assign n32817 = n32816 ^ n113 ^ 1'b0 ;
  assign n32818 = n32817 ^ n20249 ^ 1'b0 ;
  assign n32819 = n32351 & ~n32818 ;
  assign n32820 = n7596 ^ n5244 ^ 1'b0 ;
  assign n32821 = n7148 & ~n32820 ;
  assign n32822 = n31475 ^ n15327 ^ n10634 ;
  assign n32823 = n28063 ^ n16571 ^ 1'b0 ;
  assign n32824 = n32083 ^ n2494 ^ 1'b0 ;
  assign n32825 = n22338 ^ n2273 ^ 1'b0 ;
  assign n32826 = n330 | n5863 ;
  assign n32827 = n26600 & ~n32826 ;
  assign n32828 = ~n19 & n4577 ;
  assign n32829 = n10261 ^ n3549 ^ 1'b0 ;
  assign n32830 = n4511 & n32829 ;
  assign n32831 = n8990 | n14655 ;
  assign n32832 = n19475 ^ n8879 ^ 1'b0 ;
  assign n32833 = n52 & ~n32832 ;
  assign n32834 = n6933 & ~n8879 ;
  assign n32835 = n32834 ^ n7731 ^ 1'b0 ;
  assign n32836 = n6212 | n32835 ;
  assign n32837 = n6966 | n12810 ;
  assign n32838 = ~n32836 & n32837 ;
  assign n32839 = ~n9315 & n32838 ;
  assign n32840 = n23515 ^ n9410 ^ 1'b0 ;
  assign n32841 = n6849 & n26287 ;
  assign n32842 = ( ~n7134 & n7550 ) | ( ~n7134 & n18195 ) | ( n7550 & n18195 ) ;
  assign n32843 = n14455 & n32842 ;
  assign n32844 = ~n15241 & n25783 ;
  assign n32845 = n30009 & ~n32844 ;
  assign n32846 = ~n29056 & n32845 ;
  assign n32847 = n5823 & n27454 ;
  assign n32848 = n22267 & ~n32847 ;
  assign n32849 = ~n423 & n32848 ;
  assign n32850 = n5984 ^ n810 ^ 1'b0 ;
  assign n32851 = ~n2316 & n12511 ;
  assign n32852 = n475 & n32851 ;
  assign n32853 = ~n31219 & n32852 ;
  assign n32854 = ~n4396 & n9476 ;
  assign n32855 = n15576 ^ n5440 ^ 1'b0 ;
  assign n32856 = ~n1472 & n4327 ;
  assign n32857 = ~n6826 & n32856 ;
  assign n32858 = n159 | n10723 ;
  assign n32859 = n3210 | n32858 ;
  assign n32860 = n3262 | n8627 ;
  assign n32861 = n15077 ^ n7938 ^ 1'b0 ;
  assign n32862 = n5628 & n15680 ;
  assign n32863 = n32862 ^ n19333 ^ 1'b0 ;
  assign n32864 = n8771 & n32863 ;
  assign n32865 = n6081 ^ n1307 ^ n639 ;
  assign n32866 = n32865 ^ n21989 ^ n17534 ;
  assign n32867 = n14185 & ~n32866 ;
  assign n32868 = n1133 & n25766 ;
  assign n32869 = n8467 ^ n5128 ^ 1'b0 ;
  assign n32870 = ~n5059 & n32869 ;
  assign n32871 = n9586 & ~n18415 ;
  assign n32872 = n9051 & ~n32871 ;
  assign n32873 = n14130 & ~n23888 ;
  assign n32874 = n32873 ^ n14536 ^ 1'b0 ;
  assign n32875 = ~n10106 & n16387 ;
  assign n32876 = n32875 ^ n20706 ^ 1'b0 ;
  assign n32877 = n908 | n4541 ;
  assign n32878 = n21209 ^ n7955 ^ 1'b0 ;
  assign n32879 = n22628 | n25392 ;
  assign n32881 = n10392 ^ n8822 ^ 1'b0 ;
  assign n32880 = n6039 & n7702 ;
  assign n32882 = n32881 ^ n32880 ^ 1'b0 ;
  assign n32883 = n32882 ^ n6567 ^ 1'b0 ;
  assign n32884 = n1135 & n5370 ;
  assign n32885 = ~n16538 & n32884 ;
  assign n32886 = n12646 ^ n12463 ^ n12002 ;
  assign n32887 = n9354 & ~n17021 ;
  assign n32888 = n6842 & ~n25803 ;
  assign n32889 = ~n27649 & n32888 ;
  assign n32890 = ~n5779 & n7061 ;
  assign n32891 = n20336 ^ n3074 ^ 1'b0 ;
  assign n32892 = n1415 & n32891 ;
  assign n32893 = n8883 | n10427 ;
  assign n32894 = ~n4885 & n7250 ;
  assign n32895 = ~n4504 & n32894 ;
  assign n32896 = ~n12694 & n22897 ;
  assign n32897 = n32896 ^ n2270 ^ 1'b0 ;
  assign n32898 = n3477 & ~n21539 ;
  assign n32899 = ~n32897 & n32898 ;
  assign n32900 = ~n793 & n11548 ;
  assign n32901 = n5256 | n8639 ;
  assign n32902 = n13554 & n32901 ;
  assign n32903 = n32902 ^ n928 ^ 1'b0 ;
  assign n32904 = n24097 ^ n4117 ^ 1'b0 ;
  assign n32905 = n10637 & n32904 ;
  assign n32906 = ~n7641 & n18028 ;
  assign n32907 = ~n4835 & n9424 ;
  assign n32908 = ( n23980 & n24909 ) | ( n23980 & ~n32907 ) | ( n24909 & ~n32907 ) ;
  assign n32909 = n30271 ^ n16403 ^ 1'b0 ;
  assign n32910 = n16193 ^ n6444 ^ 1'b0 ;
  assign n32911 = n7998 | n12065 ;
  assign n32912 = n207 & n32911 ;
  assign n32913 = n5102 ^ n5045 ^ 1'b0 ;
  assign n32914 = n10606 & ~n32913 ;
  assign n32915 = n32914 ^ n3988 ^ 1'b0 ;
  assign n32916 = n4273 & n8525 ;
  assign n32917 = ( n29017 & ~n32915 ) | ( n29017 & n32916 ) | ( ~n32915 & n32916 ) ;
  assign n32918 = ~n32912 & n32917 ;
  assign n32919 = n7977 ^ n1193 ^ 1'b0 ;
  assign n32920 = ~n1842 & n32919 ;
  assign n32921 = n28935 | n30884 ;
  assign n32922 = n677 | n10252 ;
  assign n32923 = ( n15698 & n25241 ) | ( n15698 & ~n32922 ) | ( n25241 & ~n32922 ) ;
  assign n32924 = n2278 | n2486 ;
  assign n32925 = n32924 ^ n8876 ^ 1'b0 ;
  assign n32926 = n662 & ~n8915 ;
  assign n32927 = n1192 & n15435 ;
  assign n32928 = n7715 & n32927 ;
  assign n32929 = n32926 & n32928 ;
  assign n32930 = n32616 ^ n22080 ^ 1'b0 ;
  assign n32931 = ~n2404 & n20007 ;
  assign n32932 = n15811 & n32931 ;
  assign n32933 = n22228 & n32932 ;
  assign n32934 = n5905 & n24002 ;
  assign n32935 = ( n766 & n19758 ) | ( n766 & ~n22134 ) | ( n19758 & ~n22134 ) ;
  assign n32936 = n8109 & n32935 ;
  assign n32937 = ~n11413 & n29997 ;
  assign n32938 = n32937 ^ n37 ^ 1'b0 ;
  assign n32939 = n8077 & n10886 ;
  assign n32940 = n18205 & n25595 ;
  assign n32941 = n32940 ^ n3744 ^ 1'b0 ;
  assign n32942 = n14392 | n29475 ;
  assign n32943 = n2712 & ~n19544 ;
  assign n32944 = n4131 & n32943 ;
  assign n32945 = n1370 | n12381 ;
  assign n32946 = n2164 | n32945 ;
  assign n32947 = n32946 ^ n16752 ^ 1'b0 ;
  assign n32948 = n68 | n7264 ;
  assign n32949 = n2969 ^ n75 ^ 1'b0 ;
  assign n32950 = ( n5431 & n32948 ) | ( n5431 & ~n32949 ) | ( n32948 & ~n32949 ) ;
  assign n32951 = n32950 ^ n16010 ^ 1'b0 ;
  assign n32952 = ( ~n4258 & n15532 ) | ( ~n4258 & n19294 ) | ( n15532 & n19294 ) ;
  assign n32953 = n12487 | n15810 ;
  assign n32954 = ~n2397 & n11824 ;
  assign n32955 = n9544 & ~n32954 ;
  assign n32956 = n6144 & n10212 ;
  assign n32957 = ~n3346 & n13853 ;
  assign n32958 = ~n4591 & n32957 ;
  assign n32959 = n31087 ^ n102 ^ 1'b0 ;
  assign n32960 = n460 & n32959 ;
  assign n32961 = n23778 ^ n13800 ^ 1'b0 ;
  assign n32962 = n17988 ^ n13766 ^ 1'b0 ;
  assign n32963 = n601 & ~n2973 ;
  assign n32964 = n14182 | n21106 ;
  assign n32965 = n29276 | n32964 ;
  assign n32966 = ~n21112 & n32965 ;
  assign n32967 = n3067 & n32966 ;
  assign n32968 = n1491 | n21647 ;
  assign n32969 = n2107 & ~n7319 ;
  assign n32970 = ~n1191 & n9401 ;
  assign n32971 = n32970 ^ n30332 ^ 1'b0 ;
  assign n32972 = n15430 | n32143 ;
  assign n32973 = n6529 ^ n3674 ^ 1'b0 ;
  assign n32974 = n6454 ^ n535 ^ 1'b0 ;
  assign n32975 = n8457 & ~n12557 ;
  assign n32976 = n8312 & ~n27610 ;
  assign n32977 = n32976 ^ n29901 ^ 1'b0 ;
  assign n32978 = n197 & n32977 ;
  assign n32979 = ~n5758 & n11803 ;
  assign n32980 = n1878 & n6277 ;
  assign n32981 = n517 & n32980 ;
  assign n32982 = n27399 | n32981 ;
  assign n32983 = n7059 ^ n6046 ^ 1'b0 ;
  assign n32984 = ~n14646 & n32983 ;
  assign n32985 = ( n488 & n832 ) | ( n488 & n15672 ) | ( n832 & n15672 ) ;
  assign n32987 = ~n3251 & n25828 ;
  assign n32986 = n7579 & n11913 ;
  assign n32988 = n32987 ^ n32986 ^ 1'b0 ;
  assign n32990 = n1732 | n8226 ;
  assign n32989 = n13795 & n31109 ;
  assign n32991 = n32990 ^ n32989 ^ 1'b0 ;
  assign n32994 = n4294 ^ n835 ^ 1'b0 ;
  assign n32995 = ~n9158 & n32994 ;
  assign n32992 = ~n6212 & n16491 ;
  assign n32993 = n4453 | n32992 ;
  assign n32996 = n32995 ^ n32993 ^ 1'b0 ;
  assign n32997 = n8228 & ~n32996 ;
  assign n32998 = n19446 ^ n817 ^ 1'b0 ;
  assign n32999 = n1901 & n25457 ;
  assign n33000 = ( n8893 & ~n14551 ) | ( n8893 & n20131 ) | ( ~n14551 & n20131 ) ;
  assign n33001 = n11089 | n33000 ;
  assign n33002 = n14493 ^ n6492 ^ 1'b0 ;
  assign n33003 = n934 & n5113 ;
  assign n33004 = ~n2062 & n33003 ;
  assign n33005 = n9551 | n17239 ;
  assign n33006 = n33005 ^ n13834 ^ 1'b0 ;
  assign n33007 = n3853 & n10603 ;
  assign n33008 = n25789 ^ n116 ^ 1'b0 ;
  assign n33009 = n4830 & ~n8033 ;
  assign n33010 = n33009 ^ n1558 ^ 1'b0 ;
  assign n33011 = n10833 ^ n10175 ^ 1'b0 ;
  assign n33012 = ~n497 & n15625 ;
  assign n33013 = n30654 ^ n12932 ^ 1'b0 ;
  assign n33014 = n178 & ~n3051 ;
  assign n33015 = ~n33013 & n33014 ;
  assign n33016 = n20727 | n33015 ;
  assign n33017 = n4520 & ~n31353 ;
  assign n33018 = n3739 & ~n27158 ;
  assign n33019 = n14217 & ~n33018 ;
  assign n33020 = n33019 ^ n32770 ^ 1'b0 ;
  assign n33021 = n29973 ^ n1193 ^ 1'b0 ;
  assign n33022 = n9983 | n33021 ;
  assign n33023 = n2209 | n15526 ;
  assign n33024 = n8403 & ~n11916 ;
  assign n33025 = n4930 & n33024 ;
  assign n33026 = n24097 ^ n21418 ^ 1'b0 ;
  assign n33027 = ~n11167 & n13695 ;
  assign n33028 = ~n4967 & n27973 ;
  assign n33029 = n33028 ^ n11027 ^ 1'b0 ;
  assign n33030 = n17845 & ~n33029 ;
  assign n33031 = n2414 | n17360 ;
  assign n33032 = n33030 | n33031 ;
  assign n33033 = n22634 ^ n18556 ^ 1'b0 ;
  assign n33034 = n21476 ^ n10242 ^ 1'b0 ;
  assign n33035 = n27829 & ~n33034 ;
  assign n33036 = n33035 ^ n17029 ^ 1'b0 ;
  assign n33037 = n1463 & n18977 ;
  assign n33038 = n33037 ^ n9788 ^ 1'b0 ;
  assign n33039 = n8927 & ~n26305 ;
  assign n33040 = n20541 ^ n7179 ^ 1'b0 ;
  assign n33041 = n21843 ^ n9831 ^ 1'b0 ;
  assign n33042 = n3367 ^ n1937 ^ 1'b0 ;
  assign n33043 = n7850 ^ n3866 ^ 1'b0 ;
  assign n33044 = ~n5769 & n33043 ;
  assign n33045 = n26188 | n33044 ;
  assign n33046 = n18351 ^ n16656 ^ 1'b0 ;
  assign n33047 = n24532 ^ n10303 ^ 1'b0 ;
  assign n33048 = n962 | n10867 ;
  assign n33049 = n21237 ^ n5532 ^ 1'b0 ;
  assign n33050 = n33048 | n33049 ;
  assign n33051 = n31801 ^ n8446 ^ 1'b0 ;
  assign n33052 = n33051 ^ n31035 ^ 1'b0 ;
  assign n33053 = n3481 & ~n6081 ;
  assign n33054 = ~n4027 & n33053 ;
  assign n33055 = n24859 & n33054 ;
  assign n33056 = n1968 | n3679 ;
  assign n33057 = n20101 | n33056 ;
  assign n33058 = n33057 ^ n17839 ^ 1'b0 ;
  assign n33059 = n26283 ^ n10261 ^ 1'b0 ;
  assign n33060 = ~n6653 & n18874 ;
  assign n33061 = n10399 ^ n6170 ^ 1'b0 ;
  assign n33062 = ~n33060 & n33061 ;
  assign n33063 = n33059 | n33062 ;
  assign n33064 = n2572 & n20334 ;
  assign n33065 = ~n8763 & n33064 ;
  assign n33066 = n7455 & n33065 ;
  assign n33067 = n10891 | n27406 ;
  assign n33068 = n18564 ^ n484 ^ 1'b0 ;
  assign n33069 = n6277 & ~n33068 ;
  assign n33070 = n20848 & n33069 ;
  assign n33071 = n23848 ^ n1087 ^ 1'b0 ;
  assign n33072 = n5551 & n22580 ;
  assign n33073 = n633 ^ n315 ^ 1'b0 ;
  assign n33074 = n12489 ^ n9409 ^ 1'b0 ;
  assign n33075 = n13690 ^ n254 ^ 1'b0 ;
  assign n33076 = n4088 & n21993 ;
  assign n33077 = ~n1144 & n33076 ;
  assign n33078 = n9576 & n33077 ;
  assign n33079 = n33078 ^ n11061 ^ 1'b0 ;
  assign n33080 = ~n5655 & n33079 ;
  assign n33081 = n10243 & ~n12063 ;
  assign n33082 = ~n28137 & n33081 ;
  assign n33083 = n18590 & ~n33082 ;
  assign n33084 = n5135 & n13843 ;
  assign n33085 = n13101 | n19606 ;
  assign n33086 = n33084 & ~n33085 ;
  assign n33087 = n11929 | n33086 ;
  assign n33088 = n16007 & n33087 ;
  assign n33089 = n3836 & ~n33088 ;
  assign n33090 = n33083 | n33089 ;
  assign n33091 = n14258 ^ n3512 ^ 1'b0 ;
  assign n33092 = n20761 & ~n33091 ;
  assign n33093 = n5617 | n17561 ;
  assign n33094 = n1054 & n9058 ;
  assign n33095 = n25815 & n33094 ;
  assign n33096 = n33093 & n33095 ;
  assign n33097 = n7301 & ~n10386 ;
  assign n33098 = n33097 ^ n22112 ^ 1'b0 ;
  assign n33099 = n5749 & n33098 ;
  assign n33100 = n33099 ^ n7612 ^ 1'b0 ;
  assign n33101 = n11323 ^ n10649 ^ 1'b0 ;
  assign n33102 = n9092 | n12211 ;
  assign n33103 = n13469 & n33102 ;
  assign n33104 = n4748 | n28165 ;
  assign n33105 = n33104 ^ n22096 ^ 1'b0 ;
  assign n33106 = n14057 ^ n4153 ^ 1'b0 ;
  assign n33107 = ~n5273 & n33106 ;
  assign n33108 = n8553 ^ n236 ^ 1'b0 ;
  assign n33109 = ~n16475 & n31624 ;
  assign n33110 = n2693 | n26061 ;
  assign n33111 = n4986 | n26051 ;
  assign n33112 = n6759 & ~n33111 ;
  assign n33113 = n21875 & n33112 ;
  assign n33114 = ~n6325 & n14874 ;
  assign n33115 = n18865 | n25223 ;
  assign n33116 = n11119 ^ n4330 ^ 1'b0 ;
  assign n33117 = n33115 & n33116 ;
  assign n33118 = ~n128 & n3606 ;
  assign n33119 = ~n216 & n33118 ;
  assign n33120 = n33119 ^ n25630 ^ n5286 ;
  assign n33121 = n2072 ^ n1227 ^ 1'b0 ;
  assign n33122 = n104 & ~n33121 ;
  assign n33123 = n9275 & n16052 ;
  assign n33124 = n1676 & n33123 ;
  assign n33125 = n33122 & n33124 ;
  assign n33126 = n13196 | n33125 ;
  assign n33127 = n4133 & ~n19618 ;
  assign n33128 = n10066 ^ n7227 ^ 1'b0 ;
  assign n33129 = ~n6974 & n33128 ;
  assign n33130 = n18975 & n33129 ;
  assign n33131 = ~n33127 & n33130 ;
  assign n33132 = n33126 & ~n33131 ;
  assign n33133 = n5053 & ~n25839 ;
  assign n33134 = n20250 & n33133 ;
  assign n33135 = n596 | n14750 ;
  assign n33136 = n33134 & ~n33135 ;
  assign n33137 = n23449 ^ n14074 ^ 1'b0 ;
  assign n33138 = ~n8886 & n33137 ;
  assign n33139 = n2148 & ~n8838 ;
  assign n33140 = n814 & ~n1117 ;
  assign n33141 = n4415 ^ n452 ^ 1'b0 ;
  assign n33142 = ~n4508 & n33141 ;
  assign n33143 = ~n12678 & n33142 ;
  assign n33144 = ~n33140 & n33143 ;
  assign n33145 = ~n1083 & n15495 ;
  assign n33146 = ~n20782 & n23463 ;
  assign n33147 = n4956 ^ n4181 ^ 1'b0 ;
  assign n33148 = n28968 & n33147 ;
  assign n33149 = n7113 | n16189 ;
  assign n33150 = n33148 | n33149 ;
  assign n33151 = n33150 ^ n23636 ^ 1'b0 ;
  assign n33152 = n15670 ^ n2155 ^ 1'b0 ;
  assign n33153 = n7097 & n33152 ;
  assign n33155 = n21078 ^ n18937 ^ 1'b0 ;
  assign n33154 = n13929 & n20325 ;
  assign n33156 = n33155 ^ n33154 ^ 1'b0 ;
  assign n33157 = n3297 & ~n21412 ;
  assign n33158 = ~n21535 & n30880 ;
  assign n33159 = n33158 ^ n16822 ^ 1'b0 ;
  assign n33160 = n17963 & n29326 ;
  assign n33161 = n7952 | n14926 ;
  assign n33162 = n33088 ^ n10144 ^ 1'b0 ;
  assign n33163 = n33161 | n33162 ;
  assign n33165 = n9209 ^ n6224 ^ 1'b0 ;
  assign n33164 = ~n462 & n11800 ;
  assign n33166 = n33165 ^ n33164 ^ 1'b0 ;
  assign n33167 = n3534 & n9273 ;
  assign n33168 = ~n9273 & n33167 ;
  assign n33169 = n5760 & n29315 ;
  assign n33170 = ~n3189 & n4510 ;
  assign n33171 = ~n4510 & n33170 ;
  assign n33172 = n33171 ^ n6552 ^ 1'b0 ;
  assign n33173 = ~n28018 & n33172 ;
  assign n33174 = n1702 & n33173 ;
  assign n33175 = n1648 & n33174 ;
  assign n33176 = n33169 | n33175 ;
  assign n33177 = n33168 & ~n33176 ;
  assign n33178 = n15441 ^ n2062 ^ 1'b0 ;
  assign n33179 = n3514 ^ n1367 ^ 1'b0 ;
  assign n33180 = n30154 & ~n33179 ;
  assign n33181 = n919 | n20099 ;
  assign n33182 = n6642 & ~n17205 ;
  assign n33183 = n33182 ^ n19076 ^ 1'b0 ;
  assign n33184 = ~n8601 & n16570 ;
  assign n33185 = n33184 ^ n6078 ^ 1'b0 ;
  assign n33186 = n31919 | n33185 ;
  assign n33187 = n33186 ^ n2534 ^ 1'b0 ;
  assign n33188 = n11090 ^ n2124 ^ 1'b0 ;
  assign n33189 = n982 & n33188 ;
  assign n33190 = ( ~n12536 & n32632 ) | ( ~n12536 & n33189 ) | ( n32632 & n33189 ) ;
  assign n33191 = n10599 & ~n33190 ;
  assign n33192 = n27463 ^ n4791 ^ 1'b0 ;
  assign n33193 = n246 | n3864 ;
  assign n33194 = n33193 ^ n32079 ^ 1'b0 ;
  assign n33195 = n6527 ^ n1159 ^ 1'b0 ;
  assign n33196 = n17477 & n33195 ;
  assign n33197 = n13901 & ~n24598 ;
  assign n33198 = n20770 & ~n33197 ;
  assign n33199 = ~n22132 & n33198 ;
  assign n33200 = n10133 & n16669 ;
  assign n33201 = n12331 ^ n1658 ^ 1'b0 ;
  assign n33202 = n22426 & n33201 ;
  assign n33203 = n33202 ^ n7780 ^ 1'b0 ;
  assign n33204 = ~n33200 & n33203 ;
  assign n33205 = n4862 | n5004 ;
  assign n33206 = n33205 ^ n4668 ^ 1'b0 ;
  assign n33207 = n3861 & ~n33206 ;
  assign n33208 = n33207 ^ n29097 ^ 1'b0 ;
  assign n33209 = n1212 & ~n30477 ;
  assign n33210 = n33209 ^ n828 ^ 1'b0 ;
  assign n33211 = n22186 ^ n1438 ^ 1'b0 ;
  assign n33212 = ~n33210 & n33211 ;
  assign n33213 = n3193 & n11228 ;
  assign n33214 = n33213 ^ n28970 ^ 1'b0 ;
  assign n33215 = n6039 | n17834 ;
  assign n33216 = n33214 & ~n33215 ;
  assign n33217 = ~n7811 & n15847 ;
  assign n33218 = n26339 & n33217 ;
  assign n33219 = n20610 & ~n33218 ;
  assign n33220 = n3032 & ~n25179 ;
  assign n33221 = n33220 ^ n13456 ^ 1'b0 ;
  assign n33222 = n32685 ^ n20672 ^ 1'b0 ;
  assign n33223 = n12109 ^ n11578 ^ n5575 ;
  assign n33224 = ~n8209 & n8495 ;
  assign n33225 = n33224 ^ n11390 ^ 1'b0 ;
  assign n33226 = n9082 | n18793 ;
  assign n33227 = n2627 & ~n12255 ;
  assign n33228 = n11049 & n31837 ;
  assign n33229 = n33228 ^ n25764 ^ 1'b0 ;
  assign n33230 = n24077 ^ n2203 ^ 1'b0 ;
  assign n33231 = n33230 ^ n25806 ^ 1'b0 ;
  assign n33232 = n9718 ^ n2607 ^ 1'b0 ;
  assign n33234 = n14697 ^ n10950 ^ 1'b0 ;
  assign n33233 = ~n244 & n7510 ;
  assign n33235 = n33234 ^ n33233 ^ 1'b0 ;
  assign n33236 = n940 & n3423 ;
  assign n33237 = n26224 & ~n32940 ;
  assign n33238 = n7315 ^ n339 ^ 1'b0 ;
  assign n33239 = ~n4485 & n33238 ;
  assign n33240 = n33239 ^ n158 ^ 1'b0 ;
  assign n33241 = n12054 ^ n4966 ^ 1'b0 ;
  assign n33242 = n31418 ^ n21651 ^ 1'b0 ;
  assign n33243 = n1565 & n4350 ;
  assign n33244 = n33242 & ~n33243 ;
  assign n33245 = ~n316 & n1480 ;
  assign n33246 = n11394 & ~n33245 ;
  assign n33247 = n10216 & ~n33246 ;
  assign n33248 = n2862 & ~n33247 ;
  assign n33249 = n15752 ^ n15200 ^ 1'b0 ;
  assign n33250 = ~n30442 & n33249 ;
  assign n33251 = ~n982 & n33250 ;
  assign n33252 = n19178 ^ n5269 ^ 1'b0 ;
  assign n33253 = n7898 ^ n2344 ^ 1'b0 ;
  assign n33254 = n8046 & ~n33253 ;
  assign n33255 = n3744 & n19875 ;
  assign n33256 = n22981 | n33255 ;
  assign n33257 = n20618 | n33256 ;
  assign n33258 = n33254 | n33257 ;
  assign n33260 = ~n387 & n5226 ;
  assign n33261 = n33260 ^ n14123 ^ 1'b0 ;
  assign n33262 = n9552 & n33261 ;
  assign n33259 = n408 | n3776 ;
  assign n33263 = n33262 ^ n33259 ^ 1'b0 ;
  assign n33264 = n9084 ^ n7192 ^ 1'b0 ;
  assign n33265 = n33264 ^ n22551 ^ 1'b0 ;
  assign n33266 = n2269 ^ n1425 ^ 1'b0 ;
  assign n33267 = n33266 ^ n9898 ^ n4350 ;
  assign n33269 = n1571 ^ n397 ^ 1'b0 ;
  assign n33270 = n29465 & n33269 ;
  assign n33268 = n1458 & n16621 ;
  assign n33271 = n33270 ^ n33268 ^ 1'b0 ;
  assign n33272 = n17958 ^ n16122 ^ 1'b0 ;
  assign n33273 = n11336 ^ n3116 ^ 1'b0 ;
  assign n33274 = n794 & ~n33273 ;
  assign n33275 = ~n3054 & n33274 ;
  assign n33276 = n6062 ^ n839 ^ 1'b0 ;
  assign n33277 = ~n3690 & n33276 ;
  assign n33278 = n12293 & ~n33277 ;
  assign n33279 = n8479 | n33278 ;
  assign n33280 = n33278 & ~n33279 ;
  assign n33281 = n33280 ^ n11336 ^ 1'b0 ;
  assign n33282 = n4816 & ~n6055 ;
  assign n33283 = n10005 ^ n142 ^ 1'b0 ;
  assign n33284 = n5172 & n33283 ;
  assign n33285 = ~n4720 & n33284 ;
  assign n33286 = n28979 ^ n12422 ^ n12310 ;
  assign n33287 = n6466 ^ n917 ^ 1'b0 ;
  assign n33288 = n18460 | n33287 ;
  assign n33289 = n33286 & ~n33288 ;
  assign n33290 = n382 | n25457 ;
  assign n33291 = n33290 ^ n16349 ^ 1'b0 ;
  assign n33292 = n23753 & ~n31655 ;
  assign n33293 = n15435 & n21973 ;
  assign n33294 = n6063 & ~n9931 ;
  assign n33295 = n15111 ^ n14062 ^ 1'b0 ;
  assign n33296 = n33294 & n33295 ;
  assign n33297 = ( ~n13470 & n21221 ) | ( ~n13470 & n33296 ) | ( n21221 & n33296 ) ;
  assign n33298 = n15707 ^ n14879 ^ 1'b0 ;
  assign n33299 = n12242 | n33298 ;
  assign n33300 = n27466 | n33299 ;
  assign n33301 = n23052 ^ n139 ^ 1'b0 ;
  assign n33302 = n13795 & ~n17621 ;
  assign n33303 = ~n28712 & n33302 ;
  assign n33304 = n25689 ^ n3925 ^ 1'b0 ;
  assign n33305 = n17500 ^ n17297 ^ 1'b0 ;
  assign n33306 = n3640 | n9570 ;
  assign n33307 = n15820 | n33306 ;
  assign n33308 = n8941 & n33307 ;
  assign n33309 = n7812 & n33308 ;
  assign n33310 = n6332 ^ n4586 ^ 1'b0 ;
  assign n33311 = n5373 & ~n33310 ;
  assign n33312 = n31686 ^ n25812 ^ 1'b0 ;
  assign n33313 = ~n13869 & n33312 ;
  assign n33314 = n7610 & n33313 ;
  assign n33315 = n14105 & ~n33314 ;
  assign n33316 = n5942 & ~n28311 ;
  assign n33317 = ~n2242 & n21748 ;
  assign n33318 = n27783 & n28194 ;
  assign n33319 = n17241 | n32635 ;
  assign n33322 = n3063 & n3656 ;
  assign n33323 = n33322 ^ n484 ^ 1'b0 ;
  assign n33321 = n113 & ~n13532 ;
  assign n33324 = n33323 ^ n33321 ^ 1'b0 ;
  assign n33320 = ~n3579 & n20342 ;
  assign n33325 = n33324 ^ n33320 ^ 1'b0 ;
  assign n33326 = n8283 ^ n937 ^ 1'b0 ;
  assign n33327 = n20578 ^ n2308 ^ 1'b0 ;
  assign n33328 = n2761 | n27215 ;
  assign n33329 = n33327 & ~n33328 ;
  assign n33330 = n16730 & ~n33329 ;
  assign n33331 = n4760 & n33330 ;
  assign n33332 = n2307 & ~n33331 ;
  assign n33333 = n13453 ^ n2136 ^ 1'b0 ;
  assign n33334 = n33333 ^ n2482 ^ 1'b0 ;
  assign n33335 = ~n436 & n8429 ;
  assign n33336 = ~n19231 & n33335 ;
  assign n33337 = ( n4156 & ~n6644 ) | ( n4156 & n22219 ) | ( ~n6644 & n22219 ) ;
  assign n33338 = ( n4383 & n5725 ) | ( n4383 & n23972 ) | ( n5725 & n23972 ) ;
  assign n33339 = n5068 | n33338 ;
  assign n33340 = n30 | n33339 ;
  assign n33341 = n23306 ^ n14317 ^ 1'b0 ;
  assign n33342 = n4394 & n33341 ;
  assign n33343 = n11277 | n30144 ;
  assign n33344 = n33342 & ~n33343 ;
  assign n33345 = ~n6903 & n33344 ;
  assign n33346 = n7782 | n11583 ;
  assign n33347 = n33346 ^ n17876 ^ 1'b0 ;
  assign n33348 = n3593 | n33347 ;
  assign n33349 = n33348 ^ n3037 ^ 1'b0 ;
  assign n33350 = n2690 | n32713 ;
  assign n33351 = n4710 | n12466 ;
  assign n33352 = ~n24347 & n26617 ;
  assign n33353 = ~n14226 & n33352 ;
  assign n33354 = n24466 ^ n6375 ^ 1'b0 ;
  assign n33355 = n8025 & ~n33354 ;
  assign n33356 = n415 ^ n257 ^ 1'b0 ;
  assign n33357 = n25783 ^ n3385 ^ 1'b0 ;
  assign n33358 = n3138 & ~n16027 ;
  assign n33359 = n33358 ^ n8452 ^ 1'b0 ;
  assign n33360 = n6884 & ~n33359 ;
  assign n33361 = n12404 ^ n9821 ^ 1'b0 ;
  assign n33362 = n9201 ^ n158 ^ 1'b0 ;
  assign n33363 = n15536 ^ n1766 ^ 1'b0 ;
  assign n33364 = ~n2128 & n33363 ;
  assign n33365 = n17923 ^ n229 ^ 1'b0 ;
  assign n33366 = n33365 ^ n23389 ^ n4747 ;
  assign n33367 = n14479 & ~n18026 ;
  assign n33368 = n28424 & ~n33367 ;
  assign n33369 = n6552 ^ n4324 ^ 1'b0 ;
  assign n33370 = n6653 & n20099 ;
  assign n33371 = ~n6926 & n22338 ;
  assign n33372 = ~n22338 & n33371 ;
  assign n33373 = n33370 & ~n33372 ;
  assign n33374 = ~n33370 & n33373 ;
  assign n33375 = n20367 | n33374 ;
  assign n33376 = n33374 & ~n33375 ;
  assign n33377 = n3452 | n6853 ;
  assign n33378 = n23455 & ~n25222 ;
  assign n33379 = n33378 ^ n7160 ^ 1'b0 ;
  assign n33380 = n22702 ^ n13080 ^ 1'b0 ;
  assign n33381 = n627 & n6106 ;
  assign n33382 = n33381 ^ n2571 ^ 1'b0 ;
  assign n33383 = n20326 ^ n16853 ^ 1'b0 ;
  assign n33384 = n7700 & ~n8994 ;
  assign n33385 = n6581 & ~n17479 ;
  assign n33386 = n7603 & n33385 ;
  assign n33387 = n20576 ^ n1245 ^ 1'b0 ;
  assign n33388 = n33386 | n33387 ;
  assign n33389 = n14830 ^ n6647 ^ 1'b0 ;
  assign n33390 = n8226 & n33389 ;
  assign n33391 = n6022 ^ n1390 ^ 1'b0 ;
  assign n33392 = n22941 ^ n8351 ^ 1'b0 ;
  assign n33393 = n542 & n2780 ;
  assign n33394 = n25790 ^ n2386 ^ 1'b0 ;
  assign n33395 = n8250 & n33394 ;
  assign n33396 = n8325 ^ n5892 ^ 1'b0 ;
  assign n33397 = ~n22233 & n33396 ;
  assign n33398 = n33397 ^ n18845 ^ 1'b0 ;
  assign n33399 = n19661 ^ n4906 ^ 1'b0 ;
  assign n33400 = ~n10746 & n33399 ;
  assign n33401 = n9903 & ~n33400 ;
  assign n33402 = n15458 | n19049 ;
  assign n33403 = n15072 | n25497 ;
  assign n33404 = n17755 | n33403 ;
  assign n33405 = n16947 & n21023 ;
  assign n33406 = n10105 & n33405 ;
  assign n33407 = n24396 | n33406 ;
  assign n33408 = ( n1739 & ~n2752 ) | ( n1739 & n14066 ) | ( ~n2752 & n14066 ) ;
  assign n33409 = n9881 | n33408 ;
  assign n33410 = n3985 | n33409 ;
  assign n33411 = n46 & n33410 ;
  assign n33412 = n12339 ^ n3423 ^ 1'b0 ;
  assign n33413 = n31520 ^ n1217 ^ 1'b0 ;
  assign n33414 = n10780 & n33413 ;
  assign n33415 = n8081 ^ n7033 ^ 1'b0 ;
  assign n33416 = n7619 ^ n1867 ^ 1'b0 ;
  assign n33417 = n33415 | n33416 ;
  assign n33418 = ~n1172 & n2818 ;
  assign n33419 = ~n290 & n33418 ;
  assign n33420 = n23617 ^ n22418 ^ 1'b0 ;
  assign n33421 = n28757 ^ n25302 ^ 1'b0 ;
  assign n33422 = n30678 ^ n4015 ^ 1'b0 ;
  assign n33423 = n129 & ~n3779 ;
  assign n33424 = n33423 ^ n4320 ^ 1'b0 ;
  assign n33425 = n33422 & n33424 ;
  assign n33426 = n5733 | n13183 ;
  assign n33427 = n32580 ^ n18963 ^ 1'b0 ;
  assign n33428 = ~n5590 & n6011 ;
  assign n33429 = n545 & ~n16617 ;
  assign n33430 = n33429 ^ n7048 ^ 1'b0 ;
  assign n33431 = n32099 ^ n15200 ^ 1'b0 ;
  assign n33432 = n172 & n11691 ;
  assign n33433 = ~n7373 & n33432 ;
  assign n33434 = n7596 | n7626 ;
  assign n33435 = n4811 & ~n5443 ;
  assign n33436 = n2460 | n10916 ;
  assign n33437 = n119 | n8079 ;
  assign n33438 = n11806 & ~n33437 ;
  assign n33439 = n10992 | n33438 ;
  assign n33440 = n33439 ^ n9745 ^ 1'b0 ;
  assign n33441 = n22924 ^ n12236 ^ n5607 ;
  assign n33442 = n25589 | n33441 ;
  assign n33443 = n33440 | n33442 ;
  assign n33444 = n11317 ^ n9742 ^ 1'b0 ;
  assign n33445 = n2951 & ~n33444 ;
  assign n33446 = ~n11438 & n33445 ;
  assign n33447 = n20576 & n33446 ;
  assign n33448 = n10548 ^ n35 ^ 1'b0 ;
  assign n33449 = n33448 ^ n4344 ^ 1'b0 ;
  assign n33450 = n7310 ^ n2644 ^ 1'b0 ;
  assign n33451 = n2141 | n33450 ;
  assign n33452 = n16322 | n33451 ;
  assign n33453 = n1927 & n16291 ;
  assign n33454 = ~n13470 & n33453 ;
  assign n33455 = n26713 ^ n17973 ^ 1'b0 ;
  assign n33456 = n2825 & ~n19416 ;
  assign n33457 = n13108 ^ n8040 ^ 1'b0 ;
  assign n33458 = ~n23267 & n28903 ;
  assign n33459 = ~n12213 & n30895 ;
  assign n33460 = n33459 ^ n8958 ^ 1'b0 ;
  assign n33461 = n10430 ^ n3401 ^ 1'b0 ;
  assign n33462 = n33461 ^ n31468 ^ 1'b0 ;
  assign n33463 = n6281 | n33462 ;
  assign n33465 = n2943 & n5194 ;
  assign n33466 = n3724 & n33465 ;
  assign n33464 = n5917 | n21066 ;
  assign n33467 = n33466 ^ n33464 ^ 1'b0 ;
  assign n33468 = n3371 | n33467 ;
  assign n33469 = n15266 ^ n4485 ^ 1'b0 ;
  assign n33470 = n657 | n9172 ;
  assign n33471 = ~n323 & n13266 ;
  assign n33472 = n6414 & n33471 ;
  assign n33473 = n30914 ^ n9322 ^ 1'b0 ;
  assign n33474 = n27864 & ~n28139 ;
  assign n33475 = n18252 ^ n16273 ^ 1'b0 ;
  assign n33476 = ~n7497 & n33475 ;
  assign n33477 = n430 | n4468 ;
  assign n33478 = n931 & ~n16604 ;
  assign n33479 = ~n33477 & n33478 ;
  assign n33480 = n850 | n33479 ;
  assign n33481 = n20472 & ~n33480 ;
  assign n33482 = n32972 & ~n33481 ;
  assign n33483 = n78 & n5876 ;
  assign n33484 = ~n17921 & n33483 ;
  assign n33485 = ( n9324 & n17879 ) | ( n9324 & n33484 ) | ( n17879 & n33484 ) ;
  assign n33486 = ~n10678 & n15511 ;
  assign n33487 = n11653 ^ n4944 ^ 1'b0 ;
  assign n33488 = ~n33486 & n33487 ;
  assign n33489 = n3409 | n14515 ;
  assign n33490 = n33489 ^ n886 ^ 1'b0 ;
  assign n33491 = n11235 ^ n6903 ^ 1'b0 ;
  assign n33492 = ~n29733 & n33491 ;
  assign n33493 = ~n9534 & n23747 ;
  assign n33494 = n13165 & n14192 ;
  assign n33495 = n33494 ^ n2727 ^ 1'b0 ;
  assign n33497 = n2152 & n11218 ;
  assign n33498 = n31750 & n33497 ;
  assign n33499 = n9120 | n33498 ;
  assign n33496 = n3633 | n25485 ;
  assign n33500 = n33499 ^ n33496 ^ 1'b0 ;
  assign n33501 = n33500 ^ n5721 ^ 1'b0 ;
  assign n33502 = n16029 | n30080 ;
  assign n33503 = n33502 ^ n2221 ^ 1'b0 ;
  assign n33504 = n33503 ^ n581 ^ 1'b0 ;
  assign n33505 = n2320 & n20468 ;
  assign n33506 = ( n24573 & n29175 ) | ( n24573 & ~n29994 ) | ( n29175 & ~n29994 ) ;
  assign n33507 = ~n9540 & n10383 ;
  assign n33508 = n1425 & ~n10548 ;
  assign n33509 = ~n33507 & n33508 ;
  assign n33510 = n767 & ~n14256 ;
  assign n33511 = n33510 ^ n9885 ^ 1'b0 ;
  assign n33512 = n6496 | n13875 ;
  assign n33513 = n33511 | n33512 ;
  assign n33514 = ~n1144 & n12944 ;
  assign n33515 = n568 & ~n11827 ;
  assign n33516 = n30198 ^ n6775 ^ 1'b0 ;
  assign n33517 = n17683 & n33516 ;
  assign n33518 = ~n3938 & n4964 ;
  assign n33519 = n616 & n33518 ;
  assign n33520 = n28134 & ~n33519 ;
  assign n33521 = n12450 ^ n5060 ^ 1'b0 ;
  assign n33522 = n33521 ^ n7800 ^ 1'b0 ;
  assign n33523 = n10870 ^ n3369 ^ 1'b0 ;
  assign n33524 = n17211 & ~n19106 ;
  assign n33525 = n4859 ^ n3443 ^ 1'b0 ;
  assign n33526 = n31736 | n33525 ;
  assign n33527 = n557 & n15896 ;
  assign n33528 = n18112 | n33527 ;
  assign n33529 = n20338 & ~n33528 ;
  assign n33530 = n13702 ^ n392 ^ 1'b0 ;
  assign n33531 = n33530 ^ n5603 ^ 1'b0 ;
  assign n33532 = n6633 ^ n3291 ^ 1'b0 ;
  assign n33533 = n5391 & ~n33532 ;
  assign n33534 = n33533 ^ n1370 ^ 1'b0 ;
  assign n33535 = n13408 & n19296 ;
  assign n33536 = n20612 & n33535 ;
  assign n33537 = n17940 ^ n685 ^ 1'b0 ;
  assign n33538 = ~n227 & n33537 ;
  assign n33539 = n627 | n2283 ;
  assign n33540 = n2424 & n24667 ;
  assign n33541 = ~n33539 & n33540 ;
  assign n33542 = n33541 ^ n27842 ^ 1'b0 ;
  assign n33544 = ~n4197 & n8685 ;
  assign n33545 = n15899 & n33544 ;
  assign n33543 = n6394 & n13962 ;
  assign n33546 = n33545 ^ n33543 ^ 1'b0 ;
  assign n33547 = n4629 & ~n19716 ;
  assign n33548 = n2769 & ~n10262 ;
  assign n33549 = ~n14776 & n33548 ;
  assign n33550 = n272 & n21085 ;
  assign n33551 = n9120 & n33550 ;
  assign n33552 = n33551 ^ n6706 ^ 1'b0 ;
  assign n33553 = n5225 | n16816 ;
  assign n33554 = n33552 | n33553 ;
  assign n33556 = n7231 & ~n7520 ;
  assign n33555 = ~n8312 & n9670 ;
  assign n33557 = n33556 ^ n33555 ^ 1'b0 ;
  assign n33558 = n8138 & ~n11850 ;
  assign n33559 = n13442 & n33558 ;
  assign n33560 = n677 & n4697 ;
  assign n33561 = n10459 & n33560 ;
  assign n33562 = ( n619 & ~n8128 ) | ( n619 & n21354 ) | ( ~n8128 & n21354 ) ;
  assign n33563 = n26110 ^ n10255 ^ 1'b0 ;
  assign n33564 = n5338 | n33563 ;
  assign n33565 = n26185 & n33564 ;
  assign n33566 = n15910 ^ n14549 ^ 1'b0 ;
  assign n33567 = n16326 & ~n25095 ;
  assign n33568 = n1345 & ~n33567 ;
  assign n33569 = n33568 ^ n2828 ^ 1'b0 ;
  assign n33570 = n16910 ^ n12681 ^ 1'b0 ;
  assign n33571 = n27574 & ~n33570 ;
  assign n33572 = n1254 | n6046 ;
  assign n33573 = n1790 & ~n33572 ;
  assign n33574 = n33573 ^ n9878 ^ 1'b0 ;
  assign n33575 = ~n7550 & n17072 ;
  assign n33576 = ~n26489 & n33575 ;
  assign n33577 = n707 | n33576 ;
  assign n33578 = n31877 ^ n4214 ^ 1'b0 ;
  assign n33580 = n19330 ^ n3475 ^ 1'b0 ;
  assign n33579 = n4328 & n31024 ;
  assign n33581 = n33580 ^ n33579 ^ 1'b0 ;
  assign n33582 = n9301 & n27687 ;
  assign n33583 = n33582 ^ n10360 ^ 1'b0 ;
  assign n33585 = n29687 ^ n20103 ^ 1'b0 ;
  assign n33584 = n6897 & ~n7698 ;
  assign n33586 = n33585 ^ n33584 ^ 1'b0 ;
  assign n33587 = n1531 & n30283 ;
  assign n33588 = ~n21304 & n33587 ;
  assign n33589 = n4742 & n33588 ;
  assign n33590 = n6865 & n31061 ;
  assign n33591 = ~n9341 & n10383 ;
  assign n33592 = n33591 ^ n25031 ^ 1'b0 ;
  assign n33593 = n30458 | n31738 ;
  assign n33594 = n6493 ^ n5652 ^ 1'b0 ;
  assign n33595 = x1 & n6664 ;
  assign n33596 = n5529 | n27568 ;
  assign n33597 = n18552 & ~n33596 ;
  assign n33598 = n11061 | n31509 ;
  assign n33599 = n33598 ^ n4700 ^ 1'b0 ;
  assign n33600 = n3389 & n33599 ;
  assign n33601 = ~n809 & n33600 ;
  assign n33602 = n3449 & n33601 ;
  assign n33603 = n850 & n5330 ;
  assign n33604 = n17194 & ~n33603 ;
  assign n33605 = ~n2020 & n15012 ;
  assign n33606 = n17533 ^ n2624 ^ 1'b0 ;
  assign n33607 = n28127 & ~n33606 ;
  assign n33608 = n33607 ^ n10627 ^ n7299 ;
  assign n33610 = n7596 | n12320 ;
  assign n33609 = n9898 & ~n17755 ;
  assign n33611 = n33610 ^ n33609 ^ 1'b0 ;
  assign n33612 = n25143 ^ n3120 ^ 1'b0 ;
  assign n33613 = n8107 | n16385 ;
  assign n33614 = n8979 & ~n33613 ;
  assign n33615 = n21233 ^ n1922 ^ 1'b0 ;
  assign n33616 = n10508 & n33615 ;
  assign n33617 = n33614 & n33616 ;
  assign n33618 = n26464 ^ n5635 ^ 1'b0 ;
  assign n33619 = n33617 | n33618 ;
  assign n33620 = n20457 & n22122 ;
  assign n33621 = n10203 | n30677 ;
  assign n33622 = n4043 | n33621 ;
  assign n33623 = n5752 & ~n33622 ;
  assign n33624 = n3672 ^ n3442 ^ 1'b0 ;
  assign n33625 = n5629 & n33624 ;
  assign n33626 = n33625 ^ n3969 ^ 1'b0 ;
  assign n33627 = n15035 & n33626 ;
  assign n33628 = ~n3267 & n4334 ;
  assign n33629 = n2038 & ~n33628 ;
  assign n33630 = ~n22961 & n33629 ;
  assign n33631 = n3380 | n33630 ;
  assign n33632 = n5468 & ~n29313 ;
  assign n33633 = n33632 ^ n33342 ^ 1'b0 ;
  assign n33634 = ~n703 & n18980 ;
  assign n33635 = n1782 | n1866 ;
  assign n33636 = n26707 ^ n20104 ^ n643 ;
  assign n33637 = n33635 | n33636 ;
  assign n33638 = n427 & ~n770 ;
  assign n33639 = n33638 ^ n11359 ^ n3100 ;
  assign n33640 = n19962 ^ n12293 ^ 1'b0 ;
  assign n33641 = n33640 ^ n3360 ^ 1'b0 ;
  assign n33642 = n13810 | n33641 ;
  assign n33643 = n27757 ^ n1110 ^ 1'b0 ;
  assign n33644 = n5040 & ~n33643 ;
  assign n33647 = n19971 ^ n11471 ^ 1'b0 ;
  assign n33645 = n4920 ^ n1961 ^ 1'b0 ;
  assign n33646 = ~n813 & n33645 ;
  assign n33648 = n33647 ^ n33646 ^ 1'b0 ;
  assign n33649 = ~n2269 & n3680 ;
  assign n33650 = ~n4024 & n33649 ;
  assign n33651 = n14657 & n26948 ;
  assign n33652 = n11483 ^ n9524 ^ 1'b0 ;
  assign n33653 = n1469 | n2495 ;
  assign n33654 = n8768 & n31433 ;
  assign n33655 = n4508 & n5449 ;
  assign n33656 = n33655 ^ n17946 ^ 1'b0 ;
  assign n33657 = n33656 ^ n23461 ^ 1'b0 ;
  assign n33658 = ~n33654 & n33657 ;
  assign n33659 = n19838 ^ n12513 ^ 1'b0 ;
  assign n33660 = n3209 & ~n33659 ;
  assign n33661 = n83 & n17844 ;
  assign n33662 = ~n3318 & n33661 ;
  assign n33663 = ~n7503 & n19674 ;
  assign n33664 = n17916 & n33663 ;
  assign n33665 = ~n1164 & n19149 ;
  assign n33666 = n33664 & n33665 ;
  assign n33667 = n1070 | n17596 ;
  assign n33668 = n2141 | n33667 ;
  assign n33669 = ( n1212 & ~n10259 ) | ( n1212 & n10844 ) | ( ~n10259 & n10844 ) ;
  assign n33670 = n6825 | n33669 ;
  assign n33671 = n14614 | n33670 ;
  assign n33672 = n520 & n33671 ;
  assign n33673 = n9806 & n33672 ;
  assign n33674 = n33673 ^ n24313 ^ 1'b0 ;
  assign n33675 = n2222 & ~n14973 ;
  assign n33676 = n33675 ^ n13573 ^ 1'b0 ;
  assign n33677 = n13561 | n25012 ;
  assign n33678 = n102 & ~n17929 ;
  assign n33679 = n19803 & n33678 ;
  assign n33680 = ~n26491 & n33679 ;
  assign n33681 = n9401 & ~n19544 ;
  assign n33682 = n8008 & n33681 ;
  assign n33685 = n8370 ^ n328 ^ 1'b0 ;
  assign n33686 = n20608 ^ n20540 ^ 1'b0 ;
  assign n33687 = n33685 | n33686 ;
  assign n33688 = n12303 | n33687 ;
  assign n33689 = n33688 ^ n14833 ^ 1'b0 ;
  assign n33683 = ~n357 & n5428 ;
  assign n33684 = n2196 | n33683 ;
  assign n33690 = n33689 ^ n33684 ^ 1'b0 ;
  assign n33692 = n25114 ^ n21275 ^ 1'b0 ;
  assign n33693 = n3074 & ~n33692 ;
  assign n33694 = n27900 & n33693 ;
  assign n33695 = n33694 ^ n16292 ^ 1'b0 ;
  assign n33691 = n2595 & ~n19854 ;
  assign n33696 = n33695 ^ n33691 ^ 1'b0 ;
  assign n33697 = ~n33690 & n33696 ;
  assign n33698 = n12768 | n17583 ;
  assign n33699 = n1134 & ~n3458 ;
  assign n33700 = n33699 ^ n9108 ^ 1'b0 ;
  assign n33701 = n13073 | n33700 ;
  assign n33702 = n1010 | n33701 ;
  assign n33703 = n13815 | n14462 ;
  assign n33704 = ( ~n6249 & n19085 ) | ( ~n6249 & n21227 ) | ( n19085 & n21227 ) ;
  assign n33705 = n33704 ^ n2380 ^ 1'b0 ;
  assign n33706 = n27681 | n33705 ;
  assign n33707 = n4448 | n5284 ;
  assign n33708 = ~n6281 & n24216 ;
  assign n33709 = ~n33707 & n33708 ;
  assign n33710 = ~n2382 & n22559 ;
  assign n33711 = n33710 ^ n26340 ^ 1'b0 ;
  assign n33712 = n15876 ^ n14429 ^ 1'b0 ;
  assign n33713 = n33712 ^ n21356 ^ 1'b0 ;
  assign n33714 = n1315 | n19575 ;
  assign n33715 = n5034 & n11278 ;
  assign n33716 = n9120 & n33715 ;
  assign n33717 = n33716 ^ n3368 ^ 1'b0 ;
  assign n33718 = n33714 | n33717 ;
  assign n33719 = n8730 ^ n5294 ^ 1'b0 ;
  assign n33720 = n33719 ^ n16079 ^ n4652 ;
  assign n33721 = n15861 & n31855 ;
  assign n33722 = ~n33720 & n33721 ;
  assign n33723 = n7277 ^ n4458 ^ 1'b0 ;
  assign n33724 = n26102 ^ n4626 ^ 1'b0 ;
  assign n33725 = n23233 ^ n20497 ^ 1'b0 ;
  assign n33726 = n29568 ^ n469 ^ 1'b0 ;
  assign n33727 = ~n21124 & n33726 ;
  assign n33728 = n33727 ^ n24623 ^ n16858 ;
  assign n33729 = ~n2321 & n33728 ;
  assign n33730 = ~n7179 & n13621 ;
  assign n33731 = n33730 ^ n330 ^ 1'b0 ;
  assign n33732 = n10521 ^ n8998 ^ n2092 ;
  assign n33733 = n4210 ^ n1239 ^ 1'b0 ;
  assign n33734 = n10285 & ~n33733 ;
  assign n33735 = ~n527 & n33734 ;
  assign n33736 = n33735 ^ n25788 ^ 1'b0 ;
  assign n33737 = ~n354 & n9563 ;
  assign n33738 = n33737 ^ n5292 ^ 1'b0 ;
  assign n33739 = n25422 ^ n1254 ^ 1'b0 ;
  assign n33741 = ~n5972 & n29239 ;
  assign n33740 = ~n4747 & n8842 ;
  assign n33742 = n33741 ^ n33740 ^ 1'b0 ;
  assign n33743 = n489 & n27308 ;
  assign n33744 = ~n5140 & n33743 ;
  assign n33745 = n33744 ^ n13976 ^ 1'b0 ;
  assign n33746 = n1394 | n2154 ;
  assign n33747 = n29217 | n33746 ;
  assign n33748 = n26604 ^ n15154 ^ 1'b0 ;
  assign n33749 = n15007 & n19896 ;
  assign n33750 = n33749 ^ n9412 ^ 1'b0 ;
  assign n33751 = n290 ^ n47 ^ 1'b0 ;
  assign n33752 = n20052 ^ n15208 ^ 1'b0 ;
  assign n33753 = n9697 & ~n33752 ;
  assign n33757 = n325 & ~n8236 ;
  assign n33758 = n509 & ~n33757 ;
  assign n33754 = n2463 | n8008 ;
  assign n33755 = n33754 ^ n5084 ^ 1'b0 ;
  assign n33756 = n137 & n33755 ;
  assign n33759 = n33758 ^ n33756 ^ 1'b0 ;
  assign n33760 = n5021 | n7936 ;
  assign n33768 = n23 | n37 ;
  assign n33769 = n23 & ~n33768 ;
  assign n33770 = n382 | n33769 ;
  assign n33771 = n33769 & ~n33770 ;
  assign n33772 = n1722 | n33771 ;
  assign n33761 = n8977 & ~n19426 ;
  assign n33762 = ~n8977 & n33761 ;
  assign n33763 = n33762 ^ n16413 ^ 1'b0 ;
  assign n33764 = n4947 | n12563 ;
  assign n33765 = n7840 & n33764 ;
  assign n33766 = ~n33763 & n33765 ;
  assign n33767 = n24775 | n33766 ;
  assign n33773 = n33772 ^ n33767 ^ 1'b0 ;
  assign n33774 = n7030 ^ n5245 ^ 1'b0 ;
  assign n33775 = n869 & n3789 ;
  assign n33776 = ~n13128 & n33775 ;
  assign n33777 = n33776 ^ n27876 ^ 1'b0 ;
  assign n33778 = n33774 | n33777 ;
  assign n33779 = n3321 | n4927 ;
  assign n33780 = n33445 ^ n13951 ^ 1'b0 ;
  assign n33781 = ~n439 & n15093 ;
  assign n33782 = n26283 ^ n16653 ^ 1'b0 ;
  assign n33783 = n31166 & ~n33782 ;
  assign n33784 = n14048 ^ n2032 ^ 1'b0 ;
  assign n33785 = ( n351 & n2154 ) | ( n351 & ~n19198 ) | ( n2154 & ~n19198 ) ;
  assign n33786 = n5284 & n33785 ;
  assign n33788 = n6530 ^ n1676 ^ 1'b0 ;
  assign n33787 = n2059 & n9385 ;
  assign n33789 = n33788 ^ n33787 ^ 1'b0 ;
  assign n33790 = n8330 & n20715 ;
  assign n33791 = n33790 ^ n24512 ^ 1'b0 ;
  assign n33792 = n32598 ^ n1829 ^ 1'b0 ;
  assign n33793 = ~n33791 & n33792 ;
  assign n33794 = n8790 & n24587 ;
  assign n33795 = n1337 | n5187 ;
  assign n33796 = n5187 & ~n33795 ;
  assign n33797 = n12642 | n33796 ;
  assign n33798 = n2879 & ~n17697 ;
  assign n33799 = n33798 ^ n3916 ^ 1'b0 ;
  assign n33800 = n14 | n14936 ;
  assign n33801 = n33799 & ~n33800 ;
  assign n33802 = n13682 & ~n33801 ;
  assign n33803 = n18229 ^ n1829 ^ 1'b0 ;
  assign n33805 = ~n1154 & n1927 ;
  assign n33806 = ~n2110 & n33805 ;
  assign n33804 = n1372 & n14391 ;
  assign n33807 = n33806 ^ n33804 ^ 1'b0 ;
  assign n33808 = n2144 & ~n5265 ;
  assign n33809 = n33808 ^ n5303 ^ 1'b0 ;
  assign n33810 = n11235 ^ n7355 ^ 1'b0 ;
  assign n33811 = n20752 ^ n13791 ^ 1'b0 ;
  assign n33812 = n9633 ^ n1445 ^ 1'b0 ;
  assign n33813 = ~n2762 & n11679 ;
  assign n33814 = n23568 & ~n33813 ;
  assign n33815 = n33814 ^ n10405 ^ 1'b0 ;
  assign n33816 = n5347 & n33815 ;
  assign n33817 = n11421 ^ n364 ^ 1'b0 ;
  assign n33818 = n17891 | n33817 ;
  assign n33819 = ~n6658 & n12978 ;
  assign n33820 = n10072 & n33819 ;
  assign n33821 = n22715 ^ n7608 ^ 1'b0 ;
  assign n33822 = n16909 & n23347 ;
  assign n33824 = n11651 ^ n2936 ^ 1'b0 ;
  assign n33825 = ~n3965 & n33824 ;
  assign n33826 = ~n1673 & n33825 ;
  assign n33827 = n33826 ^ n11096 ^ 1'b0 ;
  assign n33828 = ~n325 & n33827 ;
  assign n33829 = ~n1794 & n33828 ;
  assign n33823 = n14540 ^ n1511 ^ 1'b0 ;
  assign n33830 = n33829 ^ n33823 ^ 1'b0 ;
  assign n33832 = ~n2431 & n13350 ;
  assign n33831 = ~n9104 & n29596 ;
  assign n33833 = n33832 ^ n33831 ^ 1'b0 ;
  assign n33834 = n12000 & ~n33833 ;
  assign n33835 = n4411 & n25670 ;
  assign n33836 = n33835 ^ n23098 ^ n22993 ;
  assign n33837 = n33836 ^ n25449 ^ n16576 ;
  assign n33838 = n1472 | n3085 ;
  assign n33839 = n33838 ^ n671 ^ 1'b0 ;
  assign n33840 = n26329 ^ n16156 ^ 1'b0 ;
  assign n33841 = n30131 ^ n20255 ^ 1'b0 ;
  assign n33845 = n11334 ^ n2414 ^ 1'b0 ;
  assign n33842 = n1439 & ~n1822 ;
  assign n33843 = ~n1763 & n33842 ;
  assign n33844 = n33843 ^ n18047 ^ 1'b0 ;
  assign n33846 = n33845 ^ n33844 ^ 1'b0 ;
  assign n33847 = n536 | n33846 ;
  assign n33848 = n26775 ^ n15055 ^ 1'b0 ;
  assign n33849 = n20272 & n26408 ;
  assign n33850 = ~n3112 & n27252 ;
  assign n33851 = n23894 & ~n33850 ;
  assign n33852 = n15933 ^ n4823 ^ 1'b0 ;
  assign n33853 = n33851 & n33852 ;
  assign n33854 = n4465 & ~n16441 ;
  assign n33855 = n4090 & ~n11412 ;
  assign n33856 = n4236 | n33855 ;
  assign n33857 = n3773 ^ n663 ^ 1'b0 ;
  assign n33858 = n3804 & n11961 ;
  assign n33859 = ~n33857 & n33858 ;
  assign n33860 = n159 & n3042 ;
  assign n33861 = n33629 ^ n1134 ^ 1'b0 ;
  assign n33862 = n5096 ^ n4906 ^ n4550 ;
  assign n33863 = n21525 | n33862 ;
  assign n33864 = n31079 ^ n18654 ^ 1'b0 ;
  assign n33865 = ~n6102 & n33864 ;
  assign n33866 = ~n4008 & n8721 ;
  assign n33867 = n33866 ^ n995 ^ 1'b0 ;
  assign n33868 = n33867 ^ n10362 ^ 1'b0 ;
  assign n33869 = n26756 ^ n11407 ^ n748 ;
  assign n33870 = ~n144 & n33869 ;
  assign n33871 = n495 & n802 ;
  assign n33872 = n5928 ^ n5920 ^ 1'b0 ;
  assign n33873 = n24608 ^ n553 ^ 1'b0 ;
  assign n33874 = ~n33256 & n33873 ;
  assign n33875 = n33874 ^ n5423 ^ 1'b0 ;
  assign n33876 = n6889 & ~n23030 ;
  assign n33877 = n4256 & ~n24713 ;
  assign n33878 = n29823 ^ n82 ^ 1'b0 ;
  assign n33879 = ~n4098 & n19188 ;
  assign n33880 = n164 & n33879 ;
  assign n33881 = n33880 ^ n6605 ^ 1'b0 ;
  assign n33882 = ~n1889 & n33881 ;
  assign n33884 = n1401 & ~n18016 ;
  assign n33885 = n33884 ^ n12890 ^ 1'b0 ;
  assign n33883 = n15742 | n25112 ;
  assign n33886 = n33885 ^ n33883 ^ 1'b0 ;
  assign n33887 = n29640 ^ n20474 ^ 1'b0 ;
  assign n33888 = ~n4954 & n18294 ;
  assign n33889 = n33887 & n33888 ;
  assign n33890 = ~n13808 & n26182 ;
  assign n33891 = n33890 ^ n32545 ^ 1'b0 ;
  assign n33892 = n33891 ^ n13519 ^ 1'b0 ;
  assign n33893 = ~n1650 & n3512 ;
  assign n33894 = n17800 | n20141 ;
  assign n33895 = n21722 & ~n33894 ;
  assign n33896 = n25060 ^ n5465 ^ n47 ;
  assign n33898 = n2907 & n23311 ;
  assign n33897 = n5844 & ~n7596 ;
  assign n33899 = n33898 ^ n33897 ^ n15326 ;
  assign n33900 = n33899 ^ n24544 ^ 1'b0 ;
  assign n33901 = ~n12157 & n20224 ;
  assign n33902 = n33900 & n33901 ;
  assign n33903 = n26246 ^ n10762 ^ n9800 ;
  assign n33904 = n16554 | n23753 ;
  assign n33905 = n4239 & n5790 ;
  assign n33906 = ~n1309 & n12561 ;
  assign n33907 = n3317 & n31544 ;
  assign n33908 = ~n31544 & n33907 ;
  assign n33909 = n10845 & ~n33908 ;
  assign n33912 = ( n2074 & n2891 ) | ( n2074 & n15244 ) | ( n2891 & n15244 ) ;
  assign n33910 = n10343 ^ n3859 ^ 1'b0 ;
  assign n33911 = n10438 & n33910 ;
  assign n33913 = n33912 ^ n33911 ^ 1'b0 ;
  assign n33914 = n364 | n2661 ;
  assign n33915 = n33914 ^ n27899 ^ 1'b0 ;
  assign n33916 = n11389 ^ n7406 ^ 1'b0 ;
  assign n33917 = ~n33915 & n33916 ;
  assign n33918 = ~n4726 & n13556 ;
  assign n33919 = n9750 ^ n327 ^ 1'b0 ;
  assign n33920 = n13934 & ~n33919 ;
  assign n33921 = ~n19891 & n33920 ;
  assign n33922 = n2175 ^ n1345 ^ 1'b0 ;
  assign n33923 = n2128 & ~n33922 ;
  assign n33924 = n3676 & n33923 ;
  assign n33925 = n33924 ^ n18308 ^ 1'b0 ;
  assign n33926 = n6994 & n33925 ;
  assign n33927 = n19870 | n25037 ;
  assign n33928 = n942 & n8370 ;
  assign n33929 = n33928 ^ n27162 ^ 1'b0 ;
  assign n33930 = ~n4785 & n33929 ;
  assign n33931 = n21942 & ~n33930 ;
  assign n33932 = n33931 ^ n24353 ^ 1'b0 ;
  assign n33933 = n32781 ^ n12157 ^ n1298 ;
  assign n33934 = n2523 & ~n4660 ;
  assign n33935 = ~n3483 & n12978 ;
  assign n33936 = n17785 & n33935 ;
  assign n33938 = n20314 ^ n7384 ^ 1'b0 ;
  assign n33937 = n8486 & ~n27001 ;
  assign n33939 = n33938 ^ n33937 ^ 1'b0 ;
  assign n33940 = ~n1740 & n33939 ;
  assign n33941 = n33940 ^ n6986 ^ 1'b0 ;
  assign n33942 = n29119 ^ n2933 ^ 1'b0 ;
  assign n33943 = n23217 ^ n6764 ^ 1'b0 ;
  assign n33944 = ~n25579 & n33943 ;
  assign n33945 = n10762 & ~n23140 ;
  assign n33946 = n11330 & ~n12518 ;
  assign n33947 = n7650 & ~n33946 ;
  assign n33948 = ~n4088 & n33947 ;
  assign n33949 = n26977 | n33948 ;
  assign n33950 = n16140 ^ n296 ^ 1'b0 ;
  assign n33951 = ~n9968 & n33950 ;
  assign n33952 = n5125 & n33951 ;
  assign n33953 = ~n29800 & n33952 ;
  assign n33954 = ~n8380 & n33347 ;
  assign n33955 = n2460 | n20365 ;
  assign n33956 = n33955 ^ n9903 ^ 1'b0 ;
  assign n33957 = ~n7404 & n18715 ;
  assign n33958 = n30687 ^ n24197 ^ 1'b0 ;
  assign n33959 = n2490 | n33958 ;
  assign n33960 = n684 & ~n33959 ;
  assign n33961 = ~n19211 & n33960 ;
  assign n33962 = n25223 & ~n33961 ;
  assign n33963 = n6349 & ~n8793 ;
  assign n33964 = n20189 & n33963 ;
  assign n33965 = ~n497 & n9461 ;
  assign n33966 = n4095 | n12087 ;
  assign n33967 = n33965 & ~n33966 ;
  assign n33968 = ~n11275 & n15814 ;
  assign n33969 = n9954 & ~n12495 ;
  assign n33970 = n33969 ^ n452 ^ 1'b0 ;
  assign n33971 = n33968 | n33970 ;
  assign n33972 = ~n8692 & n9668 ;
  assign n33973 = ~n582 & n6444 ;
  assign n33974 = n33973 ^ n13164 ^ n6054 ;
  assign n33975 = n33972 & ~n33974 ;
  assign n33976 = n33975 ^ n5972 ^ 1'b0 ;
  assign n33977 = n10548 ^ n2619 ^ 1'b0 ;
  assign n33978 = ~n9817 & n26420 ;
  assign n33979 = n16954 ^ n3921 ^ 1'b0 ;
  assign n33980 = n26218 ^ n10917 ^ 1'b0 ;
  assign n33981 = ~n14483 & n25184 ;
  assign n33982 = n8518 & n30625 ;
  assign n33983 = n33982 ^ n1486 ^ 1'b0 ;
  assign n33984 = n11226 | n21131 ;
  assign n33985 = ( n16904 & n20812 ) | ( n16904 & ~n33984 ) | ( n20812 & ~n33984 ) ;
  assign n33986 = ( n7269 & n18176 ) | ( n7269 & ~n28246 ) | ( n18176 & ~n28246 ) ;
  assign n33987 = n17989 & ~n33986 ;
  assign n33988 = n8886 & n33987 ;
  assign n33989 = n3885 & ~n24649 ;
  assign n33990 = n16117 | n33989 ;
  assign n33991 = n33988 & ~n33990 ;
  assign n33992 = ~n348 & n18778 ;
  assign n33993 = n33992 ^ n13833 ^ 1'b0 ;
  assign n33994 = n16492 & n29077 ;
  assign n33995 = ~n1686 & n33994 ;
  assign n33996 = n532 | n6481 ;
  assign n33997 = n33996 ^ n7612 ^ 1'b0 ;
  assign n33998 = ~n9143 & n29226 ;
  assign n33999 = n1931 & ~n11024 ;
  assign n34000 = ~n33998 & n33999 ;
  assign n34001 = n34000 ^ n14331 ^ 1'b0 ;
  assign n34002 = n8161 & n34001 ;
  assign n34003 = n14544 ^ n81 ^ 1'b0 ;
  assign n34006 = n339 | n8894 ;
  assign n34004 = n12119 | n18148 ;
  assign n34005 = n15 & ~n34004 ;
  assign n34007 = n34006 ^ n34005 ^ n7074 ;
  assign n34008 = n29072 | n34007 ;
  assign n34009 = n34008 ^ n9233 ^ 1'b0 ;
  assign n34010 = n1203 & n5749 ;
  assign n34011 = ~n17178 & n34010 ;
  assign n34012 = n3444 | n8046 ;
  assign n34013 = n34011 & ~n34012 ;
  assign n34014 = ( n940 & ~n3121 ) | ( n940 & n11483 ) | ( ~n3121 & n11483 ) ;
  assign n34015 = n461 | n34014 ;
  assign n34016 = n3208 & ~n34015 ;
  assign n34017 = n4629 ^ n196 ^ 1'b0 ;
  assign n34018 = ~n6751 & n12008 ;
  assign n34019 = ~n12339 & n34018 ;
  assign n34020 = n34019 ^ n24936 ^ 1'b0 ;
  assign n34021 = ~n376 & n11822 ;
  assign n34022 = n16011 & n34021 ;
  assign n34023 = n17560 & ~n32700 ;
  assign n34024 = ~n23805 & n24026 ;
  assign n34025 = ~n34023 & n34024 ;
  assign n34026 = n34025 ^ n16395 ^ 1'b0 ;
  assign n34027 = n6949 | n27444 ;
  assign n34028 = n34027 ^ n18735 ^ 1'b0 ;
  assign n34029 = ~n8954 & n34028 ;
  assign n34030 = n9934 & n14306 ;
  assign n34031 = n14071 | n34030 ;
  assign n34032 = n5575 | n34031 ;
  assign n34033 = n805 & ~n20510 ;
  assign n34034 = ~n7264 & n16029 ;
  assign n34035 = n34034 ^ n18538 ^ 1'b0 ;
  assign n34036 = n7904 & n9051 ;
  assign n34037 = n4409 ^ n995 ^ 1'b0 ;
  assign n34038 = n11312 ^ n10767 ^ 1'b0 ;
  assign n34039 = n34038 ^ n30653 ^ 1'b0 ;
  assign n34040 = n34037 & n34039 ;
  assign n34041 = n19359 ^ n5293 ^ 1'b0 ;
  assign n34042 = n10586 | n34041 ;
  assign n34043 = n2286 & ~n8751 ;
  assign n34044 = n8246 | n8656 ;
  assign n34045 = n34043 | n34044 ;
  assign n34046 = n34045 ^ n10201 ^ 1'b0 ;
  assign n34047 = n20951 ^ n14039 ^ 1'b0 ;
  assign n34048 = n18058 ^ n13488 ^ 1'b0 ;
  assign n34049 = n338 & n16104 ;
  assign n34050 = n34049 ^ n34007 ^ 1'b0 ;
  assign n34051 = n10544 ^ n4586 ^ 1'b0 ;
  assign n34052 = n6578 | n34051 ;
  assign n34053 = n34052 ^ n26341 ^ n5012 ;
  assign n34054 = n10736 ^ n951 ^ 1'b0 ;
  assign n34055 = n2107 | n34054 ;
  assign n34056 = ~n1015 & n34055 ;
  assign n34057 = n11735 | n31778 ;
  assign n34058 = ~n627 & n4650 ;
  assign n34059 = n14211 & n17796 ;
  assign n34060 = n8189 & ~n18970 ;
  assign n34061 = n8227 ^ n675 ^ n139 ;
  assign n34062 = n6855 & n31198 ;
  assign n34063 = ~n5971 & n34062 ;
  assign n34064 = ~n7098 & n25662 ;
  assign n34065 = n34064 ^ n1637 ^ 1'b0 ;
  assign n34069 = ~n3219 & n14410 ;
  assign n34070 = ~n2912 & n34069 ;
  assign n34066 = n17364 ^ n11525 ^ 1'b0 ;
  assign n34067 = ~n703 & n34066 ;
  assign n34068 = ~n29515 & n34067 ;
  assign n34071 = n34070 ^ n34068 ^ 1'b0 ;
  assign n34072 = ~n4258 & n5918 ;
  assign n34073 = n200 | n19896 ;
  assign n34074 = n5731 | n28537 ;
  assign n34075 = n1785 | n34074 ;
  assign n34076 = n695 & n7606 ;
  assign n34077 = n34076 ^ n504 ^ 1'b0 ;
  assign n34078 = n22422 ^ n5014 ^ 1'b0 ;
  assign n34079 = n2269 & ~n24036 ;
  assign n34080 = ~n20848 & n34079 ;
  assign n34081 = n20059 & n34080 ;
  assign n34082 = ~n3577 & n34081 ;
  assign n34083 = n34082 ^ n5575 ^ 1'b0 ;
  assign n34084 = n1683 ^ n545 ^ 1'b0 ;
  assign n34085 = ( n2512 & ~n6911 ) | ( n2512 & n12431 ) | ( ~n6911 & n12431 ) ;
  assign n34086 = ~n30837 & n34085 ;
  assign n34090 = n7260 & n8987 ;
  assign n34091 = n34090 ^ n8274 ^ 1'b0 ;
  assign n34087 = n2627 & n7767 ;
  assign n34088 = n22907 & ~n25196 ;
  assign n34089 = n34087 & n34088 ;
  assign n34092 = n34091 ^ n34089 ^ 1'b0 ;
  assign n34093 = n3702 & ~n4422 ;
  assign n34094 = n34093 ^ n1598 ^ 1'b0 ;
  assign n34095 = ~n11046 & n34094 ;
  assign n34096 = n16239 ^ n14474 ^ 1'b0 ;
  assign n34098 = ~n539 & n2438 ;
  assign n34099 = n34098 ^ n29103 ^ 1'b0 ;
  assign n34100 = n139 | n5471 ;
  assign n34101 = n34100 ^ n9390 ^ 1'b0 ;
  assign n34102 = n34099 & ~n34101 ;
  assign n34097 = n5502 | n6533 ;
  assign n34103 = n34102 ^ n34097 ^ 1'b0 ;
  assign n34104 = n2092 & n12201 ;
  assign n34105 = n34104 ^ n2515 ^ 1'b0 ;
  assign n34106 = n1117 & ~n13063 ;
  assign n34107 = ~n8389 & n34106 ;
  assign n34108 = n15711 ^ n7340 ^ 1'b0 ;
  assign n34109 = n10937 ^ n4473 ^ n1117 ;
  assign n34110 = ~n4120 & n34109 ;
  assign n34111 = n34110 ^ n4416 ^ 1'b0 ;
  assign n34112 = n34108 | n34111 ;
  assign n34113 = n34112 ^ n19375 ^ 1'b0 ;
  assign n34114 = n11299 & ~n34113 ;
  assign n34115 = n6477 ^ n462 ^ 1'b0 ;
  assign n34116 = n24125 & n34115 ;
  assign n34117 = ~n8290 & n22273 ;
  assign n34118 = n34117 ^ n24761 ^ 1'b0 ;
  assign n34119 = n7006 | n7376 ;
  assign n34120 = n851 & n34119 ;
  assign n34125 = n11027 & n15454 ;
  assign n34126 = n34125 ^ n22528 ^ 1'b0 ;
  assign n34121 = n5513 | n25868 ;
  assign n34122 = n34121 ^ n20590 ^ 1'b0 ;
  assign n34123 = ~n169 & n34122 ;
  assign n34124 = n14667 & ~n34123 ;
  assign n34127 = n34126 ^ n34124 ^ 1'b0 ;
  assign n34128 = ~n5979 & n17163 ;
  assign n34129 = n34128 ^ n7066 ^ 1'b0 ;
  assign n34130 = n1814 ^ n621 ^ 1'b0 ;
  assign n34131 = n3472 | n34130 ;
  assign n34132 = n34131 ^ n4629 ^ 1'b0 ;
  assign n34133 = n7221 | n13854 ;
  assign n34134 = n34133 ^ n26090 ^ 1'b0 ;
  assign n34135 = n7115 & ~n24859 ;
  assign n34136 = n18076 ^ n5477 ^ 1'b0 ;
  assign n34137 = n13656 ^ n11265 ^ 1'b0 ;
  assign n34138 = ~n34136 & n34137 ;
  assign n34139 = ~n2209 & n34138 ;
  assign n34140 = n4689 | n22198 ;
  assign n34141 = n34140 ^ n14955 ^ 1'b0 ;
  assign n34142 = n13877 & ~n19452 ;
  assign n34143 = n31698 ^ n8539 ^ 1'b0 ;
  assign n34144 = n33716 ^ n6230 ^ 1'b0 ;
  assign n34145 = n4793 & ~n6509 ;
  assign n34146 = n10229 & n34145 ;
  assign n34147 = n34146 ^ n7646 ^ 1'b0 ;
  assign n34148 = n29096 & n34147 ;
  assign n34149 = n3311 & ~n34148 ;
  assign n34150 = n22709 ^ n764 ^ 1'b0 ;
  assign n34151 = ~n7231 & n34150 ;
  assign n34152 = n3077 & n5370 ;
  assign n34153 = ~n419 & n34152 ;
  assign n34154 = n1571 ^ n942 ^ 1'b0 ;
  assign n34155 = n1768 | n8186 ;
  assign n34156 = n9767 | n34155 ;
  assign n34157 = n18422 ^ n11533 ^ 1'b0 ;
  assign n34158 = n7420 & ~n34157 ;
  assign n34159 = n19 & n34158 ;
  assign n34160 = n34159 ^ n9887 ^ 1'b0 ;
  assign n34161 = n9425 | n27466 ;
  assign n34162 = n12534 ^ n7574 ^ 1'b0 ;
  assign n34163 = n5793 ^ n4559 ^ n1194 ;
  assign n34164 = ~n754 & n14675 ;
  assign n34165 = n5345 ^ n4474 ^ 1'b0 ;
  assign n34166 = ~n9860 & n34165 ;
  assign n34167 = n34166 ^ n19712 ^ n11488 ;
  assign n34168 = n6822 & ~n29167 ;
  assign n34169 = n34168 ^ n33210 ^ 1'b0 ;
  assign n34170 = ~n8915 & n34169 ;
  assign n34171 = ~n504 & n34170 ;
  assign n34172 = n1248 & n5788 ;
  assign n34173 = n34172 ^ n8863 ^ 1'b0 ;
  assign n34174 = ( n30928 & n31049 ) | ( n30928 & ~n34173 ) | ( n31049 & ~n34173 ) ;
  assign n34175 = n22099 ^ n16775 ^ 1'b0 ;
  assign n34176 = n25553 ^ n2083 ^ 1'b0 ;
  assign n34177 = ~n371 & n34176 ;
  assign n34178 = ~n5388 & n16244 ;
  assign n34179 = n55 | n34178 ;
  assign n34180 = n6168 | n14437 ;
  assign n34181 = n34180 ^ n4201 ^ n578 ;
  assign n34182 = n4533 & n34181 ;
  assign n34183 = ~n4286 & n34182 ;
  assign n34184 = n1358 & n17569 ;
  assign n34185 = n34184 ^ n12115 ^ 1'b0 ;
  assign n34186 = ~n5033 & n17818 ;
  assign n34187 = n949 & n19632 ;
  assign n34188 = n1392 & n34187 ;
  assign n34189 = n13095 & ~n19064 ;
  assign n34190 = n22762 ^ n227 ^ 1'b0 ;
  assign n34191 = n34190 ^ n9925 ^ 1'b0 ;
  assign n34192 = n6043 | n15511 ;
  assign n34193 = ~n11275 & n34192 ;
  assign n34194 = n34193 ^ n16186 ^ 1'b0 ;
  assign n34195 = n34194 ^ n7948 ^ 1'b0 ;
  assign n34196 = n19760 & n27931 ;
  assign n34197 = n6089 ^ n4361 ^ 1'b0 ;
  assign n34198 = n6732 & ~n11355 ;
  assign n34199 = n4677 & ~n16928 ;
  assign n34200 = n34199 ^ n5056 ^ 1'b0 ;
  assign n34201 = n11439 ^ n7360 ^ 1'b0 ;
  assign n34202 = n947 | n2814 ;
  assign n34203 = n5364 | n12167 ;
  assign n34204 = n18434 & ~n26516 ;
  assign n34205 = n10202 ^ n9201 ^ 1'b0 ;
  assign n34206 = n15666 & n34205 ;
  assign n34207 = n12665 | n16534 ;
  assign n34211 = n5387 & ~n7340 ;
  assign n34208 = n265 & n354 ;
  assign n34209 = n2789 & n34208 ;
  assign n34210 = n17635 | n34209 ;
  assign n34212 = n34211 ^ n34210 ^ 1'b0 ;
  assign n34214 = n26598 ^ n2645 ^ 1'b0 ;
  assign n34215 = n31970 | n34214 ;
  assign n34213 = ~n3401 & n12663 ;
  assign n34216 = n34215 ^ n34213 ^ 1'b0 ;
  assign n34217 = n20556 ^ n7622 ^ 1'b0 ;
  assign n34218 = ~n10340 & n34217 ;
  assign n34219 = n13184 | n15316 ;
  assign n34220 = n5024 ^ n2842 ^ 1'b0 ;
  assign n34221 = ~n17013 & n34220 ;
  assign n34222 = n23237 ^ n596 ^ 1'b0 ;
  assign n34223 = n6929 ^ n2869 ^ 1'b0 ;
  assign n34224 = ~n10038 & n34223 ;
  assign n34225 = ~x0 & n34224 ;
  assign n34226 = n34225 ^ n3309 ^ 1'b0 ;
  assign n34227 = n13326 ^ n4710 ^ 1'b0 ;
  assign n34228 = n2790 | n34227 ;
  assign n34229 = n11087 & ~n34228 ;
  assign n34230 = n34229 ^ n2376 ^ 1'b0 ;
  assign n34231 = n15992 & ~n34230 ;
  assign n34232 = n21537 ^ n8072 ^ 1'b0 ;
  assign n34233 = ~n2594 & n34232 ;
  assign n34234 = n27355 & n34233 ;
  assign n34235 = n34234 ^ n11678 ^ 1'b0 ;
  assign n34236 = ~n1304 & n15438 ;
  assign n34237 = n24955 & n34236 ;
  assign n34238 = n34237 ^ n6351 ^ 1'b0 ;
  assign n34239 = n4479 & n34238 ;
  assign n34240 = n19479 ^ n19011 ^ 1'b0 ;
  assign n34241 = n21229 | n34240 ;
  assign n34242 = ~n7221 & n22472 ;
  assign n34243 = n21021 ^ n5059 ^ 1'b0 ;
  assign n34244 = ( ~n612 & n15810 ) | ( ~n612 & n31101 ) | ( n15810 & n31101 ) ;
  assign n34245 = n25876 ^ n15673 ^ 1'b0 ;
  assign n34246 = n9390 | n34245 ;
  assign n34247 = n25826 ^ n7328 ^ n940 ;
  assign n34248 = ~n4449 & n13576 ;
  assign n34249 = n29069 & n34248 ;
  assign n34253 = n7596 ^ n4869 ^ 1'b0 ;
  assign n34250 = n22840 ^ n7980 ^ 1'b0 ;
  assign n34251 = n11200 & n34250 ;
  assign n34252 = ~n16475 & n34251 ;
  assign n34254 = n34253 ^ n34252 ^ 1'b0 ;
  assign n34255 = ( ~n8397 & n9075 ) | ( ~n8397 & n13110 ) | ( n9075 & n13110 ) ;
  assign n34256 = n4439 | n15698 ;
  assign n34257 = n34256 ^ n7424 ^ 1'b0 ;
  assign n34260 = n17069 & ~n27746 ;
  assign n34261 = n34260 ^ n16677 ^ 1'b0 ;
  assign n34258 = n7110 ^ n4924 ^ 1'b0 ;
  assign n34259 = n25693 & n34258 ;
  assign n34262 = n34261 ^ n34259 ^ 1'b0 ;
  assign n34263 = n2955 | n6587 ;
  assign n34264 = n34263 ^ n24102 ^ 1'b0 ;
  assign n34265 = n34264 ^ n11061 ^ n5183 ;
  assign n34266 = n27165 | n34265 ;
  assign n34267 = n8757 & n11760 ;
  assign n34268 = n10996 ^ n5248 ^ 1'b0 ;
  assign n34269 = n34268 ^ n20844 ^ 1'b0 ;
  assign n34270 = n2142 & n4668 ;
  assign n34271 = n11291 & ~n21982 ;
  assign n34272 = n34271 ^ n24256 ^ 1'b0 ;
  assign n34273 = ~n18332 & n20240 ;
  assign n34274 = n16728 ^ n5418 ^ 1'b0 ;
  assign n34275 = n21436 ^ n6653 ^ 1'b0 ;
  assign n34276 = n16673 & ~n34275 ;
  assign n34277 = n27735 & n28968 ;
  assign n34278 = n25007 ^ x0 ^ 1'b0 ;
  assign n34279 = ( n5010 & n9666 ) | ( n5010 & n21752 ) | ( n9666 & n21752 ) ;
  assign n34280 = ~n557 & n34279 ;
  assign n34281 = n15543 ^ n1637 ^ 1'b0 ;
  assign n34282 = ~n5747 & n11934 ;
  assign n34283 = n5373 & ~n8358 ;
  assign n34284 = n34283 ^ n14516 ^ 1'b0 ;
  assign n34285 = n21868 | n34284 ;
  assign n34286 = n34285 ^ n3368 ^ 1'b0 ;
  assign n34287 = n1186 & n7767 ;
  assign n34288 = ~n30 & n34287 ;
  assign n34289 = n3701 & ~n9526 ;
  assign n34290 = n6519 & n34289 ;
  assign n34291 = ( n17974 & ~n34288 ) | ( n17974 & n34290 ) | ( ~n34288 & n34290 ) ;
  assign n34292 = n1135 | n4533 ;
  assign n34293 = n4759 | n34292 ;
  assign n34294 = n25634 & n26203 ;
  assign n34295 = n18534 ^ n11365 ^ 1'b0 ;
  assign n34296 = n2967 ^ n1802 ^ 1'b0 ;
  assign n34297 = ~n18735 & n34296 ;
  assign n34298 = n8138 | n34297 ;
  assign n34299 = ( n764 & ~n9805 ) | ( n764 & n16192 ) | ( ~n9805 & n16192 ) ;
  assign n34300 = n34299 ^ n26420 ^ 1'b0 ;
  assign n34301 = n6277 | n34300 ;
  assign n34302 = n3036 & n9404 ;
  assign n34303 = ~n10954 & n34302 ;
  assign n34304 = n34303 ^ n25900 ^ 1'b0 ;
  assign n34305 = n18440 & ~n34304 ;
  assign n34306 = ~n10574 & n17273 ;
  assign n34307 = n34306 ^ n18869 ^ 1'b0 ;
  assign n34308 = n17574 | n17737 ;
  assign n34309 = n2910 & n34308 ;
  assign n34310 = n34307 | n34309 ;
  assign n34311 = n12633 ^ n8865 ^ 1'b0 ;
  assign n34312 = n11722 & n13688 ;
  assign n34313 = n34312 ^ n292 ^ 1'b0 ;
  assign n34314 = n28243 & n34313 ;
  assign n34315 = ~n34311 & n34314 ;
  assign n34316 = n20118 ^ n5398 ^ 1'b0 ;
  assign n34317 = n16752 & n34316 ;
  assign n34318 = n33476 & ~n34317 ;
  assign n34319 = n5144 & n10294 ;
  assign n34320 = n34319 ^ n24232 ^ 1'b0 ;
  assign n34323 = n10937 ^ n1951 ^ 1'b0 ;
  assign n34321 = ~n726 & n6003 ;
  assign n34322 = ~n7737 & n34321 ;
  assign n34324 = n34323 ^ n34322 ^ 1'b0 ;
  assign n34325 = ~n2214 & n34324 ;
  assign n34327 = n43 & ~n2747 ;
  assign n34328 = ~n43 & n34327 ;
  assign n34329 = ~n1543 & n34328 ;
  assign n34330 = n34329 ^ n11390 ^ 1'b0 ;
  assign n34331 = n165 & ~n17849 ;
  assign n34332 = n17849 & n34331 ;
  assign n34333 = n34332 ^ n13110 ^ 1'b0 ;
  assign n34334 = n34330 & ~n34333 ;
  assign n34335 = n34334 ^ n1229 ^ 1'b0 ;
  assign n34326 = n5539 & n10794 ;
  assign n34336 = n34335 ^ n34326 ^ 1'b0 ;
  assign n34337 = n32935 | n34336 ;
  assign n34338 = n34325 & n34337 ;
  assign n34339 = n17752 ^ n6887 ^ 1'b0 ;
  assign n34340 = n24185 & n34339 ;
  assign n34341 = n34340 ^ n4133 ^ 1'b0 ;
  assign n34342 = n6377 | n11573 ;
  assign n34343 = n7039 ^ n3566 ^ 1'b0 ;
  assign n34344 = n24072 | n34343 ;
  assign n34345 = n34342 | n34344 ;
  assign n34346 = n6884 & ~n34345 ;
  assign n34347 = n34341 & n34346 ;
  assign n34348 = n29119 & ~n34347 ;
  assign n34349 = n15593 & n15667 ;
  assign n34350 = n24307 ^ n2817 ^ 1'b0 ;
  assign n34351 = n3663 | n34350 ;
  assign n34352 = n9114 ^ n618 ^ 1'b0 ;
  assign n34353 = ~n24938 & n26749 ;
  assign n34354 = ~n16746 & n23739 ;
  assign n34355 = n17349 & n34354 ;
  assign n34356 = n4381 | n6390 ;
  assign n34357 = n741 | n34356 ;
  assign n34358 = ~n5535 & n34357 ;
  assign n34359 = ~n22643 & n34358 ;
  assign n34360 = n26769 ^ n24158 ^ 1'b0 ;
  assign n34361 = ~n4893 & n34360 ;
  assign n34362 = n27080 ^ n16773 ^ 1'b0 ;
  assign n34363 = n1602 ^ n632 ^ 1'b0 ;
  assign n34364 = ~n18996 & n26129 ;
  assign n34365 = n34364 ^ n3447 ^ 1'b0 ;
  assign n34366 = n10091 & ~n14683 ;
  assign n34367 = ~n14353 & n18574 ;
  assign n34368 = n20406 & ~n28821 ;
  assign n34369 = n34368 ^ n18477 ^ 1'b0 ;
  assign n34370 = n6139 ^ n4684 ^ 1'b0 ;
  assign n34371 = ~n12228 & n34370 ;
  assign n34372 = n34371 ^ n24418 ^ 1'b0 ;
  assign n34373 = ( ~n14838 & n33862 ) | ( ~n14838 & n34372 ) | ( n33862 & n34372 ) ;
  assign n34374 = n31318 ^ n2916 ^ 1'b0 ;
  assign n34375 = n24473 ^ n5317 ^ 1'b0 ;
  assign n34376 = n33166 ^ n32082 ^ 1'b0 ;
  assign n34377 = n5400 | n34376 ;
  assign n34378 = n2269 & ~n5084 ;
  assign n34379 = n34378 ^ n297 ^ 1'b0 ;
  assign n34380 = n9302 & ~n34379 ;
  assign n34381 = n55 & n34380 ;
  assign n34382 = n8879 | n27002 ;
  assign n34383 = n2967 & ~n24380 ;
  assign n34384 = n6160 & ~n28908 ;
  assign n34385 = n34384 ^ n17730 ^ 1'b0 ;
  assign n34386 = n524 ^ n37 ^ 1'b0 ;
  assign n34387 = n24216 ^ n17914 ^ n17794 ;
  assign n34388 = ~n7056 & n34387 ;
  assign n34389 = ( n423 & n813 ) | ( n423 & n13193 ) | ( n813 & n13193 ) ;
  assign n34390 = ( n8763 & n12721 ) | ( n8763 & n34389 ) | ( n12721 & n34389 ) ;
  assign n34391 = n34390 ^ n16411 ^ 1'b0 ;
  assign n34392 = n26456 & ~n34391 ;
  assign n34393 = n11775 & ~n33640 ;
  assign n34394 = ~n34392 & n34393 ;
  assign n34395 = n8416 ^ n5084 ^ 1'b0 ;
  assign n34396 = n10571 ^ n8685 ^ n6944 ;
  assign n34397 = n7277 & n34396 ;
  assign n34398 = n11885 ^ n9228 ^ 1'b0 ;
  assign n34399 = n6627 | n34398 ;
  assign n34400 = ~n29777 & n34399 ;
  assign n34401 = n23814 ^ n11412 ^ 1'b0 ;
  assign n34402 = n907 | n34401 ;
  assign n34403 = n34400 & ~n34402 ;
  assign n34404 = n376 & ~n1659 ;
  assign n34405 = n11611 & n34404 ;
  assign n34406 = n9170 | n10219 ;
  assign n34407 = ~n8792 & n34406 ;
  assign n34408 = ~n4000 & n34407 ;
  assign n34409 = n18942 & ~n34408 ;
  assign n34410 = ~n22472 & n34409 ;
  assign n34411 = ~n8215 & n10327 ;
  assign n34412 = n26523 & n34411 ;
  assign n34413 = n34412 ^ n5280 ^ 1'b0 ;
  assign n34414 = ~n2733 & n3827 ;
  assign n34415 = ~n86 & n34414 ;
  assign n34416 = n23493 ^ n3828 ^ 1'b0 ;
  assign n34417 = n34415 | n34416 ;
  assign n34418 = n709 & ~n7718 ;
  assign n34419 = ~n1394 & n2784 ;
  assign n34420 = n28116 & n34419 ;
  assign n34421 = n5890 & n31301 ;
  assign n34422 = ~n2805 & n34421 ;
  assign n34423 = n32545 ^ n22502 ^ 1'b0 ;
  assign n34424 = n2882 & n10495 ;
  assign n34425 = n34424 ^ n13831 ^ 1'b0 ;
  assign n34426 = n34425 ^ n21456 ^ 1'b0 ;
  assign n34429 = n7872 & n15411 ;
  assign n34430 = n32409 & n34429 ;
  assign n34427 = n3487 & n5776 ;
  assign n34428 = n34427 ^ n21458 ^ 1'b0 ;
  assign n34431 = n34430 ^ n34428 ^ 1'b0 ;
  assign n34432 = ~n19263 & n19388 ;
  assign n34433 = n31774 | n34432 ;
  assign n34434 = n288 & n11827 ;
  assign n34435 = n34434 ^ n68 ^ 1'b0 ;
  assign n34436 = n8198 ^ n3263 ^ 1'b0 ;
  assign n34437 = n12676 & n34436 ;
  assign n34438 = n14887 ^ n1309 ^ 1'b0 ;
  assign n34439 = ~n5573 & n34438 ;
  assign n34440 = n34439 ^ n11332 ^ 1'b0 ;
  assign n34441 = n19066 & ~n34440 ;
  assign n34442 = n11656 ^ n11205 ^ n7390 ;
  assign n34443 = n34442 ^ n11780 ^ 1'b0 ;
  assign n34444 = n5255 ^ n2640 ^ 1'b0 ;
  assign n34445 = n12723 & ~n34444 ;
  assign n34446 = n34445 ^ n7773 ^ 1'b0 ;
  assign n34447 = n18191 & ~n22657 ;
  assign n34448 = n2874 | n2933 ;
  assign n34449 = n12364 & n34448 ;
  assign n34450 = n6748 & ~n18552 ;
  assign n34451 = n34450 ^ n20313 ^ 1'b0 ;
  assign n34452 = n1403 & ~n34451 ;
  assign n34453 = n5657 ^ n2933 ^ 1'b0 ;
  assign n34454 = n3965 & ~n7231 ;
  assign n34455 = ~n378 & n19299 ;
  assign n34456 = n2493 | n3803 ;
  assign n34457 = n27022 & ~n34456 ;
  assign n34458 = n7715 & ~n9748 ;
  assign n34459 = n1794 | n34458 ;
  assign n34460 = n34457 | n34459 ;
  assign n34461 = n33218 ^ n2567 ^ 1'b0 ;
  assign n34462 = n30431 & n34461 ;
  assign n34463 = n133 & ~n33968 ;
  assign n34464 = n22239 & ~n32306 ;
  assign n34465 = ~n2120 & n34464 ;
  assign n34466 = n5112 | n5116 ;
  assign n34467 = n34466 ^ n2303 ^ 1'b0 ;
  assign n34468 = n31091 ^ n22118 ^ 1'b0 ;
  assign n34469 = ~n7288 & n12728 ;
  assign n34472 = n1229 | n19895 ;
  assign n34473 = n9335 & ~n34472 ;
  assign n34470 = n12865 ^ n6837 ^ 1'b0 ;
  assign n34471 = n6447 & n34470 ;
  assign n34474 = n34473 ^ n34471 ^ 1'b0 ;
  assign n34475 = ~n55 & n3939 ;
  assign n34476 = ~n520 & n34475 ;
  assign n34477 = n3373 | n10038 ;
  assign n34478 = n11034 | n34477 ;
  assign n34479 = ( n4054 & n7905 ) | ( n4054 & ~n16646 ) | ( n7905 & ~n16646 ) ;
  assign n34480 = n34478 & n34479 ;
  assign n34481 = n715 & ~n30269 ;
  assign n34482 = n30625 ^ n26930 ^ 1'b0 ;
  assign n34483 = n25790 | n34482 ;
  assign n34484 = n799 & ~n15786 ;
  assign n34485 = n34484 ^ n310 ^ 1'b0 ;
  assign n34486 = n10259 & n15495 ;
  assign n34487 = n34486 ^ n12730 ^ 1'b0 ;
  assign n34488 = n33262 & n34487 ;
  assign n34489 = n18216 & n23592 ;
  assign n34490 = n461 & ~n34489 ;
  assign n34491 = n4740 & ~n34490 ;
  assign n34492 = n2491 & n7231 ;
  assign n34493 = ~n294 & n993 ;
  assign n34494 = n7480 & n34493 ;
  assign n34495 = n113 & n18439 ;
  assign n34496 = n25078 ^ n128 ^ 1'b0 ;
  assign n34497 = n34495 & ~n34496 ;
  assign n34498 = n950 & ~n963 ;
  assign n34499 = n34498 ^ n24389 ^ 1'b0 ;
  assign n34500 = n8062 ^ n302 ^ n47 ;
  assign n34501 = ~n18226 & n34500 ;
  assign n34502 = n7928 & ~n8749 ;
  assign n34503 = n12982 | n34502 ;
  assign n34504 = n34503 ^ n6958 ^ 1'b0 ;
  assign n34505 = ~n159 & n3718 ;
  assign n34506 = n1836 | n25456 ;
  assign n34507 = n18507 & ~n23290 ;
  assign n34508 = n34507 ^ n24659 ^ 1'b0 ;
  assign n34509 = n12883 & n34508 ;
  assign n34510 = n19202 | n29299 ;
  assign n34511 = n9620 & ~n25485 ;
  assign n34512 = n34511 ^ n12473 ^ 1'b0 ;
  assign n34516 = ~n1988 & n4951 ;
  assign n34513 = n18847 ^ n14701 ^ n5554 ;
  assign n34514 = n10927 & ~n34513 ;
  assign n34515 = n1833 | n34514 ;
  assign n34517 = n34516 ^ n34515 ^ 1'b0 ;
  assign n34518 = ~n24032 & n34517 ;
  assign n34519 = n5958 & n11126 ;
  assign n34520 = ~n5643 & n34519 ;
  assign n34521 = n34520 ^ n9645 ^ 1'b0 ;
  assign n34522 = n20488 | n34521 ;
  assign n34523 = n32992 | n34522 ;
  assign n34524 = ~n5675 & n22497 ;
  assign n34525 = n29175 & n34524 ;
  assign n34526 = n4797 & n16448 ;
  assign n34527 = n602 & ~n16651 ;
  assign n34529 = n6225 & ~n14907 ;
  assign n34528 = ~n10590 & n15748 ;
  assign n34530 = n34529 ^ n34528 ^ 1'b0 ;
  assign n34531 = n6364 ^ n2591 ^ 1'b0 ;
  assign n34532 = ~n21199 & n32335 ;
  assign n34533 = n34532 ^ n1555 ^ 1'b0 ;
  assign n34534 = n24232 ^ n167 ^ 1'b0 ;
  assign n34535 = n24575 & n34534 ;
  assign n34536 = n1227 & n2480 ;
  assign n34537 = n34536 ^ n4848 ^ 1'b0 ;
  assign n34538 = ~n1355 & n9304 ;
  assign n34539 = n34538 ^ n1404 ^ 1'b0 ;
  assign n34540 = ~n2556 & n34539 ;
  assign n34541 = n34540 ^ n3352 ^ 1'b0 ;
  assign n34542 = n4526 & ~n10105 ;
  assign n34543 = n8922 ^ n4010 ^ 1'b0 ;
  assign n34544 = n34543 ^ n17875 ^ 1'b0 ;
  assign n34545 = n9712 & ~n34544 ;
  assign n34546 = n16887 | n29793 ;
  assign n34547 = n5567 | n34546 ;
  assign n34548 = n31405 ^ n15989 ^ 1'b0 ;
  assign n34549 = n13034 | n34548 ;
  assign n34550 = n5102 ^ n3443 ^ n323 ;
  assign n34551 = n34550 ^ n32951 ^ 1'b0 ;
  assign n34552 = n7669 & n9349 ;
  assign n34553 = ~n2771 & n34552 ;
  assign n34554 = ~n356 & n4921 ;
  assign n34555 = ~n9461 & n33923 ;
  assign n34556 = n19716 | n23649 ;
  assign n34557 = n17750 & ~n34556 ;
  assign n34558 = n7285 & ~n17802 ;
  assign n34559 = ~n1175 & n34558 ;
  assign n34560 = ~n10447 & n34559 ;
  assign n34561 = ~n6674 & n33823 ;
  assign n34562 = n30311 & ~n34561 ;
  assign n34563 = n34562 ^ n364 ^ 1'b0 ;
  assign n34564 = n5811 & n34563 ;
  assign n34565 = n13715 | n20967 ;
  assign n34566 = n12320 ^ n142 ^ 1'b0 ;
  assign n34567 = ~n11205 & n34566 ;
  assign n34568 = n34567 ^ n27361 ^ 1'b0 ;
  assign n34569 = n34565 | n34568 ;
  assign n34570 = ~n2744 & n4531 ;
  assign n34571 = n11117 | n17118 ;
  assign n34572 = n30874 ^ n178 ^ 1'b0 ;
  assign n34573 = n8047 ^ n404 ^ 1'b0 ;
  assign n34574 = ~n6286 & n18133 ;
  assign n34575 = n34574 ^ n33585 ^ 1'b0 ;
  assign n34576 = n324 & n25472 ;
  assign n34577 = n20292 | n23217 ;
  assign n34578 = n158 & ~n34577 ;
  assign n34579 = n525 | n1135 ;
  assign n34580 = n34579 ^ n5398 ^ 1'b0 ;
  assign n34581 = n8445 | n34580 ;
  assign n34582 = n34581 ^ n15655 ^ 1'b0 ;
  assign n34583 = n27399 & n29621 ;
  assign n34584 = n37 & ~n142 ;
  assign n34585 = ~n37 & n34584 ;
  assign n34586 = n481 | n34585 ;
  assign n34587 = n34585 & ~n34586 ;
  assign n34588 = ~n296 & n2028 ;
  assign n34589 = n296 & n34588 ;
  assign n34590 = n677 | n17409 ;
  assign n34591 = n677 & ~n34590 ;
  assign n34592 = n661 | n34591 ;
  assign n34593 = n661 & ~n34592 ;
  assign n34594 = n2328 | n34593 ;
  assign n34595 = n34589 & ~n34594 ;
  assign n34596 = ~n34587 & n34595 ;
  assign n34599 = n236 & n527 ;
  assign n34600 = ~n236 & n34599 ;
  assign n34601 = n2621 & ~n34600 ;
  assign n34602 = n34600 & n34601 ;
  assign n34597 = n1937 & n6596 ;
  assign n34598 = ~n1937 & n34597 ;
  assign n34603 = n34602 ^ n34598 ^ 1'b0 ;
  assign n34604 = ~n1172 & n2670 ;
  assign n34605 = ~n34603 & n34604 ;
  assign n34606 = n34596 & n34605 ;
  assign n34607 = n34606 ^ n941 ^ 1'b0 ;
  assign n34608 = ~n5428 & n7069 ;
  assign n34609 = n19333 ^ n6102 ^ 1'b0 ;
  assign n34610 = n17879 & n34609 ;
  assign n34611 = n25455 | n34610 ;
  assign n34612 = n19639 | n34611 ;
  assign n34613 = ~n5206 & n29096 ;
  assign n34614 = n34038 ^ n10588 ^ n1765 ;
  assign n34615 = n18474 | n28341 ;
  assign n34616 = n9870 & ~n10293 ;
  assign n34617 = n4131 & n34616 ;
  assign n34618 = n11041 & n34617 ;
  assign n34621 = n13788 ^ n501 ^ 1'b0 ;
  assign n34619 = n5632 & n20255 ;
  assign n34620 = ~n1304 & n34619 ;
  assign n34622 = n34621 ^ n34620 ^ 1'b0 ;
  assign n34623 = n14433 ^ n9699 ^ 1'b0 ;
  assign n34624 = n13908 & ~n34623 ;
  assign n34625 = n34624 ^ n7523 ^ 1'b0 ;
  assign n34626 = n19838 | n34625 ;
  assign n34627 = n34622 | n34626 ;
  assign n34628 = n1708 | n2410 ;
  assign n34629 = n34628 ^ n2938 ^ 1'b0 ;
  assign n34630 = n34629 ^ n8963 ^ 1'b0 ;
  assign n34631 = ~n1078 & n34630 ;
  assign n34632 = n34631 ^ n2514 ^ 1'b0 ;
  assign n34633 = n13864 | n34632 ;
  assign n34634 = n5421 | n34633 ;
  assign n34635 = n34634 ^ n10749 ^ 1'b0 ;
  assign n34636 = n34635 ^ n258 ^ 1'b0 ;
  assign n34637 = n2991 | n11012 ;
  assign n34638 = n9709 & ~n34637 ;
  assign n34639 = ( ~n8769 & n17021 ) | ( ~n8769 & n20666 ) | ( n17021 & n20666 ) ;
  assign n34640 = ~n10083 & n34639 ;
  assign n34641 = n34640 ^ n14046 ^ 1'b0 ;
  assign n34642 = n7355 & ~n7926 ;
  assign n34643 = n34642 ^ n21481 ^ n128 ;
  assign n34644 = n34643 ^ n19258 ^ n8475 ;
  assign n34645 = n9923 ^ n3036 ^ 1'b0 ;
  assign n34646 = n34529 & n34645 ;
  assign n34647 = x3 | n25851 ;
  assign n34648 = n21529 & ~n34647 ;
  assign n34649 = n7789 ^ n2170 ^ 1'b0 ;
  assign n34650 = n8652 & ~n34649 ;
  assign n34651 = ( n1217 & ~n5443 ) | ( n1217 & n9589 ) | ( ~n5443 & n9589 ) ;
  assign n34652 = n12560 ^ n6642 ^ 1'b0 ;
  assign n34653 = n27727 | n34652 ;
  assign n34654 = ( n883 & n34651 ) | ( n883 & ~n34653 ) | ( n34651 & ~n34653 ) ;
  assign n34655 = n34650 & ~n34654 ;
  assign n34656 = n11479 ^ n11355 ^ 1'b0 ;
  assign n34657 = n31815 & ~n34656 ;
  assign n34658 = n30600 ^ n23309 ^ 1'b0 ;
  assign n34659 = n26800 ^ n10533 ^ 1'b0 ;
  assign n34660 = n17039 ^ n14378 ^ 1'b0 ;
  assign n34661 = n15066 ^ n2784 ^ 1'b0 ;
  assign n34662 = n24088 ^ n8382 ^ 1'b0 ;
  assign n34663 = n1080 ^ n462 ^ 1'b0 ;
  assign n34664 = n6031 | n34663 ;
  assign n34665 = n25202 ^ n9253 ^ 1'b0 ;
  assign n34666 = n34665 ^ n18264 ^ 1'b0 ;
  assign n34667 = n10053 & n34666 ;
  assign n34668 = n6263 ^ n1106 ^ 1'b0 ;
  assign n34669 = n14001 & n34668 ;
  assign n34670 = n34669 ^ n2597 ^ 1'b0 ;
  assign n34671 = n30078 ^ n3720 ^ 1'b0 ;
  assign n34672 = ~n4131 & n34671 ;
  assign n34673 = n3087 & n8312 ;
  assign n34674 = ~n34672 & n34673 ;
  assign n34675 = n10851 | n34674 ;
  assign n34678 = n23320 ^ n272 ^ 1'b0 ;
  assign n34679 = n1467 & n34678 ;
  assign n34676 = n1818 & n33252 ;
  assign n34677 = ~n627 & n34676 ;
  assign n34680 = n34679 ^ n34677 ^ 1'b0 ;
  assign n34681 = ~n1438 & n24271 ;
  assign n34682 = n34681 ^ n19906 ^ 1'b0 ;
  assign n34683 = n32808 & ~n34682 ;
  assign n34684 = n34683 ^ n22135 ^ 1'b0 ;
  assign n34685 = n12234 ^ n4328 ^ 1'b0 ;
  assign n34686 = n6217 & n34685 ;
  assign n34687 = n34686 ^ n98 ^ 1'b0 ;
  assign n34688 = n19716 | n24869 ;
  assign n34689 = ~n2531 & n3576 ;
  assign n34690 = ~n8657 & n34689 ;
  assign n34691 = n497 & ~n5856 ;
  assign n34692 = ~n497 & n34691 ;
  assign n34693 = n34692 ^ n16 ^ 1'b0 ;
  assign n34694 = n274 | n294 ;
  assign n34695 = n274 & ~n34694 ;
  assign n34696 = n1175 & n9947 ;
  assign n34697 = n475 & n34696 ;
  assign n34698 = n2027 & ~n34697 ;
  assign n34699 = ~n34695 & n34698 ;
  assign n34700 = n34699 ^ n9112 ^ 1'b0 ;
  assign n34701 = n34693 & ~n34700 ;
  assign n34702 = n34701 ^ n5573 ^ 1'b0 ;
  assign n34703 = n9775 & ~n34702 ;
  assign n34704 = n14232 ^ n83 ^ 1'b0 ;
  assign n34705 = n29144 & n34704 ;
  assign n34706 = n408 | n11228 ;
  assign n34707 = n33706 ^ n3014 ^ 1'b0 ;
  assign n34708 = n7797 ^ n3871 ^ 1'b0 ;
  assign n34709 = n34226 & n34708 ;
  assign n34710 = n34709 ^ n4281 ^ 1'b0 ;
  assign n34714 = n26988 ^ n7870 ^ 1'b0 ;
  assign n34715 = ~n19426 & n34714 ;
  assign n34711 = n31728 ^ n31219 ^ 1'b0 ;
  assign n34712 = n34711 ^ n8353 ^ 1'b0 ;
  assign n34713 = x0 | n34712 ;
  assign n34716 = n34715 ^ n34713 ^ 1'b0 ;
  assign n34717 = n17568 ^ n16393 ^ 1'b0 ;
  assign n34718 = n18509 & n34717 ;
  assign n34721 = n21007 ^ n4495 ^ 1'b0 ;
  assign n34722 = n21303 | n34721 ;
  assign n34723 = n8446 ^ n8000 ^ 1'b0 ;
  assign n34724 = n34722 | n34723 ;
  assign n34725 = n34724 ^ n1666 ^ 1'b0 ;
  assign n34726 = n15808 & ~n34725 ;
  assign n34719 = n26415 ^ n231 ^ 1'b0 ;
  assign n34720 = n11348 & ~n34719 ;
  assign n34727 = n34726 ^ n34720 ^ 1'b0 ;
  assign n34728 = n319 & ~n4703 ;
  assign n34729 = n779 | n1467 ;
  assign n34730 = n13159 & ~n34729 ;
  assign n34731 = n34730 ^ n5771 ^ 1'b0 ;
  assign n34732 = ~n34728 & n34731 ;
  assign n34733 = n34280 ^ n6670 ^ 1'b0 ;
  assign n34734 = n6323 | n34733 ;
  assign n34735 = n6356 & ~n21354 ;
  assign n34736 = ~n14235 & n34711 ;
  assign n34737 = n19012 & n31637 ;
  assign n34738 = n34737 ^ n3146 ^ 1'b0 ;
  assign n34739 = n12347 & n34738 ;
  assign n34740 = n34739 ^ n10346 ^ 1'b0 ;
  assign n34741 = n142 & ~n15366 ;
  assign n34742 = ~n10486 & n34741 ;
  assign n34743 = n34742 ^ n2699 ^ 1'b0 ;
  assign n34744 = n255 & ~n34743 ;
  assign n34745 = n21774 & ~n33294 ;
  assign n34746 = ( n18192 & n27223 ) | ( n18192 & ~n34745 ) | ( n27223 & ~n34745 ) ;
  assign n34747 = n1718 | n18274 ;
  assign n34748 = n17563 ^ n8099 ^ 1'b0 ;
  assign n34749 = n34748 ^ n489 ^ 1'b0 ;
  assign n34750 = ( n823 & n6933 ) | ( n823 & n34749 ) | ( n6933 & n34749 ) ;
  assign n34751 = ~n3280 & n24567 ;
  assign n34752 = n34751 ^ n3247 ^ 1'b0 ;
  assign n34753 = n19257 ^ n2594 ^ 1'b0 ;
  assign n34754 = ~n8139 & n34091 ;
  assign n34755 = n3291 & n13118 ;
  assign n34756 = n2456 & n34755 ;
  assign n34757 = n10527 | n16635 ;
  assign n34758 = n34757 ^ n5933 ^ 1'b0 ;
  assign n34759 = n34758 ^ n10813 ^ 1'b0 ;
  assign n34760 = n533 & n34759 ;
  assign n34761 = n34756 & n34760 ;
  assign n34762 = n34754 | n34761 ;
  assign n34763 = n2199 | n16195 ;
  assign n34764 = n9552 & n18003 ;
  assign n34765 = n8047 | n12207 ;
  assign n34766 = n34765 ^ n417 ^ 1'b0 ;
  assign n34767 = n3118 & ~n9758 ;
  assign n34768 = ~n1976 & n2034 ;
  assign n34769 = n142 & n34768 ;
  assign n34770 = ( n9775 & n27497 ) | ( n9775 & ~n34769 ) | ( n27497 & ~n34769 ) ;
  assign n34771 = n5643 & n6249 ;
  assign n34772 = n34771 ^ n4036 ^ 1'b0 ;
  assign n34773 = n21221 | n26777 ;
  assign n34774 = n34773 ^ n1598 ^ 1'b0 ;
  assign n34775 = n18435 | n28808 ;
  assign n34776 = n34775 ^ n14253 ^ 1'b0 ;
  assign n34777 = ~n5714 & n34776 ;
  assign n34778 = n15866 ^ n13110 ^ 1'b0 ;
  assign n34779 = n8914 | n34778 ;
  assign n34780 = n23611 ^ n22163 ^ 1'b0 ;
  assign n34781 = ( ~n5087 & n5685 ) | ( ~n5087 & n28114 ) | ( n5685 & n28114 ) ;
  assign n34782 = n17733 & ~n34781 ;
  assign n34783 = n1774 ^ n497 ^ 1'b0 ;
  assign n34784 = n34783 ^ n12867 ^ 1'b0 ;
  assign n34785 = n8282 & n34784 ;
  assign n34786 = n34785 ^ n25414 ^ 1'b0 ;
  assign n34787 = ~n13574 & n34786 ;
  assign n34788 = n294 & n22733 ;
  assign n34789 = ~n4098 & n5125 ;
  assign n34790 = n713 | n18912 ;
  assign n34791 = ~n13310 & n34790 ;
  assign n34792 = n34514 ^ n3178 ^ 1'b0 ;
  assign n34793 = n609 & n9231 ;
  assign n34794 = n34792 & n34793 ;
  assign n34795 = n26381 ^ n11659 ^ 1'b0 ;
  assign n34796 = n13751 & n26711 ;
  assign n34797 = n18490 & n34796 ;
  assign n34798 = ~n158 & n30750 ;
  assign n34799 = n34798 ^ n28936 ^ 1'b0 ;
  assign n34800 = ~n4419 & n34799 ;
  assign n34801 = n15526 & n22835 ;
  assign n34802 = ~n627 & n34801 ;
  assign n34803 = n1052 & ~n8218 ;
  assign n34804 = ~n17502 & n34803 ;
  assign n34805 = n1814 | n34804 ;
  assign n34806 = n25506 ^ n13727 ^ 1'b0 ;
  assign n34807 = n6200 | n34806 ;
  assign n34808 = n34805 & n34807 ;
  assign n34809 = n24635 ^ n14808 ^ 1'b0 ;
  assign n34810 = n7380 & n22912 ;
  assign n34811 = n20017 ^ n15179 ^ 1'b0 ;
  assign n34812 = n1246 ^ n364 ^ 1'b0 ;
  assign n34813 = n25510 | n34812 ;
  assign n34814 = n2018 & ~n13199 ;
  assign n34815 = n7520 | n16006 ;
  assign n34816 = n34814 & ~n34815 ;
  assign n34817 = ~n8460 & n11180 ;
  assign n34818 = n34817 ^ n27856 ^ 1'b0 ;
  assign n34819 = n6689 & ~n34818 ;
  assign n34820 = n34819 ^ n9733 ^ 1'b0 ;
  assign n34821 = n14911 & n29852 ;
  assign n34822 = n31757 ^ n29116 ^ 1'b0 ;
  assign n34823 = n6667 & n24406 ;
  assign n34824 = n34823 ^ n8714 ^ 1'b0 ;
  assign n34825 = n12383 ^ n1593 ^ 1'b0 ;
  assign n34826 = n34824 & n34825 ;
  assign n34827 = ~n3437 & n3671 ;
  assign n34828 = ( ~n1631 & n7391 ) | ( ~n1631 & n34827 ) | ( n7391 & n34827 ) ;
  assign n34829 = n1565 | n12345 ;
  assign n34830 = ~n175 & n581 ;
  assign n34831 = n3339 & n34830 ;
  assign n34832 = n2719 | n34831 ;
  assign n34833 = n2757 | n34832 ;
  assign n34834 = n709 & n34833 ;
  assign n34835 = n34834 ^ n500 ^ 1'b0 ;
  assign n34836 = ~n26735 & n34835 ;
  assign n34837 = n1550 & n29856 ;
  assign n34838 = n25063 & n34837 ;
  assign n34839 = n29345 ^ n8279 ^ 1'b0 ;
  assign n34840 = n7581 | n26207 ;
  assign n34841 = n9934 | n34840 ;
  assign n34842 = n34841 ^ n9242 ^ 1'b0 ;
  assign n34843 = n1992 & ~n14970 ;
  assign n34844 = n34843 ^ n24164 ^ 1'b0 ;
  assign n34845 = n21049 ^ n19304 ^ n10879 ;
  assign n34846 = ~n33123 & n34845 ;
  assign n34847 = n4482 & n16906 ;
  assign n34848 = ~n34755 & n34847 ;
  assign n34849 = n10589 | n33823 ;
  assign n34850 = n21145 | n31049 ;
  assign n34851 = n34850 ^ n18385 ^ 1'b0 ;
  assign n34852 = n2509 | n34851 ;
  assign n34853 = n27715 ^ n947 ^ 1'b0 ;
  assign n34854 = n3262 | n34853 ;
  assign n34855 = ( ~n7548 & n14056 ) | ( ~n7548 & n15883 ) | ( n14056 & n15883 ) ;
  assign n34856 = n11775 & ~n34855 ;
  assign n34857 = n14902 ^ n12679 ^ 1'b0 ;
  assign n34858 = n14001 & ~n34857 ;
  assign n34859 = ~n1315 & n5317 ;
  assign n34860 = n9727 ^ n2041 ^ 1'b0 ;
  assign n34861 = n16906 ^ n3804 ^ 1'b0 ;
  assign n34862 = ~n1763 & n13752 ;
  assign n34863 = n4970 & n34862 ;
  assign n34864 = n9492 & ~n34863 ;
  assign n34865 = n34864 ^ n25416 ^ n23788 ;
  assign n34866 = n14184 ^ n1885 ^ 1'b0 ;
  assign n34867 = ~n62 & n25951 ;
  assign n34868 = n34867 ^ n12455 ^ 1'b0 ;
  assign n34869 = n29903 ^ n6023 ^ n3374 ;
  assign n34870 = n12303 ^ n5934 ^ 1'b0 ;
  assign n34871 = n11283 & ~n34870 ;
  assign n34872 = n26602 ^ n24353 ^ 1'b0 ;
  assign n34873 = ~n3990 & n34872 ;
  assign n34874 = n4334 | n10547 ;
  assign n34875 = n13859 ^ n1587 ^ 1'b0 ;
  assign n34876 = n2470 & n14645 ;
  assign n34877 = n9340 ^ n4855 ^ 1'b0 ;
  assign n34878 = n185 & ~n11882 ;
  assign n34879 = n34878 ^ n318 ^ 1'b0 ;
  assign n34880 = n34879 ^ n1399 ^ 1'b0 ;
  assign n34881 = n34877 & n34880 ;
  assign n34882 = n19438 ^ n17891 ^ 1'b0 ;
  assign n34883 = n50 & n2403 ;
  assign n34884 = n34882 & n34883 ;
  assign n34885 = n322 ^ n213 ^ 1'b0 ;
  assign n34886 = n756 & n27943 ;
  assign n34887 = n34886 ^ n213 ^ 1'b0 ;
  assign n34888 = n22387 | n34887 ;
  assign n34889 = n34888 ^ n31946 ^ 1'b0 ;
  assign n34890 = n1370 & n28734 ;
  assign n34891 = n17794 ^ n15426 ^ 1'b0 ;
  assign n34892 = n2059 | n34891 ;
  assign n34893 = ~n12444 & n24287 ;
  assign n34894 = n34893 ^ n33060 ^ n4668 ;
  assign n34896 = n1086 & ~n26453 ;
  assign n34897 = n34896 ^ n22556 ^ n14713 ;
  assign n34898 = n3974 & n34897 ;
  assign n34899 = n7523 & n34898 ;
  assign n34900 = n34899 ^ n24720 ^ 1'b0 ;
  assign n34895 = ~n19761 & n30750 ;
  assign n34901 = n34900 ^ n34895 ^ 1'b0 ;
  assign n34902 = n17039 ^ n11977 ^ 1'b0 ;
  assign n34903 = n19050 ^ n758 ^ 1'b0 ;
  assign n34904 = n29096 ^ n23218 ^ 1'b0 ;
  assign n34905 = n4306 ^ n183 ^ 1'b0 ;
  assign n34906 = n26504 ^ n23229 ^ 1'b0 ;
  assign n34907 = n12295 ^ n1425 ^ 1'b0 ;
  assign n34908 = ~n10470 & n13841 ;
  assign n34909 = n34908 ^ n9853 ^ 1'b0 ;
  assign n34910 = n34909 ^ n34178 ^ 1'b0 ;
  assign n34911 = n29437 & ~n30269 ;
  assign n34912 = ~n9906 & n34911 ;
  assign n34913 = n30952 ^ n29480 ^ 1'b0 ;
  assign n34933 = n7377 & n25526 ;
  assign n34934 = ~n7377 & n34933 ;
  assign n34932 = n26405 | n29359 ;
  assign n34935 = n34934 ^ n34932 ^ 1'b0 ;
  assign n34914 = n2587 & n5846 ;
  assign n34915 = ~n5846 & n34914 ;
  assign n34916 = ~n9008 & n34915 ;
  assign n34917 = n58 & n9046 ;
  assign n34918 = n2800 | n34917 ;
  assign n34919 = n34917 & ~n34918 ;
  assign n34920 = ~n1112 & n1345 ;
  assign n34921 = ~n1345 & n34920 ;
  assign n34922 = n2092 & n8622 ;
  assign n34923 = ~n2092 & n34922 ;
  assign n34924 = n5535 | n34923 ;
  assign n34925 = n5535 & ~n34924 ;
  assign n34926 = n34921 & ~n34925 ;
  assign n34927 = ~n34919 & n34926 ;
  assign n34928 = n13461 & n34927 ;
  assign n34929 = n34928 ^ n4544 ^ 1'b0 ;
  assign n34930 = ~n34916 & n34929 ;
  assign n34931 = ~n24891 & n34930 ;
  assign n34936 = n34935 ^ n34931 ^ 1'b0 ;
  assign n34937 = n13463 ^ n1036 ^ 1'b0 ;
  assign n34938 = n169 | n34937 ;
  assign n34939 = n179 | n16981 ;
  assign n34940 = n3001 | n32770 ;
  assign n34941 = n17814 | n34940 ;
  assign n34942 = n8409 ^ n241 ^ 1'b0 ;
  assign n34943 = n34941 & n34942 ;
  assign n34944 = n684 | n1707 ;
  assign n34945 = n34944 ^ n13688 ^ 1'b0 ;
  assign n34946 = n4799 ^ n165 ^ 1'b0 ;
  assign n34947 = n1888 | n5974 ;
  assign n34948 = n34947 ^ n13967 ^ 1'b0 ;
  assign n34949 = n18014 ^ n2220 ^ 1'b0 ;
  assign n34950 = ~n34948 & n34949 ;
  assign n34951 = ~n2321 & n6476 ;
  assign n34952 = n24300 & n34951 ;
  assign n34953 = ~n8653 & n28848 ;
  assign n34954 = n34953 ^ n1518 ^ 1'b0 ;
  assign n34955 = n2060 ^ n83 ^ 1'b0 ;
  assign n34956 = n27504 & n34955 ;
  assign n34957 = n4883 | n5144 ;
  assign n34958 = n541 & ~n15814 ;
  assign n34959 = n19332 & n34958 ;
  assign n34960 = n34959 ^ n2140 ^ 1'b0 ;
  assign n34961 = n5053 & ~n34447 ;
  assign n34962 = n5330 ^ n3333 ^ 1'b0 ;
  assign n34963 = n34962 ^ n17135 ^ 1'b0 ;
  assign n34964 = n4303 & n34963 ;
  assign n34965 = n17737 & n19681 ;
  assign n34966 = n30507 ^ n22485 ^ 1'b0 ;
  assign n34967 = n364 & n34966 ;
  assign n34968 = n18278 ^ n14455 ^ 1'b0 ;
  assign n34969 = n29022 & n34968 ;
  assign n34970 = ~n12194 & n34969 ;
  assign n34971 = n10239 & n12502 ;
  assign n34972 = n34971 ^ n21444 ^ 1'b0 ;
  assign n34973 = n25079 ^ n16102 ^ 1'b0 ;
  assign n34974 = n5972 & ~n11333 ;
  assign n34975 = n16728 & n29154 ;
  assign n34976 = n2541 & n34975 ;
  assign n34977 = n34976 ^ n26419 ^ 1'b0 ;
  assign n34978 = n4210 & ~n34977 ;
  assign n34979 = n522 & n9004 ;
  assign n34980 = n4349 | n34979 ;
  assign n34981 = n34980 ^ n2792 ^ 1'b0 ;
  assign n34982 = n11768 | n34981 ;
  assign n34983 = n17583 & ~n34982 ;
  assign n34984 = n3038 & ~n3520 ;
  assign n34985 = n34984 ^ n2865 ^ 1'b0 ;
  assign n34986 = n10660 | n34985 ;
  assign n34987 = ~n64 & n15729 ;
  assign n34988 = ~n3081 & n34987 ;
  assign n34989 = ~n2410 & n34988 ;
  assign n34990 = n2410 & n34989 ;
  assign n34991 = n34990 ^ n7497 ^ n2339 ;
  assign n34992 = n34991 ^ n10433 ^ 1'b0 ;
  assign n34993 = ~n8363 & n9216 ;
  assign n34994 = ~n34992 & n34993 ;
  assign n34995 = n7301 & n13168 ;
  assign n34996 = n4572 & n34995 ;
  assign n34997 = n34996 ^ n5256 ^ 1'b0 ;
  assign n34998 = n34997 ^ n16782 ^ 1'b0 ;
  assign n34999 = n22497 & n34998 ;
  assign n35000 = n34999 ^ n24857 ^ 1'b0 ;
  assign n35001 = ~n3085 & n14125 ;
  assign n35002 = n35001 ^ n743 ^ 1'b0 ;
  assign n35003 = n5700 & n35002 ;
  assign n35004 = n1867 | n1935 ;
  assign n35005 = n16703 | n35004 ;
  assign n35006 = n35003 | n35005 ;
  assign n35007 = n142 | n35006 ;
  assign n35008 = n5393 & ~n24315 ;
  assign n35009 = ~n4273 & n23400 ;
  assign n35010 = n21805 ^ n19159 ^ 1'b0 ;
  assign n35011 = n27911 ^ n13165 ^ 1'b0 ;
  assign n35012 = ~n35010 & n35011 ;
  assign n35013 = n3436 & n12205 ;
  assign n35014 = ~n19163 & n35013 ;
  assign n35015 = n5241 | n19179 ;
  assign n35016 = n25241 & n27722 ;
  assign n35017 = ~n13252 & n35016 ;
  assign n35018 = n2078 & n32080 ;
  assign n35019 = n19363 ^ n6322 ^ 1'b0 ;
  assign n35020 = n4019 & n20796 ;
  assign n35021 = n5399 & n35020 ;
  assign n35022 = n804 & ~n35021 ;
  assign n35023 = n1355 & ~n16945 ;
  assign n35024 = n5790 ^ n599 ^ 1'b0 ;
  assign n35025 = n19534 & ~n35024 ;
  assign n35026 = n25671 ^ n16532 ^ 1'b0 ;
  assign n35027 = n19136 ^ n5726 ^ 1'b0 ;
  assign n35028 = ~n4449 & n30107 ;
  assign n35029 = n5726 | n35028 ;
  assign n35030 = n9046 ^ n963 ^ 1'b0 ;
  assign n35031 = n33825 ^ n7927 ^ 1'b0 ;
  assign n35032 = n737 & ~n35031 ;
  assign n35033 = ~n4924 & n8068 ;
  assign n35034 = ~n3279 & n35033 ;
  assign n35035 = ( ~n227 & n9341 ) | ( ~n227 & n21584 ) | ( n9341 & n21584 ) ;
  assign n35036 = n2027 & n3957 ;
  assign n35037 = n35036 ^ n14141 ^ n4084 ;
  assign n35038 = ~n2341 & n35037 ;
  assign n35039 = n6185 | n19124 ;
  assign n35040 = ~n9811 & n12646 ;
  assign n35041 = ( n20005 & n20052 ) | ( n20005 & n35040 ) | ( n20052 & n35040 ) ;
  assign n35042 = n10239 ^ n2047 ^ 1'b0 ;
  assign n35043 = n35042 ^ n10444 ^ 1'b0 ;
  assign n35044 = ~n1337 & n16607 ;
  assign n35045 = n35044 ^ n23525 ^ 1'b0 ;
  assign n35046 = n9727 ^ n8282 ^ 1'b0 ;
  assign n35047 = ~n1827 & n7899 ;
  assign n35048 = n8230 | n35047 ;
  assign n35049 = n13724 | n19712 ;
  assign n35050 = n16972 ^ n2564 ^ 1'b0 ;
  assign n35051 = n11707 | n35050 ;
  assign n35052 = n16013 & n35051 ;
  assign n35053 = n35052 ^ n1555 ^ 1'b0 ;
  assign n35054 = n1887 & n35053 ;
  assign n35055 = n28838 ^ n23751 ^ 1'b0 ;
  assign n35056 = n1681 & ~n35055 ;
  assign n35057 = n3485 ^ n800 ^ 1'b0 ;
  assign n35058 = n107 & ~n13092 ;
  assign n35059 = n1051 & ~n20415 ;
  assign n35060 = n32436 & n35059 ;
  assign n35061 = n776 & n19882 ;
  assign n35062 = n35061 ^ n23551 ^ 1'b0 ;
  assign n35063 = n35060 & ~n35062 ;
  assign n35064 = n8299 & ~n20517 ;
  assign n35065 = n35064 ^ n8703 ^ 1'b0 ;
  assign n35066 = n6106 & ~n12728 ;
  assign n35067 = n5334 & ~n8175 ;
  assign n35068 = n13538 ^ n2283 ^ n1362 ;
  assign n35069 = n849 & ~n35068 ;
  assign n35070 = n3246 & ~n9492 ;
  assign n35071 = n5154 ^ n4903 ^ 1'b0 ;
  assign n35072 = n32492 | n35071 ;
  assign n35073 = n5045 ^ n799 ^ 1'b0 ;
  assign n35074 = n2573 & ~n35073 ;
  assign n35075 = n24889 & n28232 ;
  assign n35076 = n21525 & ~n26707 ;
  assign n35077 = ~n6338 & n19555 ;
  assign n35078 = ~n1149 & n35077 ;
  assign n35079 = ~n8022 & n22284 ;
  assign n35080 = ~n29882 & n35079 ;
  assign n35081 = n3935 | n23888 ;
  assign n35082 = n35081 ^ n12730 ^ 1'b0 ;
  assign n35083 = n5832 | n6072 ;
  assign n35084 = n35083 ^ n2612 ^ 1'b0 ;
  assign n35085 = n13073 ^ n4499 ^ n3638 ;
  assign n35086 = n35085 ^ n25638 ^ 1'b0 ;
  assign n35087 = n35084 | n35086 ;
  assign n35088 = n10022 ^ n4895 ^ 1'b0 ;
  assign n35089 = n1366 & ~n5573 ;
  assign n35090 = n26297 | n27723 ;
  assign n35091 = n35090 ^ n26635 ^ 1'b0 ;
  assign n35092 = n3801 ^ n37 ^ 1'b0 ;
  assign n35093 = n13194 & n24905 ;
  assign n35094 = n35093 ^ n10395 ^ 1'b0 ;
  assign n35095 = ~n3909 & n12219 ;
  assign n35096 = n35095 ^ n9120 ^ 1'b0 ;
  assign n35097 = n9619 | n13439 ;
  assign n35098 = n35096 | n35097 ;
  assign n35099 = n16017 | n32802 ;
  assign n35100 = n18387 ^ n14734 ^ 1'b0 ;
  assign n35101 = n14075 | n15983 ;
  assign n35102 = n17287 | n35101 ;
  assign n35103 = n30252 ^ n29161 ^ n23535 ;
  assign n35104 = n2185 | n21724 ;
  assign n35105 = n35104 ^ n4227 ^ 1'b0 ;
  assign n35106 = n142 & ~n12113 ;
  assign n35107 = n11539 & n35106 ;
  assign n35108 = ~n3670 & n17961 ;
  assign n35109 = n7940 | n35108 ;
  assign n35110 = n1000 | n23045 ;
  assign n35111 = n33832 | n35110 ;
  assign n35112 = n2782 ^ n116 ^ 1'b0 ;
  assign n35113 = n24769 & ~n35112 ;
  assign n35114 = n419 | n27371 ;
  assign n35115 = n3965 & ~n12039 ;
  assign n35116 = n11201 & n18729 ;
  assign n35117 = n703 & n16104 ;
  assign n35118 = n35117 ^ n13256 ^ 1'b0 ;
  assign n35120 = n11843 | n12519 ;
  assign n35119 = n342 & n1870 ;
  assign n35121 = n35120 ^ n35119 ^ 1'b0 ;
  assign n35122 = n35121 ^ n16320 ^ n9884 ;
  assign n35123 = n13034 ^ n556 ^ 1'b0 ;
  assign n35124 = ~n8067 & n10636 ;
  assign n35125 = ~n5462 & n35124 ;
  assign n35126 = n25025 ^ n3724 ^ 1'b0 ;
  assign n35127 = n11106 & n35126 ;
  assign n35128 = n2292 | n6906 ;
  assign n35129 = n6906 & ~n35128 ;
  assign n35130 = n5032 & ~n35129 ;
  assign n35131 = ~n5032 & n35130 ;
  assign n35132 = ~n16671 & n35131 ;
  assign n35133 = n684 & n8350 ;
  assign n35134 = n35132 & n35133 ;
  assign n35135 = n10608 ^ n1707 ^ 1'b0 ;
  assign n35136 = n7090 ^ n3304 ^ 1'b0 ;
  assign n35137 = n35135 & ~n35136 ;
  assign n35138 = n13640 & ~n34371 ;
  assign n35139 = n35138 ^ n2644 ^ 1'b0 ;
  assign n35140 = ~n26012 & n35139 ;
  assign n35141 = n21607 ^ n20894 ^ 1'b0 ;
  assign n35142 = ( n14714 & ~n24759 ) | ( n14714 & n25614 ) | ( ~n24759 & n25614 ) ;
  assign n35145 = n13573 ^ n2414 ^ 1'b0 ;
  assign n35146 = n7917 & n35145 ;
  assign n35147 = n35146 ^ n7055 ^ n6809 ;
  assign n35144 = ~n13167 & n15473 ;
  assign n35148 = n35147 ^ n35144 ^ 1'b0 ;
  assign n35143 = n5431 | n23449 ;
  assign n35149 = n35148 ^ n35143 ^ 1'b0 ;
  assign n35150 = n16007 & n35149 ;
  assign n35151 = n17962 ^ n17031 ^ 1'b0 ;
  assign n35152 = n29693 ^ n11334 ^ 1'b0 ;
  assign n35153 = n7504 | n35152 ;
  assign n35154 = n12295 ^ n1245 ^ 1'b0 ;
  assign n35155 = n26088 ^ n963 ^ 1'b0 ;
  assign n35156 = n4261 & n35155 ;
  assign n35157 = n35156 ^ n4295 ^ 1'b0 ;
  assign n35158 = n17078 ^ n6920 ^ 1'b0 ;
  assign n35159 = n35157 & ~n35158 ;
  assign n35160 = n8787 & n35159 ;
  assign n35161 = n12498 ^ n3530 ^ n847 ;
  assign n35162 = n16895 ^ n2068 ^ 1'b0 ;
  assign n35163 = n11235 | n19091 ;
  assign n35164 = n14813 | n35163 ;
  assign n35165 = n11451 ^ n10259 ^ n8611 ;
  assign n35166 = n6930 ^ n3110 ^ 1'b0 ;
  assign n35167 = n1847 & n35166 ;
  assign n35168 = n30664 & n35167 ;
  assign n35169 = n28622 ^ n17182 ^ 1'b0 ;
  assign n35170 = n18494 & n35169 ;
  assign n35171 = n29252 ^ n13960 ^ 1'b0 ;
  assign n35172 = n26634 ^ n4481 ^ 1'b0 ;
  assign n35173 = ~n1902 & n35172 ;
  assign n35174 = n28036 ^ n8349 ^ n2090 ;
  assign n35175 = n14232 ^ n2039 ^ 1'b0 ;
  assign n35176 = n7088 | n8047 ;
  assign n35177 = ~n1718 & n2701 ;
  assign n35178 = n19420 ^ n4906 ^ n1685 ;
  assign n35179 = n35178 ^ n6471 ^ 1'b0 ;
  assign n35180 = n22700 ^ n1118 ^ 1'b0 ;
  assign n35181 = n8675 ^ n6527 ^ 1'b0 ;
  assign n35182 = ~n724 & n13946 ;
  assign n35183 = n35182 ^ n7079 ^ 1'b0 ;
  assign n35184 = n24418 | n35183 ;
  assign n35185 = ( n11439 & n35181 ) | ( n11439 & ~n35184 ) | ( n35181 & ~n35184 ) ;
  assign n35186 = n35185 ^ n14190 ^ 1'b0 ;
  assign n35188 = n29918 ^ n9651 ^ 1'b0 ;
  assign n35187 = n14696 & n27424 ;
  assign n35189 = n35188 ^ n35187 ^ 1'b0 ;
  assign n35190 = n26609 & n29863 ;
  assign n35191 = n10470 ^ n2584 ^ n440 ;
  assign n35192 = n35191 ^ n3583 ^ 1'b0 ;
  assign n35193 = n5314 & ~n15252 ;
  assign n35194 = ~n1934 & n19450 ;
  assign n35195 = n184 & n9333 ;
  assign n35196 = n35195 ^ n14462 ^ 1'b0 ;
  assign n35197 = n16589 & n27412 ;
  assign n35198 = ~n35196 & n35197 ;
  assign n35199 = ~n4550 & n9401 ;
  assign n35200 = n16506 & n35199 ;
  assign n35201 = n35198 & n35200 ;
  assign n35202 = n34109 ^ n24308 ^ 1'b0 ;
  assign n35203 = n14513 & ~n25941 ;
  assign n35204 = n35203 ^ n6194 ^ 1'b0 ;
  assign n35205 = ~n13688 & n28139 ;
  assign n35206 = n20454 ^ n748 ^ 1'b0 ;
  assign n35207 = n16296 & n24090 ;
  assign n35208 = n35207 ^ n23381 ^ 1'b0 ;
  assign n35209 = n3258 & n14793 ;
  assign n35210 = n35209 ^ n1633 ^ 1'b0 ;
  assign n35211 = n6399 & n35210 ;
  assign n35212 = n8841 & ~n8999 ;
  assign n35213 = n9242 & n35212 ;
  assign n35214 = n35213 ^ n6176 ^ 1'b0 ;
  assign n35215 = n11950 & n35214 ;
  assign n35216 = n8171 & ~n31962 ;
  assign n35217 = n5338 & n35216 ;
  assign n35218 = n11122 | n19333 ;
  assign n35219 = n3533 | n35218 ;
  assign n35220 = n4706 & n14724 ;
  assign n35221 = n582 | n35220 ;
  assign n35222 = n2853 ^ n300 ^ 1'b0 ;
  assign n35223 = n1714 | n35222 ;
  assign n35224 = n3776 & ~n35223 ;
  assign n35225 = n30565 ^ n17013 ^ 1'b0 ;
  assign n35226 = n17163 & ~n35225 ;
  assign n35227 = n7844 ^ n2728 ^ 1'b0 ;
  assign n35228 = n5970 & n26110 ;
  assign n35229 = n35228 ^ n414 ^ 1'b0 ;
  assign n35230 = n33874 ^ n11042 ^ 1'b0 ;
  assign n35231 = n12646 & n35230 ;
  assign n35232 = n6349 | n9357 ;
  assign n35233 = n6349 & ~n35232 ;
  assign n35234 = n2945 | n35233 ;
  assign n35235 = n2945 & ~n35234 ;
  assign n35236 = n33108 & ~n35235 ;
  assign n35237 = n35236 ^ n31079 ^ n24036 ;
  assign n35238 = ~n4406 & n15072 ;
  assign n35239 = n187 & ~n6145 ;
  assign n35240 = n5045 & ~n5982 ;
  assign n35241 = ~n35239 & n35240 ;
  assign n35242 = n24404 & n35241 ;
  assign n35243 = ( n5542 & n16274 ) | ( n5542 & ~n23158 ) | ( n16274 & ~n23158 ) ;
  assign n35244 = n11047 & ~n11797 ;
  assign n35245 = n9709 | n19175 ;
  assign n35246 = n33720 ^ n3843 ^ 1'b0 ;
  assign n35247 = ~n35245 & n35246 ;
  assign n35249 = n3295 & n10971 ;
  assign n35248 = ~n1112 & n1370 ;
  assign n35250 = n35249 ^ n35248 ^ n27234 ;
  assign n35251 = n1048 & n3812 ;
  assign n35252 = ~n1486 & n35251 ;
  assign n35253 = n15368 | n19968 ;
  assign n35254 = ~n3718 & n8657 ;
  assign n35255 = n28584 & n35254 ;
  assign n35256 = ~n1611 & n6713 ;
  assign n35257 = ~n1947 & n3744 ;
  assign n35258 = n35256 & n35257 ;
  assign n35259 = ~n1065 & n31101 ;
  assign n35260 = n11840 & n14212 ;
  assign n35261 = n32275 & n35260 ;
  assign n35262 = ~n20270 & n35261 ;
  assign n35263 = n34408 & ~n35262 ;
  assign n35264 = n191 & ~n9840 ;
  assign n35265 = n33256 ^ n3853 ^ 1'b0 ;
  assign n35266 = n19356 & ~n35265 ;
  assign n35267 = n3464 & n12676 ;
  assign n35268 = n7784 ^ n4918 ^ 1'b0 ;
  assign n35269 = n13878 | n16525 ;
  assign n35270 = ~n1465 & n17019 ;
  assign n35271 = ~n21937 & n35270 ;
  assign n35272 = n35271 ^ n20478 ^ 1'b0 ;
  assign n35273 = ~n3589 & n3925 ;
  assign n35275 = n16529 & n35002 ;
  assign n35274 = n12672 & ~n31657 ;
  assign n35276 = n35275 ^ n35274 ^ 1'b0 ;
  assign n35277 = n18181 & n23616 ;
  assign n35278 = n415 | n35277 ;
  assign n35279 = n18181 & ~n33850 ;
  assign n35280 = n24428 ^ n5543 ^ 1'b0 ;
  assign n35281 = ~n17935 & n35280 ;
  assign n35282 = n29629 ^ n21204 ^ 1'b0 ;
  assign n35283 = n1090 & ~n35282 ;
  assign n35284 = ~n837 & n14622 ;
  assign n35285 = n22597 & ~n24049 ;
  assign n35286 = n8690 & n35285 ;
  assign n35287 = ~n117 & n27422 ;
  assign n35288 = n35287 ^ n24547 ^ 1'b0 ;
  assign n35289 = n15191 & n32246 ;
  assign n35290 = n4968 & ~n35289 ;
  assign n35291 = n35290 ^ n18624 ^ 1'b0 ;
  assign n35292 = n29882 ^ n19908 ^ 1'b0 ;
  assign n35293 = n963 | n35292 ;
  assign n35294 = n25051 ^ n17100 ^ 1'b0 ;
  assign n35295 = n29150 & n35294 ;
  assign n35296 = n661 | n800 ;
  assign n35297 = n178 | n310 ;
  assign n35298 = n35297 ^ n6642 ^ 1'b0 ;
  assign n35299 = n2948 & n19712 ;
  assign n35300 = n35299 ^ n2545 ^ 1'b0 ;
  assign n35301 = n6695 & ~n35300 ;
  assign n35302 = n3423 & ~n6926 ;
  assign n35303 = n4845 & n35302 ;
  assign n35304 = n35303 ^ n2022 ^ 1'b0 ;
  assign n35305 = n7186 & n8789 ;
  assign n35306 = n1406 | n17961 ;
  assign n35307 = n35306 ^ n19091 ^ 1'b0 ;
  assign n35308 = ~n34347 & n35307 ;
  assign n35309 = n3512 & n24244 ;
  assign n35310 = ~n2506 & n35309 ;
  assign n35311 = ~n321 & n3506 ;
  assign n35312 = ~n12049 & n35311 ;
  assign n35313 = n2825 & n2987 ;
  assign n35314 = n35313 ^ n15200 ^ 1'b0 ;
  assign n35315 = n35314 ^ n7327 ^ 1'b0 ;
  assign n35316 = ~n12291 & n35315 ;
  assign n35317 = n14840 & ~n17259 ;
  assign n35318 = ~n35316 & n35317 ;
  assign n35319 = ~n1699 & n35318 ;
  assign n35320 = n35312 & n35319 ;
  assign n35321 = n2027 ^ n1502 ^ 1'b0 ;
  assign n35322 = n13564 | n35321 ;
  assign n35323 = n2888 ^ n1761 ^ 1'b0 ;
  assign n35324 = n2463 | n35323 ;
  assign n35325 = n8851 & n17627 ;
  assign n35326 = n4120 | n14938 ;
  assign n35327 = n35325 | n35326 ;
  assign n35328 = n1237 & n6587 ;
  assign n35329 = n7038 & n16969 ;
  assign n35330 = n17953 | n35329 ;
  assign n35331 = n26114 ^ n10390 ^ 1'b0 ;
  assign n35332 = n1426 & ~n35331 ;
  assign n35333 = n5609 & n9364 ;
  assign n35334 = n25551 | n31237 ;
  assign n35335 = n14083 & n35334 ;
  assign n35336 = n7236 ^ n6356 ^ n1300 ;
  assign n35337 = n9126 & ~n35336 ;
  assign n35338 = ~n32176 & n35337 ;
  assign n35339 = n23054 & ~n34230 ;
  assign n35340 = n35339 ^ n11648 ^ 1'b0 ;
  assign n35341 = ~n492 & n7688 ;
  assign n35342 = ~n2955 & n35341 ;
  assign n35343 = n18226 & ~n35342 ;
  assign n35344 = n35340 & n35343 ;
  assign n35345 = n345 | n8705 ;
  assign n35346 = n5501 | n35345 ;
  assign n35347 = n24640 & n35346 ;
  assign n35348 = n31181 | n31293 ;
  assign n35349 = n35348 ^ n26303 ^ 1'b0 ;
  assign n35350 = n35349 ^ n4021 ^ 1'b0 ;
  assign n35351 = n17647 & ~n31627 ;
  assign n35352 = n22598 | n27470 ;
  assign n35353 = n6826 & n33150 ;
  assign n35354 = ( ~n3681 & n4042 ) | ( ~n3681 & n16821 ) | ( n4042 & n16821 ) ;
  assign n35355 = ( ~n13993 & n23267 ) | ( ~n13993 & n35354 ) | ( n23267 & n35354 ) ;
  assign n35356 = n508 & n26513 ;
  assign n35357 = n35356 ^ n1078 ^ 1'b0 ;
  assign n35358 = n6822 ^ n685 ^ 1'b0 ;
  assign n35359 = n321 | n35358 ;
  assign n35360 = n19610 & n35359 ;
  assign n35361 = n10175 ^ n6488 ^ 1'b0 ;
  assign n35362 = n16835 & n35361 ;
  assign n35363 = ~n2353 & n35362 ;
  assign n35364 = ( ~n4437 & n12255 ) | ( ~n4437 & n23310 ) | ( n12255 & n23310 ) ;
  assign n35365 = n18711 | n18921 ;
  assign n35366 = n14987 ^ n9873 ^ 1'b0 ;
  assign n35367 = n2472 | n13132 ;
  assign n35368 = n35367 ^ n19906 ^ 1'b0 ;
  assign n35369 = n66 & ~n1742 ;
  assign n35370 = n35369 ^ n3791 ^ 1'b0 ;
  assign n35371 = n12388 & ~n35370 ;
  assign n35372 = n35371 ^ n4347 ^ 1'b0 ;
  assign n35373 = n9925 ^ n979 ^ 1'b0 ;
  assign n35374 = n24023 ^ n3221 ^ 1'b0 ;
  assign n35375 = n35373 & ~n35374 ;
  assign n35376 = n19588 ^ n12040 ^ n8234 ;
  assign n35377 = n2284 & n29437 ;
  assign n35378 = n5945 & ~n14164 ;
  assign n35379 = ~n30416 & n35378 ;
  assign n35380 = n35379 ^ n5642 ^ 1'b0 ;
  assign n35381 = n9263 ^ n3262 ^ 1'b0 ;
  assign n35382 = n19773 | n33392 ;
  assign n35383 = n23057 | n23771 ;
  assign n35384 = n35383 ^ n5394 ^ 1'b0 ;
  assign n35385 = n35384 ^ n4995 ^ 1'b0 ;
  assign n35386 = n15074 ^ n8375 ^ 1'b0 ;
  assign n35387 = n10543 & ~n35386 ;
  assign n35388 = n14624 ^ n9935 ^ 1'b0 ;
  assign n35389 = n532 & n35388 ;
  assign n35390 = n19825 ^ n6578 ^ 1'b0 ;
  assign n35391 = n9611 & ~n35390 ;
  assign n35392 = ~n14278 & n17508 ;
  assign n35393 = n35391 & ~n35392 ;
  assign n35394 = ~n542 & n7641 ;
  assign n35395 = n35394 ^ n27509 ^ 1'b0 ;
  assign n35396 = n16582 & ~n25872 ;
  assign n35397 = n32952 ^ n17473 ^ 1'b0 ;
  assign n35398 = ~n80 & n35397 ;
  assign n35399 = n29565 ^ n3152 ^ 1'b0 ;
  assign n35400 = n22619 | n35399 ;
  assign n35401 = n35400 ^ n495 ^ 1'b0 ;
  assign n35402 = n19660 ^ n3576 ^ 1'b0 ;
  assign n35403 = n24116 & n29508 ;
  assign n35404 = n6033 & ~n27623 ;
  assign n35405 = n30675 | n35404 ;
  assign n35406 = ~n11067 & n16301 ;
  assign n35407 = n5758 & n35406 ;
  assign n35408 = n17186 | n28266 ;
  assign n35409 = n32482 | n35408 ;
  assign n35412 = n5187 | n5882 ;
  assign n35413 = n1893 & n35412 ;
  assign n35410 = n114 & ~n14605 ;
  assign n35411 = n2644 & n35410 ;
  assign n35414 = n35413 ^ n35411 ^ 1'b0 ;
  assign n35415 = n24462 | n35414 ;
  assign n35416 = n1368 | n1692 ;
  assign n35417 = n35415 & ~n35416 ;
  assign n35418 = n653 & ~n19875 ;
  assign n35419 = n9901 & ~n35418 ;
  assign n35420 = n6846 & ~n35419 ;
  assign n35421 = n24500 ^ n11389 ^ 1'b0 ;
  assign n35422 = n2984 & ~n4611 ;
  assign n35423 = ~n2283 & n35422 ;
  assign n35424 = n35423 ^ n14998 ^ 1'b0 ;
  assign n35425 = ~n1525 & n3818 ;
  assign n35426 = n26733 & n35425 ;
  assign n35427 = n19131 ^ n10586 ^ 1'b0 ;
  assign n35428 = n32852 ^ n11931 ^ 1'b0 ;
  assign n35429 = n35427 & ~n35428 ;
  assign n35430 = ~n1077 & n35429 ;
  assign n35431 = n1303 & n35430 ;
  assign n35432 = n4866 | n35431 ;
  assign n35433 = n18858 ^ n2235 ^ 1'b0 ;
  assign n35434 = ~n5794 & n28122 ;
  assign n35435 = n1538 | n3719 ;
  assign n35436 = n3719 & ~n35435 ;
  assign n35437 = n35436 ^ n364 ^ 1'b0 ;
  assign n35438 = n3131 & ~n35437 ;
  assign n35439 = n35438 ^ n5780 ^ 1'b0 ;
  assign n35440 = n18719 ^ n184 ^ 1'b0 ;
  assign n35441 = n13694 & n35440 ;
  assign n35442 = n17323 & n20059 ;
  assign n35443 = ( n7102 & n17350 ) | ( n7102 & ~n35442 ) | ( n17350 & ~n35442 ) ;
  assign n35444 = n3033 | n3744 ;
  assign n35445 = n35444 ^ n5024 ^ 1'b0 ;
  assign n35446 = ~n35443 & n35445 ;
  assign n35447 = ~n11078 & n25863 ;
  assign n35448 = n32247 ^ n3670 ^ 1'b0 ;
  assign n35449 = ~n11573 & n35448 ;
  assign n35450 = n23605 ^ n18530 ^ 1'b0 ;
  assign n35451 = n9105 ^ n838 ^ 1'b0 ;
  assign n35452 = ~n325 & n3814 ;
  assign n35453 = ~n3814 & n35452 ;
  assign n35454 = n35453 ^ n27936 ^ 1'b0 ;
  assign n35455 = n29474 ^ n27066 ^ 1'b0 ;
  assign n35456 = n942 & n21033 ;
  assign n35457 = n35456 ^ n10507 ^ 1'b0 ;
  assign n35458 = ~n1891 & n35457 ;
  assign n35459 = n12539 | n28784 ;
  assign n35460 = n35459 ^ n12770 ^ 1'b0 ;
  assign n35461 = ~n1679 & n12125 ;
  assign n35462 = n2885 | n7179 ;
  assign n35463 = n35462 ^ n2220 ^ 1'b0 ;
  assign n35464 = n4449 | n35463 ;
  assign n35465 = n35461 | n35464 ;
  assign n35466 = ~n10009 & n13929 ;
  assign n35467 = ( ~n501 & n1629 ) | ( ~n501 & n14618 ) | ( n1629 & n14618 ) ;
  assign n35468 = n34123 | n35467 ;
  assign n35469 = n5846 | n35468 ;
  assign n35470 = n20487 & ~n27762 ;
  assign n35471 = ~n9038 & n9574 ;
  assign n35472 = n13324 | n35471 ;
  assign n35473 = ~n2067 & n22897 ;
  assign n35474 = n27461 ^ n27287 ^ 1'b0 ;
  assign n35475 = n24310 ^ n13137 ^ 1'b0 ;
  assign n35477 = n12948 & ~n30519 ;
  assign n35476 = n7181 | n7915 ;
  assign n35478 = n35477 ^ n35476 ^ 1'b0 ;
  assign n35479 = n28347 ^ n4193 ^ 1'b0 ;
  assign n35480 = n16345 | n20619 ;
  assign n35481 = n9688 ^ n832 ^ 1'b0 ;
  assign n35482 = n17632 ^ n2510 ^ 1'b0 ;
  assign n35483 = ~n35481 & n35482 ;
  assign n35484 = n30609 ^ n1152 ^ 1'b0 ;
  assign n35485 = n35483 & n35484 ;
  assign n35486 = n4023 | n5724 ;
  assign n35487 = ( n6810 & n13055 ) | ( n6810 & ~n35486 ) | ( n13055 & ~n35486 ) ;
  assign n35488 = n27530 & ~n35487 ;
  assign n35489 = n8220 & n35488 ;
  assign n35490 = n483 | n4516 ;
  assign n35491 = n11597 | n35490 ;
  assign n35492 = n35491 ^ n20094 ^ 1'b0 ;
  assign n35493 = n8551 & n35492 ;
  assign n35494 = n18069 ^ n253 ^ 1'b0 ;
  assign n35495 = n3939 & n13361 ;
  assign n35496 = n18975 | n35495 ;
  assign n35497 = ~n15652 & n17592 ;
  assign n35498 = n35496 & n35497 ;
  assign n35499 = n6764 ^ n4469 ^ 1'b0 ;
  assign n35500 = n32416 & ~n35499 ;
  assign n35501 = n20190 ^ n14838 ^ 1'b0 ;
  assign n35502 = n29585 ^ n16478 ^ 1'b0 ;
  assign n35503 = ~n8730 & n18808 ;
  assign n35504 = n20325 & n35503 ;
  assign n35505 = n35504 ^ n15617 ^ 1'b0 ;
  assign n35506 = n5402 & n17862 ;
  assign n35507 = n35506 ^ n7272 ^ 1'b0 ;
  assign n35508 = n12224 ^ n3258 ^ 1'b0 ;
  assign n35509 = n35507 & ~n35508 ;
  assign n35510 = n22991 ^ n6558 ^ 1'b0 ;
  assign n35511 = ( n605 & n11281 ) | ( n605 & ~n35510 ) | ( n11281 & ~n35510 ) ;
  assign n35512 = ~n7448 & n16020 ;
  assign n35513 = n10195 & ~n35512 ;
  assign n35514 = n35513 ^ n15911 ^ 1'b0 ;
  assign n35515 = n81 & n14217 ;
  assign n35516 = n35515 ^ n6094 ^ 1'b0 ;
  assign n35517 = n35516 ^ n24394 ^ n13590 ;
  assign n35518 = n21392 | n30506 ;
  assign n35519 = n2543 | n4166 ;
  assign n35520 = n6384 | n35519 ;
  assign n35521 = n35520 ^ n1546 ^ 1'b0 ;
  assign n35522 = n624 & n2744 ;
  assign n35523 = n35522 ^ n4823 ^ 1'b0 ;
  assign n35524 = n35523 ^ n16479 ^ 1'b0 ;
  assign n35525 = ( ~n6432 & n21083 ) | ( ~n6432 & n22647 ) | ( n21083 & n22647 ) ;
  assign n35526 = n8442 & ~n20580 ;
  assign n35527 = n17113 & n35526 ;
  assign n35528 = n4365 & ~n16362 ;
  assign n35529 = n35527 & n35528 ;
  assign n35530 = n19190 ^ n2344 ^ 1'b0 ;
  assign n35531 = n24387 ^ n21988 ^ 1'b0 ;
  assign n35533 = n7528 ^ n4629 ^ n1178 ;
  assign n35534 = ~n2933 & n35533 ;
  assign n35535 = n10691 & n35534 ;
  assign n35532 = n412 & n7031 ;
  assign n35536 = n35535 ^ n35532 ^ n707 ;
  assign n35537 = n35531 | n35536 ;
  assign n35541 = n9606 ^ n216 ^ 1'b0 ;
  assign n35542 = n7378 & n35541 ;
  assign n35538 = n6411 & ~n17833 ;
  assign n35539 = n35538 ^ n1390 ^ 1'b0 ;
  assign n35540 = n31805 & ~n35539 ;
  assign n35543 = n35542 ^ n35540 ^ 1'b0 ;
  assign n35544 = n2566 & ~n17055 ;
  assign n35545 = n7805 ^ n310 ^ 1'b0 ;
  assign n35546 = n11229 | n35545 ;
  assign n35547 = n9052 & ~n35546 ;
  assign n35548 = n35519 & n35547 ;
  assign n35549 = n35548 ^ n5015 ^ 1'b0 ;
  assign n35550 = n1840 ^ n102 ^ 1'b0 ;
  assign n35551 = n15617 ^ n14218 ^ 1'b0 ;
  assign n35552 = n5271 & n33898 ;
  assign n35553 = n18873 & n23379 ;
  assign n35554 = n34708 ^ n15577 ^ 1'b0 ;
  assign n35555 = n24912 ^ n12123 ^ 1'b0 ;
  assign n35556 = ~n16130 & n21075 ;
  assign n35560 = n12788 ^ n2003 ^ 1'b0 ;
  assign n35561 = n6194 & n35560 ;
  assign n35557 = n33716 ^ n3211 ^ 1'b0 ;
  assign n35558 = n79 | n35557 ;
  assign n35559 = n11003 | n35558 ;
  assign n35562 = n35561 ^ n35559 ^ n4903 ;
  assign n35563 = n3226 & ~n25943 ;
  assign n35564 = n26222 ^ n11755 ^ 1'b0 ;
  assign n35565 = n5513 | n35564 ;
  assign n35566 = ~n22348 & n35565 ;
  assign n35567 = n9099 ^ n833 ^ 1'b0 ;
  assign n35568 = n13493 & n35567 ;
  assign n35569 = n2288 & n11709 ;
  assign n35570 = ~n4122 & n24759 ;
  assign n35571 = n11641 | n18767 ;
  assign n35572 = n3830 | n29372 ;
  assign n35573 = n35571 & ~n35572 ;
  assign n35574 = n300 & ~n12303 ;
  assign n35575 = ~n2846 & n35574 ;
  assign n35576 = n2023 | n10481 ;
  assign n35577 = n1396 | n2553 ;
  assign n35578 = ~n13519 & n34686 ;
  assign n35579 = n29290 ^ n28253 ^ 1'b0 ;
  assign n35580 = n16292 & n20373 ;
  assign n35581 = n4898 | n5650 ;
  assign n35582 = n35581 ^ n18458 ^ 1'b0 ;
  assign n35583 = ~n2342 & n35582 ;
  assign n35584 = n6477 & n24172 ;
  assign n35585 = ~n5736 & n35584 ;
  assign n35586 = n2022 & ~n35585 ;
  assign n35587 = n2216 & ~n17460 ;
  assign n35588 = n35587 ^ n3162 ^ 1'b0 ;
  assign n35589 = ~n12857 & n25429 ;
  assign n35590 = n35589 ^ n856 ^ 1'b0 ;
  assign n35591 = n21961 ^ n6325 ^ 1'b0 ;
  assign n35592 = n9580 | n35591 ;
  assign n35593 = n23299 & ~n29585 ;
  assign n35594 = n19043 & ~n35593 ;
  assign n35595 = n4570 | n35594 ;
  assign n35596 = n35595 ^ n5310 ^ 1'b0 ;
  assign n35597 = n31403 ^ n14224 ^ 1'b0 ;
  assign n35598 = n4249 & n13102 ;
  assign n35599 = n27981 & ~n35598 ;
  assign n35600 = n654 & n35599 ;
  assign n35601 = ~n12649 & n14759 ;
  assign n35602 = n2209 & ~n7350 ;
  assign n35603 = n35602 ^ n1381 ^ 1'b0 ;
  assign n35604 = n3793 & ~n35603 ;
  assign n35609 = n294 & ~n2378 ;
  assign n35605 = n2477 & n5952 ;
  assign n35606 = n14114 & n35605 ;
  assign n35607 = n10889 | n35606 ;
  assign n35608 = n8106 & n35607 ;
  assign n35610 = n35609 ^ n35608 ^ 1'b0 ;
  assign n35611 = n34629 ^ n31362 ^ 1'b0 ;
  assign n35612 = n2659 | n10096 ;
  assign n35613 = n35611 & ~n35612 ;
  assign n35614 = n35613 ^ n7110 ^ 1'b0 ;
  assign n35615 = n24782 & n35614 ;
  assign n35616 = n5999 & n35615 ;
  assign n35617 = n35616 ^ n15313 ^ 1'b0 ;
  assign n35618 = n3122 | n15414 ;
  assign n35619 = n35618 ^ n6438 ^ 1'b0 ;
  assign n35620 = n9335 & n28123 ;
  assign n35621 = ~n35619 & n35620 ;
  assign n35622 = n8756 ^ n2142 ^ 1'b0 ;
  assign n35623 = n8158 & n35622 ;
  assign n35624 = ~n3509 & n35623 ;
  assign n35625 = ~n1994 & n35624 ;
  assign n35626 = n825 & n5271 ;
  assign n35627 = n5012 & n35626 ;
  assign n35628 = n30522 | n35627 ;
  assign n35629 = n25143 & ~n35628 ;
  assign n35631 = n26824 ^ n18736 ^ 1'b0 ;
  assign n35630 = n200 & n27985 ;
  assign n35632 = n35631 ^ n35630 ^ 1'b0 ;
  assign n35633 = n6785 ^ n2136 ^ 1'b0 ;
  assign n35634 = n18002 & ~n35633 ;
  assign n35635 = ~n2757 & n5124 ;
  assign n35636 = n35635 ^ n7818 ^ 1'b0 ;
  assign n35637 = n5458 & n35636 ;
  assign n35638 = ~n12432 & n35637 ;
  assign n35639 = n16355 & n26620 ;
  assign n35640 = n23698 ^ n11329 ^ 1'b0 ;
  assign n35641 = n2260 | n13813 ;
  assign n35642 = n35641 ^ n980 ^ 1'b0 ;
  assign n35643 = n3280 | n35642 ;
  assign n35644 = n292 | n23948 ;
  assign n35645 = n20135 ^ n5190 ^ 1'b0 ;
  assign n35646 = n4186 & n35645 ;
  assign n35647 = n35644 & ~n35646 ;
  assign n35648 = n14948 & n29159 ;
  assign n35649 = n35648 ^ n21140 ^ 1'b0 ;
  assign n35650 = n22668 & ~n33451 ;
  assign n35651 = ~n19377 & n35650 ;
  assign n35652 = ~n11796 & n33234 ;
  assign n35653 = n15907 ^ n2607 ^ 1'b0 ;
  assign n35654 = n35652 & n35653 ;
  assign n35655 = n1683 & n1867 ;
  assign n35656 = n6770 & ~n35655 ;
  assign n35657 = n2426 & n3196 ;
  assign n35658 = n17119 & n35657 ;
  assign n35659 = n35658 ^ n432 ^ 1'b0 ;
  assign n35660 = ~n2478 & n3037 ;
  assign n35661 = ( n210 & n495 ) | ( n210 & n1705 ) | ( n495 & n1705 ) ;
  assign n35662 = n9417 | n10926 ;
  assign n35663 = n35662 ^ n36 ^ 1'b0 ;
  assign n35664 = n35663 ^ n23843 ^ n19844 ;
  assign n35665 = ~n11117 & n26100 ;
  assign n35666 = n7607 & n29798 ;
  assign n35667 = n8870 | n11563 ;
  assign n35668 = n22993 ^ n4911 ^ 1'b0 ;
  assign n35669 = n1718 | n6074 ;
  assign n35670 = n16136 | n35669 ;
  assign n35671 = n9649 | n27683 ;
  assign n35672 = n13752 ^ n191 ^ 1'b0 ;
  assign n35673 = ( n10785 & n15588 ) | ( n10785 & ~n35672 ) | ( n15588 & ~n35672 ) ;
  assign n35674 = n29753 & ~n35673 ;
  assign n35675 = n35674 ^ n30687 ^ n20540 ;
  assign n35676 = n6114 | n7767 ;
  assign n35677 = n4951 ^ n1814 ^ 1'b0 ;
  assign n35678 = n35676 & n35677 ;
  assign n35679 = n9128 & n12073 ;
  assign n35680 = n16318 & n35679 ;
  assign n35681 = n2317 & ~n18308 ;
  assign n35682 = n35681 ^ n33243 ^ 1'b0 ;
  assign n35683 = n11784 ^ n9105 ^ 1'b0 ;
  assign n35684 = ~n233 & n35683 ;
  assign n35685 = n35684 ^ n18578 ^ 1'b0 ;
  assign n35686 = n3509 & ~n19068 ;
  assign n35687 = n5161 & n10005 ;
  assign n35688 = n31351 ^ n16307 ^ 1'b0 ;
  assign n35689 = ~n6633 & n10799 ;
  assign n35690 = ( n670 & ~n9703 ) | ( n670 & n35689 ) | ( ~n9703 & n35689 ) ;
  assign n35691 = n15582 & ~n35690 ;
  assign n35692 = ~n19330 & n24045 ;
  assign n35693 = n8011 ^ n3579 ^ 1'b0 ;
  assign n35694 = n10545 & ~n35693 ;
  assign n35695 = n8416 & ~n35694 ;
  assign n35696 = n1102 & ~n35695 ;
  assign n35697 = n34445 ^ n274 ^ 1'b0 ;
  assign n35698 = n7159 & n30492 ;
  assign n35699 = n35697 & n35698 ;
  assign n35700 = n11846 ^ n5914 ^ 1'b0 ;
  assign n35701 = n7203 & ~n35700 ;
  assign n35702 = n35701 ^ n13842 ^ n4840 ;
  assign n35703 = ~x0 & n13953 ;
  assign n35704 = ~n35702 & n35703 ;
  assign n35705 = ~n20547 & n29196 ;
  assign n35706 = n3589 ^ n1909 ^ 1'b0 ;
  assign n35707 = n1096 ^ n153 ^ 1'b0 ;
  assign n35708 = n35706 & n35707 ;
  assign n35709 = ~n4061 & n10277 ;
  assign n35710 = n20559 ^ n7040 ^ 1'b0 ;
  assign n35711 = n2697 & ~n35710 ;
  assign n35712 = n8081 | n29785 ;
  assign n35713 = n18033 ^ n4606 ^ 1'b0 ;
  assign n35714 = ~n1990 & n35713 ;
  assign n35715 = n2912 ^ n105 ^ 1'b0 ;
  assign n35716 = n5143 & n13660 ;
  assign n35717 = n10031 ^ n3820 ^ 1'b0 ;
  assign n35718 = n11803 | n11876 ;
  assign n35719 = n35718 ^ n23605 ^ 1'b0 ;
  assign n35720 = n6669 ^ n4419 ^ 1'b0 ;
  assign n35721 = n3988 & n35720 ;
  assign n35722 = n4491 & n35721 ;
  assign n35723 = n35075 ^ n16491 ^ 1'b0 ;
  assign n35724 = ~n29163 & n35723 ;
  assign n35726 = n6826 | n16413 ;
  assign n35727 = ~n24573 & n35726 ;
  assign n35725 = n25380 & n25529 ;
  assign n35728 = n35727 ^ n35725 ^ 1'b0 ;
  assign n35729 = n7607 & ~n10777 ;
  assign n35730 = n6150 | n35729 ;
  assign n35731 = n14946 ^ n4437 ^ 1'b0 ;
  assign n35732 = n20094 | n35731 ;
  assign n35733 = n35730 | n35732 ;
  assign n35734 = n1931 & ~n28194 ;
  assign n35735 = n9176 | n35734 ;
  assign n35736 = n7341 & n35735 ;
  assign n35737 = n35736 ^ n16803 ^ 1'b0 ;
  assign n35738 = n3843 | n5481 ;
  assign n35739 = n35738 ^ n10928 ^ 1'b0 ;
  assign n35740 = n35739 ^ n21379 ^ n6849 ;
  assign n35741 = ~n6159 & n10708 ;
  assign n35742 = n3431 & ~n10743 ;
  assign n35743 = n23108 ^ n7554 ^ 1'b0 ;
  assign n35744 = n4202 & n4332 ;
  assign n35745 = n8128 & ~n16528 ;
  assign n35746 = n10763 & ~n22551 ;
  assign n35747 = n35746 ^ n29231 ^ 1'b0 ;
  assign n35748 = n19715 & n24349 ;
  assign n35749 = n23337 ^ n556 ^ 1'b0 ;
  assign n35750 = n35749 ^ n1750 ^ 1'b0 ;
  assign n35751 = ~n2536 & n35750 ;
  assign n35752 = n11848 ^ n191 ^ 1'b0 ;
  assign n35753 = n18058 & ~n35752 ;
  assign n35754 = n1687 & n8896 ;
  assign n35755 = n35754 ^ n4324 ^ 1'b0 ;
  assign n35756 = n1511 & n1520 ;
  assign n35757 = n544 & ~n35756 ;
  assign n35758 = ~n35755 & n35757 ;
  assign n35759 = n7442 & n9012 ;
  assign n35760 = n35759 ^ n23633 ^ 1'b0 ;
  assign n35761 = n13376 ^ n592 ^ 1'b0 ;
  assign n35762 = n35761 ^ n11981 ^ 1'b0 ;
  assign n35763 = ~n28864 & n35762 ;
  assign n35764 = n30757 ^ n1065 ^ 1'b0 ;
  assign n35765 = n35763 & ~n35764 ;
  assign n35766 = ~n216 & n6084 ;
  assign n35767 = n2482 & ~n2947 ;
  assign n35768 = n35767 ^ n14080 ^ 1'b0 ;
  assign n35769 = n28526 & n35768 ;
  assign n35770 = n17743 & ~n35769 ;
  assign n35771 = ~n3924 & n30819 ;
  assign n35772 = n102 & n8042 ;
  assign n35773 = ~n1704 & n34312 ;
  assign n35774 = n13554 ^ n13167 ^ 1'b0 ;
  assign n35775 = n8551 ^ n7678 ^ 1'b0 ;
  assign n35776 = n14432 & ~n35775 ;
  assign n35777 = n26481 | n28063 ;
  assign n35778 = n11802 | n35777 ;
  assign n35779 = n8770 ^ n812 ^ 1'b0 ;
  assign n35780 = n2203 & ~n34490 ;
  assign n35781 = n6149 | n6742 ;
  assign n35782 = n35781 ^ n17841 ^ 1'b0 ;
  assign n35783 = n18856 & n35782 ;
  assign n35784 = n18548 | n27766 ;
  assign n35785 = n35784 ^ n32387 ^ 1'b0 ;
  assign n35786 = n2613 & ~n27522 ;
  assign n35787 = n16263 & ~n31358 ;
  assign n35788 = n5201 & n35787 ;
  assign n35789 = n8508 & n29960 ;
  assign n35790 = ~n4400 & n22967 ;
  assign n35791 = n3305 & n35790 ;
  assign n35792 = n35791 ^ n3707 ^ 1'b0 ;
  assign n35793 = n16893 & n35792 ;
  assign n35794 = n587 & ~n11529 ;
  assign n35795 = n2116 | n35794 ;
  assign n35796 = n9899 | n35795 ;
  assign n35797 = n35793 | n35796 ;
  assign n35798 = n32649 ^ n14694 ^ 1'b0 ;
  assign n35799 = n9164 ^ n2436 ^ 1'b0 ;
  assign n35800 = n35799 ^ n9935 ^ 1'b0 ;
  assign n35801 = n22916 ^ n2260 ^ 1'b0 ;
  assign n35802 = n12793 & n35801 ;
  assign n35803 = n4256 ^ n640 ^ 1'b0 ;
  assign n35804 = n20700 & ~n35803 ;
  assign n35805 = n9434 ^ n1959 ^ n1344 ;
  assign n35806 = ~n3133 & n35805 ;
  assign n35809 = n1164 | n15439 ;
  assign n35810 = n1164 & ~n35809 ;
  assign n35811 = n26287 | n35810 ;
  assign n35808 = ~n941 & n33400 ;
  assign n35812 = n35811 ^ n35808 ^ 1'b0 ;
  assign n35807 = n11120 & n33009 ;
  assign n35813 = n35812 ^ n35807 ^ 1'b0 ;
  assign n35814 = n4843 ^ n2514 ^ 1'b0 ;
  assign n35815 = n1617 | n2681 ;
  assign n35816 = n592 | n23392 ;
  assign n35817 = n35816 ^ n22239 ^ 1'b0 ;
  assign n35819 = n1690 & n2391 ;
  assign n35820 = ~n27798 & n35819 ;
  assign n35818 = n6950 | n29101 ;
  assign n35821 = n35820 ^ n35818 ^ 1'b0 ;
  assign n35822 = n6493 | n23589 ;
  assign n35823 = n17180 ^ n4775 ^ 1'b0 ;
  assign n35824 = n14731 ^ n4687 ^ 1'b0 ;
  assign n35825 = n35823 | n35824 ;
  assign n35826 = n15528 & n19411 ;
  assign n35827 = n20713 ^ n6236 ^ 1'b0 ;
  assign n35828 = n497 & n13841 ;
  assign n35829 = n35827 & n35828 ;
  assign n35830 = n16418 | n19830 ;
  assign n35831 = n159 & n15098 ;
  assign n35832 = n5046 & ~n35831 ;
  assign n35833 = ~n159 & n16422 ;
  assign n35834 = n35833 ^ n7007 ^ 1'b0 ;
  assign n35835 = n652 & n28881 ;
  assign n35836 = n11439 ^ n713 ^ n243 ;
  assign n35837 = n10061 ^ n5178 ^ 1'b0 ;
  assign n35838 = n1994 & ~n35837 ;
  assign n35839 = n24154 ^ n3692 ^ 1'b0 ;
  assign n35840 = n1975 & ~n35839 ;
  assign n35841 = n35838 & ~n35840 ;
  assign n35842 = n9662 ^ n133 ^ 1'b0 ;
  assign n35843 = ~n1900 & n35842 ;
  assign n35844 = ~n13947 & n28260 ;
  assign n35845 = ~n3739 & n15549 ;
  assign n35847 = n310 | n5823 ;
  assign n35848 = n35847 ^ n11915 ^ 1'b0 ;
  assign n35846 = n1622 | n16952 ;
  assign n35849 = n35848 ^ n35846 ^ 1'b0 ;
  assign n35850 = n419 | n616 ;
  assign n35851 = n34609 ^ n9765 ^ 1'b0 ;
  assign n35852 = n8894 | n35851 ;
  assign n35853 = n31837 ^ n5924 ^ 1'b0 ;
  assign n35854 = n14895 ^ n290 ^ 1'b0 ;
  assign n35855 = n25188 ^ n16413 ^ 1'b0 ;
  assign n35856 = n8568 | n20696 ;
  assign n35857 = n1463 & ~n35856 ;
  assign n35858 = n596 | n11187 ;
  assign n35859 = n4635 | n11095 ;
  assign n35861 = n1663 | n4441 ;
  assign n35862 = n31021 | n35861 ;
  assign n35860 = ~n3561 & n19400 ;
  assign n35863 = n35862 ^ n35860 ^ 1'b0 ;
  assign n35864 = n32299 ^ n18319 ^ 1'b0 ;
  assign n35865 = n2607 | n4422 ;
  assign n35866 = n20095 ^ n8079 ^ 1'b0 ;
  assign n35867 = n9580 ^ n1179 ^ 1'b0 ;
  assign n35868 = ~n2494 & n5074 ;
  assign n35869 = ~n9586 & n35868 ;
  assign n35870 = n24378 ^ n9523 ^ 1'b0 ;
  assign n35871 = n16962 & n35870 ;
  assign n35872 = n9619 & n13996 ;
  assign n35873 = n22309 & ~n35872 ;
  assign n35874 = n21399 ^ n17117 ^ 1'b0 ;
  assign n35875 = n35146 ^ n2060 ^ 1'b0 ;
  assign n35876 = n2414 & n35875 ;
  assign n35877 = ~n35874 & n35876 ;
  assign n35878 = n7301 & ~n26887 ;
  assign n35879 = n7247 & n8242 ;
  assign n35880 = n27573 ^ n21326 ^ 1'b0 ;
  assign n35881 = n35879 | n35880 ;
  assign n35883 = n7056 | n21424 ;
  assign n35882 = ~n499 & n29453 ;
  assign n35884 = n35883 ^ n35882 ^ 1'b0 ;
  assign n35885 = n1950 & n6371 ;
  assign n35886 = n3529 & n35885 ;
  assign n35887 = ~n10895 & n11112 ;
  assign n35888 = n35887 ^ n8980 ^ 1'b0 ;
  assign n35889 = n28512 ^ n3668 ^ 1'b0 ;
  assign n35890 = ~n10618 & n35889 ;
  assign n35891 = n8916 ^ n1456 ^ 1'b0 ;
  assign n35892 = n884 | n35891 ;
  assign n35893 = n3260 | n35892 ;
  assign n35894 = n35893 ^ n21167 ^ 1'b0 ;
  assign n35895 = n13864 | n29069 ;
  assign n35896 = n757 | n3088 ;
  assign n35897 = n35896 ^ n7310 ^ 1'b0 ;
  assign n35898 = n33273 ^ n11205 ^ n6566 ;
  assign n35899 = n11865 & n17879 ;
  assign n35900 = n13690 & ~n35899 ;
  assign n35901 = n954 | n9080 ;
  assign n35902 = n12217 | n31947 ;
  assign n35903 = n2073 | n22276 ;
  assign n35904 = n35902 & ~n35903 ;
  assign n35905 = n35904 ^ n15903 ^ 1'b0 ;
  assign n35906 = ~n8397 & n35905 ;
  assign n35907 = n17174 ^ n8102 ^ 1'b0 ;
  assign n35908 = n1304 & ~n16338 ;
  assign n35909 = n35908 ^ n4439 ^ 1'b0 ;
  assign n35910 = n26839 ^ n1495 ^ 1'b0 ;
  assign n35911 = n17008 & n20948 ;
  assign n35912 = n12044 & n35911 ;
  assign n35913 = n35910 & ~n35912 ;
  assign n35914 = n1928 & ~n18244 ;
  assign n35915 = n378 & n33392 ;
  assign n35916 = ~n9439 & n35915 ;
  assign n35917 = ( ~n174 & n513 ) | ( ~n174 & n4998 ) | ( n513 & n4998 ) ;
  assign n35918 = n10996 & n35917 ;
  assign n35919 = n35918 ^ n16441 ^ 1'b0 ;
  assign n35920 = n35919 ^ n18434 ^ n3413 ;
  assign n35921 = n35920 ^ n25876 ^ 1'b0 ;
  assign n35922 = n35921 ^ n169 ^ 1'b0 ;
  assign n35923 = n2842 ^ n200 ^ 1'b0 ;
  assign n35924 = ~n7383 & n17733 ;
  assign n35925 = n1838 & ~n35924 ;
  assign n35926 = n5013 & ~n12804 ;
  assign n35927 = n9702 | n21856 ;
  assign n35928 = n5427 & ~n35927 ;
  assign n35929 = n21795 ^ n14226 ^ 1'b0 ;
  assign n35930 = ~n29350 & n35929 ;
  assign n35931 = ( n9780 & n27384 ) | ( n9780 & ~n35930 ) | ( n27384 & ~n35930 ) ;
  assign n35932 = n35931 ^ n19041 ^ n12525 ;
  assign n35933 = n6950 ^ n384 ^ 1'b0 ;
  assign n35934 = n2562 & n35933 ;
  assign n35935 = n2362 | n4207 ;
  assign n35936 = n35934 | n35935 ;
  assign n35937 = ~n899 & n4925 ;
  assign n35938 = n10053 ^ n1552 ^ 1'b0 ;
  assign n35939 = ~n35937 & n35938 ;
  assign n35940 = n32600 ^ n13364 ^ 1'b0 ;
  assign n35941 = n19794 | n33406 ;
  assign n35942 = n4976 & ~n35941 ;
  assign n35943 = n5218 & ~n35942 ;
  assign n35944 = n10007 | n20377 ;
  assign n35945 = n35944 ^ n21509 ^ 1'b0 ;
  assign n35946 = n120 | n21043 ;
  assign n35947 = n35946 ^ n15468 ^ n10219 ;
  assign n35948 = ~n6695 & n8639 ;
  assign n35949 = n14984 ^ n2721 ^ 1'b0 ;
  assign n35950 = n853 | n4824 ;
  assign n35951 = n35950 ^ n13585 ^ 1'b0 ;
  assign n35952 = n27489 ^ n9894 ^ 1'b0 ;
  assign n35953 = ~n6863 & n17987 ;
  assign n35954 = ~n12469 & n35953 ;
  assign n35966 = ~n92 & n20921 ;
  assign n35967 = n878 & ~n35966 ;
  assign n35968 = n35966 & n35967 ;
  assign n35969 = n542 | n35968 ;
  assign n35970 = n35968 & ~n35969 ;
  assign n35971 = n1852 & n35970 ;
  assign n35955 = n928 & n7412 ;
  assign n35961 = n18692 & n30248 ;
  assign n35956 = n855 | n22513 ;
  assign n35957 = n22513 & ~n35956 ;
  assign n35958 = n952 & n35957 ;
  assign n35959 = n10461 & n35958 ;
  assign n35960 = n24788 | n35959 ;
  assign n35962 = n35961 ^ n35960 ^ 1'b0 ;
  assign n35963 = n23652 | n35962 ;
  assign n35964 = n35955 | n35963 ;
  assign n35965 = ~n27852 & n35964 ;
  assign n35972 = n35971 ^ n35965 ^ 1'b0 ;
  assign n35973 = n28308 ^ n1810 ^ 1'b0 ;
  assign n35974 = n8827 & ~n35973 ;
  assign n35975 = n9402 & n14195 ;
  assign n35976 = n13042 | n35975 ;
  assign n35977 = n9839 ^ n7767 ^ n6777 ;
  assign n35978 = n35275 ^ n13242 ^ 1'b0 ;
  assign n35979 = n1020 & n24343 ;
  assign n35980 = n35979 ^ n29426 ^ 1'b0 ;
  assign n35981 = n35978 & n35980 ;
  assign n35982 = n8418 & n26529 ;
  assign n35983 = n2910 & ~n16853 ;
  assign n35984 = n4321 & n5183 ;
  assign n35985 = n6567 & n35984 ;
  assign n35986 = n3960 & ~n35985 ;
  assign n35987 = n5205 | n12504 ;
  assign n35988 = n18555 | n35987 ;
  assign n35989 = n25260 ^ n12395 ^ 1'b0 ;
  assign n35990 = n11131 | n35989 ;
  assign n35991 = n35990 ^ n4742 ^ 1'b0 ;
  assign n35992 = n14838 & ~n23108 ;
  assign n35993 = n19575 | n35992 ;
  assign n35994 = n5393 & ~n9614 ;
  assign n35995 = ~n4556 & n35994 ;
  assign n35996 = n35995 ^ n14256 ^ 1'b0 ;
  assign n35997 = ~n7135 & n35996 ;
  assign n35998 = n776 & n15117 ;
  assign n35999 = ~n682 & n35998 ;
  assign n36000 = ~n3244 & n19370 ;
  assign n36001 = n21121 & n36000 ;
  assign n36002 = n18594 ^ n6041 ^ 1'b0 ;
  assign n36003 = ~n7614 & n36002 ;
  assign n36004 = n36003 ^ n190 ^ 1'b0 ;
  assign n36005 = n18657 | n36004 ;
  assign n36006 = n6666 & n17862 ;
  assign n36007 = n36006 ^ n6866 ^ 1'b0 ;
  assign n36008 = n36005 | n36007 ;
  assign n36009 = ~n1339 & n21875 ;
  assign n36010 = ~n5330 & n36009 ;
  assign n36011 = n36010 ^ n8891 ^ 1'b0 ;
  assign n36012 = ~n36008 & n36011 ;
  assign n36013 = n13701 ^ n11192 ^ 1'b0 ;
  assign n36014 = n6272 | n36013 ;
  assign n36015 = n35325 & ~n36014 ;
  assign n36016 = n2264 & n4485 ;
  assign n36017 = n36016 ^ n83 ^ 1'b0 ;
  assign n36018 = n8232 & n8524 ;
  assign n36019 = n36018 ^ n22254 ^ n6610 ;
  assign n36020 = n18195 & ~n22198 ;
  assign n36021 = n36020 ^ n5468 ^ 1'b0 ;
  assign n36022 = ~n7079 & n25952 ;
  assign n36023 = n36022 ^ n7745 ^ 1'b0 ;
  assign n36024 = n3500 & ~n7106 ;
  assign n36025 = n27073 & n36024 ;
  assign n36026 = n36025 ^ n8429 ^ 1'b0 ;
  assign n36027 = n36023 & ~n36026 ;
  assign n36028 = n9619 & ~n9983 ;
  assign n36029 = n32096 & n36028 ;
  assign n36030 = n22850 & n36029 ;
  assign n36031 = n3112 | n11203 ;
  assign n36032 = n21850 ^ n609 ^ 1'b0 ;
  assign n36033 = n1347 | n8693 ;
  assign n36034 = n36033 ^ n17901 ^ 1'b0 ;
  assign n36035 = n7596 | n36034 ;
  assign n36036 = n6764 | n26112 ;
  assign n36037 = n6165 ^ n683 ^ 1'b0 ;
  assign n36038 = n27206 | n36037 ;
  assign n36039 = ~n2933 & n31330 ;
  assign n36040 = n2820 & ~n3295 ;
  assign n36041 = n30154 | n34052 ;
  assign n36042 = ~n310 & n26761 ;
  assign n36043 = n1480 | n8856 ;
  assign n36044 = n36042 & ~n36043 ;
  assign n36045 = n5458 & n36044 ;
  assign n36046 = n8442 & n19000 ;
  assign n36047 = n36046 ^ n33977 ^ 1'b0 ;
  assign n36048 = n6878 & n15154 ;
  assign n36049 = n32778 ^ n25055 ^ 1'b0 ;
  assign n36050 = n3498 & n36049 ;
  assign n36051 = ( n15756 & ~n27198 ) | ( n15756 & n36050 ) | ( ~n27198 & n36050 ) ;
  assign n36052 = ~n21887 & n28430 ;
  assign n36053 = ~n35276 & n36052 ;
  assign n36054 = n6351 & n36053 ;
  assign n36055 = n14684 & ~n36054 ;
  assign n36056 = n2751 & n36055 ;
  assign n36057 = n11172 & ~n18741 ;
  assign n36058 = ~n1440 & n10174 ;
  assign n36059 = n11922 & n36058 ;
  assign n36060 = ( n78 & n2245 ) | ( n78 & n16342 ) | ( n2245 & n16342 ) ;
  assign n36061 = n21753 ^ n5533 ^ 1'b0 ;
  assign n36062 = n3416 | n36061 ;
  assign n36063 = n12046 | n17356 ;
  assign n36064 = n11521 | n36063 ;
  assign n36065 = n1927 & ~n5957 ;
  assign n36067 = n4650 ^ n2288 ^ 1'b0 ;
  assign n36068 = n4766 | n36067 ;
  assign n36066 = n21394 ^ n21199 ^ 1'b0 ;
  assign n36069 = n36068 ^ n36066 ^ 1'b0 ;
  assign n36070 = ~n3374 & n8028 ;
  assign n36071 = n10794 & n36070 ;
  assign n36072 = ~n17692 & n25868 ;
  assign n36073 = n13459 ^ n7491 ^ 1'b0 ;
  assign n36074 = ~n5050 & n36073 ;
  assign n36075 = n16916 & n21114 ;
  assign n36076 = n36075 ^ n24127 ^ 1'b0 ;
  assign n36077 = n36076 ^ n26350 ^ 1'b0 ;
  assign n36078 = n3535 & n10259 ;
  assign n36079 = n36078 ^ n470 ^ 1'b0 ;
  assign n36080 = n3221 & n3817 ;
  assign n36081 = ~n10751 & n36080 ;
  assign n36082 = n710 & ~n36081 ;
  assign n36083 = n20780 & n36082 ;
  assign n36084 = n36083 ^ n23860 ^ 1'b0 ;
  assign n36085 = n7040 & n19311 ;
  assign n36086 = n6922 ^ n4857 ^ 1'b0 ;
  assign n36087 = ~n36085 & n36086 ;
  assign n36088 = n26802 ^ n21298 ^ n11684 ;
  assign n36090 = n104 & ~n1138 ;
  assign n36091 = ~n9539 & n10433 ;
  assign n36092 = n36090 & ~n36091 ;
  assign n36093 = ~n8583 & n36092 ;
  assign n36089 = ~n2572 & n13354 ;
  assign n36094 = n36093 ^ n36089 ^ 1'b0 ;
  assign n36095 = n1350 & ~n15620 ;
  assign n36096 = n36095 ^ n11611 ^ n5466 ;
  assign n36097 = ~n14961 & n30896 ;
  assign n36098 = n26131 ^ n4661 ^ 1'b0 ;
  assign n36099 = n10484 | n36098 ;
  assign n36100 = n13782 & ~n15723 ;
  assign n36101 = n36100 ^ n18035 ^ 1'b0 ;
  assign n36102 = ~n14665 & n33900 ;
  assign n36103 = n24662 ^ n3032 ^ 1'b0 ;
  assign n36104 = n8599 ^ n8473 ^ n4183 ;
  assign n36105 = n5032 & n20347 ;
  assign n36106 = n4688 & n6664 ;
  assign n36107 = n1480 & n36106 ;
  assign n36108 = n33075 | n36107 ;
  assign n36109 = n36105 | n36108 ;
  assign n36110 = n16580 ^ n8568 ^ 1'b0 ;
  assign n36111 = n30131 ^ n12496 ^ 1'b0 ;
  assign n36112 = n36110 & ~n36111 ;
  assign n36113 = n7193 ^ n3524 ^ 1'b0 ;
  assign n36114 = n4568 & ~n36113 ;
  assign n36115 = n14495 & ~n35645 ;
  assign n36125 = n14932 ^ n4493 ^ 1'b0 ;
  assign n36116 = n3415 ^ n2136 ^ 1'b0 ;
  assign n36117 = n5836 | n36116 ;
  assign n36118 = n18110 | n36117 ;
  assign n36119 = n36118 ^ n21078 ^ 1'b0 ;
  assign n36120 = n19228 ^ n11201 ^ 1'b0 ;
  assign n36121 = n2317 & ~n36120 ;
  assign n36122 = n36121 ^ n2849 ^ 1'b0 ;
  assign n36123 = ~n3609 & n36122 ;
  assign n36124 = ~n36119 & n36123 ;
  assign n36126 = n36125 ^ n36124 ^ 1'b0 ;
  assign n36127 = ~n16049 & n36126 ;
  assign n36128 = n6646 ^ n2352 ^ 1'b0 ;
  assign n36129 = ~n34719 & n36128 ;
  assign n36130 = n8977 ^ n4268 ^ 1'b0 ;
  assign n36131 = n16143 ^ n3871 ^ 1'b0 ;
  assign n36132 = n36130 & ~n36131 ;
  assign n36133 = n36129 & ~n36132 ;
  assign n36134 = n14678 & ~n27004 ;
  assign n36135 = ( ~n16259 & n26142 ) | ( ~n16259 & n36134 ) | ( n26142 & n36134 ) ;
  assign n36136 = n4348 & ~n31459 ;
  assign n36137 = n21498 ^ n19876 ^ 1'b0 ;
  assign n36138 = ~n4360 & n21997 ;
  assign n36139 = ~n3762 & n36138 ;
  assign n36140 = n5559 ^ n2914 ^ 1'b0 ;
  assign n36141 = ~n36139 & n36140 ;
  assign n36142 = n17207 ^ n7429 ^ 1'b0 ;
  assign n36143 = n1135 & ~n6514 ;
  assign n36144 = n36142 & n36143 ;
  assign n36145 = n4097 & n26802 ;
  assign n36146 = n36145 ^ n13891 ^ 1'b0 ;
  assign n36147 = ~n1933 & n7678 ;
  assign n36148 = n3546 | n31936 ;
  assign n36149 = n36148 ^ n6197 ^ 1'b0 ;
  assign n36150 = n9752 & ~n18943 ;
  assign n36151 = n29613 | n36150 ;
  assign n36152 = ( n8319 & n14802 ) | ( n8319 & ~n30875 ) | ( n14802 & ~n30875 ) ;
  assign n36153 = n25027 ^ n5663 ^ 1'b0 ;
  assign n36154 = n19109 | n36153 ;
  assign n36155 = n36152 | n36154 ;
  assign n36171 = n89 & ~n255 ;
  assign n36172 = n12620 & n36171 ;
  assign n36173 = n223 & ~n36172 ;
  assign n36174 = ~n223 & n36173 ;
  assign n36175 = n17083 | n36174 ;
  assign n36176 = n17083 & ~n36175 ;
  assign n36156 = n1345 & ~n2517 ;
  assign n36157 = n18902 & n36156 ;
  assign n36158 = ~n18095 & n36157 ;
  assign n36159 = n1191 & ~n15935 ;
  assign n36160 = n512 & ~n28456 ;
  assign n36161 = n28456 & n36160 ;
  assign n36162 = n32 | n36161 ;
  assign n36163 = n36161 & ~n36162 ;
  assign n36164 = n638 & n942 ;
  assign n36165 = ~n638 & n36164 ;
  assign n36166 = n276 & n36165 ;
  assign n36167 = n36163 & ~n36166 ;
  assign n36168 = ~n36159 & n36167 ;
  assign n36169 = n36158 & n36168 ;
  assign n36170 = n36169 ^ n15387 ^ 1'b0 ;
  assign n36177 = n36176 ^ n36170 ^ 1'b0 ;
  assign n36178 = n7247 & n7915 ;
  assign n36179 = n36178 ^ n2364 ^ 1'b0 ;
  assign n36180 = n5831 | n36179 ;
  assign n36181 = n36180 ^ n6332 ^ 1'b0 ;
  assign n36182 = n36181 ^ n11961 ^ 1'b0 ;
  assign n36183 = n36177 & n36182 ;
  assign n36184 = n28062 ^ n10607 ^ 1'b0 ;
  assign n36185 = n13125 | n19922 ;
  assign n36186 = n4851 & ~n16979 ;
  assign n36187 = n11533 & n36186 ;
  assign n36188 = n9931 ^ n6808 ^ 1'b0 ;
  assign n36189 = ~n36187 & n36188 ;
  assign n36190 = n34643 & n36189 ;
  assign n36191 = n284 & n4818 ;
  assign n36192 = ~n2774 & n36191 ;
  assign n36193 = ~n32389 & n36192 ;
  assign n36194 = n10347 ^ n5747 ^ 1'b0 ;
  assign n36195 = n33695 & n36194 ;
  assign n36196 = n34207 ^ n3050 ^ 1'b0 ;
  assign n36197 = n6703 ^ n5846 ^ 1'b0 ;
  assign n36198 = ~n33960 & n36197 ;
  assign n36199 = n32092 & ~n35372 ;
  assign n36200 = n22978 ^ n18298 ^ n9343 ;
  assign n36201 = n2610 & ~n8976 ;
  assign n36202 = n36201 ^ n2910 ^ 1'b0 ;
  assign n36203 = ~n6349 & n20828 ;
  assign n36204 = ~n36202 & n36203 ;
  assign n36205 = n5863 & n16862 ;
  assign n36206 = ~n2722 & n14734 ;
  assign n36207 = ~n2789 & n16321 ;
  assign n36208 = ~n33422 & n36207 ;
  assign n36209 = n8091 | n15585 ;
  assign n36210 = ( n2212 & n3535 ) | ( n2212 & n30639 ) | ( n3535 & n30639 ) ;
  assign n36211 = ~n2260 & n10512 ;
  assign n36212 = ~n501 & n36211 ;
  assign n36213 = ~n20201 & n34650 ;
  assign n36214 = n18214 ^ n6493 ^ 1'b0 ;
  assign n36215 = n7096 & n36214 ;
  assign n36216 = n4645 ^ n4041 ^ 1'b0 ;
  assign n36217 = n22621 ^ n83 ^ 1'b0 ;
  assign n36218 = n36216 & ~n36217 ;
  assign n36219 = n36218 ^ n25197 ^ 1'b0 ;
  assign n36220 = n7973 ^ n4448 ^ 1'b0 ;
  assign n36221 = ~n12407 & n36220 ;
  assign n36222 = n36221 ^ n21351 ^ 1'b0 ;
  assign n36223 = ~n7132 & n36222 ;
  assign n36224 = n7913 ^ n775 ^ 1'b0 ;
  assign n36225 = n36224 ^ n2785 ^ 1'b0 ;
  assign n36226 = ~n135 & n4798 ;
  assign n36227 = n36226 ^ n28379 ^ 1'b0 ;
  assign n36228 = ~n793 & n26813 ;
  assign n36229 = ~n28793 & n36228 ;
  assign n36230 = n582 & ~n7825 ;
  assign n36231 = n36229 & n36230 ;
  assign n36232 = n36231 ^ n582 ^ 1'b0 ;
  assign n36233 = n10584 ^ n246 ^ 1'b0 ;
  assign n36234 = n36232 & n36233 ;
  assign n36235 = n4504 ^ n1243 ^ 1'b0 ;
  assign n36236 = n16417 & n36235 ;
  assign n36237 = n879 & n6588 ;
  assign n36238 = ~n10909 & n36237 ;
  assign n36239 = n27943 & ~n36238 ;
  assign n36240 = n24701 | n36239 ;
  assign n36241 = n13726 ^ n2642 ^ n758 ;
  assign n36242 = n20723 ^ n1096 ^ n300 ;
  assign n36243 = n36242 ^ n20086 ^ 1'b0 ;
  assign n36244 = ~n1326 & n20487 ;
  assign n36245 = n6551 & ~n23619 ;
  assign n36246 = n11777 & ~n33353 ;
  assign n36247 = n36246 ^ n2148 ^ 1'b0 ;
  assign n36248 = n7376 | n12504 ;
  assign n36249 = n14476 & n36248 ;
  assign n36250 = n27501 ^ n11833 ^ 1'b0 ;
  assign n36251 = ~n36249 & n36250 ;
  assign n36252 = n36251 ^ n10145 ^ 1'b0 ;
  assign n36253 = n28881 ^ n23001 ^ 1'b0 ;
  assign n36254 = n8319 ^ n6357 ^ 1'b0 ;
  assign n36255 = n3356 & n3477 ;
  assign n36256 = n403 & n9414 ;
  assign n36257 = n3570 | n36256 ;
  assign n36258 = n10544 | n12457 ;
  assign n36259 = n20872 & ~n26972 ;
  assign n36260 = n20531 ^ n748 ^ 1'b0 ;
  assign n36261 = n36259 & ~n36260 ;
  assign n36262 = n10293 | n10653 ;
  assign n36263 = n22998 & ~n36262 ;
  assign n36264 = n8283 & ~n22496 ;
  assign n36265 = n17112 & n27228 ;
  assign n36266 = n36265 ^ n2431 ^ 1'b0 ;
  assign n36267 = n33884 ^ n9036 ^ 1'b0 ;
  assign n36268 = n8342 & n36267 ;
  assign n36269 = n36268 ^ n15775 ^ 1'b0 ;
  assign n36270 = n3595 | n15965 ;
  assign n36271 = n11079 ^ n2302 ^ 1'b0 ;
  assign n36272 = n10831 & n36271 ;
  assign n36273 = n336 & ~n36272 ;
  assign n36274 = n20750 & n27192 ;
  assign n36275 = n22213 ^ n18205 ^ 1'b0 ;
  assign n36276 = ~n3283 & n36275 ;
  assign n36280 = n5463 & ~n11197 ;
  assign n36277 = n2420 | n6100 ;
  assign n36278 = n36277 ^ n11923 ^ 1'b0 ;
  assign n36279 = n709 & n36278 ;
  assign n36281 = n36280 ^ n36279 ^ 1'b0 ;
  assign n36282 = ~n2362 & n7627 ;
  assign n36283 = n36282 ^ n9082 ^ 1'b0 ;
  assign n36284 = n6880 & n36283 ;
  assign n36285 = n30196 | n31746 ;
  assign n36286 = n36285 ^ n3640 ^ 1'b0 ;
  assign n36287 = n36286 ^ n456 ^ 1'b0 ;
  assign n36288 = n142 & ~n15329 ;
  assign n36290 = n8897 | n12501 ;
  assign n36291 = n5538 & ~n36290 ;
  assign n36289 = n1000 & n5880 ;
  assign n36292 = n36291 ^ n36289 ^ 1'b0 ;
  assign n36293 = n10133 & ~n18016 ;
  assign n36294 = n1880 & n12454 ;
  assign n36295 = n36294 ^ n4139 ^ 1'b0 ;
  assign n36296 = n18207 & n25348 ;
  assign n36297 = n1785 & ~n36296 ;
  assign n36298 = n12280 | n36297 ;
  assign n36299 = ~n8393 & n25118 ;
  assign n36300 = n36298 & n36299 ;
  assign n36301 = n14532 ^ n2456 ^ 1'b0 ;
  assign n36302 = n10420 & n36301 ;
  assign n36303 = n6622 & ~n36302 ;
  assign n36304 = n7497 & n35461 ;
  assign n36305 = n36304 ^ n11934 ^ 1'b0 ;
  assign n36306 = n31432 ^ n2431 ^ 1'b0 ;
  assign n36307 = ~n8967 & n16972 ;
  assign n36308 = ~n10682 & n36307 ;
  assign n36309 = n30528 ^ n29685 ^ 1'b0 ;
  assign n36310 = ~n4904 & n8442 ;
  assign n36311 = n35603 ^ n9848 ^ 1'b0 ;
  assign n36312 = n21199 ^ n13080 ^ 1'b0 ;
  assign n36313 = n568 & n18384 ;
  assign n36314 = n13683 ^ n10343 ^ 1'b0 ;
  assign n36315 = n19788 | n36314 ;
  assign n36316 = n18715 & n21565 ;
  assign n36317 = ~n390 & n1704 ;
  assign n36318 = ~n3214 & n36317 ;
  assign n36319 = ~n1113 & n2399 ;
  assign n36320 = n36319 ^ n16577 ^ 1'b0 ;
  assign n36321 = n465 | n9933 ;
  assign n36322 = ~n21242 & n36321 ;
  assign n36323 = ~n17934 & n36322 ;
  assign n36324 = n10923 ^ n3919 ^ 1'b0 ;
  assign n36325 = n14659 & ~n16558 ;
  assign n36326 = ~n36324 & n36325 ;
  assign n36327 = n16491 & ~n23945 ;
  assign n36328 = n36327 ^ n25052 ^ n2235 ;
  assign n36329 = n1878 & ~n5914 ;
  assign n36330 = n32138 & n36329 ;
  assign n36331 = n18564 & n22450 ;
  assign n36332 = n18647 & n36331 ;
  assign n36333 = n36332 ^ n5971 ^ 1'b0 ;
  assign n36334 = n987 | n15042 ;
  assign n36335 = n36334 ^ n8889 ^ 1'b0 ;
  assign n36336 = n1790 & ~n24831 ;
  assign n36337 = n24970 ^ n3427 ^ 1'b0 ;
  assign n36338 = n33816 ^ n29860 ^ 1'b0 ;
  assign n36339 = n34538 ^ n7952 ^ 1'b0 ;
  assign n36340 = ~n5190 & n13842 ;
  assign n36341 = n36340 ^ n9636 ^ 1'b0 ;
  assign n36342 = n7523 & n26234 ;
  assign n36343 = n27489 ^ n13695 ^ 1'b0 ;
  assign n36344 = n9501 | n22124 ;
  assign n36345 = n36344 ^ n29109 ^ 1'b0 ;
  assign n36346 = n8401 & ~n34431 ;
  assign n36347 = n11083 & n36346 ;
  assign n36348 = ~n5744 & n26331 ;
  assign n36349 = n6196 & n36348 ;
  assign n36350 = n3382 & ~n36349 ;
  assign n36351 = n7690 & ~n11777 ;
  assign n36352 = ( n722 & n31778 ) | ( n722 & ~n36351 ) | ( n31778 & ~n36351 ) ;
  assign n36353 = n31505 ^ n30794 ^ 1'b0 ;
  assign n36354 = n4563 ^ n2843 ^ 1'b0 ;
  assign n36355 = n1437 | n36354 ;
  assign n36356 = n36355 ^ n3354 ^ 1'b0 ;
  assign n36357 = n18953 ^ n1435 ^ 1'b0 ;
  assign n36358 = n10420 & n32276 ;
  assign n36359 = n23910 ^ n1981 ^ 1'b0 ;
  assign n36361 = n19584 ^ n3346 ^ 1'b0 ;
  assign n36362 = n86 & ~n36361 ;
  assign n36360 = n38 & ~n8632 ;
  assign n36363 = n36362 ^ n36360 ^ 1'b0 ;
  assign n36364 = ( n1210 & n1469 ) | ( n1210 & n14587 ) | ( n1469 & n14587 ) ;
  assign n36365 = n15790 & n26791 ;
  assign n36366 = n32487 & n36365 ;
  assign n36367 = n2326 | n8643 ;
  assign n36368 = n34251 | n36367 ;
  assign n36369 = n6922 ^ n4591 ^ 1'b0 ;
  assign n36370 = n37 | n36369 ;
  assign n36371 = n1887 & ~n36370 ;
  assign n36372 = n36371 ^ n21136 ^ 1'b0 ;
  assign n36373 = n177 & ~n36372 ;
  assign n36374 = n11350 & ~n32690 ;
  assign n36375 = n20426 & ~n36187 ;
  assign n36376 = n22085 ^ n7860 ^ 1'b0 ;
  assign n36377 = n294 & n7395 ;
  assign n36378 = ~n27565 & n36377 ;
  assign n36379 = n7214 | n28879 ;
  assign n36380 = ~n3719 & n28198 ;
  assign n36381 = n1759 & ~n8990 ;
  assign n36382 = n17339 & n36381 ;
  assign n36383 = ~n10020 & n36068 ;
  assign n36384 = n34980 ^ n34854 ^ 1'b0 ;
  assign n36385 = n1040 & ~n36384 ;
  assign n36386 = ~n5205 & n14157 ;
  assign n36387 = n6376 & n23882 ;
  assign n36388 = n13682 & n36387 ;
  assign n36389 = n36388 ^ n33930 ^ 1'b0 ;
  assign n36390 = n2898 | n7424 ;
  assign n36391 = n14109 | n36390 ;
  assign n36392 = n4466 | n11573 ;
  assign n36393 = n4635 ^ n1444 ^ 1'b0 ;
  assign n36394 = n3523 | n36393 ;
  assign n36395 = n21683 | n36394 ;
  assign n36396 = n17096 & ~n36395 ;
  assign n36397 = n14383 | n32881 ;
  assign n36398 = n20929 ^ n5684 ^ 1'b0 ;
  assign n36399 = n3527 | n36398 ;
  assign n36400 = n16072 & ~n36399 ;
  assign n36401 = ~n8289 & n9227 ;
  assign n36402 = n36401 ^ n7870 ^ 1'b0 ;
  assign n36403 = n36402 ^ n14976 ^ 1'b0 ;
  assign n36404 = n36400 | n36403 ;
  assign n36405 = n34668 | n35109 ;
  assign n36406 = n36404 & ~n36405 ;
  assign n36407 = ~n76 & n5914 ;
  assign n36408 = n15305 & ~n36407 ;
  assign n36409 = n4202 & ~n20364 ;
  assign n36410 = n5823 & n9781 ;
  assign n36411 = n21136 ^ n8422 ^ 1'b0 ;
  assign n36412 = n13068 | n36411 ;
  assign n36413 = n9592 ^ n1443 ^ 1'b0 ;
  assign n36414 = n15770 & ~n36413 ;
  assign n36415 = n36412 | n36414 ;
  assign n36416 = ~n25790 & n33972 ;
  assign n36417 = ~n4093 & n36416 ;
  assign n36418 = n34146 & ~n36417 ;
  assign n36419 = n33084 ^ n18392 ^ 1'b0 ;
  assign n36420 = n8970 & n10747 ;
  assign n36421 = n23328 & n36420 ;
  assign n36422 = n20185 ^ n11266 ^ 1'b0 ;
  assign n36423 = ~n22213 & n29300 ;
  assign n36424 = n23397 ^ n15086 ^ 1'b0 ;
  assign n36425 = n21225 | n36424 ;
  assign n36426 = n6463 | n20695 ;
  assign n36427 = n12969 | n36426 ;
  assign n36428 = n36427 ^ n33638 ^ n1922 ;
  assign n36429 = n5761 & n14941 ;
  assign n36430 = n36429 ^ n26737 ^ 1'b0 ;
  assign n36431 = n17907 & ~n35276 ;
  assign n36432 = n36431 ^ n2856 ^ 1'b0 ;
  assign n36433 = ~n624 & n6444 ;
  assign n36434 = n8056 ^ n4299 ^ 1'b0 ;
  assign n36435 = n1851 | n36434 ;
  assign n36436 = n158 | n6174 ;
  assign n36437 = n1227 & ~n36436 ;
  assign n36438 = n36437 ^ n10617 ^ 1'b0 ;
  assign n36439 = n14469 & ~n36438 ;
  assign n36440 = n36439 ^ n12114 ^ 1'b0 ;
  assign n36441 = n27434 ^ n24343 ^ 1'b0 ;
  assign n36442 = n2542 ^ n1214 ^ 1'b0 ;
  assign n36443 = n36442 ^ n24869 ^ 1'b0 ;
  assign n36444 = n9299 & n36443 ;
  assign n36446 = n12661 ^ n193 ^ 1'b0 ;
  assign n36445 = n1591 & ~n13868 ;
  assign n36447 = n36446 ^ n36445 ^ 1'b0 ;
  assign n36448 = n998 & n1031 ;
  assign n36449 = n36448 ^ n7920 ^ 1'b0 ;
  assign n36450 = ~n26264 & n36449 ;
  assign n36451 = n14209 | n15283 ;
  assign n36452 = n24651 ^ n497 ^ 1'b0 ;
  assign n36453 = n8408 & ~n36452 ;
  assign n36454 = n18976 ^ n9911 ^ 1'b0 ;
  assign n36455 = n1523 & n36454 ;
  assign n36456 = n6834 & n36455 ;
  assign n36457 = n164 | n9775 ;
  assign n36458 = n5050 & n8563 ;
  assign n36459 = n6731 ^ n1849 ^ 1'b0 ;
  assign n36460 = ~n2593 & n36066 ;
  assign n36461 = n8268 & n13529 ;
  assign n36462 = ~n29175 & n36461 ;
  assign n36463 = n25075 & n29035 ;
  assign n36464 = n36463 ^ n1437 ^ 1'b0 ;
  assign n36465 = n31108 & n36464 ;
  assign n36466 = n5148 ^ n758 ^ 1'b0 ;
  assign n36467 = n28345 ^ n17502 ^ n339 ;
  assign n36473 = ~n212 & n10987 ;
  assign n36468 = n5045 ^ n255 ^ 1'b0 ;
  assign n36469 = n7815 | n36468 ;
  assign n36470 = n36469 ^ n9539 ^ 1'b0 ;
  assign n36471 = n15521 & n36470 ;
  assign n36472 = ~n2497 & n36471 ;
  assign n36474 = n36473 ^ n36472 ^ 1'b0 ;
  assign n36475 = n27648 ^ n19413 ^ 1'b0 ;
  assign n36476 = n25655 | n31428 ;
  assign n36477 = n1677 ^ n1087 ^ 1'b0 ;
  assign n36478 = n36477 ^ n4963 ^ 1'b0 ;
  assign n36479 = n3882 & ~n8024 ;
  assign n36480 = n36479 ^ n17003 ^ 1'b0 ;
  assign n36481 = n36480 ^ n4933 ^ 1'b0 ;
  assign n36482 = n10459 & ~n15448 ;
  assign n36483 = n29180 & n36482 ;
  assign n36484 = n19854 | n24689 ;
  assign n36485 = n1604 ^ n210 ^ 1'b0 ;
  assign n36486 = n32349 & ~n36485 ;
  assign n36487 = n1845 | n20058 ;
  assign n36488 = n36486 | n36487 ;
  assign n36491 = n17684 ^ n3226 ^ 1'b0 ;
  assign n36492 = n22122 & n36491 ;
  assign n36489 = n21942 & ~n30956 ;
  assign n36490 = n36489 ^ n21793 ^ 1'b0 ;
  assign n36493 = n36492 ^ n36490 ^ 1'b0 ;
  assign n36494 = n19390 & ~n27151 ;
  assign n36495 = n7902 & n36098 ;
  assign n36496 = n36495 ^ n18927 ^ 1'b0 ;
  assign n36497 = ~n2943 & n22890 ;
  assign n36498 = n11130 & ~n16173 ;
  assign n36499 = n1050 | n11680 ;
  assign n36500 = n36499 ^ n2552 ^ 1'b0 ;
  assign n36501 = n36500 ^ n34041 ^ 1'b0 ;
  assign n36502 = n4334 & ~n13275 ;
  assign n36503 = n36502 ^ n13003 ^ 1'b0 ;
  assign n36504 = n229 & n35917 ;
  assign n36505 = n36503 & n36504 ;
  assign n36506 = n15769 ^ n10587 ^ 1'b0 ;
  assign n36507 = n16677 ^ n4706 ^ 1'b0 ;
  assign n36508 = n15775 ^ n13341 ^ 1'b0 ;
  assign n36509 = n36507 | n36508 ;
  assign n36510 = n16724 | n36509 ;
  assign n36511 = n741 | n36510 ;
  assign n36512 = n670 & ~n8518 ;
  assign n36513 = n36512 ^ n12737 ^ 1'b0 ;
  assign n36514 = n28011 & ~n36513 ;
  assign n36515 = n36514 ^ n36509 ^ 1'b0 ;
  assign n36516 = n2774 ^ n1396 ^ 1'b0 ;
  assign n36517 = ~n4853 & n36516 ;
  assign n36518 = ~n10265 & n26027 ;
  assign n36519 = n6651 & n36518 ;
  assign n36520 = n3433 ^ n148 ^ 1'b0 ;
  assign n36521 = n25271 & n36520 ;
  assign n36522 = n36521 ^ n16395 ^ n14748 ;
  assign n36523 = n12109 & ~n17616 ;
  assign n36524 = n12801 & n13611 ;
  assign n36525 = n17560 & ~n25025 ;
  assign n36526 = n36525 ^ n1109 ^ 1'b0 ;
  assign n36528 = n5755 | n11044 ;
  assign n36529 = n8590 | n36528 ;
  assign n36527 = ~n18026 & n19236 ;
  assign n36530 = n36529 ^ n36527 ^ 1'b0 ;
  assign n36531 = ~n158 & n36530 ;
  assign n36532 = n964 | n15066 ;
  assign n36533 = n9136 & ~n36532 ;
  assign n36534 = n2034 ^ n612 ^ 1'b0 ;
  assign n36535 = n30606 ^ n1658 ^ 1'b0 ;
  assign n36536 = n16070 & ~n36535 ;
  assign n36537 = ( n4415 & n12519 ) | ( n4415 & ~n35955 ) | ( n12519 & ~n35955 ) ;
  assign n36538 = n12664 | n28751 ;
  assign n36539 = n1368 | n36538 ;
  assign n36540 = n8129 & n29780 ;
  assign n36541 = n6226 & n36540 ;
  assign n36542 = n36541 ^ n177 ^ 1'b0 ;
  assign n36544 = n4430 ^ n2687 ^ 1'b0 ;
  assign n36545 = n669 | n21778 ;
  assign n36546 = n36544 & ~n36545 ;
  assign n36543 = n1880 & ~n21651 ;
  assign n36547 = n36546 ^ n36543 ^ 1'b0 ;
  assign n36548 = ~n1662 & n36268 ;
  assign n36549 = n14401 & n36548 ;
  assign n36550 = n36549 ^ n35350 ^ 1'b0 ;
  assign n36551 = n21476 & n36550 ;
  assign n36552 = ~n2642 & n13585 ;
  assign n36553 = n36552 ^ n16925 ^ 1'b0 ;
  assign n36554 = n3440 | n36553 ;
  assign n36555 = n17490 ^ n3875 ^ 1'b0 ;
  assign n36556 = n11003 ^ n851 ^ 1'b0 ;
  assign n36557 = n21683 ^ n9845 ^ 1'b0 ;
  assign n36558 = n9085 ^ n5537 ^ 1'b0 ;
  assign n36559 = ~n2833 & n36558 ;
  assign n36560 = n2862 & ~n25839 ;
  assign n36561 = n26499 & n36560 ;
  assign n36562 = n24833 | n36561 ;
  assign n36564 = n5024 ^ n23 ^ 1'b0 ;
  assign n36563 = n247 & n26363 ;
  assign n36565 = n36564 ^ n36563 ^ 1'b0 ;
  assign n36566 = n36565 ^ n3247 ^ 1'b0 ;
  assign n36567 = n30914 ^ n13930 ^ 1'b0 ;
  assign n36568 = n11874 ^ n2484 ^ 1'b0 ;
  assign n36569 = n713 & n23119 ;
  assign n36570 = ~n5406 & n33278 ;
  assign n36571 = n36570 ^ n18223 ^ 1'b0 ;
  assign n36572 = ~n10156 & n13588 ;
  assign n36573 = ~n19466 & n36572 ;
  assign n36574 = n5661 & n36573 ;
  assign n36575 = n7109 & ~n19217 ;
  assign n36576 = ~n5070 & n8571 ;
  assign n36577 = ~n10517 & n36576 ;
  assign n36578 = n7673 ^ n6544 ^ 1'b0 ;
  assign n36579 = n553 & ~n36578 ;
  assign n36580 = ~n2534 & n16431 ;
  assign n36581 = ( n612 & n9687 ) | ( n612 & ~n36580 ) | ( n9687 & ~n36580 ) ;
  assign n36582 = n843 & ~n4536 ;
  assign n36583 = ~n1768 & n36582 ;
  assign n36584 = n2639 | n7932 ;
  assign n36585 = n1175 & ~n36584 ;
  assign n36586 = ~n1469 & n15979 ;
  assign n36587 = n20107 ^ n185 ^ 1'b0 ;
  assign n36588 = n36586 & n36587 ;
  assign n36589 = n24008 ^ n8044 ^ 1'b0 ;
  assign n36590 = ~n19730 & n36589 ;
  assign n36591 = n15536 ^ n10177 ^ 1'b0 ;
  assign n36592 = n930 & n36591 ;
  assign n36593 = n22536 ^ n1392 ^ 1'b0 ;
  assign n36594 = n9215 | n16645 ;
  assign n36595 = n36593 & ~n36594 ;
  assign n36596 = n17705 | n36595 ;
  assign n36597 = n36596 ^ n2640 ^ 1'b0 ;
  assign n36598 = n1445 & n36597 ;
  assign n36599 = n36598 ^ n19356 ^ 1'b0 ;
  assign n36600 = n11359 ^ n4037 ^ 1'b0 ;
  assign n36601 = ~n964 & n32175 ;
  assign n36602 = ~n13039 & n36601 ;
  assign n36603 = n14920 ^ n7397 ^ 1'b0 ;
  assign n36604 = n13654 ^ n3886 ^ 1'b0 ;
  assign n36605 = ~n36603 & n36604 ;
  assign n36606 = n25533 ^ n20847 ^ 1'b0 ;
  assign n36607 = n21199 | n28284 ;
  assign n36608 = n8489 ^ n520 ^ 1'b0 ;
  assign n36609 = n495 & ~n36608 ;
  assign n36610 = n294 & n3584 ;
  assign n36611 = n36610 ^ n19095 ^ 1'b0 ;
  assign n36612 = ( n412 & n36609 ) | ( n412 & ~n36611 ) | ( n36609 & ~n36611 ) ;
  assign n36613 = n5180 ^ n2073 ^ 1'b0 ;
  assign n36614 = n16158 & ~n36613 ;
  assign n36615 = ~n3862 & n36614 ;
  assign n36616 = n36615 ^ n642 ^ n616 ;
  assign n36617 = ~n3415 & n36616 ;
  assign n36618 = n1870 & ~n18028 ;
  assign n36619 = n15481 | n36618 ;
  assign n36620 = n14694 | n19627 ;
  assign n36621 = n36620 ^ n36273 ^ 1'b0 ;
  assign n36622 = n16195 & ~n26184 ;
  assign n36623 = n2792 & n36622 ;
  assign n36624 = n748 & n24714 ;
  assign n36625 = n36624 ^ n22590 ^ n5241 ;
  assign n36626 = n9966 ^ n2157 ^ 1'b0 ;
  assign n36627 = n4171 | n14737 ;
  assign n36628 = n36626 & ~n36627 ;
  assign n36629 = ~n4700 & n34604 ;
  assign n36630 = ~n19830 & n36629 ;
  assign n36631 = n13547 & ~n21959 ;
  assign n36632 = n36631 ^ n22410 ^ 1'b0 ;
  assign n36633 = n15824 ^ n13691 ^ 1'b0 ;
  assign n36634 = ~n2512 & n36633 ;
  assign n36635 = n9714 & n36268 ;
  assign n36636 = n1518 | n14450 ;
  assign n36637 = n13930 | n36636 ;
  assign n36638 = n11585 ^ n3885 ^ 1'b0 ;
  assign n36639 = n10705 ^ n1339 ^ 1'b0 ;
  assign n36640 = n36638 & n36639 ;
  assign n36641 = n7901 | n16505 ;
  assign n36642 = n23678 & n36641 ;
  assign n36643 = ~n25697 & n36642 ;
  assign n36644 = n776 & n12357 ;
  assign n36645 = n36643 & n36644 ;
  assign n36646 = n2083 & n34500 ;
  assign n36647 = n11479 & ~n36646 ;
  assign n36648 = n1388 | n26452 ;
  assign n36649 = n23025 & n36648 ;
  assign n36650 = n3221 & ~n9353 ;
  assign n36651 = n17667 & n36650 ;
  assign n36652 = n3962 & n21878 ;
  assign n36657 = n1462 | n17774 ;
  assign n36658 = n5516 & n36657 ;
  assign n36653 = n1707 & ~n3208 ;
  assign n36654 = n36653 ^ n6849 ^ 1'b0 ;
  assign n36655 = n8893 | n14730 ;
  assign n36656 = n36654 | n36655 ;
  assign n36659 = n36658 ^ n36656 ^ n4211 ;
  assign n36660 = n528 & n1530 ;
  assign n36661 = ~n10743 & n27201 ;
  assign n36662 = ( n10131 & ~n14111 ) | ( n10131 & n26552 ) | ( ~n14111 & n26552 ) ;
  assign n36663 = ~n21464 & n36662 ;
  assign n36664 = n36663 ^ n31559 ^ 1'b0 ;
  assign n36665 = n1132 & ~n36664 ;
  assign n36666 = n11592 ^ n10942 ^ 1'b0 ;
  assign n36667 = ~n19776 & n36666 ;
  assign n36668 = n24047 ^ n1904 ^ 1'b0 ;
  assign n36669 = ~n30025 & n36668 ;
  assign n36670 = n13981 ^ n6300 ^ 1'b0 ;
  assign n36671 = n36670 ^ n12649 ^ 1'b0 ;
  assign n36672 = n36669 & ~n36671 ;
  assign n36673 = n4288 & ~n18655 ;
  assign n36674 = n36673 ^ n3757 ^ 1'b0 ;
  assign n36675 = n6419 & ~n7872 ;
  assign n36676 = n3068 & n9756 ;
  assign n36677 = ( ~n2754 & n36675 ) | ( ~n2754 & n36676 ) | ( n36675 & n36676 ) ;
  assign n36678 = n977 & n2310 ;
  assign n36679 = n15901 ^ n7008 ^ 1'b0 ;
  assign n36680 = n36678 | n36679 ;
  assign n36681 = n1602 | n5634 ;
  assign n36682 = n6298 & n31219 ;
  assign n36683 = n36681 & n36682 ;
  assign n36684 = n5696 | n28750 ;
  assign n36685 = n3646 | n11837 ;
  assign n36686 = n14388 | n36685 ;
  assign n36687 = n30549 ^ n1936 ^ 1'b0 ;
  assign n36688 = n8770 & n36687 ;
  assign n36689 = n28944 ^ n6016 ^ 1'b0 ;
  assign n36691 = n5530 & ~n8570 ;
  assign n36690 = n12421 & ~n20215 ;
  assign n36692 = n36691 ^ n36690 ^ 1'b0 ;
  assign n36693 = n36692 ^ n6181 ^ n296 ;
  assign n36694 = n16296 ^ n3471 ^ 1'b0 ;
  assign n36695 = n10527 | n36694 ;
  assign n36696 = n36695 ^ n22471 ^ 1'b0 ;
  assign n36697 = n14941 ^ n9023 ^ 1'b0 ;
  assign n36698 = n3950 | n13775 ;
  assign n36699 = ~n36697 & n36698 ;
  assign n36700 = n322 & n36699 ;
  assign n36701 = n36700 ^ n15983 ^ 1'b0 ;
  assign n36702 = n27433 ^ n21584 ^ 1'b0 ;
  assign n36703 = n36702 ^ n18007 ^ 1'b0 ;
  assign n36704 = n10099 ^ n183 ^ 1'b0 ;
  assign n36705 = n26741 | n36704 ;
  assign n36706 = n2983 | n20339 ;
  assign n36707 = n36705 & ~n36706 ;
  assign n36708 = n8995 ^ n690 ^ 1'b0 ;
  assign n36709 = n8458 & n10393 ;
  assign n36710 = n36709 ^ n7221 ^ 1'b0 ;
  assign n36711 = n1528 | n16333 ;
  assign n36712 = n6094 ^ n1884 ^ 1'b0 ;
  assign n36713 = n36711 & n36712 ;
  assign n36714 = ~n866 & n8002 ;
  assign n36715 = n22850 ^ n17473 ^ 1'b0 ;
  assign n36716 = n13747 | n22487 ;
  assign n36717 = n36715 & ~n36716 ;
  assign n36718 = n36714 & ~n36717 ;
  assign n36719 = n36718 ^ n20027 ^ 1'b0 ;
  assign n36720 = n10390 & ~n14759 ;
  assign n36721 = n36720 ^ n4791 ^ 1'b0 ;
  assign n36722 = n10663 ^ n1202 ^ 1'b0 ;
  assign n36723 = n36722 ^ n14236 ^ n12663 ;
  assign n36724 = n35427 & ~n36723 ;
  assign n36725 = n13237 | n16182 ;
  assign n36726 = n10438 | n36725 ;
  assign n36727 = n28822 | n36726 ;
  assign n36728 = n14558 ^ n8740 ^ 1'b0 ;
  assign n36729 = n34111 | n36728 ;
  assign n36730 = n512 | n36729 ;
  assign n36731 = n36730 ^ n14731 ^ 1'b0 ;
  assign n36733 = n23197 ^ n2517 ^ 1'b0 ;
  assign n36732 = n1732 & ~n5749 ;
  assign n36734 = n36733 ^ n36732 ^ n10674 ;
  assign n36735 = n36734 ^ n958 ^ 1'b0 ;
  assign n36736 = ( n7460 & ~n14447 ) | ( n7460 & n27666 ) | ( ~n14447 & n27666 ) ;
  assign n36737 = n5309 ^ n561 ^ 1'b0 ;
  assign n36738 = ~n5994 & n36737 ;
  assign n36739 = n36738 ^ n6447 ^ 1'b0 ;
  assign n36740 = n506 & n9498 ;
  assign n36741 = n28396 ^ n28357 ^ 1'b0 ;
  assign n36743 = n18963 ^ n1375 ^ 1'b0 ;
  assign n36742 = n12982 ^ n7192 ^ 1'b0 ;
  assign n36744 = n36743 ^ n36742 ^ 1'b0 ;
  assign n36745 = n22610 & n36744 ;
  assign n36746 = n29077 & n36745 ;
  assign n36747 = n9309 & ~n13099 ;
  assign n36748 = n8877 & n20833 ;
  assign n36749 = n16072 & n36748 ;
  assign n36750 = n26441 ^ n14844 ^ 1'b0 ;
  assign n36751 = ~n36749 & n36750 ;
  assign n36752 = ~n24553 & n25274 ;
  assign n36753 = ~n6023 & n20576 ;
  assign n36754 = n1435 | n27286 ;
  assign n36755 = n21037 & n32534 ;
  assign n36756 = n6700 ^ n5397 ^ 1'b0 ;
  assign n36757 = n6242 | n36756 ;
  assign n36758 = n812 & n2517 ;
  assign n36759 = n36758 ^ n815 ^ 1'b0 ;
  assign n36760 = ~n6028 & n36759 ;
  assign n36761 = n2252 & ~n32524 ;
  assign n36762 = n36761 ^ n11167 ^ 1'b0 ;
  assign n36763 = n14845 & n23035 ;
  assign n36764 = n36763 ^ n89 ^ 1'b0 ;
  assign n36765 = n688 | n3514 ;
  assign n36766 = n2684 ^ n1659 ^ 1'b0 ;
  assign n36767 = n36765 & ~n36766 ;
  assign n36768 = ~n354 & n9252 ;
  assign n36769 = n11061 ^ n6933 ^ 1'b0 ;
  assign n36770 = n2511 | n36769 ;
  assign n36771 = n36768 | n36770 ;
  assign n36772 = n23683 ^ n15400 ^ 1'b0 ;
  assign n36773 = n395 | n36772 ;
  assign n36774 = n3988 & n35185 ;
  assign n36775 = n36773 & n36774 ;
  assign n36776 = ( n3653 & n5099 ) | ( n3653 & n5135 ) | ( n5099 & n5135 ) ;
  assign n36777 = n6904 & n36776 ;
  assign n36778 = n9732 & n36777 ;
  assign n36779 = n2694 & ~n22186 ;
  assign n36780 = n36779 ^ n6154 ^ 1'b0 ;
  assign n36781 = ~n13073 & n36220 ;
  assign n36782 = n36471 ^ n3599 ^ n2495 ;
  assign n36783 = n30606 & ~n34446 ;
  assign n36784 = n36783 ^ n12206 ^ 1'b0 ;
  assign n36785 = n148 & n15769 ;
  assign n36786 = ~n13110 & n36785 ;
  assign n36787 = n15925 ^ n14906 ^ n9630 ;
  assign n36788 = ~n36786 & n36787 ;
  assign n36789 = n4307 & n21131 ;
  assign n36790 = n2767 | n36789 ;
  assign n36791 = n36790 ^ n6295 ^ 1'b0 ;
  assign n36793 = n13171 ^ n3664 ^ 1'b0 ;
  assign n36792 = n3107 & ~n20197 ;
  assign n36794 = n36793 ^ n36792 ^ 1'b0 ;
  assign n36795 = ~n24353 & n31488 ;
  assign n36796 = ~n16406 & n36795 ;
  assign n36797 = n2978 | n36623 ;
  assign n36798 = n36797 ^ n26240 ^ 1'b0 ;
  assign n36799 = n18530 ^ n8169 ^ 1'b0 ;
  assign n36800 = n2348 & n36799 ;
  assign n36801 = ~n12939 & n36800 ;
  assign n36802 = n12271 ^ n7904 ^ 1'b0 ;
  assign n36803 = ~n36801 & n36802 ;
  assign n36804 = n22792 ^ n20531 ^ 1'b0 ;
  assign n36805 = n5956 | n36804 ;
  assign n36806 = ~n3921 & n35238 ;
  assign n36807 = n17066 ^ n15769 ^ 1'b0 ;
  assign n36808 = n3467 | n5535 ;
  assign n36809 = n36808 ^ n5359 ^ 1'b0 ;
  assign n36810 = n36809 ^ n3080 ^ 1'b0 ;
  assign n36811 = n36810 ^ n16762 ^ n8788 ;
  assign n36812 = n15625 & ~n20824 ;
  assign n36813 = ~n5473 & n15196 ;
  assign n36814 = n30011 & n36813 ;
  assign n36815 = n1105 ^ n164 ^ 1'b0 ;
  assign n36816 = ~n7360 & n36815 ;
  assign n36817 = n8652 & n36816 ;
  assign n36818 = ~n14884 & n36817 ;
  assign n36819 = n4336 & n35692 ;
  assign n36820 = n36819 ^ n22967 ^ 1'b0 ;
  assign n36821 = n13778 ^ n649 ^ 1'b0 ;
  assign n36822 = n2456 | n24313 ;
  assign n36823 = n36822 ^ n13330 ^ 1'b0 ;
  assign n36824 = n34188 ^ n11079 ^ 1'b0 ;
  assign n36825 = ~n35508 & n36824 ;
  assign n36826 = ~n21506 & n33489 ;
  assign n36827 = n17532 ^ n4485 ^ n3648 ;
  assign n36828 = n14085 ^ n9596 ^ 1'b0 ;
  assign n36829 = n23802 | n36468 ;
  assign n36830 = n19181 ^ n12892 ^ 1'b0 ;
  assign n36831 = n14158 & ~n28607 ;
  assign n36832 = n36831 ^ n10882 ^ 1'b0 ;
  assign n36833 = n599 | n12982 ;
  assign n36834 = n3558 | n36833 ;
  assign n36835 = n9344 & ~n36834 ;
  assign n36836 = n2672 ^ n1220 ^ 1'b0 ;
  assign n36837 = n7126 & n36836 ;
  assign n36838 = n36837 ^ n34583 ^ 1'b0 ;
  assign n36840 = n17705 ^ n757 ^ 1'b0 ;
  assign n36841 = n33492 & n36840 ;
  assign n36839 = n26733 & n33845 ;
  assign n36842 = n36841 ^ n36839 ^ 1'b0 ;
  assign n36843 = n7791 | n31234 ;
  assign n36844 = n13792 & ~n31107 ;
  assign n36845 = n36844 ^ n5927 ^ 1'b0 ;
  assign n36846 = n35062 ^ n4396 ^ n1388 ;
  assign n36847 = n687 | n13713 ;
  assign n36848 = n36847 ^ n33142 ^ 1'b0 ;
  assign n36849 = n36848 ^ n12537 ^ 1'b0 ;
  assign n36850 = n2209 | n9171 ;
  assign n36851 = n2373 & ~n19826 ;
  assign n36852 = ~n3600 & n31108 ;
  assign n36853 = n36852 ^ n7489 ^ 1'b0 ;
  assign n36854 = ~n34756 & n35084 ;
  assign n36855 = n23108 ^ n13892 ^ 1'b0 ;
  assign n36856 = ~n14333 & n36855 ;
  assign n36857 = n36856 ^ n19124 ^ 1'b0 ;
  assign n36858 = ( n8148 & ~n10395 ) | ( n8148 & n18353 ) | ( ~n10395 & n18353 ) ;
  assign n36859 = ~n7580 & n11036 ;
  assign n36860 = n6015 | n8210 ;
  assign n36861 = n3061 & ~n8248 ;
  assign n36862 = n36861 ^ n10652 ^ 1'b0 ;
  assign n36863 = n28810 ^ n12289 ^ 1'b0 ;
  assign n36864 = n22676 ^ n5182 ^ 1'b0 ;
  assign n36865 = n11483 ^ n37 ^ 1'b0 ;
  assign n36866 = ~n13752 & n14328 ;
  assign n36867 = n2059 & ~n10753 ;
  assign n36868 = ~n13111 & n36867 ;
  assign n36869 = n7005 & n33533 ;
  assign n36870 = n36869 ^ n5024 ^ 1'b0 ;
  assign n36871 = n12324 & n13011 ;
  assign n36872 = n9833 ^ n1057 ^ 1'b0 ;
  assign n36873 = n2301 & n36872 ;
  assign n36874 = n36873 ^ n21399 ^ 1'b0 ;
  assign n36875 = n25766 ^ n1210 ^ 1'b0 ;
  assign n36876 = ~n1793 & n19961 ;
  assign n36877 = ~n6764 & n16509 ;
  assign n36878 = ~n6841 & n36877 ;
  assign n36881 = n11556 & n24370 ;
  assign n36879 = n5830 | n9834 ;
  assign n36880 = n5378 & ~n36879 ;
  assign n36882 = n36881 ^ n36880 ^ n6443 ;
  assign n36883 = n4919 & ~n36882 ;
  assign n36884 = n25488 | n36883 ;
  assign n36885 = n22052 ^ n3138 ^ 1'b0 ;
  assign n36886 = n24615 | n35672 ;
  assign n36887 = n36886 ^ n879 ^ 1'b0 ;
  assign n36888 = ( ~n8946 & n10763 ) | ( ~n8946 & n36887 ) | ( n10763 & n36887 ) ;
  assign n36889 = n14255 | n36888 ;
  assign n36890 = n36889 ^ n1431 ^ 1'b0 ;
  assign n36891 = n16157 ^ n582 ^ 1'b0 ;
  assign n36892 = ~n7589 & n36891 ;
  assign n36893 = n15843 ^ n1447 ^ 1'b0 ;
  assign n36894 = n1870 & ~n36893 ;
  assign n36895 = n18091 | n21604 ;
  assign n36896 = n2018 | n36895 ;
  assign n36897 = n36896 ^ n18096 ^ 1'b0 ;
  assign n36898 = n7920 & n36897 ;
  assign n36899 = n5830 ^ n3897 ^ 1'b0 ;
  assign n36900 = n18308 | n36899 ;
  assign n36901 = n36900 ^ n6207 ^ n278 ;
  assign n36902 = n6141 ^ n4264 ^ 1'b0 ;
  assign n36903 = n36902 ^ n3265 ^ 1'b0 ;
  assign n36904 = n4449 ^ n1893 ^ 1'b0 ;
  assign n36905 = ~n4037 & n36904 ;
  assign n36906 = n11837 ^ n11409 ^ 1'b0 ;
  assign n36907 = n16280 ^ n1029 ^ 1'b0 ;
  assign n36908 = ~n677 & n4186 ;
  assign n36909 = n5172 & n36908 ;
  assign n36914 = n4004 | n12605 ;
  assign n36915 = n4004 & ~n36914 ;
  assign n36916 = n1541 & ~n31397 ;
  assign n36917 = ~n1541 & n36916 ;
  assign n36918 = n4281 & ~n36917 ;
  assign n36919 = ~n4281 & n36918 ;
  assign n36920 = n4689 | n36919 ;
  assign n36921 = n36915 & ~n36920 ;
  assign n36913 = n3183 & n26780 ;
  assign n36922 = n36921 ^ n36913 ^ 1'b0 ;
  assign n36910 = n861 & ~n3985 ;
  assign n36911 = n3985 & n36910 ;
  assign n36912 = n31418 & ~n36911 ;
  assign n36923 = n36922 ^ n36912 ^ 1'b0 ;
  assign n36924 = n23929 & ~n36923 ;
  assign n36925 = n18594 & n36924 ;
  assign n36926 = n2733 & n12418 ;
  assign n36927 = n36926 ^ n2128 ^ 1'b0 ;
  assign n36928 = n5507 | n8321 ;
  assign n36929 = n36928 ^ n4774 ^ 1'b0 ;
  assign n36930 = n36929 ^ n20697 ^ n6566 ;
  assign n36931 = n23655 & ~n36930 ;
  assign n36932 = n1246 & n36931 ;
  assign n36933 = n15921 ^ n253 ^ 1'b0 ;
  assign n36934 = n36932 | n36933 ;
  assign n36935 = n2346 | n36934 ;
  assign n36936 = n1295 & ~n8688 ;
  assign n36937 = n9922 | n36936 ;
  assign n36938 = n1585 | n36937 ;
  assign n36939 = ~n16760 & n25946 ;
  assign n36940 = n36939 ^ n9570 ^ 1'b0 ;
  assign n36941 = n29943 ^ n26945 ^ 1'b0 ;
  assign n36942 = n25872 & ~n36941 ;
  assign n36943 = n15604 & n36942 ;
  assign n36944 = n6629 & n19915 ;
  assign n36945 = n36944 ^ n1003 ^ 1'b0 ;
  assign n36946 = n2433 & n36218 ;
  assign n36947 = ~n36133 & n36946 ;
  assign n36948 = ~n3523 & n4850 ;
  assign n36949 = n9918 ^ n1057 ^ 1'b0 ;
  assign n36950 = ~n32944 & n36949 ;
  assign n36951 = n9086 & n19954 ;
  assign n36952 = n36951 ^ n182 ^ 1'b0 ;
  assign n36953 = ~n18396 & n27244 ;
  assign n36954 = ( n4644 & n7069 ) | ( n4644 & n25922 ) | ( n7069 & n25922 ) ;
  assign n36955 = n31301 ^ n647 ^ 1'b0 ;
  assign n36956 = n9381 & ~n28446 ;
  assign n36957 = n36956 ^ n34470 ^ 1'b0 ;
  assign n36958 = n24204 & n27435 ;
  assign n36959 = n20520 ^ n8141 ^ 1'b0 ;
  assign n36960 = n23222 ^ n18370 ^ 1'b0 ;
  assign n36961 = n4072 ^ n288 ^ 1'b0 ;
  assign n36962 = ~n8981 & n36961 ;
  assign n36963 = n36960 & ~n36962 ;
  assign n36964 = n689 & n2903 ;
  assign n36965 = n4078 | n9809 ;
  assign n36966 = n36964 | n36965 ;
  assign n36967 = n330 | n17607 ;
  assign n36968 = ( ~n14753 & n16454 ) | ( ~n14753 & n36967 ) | ( n16454 & n36967 ) ;
  assign n36969 = n602 & ~n10346 ;
  assign n36970 = ~n122 & n2881 ;
  assign n36971 = n2349 & n36970 ;
  assign n36972 = n20263 | n36971 ;
  assign n36973 = n36969 & ~n36972 ;
  assign n36974 = ~n960 & n20189 ;
  assign n36975 = n4662 & n19610 ;
  assign n36976 = n36975 ^ n9917 ^ 1'b0 ;
  assign n36977 = n1151 & ~n36976 ;
  assign n36978 = n759 & n1948 ;
  assign n36979 = n36978 ^ n14587 ^ 1'b0 ;
  assign n36980 = n23137 | n33233 ;
  assign n36981 = n36979 & ~n36980 ;
  assign n36982 = n23463 | n35611 ;
  assign n36983 = ~n36981 & n36982 ;
  assign n36984 = n5588 & n28745 ;
  assign n36985 = ~n25952 & n36984 ;
  assign n36986 = n7526 & ~n36985 ;
  assign n36987 = n33788 ^ n20330 ^ n4673 ;
  assign n36988 = n32759 & n36987 ;
  assign n36989 = ~n25867 & n29803 ;
  assign n36990 = n5438 | n7056 ;
  assign n36991 = n1315 & ~n34514 ;
  assign n36992 = n36991 ^ n2185 ^ 1'b0 ;
  assign n36993 = n5942 & n36992 ;
  assign n36994 = ~n36990 & n36993 ;
  assign n36995 = ~n632 & n19575 ;
  assign n36996 = ~n7105 & n36995 ;
  assign n36997 = n1920 | n36996 ;
  assign n36998 = n31903 ^ n18104 ^ 1'b0 ;
  assign n36999 = ~n36997 & n36998 ;
  assign n37000 = n3371 & ~n20747 ;
  assign n37001 = n11063 & ~n13600 ;
  assign n37002 = n6371 ^ n4604 ^ 1'b0 ;
  assign n37003 = n7882 | n37002 ;
  assign n37004 = n37003 ^ n3346 ^ 1'b0 ;
  assign n37005 = ~n5176 & n37004 ;
  assign n37006 = ( n9081 & n25417 ) | ( n9081 & ~n37005 ) | ( n25417 & ~n37005 ) ;
  assign n37007 = n37006 ^ n36689 ^ 1'b0 ;
  assign n37008 = n7205 | n19654 ;
  assign n37009 = n12241 ^ n2829 ^ 1'b0 ;
  assign n37010 = ~n9394 & n37009 ;
  assign n37011 = ~n10349 & n37010 ;
  assign n37012 = n19131 | n35322 ;
  assign n37013 = n12316 | n37012 ;
  assign n37014 = n21063 ^ n4419 ^ 1'b0 ;
  assign n37015 = n602 & ~n37014 ;
  assign n37016 = n37015 ^ n22118 ^ 1'b0 ;
  assign n37020 = n5908 & n11868 ;
  assign n37021 = n7299 & n37020 ;
  assign n37022 = n7609 & ~n37021 ;
  assign n37019 = n9898 & ~n12402 ;
  assign n37017 = n10768 & ~n21976 ;
  assign n37018 = n37017 ^ n22593 ^ 1'b0 ;
  assign n37023 = n37022 ^ n37019 ^ n37018 ;
  assign n37025 = n6061 ^ n1315 ^ 1'b0 ;
  assign n37024 = ~n30691 & n30991 ;
  assign n37026 = n37025 ^ n37024 ^ 1'b0 ;
  assign n37027 = n14142 ^ n4631 ^ 1'b0 ;
  assign n37028 = n1847 & ~n37027 ;
  assign n37029 = n2917 & ~n4776 ;
  assign n37030 = n24637 ^ n8869 ^ 1'b0 ;
  assign n37031 = n26965 & n37030 ;
  assign n37032 = n23390 ^ n7456 ^ n928 ;
  assign n37033 = n27991 ^ n4093 ^ 1'b0 ;
  assign n37034 = n15986 ^ n10470 ^ n4209 ;
  assign n37035 = n32472 & ~n37034 ;
  assign n37036 = n5603 ^ n3584 ^ 1'b0 ;
  assign n37037 = n9451 & n37036 ;
  assign n37038 = n847 | n10025 ;
  assign n37039 = n184 & ~n37038 ;
  assign n37040 = n37039 ^ n17205 ^ 1'b0 ;
  assign n37041 = n17058 & n37040 ;
  assign n37042 = ~n26537 & n36202 ;
  assign n37043 = n37042 ^ n1907 ^ 1'b0 ;
  assign n37044 = n13135 | n25315 ;
  assign n37045 = n8463 & n24512 ;
  assign n37046 = n37045 ^ n1859 ^ 1'b0 ;
  assign n37049 = n25537 ^ n3137 ^ 1'b0 ;
  assign n37047 = n32482 ^ n6510 ^ 1'b0 ;
  assign n37048 = x0 & ~n37047 ;
  assign n37050 = n37049 ^ n37048 ^ 1'b0 ;
  assign n37051 = n633 & ~n5790 ;
  assign n37052 = n2642 ^ n984 ^ 1'b0 ;
  assign n37053 = n4848 & n37052 ;
  assign n37054 = n37053 ^ n13198 ^ 1'b0 ;
  assign n37055 = ~n37051 & n37054 ;
  assign n37056 = n37055 ^ n36242 ^ n14924 ;
  assign n37057 = n3399 | n24825 ;
  assign n37058 = n31715 | n37057 ;
  assign n37059 = ~n2595 & n6466 ;
  assign n37060 = n23302 ^ n10036 ^ 1'b0 ;
  assign n37061 = n37059 | n37060 ;
  assign n37062 = ( n4770 & n23589 ) | ( n4770 & ~n35893 ) | ( n23589 & ~n35893 ) ;
  assign n37063 = n31215 ^ n15468 ^ 1'b0 ;
  assign n37064 = n33121 & n37063 ;
  assign n37065 = n3194 & ~n13855 ;
  assign n37066 = n3238 & ~n3409 ;
  assign n37067 = n3409 & n37066 ;
  assign n37068 = n5380 & ~n20207 ;
  assign n37069 = n37067 & n37068 ;
  assign n37070 = ~n8141 & n28543 ;
  assign n37071 = ~n28543 & n37070 ;
  assign n37072 = n29144 & ~n37071 ;
  assign n37073 = ~n37069 & n37072 ;
  assign n37074 = n37069 & n37073 ;
  assign n37075 = n2577 | n21225 ;
  assign n37076 = n12436 ^ n7491 ^ 1'b0 ;
  assign n37077 = n7143 & ~n37076 ;
  assign n37078 = n2283 & ~n37077 ;
  assign n37079 = ~n10584 & n16088 ;
  assign n37080 = n37079 ^ n17486 ^ 1'b0 ;
  assign n37081 = n196 & ~n10255 ;
  assign n37082 = n1144 & ~n19158 ;
  assign n37083 = n2072 & n16417 ;
  assign n37084 = ~n1438 & n10230 ;
  assign n37085 = n6611 ^ n1219 ^ 1'b0 ;
  assign n37086 = ~n2629 & n8594 ;
  assign n37087 = n9130 | n18003 ;
  assign n37088 = ( n9699 & ~n15015 ) | ( n9699 & n37087 ) | ( ~n15015 & n37087 ) ;
  assign n37089 = n736 & ~n10819 ;
  assign n37090 = ~n7981 & n8171 ;
  assign n37091 = ~n185 & n37090 ;
  assign n37092 = n3437 & ~n37091 ;
  assign n37093 = n7272 & n11917 ;
  assign n37094 = n1516 & n9619 ;
  assign n37095 = ~n37093 & n37094 ;
  assign n37096 = n31779 ^ n5284 ^ 1'b0 ;
  assign n37097 = n175 | n37096 ;
  assign n37098 = n37097 ^ n10731 ^ 1'b0 ;
  assign n37099 = n20697 ^ n3423 ^ 1'b0 ;
  assign n37100 = n15721 ^ n10367 ^ 1'b0 ;
  assign n37101 = n367 & n37100 ;
  assign n37102 = n1900 & ~n16700 ;
  assign n37103 = ~n37101 & n37102 ;
  assign n37104 = ~n4655 & n31070 ;
  assign n37105 = n37104 ^ n4000 ^ 1'b0 ;
  assign n37106 = n37103 | n37105 ;
  assign n37107 = n37106 ^ n23910 ^ 1'b0 ;
  assign n37108 = n12292 ^ n5809 ^ 1'b0 ;
  assign n37109 = n29358 & ~n37108 ;
  assign n37110 = n1626 & n28239 ;
  assign n37111 = ~n37109 & n37110 ;
  assign n37112 = n16198 ^ n2996 ^ 1'b0 ;
  assign n37113 = n627 & ~n14552 ;
  assign n37114 = ~n37112 & n37113 ;
  assign n37115 = ~n14590 & n14990 ;
  assign n37116 = n37115 ^ n27148 ^ 1'b0 ;
  assign n37117 = n37116 ^ n22542 ^ 1'b0 ;
  assign n37118 = n27 & n37117 ;
  assign n37119 = n37114 & n37118 ;
  assign n37120 = n24032 ^ n6408 ^ 1'b0 ;
  assign n37121 = ~n14815 & n18733 ;
  assign n37122 = n10265 ^ n8747 ^ 1'b0 ;
  assign n37123 = ~n37121 & n37122 ;
  assign n37124 = n23473 ^ n11723 ^ 1'b0 ;
  assign n37125 = n977 | n7264 ;
  assign n37126 = n29719 | n37125 ;
  assign n37127 = n3682 & n11957 ;
  assign n37128 = ~n7792 & n37127 ;
  assign n37129 = n18962 ^ n4917 ^ 1'b0 ;
  assign n37130 = n7449 & n8099 ;
  assign n37131 = n15297 & n37130 ;
  assign n37132 = n1474 | n37131 ;
  assign n37133 = n11641 ^ n6595 ^ 1'b0 ;
  assign n37134 = n3725 & n37133 ;
  assign n37135 = n18765 & n37134 ;
  assign n37136 = n37135 ^ n5469 ^ 1'b0 ;
  assign n37137 = n3068 & ~n37136 ;
  assign n37138 = n1928 & n2218 ;
  assign n37139 = ~n7309 & n37138 ;
  assign n37140 = n17528 & ~n37139 ;
  assign n37141 = n37140 ^ n1226 ^ 1'b0 ;
  assign n37142 = n24937 ^ n1513 ^ 1'b0 ;
  assign n37143 = n367 & ~n37142 ;
  assign n37147 = n2027 | n32096 ;
  assign n37148 = n27219 | n37147 ;
  assign n37144 = n4022 & ~n4552 ;
  assign n37145 = n37144 ^ n17257 ^ 1'b0 ;
  assign n37146 = n8262 & ~n37145 ;
  assign n37149 = n37148 ^ n37146 ^ 1'b0 ;
  assign n37150 = ~n5380 & n16810 ;
  assign n37151 = n5538 & n8046 ;
  assign n37152 = n13548 ^ n5495 ^ 1'b0 ;
  assign n37153 = n9698 | n37152 ;
  assign n37154 = ~n14376 & n27240 ;
  assign n37155 = ~n14991 & n24081 ;
  assign n37156 = n33200 ^ n18537 ^ 1'b0 ;
  assign n37157 = n86 | n37156 ;
  assign n37158 = n3434 | n37157 ;
  assign n37160 = n14142 | n26570 ;
  assign n37159 = n30956 ^ n2292 ^ 1'b0 ;
  assign n37161 = n37160 ^ n37159 ^ 1'b0 ;
  assign n37162 = n14614 & ~n28347 ;
  assign n37163 = ~n30985 & n37162 ;
  assign n37164 = n246 | n34111 ;
  assign n37165 = n20025 & ~n37164 ;
  assign n37166 = n1879 & n11643 ;
  assign n37167 = ~n15261 & n37166 ;
  assign n37168 = n37167 ^ n10078 ^ 1'b0 ;
  assign n37169 = n17675 & ~n37168 ;
  assign n37170 = n1112 | n37169 ;
  assign n37171 = n5812 ^ n4061 ^ 1'b0 ;
  assign n37172 = ~n954 & n12411 ;
  assign n37173 = n12552 | n22616 ;
  assign n37174 = n18207 ^ n55 ^ 1'b0 ;
  assign n37175 = ~n33699 & n37174 ;
  assign n37176 = ~n5096 & n27876 ;
  assign n37177 = n3668 ^ n340 ^ 1'b0 ;
  assign n37178 = n3417 ^ n818 ^ 1'b0 ;
  assign n37179 = n10141 & ~n37178 ;
  assign n37180 = n20585 & n37179 ;
  assign n37181 = n1535 | n8312 ;
  assign n37182 = ~n5323 & n24516 ;
  assign n37183 = n37182 ^ n33695 ^ 1'b0 ;
  assign n37184 = n1287 & ~n13244 ;
  assign n37185 = n1243 & n37184 ;
  assign n37186 = n8158 | n18484 ;
  assign n37187 = n37185 & ~n37186 ;
  assign n37188 = n8189 & ~n37187 ;
  assign n37189 = ~n5398 & n37188 ;
  assign n37190 = n3019 ^ n2127 ^ 1'b0 ;
  assign n37191 = n16853 ^ n1181 ^ 1'b0 ;
  assign n37192 = n21173 | n37191 ;
  assign n37194 = n3151 ^ n1582 ^ 1'b0 ;
  assign n37193 = n3498 & ~n13755 ;
  assign n37195 = n37194 ^ n37193 ^ 1'b0 ;
  assign n37197 = ~n2608 & n35535 ;
  assign n37196 = n5793 | n37051 ;
  assign n37198 = n37197 ^ n37196 ^ 1'b0 ;
  assign n37199 = n553 ^ n60 ^ 1'b0 ;
  assign n37200 = n37198 & ~n37199 ;
  assign n37201 = n16700 ^ n14556 ^ 1'b0 ;
  assign n37202 = ~n1309 & n25620 ;
  assign n37203 = n14975 ^ n11902 ^ 1'b0 ;
  assign n37204 = n28399 ^ n17052 ^ 1'b0 ;
  assign n37205 = n12563 & ~n15166 ;
  assign n37206 = n37205 ^ n32572 ^ 1'b0 ;
  assign n37207 = n19530 & n37206 ;
  assign n37208 = n16302 | n30120 ;
  assign n37210 = n7268 & n8039 ;
  assign n37209 = n17487 | n21788 ;
  assign n37211 = n37210 ^ n37209 ^ 1'b0 ;
  assign n37212 = n270 & ~n37211 ;
  assign n37213 = n11375 ^ n614 ^ 1'b0 ;
  assign n37214 = n27504 & n37213 ;
  assign n37215 = ~n4432 & n22482 ;
  assign n37216 = n37215 ^ n10364 ^ 1'b0 ;
  assign n37217 = n528 | n3244 ;
  assign n37218 = n6601 | n37217 ;
  assign n37219 = n20432 | n37218 ;
  assign n37220 = n38 | n8561 ;
  assign n37221 = ~n13556 & n37220 ;
  assign n37222 = ( n7896 & n32700 ) | ( n7896 & ~n37221 ) | ( n32700 & ~n37221 ) ;
  assign n37223 = n29175 | n32008 ;
  assign n37224 = n3887 & n4329 ;
  assign n37225 = n60 & n37224 ;
  assign n37226 = ~n20201 & n37225 ;
  assign n37227 = n11234 | n24437 ;
  assign n37232 = n23775 ^ n17892 ^ 1'b0 ;
  assign n37228 = n715 & ~n7568 ;
  assign n37229 = n6752 & n37228 ;
  assign n37230 = n37229 ^ n5471 ^ 1'b0 ;
  assign n37231 = ~n10117 & n37230 ;
  assign n37233 = n37232 ^ n37231 ^ 1'b0 ;
  assign n37234 = n2361 & ~n20691 ;
  assign n37235 = ~n3141 & n12436 ;
  assign n37236 = n7480 & n37235 ;
  assign n37237 = n21975 ^ n3485 ^ 1'b0 ;
  assign n37238 = n7596 & n34254 ;
  assign n37239 = n37238 ^ n14736 ^ 1'b0 ;
  assign n37240 = n23838 ^ n11252 ^ 1'b0 ;
  assign n37241 = ~n183 & n4419 ;
  assign n37242 = n10905 | n37241 ;
  assign n37243 = n6263 | n37242 ;
  assign n37244 = n18438 ^ n2185 ^ 1'b0 ;
  assign n37245 = n4607 ^ n507 ^ 1'b0 ;
  assign n37246 = n37244 & n37245 ;
  assign n37247 = n19475 ^ n4010 ^ 1'b0 ;
  assign n37248 = n32823 & n37247 ;
  assign n37249 = n22487 ^ n21958 ^ 1'b0 ;
  assign n37250 = n22273 ^ n9245 ^ 1'b0 ;
  assign n37251 = n4131 | n37250 ;
  assign n37252 = ~n18026 & n23438 ;
  assign n37253 = ~n3878 & n37252 ;
  assign n37254 = n22111 & ~n37253 ;
  assign n37255 = ~n7304 & n37254 ;
  assign n37256 = n22261 ^ n17021 ^ 1'b0 ;
  assign n37257 = n5169 & n37256 ;
  assign n37258 = n37257 ^ n7679 ^ 1'b0 ;
  assign n37259 = n7443 | n37258 ;
  assign n37260 = n21216 ^ n7384 ^ 1'b0 ;
  assign n37261 = n16762 | n37260 ;
  assign n37262 = n2446 | n13911 ;
  assign n37263 = n37261 & ~n37262 ;
  assign n37264 = n2073 | n9507 ;
  assign n37265 = n37264 ^ n4277 ^ 1'b0 ;
  assign n37266 = ( ~n6753 & n12364 ) | ( ~n6753 & n37265 ) | ( n12364 & n37265 ) ;
  assign n37267 = ( n6365 & n9311 ) | ( n6365 & n37266 ) | ( n9311 & n37266 ) ;
  assign n37268 = n30061 & ~n37267 ;
  assign n37269 = n11378 ^ n1693 ^ 1'b0 ;
  assign n37270 = n26346 ^ n10078 ^ 1'b0 ;
  assign n37271 = n12321 ^ n1246 ^ 1'b0 ;
  assign n37272 = ~n37270 & n37271 ;
  assign n37273 = n33777 ^ n25709 ^ 1'b0 ;
  assign n37274 = ~n1151 & n25385 ;
  assign n37275 = n36933 ^ n32192 ^ 1'b0 ;
  assign n37276 = n5101 | n37275 ;
  assign n37277 = n35893 ^ n15367 ^ 1'b0 ;
  assign n37278 = n3074 & n21257 ;
  assign n37279 = ~n8720 & n37278 ;
  assign n37280 = n649 & n37279 ;
  assign n37281 = n1523 | n9925 ;
  assign n37282 = ~n3267 & n37281 ;
  assign n37283 = n17581 | n37282 ;
  assign n37284 = ~n4436 & n20749 ;
  assign n37285 = n385 & ~n7501 ;
  assign n37286 = n37285 ^ n36558 ^ 1'b0 ;
  assign n37287 = n37286 ^ n2047 ^ 1'b0 ;
  assign n37288 = n24595 & ~n37287 ;
  assign n37289 = n101 | n4931 ;
  assign n37290 = n24890 ^ n323 ^ 1'b0 ;
  assign n37291 = ~n375 & n10014 ;
  assign n37292 = n228 & n11631 ;
  assign n37293 = ~n37291 & n37292 ;
  assign n37294 = ( n4307 & n35359 ) | ( n4307 & n37293 ) | ( n35359 & n37293 ) ;
  assign n37295 = n19621 & ~n37294 ;
  assign n37296 = n37290 & n37295 ;
  assign n37297 = n23023 ^ n16382 ^ 1'b0 ;
  assign n37298 = n4166 & n8430 ;
  assign n37299 = n1907 | n37298 ;
  assign n37300 = n310 & ~n14713 ;
  assign n37301 = n37300 ^ n14546 ^ 1'b0 ;
  assign n37302 = n31744 & ~n37301 ;
  assign n37303 = n3361 & n6515 ;
  assign n37304 = n37303 ^ n8226 ^ 1'b0 ;
  assign n37305 = n18789 & n28249 ;
  assign n37306 = n37304 & n37305 ;
  assign n37308 = n575 | n34123 ;
  assign n37307 = n19781 ^ n11905 ^ 1'b0 ;
  assign n37309 = n37308 ^ n37307 ^ 1'b0 ;
  assign n37310 = n6274 | n8665 ;
  assign n37311 = n6333 | n37310 ;
  assign n37312 = n5231 & n17248 ;
  assign n37313 = n24847 & n37312 ;
  assign n37314 = n6308 | n14734 ;
  assign n37315 = ~n472 & n3107 ;
  assign n37316 = ~n4353 & n37315 ;
  assign n37317 = n6590 & n8667 ;
  assign n37318 = n37316 & n37317 ;
  assign n37319 = n1645 & n21231 ;
  assign n37320 = n37319 ^ n11122 ^ 1'b0 ;
  assign n37321 = n37320 ^ n35799 ^ 1'b0 ;
  assign n37322 = n13634 | n37321 ;
  assign n37323 = n14184 ^ n7378 ^ 1'b0 ;
  assign n37324 = n675 | n15725 ;
  assign n37325 = n18004 ^ n12997 ^ 1'b0 ;
  assign n37326 = n37324 & ~n37325 ;
  assign n37327 = n28972 ^ n14488 ^ 1'b0 ;
  assign n37328 = n32763 ^ n26489 ^ 1'b0 ;
  assign n37329 = n12062 & ~n30922 ;
  assign n37330 = n26420 & n37329 ;
  assign n37331 = n6367 & n33923 ;
  assign n37332 = ~n4077 & n37331 ;
  assign n37333 = n7371 | n37332 ;
  assign n37334 = n37330 & ~n37333 ;
  assign n37335 = ~n3540 & n3645 ;
  assign n37336 = ~n3371 & n37335 ;
  assign n37337 = n8107 | n14935 ;
  assign n37338 = n310 & ~n37337 ;
  assign n37339 = n5064 ^ n300 ^ 1'b0 ;
  assign n37340 = n23475 | n27466 ;
  assign n37341 = n37340 ^ n8329 ^ 1'b0 ;
  assign n37342 = n17526 & ~n20514 ;
  assign n37343 = ~n47 & n37342 ;
  assign n37344 = ~n22413 & n25439 ;
  assign n37345 = n37344 ^ n11865 ^ 1'b0 ;
  assign n37346 = ~n8504 & n10594 ;
  assign n37347 = ~n37345 & n37346 ;
  assign n37348 = ~n28348 & n37347 ;
  assign n37349 = ~n31807 & n37348 ;
  assign n37350 = n8175 | n33233 ;
  assign n37351 = ~n339 & n7439 ;
  assign n37352 = n3917 | n6953 ;
  assign n37353 = n37352 ^ n6114 ^ 1'b0 ;
  assign n37354 = n2104 & n3597 ;
  assign n37355 = n8034 ^ n753 ^ 1'b0 ;
  assign n37356 = n19491 & ~n37355 ;
  assign n37357 = n20070 ^ n5914 ^ 1'b0 ;
  assign n37358 = n37357 ^ n8552 ^ 1'b0 ;
  assign n37359 = n11090 ^ n2101 ^ 1'b0 ;
  assign n37360 = n7259 ^ n1065 ^ 1'b0 ;
  assign n37361 = n37359 & n37360 ;
  assign n37362 = n9884 & n23965 ;
  assign n37363 = n1997 & ~n8132 ;
  assign n37364 = n37363 ^ n611 ^ 1'b0 ;
  assign n37365 = n508 | n6093 ;
  assign n37366 = n1845 & n6048 ;
  assign n37367 = n5445 | n37366 ;
  assign n37368 = n1672 | n12540 ;
  assign n37369 = n37368 ^ n3271 ^ 1'b0 ;
  assign n37370 = n37369 ^ n2269 ^ 1'b0 ;
  assign n37372 = n3007 & n18477 ;
  assign n37373 = ~n3974 & n37372 ;
  assign n37371 = n1771 | n8653 ;
  assign n37374 = n37373 ^ n37371 ^ n10824 ;
  assign n37375 = ~n9719 & n14143 ;
  assign n37376 = ~n28390 & n37375 ;
  assign n37377 = n3282 & ~n13167 ;
  assign n37378 = ~n3177 & n37377 ;
  assign n37381 = n1194 | n3260 ;
  assign n37379 = ( n5074 & ~n7369 ) | ( n5074 & n11515 ) | ( ~n7369 & n11515 ) ;
  assign n37380 = n31350 & ~n37379 ;
  assign n37382 = n37381 ^ n37380 ^ 1'b0 ;
  assign n37383 = n27712 ^ n25746 ^ 1'b0 ;
  assign n37384 = n30500 | n37383 ;
  assign n37385 = n10029 & n21820 ;
  assign n37386 = n26581 & n37385 ;
  assign n37387 = n20342 | n37386 ;
  assign n37388 = ~n6133 & n11267 ;
  assign n37389 = n5338 | n7596 ;
  assign n37390 = n37389 ^ n12088 ^ 1'b0 ;
  assign n37391 = n37390 ^ n36103 ^ 1'b0 ;
  assign n37392 = n10836 ^ n3162 ^ 1'b0 ;
  assign n37393 = ~n26761 & n37392 ;
  assign n37394 = n37393 ^ n1394 ^ 1'b0 ;
  assign n37395 = ~n4449 & n37394 ;
  assign n37396 = n37395 ^ n1467 ^ 1'b0 ;
  assign n37397 = n3108 | n3613 ;
  assign n37398 = n23317 ^ n4271 ^ 1'b0 ;
  assign n37399 = n22478 ^ n10709 ^ 1'b0 ;
  assign n37400 = n9752 & n37399 ;
  assign n37401 = n19 | n34944 ;
  assign n37402 = n24577 | n37401 ;
  assign n37403 = n12540 ^ n3941 ^ 1'b0 ;
  assign n37404 = n12396 | n37403 ;
  assign n37405 = n37404 ^ n13793 ^ 1'b0 ;
  assign n37406 = ~n9142 & n16742 ;
  assign n37407 = n37406 ^ n18899 ^ 1'b0 ;
  assign n37408 = ~n6228 & n37407 ;
  assign n37412 = n10578 | n25714 ;
  assign n37413 = n7744 & ~n37412 ;
  assign n37410 = n1976 ^ n227 ^ 1'b0 ;
  assign n37411 = n31837 | n37410 ;
  assign n37409 = ~n11827 & n32025 ;
  assign n37414 = n37413 ^ n37411 ^ n37409 ;
  assign n37415 = n7214 ^ n213 ^ 1'b0 ;
  assign n37416 = n23498 | n37415 ;
  assign n37419 = n346 & ~n2004 ;
  assign n37420 = n37419 ^ n3056 ^ 1'b0 ;
  assign n37421 = ~n5752 & n37420 ;
  assign n37417 = n12654 ^ n1165 ^ 1'b0 ;
  assign n37418 = n25137 | n37417 ;
  assign n37422 = n37421 ^ n37418 ^ 1'b0 ;
  assign n37423 = n3940 | n5697 ;
  assign n37424 = n279 & ~n33266 ;
  assign n37425 = n21321 & n37424 ;
  assign n37426 = n37425 ^ n23066 ^ n8705 ;
  assign n37427 = n37426 ^ n9851 ^ 1'b0 ;
  assign n37428 = ~n37423 & n37427 ;
  assign n37429 = n2929 | n17111 ;
  assign n37430 = n8284 ^ n6157 ^ 1'b0 ;
  assign n37431 = ~n37429 & n37430 ;
  assign n37432 = n37431 ^ n33629 ^ 1'b0 ;
  assign n37433 = ~n14760 & n37432 ;
  assign n37434 = n26740 & n37433 ;
  assign n37435 = n35360 ^ n35023 ^ 1'b0 ;
  assign n37436 = ~n4163 & n31051 ;
  assign n37437 = n4668 | n8848 ;
  assign n37438 = n3061 & n37437 ;
  assign n37439 = n1287 & ~n20272 ;
  assign n37440 = n37439 ^ n34759 ^ 1'b0 ;
  assign n37441 = n6865 & n20698 ;
  assign n37442 = n20334 & ~n37441 ;
  assign n37443 = n37442 ^ n10650 ^ 1'b0 ;
  assign n37444 = n1924 & ~n37443 ;
  assign n37445 = n5732 | n12492 ;
  assign n37446 = n37445 ^ n1373 ^ 1'b0 ;
  assign n37447 = n26741 ^ n16568 ^ 1'b0 ;
  assign n37448 = n18039 | n37447 ;
  assign n37449 = n4319 ^ n1396 ^ 1'b0 ;
  assign n37450 = n6001 & n10435 ;
  assign n37451 = ~n10435 & n37450 ;
  assign n37452 = ~n5706 & n9088 ;
  assign n37453 = n1358 & n25302 ;
  assign n37454 = n4036 ^ n3162 ^ 1'b0 ;
  assign n37455 = n37453 & ~n37454 ;
  assign n37456 = n5092 | n7779 ;
  assign n37457 = n34950 ^ n13974 ^ 1'b0 ;
  assign n37458 = n1350 | n20541 ;
  assign n37460 = n9175 ^ n1263 ^ 1'b0 ;
  assign n37461 = n1118 | n37460 ;
  assign n37459 = n1250 & n10729 ;
  assign n37462 = n37461 ^ n37459 ^ 1'b0 ;
  assign n37463 = n37462 ^ n25195 ^ 1'b0 ;
  assign n37464 = n2695 & n13717 ;
  assign n37465 = n17316 ^ n6755 ^ 1'b0 ;
  assign n37466 = n4284 & n37465 ;
  assign n37467 = n83 & ~n9201 ;
  assign n37468 = n18463 ^ n7440 ^ 1'b0 ;
  assign n37469 = ~n21658 & n37468 ;
  assign n37470 = ~n12734 & n33995 ;
  assign n37471 = n8993 & n14159 ;
  assign n37472 = n37471 ^ n3722 ^ 1'b0 ;
  assign n37473 = n12457 | n37270 ;
  assign n37474 = n37472 & ~n37473 ;
  assign n37475 = n32537 | n37474 ;
  assign n37476 = n37475 ^ n35519 ^ 1'b0 ;
  assign n37478 = n2410 ^ n1785 ^ 1'b0 ;
  assign n37479 = n4568 ^ n4219 ^ 1'b0 ;
  assign n37480 = n37478 & ~n37479 ;
  assign n37481 = ~n1828 & n7030 ;
  assign n37482 = ~n37480 & n37481 ;
  assign n37477 = n11521 & n16491 ;
  assign n37483 = n37482 ^ n37477 ^ 1'b0 ;
  assign n37484 = n7353 ^ n2788 ^ 1'b0 ;
  assign n37485 = n37484 ^ n8317 ^ n1257 ;
  assign n37486 = ~n4676 & n9586 ;
  assign n37487 = n20618 & ~n24376 ;
  assign n37488 = n20838 ^ n1632 ^ 1'b0 ;
  assign n37489 = ~n37487 & n37488 ;
  assign n37491 = n4993 ^ n3369 ^ 1'b0 ;
  assign n37490 = n20902 & ~n35944 ;
  assign n37492 = n37491 ^ n37490 ^ 1'b0 ;
  assign n37493 = n36010 & ~n37492 ;
  assign n37494 = n1754 | n14789 ;
  assign n37495 = n15081 ^ n7860 ^ 1'b0 ;
  assign n37496 = ~n798 & n9667 ;
  assign n37497 = n13251 & n37496 ;
  assign n37498 = n28610 ^ n21944 ^ 1'b0 ;
  assign n37499 = n11643 & n37498 ;
  assign n37500 = n37497 & n37499 ;
  assign n37501 = n37500 ^ n29242 ^ 1'b0 ;
  assign n37502 = n15408 & ~n19744 ;
  assign n37503 = n37502 ^ n11229 ^ 1'b0 ;
  assign n37504 = n8262 ^ n3077 ^ 1'b0 ;
  assign n37505 = ~n4311 & n37504 ;
  assign n37506 = n37505 ^ n3890 ^ 1'b0 ;
  assign n37507 = n37503 & n37506 ;
  assign n37508 = n37507 ^ n8206 ^ 1'b0 ;
  assign n37509 = n22961 ^ n20837 ^ 1'b0 ;
  assign n37510 = n4193 & ~n37509 ;
  assign n37511 = ~n18201 & n37510 ;
  assign n37512 = n37511 ^ n21534 ^ 1'b0 ;
  assign n37513 = ~n113 & n7612 ;
  assign n37514 = ~n4246 & n37513 ;
  assign n37515 = n11554 ^ n4984 ^ 1'b0 ;
  assign n37516 = ~n21360 & n37515 ;
  assign n37517 = n6184 ^ n120 ^ 1'b0 ;
  assign n37518 = n34612 & n37517 ;
  assign n37519 = n18847 & n37518 ;
  assign n37522 = n1802 & ~n14416 ;
  assign n37523 = ~n4700 & n37522 ;
  assign n37520 = n6256 | n36150 ;
  assign n37521 = n10286 & ~n37520 ;
  assign n37524 = n37523 ^ n37521 ^ 1'b0 ;
  assign n37525 = n37524 ^ n2090 ^ 1'b0 ;
  assign n37526 = n4247 & ~n10930 ;
  assign n37527 = n37526 ^ n19138 ^ 1'b0 ;
  assign n37528 = n21424 ^ n4473 ^ 1'b0 ;
  assign n37529 = n18093 ^ n34 ^ 1'b0 ;
  assign n37530 = n1227 & ~n37529 ;
  assign n37531 = n36314 ^ n19779 ^ n11606 ;
  assign n37532 = ~n10992 & n11535 ;
  assign n37533 = n37531 & n37532 ;
  assign n37534 = n31744 ^ n20301 ^ 1'b0 ;
  assign n37535 = n427 | n11076 ;
  assign n37536 = n11698 & n18468 ;
  assign n37537 = n995 & n37536 ;
  assign n37538 = n25137 & n37537 ;
  assign n37539 = ( n6524 & n11758 ) | ( n6524 & ~n21468 ) | ( n11758 & ~n21468 ) ;
  assign n37540 = n10785 & n37539 ;
  assign n37541 = ~n19776 & n37540 ;
  assign n37542 = n14824 ^ n11626 ^ 1'b0 ;
  assign n37543 = n4638 & n15763 ;
  assign n37544 = n37543 ^ n21481 ^ 1'b0 ;
  assign n37545 = n13719 ^ n6907 ^ 1'b0 ;
  assign n37546 = n406 & n37545 ;
  assign n37547 = ~n22135 & n37089 ;
  assign n37548 = n6281 & n19389 ;
  assign n37549 = n1167 & n37548 ;
  assign n37550 = n18462 & n27009 ;
  assign n37551 = n7594 | n33161 ;
  assign n37552 = n37551 ^ n14474 ^ 1'b0 ;
  assign n37553 = ~n14316 & n37552 ;
  assign n37554 = n37553 ^ n3301 ^ 1'b0 ;
  assign n37555 = n13700 ^ n4428 ^ 1'b0 ;
  assign n37558 = n7594 & n16124 ;
  assign n37556 = n9208 & n10427 ;
  assign n37557 = n1344 & ~n37556 ;
  assign n37559 = n37558 ^ n37557 ^ 1'b0 ;
  assign n37560 = n28300 ^ n24561 ^ 1'b0 ;
  assign n37562 = n3981 & ~n20782 ;
  assign n37561 = n8409 & n10736 ;
  assign n37563 = n37562 ^ n37561 ^ 1'b0 ;
  assign n37564 = ~n13846 & n37563 ;
  assign n37565 = n37564 ^ n18102 ^ 1'b0 ;
  assign n37566 = n2148 | n14316 ;
  assign n37567 = n37566 ^ n16749 ^ 1'b0 ;
  assign n37568 = n7487 & ~n29690 ;
  assign n37569 = n34913 | n36437 ;
  assign n37570 = n3211 & ~n37569 ;
  assign n37571 = n24655 ^ n10021 ^ 1'b0 ;
  assign n37572 = n632 | n6209 ;
  assign n37573 = n19720 ^ n3295 ^ 1'b0 ;
  assign n37574 = n4216 | n15288 ;
  assign n37575 = n37574 ^ n13389 ^ 1'b0 ;
  assign n37576 = n3125 & n37575 ;
  assign n37577 = ~n1205 & n7056 ;
  assign n37578 = n564 & n18761 ;
  assign n37579 = n37578 ^ n3640 ^ 1'b0 ;
  assign n37580 = n37577 & ~n37579 ;
  assign n37581 = n653 & n949 ;
  assign n37582 = ~n2439 & n37581 ;
  assign n37583 = n2159 & ~n37582 ;
  assign n37584 = n3826 | n15637 ;
  assign n37585 = n36876 & n37584 ;
  assign n37586 = n627 & n1790 ;
  assign n37587 = n37586 ^ n24326 ^ n22727 ;
  assign n37588 = ~n2318 & n5369 ;
  assign n37589 = n1771 | n37588 ;
  assign n37590 = n20101 & n23894 ;
  assign n37591 = n37590 ^ n7352 ^ 1'b0 ;
  assign n37592 = n32774 & ~n37591 ;
  assign n37593 = n9478 ^ n259 ^ 1'b0 ;
  assign n37594 = n28268 & ~n37593 ;
  assign n37595 = n24146 & n37594 ;
  assign n37597 = n20829 | n23262 ;
  assign n37596 = n1885 & ~n2011 ;
  assign n37598 = n37597 ^ n37596 ^ 1'b0 ;
  assign n37599 = n3992 & n7650 ;
  assign n37600 = n37599 ^ n30078 ^ 1'b0 ;
  assign n37601 = n9491 & ~n30098 ;
  assign n37602 = n37601 ^ n4358 ^ 1'b0 ;
  assign n37603 = n2012 & n26944 ;
  assign n37604 = n3465 & n15761 ;
  assign n37605 = ~n22790 & n37604 ;
  assign n37606 = ~n33477 & n33816 ;
  assign n37607 = n6021 ^ n2029 ^ 1'b0 ;
  assign n37608 = n34162 ^ n31973 ^ 1'b0 ;
  assign n37609 = ~n17263 & n19626 ;
  assign n37610 = n37609 ^ n4609 ^ 1'b0 ;
  assign n37611 = n13972 ^ n477 ^ 1'b0 ;
  assign n37612 = ~n14901 & n37611 ;
  assign n37613 = n3877 & ~n6543 ;
  assign n37614 = n12363 ^ n9883 ^ 1'b0 ;
  assign n37615 = n4133 & n33060 ;
  assign n37616 = n37615 ^ n23139 ^ 1'b0 ;
  assign n37619 = n20409 & ~n25091 ;
  assign n37617 = ~n21653 & n29722 ;
  assign n37618 = n37617 ^ n22338 ^ 1'b0 ;
  assign n37620 = n37619 ^ n37618 ^ n37357 ;
  assign n37621 = n26611 ^ n3679 ^ 1'b0 ;
  assign n37623 = n323 & n8517 ;
  assign n37624 = n37623 ^ n21759 ^ 1'b0 ;
  assign n37622 = n9695 | n13165 ;
  assign n37625 = n37624 ^ n37622 ^ 1'b0 ;
  assign n37626 = n10600 | n15294 ;
  assign n37627 = n37625 | n37626 ;
  assign n37628 = n3592 & n5806 ;
  assign n37629 = n9463 | n37628 ;
  assign n37630 = n6028 | n37629 ;
  assign n37631 = n37112 | n37630 ;
  assign n37632 = n339 & n21276 ;
  assign n37635 = n14464 & n35467 ;
  assign n37633 = n2205 & n7334 ;
  assign n37634 = n37633 ^ n14558 ^ 1'b0 ;
  assign n37636 = n37635 ^ n37634 ^ 1'b0 ;
  assign n37637 = ~n2872 & n7593 ;
  assign n37638 = n7003 & n37637 ;
  assign n37639 = n486 & n5752 ;
  assign n37640 = n37639 ^ n7863 ^ 1'b0 ;
  assign n37641 = n4956 & ~n27156 ;
  assign n37642 = n25385 ^ n18123 ^ 1'b0 ;
  assign n37643 = ~n2984 & n13206 ;
  assign n37644 = n10824 ^ n2542 ^ 1'b0 ;
  assign n37645 = ( n12489 & ~n37643 ) | ( n12489 & n37644 ) | ( ~n37643 & n37644 ) ;
  assign n37646 = n24649 ^ n19792 ^ n534 ;
  assign n37647 = n1681 ^ n836 ^ 1'b0 ;
  assign n37648 = n21506 & n32083 ;
  assign n37649 = ~n14175 & n37648 ;
  assign n37650 = n6919 ^ n5011 ^ 1'b0 ;
  assign n37651 = n4469 & ~n11405 ;
  assign n37652 = n37651 ^ n1957 ^ 1'b0 ;
  assign n37653 = n37652 ^ n3447 ^ 1'b0 ;
  assign n37654 = n37650 | n37653 ;
  assign n37655 = ~n25719 & n37654 ;
  assign n37656 = n18001 ^ n630 ^ 1'b0 ;
  assign n37657 = n23349 & n37656 ;
  assign n37658 = n27067 ^ n10249 ^ 1'b0 ;
  assign n37659 = n302 & ~n5913 ;
  assign n37660 = n3774 ^ n799 ^ 1'b0 ;
  assign n37661 = n27220 & ~n37660 ;
  assign n37662 = n423 & n34313 ;
  assign n37663 = n37662 ^ n20486 ^ 1'b0 ;
  assign n37664 = n37663 ^ n5367 ^ 1'b0 ;
  assign n37665 = n13981 | n37664 ;
  assign n37666 = n19138 ^ n6986 ^ 1'b0 ;
  assign n37667 = n37666 ^ n6397 ^ 1'b0 ;
  assign n37668 = n16011 | n19825 ;
  assign n37669 = ~n3594 & n15117 ;
  assign n37670 = ~n3516 & n14678 ;
  assign n37671 = n4811 | n8108 ;
  assign n37672 = n37671 ^ n5532 ^ 1'b0 ;
  assign n37673 = n29039 ^ n5308 ^ 1'b0 ;
  assign n37674 = n37672 & ~n37673 ;
  assign n37675 = n8263 & n37674 ;
  assign n37676 = n2884 | n31907 ;
  assign n37678 = n11771 ^ n8156 ^ 1'b0 ;
  assign n37679 = n7477 | n37678 ;
  assign n37677 = n2759 ^ n1081 ^ 1'b0 ;
  assign n37680 = n37679 ^ n37677 ^ 1'b0 ;
  assign n37681 = ~n11619 & n14645 ;
  assign n37682 = n27725 ^ n8197 ^ 1'b0 ;
  assign n37683 = n37681 & n37682 ;
  assign n37684 = n22990 ^ n1802 ^ 1'b0 ;
  assign n37685 = n216 | n963 ;
  assign n37686 = n4904 ^ n1328 ^ 1'b0 ;
  assign n37687 = n9126 & n37686 ;
  assign n37688 = n20149 & n37687 ;
  assign n37689 = n37688 ^ n17959 ^ 1'b0 ;
  assign n37690 = n37689 ^ n21077 ^ n62 ;
  assign n37691 = n7229 & n25095 ;
  assign n37692 = n37691 ^ n11409 ^ 1'b0 ;
  assign n37693 = n22472 ^ n14696 ^ 1'b0 ;
  assign n37694 = ( ~n2660 & n10611 ) | ( ~n2660 & n22213 ) | ( n10611 & n22213 ) ;
  assign n37695 = n37694 ^ n32403 ^ 1'b0 ;
  assign n37696 = ~n14483 & n37695 ;
  assign n37697 = n20496 ^ n12178 ^ 1'b0 ;
  assign n37698 = n5174 & n11585 ;
  assign n37699 = n12665 | n23794 ;
  assign n37700 = n3194 | n37699 ;
  assign n37701 = ~n2973 & n5747 ;
  assign n37702 = n477 & ~n2627 ;
  assign n37703 = n4280 & ~n7263 ;
  assign n37704 = n37703 ^ n12171 ^ 1'b0 ;
  assign n37705 = n2067 & ~n37704 ;
  assign n37706 = n37702 & n37705 ;
  assign n37707 = n23948 ^ n11624 ^ 1'b0 ;
  assign n37708 = n12172 & ~n24069 ;
  assign n37709 = n12019 ^ n5193 ^ 1'b0 ;
  assign n37710 = ~n1763 & n37709 ;
  assign n37711 = ~n33823 & n37710 ;
  assign n37712 = ~n37708 & n37711 ;
  assign n37713 = ( n2008 & ~n3679 ) | ( n2008 & n14411 ) | ( ~n3679 & n14411 ) ;
  assign n37714 = n4109 & n4193 ;
  assign n37715 = ~n37713 & n37714 ;
  assign n37716 = n19073 ^ n9880 ^ 1'b0 ;
  assign n37717 = n32061 ^ n1329 ^ 1'b0 ;
  assign n37718 = n10877 ^ n938 ^ 1'b0 ;
  assign n37719 = n20330 & ~n37718 ;
  assign n37720 = ~n5465 & n6775 ;
  assign n37721 = n17386 ^ n4581 ^ 1'b0 ;
  assign n37722 = n20846 & n37721 ;
  assign n37723 = ~n5926 & n37722 ;
  assign n37724 = n11409 & n14544 ;
  assign n37725 = n37724 ^ n25633 ^ 1'b0 ;
  assign n37726 = n16271 ^ n5556 ^ 1'b0 ;
  assign n37727 = n11129 ^ n1249 ^ 1'b0 ;
  assign n37728 = n25831 ^ n21219 ^ 1'b0 ;
  assign n37729 = ~n8508 & n9544 ;
  assign n37730 = ~n5111 & n18650 ;
  assign n37731 = ( n10363 & n14109 ) | ( n10363 & n18387 ) | ( n14109 & n18387 ) ;
  assign n37732 = n9770 & ~n25029 ;
  assign n37733 = n9074 & n37732 ;
  assign n37734 = n540 ^ n68 ^ 1'b0 ;
  assign n37735 = n29027 & n37734 ;
  assign n37736 = n37733 & n37735 ;
  assign n37737 = n23035 ^ n2785 ^ 1'b0 ;
  assign n37738 = n37736 | n37737 ;
  assign n37739 = n6361 | n30415 ;
  assign n37740 = n33733 | n37739 ;
  assign n37741 = n3981 & ~n26966 ;
  assign n37742 = n2266 & ~n2789 ;
  assign n37743 = n37742 ^ n19 ^ 1'b0 ;
  assign n37744 = n928 | n24972 ;
  assign n37745 = n4590 & ~n19540 ;
  assign n37746 = n25803 & n37745 ;
  assign n37747 = n1995 & ~n6960 ;
  assign n37748 = n2439 & n23841 ;
  assign n37749 = n37748 ^ n6608 ^ 1'b0 ;
  assign n37750 = n37749 ^ n22219 ^ 1'b0 ;
  assign n37751 = n37747 | n37750 ;
  assign n37755 = ~n2684 & n3456 ;
  assign n37756 = ~n3456 & n37755 ;
  assign n37757 = n4019 & ~n37756 ;
  assign n37758 = ~n4019 & n37757 ;
  assign n37759 = n15739 & ~n37758 ;
  assign n37760 = n5021 & n37759 ;
  assign n37752 = n1664 & ~n34342 ;
  assign n37753 = ~n1664 & n37752 ;
  assign n37754 = n5957 | n37753 ;
  assign n37761 = n37760 ^ n37754 ^ 1'b0 ;
  assign n37762 = n2483 | n37761 ;
  assign n37763 = n37762 ^ n11286 ^ 1'b0 ;
  assign n37764 = n19826 ^ n8031 ^ 1'b0 ;
  assign n37765 = ~n19359 & n37764 ;
  assign n37766 = n17016 ^ n4273 ^ 1'b0 ;
  assign n37768 = ~n13997 & n16124 ;
  assign n37769 = n7744 | n37768 ;
  assign n37767 = n251 & n1852 ;
  assign n37770 = n37769 ^ n37767 ^ 1'b0 ;
  assign n37771 = n27198 ^ n9918 ^ 1'b0 ;
  assign n37772 = n15261 & ~n20480 ;
  assign n37773 = n2792 & n37772 ;
  assign n37774 = n34576 | n37773 ;
  assign n37775 = ~n8079 & n31654 ;
  assign n37777 = n440 | n7744 ;
  assign n37778 = n32927 | n37777 ;
  assign n37776 = n1210 & n13326 ;
  assign n37779 = n37778 ^ n37776 ^ 1'b0 ;
  assign n37780 = n879 & n25867 ;
  assign n37781 = n3676 & n4097 ;
  assign n37783 = n8532 ^ n2967 ^ 1'b0 ;
  assign n37782 = ~n16741 & n21111 ;
  assign n37784 = n37783 ^ n37782 ^ 1'b0 ;
  assign n37785 = n6102 ^ n3231 ^ 1'b0 ;
  assign n37786 = n13165 | n37785 ;
  assign n37787 = n666 | n37786 ;
  assign n37788 = n15273 ^ n12354 ^ 1'b0 ;
  assign n37789 = n37787 & n37788 ;
  assign n37790 = n6174 | n8713 ;
  assign n37791 = n37790 ^ n3990 ^ 1'b0 ;
  assign n37792 = n37791 ^ n30842 ^ 1'b0 ;
  assign n37793 = n8014 & n33246 ;
  assign n37794 = n4034 & n22491 ;
  assign n37795 = n6157 ^ n2476 ^ 1'b0 ;
  assign n37796 = n1834 & ~n37795 ;
  assign n37797 = n37796 ^ n24204 ^ 1'b0 ;
  assign n37798 = n129 & ~n10470 ;
  assign n37799 = n37798 ^ n16956 ^ 1'b0 ;
  assign n37800 = n1968 ^ n226 ^ 1'b0 ;
  assign n37801 = n13537 & n13679 ;
  assign n37802 = ~n1086 & n37801 ;
  assign n37803 = n24838 ^ n6776 ^ 1'b0 ;
  assign n37804 = n16660 ^ n9574 ^ n8876 ;
  assign n37805 = n16465 | n37804 ;
  assign n37806 = n30192 & ~n37805 ;
  assign n37807 = n37806 ^ n35763 ^ 1'b0 ;
  assign n37808 = n15694 | n23624 ;
  assign n37809 = n28283 & ~n37808 ;
  assign n37810 = ~n18282 & n27145 ;
  assign n37811 = n29080 & n37810 ;
  assign n37812 = n2047 & ~n5923 ;
  assign n37813 = n37812 ^ n10421 ^ 1'b0 ;
  assign n37814 = n28942 ^ n2859 ^ 1'b0 ;
  assign n37815 = ~n34094 & n37814 ;
  assign n37816 = n5950 & ~n37815 ;
  assign n37817 = n33920 ^ n17999 ^ 1'b0 ;
  assign n37818 = n12657 & n19946 ;
  assign n37819 = n37818 ^ n175 ^ 1'b0 ;
  assign n37820 = n29342 & n37819 ;
  assign n37821 = n37820 ^ n2936 ^ 1'b0 ;
  assign n37822 = n3584 & ~n37821 ;
  assign n37823 = n2403 & n37822 ;
  assign n37824 = ~n4532 & n8624 ;
  assign n37825 = n7662 & n25382 ;
  assign n37826 = n11702 | n37332 ;
  assign n37827 = n37826 ^ n1945 ^ 1'b0 ;
  assign n37828 = n8518 | n14991 ;
  assign n37829 = n8479 & ~n37828 ;
  assign n37830 = n20004 | n37829 ;
  assign n37831 = n11859 | n21943 ;
  assign n37832 = n3965 & n15792 ;
  assign n37833 = n26461 & n37832 ;
  assign n37834 = n37833 ^ n673 ^ 1'b0 ;
  assign n37835 = n37831 | n37834 ;
  assign n37836 = n23177 ^ n817 ^ 1'b0 ;
  assign n37837 = n19414 ^ n14325 ^ 1'b0 ;
  assign n37838 = n37836 & ~n37837 ;
  assign n37839 = n1721 & ~n27580 ;
  assign n37840 = ~n26048 & n37839 ;
  assign n37841 = n24403 ^ n9873 ^ 1'b0 ;
  assign n37842 = n1358 & n10374 ;
  assign n37843 = n13478 & ~n15191 ;
  assign n37844 = n29022 ^ n592 ^ 1'b0 ;
  assign n37845 = n599 & n624 ;
  assign n37846 = n30163 ^ n21464 ^ 1'b0 ;
  assign n37847 = n6135 ^ n185 ^ 1'b0 ;
  assign n37848 = n20667 | n37847 ;
  assign n37850 = n2835 | n14321 ;
  assign n37851 = n17445 | n37850 ;
  assign n37849 = n20808 ^ n15668 ^ 1'b0 ;
  assign n37852 = n37851 ^ n37849 ^ n3846 ;
  assign n37853 = n22966 ^ n18937 ^ 1'b0 ;
  assign n37854 = n6849 & ~n37853 ;
  assign n37855 = n1577 & n8624 ;
  assign n37856 = n37855 ^ n7330 ^ 1'b0 ;
  assign n37857 = n37856 ^ n13536 ^ 1'b0 ;
  assign n37859 = n5522 | n11674 ;
  assign n37858 = ~n5942 & n26313 ;
  assign n37860 = n37859 ^ n37858 ^ 1'b0 ;
  assign n37861 = n33699 ^ n12125 ^ n1492 ;
  assign n37863 = n13163 & n23306 ;
  assign n37862 = n12238 ^ n10018 ^ 1'b0 ;
  assign n37864 = n37863 ^ n37862 ^ n36662 ;
  assign n37865 = n79 & ~n19867 ;
  assign n37866 = n37865 ^ n17695 ^ 1'b0 ;
  assign n37867 = n253 & n10184 ;
  assign n37868 = n11447 & ~n37867 ;
  assign n37869 = n6644 & n28297 ;
  assign n37870 = n467 | n512 ;
  assign n37871 = n5554 & n14329 ;
  assign n37872 = n37871 ^ n5124 ^ 1'b0 ;
  assign n37873 = n2808 | n37872 ;
  assign n37875 = ~n11624 & n14128 ;
  assign n37876 = n16617 & n37875 ;
  assign n37874 = n169 | n25110 ;
  assign n37877 = n37876 ^ n37874 ^ 1'b0 ;
  assign n37878 = n2460 ^ n973 ^ n895 ;
  assign n37879 = n1802 & ~n14552 ;
  assign n37880 = n37879 ^ n8627 ^ 1'b0 ;
  assign n37881 = n22947 & n37880 ;
  assign n37882 = n22686 ^ n13238 ^ 1'b0 ;
  assign n37883 = n12685 | n37882 ;
  assign n37884 = n2542 ^ n257 ^ 1'b0 ;
  assign n37885 = n16288 & n37884 ;
  assign n37886 = n37885 ^ n4074 ^ 1'b0 ;
  assign n37887 = n37886 ^ n31946 ^ 1'b0 ;
  assign n37888 = ~n5794 & n13293 ;
  assign n37889 = n37888 ^ n1533 ^ 1'b0 ;
  assign n37890 = n6039 & ~n37889 ;
  assign n37891 = n558 & n37890 ;
  assign n37892 = n11653 ^ n2826 ^ 1'b0 ;
  assign n37893 = n32535 ^ n6162 ^ 1'b0 ;
  assign n37894 = ~n4531 & n10837 ;
  assign n37896 = ~n6892 & n10897 ;
  assign n37895 = n642 | n26924 ;
  assign n37897 = n37896 ^ n37895 ^ n929 ;
  assign n37898 = n33911 ^ n8092 ^ 1'b0 ;
  assign n37899 = ~n4465 & n10855 ;
  assign n37900 = n37899 ^ x0 ^ 1'b0 ;
  assign n37901 = n14164 ^ n2282 ^ 1'b0 ;
  assign n37902 = n2070 | n37901 ;
  assign n37903 = n37902 ^ n19546 ^ 1'b0 ;
  assign n37904 = ( n2800 & n13872 ) | ( n2800 & n33912 ) | ( n13872 & n33912 ) ;
  assign n37905 = n10833 & n37904 ;
  assign n37906 = ~n37903 & n37905 ;
  assign n37907 = n2316 | n16109 ;
  assign n37908 = n35373 & n36273 ;
  assign n37909 = n20111 ^ n2535 ^ 1'b0 ;
  assign n37910 = n3593 ^ n56 ^ 1'b0 ;
  assign n37911 = ~n21594 & n37910 ;
  assign n37912 = ~n1695 & n10383 ;
  assign n37913 = n34631 ^ n15631 ^ n13685 ;
  assign n37914 = n26287 ^ n3088 ^ 1'b0 ;
  assign n37915 = n7701 & ~n37914 ;
  assign n37916 = n2348 | n11931 ;
  assign n37917 = ~n1598 & n37916 ;
  assign n37918 = n30255 ^ n23024 ^ 1'b0 ;
  assign n37919 = n8543 | n37918 ;
  assign n37920 = n10740 ^ n8677 ^ 1'b0 ;
  assign n37921 = n34263 ^ n12482 ^ 1'b0 ;
  assign n37922 = n37920 | n37921 ;
  assign n37923 = n37922 ^ n25043 ^ 1'b0 ;
  assign n37925 = n200 & ~n6611 ;
  assign n37924 = ~n7179 & n11703 ;
  assign n37926 = n37925 ^ n37924 ^ 1'b0 ;
  assign n37927 = n20131 ^ n7675 ^ n1403 ;
  assign n37928 = n37927 ^ n34567 ^ n29859 ;
  assign n37929 = n4202 & n8613 ;
  assign n37930 = n24938 ^ n5513 ^ n1895 ;
  assign n37931 = n8864 ^ n1945 ^ 1'b0 ;
  assign n37932 = n14177 ^ n2155 ^ 1'b0 ;
  assign n37933 = n24024 & n37932 ;
  assign n37934 = n37931 & n37933 ;
  assign n37937 = ~n10934 & n13730 ;
  assign n37935 = n3167 ^ n581 ^ 1'b0 ;
  assign n37936 = n8984 | n37935 ;
  assign n37938 = n37937 ^ n37936 ^ 1'b0 ;
  assign n37939 = n32204 & ~n37938 ;
  assign n37940 = n37939 ^ n31162 ^ 1'b0 ;
  assign n37941 = ~n567 & n6335 ;
  assign n37942 = n6732 | n10284 ;
  assign n37943 = n37941 | n37942 ;
  assign n37944 = ( n11071 & n24256 ) | ( n11071 & n37049 ) | ( n24256 & n37049 ) ;
  assign n37945 = n14088 & ~n37944 ;
  assign n37946 = n12000 ^ n2545 ^ 1'b0 ;
  assign n37947 = n32550 ^ n27377 ^ 1'b0 ;
  assign n37948 = ~n20507 & n37947 ;
  assign n37949 = n12563 ^ n1048 ^ 1'b0 ;
  assign n37950 = n29476 ^ n4022 ^ 1'b0 ;
  assign n37951 = n2205 & ~n37950 ;
  assign n37952 = n30636 ^ n807 ^ 1'b0 ;
  assign n37953 = n15543 | n37952 ;
  assign n37954 = n1693 | n37953 ;
  assign n37955 = n37951 | n37954 ;
  assign n37956 = n15646 & n26735 ;
  assign n37957 = n4913 & ~n37956 ;
  assign n37958 = n3559 & n37957 ;
  assign n37959 = n31147 ^ n13985 ^ n2807 ;
  assign n37960 = ~n8142 & n20131 ;
  assign n37961 = n35256 ^ n6617 ^ 1'b0 ;
  assign n37962 = ~n2843 & n37961 ;
  assign n37963 = n15109 & n37962 ;
  assign n37964 = n6197 | n37963 ;
  assign n37965 = n37964 ^ n2214 ^ 1'b0 ;
  assign n37966 = n11098 | n12034 ;
  assign n37967 = n25824 ^ n21227 ^ 1'b0 ;
  assign n37968 = n37966 & ~n37967 ;
  assign n37969 = n3227 | n5158 ;
  assign n37970 = ~n11826 & n37969 ;
  assign n37971 = ~n16607 & n37970 ;
  assign n37972 = n8817 & ~n15901 ;
  assign n37973 = n9659 & ~n21392 ;
  assign n37974 = n37973 ^ n32771 ^ 1'b0 ;
  assign n37975 = n28942 ^ n21521 ^ 1'b0 ;
  assign n37976 = n1435 & ~n37975 ;
  assign n37977 = n3260 | n28134 ;
  assign n37992 = ~n180 & n1166 ;
  assign n37993 = n180 & n37992 ;
  assign n37978 = n37 & ~n397 ;
  assign n37979 = n16 & ~n37978 ;
  assign n37980 = n12620 | n30359 ;
  assign n37981 = n30359 & ~n37980 ;
  assign n37982 = n119 | n37981 ;
  assign n37983 = n119 & ~n37982 ;
  assign n37984 = n37979 & ~n37983 ;
  assign n37985 = ~n37979 & n37984 ;
  assign n37986 = n18165 | n37985 ;
  assign n37987 = n18165 & ~n37986 ;
  assign n37988 = n216 & n2634 ;
  assign n37989 = ~n2634 & n37988 ;
  assign n37990 = n37989 ^ n1441 ^ 1'b0 ;
  assign n37991 = n37987 | n37990 ;
  assign n37994 = n37993 ^ n37991 ^ 1'b0 ;
  assign n37995 = n321 & ~n37994 ;
  assign n37996 = ~n3122 & n32143 ;
  assign n37997 = n6874 & ~n15582 ;
  assign n37998 = ~n3653 & n37997 ;
  assign n37999 = n31492 & n37998 ;
  assign n38000 = n19117 & n34294 ;
  assign n38001 = n3663 ^ n168 ^ 1'b0 ;
  assign n38002 = n34 & ~n38001 ;
  assign n38003 = ~n9521 & n38002 ;
  assign n38004 = n38003 ^ n11319 ^ 1'b0 ;
  assign n38005 = n16226 ^ n12743 ^ 1'b0 ;
  assign n38006 = ~n4594 & n11629 ;
  assign n38007 = n2826 | n6297 ;
  assign n38008 = ( ~n8473 & n25104 ) | ( ~n8473 & n38007 ) | ( n25104 & n38007 ) ;
  assign n38009 = n11643 & ~n38008 ;
  assign n38010 = n38006 & n38009 ;
  assign n38011 = n1593 & ~n10014 ;
  assign n38012 = n38011 ^ n1154 ^ 1'b0 ;
  assign n38013 = ~n6940 & n23166 ;
  assign n38014 = ~n38012 & n38013 ;
  assign n38015 = n19633 & n38014 ;
  assign n38016 = n4314 & n27435 ;
  assign n38017 = n3177 | n38016 ;
  assign n38018 = n5914 & ~n20555 ;
  assign n38019 = n38018 ^ n7321 ^ 1'b0 ;
  assign n38021 = n9337 ^ n5237 ^ 1'b0 ;
  assign n38020 = ~n9134 & n10785 ;
  assign n38022 = n38021 ^ n38020 ^ 1'b0 ;
  assign n38023 = n28049 | n30551 ;
  assign n38024 = n17395 ^ n13979 ^ 1'b0 ;
  assign n38025 = n14055 & ~n38024 ;
  assign n38026 = n9011 | n25108 ;
  assign n38027 = n38026 ^ n9434 ^ n1565 ;
  assign n38028 = ~n11893 & n22461 ;
  assign n38030 = n18333 ^ n2441 ^ 1'b0 ;
  assign n38029 = ~n8969 & n9890 ;
  assign n38031 = n38030 ^ n38029 ^ 1'b0 ;
  assign n38032 = n3452 | n38031 ;
  assign n38033 = n38032 ^ n23390 ^ 1'b0 ;
  assign n38034 = n9474 & n37611 ;
  assign n38035 = n38034 ^ n12934 ^ 1'b0 ;
  assign n38036 = ~n38033 & n38035 ;
  assign n38037 = n3671 ^ n1061 ^ 1'b0 ;
  assign n38038 = n2342 & n38037 ;
  assign n38039 = ( n5685 & n22611 ) | ( n5685 & n24179 ) | ( n22611 & n24179 ) ;
  assign n38040 = n811 | n23338 ;
  assign n38041 = n26303 ^ n4082 ^ 1'b0 ;
  assign n38042 = ~n19 & n1874 ;
  assign n38043 = n38042 ^ n20573 ^ 1'b0 ;
  assign n38044 = n13179 & n38043 ;
  assign n38045 = n1441 ^ n1417 ^ 1'b0 ;
  assign n38046 = n29594 & n38045 ;
  assign n38047 = n29882 & n36427 ;
  assign n38048 = ~n38046 & n38047 ;
  assign n38049 = n3901 & ~n24006 ;
  assign n38050 = n38049 ^ n12798 ^ 1'b0 ;
  assign n38051 = ( n856 & n9352 ) | ( n856 & ~n38050 ) | ( n9352 & ~n38050 ) ;
  assign n38052 = n35036 & ~n38051 ;
  assign n38053 = n11374 & n38052 ;
  assign n38054 = n908 & ~n38053 ;
  assign n38055 = n38048 & n38054 ;
  assign n38056 = n610 & ~n3279 ;
  assign n38057 = n14265 ^ n10303 ^ 1'b0 ;
  assign n38058 = ( n12206 & n12661 ) | ( n12206 & ~n38057 ) | ( n12661 & ~n38057 ) ;
  assign n38059 = n7483 ^ n7373 ^ 1'b0 ;
  assign n38060 = n4619 | n38059 ;
  assign n38061 = n3756 | n38060 ;
  assign n38062 = n1637 | n7231 ;
  assign n38063 = n38061 | n38062 ;
  assign n38064 = n15836 ^ n9646 ^ 1'b0 ;
  assign n38065 = n1409 & n38064 ;
  assign n38066 = n26224 ^ n1173 ^ 1'b0 ;
  assign n38067 = ~n11291 & n14710 ;
  assign n38068 = n1154 | n31648 ;
  assign n38069 = n38068 ^ n30563 ^ 1'b0 ;
  assign n38071 = n15771 ^ n2268 ^ 1'b0 ;
  assign n38070 = n12720 & ~n16459 ;
  assign n38072 = n38071 ^ n38070 ^ 1'b0 ;
  assign n38073 = n38072 ^ n8250 ^ 1'b0 ;
  assign n38074 = ~n3286 & n5716 ;
  assign n38075 = ~n938 & n38074 ;
  assign n38076 = n947 & n8619 ;
  assign n38077 = n4797 & n7803 ;
  assign n38078 = ~n16178 & n38077 ;
  assign n38079 = n26574 ^ n23814 ^ 1'b0 ;
  assign n38080 = n8368 ^ n6307 ^ 1'b0 ;
  assign n38081 = n4274 | n4747 ;
  assign n38082 = n4747 & ~n38081 ;
  assign n38083 = n13009 | n38082 ;
  assign n38084 = ~n5570 & n9954 ;
  assign n38085 = n5570 & n38084 ;
  assign n38086 = n38085 ^ n31916 ^ 1'b0 ;
  assign n38087 = n38083 | n38086 ;
  assign n38088 = n20961 & ~n38087 ;
  assign n38089 = n38087 & n38088 ;
  assign n38090 = ~n15457 & n32602 ;
  assign n38091 = n3826 & ~n8948 ;
  assign n38092 = n38091 ^ n9069 ^ 1'b0 ;
  assign n38093 = n10201 & ~n38092 ;
  assign n38094 = n274 & n2436 ;
  assign n38095 = n428 | n8030 ;
  assign n38096 = n38094 & ~n38095 ;
  assign n38097 = n5532 & n8292 ;
  assign n38098 = n38097 ^ n23826 ^ 1'b0 ;
  assign n38100 = n5420 & ~n35260 ;
  assign n38099 = n3271 & n14398 ;
  assign n38101 = n38100 ^ n38099 ^ 1'b0 ;
  assign n38102 = n8269 | n14187 ;
  assign n38103 = n2850 | n38102 ;
  assign n38104 = n3141 & n38103 ;
  assign n38105 = n21423 ^ n12534 ^ 1'b0 ;
  assign n38106 = n23186 & n38105 ;
  assign n38107 = ( ~n5180 & n7848 ) | ( ~n5180 & n34500 ) | ( n7848 & n34500 ) ;
  assign n38108 = n1414 & n38107 ;
  assign n38109 = ( n840 & n1745 ) | ( n840 & n9540 ) | ( n1745 & n9540 ) ;
  assign n38110 = ~n8463 & n38109 ;
  assign n38111 = ~n22342 & n38110 ;
  assign n38112 = n17 | n8130 ;
  assign n38114 = ~n5691 & n18029 ;
  assign n38115 = n38114 ^ n5948 ^ 1'b0 ;
  assign n38113 = n21298 & n31007 ;
  assign n38116 = n38115 ^ n38113 ^ n8751 ;
  assign n38117 = ~n4855 & n26684 ;
  assign n38118 = n715 & ~n32628 ;
  assign n38119 = ~n19128 & n38118 ;
  assign n38120 = ~n4527 & n6192 ;
  assign n38121 = x8 & ~n5018 ;
  assign n38122 = n2414 | n9934 ;
  assign n38123 = ~n5856 & n20248 ;
  assign n38124 = ~n19144 & n38123 ;
  assign n38125 = n38124 ^ n15985 ^ 1'b0 ;
  assign n38126 = n8317 | n38125 ;
  assign n38127 = n1820 & ~n8107 ;
  assign n38128 = ~n710 & n38127 ;
  assign n38129 = ~n4360 & n38128 ;
  assign n38130 = ~n3594 & n12100 ;
  assign n38131 = ~n19072 & n21444 ;
  assign n38132 = n12534 ^ n3260 ^ 1'b0 ;
  assign n38133 = n15593 ^ n8181 ^ 1'b0 ;
  assign n38135 = ~n7136 & n8931 ;
  assign n38134 = ~n14779 & n31500 ;
  assign n38136 = n38135 ^ n38134 ^ 1'b0 ;
  assign n38137 = n37826 ^ n24900 ^ 1'b0 ;
  assign n38138 = n11388 & n38137 ;
  assign n38139 = n8461 | n17090 ;
  assign n38140 = ~n1263 & n2261 ;
  assign n38141 = n12087 | n32945 ;
  assign n38142 = ~n713 & n9354 ;
  assign n38143 = n1687 | n38142 ;
  assign n38144 = n38143 ^ n27640 ^ 1'b0 ;
  assign n38145 = n15134 ^ n12898 ^ 1'b0 ;
  assign n38146 = n8581 | n38145 ;
  assign n38147 = n1637 & ~n16527 ;
  assign n38148 = n38147 ^ n4440 ^ 1'b0 ;
  assign n38149 = n25361 | n38148 ;
  assign n38150 = n5871 | n8125 ;
  assign n38151 = n32563 ^ n17281 ^ 1'b0 ;
  assign n38153 = n7056 & ~n10257 ;
  assign n38154 = ~n596 & n38153 ;
  assign n38152 = n6400 & ~n11588 ;
  assign n38155 = n38154 ^ n38152 ^ 1'b0 ;
  assign n38156 = n5194 ^ n2168 ^ 1'b0 ;
  assign n38157 = n30783 & n38156 ;
  assign n38158 = n38157 ^ n28856 ^ 1'b0 ;
  assign n38159 = n21638 | n31752 ;
  assign n38160 = n38158 | n38159 ;
  assign n38161 = n2529 | n6809 ;
  assign n38162 = n438 | n38161 ;
  assign n38163 = n14646 ^ n8246 ^ 1'b0 ;
  assign n38164 = n10377 & ~n24531 ;
  assign n38165 = n37417 ^ n3312 ^ 1'b0 ;
  assign n38166 = n12104 & n38165 ;
  assign n38167 = n38166 ^ n33202 ^ 1'b0 ;
  assign n38168 = n32321 ^ n2968 ^ 1'b0 ;
  assign n38169 = n2093 | n9535 ;
  assign n38170 = n8520 | n10294 ;
  assign n38171 = n15832 ^ n9036 ^ 1'b0 ;
  assign n38172 = n2212 | n2328 ;
  assign n38173 = n2328 & ~n38172 ;
  assign n38174 = n653 | n38173 ;
  assign n38175 = n907 | n3779 ;
  assign n38176 = n907 & ~n38175 ;
  assign n38177 = n38174 & ~n38176 ;
  assign n38178 = n38177 ^ n12636 ^ 1'b0 ;
  assign n38179 = n26052 & n38178 ;
  assign n38180 = n497 | n13830 ;
  assign n38181 = n36137 ^ n10475 ^ 1'b0 ;
  assign n38183 = n3777 | n12871 ;
  assign n38184 = n38183 ^ n10973 ^ 1'b0 ;
  assign n38182 = ~n12749 & n27676 ;
  assign n38185 = n38184 ^ n38182 ^ n14670 ;
  assign n38186 = n19239 ^ n1961 ^ 1'b0 ;
  assign n38187 = n14454 & n38186 ;
  assign n38188 = n33083 ^ n21545 ^ 1'b0 ;
  assign n38189 = n16567 | n38188 ;
  assign n38190 = ~n84 & n28088 ;
  assign n38191 = n38190 ^ n14339 ^ 1'b0 ;
  assign n38192 = n13691 | n35621 ;
  assign n38193 = n3939 & ~n38192 ;
  assign n38194 = n24930 ^ n15015 ^ 1'b0 ;
  assign n38195 = n2842 ^ n2012 ^ 1'b0 ;
  assign n38196 = n2219 & n38195 ;
  assign n38197 = n14236 | n38196 ;
  assign n38198 = n25273 | n27570 ;
  assign n38199 = n8409 ^ n4639 ^ 1'b0 ;
  assign n38200 = n38199 ^ n11266 ^ 1'b0 ;
  assign n38201 = ~n37131 & n38200 ;
  assign n38202 = n33712 ^ n4899 ^ n1124 ;
  assign n38203 = n6921 & ~n28255 ;
  assign n38204 = n10261 & n38203 ;
  assign n38205 = n7247 & n37584 ;
  assign n38206 = n38205 ^ n20327 ^ 1'b0 ;
  assign n38207 = n9751 ^ n6501 ^ 1'b0 ;
  assign n38208 = n14662 & ~n38207 ;
  assign n38209 = n11338 | n38208 ;
  assign n38210 = n21785 & n33539 ;
  assign n38211 = ~n1177 & n20213 ;
  assign n38212 = n12325 ^ n6715 ^ 1'b0 ;
  assign n38213 = n28682 & n38212 ;
  assign n38214 = n340 & n1375 ;
  assign n38215 = ~n38213 & n38214 ;
  assign n38216 = n13293 & ~n32085 ;
  assign n38217 = n2566 & n38216 ;
  assign n38218 = ~n31007 & n38217 ;
  assign n38219 = n26129 ^ n5657 ^ 1'b0 ;
  assign n38220 = n16263 & ~n38219 ;
  assign n38221 = n246 & ~n10035 ;
  assign n38222 = n23758 & ~n38221 ;
  assign n38223 = ~n38220 & n38222 ;
  assign n38225 = n20612 & ~n21360 ;
  assign n38226 = n38225 ^ n2394 ^ 1'b0 ;
  assign n38227 = ~n12402 & n38226 ;
  assign n38224 = n717 & n10541 ;
  assign n38228 = n38227 ^ n38224 ^ 1'b0 ;
  assign n38229 = ~n25053 & n37783 ;
  assign n38230 = n30701 & n38229 ;
  assign n38231 = n2953 | n4947 ;
  assign n38232 = ~n9733 & n38231 ;
  assign n38233 = n32668 & n37031 ;
  assign n38234 = n21669 & ~n28862 ;
  assign n38235 = ~n12160 & n34211 ;
  assign n38236 = n38235 ^ n690 ^ 1'b0 ;
  assign n38237 = n15615 & n38236 ;
  assign n38238 = n38237 ^ n941 ^ 1'b0 ;
  assign n38239 = n8990 & ~n12002 ;
  assign n38240 = n38239 ^ n36125 ^ 1'b0 ;
  assign n38241 = n10153 ^ n6890 ^ 1'b0 ;
  assign n38242 = ( n13197 & n15204 ) | ( n13197 & n38241 ) | ( n15204 & n38241 ) ;
  assign n38243 = ~n10687 & n37666 ;
  assign n38244 = ~n1213 & n38243 ;
  assign n38245 = n38244 ^ n16307 ^ 1'b0 ;
  assign n38246 = n37512 & n38245 ;
  assign n38247 = ~n2762 & n38246 ;
  assign n38248 = ~n169 & n35094 ;
  assign n38250 = n293 & n315 ;
  assign n38251 = n12855 ^ n1591 ^ 1'b0 ;
  assign n38252 = n16418 | n38251 ;
  assign n38253 = n5131 & ~n38252 ;
  assign n38254 = n38250 & n38253 ;
  assign n38249 = n514 & ~n6916 ;
  assign n38255 = n38254 ^ n38249 ^ 1'b0 ;
  assign n38256 = ~n1229 & n38255 ;
  assign n38257 = n38256 ^ n6738 ^ 1'b0 ;
  assign n38258 = n38257 ^ n28810 ^ 1'b0 ;
  assign n38259 = ~n6521 & n22531 ;
  assign n38260 = ~n26776 & n38259 ;
  assign n38261 = n8970 & n38260 ;
  assign n38262 = ~n3773 & n15781 ;
  assign n38264 = n20578 ^ n5061 ^ 1'b0 ;
  assign n38263 = n7640 & ~n16695 ;
  assign n38265 = n38264 ^ n38263 ^ 1'b0 ;
  assign n38266 = n776 & n15792 ;
  assign n38267 = n1202 | n20862 ;
  assign n38268 = n1202 & ~n38267 ;
  assign n38269 = n2481 & n2512 ;
  assign n38270 = ~n2481 & n38269 ;
  assign n38271 = n38268 | n38270 ;
  assign n38272 = n12266 & ~n38271 ;
  assign n38273 = n38272 ^ n10902 ^ 1'b0 ;
  assign n38274 = ~n38266 & n38273 ;
  assign n38275 = n11592 & ~n22707 ;
  assign n38277 = n1950 & n17690 ;
  assign n38278 = ~n8513 & n38277 ;
  assign n38276 = n378 & n6079 ;
  assign n38279 = n38278 ^ n38276 ^ 1'b0 ;
  assign n38280 = n4522 ^ n2358 ^ 1'b0 ;
  assign n38281 = n17631 ^ n15414 ^ 1'b0 ;
  assign n38282 = n18373 & ~n38281 ;
  assign n38283 = ~n6159 & n38282 ;
  assign n38284 = ~n35718 & n38283 ;
  assign n38285 = n17445 & ~n27936 ;
  assign n38286 = n38284 & n38285 ;
  assign n38287 = n2027 | n8660 ;
  assign n38289 = ~n6974 & n10635 ;
  assign n38290 = ~n21811 & n38289 ;
  assign n38288 = n2963 | n33832 ;
  assign n38291 = n38290 ^ n38288 ^ 1'b0 ;
  assign n38292 = ~n1110 & n36529 ;
  assign n38293 = n1438 | n8264 ;
  assign n38294 = n38293 ^ n13488 ^ 1'b0 ;
  assign n38295 = n6874 | n18580 ;
  assign n38296 = n18833 & n33125 ;
  assign n38297 = ~n38295 & n38296 ;
  assign n38298 = n3631 & n11851 ;
  assign n38299 = n38298 ^ n10025 ^ 1'b0 ;
  assign n38300 = ~n7915 & n24569 ;
  assign n38302 = n33408 ^ n14106 ^ 1'b0 ;
  assign n38301 = n16150 | n22762 ;
  assign n38303 = n38302 ^ n38301 ^ 1'b0 ;
  assign n38304 = n30916 & n31643 ;
  assign n38305 = n24370 ^ n19408 ^ 1'b0 ;
  assign n38306 = n22899 & ~n23796 ;
  assign n38307 = n1933 & ~n9851 ;
  assign n38308 = n25711 & ~n38307 ;
  assign n38309 = ~n3546 & n13007 ;
  assign n38310 = n34749 & n38309 ;
  assign n38311 = n35917 ^ n435 ^ 1'b0 ;
  assign n38312 = n31231 & ~n38311 ;
  assign n38313 = n38312 ^ n7265 ^ 1'b0 ;
  assign n38314 = n5872 & n13679 ;
  assign n38315 = n38314 ^ n6424 ^ 1'b0 ;
  assign n38316 = n38315 ^ n15796 ^ 1'b0 ;
  assign n38317 = n25239 & n38316 ;
  assign n38318 = n38317 ^ n19068 ^ 1'b0 ;
  assign n38319 = n19568 ^ n5535 ^ 1'b0 ;
  assign n38320 = n7938 | n38319 ;
  assign n38321 = n38320 ^ n7355 ^ 1'b0 ;
  assign n38322 = ~n2987 & n13639 ;
  assign n38323 = n530 & n9794 ;
  assign n38324 = n2655 & n38323 ;
  assign n38325 = n38324 ^ n3028 ^ 1'b0 ;
  assign n38326 = n6170 | n21788 ;
  assign n38327 = n38326 ^ n1889 ^ 1'b0 ;
  assign n38328 = n38327 ^ n616 ^ 1'b0 ;
  assign n38329 = n5354 & ~n6390 ;
  assign n38330 = ~n6325 & n11615 ;
  assign n38331 = n38330 ^ n6580 ^ 1'b0 ;
  assign n38332 = n2578 & ~n16263 ;
  assign n38333 = n299 & ~n37436 ;
  assign n38334 = n12046 & n38333 ;
  assign n38335 = n5148 & ~n7815 ;
  assign n38336 = n38335 ^ n33029 ^ n17192 ;
  assign n38337 = n14351 ^ n931 ^ 1'b0 ;
  assign n38338 = n21152 | n38337 ;
  assign n38339 = n38338 ^ n5817 ^ 1'b0 ;
  assign n38340 = n12982 & ~n13790 ;
  assign n38341 = n38340 ^ n18065 ^ 1'b0 ;
  assign n38342 = n23206 ^ n4243 ^ 1'b0 ;
  assign n38343 = n4112 & ~n17001 ;
  assign n38344 = n36068 ^ n7972 ^ 1'b0 ;
  assign n38345 = n28442 & n38344 ;
  assign n38347 = n2567 & n5995 ;
  assign n38348 = n7745 | n16079 ;
  assign n38349 = n23037 & n38348 ;
  assign n38350 = n38347 & n38349 ;
  assign n38346 = n11260 & n16461 ;
  assign n38351 = n38350 ^ n38346 ^ 1'b0 ;
  assign n38352 = n3679 | n38351 ;
  assign n38353 = n7582 | n20696 ;
  assign n38354 = n1254 & ~n38353 ;
  assign n38355 = ~n9742 & n14135 ;
  assign n38356 = n38355 ^ n2410 ^ 1'b0 ;
  assign n38357 = n17947 | n23772 ;
  assign n38358 = n5362 & ~n38357 ;
  assign n38359 = n7269 & ~n35103 ;
  assign n38360 = n11917 & n30003 ;
  assign n38363 = n7425 & ~n25674 ;
  assign n38361 = n536 | n1785 ;
  assign n38362 = n35913 | n38361 ;
  assign n38364 = n38363 ^ n38362 ^ 1'b0 ;
  assign n38365 = n4700 & n13896 ;
  assign n38366 = n38365 ^ n5013 ^ 1'b0 ;
  assign n38367 = n9934 & ~n38366 ;
  assign n38368 = n16882 ^ n2313 ^ 1'b0 ;
  assign n38369 = n21232 & ~n38368 ;
  assign n38371 = x9 & ~n991 ;
  assign n38370 = n3928 & n15321 ;
  assign n38372 = n38371 ^ n38370 ^ 1'b0 ;
  assign n38373 = n38369 & ~n38372 ;
  assign n38374 = n4650 ^ n2430 ^ 1'b0 ;
  assign n38375 = n38373 & n38374 ;
  assign n38376 = n1772 & n5324 ;
  assign n38377 = n38376 ^ n36247 ^ 1'b0 ;
  assign n38378 = n5802 & ~n12664 ;
  assign n38379 = n2517 | n27870 ;
  assign n38380 = n25527 & ~n32167 ;
  assign n38381 = n8887 & ~n15623 ;
  assign n38382 = n6655 & n7808 ;
  assign n38383 = n14848 & n38382 ;
  assign n38384 = n35172 ^ n31776 ^ 1'b0 ;
  assign n38385 = n25652 ^ n19315 ^ 1'b0 ;
  assign n38386 = n1880 & n20406 ;
  assign n38387 = n38386 ^ n30890 ^ 1'b0 ;
  assign n38388 = n37916 | n38387 ;
  assign n38389 = n375 | n7442 ;
  assign n38390 = n18580 & ~n38389 ;
  assign n38391 = ~n9240 & n32940 ;
  assign n38392 = n17892 ^ n530 ^ 1'b0 ;
  assign n38393 = ~n27822 & n38392 ;
  assign n38394 = n3883 | n5575 ;
  assign n38395 = n5575 & ~n38394 ;
  assign n38396 = n3008 | n38395 ;
  assign n38397 = ( ~n12862 & n14405 ) | ( ~n12862 & n38396 ) | ( n14405 & n38396 ) ;
  assign n38398 = ~n23302 & n33397 ;
  assign n38399 = n7029 & n29685 ;
  assign n38400 = n38399 ^ n35838 ^ 1'b0 ;
  assign n38401 = n31465 ^ n25508 ^ 1'b0 ;
  assign n38402 = n20301 ^ n1848 ^ 1'b0 ;
  assign n38403 = ~n38401 & n38402 ;
  assign n38404 = n29551 ^ n27504 ^ 1'b0 ;
  assign n38405 = ~n3411 & n10658 ;
  assign n38406 = n1472 & n16138 ;
  assign n38407 = n5845 & ~n9758 ;
  assign n38408 = n7810 & n27221 ;
  assign n38409 = n4904 | n35213 ;
  assign n38410 = n9717 ^ n1089 ^ 1'b0 ;
  assign n38411 = n5656 & n38410 ;
  assign n38412 = n8950 ^ n3406 ^ 1'b0 ;
  assign n38413 = n6587 ^ n915 ^ 1'b0 ;
  assign n38414 = ~n38412 & n38413 ;
  assign n38415 = n1571 | n3088 ;
  assign n38416 = ~n22483 & n38415 ;
  assign n38417 = n22856 ^ n6072 ^ 1'b0 ;
  assign n38418 = ~n12171 & n38417 ;
  assign n38419 = n3331 ^ n133 ^ 1'b0 ;
  assign n38420 = n17397 & ~n38419 ;
  assign n38421 = ~n29447 & n38420 ;
  assign n38422 = n5382 & n16251 ;
  assign n38423 = n17003 & n25118 ;
  assign n38424 = n8262 | n8756 ;
  assign n38425 = n15456 ^ n8460 ^ 1'b0 ;
  assign n38426 = n20342 | n38425 ;
  assign n38427 = n26986 ^ n7546 ^ x5 ;
  assign n38428 = n11690 | n35633 ;
  assign n38429 = n18982 ^ n14992 ^ n3025 ;
  assign n38430 = n25773 ^ n18349 ^ 1'b0 ;
  assign n38431 = n37771 ^ n29074 ^ 1'b0 ;
  assign n38432 = n3318 | n36657 ;
  assign n38433 = n3431 | n38432 ;
  assign n38434 = n663 & ~n33126 ;
  assign n38435 = n38434 ^ n25751 ^ 1'b0 ;
  assign n38436 = n38433 & ~n38435 ;
  assign n38437 = ~n2789 & n12205 ;
  assign n38438 = n32587 & n38437 ;
  assign n38439 = n31829 ^ n1825 ^ 1'b0 ;
  assign n38440 = ~n5857 & n38439 ;
  assign n38441 = n30667 ^ n1406 ^ 1'b0 ;
  assign n38442 = n16311 ^ n4365 ^ 1'b0 ;
  assign n38443 = n8707 ^ n5278 ^ 1'b0 ;
  assign n38444 = n1337 | n38443 ;
  assign n38445 = ~n988 & n37916 ;
  assign n38446 = n3378 & n38445 ;
  assign n38447 = n38444 & ~n38446 ;
  assign n38448 = ~n669 & n20625 ;
  assign n38449 = n6519 | n9672 ;
  assign n38450 = n38449 ^ n4375 ^ 1'b0 ;
  assign n38451 = n11239 ^ n4733 ^ 1'b0 ;
  assign n38452 = n8542 & n38451 ;
  assign n38453 = n19406 & ~n38452 ;
  assign n38454 = n135 & ~n38453 ;
  assign n38455 = n1484 | n38454 ;
  assign n38458 = n29441 ^ n16636 ^ 1'b0 ;
  assign n38459 = ~n14893 & n38458 ;
  assign n38456 = n6022 | n16393 ;
  assign n38457 = n15426 & ~n38456 ;
  assign n38460 = n38459 ^ n38457 ^ 1'b0 ;
  assign n38461 = ~n25119 & n27773 ;
  assign n38462 = n37805 & n38461 ;
  assign n38463 = n3311 & ~n38462 ;
  assign n38464 = n24378 | n33091 ;
  assign n38465 = n31807 & ~n38464 ;
  assign n38466 = ~n10718 & n32051 ;
  assign n38467 = ~n3472 & n38466 ;
  assign n38468 = n12969 & n23329 ;
  assign n38469 = ~n3096 & n38468 ;
  assign n38470 = n8744 | n18488 ;
  assign n38471 = n2875 ^ n316 ^ 1'b0 ;
  assign n38472 = ~n23737 & n38471 ;
  assign n38473 = n38470 & n38472 ;
  assign n38474 = n542 | n1759 ;
  assign n38475 = n3056 & n6249 ;
  assign n38476 = n6493 & ~n15297 ;
  assign n38477 = ~n38475 & n38476 ;
  assign n38478 = n3939 & n4508 ;
  assign n38479 = ~n24722 & n34414 ;
  assign n38480 = n6383 & ~n38479 ;
  assign n38481 = n677 | n38480 ;
  assign n38482 = n38481 ^ n6822 ^ 1'b0 ;
  assign n38483 = n11821 & n38482 ;
  assign n38484 = ~n18624 & n20284 ;
  assign n38485 = n38484 ^ n4742 ^ 1'b0 ;
  assign n38486 = ~n11622 & n38485 ;
  assign n38487 = ~n15029 & n20348 ;
  assign n38490 = n2652 & ~n27555 ;
  assign n38491 = n38490 ^ n33018 ^ n962 ;
  assign n38492 = n15146 & n38491 ;
  assign n38488 = ~n2141 & n14768 ;
  assign n38489 = n38488 ^ n2410 ^ 1'b0 ;
  assign n38493 = n38492 ^ n38489 ^ n25954 ;
  assign n38494 = n12170 | n15167 ;
  assign n38495 = n1226 & n38494 ;
  assign n38496 = ~n8804 & n38495 ;
  assign n38497 = x2 & ~n38496 ;
  assign n38498 = n38497 ^ n25574 ^ 1'b0 ;
  assign n38499 = n10521 ^ n10059 ^ n1672 ;
  assign n38500 = n13429 & ~n38499 ;
  assign n38501 = n19128 ^ n10572 ^ 1'b0 ;
  assign n38502 = ~n2212 & n38501 ;
  assign n38503 = n38502 ^ n17360 ^ 1'b0 ;
  assign n38504 = n38503 ^ n36658 ^ 1'b0 ;
  assign n38505 = n23692 & n26065 ;
  assign n38506 = n38505 ^ n33910 ^ 1'b0 ;
  assign n38507 = n7977 & n24215 ;
  assign n38508 = n38507 ^ n19862 ^ 1'b0 ;
  assign n38509 = n22958 ^ n14569 ^ 1'b0 ;
  assign n38510 = n1276 ^ n278 ^ 1'b0 ;
  assign n38511 = n37422 & ~n38510 ;
  assign n38512 = ~n475 & n38511 ;
  assign n38517 = n1350 & n2060 ;
  assign n38518 = n38517 ^ n3603 ^ 1'b0 ;
  assign n38513 = ~n381 & n5694 ;
  assign n38514 = n38513 ^ n10624 ^ 1'b0 ;
  assign n38515 = n7880 | n38514 ;
  assign n38516 = ~n1565 & n38515 ;
  assign n38519 = n38518 ^ n38516 ^ 1'b0 ;
  assign n38520 = n1961 | n28233 ;
  assign n38521 = n14177 & ~n18558 ;
  assign n38522 = n3221 & n38521 ;
  assign n38523 = n26464 ^ n11624 ^ 1'b0 ;
  assign n38524 = n713 ^ n678 ^ 1'b0 ;
  assign n38525 = n22864 | n38524 ;
  assign n38526 = n12236 ^ n9376 ^ n3211 ;
  assign n38527 = n13690 ^ n10996 ^ 1'b0 ;
  assign n38528 = n16476 & ~n19466 ;
  assign n38529 = n38528 ^ n3720 ^ 1'b0 ;
  assign n38530 = n38527 & n38529 ;
  assign n38531 = n38530 ^ n1452 ^ 1'b0 ;
  assign n38532 = n18888 | n20994 ;
  assign n38533 = ~n339 & n2900 ;
  assign n38534 = n38533 ^ n20384 ^ 1'b0 ;
  assign n38535 = n2185 & ~n38534 ;
  assign n38536 = n38535 ^ n31412 ^ 1'b0 ;
  assign n38537 = n4022 & n38536 ;
  assign n38538 = n756 & ~n38537 ;
  assign n38539 = n30999 ^ n8594 ^ 1'b0 ;
  assign n38540 = n10876 | n38539 ;
  assign n38541 = ~n21372 & n21408 ;
  assign n38542 = ~n6951 & n38541 ;
  assign n38544 = n34804 ^ n1081 ^ 1'b0 ;
  assign n38543 = n5739 | n10007 ;
  assign n38545 = n38544 ^ n38543 ^ 1'b0 ;
  assign n38546 = ~n9184 & n31891 ;
  assign n38547 = n1031 & ~n16156 ;
  assign n38548 = n26418 & n38547 ;
  assign n38550 = n3182 | n5167 ;
  assign n38551 = n8461 | n38550 ;
  assign n38549 = n2905 & n13906 ;
  assign n38552 = n38551 ^ n38549 ^ 1'b0 ;
  assign n38553 = ~n2919 & n17159 ;
  assign n38554 = n38553 ^ n3074 ^ 1'b0 ;
  assign n38555 = n7755 & ~n19619 ;
  assign n38556 = ~n8751 & n38555 ;
  assign n38557 = ~n20890 & n38556 ;
  assign n38558 = n13094 ^ n11329 ^ 1'b0 ;
  assign n38559 = n20838 | n38558 ;
  assign n38560 = n206 | n38559 ;
  assign n38561 = n16979 & ~n38560 ;
  assign n38562 = ( n9504 & n13847 ) | ( n9504 & n27522 ) | ( n13847 & n27522 ) ;
  assign n38563 = ~n7676 & n38562 ;
  assign n38565 = n14784 ^ n11726 ^ 1'b0 ;
  assign n38566 = n1922 | n38565 ;
  assign n38564 = n1194 & ~n12743 ;
  assign n38567 = n38566 ^ n38564 ^ 1'b0 ;
  assign n38568 = ~n18384 & n38567 ;
  assign n38569 = n38568 ^ n13723 ^ 1'b0 ;
  assign n38570 = n1175 & ~n2956 ;
  assign n38571 = n19444 ^ n12639 ^ 1'b0 ;
  assign n38572 = ~n10020 & n17765 ;
  assign n38573 = ( n1349 & n11463 ) | ( n1349 & n14168 ) | ( n11463 & n14168 ) ;
  assign n38574 = n601 & ~n17270 ;
  assign n38575 = ~n38265 & n38574 ;
  assign n38576 = n38575 ^ n8697 ^ 1'b0 ;
  assign n38577 = n26095 ^ n9067 ^ 1'b0 ;
  assign n38578 = ~n15838 & n23322 ;
  assign n38579 = n12407 & n38578 ;
  assign n38580 = n5537 & n9703 ;
  assign n38581 = ~n17508 & n38580 ;
  assign n38582 = n2137 & ~n9118 ;
  assign n38583 = ~n25984 & n38582 ;
  assign n38584 = ~n24991 & n38583 ;
  assign n38585 = n33197 ^ n8885 ^ 1'b0 ;
  assign n38586 = n17969 & n38585 ;
  assign n38587 = n3804 & ~n7007 ;
  assign n38588 = n38587 ^ n3331 ^ 1'b0 ;
  assign n38589 = n30552 ^ n246 ^ 1'b0 ;
  assign n38590 = ~n2912 & n18832 ;
  assign n38591 = n38590 ^ n10582 ^ 1'b0 ;
  assign n38592 = n29166 ^ n3820 ^ 1'b0 ;
  assign n38593 = n28674 | n38592 ;
  assign n38594 = n38593 ^ n33602 ^ 1'b0 ;
  assign n38595 = n957 & ~n38594 ;
  assign n38596 = n4117 | n37533 ;
  assign n38597 = n38596 ^ n24970 ^ 1'b0 ;
  assign n38598 = ~n10233 & n36018 ;
  assign n38599 = n38598 ^ n20830 ^ 1'b0 ;
  assign n38600 = n36259 ^ n24008 ^ n8843 ;
  assign n38601 = n9780 ^ n107 ^ 1'b0 ;
  assign n38602 = n5452 ^ n2665 ^ 1'b0 ;
  assign n38603 = n4012 | n17871 ;
  assign n38604 = n38603 ^ n17291 ^ 1'b0 ;
  assign n38605 = n6492 & n7450 ;
  assign n38606 = ~n29359 & n38605 ;
  assign n38607 = n5067 | n20723 ;
  assign n38608 = ( n495 & n38606 ) | ( n495 & n38607 ) | ( n38606 & n38607 ) ;
  assign n38609 = n16397 ^ n175 ^ 1'b0 ;
  assign n38610 = ~n4022 & n38609 ;
  assign n38611 = n5814 ^ n3311 ^ 1'b0 ;
  assign n38612 = n38611 ^ n27435 ^ n2830 ;
  assign n38613 = n456 | n38612 ;
  assign n38614 = n38610 | n38613 ;
  assign n38615 = ~n4163 & n7850 ;
  assign n38616 = n4129 & n38615 ;
  assign n38617 = n3844 | n16799 ;
  assign n38618 = n4712 & n38617 ;
  assign n38619 = n8000 ^ n754 ^ 1'b0 ;
  assign n38620 = ~n5733 & n14805 ;
  assign n38621 = n38620 ^ n5716 ^ 1'b0 ;
  assign n38622 = n25637 & ~n38621 ;
  assign n38623 = n7237 & ~n38622 ;
  assign n38624 = n9931 ^ n741 ^ 1'b0 ;
  assign n38625 = n547 & ~n38624 ;
  assign n38626 = n18471 ^ n12190 ^ 1'b0 ;
  assign n38627 = n33669 & n34863 ;
  assign n38628 = n12404 & ~n37304 ;
  assign n38629 = n9697 & n38628 ;
  assign n38630 = n4105 & n8457 ;
  assign n38631 = n6492 | n22207 ;
  assign n38632 = n38630 | n38631 ;
  assign n38633 = n38632 ^ n18320 ^ 1'b0 ;
  assign n38634 = n15522 ^ n9023 ^ 1'b0 ;
  assign n38635 = n38633 | n38634 ;
  assign n38636 = n13960 ^ n7975 ^ 1'b0 ;
  assign n38637 = ~n28068 & n38636 ;
  assign n38638 = n13629 & n38637 ;
  assign n38639 = n30898 ^ n13606 ^ n3527 ;
  assign n38640 = ~n3606 & n38639 ;
  assign n38641 = n38640 ^ n4374 ^ 1'b0 ;
  assign n38643 = n15905 | n20222 ;
  assign n38642 = n1611 & ~n32169 ;
  assign n38644 = n38643 ^ n38642 ^ 1'b0 ;
  assign n38645 = n2575 & n9592 ;
  assign n38646 = n23510 & ~n38645 ;
  assign n38647 = n6074 | n30616 ;
  assign n38648 = n37075 & ~n38647 ;
  assign n38649 = ~n6777 & n10138 ;
  assign n38650 = n38649 ^ n21537 ^ 1'b0 ;
  assign n38651 = n9719 | n38650 ;
  assign n38652 = ~n38648 & n38651 ;
  assign n38653 = n295 | n1472 ;
  assign n38654 = n9625 & n25118 ;
  assign n38655 = n13853 & ~n27188 ;
  assign n38656 = ~n2484 & n2549 ;
  assign n38657 = n4872 & ~n20640 ;
  assign n38658 = ~n38656 & n38657 ;
  assign n38659 = n6990 & n35575 ;
  assign n38660 = n512 ^ n232 ^ 1'b0 ;
  assign n38661 = n38660 ^ n5076 ^ 1'b0 ;
  assign n38662 = ~n4613 & n38661 ;
  assign n38663 = n4294 ^ n2028 ^ 1'b0 ;
  assign n38664 = n87 | n38663 ;
  assign n38665 = n38664 ^ n6596 ^ 1'b0 ;
  assign n38666 = n15497 & ~n24435 ;
  assign n38667 = n22868 & n38666 ;
  assign n38668 = n30444 ^ n2549 ^ 1'b0 ;
  assign n38669 = n5856 ^ n86 ^ 1'b0 ;
  assign n38672 = n21982 ^ n9340 ^ 1'b0 ;
  assign n38673 = n10624 | n38672 ;
  assign n38671 = ~n6442 & n6573 ;
  assign n38674 = n38673 ^ n38671 ^ 1'b0 ;
  assign n38670 = n1957 | n26082 ;
  assign n38675 = n38674 ^ n38670 ^ 1'b0 ;
  assign n38676 = n10490 & ~n38675 ;
  assign n38677 = n17974 ^ n3008 ^ 1'b0 ;
  assign n38678 = n10785 ^ n218 ^ 1'b0 ;
  assign n38679 = n9322 ^ n2771 ^ 1'b0 ;
  assign n38681 = n22363 ^ n10161 ^ 1'b0 ;
  assign n38682 = n7214 | n38681 ;
  assign n38680 = ~n11831 & n35018 ;
  assign n38683 = n38682 ^ n38680 ^ 1'b0 ;
  assign n38684 = n17004 ^ n7304 ^ 1'b0 ;
  assign n38685 = n4320 | n24149 ;
  assign n38686 = n20224 & ~n24506 ;
  assign n38687 = n38686 ^ n15711 ^ 1'b0 ;
  assign n38688 = n3459 | n5158 ;
  assign n38689 = n5158 & ~n38688 ;
  assign n38690 = n3539 | n38689 ;
  assign n38691 = n3539 & ~n38690 ;
  assign n38704 = n271 & n524 ;
  assign n38705 = ~n524 & n38704 ;
  assign n38706 = n8986 & ~n38705 ;
  assign n38699 = n677 | n2124 ;
  assign n38700 = n677 & ~n38699 ;
  assign n38701 = n5012 | n38700 ;
  assign n38702 = n5012 & ~n38701 ;
  assign n38692 = n268 ^ n267 ^ 1'b0 ;
  assign n38693 = n14365 | n38692 ;
  assign n38694 = n14365 & ~n38693 ;
  assign n38695 = n2694 & ~n3757 ;
  assign n38696 = ~n2694 & n38695 ;
  assign n38697 = n38694 & ~n38696 ;
  assign n38698 = n9950 & n38697 ;
  assign n38703 = n38702 ^ n38698 ^ 1'b0 ;
  assign n38707 = n38706 ^ n38703 ^ 1'b0 ;
  assign n38708 = n38691 | n38707 ;
  assign n38709 = n13266 & ~n38708 ;
  assign n38710 = n38709 ^ n2386 ^ 1'b0 ;
  assign n38711 = n23718 & n38710 ;
  assign n38712 = n4916 & n12205 ;
  assign n38713 = n38712 ^ n231 ^ 1'b0 ;
  assign n38714 = n23644 & ~n38713 ;
  assign n38715 = n21685 ^ n16440 ^ 1'b0 ;
  assign n38716 = n5232 & ~n38715 ;
  assign n38717 = n12159 ^ n8602 ^ 1'b0 ;
  assign n38718 = n19232 ^ n324 ^ 1'b0 ;
  assign n38719 = n15174 & n38718 ;
  assign n38720 = n17783 ^ n4882 ^ 1'b0 ;
  assign n38721 = n15706 & n38720 ;
  assign n38722 = n38721 ^ n35902 ^ 1'b0 ;
  assign n38723 = n3530 ^ n2923 ^ 1'b0 ;
  assign n38724 = n26161 | n38723 ;
  assign n38725 = n22890 ^ n10942 ^ 1'b0 ;
  assign n38726 = n3484 & n38725 ;
  assign n38727 = n6376 & ~n38726 ;
  assign n38728 = n35278 ^ n32957 ^ 1'b0 ;
  assign n38729 = ~n12498 & n38307 ;
  assign n38730 = n38729 ^ n13678 ^ 1'b0 ;
  assign n38731 = n38730 ^ n26453 ^ n2604 ;
  assign n38732 = n32263 ^ n785 ^ 1'b0 ;
  assign n38733 = n3385 | n21384 ;
  assign n38734 = n27774 | n38733 ;
  assign n38735 = n18993 | n35158 ;
  assign n38736 = n27016 ^ n1469 ^ 1'b0 ;
  assign n38737 = n29319 | n34893 ;
  assign n38738 = n1836 & n13314 ;
  assign n38739 = n904 | n38738 ;
  assign n38740 = n904 & ~n38739 ;
  assign n38741 = n14712 | n38740 ;
  assign n38742 = n14712 & ~n38741 ;
  assign n38746 = n56 & n75 ;
  assign n38743 = ~n1001 & n5083 ;
  assign n38744 = ~n5083 & n38743 ;
  assign n38745 = n7060 | n38744 ;
  assign n38747 = n38746 ^ n38745 ^ 1'b0 ;
  assign n38748 = n38742 & ~n38747 ;
  assign n38749 = n958 & ~n2875 ;
  assign n38750 = ~n958 & n38749 ;
  assign n38751 = ~n2896 & n38750 ;
  assign n38752 = n129 & ~n38751 ;
  assign n38753 = n853 | n1329 ;
  assign n38754 = n853 & ~n38753 ;
  assign n38755 = ~n1170 & n38754 ;
  assign n38756 = n38752 & ~n38755 ;
  assign n38757 = ~n38752 & n38756 ;
  assign n38758 = n38757 ^ n66 ^ 1'b0 ;
  assign n38759 = n38748 & ~n38758 ;
  assign n38761 = ~n1473 & n10615 ;
  assign n38762 = n1473 & n38761 ;
  assign n38760 = n596 & n9206 ;
  assign n38763 = n38762 ^ n38760 ^ 1'b0 ;
  assign n38764 = n38759 & ~n38763 ;
  assign n38765 = ~n16669 & n38764 ;
  assign n38766 = n16669 & n38765 ;
  assign n38767 = n12479 ^ n6370 ^ 1'b0 ;
  assign n38768 = n174 | n2001 ;
  assign n38769 = n18022 & ~n38768 ;
  assign n38770 = ~n782 & n866 ;
  assign n38771 = n18438 & n38770 ;
  assign n38772 = n38771 ^ n31417 ^ 1'b0 ;
  assign n38773 = n34309 ^ n4749 ^ 1'b0 ;
  assign n38774 = ~n38772 & n38773 ;
  assign n38775 = n13947 | n24487 ;
  assign n38776 = n726 & ~n10412 ;
  assign n38777 = ~n6882 & n38776 ;
  assign n38778 = n23455 ^ n15794 ^ 1'b0 ;
  assign n38779 = n15198 ^ n13397 ^ 1'b0 ;
  assign n38780 = ~n14573 & n38779 ;
  assign n38781 = n16423 & ~n23281 ;
  assign n38782 = ~n708 & n32114 ;
  assign n38783 = n32471 ^ n27468 ^ 1'b0 ;
  assign n38784 = n1316 & ~n10674 ;
  assign n38785 = n38784 ^ n8646 ^ 1'b0 ;
  assign n38786 = ~n5201 & n24733 ;
  assign n38787 = n36060 ^ n10891 ^ 1'b0 ;
  assign n38788 = n8951 | n10118 ;
  assign n38789 = n29480 ^ n4171 ^ 1'b0 ;
  assign n38790 = n28956 ^ n22107 ^ 1'b0 ;
  assign n38791 = n144 | n5169 ;
  assign n38792 = n38791 ^ n13631 ^ 1'b0 ;
  assign n38793 = n4474 & ~n5057 ;
  assign n38794 = ~n7697 & n38793 ;
  assign n38795 = n26732 | n38794 ;
  assign n38796 = n38792 & ~n38795 ;
  assign n38797 = n1177 | n22504 ;
  assign n38798 = n7543 | n23999 ;
  assign n38799 = n38798 ^ n5481 ^ 1'b0 ;
  assign n38800 = ~n22464 & n25625 ;
  assign n38801 = n532 & n38800 ;
  assign n38802 = n19841 ^ n8114 ^ 1'b0 ;
  assign n38803 = ~n38801 & n38802 ;
  assign n38804 = n7420 ^ n2872 ^ 1'b0 ;
  assign n38805 = n38462 ^ n2233 ^ 1'b0 ;
  assign n38806 = n8350 & ~n19138 ;
  assign n38807 = n21568 & ~n38806 ;
  assign n38808 = ~n7918 & n38807 ;
  assign n38809 = n28462 ^ n4589 ^ 1'b0 ;
  assign n38816 = n270 & ~n9184 ;
  assign n38817 = ~n270 & n38816 ;
  assign n38818 = n506 | n38817 ;
  assign n38810 = n653 & n4355 ;
  assign n38811 = ~n653 & n38810 ;
  assign n38812 = ~n37 & n38811 ;
  assign n38813 = ~n19 & n38812 ;
  assign n38814 = n19 & n38813 ;
  assign n38815 = n38814 ^ n4077 ^ 1'b0 ;
  assign n38819 = n38818 ^ n38815 ^ 1'b0 ;
  assign n38820 = n38809 & ~n38819 ;
  assign n38821 = n38820 ^ n9134 ^ 1'b0 ;
  assign n38822 = n38135 & n38821 ;
  assign n38823 = n6700 & n21985 ;
  assign n38824 = n38823 ^ n30662 ^ 1'b0 ;
  assign n38825 = n6981 & ~n33330 ;
  assign n38826 = n38825 ^ n22426 ^ 1'b0 ;
  assign n38827 = n38826 ^ n29566 ^ 1'b0 ;
  assign n38828 = n6658 ^ n4436 ^ 1'b0 ;
  assign n38829 = n38827 & n38828 ;
  assign n38830 = n16346 ^ n336 ^ 1'b0 ;
  assign n38835 = n36670 ^ n20522 ^ 1'b0 ;
  assign n38836 = n4229 | n38835 ;
  assign n38837 = n14059 & n38836 ;
  assign n38838 = n38837 ^ n4535 ^ 1'b0 ;
  assign n38839 = n17580 | n38838 ;
  assign n38831 = n4850 & ~n19719 ;
  assign n38832 = n38831 ^ n311 ^ 1'b0 ;
  assign n38833 = n15485 & n38832 ;
  assign n38834 = ~n1469 & n38833 ;
  assign n38840 = n38839 ^ n38834 ^ 1'b0 ;
  assign n38841 = n18977 & n20382 ;
  assign n38842 = n38841 ^ n24122 ^ 1'b0 ;
  assign n38843 = ~n14730 & n35534 ;
  assign n38844 = ~n38842 & n38843 ;
  assign n38845 = n29469 & ~n38844 ;
  assign n38846 = n3268 | n14886 ;
  assign n38847 = n484 | n38846 ;
  assign n38848 = n3440 & n6265 ;
  assign n38849 = n38848 ^ n8092 ^ 1'b0 ;
  assign n38850 = ~n813 & n38849 ;
  assign n38851 = n19629 & n30021 ;
  assign n38852 = n24300 ^ n4761 ^ 1'b0 ;
  assign n38853 = ~n9342 & n38852 ;
  assign n38855 = n11640 & ~n14343 ;
  assign n38856 = n38855 ^ n31117 ^ 1'b0 ;
  assign n38854 = n24507 & n29669 ;
  assign n38857 = n38856 ^ n38854 ^ 1'b0 ;
  assign n38858 = n8922 | n12681 ;
  assign n38860 = ~n4075 & n19158 ;
  assign n38861 = n38860 ^ n26802 ^ 1'b0 ;
  assign n38859 = n1003 | n19539 ;
  assign n38862 = n38861 ^ n38859 ^ 1'b0 ;
  assign n38863 = n38858 & n38862 ;
  assign n38864 = n11582 | n18899 ;
  assign n38865 = n38864 ^ n340 ^ 1'b0 ;
  assign n38866 = n2668 & n29259 ;
  assign n38867 = n38866 ^ n19419 ^ 1'b0 ;
  assign n38868 = n1602 | n3583 ;
  assign n38869 = n1602 & ~n38868 ;
  assign n38870 = n38057 & ~n38869 ;
  assign n38871 = n24 | n12291 ;
  assign n38872 = n24 & ~n38871 ;
  assign n38880 = n459 & ~n542 ;
  assign n38881 = n542 & n38880 ;
  assign n38882 = n10851 & ~n38881 ;
  assign n38873 = n806 & n1564 ;
  assign n38874 = ~n1564 & n38873 ;
  assign n38875 = n1304 & ~n38874 ;
  assign n38876 = ~n1304 & n38875 ;
  assign n38877 = n1496 & n38876 ;
  assign n38878 = ~n3080 & n5764 ;
  assign n38879 = n38877 & n38878 ;
  assign n38883 = n38882 ^ n38879 ^ 1'b0 ;
  assign n38884 = n38872 | n38883 ;
  assign n38885 = n38870 & ~n38884 ;
  assign n38886 = n38885 ^ n29695 ^ 1'b0 ;
  assign n38887 = n2730 | n38886 ;
  assign n38888 = n30947 | n38887 ;
  assign n38889 = n27820 | n36733 ;
  assign n38890 = n9273 & n27532 ;
  assign n38891 = ~n292 & n38890 ;
  assign n38892 = n30248 ^ n25987 ^ 1'b0 ;
  assign n38894 = n12457 | n16983 ;
  assign n38895 = n23981 & ~n38894 ;
  assign n38893 = n785 & ~n2812 ;
  assign n38896 = n38895 ^ n38893 ^ 1'b0 ;
  assign n38897 = n6376 & ~n30677 ;
  assign n38898 = n2481 & n35791 ;
  assign n38899 = n33631 | n38898 ;
  assign n38900 = n18936 ^ n4018 ^ 1'b0 ;
  assign n38901 = n4951 & n38900 ;
  assign n38902 = n38901 ^ n14522 ^ 1'b0 ;
  assign n38903 = n22768 ^ n14964 ^ 1'b0 ;
  assign n38904 = n12661 ^ n942 ^ 1'b0 ;
  assign n38905 = n32916 | n38904 ;
  assign n38906 = n4933 | n7814 ;
  assign n38907 = n3965 & ~n38906 ;
  assign n38908 = n35731 & n38907 ;
  assign n38909 = ( n1286 & n1982 ) | ( n1286 & ~n5187 ) | ( n1982 & ~n5187 ) ;
  assign n38910 = n3118 | n38909 ;
  assign n38911 = n15124 | n34912 ;
  assign n38912 = n4294 & ~n38911 ;
  assign n38914 = n4917 | n19070 ;
  assign n38913 = n23278 & ~n29687 ;
  assign n38915 = n38914 ^ n38913 ^ n7759 ;
  assign n38916 = n2189 & n8997 ;
  assign n38917 = n27568 ^ n14539 ^ 1'b0 ;
  assign n38918 = n14117 & ~n38917 ;
  assign n38919 = n17893 ^ n10600 ^ 1'b0 ;
  assign n38920 = n9638 & n23438 ;
  assign n38921 = n33287 ^ n2644 ^ 1'b0 ;
  assign n38922 = n38920 & ~n38921 ;
  assign n38923 = n38922 ^ n8888 ^ 1'b0 ;
  assign n38924 = n38923 ^ n6583 ^ 1'b0 ;
  assign n38925 = n9211 & n9490 ;
  assign n38926 = x2 | n38925 ;
  assign n38927 = n24225 ^ n7998 ^ 1'b0 ;
  assign n38928 = n24310 & ~n38927 ;
  assign n38929 = n38928 ^ n24322 ^ 1'b0 ;
  assign n38930 = n15115 ^ n4292 ^ 1'b0 ;
  assign n38931 = ~n1106 & n38930 ;
  assign n38932 = n7245 & n7550 ;
  assign n38933 = n764 & n38932 ;
  assign n38934 = ~n7424 & n38933 ;
  assign n38935 = n26899 ^ n15441 ^ 1'b0 ;
  assign n38937 = n1250 & n13856 ;
  assign n38938 = n461 | n3894 ;
  assign n38939 = n7136 & n38938 ;
  assign n38940 = ~n38937 & n38939 ;
  assign n38936 = n83 | n14219 ;
  assign n38941 = n38940 ^ n38936 ^ 1'b0 ;
  assign n38942 = ~n636 & n2969 ;
  assign n38943 = ~n6438 & n38942 ;
  assign n38944 = n6818 | n38943 ;
  assign n38945 = n38941 & ~n38944 ;
  assign n38946 = n1256 & ~n1394 ;
  assign n38947 = n3981 | n10080 ;
  assign n38948 = ~n38946 & n38947 ;
  assign n38949 = n8430 ^ n5574 ^ 1'b0 ;
  assign n38951 = n22981 ^ n367 ^ n32 ;
  assign n38950 = ~n7486 & n33984 ;
  assign n38952 = n38951 ^ n38950 ^ 1'b0 ;
  assign n38953 = n38952 ^ n4895 ^ 1'b0 ;
  assign n38954 = ~n37413 & n38953 ;
  assign n38955 = n13052 & n19639 ;
  assign n38956 = n38955 ^ n3260 ^ 1'b0 ;
  assign n38957 = n4904 & ~n18663 ;
  assign n38958 = ~n25951 & n38957 ;
  assign n38959 = n35483 & ~n38958 ;
  assign n38960 = ~n3426 & n38959 ;
  assign n38961 = ~n24779 & n38960 ;
  assign n38962 = n16309 ^ n7369 ^ 1'b0 ;
  assign n38963 = n1174 & ~n8519 ;
  assign n38964 = n30445 ^ n19904 ^ 1'b0 ;
  assign n38965 = n15521 | n18725 ;
  assign n38966 = n2130 & ~n2212 ;
  assign n38967 = n38966 ^ n3219 ^ 1'b0 ;
  assign n38968 = n13108 ^ n1214 ^ 1'b0 ;
  assign n38969 = n35644 & ~n38968 ;
  assign n38970 = n7109 & n17139 ;
  assign n38971 = n6094 & ~n20890 ;
  assign n38972 = n38970 & n38971 ;
  assign n38973 = n15851 | n19776 ;
  assign n38974 = n38973 ^ n8508 ^ 1'b0 ;
  assign n38975 = n21796 & n38974 ;
  assign n38976 = ~n5386 & n38975 ;
  assign n38977 = n9424 & n38976 ;
  assign n38978 = n4424 | n10375 ;
  assign n38979 = n38977 & ~n38978 ;
  assign n38980 = n29206 ^ n13091 ^ 1'b0 ;
  assign n38981 = n38980 ^ n5293 ^ 1'b0 ;
  assign n38982 = n20446 | n38981 ;
  assign n38983 = n11609 | n31068 ;
  assign n38984 = n28363 ^ n8360 ^ 1'b0 ;
  assign n38985 = ~n15551 & n38984 ;
  assign n38986 = n10078 & ~n38985 ;
  assign n38987 = n29878 ^ n24089 ^ 1'b0 ;
  assign n38988 = n17247 & ~n38987 ;
  assign n38989 = ~n7601 & n38988 ;
  assign n38990 = n13592 ^ n3290 ^ 1'b0 ;
  assign n38991 = n2707 & ~n38990 ;
  assign n38992 = n38991 ^ n10635 ^ 1'b0 ;
  assign n38993 = n2738 | n2881 ;
  assign n38994 = n11289 | n38993 ;
  assign n38995 = n38994 ^ n228 ^ 1'b0 ;
  assign n38996 = n31988 ^ n8489 ^ 1'b0 ;
  assign n38997 = n38995 & ~n38996 ;
  assign n38998 = n38997 ^ n12309 ^ 1'b0 ;
  assign n38999 = ~n1437 & n29091 ;
  assign n39000 = n38999 ^ n13766 ^ 1'b0 ;
  assign n39002 = n30010 ^ n10505 ^ 1'b0 ;
  assign n39003 = n37152 & ~n39002 ;
  assign n39001 = n12472 | n25081 ;
  assign n39004 = n39003 ^ n39001 ^ 1'b0 ;
  assign n39005 = n8829 & n37524 ;
  assign n39006 = ~n31914 & n39005 ;
  assign n39007 = n7589 ^ n7510 ^ 1'b0 ;
  assign n39008 = n39007 ^ n32935 ^ 1'b0 ;
  assign n39009 = n18937 & ~n39008 ;
  assign n39010 = n297 & ~n12395 ;
  assign n39011 = ~n39009 & n39010 ;
  assign n39012 = n15876 ^ n14043 ^ n2568 ;
  assign n39013 = n16529 & ~n18030 ;
  assign n39014 = n15117 ^ n8053 ^ 1'b0 ;
  assign n39015 = n20625 & n39014 ;
  assign n39016 = n4924 ^ n2096 ^ 1'b0 ;
  assign n39017 = n39016 ^ n38986 ^ 1'b0 ;
  assign n39018 = n27151 & n39017 ;
  assign n39019 = n1192 | n3447 ;
  assign n39020 = n5231 & ~n13068 ;
  assign n39021 = n345 & n39020 ;
  assign n39022 = ~n3941 & n39021 ;
  assign n39023 = n39022 ^ n18314 ^ 1'b0 ;
  assign n39024 = ( n14902 & n27406 ) | ( n14902 & ~n28407 ) | ( n27406 & ~n28407 ) ;
  assign n39025 = n39024 ^ n13197 ^ 1'b0 ;
  assign n39026 = n3123 | n33933 ;
  assign n39027 = n3793 ^ n1539 ^ 1'b0 ;
  assign n39028 = ~n36370 & n39027 ;
  assign n39029 = n30682 & n39028 ;
  assign n39030 = ~n39028 & n39029 ;
  assign n39031 = ~n7819 & n29109 ;
  assign n39032 = n1793 ^ n279 ^ 1'b0 ;
  assign n39033 = n12888 & ~n39032 ;
  assign n39034 = n33644 & n39033 ;
  assign n39035 = n3527 & n39034 ;
  assign n39039 = n10984 & n20373 ;
  assign n39036 = n977 & n5180 ;
  assign n39037 = n13634 & n39036 ;
  assign n39038 = n84 | n39037 ;
  assign n39040 = n39039 ^ n39038 ^ 1'b0 ;
  assign n39041 = n2923 | n36626 ;
  assign n39042 = n33397 | n39041 ;
  assign n39043 = ~n5923 & n19921 ;
  assign n39044 = ~n13204 & n39043 ;
  assign n39045 = n5046 & ~n39044 ;
  assign n39046 = ~n39042 & n39045 ;
  assign n39047 = n14554 & ~n27869 ;
  assign n39048 = n39047 ^ n16289 ^ 1'b0 ;
  assign n39049 = ~n10191 & n39048 ;
  assign n39050 = ~n21423 & n39049 ;
  assign n39051 = n39050 ^ n16487 ^ 1'b0 ;
  assign n39052 = n26787 ^ n10729 ^ 1'b0 ;
  assign n39053 = n1470 & ~n2825 ;
  assign n39054 = ~n18624 & n32979 ;
  assign n39055 = ~n27755 & n39054 ;
  assign n39056 = n9838 | n15279 ;
  assign n39057 = n39056 ^ n7442 ^ 1'b0 ;
  assign n39058 = n7155 | n33794 ;
  assign n39059 = ~n506 & n11158 ;
  assign n39060 = n1235 & n1950 ;
  assign n39061 = n39060 ^ n880 ^ 1'b0 ;
  assign n39062 = n5747 | n16231 ;
  assign n39063 = n39062 ^ n68 ^ 1'b0 ;
  assign n39064 = ~n374 & n10357 ;
  assign n39065 = n39064 ^ n4191 ^ 1'b0 ;
  assign n39066 = n10603 | n27495 ;
  assign n39067 = n26283 ^ n12225 ^ 1'b0 ;
  assign n39068 = n9120 & n39067 ;
  assign n39069 = n38479 ^ n24101 ^ 1'b0 ;
  assign n39070 = n34419 & ~n38582 ;
  assign n39071 = n9344 ^ n1937 ^ 1'b0 ;
  assign n39072 = ~n8475 & n39071 ;
  assign n39073 = n39072 ^ n19745 ^ 1'b0 ;
  assign n39074 = n3698 | n27100 ;
  assign n39075 = n39073 | n39074 ;
  assign n39076 = n125 | n984 ;
  assign n39077 = n36670 ^ n11065 ^ 1'b0 ;
  assign n39078 = n4652 & ~n39077 ;
  assign n39079 = n19145 ^ n1497 ^ 1'b0 ;
  assign n39080 = n6019 & n39079 ;
  assign n39081 = n2506 & ~n11622 ;
  assign n39082 = n20570 & n39081 ;
  assign n39083 = n1310 & n10959 ;
  assign n39084 = n488 & n37027 ;
  assign n39085 = n7540 & ~n34447 ;
  assign n39086 = n11288 ^ n5043 ^ 1'b0 ;
  assign n39087 = n24776 & ~n39086 ;
  assign n39088 = n17284 ^ n5894 ^ 1'b0 ;
  assign n39089 = n5701 & n39088 ;
  assign n39090 = n22601 ^ n10257 ^ 1'b0 ;
  assign n39091 = n35021 | n39090 ;
  assign n39092 = n3032 & ~n26725 ;
  assign n39093 = n39092 ^ n1863 ^ 1'b0 ;
  assign n39094 = n35791 ^ n20674 ^ 1'b0 ;
  assign n39095 = n12992 | n39094 ;
  assign n39096 = n88 | n39095 ;
  assign n39097 = ~n977 & n39096 ;
  assign n39098 = n26110 & n37000 ;
  assign n39099 = n39098 ^ n33484 ^ 1'b0 ;
  assign n39100 = n419 & ~n1954 ;
  assign n39101 = n382 & ~n33467 ;
  assign n39102 = n7876 | n39101 ;
  assign n39104 = n6687 & ~n22453 ;
  assign n39103 = n1430 | n15475 ;
  assign n39105 = n39104 ^ n39103 ^ 1'b0 ;
  assign n39106 = n21421 ^ n16646 ^ 1'b0 ;
  assign n39107 = n39105 | n39106 ;
  assign n39108 = n17385 ^ n5465 ^ 1'b0 ;
  assign n39109 = ~n22823 & n39108 ;
  assign n39110 = n1778 & n39109 ;
  assign n39111 = n1458 & n5826 ;
  assign n39112 = n15502 & n39111 ;
  assign n39113 = n39112 ^ n16454 ^ 1'b0 ;
  assign n39115 = n3459 & ~n37539 ;
  assign n39114 = n29066 & n30681 ;
  assign n39116 = n39115 ^ n39114 ^ n33499 ;
  assign n39117 = n4319 & ~n17791 ;
  assign n39118 = n12967 ^ n2433 ^ 1'b0 ;
  assign n39119 = ~n15326 & n39118 ;
  assign n39120 = ~n22851 & n39119 ;
  assign n39121 = n39120 ^ n28833 ^ 1'b0 ;
  assign n39126 = n517 & n7721 ;
  assign n39127 = n6595 & n39126 ;
  assign n39128 = n29684 & ~n39127 ;
  assign n39129 = n6280 | n39128 ;
  assign n39130 = n39129 ^ n20035 ^ 1'b0 ;
  assign n39122 = n2900 & n3408 ;
  assign n39123 = n39122 ^ n6445 ^ 1'b0 ;
  assign n39124 = ~n7118 & n39123 ;
  assign n39125 = n39124 ^ n2136 ^ 1'b0 ;
  assign n39131 = n39130 ^ n39125 ^ 1'b0 ;
  assign n39132 = n39131 ^ n21883 ^ 1'b0 ;
  assign n39133 = n16217 ^ n1600 ^ 1'b0 ;
  assign n39134 = n19088 ^ n17787 ^ 1'b0 ;
  assign n39135 = n39133 | n39134 ;
  assign n39136 = n39135 ^ n1764 ^ 1'b0 ;
  assign n39137 = n26426 ^ n2851 ^ n364 ;
  assign n39138 = n19107 & ~n22702 ;
  assign n39139 = n405 | n39138 ;
  assign n39140 = ~n23093 & n39139 ;
  assign n39141 = n3423 & ~n14333 ;
  assign n39142 = n39141 ^ n1195 ^ 1'b0 ;
  assign n39143 = n1754 | n12200 ;
  assign n39144 = n12758 & n39143 ;
  assign n39145 = n39144 ^ n2751 ^ 1'b0 ;
  assign n39146 = n3251 & n8829 ;
  assign n39147 = n8598 ^ n8408 ^ 1'b0 ;
  assign n39148 = n749 & ~n39147 ;
  assign n39149 = n39148 ^ n19642 ^ 1'b0 ;
  assign n39150 = n21217 ^ n2095 ^ 1'b0 ;
  assign n39151 = ~n364 & n20484 ;
  assign n39152 = n11849 & ~n16990 ;
  assign n39157 = n6256 ^ n3719 ^ 1'b0 ;
  assign n39158 = n8215 | n39157 ;
  assign n39153 = n7844 ^ n757 ^ 1'b0 ;
  assign n39154 = ~n25987 & n39153 ;
  assign n39155 = ~n14444 & n39154 ;
  assign n39156 = n1300 & ~n39155 ;
  assign n39159 = n39158 ^ n39156 ^ 1'b0 ;
  assign n39160 = n12709 | n22479 ;
  assign n39161 = n34397 ^ n3134 ^ 1'b0 ;
  assign n39162 = n14657 ^ n5549 ^ 1'b0 ;
  assign n39163 = ~n9399 & n39162 ;
  assign n39164 = n6698 | n14946 ;
  assign n39165 = n39164 ^ n2394 ^ 1'b0 ;
  assign n39166 = n495 & ~n39165 ;
  assign n39167 = n10123 | n32346 ;
  assign n39168 = n39167 ^ n28613 ^ n12951 ;
  assign n39169 = n17495 ^ n2795 ^ 1'b0 ;
  assign n39170 = n25719 ^ n11882 ^ 1'b0 ;
  assign n39171 = ~n39169 & n39170 ;
  assign n39172 = n257 & n34953 ;
  assign n39173 = n39172 ^ n7679 ^ 1'b0 ;
  assign n39174 = ~n14 & n39173 ;
  assign n39175 = ~n38651 & n39174 ;
  assign n39176 = n21376 ^ n13156 ^ 1'b0 ;
  assign n39177 = n8720 & ~n39176 ;
  assign n39178 = n17717 ^ n7189 ^ 1'b0 ;
  assign n39179 = n22387 ^ n2432 ^ 1'b0 ;
  assign n39180 = n39178 | n39179 ;
  assign n39181 = n20362 ^ n5200 ^ 1'b0 ;
  assign n39182 = n5135 & n8589 ;
  assign n39183 = ~n37359 & n39182 ;
  assign n39184 = n39183 ^ n18049 ^ 1'b0 ;
  assign n39185 = n6649 & n39184 ;
  assign n39186 = n3481 | n39185 ;
  assign n39187 = ~n3964 & n9091 ;
  assign n39188 = n39187 ^ n34979 ^ 1'b0 ;
  assign n39189 = n5802 & ~n30080 ;
  assign n39190 = n39189 ^ n748 ^ 1'b0 ;
  assign n39191 = n23913 & ~n29503 ;
  assign n39192 = n28115 ^ n24439 ^ 1'b0 ;
  assign n39194 = n19484 ^ n1704 ^ 1'b0 ;
  assign n39193 = ~n32646 & n34038 ;
  assign n39195 = n39194 ^ n39193 ^ 1'b0 ;
  assign n39196 = ~n5819 & n19149 ;
  assign n39197 = n9231 & n17974 ;
  assign n39198 = n39197 ^ n5456 ^ 1'b0 ;
  assign n39199 = n13554 | n32103 ;
  assign n39200 = ~n19990 & n31200 ;
  assign n39201 = n15591 & ~n16906 ;
  assign n39202 = ~n3633 & n7299 ;
  assign n39203 = ~n16102 & n39202 ;
  assign n39204 = n39203 ^ n7617 ^ 1'b0 ;
  assign n39205 = n227 & n4740 ;
  assign n39206 = ~n19364 & n27435 ;
  assign n39207 = ~n924 & n16791 ;
  assign n39208 = n10174 ^ n8690 ^ n3692 ;
  assign n39209 = n26785 & ~n39208 ;
  assign n39210 = n7773 ^ n6392 ^ n1227 ;
  assign n39211 = n13163 ^ n10621 ^ n7805 ;
  assign n39212 = n39210 & ~n39211 ;
  assign n39213 = n4791 ^ n2853 ^ 1'b0 ;
  assign n39214 = ~n1283 & n2984 ;
  assign n39215 = ~n11155 & n39214 ;
  assign n39216 = ~n34192 & n39215 ;
  assign n39217 = ~n291 & n560 ;
  assign n39218 = ~n39216 & n39217 ;
  assign n39219 = n8559 & n25795 ;
  assign n39220 = n10009 & n39219 ;
  assign n39221 = n1822 | n31045 ;
  assign n39222 = n14701 & ~n32615 ;
  assign n39223 = n39222 ^ n895 ^ 1'b0 ;
  assign n39224 = n12804 ^ n6521 ^ 1'b0 ;
  assign n39225 = n36702 ^ n32114 ^ n6247 ;
  assign n39226 = n14960 & n21395 ;
  assign n39228 = n11479 ^ n942 ^ 1'b0 ;
  assign n39229 = n501 & ~n39228 ;
  assign n39230 = ( n10219 & n29155 ) | ( n10219 & n39229 ) | ( n29155 & n39229 ) ;
  assign n39227 = n20649 & ~n33088 ;
  assign n39231 = n39230 ^ n39227 ^ 1'b0 ;
  assign n39233 = n18423 ^ n10443 ^ 1'b0 ;
  assign n39234 = n29647 & n39233 ;
  assign n39232 = n24404 ^ n16283 ^ 1'b0 ;
  assign n39235 = n39234 ^ n39232 ^ 1'b0 ;
  assign n39236 = n5936 | n9437 ;
  assign n39237 = n14955 | n30920 ;
  assign n39238 = n64 | n684 ;
  assign n39239 = n9737 & ~n16370 ;
  assign n39240 = n39239 ^ n912 ^ 1'b0 ;
  assign n39241 = n29268 & n39240 ;
  assign n39242 = ~n3447 & n20192 ;
  assign n39243 = n39242 ^ n23149 ^ 1'b0 ;
  assign n39244 = n38097 ^ n410 ^ 1'b0 ;
  assign n39245 = n39243 & n39244 ;
  assign n39246 = n9281 & ~n21569 ;
  assign n39247 = n1370 ^ n292 ^ 1'b0 ;
  assign n39248 = n7917 & ~n39247 ;
  assign n39249 = n804 & ~n2394 ;
  assign n39250 = n39249 ^ n24142 ^ 1'b0 ;
  assign n39251 = n22185 & ~n39250 ;
  assign n39252 = n13678 ^ n5400 ^ n1732 ;
  assign n39253 = n15582 & ~n39252 ;
  assign n39254 = ~n4769 & n14311 ;
  assign n39255 = ~n977 & n14155 ;
  assign n39256 = n39255 ^ n3389 ^ 1'b0 ;
  assign n39257 = n4543 | n39256 ;
  assign n39258 = n39257 ^ n1455 ^ 1'b0 ;
  assign n39259 = n9163 | n39258 ;
  assign n39260 = n26316 ^ n19158 ^ 1'b0 ;
  assign n39261 = ~n741 & n3131 ;
  assign n39262 = n17844 ^ n7590 ^ 1'b0 ;
  assign n39263 = ~n888 & n39262 ;
  assign n39266 = n6508 ^ n1742 ^ 1'b0 ;
  assign n39267 = n2552 | n39266 ;
  assign n39264 = ~n385 & n20116 ;
  assign n39265 = ~n6286 & n39264 ;
  assign n39268 = n39267 ^ n39265 ^ 1'b0 ;
  assign n39269 = n32778 ^ n9051 ^ 1'b0 ;
  assign n39270 = n4636 | n5856 ;
  assign n39271 = n39270 ^ n3698 ^ 1'b0 ;
  assign n39272 = n34859 ^ n5241 ^ 1'b0 ;
  assign n39273 = n39271 | n39272 ;
  assign n39274 = n29037 ^ n8869 ^ 1'b0 ;
  assign n39275 = n4751 | n37253 ;
  assign n39276 = n39275 ^ n18205 ^ 1'b0 ;
  assign n39277 = n39276 ^ n12540 ^ 1'b0 ;
  assign n39278 = n19625 ^ n10309 ^ 1'b0 ;
  assign n39279 = n278 & n23599 ;
  assign n39280 = n26202 & n39279 ;
  assign n39281 = ~n11735 & n37961 ;
  assign n39282 = n241 | n758 ;
  assign n39283 = n39282 ^ n27923 ^ 1'b0 ;
  assign n39284 = n21535 | n30933 ;
  assign n39285 = n39283 & ~n39284 ;
  assign n39286 = n11028 & n19158 ;
  assign n39287 = n722 & n29159 ;
  assign n39288 = n39286 & n39287 ;
  assign n39289 = ~n2490 & n26360 ;
  assign n39290 = n2613 | n2617 ;
  assign n39294 = n7368 & n18798 ;
  assign n39295 = ~n1571 & n39294 ;
  assign n39291 = n1218 & n3036 ;
  assign n39292 = n14151 & n39291 ;
  assign n39293 = n8453 | n39292 ;
  assign n39296 = n39295 ^ n39293 ^ 1'b0 ;
  assign n39297 = n8291 & ~n11095 ;
  assign n39298 = n31070 & ~n32317 ;
  assign n39299 = ~n1137 & n11222 ;
  assign n39300 = n17484 | n39299 ;
  assign n39302 = ~n20269 & n25273 ;
  assign n39301 = ~n7667 & n8760 ;
  assign n39303 = n39302 ^ n39301 ^ 1'b0 ;
  assign n39304 = n35384 ^ n10145 ^ 1'b0 ;
  assign n39305 = n34942 & ~n39304 ;
  assign n39306 = n12808 & n33286 ;
  assign n39307 = n39306 ^ n8155 ^ 1'b0 ;
  assign n39308 = n4126 ^ n804 ^ 1'b0 ;
  assign n39309 = n36698 ^ n7676 ^ 1'b0 ;
  assign n39310 = n16913 | n27434 ;
  assign n39311 = n7194 | n21086 ;
  assign n39312 = n34100 ^ n29937 ^ 1'b0 ;
  assign n39313 = ~n39311 & n39312 ;
  assign n39314 = ~n7596 & n14955 ;
  assign n39315 = ( n5903 & n6728 ) | ( n5903 & ~n9693 ) | ( n6728 & ~n9693 ) ;
  assign n39316 = n1774 & ~n39315 ;
  assign n39317 = ~n25388 & n39316 ;
  assign n39318 = n1887 & n25711 ;
  assign n39319 = n4716 & n12095 ;
  assign n39320 = n32105 ^ n28103 ^ 1'b0 ;
  assign n39321 = ~n27742 & n39320 ;
  assign n39322 = n2288 | n6434 ;
  assign n39323 = n22733 ^ n13760 ^ 1'b0 ;
  assign n39324 = n10598 | n19202 ;
  assign n39325 = n39324 ^ n13425 ^ 1'b0 ;
  assign n39326 = ~n30978 & n39325 ;
  assign n39327 = ~n1226 & n39326 ;
  assign n39329 = ~n508 & n1523 ;
  assign n39328 = n13120 & ~n22348 ;
  assign n39330 = n39329 ^ n39328 ^ 1'b0 ;
  assign n39331 = n39330 ^ n14683 ^ 1'b0 ;
  assign n39332 = n14172 & n39331 ;
  assign n39333 = n1724 ^ n583 ^ 1'b0 ;
  assign n39334 = ~n37 & n39333 ;
  assign n39335 = n14394 & n39334 ;
  assign n39336 = ~n26287 & n39335 ;
  assign n39337 = ~n6272 & n17463 ;
  assign n39338 = n25118 & n29619 ;
  assign n39339 = n9504 ^ n2263 ^ 1'b0 ;
  assign n39340 = n29476 & n39339 ;
  assign n39341 = n2986 & n13158 ;
  assign n39342 = ~n39340 & n39341 ;
  assign n39343 = n31679 ^ n20512 ^ 1'b0 ;
  assign n39344 = n24125 & n39343 ;
  assign n39345 = n39344 ^ n6254 ^ 1'b0 ;
  assign n39346 = n6194 & ~n11178 ;
  assign n39347 = n22185 & n39346 ;
  assign n39348 = n958 ^ n509 ^ 1'b0 ;
  assign n39349 = ~n10603 & n27133 ;
  assign n39350 = n39348 & n39349 ;
  assign n39351 = n13909 ^ n661 ^ 1'b0 ;
  assign n39352 = n6846 & n39351 ;
  assign n39353 = ~n5688 & n39352 ;
  assign n39354 = n30711 ^ n228 ^ 1'b0 ;
  assign n39355 = ~n9419 & n32138 ;
  assign n39356 = n2018 | n33102 ;
  assign n39357 = n39356 ^ n32904 ^ 1'b0 ;
  assign n39358 = n32622 ^ n26203 ^ n158 ;
  assign n39359 = n13327 ^ n4823 ^ 1'b0 ;
  assign n39360 = n2865 & ~n21751 ;
  assign n39361 = n7144 & ~n17172 ;
  assign n39362 = n39361 ^ n9417 ^ 1'b0 ;
  assign n39363 = n9952 | n11308 ;
  assign n39364 = ~n5040 & n39363 ;
  assign n39365 = n958 & n6788 ;
  assign n39366 = n39365 ^ n1572 ^ 1'b0 ;
  assign n39367 = ~n6006 & n39366 ;
  assign n39368 = ~n16097 & n39367 ;
  assign n39369 = n3297 & ~n8135 ;
  assign n39370 = n39369 ^ n37282 ^ n23177 ;
  assign n39371 = n3071 & ~n10395 ;
  assign n39372 = n11604 | n39371 ;
  assign n39373 = n205 & n19854 ;
  assign n39374 = n39373 ^ n694 ^ 1'b0 ;
  assign n39375 = n39374 ^ n1418 ^ 1'b0 ;
  assign n39376 = n39375 ^ n1385 ^ 1'b0 ;
  assign n39377 = n35683 & n39376 ;
  assign n39378 = n39377 ^ n9384 ^ 1'b0 ;
  assign n39379 = n37382 ^ n22693 ^ 1'b0 ;
  assign n39380 = ~n2469 & n39379 ;
  assign n39382 = n20218 ^ n3423 ^ 1'b0 ;
  assign n39381 = n1431 & ~n8262 ;
  assign n39383 = n39382 ^ n39381 ^ 1'b0 ;
  assign n39384 = ~n2547 & n39383 ;
  assign n39385 = n28762 ^ n22832 ^ 1'b0 ;
  assign n39386 = n3260 & ~n39385 ;
  assign n39387 = n1070 | n35191 ;
  assign n39388 = n39387 ^ n2086 ^ 1'b0 ;
  assign n39389 = n21078 & n39388 ;
  assign n39390 = n13847 & n39389 ;
  assign n39391 = ~n8628 & n39390 ;
  assign n39392 = ~n6174 & n15197 ;
  assign n39393 = n37769 ^ n6190 ^ 1'b0 ;
  assign n39394 = n13204 | n39393 ;
  assign n39395 = n7685 | n8715 ;
  assign n39396 = n14235 ^ n2983 ^ 1'b0 ;
  assign n39397 = n39395 | n39396 ;
  assign n39398 = ~n21519 & n37053 ;
  assign n39399 = n39398 ^ n37031 ^ 1'b0 ;
  assign n39400 = n10675 ^ n9375 ^ 1'b0 ;
  assign n39401 = n11932 | n39400 ;
  assign n39402 = n8525 | n39401 ;
  assign n39403 = n39402 ^ n2122 ^ 1'b0 ;
  assign n39404 = ~n6419 & n39403 ;
  assign n39405 = n4448 | n10846 ;
  assign n39406 = n39405 ^ n2947 ^ 1'b0 ;
  assign n39407 = n35826 | n39406 ;
  assign n39408 = n34345 & ~n39407 ;
  assign n39409 = n1655 & ~n39408 ;
  assign n39410 = n10589 & n39409 ;
  assign n39411 = n10037 & ~n10728 ;
  assign n39412 = n9933 & ~n11071 ;
  assign n39413 = n39412 ^ n14572 ^ 1'b0 ;
  assign n39414 = n5206 | n36570 ;
  assign n39415 = n39414 ^ n14233 ^ 1'b0 ;
  assign n39416 = n39415 ^ n3591 ^ 1'b0 ;
  assign n39417 = n2975 & n13134 ;
  assign n39418 = n39417 ^ n8693 ^ 1'b0 ;
  assign n39419 = n4155 & ~n7289 ;
  assign n39420 = n6098 & n39419 ;
  assign n39421 = n2722 | n23197 ;
  assign n39422 = ~n227 & n3742 ;
  assign n39423 = n3663 & n39422 ;
  assign n39424 = n9053 | n39423 ;
  assign n39425 = n3164 | n31887 ;
  assign n39426 = n24228 ^ n1887 ^ 1'b0 ;
  assign n39427 = ~n596 & n5412 ;
  assign n39428 = n39426 & n39427 ;
  assign n39429 = n2031 | n39428 ;
  assign n39430 = n39429 ^ n11308 ^ 1'b0 ;
  assign n39431 = n9387 & n26596 ;
  assign n39432 = n24109 ^ n16746 ^ 1'b0 ;
  assign n39433 = n13964 ^ n2436 ^ 1'b0 ;
  assign n39434 = n23894 ^ n6758 ^ 1'b0 ;
  assign n39435 = n13730 | n39434 ;
  assign n39437 = n23152 ^ n8995 ^ 1'b0 ;
  assign n39438 = n21597 | n39437 ;
  assign n39436 = n52 & n31858 ;
  assign n39439 = n39438 ^ n39436 ^ 1'b0 ;
  assign n39440 = n235 & n3255 ;
  assign n39441 = n12034 ^ n1410 ^ 1'b0 ;
  assign n39442 = n547 & ~n39441 ;
  assign n39443 = n820 | n22561 ;
  assign n39444 = n13070 & ~n39443 ;
  assign n39445 = n39442 | n39444 ;
  assign n39446 = n18083 ^ n6644 ^ 1'b0 ;
  assign n39447 = n86 & n5152 ;
  assign n39448 = n17395 & n19921 ;
  assign n39449 = n44 & n7328 ;
  assign n39450 = ~n435 & n39449 ;
  assign n39451 = n32534 & ~n39450 ;
  assign n39452 = n4923 ^ n691 ^ 1'b0 ;
  assign n39453 = n9539 & n21614 ;
  assign n39454 = n7606 & n39453 ;
  assign n39455 = n39452 & n39454 ;
  assign n39456 = n6990 & n21066 ;
  assign n39457 = n15643 & n39456 ;
  assign n39458 = n11556 ^ n1053 ^ 1'b0 ;
  assign n39459 = n18780 & n39458 ;
  assign n39460 = n1987 & n39459 ;
  assign n39461 = n39460 ^ n29800 ^ 1'b0 ;
  assign n39462 = n6646 & ~n39461 ;
  assign n39463 = n22309 & ~n31556 ;
  assign n39464 = n8199 & ~n27964 ;
  assign n39465 = ~n2017 & n11920 ;
  assign n39466 = n39465 ^ n867 ^ 1'b0 ;
  assign n39467 = ~n228 & n17607 ;
  assign n39468 = n26235 & n39467 ;
  assign n39469 = n7191 ^ n1956 ^ 1'b0 ;
  assign n39470 = n39469 ^ n7153 ^ 1'b0 ;
  assign n39471 = ~n14774 & n28274 ;
  assign n39472 = n30662 & n39471 ;
  assign n39473 = n14901 & ~n39472 ;
  assign n39474 = n10971 ^ n945 ^ 1'b0 ;
  assign n39475 = n3194 & n39474 ;
  assign n39476 = n33720 ^ n17303 ^ 1'b0 ;
  assign n39477 = n17912 ^ n1936 ^ 1'b0 ;
  assign n39478 = n6440 & n39477 ;
  assign n39479 = ~n6610 & n38518 ;
  assign n39480 = n1375 & n7390 ;
  assign n39481 = ~n27870 & n39480 ;
  assign n39482 = ~n13139 & n39481 ;
  assign n39483 = n22118 ^ n18350 ^ 1'b0 ;
  assign n39484 = n9851 | n39483 ;
  assign n39485 = n18845 ^ n169 ^ 1'b0 ;
  assign n39486 = n39484 | n39485 ;
  assign n39487 = n21489 ^ n9424 ^ 1'b0 ;
  assign n39488 = n274 & n1979 ;
  assign n39489 = n14432 | n39488 ;
  assign n39490 = n8325 & ~n27870 ;
  assign n39491 = n5930 ^ n1285 ^ 1'b0 ;
  assign n39492 = n10731 & n12039 ;
  assign n39493 = n3080 | n4294 ;
  assign n39494 = n11421 | n39493 ;
  assign n39495 = n39494 ^ n18205 ^ 1'b0 ;
  assign n39496 = n2388 & n9240 ;
  assign n39497 = ~n3717 & n15632 ;
  assign n39498 = n39497 ^ n25012 ^ n3692 ;
  assign n39499 = n39498 ^ n22365 ^ 1'b0 ;
  assign n39500 = n2067 ^ n1946 ^ 1'b0 ;
  assign n39501 = n24106 | n39500 ;
  assign n39502 = n39501 ^ n6218 ^ 1'b0 ;
  assign n39503 = ~n15108 & n23105 ;
  assign n39504 = n16226 ^ n15595 ^ 1'b0 ;
  assign n39505 = n27085 | n39504 ;
  assign n39506 = n9989 | n36224 ;
  assign n39507 = n5228 & n39506 ;
  assign n39508 = n6644 & n21090 ;
  assign n39509 = n989 | n20255 ;
  assign n39510 = n39509 ^ n175 ^ 1'b0 ;
  assign n39511 = ~n14203 & n39510 ;
  assign n39512 = n2311 | n36192 ;
  assign n39513 = ~n10924 & n28282 ;
  assign n39514 = n39513 ^ n6417 ^ 1'b0 ;
  assign n39515 = n37405 & ~n38305 ;
  assign n39516 = n39514 & n39515 ;
  assign n39517 = n12028 | n19896 ;
  assign n39518 = n39517 ^ n32366 ^ 1'b0 ;
  assign n39519 = n38491 ^ n1254 ^ 1'b0 ;
  assign n39520 = ~n83 & n13414 ;
  assign n39521 = n3997 & ~n10303 ;
  assign n39522 = n12366 & n39521 ;
  assign n39523 = n1081 | n39522 ;
  assign n39524 = n5138 & n37936 ;
  assign n39525 = n39524 ^ n35296 ^ n19127 ;
  assign n39526 = n39525 ^ n29730 ^ 1'b0 ;
  assign n39527 = n15082 ^ n9416 ^ 1'b0 ;
  assign n39528 = n2917 | n8067 ;
  assign n39529 = n39528 ^ n13599 ^ 1'b0 ;
  assign n39530 = ( n3074 & ~n39527 ) | ( n3074 & n39529 ) | ( ~n39527 & n39529 ) ;
  assign n39531 = n1990 | n9096 ;
  assign n39532 = n39531 ^ n17175 ^ 1'b0 ;
  assign n39533 = ~n13056 & n14535 ;
  assign n39534 = n39533 ^ n6992 ^ 1'b0 ;
  assign n39535 = n3646 | n39534 ;
  assign n39536 = n1469 & n12325 ;
  assign n39537 = n1910 & ~n3631 ;
  assign n39538 = n39537 ^ n5561 ^ 1'b0 ;
  assign n39539 = n4724 | n39538 ;
  assign n39540 = n39539 ^ n13011 ^ 1'b0 ;
  assign n39541 = n2269 | n37657 ;
  assign n39542 = n17176 ^ n988 ^ 1'b0 ;
  assign n39543 = ~n9184 & n39542 ;
  assign n39544 = n39543 ^ n11476 ^ n8453 ;
  assign n39545 = n5927 & ~n33829 ;
  assign n39546 = n7944 & n39545 ;
  assign n39547 = n8179 | n39546 ;
  assign n39548 = n39547 ^ n4424 ^ 1'b0 ;
  assign n39549 = n39548 ^ n16162 ^ 1'b0 ;
  assign n39550 = ~n1112 & n21167 ;
  assign n39551 = n10357 ^ n556 ^ 1'b0 ;
  assign n39552 = ~n1789 & n3634 ;
  assign n39553 = n13682 | n39552 ;
  assign n39554 = n39553 ^ n6476 ^ 1'b0 ;
  assign n39555 = n37136 & ~n39554 ;
  assign n39556 = n2156 ^ n1786 ^ 1'b0 ;
  assign n39557 = n4983 & ~n39556 ;
  assign n39558 = n39557 ^ n16021 ^ 1'b0 ;
  assign n39559 = n11265 ^ n2776 ^ 1'b0 ;
  assign n39560 = n39559 ^ n31515 ^ n5775 ;
  assign n39562 = n12100 ^ n4204 ^ 1'b0 ;
  assign n39563 = ~n10583 & n39562 ;
  assign n39561 = ~n5583 & n6875 ;
  assign n39564 = n39563 ^ n39561 ^ 1'b0 ;
  assign n39565 = n11619 & n14719 ;
  assign n39566 = n792 ^ n34 ^ 1'b0 ;
  assign n39567 = n276 & ~n39566 ;
  assign n39568 = n1633 & n39567 ;
  assign n39569 = ~n20623 & n39568 ;
  assign n39570 = n7668 ^ n2107 ^ 1'b0 ;
  assign n39571 = n39570 ^ n8764 ^ 1'b0 ;
  assign n39572 = ~n39569 & n39571 ;
  assign n39573 = n39572 ^ n22301 ^ 1'b0 ;
  assign n39574 = ~n4025 & n39573 ;
  assign n39575 = n14609 ^ n3398 ^ 1'b0 ;
  assign n39576 = n68 | n22205 ;
  assign n39577 = ~n35652 & n39576 ;
  assign n39578 = n39575 & ~n39577 ;
  assign n39579 = ( n123 & n2696 ) | ( n123 & n38051 ) | ( n2696 & n38051 ) ;
  assign n39580 = n21613 & ~n38859 ;
  assign n39581 = ~n39579 & n39580 ;
  assign n39582 = ~n3311 & n3810 ;
  assign n39583 = n23913 & n39582 ;
  assign n39584 = ~n3137 & n16119 ;
  assign n39585 = n13644 ^ n11305 ^ 1'b0 ;
  assign n39586 = n3081 & n9801 ;
  assign n39587 = ~n25670 & n39586 ;
  assign n39590 = ~n832 & n36121 ;
  assign n39591 = n39590 ^ n9737 ^ 1'b0 ;
  assign n39588 = n20276 ^ n12331 ^ 1'b0 ;
  assign n39589 = n102 & n39588 ;
  assign n39592 = n39591 ^ n39589 ^ 1'b0 ;
  assign n39593 = n4969 & n16906 ;
  assign n39594 = n39593 ^ n19367 ^ 1'b0 ;
  assign n39595 = n1118 ^ n1048 ^ 1'b0 ;
  assign n39596 = ~n1718 & n39595 ;
  assign n39597 = n22711 ^ n492 ^ 1'b0 ;
  assign n39598 = n1896 & n21953 ;
  assign n39599 = n6120 | n6527 ;
  assign n39600 = n9747 & ~n39599 ;
  assign n39601 = n13295 & n39600 ;
  assign n39602 = ~n5317 & n12704 ;
  assign n39603 = ~n7770 & n39602 ;
  assign n39604 = n39601 & n39603 ;
  assign n39605 = n39604 ^ n1676 ^ 1'b0 ;
  assign n39606 = n1742 | n39605 ;
  assign n39607 = n18209 & n20467 ;
  assign n39608 = n39607 ^ n832 ^ 1'b0 ;
  assign n39609 = ( ~n4088 & n8917 ) | ( ~n4088 & n38031 ) | ( n8917 & n38031 ) ;
  assign n39610 = n21571 ^ n15901 ^ 1'b0 ;
  assign n39614 = n15426 ^ n1774 ^ 1'b0 ;
  assign n39615 = n8630 & n39614 ;
  assign n39611 = n3118 & ~n15779 ;
  assign n39612 = n39611 ^ n27595 ^ 1'b0 ;
  assign n39613 = ~n29650 & n39612 ;
  assign n39616 = n39615 ^ n39613 ^ 1'b0 ;
  assign n39617 = n22097 ^ n14970 ^ 1'b0 ;
  assign n39618 = ~n30196 & n39617 ;
  assign n39619 = n29693 & ~n37523 ;
  assign n39620 = n26220 ^ n3032 ^ 1'b0 ;
  assign n39622 = n12054 ^ n8991 ^ 1'b0 ;
  assign n39621 = n8876 & ~n36570 ;
  assign n39623 = n39622 ^ n39621 ^ 1'b0 ;
  assign n39624 = n325 | n39623 ;
  assign n39625 = n8630 | n39624 ;
  assign n39626 = n39625 ^ n12160 ^ 1'b0 ;
  assign n39627 = ( ~n9594 & n21810 ) | ( ~n9594 & n34440 ) | ( n21810 & n34440 ) ;
  assign n39628 = n5551 | n25197 ;
  assign n39629 = n22248 & ~n22783 ;
  assign n39630 = n39629 ^ n34069 ^ n14388 ;
  assign n39631 = n39630 ^ n31417 ^ 1'b0 ;
  assign n39632 = n26741 ^ n759 ^ 1'b0 ;
  assign n39633 = n26142 ^ n14483 ^ n3784 ;
  assign n39634 = n20568 ^ n17008 ^ n5846 ;
  assign n39635 = n39576 ^ n2948 ^ 1'b0 ;
  assign n39636 = n19831 ^ n883 ^ 1'b0 ;
  assign n39637 = n3277 & ~n16072 ;
  assign n39638 = ~n8639 & n20021 ;
  assign n39639 = ~n6419 & n39638 ;
  assign n39640 = n1571 | n39639 ;
  assign n39641 = n39640 ^ n11923 ^ 1'b0 ;
  assign n39642 = ~n23582 & n29950 ;
  assign n39643 = n1577 & ~n17572 ;
  assign n39644 = n10095 & n32418 ;
  assign n39645 = n5727 & ~n24056 ;
  assign n39646 = n83 & n2303 ;
  assign n39647 = n1722 & ~n39646 ;
  assign n39648 = n8316 & ~n15147 ;
  assign n39649 = ~n12628 & n39648 ;
  assign n39650 = n34901 & ~n39649 ;
  assign n39651 = ~n31108 & n39650 ;
  assign n39652 = ~n7449 & n29290 ;
  assign n39653 = n39652 ^ n7508 ^ 1'b0 ;
  assign n39654 = ~n11204 & n27665 ;
  assign n39655 = n39654 ^ n17542 ^ 1'b0 ;
  assign n39656 = n4505 & n9461 ;
  assign n39657 = n15864 | n39656 ;
  assign n39658 = n39657 ^ n6709 ^ 1'b0 ;
  assign n39659 = n18621 ^ n2304 ^ 1'b0 ;
  assign n39660 = ~n2125 & n25121 ;
  assign n39661 = n19654 ^ n10124 ^ 1'b0 ;
  assign n39662 = ~n32461 & n39661 ;
  assign n39666 = ~n3337 & n7001 ;
  assign n39667 = n3337 & n39666 ;
  assign n39668 = n39667 ^ n688 ^ 1'b0 ;
  assign n39663 = ~n294 & n2953 ;
  assign n39664 = n294 & n39663 ;
  assign n39665 = n39664 ^ n294 ^ 1'b0 ;
  assign n39669 = n39668 ^ n39665 ^ 1'b0 ;
  assign n39670 = n31433 & n39669 ;
  assign n39671 = n24661 ^ n23228 ^ n3576 ;
  assign n39672 = n39670 & n39671 ;
  assign n39673 = n17283 ^ n12877 ^ n6383 ;
  assign n39674 = n14398 | n30433 ;
  assign n39675 = n39674 ^ n9835 ^ 1'b0 ;
  assign n39676 = n15309 | n21535 ;
  assign n39677 = n5660 & n7907 ;
  assign n39678 = ~n35239 & n37320 ;
  assign n39679 = n8389 ^ n646 ^ 1'b0 ;
  assign n39680 = n7353 & n39679 ;
  assign n39681 = n20954 ^ n2109 ^ 1'b0 ;
  assign n39682 = n29373 & n30498 ;
  assign n39683 = ~n307 & n16099 ;
  assign n39684 = n15967 & n36133 ;
  assign n39685 = ~n31935 & n39684 ;
  assign n39686 = ~n3822 & n8312 ;
  assign n39687 = n39686 ^ n719 ^ 1'b0 ;
  assign n39688 = n4400 & ~n17807 ;
  assign n39689 = n38608 ^ n19064 ^ 1'b0 ;
  assign n39690 = n8281 | n39689 ;
  assign n39691 = n11804 & ~n21167 ;
  assign n39692 = n39691 ^ n24008 ^ 1'b0 ;
  assign n39693 = n27392 ^ n6610 ^ 1'b0 ;
  assign n39694 = n9079 & ~n30061 ;
  assign n39695 = n310 & n11808 ;
  assign n39696 = n4197 | n27491 ;
  assign n39697 = n17694 & ~n39696 ;
  assign n39698 = n11429 & ~n39697 ;
  assign n39699 = n33751 ^ n9422 ^ 1'b0 ;
  assign n39700 = ~n22085 & n27546 ;
  assign n39701 = n12692 & n16199 ;
  assign n39702 = n39701 ^ n2018 ^ 1'b0 ;
  assign n39703 = n26595 ^ n3150 ^ 1'b0 ;
  assign n39704 = n39702 & n39703 ;
  assign n39705 = n4210 & ~n5317 ;
  assign n39706 = ~n6667 & n39705 ;
  assign n39707 = n39706 ^ n29231 ^ 1'b0 ;
  assign n39708 = n9675 & n33521 ;
  assign n39709 = ~n6462 & n25197 ;
  assign n39710 = n12754 & ~n36495 ;
  assign n39711 = n1449 | n14549 ;
  assign n39712 = ~n11245 & n35661 ;
  assign n39713 = n39712 ^ n10851 ^ 1'b0 ;
  assign n39714 = n39713 ^ n28970 ^ 1'b0 ;
  assign n39715 = n39714 ^ n34839 ^ 1'b0 ;
  assign n39716 = ~n4029 & n39715 ;
  assign n39717 = n14590 | n35121 ;
  assign n39718 = n5024 ^ n294 ^ 1'b0 ;
  assign n39719 = n5872 & ~n39718 ;
  assign n39720 = n39719 ^ n21349 ^ 1'b0 ;
  assign n39722 = n227 & n25337 ;
  assign n39721 = n16377 | n35306 ;
  assign n39723 = n39722 ^ n39721 ^ 1'b0 ;
  assign n39724 = n2546 & ~n39723 ;
  assign n39725 = n18654 ^ n13807 ^ n5083 ;
  assign n39726 = n39725 ^ n534 ^ 1'b0 ;
  assign n39727 = n17477 & n17557 ;
  assign n39728 = ~n10282 & n39727 ;
  assign n39729 = ~n33619 & n39728 ;
  assign n39730 = ~n11192 & n39729 ;
  assign n39731 = n12954 | n23076 ;
  assign n39732 = n15121 & ~n39731 ;
  assign n39733 = n16898 ^ n10382 ^ 1'b0 ;
  assign n39734 = ~n6159 & n39733 ;
  assign n39735 = n11415 ^ n5394 ^ 1'b0 ;
  assign n39736 = n25027 ^ n185 ^ 1'b0 ;
  assign n39737 = ~n15081 & n39736 ;
  assign n39738 = ~n9891 & n12899 ;
  assign n39739 = ~n5892 & n39738 ;
  assign n39740 = n28833 ^ n4966 ^ 1'b0 ;
  assign n39741 = n5286 & ~n39740 ;
  assign n39742 = ~n10403 & n39741 ;
  assign n39743 = n39742 ^ n1080 ^ 1'b0 ;
  assign n39744 = n39739 & ~n39743 ;
  assign n39745 = n39602 ^ n19332 ^ 1'b0 ;
  assign n39746 = ~n31651 & n35635 ;
  assign n39747 = ~n13892 & n39746 ;
  assign n39748 = n14464 ^ n3262 ^ 1'b0 ;
  assign n39749 = n32357 & n39748 ;
  assign n39750 = n39749 ^ n29267 ^ 1'b0 ;
  assign n39751 = ~n25175 & n39750 ;
  assign n39752 = ~n2829 & n23819 ;
  assign n39753 = n23401 & n39752 ;
  assign n39754 = n3688 | n23012 ;
  assign n39755 = n38928 & ~n39754 ;
  assign n39756 = n39755 ^ n4840 ^ 1'b0 ;
  assign n39757 = n34909 ^ n1818 ^ 1'b0 ;
  assign n39758 = n6185 | n39757 ;
  assign n39763 = n784 | n3311 ;
  assign n39759 = n5990 & n14123 ;
  assign n39760 = n39759 ^ n15183 ^ 1'b0 ;
  assign n39761 = n39760 ^ n98 ^ 1'b0 ;
  assign n39762 = n5270 | n39761 ;
  assign n39764 = n39763 ^ n39762 ^ 1'b0 ;
  assign n39765 = n39764 ^ n39215 ^ 1'b0 ;
  assign n39766 = n1385 & n7472 ;
  assign n39767 = n39766 ^ n1520 ^ 1'b0 ;
  assign n39768 = n38567 | n39767 ;
  assign n39769 = n17269 ^ n6916 ^ 1'b0 ;
  assign n39770 = n13760 ^ n12709 ^ 1'b0 ;
  assign n39771 = ~n13735 & n39770 ;
  assign n39772 = n4010 & n39771 ;
  assign n39773 = ~n39769 & n39772 ;
  assign n39774 = n290 | n16013 ;
  assign n39775 = n18276 ^ n832 ^ 1'b0 ;
  assign n39776 = n23507 | n39775 ;
  assign n39777 = n39776 ^ n7483 ^ 1'b0 ;
  assign n39778 = n13791 ^ n9425 ^ 1'b0 ;
  assign n39779 = n4029 | n7845 ;
  assign n39780 = n3249 | n39779 ;
  assign n39781 = ~n34846 & n39780 ;
  assign n39782 = n20278 & n21075 ;
  assign n39783 = n39782 ^ n36203 ^ 1'b0 ;
  assign n39784 = n16024 ^ n330 ^ 1'b0 ;
  assign n39786 = n508 & n17506 ;
  assign n39785 = ~n7128 & n38975 ;
  assign n39787 = n39786 ^ n39785 ^ 1'b0 ;
  assign n39788 = n8749 | n16424 ;
  assign n39789 = n6608 & ~n6709 ;
  assign n39790 = n18962 & n39253 ;
  assign n39791 = n21029 | n36509 ;
  assign n39792 = n18531 & ~n39791 ;
  assign n39793 = n13930 ^ n4377 ^ 1'b0 ;
  assign n39794 = n19933 | n39793 ;
  assign n39796 = n6024 | n9139 ;
  assign n39797 = n18314 & n39796 ;
  assign n39795 = ~n5011 & n20780 ;
  assign n39798 = n39797 ^ n39795 ^ 1'b0 ;
  assign n39799 = ~n937 & n1205 ;
  assign n39800 = n39799 ^ n2717 ^ 1'b0 ;
  assign n39801 = n17583 & ~n36223 ;
  assign n39802 = ~n4833 & n33836 ;
  assign n39803 = n14813 ^ n10394 ^ n2426 ;
  assign n39804 = n22148 ^ n19822 ^ 1'b0 ;
  assign n39805 = n39804 ^ n445 ^ 1'b0 ;
  assign n39806 = n14647 & ~n34278 ;
  assign n39807 = n39806 ^ n22790 ^ 1'b0 ;
  assign n39808 = n6166 ^ n1178 ^ 1'b0 ;
  assign n39809 = n4797 & n39808 ;
  assign n39810 = n7739 & n13541 ;
  assign n39811 = ~n128 & n39810 ;
  assign n39812 = n15583 & ~n39811 ;
  assign n39813 = n11897 & ~n36984 ;
  assign n39814 = n39813 ^ n1792 ^ 1'b0 ;
  assign n39815 = n8777 | n11267 ;
  assign n39816 = n39815 ^ n36387 ^ 1'b0 ;
  assign n39817 = n7796 | n37822 ;
  assign n39818 = ~n3905 & n28535 ;
  assign n39819 = ~n5846 & n39818 ;
  assign n39820 = n2260 & n33760 ;
  assign n39821 = n22329 ^ n22134 ^ 1'b0 ;
  assign n39822 = ~n23450 & n39821 ;
  assign n39823 = ~n1467 & n22597 ;
  assign n39824 = n38535 ^ n14557 ^ 1'b0 ;
  assign n39825 = n3182 | n39824 ;
  assign n39826 = n21482 & n24573 ;
  assign n39827 = n5362 & n39826 ;
  assign n39828 = n2307 & ~n21766 ;
  assign n39829 = n39828 ^ n8887 ^ 1'b0 ;
  assign n39830 = n23982 | n39829 ;
  assign n39831 = n39830 ^ n11973 ^ 1'b0 ;
  assign n39832 = n1358 & n39831 ;
  assign n39833 = ~n13618 & n16262 ;
  assign n39834 = n3089 & n6389 ;
  assign n39835 = n39833 & ~n39834 ;
  assign n39836 = n4185 & n29717 ;
  assign n39837 = n39836 ^ n4281 ^ 1'b0 ;
  assign n39838 = n39837 ^ n33918 ^ 1'b0 ;
  assign n39839 = n3407 & ~n39838 ;
  assign n39840 = n28028 ^ n467 ^ 1'b0 ;
  assign n39841 = n26114 ^ n729 ^ 1'b0 ;
  assign n39842 = ~x11 & n28016 ;
  assign n39843 = n8106 | n37820 ;
  assign n39844 = n39843 ^ n21404 ^ 1'b0 ;
  assign n39845 = ~n9557 & n24443 ;
  assign n39846 = n39845 ^ n717 ^ 1'b0 ;
  assign n39847 = n23761 ^ n9329 ^ 1'b0 ;
  assign n39848 = n39846 | n39847 ;
  assign n39849 = ~n10930 & n11937 ;
  assign n39850 = n7449 & ~n13853 ;
  assign n39851 = n2969 | n4546 ;
  assign n39852 = n2572 & n39851 ;
  assign n39853 = n9010 & ~n19347 ;
  assign n39854 = n4193 & n20761 ;
  assign n39855 = n5194 ^ n2694 ^ 1'b0 ;
  assign n39856 = n39854 | n39855 ;
  assign n39857 = n5867 | n6492 ;
  assign n39858 = n36154 ^ n28306 ^ 1'b0 ;
  assign n39860 = n928 & n14608 ;
  assign n39861 = n39860 ^ n6371 ^ 1'b0 ;
  assign n39859 = n727 & ~n11621 ;
  assign n39862 = n39861 ^ n39859 ^ 1'b0 ;
  assign n39864 = ~n683 & n33695 ;
  assign n39865 = ~n13579 & n39864 ;
  assign n39863 = ~n3354 & n12102 ;
  assign n39866 = n39865 ^ n39863 ^ 1'b0 ;
  assign n39867 = n30544 ^ n8841 ^ 1'b0 ;
  assign n39868 = n16410 ^ n1626 ^ 1'b0 ;
  assign n39869 = ~n26776 & n39868 ;
  assign n39870 = n16424 ^ n11078 ^ 1'b0 ;
  assign n39877 = ~n244 & n4497 ;
  assign n39878 = n13613 & n39877 ;
  assign n39879 = n2117 & n39878 ;
  assign n39880 = n2424 & n17685 ;
  assign n39881 = ~n39879 & n39880 ;
  assign n39871 = n1205 & ~n11568 ;
  assign n39872 = n39871 ^ n20377 ^ 1'b0 ;
  assign n39873 = ~n1020 & n39872 ;
  assign n39874 = n20312 ^ n6944 ^ 1'b0 ;
  assign n39875 = ( n2455 & ~n39873 ) | ( n2455 & n39874 ) | ( ~n39873 & n39874 ) ;
  assign n39876 = n23975 & n39875 ;
  assign n39882 = n39881 ^ n39876 ^ 1'b0 ;
  assign n39883 = ~n15441 & n39882 ;
  assign n39884 = ~n30464 & n39524 ;
  assign n39885 = ~n36076 & n39884 ;
  assign n39886 = n6962 | n24338 ;
  assign n39887 = n39886 ^ n8497 ^ 1'b0 ;
  assign n39888 = n15056 & n23171 ;
  assign n39889 = n39888 ^ n16391 ^ 1'b0 ;
  assign n39890 = n5537 & n6776 ;
  assign n39891 = n39890 ^ n1011 ^ 1'b0 ;
  assign n39892 = n675 & n39891 ;
  assign n39893 = n16746 & ~n39892 ;
  assign n39894 = ~n10258 & n21069 ;
  assign n39895 = n39894 ^ n8518 ^ 1'b0 ;
  assign n39896 = ~n273 & n3997 ;
  assign n39897 = ~n2607 & n39896 ;
  assign n39898 = n21718 | n39897 ;
  assign n39899 = n26802 | n27228 ;
  assign n39900 = n39899 ^ n22201 ^ 1'b0 ;
  assign n39901 = n9596 ^ n7543 ^ 1'b0 ;
  assign n39902 = n13872 & n39901 ;
  assign n39903 = n21210 ^ n13778 ^ 1'b0 ;
  assign n39904 = n13263 & ~n30242 ;
  assign n39905 = ~n30808 & n39904 ;
  assign n39906 = n252 & ~n5917 ;
  assign n39907 = n8904 & ~n39906 ;
  assign n39908 = ~n16 & n292 ;
  assign n39909 = ( n6849 & n14991 ) | ( n6849 & n39908 ) | ( n14991 & n39908 ) ;
  assign n39910 = ~n13756 & n28525 ;
  assign n39911 = n39910 ^ n1958 ^ 1'b0 ;
  assign n39912 = n39911 ^ n2277 ^ 1'b0 ;
  assign n39913 = n29752 | n39912 ;
  assign n39914 = n34058 | n39913 ;
  assign n39915 = n2900 & ~n39914 ;
  assign n39916 = ~n39909 & n39915 ;
  assign n39917 = n7237 & n28306 ;
  assign n39918 = n10200 & n16296 ;
  assign n39919 = n11241 & n39918 ;
  assign n39920 = n25379 & n27687 ;
  assign n39921 = n39919 & n39920 ;
  assign n39922 = n16733 | n39921 ;
  assign n39923 = n2120 & n37229 ;
  assign n39924 = n11691 & n17069 ;
  assign n39925 = n8532 & n39924 ;
  assign n39926 = n3841 & n28697 ;
  assign n39927 = n3660 & n39926 ;
  assign n39928 = n814 & n6653 ;
  assign n39929 = n32389 ^ n3670 ^ 1'b0 ;
  assign n39930 = n4395 | n9392 ;
  assign n39931 = n14659 & n24260 ;
  assign n39932 = n5111 & n5948 ;
  assign n39933 = ~n24055 & n39932 ;
  assign n39934 = n39933 ^ n22119 ^ 1'b0 ;
  assign n39935 = n34131 ^ n1848 ^ 1'b0 ;
  assign n39936 = n39935 ^ n14064 ^ n11971 ;
  assign n39937 = n17610 & n36224 ;
  assign n39938 = ~n39936 & n39937 ;
  assign n39939 = ~n18065 & n28781 ;
  assign n39940 = n29237 ^ n8753 ^ 1'b0 ;
  assign n39941 = n1772 | n39940 ;
  assign n39942 = n1070 & ~n39941 ;
  assign n39943 = n39942 ^ n4231 ^ 1'b0 ;
  assign n39944 = ~n736 & n11680 ;
  assign n39945 = n39944 ^ n7208 ^ 1'b0 ;
  assign n39946 = n18264 ^ n10509 ^ n9682 ;
  assign n39947 = n8430 & ~n14736 ;
  assign n39948 = n39947 ^ n31935 ^ 1'b0 ;
  assign n39949 = n25095 ^ n185 ^ 1'b0 ;
  assign n39950 = n32037 & n39949 ;
  assign n39951 = n39950 ^ n17274 ^ 1'b0 ;
  assign n39952 = n9732 ^ n2122 ^ 1'b0 ;
  assign n39953 = n7734 & ~n36238 ;
  assign n39954 = n39953 ^ n24109 ^ 1'b0 ;
  assign n39955 = n35369 ^ n32195 ^ 1'b0 ;
  assign n39956 = n28543 & ~n39955 ;
  assign n39957 = n13635 & ~n34028 ;
  assign n39958 = n144 | n1793 ;
  assign n39959 = n39958 ^ n25763 ^ 1'b0 ;
  assign n39960 = n12497 & ~n13967 ;
  assign n39961 = n39960 ^ n14045 ^ n7554 ;
  assign n39962 = n1194 | n39961 ;
  assign n39963 = ~n8278 & n39962 ;
  assign n39964 = n4927 & ~n39963 ;
  assign n39965 = n9719 ^ n7548 ^ 1'b0 ;
  assign n39966 = n7578 & ~n39965 ;
  assign n39967 = n4158 & n39966 ;
  assign n39968 = n495 & ~n36414 ;
  assign n39969 = n21763 ^ n1899 ^ 1'b0 ;
  assign n39970 = n1255 & n39969 ;
  assign n39971 = n39970 ^ n8317 ^ 1'b0 ;
  assign n39972 = n39968 | n39971 ;
  assign n39973 = n745 | n39972 ;
  assign n39974 = n5637 & ~n20078 ;
  assign n39975 = n26593 & ~n39970 ;
  assign n39976 = n1842 ^ n748 ^ 1'b0 ;
  assign n39977 = n6315 & n19962 ;
  assign n39978 = n39977 ^ n16367 ^ 1'b0 ;
  assign n39979 = n34954 & n39978 ;
  assign n39980 = ~n21340 & n32676 ;
  assign n39981 = n39980 ^ n15390 ^ 1'b0 ;
  assign n39982 = n33046 ^ n26955 ^ 1'b0 ;
  assign n39983 = ~n144 & n39982 ;
  assign n39984 = n39983 ^ n7135 ^ 1'b0 ;
  assign n39985 = n4591 & ~n11122 ;
  assign n39986 = n14165 ^ n13608 ^ 1'b0 ;
  assign n39987 = n39985 & ~n39986 ;
  assign n39988 = n1311 & ~n8158 ;
  assign n39989 = ~n9659 & n39988 ;
  assign n39990 = n13043 ^ n5723 ^ 1'b0 ;
  assign n39991 = n13132 & ~n39990 ;
  assign n39992 = n23256 ^ n21870 ^ 1'b0 ;
  assign n39993 = n34876 & n39992 ;
  assign n39994 = n39993 ^ n37916 ^ 1'b0 ;
  assign n39995 = n31511 | n39994 ;
  assign n39996 = n20011 ^ n968 ^ 1'b0 ;
  assign n39997 = n799 & n39996 ;
  assign n39998 = ~n5597 & n39997 ;
  assign n39999 = n12345 ^ n6731 ^ 1'b0 ;
  assign n40000 = n19546 & n39999 ;
  assign n40001 = n3345 & ~n15598 ;
  assign n40002 = ( n113 & n4351 ) | ( n113 & ~n40001 ) | ( n4351 & ~n40001 ) ;
  assign n40003 = n17383 | n28687 ;
  assign n40004 = n40002 | n40003 ;
  assign n40008 = n2905 & ~n9286 ;
  assign n40005 = ~n1339 & n9560 ;
  assign n40006 = n26078 | n40005 ;
  assign n40007 = ~n29753 & n40006 ;
  assign n40009 = n40008 ^ n40007 ^ 1'b0 ;
  assign n40010 = ~n5923 & n14964 ;
  assign n40011 = ~n670 & n9245 ;
  assign n40012 = n7977 ^ n1428 ^ 1'b0 ;
  assign n40013 = n20556 & n40012 ;
  assign n40014 = n40013 ^ n34154 ^ 1'b0 ;
  assign n40015 = n4510 & n40014 ;
  assign n40016 = n5084 & ~n18716 ;
  assign n40017 = n40016 ^ n13330 ^ 1'b0 ;
  assign n40018 = n7269 & n27871 ;
  assign n40019 = n23463 & n23977 ;
  assign n40020 = n1893 & n40019 ;
  assign n40021 = n17574 | n26547 ;
  assign n40022 = n40021 ^ n26287 ^ 1'b0 ;
  assign n40023 = n1283 | n6466 ;
  assign n40024 = ~n40022 & n40023 ;
  assign n40025 = ~n128 & n4243 ;
  assign n40026 = ~n14622 & n40025 ;
  assign n40027 = n40026 ^ n18966 ^ 1'b0 ;
  assign n40028 = n24573 & n30749 ;
  assign n40029 = n8705 & n40028 ;
  assign n40030 = n24251 ^ n13483 ^ 1'b0 ;
  assign n40031 = n12186 ^ n1888 ^ 1'b0 ;
  assign n40032 = n28857 & ~n40031 ;
  assign n40033 = ( n3182 & ~n16703 ) | ( n3182 & n40032 ) | ( ~n16703 & n40032 ) ;
  assign n40034 = ~n7237 & n27255 ;
  assign n40035 = n3378 | n37048 ;
  assign n40036 = n6023 & n9661 ;
  assign n40037 = n12054 ^ n2261 ^ 1'b0 ;
  assign n40038 = n33898 ^ n7338 ^ 1'b0 ;
  assign n40039 = n37 & ~n40038 ;
  assign n40040 = ~n1421 & n40039 ;
  assign n40041 = n10069 & n25685 ;
  assign n40042 = n2738 & n40041 ;
  assign n40043 = n36656 ^ n5363 ^ n1212 ;
  assign n40044 = n2938 & n19561 ;
  assign n40045 = n20108 & n40044 ;
  assign n40046 = n40045 ^ n1357 ^ 1'b0 ;
  assign n40047 = ~n39133 & n40046 ;
  assign n40048 = n14954 ^ n3821 ^ 1'b0 ;
  assign n40049 = n20541 | n24631 ;
  assign n40050 = n32150 & ~n40049 ;
  assign n40051 = n12000 & ~n12349 ;
  assign n40052 = n11485 & n40051 ;
  assign n40053 = n23075 | n40052 ;
  assign n40054 = ~n7589 & n20401 ;
  assign n40055 = n40054 ^ n89 ^ 1'b0 ;
  assign n40056 = n18058 ^ n556 ^ 1'b0 ;
  assign n40057 = n40056 ^ n1426 ^ 1'b0 ;
  assign n40058 = n8843 & ~n39382 ;
  assign n40059 = n28087 ^ n25756 ^ n8628 ;
  assign n40060 = n30798 ^ n11123 ^ 1'b0 ;
  assign n40061 = n35769 & n40060 ;
  assign n40062 = ~n9169 & n39249 ;
  assign n40063 = n23297 ^ n15304 ^ n488 ;
  assign n40064 = n15200 & n40063 ;
  assign n40065 = n11116 & ~n30678 ;
  assign n40066 = n802 & n40065 ;
  assign n40067 = n38393 & ~n40066 ;
  assign n40068 = n2907 ^ n1593 ^ 1'b0 ;
  assign n40069 = n2155 & n40068 ;
  assign n40070 = n2723 & n8262 ;
  assign n40071 = n33125 & n37521 ;
  assign n40072 = n20348 | n24654 ;
  assign n40073 = n16987 | n40072 ;
  assign n40074 = n16365 & ~n40073 ;
  assign n40075 = n1598 | n37326 ;
  assign n40076 = n39148 ^ n2301 ^ 1'b0 ;
  assign n40077 = n11095 ^ n5336 ^ n340 ;
  assign n40078 = n20695 ^ n8326 ^ 1'b0 ;
  assign n40079 = n3374 ^ n1722 ^ 1'b0 ;
  assign n40080 = n8990 | n40079 ;
  assign n40081 = n8375 | n40080 ;
  assign n40082 = n767 ^ n77 ^ 1'b0 ;
  assign n40083 = n40082 ^ n16260 ^ 1'b0 ;
  assign n40084 = n7875 & n40083 ;
  assign n40085 = n1081 | n6721 ;
  assign n40086 = n40085 ^ n17117 ^ 1'b0 ;
  assign n40087 = n4093 & n8639 ;
  assign n40088 = n40087 ^ n7383 ^ 1'b0 ;
  assign n40089 = n60 | n40088 ;
  assign n40090 = n685 & ~n40089 ;
  assign n40091 = n31715 ^ n12873 ^ 1'b0 ;
  assign n40092 = n8069 | n40091 ;
  assign n40093 = n2785 | n40092 ;
  assign n40094 = n973 & ~n7933 ;
  assign n40095 = n729 | n40094 ;
  assign n40096 = n15956 ^ n4189 ^ 1'b0 ;
  assign n40097 = n3583 & n27165 ;
  assign n40098 = n40097 ^ n10320 ^ 1'b0 ;
  assign n40099 = n8181 & ~n40098 ;
  assign n40100 = n11997 ^ n10551 ^ 1'b0 ;
  assign n40101 = n530 | n1159 ;
  assign n40102 = n40101 ^ n5751 ^ 1'b0 ;
  assign n40103 = n14683 & ~n40102 ;
  assign n40104 = n20798 ^ n8664 ^ 1'b0 ;
  assign n40105 = n35371 & n40104 ;
  assign n40106 = n627 & ~n26342 ;
  assign n40107 = n20216 ^ n3738 ^ 1'b0 ;
  assign n40108 = n25387 ^ n20190 ^ 1'b0 ;
  assign n40109 = ~n40107 & n40108 ;
  assign n40110 = n1812 | n12163 ;
  assign n40111 = n10925 ^ n9952 ^ 1'b0 ;
  assign n40112 = ~n3509 & n40111 ;
  assign n40113 = n19323 ^ n13429 ^ 1'b0 ;
  assign n40114 = n3305 & n40113 ;
  assign n40115 = n11322 & ~n35523 ;
  assign n40116 = n6207 & n30102 ;
  assign n40117 = n4448 | n27414 ;
  assign n40118 = n7221 ^ n7185 ^ n6444 ;
  assign n40119 = n40117 | n40118 ;
  assign n40120 = n6376 & n31097 ;
  assign n40121 = n2403 & n40120 ;
  assign n40122 = n2955 | n30462 ;
  assign n40123 = n9442 | n40122 ;
  assign n40124 = n5187 & n10132 ;
  assign n40125 = n10481 | n10519 ;
  assign n40126 = n15266 ^ n14723 ^ n3318 ;
  assign n40127 = n4545 & ~n33455 ;
  assign n40128 = n2109 & ~n16020 ;
  assign n40129 = n5465 & n40128 ;
  assign n40130 = n6141 & n14824 ;
  assign n40131 = n24037 & ~n40130 ;
  assign n40132 = n4361 | n7051 ;
  assign n40133 = n941 ^ n878 ^ 1'b0 ;
  assign n40135 = n14520 & ~n29770 ;
  assign n40136 = n1619 & n40135 ;
  assign n40134 = n8957 & ~n19315 ;
  assign n40137 = n40136 ^ n40134 ^ 1'b0 ;
  assign n40138 = n31824 ^ n18158 ^ 1'b0 ;
  assign n40139 = n5756 | n35588 ;
  assign n40140 = n520 & n31639 ;
  assign n40141 = n40140 ^ n11740 ^ 1'b0 ;
  assign n40142 = ~n36649 & n40141 ;
  assign n40143 = ~n3466 & n38988 ;
  assign n40145 = n2080 & n5995 ;
  assign n40144 = n1233 | n2270 ;
  assign n40146 = n40145 ^ n40144 ^ 1'b0 ;
  assign n40147 = ( n212 & n1178 ) | ( n212 & n17749 ) | ( n1178 & n17749 ) ;
  assign n40148 = ~n5663 & n15302 ;
  assign n40149 = ~n3941 & n40148 ;
  assign n40150 = n2038 | n18646 ;
  assign n40151 = n17708 & ~n40150 ;
  assign n40152 = ~n40149 & n40151 ;
  assign n40153 = n6476 ^ n2687 ^ 1'b0 ;
  assign n40154 = n27489 & n40153 ;
  assign n40155 = ~n11875 & n40154 ;
  assign n40156 = n8092 & ~n29161 ;
  assign n40157 = n40156 ^ n1602 ^ 1'b0 ;
  assign n40158 = ~n7487 & n11798 ;
  assign n40159 = n27804 & n40158 ;
  assign n40160 = n40159 ^ n40078 ^ 1'b0 ;
  assign n40161 = n17834 & ~n18782 ;
  assign n40162 = n21275 & ~n37833 ;
  assign n40163 = n40162 ^ n7479 ^ 1'b0 ;
  assign n40164 = n32306 ^ n10026 ^ 1'b0 ;
  assign n40165 = n34180 ^ n10358 ^ 1'b0 ;
  assign n40166 = n11672 & ~n40165 ;
  assign n40167 = n22641 ^ n13108 ^ 1'b0 ;
  assign n40168 = n25378 | n35094 ;
  assign n40169 = n1455 | n40168 ;
  assign n40170 = n8597 | n40169 ;
  assign n40171 = ( n14476 & ~n14535 ) | ( n14476 & n25488 ) | ( ~n14535 & n25488 ) ;
  assign n40172 = n13742 ^ n781 ^ 1'b0 ;
  assign n40173 = n28015 & n40172 ;
  assign n40174 = n35367 & n40173 ;
  assign n40175 = n4578 & ~n23881 ;
  assign n40176 = n9591 ^ n3798 ^ 1'b0 ;
  assign n40177 = n1406 & ~n40176 ;
  assign n40178 = n29977 & n40177 ;
  assign n40179 = n40178 ^ n3939 ^ 1'b0 ;
  assign n40180 = n27026 ^ n561 ^ 1'b0 ;
  assign n40181 = n14523 & n40180 ;
  assign n40182 = n40181 ^ n24725 ^ 1'b0 ;
  assign n40183 = ~n4131 & n24661 ;
  assign n40187 = ~n1401 & n5868 ;
  assign n40188 = n40187 ^ n3706 ^ 1'b0 ;
  assign n40189 = n16619 & n40188 ;
  assign n40184 = n39104 ^ n3449 ^ 1'b0 ;
  assign n40185 = n40184 ^ n24513 ^ 1'b0 ;
  assign n40186 = n3532 & ~n40185 ;
  assign n40190 = n40189 ^ n40186 ^ 1'b0 ;
  assign n40191 = n40190 ^ n22590 ^ 1'b0 ;
  assign n40192 = n3312 ^ n666 ^ 1'b0 ;
  assign n40193 = ~n7596 & n11680 ;
  assign n40194 = n32493 | n40193 ;
  assign n40195 = n2361 & ~n3280 ;
  assign n40196 = n921 & n10433 ;
  assign n40197 = n40196 ^ n4545 ^ 1'b0 ;
  assign n40198 = n726 | n22061 ;
  assign n40199 = ( ~n19580 & n29797 ) | ( ~n19580 & n34128 ) | ( n29797 & n34128 ) ;
  assign n40200 = n40199 ^ n31684 ^ 1'b0 ;
  assign n40201 = n28371 ^ n5269 ^ 1'b0 ;
  assign n40202 = n175 | n31278 ;
  assign n40203 = n24611 | n40202 ;
  assign n40204 = n2162 | n14440 ;
  assign n40205 = n40204 ^ n3516 ^ 1'b0 ;
  assign n40206 = n883 | n40205 ;
  assign n40207 = n32133 ^ n2725 ^ n2076 ;
  assign n40208 = n40207 ^ n3589 ^ 1'b0 ;
  assign n40209 = ~n39469 & n40208 ;
  assign n40210 = n10389 & n40209 ;
  assign n40211 = n14443 | n40210 ;
  assign n40212 = n40211 ^ n10421 ^ 1'b0 ;
  assign n40213 = n16108 ^ n15913 ^ 1'b0 ;
  assign n40214 = ~n685 & n22663 ;
  assign n40215 = n32429 ^ n17569 ^ 1'b0 ;
  assign n40216 = n13784 & n18064 ;
  assign n40217 = n10780 & n40216 ;
  assign n40218 = n14054 & ~n21168 ;
  assign n40219 = n37743 ^ n12393 ^ 1'b0 ;
  assign n40220 = n8828 & n40219 ;
  assign n40221 = n2252 & ~n22417 ;
  assign n40222 = n23486 & n40221 ;
  assign n40223 = n5005 & n14226 ;
  assign n40224 = ~n38316 & n40223 ;
  assign n40225 = ~n24060 & n32616 ;
  assign n40226 = n17776 ^ n7358 ^ 1'b0 ;
  assign n40231 = n18302 & n18963 ;
  assign n40227 = ~n4367 & n8823 ;
  assign n40228 = n40227 ^ x3 ^ 1'b0 ;
  assign n40229 = n39782 | n40228 ;
  assign n40230 = n40229 ^ n26161 ^ 1'b0 ;
  assign n40232 = n40231 ^ n40230 ^ 1'b0 ;
  assign n40233 = n4760 & n12010 ;
  assign n40234 = n21126 & n40233 ;
  assign n40235 = n14259 ^ n7652 ^ 1'b0 ;
  assign n40236 = n85 | n1377 ;
  assign n40237 = n40235 & ~n40236 ;
  assign n40238 = ~n4840 & n14824 ;
  assign n40239 = n6349 & n40238 ;
  assign n40240 = n32451 ^ n13170 ^ n9079 ;
  assign n40241 = n13772 | n22059 ;
  assign n40242 = n40241 ^ n5929 ^ 1'b0 ;
  assign n40243 = n21059 & ~n40242 ;
  assign n40244 = n36956 ^ n22771 ^ n6453 ;
  assign n40245 = n3960 & ~n40244 ;
  assign n40246 = n2842 ^ n68 ^ 1'b0 ;
  assign n40247 = n35296 ^ n7060 ^ 1'b0 ;
  assign n40248 = n5551 | n34665 ;
  assign n40249 = n32424 ^ n2082 ^ 1'b0 ;
  assign n40250 = n378 & ~n40249 ;
  assign n40251 = n17999 ^ n2757 ^ 1'b0 ;
  assign n40252 = n40251 ^ n14792 ^ 1'b0 ;
  assign n40253 = n5642 & n12908 ;
  assign n40254 = ~n26707 & n40253 ;
  assign n40255 = n40254 ^ n31201 ^ 1'b0 ;
  assign n40256 = n40255 ^ n35717 ^ 1'b0 ;
  assign n40257 = n35721 ^ n6281 ^ 1'b0 ;
  assign n40258 = n9100 & n18956 ;
  assign n40260 = n29639 ^ n185 ^ 1'b0 ;
  assign n40261 = n2220 & n40260 ;
  assign n40259 = n4700 & n16130 ;
  assign n40262 = n40261 ^ n40259 ^ 1'b0 ;
  assign n40263 = n2335 | n8172 ;
  assign n40264 = n14381 & n40263 ;
  assign n40265 = n979 & n35444 ;
  assign n40266 = n38956 | n40265 ;
  assign n40267 = n34976 & ~n40266 ;
  assign n40268 = n9606 ^ n2040 ^ 1'b0 ;
  assign n40269 = n9461 & n40268 ;
  assign n40270 = ~n3095 & n13868 ;
  assign n40271 = n31418 ^ n24602 ^ 1'b0 ;
  assign n40272 = n40271 ^ n18316 ^ 1'b0 ;
  assign n40273 = ~n3237 & n4096 ;
  assign n40274 = n40273 ^ n16706 ^ 1'b0 ;
  assign n40275 = n4840 & n40274 ;
  assign n40276 = n14591 | n16704 ;
  assign n40277 = n40276 ^ n25333 ^ 1'b0 ;
  assign n40278 = n5245 ^ n4367 ^ 1'b0 ;
  assign n40279 = n40278 ^ n19875 ^ n7095 ;
  assign n40280 = ~n722 & n40279 ;
  assign n40281 = ~n5094 & n31998 ;
  assign n40282 = ~n24590 & n40281 ;
  assign n40283 = n22375 & ~n31962 ;
  assign n40284 = n757 | n4807 ;
  assign n40285 = n7860 ^ n2462 ^ 1'b0 ;
  assign n40286 = n7118 ^ n2419 ^ 1'b0 ;
  assign n40287 = n32713 ^ n5970 ^ 1'b0 ;
  assign n40288 = n4606 & ~n21849 ;
  assign n40289 = n184 & ~n35795 ;
  assign n40290 = n22329 ^ n10492 ^ 1'b0 ;
  assign n40291 = n38675 & n40290 ;
  assign n40292 = ~n148 & n3040 ;
  assign n40293 = n24569 & n40292 ;
  assign n40294 = n38113 ^ n8897 ^ 1'b0 ;
  assign n40295 = n30280 & n40294 ;
  assign n40296 = n2841 & ~n17913 ;
  assign n40297 = n40296 ^ n8347 ^ 1'b0 ;
  assign n40298 = ~n11574 & n40297 ;
  assign n40299 = n4137 | n27626 ;
  assign n40300 = n10828 & ~n40299 ;
  assign n40301 = n15188 ^ n8373 ^ 1'b0 ;
  assign n40302 = n4045 ^ n986 ^ 1'b0 ;
  assign n40303 = n40302 ^ n2068 ^ 1'b0 ;
  assign n40304 = ( n3968 & n18121 ) | ( n3968 & ~n24122 ) | ( n18121 & ~n24122 ) ;
  assign n40305 = n8656 & n40304 ;
  assign n40306 = ~n5789 & n40305 ;
  assign n40307 = ~n5973 & n15247 ;
  assign n40308 = n12371 & n40307 ;
  assign n40309 = n381 | n40308 ;
  assign n40310 = n40309 ^ n15255 ^ 1'b0 ;
  assign n40311 = n4193 & n21735 ;
  assign n40312 = n40311 ^ n2792 ^ 1'b0 ;
  assign n40313 = n19225 ^ n7670 ^ 1'b0 ;
  assign n40314 = n15438 ^ n12328 ^ 1'b0 ;
  assign n40315 = n2454 | n19333 ;
  assign n40316 = n7959 ^ n354 ^ 1'b0 ;
  assign n40317 = n15407 & n40316 ;
  assign n40318 = n40317 ^ n1070 ^ 1'b0 ;
  assign n40319 = n512 & n28044 ;
  assign n40320 = ~n488 & n2917 ;
  assign n40321 = ~n27257 & n40320 ;
  assign n40322 = n40321 ^ n8382 ^ 1'b0 ;
  assign n40323 = ~n22683 & n36469 ;
  assign n40324 = ~n14520 & n40323 ;
  assign n40325 = n23198 ^ n12877 ^ 1'b0 ;
  assign n40326 = n6296 & ~n12213 ;
  assign n40327 = ~n16225 & n40326 ;
  assign n40328 = n1235 & ~n40327 ;
  assign n40329 = n22438 & n40328 ;
  assign n40330 = n40329 ^ n4774 ^ 1'b0 ;
  assign n40331 = n25749 & ~n40330 ;
  assign n40332 = ~n12984 & n36743 ;
  assign n40333 = ~n6876 & n7143 ;
  assign n40334 = n40333 ^ n13559 ^ 1'b0 ;
  assign n40335 = n13000 ^ n2194 ^ 1'b0 ;
  assign n40336 = ~n28587 & n40335 ;
  assign n40337 = ~n8868 & n31109 ;
  assign n40338 = n36662 ^ n13691 ^ n10990 ;
  assign n40339 = ~n5801 & n18013 ;
  assign n40340 = n10431 | n28445 ;
  assign n40341 = n40339 | n40340 ;
  assign n40342 = n2476 & n25763 ;
  assign n40343 = n24246 ^ n13819 ^ 1'b0 ;
  assign n40344 = n25203 ^ n23457 ^ 1'b0 ;
  assign n40345 = n8562 & ~n10930 ;
  assign n40346 = n40345 ^ n7545 ^ 1'b0 ;
  assign n40347 = n30041 ^ n28979 ^ 1'b0 ;
  assign n40348 = ~n19128 & n40347 ;
  assign n40349 = n25576 ^ n21123 ^ 1'b0 ;
  assign n40350 = n12159 ^ n10035 ^ 1'b0 ;
  assign n40351 = n2342 & ~n40350 ;
  assign n40352 = n23493 ^ n768 ^ 1'b0 ;
  assign n40353 = n24304 ^ n6272 ^ 1'b0 ;
  assign n40354 = n159 | n40353 ;
  assign n40355 = n6711 ^ n5049 ^ 1'b0 ;
  assign n40356 = ~n13009 & n14874 ;
  assign n40357 = ~n30675 & n40356 ;
  assign n40358 = n7753 & n40357 ;
  assign n40359 = n5452 & ~n29597 ;
  assign n40360 = n404 | n40359 ;
  assign n40362 = n9213 ^ n6616 ^ 1'b0 ;
  assign n40363 = n7459 & n40362 ;
  assign n40361 = x0 & n38669 ;
  assign n40364 = n40363 ^ n40361 ^ 1'b0 ;
  assign n40368 = n13837 & ~n16047 ;
  assign n40365 = n675 | n3386 ;
  assign n40366 = ~n3030 & n40365 ;
  assign n40367 = n16346 | n40366 ;
  assign n40369 = n40368 ^ n40367 ^ 1'b0 ;
  assign n40370 = n8209 | n11177 ;
  assign n40371 = n40370 ^ n14586 ^ 1'b0 ;
  assign n40372 = n26130 & n40371 ;
  assign n40373 = ~n9036 & n14432 ;
  assign n40374 = ~n23862 & n40373 ;
  assign n40375 = ( ~n17073 & n34561 ) | ( ~n17073 & n40374 ) | ( n34561 & n40374 ) ;
  assign n40376 = ~n21820 & n32759 ;
  assign n40377 = n38265 ^ n4210 ^ 1'b0 ;
  assign n40378 = n17827 & ~n40377 ;
  assign n40379 = ~n5389 & n10044 ;
  assign n40380 = n40379 ^ n1404 ^ 1'b0 ;
  assign n40381 = ~n1637 & n37078 ;
  assign n40382 = n15443 ^ n351 ^ 1'b0 ;
  assign n40383 = n7091 | n31085 ;
  assign n40384 = n806 & ~n24349 ;
  assign n40385 = n40384 ^ n8353 ^ 1'b0 ;
  assign n40386 = n8472 & ~n20696 ;
  assign n40387 = ~n18181 & n40386 ;
  assign n40388 = n40387 ^ n23009 ^ 1'b0 ;
  assign n40389 = n26991 | n35311 ;
  assign n40390 = n40389 ^ n2105 ^ 1'b0 ;
  assign n40391 = n40390 ^ n8775 ^ 1'b0 ;
  assign n40392 = n34265 & ~n40391 ;
  assign n40394 = n13109 ^ n1669 ^ 1'b0 ;
  assign n40395 = n7693 & n40394 ;
  assign n40393 = ~n6256 & n8207 ;
  assign n40396 = n40395 ^ n40393 ^ n30532 ;
  assign n40398 = ( n4556 & n7920 ) | ( n4556 & ~n10398 ) | ( n7920 & ~n10398 ) ;
  assign n40399 = n9120 | n40398 ;
  assign n40397 = n297 & ~n6979 ;
  assign n40400 = n40399 ^ n40397 ^ 1'b0 ;
  assign n40401 = n40400 ^ n13121 ^ 1'b0 ;
  assign n40402 = n3589 & ~n4923 ;
  assign n40403 = ~n4906 & n40402 ;
  assign n40404 = n10191 & ~n40403 ;
  assign n40405 = n40404 ^ n32721 ^ 1'b0 ;
  assign n40406 = n5336 ^ n618 ^ 1'b0 ;
  assign n40407 = n36836 & ~n40406 ;
  assign n40408 = n26494 ^ n9507 ^ 1'b0 ;
  assign n40409 = n37819 | n40408 ;
  assign n40410 = n40407 & ~n40409 ;
  assign n40411 = n40410 ^ n25868 ^ 1'b0 ;
  assign n40412 = ~n11900 & n14083 ;
  assign n40413 = n29231 ^ n14926 ^ n12304 ;
  assign n40414 = n1992 | n9111 ;
  assign n40415 = n29951 ^ n3074 ^ 1'b0 ;
  assign n40416 = n40414 & n40415 ;
  assign n40418 = n9803 ^ n8857 ^ 1'b0 ;
  assign n40417 = n9655 & ~n12302 ;
  assign n40419 = n40418 ^ n40417 ^ 1'b0 ;
  assign n40420 = n9070 ^ n7223 ^ 1'b0 ;
  assign n40421 = n38980 ^ n30448 ^ 1'b0 ;
  assign n40422 = n19779 | n40421 ;
  assign n40423 = n2774 | n7786 ;
  assign n40424 = n40423 ^ n1512 ^ 1'b0 ;
  assign n40425 = ~n7079 & n30856 ;
  assign n40426 = n14918 ^ n13258 ^ 1'b0 ;
  assign n40427 = n29753 ^ n15770 ^ 1'b0 ;
  assign n40428 = n14908 | n40427 ;
  assign n40429 = n622 & n19420 ;
  assign n40430 = n29146 ^ n5583 ^ 1'b0 ;
  assign n40431 = n40429 & n40430 ;
  assign n40432 = n23948 ^ n2862 ^ 1'b0 ;
  assign n40433 = n1409 & n11460 ;
  assign n40434 = ~n1748 & n2636 ;
  assign n40435 = ~n23636 & n40434 ;
  assign n40436 = n10780 & n40435 ;
  assign n40438 = n4883 & ~n25538 ;
  assign n40437 = ~n32517 & n37282 ;
  assign n40439 = n40438 ^ n40437 ^ 1'b0 ;
  assign n40440 = n9823 ^ n6484 ^ 1'b0 ;
  assign n40441 = n7784 & n40440 ;
  assign n40442 = n25276 & n40441 ;
  assign n40443 = n18179 ^ n5747 ^ n2148 ;
  assign n40444 = n40443 ^ n29107 ^ 1'b0 ;
  assign n40446 = ~n5990 & n23678 ;
  assign n40445 = n10399 | n27627 ;
  assign n40447 = n40446 ^ n40445 ^ 1'b0 ;
  assign n40448 = n17024 ^ n10559 ^ 1'b0 ;
  assign n40449 = n8031 & ~n12316 ;
  assign n40450 = n39366 | n40449 ;
  assign n40451 = n12657 & n40450 ;
  assign n40452 = n40451 ^ n2813 ^ 1'b0 ;
  assign n40453 = n18588 | n37039 ;
  assign n40454 = n5302 | n33573 ;
  assign n40455 = n40453 & ~n40454 ;
  assign n40456 = n11501 ^ n2064 ^ 1'b0 ;
  assign n40457 = n36202 & n40456 ;
  assign n40458 = n35769 ^ n21532 ^ 1'b0 ;
  assign n40459 = n1310 & ~n29075 ;
  assign n40460 = n40458 & ~n40459 ;
  assign n40461 = n11209 ^ n6644 ^ 1'b0 ;
  assign n40462 = n4307 & n40461 ;
  assign n40463 = ~n37117 & n40462 ;
  assign n40464 = n8896 | n40463 ;
  assign n40465 = n2568 | n40464 ;
  assign n40466 = n11714 & ~n40465 ;
  assign n40467 = n40466 ^ n16344 ^ 1'b0 ;
  assign n40468 = n4931 & ~n28376 ;
  assign n40469 = ~n4062 & n10835 ;
  assign n40470 = ~n10517 & n40469 ;
  assign n40471 = ~n16013 & n40470 ;
  assign n40472 = n4749 & ~n12049 ;
  assign n40473 = ~n22374 & n40472 ;
  assign n40478 = n11502 ^ n1075 ^ 1'b0 ;
  assign n40476 = n7767 | n25159 ;
  assign n40477 = n40476 ^ n8405 ^ 1'b0 ;
  assign n40474 = n19445 | n25131 ;
  assign n40475 = n4616 & ~n40474 ;
  assign n40479 = n40478 ^ n40477 ^ n40475 ;
  assign n40480 = n11405 ^ n5227 ^ 1'b0 ;
  assign n40481 = n8689 | n40480 ;
  assign n40482 = n4780 | n40481 ;
  assign n40483 = n5677 & ~n40482 ;
  assign n40484 = n12234 ^ n6775 ^ n4328 ;
  assign n40485 = n33230 | n40484 ;
  assign n40486 = ~n6326 & n12540 ;
  assign n40487 = n23233 ^ n9747 ^ 1'b0 ;
  assign n40488 = n29973 ^ n15694 ^ 1'b0 ;
  assign n40489 = n24816 | n36858 ;
  assign n40495 = n626 & ~n6080 ;
  assign n40490 = n23652 ^ n865 ^ 1'b0 ;
  assign n40491 = n17910 & n27733 ;
  assign n40492 = n40491 ^ n39706 ^ 1'b0 ;
  assign n40493 = n40490 & ~n40492 ;
  assign n40494 = n40493 ^ n14984 ^ 1'b0 ;
  assign n40496 = n40495 ^ n40494 ^ n9337 ;
  assign n40497 = n38988 ^ n615 ^ 1'b0 ;
  assign n40498 = n466 & n29870 ;
  assign n40499 = n3692 | n14790 ;
  assign n40500 = n36770 ^ n1800 ^ 1'b0 ;
  assign n40501 = ~n40499 & n40500 ;
  assign n40502 = n8891 & n22643 ;
  assign n40503 = n31270 | n40502 ;
  assign n40504 = n40503 ^ n9032 ^ 1'b0 ;
  assign n40505 = n9233 | n12290 ;
  assign n40506 = n15398 ^ n1051 ^ 1'b0 ;
  assign n40507 = n4040 & ~n40506 ;
  assign n40508 = ~n4644 & n32988 ;
  assign n40509 = ~n10224 & n24156 ;
  assign n40510 = n159 & ~n4594 ;
  assign n40511 = n40509 & n40510 ;
  assign n40512 = ~n2295 & n32837 ;
  assign n40513 = n5684 | n15395 ;
  assign n40514 = n11707 & ~n40513 ;
  assign n40515 = n29664 ^ n27454 ^ 1'b0 ;
  assign n40516 = ~n31654 & n40515 ;
  assign n40517 = n3123 & ~n5551 ;
  assign n40518 = n40517 ^ n30791 ^ 1'b0 ;
  assign n40519 = n1008 | n4120 ;
  assign n40520 = n4620 & ~n40519 ;
  assign n40521 = n40269 & ~n40520 ;
  assign n40522 = ~n40518 & n40521 ;
  assign n40523 = n16184 | n22908 ;
  assign n40524 = n40523 ^ n12539 ^ 1'b0 ;
  assign n40525 = ( n6878 & ~n15132 ) | ( n6878 & n40524 ) | ( ~n15132 & n40524 ) ;
  assign n40526 = n9625 & n40525 ;
  assign n40527 = n29128 ^ n9903 ^ 1'b0 ;
  assign n40528 = n5894 & n10202 ;
  assign n40529 = ~n18494 & n40528 ;
  assign n40530 = ( n685 & n22649 ) | ( n685 & n40529 ) | ( n22649 & n40529 ) ;
  assign n40531 = n28077 & ~n40530 ;
  assign n40532 = n23506 & n40531 ;
  assign n40533 = n9490 | n11583 ;
  assign n40534 = n1790 & ~n40533 ;
  assign n40535 = n144 & ~n40534 ;
  assign n40536 = n40535 ^ n20683 ^ 1'b0 ;
  assign n40537 = x3 | n30875 ;
  assign n40538 = n4580 & ~n40537 ;
  assign n40539 = n1914 & n23065 ;
  assign n40540 = n40539 ^ n34470 ^ 1'b0 ;
  assign n40545 = ~n8121 & n26125 ;
  assign n40546 = ~n10676 & n40545 ;
  assign n40541 = n28438 ^ n6725 ^ 1'b0 ;
  assign n40542 = n17066 & ~n40541 ;
  assign n40543 = n40542 ^ n12697 ^ n8283 ;
  assign n40544 = ~n36447 & n40543 ;
  assign n40547 = n40546 ^ n40544 ^ 1'b0 ;
  assign n40548 = ( n2430 & n2929 ) | ( n2430 & n17550 ) | ( n2929 & n17550 ) ;
  assign n40549 = n7656 | n9705 ;
  assign n40550 = n40549 ^ n5731 ^ 1'b0 ;
  assign n40551 = n38245 & n40257 ;
  assign n40552 = n40550 & n40551 ;
  assign n40553 = ~n2680 & n37442 ;
  assign n40554 = n25153 ^ n21808 ^ 1'b0 ;
  assign n40555 = n23455 & ~n28871 ;
  assign n40556 = n40555 ^ n1739 ^ 1'b0 ;
  assign n40557 = n30708 ^ n29483 ^ 1'b0 ;
  assign n40558 = n5518 & ~n17467 ;
  assign n40559 = n24599 ^ n4552 ^ 1'b0 ;
  assign n40560 = ~n9488 & n31741 ;
  assign n40561 = ~n2761 & n5915 ;
  assign n40562 = n29072 & n40561 ;
  assign n40563 = n6332 & ~n37733 ;
  assign n40564 = ~n5706 & n40563 ;
  assign n40569 = n18223 ^ n6878 ^ n865 ;
  assign n40565 = n1887 & n7319 ;
  assign n40566 = n40565 ^ n2443 ^ 1'b0 ;
  assign n40567 = ~n1341 & n21495 ;
  assign n40568 = ( ~n17273 & n40566 ) | ( ~n17273 & n40567 ) | ( n40566 & n40567 ) ;
  assign n40570 = n40569 ^ n40568 ^ n22841 ;
  assign n40571 = n11057 & n14469 ;
  assign n40572 = n40571 ^ n3663 ^ 1'b0 ;
  assign n40573 = n9136 ^ n1653 ^ 1'b0 ;
  assign n40574 = n21076 & ~n40573 ;
  assign n40575 = ~n3681 & n11133 ;
  assign n40576 = n29579 ^ n23784 ^ 1'b0 ;
  assign n40577 = n32009 ^ n25307 ^ 1'b0 ;
  assign n40578 = n13094 ^ n10118 ^ 1'b0 ;
  assign n40579 = n12628 & n13537 ;
  assign n40580 = ~n26443 & n40579 ;
  assign n40581 = n40580 ^ n32018 ^ 1'b0 ;
  assign n40582 = ~n17763 & n23952 ;
  assign n40583 = ~n29872 & n40582 ;
  assign n40584 = n4968 | n15329 ;
  assign n40585 = n40584 ^ n79 ^ 1'b0 ;
  assign n40586 = n13354 | n31509 ;
  assign n40587 = ~n27364 & n36700 ;
  assign n40588 = n11590 & n39527 ;
  assign n40589 = n4504 & n34646 ;
  assign n40590 = ~n6250 & n40589 ;
  assign n40591 = n16687 ^ n2839 ^ 1'b0 ;
  assign n40592 = n22110 ^ n14786 ^ 1'b0 ;
  assign n40593 = n17717 & n32114 ;
  assign n40594 = n10280 | n40593 ;
  assign n40595 = n21066 ^ n9227 ^ 1'b0 ;
  assign n40596 = ~n26453 & n36238 ;
  assign n40597 = n21072 ^ n11585 ^ 1'b0 ;
  assign n40598 = n1525 & ~n8261 ;
  assign n40599 = ~n1660 & n40598 ;
  assign n40600 = n30487 ^ n19894 ^ 1'b0 ;
  assign n40601 = x1 & ~n40600 ;
  assign n40602 = n38252 ^ n17484 ^ 1'b0 ;
  assign n40603 = n2269 & ~n40602 ;
  assign n40604 = n39823 ^ n12899 ^ 1'b0 ;
  assign n40605 = n122 & ~n40604 ;
  assign n40606 = n27355 & ~n38891 ;
  assign n40607 = ~n11260 & n40606 ;
  assign n40608 = n3211 | n13877 ;
  assign n40609 = n18532 & ~n40608 ;
  assign n40610 = n6766 ^ n2849 ^ 1'b0 ;
  assign n40613 = ~n2979 & n28935 ;
  assign n40614 = ~n246 & n40613 ;
  assign n40615 = n21970 & n40614 ;
  assign n40611 = n1106 & n4991 ;
  assign n40612 = n14166 & n40611 ;
  assign n40616 = n40615 ^ n40612 ^ 1'b0 ;
  assign n40617 = n40616 ^ n17176 ^ 1'b0 ;
  assign n40618 = n34478 ^ n15574 ^ 1'b0 ;
  assign n40619 = ~n10925 & n15672 ;
  assign n40620 = n1520 & ~n40133 ;
  assign n40621 = n984 & n7345 ;
  assign n40622 = n40621 ^ n7920 ^ 1'b0 ;
  assign n40623 = ( n4742 & ~n37187 ) | ( n4742 & n40622 ) | ( ~n37187 & n40622 ) ;
  assign n40624 = n35442 ^ n1206 ^ 1'b0 ;
  assign n40625 = n28734 ^ n15655 ^ 1'b0 ;
  assign n40626 = n6187 | n20792 ;
  assign n40627 = ~n3779 & n29930 ;
  assign n40628 = n33484 ^ n9195 ^ n2734 ;
  assign n40629 = n2185 & n21325 ;
  assign n40630 = n156 | n25542 ;
  assign n40631 = n13470 | n40630 ;
  assign n40632 = n7612 | n15066 ;
  assign n40633 = n40632 ^ n25384 ^ n23987 ;
  assign n40634 = n6890 & n23512 ;
  assign n40635 = ~n5655 & n6084 ;
  assign n40636 = n40635 ^ n5043 ^ 1'b0 ;
  assign n40637 = n6071 | n17349 ;
  assign n40638 = n40637 ^ n1760 ^ 1'b0 ;
  assign n40639 = n5204 ^ n3158 ^ 1'b0 ;
  assign n40640 = n9197 & n10673 ;
  assign n40641 = n12649 ^ n8963 ^ 1'b0 ;
  assign n40642 = n23947 ^ n55 ^ 1'b0 ;
  assign n40643 = n294 & n10587 ;
  assign n40644 = n40643 ^ n2959 ^ 1'b0 ;
  assign n40645 = n37234 | n40644 ;
  assign n40646 = n1707 | n16947 ;
  assign n40647 = n20599 | n40646 ;
  assign n40648 = n2694 ^ n2585 ^ 1'b0 ;
  assign n40649 = n11907 & ~n16475 ;
  assign n40650 = n40649 ^ n2637 ^ 1'b0 ;
  assign n40651 = n5180 & ~n9193 ;
  assign n40652 = n28886 & n40651 ;
  assign n40653 = ~n7265 & n12274 ;
  assign n40654 = n12381 & n40653 ;
  assign n40655 = n2481 & n40654 ;
  assign n40656 = ~n1396 & n9425 ;
  assign n40657 = n40656 ^ n5284 ^ 1'b0 ;
  assign n40658 = n257 & ~n40657 ;
  assign n40659 = n1119 & n25953 ;
  assign n40660 = n37481 ^ n3116 ^ 1'b0 ;
  assign n40661 = n11833 & n29596 ;
  assign n40662 = n3008 | n38905 ;
  assign n40663 = n1141 ^ x4 ^ 1'b0 ;
  assign n40664 = n14245 ^ n1362 ^ 1'b0 ;
  assign n40665 = n19565 | n36900 ;
  assign n40666 = n40665 ^ n24336 ^ 1'b0 ;
  assign n40667 = n3146 & n40666 ;
  assign n40668 = n22397 ^ n11229 ^ 1'b0 ;
  assign n40669 = n9032 & ~n40668 ;
  assign n40670 = ~n352 & n40669 ;
  assign n40671 = n40670 ^ n7192 ^ 1'b0 ;
  assign n40672 = n18803 ^ n8874 ^ 1'b0 ;
  assign n40673 = n36362 ^ n30165 ^ 1'b0 ;
  assign n40674 = n40672 & n40673 ;
  assign n40675 = n5180 & n26313 ;
  assign n40676 = n2705 & ~n34307 ;
  assign n40677 = n2455 & n19944 ;
  assign n40678 = n10487 ^ n1027 ^ 1'b0 ;
  assign n40679 = n6200 | n19854 ;
  assign n40680 = n4320 ^ n3028 ^ 1'b0 ;
  assign n40681 = n9298 | n40680 ;
  assign n40682 = n17601 ^ n4882 ^ 1'b0 ;
  assign n40683 = n36859 ^ n3452 ^ 1'b0 ;
  assign n40684 = n1851 & ~n36152 ;
  assign n40685 = ~n47 & n40684 ;
  assign n40686 = n1860 | n10355 ;
  assign n40687 = n40686 ^ n22794 ^ 1'b0 ;
  assign n40688 = n40687 ^ n14046 ^ 1'b0 ;
  assign n40689 = n37087 ^ n14535 ^ 1'b0 ;
  assign n40690 = n1531 | n3452 ;
  assign n40691 = ~n556 & n828 ;
  assign n40692 = ~n40690 & n40691 ;
  assign n40693 = n5904 & n32436 ;
  assign n40694 = n8186 | n36270 ;
  assign n40695 = n40694 ^ n2314 ^ 1'b0 ;
  assign n40696 = n11037 & n25858 ;
  assign n40697 = n14245 ^ n2573 ^ n2431 ;
  assign n40698 = n38444 ^ n5562 ^ 1'b0 ;
  assign n40699 = ~n6434 & n19390 ;
  assign n40700 = n23099 ^ n14380 ^ 1'b0 ;
  assign n40703 = n5880 & n25250 ;
  assign n40701 = ~n8540 & n29132 ;
  assign n40702 = n32899 | n40701 ;
  assign n40704 = n40703 ^ n40702 ^ 1'b0 ;
  assign n40705 = n39754 ^ n20274 ^ 1'b0 ;
  assign n40706 = n16929 & ~n40705 ;
  assign n40707 = n40706 ^ n26385 ^ 1'b0 ;
  assign n40708 = n7376 | n7789 ;
  assign n40709 = n9009 | n14572 ;
  assign n40710 = n40708 | n40709 ;
  assign n40711 = ~n11448 & n11548 ;
  assign n40712 = n40711 ^ n867 ^ 1'b0 ;
  assign n40713 = ~n403 & n35907 ;
  assign n40714 = n3889 | n40713 ;
  assign n40715 = n20058 ^ n12175 ^ 1'b0 ;
  assign n40716 = ~n11245 & n18412 ;
  assign n40717 = n158 & ~n5270 ;
  assign n40718 = n128 & n40717 ;
  assign n40719 = n21363 & n40718 ;
  assign n40720 = ~n5121 & n40719 ;
  assign n40721 = ( n662 & ~n2913 ) | ( n662 & n8766 ) | ( ~n2913 & n8766 ) ;
  assign n40722 = n40721 ^ n38597 ^ 1'b0 ;
  assign n40723 = ~n7698 & n40722 ;
  assign n40724 = ~n23231 & n25796 ;
  assign n40725 = ~n1979 & n18833 ;
  assign n40726 = n26465 ^ n5094 ^ 1'b0 ;
  assign n40728 = n16438 & n17618 ;
  assign n40727 = ~n182 & n23990 ;
  assign n40729 = n40728 ^ n40727 ^ 1'b0 ;
  assign n40730 = n11618 | n25831 ;
  assign n40731 = n2238 & n2511 ;
  assign n40732 = n15626 & ~n40731 ;
  assign n40733 = ~n11464 & n40732 ;
  assign n40734 = n16819 ^ n12293 ^ 1'b0 ;
  assign n40735 = n33179 ^ n22140 ^ 1'b0 ;
  assign n40736 = n8169 ^ n353 ^ 1'b0 ;
  assign n40737 = ~n6603 & n40736 ;
  assign n40738 = n6107 & n40737 ;
  assign n40739 = n198 & n40738 ;
  assign n40740 = n15686 | n28363 ;
  assign n40741 = ~n590 & n1631 ;
  assign n40742 = ~n1874 & n30671 ;
  assign n40743 = n40742 ^ n15098 ^ 1'b0 ;
  assign n40744 = n34734 ^ n11740 ^ n4400 ;
  assign n40745 = n9524 ^ n8401 ^ 1'b0 ;
  assign n40746 = n8387 | n40745 ;
  assign n40747 = n24719 & ~n33700 ;
  assign n40748 = n40747 ^ n35627 ^ 1'b0 ;
  assign n40749 = n23538 ^ n10119 ^ n2082 ;
  assign n40750 = n12920 & n22976 ;
  assign n40751 = n6785 & n16212 ;
  assign n40752 = n5218 & n40751 ;
  assign n40753 = n40750 & n40752 ;
  assign n40754 = ( ~n1953 & n5635 ) | ( ~n1953 & n16367 ) | ( n5635 & n16367 ) ;
  assign n40755 = n5721 & n12238 ;
  assign n40756 = ~n12652 & n40755 ;
  assign n40757 = n40756 ^ n23948 ^ 1'b0 ;
  assign n40758 = n18186 ^ n4000 ^ 1'b0 ;
  assign n40759 = n27624 & n40758 ;
  assign n40760 = n17741 ^ n3408 ^ 1'b0 ;
  assign n40761 = n40760 ^ n9353 ^ 1'b0 ;
  assign n40762 = n37234 ^ n7269 ^ 1'b0 ;
  assign n40763 = n10878 | n40762 ;
  assign n40764 = n966 & n15090 ;
  assign n40765 = n40764 ^ n7936 ^ 1'b0 ;
  assign n40766 = n18224 | n20990 ;
  assign n40767 = n816 & ~n5319 ;
  assign n40768 = n7674 | n40767 ;
  assign n40769 = n10662 | n25512 ;
  assign n40770 = n40769 ^ n31774 ^ 1'b0 ;
  assign n40771 = ~n1491 & n4024 ;
  assign n40772 = n11373 ^ n5466 ^ 1'b0 ;
  assign n40773 = ~n10877 & n40772 ;
  assign n40774 = n40773 ^ n27362 ^ 1'b0 ;
  assign n40775 = n34781 & ~n40774 ;
  assign n40776 = n22055 & n40775 ;
  assign n40777 = ~n3025 & n10656 ;
  assign n40778 = ~n3116 & n40777 ;
  assign n40779 = n101 & ~n40778 ;
  assign n40780 = n40779 ^ n8548 ^ 1'b0 ;
  assign n40781 = n40780 ^ n14767 ^ 1'b0 ;
  assign n40782 = n32867 & ~n40781 ;
  assign n40783 = ~n20099 & n22239 ;
  assign n40784 = ~n982 & n32048 ;
  assign n40785 = n40784 ^ n962 ^ 1'b0 ;
  assign n40786 = n1165 | n32030 ;
  assign n40787 = ~n3408 & n14986 ;
  assign n40788 = n40787 ^ n2880 ^ 1'b0 ;
  assign n40789 = ~n7040 & n32367 ;
  assign n40790 = n19830 & n27740 ;
  assign n40791 = n40790 ^ n40569 ^ 1'b0 ;
  assign n40792 = ~n7110 & n26680 ;
  assign n40793 = n18041 | n19363 ;
  assign n40794 = n36689 ^ n19550 ^ 1'b0 ;
  assign n40795 = ~n371 & n40794 ;
  assign n40796 = ~n21232 & n27778 ;
  assign n40797 = n21639 | n27578 ;
  assign n40798 = n9959 & n40797 ;
  assign n40799 = n40798 ^ n27891 ^ 1'b0 ;
  assign n40800 = n26146 ^ n8840 ^ 1'b0 ;
  assign n40801 = n3524 | n23074 ;
  assign n40802 = n40801 ^ n14946 ^ 1'b0 ;
  assign n40803 = n13885 ^ n8637 ^ 1'b0 ;
  assign n40804 = n10477 & ~n40803 ;
  assign n40805 = ~n872 & n40804 ;
  assign n40806 = n15713 ^ n2004 ^ 1'b0 ;
  assign n40807 = ~n1379 & n24497 ;
  assign n40808 = ~n40806 & n40807 ;
  assign n40809 = n8185 ^ n1976 ^ 1'b0 ;
  assign n40810 = n1403 & n40809 ;
  assign n40811 = n7596 & n23691 ;
  assign n40812 = ~n8251 & n40811 ;
  assign n40813 = n26259 ^ n22291 ^ 1'b0 ;
  assign n40814 = ~n40812 & n40813 ;
  assign n40817 = n7679 ^ n2773 ^ 1'b0 ;
  assign n40815 = n27686 ^ n15810 ^ 1'b0 ;
  assign n40816 = n33735 | n40815 ;
  assign n40818 = n40817 ^ n40816 ^ 1'b0 ;
  assign n40819 = n2992 ^ n1893 ^ 1'b0 ;
  assign n40820 = n36123 ^ n25558 ^ 1'b0 ;
  assign n40821 = ~n108 & n302 ;
  assign n40822 = n40821 ^ n31794 ^ 1'b0 ;
  assign n40823 = n22699 ^ n5985 ^ 1'b0 ;
  assign n40824 = n6363 ^ n129 ^ 1'b0 ;
  assign n40825 = n8306 ^ n1914 ^ 1'b0 ;
  assign n40826 = n11436 ^ n929 ^ 1'b0 ;
  assign n40827 = n8461 & n22457 ;
  assign n40828 = n24689 ^ n3091 ^ 1'b0 ;
  assign n40829 = n5400 & n40828 ;
  assign n40830 = n40827 & n40829 ;
  assign n40831 = n40748 ^ n2910 ^ 1'b0 ;
  assign n40832 = n8321 & ~n39089 ;
  assign n40833 = ~n2342 & n15764 ;
  assign n40834 = n40833 ^ n1840 ^ 1'b0 ;
  assign n40835 = ~n17126 & n37643 ;
  assign n40836 = n40835 ^ n27820 ^ 1'b0 ;
  assign n40837 = n236 | n40836 ;
  assign n40838 = n7797 & ~n15098 ;
  assign n40839 = n9682 ^ n7927 ^ 1'b0 ;
  assign n40840 = ~n11787 & n40839 ;
  assign n40841 = ~n10156 & n40840 ;
  assign n40842 = n40841 ^ n727 ^ 1'b0 ;
  assign n40843 = n14701 ^ n5554 ^ 1'b0 ;
  assign n40844 = n40843 ^ n22134 ^ n10145 ;
  assign n40845 = n3853 & n9691 ;
  assign n40846 = n14128 & n28224 ;
  assign n40847 = n40846 ^ n2334 ^ 1'b0 ;
  assign n40848 = n520 ^ n55 ^ 1'b0 ;
  assign n40849 = n38630 & n40848 ;
  assign n40850 = ~n10349 & n40849 ;
  assign n40851 = x2 | n6691 ;
  assign n40852 = n40851 ^ n6998 ^ 1'b0 ;
  assign n40853 = n18818 | n24182 ;
  assign n40854 = n40853 ^ n28324 ^ 1'b0 ;
  assign n40855 = n40852 | n40854 ;
  assign n40856 = n9667 & n18062 ;
  assign n40857 = n4320 ^ n745 ^ 1'b0 ;
  assign n40858 = n3278 & n6365 ;
  assign n40859 = n12898 ^ n823 ^ 1'b0 ;
  assign n40860 = n15481 & n40859 ;
  assign n40861 = n8842 & ~n13164 ;
  assign n40862 = n12871 & n40861 ;
  assign n40863 = n26656 ^ n588 ^ 1'b0 ;
  assign n40864 = n2160 & n40863 ;
  assign n40865 = n3919 & n40864 ;
  assign n40866 = n14789 ^ n13612 ^ 1'b0 ;
  assign n40867 = n5034 | n40866 ;
  assign n40868 = n4231 | n40867 ;
  assign n40869 = ~n10056 & n14109 ;
  assign n40870 = n19330 | n22193 ;
  assign n40871 = n19964 | n23283 ;
  assign n40872 = n16040 ^ n1701 ^ 1'b0 ;
  assign n40873 = ~n215 & n40872 ;
  assign n40874 = n40871 & n40873 ;
  assign n40875 = n3542 & n17914 ;
  assign n40876 = n40875 ^ n22132 ^ 1'b0 ;
  assign n40877 = n1038 | n3141 ;
  assign n40878 = n23450 | n40877 ;
  assign n40879 = n31810 | n40878 ;
  assign n40880 = n18156 ^ n814 ^ 1'b0 ;
  assign n40881 = n387 | n40880 ;
  assign n40882 = n22422 ^ n18963 ^ 1'b0 ;
  assign n40883 = n27124 ^ n9483 ^ 1'b0 ;
  assign n40884 = ~n4545 & n40883 ;
  assign n40885 = n22215 ^ n3732 ^ 1'b0 ;
  assign n40886 = n11479 | n40885 ;
  assign n40887 = n412 & ~n584 ;
  assign n40888 = ~n2991 & n17994 ;
  assign n40889 = n14571 & ~n40888 ;
  assign n40890 = n13128 ^ n12995 ^ n1212 ;
  assign n40891 = n17635 ^ n16803 ^ 1'b0 ;
  assign n40892 = ~n40890 & n40891 ;
  assign n40893 = ~n14259 & n19099 ;
  assign n40894 = n34743 & n40893 ;
  assign n40895 = n2757 & n27778 ;
  assign n40896 = n27572 ^ n3477 ^ 1'b0 ;
  assign n40897 = n9796 ^ n2458 ^ 1'b0 ;
  assign n40898 = n2233 & ~n14544 ;
  assign n40899 = n40898 ^ n7888 ^ 1'b0 ;
  assign n40900 = n40899 ^ n1950 ^ 1'b0 ;
  assign n40901 = n12293 & n38241 ;
  assign n40902 = n16667 & ~n34288 ;
  assign n40903 = ~n3442 & n20847 ;
  assign n40904 = n30555 | n36035 ;
  assign n40905 = n14246 & ~n25704 ;
  assign n40906 = ~n12659 & n40905 ;
  assign n40907 = n27190 ^ n10459 ^ 1'b0 ;
  assign n40908 = n6141 ^ n3490 ^ 1'b0 ;
  assign n40909 = ~n33323 & n40908 ;
  assign n40911 = n7003 ^ n5180 ^ 1'b0 ;
  assign n40910 = n1947 | n9162 ;
  assign n40912 = n40911 ^ n40910 ^ 1'b0 ;
  assign n40913 = n19430 & n34408 ;
  assign n40914 = ~n6619 & n11158 ;
  assign n40915 = ~n28320 & n40914 ;
  assign n40916 = ~n33333 & n40915 ;
  assign n40919 = n10808 ^ n5068 ^ 1'b0 ;
  assign n40917 = n5727 ^ n646 ^ 1'b0 ;
  assign n40918 = ~n86 & n40917 ;
  assign n40920 = n40919 ^ n40918 ^ 1'b0 ;
  assign n40921 = n8158 ^ n7439 ^ 1'b0 ;
  assign n40922 = n15570 & n40921 ;
  assign n40923 = n2289 & n8295 ;
  assign n40924 = n5702 & n40923 ;
  assign n40925 = n40924 ^ n16687 ^ 1'b0 ;
  assign n40926 = n3032 | n40925 ;
  assign n40928 = n4365 ^ n191 ^ 1'b0 ;
  assign n40927 = ~n9377 & n14606 ;
  assign n40929 = n40928 ^ n40927 ^ 1'b0 ;
  assign n40930 = n20610 & n40929 ;
  assign n40931 = n11514 | n19776 ;
  assign n40932 = n40931 ^ n8330 ^ 1'b0 ;
  assign n40933 = n36220 ^ n24902 ^ n18342 ;
  assign n40934 = n836 & ~n1096 ;
  assign n40935 = ~n836 & n40934 ;
  assign n40936 = n2268 | n4578 ;
  assign n40937 = n40935 & ~n40936 ;
  assign n40938 = ~n1794 & n40937 ;
  assign n40939 = n5089 & n8589 ;
  assign n40940 = n40938 & n40939 ;
  assign n40941 = n4746 & ~n40940 ;
  assign n40942 = n40941 ^ n13229 ^ 1'b0 ;
  assign n40943 = n283 ^ n129 ^ 1'b0 ;
  assign n40944 = n40942 & n40943 ;
  assign n40945 = n40944 ^ n19227 ^ 1'b0 ;
  assign n40946 = n21449 ^ n97 ^ 1'b0 ;
  assign n40947 = n20044 & n40946 ;
  assign n40948 = n40947 ^ n24382 ^ 1'b0 ;
  assign n40949 = n40945 & ~n40948 ;
  assign n40950 = n29771 ^ n11323 ^ 1'b0 ;
  assign n40951 = n528 & n5688 ;
  assign n40952 = n40951 ^ n27423 ^ 1'b0 ;
  assign n40953 = n708 & n17530 ;
  assign n40954 = ~n22373 & n22623 ;
  assign n40955 = n40953 & n40954 ;
  assign n40956 = n22624 & n25212 ;
  assign n40957 = n40956 ^ n13841 ^ 1'b0 ;
  assign n40958 = ~n7676 & n12641 ;
  assign n40960 = n13174 ^ n713 ^ 1'b0 ;
  assign n40959 = n6289 & ~n13108 ;
  assign n40961 = n40960 ^ n40959 ^ 1'b0 ;
  assign n40962 = n22614 ^ n14194 ^ 1'b0 ;
  assign n40963 = n8181 & n40962 ;
  assign n40964 = n4809 ^ n3188 ^ 1'b0 ;
  assign n40965 = n3203 | n6926 ;
  assign n40966 = n20555 & ~n40965 ;
  assign n40967 = n40966 ^ n14483 ^ 1'b0 ;
  assign n40968 = n743 & n23633 ;
  assign n40969 = n7181 | n40968 ;
  assign n40970 = n5543 & ~n40969 ;
  assign n40971 = n40970 ^ n29899 ^ n12723 ;
  assign n40972 = n153 & ~n25519 ;
  assign n40973 = n38209 & n40972 ;
  assign n40974 = n25382 ^ n8503 ^ 1'b0 ;
  assign n40975 = n29579 | n40974 ;
  assign n40976 = n3472 & ~n40929 ;
  assign n40977 = n40976 ^ n9592 ^ 1'b0 ;
  assign n40978 = n40977 ^ n246 ^ 1'b0 ;
  assign n40979 = n40978 ^ n24938 ^ 1'b0 ;
  assign n40980 = ~n30070 & n30565 ;
  assign n40981 = ~n9354 & n23304 ;
  assign n40982 = n36856 ^ n36641 ^ 1'b0 ;
  assign n40983 = n16255 & ~n40982 ;
  assign n40984 = n40983 ^ n19146 ^ 1'b0 ;
  assign n40985 = n40981 | n40984 ;
  assign n40986 = n2613 | n15631 ;
  assign n40987 = n1310 & n16483 ;
  assign n40988 = n40987 ^ n3693 ^ 1'b0 ;
  assign n40989 = n1652 | n4907 ;
  assign n40990 = n4907 & ~n40989 ;
  assign n40991 = n7851 & n40990 ;
  assign n40992 = n12801 & n40991 ;
  assign n40993 = ~n12801 & n40992 ;
  assign n40994 = n40988 | n40993 ;
  assign n40995 = n40994 ^ n18276 ^ 1'b0 ;
  assign n40996 = ~n2873 & n40995 ;
  assign n40997 = n17449 ^ n7707 ^ 1'b0 ;
  assign n40998 = n4549 & n40997 ;
  assign n40999 = n10740 & n22464 ;
  assign n41000 = n7061 ^ n433 ^ 1'b0 ;
  assign n41001 = n4991 & n41000 ;
  assign n41002 = n37282 ^ n18831 ^ 1'b0 ;
  assign n41003 = n24470 ^ n7193 ^ 1'b0 ;
  assign n41004 = n15576 ^ n8564 ^ 1'b0 ;
  assign n41005 = ~n41003 & n41004 ;
  assign n41006 = n7998 ^ n7599 ^ 1'b0 ;
  assign n41007 = ~n16027 & n41006 ;
  assign n41008 = ~n4923 & n13453 ;
  assign n41009 = ~n19627 & n21572 ;
  assign n41010 = n957 & n14051 ;
  assign n41011 = ~n39325 & n41010 ;
  assign n41012 = n246 | n14272 ;
  assign n41013 = n41012 ^ n1933 ^ 1'b0 ;
  assign n41014 = n41013 ^ n18735 ^ 1'b0 ;
  assign n41015 = ~n1555 & n3537 ;
  assign n41016 = n41015 ^ n25965 ^ 1'b0 ;
  assign n41017 = n14440 & n24483 ;
  assign n41018 = n41017 ^ n32133 ^ 1'b0 ;
  assign n41019 = n17356 & n41018 ;
  assign n41020 = ( n3084 & ~n5270 ) | ( n3084 & n11629 ) | ( ~n5270 & n11629 ) ;
  assign n41021 = ~n1693 & n2101 ;
  assign n41022 = n41020 & ~n41021 ;
  assign n41023 = ~n4917 & n41022 ;
  assign n41024 = n8877 & ~n41023 ;
  assign n41025 = ( n31377 & n31630 ) | ( n31377 & ~n34477 ) | ( n31630 & ~n34477 ) ;
  assign n41026 = n5860 & ~n12325 ;
  assign n41027 = n13827 & n18223 ;
  assign n41028 = n14935 & n41027 ;
  assign n41029 = n2714 ^ n899 ^ 1'b0 ;
  assign n41030 = ~n2751 & n41029 ;
  assign n41031 = ~n495 & n41030 ;
  assign n41032 = n25195 & n27555 ;
  assign n41033 = n3808 & n24403 ;
  assign n41034 = n3264 | n3928 ;
  assign n41035 = n41034 ^ n34659 ^ 1'b0 ;
  assign n41036 = n41033 & ~n41035 ;
  assign n41037 = n21837 ^ n817 ^ 1'b0 ;
  assign n41038 = n3012 | n41037 ;
  assign n41040 = n26177 | n26185 ;
  assign n41039 = n1587 & ~n27313 ;
  assign n41041 = n41040 ^ n41039 ^ 1'b0 ;
  assign n41043 = ~n1947 & n28364 ;
  assign n41042 = n29977 & ~n34952 ;
  assign n41044 = n41043 ^ n41042 ^ 1'b0 ;
  assign n41045 = n14233 ^ n13038 ^ 1'b0 ;
  assign n41048 = n5732 | n16501 ;
  assign n41049 = n41048 ^ n1192 ^ 1'b0 ;
  assign n41046 = n1597 | n14278 ;
  assign n41047 = n41046 ^ n10931 ^ 1'b0 ;
  assign n41050 = n41049 ^ n41047 ^ 1'b0 ;
  assign n41051 = n9800 | n12343 ;
  assign n41052 = n1622 & ~n41051 ;
  assign n41053 = n34885 | n41052 ;
  assign n41054 = n33958 ^ n24391 ^ 1'b0 ;
  assign n41055 = n21754 & ~n24898 ;
  assign n41056 = n25564 ^ n3219 ^ 1'b0 ;
  assign n41057 = n22998 ^ n5905 ^ 1'b0 ;
  assign n41058 = n2109 & n41057 ;
  assign n41059 = n104 & ~n1929 ;
  assign n41060 = n10038 & ~n41059 ;
  assign n41061 = n30152 ^ n25239 ^ 1'b0 ;
  assign n41062 = ( n177 & n6770 ) | ( n177 & ~n41061 ) | ( n6770 & ~n41061 ) ;
  assign n41063 = n1007 & n12939 ;
  assign n41064 = n41063 ^ n235 ^ 1'b0 ;
  assign n41065 = n41062 | n41064 ;
  assign n41066 = n35448 ^ n19565 ^ 1'b0 ;
  assign n41067 = n5232 & n28899 ;
  assign n41068 = n22634 ^ n159 ^ 1'b0 ;
  assign n41069 = n19025 | n41068 ;
  assign n41070 = n1025 | n9760 ;
  assign n41071 = ~n10366 & n41070 ;
  assign n41072 = ( n2185 & n2969 ) | ( n2185 & n4830 ) | ( n2969 & n4830 ) ;
  assign n41073 = n10180 | n22697 ;
  assign n41074 = n41073 ^ n4254 ^ 1'b0 ;
  assign n41075 = n39773 & ~n41074 ;
  assign n41081 = n530 & n4845 ;
  assign n41079 = n8033 & n9370 ;
  assign n41076 = n16120 & ~n34633 ;
  assign n41077 = n41076 ^ n1505 ^ 1'b0 ;
  assign n41078 = n1800 | n41077 ;
  assign n41080 = n41079 ^ n41078 ^ 1'b0 ;
  assign n41082 = n41081 ^ n41080 ^ 1'b0 ;
  assign n41083 = n198 | n7814 ;
  assign n41084 = n27384 & n41083 ;
  assign n41085 = n34235 ^ n3221 ^ 1'b0 ;
  assign n41086 = n17592 & ~n41085 ;
  assign n41087 = ~n18047 & n29808 ;
  assign n41088 = n9499 & ~n35004 ;
  assign n41089 = n16391 & n25138 ;
  assign n41091 = n938 & n9359 ;
  assign n41092 = n41091 ^ n10288 ^ 1'b0 ;
  assign n41090 = n14472 & n24361 ;
  assign n41093 = n41092 ^ n41090 ^ 1'b0 ;
  assign n41094 = n7634 ^ n5084 ^ 1'b0 ;
  assign n41095 = n30240 & n41094 ;
  assign n41096 = n13174 | n27362 ;
  assign n41097 = n40888 & ~n41096 ;
  assign n41098 = n27885 ^ n8185 ^ 1'b0 ;
  assign n41099 = n36691 & ~n41098 ;
  assign n41100 = n33697 ^ n290 ^ 1'b0 ;
  assign n41101 = n3706 & ~n28757 ;
  assign n41102 = n41101 ^ n3235 ^ 1'b0 ;
  assign n41103 = n18995 ^ n2889 ^ 1'b0 ;
  assign n41104 = n27743 ^ n16031 ^ 1'b0 ;
  assign n41105 = n41103 | n41104 ;
  assign n41106 = n41105 ^ n36121 ^ 1'b0 ;
  assign n41107 = n3499 & ~n23553 ;
  assign n41108 = n41107 ^ n6819 ^ 1'b0 ;
  assign n41109 = n470 & ~n41108 ;
  assign n41110 = n22790 & n41109 ;
  assign n41111 = n665 & n13054 ;
  assign n41112 = ~n5981 & n8458 ;
  assign n41113 = ~n4779 & n41112 ;
  assign n41114 = n41113 ^ n29508 ^ n20014 ;
  assign n41115 = ~n25208 & n40516 ;
  assign n41116 = ( n7056 & ~n41114 ) | ( n7056 & n41115 ) | ( ~n41114 & n41115 ) ;
  assign n41117 = n4320 | n23718 ;
  assign n41118 = n11328 ^ n290 ^ 1'b0 ;
  assign n41119 = n5461 & ~n41118 ;
  assign n41120 = ~n190 & n10083 ;
  assign n41121 = n41030 ^ n41020 ^ 1'b0 ;
  assign n41123 = n24106 ^ n1184 ^ 1'b0 ;
  assign n41122 = n5746 | n31049 ;
  assign n41124 = n41123 ^ n41122 ^ 1'b0 ;
  assign n41125 = n818 & n16981 ;
  assign n41126 = n2761 & ~n41125 ;
  assign n41127 = n12935 & n30770 ;
  assign n41128 = ~n14808 & n41127 ;
  assign n41129 = n19055 & n26670 ;
  assign n41131 = n26966 & ~n35418 ;
  assign n41132 = n7188 & n41131 ;
  assign n41133 = n337 & n41132 ;
  assign n41130 = n11895 & n30004 ;
  assign n41134 = n41133 ^ n41130 ^ 1'b0 ;
  assign n41135 = n12293 & ~n17961 ;
  assign n41136 = n41135 ^ n3522 ^ 1'b0 ;
  assign n41137 = ~n10426 & n41136 ;
  assign n41138 = n31709 & n41137 ;
  assign n41139 = n37060 & n41138 ;
  assign n41140 = ~n9344 & n29447 ;
  assign n41141 = n11084 | n15925 ;
  assign n41142 = n622 & n20507 ;
  assign n41143 = n5574 ^ n1564 ^ 1'b0 ;
  assign n41144 = ~n41142 & n41143 ;
  assign n41145 = n770 & n4257 ;
  assign n41146 = ( n310 & n517 ) | ( n310 & n41145 ) | ( n517 & n41145 ) ;
  assign n41147 = ~n4981 & n6620 ;
  assign n41148 = n41147 ^ n4840 ^ 1'b0 ;
  assign n41149 = n41148 ^ n3452 ^ 1'b0 ;
  assign n41150 = n41146 | n41149 ;
  assign n41151 = n16923 | n41150 ;
  assign n41152 = n15902 ^ n984 ^ 1'b0 ;
  assign n41153 = n41152 ^ n16512 ^ 1'b0 ;
  assign n41154 = n41151 | n41153 ;
  assign n41155 = n472 | n6242 ;
  assign n41156 = n3742 ^ n2751 ^ 1'b0 ;
  assign n41157 = n4062 | n41156 ;
  assign n41158 = n41157 ^ n21167 ^ 1'b0 ;
  assign n41159 = ~n1771 & n24962 ;
  assign n41160 = n41159 ^ n28137 ^ 1'b0 ;
  assign n41161 = n16972 ^ n3589 ^ 1'b0 ;
  assign n41162 = n11434 ^ n5264 ^ 1'b0 ;
  assign n41163 = n5542 | n41162 ;
  assign n41164 = n25965 & ~n31280 ;
  assign n41165 = n33207 & n41164 ;
  assign n41166 = ~n1197 & n33720 ;
  assign n41167 = n41166 ^ n26495 ^ 1'b0 ;
  assign n41168 = n31818 ^ n5731 ^ 1'b0 ;
  assign n41169 = n11714 ^ n1235 ^ 1'b0 ;
  assign n41170 = n1683 | n28881 ;
  assign n41171 = n36654 ^ n21303 ^ 1'b0 ;
  assign n41172 = ~n20434 & n34624 ;
  assign n41173 = ~n40751 & n41172 ;
  assign n41174 = n28088 ^ n4193 ^ 1'b0 ;
  assign n41175 = ( n434 & ~n18609 ) | ( n434 & n19964 ) | ( ~n18609 & n19964 ) ;
  assign n41176 = n1891 | n41175 ;
  assign n41177 = n1268 & n2816 ;
  assign n41178 = n41177 ^ n12119 ^ 1'b0 ;
  assign n41179 = ~n12669 & n39624 ;
  assign n41180 = n14983 & ~n17546 ;
  assign n41181 = n41180 ^ n22762 ^ 1'b0 ;
  assign n41187 = n3300 | n12557 ;
  assign n41188 = n41187 ^ n16926 ^ 1'b0 ;
  assign n41182 = n5775 | n6463 ;
  assign n41183 = ~n1325 & n41182 ;
  assign n41184 = n21395 & n41183 ;
  assign n41185 = n41184 ^ n25861 ^ 1'b0 ;
  assign n41186 = ~n9070 & n41185 ;
  assign n41189 = n41188 ^ n41186 ^ 1'b0 ;
  assign n41190 = n178 & n3028 ;
  assign n41191 = n41190 ^ n1585 ^ 1'b0 ;
  assign n41192 = n23322 ^ n9384 ^ n2615 ;
  assign n41193 = n3040 | n41192 ;
  assign n41194 = n41193 ^ n3637 ^ 1'b0 ;
  assign n41195 = n16116 ^ n830 ^ 1'b0 ;
  assign n41196 = n5942 & ~n41195 ;
  assign n41197 = n36669 ^ n15745 ^ 1'b0 ;
  assign n41198 = n14383 ^ n1100 ^ 1'b0 ;
  assign n41199 = n748 | n41198 ;
  assign n41200 = n26287 ^ n24182 ^ n12028 ;
  assign n41201 = n15792 & n41200 ;
  assign n41202 = n23181 | n41201 ;
  assign n41203 = n41202 ^ n1057 ^ 1'b0 ;
  assign n41205 = n26221 ^ n6189 ^ 1'b0 ;
  assign n41204 = ~n11578 & n22052 ;
  assign n41206 = n41205 ^ n41204 ^ 1'b0 ;
  assign n41207 = ~n7819 & n37832 ;
  assign n41208 = n10638 & n41207 ;
  assign n41209 = ~n3007 & n13438 ;
  assign n41210 = n41208 & n41209 ;
  assign n41211 = n9213 ^ n6809 ^ n4899 ;
  assign n41212 = n41211 ^ n15668 ^ n2497 ;
  assign n41213 = n8090 | n33131 ;
  assign n41214 = n25439 ^ n1629 ^ 1'b0 ;
  assign n41215 = ~n16821 & n41214 ;
  assign n41216 = n41215 ^ n22363 ^ n20738 ;
  assign n41217 = n3321 & ~n41216 ;
  assign n41218 = ~n10194 & n41217 ;
  assign n41219 = n13381 ^ n12445 ^ 1'b0 ;
  assign n41220 = n7416 & ~n21804 ;
  assign n41221 = ~n12418 & n41220 ;
  assign n41222 = n4279 ^ n1286 ^ 1'b0 ;
  assign n41223 = n8209 & ~n22097 ;
  assign n41224 = n2249 & ~n15896 ;
  assign n41225 = n10113 ^ n7126 ^ 1'b0 ;
  assign n41226 = ~n17044 & n41225 ;
  assign n41227 = n39375 ^ n28285 ^ 1'b0 ;
  assign n41228 = n7626 & ~n18449 ;
  assign n41229 = n3149 & n23997 ;
  assign n41230 = n41229 ^ n6529 ^ 1'b0 ;
  assign n41231 = ~n41228 & n41230 ;
  assign n41232 = n41231 ^ n412 ^ 1'b0 ;
  assign n41234 = n1418 | n25871 ;
  assign n41235 = n8046 & ~n41234 ;
  assign n41233 = n55 & n27755 ;
  assign n41236 = n41235 ^ n41233 ^ 1'b0 ;
  assign n41237 = n41236 ^ n9292 ^ 1'b0 ;
  assign n41238 = n16535 | n41237 ;
  assign n41239 = ~n9524 & n19138 ;
  assign n41240 = n41239 ^ n19165 ^ 1'b0 ;
  assign n41241 = n12000 & ~n18636 ;
  assign n41242 = n23150 & ~n26439 ;
  assign n41243 = n17948 & n35381 ;
  assign n41244 = ~n34258 & n41243 ;
  assign n41245 = n33911 ^ n6944 ^ 1'b0 ;
  assign n41246 = ~n1958 & n13073 ;
  assign n41247 = n8885 & ~n10685 ;
  assign n41248 = n41247 ^ n10159 ^ 1'b0 ;
  assign n41249 = n41246 & ~n41248 ;
  assign n41250 = n2330 & ~n16072 ;
  assign n41251 = ~n3718 & n41250 ;
  assign n41252 = n41251 ^ n25976 ^ 1'b0 ;
  assign n41253 = n4640 | n5338 ;
  assign n41254 = n1314 & ~n12325 ;
  assign n41255 = n32963 ^ n16738 ^ 1'b0 ;
  assign n41256 = n7782 | n32997 ;
  assign n41257 = n19136 ^ n766 ^ 1'b0 ;
  assign n41258 = n16288 & n41257 ;
  assign n41259 = ~n23108 & n34018 ;
  assign n41260 = ~n41258 & n41259 ;
  assign n41261 = n21720 & n31973 ;
  assign n41262 = ~n8889 & n16344 ;
  assign n41263 = n6543 & n21597 ;
  assign n41264 = n470 & n1491 ;
  assign n41265 = n6058 & n41264 ;
  assign n41266 = n3585 | n14704 ;
  assign n41267 = n6336 ^ n2610 ^ 1'b0 ;
  assign n41268 = n29226 & ~n41267 ;
  assign n41269 = n41143 ^ n25709 ^ 1'b0 ;
  assign n41270 = n41268 & n41269 ;
  assign n41271 = n532 | n41270 ;
  assign n41272 = n7646 | n10098 ;
  assign n41273 = n12337 | n41272 ;
  assign n41274 = n18187 & ~n38338 ;
  assign n41275 = n5199 | n12721 ;
  assign n41276 = n41275 ^ n3021 ^ 1'b0 ;
  assign n41277 = n37210 ^ n25333 ^ 1'b0 ;
  assign n41278 = n2095 ^ n628 ^ n137 ;
  assign n41279 = n809 & ~n41278 ;
  assign n41280 = n891 | n16251 ;
  assign n41281 = n7654 | n30677 ;
  assign n41282 = n41281 ^ n27001 ^ 1'b0 ;
  assign n41283 = n41282 ^ n40146 ^ 1'b0 ;
  assign n41284 = ~n41280 & n41283 ;
  assign n41285 = n19410 | n25997 ;
  assign n41286 = n41285 ^ n5162 ^ 1'b0 ;
  assign n41287 = n6530 & ~n19713 ;
  assign n41288 = ~n41286 & n41287 ;
  assign n41289 = n32734 ^ n31839 ^ 1'b0 ;
  assign n41290 = n1847 ^ n371 ^ 1'b0 ;
  assign n41291 = ( ~n21475 & n27674 ) | ( ~n21475 & n41290 ) | ( n27674 & n41290 ) ;
  assign n41292 = ( n2995 & n10477 ) | ( n2995 & ~n11915 ) | ( n10477 & ~n11915 ) ;
  assign n41293 = n10346 ^ n1287 ^ 1'b0 ;
  assign n41294 = n13204 ^ n11437 ^ 1'b0 ;
  assign n41295 = ~n23764 & n41294 ;
  assign n41296 = n4155 & ~n24389 ;
  assign n41297 = ~n11319 & n41296 ;
  assign n41298 = ~n179 & n3370 ;
  assign n41299 = n4724 | n41298 ;
  assign n41300 = n41299 ^ n17075 ^ 1'b0 ;
  assign n41301 = n3178 | n41300 ;
  assign n41304 = n16137 & n23231 ;
  assign n41302 = ~n6090 & n7792 ;
  assign n41303 = n24254 | n41302 ;
  assign n41305 = n41304 ^ n41303 ^ 1'b0 ;
  assign n41306 = n22355 ^ n14924 ^ 1'b0 ;
  assign n41307 = ~n6442 & n9362 ;
  assign n41308 = ~n914 & n41307 ;
  assign n41309 = n4969 & n13433 ;
  assign n41310 = ~n4774 & n11160 ;
  assign n41311 = n41310 ^ n8210 ^ 1'b0 ;
  assign n41312 = n23754 ^ n19371 ^ 1'b0 ;
  assign n41313 = n6830 | n41312 ;
  assign n41314 = n27523 | n41313 ;
  assign n41315 = n41314 ^ n26303 ^ 1'b0 ;
  assign n41317 = n1137 | n1961 ;
  assign n41318 = n1137 & ~n41317 ;
  assign n41319 = n6133 & ~n41318 ;
  assign n41316 = n2166 & ~n27292 ;
  assign n41320 = n41319 ^ n41316 ^ 1'b0 ;
  assign n41321 = n527 & n20130 ;
  assign n41322 = n27414 & n41321 ;
  assign n41323 = ( n748 & n6713 ) | ( n748 & n8843 ) | ( n6713 & n8843 ) ;
  assign n41324 = ~n22701 & n24490 ;
  assign n41325 = n23635 & ~n29713 ;
  assign n41326 = n41325 ^ n13717 ^ 1'b0 ;
  assign n41327 = n7824 ^ n7273 ^ 1'b0 ;
  assign n41328 = n13085 ^ n7681 ^ 1'b0 ;
  assign n41329 = ~n14612 & n21988 ;
  assign n41330 = n41329 ^ n13380 ^ 1'b0 ;
  assign n41331 = n41328 | n41330 ;
  assign n41332 = n3701 & ~n5823 ;
  assign n41333 = n41332 ^ n38920 ^ 1'b0 ;
  assign n41334 = n2983 | n12678 ;
  assign n41335 = ( n1073 & ~n3801 ) | ( n1073 & n41334 ) | ( ~n3801 & n41334 ) ;
  assign n41336 = n8755 | n16421 ;
  assign n41337 = n12073 | n29307 ;
  assign n41338 = n5284 & ~n41337 ;
  assign n41339 = n3656 & n35554 ;
  assign n41340 = n41339 ^ n659 ^ 1'b0 ;
  assign n41341 = ~n525 & n34041 ;
  assign n41342 = ~n2558 & n41341 ;
  assign n41343 = n41342 ^ n618 ^ 1'b0 ;
  assign n41344 = n41340 | n41343 ;
  assign n41345 = n2883 | n33519 ;
  assign n41346 = n31919 ^ n7455 ^ 1'b0 ;
  assign n41347 = n12199 | n41346 ;
  assign n41348 = n20395 ^ n10190 ^ 1'b0 ;
  assign n41349 = n41348 ^ n20649 ^ n17371 ;
  assign n41350 = n17796 ^ n2356 ^ 1'b0 ;
  assign n41351 = n41350 ^ n35042 ^ 1'b0 ;
  assign n41352 = n6270 & n8128 ;
  assign n41353 = n41352 ^ n745 ^ 1'b0 ;
  assign n41354 = ~n9954 & n39376 ;
  assign n41355 = n4779 & ~n10255 ;
  assign n41356 = n10784 & n41355 ;
  assign n41357 = n41356 ^ n24930 ^ 1'b0 ;
  assign n41358 = n41357 ^ n17934 ^ 1'b0 ;
  assign n41359 = n2611 & n5977 ;
  assign n41360 = n41359 ^ n23003 ^ n3370 ;
  assign n41361 = n7117 & ~n15958 ;
  assign n41362 = n41361 ^ n4394 ^ 1'b0 ;
  assign n41363 = n18387 & ~n41362 ;
  assign n41364 = n8071 | n12310 ;
  assign n41365 = n41363 & ~n41364 ;
  assign n41366 = n5826 | n41365 ;
  assign n41367 = n11827 | n36357 ;
  assign n41368 = n41367 ^ n24782 ^ 1'b0 ;
  assign n41369 = n532 | n32154 ;
  assign n41370 = n8625 & n15693 ;
  assign n41371 = n9086 & ~n29963 ;
  assign n41372 = n41370 & n41371 ;
  assign n41373 = n38771 ^ n15023 ^ n13588 ;
  assign n41374 = ~n14792 & n15322 ;
  assign n41375 = ~n737 & n9512 ;
  assign n41376 = ~n27774 & n41375 ;
  assign n41377 = n41374 & ~n41376 ;
  assign n41378 = n4000 | n8397 ;
  assign n41379 = n1550 & ~n1753 ;
  assign n41380 = n41379 ^ n2426 ^ 1'b0 ;
  assign n41381 = n41380 ^ n38847 ^ n24393 ;
  assign n41382 = n7338 | n17816 ;
  assign n41383 = n41247 & ~n41382 ;
  assign n41384 = n10966 ^ n2939 ^ 1'b0 ;
  assign n41385 = n8139 | n41384 ;
  assign n41386 = n857 | n8034 ;
  assign n41387 = n3363 & n13691 ;
  assign n41388 = ~n41386 & n41387 ;
  assign n41389 = n13577 & ~n35625 ;
  assign n41390 = n31695 & n41389 ;
  assign n41391 = n36427 ^ n18820 ^ 1'b0 ;
  assign n41392 = n6885 | n12887 ;
  assign n41393 = n28992 ^ n8567 ^ 1'b0 ;
  assign n41394 = n41392 | n41393 ;
  assign n41395 = n36529 ^ n15546 ^ 1'b0 ;
  assign n41396 = n5152 & ~n16124 ;
  assign n41397 = ~n41395 & n41396 ;
  assign n41398 = n7910 ^ n16 ^ 1'b0 ;
  assign n41399 = n35749 ^ n20501 ^ 1'b0 ;
  assign n41400 = n37 | n41399 ;
  assign n41401 = n14123 ^ n182 ^ 1'b0 ;
  assign n41402 = n41400 | n41401 ;
  assign n41403 = n13453 ^ n3717 ^ 1'b0 ;
  assign n41404 = n33733 & n41403 ;
  assign n41405 = ~n2822 & n41404 ;
  assign n41406 = n41405 ^ n5953 ^ 1'b0 ;
  assign n41407 = n41402 | n41406 ;
  assign n41408 = n32136 ^ n1277 ^ 1'b0 ;
  assign n41409 = ~n3764 & n4120 ;
  assign n41410 = n41409 ^ n37658 ^ 1'b0 ;
  assign n41412 = n10978 | n17764 ;
  assign n41413 = n41412 ^ n32624 ^ 1'b0 ;
  assign n41411 = n16176 | n20619 ;
  assign n41414 = n41413 ^ n41411 ^ 1'b0 ;
  assign n41415 = n5152 & n33423 ;
  assign n41416 = n41415 ^ n24609 ^ 1'b0 ;
  assign n41417 = n32578 ^ n23564 ^ 1'b0 ;
  assign n41418 = ~n1331 & n8667 ;
  assign n41419 = ~n6967 & n41418 ;
  assign n41420 = n41419 ^ n393 ^ 1'b0 ;
  assign n41421 = n33545 ^ n9997 ^ 1'b0 ;
  assign n41422 = ~n7290 & n9335 ;
  assign n41423 = n28343 & n41422 ;
  assign n41424 = n2251 | n11646 ;
  assign n41425 = n41423 & ~n41424 ;
  assign n41426 = n6907 | n41425 ;
  assign n41427 = n41426 ^ n883 ^ 1'b0 ;
  assign n41428 = n20225 & ~n38008 ;
  assign n41429 = n5981 & n41428 ;
  assign n41430 = n36245 ^ n31618 ^ 1'b0 ;
  assign n41431 = n29035 ^ n2923 ^ 1'b0 ;
  assign n41432 = n19102 | n41431 ;
  assign n41433 = n10930 | n29097 ;
  assign n41434 = n6847 & ~n11623 ;
  assign n41436 = n1533 | n4969 ;
  assign n41435 = n2727 | n32248 ;
  assign n41437 = n41436 ^ n41435 ^ 1'b0 ;
  assign n41438 = n25694 ^ n4159 ^ 1'b0 ;
  assign n41440 = n22770 ^ n1645 ^ 1'b0 ;
  assign n41439 = n9449 & ~n30951 ;
  assign n41441 = n41440 ^ n41439 ^ 1'b0 ;
  assign n41442 = n4182 | n5227 ;
  assign n41445 = n12799 ^ n6304 ^ n2843 ;
  assign n41446 = n1106 & n41445 ;
  assign n41447 = n41446 ^ n24006 ^ 1'b0 ;
  assign n41448 = n2807 ^ n1598 ^ 1'b0 ;
  assign n41449 = n41447 & n41448 ;
  assign n41443 = n4209 ^ n3095 ^ 1'b0 ;
  assign n41444 = n29169 & ~n41443 ;
  assign n41450 = n41449 ^ n41444 ^ 1'b0 ;
  assign n41451 = n363 | n6192 ;
  assign n41452 = ( n28556 & ~n32201 ) | ( n28556 & n41451 ) | ( ~n32201 & n41451 ) ;
  assign n41453 = ~n3743 & n26509 ;
  assign n41454 = n5872 & n16925 ;
  assign n41455 = n41454 ^ n5212 ^ 1'b0 ;
  assign n41456 = n2538 | n7360 ;
  assign n41457 = n41456 ^ n7495 ^ 1'b0 ;
  assign n41458 = n27708 & ~n41457 ;
  assign n41459 = ~n41455 & n41458 ;
  assign n41460 = n8953 | n11670 ;
  assign n41461 = ( n5747 & n39216 ) | ( n5747 & n41460 ) | ( n39216 & n41460 ) ;
  assign n41462 = n41461 ^ n15981 ^ 1'b0 ;
  assign n41463 = n7192 | n10725 ;
  assign n41464 = n11917 | n41463 ;
  assign n41465 = n41464 ^ n30269 ^ 1'b0 ;
  assign n41466 = ~n2686 & n29254 ;
  assign n41467 = n6441 & n12991 ;
  assign n41468 = ~n16473 & n41467 ;
  assign n41469 = n10762 & n26733 ;
  assign n41470 = n7707 | n35306 ;
  assign n41471 = n41469 | n41470 ;
  assign n41472 = n9461 ^ n2909 ^ 1'b0 ;
  assign n41473 = n13281 & ~n41472 ;
  assign n41474 = n13174 | n41473 ;
  assign n41475 = n41474 ^ n35657 ^ n98 ;
  assign n41476 = n1634 | n2661 ;
  assign n41477 = n10726 & ~n41476 ;
  assign n41478 = n27510 & ~n41477 ;
  assign n41479 = n19630 & n40251 ;
  assign n41480 = ~n627 & n41479 ;
  assign n41481 = n4525 | n11808 ;
  assign n41482 = n41481 ^ n21753 ^ 1'b0 ;
  assign n41483 = n10215 | n19566 ;
  assign n41484 = n12090 | n41483 ;
  assign n41485 = n26796 ^ n15777 ^ 1'b0 ;
  assign n41486 = n41484 & n41485 ;
  assign n41487 = n11803 & ~n14105 ;
  assign n41489 = n24839 ^ n7003 ^ 1'b0 ;
  assign n41488 = n21288 | n27198 ;
  assign n41490 = n41489 ^ n41488 ^ 1'b0 ;
  assign n41491 = n5518 ^ n1602 ^ 1'b0 ;
  assign n41492 = n6079 & ~n41491 ;
  assign n41493 = n30289 ^ n28684 ^ 1'b0 ;
  assign n41494 = n12169 ^ n6219 ^ 1'b0 ;
  assign n41495 = ~n5423 & n36015 ;
  assign n41496 = n5119 & ~n8056 ;
  assign n41497 = n5779 | n6464 ;
  assign n41498 = ~n30429 & n35140 ;
  assign n41499 = ~n41497 & n41498 ;
  assign n41505 = ~n1038 & n20437 ;
  assign n41506 = n37523 & n41505 ;
  assign n41503 = n18047 ^ n657 ^ 1'b0 ;
  assign n41504 = ~n28323 & n41503 ;
  assign n41507 = n41506 ^ n41504 ^ 1'b0 ;
  assign n41500 = n33844 ^ n25190 ^ 1'b0 ;
  assign n41501 = n6534 & n41500 ;
  assign n41502 = n17445 & n41501 ;
  assign n41508 = n41507 ^ n41502 ^ 1'b0 ;
  assign n41509 = n13044 ^ n10025 ^ 1'b0 ;
  assign n41510 = n1825 ^ n395 ^ 1'b0 ;
  assign n41511 = ~n21976 & n41510 ;
  assign n41512 = n41511 ^ n13092 ^ 1'b0 ;
  assign n41513 = ~n23978 & n29973 ;
  assign n41514 = n30922 ^ n1865 ^ 1'b0 ;
  assign n41515 = n2558 & n14094 ;
  assign n41516 = ~n1106 & n7247 ;
  assign n41517 = n38617 ^ n29175 ^ 1'b0 ;
  assign n41518 = n6619 & ~n14114 ;
  assign n41519 = n259 | n6284 ;
  assign n41520 = ~n7383 & n41519 ;
  assign n41521 = n18894 ^ n16840 ^ 1'b0 ;
  assign n41522 = n24089 ^ n21742 ^ 1'b0 ;
  assign n41523 = ~n4729 & n5763 ;
  assign n41524 = n23142 & n41523 ;
  assign n41525 = n17800 ^ n13042 ^ 1'b0 ;
  assign n41526 = ~n12750 & n26742 ;
  assign n41527 = n41526 ^ n2203 ^ 1'b0 ;
  assign n41528 = n33479 | n37819 ;
  assign n41529 = n41528 ^ n9800 ^ 1'b0 ;
  assign n41530 = n26600 & n34479 ;
  assign n41531 = n41530 ^ n9004 ^ 1'b0 ;
  assign n41532 = n12738 & n38053 ;
  assign n41533 = n30781 & ~n41532 ;
  assign n41534 = n41531 & n41533 ;
  assign n41535 = n16760 ^ n323 ^ 1'b0 ;
  assign n41536 = n117 & ~n1456 ;
  assign n41537 = n39374 ^ n3154 ^ 1'b0 ;
  assign n41538 = n7674 & ~n41537 ;
  assign n41539 = n11235 & n41538 ;
  assign n41540 = ~n8151 & n12446 ;
  assign n41541 = n18630 & ~n41540 ;
  assign n41542 = ( ~n7678 & n25091 ) | ( ~n7678 & n29592 ) | ( n25091 & n29592 ) ;
  assign n41543 = n36218 ^ n2731 ^ 1'b0 ;
  assign n41544 = n41542 & ~n41543 ;
  assign n41545 = ~n20517 & n22148 ;
  assign n41546 = n3922 & n5199 ;
  assign n41547 = n8539 ^ n1491 ^ 1'b0 ;
  assign n41548 = ~n3299 & n41547 ;
  assign n41549 = n15759 ^ n15111 ^ n9512 ;
  assign n41550 = n129 & n13608 ;
  assign n41551 = n4186 & ~n28497 ;
  assign n41552 = n1528 & ~n3416 ;
  assign n41553 = n3637 | n41552 ;
  assign n41554 = ( n3601 & n7403 ) | ( n3601 & n18205 ) | ( n7403 & n18205 ) ;
  assign n41555 = n9169 | n27964 ;
  assign n41556 = n32487 & ~n41555 ;
  assign n41557 = ~n11427 & n12529 ;
  assign n41558 = ~n4139 & n13469 ;
  assign n41559 = n2837 & ~n40853 ;
  assign n41560 = n23412 & n41559 ;
  assign n41561 = n7775 | n20730 ;
  assign n41562 = n1209 ^ n556 ^ 1'b0 ;
  assign n41563 = n38061 & ~n41562 ;
  assign n41564 = n12185 & ~n21091 ;
  assign n41565 = ~n38015 & n41564 ;
  assign n41566 = n36697 & n41565 ;
  assign n41567 = n25344 | n41477 ;
  assign n41572 = n12672 ^ n10166 ^ 1'b0 ;
  assign n41573 = n6161 & n41572 ;
  assign n41568 = n15512 ^ n5018 ^ 1'b0 ;
  assign n41569 = n23316 & ~n41568 ;
  assign n41570 = n41569 ^ n2699 ^ 1'b0 ;
  assign n41571 = n25315 & n41570 ;
  assign n41574 = n41573 ^ n41571 ^ 1'b0 ;
  assign n41575 = ~n30744 & n31964 ;
  assign n41576 = n41575 ^ n13844 ^ 1'b0 ;
  assign n41577 = n715 & ~n24859 ;
  assign n41578 = n29641 ^ n7749 ^ 1'b0 ;
  assign n41579 = n41577 & n41578 ;
  assign n41580 = ~n25220 & n41579 ;
  assign n41581 = n35774 & n35931 ;
  assign n41582 = n41581 ^ n31964 ^ 1'b0 ;
  assign n41583 = n33051 ^ n31484 ^ 1'b0 ;
  assign n41584 = n7894 ^ n7135 ^ 1'b0 ;
  assign n41585 = ~n10836 & n16714 ;
  assign n41586 = n1759 | n37056 ;
  assign n41587 = ~n10655 & n11798 ;
  assign n41588 = ~n20255 & n41587 ;
  assign n41589 = n6454 & n7803 ;
  assign n41590 = n41589 ^ n7853 ^ 1'b0 ;
  assign n41591 = ~n2148 & n16336 ;
  assign n41592 = n41591 ^ n6834 ^ 1'b0 ;
  assign n41593 = ~n25510 & n41592 ;
  assign n41594 = n31986 ^ n17191 ^ 1'b0 ;
  assign n41595 = n1207 & ~n24914 ;
  assign n41596 = n18997 & n41595 ;
  assign n41597 = n41596 ^ n23843 ^ 1'b0 ;
  assign n41598 = n2521 | n18028 ;
  assign n41599 = ~n4111 & n16322 ;
  assign n41600 = n2615 & n39319 ;
  assign n41601 = n41600 ^ n2150 ^ 1'b0 ;
  assign n41602 = n2303 | n5495 ;
  assign n41603 = n41602 ^ n10047 ^ 1'b0 ;
  assign n41604 = n128 & n17169 ;
  assign n41605 = n532 | n19350 ;
  assign n41606 = n412 | n41605 ;
  assign n41607 = ~n3089 & n8257 ;
  assign n41608 = n403 & n41607 ;
  assign n41609 = n24784 ^ n22214 ^ 1'b0 ;
  assign n41610 = n8817 & ~n41609 ;
  assign n41611 = ~n17895 & n41610 ;
  assign n41612 = n7383 & n8990 ;
  assign n41613 = n10268 | n10952 ;
  assign n41614 = n3093 & n35673 ;
  assign n41615 = ~n41613 & n41614 ;
  assign n41616 = n3314 ^ n177 ^ 1'b0 ;
  assign n41617 = n25514 | n41616 ;
  assign n41618 = n21299 & n40928 ;
  assign n41619 = n33929 ^ n1270 ^ 1'b0 ;
  assign n41620 = ~n8061 & n41619 ;
  assign n41621 = n310 | n17104 ;
  assign n41622 = n41621 ^ n32863 ^ 1'b0 ;
  assign n41623 = n1469 | n37003 ;
  assign n41624 = n31231 & n39094 ;
  assign n41625 = ~n191 & n11308 ;
  assign n41626 = n41625 ^ n17460 ^ 1'b0 ;
  assign n41627 = n3378 | n13838 ;
  assign n41628 = n25560 ^ n8081 ^ 1'b0 ;
  assign n41629 = n7319 & ~n41628 ;
  assign n41630 = n7197 | n39397 ;
  assign n41631 = n1065 & ~n41630 ;
  assign n41633 = n10439 & ~n10879 ;
  assign n41634 = n41633 ^ n11277 ^ 1'b0 ;
  assign n41632 = n6017 ^ n3606 ^ 1'b0 ;
  assign n41635 = n41634 ^ n41632 ^ n32995 ;
  assign n41636 = n19832 & ~n24419 ;
  assign n41637 = n14086 & n22097 ;
  assign n41638 = n39987 & n41637 ;
  assign n41639 = n41638 ^ n5854 ^ 1'b0 ;
  assign n41640 = n30500 ^ n18979 ^ 1'b0 ;
  assign n41641 = n34792 | n41640 ;
  assign n41642 = n10233 ^ n2714 ^ 1'b0 ;
  assign n41643 = n4937 & ~n41642 ;
  assign n41644 = ~n1878 & n41643 ;
  assign n41645 = n2767 | n8309 ;
  assign n41646 = n321 & n31209 ;
  assign n41647 = ~n8692 & n9312 ;
  assign n41648 = n11907 & n39617 ;
  assign n41649 = n20575 ^ n5067 ^ 1'b0 ;
  assign n41650 = n2476 & ~n41649 ;
  assign n41651 = n12361 & n41650 ;
  assign n41652 = n30471 ^ n484 ^ 1'b0 ;
  assign n41653 = n3900 & n41652 ;
  assign n41654 = n22401 | n27031 ;
  assign n41655 = ~n2288 & n7563 ;
  assign n41656 = ~n23580 & n41655 ;
  assign n41657 = n16356 | n41656 ;
  assign n41658 = n35256 ^ n30956 ^ 1'b0 ;
  assign n41659 = ~n7612 & n41658 ;
  assign n41660 = n37507 ^ n7265 ^ 1'b0 ;
  assign n41661 = n30100 ^ n20289 ^ 1'b0 ;
  assign n41662 = ( n6365 & ~n14441 ) | ( n6365 & n41661 ) | ( ~n14441 & n41661 ) ;
  assign n41663 = ~n18144 & n35542 ;
  assign n41664 = ~n6822 & n41663 ;
  assign n41665 = ~n7537 & n10425 ;
  assign n41666 = n15244 & n22348 ;
  assign n41667 = n3784 & n7924 ;
  assign n41668 = n41667 ^ n16645 ^ 1'b0 ;
  assign n41669 = n4228 & n41668 ;
  assign n41670 = n33895 ^ n7749 ^ 1'b0 ;
  assign n41671 = n41669 & n41670 ;
  assign n41672 = ~n4688 & n9085 ;
  assign n41673 = n41672 ^ n993 ^ 1'b0 ;
  assign n41674 = n4924 & n31574 ;
  assign n41675 = n41674 ^ n40231 ^ 1'b0 ;
  assign n41676 = n1523 & ~n39053 ;
  assign n41677 = n41676 ^ n791 ^ 1'b0 ;
  assign n41678 = n3779 ^ n2112 ^ 1'b0 ;
  assign n41679 = n12526 & ~n41678 ;
  assign n41680 = n3713 ^ n2435 ^ 1'b0 ;
  assign n41681 = n38975 ^ n2156 ^ 1'b0 ;
  assign n41682 = n5409 & n26205 ;
  assign n41690 = ~n5637 & n26341 ;
  assign n41683 = n513 & ~n1794 ;
  assign n41684 = n1794 & n41683 ;
  assign n41685 = n7817 ^ n1552 ^ 1'b0 ;
  assign n41686 = ~n41684 & n41685 ;
  assign n41687 = n8292 & n41686 ;
  assign n41688 = n5128 & n41687 ;
  assign n41689 = n41688 ^ n35336 ^ n15544 ;
  assign n41691 = n41690 ^ n41689 ^ 1'b0 ;
  assign n41692 = n378 & ~n16673 ;
  assign n41693 = ~n21522 & n41692 ;
  assign n41694 = n3104 & ~n23197 ;
  assign n41695 = n7148 & n7516 ;
  assign n41696 = n41695 ^ n33639 ^ 1'b0 ;
  assign n41697 = n1179 | n41696 ;
  assign n41698 = n19554 ^ n18387 ^ n3139 ;
  assign n41699 = n18229 & ~n41698 ;
  assign n41700 = n984 | n2005 ;
  assign n41701 = n41700 ^ n21989 ^ 1'b0 ;
  assign n41702 = n41275 ^ n11669 ^ 1'b0 ;
  assign n41703 = n6178 | n41702 ;
  assign n41704 = ~n280 & n35302 ;
  assign n41705 = ~n741 & n41704 ;
  assign n41706 = n11430 ^ n8548 ^ 1'b0 ;
  assign n41707 = n22687 | n30085 ;
  assign n41708 = n1096 | n29292 ;
  assign n41709 = ~n2318 & n41708 ;
  assign n41710 = n24329 & ~n30616 ;
  assign n41711 = n7348 & n13242 ;
  assign n41712 = n30536 ^ n246 ^ 1'b0 ;
  assign n41713 = n41711 & n41712 ;
  assign n41714 = n18517 ^ n9880 ^ 1'b0 ;
  assign n41715 = ( n15655 & n39249 ) | ( n15655 & n41714 ) | ( n39249 & n41714 ) ;
  assign n41716 = ~n1649 & n5616 ;
  assign n41717 = n1000 & n41716 ;
  assign n41718 = n13453 | n29976 ;
  assign n41719 = n4037 & n5245 ;
  assign n41720 = n29164 & n41719 ;
  assign n41721 = n573 | n2538 ;
  assign n41722 = ( n8189 & n35036 ) | ( n8189 & n41721 ) | ( n35036 & n41721 ) ;
  assign n41723 = n10058 & ~n17445 ;
  assign n41724 = n6863 | n41723 ;
  assign n41725 = n5330 | n21778 ;
  assign n41726 = n41725 ^ n940 ^ 1'b0 ;
  assign n41727 = n774 & ~n1025 ;
  assign n41728 = n1025 & n41727 ;
  assign n41729 = n41728 ^ n1491 ^ 1'b0 ;
  assign n41730 = n3186 | n41729 ;
  assign n41731 = n41730 ^ n27764 ^ 1'b0 ;
  assign n41732 = n36561 | n41731 ;
  assign n41733 = n9902 ^ n7336 ^ 1'b0 ;
  assign n41734 = n5716 & ~n41733 ;
  assign n41735 = n10266 & ~n41734 ;
  assign n41740 = n29019 & ~n41370 ;
  assign n41737 = n5018 & ~n5583 ;
  assign n41736 = n16300 | n30251 ;
  assign n41738 = n41737 ^ n41736 ^ 1'b0 ;
  assign n41739 = n41738 ^ n16826 ^ n6316 ;
  assign n41741 = n41740 ^ n41739 ^ n1887 ;
  assign n41742 = n7102 | n25186 ;
  assign n41743 = ~n5138 & n41742 ;
  assign y0 = x1 ;
  assign y1 = x2 ;
  assign y2 = x7 ;
  assign y3 = x8 ;
  assign y4 = x9 ;
  assign y5 = x11 ;
  assign y6 = ~1'b0 ;
  assign y7 = ~n14 ;
  assign y8 = n16 ;
  assign y9 = ~n17 ;
  assign y10 = ~1'b0 ;
  assign y11 = ~1'b0 ;
  assign y12 = 1'b0 ;
  assign y13 = ~1'b0 ;
  assign y14 = ~n19 ;
  assign y15 = ~1'b0 ;
  assign y16 = ~n25 ;
  assign y17 = n27 ;
  assign y18 = n28 ;
  assign y19 = ~1'b0 ;
  assign y20 = n36 ;
  assign y21 = ~n37 ;
  assign y22 = ~x8 ;
  assign y23 = ~1'b0 ;
  assign y24 = ~1'b0 ;
  assign y25 = ~n42 ;
  assign y26 = n44 ;
  assign y27 = n46 ;
  assign y28 = ~n48 ;
  assign y29 = n51 ;
  assign y30 = ~n53 ;
  assign y31 = n55 ;
  assign y32 = ~1'b0 ;
  assign y33 = ~1'b0 ;
  assign y34 = ~n58 ;
  assign y35 = ~n62 ;
  assign y36 = ~n70 ;
  assign y37 = n72 ;
  assign y38 = ~n76 ;
  assign y39 = ~n79 ;
  assign y40 = ~1'b0 ;
  assign y41 = ~1'b0 ;
  assign y42 = ~1'b0 ;
  assign y43 = n81 ;
  assign y44 = n82 ;
  assign y45 = ~n85 ;
  assign y46 = n87 ;
  assign y47 = ~n96 ;
  assign y48 = ~1'b0 ;
  assign y49 = n98 ;
  assign y50 = n104 ;
  assign y51 = n105 ;
  assign y52 = ~n106 ;
  assign y53 = n109 ;
  assign y54 = n111 ;
  assign y55 = n113 ;
  assign y56 = n114 ;
  assign y57 = ~n116 ;
  assign y58 = ~n117 ;
  assign y59 = ~n120 ;
  assign y60 = ~n125 ;
  assign y61 = ~1'b0 ;
  assign y62 = n129 ;
  assign y63 = ~n130 ;
  assign y64 = ~n131 ;
  assign y65 = ~1'b0 ;
  assign y66 = ~1'b0 ;
  assign y67 = ~n133 ;
  assign y68 = ~1'b0 ;
  assign y69 = ~n64 ;
  assign y70 = ~1'b0 ;
  assign y71 = ~n139 ;
  assign y72 = ~n142 ;
  assign y73 = ~1'b0 ;
  assign y74 = ~n146 ;
  assign y75 = ~n148 ;
  assign y76 = ~1'b0 ;
  assign y77 = n154 ;
  assign y78 = n155 ;
  assign y79 = n156 ;
  assign y80 = ~1'b0 ;
  assign y81 = ~1'b0 ;
  assign y82 = n157 ;
  assign y83 = ~n158 ;
  assign y84 = ~n163 ;
  assign y85 = ~1'b0 ;
  assign y86 = ~1'b0 ;
  assign y87 = ~1'b0 ;
  assign y88 = ~1'b0 ;
  assign y89 = ~1'b0 ;
  assign y90 = 1'b0 ;
  assign y91 = ~1'b0 ;
  assign y92 = 1'b0 ;
  assign y93 = ~n164 ;
  assign y94 = n165 ;
  assign y95 = ~n167 ;
  assign y96 = ~1'b0 ;
  assign y97 = ~1'b0 ;
  assign y98 = ~1'b0 ;
  assign y99 = n168 ;
  assign y100 = n139 ;
  assign y101 = ~n55 ;
  assign y102 = n170 ;
  assign y103 = ~1'b0 ;
  assign y104 = ~n174 ;
  assign y105 = ~1'b0 ;
  assign y106 = ~n175 ;
  assign y107 = ~1'b0 ;
  assign y108 = n178 ;
  assign y109 = ~n180 ;
  assign y110 = n182 ;
  assign y111 = n185 ;
  assign y112 = n186 ;
  assign y113 = ~1'b0 ;
  assign y114 = n188 ;
  assign y115 = ~1'b0 ;
  assign y116 = ~n190 ;
  assign y117 = 1'b0 ;
  assign y118 = ~1'b0 ;
  assign y119 = ~1'b0 ;
  assign y120 = ~n192 ;
  assign y121 = ~1'b0 ;
  assign y122 = n193 ;
  assign y123 = ~1'b0 ;
  assign y124 = n196 ;
  assign y125 = n197 ;
  assign y126 = ~1'b0 ;
  assign y127 = ~n198 ;
  assign y128 = n205 ;
  assign y129 = n185 ;
  assign y130 = ~1'b0 ;
  assign y131 = ~n206 ;
  assign y132 = n208 ;
  assign y133 = ~1'b0 ;
  assign y134 = ~1'b0 ;
  assign y135 = ~n210 ;
  assign y136 = ~1'b0 ;
  assign y137 = ~n212 ;
  assign y138 = ~1'b0 ;
  assign y139 = ~n215 ;
  assign y140 = ~n227 ;
  assign y141 = ~1'b0 ;
  assign y142 = ~n228 ;
  assign y143 = ~1'b0 ;
  assign y144 = ~1'b0 ;
  assign y145 = ~1'b0 ;
  assign y146 = n229 ;
  assign y147 = ~1'b0 ;
  assign y148 = ~n231 ;
  assign y149 = ~n23 ;
  assign y150 = ~n148 ;
  assign y151 = n233 ;
  assign y152 = ~n234 ;
  assign y153 = ~n161 ;
  assign y154 = ~1'b0 ;
  assign y155 = n235 ;
  assign y156 = ~n241 ;
  assign y157 = ~n244 ;
  assign y158 = ~n246 ;
  assign y159 = n247 ;
  assign y160 = ~n55 ;
  assign y161 = ~1'b0 ;
  assign y162 = ~1'b0 ;
  assign y163 = n251 ;
  assign y164 = n252 ;
  assign y165 = ~1'b0 ;
  assign y166 = n253 ;
  assign y167 = n254 ;
  assign y168 = ~n261 ;
  assign y169 = n265 ;
  assign y170 = ~n55 ;
  assign y171 = ~n270 ;
  assign y172 = n271 ;
  assign y173 = n272 ;
  assign y174 = ~x0 ;
  assign y175 = n273 ;
  assign y176 = n17 ;
  assign y177 = ~n277 ;
  assign y178 = ~1'b0 ;
  assign y179 = 1'b0 ;
  assign y180 = n278 ;
  assign y181 = ~n279 ;
  assign y182 = n283 ;
  assign y183 = ~x1 ;
  assign y184 = ~1'b0 ;
  assign y185 = ~1'b0 ;
  assign y186 = ~n284 ;
  assign y187 = ~1'b0 ;
  assign y188 = ~n286 ;
  assign y189 = n288 ;
  assign y190 = n291 ;
  assign y191 = ~x0 ;
  assign y192 = ~n293 ;
  assign y193 = ~n294 ;
  assign y194 = ~n295 ;
  assign y195 = ~n302 ;
  assign y196 = n309 ;
  assign y197 = ~n68 ;
  assign y198 = ~n310 ;
  assign y199 = ~1'b0 ;
  assign y200 = 1'b0 ;
  assign y201 = ~1'b0 ;
  assign y202 = n16 ;
  assign y203 = ~1'b0 ;
  assign y204 = n236 ;
  assign y205 = n311 ;
  assign y206 = ~1'b0 ;
  assign y207 = ~n313 ;
  assign y208 = n86 ;
  assign y209 = ~1'b0 ;
  assign y210 = ~1'b0 ;
  assign y211 = n102 ;
  assign y212 = n315 ;
  assign y213 = ~n316 ;
  assign y214 = ~1'b0 ;
  assign y215 = n114 ;
  assign y216 = ~1'b0 ;
  assign y217 = n268 ;
  assign y218 = n321 ;
  assign y219 = ~1'b0 ;
  assign y220 = ~n286 ;
  assign y221 = ~n322 ;
  assign y222 = ~n323 ;
  assign y223 = n327 ;
  assign y224 = ~1'b0 ;
  assign y225 = n328 ;
  assign y226 = ~1'b0 ;
  assign y227 = n333 ;
  assign y228 = ~n294 ;
  assign y229 = n335 ;
  assign y230 = ~1'b0 ;
  assign y231 = n337 ;
  assign y232 = n338 ;
  assign y233 = ~1'b0 ;
  assign y234 = n258 ;
  assign y235 = ~1'b0 ;
  assign y236 = n339 ;
  assign y237 = ~n340 ;
  assign y238 = n342 ;
  assign y239 = ~1'b0 ;
  assign y240 = ~n343 ;
  assign y241 = ~1'b0 ;
  assign y242 = ~n345 ;
  assign y243 = ~1'b0 ;
  assign y244 = ~n83 ;
  assign y245 = n350 ;
  assign y246 = ~n352 ;
  assign y247 = ~1'b0 ;
  assign y248 = ~1'b0 ;
  assign y249 = n359 ;
  assign y250 = ~1'b0 ;
  assign y251 = 1'b0 ;
  assign y252 = n361 ;
  assign y253 = ~n364 ;
  assign y254 = n366 ;
  assign y255 = ~1'b0 ;
  assign y256 = ~n374 ;
  assign y257 = ~1'b0 ;
  assign y258 = ~n375 ;
  assign y259 = ~n376 ;
  assign y260 = n142 ;
  assign y261 = ~1'b0 ;
  assign y262 = ~n133 ;
  assign y263 = 1'b0 ;
  assign y264 = n328 ;
  assign y265 = ~1'b0 ;
  assign y266 = n79 ;
  assign y267 = ~1'b0 ;
  assign y268 = n378 ;
  assign y269 = ~n381 ;
  assign y270 = ~n385 ;
  assign y271 = n389 ;
  assign y272 = ~1'b0 ;
  assign y273 = ~n169 ;
  assign y274 = ~n393 ;
  assign y275 = ~n395 ;
  assign y276 = n398 ;
  assign y277 = ~1'b0 ;
  assign y278 = 1'b0 ;
  assign y279 = ~1'b0 ;
  assign y280 = ~x3 ;
  assign y281 = ~1'b0 ;
  assign y282 = ~n405 ;
  assign y283 = ~1'b0 ;
  assign y284 = ~1'b0 ;
  assign y285 = ~1'b0 ;
  assign y286 = n37 ;
  assign y287 = ~n408 ;
  assign y288 = ~1'b0 ;
  assign y289 = ~n410 ;
  assign y290 = ~1'b0 ;
  assign y291 = n412 ;
  assign y292 = n415 ;
  assign y293 = ~n418 ;
  assign y294 = ~n419 ;
  assign y295 = ~1'b0 ;
  assign y296 = ~n425 ;
  assign y297 = n354 ;
  assign y298 = ~1'b0 ;
  assign y299 = 1'b0 ;
  assign y300 = ~1'b0 ;
  assign y301 = n427 ;
  assign y302 = ~n428 ;
  assign y303 = ~1'b0 ;
  assign y304 = ~n60 ;
  assign y305 = ~n432 ;
  assign y306 = ~1'b0 ;
  assign y307 = n433 ;
  assign y308 = ~1'b0 ;
  assign y309 = ~n434 ;
  assign y310 = n435 ;
  assign y311 = n437 ;
  assign y312 = ~n441 ;
  assign y313 = ~n442 ;
  assign y314 = ~n445 ;
  assign y315 = n205 ;
  assign y316 = 1'b0 ;
  assign y317 = ~n43 ;
  assign y318 = n448 ;
  assign y319 = ~1'b0 ;
  assign y320 = n450 ;
  assign y321 = ~1'b0 ;
  assign y322 = ~n455 ;
  assign y323 = ~n458 ;
  assign y324 = ~1'b0 ;
  assign y325 = ~n459 ;
  assign y326 = ~n461 ;
  assign y327 = 1'b0 ;
  assign y328 = 1'b0 ;
  assign y329 = n83 ;
  assign y330 = ~n462 ;
  assign y331 = n466 ;
  assign y332 = n468 ;
  assign y333 = ~n471 ;
  assign y334 = ~1'b0 ;
  assign y335 = 1'b0 ;
  assign y336 = ~n474 ;
  assign y337 = ~n475 ;
  assign y338 = n477 ;
  assign y339 = ~n294 ;
  assign y340 = ~1'b0 ;
  assign y341 = ~n478 ;
  assign y342 = ~n479 ;
  assign y343 = n482 ;
  assign y344 = n487 ;
  assign y345 = n488 ;
  assign y346 = ~1'b0 ;
  assign y347 = n489 ;
  assign y348 = ~n492 ;
  assign y349 = 1'b0 ;
  assign y350 = ~1'b0 ;
  assign y351 = ~1'b0 ;
  assign y352 = ~n493 ;
  assign y353 = ~1'b0 ;
  assign y354 = ~1'b0 ;
  assign y355 = ~1'b0 ;
  assign y356 = n495 ;
  assign y357 = n497 ;
  assign y358 = ~n500 ;
  assign y359 = ~n508 ;
  assign y360 = ~1'b0 ;
  assign y361 = ~n509 ;
  assign y362 = ~n510 ;
  assign y363 = ~1'b0 ;
  assign y364 = n233 ;
  assign y365 = n514 ;
  assign y366 = n518 ;
  assign y367 = ~n520 ;
  assign y368 = n524 ;
  assign y369 = ~1'b0 ;
  assign y370 = ~1'b0 ;
  assign y371 = ~1'b0 ;
  assign y372 = n526 ;
  assign y373 = n527 ;
  assign y374 = ~n528 ;
  assign y375 = ~1'b0 ;
  assign y376 = n532 ;
  assign y377 = ~n534 ;
  assign y378 = n535 ;
  assign y379 = ~n538 ;
  assign y380 = ~n169 ;
  assign y381 = ~n539 ;
  assign y382 = ~n540 ;
  assign y383 = n541 ;
  assign y384 = ~n177 ;
  assign y385 = ~1'b0 ;
  assign y386 = ~n542 ;
  assign y387 = ~1'b0 ;
  assign y388 = n544 ;
  assign y389 = ~n551 ;
  assign y390 = ~n390 ;
  assign y391 = n552 ;
  assign y392 = ~1'b0 ;
  assign y393 = ~1'b0 ;
  assign y394 = ~1'b0 ;
  assign y395 = n384 ;
  assign y396 = n555 ;
  assign y397 = ~n532 ;
  assign y398 = n66 ;
  assign y399 = ~n561 ;
  assign y400 = ~n562 ;
  assign y401 = ~1'b0 ;
  assign y402 = n564 ;
  assign y403 = ~1'b0 ;
  assign y404 = ~1'b0 ;
  assign y405 = ~n565 ;
  assign y406 = n489 ;
  assign y407 = ~n567 ;
  assign y408 = ~n158 ;
  assign y409 = n568 ;
  assign y410 = ~1'b0 ;
  assign y411 = n509 ;
  assign y412 = ~1'b0 ;
  assign y413 = n573 ;
  assign y414 = ~n575 ;
  assign y415 = ~n576 ;
  assign y416 = n580 ;
  assign y417 = ~1'b0 ;
  assign y418 = n582 ;
  assign y419 = n584 ;
  assign y420 = ~1'b0 ;
  assign y421 = ~n585 ;
  assign y422 = ~n588 ;
  assign y423 = ~n591 ;
  assign y424 = ~1'b0 ;
  assign y425 = 1'b0 ;
  assign y426 = n593 ;
  assign y427 = n596 ;
  assign y428 = ~n601 ;
  assign y429 = ~1'b0 ;
  assign y430 = 1'b0 ;
  assign y431 = n602 ;
  assign y432 = ~1'b0 ;
  assign y433 = n603 ;
  assign y434 = ~n608 ;
  assign y435 = ~1'b0 ;
  assign y436 = ~n609 ;
  assign y437 = ~1'b0 ;
  assign y438 = ~1'b0 ;
  assign y439 = ~1'b0 ;
  assign y440 = ~n615 ;
  assign y441 = n619 ;
  assign y442 = ~n621 ;
  assign y443 = ~1'b0 ;
  assign y444 = n622 ;
  assign y445 = n624 ;
  assign y446 = ~1'b0 ;
  assign y447 = ~n626 ;
  assign y448 = ~n627 ;
  assign y449 = ~n632 ;
  assign y450 = n634 ;
  assign y451 = ~n637 ;
  assign y452 = ~1'b0 ;
  assign y453 = ~1'b0 ;
  assign y454 = n638 ;
  assign y455 = n639 ;
  assign y456 = ~n640 ;
  assign y457 = ~n643 ;
  assign y458 = n456 ;
  assign y459 = ~1'b0 ;
  assign y460 = ~n644 ;
  assign y461 = ~n384 ;
  assign y462 = n647 ;
  assign y463 = ~n649 ;
  assign y464 = ~1'b0 ;
  assign y465 = ~1'b0 ;
  assign y466 = n653 ;
  assign y467 = ~n656 ;
  assign y468 = ~n68 ;
  assign y469 = ~1'b0 ;
  assign y470 = n659 ;
  assign y471 = n662 ;
  assign y472 = ~n663 ;
  assign y473 = ~n664 ;
  assign y474 = ~n665 ;
  assign y475 = n667 ;
  assign y476 = n670 ;
  assign y477 = n671 ;
  assign y478 = n400 ;
  assign y479 = n673 ;
  assign y480 = ~1'b0 ;
  assign y481 = ~n675 ;
  assign y482 = ~n678 ;
  assign y483 = n679 ;
  assign y484 = ~1'b0 ;
  assign y485 = ~1'b0 ;
  assign y486 = ~1'b0 ;
  assign y487 = n271 ;
  assign y488 = ~1'b0 ;
  assign y489 = ~n643 ;
  assign y490 = ~n681 ;
  assign y491 = ~1'b0 ;
  assign y492 = ~n683 ;
  assign y493 = ~n688 ;
  assign y494 = ~n689 ;
  assign y495 = n412 ;
  assign y496 = n697 ;
  assign y497 = ~1'b0 ;
  assign y498 = ~1'b0 ;
  assign y499 = 1'b0 ;
  assign y500 = ~1'b0 ;
  assign y501 = ~1'b0 ;
  assign y502 = ~n698 ;
  assign y503 = ~1'b0 ;
  assign y504 = ~1'b0 ;
  assign y505 = n699 ;
  assign y506 = n700 ;
  assign y507 = ~n78 ;
  assign y508 = ~n702 ;
  assign y509 = ~1'b0 ;
  assign y510 = n703 ;
  assign y511 = n704 ;
  assign y512 = ~n705 ;
  assign y513 = ~1'b0 ;
  assign y514 = n707 ;
  assign y515 = ~1'b0 ;
  assign y516 = ~1'b0 ;
  assign y517 = 1'b0 ;
  assign y518 = ~1'b0 ;
  assign y519 = ~1'b0 ;
  assign y520 = ~1'b0 ;
  assign y521 = ~n708 ;
  assign y522 = n113 ;
  assign y523 = n709 ;
  assign y524 = ~n60 ;
  assign y525 = n710 ;
  assign y526 = ~1'b0 ;
  assign y527 = ~1'b0 ;
  assign y528 = ~n712 ;
  assign y529 = ~n713 ;
  assign y530 = ~n608 ;
  assign y531 = n714 ;
  assign y532 = ~1'b0 ;
  assign y533 = ~n729 ;
  assign y534 = ~n330 ;
  assign y535 = ~1'b0 ;
  assign y536 = ~1'b0 ;
  assign y537 = n732 ;
  assign y538 = ~n740 ;
  assign y539 = ~n743 ;
  assign y540 = ~n744 ;
  assign y541 = ~1'b0 ;
  assign y542 = ~1'b0 ;
  assign y543 = ~n302 ;
  assign y544 = ~n747 ;
  assign y545 = ~n754 ;
  assign y546 = ~1'b0 ;
  assign y547 = ~1'b0 ;
  assign y548 = ~1'b0 ;
  assign y549 = ~1'b0 ;
  assign y550 = ~n508 ;
  assign y551 = ~n757 ;
  assign y552 = n760 ;
  assign y553 = n763 ;
  assign y554 = ~1'b0 ;
  assign y555 = ~1'b0 ;
  assign y556 = n765 ;
  assign y557 = n767 ;
  assign y558 = ~1'b0 ;
  assign y559 = ~1'b0 ;
  assign y560 = n770 ;
  assign y561 = ~1'b0 ;
  assign y562 = 1'b0 ;
  assign y563 = ~n772 ;
  assign y564 = ~1'b0 ;
  assign y565 = 1'b0 ;
  assign y566 = ~n773 ;
  assign y567 = n774 ;
  assign y568 = ~1'b0 ;
  assign y569 = ~1'b0 ;
  assign y570 = ~1'b0 ;
  assign y571 = ~1'b0 ;
  assign y572 = ~n782 ;
  assign y573 = ~n785 ;
  assign y574 = ~1'b0 ;
  assign y575 = n787 ;
  assign y576 = ~n792 ;
  assign y577 = ~1'b0 ;
  assign y578 = ~n794 ;
  assign y579 = ~n191 ;
  assign y580 = n798 ;
  assign y581 = n799 ;
  assign y582 = ~1'b0 ;
  assign y583 = ~1'b0 ;
  assign y584 = ~1'b0 ;
  assign y585 = n804 ;
  assign y586 = n806 ;
  assign y587 = ~n807 ;
  assign y588 = n810 ;
  assign y589 = ~n812 ;
  assign y590 = n364 ;
  assign y591 = ~n58 ;
  assign y592 = ~n813 ;
  assign y593 = n815 ;
  assign y594 = ~n817 ;
  assign y595 = ~n52 ;
  assign y596 = ~1'b0 ;
  assign y597 = ~n820 ;
  assign y598 = ~1'b0 ;
  assign y599 = n825 ;
  assign y600 = ~1'b0 ;
  assign y601 = ~1'b0 ;
  assign y602 = ~1'b0 ;
  assign y603 = n828 ;
  assign y604 = ~1'b0 ;
  assign y605 = n830 ;
  assign y606 = ~1'b0 ;
  assign y607 = ~n833 ;
  assign y608 = n839 ;
  assign y609 = ~n841 ;
  assign y610 = ~n843 ;
  assign y611 = ~n846 ;
  assign y612 = ~1'b0 ;
  assign y613 = ~1'b0 ;
  assign y614 = ~1'b0 ;
  assign y615 = ~1'b0 ;
  assign y616 = n688 ;
  assign y617 = ~n847 ;
  assign y618 = ~n853 ;
  assign y619 = ~n859 ;
  assign y620 = ~1'b0 ;
  assign y621 = ~1'b0 ;
  assign y622 = n861 ;
  assign y623 = ~1'b0 ;
  assign y624 = ~1'b0 ;
  assign y625 = n862 ;
  assign y626 = n869 ;
  assign y627 = 1'b0 ;
  assign y628 = n788 ;
  assign y629 = ~1'b0 ;
  assign y630 = ~n870 ;
  assign y631 = ~n273 ;
  assign y632 = n874 ;
  assign y633 = ~1'b0 ;
  assign y634 = ~n876 ;
  assign y635 = n878 ;
  assign y636 = ~n879 ;
  assign y637 = ~n882 ;
  assign y638 = ~n128 ;
  assign y639 = ~1'b0 ;
  assign y640 = ~n812 ;
  assign y641 = n883 ;
  assign y642 = ~1'b0 ;
  assign y643 = ~n890 ;
  assign y644 = n549 ;
  assign y645 = ~1'b0 ;
  assign y646 = ~1'b0 ;
  assign y647 = ~1'b0 ;
  assign y648 = n892 ;
  assign y649 = ~n153 ;
  assign y650 = n894 ;
  assign y651 = ~1'b0 ;
  assign y652 = ~1'b0 ;
  assign y653 = ~1'b0 ;
  assign y654 = n896 ;
  assign y655 = ~1'b0 ;
  assign y656 = ~1'b0 ;
  assign y657 = ~n906 ;
  assign y658 = ~1'b0 ;
  assign y659 = ~1'b0 ;
  assign y660 = ~n907 ;
  assign y661 = ~n833 ;
  assign y662 = n908 ;
  assign y663 = ~1'b0 ;
  assign y664 = ~n910 ;
  assign y665 = ~1'b0 ;
  assign y666 = ~n912 ;
  assign y667 = ~n683 ;
  assign y668 = n914 ;
  assign y669 = n921 ;
  assign y670 = ~n924 ;
  assign y671 = ~n927 ;
  assign y672 = ~1'b0 ;
  assign y673 = n83 ;
  assign y674 = ~1'b0 ;
  assign y675 = ~1'b0 ;
  assign y676 = ~1'b0 ;
  assign y677 = ~1'b0 ;
  assign y678 = ~n835 ;
  assign y679 = ~1'b0 ;
  assign y680 = n929 ;
  assign y681 = ~n932 ;
  assign y682 = ~n456 ;
  assign y683 = ~n694 ;
  assign y684 = ~n934 ;
  assign y685 = ~n935 ;
  assign y686 = ~1'b0 ;
  assign y687 = ~1'b0 ;
  assign y688 = ~1'b0 ;
  assign y689 = ~n940 ;
  assign y690 = ~1'b0 ;
  assign y691 = n944 ;
  assign y692 = n949 ;
  assign y693 = ~n951 ;
  assign y694 = ~1'b0 ;
  assign y695 = n955 ;
  assign y696 = n296 ;
  assign y697 = n553 ;
  assign y698 = ~n958 ;
  assign y699 = n960 ;
  assign y700 = ~n961 ;
  assign y701 = ~n963 ;
  assign y702 = ~n964 ;
  assign y703 = n966 ;
  assign y704 = ~n158 ;
  assign y705 = ~1'b0 ;
  assign y706 = 1'b0 ;
  assign y707 = n973 ;
  assign y708 = ~1'b0 ;
  assign y709 = 1'b0 ;
  assign y710 = ~n974 ;
  assign y711 = ~1'b0 ;
  assign y712 = n975 ;
  assign y713 = n977 ;
  assign y714 = ~1'b0 ;
  assign y715 = ~1'b0 ;
  assign y716 = n980 ;
  assign y717 = ~n983 ;
  assign y718 = n984 ;
  assign y719 = 1'b0 ;
  assign y720 = ~n986 ;
  assign y721 = ~n988 ;
  assign y722 = ~1'b0 ;
  assign y723 = ~1'b0 ;
  assign y724 = ~1'b0 ;
  assign y725 = ~1'b0 ;
  assign y726 = n993 ;
  assign y727 = 1'b0 ;
  assign y728 = n998 ;
  assign y729 = n1000 ;
  assign y730 = n938 ;
  assign y731 = ~n1001 ;
  assign y732 = ~n1002 ;
  assign y733 = ~1'b0 ;
  assign y734 = ~n1003 ;
  assign y735 = ~1'b0 ;
  assign y736 = n1005 ;
  assign y737 = ~1'b0 ;
  assign y738 = n1008 ;
  assign y739 = n1013 ;
  assign y740 = ~n1015 ;
  assign y741 = ~n1016 ;
  assign y742 = ~1'b0 ;
  assign y743 = ~n1020 ;
  assign y744 = ~1'b0 ;
  assign y745 = n618 ;
  assign y746 = n1022 ;
  assign y747 = n1024 ;
  assign y748 = ~1'b0 ;
  assign y749 = ~n1025 ;
  assign y750 = n1031 ;
  assign y751 = ~1'b0 ;
  assign y752 = ~1'b0 ;
  assign y753 = ~n1034 ;
  assign y754 = ~n1036 ;
  assign y755 = ~n1039 ;
  assign y756 = ~1'b0 ;
  assign y757 = n1041 ;
  assign y758 = ~n1043 ;
  assign y759 = ~n1047 ;
  assign y760 = ~1'b0 ;
  assign y761 = ~n833 ;
  assign y762 = ~n1048 ;
  assign y763 = ~1'b0 ;
  assign y764 = n1049 ;
  assign y765 = ~n1050 ;
  assign y766 = ~1'b0 ;
  assign y767 = ~1'b0 ;
  assign y768 = ~1'b0 ;
  assign y769 = 1'b0 ;
  assign y770 = ~1'b0 ;
  assign y771 = n1051 ;
  assign y772 = n1052 ;
  assign y773 = ~n322 ;
  assign y774 = ~1'b0 ;
  assign y775 = n1053 ;
  assign y776 = ~n1054 ;
  assign y777 = ~n622 ;
  assign y778 = ~n1056 ;
  assign y779 = ~n1058 ;
  assign y780 = ~1'b0 ;
  assign y781 = ~1'b0 ;
  assign y782 = ~1'b0 ;
  assign y783 = ~1'b0 ;
  assign y784 = ~n1059 ;
  assign y785 = ~1'b0 ;
  assign y786 = n530 ;
  assign y787 = ~n1066 ;
  assign y788 = ~1'b0 ;
  assign y789 = ~n1067 ;
  assign y790 = ~1'b0 ;
  assign y791 = n1069 ;
  assign y792 = ~1'b0 ;
  assign y793 = ~n1077 ;
  assign y794 = ~n1078 ;
  assign y795 = n1079 ;
  assign y796 = ~1'b0 ;
  assign y797 = ~n325 ;
  assign y798 = n1083 ;
  assign y799 = ~n1086 ;
  assign y800 = 1'b0 ;
  assign y801 = ~n1088 ;
  assign y802 = n1089 ;
  assign y803 = n1096 ;
  assign y804 = ~n1097 ;
  assign y805 = ~n1098 ;
  assign y806 = ~1'b0 ;
  assign y807 = ~n1103 ;
  assign y808 = n1106 ;
  assign y809 = ~n1109 ;
  assign y810 = ~1'b0 ;
  assign y811 = n1110 ;
  assign y812 = ~n158 ;
  assign y813 = n1112 ;
  assign y814 = ~n1113 ;
  assign y815 = ~n1115 ;
  assign y816 = ~n1117 ;
  assign y817 = ~n1118 ;
  assign y818 = 1'b0 ;
  assign y819 = n1119 ;
  assign y820 = 1'b0 ;
  assign y821 = 1'b0 ;
  assign y822 = 1'b0 ;
  assign y823 = ~1'b0 ;
  assign y824 = ~n1089 ;
  assign y825 = ~1'b0 ;
  assign y826 = n1121 ;
  assign y827 = ~1'b0 ;
  assign y828 = n1129 ;
  assign y829 = n1130 ;
  assign y830 = ~1'b0 ;
  assign y831 = ~n1132 ;
  assign y832 = n1134 ;
  assign y833 = ~1'b0 ;
  assign y834 = 1'b0 ;
  assign y835 = ~1'b0 ;
  assign y836 = ~n1138 ;
  assign y837 = ~n1139 ;
  assign y838 = n1141 ;
  assign y839 = ~n1143 ;
  assign y840 = ~1'b0 ;
  assign y841 = ~1'b0 ;
  assign y842 = ~1'b0 ;
  assign y843 = n1144 ;
  assign y844 = ~n1148 ;
  assign y845 = ~1'b0 ;
  assign y846 = ~1'b0 ;
  assign y847 = ~1'b0 ;
  assign y848 = ~1'b0 ;
  assign y849 = n1151 ;
  assign y850 = ~1'b0 ;
  assign y851 = ~n599 ;
  assign y852 = ~1'b0 ;
  assign y853 = ~1'b0 ;
  assign y854 = 1'b0 ;
  assign y855 = n1152 ;
  assign y856 = n1157 ;
  assign y857 = ~1'b0 ;
  assign y858 = n1161 ;
  assign y859 = ~1'b0 ;
  assign y860 = ~n1162 ;
  assign y861 = ~1'b0 ;
  assign y862 = ~1'b0 ;
  assign y863 = ~n1163 ;
  assign y864 = ~1'b0 ;
  assign y865 = ~1'b0 ;
  assign y866 = ~n1164 ;
  assign y867 = 1'b0 ;
  assign y868 = n1166 ;
  assign y869 = ~1'b0 ;
  assign y870 = ~n1170 ;
  assign y871 = n1179 ;
  assign y872 = n1133 ;
  assign y873 = ~1'b0 ;
  assign y874 = ~n1183 ;
  assign y875 = ~1'b0 ;
  assign y876 = ~n1184 ;
  assign y877 = ~1'b0 ;
  assign y878 = ~1'b0 ;
  assign y879 = ~1'b0 ;
  assign y880 = ~n1185 ;
  assign y881 = ~1'b0 ;
  assign y882 = ~1'b0 ;
  assign y883 = n1192 ;
  assign y884 = ~n1193 ;
  assign y885 = ~1'b0 ;
  assign y886 = n1194 ;
  assign y887 = ~n1197 ;
  assign y888 = ~n1201 ;
  assign y889 = 1'b0 ;
  assign y890 = n1202 ;
  assign y891 = ~1'b0 ;
  assign y892 = ~1'b0 ;
  assign y893 = ~n1206 ;
  assign y894 = ~1'b0 ;
  assign y895 = ~1'b0 ;
  assign y896 = ~n1208 ;
  assign y897 = n1209 ;
  assign y898 = n1210 ;
  assign y899 = ~n1212 ;
  assign y900 = ~n1213 ;
  assign y901 = n1214 ;
  assign y902 = n1218 ;
  assign y903 = ~1'b0 ;
  assign y904 = ~1'b0 ;
  assign y905 = n1220 ;
  assign y906 = n1222 ;
  assign y907 = ~1'b0 ;
  assign y908 = ~1'b0 ;
  assign y909 = ~1'b0 ;
  assign y910 = ~1'b0 ;
  assign y911 = ~1'b0 ;
  assign y912 = ~1'b0 ;
  assign y913 = n1223 ;
  assign y914 = n1224 ;
  assign y915 = n1226 ;
  assign y916 = ~n1229 ;
  assign y917 = ~1'b0 ;
  assign y918 = n229 ;
  assign y919 = n1230 ;
  assign y920 = ~n1231 ;
  assign y921 = ~n1232 ;
  assign y922 = ~1'b0 ;
  assign y923 = ~1'b0 ;
  assign y924 = ~n1239 ;
  assign y925 = 1'b0 ;
  assign y926 = n1246 ;
  assign y927 = ~n1249 ;
  assign y928 = n1250 ;
  assign y929 = ~n1257 ;
  assign y930 = n1260 ;
  assign y931 = ~n1262 ;
  assign y932 = ~1'b0 ;
  assign y933 = ~n1264 ;
  assign y934 = ~1'b0 ;
  assign y935 = ~1'b0 ;
  assign y936 = n1267 ;
  assign y937 = n1268 ;
  assign y938 = ~n1270 ;
  assign y939 = n1276 ;
  assign y940 = n1277 ;
  assign y941 = ~1'b0 ;
  assign y942 = ~1'b0 ;
  assign y943 = 1'b0 ;
  assign y944 = ~1'b0 ;
  assign y945 = n1280 ;
  assign y946 = ~1'b0 ;
  assign y947 = ~n1284 ;
  assign y948 = n1285 ;
  assign y949 = n1287 ;
  assign y950 = ~n1289 ;
  assign y951 = n1291 ;
  assign y952 = n1292 ;
  assign y953 = ~n1297 ;
  assign y954 = ~1'b0 ;
  assign y955 = ~1'b0 ;
  assign y956 = n1298 ;
  assign y957 = ~1'b0 ;
  assign y958 = ~1'b0 ;
  assign y959 = n1192 ;
  assign y960 = ~1'b0 ;
  assign y961 = n1302 ;
  assign y962 = ~1'b0 ;
  assign y963 = ~n1303 ;
  assign y964 = ~1'b0 ;
  assign y965 = ~1'b0 ;
  assign y966 = ~n310 ;
  assign y967 = 1'b0 ;
  assign y968 = ~n1307 ;
  assign y969 = ~1'b0 ;
  assign y970 = ~n1308 ;
  assign y971 = ~n1318 ;
  assign y972 = ~1'b0 ;
  assign y973 = ~n1322 ;
  assign y974 = ~1'b0 ;
  assign y975 = ~1'b0 ;
  assign y976 = ~1'b0 ;
  assign y977 = ~1'b0 ;
  assign y978 = ~1'b0 ;
  assign y979 = ~1'b0 ;
  assign y980 = 1'b0 ;
  assign y981 = ~n1325 ;
  assign y982 = ~1'b0 ;
  assign y983 = n1326 ;
  assign y984 = ~n1329 ;
  assign y985 = n1331 ;
  assign y986 = n1332 ;
  assign y987 = n1334 ;
  assign y988 = ~x5 ;
  assign y989 = ~1'b0 ;
  assign y990 = n1335 ;
  assign y991 = ~n1337 ;
  assign y992 = ~1'b0 ;
  assign y993 = n1341 ;
  assign y994 = n1345 ;
  assign y995 = n1346 ;
  assign y996 = ~1'b0 ;
  assign y997 = ~n1347 ;
  assign y998 = ~n1349 ;
  assign y999 = 1'b0 ;
  assign y1000 = n1354 ;
  assign y1001 = ~n1357 ;
  assign y1002 = n1359 ;
  assign y1003 = ~n19 ;
  assign y1004 = ~n1360 ;
  assign y1005 = 1'b0 ;
  assign y1006 = n1367 ;
  assign y1007 = ~1'b0 ;
  assign y1008 = ~1'b0 ;
  assign y1009 = n1368 ;
  assign y1010 = ~1'b0 ;
  assign y1011 = n216 ;
  assign y1012 = n157 ;
  assign y1013 = n1370 ;
  assign y1014 = ~1'b0 ;
  assign y1015 = n1377 ;
  assign y1016 = ~n1379 ;
  assign y1017 = ~1'b0 ;
  assign y1018 = n1384 ;
  assign y1019 = n1385 ;
  assign y1020 = ~n1044 ;
  assign y1021 = ~n1388 ;
  assign y1022 = ~1'b0 ;
  assign y1023 = ~1'b0 ;
  assign y1024 = ~1'b0 ;
  assign y1025 = ~n1392 ;
  assign y1026 = ~1'b0 ;
  assign y1027 = ~n1401 ;
  assign y1028 = n1406 ;
  assign y1029 = 1'b0 ;
  assign y1030 = ~1'b0 ;
  assign y1031 = n1161 ;
  assign y1032 = ~n1410 ;
  assign y1033 = ~n566 ;
  assign y1034 = n1411 ;
  assign y1035 = n1414 ;
  assign y1036 = ~1'b0 ;
  assign y1037 = ~n1416 ;
  assign y1038 = ~n1418 ;
  assign y1039 = ~n38 ;
  assign y1040 = ~1'b0 ;
  assign y1041 = ~n1428 ;
  assign y1042 = ~n1429 ;
  assign y1043 = ~n1431 ;
  assign y1044 = ~1'b0 ;
  assign y1045 = ~n1437 ;
  assign y1046 = 1'b0 ;
  assign y1047 = 1'b0 ;
  assign y1048 = ~n1438 ;
  assign y1049 = n1439 ;
  assign y1050 = ~1'b0 ;
  assign y1051 = ~1'b0 ;
  assign y1052 = ~n1130 ;
  assign y1053 = ~n1440 ;
  assign y1054 = ~1'b0 ;
  assign y1055 = ~n1445 ;
  assign y1056 = ~1'b0 ;
  assign y1057 = n1447 ;
  assign y1058 = ~n1450 ;
  assign y1059 = n671 ;
  assign y1060 = ~1'b0 ;
  assign y1061 = 1'b0 ;
  assign y1062 = ~1'b0 ;
  assign y1063 = n1455 ;
  assign y1064 = ~n1462 ;
  assign y1065 = ~n977 ;
  assign y1066 = ~1'b0 ;
  assign y1067 = n1463 ;
  assign y1068 = ~n1464 ;
  assign y1069 = ~n1465 ;
  assign y1070 = ~n1472 ;
  assign y1071 = ~1'b0 ;
  assign y1072 = n1475 ;
  assign y1073 = n1477 ;
  assign y1074 = ~1'b0 ;
  assign y1075 = 1'b0 ;
  assign y1076 = ~1'b0 ;
  assign y1077 = ~n1478 ;
  assign y1078 = ~n257 ;
  assign y1079 = ~n1480 ;
  assign y1080 = ~n1484 ;
  assign y1081 = ~1'b0 ;
  assign y1082 = ~1'b0 ;
  assign y1083 = n1487 ;
  assign y1084 = ~1'b0 ;
  assign y1085 = ~n1492 ;
  assign y1086 = n1493 ;
  assign y1087 = ~1'b0 ;
  assign y1088 = 1'b0 ;
  assign y1089 = ~n1496 ;
  assign y1090 = ~n1497 ;
  assign y1091 = 1'b0 ;
  assign y1092 = n1504 ;
  assign y1093 = 1'b0 ;
  assign y1094 = ~n1505 ;
  assign y1095 = ~1'b0 ;
  assign y1096 = ~1'b0 ;
  assign y1097 = ~1'b0 ;
  assign y1098 = ~1'b0 ;
  assign y1099 = ~1'b0 ;
  assign y1100 = ~n1508 ;
  assign y1101 = ~1'b0 ;
  assign y1102 = ~1'b0 ;
  assign y1103 = ~1'b0 ;
  assign y1104 = ~1'b0 ;
  assign y1105 = ~n1511 ;
  assign y1106 = n1512 ;
  assign y1107 = ~n1513 ;
  assign y1108 = 1'b0 ;
  assign y1109 = ~1'b0 ;
  assign y1110 = ~1'b0 ;
  assign y1111 = ~n1515 ;
  assign y1112 = ~1'b0 ;
  assign y1113 = ~1'b0 ;
  assign y1114 = n1516 ;
  assign y1115 = ~n164 ;
  assign y1116 = ~1'b0 ;
  assign y1117 = n1518 ;
  assign y1118 = n470 ;
  assign y1119 = n1519 ;
  assign y1120 = ~n1523 ;
  assign y1121 = n228 ;
  assign y1122 = ~n1526 ;
  assign y1123 = n1527 ;
  assign y1124 = ~1'b0 ;
  assign y1125 = n1529 ;
  assign y1126 = ~1'b0 ;
  assign y1127 = n663 ;
  assign y1128 = n1530 ;
  assign y1129 = n1537 ;
  assign y1130 = ~n1538 ;
  assign y1131 = ~1'b0 ;
  assign y1132 = ~n1539 ;
  assign y1133 = n1227 ;
  assign y1134 = ~1'b0 ;
  assign y1135 = n1541 ;
  assign y1136 = ~n1545 ;
  assign y1137 = ~1'b0 ;
  assign y1138 = n1550 ;
  assign y1139 = ~1'b0 ;
  assign y1140 = ~n1552 ;
  assign y1141 = ~n1559 ;
  assign y1142 = ~1'b0 ;
  assign y1143 = ~n1560 ;
  assign y1144 = n1566 ;
  assign y1145 = ~n1571 ;
  assign y1146 = n1579 ;
  assign y1147 = ~n1581 ;
  assign y1148 = ~n1582 ;
  assign y1149 = 1'b0 ;
  assign y1150 = ~1'b0 ;
  assign y1151 = ~1'b0 ;
  assign y1152 = ~1'b0 ;
  assign y1153 = ~n616 ;
  assign y1154 = ~n1588 ;
  assign y1155 = n1591 ;
  assign y1156 = n337 ;
  assign y1157 = n1593 ;
  assign y1158 = ~1'b0 ;
  assign y1159 = ~1'b0 ;
  assign y1160 = ~1'b0 ;
  assign y1161 = ~1'b0 ;
  assign y1162 = ~n1597 ;
  assign y1163 = n1599 ;
  assign y1164 = ~n1602 ;
  assign y1165 = n1604 ;
  assign y1166 = ~1'b0 ;
  assign y1167 = ~1'b0 ;
  assign y1168 = n1609 ;
  assign y1169 = ~1'b0 ;
  assign y1170 = ~1'b0 ;
  assign y1171 = n1615 ;
  assign y1172 = ~n1622 ;
  assign y1173 = ~1'b0 ;
  assign y1174 = n1624 ;
  assign y1175 = 1'b0 ;
  assign y1176 = ~1'b0 ;
  assign y1177 = ~1'b0 ;
  assign y1178 = n1626 ;
  assign y1179 = ~1'b0 ;
  assign y1180 = n1627 ;
  assign y1181 = n1629 ;
  assign y1182 = n1630 ;
  assign y1183 = n336 ;
  assign y1184 = n715 ;
  assign y1185 = n1631 ;
  assign y1186 = ~1'b0 ;
  assign y1187 = ~n1632 ;
  assign y1188 = ~n1634 ;
  assign y1189 = ~1'b0 ;
  assign y1190 = ~1'b0 ;
  assign y1191 = ~n1159 ;
  assign y1192 = ~n1635 ;
  assign y1193 = ~n1638 ;
  assign y1194 = n1640 ;
  assign y1195 = 1'b0 ;
  assign y1196 = ~1'b0 ;
  assign y1197 = n1642 ;
  assign y1198 = ~1'b0 ;
  assign y1199 = n1645 ;
  assign y1200 = n1649 ;
  assign y1201 = ~1'b0 ;
  assign y1202 = ~n776 ;
  assign y1203 = ~1'b0 ;
  assign y1204 = ~n1650 ;
  assign y1205 = n1655 ;
  assign y1206 = n1656 ;
  assign y1207 = n1658 ;
  assign y1208 = ~n290 ;
  assign y1209 = ~n1660 ;
  assign y1210 = n1664 ;
  assign y1211 = n1666 ;
  assign y1212 = ~1'b0 ;
  assign y1213 = n1669 ;
  assign y1214 = 1'b0 ;
  assign y1215 = ~1'b0 ;
  assign y1216 = ~1'b0 ;
  assign y1217 = ~n1671 ;
  assign y1218 = ~1'b0 ;
  assign y1219 = ~1'b0 ;
  assign y1220 = ~n1676 ;
  assign y1221 = ~1'b0 ;
  assign y1222 = n1681 ;
  assign y1223 = ~1'b0 ;
  assign y1224 = ~1'b0 ;
  assign y1225 = 1'b0 ;
  assign y1226 = n1683 ;
  assign y1227 = n1687 ;
  assign y1228 = ~1'b0 ;
  assign y1229 = n1663 ;
  assign y1230 = ~n1688 ;
  assign y1231 = ~n1691 ;
  assign y1232 = ~n1692 ;
  assign y1233 = 1'b0 ;
  assign y1234 = ~n1693 ;
  assign y1235 = ~1'b0 ;
  assign y1236 = ~1'b0 ;
  assign y1237 = 1'b0 ;
  assign y1238 = ~1'b0 ;
  assign y1239 = ~1'b0 ;
  assign y1240 = ~n119 ;
  assign y1241 = ~1'b0 ;
  assign y1242 = ~1'b0 ;
  assign y1243 = ~n158 ;
  assign y1244 = n1695 ;
  assign y1245 = n1697 ;
  assign y1246 = n1699 ;
  assign y1247 = ~1'b0 ;
  assign y1248 = n1701 ;
  assign y1249 = ~1'b0 ;
  assign y1250 = n1702 ;
  assign y1251 = ~1'b0 ;
  assign y1252 = ~n1705 ;
  assign y1253 = ~n1708 ;
  assign y1254 = ~n1709 ;
  assign y1255 = ~n1710 ;
  assign y1256 = ~1'b0 ;
  assign y1257 = ~n1711 ;
  assign y1258 = ~1'b0 ;
  assign y1259 = ~n1712 ;
  assign y1260 = n1713 ;
  assign y1261 = ~1'b0 ;
  assign y1262 = n94 ;
  assign y1263 = 1'b0 ;
  assign y1264 = n1715 ;
  assign y1265 = ~n1720 ;
  assign y1266 = ~1'b0 ;
  assign y1267 = n1721 ;
  assign y1268 = ~n1722 ;
  assign y1269 = n1728 ;
  assign y1270 = ~n1730 ;
  assign y1271 = ~1'b0 ;
  assign y1272 = ~n1732 ;
  assign y1273 = ~n1662 ;
  assign y1274 = n1734 ;
  assign y1275 = ~1'b0 ;
  assign y1276 = ~n68 ;
  assign y1277 = ~1'b0 ;
  assign y1278 = n1688 ;
  assign y1279 = n1736 ;
  assign y1280 = ~1'b0 ;
  assign y1281 = ~1'b0 ;
  assign y1282 = ~1'b0 ;
  assign y1283 = ~n1737 ;
  assign y1284 = ~1'b0 ;
  assign y1285 = ~n1740 ;
  assign y1286 = ~n1743 ;
  assign y1287 = n1745 ;
  assign y1288 = ~1'b0 ;
  assign y1289 = ~1'b0 ;
  assign y1290 = ~1'b0 ;
  assign y1291 = ~1'b0 ;
  assign y1292 = ~1'b0 ;
  assign y1293 = n1747 ;
  assign y1294 = n1750 ;
  assign y1295 = ~n1751 ;
  assign y1296 = 1'b0 ;
  assign y1297 = n1756 ;
  assign y1298 = n1757 ;
  assign y1299 = n1759 ;
  assign y1300 = ~n1764 ;
  assign y1301 = ~1'b0 ;
  assign y1302 = n1765 ;
  assign y1303 = ~1'b0 ;
  assign y1304 = ~1'b0 ;
  assign y1305 = ~1'b0 ;
  assign y1306 = ~n1766 ;
  assign y1307 = ~1'b0 ;
  assign y1308 = ~1'b0 ;
  assign y1309 = n1768 ;
  assign y1310 = ~1'b0 ;
  assign y1311 = ~1'b0 ;
  assign y1312 = ~1'b0 ;
  assign y1313 = n1770 ;
  assign y1314 = n1774 ;
  assign y1315 = ~1'b0 ;
  assign y1316 = ~1'b0 ;
  assign y1317 = ~n1779 ;
  assign y1318 = ~1'b0 ;
  assign y1319 = ~1'b0 ;
  assign y1320 = n1783 ;
  assign y1321 = n1786 ;
  assign y1322 = ~1'b0 ;
  assign y1323 = ~n15 ;
  assign y1324 = ~n1790 ;
  assign y1325 = ~n1791 ;
  assign y1326 = ~n1792 ;
  assign y1327 = 1'b0 ;
  assign y1328 = ~n1794 ;
  assign y1329 = n1800 ;
  assign y1330 = n1802 ;
  assign y1331 = ~n1807 ;
  assign y1332 = ~1'b0 ;
  assign y1333 = ~n1811 ;
  assign y1334 = ~1'b0 ;
  assign y1335 = n1815 ;
  assign y1336 = ~1'b0 ;
  assign y1337 = n1816 ;
  assign y1338 = ~n1817 ;
  assign y1339 = n1818 ;
  assign y1340 = ~1'b0 ;
  assign y1341 = n1820 ;
  assign y1342 = n1821 ;
  assign y1343 = n159 ;
  assign y1344 = ~1'b0 ;
  assign y1345 = ~1'b0 ;
  assign y1346 = n1826 ;
  assign y1347 = n628 ;
  assign y1348 = n1827 ;
  assign y1349 = ~n1828 ;
  assign y1350 = ~1'b0 ;
  assign y1351 = ~n1829 ;
  assign y1352 = n1831 ;
  assign y1353 = ~n1832 ;
  assign y1354 = ~n1833 ;
  assign y1355 = n1838 ;
  assign y1356 = ~n1839 ;
  assign y1357 = ~n1840 ;
  assign y1358 = ~1'b0 ;
  assign y1359 = ~1'b0 ;
  assign y1360 = n1841 ;
  assign y1361 = ~n1844 ;
  assign y1362 = ~1'b0 ;
  assign y1363 = ~n1845 ;
  assign y1364 = n1847 ;
  assign y1365 = 1'b0 ;
  assign y1366 = n1851 ;
  assign y1367 = ~1'b0 ;
  assign y1368 = n1852 ;
  assign y1369 = ~1'b0 ;
  assign y1370 = ~1'b0 ;
  assign y1371 = n1856 ;
  assign y1372 = n1857 ;
  assign y1373 = ~n1858 ;
  assign y1374 = n1859 ;
  assign y1375 = ~1'b0 ;
  assign y1376 = ~n1864 ;
  assign y1377 = n86 ;
  assign y1378 = ~n1867 ;
  assign y1379 = ~1'b0 ;
  assign y1380 = n246 ;
  assign y1381 = ~1'b0 ;
  assign y1382 = ~1'b0 ;
  assign y1383 = ~1'b0 ;
  assign y1384 = ~1'b0 ;
  assign y1385 = n1868 ;
  assign y1386 = n832 ;
  assign y1387 = n1873 ;
  assign y1388 = n1874 ;
  assign y1389 = ~n1875 ;
  assign y1390 = ~1'b0 ;
  assign y1391 = ~n1878 ;
  assign y1392 = n1491 ;
  assign y1393 = ~1'b0 ;
  assign y1394 = ~1'b0 ;
  assign y1395 = ~1'b0 ;
  assign y1396 = ~1'b0 ;
  assign y1397 = ~n1880 ;
  assign y1398 = 1'b0 ;
  assign y1399 = ~1'b0 ;
  assign y1400 = n1883 ;
  assign y1401 = ~1'b0 ;
  assign y1402 = 1'b0 ;
  assign y1403 = ~1'b0 ;
  assign y1404 = ~1'b0 ;
  assign y1405 = ~1'b0 ;
  assign y1406 = ~n1884 ;
  assign y1407 = ~n1866 ;
  assign y1408 = ~1'b0 ;
  assign y1409 = ~1'b0 ;
  assign y1410 = ~1'b0 ;
  assign y1411 = ~n1885 ;
  assign y1412 = n1887 ;
  assign y1413 = ~n1888 ;
  assign y1414 = ~1'b0 ;
  assign y1415 = ~1'b0 ;
  assign y1416 = ~1'b0 ;
  assign y1417 = ~n1893 ;
  assign y1418 = 1'b0 ;
  assign y1419 = ~1'b0 ;
  assign y1420 = ~n1895 ;
  assign y1421 = ~1'b0 ;
  assign y1422 = n1899 ;
  assign y1423 = n1901 ;
  assign y1424 = ~n1902 ;
  assign y1425 = ~n1112 ;
  assign y1426 = 1'b0 ;
  assign y1427 = ~n1906 ;
  assign y1428 = ~n1907 ;
  assign y1429 = ~n1909 ;
  assign y1430 = ~n1918 ;
  assign y1431 = ~n587 ;
  assign y1432 = n1668 ;
  assign y1433 = ~n1008 ;
  assign y1434 = n1926 ;
  assign y1435 = n1927 ;
  assign y1436 = n1928 ;
  assign y1437 = n1931 ;
  assign y1438 = ~1'b0 ;
  assign y1439 = n954 ;
  assign y1440 = ~n1192 ;
  assign y1441 = n1932 ;
  assign y1442 = ~n469 ;
  assign y1443 = ~1'b0 ;
  assign y1444 = n1710 ;
  assign y1445 = ~1'b0 ;
  assign y1446 = n1933 ;
  assign y1447 = ~n1935 ;
  assign y1448 = ~1'b0 ;
  assign y1449 = ~n1936 ;
  assign y1450 = ~1'b0 ;
  assign y1451 = ~n184 ;
  assign y1452 = ~1'b0 ;
  assign y1453 = ~n1939 ;
  assign y1454 = ~n175 ;
  assign y1455 = n1940 ;
  assign y1456 = ~1'b0 ;
  assign y1457 = n1943 ;
  assign y1458 = ~1'b0 ;
  assign y1459 = ~1'b0 ;
  assign y1460 = n1944 ;
  assign y1461 = ~n1946 ;
  assign y1462 = ~n1947 ;
  assign y1463 = n1949 ;
  assign y1464 = ~1'b0 ;
  assign y1465 = ~1'b0 ;
  assign y1466 = n1950 ;
  assign y1467 = n1954 ;
  assign y1468 = ~1'b0 ;
  assign y1469 = ~n1956 ;
  assign y1470 = n1957 ;
  assign y1471 = n1959 ;
  assign y1472 = ~1'b0 ;
  assign y1473 = n1960 ;
  assign y1474 = n1963 ;
  assign y1475 = ~n1964 ;
  assign y1476 = ~1'b0 ;
  assign y1477 = ~1'b0 ;
  assign y1478 = ~1'b0 ;
  assign y1479 = ~n1966 ;
  assign y1480 = n1970 ;
  assign y1481 = ~n1246 ;
  assign y1482 = ~n832 ;
  assign y1483 = ~n1971 ;
  assign y1484 = ~1'b0 ;
  assign y1485 = ~1'b0 ;
  assign y1486 = ~n1976 ;
  assign y1487 = n1984 ;
  assign y1488 = ~n1986 ;
  assign y1489 = ~1'b0 ;
  assign y1490 = ~n1990 ;
  assign y1491 = n1992 ;
  assign y1492 = n1994 ;
  assign y1493 = ~n1097 ;
  assign y1494 = n1997 ;
  assign y1495 = ~1'b0 ;
  assign y1496 = n2004 ;
  assign y1497 = ~n2005 ;
  assign y1498 = n2007 ;
  assign y1499 = ~1'b0 ;
  assign y1500 = ~1'b0 ;
  assign y1501 = ~n2010 ;
  assign y1502 = ~1'b0 ;
  assign y1503 = ~1'b0 ;
  assign y1504 = ~n2011 ;
  assign y1505 = ~n2012 ;
  assign y1506 = ~n2014 ;
  assign y1507 = n2017 ;
  assign y1508 = ~n2018 ;
  assign y1509 = n2027 ;
  assign y1510 = n2012 ;
  assign y1511 = ~n2031 ;
  assign y1512 = n2032 ;
  assign y1513 = 1'b0 ;
  assign y1514 = n2034 ;
  assign y1515 = n2041 ;
  assign y1516 = ~n2044 ;
  assign y1517 = n2049 ;
  assign y1518 = n2050 ;
  assign y1519 = ~1'b0 ;
  assign y1520 = ~1'b0 ;
  assign y1521 = ~1'b0 ;
  assign y1522 = ~1'b0 ;
  assign y1523 = n2058 ;
  assign y1524 = ~1'b0 ;
  assign y1525 = n2059 ;
  assign y1526 = ~1'b0 ;
  assign y1527 = n423 ;
  assign y1528 = ~1'b0 ;
  assign y1529 = n2060 ;
  assign y1530 = n2062 ;
  assign y1531 = n1441 ;
  assign y1532 = ~1'b0 ;
  assign y1533 = n2063 ;
  assign y1534 = 1'b0 ;
  assign y1535 = n2065 ;
  assign y1536 = n2067 ;
  assign y1537 = ~1'b0 ;
  assign y1538 = ~n2072 ;
  assign y1539 = ~n1368 ;
  assign y1540 = n2075 ;
  assign y1541 = ~1'b0 ;
  assign y1542 = ~n2083 ;
  assign y1543 = n2087 ;
  assign y1544 = n2096 ;
  assign y1545 = ~n1593 ;
  assign y1546 = n2099 ;
  assign y1547 = ~n2100 ;
  assign y1548 = ~1'b0 ;
  assign y1549 = n2102 ;
  assign y1550 = n804 ;
  assign y1551 = ~n506 ;
  assign y1552 = n2103 ;
  assign y1553 = ~1'b0 ;
  assign y1554 = n2104 ;
  assign y1555 = n2106 ;
  assign y1556 = n2108 ;
  assign y1557 = ~1'b0 ;
  assign y1558 = ~1'b0 ;
  assign y1559 = 1'b0 ;
  assign y1560 = ~n472 ;
  assign y1561 = ~1'b0 ;
  assign y1562 = n2109 ;
  assign y1563 = n2112 ;
  assign y1564 = ~n2114 ;
  assign y1565 = n2119 ;
  assign y1566 = ~1'b0 ;
  assign y1567 = ~1'b0 ;
  assign y1568 = n2122 ;
  assign y1569 = ~n2124 ;
  assign y1570 = n2128 ;
  assign y1571 = ~1'b0 ;
  assign y1572 = 1'b0 ;
  assign y1573 = n2130 ;
  assign y1574 = 1'b0 ;
  assign y1575 = ~n2131 ;
  assign y1576 = ~n2133 ;
  assign y1577 = n2134 ;
  assign y1578 = ~n2135 ;
  assign y1579 = 1'b0 ;
  assign y1580 = ~n2065 ;
  assign y1581 = ~1'b0 ;
  assign y1582 = n2136 ;
  assign y1583 = n1048 ;
  assign y1584 = ~n2140 ;
  assign y1585 = ~1'b0 ;
  assign y1586 = ~n2141 ;
  assign y1587 = n2142 ;
  assign y1588 = ~n246 ;
  assign y1589 = 1'b0 ;
  assign y1590 = ~n2145 ;
  assign y1591 = ~1'b0 ;
  assign y1592 = ~n2148 ;
  assign y1593 = n2150 ;
  assign y1594 = n2152 ;
  assign y1595 = ~n2155 ;
  assign y1596 = n477 ;
  assign y1597 = 1'b0 ;
  assign y1598 = n2159 ;
  assign y1599 = ~1'b0 ;
  assign y1600 = ~1'b0 ;
  assign y1601 = n2160 ;
  assign y1602 = ~n2162 ;
  assign y1603 = ~n2164 ;
  assign y1604 = n2167 ;
  assign y1605 = n2170 ;
  assign y1606 = n2172 ;
  assign y1607 = ~n2175 ;
  assign y1608 = ~1'b0 ;
  assign y1609 = n294 ;
  assign y1610 = ~n2176 ;
  assign y1611 = ~n2178 ;
  assign y1612 = ~1'b0 ;
  assign y1613 = ~1'b0 ;
  assign y1614 = ~1'b0 ;
  assign y1615 = ~n2180 ;
  assign y1616 = ~1'b0 ;
  assign y1617 = n2181 ;
  assign y1618 = ~1'b0 ;
  assign y1619 = n2183 ;
  assign y1620 = n2186 ;
  assign y1621 = ~n2188 ;
  assign y1622 = n2199 ;
  assign y1623 = n2200 ;
  assign y1624 = ~1'b0 ;
  assign y1625 = ~1'b0 ;
  assign y1626 = n2203 ;
  assign y1627 = n2204 ;
  assign y1628 = ~1'b0 ;
  assign y1629 = ~1'b0 ;
  assign y1630 = ~n2097 ;
  assign y1631 = ~1'b0 ;
  assign y1632 = ~n2209 ;
  assign y1633 = n2210 ;
  assign y1634 = n2216 ;
  assign y1635 = ~1'b0 ;
  assign y1636 = n2218 ;
  assign y1637 = ~1'b0 ;
  assign y1638 = n2219 ;
  assign y1639 = 1'b0 ;
  assign y1640 = 1'b0 ;
  assign y1641 = n2220 ;
  assign y1642 = ~1'b0 ;
  assign y1643 = ~1'b0 ;
  assign y1644 = n2222 ;
  assign y1645 = 1'b0 ;
  assign y1646 = n2227 ;
  assign y1647 = n2228 ;
  assign y1648 = ~1'b0 ;
  assign y1649 = ~1'b0 ;
  assign y1650 = ~1'b0 ;
  assign y1651 = n2231 ;
  assign y1652 = n2235 ;
  assign y1653 = n2238 ;
  assign y1654 = ~1'b0 ;
  assign y1655 = n2239 ;
  assign y1656 = ~n2240 ;
  assign y1657 = ~1'b0 ;
  assign y1658 = ~n2242 ;
  assign y1659 = ~n2243 ;
  assign y1660 = ~1'b0 ;
  assign y1661 = ~n2244 ;
  assign y1662 = ~n2245 ;
  assign y1663 = n2248 ;
  assign y1664 = ~1'b0 ;
  assign y1665 = ~1'b0 ;
  assign y1666 = ~1'b0 ;
  assign y1667 = ~1'b0 ;
  assign y1668 = ~1'b0 ;
  assign y1669 = ~n2251 ;
  assign y1670 = n2252 ;
  assign y1671 = ~n2257 ;
  assign y1672 = n2261 ;
  assign y1673 = ~1'b0 ;
  assign y1674 = ~n439 ;
  assign y1675 = 1'b0 ;
  assign y1676 = n2101 ;
  assign y1677 = n2266 ;
  assign y1678 = ~n2267 ;
  assign y1679 = ~1'b0 ;
  assign y1680 = ~1'b0 ;
  assign y1681 = ~1'b0 ;
  assign y1682 = ~n2270 ;
  assign y1683 = ~n2277 ;
  assign y1684 = n2279 ;
  assign y1685 = n128 ;
  assign y1686 = ~1'b0 ;
  assign y1687 = n2280 ;
  assign y1688 = ~1'b0 ;
  assign y1689 = n2281 ;
  assign y1690 = ~1'b0 ;
  assign y1691 = ~1'b0 ;
  assign y1692 = ~n2282 ;
  assign y1693 = n2283 ;
  assign y1694 = 1'b0 ;
  assign y1695 = ~n2288 ;
  assign y1696 = ~n2301 ;
  assign y1697 = n2302 ;
  assign y1698 = n2303 ;
  assign y1699 = ~1'b0 ;
  assign y1700 = ~n2304 ;
  assign y1701 = ~n2307 ;
  assign y1702 = ~1'b0 ;
  assign y1703 = n2308 ;
  assign y1704 = n630 ;
  assign y1705 = ~1'b0 ;
  assign y1706 = ~1'b0 ;
  assign y1707 = ~1'b0 ;
  assign y1708 = ~1'b0 ;
  assign y1709 = n2310 ;
  assign y1710 = ~1'b0 ;
  assign y1711 = ~1'b0 ;
  assign y1712 = ~n2311 ;
  assign y1713 = ~n2313 ;
  assign y1714 = ~1'b0 ;
  assign y1715 = ~1'b0 ;
  assign y1716 = ~n122 ;
  assign y1717 = ~1'b0 ;
  assign y1718 = n2317 ;
  assign y1719 = ~1'b0 ;
  assign y1720 = n2322 ;
  assign y1721 = ~1'b0 ;
  assign y1722 = n1358 ;
  assign y1723 = ~1'b0 ;
  assign y1724 = ~n2324 ;
  assign y1725 = n2254 ;
  assign y1726 = ~1'b0 ;
  assign y1727 = ~1'b0 ;
  assign y1728 = ~1'b0 ;
  assign y1729 = ~1'b0 ;
  assign y1730 = ~n461 ;
  assign y1731 = ~n827 ;
  assign y1732 = n2330 ;
  assign y1733 = n2331 ;
  assign y1734 = n2332 ;
  assign y1735 = ~1'b0 ;
  assign y1736 = n2333 ;
  assign y1737 = n1968 ;
  assign y1738 = ~n2335 ;
  assign y1739 = ~1'b0 ;
  assign y1740 = n2342 ;
  assign y1741 = ~1'b0 ;
  assign y1742 = n2344 ;
  assign y1743 = ~n2348 ;
  assign y1744 = ~n2349 ;
  assign y1745 = n2351 ;
  assign y1746 = n2353 ;
  assign y1747 = ~n2356 ;
  assign y1748 = ~1'b0 ;
  assign y1749 = n2360 ;
  assign y1750 = n960 ;
  assign y1751 = ~1'b0 ;
  assign y1752 = n2361 ;
  assign y1753 = ~1'b0 ;
  assign y1754 = ~1'b0 ;
  assign y1755 = ~n2366 ;
  assign y1756 = n2209 ;
  assign y1757 = ~n2369 ;
  assign y1758 = n2370 ;
  assign y1759 = n2373 ;
  assign y1760 = ~n2375 ;
  assign y1761 = ~1'b0 ;
  assign y1762 = n2377 ;
  assign y1763 = ~n2378 ;
  assign y1764 = ~1'b0 ;
  assign y1765 = n2380 ;
  assign y1766 = n553 ;
  assign y1767 = ~n2382 ;
  assign y1768 = ~1'b0 ;
  assign y1769 = n2384 ;
  assign y1770 = ~1'b0 ;
  assign y1771 = ~n2386 ;
  assign y1772 = ~1'b0 ;
  assign y1773 = ~n1441 ;
  assign y1774 = n2394 ;
  assign y1775 = ~n520 ;
  assign y1776 = ~1'b0 ;
  assign y1777 = n52 ;
  assign y1778 = ~1'b0 ;
  assign y1779 = ~1'b0 ;
  assign y1780 = ~n2395 ;
  assign y1781 = n2399 ;
  assign y1782 = ~n2401 ;
  assign y1783 = n2403 ;
  assign y1784 = ~1'b0 ;
  assign y1785 = n1848 ;
  assign y1786 = n2404 ;
  assign y1787 = ~n2410 ;
  assign y1788 = ~1'b0 ;
  assign y1789 = ~1'b0 ;
  assign y1790 = ~1'b0 ;
  assign y1791 = ~1'b0 ;
  assign y1792 = 1'b0 ;
  assign y1793 = ~n2412 ;
  assign y1794 = ~1'b0 ;
  assign y1795 = ~1'b0 ;
  assign y1796 = n2415 ;
  assign y1797 = n2418 ;
  assign y1798 = n2419 ;
  assign y1799 = 1'b0 ;
  assign y1800 = ~1'b0 ;
  assign y1801 = ~1'b0 ;
  assign y1802 = n2424 ;
  assign y1803 = ~n879 ;
  assign y1804 = ~1'b0 ;
  assign y1805 = ~1'b0 ;
  assign y1806 = n2425 ;
  assign y1807 = ~1'b0 ;
  assign y1808 = n2430 ;
  assign y1809 = 1'b0 ;
  assign y1810 = ~1'b0 ;
  assign y1811 = n2431 ;
  assign y1812 = ~1'b0 ;
  assign y1813 = ~1'b0 ;
  assign y1814 = n2432 ;
  assign y1815 = ~1'b0 ;
  assign y1816 = n2433 ;
  assign y1817 = n2086 ;
  assign y1818 = 1'b0 ;
  assign y1819 = ~1'b0 ;
  assign y1820 = ~1'b0 ;
  assign y1821 = ~n2435 ;
  assign y1822 = ~n2436 ;
  assign y1823 = ~n2437 ;
  assign y1824 = ~1'b0 ;
  assign y1825 = n823 ;
  assign y1826 = ~1'b0 ;
  assign y1827 = n2438 ;
  assign y1828 = ~n2440 ;
  assign y1829 = ~n2443 ;
  assign y1830 = n2446 ;
  assign y1831 = 1'b0 ;
  assign y1832 = n2448 ;
  assign y1833 = n2452 ;
  assign y1834 = n1227 ;
  assign y1835 = ~n2454 ;
  assign y1836 = ~n2455 ;
  assign y1837 = ~n2460 ;
  assign y1838 = n2064 ;
  assign y1839 = ~n2465 ;
  assign y1840 = ~n2472 ;
  assign y1841 = ~n2477 ;
  assign y1842 = n2481 ;
  assign y1843 = ~n2483 ;
  assign y1844 = ~1'b0 ;
  assign y1845 = n2484 ;
  assign y1846 = ~n2485 ;
  assign y1847 = ~1'b0 ;
  assign y1848 = ~n2486 ;
  assign y1849 = ~1'b0 ;
  assign y1850 = n2487 ;
  assign y1851 = n2493 ;
  assign y1852 = x0 ;
  assign y1853 = ~1'b0 ;
  assign y1854 = ~n2494 ;
  assign y1855 = ~1'b0 ;
  assign y1856 = ~1'b0 ;
  assign y1857 = 1'b0 ;
  assign y1858 = ~n2495 ;
  assign y1859 = ~1'b0 ;
  assign y1860 = ~n2496 ;
  assign y1861 = n2499 ;
  assign y1862 = ~n2501 ;
  assign y1863 = ~n2502 ;
  assign y1864 = n2506 ;
  assign y1865 = n2508 ;
  assign y1866 = n2509 ;
  assign y1867 = n2510 ;
  assign y1868 = n1447 ;
  assign y1869 = n2513 ;
  assign y1870 = ~1'b0 ;
  assign y1871 = ~n2514 ;
  assign y1872 = n2515 ;
  assign y1873 = ~1'b0 ;
  assign y1874 = ~1'b0 ;
  assign y1875 = ~n2517 ;
  assign y1876 = ~1'b0 ;
  assign y1877 = n2523 ;
  assign y1878 = n2526 ;
  assign y1879 = ~1'b0 ;
  assign y1880 = ~n2529 ;
  assign y1881 = ~1'b0 ;
  assign y1882 = n2533 ;
  assign y1883 = 1'b0 ;
  assign y1884 = n2535 ;
  assign y1885 = ~1'b0 ;
  assign y1886 = n2537 ;
  assign y1887 = ~1'b0 ;
  assign y1888 = ~n2541 ;
  assign y1889 = ~1'b0 ;
  assign y1890 = ~1'b0 ;
  assign y1891 = ~1'b0 ;
  assign y1892 = ~1'b0 ;
  assign y1893 = ~n2543 ;
  assign y1894 = n2546 ;
  assign y1895 = ~1'b0 ;
  assign y1896 = n2549 ;
  assign y1897 = n2550 ;
  assign y1898 = n2551 ;
  assign y1899 = ~n2553 ;
  assign y1900 = ~n2560 ;
  assign y1901 = n2565 ;
  assign y1902 = n2566 ;
  assign y1903 = ~n2568 ;
  assign y1904 = n2569 ;
  assign y1905 = 1'b0 ;
  assign y1906 = ~n2572 ;
  assign y1907 = ~1'b0 ;
  assign y1908 = ~n2575 ;
  assign y1909 = ~n2576 ;
  assign y1910 = 1'b0 ;
  assign y1911 = 1'b0 ;
  assign y1912 = n2578 ;
  assign y1913 = ~n2581 ;
  assign y1914 = n2584 ;
  assign y1915 = ~n2260 ;
  assign y1916 = ~n2585 ;
  assign y1917 = ~1'b0 ;
  assign y1918 = ~1'b0 ;
  assign y1919 = n2587 ;
  assign y1920 = n1007 ;
  assign y1921 = ~1'b0 ;
  assign y1922 = ~n2594 ;
  assign y1923 = ~1'b0 ;
  assign y1924 = n2595 ;
  assign y1925 = ~1'b0 ;
  assign y1926 = ~1'b0 ;
  assign y1927 = ~n2599 ;
  assign y1928 = 1'b0 ;
  assign y1929 = ~1'b0 ;
  assign y1930 = ~n2601 ;
  assign y1931 = ~1'b0 ;
  assign y1932 = n2606 ;
  assign y1933 = ~n2608 ;
  assign y1934 = n2611 ;
  assign y1935 = ~n2612 ;
  assign y1936 = ~n2617 ;
  assign y1937 = n2618 ;
  assign y1938 = ~1'b0 ;
  assign y1939 = ~1'b0 ;
  assign y1940 = ~1'b0 ;
  assign y1941 = ~1'b0 ;
  assign y1942 = n2623 ;
  assign y1943 = n1096 ;
  assign y1944 = ~1'b0 ;
  assign y1945 = n2185 ;
  assign y1946 = ~n2497 ;
  assign y1947 = n2627 ;
  assign y1948 = ~1'b0 ;
  assign y1949 = ~1'b0 ;
  assign y1950 = ~1'b0 ;
  assign y1951 = ~n2630 ;
  assign y1952 = ~n2631 ;
  assign y1953 = ~1'b0 ;
  assign y1954 = ~1'b0 ;
  assign y1955 = ~1'b0 ;
  assign y1956 = ~1'b0 ;
  assign y1957 = n2637 ;
  assign y1958 = ~n2639 ;
  assign y1959 = n2647 ;
  assign y1960 = n290 ;
  assign y1961 = ~1'b0 ;
  assign y1962 = n799 ;
  assign y1963 = n2652 ;
  assign y1964 = n1810 ;
  assign y1965 = ~1'b0 ;
  assign y1966 = ~1'b0 ;
  assign y1967 = n2655 ;
  assign y1968 = n2658 ;
  assign y1969 = ~1'b0 ;
  assign y1970 = ~1'b0 ;
  assign y1971 = ~1'b0 ;
  assign y1972 = ~n626 ;
  assign y1973 = ~1'b0 ;
  assign y1974 = n2659 ;
  assign y1975 = ~n2660 ;
  assign y1976 = n685 ;
  assign y1977 = ~1'b0 ;
  assign y1978 = n2662 ;
  assign y1979 = ~n2665 ;
  assign y1980 = ~1'b0 ;
  assign y1981 = n2674 ;
  assign y1982 = ~n2676 ;
  assign y1983 = n2677 ;
  assign y1984 = ~1'b0 ;
  assign y1985 = ~1'b0 ;
  assign y1986 = n2682 ;
  assign y1987 = n2686 ;
  assign y1988 = ~n1406 ;
  assign y1989 = n2689 ;
  assign y1990 = 1'b0 ;
  assign y1991 = ~1'b0 ;
  assign y1992 = ~1'b0 ;
  assign y1993 = ~1'b0 ;
  assign y1994 = n2690 ;
  assign y1995 = ~1'b0 ;
  assign y1996 = n2695 ;
  assign y1997 = ~1'b0 ;
  assign y1998 = ~n149 ;
  assign y1999 = n2699 ;
  assign y2000 = ~1'b0 ;
  assign y2001 = ~n2702 ;
  assign y2002 = n2705 ;
  assign y2003 = ~1'b0 ;
  assign y2004 = ~1'b0 ;
  assign y2005 = 1'b0 ;
  assign y2006 = ~1'b0 ;
  assign y2007 = ~n2591 ;
  assign y2008 = ~1'b0 ;
  assign y2009 = n2607 ;
  assign y2010 = n2707 ;
  assign y2011 = ~1'b0 ;
  assign y2012 = n2074 ;
  assign y2013 = ~n2709 ;
  assign y2014 = n2712 ;
  assign y2015 = 1'b0 ;
  assign y2016 = ~1'b0 ;
  assign y2017 = n2721 ;
  assign y2018 = n2307 ;
  assign y2019 = ~n2722 ;
  assign y2020 = ~n2723 ;
  assign y2021 = ~n2726 ;
  assign y2022 = ~1'b0 ;
  assign y2023 = n2728 ;
  assign y2024 = ~n2730 ;
  assign y2025 = ~1'b0 ;
  assign y2026 = ~n2731 ;
  assign y2027 = 1'b0 ;
  assign y2028 = ~1'b0 ;
  assign y2029 = n2744 ;
  assign y2030 = ~1'b0 ;
  assign y2031 = ~1'b0 ;
  assign y2032 = n2745 ;
  assign y2033 = n2747 ;
  assign y2034 = 1'b0 ;
  assign y2035 = n2753 ;
  assign y2036 = ~1'b0 ;
  assign y2037 = ~n2760 ;
  assign y2038 = ~n2761 ;
  assign y2039 = ~n2764 ;
  assign y2040 = n2769 ;
  assign y2041 = n395 ;
  assign y2042 = n2770 ;
  assign y2043 = ~1'b0 ;
  assign y2044 = ~n2771 ;
  assign y2045 = n2773 ;
  assign y2046 = ~n2774 ;
  assign y2047 = ~n1019 ;
  assign y2048 = n2779 ;
  assign y2049 = ~n2784 ;
  assign y2050 = ~n2785 ;
  assign y2051 = ~n2786 ;
  assign y2052 = ~n2577 ;
  assign y2053 = ~n2787 ;
  assign y2054 = ~n2788 ;
  assign y2055 = ~n1341 ;
  assign y2056 = ~1'b0 ;
  assign y2057 = ~n2789 ;
  assign y2058 = ~1'b0 ;
  assign y2059 = ~1'b0 ;
  assign y2060 = 1'b0 ;
  assign y2061 = n2796 ;
  assign y2062 = ~1'b0 ;
  assign y2063 = ~1'b0 ;
  assign y2064 = ~1'b0 ;
  assign y2065 = n1931 ;
  assign y2066 = n2797 ;
  assign y2067 = n2799 ;
  assign y2068 = n2802 ;
  assign y2069 = ~1'b0 ;
  assign y2070 = ~1'b0 ;
  assign y2071 = n2809 ;
  assign y2072 = 1'b0 ;
  assign y2073 = n356 ;
  assign y2074 = ~1'b0 ;
  assign y2075 = ~n2810 ;
  assign y2076 = ~1'b0 ;
  assign y2077 = n2811 ;
  assign y2078 = n268 ;
  assign y2079 = ~n2814 ;
  assign y2080 = ~1'b0 ;
  assign y2081 = ~1'b0 ;
  assign y2082 = n1051 ;
  assign y2083 = ~n2817 ;
  assign y2084 = ~1'b0 ;
  assign y2085 = ~1'b0 ;
  assign y2086 = ~1'b0 ;
  assign y2087 = ~1'b0 ;
  assign y2088 = ~1'b0 ;
  assign y2089 = ~1'b0 ;
  assign y2090 = n2818 ;
  assign y2091 = ~n2819 ;
  assign y2092 = n2822 ;
  assign y2093 = ~n2829 ;
  assign y2094 = n2830 ;
  assign y2095 = n144 ;
  assign y2096 = ~1'b0 ;
  assign y2097 = n2831 ;
  assign y2098 = ~n2834 ;
  assign y2099 = ~1'b0 ;
  assign y2100 = ~1'b0 ;
  assign y2101 = n366 ;
  assign y2102 = n2836 ;
  assign y2103 = n2837 ;
  assign y2104 = ~n1258 ;
  assign y2105 = n2840 ;
  assign y2106 = n1430 ;
  assign y2107 = n2841 ;
  assign y2108 = ~n2110 ;
  assign y2109 = ~n2842 ;
  assign y2110 = ~1'b0 ;
  assign y2111 = ~n2844 ;
  assign y2112 = ~1'b0 ;
  assign y2113 = ~1'b0 ;
  assign y2114 = ~1'b0 ;
  assign y2115 = ~1'b0 ;
  assign y2116 = ~n2847 ;
  assign y2117 = ~1'b0 ;
  assign y2118 = ~n2848 ;
  assign y2119 = n2850 ;
  assign y2120 = 1'b0 ;
  assign y2121 = ~n2853 ;
  assign y2122 = ~n2531 ;
  assign y2123 = ~n2855 ;
  assign y2124 = ~1'b0 ;
  assign y2125 = ~1'b0 ;
  assign y2126 = ~n2858 ;
  assign y2127 = ~n2859 ;
  assign y2128 = ~n2860 ;
  assign y2129 = n2861 ;
  assign y2130 = ~1'b0 ;
  assign y2131 = n2862 ;
  assign y2132 = n1431 ;
  assign y2133 = ~n2864 ;
  assign y2134 = ~n246 ;
  assign y2135 = ~n2866 ;
  assign y2136 = ~n2867 ;
  assign y2137 = ~1'b0 ;
  assign y2138 = ~n2869 ;
  assign y2139 = ~1'b0 ;
  assign y2140 = ~1'b0 ;
  assign y2141 = n2870 ;
  assign y2142 = ~1'b0 ;
  assign y2143 = ~1'b0 ;
  assign y2144 = ~1'b0 ;
  assign y2145 = ~1'b0 ;
  assign y2146 = n2872 ;
  assign y2147 = n2873 ;
  assign y2148 = n2880 ;
  assign y2149 = n1920 ;
  assign y2150 = ~1'b0 ;
  assign y2151 = ~n2891 ;
  assign y2152 = ~1'b0 ;
  assign y2153 = n2893 ;
  assign y2154 = ~n2894 ;
  assign y2155 = ~1'b0 ;
  assign y2156 = ~1'b0 ;
  assign y2157 = ~n2898 ;
  assign y2158 = n2899 ;
  assign y2159 = n2348 ;
  assign y2160 = ~1'b0 ;
  assign y2161 = n2900 ;
  assign y2162 = ~n2902 ;
  assign y2163 = ~n2903 ;
  assign y2164 = ~n2848 ;
  assign y2165 = ~1'b0 ;
  assign y2166 = n2906 ;
  assign y2167 = ~n2907 ;
  assign y2168 = ~n2908 ;
  assign y2169 = ~1'b0 ;
  assign y2170 = ~1'b0 ;
  assign y2171 = ~1'b0 ;
  assign y2172 = ~1'b0 ;
  assign y2173 = ~1'b0 ;
  assign y2174 = n2910 ;
  assign y2175 = ~n2911 ;
  assign y2176 = n2913 ;
  assign y2177 = ~1'b0 ;
  assign y2178 = ~n2914 ;
  assign y2179 = 1'b0 ;
  assign y2180 = n2915 ;
  assign y2181 = ~1'b0 ;
  assign y2182 = ~n2916 ;
  assign y2183 = 1'b0 ;
  assign y2184 = ~n2917 ;
  assign y2185 = ~n2923 ;
  assign y2186 = ~n2924 ;
  assign y2187 = 1'b0 ;
  assign y2188 = ~1'b0 ;
  assign y2189 = n2929 ;
  assign y2190 = ~1'b0 ;
  assign y2191 = ~1'b0 ;
  assign y2192 = n302 ;
  assign y2193 = ~1'b0 ;
  assign y2194 = ~1'b0 ;
  assign y2195 = ~n2933 ;
  assign y2196 = n2936 ;
  assign y2197 = x11 ;
  assign y2198 = ~1'b0 ;
  assign y2199 = n2938 ;
  assign y2200 = ~n2943 ;
  assign y2201 = ~n2945 ;
  assign y2202 = ~1'b0 ;
  assign y2203 = ~n2946 ;
  assign y2204 = ~1'b0 ;
  assign y2205 = ~n2947 ;
  assign y2206 = n2953 ;
  assign y2207 = ~1'b0 ;
  assign y2208 = ~n310 ;
  assign y2209 = ~n2959 ;
  assign y2210 = ~1'b0 ;
  assign y2211 = ~n2963 ;
  assign y2212 = 1'b0 ;
  assign y2213 = n2967 ;
  assign y2214 = n2968 ;
  assign y2215 = n2969 ;
  assign y2216 = n2971 ;
  assign y2217 = ~1'b0 ;
  assign y2218 = ~1'b0 ;
  assign y2219 = ~1'b0 ;
  assign y2220 = ~n2973 ;
  assign y2221 = n2975 ;
  assign y2222 = ~1'b0 ;
  assign y2223 = ~n2978 ;
  assign y2224 = 1'b0 ;
  assign y2225 = ~1'b0 ;
  assign y2226 = ~1'b0 ;
  assign y2227 = ~1'b0 ;
  assign y2228 = ~n2979 ;
  assign y2229 = n2982 ;
  assign y2230 = ~n2020 ;
  assign y2231 = ~n724 ;
  assign y2232 = ~1'b0 ;
  assign y2233 = ~n158 ;
  assign y2234 = ~1'b0 ;
  assign y2235 = n1300 ;
  assign y2236 = n2986 ;
  assign y2237 = ~n2988 ;
  assign y2238 = n2990 ;
  assign y2239 = ~n2991 ;
  assign y2240 = ~n2999 ;
  assign y2241 = ~1'b0 ;
  assign y2242 = ~n3001 ;
  assign y2243 = ~1'b0 ;
  assign y2244 = ~1'b0 ;
  assign y2245 = n489 ;
  assign y2246 = ~1'b0 ;
  assign y2247 = n1152 ;
  assign y2248 = ~1'b0 ;
  assign y2249 = n3002 ;
  assign y2250 = ~1'b0 ;
  assign y2251 = ~1'b0 ;
  assign y2252 = n1425 ;
  assign y2253 = ~n3007 ;
  assign y2254 = n3009 ;
  assign y2255 = ~n3010 ;
  assign y2256 = n3014 ;
  assign y2257 = n512 ;
  assign y2258 = n1851 ;
  assign y2259 = n3022 ;
  assign y2260 = n3023 ;
  assign y2261 = ~1'b0 ;
  assign y2262 = ~n3024 ;
  assign y2263 = x11 ;
  assign y2264 = ~n907 ;
  assign y2265 = ~n3027 ;
  assign y2266 = ~1'b0 ;
  assign y2267 = n3028 ;
  assign y2268 = ~1'b0 ;
  assign y2269 = ~1'b0 ;
  assign y2270 = ~n1591 ;
  assign y2271 = n1918 ;
  assign y2272 = ~n3030 ;
  assign y2273 = n3037 ;
  assign y2274 = n3040 ;
  assign y2275 = n3042 ;
  assign y2276 = n3044 ;
  assign y2277 = ~n754 ;
  assign y2278 = ~1'b0 ;
  assign y2279 = n3049 ;
  assign y2280 = n3050 ;
  assign y2281 = ~1'b0 ;
  assign y2282 = ~n3051 ;
  assign y2283 = 1'b0 ;
  assign y2284 = ~n3053 ;
  assign y2285 = n3054 ;
  assign y2286 = ~n3056 ;
  assign y2287 = n3057 ;
  assign y2288 = ~1'b0 ;
  assign y2289 = n3061 ;
  assign y2290 = ~1'b0 ;
  assign y2291 = ~n3064 ;
  assign y2292 = ~n3067 ;
  assign y2293 = ~n3069 ;
  assign y2294 = ~n820 ;
  assign y2295 = n3075 ;
  assign y2296 = n3077 ;
  assign y2297 = ~1'b0 ;
  assign y2298 = n3078 ;
  assign y2299 = ~1'b0 ;
  assign y2300 = ~n3080 ;
  assign y2301 = ~n3083 ;
  assign y2302 = ~n1471 ;
  assign y2303 = ~1'b0 ;
  assign y2304 = ~n3085 ;
  assign y2305 = n3089 ;
  assign y2306 = ~n1688 ;
  assign y2307 = ~1'b0 ;
  assign y2308 = ~1'b0 ;
  assign y2309 = ~n3091 ;
  assign y2310 = n3093 ;
  assign y2311 = ~n3098 ;
  assign y2312 = ~n2446 ;
  assign y2313 = n3099 ;
  assign y2314 = ~n3103 ;
  assign y2315 = ~n3104 ;
  assign y2316 = n3106 ;
  assign y2317 = ~n1802 ;
  assign y2318 = n1474 ;
  assign y2319 = n3107 ;
  assign y2320 = n3114 ;
  assign y2321 = ~n3115 ;
  assign y2322 = ~n3116 ;
  assign y2323 = ~1'b0 ;
  assign y2324 = ~1'b0 ;
  assign y2325 = ~1'b0 ;
  assign y2326 = n581 ;
  assign y2327 = ~1'b0 ;
  assign y2328 = n995 ;
  assign y2329 = ~1'b0 ;
  assign y2330 = n3120 ;
  assign y2331 = ~1'b0 ;
  assign y2332 = ~n3122 ;
  assign y2333 = n3123 ;
  assign y2334 = n3126 ;
  assign y2335 = ~n3127 ;
  assign y2336 = ~n3131 ;
  assign y2337 = ~1'b0 ;
  assign y2338 = ~1'b0 ;
  assign y2339 = n3135 ;
  assign y2340 = n3137 ;
  assign y2341 = ~1'b0 ;
  assign y2342 = ~1'b0 ;
  assign y2343 = n3146 ;
  assign y2344 = n3152 ;
  assign y2345 = ~1'b0 ;
  assign y2346 = n3154 ;
  assign y2347 = ~n3156 ;
  assign y2348 = 1'b0 ;
  assign y2349 = ~1'b0 ;
  assign y2350 = ~n3158 ;
  assign y2351 = n3160 ;
  assign y2352 = n3162 ;
  assign y2353 = ~1'b0 ;
  assign y2354 = ~1'b0 ;
  assign y2355 = ~1'b0 ;
  assign y2356 = ~1'b0 ;
  assign y2357 = n3166 ;
  assign y2358 = n3167 ;
  assign y2359 = n3173 ;
  assign y2360 = n3175 ;
  assign y2361 = ~n1370 ;
  assign y2362 = ~1'b0 ;
  assign y2363 = ~n3177 ;
  assign y2364 = ~n3179 ;
  assign y2365 = ~n3180 ;
  assign y2366 = n3185 ;
  assign y2367 = ~n3186 ;
  assign y2368 = n3191 ;
  assign y2369 = n3192 ;
  assign y2370 = ~n3193 ;
  assign y2371 = n3197 ;
  assign y2372 = ~n3199 ;
  assign y2373 = ~1'b0 ;
  assign y2374 = ~1'b0 ;
  assign y2375 = ~n3202 ;
  assign y2376 = ~1'b0 ;
  assign y2377 = ~1'b0 ;
  assign y2378 = ~1'b0 ;
  assign y2379 = ~1'b0 ;
  assign y2380 = ~1'b0 ;
  assign y2381 = ~n3203 ;
  assign y2382 = ~1'b0 ;
  assign y2383 = ~n3207 ;
  assign y2384 = n495 ;
  assign y2385 = ~1'b0 ;
  assign y2386 = ~n3211 ;
  assign y2387 = ~1'b0 ;
  assign y2388 = n3212 ;
  assign y2389 = n3214 ;
  assign y2390 = ~n3216 ;
  assign y2391 = n3217 ;
  assign y2392 = n3218 ;
  assign y2393 = ~1'b0 ;
  assign y2394 = n3219 ;
  assign y2395 = ~n3220 ;
  assign y2396 = ~1'b0 ;
  assign y2397 = 1'b0 ;
  assign y2398 = n3221 ;
  assign y2399 = ~1'b0 ;
  assign y2400 = ~n3225 ;
  assign y2401 = ~1'b0 ;
  assign y2402 = n3226 ;
  assign y2403 = ~1'b0 ;
  assign y2404 = ~n3227 ;
  assign y2405 = ~1'b0 ;
  assign y2406 = ~n3228 ;
  assign y2407 = ~1'b0 ;
  assign y2408 = ~n1584 ;
  assign y2409 = ~1'b0 ;
  assign y2410 = ~1'b0 ;
  assign y2411 = ~n3229 ;
  assign y2412 = 1'b0 ;
  assign y2413 = ~n3231 ;
  assign y2414 = ~1'b0 ;
  assign y2415 = ~1'b0 ;
  assign y2416 = ~n3233 ;
  assign y2417 = n3238 ;
  assign y2418 = n3239 ;
  assign y2419 = ~1'b0 ;
  assign y2420 = ~1'b0 ;
  assign y2421 = ~n3240 ;
  assign y2422 = n3242 ;
  assign y2423 = ~1'b0 ;
  assign y2424 = n3243 ;
  assign y2425 = n3244 ;
  assign y2426 = n3245 ;
  assign y2427 = ~1'b0 ;
  assign y2428 = ~1'b0 ;
  assign y2429 = n3246 ;
  assign y2430 = ~1'b0 ;
  assign y2431 = ~1'b0 ;
  assign y2432 = ~n3248 ;
  assign y2433 = ~1'b0 ;
  assign y2434 = n3254 ;
  assign y2435 = n3255 ;
  assign y2436 = n3265 ;
  assign y2437 = n3266 ;
  assign y2438 = ~1'b0 ;
  assign y2439 = ~1'b0 ;
  assign y2440 = ~1'b0 ;
  assign y2441 = ~n986 ;
  assign y2442 = ~1'b0 ;
  assign y2443 = ~n1310 ;
  assign y2444 = n3267 ;
  assign y2445 = ~1'b0 ;
  assign y2446 = ~1'b0 ;
  assign y2447 = n101 ;
  assign y2448 = ~n3268 ;
  assign y2449 = ~1'b0 ;
  assign y2450 = ~1'b0 ;
  assign y2451 = n3269 ;
  assign y2452 = ~n3274 ;
  assign y2453 = ~n3277 ;
  assign y2454 = n3278 ;
  assign y2455 = ~n3280 ;
  assign y2456 = ~1'b0 ;
  assign y2457 = 1'b0 ;
  assign y2458 = ~1'b0 ;
  assign y2459 = n3282 ;
  assign y2460 = ~n3284 ;
  assign y2461 = n3285 ;
  assign y2462 = ~n3286 ;
  assign y2463 = ~n3287 ;
  assign y2464 = ~1'b0 ;
  assign y2465 = ~n3289 ;
  assign y2466 = n3295 ;
  assign y2467 = n3299 ;
  assign y2468 = ~n3303 ;
  assign y2469 = n3304 ;
  assign y2470 = ~1'b0 ;
  assign y2471 = 1'b0 ;
  assign y2472 = ~n1396 ;
  assign y2473 = n3305 ;
  assign y2474 = n3306 ;
  assign y2475 = n3307 ;
  assign y2476 = ~1'b0 ;
  assign y2477 = n154 ;
  assign y2478 = ~1'b0 ;
  assign y2479 = ~1'b0 ;
  assign y2480 = ~n3309 ;
  assign y2481 = ~n3314 ;
  assign y2482 = n3320 ;
  assign y2483 = n3321 ;
  assign y2484 = ~n2882 ;
  assign y2485 = n3325 ;
  assign y2486 = n3327 ;
  assign y2487 = n3329 ;
  assign y2488 = ~n3334 ;
  assign y2489 = n3335 ;
  assign y2490 = ~1'b0 ;
  assign y2491 = ~n3337 ;
  assign y2492 = n1693 ;
  assign y2493 = n3338 ;
  assign y2494 = ~n3341 ;
  assign y2495 = n3345 ;
  assign y2496 = 1'b0 ;
  assign y2497 = ~n3347 ;
  assign y2498 = n3348 ;
  assign y2499 = ~n520 ;
  assign y2500 = ~1'b0 ;
  assign y2501 = ~n2294 ;
  assign y2502 = ~1'b0 ;
  assign y2503 = n3353 ;
  assign y2504 = ~1'b0 ;
  assign y2505 = ~1'b0 ;
  assign y2506 = ~n3354 ;
  assign y2507 = ~n3355 ;
  assign y2508 = n3356 ;
  assign y2509 = ~n3359 ;
  assign y2510 = n3361 ;
  assign y2511 = n3363 ;
  assign y2512 = n3368 ;
  assign y2513 = ~1'b0 ;
  assign y2514 = ~n3371 ;
  assign y2515 = ~1'b0 ;
  assign y2516 = n3374 ;
  assign y2517 = 1'b0 ;
  assign y2518 = n3377 ;
  assign y2519 = ~1'b0 ;
  assign y2520 = n187 ;
  assign y2521 = ~n3378 ;
  assign y2522 = ~1'b0 ;
  assign y2523 = ~n3380 ;
  assign y2524 = n3384 ;
  assign y2525 = ~1'b0 ;
  assign y2526 = ~1'b0 ;
  assign y2527 = 1'b0 ;
  assign y2528 = ~1'b0 ;
  assign y2529 = ~1'b0 ;
  assign y2530 = ~1'b0 ;
  assign y2531 = ~1'b0 ;
  assign y2532 = ~n3385 ;
  assign y2533 = ~n1089 ;
  assign y2534 = n3386 ;
  assign y2535 = ~1'b0 ;
  assign y2536 = n3389 ;
  assign y2537 = n3390 ;
  assign y2538 = ~n3392 ;
  assign y2539 = n3394 ;
  assign y2540 = ~n3395 ;
  assign y2541 = n3398 ;
  assign y2542 = ~1'b0 ;
  assign y2543 = ~1'b0 ;
  assign y2544 = n3399 ;
  assign y2545 = ~1'b0 ;
  assign y2546 = ~n3401 ;
  assign y2547 = n3402 ;
  assign y2548 = n3403 ;
  assign y2549 = ~n1822 ;
  assign y2550 = ~n3405 ;
  assign y2551 = 1'b0 ;
  assign y2552 = ~1'b0 ;
  assign y2553 = ~1'b0 ;
  assign y2554 = ~1'b0 ;
  assign y2555 = ~1'b0 ;
  assign y2556 = n3407 ;
  assign y2557 = ~1'b0 ;
  assign y2558 = ~n3411 ;
  assign y2559 = ~1'b0 ;
  assign y2560 = ~1'b0 ;
  assign y2561 = ~n3412 ;
  assign y2562 = 1'b0 ;
  assign y2563 = ~1'b0 ;
  assign y2564 = n3414 ;
  assign y2565 = n3415 ;
  assign y2566 = n3418 ;
  assign y2567 = ~1'b0 ;
  assign y2568 = ~n3422 ;
  assign y2569 = n3423 ;
  assign y2570 = n3426 ;
  assign y2571 = n3427 ;
  assign y2572 = ~1'b0 ;
  assign y2573 = n3428 ;
  assign y2574 = 1'b0 ;
  assign y2575 = ~1'b0 ;
  assign y2576 = n724 ;
  assign y2577 = ~n3429 ;
  assign y2578 = n3431 ;
  assign y2579 = ~n3435 ;
  assign y2580 = n3436 ;
  assign y2581 = n3437 ;
  assign y2582 = ~1'b0 ;
  assign y2583 = n3440 ;
  assign y2584 = ~n3444 ;
  assign y2585 = ~1'b0 ;
  assign y2586 = n1496 ;
  assign y2587 = ~n3446 ;
  assign y2588 = 1'b0 ;
  assign y2589 = n3456 ;
  assign y2590 = n3457 ;
  assign y2591 = n3458 ;
  assign y2592 = ~1'b0 ;
  assign y2593 = n3461 ;
  assign y2594 = ~n3464 ;
  assign y2595 = ~1'b0 ;
  assign y2596 = n3465 ;
  assign y2597 = ~1'b0 ;
  assign y2598 = ~1'b0 ;
  assign y2599 = n3466 ;
  assign y2600 = ~n3469 ;
  assign y2601 = n3472 ;
  assign y2602 = 1'b0 ;
  assign y2603 = n3473 ;
  assign y2604 = 1'b0 ;
  assign y2605 = n3475 ;
  assign y2606 = ~n1693 ;
  assign y2607 = ~1'b0 ;
  assign y2608 = ~1'b0 ;
  assign y2609 = ~1'b0 ;
  assign y2610 = n3477 ;
  assign y2611 = n1874 ;
  assign y2612 = ~1'b0 ;
  assign y2613 = ~n3481 ;
  assign y2614 = ~1'b0 ;
  assign y2615 = n3483 ;
  assign y2616 = ~1'b0 ;
  assign y2617 = n3487 ;
  assign y2618 = ~1'b0 ;
  assign y2619 = ~n3489 ;
  assign y2620 = 1'b0 ;
  assign y2621 = ~n1785 ;
  assign y2622 = ~1'b0 ;
  assign y2623 = n3443 ;
  assign y2624 = ~1'b0 ;
  assign y2625 = ~n3490 ;
  assign y2626 = n3493 ;
  assign y2627 = ~1'b0 ;
  assign y2628 = ~1'b0 ;
  assign y2629 = ~n3495 ;
  assign y2630 = ~1'b0 ;
  assign y2631 = ~1'b0 ;
  assign y2632 = n3498 ;
  assign y2633 = ~n3501 ;
  assign y2634 = ~n3503 ;
  assign y2635 = ~1'b0 ;
  assign y2636 = ~1'b0 ;
  assign y2637 = ~n3506 ;
  assign y2638 = ~n3509 ;
  assign y2639 = n3512 ;
  assign y2640 = ~1'b0 ;
  assign y2641 = ~n3513 ;
  assign y2642 = ~1'b0 ;
  assign y2643 = ~1'b0 ;
  assign y2644 = ~n1127 ;
  assign y2645 = ~n3514 ;
  assign y2646 = ~1'b0 ;
  assign y2647 = ~1'b0 ;
  assign y2648 = n3516 ;
  assign y2649 = ~1'b0 ;
  assign y2650 = ~n3522 ;
  assign y2651 = n1961 ;
  assign y2652 = ~n3527 ;
  assign y2653 = n3532 ;
  assign y2654 = ~n3533 ;
  assign y2655 = n2532 ;
  assign y2656 = ~1'b0 ;
  assign y2657 = ~1'b0 ;
  assign y2658 = n3534 ;
  assign y2659 = 1'b0 ;
  assign y2660 = n3537 ;
  assign y2661 = ~n3540 ;
  assign y2662 = ~1'b0 ;
  assign y2663 = ~1'b0 ;
  assign y2664 = n3542 ;
  assign y2665 = ~n3546 ;
  assign y2666 = n3548 ;
  assign y2667 = n3556 ;
  assign y2668 = ~1'b0 ;
  assign y2669 = ~n3559 ;
  assign y2670 = ~1'b0 ;
  assign y2671 = ~1'b0 ;
  assign y2672 = ~1'b0 ;
  assign y2673 = n3472 ;
  assign y2674 = ~1'b0 ;
  assign y2675 = ~n3564 ;
  assign y2676 = ~n3567 ;
  assign y2677 = n3571 ;
  assign y2678 = n3574 ;
  assign y2679 = ~n1026 ;
  assign y2680 = n3576 ;
  assign y2681 = ~n594 ;
  assign y2682 = ~n3577 ;
  assign y2683 = ~1'b0 ;
  assign y2684 = ~1'b0 ;
  assign y2685 = n3579 ;
  assign y2686 = ~1'b0 ;
  assign y2687 = ~1'b0 ;
  assign y2688 = ~1'b0 ;
  assign y2689 = n3580 ;
  assign y2690 = ~1'b0 ;
  assign y2691 = ~1'b0 ;
  assign y2692 = ~n3581 ;
  assign y2693 = n3583 ;
  assign y2694 = ~1'b0 ;
  assign y2695 = ~1'b0 ;
  assign y2696 = n3584 ;
  assign y2697 = ~n3585 ;
  assign y2698 = n3592 ;
  assign y2699 = ~1'b0 ;
  assign y2700 = ~n3593 ;
  assign y2701 = ~n3597 ;
  assign y2702 = ~1'b0 ;
  assign y2703 = ~1'b0 ;
  assign y2704 = ~1'b0 ;
  assign y2705 = ~n3599 ;
  assign y2706 = 1'b0 ;
  assign y2707 = ~1'b0 ;
  assign y2708 = 1'b0 ;
  assign y2709 = n3600 ;
  assign y2710 = ~n3603 ;
  assign y2711 = n3604 ;
  assign y2712 = ~1'b0 ;
  assign y2713 = ~1'b0 ;
  assign y2714 = 1'b0 ;
  assign y2715 = ~1'b0 ;
  assign y2716 = n3606 ;
  assign y2717 = ~n2512 ;
  assign y2718 = ~n3616 ;
  assign y2719 = ~n3617 ;
  assign y2720 = ~1'b0 ;
  assign y2721 = ~1'b0 ;
  assign y2722 = ~1'b0 ;
  assign y2723 = ~n3622 ;
  assign y2724 = ~1'b0 ;
  assign y2725 = 1'b0 ;
  assign y2726 = ~n3632 ;
  assign y2727 = ~1'b0 ;
  assign y2728 = ~1'b0 ;
  assign y2729 = n3635 ;
  assign y2730 = ~n3636 ;
  assign y2731 = n3637 ;
  assign y2732 = ~n3640 ;
  assign y2733 = ~1'b0 ;
  assign y2734 = ~n3641 ;
  assign y2735 = ~1'b0 ;
  assign y2736 = n3643 ;
  assign y2737 = ~1'b0 ;
  assign y2738 = ~n3646 ;
  assign y2739 = ~1'b0 ;
  assign y2740 = ~1'b0 ;
  assign y2741 = ~1'b0 ;
  assign y2742 = n3648 ;
  assign y2743 = ~1'b0 ;
  assign y2744 = ~n3650 ;
  assign y2745 = ~n1748 ;
  assign y2746 = n3655 ;
  assign y2747 = n507 ;
  assign y2748 = ~n3659 ;
  assign y2749 = n3665 ;
  assign y2750 = ~1'b0 ;
  assign y2751 = ~1'b0 ;
  assign y2752 = ~1'b0 ;
  assign y2753 = n3668 ;
  assign y2754 = ~n3670 ;
  assign y2755 = ~n3671 ;
  assign y2756 = n3676 ;
  assign y2757 = ~n3678 ;
  assign y2758 = n3680 ;
  assign y2759 = n3681 ;
  assign y2760 = ~n3688 ;
  assign y2761 = ~1'b0 ;
  assign y2762 = ~n3696 ;
  assign y2763 = ~n1933 ;
  assign y2764 = ~1'b0 ;
  assign y2765 = ~n3698 ;
  assign y2766 = ~n3040 ;
  assign y2767 = ~1'b0 ;
  assign y2768 = ~1'b0 ;
  assign y2769 = n2933 ;
  assign y2770 = ~1'b0 ;
  assign y2771 = ~1'b0 ;
  assign y2772 = n3087 ;
  assign y2773 = n3701 ;
  assign y2774 = ~1'b0 ;
  assign y2775 = n3702 ;
  assign y2776 = n3704 ;
  assign y2777 = n3706 ;
  assign y2778 = ~n2519 ;
  assign y2779 = n3707 ;
  assign y2780 = ~n3708 ;
  assign y2781 = ~n1505 ;
  assign y2782 = n2436 ;
  assign y2783 = ~1'b0 ;
  assign y2784 = ~n3709 ;
  assign y2785 = ~1'b0 ;
  assign y2786 = x6 ;
  assign y2787 = n3718 ;
  assign y2788 = 1'b0 ;
  assign y2789 = ~n3724 ;
  assign y2790 = ~n3727 ;
  assign y2791 = n3282 ;
  assign y2792 = ~1'b0 ;
  assign y2793 = ~n3732 ;
  assign y2794 = ~1'b0 ;
  assign y2795 = ~1'b0 ;
  assign y2796 = ~1'b0 ;
  assign y2797 = ~1'b0 ;
  assign y2798 = ~1'b0 ;
  assign y2799 = ~1'b0 ;
  assign y2800 = 1'b0 ;
  assign y2801 = ~1'b0 ;
  assign y2802 = n3737 ;
  assign y2803 = 1'b0 ;
  assign y2804 = ~1'b0 ;
  assign y2805 = ~1'b0 ;
  assign y2806 = ~n3738 ;
  assign y2807 = ~1'b0 ;
  assign y2808 = n3741 ;
  assign y2809 = ~1'b0 ;
  assign y2810 = n3744 ;
  assign y2811 = ~1'b0 ;
  assign y2812 = ~1'b0 ;
  assign y2813 = ~n3103 ;
  assign y2814 = ~1'b0 ;
  assign y2815 = n3746 ;
  assign y2816 = ~1'b0 ;
  assign y2817 = ~n3748 ;
  assign y2818 = ~1'b0 ;
  assign y2819 = ~n216 ;
  assign y2820 = ~n3749 ;
  assign y2821 = n3750 ;
  assign y2822 = n3752 ;
  assign y2823 = ~1'b0 ;
  assign y2824 = n3753 ;
  assign y2825 = ~1'b0 ;
  assign y2826 = ~n3542 ;
  assign y2827 = ~n3758 ;
  assign y2828 = n3761 ;
  assign y2829 = ~n3589 ;
  assign y2830 = n3762 ;
  assign y2831 = ~n3080 ;
  assign y2832 = ~1'b0 ;
  assign y2833 = ~1'b0 ;
  assign y2834 = 1'b0 ;
  assign y2835 = n879 ;
  assign y2836 = ~1'b0 ;
  assign y2837 = ~1'b0 ;
  assign y2838 = ~n741 ;
  assign y2839 = ~1'b0 ;
  assign y2840 = ~n954 ;
  assign y2841 = ~1'b0 ;
  assign y2842 = ~n3764 ;
  assign y2843 = ~n3766 ;
  assign y2844 = n3769 ;
  assign y2845 = ~1'b0 ;
  assign y2846 = ~1'b0 ;
  assign y2847 = ~n3775 ;
  assign y2848 = ~n3777 ;
  assign y2849 = n3778 ;
  assign y2850 = ~n3779 ;
  assign y2851 = ~n3270 ;
  assign y2852 = ~1'b0 ;
  assign y2853 = ~1'b0 ;
  assign y2854 = ~1'b0 ;
  assign y2855 = ~1'b0 ;
  assign y2856 = ~1'b0 ;
  assign y2857 = n3780 ;
  assign y2858 = ~1'b0 ;
  assign y2859 = ~1'b0 ;
  assign y2860 = ~1'b0 ;
  assign y2861 = ~1'b0 ;
  assign y2862 = n3781 ;
  assign y2863 = ~n3782 ;
  assign y2864 = ~1'b0 ;
  assign y2865 = ~1'b0 ;
  assign y2866 = n3784 ;
  assign y2867 = n3785 ;
  assign y2868 = ~n3786 ;
  assign y2869 = ~1'b0 ;
  assign y2870 = ~1'b0 ;
  assign y2871 = ~n3789 ;
  assign y2872 = ~n3791 ;
  assign y2873 = ~n3792 ;
  assign y2874 = n3796 ;
  assign y2875 = 1'b0 ;
  assign y2876 = n3797 ;
  assign y2877 = ~n141 ;
  assign y2878 = n3798 ;
  assign y2879 = ~1'b0 ;
  assign y2880 = ~1'b0 ;
  assign y2881 = n3799 ;
  assign y2882 = ~n3800 ;
  assign y2883 = ~n3802 ;
  assign y2884 = ~1'b0 ;
  assign y2885 = ~1'b0 ;
  assign y2886 = n3804 ;
  assign y2887 = ~n3805 ;
  assign y2888 = ~n3806 ;
  assign y2889 = ~n636 ;
  assign y2890 = n3807 ;
  assign y2891 = ~1'b0 ;
  assign y2892 = ~1'b0 ;
  assign y2893 = ~n3808 ;
  assign y2894 = ~1'b0 ;
  assign y2895 = n3810 ;
  assign y2896 = ~n3509 ;
  assign y2897 = n3812 ;
  assign y2898 = n3813 ;
  assign y2899 = n3814 ;
  assign y2900 = n3817 ;
  assign y2901 = ~1'b0 ;
  assign y2902 = n3818 ;
  assign y2903 = ~1'b0 ;
  assign y2904 = ~n3821 ;
  assign y2905 = ~1'b0 ;
  assign y2906 = n227 ;
  assign y2907 = n3823 ;
  assign y2908 = ~1'b0 ;
  assign y2909 = n3826 ;
  assign y2910 = ~n3828 ;
  assign y2911 = ~n3832 ;
  assign y2912 = n3835 ;
  assign y2913 = ~n3836 ;
  assign y2914 = n1174 ;
  assign y2915 = ~n3839 ;
  assign y2916 = n3841 ;
  assign y2917 = ~n175 ;
  assign y2918 = ~1'b0 ;
  assign y2919 = ~1'b0 ;
  assign y2920 = ~n3843 ;
  assign y2921 = n37 ;
  assign y2922 = ~1'b0 ;
  assign y2923 = n3844 ;
  assign y2924 = ~1'b0 ;
  assign y2925 = ~n3845 ;
  assign y2926 = ~n3848 ;
  assign y2927 = ~1'b0 ;
  assign y2928 = ~1'b0 ;
  assign y2929 = ~1'b0 ;
  assign y2930 = 1'b0 ;
  assign y2931 = ~n3850 ;
  assign y2932 = ~1'b0 ;
  assign y2933 = ~n3851 ;
  assign y2934 = n3791 ;
  assign y2935 = n300 ;
  assign y2936 = n3854 ;
  assign y2937 = ~n3856 ;
  assign y2938 = n1982 ;
  assign y2939 = n3858 ;
  assign y2940 = ~1'b0 ;
  assign y2941 = n3859 ;
  assign y2942 = ~n3862 ;
  assign y2943 = ~1'b0 ;
  assign y2944 = n3866 ;
  assign y2945 = n3868 ;
  assign y2946 = n2414 ;
  assign y2947 = n3871 ;
  assign y2948 = 1'b0 ;
  assign y2949 = ~n310 ;
  assign y2950 = ~n3874 ;
  assign y2951 = ~n3877 ;
  assign y2952 = n3878 ;
  assign y2953 = n3882 ;
  assign y2954 = ~1'b0 ;
  assign y2955 = ~1'b0 ;
  assign y2956 = n3885 ;
  assign y2957 = n3886 ;
  assign y2958 = ~1'b0 ;
  assign y2959 = ~1'b0 ;
  assign y2960 = n3888 ;
  assign y2961 = n3890 ;
  assign y2962 = ~1'b0 ;
  assign y2963 = ~n3891 ;
  assign y2964 = ~n3892 ;
  assign y2965 = ~n3893 ;
  assign y2966 = ~n3899 ;
  assign y2967 = ~n3905 ;
  assign y2968 = ~n3908 ;
  assign y2969 = n3909 ;
  assign y2970 = ~1'b0 ;
  assign y2971 = n3914 ;
  assign y2972 = n963 ;
  assign y2973 = n3916 ;
  assign y2974 = ~n3919 ;
  assign y2975 = n3921 ;
  assign y2976 = ~n3928 ;
  assign y2977 = ~1'b0 ;
  assign y2978 = ~1'b0 ;
  assign y2979 = ~n3929 ;
  assign y2980 = n2930 ;
  assign y2981 = ~1'b0 ;
  assign y2982 = ~1'b0 ;
  assign y2983 = ~n3931 ;
  assign y2984 = ~1'b0 ;
  assign y2985 = n3933 ;
  assign y2986 = n3939 ;
  assign y2987 = ~1'b0 ;
  assign y2988 = ~1'b0 ;
  assign y2989 = n3941 ;
  assign y2990 = ~1'b0 ;
  assign y2991 = ~n3945 ;
  assign y2992 = ~n3947 ;
  assign y2993 = ~n3949 ;
  assign y2994 = ~1'b0 ;
  assign y2995 = n3953 ;
  assign y2996 = ~1'b0 ;
  assign y2997 = ~1'b0 ;
  assign y2998 = n3954 ;
  assign y2999 = n3962 ;
  assign y3000 = ~1'b0 ;
  assign y3001 = ~1'b0 ;
  assign y3002 = ~1'b0 ;
  assign y3003 = ~1'b0 ;
  assign y3004 = ~n3964 ;
  assign y3005 = n3965 ;
  assign y3006 = n1133 ;
  assign y3007 = n3966 ;
  assign y3008 = n3969 ;
  assign y3009 = n3971 ;
  assign y3010 = n2235 ;
  assign y3011 = n1739 ;
  assign y3012 = ~1'b0 ;
  assign y3013 = ~1'b0 ;
  assign y3014 = ~n3589 ;
  assign y3015 = ~n3974 ;
  assign y3016 = ~1'b0 ;
  assign y3017 = ~n3978 ;
  assign y3018 = ~1'b0 ;
  assign y3019 = ~n3980 ;
  assign y3020 = ~1'b0 ;
  assign y3021 = n2837 ;
  assign y3022 = ~1'b0 ;
  assign y3023 = ~n3981 ;
  assign y3024 = n3604 ;
  assign y3025 = ~n3983 ;
  assign y3026 = n3992 ;
  assign y3027 = n3998 ;
  assign y3028 = ~1'b0 ;
  assign y3029 = ~n3999 ;
  assign y3030 = n2273 ;
  assign y3031 = n4003 ;
  assign y3032 = ~1'b0 ;
  assign y3033 = ~n4008 ;
  assign y3034 = ~n3803 ;
  assign y3035 = n4009 ;
  assign y3036 = n4010 ;
  assign y3037 = ~1'b0 ;
  assign y3038 = ~1'b0 ;
  assign y3039 = 1'b0 ;
  assign y3040 = ~1'b0 ;
  assign y3041 = ~n4012 ;
  assign y3042 = ~n636 ;
  assign y3043 = ~n3626 ;
  assign y3044 = ~1'b0 ;
  assign y3045 = ~n4018 ;
  assign y3046 = n4020 ;
  assign y3047 = n4021 ;
  assign y3048 = ~1'b0 ;
  assign y3049 = ~1'b0 ;
  assign y3050 = ~1'b0 ;
  assign y3051 = 1'b0 ;
  assign y3052 = ~n4023 ;
  assign y3053 = n4026 ;
  assign y3054 = ~1'b0 ;
  assign y3055 = ~1'b0 ;
  assign y3056 = ~n4027 ;
  assign y3057 = ~n4033 ;
  assign y3058 = ~x0 ;
  assign y3059 = ~n3339 ;
  assign y3060 = n4039 ;
  assign y3061 = n4042 ;
  assign y3062 = ~1'b0 ;
  assign y3063 = n4043 ;
  assign y3064 = ~n1550 ;
  assign y3065 = n4049 ;
  assign y3066 = n2850 ;
  assign y3067 = 1'b0 ;
  assign y3068 = ~1'b0 ;
  assign y3069 = n4051 ;
  assign y3070 = 1'b0 ;
  assign y3071 = n4053 ;
  assign y3072 = ~n4054 ;
  assign y3073 = n817 ;
  assign y3074 = ~n4057 ;
  assign y3075 = ~1'b0 ;
  assign y3076 = ~n4059 ;
  assign y3077 = ~n4060 ;
  assign y3078 = n4061 ;
  assign y3079 = n4068 ;
  assign y3080 = ~1'b0 ;
  assign y3081 = n2003 ;
  assign y3082 = ~n4069 ;
  assign y3083 = n4070 ;
  assign y3084 = n4075 ;
  assign y3085 = n4076 ;
  assign y3086 = ~n4078 ;
  assign y3087 = ~1'b0 ;
  assign y3088 = ~1'b0 ;
  assign y3089 = ~n4084 ;
  assign y3090 = ~1'b0 ;
  assign y3091 = ~1'b0 ;
  assign y3092 = ~1'b0 ;
  assign y3093 = ~1'b0 ;
  assign y3094 = n4088 ;
  assign y3095 = ~n987 ;
  assign y3096 = ~n4091 ;
  assign y3097 = ~n4092 ;
  assign y3098 = ~1'b0 ;
  assign y3099 = ~1'b0 ;
  assign y3100 = 1'b0 ;
  assign y3101 = ~n4095 ;
  assign y3102 = n4096 ;
  assign y3103 = ~1'b0 ;
  assign y3104 = ~1'b0 ;
  assign y3105 = ~1'b0 ;
  assign y3106 = ~1'b0 ;
  assign y3107 = n4097 ;
  assign y3108 = n4100 ;
  assign y3109 = ~n4102 ;
  assign y3110 = n4104 ;
  assign y3111 = n4105 ;
  assign y3112 = ~n460 ;
  assign y3113 = ~n4106 ;
  assign y3114 = ~1'b0 ;
  assign y3115 = n4108 ;
  assign y3116 = ~n4109 ;
  assign y3117 = ~n4111 ;
  assign y3118 = n4115 ;
  assign y3119 = n4117 ;
  assign y3120 = ~n4118 ;
  assign y3121 = ~n236 ;
  assign y3122 = ~n4120 ;
  assign y3123 = ~n4123 ;
  assign y3124 = ~1'b0 ;
  assign y3125 = ~1'b0 ;
  assign y3126 = ~n2774 ;
  assign y3127 = ~n4127 ;
  assign y3128 = n4132 ;
  assign y3129 = n4133 ;
  assign y3130 = ~n4139 ;
  assign y3131 = ~n3679 ;
  assign y3132 = n4140 ;
  assign y3133 = ~n4148 ;
  assign y3134 = ~1'b0 ;
  assign y3135 = ~1'b0 ;
  assign y3136 = n4152 ;
  assign y3137 = n4153 ;
  assign y3138 = ~1'b0 ;
  assign y3139 = 1'b0 ;
  assign y3140 = 1'b0 ;
  assign y3141 = ~n4158 ;
  assign y3142 = ~n4161 ;
  assign y3143 = ~n4165 ;
  assign y3144 = ~1'b0 ;
  assign y3145 = ~n4166 ;
  assign y3146 = n4167 ;
  assign y3147 = ~n4171 ;
  assign y3148 = ~n4174 ;
  assign y3149 = ~n4182 ;
  assign y3150 = n3177 ;
  assign y3151 = n627 ;
  assign y3152 = ~1'b0 ;
  assign y3153 = n4185 ;
  assign y3154 = n4189 ;
  assign y3155 = n4192 ;
  assign y3156 = n4194 ;
  assign y3157 = ~1'b0 ;
  assign y3158 = ~n4195 ;
  assign y3159 = n4196 ;
  assign y3160 = ~1'b0 ;
  assign y3161 = n4198 ;
  assign y3162 = ~1'b0 ;
  assign y3163 = ~1'b0 ;
  assign y3164 = n4202 ;
  assign y3165 = n4207 ;
  assign y3166 = ~1'b0 ;
  assign y3167 = n4210 ;
  assign y3168 = ~1'b0 ;
  assign y3169 = ~1'b0 ;
  assign y3170 = ~n4212 ;
  assign y3171 = ~1'b0 ;
  assign y3172 = ~n4216 ;
  assign y3173 = ~n4219 ;
  assign y3174 = ~1'b0 ;
  assign y3175 = ~1'b0 ;
  assign y3176 = ~1'b0 ;
  assign y3177 = n4221 ;
  assign y3178 = n4223 ;
  assign y3179 = n4228 ;
  assign y3180 = n4239 ;
  assign y3181 = ~n4246 ;
  assign y3182 = ~1'b0 ;
  assign y3183 = n4249 ;
  assign y3184 = ~1'b0 ;
  assign y3185 = n4251 ;
  assign y3186 = ~n4188 ;
  assign y3187 = ~1'b0 ;
  assign y3188 = ~n4254 ;
  assign y3189 = n4259 ;
  assign y3190 = n4261 ;
  assign y3191 = ~n4263 ;
  assign y3192 = n4264 ;
  assign y3193 = ~1'b0 ;
  assign y3194 = ~1'b0 ;
  assign y3195 = ~1'b0 ;
  assign y3196 = ~1'b0 ;
  assign y3197 = 1'b0 ;
  assign y3198 = ~n4269 ;
  assign y3199 = ~1'b0 ;
  assign y3200 = n4271 ;
  assign y3201 = ~1'b0 ;
  assign y3202 = 1'b0 ;
  assign y3203 = n4275 ;
  assign y3204 = ~1'b0 ;
  assign y3205 = ~n4278 ;
  assign y3206 = ~1'b0 ;
  assign y3207 = ~1'b0 ;
  assign y3208 = n2722 ;
  assign y3209 = n4279 ;
  assign y3210 = n1255 ;
  assign y3211 = ~1'b0 ;
  assign y3212 = n4280 ;
  assign y3213 = ~1'b0 ;
  assign y3214 = n2604 ;
  assign y3215 = ~n4285 ;
  assign y3216 = n4286 ;
  assign y3217 = n4291 ;
  assign y3218 = ~n4292 ;
  assign y3219 = ~1'b0 ;
  assign y3220 = n4293 ;
  assign y3221 = ~n4295 ;
  assign y3222 = n4296 ;
  assign y3223 = ~n4298 ;
  assign y3224 = ~1'b0 ;
  assign y3225 = ~1'b0 ;
  assign y3226 = ~1'b0 ;
  assign y3227 = ~n4299 ;
  assign y3228 = n4300 ;
  assign y3229 = n4303 ;
  assign y3230 = ~1'b0 ;
  assign y3231 = ~1'b0 ;
  assign y3232 = 1'b0 ;
  assign y3233 = ~n1772 ;
  assign y3234 = ~1'b0 ;
  assign y3235 = ~1'b0 ;
  assign y3236 = ~n532 ;
  assign y3237 = n4306 ;
  assign y3238 = ~1'b0 ;
  assign y3239 = ~n4308 ;
  assign y3240 = ~1'b0 ;
  assign y3241 = ~1'b0 ;
  assign y3242 = ~1'b0 ;
  assign y3243 = n4313 ;
  assign y3244 = ~1'b0 ;
  assign y3245 = n1707 ;
  assign y3246 = 1'b0 ;
  assign y3247 = n4314 ;
  assign y3248 = ~1'b0 ;
  assign y3249 = n4317 ;
  assign y3250 = n4318 ;
  assign y3251 = ~1'b0 ;
  assign y3252 = n4319 ;
  assign y3253 = n4321 ;
  assign y3254 = n4328 ;
  assign y3255 = n4329 ;
  assign y3256 = ~1'b0 ;
  assign y3257 = ~1'b0 ;
  assign y3258 = ~1'b0 ;
  assign y3259 = ~n4330 ;
  assign y3260 = n4337 ;
  assign y3261 = ~1'b0 ;
  assign y3262 = n4342 ;
  assign y3263 = n2594 ;
  assign y3264 = n3427 ;
  assign y3265 = ~1'b0 ;
  assign y3266 = ~n4346 ;
  assign y3267 = ~n4347 ;
  assign y3268 = n4348 ;
  assign y3269 = ~1'b0 ;
  assign y3270 = 1'b0 ;
  assign y3271 = ~1'b0 ;
  assign y3272 = n4353 ;
  assign y3273 = ~1'b0 ;
  assign y3274 = ~1'b0 ;
  assign y3275 = n4354 ;
  assign y3276 = n4356 ;
  assign y3277 = ~1'b0 ;
  assign y3278 = ~n4360 ;
  assign y3279 = 1'b0 ;
  assign y3280 = ~1'b0 ;
  assign y3281 = ~n4363 ;
  assign y3282 = 1'b0 ;
  assign y3283 = n4368 ;
  assign y3284 = n4369 ;
  assign y3285 = n4374 ;
  assign y3286 = ~1'b0 ;
  assign y3287 = ~1'b0 ;
  assign y3288 = ~1'b0 ;
  assign y3289 = ~n4378 ;
  assign y3290 = ~n4379 ;
  assign y3291 = ~n4381 ;
  assign y3292 = n4383 ;
  assign y3293 = ~n4389 ;
  assign y3294 = n4392 ;
  assign y3295 = n4394 ;
  assign y3296 = ~1'b0 ;
  assign y3297 = ~n4395 ;
  assign y3298 = n2964 ;
  assign y3299 = ~n4396 ;
  assign y3300 = ~n4398 ;
  assign y3301 = ~1'b0 ;
  assign y3302 = ~1'b0 ;
  assign y3303 = n4349 ;
  assign y3304 = ~n4400 ;
  assign y3305 = ~1'b0 ;
  assign y3306 = n4401 ;
  assign y3307 = n4403 ;
  assign y3308 = n4404 ;
  assign y3309 = n4406 ;
  assign y3310 = ~n4409 ;
  assign y3311 = n4411 ;
  assign y3312 = ~1'b0 ;
  assign y3313 = n4412 ;
  assign y3314 = n4416 ;
  assign y3315 = ~1'b0 ;
  assign y3316 = 1'b0 ;
  assign y3317 = n4419 ;
  assign y3318 = ~n4420 ;
  assign y3319 = ~n4421 ;
  assign y3320 = ~1'b0 ;
  assign y3321 = ~n4424 ;
  assign y3322 = ~1'b0 ;
  assign y3323 = n520 ;
  assign y3324 = ~n4430 ;
  assign y3325 = ~1'b0 ;
  assign y3326 = ~1'b0 ;
  assign y3327 = n4431 ;
  assign y3328 = ~1'b0 ;
  assign y3329 = n4436 ;
  assign y3330 = n4440 ;
  assign y3331 = n4441 ;
  assign y3332 = ~1'b0 ;
  assign y3333 = ~1'b0 ;
  assign y3334 = ~n4443 ;
  assign y3335 = n3415 ;
  assign y3336 = ~1'b0 ;
  assign y3337 = n4446 ;
  assign y3338 = ~n4449 ;
  assign y3339 = ~n4450 ;
  assign y3340 = ~1'b0 ;
  assign y3341 = ~1'b0 ;
  assign y3342 = ~n1699 ;
  assign y3343 = 1'b0 ;
  assign y3344 = ~1'b0 ;
  assign y3345 = ~n2027 ;
  assign y3346 = ~n4451 ;
  assign y3347 = n4456 ;
  assign y3348 = ~1'b0 ;
  assign y3349 = ~n4463 ;
  assign y3350 = ~1'b0 ;
  assign y3351 = ~1'b0 ;
  assign y3352 = ~n4465 ;
  assign y3353 = ~1'b0 ;
  assign y3354 = ~n4466 ;
  assign y3355 = ~n4468 ;
  assign y3356 = ~n4471 ;
  assign y3357 = n4473 ;
  assign y3358 = n4474 ;
  assign y3359 = n4479 ;
  assign y3360 = ~n4481 ;
  assign y3361 = n4482 ;
  assign y3362 = ~1'b0 ;
  assign y3363 = n4485 ;
  assign y3364 = ~n4400 ;
  assign y3365 = ~1'b0 ;
  assign y3366 = ~n4492 ;
  assign y3367 = ~n4497 ;
  assign y3368 = 1'b0 ;
  assign y3369 = ~1'b0 ;
  assign y3370 = ~1'b0 ;
  assign y3371 = n4499 ;
  assign y3372 = n4506 ;
  assign y3373 = ~1'b0 ;
  assign y3374 = ~n4508 ;
  assign y3375 = n4509 ;
  assign y3376 = ~n4513 ;
  assign y3377 = n4516 ;
  assign y3378 = 1'b0 ;
  assign y3379 = 1'b0 ;
  assign y3380 = ~1'b0 ;
  assign y3381 = ~n1469 ;
  assign y3382 = 1'b0 ;
  assign y3383 = ~n4519 ;
  assign y3384 = n4520 ;
  assign y3385 = ~n4521 ;
  assign y3386 = 1'b0 ;
  assign y3387 = n4522 ;
  assign y3388 = ~1'b0 ;
  assign y3389 = ~n4526 ;
  assign y3390 = ~1'b0 ;
  assign y3391 = n2380 ;
  assign y3392 = ~1'b0 ;
  assign y3393 = ~1'b0 ;
  assign y3394 = ~n4528 ;
  assign y3395 = ~n2546 ;
  assign y3396 = ~n4537 ;
  assign y3397 = ~n4538 ;
  assign y3398 = n4540 ;
  assign y3399 = ~n4541 ;
  assign y3400 = ~n4543 ;
  assign y3401 = ~1'b0 ;
  assign y3402 = ~n4544 ;
  assign y3403 = ~1'b0 ;
  assign y3404 = n4546 ;
  assign y3405 = ~1'b0 ;
  assign y3406 = ~1'b0 ;
  assign y3407 = ~n4548 ;
  assign y3408 = ~1'b0 ;
  assign y3409 = n4549 ;
  assign y3410 = ~1'b0 ;
  assign y3411 = n715 ;
  assign y3412 = ~1'b0 ;
  assign y3413 = ~1'b0 ;
  assign y3414 = ~n4551 ;
  assign y3415 = ~1'b0 ;
  assign y3416 = n4552 ;
  assign y3417 = n4556 ;
  assign y3418 = 1'b0 ;
  assign y3419 = n2695 ;
  assign y3420 = ~n4557 ;
  assign y3421 = ~n4565 ;
  assign y3422 = n4567 ;
  assign y3423 = ~1'b0 ;
  assign y3424 = ~n3371 ;
  assign y3425 = n4569 ;
  assign y3426 = ~n4570 ;
  assign y3427 = n4573 ;
  assign y3428 = ~n4575 ;
  assign y3429 = n4582 ;
  assign y3430 = ~n4585 ;
  assign y3431 = ~1'b0 ;
  assign y3432 = ~1'b0 ;
  assign y3433 = 1'b0 ;
  assign y3434 = ~n4588 ;
  assign y3435 = ~1'b0 ;
  assign y3436 = ~1'b0 ;
  assign y3437 = n4600 ;
  assign y3438 = n4604 ;
  assign y3439 = ~n4609 ;
  assign y3440 = ~1'b0 ;
  assign y3441 = ~n613 ;
  assign y3442 = n4610 ;
  assign y3443 = ~n4618 ;
  assign y3444 = ~1'b0 ;
  assign y3445 = ~1'b0 ;
  assign y3446 = ~n4619 ;
  assign y3447 = ~1'b0 ;
  assign y3448 = ~1'b0 ;
  assign y3449 = ~1'b0 ;
  assign y3450 = ~n4620 ;
  assign y3451 = ~n4623 ;
  assign y3452 = ~1'b0 ;
  assign y3453 = n4628 ;
  assign y3454 = n4634 ;
  assign y3455 = ~1'b0 ;
  assign y3456 = ~n4636 ;
  assign y3457 = ~n613 ;
  assign y3458 = n4638 ;
  assign y3459 = ~1'b0 ;
  assign y3460 = ~1'b0 ;
  assign y3461 = n4640 ;
  assign y3462 = ~1'b0 ;
  assign y3463 = n1112 ;
  assign y3464 = n270 ;
  assign y3465 = n1385 ;
  assign y3466 = n4643 ;
  assign y3467 = ~n4645 ;
  assign y3468 = ~n36 ;
  assign y3469 = ~n4646 ;
  assign y3470 = ~1'b0 ;
  assign y3471 = n4647 ;
  assign y3472 = n4654 ;
  assign y3473 = ~n4655 ;
  assign y3474 = ~n4657 ;
  assign y3475 = 1'b0 ;
  assign y3476 = ~1'b0 ;
  assign y3477 = ~n4659 ;
  assign y3478 = n4661 ;
  assign y3479 = n4662 ;
  assign y3480 = ~1'b0 ;
  assign y3481 = ~n4664 ;
  assign y3482 = ~n4666 ;
  assign y3483 = ~n4667 ;
  assign y3484 = 1'b0 ;
  assign y3485 = 1'b0 ;
  assign y3486 = n4668 ;
  assign y3487 = n1878 ;
  assign y3488 = ~n4671 ;
  assign y3489 = ~1'b0 ;
  assign y3490 = 1'b0 ;
  assign y3491 = ~n4673 ;
  assign y3492 = 1'b0 ;
  assign y3493 = 1'b0 ;
  assign y3494 = ~n4674 ;
  assign y3495 = ~1'b0 ;
  assign y3496 = ~1'b0 ;
  assign y3497 = ~1'b0 ;
  assign y3498 = ~n4679 ;
  assign y3499 = ~1'b0 ;
  assign y3500 = 1'b0 ;
  assign y3501 = ~1'b0 ;
  assign y3502 = ~1'b0 ;
  assign y3503 = ~n4687 ;
  assign y3504 = ~1'b0 ;
  assign y3505 = n4690 ;
  assign y3506 = ~n4694 ;
  assign y3507 = ~1'b0 ;
  assign y3508 = ~1'b0 ;
  assign y3509 = ~n4695 ;
  assign y3510 = ~1'b0 ;
  assign y3511 = n4698 ;
  assign y3512 = 1'b0 ;
  assign y3513 = ~1'b0 ;
  assign y3514 = n4700 ;
  assign y3515 = ~n1000 ;
  assign y3516 = ~n4701 ;
  assign y3517 = n4703 ;
  assign y3518 = n1668 ;
  assign y3519 = n4704 ;
  assign y3520 = n4706 ;
  assign y3521 = ~1'b0 ;
  assign y3522 = n4708 ;
  assign y3523 = ~1'b0 ;
  assign y3524 = n4712 ;
  assign y3525 = n4714 ;
  assign y3526 = ~n3037 ;
  assign y3527 = ~n4716 ;
  assign y3528 = ~n4718 ;
  assign y3529 = n4722 ;
  assign y3530 = ~n4724 ;
  assign y3531 = n4726 ;
  assign y3532 = ~n4729 ;
  assign y3533 = n4731 ;
  assign y3534 = ~1'b0 ;
  assign y3535 = ~n4735 ;
  assign y3536 = ~1'b0 ;
  assign y3537 = n4740 ;
  assign y3538 = n1602 ;
  assign y3539 = n4742 ;
  assign y3540 = ~n4743 ;
  assign y3541 = ~n4747 ;
  assign y3542 = n4750 ;
  assign y3543 = ~n4751 ;
  assign y3544 = ~1'b0 ;
  assign y3545 = n4752 ;
  assign y3546 = n4754 ;
  assign y3547 = n4756 ;
  assign y3548 = n4759 ;
  assign y3549 = n4760 ;
  assign y3550 = 1'b0 ;
  assign y3551 = n4761 ;
  assign y3552 = ~n813 ;
  assign y3553 = n4764 ;
  assign y3554 = n4765 ;
  assign y3555 = ~1'b0 ;
  assign y3556 = ~n4767 ;
  assign y3557 = ~n4770 ;
  assign y3558 = n4772 ;
  assign y3559 = ~n4775 ;
  assign y3560 = n4776 ;
  assign y3561 = n3477 ;
  assign y3562 = n4777 ;
  assign y3563 = n68 ;
  assign y3564 = n4778 ;
  assign y3565 = ~1'b0 ;
  assign y3566 = n4780 ;
  assign y3567 = n4781 ;
  assign y3568 = ~n4784 ;
  assign y3569 = ~1'b0 ;
  assign y3570 = ~n4787 ;
  assign y3571 = n4788 ;
  assign y3572 = n321 ;
  assign y3573 = 1'b0 ;
  assign y3574 = ~n281 ;
  assign y3575 = ~n4796 ;
  assign y3576 = ~1'b0 ;
  assign y3577 = ~1'b0 ;
  assign y3578 = n4798 ;
  assign y3579 = ~1'b0 ;
  assign y3580 = ~n4800 ;
  assign y3581 = ~1'b0 ;
  assign y3582 = ~1'b0 ;
  assign y3583 = ~n4803 ;
  assign y3584 = ~n4809 ;
  assign y3585 = ~1'b0 ;
  assign y3586 = ~n4813 ;
  assign y3587 = n4814 ;
  assign y3588 = ~n4816 ;
  assign y3589 = n4817 ;
  assign y3590 = n4823 ;
  assign y3591 = ~n4824 ;
  assign y3592 = n4825 ;
  assign y3593 = ~n4827 ;
  assign y3594 = n4836 ;
  assign y3595 = ~1'b0 ;
  assign y3596 = n1388 ;
  assign y3597 = ~1'b0 ;
  assign y3598 = ~1'b0 ;
  assign y3599 = ~n4842 ;
  assign y3600 = ~n4843 ;
  assign y3601 = ~1'b0 ;
  assign y3602 = ~n4844 ;
  assign y3603 = n4845 ;
  assign y3604 = ~n3744 ;
  assign y3605 = n4851 ;
  assign y3606 = n469 ;
  assign y3607 = ~n4853 ;
  assign y3608 = ~1'b0 ;
  assign y3609 = ~1'b0 ;
  assign y3610 = n636 ;
  assign y3611 = ~n4856 ;
  assign y3612 = ~n4859 ;
  assign y3613 = n4862 ;
  assign y3614 = ~1'b0 ;
  assign y3615 = ~1'b0 ;
  assign y3616 = n4865 ;
  assign y3617 = ~1'b0 ;
  assign y3618 = n4867 ;
  assign y3619 = n4869 ;
  assign y3620 = ~1'b0 ;
  assign y3621 = ~1'b0 ;
  assign y3622 = ~n4873 ;
  assign y3623 = ~n4874 ;
  assign y3624 = n4875 ;
  assign y3625 = n4877 ;
  assign y3626 = ~n653 ;
  assign y3627 = n4878 ;
  assign y3628 = ~1'b0 ;
  assign y3629 = ~1'b0 ;
  assign y3630 = ~n4880 ;
  assign y3631 = ~1'b0 ;
  assign y3632 = n3378 ;
  assign y3633 = ~1'b0 ;
  assign y3634 = ~1'b0 ;
  assign y3635 = n4884 ;
  assign y3636 = ~1'b0 ;
  assign y3637 = ~n4885 ;
  assign y3638 = n4887 ;
  assign y3639 = ~1'b0 ;
  assign y3640 = ~1'b0 ;
  assign y3641 = ~1'b0 ;
  assign y3642 = ~1'b0 ;
  assign y3643 = n4890 ;
  assign y3644 = ~n4891 ;
  assign y3645 = n4893 ;
  assign y3646 = n4897 ;
  assign y3647 = ~n4898 ;
  assign y3648 = ~1'b0 ;
  assign y3649 = ~n4899 ;
  assign y3650 = n4900 ;
  assign y3651 = ~1'b0 ;
  assign y3652 = ~n4904 ;
  assign y3653 = ~n4907 ;
  assign y3654 = ~n4320 ;
  assign y3655 = ~n4909 ;
  assign y3656 = ~n4533 ;
  assign y3657 = n2263 ;
  assign y3658 = ~1'b0 ;
  assign y3659 = n4911 ;
  assign y3660 = ~1'b0 ;
  assign y3661 = ~1'b0 ;
  assign y3662 = n4913 ;
  assign y3663 = ~n3598 ;
  assign y3664 = n4916 ;
  assign y3665 = n4917 ;
  assign y3666 = ~1'b0 ;
  assign y3667 = n4921 ;
  assign y3668 = ~n4923 ;
  assign y3669 = ~1'b0 ;
  assign y3670 = n4924 ;
  assign y3671 = ~1'b0 ;
  assign y3672 = ~n4926 ;
  assign y3673 = ~1'b0 ;
  assign y3674 = ~n4929 ;
  assign y3675 = n4931 ;
  assign y3676 = ~1'b0 ;
  assign y3677 = ~n4933 ;
  assign y3678 = n4936 ;
  assign y3679 = ~n4938 ;
  assign y3680 = ~1'b0 ;
  assign y3681 = ~n4942 ;
  assign y3682 = n4943 ;
  assign y3683 = ~n4947 ;
  assign y3684 = ~n3366 ;
  assign y3685 = ~1'b0 ;
  assign y3686 = n4951 ;
  assign y3687 = ~n4955 ;
  assign y3688 = ~n4956 ;
  assign y3689 = n4965 ;
  assign y3690 = ~n4967 ;
  assign y3691 = ~n2799 ;
  assign y3692 = n4969 ;
  assign y3693 = ~n4972 ;
  assign y3694 = ~n4974 ;
  assign y3695 = ~1'b0 ;
  assign y3696 = ~n4976 ;
  assign y3697 = ~n4977 ;
  assign y3698 = 1'b0 ;
  assign y3699 = ~n2849 ;
  assign y3700 = ~1'b0 ;
  assign y3701 = ~1'b0 ;
  assign y3702 = ~1'b0 ;
  assign y3703 = ~1'b0 ;
  assign y3704 = ~n4986 ;
  assign y3705 = ~1'b0 ;
  assign y3706 = ~n4988 ;
  assign y3707 = ~1'b0 ;
  assign y3708 = ~1'b0 ;
  assign y3709 = n4991 ;
  assign y3710 = n4993 ;
  assign y3711 = n4995 ;
  assign y3712 = ~n4996 ;
  assign y3713 = ~1'b0 ;
  assign y3714 = ~n4998 ;
  assign y3715 = ~n5000 ;
  assign y3716 = ~n5004 ;
  assign y3717 = n5005 ;
  assign y3718 = ~n5008 ;
  assign y3719 = n1632 ;
  assign y3720 = ~1'b0 ;
  assign y3721 = 1'b0 ;
  assign y3722 = ~1'b0 ;
  assign y3723 = ~n5011 ;
  assign y3724 = 1'b0 ;
  assign y3725 = ~1'b0 ;
  assign y3726 = n5013 ;
  assign y3727 = ~n5023 ;
  assign y3728 = n5025 ;
  assign y3729 = ~1'b0 ;
  assign y3730 = n5026 ;
  assign y3731 = n5028 ;
  assign y3732 = ~1'b0 ;
  assign y3733 = ~1'b0 ;
  assign y3734 = n5030 ;
  assign y3735 = ~1'b0 ;
  assign y3736 = n5031 ;
  assign y3737 = n5032 ;
  assign y3738 = n726 ;
  assign y3739 = n5034 ;
  assign y3740 = ~n4439 ;
  assign y3741 = ~1'b0 ;
  assign y3742 = ~1'b0 ;
  assign y3743 = ~1'b0 ;
  assign y3744 = n5039 ;
  assign y3745 = ~1'b0 ;
  assign y3746 = ~n354 ;
  assign y3747 = n5043 ;
  assign y3748 = n5046 ;
  assign y3749 = 1'b0 ;
  assign y3750 = n5050 ;
  assign y3751 = n5051 ;
  assign y3752 = n5053 ;
  assign y3753 = ~1'b0 ;
  assign y3754 = n5056 ;
  assign y3755 = ~n5059 ;
  assign y3756 = ~n5060 ;
  assign y3757 = ~1'b0 ;
  assign y3758 = n5066 ;
  assign y3759 = ~1'b0 ;
  assign y3760 = ~1'b0 ;
  assign y3761 = ~n5067 ;
  assign y3762 = ~1'b0 ;
  assign y3763 = ~n5068 ;
  assign y3764 = ~n5074 ;
  assign y3765 = ~1'b0 ;
  assign y3766 = n5076 ;
  assign y3767 = ~n5078 ;
  assign y3768 = ~n5084 ;
  assign y3769 = ~n5095 ;
  assign y3770 = 1'b0 ;
  assign y3771 = ~1'b0 ;
  assign y3772 = ~n5101 ;
  assign y3773 = ~1'b0 ;
  assign y3774 = n5102 ;
  assign y3775 = ~1'b0 ;
  assign y3776 = n3890 ;
  assign y3777 = n5103 ;
  assign y3778 = ~n5104 ;
  assign y3779 = ~n4407 ;
  assign y3780 = ~1'b0 ;
  assign y3781 = 1'b0 ;
  assign y3782 = n5106 ;
  assign y3783 = ~n5110 ;
  assign y3784 = ~1'b0 ;
  assign y3785 = ~1'b0 ;
  assign y3786 = ~1'b0 ;
  assign y3787 = ~n5116 ;
  assign y3788 = ~1'b0 ;
  assign y3789 = ~n5118 ;
  assign y3790 = n246 ;
  assign y3791 = ~1'b0 ;
  assign y3792 = n5119 ;
  assign y3793 = ~1'b0 ;
  assign y3794 = n785 ;
  assign y3795 = ~n5121 ;
  assign y3796 = ~n5123 ;
  assign y3797 = ~1'b0 ;
  assign y3798 = n366 ;
  assign y3799 = n5125 ;
  assign y3800 = n5126 ;
  assign y3801 = n375 ;
  assign y3802 = n5127 ;
  assign y3803 = ~n5128 ;
  assign y3804 = n5130 ;
  assign y3805 = ~1'b0 ;
  assign y3806 = ~1'b0 ;
  assign y3807 = ~n5133 ;
  assign y3808 = n1655 ;
  assign y3809 = ~1'b0 ;
  assign y3810 = ~n2988 ;
  assign y3811 = ~1'b0 ;
  assign y3812 = n5134 ;
  assign y3813 = ~1'b0 ;
  assign y3814 = n4653 ;
  assign y3815 = n5135 ;
  assign y3816 = ~1'b0 ;
  assign y3817 = n5136 ;
  assign y3818 = ~1'b0 ;
  assign y3819 = ~n5138 ;
  assign y3820 = ~1'b0 ;
  assign y3821 = ~1'b0 ;
  assign y3822 = ~1'b0 ;
  assign y3823 = ~n5140 ;
  assign y3824 = ~n5141 ;
  assign y3825 = ~1'b0 ;
  assign y3826 = n5142 ;
  assign y3827 = ~n5143 ;
  assign y3828 = n5145 ;
  assign y3829 = n5146 ;
  assign y3830 = ~n3845 ;
  assign y3831 = ~1'b0 ;
  assign y3832 = n5149 ;
  assign y3833 = ~1'b0 ;
  assign y3834 = n5152 ;
  assign y3835 = ~1'b0 ;
  assign y3836 = n5154 ;
  assign y3837 = ~1'b0 ;
  assign y3838 = n3477 ;
  assign y3839 = ~1'b0 ;
  assign y3840 = ~1'b0 ;
  assign y3841 = ~n5155 ;
  assign y3842 = ~1'b0 ;
  assign y3843 = ~1'b0 ;
  assign y3844 = ~1'b0 ;
  assign y3845 = ~1'b0 ;
  assign y3846 = ~1'b0 ;
  assign y3847 = ~n1159 ;
  assign y3848 = ~n5156 ;
  assign y3849 = ~n573 ;
  assign y3850 = n5162 ;
  assign y3851 = ~n5164 ;
  assign y3852 = ~1'b0 ;
  assign y3853 = ~1'b0 ;
  assign y3854 = ~n5167 ;
  assign y3855 = ~1'b0 ;
  assign y3856 = ~n4349 ;
  assign y3857 = n5172 ;
  assign y3858 = n5174 ;
  assign y3859 = ~n5176 ;
  assign y3860 = n5178 ;
  assign y3861 = n1763 ;
  assign y3862 = n5179 ;
  assign y3863 = ~1'b0 ;
  assign y3864 = n5183 ;
  assign y3865 = ~n2751 ;
  assign y3866 = ~1'b0 ;
  assign y3867 = ~n532 ;
  assign y3868 = ~n5185 ;
  assign y3869 = ~n1226 ;
  assign y3870 = ~1'b0 ;
  assign y3871 = n5192 ;
  assign y3872 = n5194 ;
  assign y3873 = ~1'b0 ;
  assign y3874 = ~1'b0 ;
  assign y3875 = ~n5199 ;
  assign y3876 = ~n339 ;
  assign y3877 = n5204 ;
  assign y3878 = ~n2843 ;
  assign y3879 = n616 ;
  assign y3880 = n5208 ;
  assign y3881 = ~n5209 ;
  assign y3882 = n5187 ;
  assign y3883 = ~1'b0 ;
  assign y3884 = n5210 ;
  assign y3885 = ~n1768 ;
  assign y3886 = ~n5212 ;
  assign y3887 = ~n5214 ;
  assign y3888 = ~n5215 ;
  assign y3889 = n2148 ;
  assign y3890 = ~n5217 ;
  assign y3891 = n1431 ;
  assign y3892 = n5218 ;
  assign y3893 = n2203 ;
  assign y3894 = ~n726 ;
  assign y3895 = ~n5219 ;
  assign y3896 = ~1'b0 ;
  assign y3897 = ~1'b0 ;
  assign y3898 = ~1'b0 ;
  assign y3899 = n5225 ;
  assign y3900 = ~1'b0 ;
  assign y3901 = n5226 ;
  assign y3902 = n5231 ;
  assign y3903 = n759 ;
  assign y3904 = ~n5232 ;
  assign y3905 = n5234 ;
  assign y3906 = n4319 ;
  assign y3907 = ~n5235 ;
  assign y3908 = ~1'b0 ;
  assign y3909 = ~n5237 ;
  assign y3910 = ~1'b0 ;
  assign y3911 = ~1'b0 ;
  assign y3912 = n5238 ;
  assign y3913 = 1'b0 ;
  assign y3914 = ~n5239 ;
  assign y3915 = 1'b0 ;
  assign y3916 = ~n5241 ;
  assign y3917 = ~n5247 ;
  assign y3918 = n4311 ;
  assign y3919 = 1'b0 ;
  assign y3920 = n5248 ;
  assign y3921 = 1'b0 ;
  assign y3922 = ~1'b0 ;
  assign y3923 = ~1'b0 ;
  assign y3924 = n5252 ;
  assign y3925 = ~n5256 ;
  assign y3926 = n5258 ;
  assign y3927 = ~n5265 ;
  assign y3928 = ~n5267 ;
  assign y3929 = ~1'b0 ;
  assign y3930 = ~n5269 ;
  assign y3931 = 1'b0 ;
  assign y3932 = ~n5270 ;
  assign y3933 = n5275 ;
  assign y3934 = ~1'b0 ;
  assign y3935 = ~n3640 ;
  assign y3936 = ~1'b0 ;
  assign y3937 = ~n5277 ;
  assign y3938 = ~n5278 ;
  assign y3939 = ~1'b0 ;
  assign y3940 = n5280 ;
  assign y3941 = ~1'b0 ;
  assign y3942 = n5282 ;
  assign y3943 = ~n1714 ;
  assign y3944 = ~n5283 ;
  assign y3945 = ~1'b0 ;
  assign y3946 = ~1'b0 ;
  assign y3947 = n5284 ;
  assign y3948 = ~n5287 ;
  assign y3949 = ~n5289 ;
  assign y3950 = 1'b0 ;
  assign y3951 = n5290 ;
  assign y3952 = 1'b0 ;
  assign y3953 = ~n5293 ;
  assign y3954 = ~1'b0 ;
  assign y3955 = ~1'b0 ;
  assign y3956 = n5294 ;
  assign y3957 = n899 ;
  assign y3958 = n5295 ;
  assign y3959 = n5297 ;
  assign y3960 = 1'b0 ;
  assign y3961 = ~n5302 ;
  assign y3962 = ~1'b0 ;
  assign y3963 = ~1'b0 ;
  assign y3964 = n5309 ;
  assign y3965 = ~n5312 ;
  assign y3966 = n5316 ;
  assign y3967 = ~n1951 ;
  assign y3968 = n5319 ;
  assign y3969 = ~n5321 ;
  assign y3970 = ~1'b0 ;
  assign y3971 = ~n5323 ;
  assign y3972 = n5324 ;
  assign y3973 = n5325 ;
  assign y3974 = ~1'b0 ;
  assign y3975 = ~n5327 ;
  assign y3976 = ~1'b0 ;
  assign y3977 = ~n5328 ;
  assign y3978 = ~1'b0 ;
  assign y3979 = ~1'b0 ;
  assign y3980 = ~1'b0 ;
  assign y3981 = ~1'b0 ;
  assign y3982 = ~n5330 ;
  assign y3983 = ~n5331 ;
  assign y3984 = n1856 ;
  assign y3985 = n5332 ;
  assign y3986 = ~1'b0 ;
  assign y3987 = ~n5334 ;
  assign y3988 = n5335 ;
  assign y3989 = ~1'b0 ;
  assign y3990 = ~n5336 ;
  assign y3991 = ~1'b0 ;
  assign y3992 = ~1'b0 ;
  assign y3993 = n5344 ;
  assign y3994 = ~1'b0 ;
  assign y3995 = ~1'b0 ;
  assign y3996 = n5345 ;
  assign y3997 = ~1'b0 ;
  assign y3998 = n5347 ;
  assign y3999 = ~1'b0 ;
  assign y4000 = n4419 ;
  assign y4001 = n5348 ;
  assign y4002 = ~1'b0 ;
  assign y4003 = n5350 ;
  assign y4004 = ~n5357 ;
  assign y4005 = ~1'b0 ;
  assign y4006 = ~1'b0 ;
  assign y4007 = ~1'b0 ;
  assign y4008 = 1'b0 ;
  assign y4009 = n5358 ;
  assign y4010 = n2849 ;
  assign y4011 = ~n5360 ;
  assign y4012 = n3584 ;
  assign y4013 = ~1'b0 ;
  assign y4014 = ~1'b0 ;
  assign y4015 = n5361 ;
  assign y4016 = n5366 ;
  assign y4017 = n5367 ;
  assign y4018 = n5368 ;
  assign y4019 = n5370 ;
  assign y4020 = 1'b0 ;
  assign y4021 = ~1'b0 ;
  assign y4022 = ~n5372 ;
  assign y4023 = n5373 ;
  assign y4024 = ~1'b0 ;
  assign y4025 = ~1'b0 ;
  assign y4026 = ~1'b0 ;
  assign y4027 = ~n982 ;
  assign y4028 = ~n5377 ;
  assign y4029 = n5383 ;
  assign y4030 = ~1'b0 ;
  assign y4031 = ~1'b0 ;
  assign y4032 = ~1'b0 ;
  assign y4033 = ~1'b0 ;
  assign y4034 = ~n5385 ;
  assign y4035 = ~n5386 ;
  assign y4036 = 1'b0 ;
  assign y4037 = n5387 ;
  assign y4038 = ~n3742 ;
  assign y4039 = n5391 ;
  assign y4040 = ~1'b0 ;
  assign y4041 = n5397 ;
  assign y4042 = ~n5399 ;
  assign y4043 = ~n5401 ;
  assign y4044 = ~1'b0 ;
  assign y4045 = n5402 ;
  assign y4046 = n5404 ;
  assign y4047 = 1'b0 ;
  assign y4048 = ~n5408 ;
  assign y4049 = ~1'b0 ;
  assign y4050 = n5413 ;
  assign y4051 = ~n5416 ;
  assign y4052 = ~n5418 ;
  assign y4053 = ~1'b0 ;
  assign y4054 = ~n5419 ;
  assign y4055 = ~1'b0 ;
  assign y4056 = ~n2909 ;
  assign y4057 = n73 ;
  assign y4058 = ~1'b0 ;
  assign y4059 = n5420 ;
  assign y4060 = ~n5421 ;
  assign y4061 = ~1'b0 ;
  assign y4062 = n5424 ;
  assign y4063 = ~1'b0 ;
  assign y4064 = ~1'b0 ;
  assign y4065 = ~1'b0 ;
  assign y4066 = ~1'b0 ;
  assign y4067 = ~1'b0 ;
  assign y4068 = ~n5427 ;
  assign y4069 = ~n5433 ;
  assign y4070 = ~n5437 ;
  assign y4071 = ~1'b0 ;
  assign y4072 = n5439 ;
  assign y4073 = ~n5442 ;
  assign y4074 = n5443 ;
  assign y4075 = ~n5444 ;
  assign y4076 = ~1'b0 ;
  assign y4077 = n5451 ;
  assign y4078 = ~1'b0 ;
  assign y4079 = ~1'b0 ;
  assign y4080 = ~n5455 ;
  assign y4081 = n5458 ;
  assign y4082 = ~1'b0 ;
  assign y4083 = n4093 ;
  assign y4084 = ~1'b0 ;
  assign y4085 = ~n5463 ;
  assign y4086 = n3019 ;
  assign y4087 = ~1'b0 ;
  assign y4088 = ~1'b0 ;
  assign y4089 = 1'b0 ;
  assign y4090 = ~n5465 ;
  assign y4091 = n5466 ;
  assign y4092 = ~n5469 ;
  assign y4093 = n2176 ;
  assign y4094 = ~n5470 ;
  assign y4095 = ~n5471 ;
  assign y4096 = ~n5473 ;
  assign y4097 = ~n5492 ;
  assign y4098 = ~n5493 ;
  assign y4099 = n5501 ;
  assign y4100 = ~1'b0 ;
  assign y4101 = ~n5505 ;
  assign y4102 = n3988 ;
  assign y4103 = ~1'b0 ;
  assign y4104 = ~n5513 ;
  assign y4105 = ~n5514 ;
  assign y4106 = ~1'b0 ;
  assign y4107 = ~1'b0 ;
  assign y4108 = n5517 ;
  assign y4109 = n5520 ;
  assign y4110 = ~1'b0 ;
  assign y4111 = ~n5524 ;
  assign y4112 = n5527 ;
  assign y4113 = n5529 ;
  assign y4114 = ~1'b0 ;
  assign y4115 = ~1'b0 ;
  assign y4116 = n5532 ;
  assign y4117 = ~n5535 ;
  assign y4118 = n688 ;
  assign y4119 = ~1'b0 ;
  assign y4120 = n5539 ;
  assign y4121 = ~1'b0 ;
  assign y4122 = ~1'b0 ;
  assign y4123 = n5541 ;
  assign y4124 = ~1'b0 ;
  assign y4125 = ~n5543 ;
  assign y4126 = n653 ;
  assign y4127 = ~1'b0 ;
  assign y4128 = ~1'b0 ;
  assign y4129 = n5544 ;
  assign y4130 = ~1'b0 ;
  assign y4131 = ~n5550 ;
  assign y4132 = n5554 ;
  assign y4133 = ~n5555 ;
  assign y4134 = ~1'b0 ;
  assign y4135 = n5557 ;
  assign y4136 = ~n5559 ;
  assign y4137 = n5560 ;
  assign y4138 = ~n5561 ;
  assign y4139 = ~1'b0 ;
  assign y4140 = n5564 ;
  assign y4141 = ~n5566 ;
  assign y4142 = n3767 ;
  assign y4143 = ~n5570 ;
  assign y4144 = ~n5571 ;
  assign y4145 = ~n5573 ;
  assign y4146 = ~1'b0 ;
  assign y4147 = 1'b0 ;
  assign y4148 = n5579 ;
  assign y4149 = ~n5586 ;
  assign y4150 = ~n5590 ;
  assign y4151 = ~n5601 ;
  assign y4152 = n5605 ;
  assign y4153 = ~1'b0 ;
  assign y4154 = ~n5606 ;
  assign y4155 = n5610 ;
  assign y4156 = ~1'b0 ;
  assign y4157 = ~1'b0 ;
  assign y4158 = n4531 ;
  assign y4159 = ~1'b0 ;
  assign y4160 = ~n5612 ;
  assign y4161 = ~1'b0 ;
  assign y4162 = ~1'b0 ;
  assign y4163 = ~1'b0 ;
  assign y4164 = 1'b0 ;
  assign y4165 = n5615 ;
  assign y4166 = ~1'b0 ;
  assign y4167 = ~1'b0 ;
  assign y4168 = n5617 ;
  assign y4169 = ~1'b0 ;
  assign y4170 = n4668 ;
  assign y4171 = ~n5622 ;
  assign y4172 = n5623 ;
  assign y4173 = ~n1800 ;
  assign y4174 = 1'b0 ;
  assign y4175 = ~n4169 ;
  assign y4176 = ~n5624 ;
  assign y4177 = n5628 ;
  assign y4178 = ~n395 ;
  assign y4179 = ~n5630 ;
  assign y4180 = ~n5638 ;
  assign y4181 = ~n234 ;
  assign y4182 = n5639 ;
  assign y4183 = ~n5643 ;
  assign y4184 = ~1'b0 ;
  assign y4185 = ~1'b0 ;
  assign y4186 = ~1'b0 ;
  assign y4187 = n5649 ;
  assign y4188 = ~1'b0 ;
  assign y4189 = ~n5652 ;
  assign y4190 = n861 ;
  assign y4191 = ~n5657 ;
  assign y4192 = ~n5659 ;
  assign y4193 = ~1'b0 ;
  assign y4194 = ~n5660 ;
  assign y4195 = ~1'b0 ;
  assign y4196 = ~n5663 ;
  assign y4197 = ~n5665 ;
  assign y4198 = ~1'b0 ;
  assign y4199 = n5668 ;
  assign y4200 = ~n5677 ;
  assign y4201 = 1'b0 ;
  assign y4202 = ~1'b0 ;
  assign y4203 = ~n5681 ;
  assign y4204 = 1'b0 ;
  assign y4205 = ~n5684 ;
  assign y4206 = ~n1438 ;
  assign y4207 = n5690 ;
  assign y4208 = n5694 ;
  assign y4209 = ~n2124 ;
  assign y4210 = n5696 ;
  assign y4211 = ~1'b0 ;
  assign y4212 = n5698 ;
  assign y4213 = ~1'b0 ;
  assign y4214 = ~1'b0 ;
  assign y4215 = n5700 ;
  assign y4216 = n5704 ;
  assign y4217 = 1'b0 ;
  assign y4218 = ~1'b0 ;
  assign y4219 = n5707 ;
  assign y4220 = n5708 ;
  assign y4221 = n5711 ;
  assign y4222 = ~1'b0 ;
  assign y4223 = n5713 ;
  assign y4224 = ~1'b0 ;
  assign y4225 = ~1'b0 ;
  assign y4226 = ~n5205 ;
  assign y4227 = n4969 ;
  assign y4228 = ~n5714 ;
  assign y4229 = n5716 ;
  assign y4230 = ~1'b0 ;
  assign y4231 = ~1'b0 ;
  assign y4232 = n5719 ;
  assign y4233 = n5720 ;
  assign y4234 = ~1'b0 ;
  assign y4235 = ~1'b0 ;
  assign y4236 = n5721 ;
  assign y4237 = n5722 ;
  assign y4238 = n5725 ;
  assign y4239 = n5726 ;
  assign y4240 = n5729 ;
  assign y4241 = ~n5730 ;
  assign y4242 = n5736 ;
  assign y4243 = n5428 ;
  assign y4244 = ~1'b0 ;
  assign y4245 = ~1'b0 ;
  assign y4246 = ~1'b0 ;
  assign y4247 = ~1'b0 ;
  assign y4248 = ~1'b0 ;
  assign y4249 = ~n5740 ;
  assign y4250 = ~n5746 ;
  assign y4251 = n5747 ;
  assign y4252 = n1219 ;
  assign y4253 = n5752 ;
  assign y4254 = ~1'b0 ;
  assign y4255 = ~n5753 ;
  assign y4256 = ~n5754 ;
  assign y4257 = ~1'b0 ;
  assign y4258 = n3773 ;
  assign y4259 = ~n5755 ;
  assign y4260 = ~1'b0 ;
  assign y4261 = ~1'b0 ;
  assign y4262 = ~1'b0 ;
  assign y4263 = n5758 ;
  assign y4264 = n5761 ;
  assign y4265 = n5768 ;
  assign y4266 = n5771 ;
  assign y4267 = n5772 ;
  assign y4268 = ~n5774 ;
  assign y4269 = ~1'b0 ;
  assign y4270 = 1'b0 ;
  assign y4271 = ~n5778 ;
  assign y4272 = ~1'b0 ;
  assign y4273 = 1'b0 ;
  assign y4274 = n5782 ;
  assign y4275 = 1'b0 ;
  assign y4276 = ~1'b0 ;
  assign y4277 = ~n5783 ;
  assign y4278 = n5784 ;
  assign y4279 = n5785 ;
  assign y4280 = ~1'b0 ;
  assign y4281 = ~n1304 ;
  assign y4282 = n5788 ;
  assign y4283 = ~1'b0 ;
  assign y4284 = ~1'b0 ;
  assign y4285 = ~n5792 ;
  assign y4286 = ~n2769 ;
  assign y4287 = ~n5793 ;
  assign y4288 = ~1'b0 ;
  assign y4289 = n5795 ;
  assign y4290 = ~n5797 ;
  assign y4291 = n5798 ;
  assign y4292 = ~1'b0 ;
  assign y4293 = ~1'b0 ;
  assign y4294 = 1'b0 ;
  assign y4295 = 1'b0 ;
  assign y4296 = 1'b0 ;
  assign y4297 = ~n5800 ;
  assign y4298 = ~1'b0 ;
  assign y4299 = ~n5808 ;
  assign y4300 = n5809 ;
  assign y4301 = ~n5812 ;
  assign y4302 = n2075 ;
  assign y4303 = n5813 ;
  assign y4304 = ~n5817 ;
  assign y4305 = n5818 ;
  assign y4306 = ~n5819 ;
  assign y4307 = ~1'b0 ;
  assign y4308 = ~n5820 ;
  assign y4309 = ~n5821 ;
  assign y4310 = ~1'b0 ;
  assign y4311 = ~n5825 ;
  assign y4312 = n5826 ;
  assign y4313 = ~1'b0 ;
  assign y4314 = ~n5828 ;
  assign y4315 = ~n5831 ;
  assign y4316 = ~n5832 ;
  assign y4317 = ~n5835 ;
  assign y4318 = ~n5629 ;
  assign y4319 = ~n5836 ;
  assign y4320 = ~1'b0 ;
  assign y4321 = ~1'b0 ;
  assign y4322 = ~1'b0 ;
  assign y4323 = ~1'b0 ;
  assign y4324 = ~1'b0 ;
  assign y4325 = ~n5841 ;
  assign y4326 = ~1'b0 ;
  assign y4327 = ~1'b0 ;
  assign y4328 = ~1'b0 ;
  assign y4329 = n5842 ;
  assign y4330 = n3249 ;
  assign y4331 = n653 ;
  assign y4332 = ~1'b0 ;
  assign y4333 = n5849 ;
  assign y4334 = ~n5850 ;
  assign y4335 = ~n5851 ;
  assign y4336 = ~n5854 ;
  assign y4337 = 1'b0 ;
  assign y4338 = ~n5860 ;
  assign y4339 = n5862 ;
  assign y4340 = 1'b0 ;
  assign y4341 = 1'b0 ;
  assign y4342 = ~n5863 ;
  assign y4343 = ~1'b0 ;
  assign y4344 = ~1'b0 ;
  assign y4345 = n5864 ;
  assign y4346 = n5868 ;
  assign y4347 = ~n5871 ;
  assign y4348 = ~n5873 ;
  assign y4349 = n5877 ;
  assign y4350 = n5880 ;
  assign y4351 = ~1'b0 ;
  assign y4352 = ~1'b0 ;
  assign y4353 = ~1'b0 ;
  assign y4354 = ~1'b0 ;
  assign y4355 = ~1'b0 ;
  assign y4356 = ~n5885 ;
  assign y4357 = ~n294 ;
  assign y4358 = ~1'b0 ;
  assign y4359 = n3037 ;
  assign y4360 = 1'b0 ;
  assign y4361 = n5889 ;
  assign y4362 = ~1'b0 ;
  assign y4363 = 1'b0 ;
  assign y4364 = ~n5890 ;
  assign y4365 = n5895 ;
  assign y4366 = n5899 ;
  assign y4367 = ~n5900 ;
  assign y4368 = n832 ;
  assign y4369 = ~n3405 ;
  assign y4370 = ~n4677 ;
  assign y4371 = ~n5902 ;
  assign y4372 = n2724 ;
  assign y4373 = ~1'b0 ;
  assign y4374 = ~n5903 ;
  assign y4375 = n5905 ;
  assign y4376 = ~1'b0 ;
  assign y4377 = n83 ;
  assign y4378 = n5907 ;
  assign y4379 = ~1'b0 ;
  assign y4380 = ~n5909 ;
  assign y4381 = n5910 ;
  assign y4382 = n5912 ;
  assign y4383 = ~1'b0 ;
  assign y4384 = n5914 ;
  assign y4385 = n5915 ;
  assign y4386 = ~n4533 ;
  assign y4387 = ~n5917 ;
  assign y4388 = ~1'b0 ;
  assign y4389 = n5920 ;
  assign y4390 = n618 ;
  assign y4391 = ~n5922 ;
  assign y4392 = 1'b0 ;
  assign y4393 = ~1'b0 ;
  assign y4394 = ~1'b0 ;
  assign y4395 = ~1'b0 ;
  assign y4396 = ~n5923 ;
  assign y4397 = 1'b0 ;
  assign y4398 = n5924 ;
  assign y4399 = ~1'b0 ;
  assign y4400 = ~1'b0 ;
  assign y4401 = ~n5929 ;
  assign y4402 = ~n2846 ;
  assign y4403 = ~n5936 ;
  assign y4404 = ~n5939 ;
  assign y4405 = ~1'b0 ;
  assign y4406 = ~n5942 ;
  assign y4407 = ~1'b0 ;
  assign y4408 = n5945 ;
  assign y4409 = n5947 ;
  assign y4410 = 1'b0 ;
  assign y4411 = n5948 ;
  assign y4412 = 1'b0 ;
  assign y4413 = ~n2303 ;
  assign y4414 = ~1'b0 ;
  assign y4415 = n5949 ;
  assign y4416 = ~n5952 ;
  assign y4417 = ~n5953 ;
  assign y4418 = ~1'b0 ;
  assign y4419 = ~n5955 ;
  assign y4420 = ~1'b0 ;
  assign y4421 = n5956 ;
  assign y4422 = ~1'b0 ;
  assign y4423 = 1'b0 ;
  assign y4424 = ~1'b0 ;
  assign y4425 = ~n5957 ;
  assign y4426 = ~n1718 ;
  assign y4427 = n5958 ;
  assign y4428 = ~1'b0 ;
  assign y4429 = n5961 ;
  assign y4430 = ~1'b0 ;
  assign y4431 = ~1'b0 ;
  assign y4432 = n532 ;
  assign y4433 = ~1'b0 ;
  assign y4434 = n5967 ;
  assign y4435 = ~1'b0 ;
  assign y4436 = ~1'b0 ;
  assign y4437 = ~1'b0 ;
  assign y4438 = ~1'b0 ;
  assign y4439 = ~1'b0 ;
  assign y4440 = ~1'b0 ;
  assign y4441 = n5970 ;
  assign y4442 = ~n3995 ;
  assign y4443 = ~1'b0 ;
  assign y4444 = ~1'b0 ;
  assign y4445 = n5971 ;
  assign y4446 = ~1'b0 ;
  assign y4447 = ~n5972 ;
  assign y4448 = ~n5974 ;
  assign y4449 = ~n5975 ;
  assign y4450 = ~n2163 ;
  assign y4451 = ~n5979 ;
  assign y4452 = ~n178 ;
  assign y4453 = ~n5981 ;
  assign y4454 = ~n5982 ;
  assign y4455 = ~1'b0 ;
  assign y4456 = n5986 ;
  assign y4457 = ~n5989 ;
  assign y4458 = n30 ;
  assign y4459 = n1771 ;
  assign y4460 = ~1'b0 ;
  assign y4461 = n5990 ;
  assign y4462 = ~1'b0 ;
  assign y4463 = ~n5994 ;
  assign y4464 = n5995 ;
  assign y4465 = ~n5996 ;
  assign y4466 = ~n5998 ;
  assign y4467 = n5999 ;
  assign y4468 = ~1'b0 ;
  assign y4469 = n6003 ;
  assign y4470 = ~1'b0 ;
  assign y4471 = 1'b0 ;
  assign y4472 = n6005 ;
  assign y4473 = ~1'b0 ;
  assign y4474 = ~n6006 ;
  assign y4475 = n6009 ;
  assign y4476 = n6010 ;
  assign y4477 = ~1'b0 ;
  assign y4478 = ~1'b0 ;
  assign y4479 = ~n6015 ;
  assign y4480 = ~1'b0 ;
  assign y4481 = ~n6016 ;
  assign y4482 = ~1'b0 ;
  assign y4483 = n6019 ;
  assign y4484 = ~n6021 ;
  assign y4485 = ~n6022 ;
  assign y4486 = ~n6025 ;
  assign y4487 = ~1'b0 ;
  assign y4488 = n6026 ;
  assign y4489 = ~n6027 ;
  assign y4490 = n4155 ;
  assign y4491 = ~n6028 ;
  assign y4492 = ~1'b0 ;
  assign y4493 = ~n6031 ;
  assign y4494 = ~n6033 ;
  assign y4495 = ~n6036 ;
  assign y4496 = ~n6039 ;
  assign y4497 = ~1'b0 ;
  assign y4498 = ~n6040 ;
  assign y4499 = n5412 ;
  assign y4500 = 1'b0 ;
  assign y4501 = ~1'b0 ;
  assign y4502 = ~1'b0 ;
  assign y4503 = ~1'b0 ;
  assign y4504 = ~n6041 ;
  assign y4505 = 1'b0 ;
  assign y4506 = ~1'b0 ;
  assign y4507 = n6043 ;
  assign y4508 = ~1'b0 ;
  assign y4509 = ~1'b0 ;
  assign y4510 = n6046 ;
  assign y4511 = ~1'b0 ;
  assign y4512 = n6048 ;
  assign y4513 = ~1'b0 ;
  assign y4514 = ~n6049 ;
  assign y4515 = ~1'b0 ;
  assign y4516 = ~1'b0 ;
  assign y4517 = n6050 ;
  assign y4518 = n6051 ;
  assign y4519 = ~1'b0 ;
  assign y4520 = n6057 ;
  assign y4521 = ~1'b0 ;
  assign y4522 = 1'b0 ;
  assign y4523 = ~1'b0 ;
  assign y4524 = n6060 ;
  assign y4525 = n6061 ;
  assign y4526 = ~n6068 ;
  assign y4527 = ~1'b0 ;
  assign y4528 = ~n6070 ;
  assign y4529 = ~n6071 ;
  assign y4530 = n5905 ;
  assign y4531 = ~1'b0 ;
  assign y4532 = ~n1947 ;
  assign y4533 = ~1'b0 ;
  assign y4534 = n6077 ;
  assign y4535 = 1'b0 ;
  assign y4536 = ~1'b0 ;
  assign y4537 = ~n6080 ;
  assign y4538 = ~1'b0 ;
  assign y4539 = n6082 ;
  assign y4540 = n6084 ;
  assign y4541 = ~n6087 ;
  assign y4542 = n6094 ;
  assign y4543 = n6095 ;
  assign y4544 = ~n6096 ;
  assign y4545 = n6099 ;
  assign y4546 = ~1'b0 ;
  assign y4547 = ~1'b0 ;
  assign y4548 = n6104 ;
  assign y4549 = n622 ;
  assign y4550 = ~1'b0 ;
  assign y4551 = ~1'b0 ;
  assign y4552 = ~1'b0 ;
  assign y4553 = ~n5434 ;
  assign y4554 = n6109 ;
  assign y4555 = ~1'b0 ;
  assign y4556 = ~1'b0 ;
  assign y4557 = ~1'b0 ;
  assign y4558 = n5364 ;
  assign y4559 = ~n6111 ;
  assign y4560 = ~n6117 ;
  assign y4561 = ~n6128 ;
  assign y4562 = ~n6131 ;
  assign y4563 = ~n6134 ;
  assign y4564 = ~1'b0 ;
  assign y4565 = n6135 ;
  assign y4566 = n2063 ;
  assign y4567 = ~1'b0 ;
  assign y4568 = n2463 ;
  assign y4569 = ~n6139 ;
  assign y4570 = ~n1245 ;
  assign y4571 = ~1'b0 ;
  assign y4572 = n6143 ;
  assign y4573 = n6144 ;
  assign y4574 = n6145 ;
  assign y4575 = n3267 ;
  assign y4576 = ~1'b0 ;
  assign y4577 = ~n6146 ;
  assign y4578 = n6148 ;
  assign y4579 = n6149 ;
  assign y4580 = ~n6151 ;
  assign y4581 = ~n2239 ;
  assign y4582 = n6159 ;
  assign y4583 = n5533 ;
  assign y4584 = ~1'b0 ;
  assign y4585 = ~1'b0 ;
  assign y4586 = n6162 ;
  assign y4587 = n6166 ;
  assign y4588 = ~n6167 ;
  assign y4589 = n6169 ;
  assign y4590 = ~n6172 ;
  assign y4591 = ~n6173 ;
  assign y4592 = n6176 ;
  assign y4593 = ~n5454 ;
  assign y4594 = ~1'b0 ;
  assign y4595 = ~1'b0 ;
  assign y4596 = ~1'b0 ;
  assign y4597 = ~1'b0 ;
  assign y4598 = n880 ;
  assign y4599 = n6179 ;
  assign y4600 = ~n6182 ;
  assign y4601 = n6186 ;
  assign y4602 = ~n6187 ;
  assign y4603 = n6189 ;
  assign y4604 = 1'b0 ;
  assign y4605 = n6190 ;
  assign y4606 = ~n6196 ;
  assign y4607 = ~n6197 ;
  assign y4608 = ~1'b0 ;
  assign y4609 = ~n2819 ;
  assign y4610 = n163 ;
  assign y4611 = ~n6198 ;
  assign y4612 = ~n6204 ;
  assign y4613 = ~n6206 ;
  assign y4614 = ~n6209 ;
  assign y4615 = ~n6211 ;
  assign y4616 = ~n3533 ;
  assign y4617 = ~1'b0 ;
  assign y4618 = ~n553 ;
  assign y4619 = ~1'b0 ;
  assign y4620 = ~n6213 ;
  assign y4621 = ~n6218 ;
  assign y4622 = n6222 ;
  assign y4623 = ~n6224 ;
  assign y4624 = 1'b0 ;
  assign y4625 = n6225 ;
  assign y4626 = ~1'b0 ;
  assign y4627 = ~1'b0 ;
  assign y4628 = ~n6226 ;
  assign y4629 = ~1'b0 ;
  assign y4630 = ~n6228 ;
  assign y4631 = ~1'b0 ;
  assign y4632 = n6234 ;
  assign y4633 = ~1'b0 ;
  assign y4634 = n6235 ;
  assign y4635 = ~n6236 ;
  assign y4636 = ~n6238 ;
  assign y4637 = n6240 ;
  assign y4638 = ~n5076 ;
  assign y4639 = ~1'b0 ;
  assign y4640 = ~1'b0 ;
  assign y4641 = ~1'b0 ;
  assign y4642 = ~1'b0 ;
  assign y4643 = n6245 ;
  assign y4644 = ~1'b0 ;
  assign y4645 = ~1'b0 ;
  assign y4646 = 1'b0 ;
  assign y4647 = n310 ;
  assign y4648 = n6249 ;
  assign y4649 = n6253 ;
  assign y4650 = ~n6256 ;
  assign y4651 = ~n6258 ;
  assign y4652 = 1'b0 ;
  assign y4653 = n6263 ;
  assign y4654 = ~1'b0 ;
  assign y4655 = n6270 ;
  assign y4656 = n6272 ;
  assign y4657 = ~1'b0 ;
  assign y4658 = 1'b0 ;
  assign y4659 = ~1'b0 ;
  assign y4660 = n570 ;
  assign y4661 = ~1'b0 ;
  assign y4662 = ~n6274 ;
  assign y4663 = ~n6278 ;
  assign y4664 = ~n6279 ;
  assign y4665 = ~n6281 ;
  assign y4666 = ~n6285 ;
  assign y4667 = n3542 ;
  assign y4668 = ~n6286 ;
  assign y4669 = ~1'b0 ;
  assign y4670 = n1924 ;
  assign y4671 = n6287 ;
  assign y4672 = n6289 ;
  assign y4673 = n6290 ;
  assign y4674 = n6291 ;
  assign y4675 = n6292 ;
  assign y4676 = ~n6295 ;
  assign y4677 = ~1'b0 ;
  assign y4678 = ~1'b0 ;
  assign y4679 = ~1'b0 ;
  assign y4680 = ~1'b0 ;
  assign y4681 = ~1'b0 ;
  assign y4682 = n6298 ;
  assign y4683 = ~1'b0 ;
  assign y4684 = ~1'b0 ;
  assign y4685 = ~1'b0 ;
  assign y4686 = ~n3527 ;
  assign y4687 = ~n6300 ;
  assign y4688 = ~n6301 ;
  assign y4689 = ~1'b0 ;
  assign y4690 = n6303 ;
  assign y4691 = n1080 ;
  assign y4692 = ~1'b0 ;
  assign y4693 = ~1'b0 ;
  assign y4694 = ~n6304 ;
  assign y4695 = n6308 ;
  assign y4696 = ~1'b0 ;
  assign y4697 = n6313 ;
  assign y4698 = n6315 ;
  assign y4699 = ~1'b0 ;
  assign y4700 = ~1'b0 ;
  assign y4701 = ~n5981 ;
  assign y4702 = ~1'b0 ;
  assign y4703 = n6318 ;
  assign y4704 = ~n6321 ;
  assign y4705 = n6322 ;
  assign y4706 = ~n6323 ;
  assign y4707 = ~n6327 ;
  assign y4708 = ~n4784 ;
  assign y4709 = ~1'b0 ;
  assign y4710 = ~1'b0 ;
  assign y4711 = ~1'b0 ;
  assign y4712 = ~n6332 ;
  assign y4713 = n6336 ;
  assign y4714 = ~1'b0 ;
  assign y4715 = n6337 ;
  assign y4716 = ~1'b0 ;
  assign y4717 = ~1'b0 ;
  assign y4718 = ~1'b0 ;
  assign y4719 = ~n6338 ;
  assign y4720 = ~n6339 ;
  assign y4721 = ~1'b0 ;
  assign y4722 = n6340 ;
  assign y4723 = ~1'b0 ;
  assign y4724 = ~n6345 ;
  assign y4725 = ~1'b0 ;
  assign y4726 = ~1'b0 ;
  assign y4727 = ~n6351 ;
  assign y4728 = ~n6355 ;
  assign y4729 = ~1'b0 ;
  assign y4730 = n6357 ;
  assign y4731 = ~1'b0 ;
  assign y4732 = 1'b0 ;
  assign y4733 = ~n6359 ;
  assign y4734 = ~n4365 ;
  assign y4735 = ~n6363 ;
  assign y4736 = n6365 ;
  assign y4737 = n6366 ;
  assign y4738 = ~n6373 ;
  assign y4739 = ~1'b0 ;
  assign y4740 = ~n6375 ;
  assign y4741 = ~1'b0 ;
  assign y4742 = n6376 ;
  assign y4743 = ~1'b0 ;
  assign y4744 = ~1'b0 ;
  assign y4745 = ~1'b0 ;
  assign y4746 = n6377 ;
  assign y4747 = ~1'b0 ;
  assign y4748 = ~1'b0 ;
  assign y4749 = ~1'b0 ;
  assign y4750 = ~n6378 ;
  assign y4751 = n6379 ;
  assign y4752 = ~1'b0 ;
  assign y4753 = 1'b0 ;
  assign y4754 = 1'b0 ;
  assign y4755 = ~1'b0 ;
  assign y4756 = ~1'b0 ;
  assign y4757 = ~n6381 ;
  assign y4758 = ~n6384 ;
  assign y4759 = ~n3318 ;
  assign y4760 = ~1'b0 ;
  assign y4761 = n257 ;
  assign y4762 = ~1'b0 ;
  assign y4763 = ~n6387 ;
  assign y4764 = ~1'b0 ;
  assign y4765 = ~1'b0 ;
  assign y4766 = ~n6390 ;
  assign y4767 = ~1'b0 ;
  assign y4768 = ~n6392 ;
  assign y4769 = ~n6395 ;
  assign y4770 = ~1'b0 ;
  assign y4771 = ~1'b0 ;
  assign y4772 = ~1'b0 ;
  assign y4773 = n6401 ;
  assign y4774 = ~1'b0 ;
  assign y4775 = ~1'b0 ;
  assign y4776 = n6402 ;
  assign y4777 = ~1'b0 ;
  assign y4778 = n6403 ;
  assign y4779 = n6406 ;
  assign y4780 = ~1'b0 ;
  assign y4781 = ~n6407 ;
  assign y4782 = n6411 ;
  assign y4783 = ~1'b0 ;
  assign y4784 = 1'b0 ;
  assign y4785 = ~n2785 ;
  assign y4786 = ~n6412 ;
  assign y4787 = ~1'b0 ;
  assign y4788 = ~1'b0 ;
  assign y4789 = ~n6414 ;
  assign y4790 = ~n6419 ;
  assign y4791 = ~n3411 ;
  assign y4792 = ~n6420 ;
  assign y4793 = n6421 ;
  assign y4794 = ~n6422 ;
  assign y4795 = ~n6427 ;
  assign y4796 = ~1'b0 ;
  assign y4797 = ~1'b0 ;
  assign y4798 = ~n6429 ;
  assign y4799 = n6430 ;
  assign y4800 = ~n6433 ;
  assign y4801 = ~1'b0 ;
  assign y4802 = n6439 ;
  assign y4803 = ~1'b0 ;
  assign y4804 = ~n6440 ;
  assign y4805 = n6441 ;
  assign y4806 = ~n6443 ;
  assign y4807 = ~n5194 ;
  assign y4808 = ~1'b0 ;
  assign y4809 = n6444 ;
  assign y4810 = n6450 ;
  assign y4811 = ~1'b0 ;
  assign y4812 = n270 ;
  assign y4813 = ~1'b0 ;
  assign y4814 = n4448 ;
  assign y4815 = n6451 ;
  assign y4816 = ~n6454 ;
  assign y4817 = ~1'b0 ;
  assign y4818 = ~n6456 ;
  assign y4819 = ~n6459 ;
  assign y4820 = ~1'b0 ;
  assign y4821 = ~1'b0 ;
  assign y4822 = 1'b0 ;
  assign y4823 = ~n6461 ;
  assign y4824 = ~n274 ;
  assign y4825 = ~1'b0 ;
  assign y4826 = ~n6462 ;
  assign y4827 = 1'b0 ;
  assign y4828 = ~1'b0 ;
  assign y4829 = ~n6463 ;
  assign y4830 = ~1'b0 ;
  assign y4831 = ~1'b0 ;
  assign y4832 = ~n6469 ;
  assign y4833 = ~n246 ;
  assign y4834 = ~1'b0 ;
  assign y4835 = ~n6472 ;
  assign y4836 = n6476 ;
  assign y4837 = n6477 ;
  assign y4838 = ~n6479 ;
  assign y4839 = ~n6481 ;
  assign y4840 = ~1'b0 ;
  assign y4841 = ~n6482 ;
  assign y4842 = ~n6485 ;
  assign y4843 = ~1'b0 ;
  assign y4844 = ~1'b0 ;
  assign y4845 = n6486 ;
  assign y4846 = 1'b0 ;
  assign y4847 = n6488 ;
  assign y4848 = ~n6492 ;
  assign y4849 = ~n6502 ;
  assign y4850 = ~1'b0 ;
  assign y4851 = ~1'b0 ;
  assign y4852 = ~n6504 ;
  assign y4853 = n6508 ;
  assign y4854 = n1106 ;
  assign y4855 = ~n6509 ;
  assign y4856 = ~1'b0 ;
  assign y4857 = ~1'b0 ;
  assign y4858 = ~n6510 ;
  assign y4859 = ~n6514 ;
  assign y4860 = n6515 ;
  assign y4861 = ~n6518 ;
  assign y4862 = ~n6519 ;
  assign y4863 = ~n6523 ;
  assign y4864 = n6525 ;
  assign y4865 = 1'b0 ;
  assign y4866 = ~1'b0 ;
  assign y4867 = ~n6526 ;
  assign y4868 = ~n6529 ;
  assign y4869 = ~1'b0 ;
  assign y4870 = n6530 ;
  assign y4871 = ~n6531 ;
  assign y4872 = ~n1219 ;
  assign y4873 = ~1'b0 ;
  assign y4874 = ~1'b0 ;
  assign y4875 = ~n6533 ;
  assign y4876 = n6536 ;
  assign y4877 = n6537 ;
  assign y4878 = ~n1208 ;
  assign y4879 = 1'b0 ;
  assign y4880 = ~1'b0 ;
  assign y4881 = ~n1560 ;
  assign y4882 = ~1'b0 ;
  assign y4883 = ~n6539 ;
  assign y4884 = n1108 ;
  assign y4885 = n6540 ;
  assign y4886 = ~n142 ;
  assign y4887 = n6543 ;
  assign y4888 = n6546 ;
  assign y4889 = ~n6547 ;
  assign y4890 = ~1'b0 ;
  assign y4891 = n6551 ;
  assign y4892 = n6565 ;
  assign y4893 = ~n6566 ;
  assign y4894 = ~1'b0 ;
  assign y4895 = ~1'b0 ;
  assign y4896 = ~n6567 ;
  assign y4897 = ~1'b0 ;
  assign y4898 = n6569 ;
  assign y4899 = ~n6578 ;
  assign y4900 = ~1'b0 ;
  assign y4901 = ~1'b0 ;
  assign y4902 = ~n6583 ;
  assign y4903 = 1'b0 ;
  assign y4904 = ~n6584 ;
  assign y4905 = ~n6587 ;
  assign y4906 = ~1'b0 ;
  assign y4907 = 1'b0 ;
  assign y4908 = ~n153 ;
  assign y4909 = n6588 ;
  assign y4910 = ~n6592 ;
  assign y4911 = ~n6595 ;
  assign y4912 = ~1'b0 ;
  assign y4913 = ~n5317 ;
  assign y4914 = n6601 ;
  assign y4915 = ~n6605 ;
  assign y4916 = n1676 ;
  assign y4917 = n6607 ;
  assign y4918 = ~n6610 ;
  assign y4919 = n6616 ;
  assign y4920 = ~1'b0 ;
  assign y4921 = 1'b0 ;
  assign y4922 = ~n4660 ;
  assign y4923 = n6617 ;
  assign y4924 = ~n6619 ;
  assign y4925 = ~1'b0 ;
  assign y4926 = n6623 ;
  assign y4927 = ~1'b0 ;
  assign y4928 = ~1'b0 ;
  assign y4929 = ~n6627 ;
  assign y4930 = n6629 ;
  assign y4931 = ~n6640 ;
  assign y4932 = ~1'b0 ;
  assign y4933 = ~1'b0 ;
  assign y4934 = n6643 ;
  assign y4935 = n6644 ;
  assign y4936 = n2031 ;
  assign y4937 = n6646 ;
  assign y4938 = ~1'b0 ;
  assign y4939 = n865 ;
  assign y4940 = n6653 ;
  assign y4941 = ~n6656 ;
  assign y4942 = ~1'b0 ;
  assign y4943 = ~1'b0 ;
  assign y4944 = ~n6658 ;
  assign y4945 = ~1'b0 ;
  assign y4946 = ~n6660 ;
  assign y4947 = ~n3333 ;
  assign y4948 = ~1'b0 ;
  assign y4949 = n6663 ;
  assign y4950 = ~1'b0 ;
  assign y4951 = ~1'b0 ;
  assign y4952 = ~1'b0 ;
  assign y4953 = n6665 ;
  assign y4954 = n6667 ;
  assign y4955 = n6671 ;
  assign y4956 = ~n6672 ;
  assign y4957 = n6673 ;
  assign y4958 = ~1'b0 ;
  assign y4959 = n1789 ;
  assign y4960 = n6674 ;
  assign y4961 = ~1'b0 ;
  assign y4962 = n6676 ;
  assign y4963 = 1'b0 ;
  assign y4964 = ~n6677 ;
  assign y4965 = ~n6681 ;
  assign y4966 = n6682 ;
  assign y4967 = ~n6683 ;
  assign y4968 = n6687 ;
  assign y4969 = ~n6691 ;
  assign y4970 = n6697 ;
  assign y4971 = n6698 ;
  assign y4972 = ~1'b0 ;
  assign y4973 = n3512 ;
  assign y4974 = ~1'b0 ;
  assign y4975 = ~1'b0 ;
  assign y4976 = n6702 ;
  assign y4977 = ~n6705 ;
  assign y4978 = ~1'b0 ;
  assign y4979 = ~n6707 ;
  assign y4980 = ~n6710 ;
  assign y4981 = n6715 ;
  assign y4982 = n6719 ;
  assign y4983 = ~n6720 ;
  assign y4984 = n6723 ;
  assign y4985 = ~1'b0 ;
  assign y4986 = ~1'b0 ;
  assign y4987 = n6726 ;
  assign y4988 = ~n2107 ;
  assign y4989 = n6728 ;
  assign y4990 = n1052 ;
  assign y4991 = ~1'b0 ;
  assign y4992 = ~1'b0 ;
  assign y4993 = ~1'b0 ;
  assign y4994 = ~1'b0 ;
  assign y4995 = ~1'b0 ;
  assign y4996 = ~n6729 ;
  assign y4997 = ~1'b0 ;
  assign y4998 = n6732 ;
  assign y4999 = ~1'b0 ;
  assign y5000 = 1'b0 ;
  assign y5001 = ~1'b0 ;
  assign y5002 = n6734 ;
  assign y5003 = n6739 ;
  assign y5004 = ~1'b0 ;
  assign y5005 = ~1'b0 ;
  assign y5006 = ~n2107 ;
  assign y5007 = ~1'b0 ;
  assign y5008 = ~n6743 ;
  assign y5009 = ~n6749 ;
  assign y5010 = ~n6757 ;
  assign y5011 = n6762 ;
  assign y5012 = ~1'b0 ;
  assign y5013 = ~1'b0 ;
  assign y5014 = ~n6764 ;
  assign y5015 = ~n6766 ;
  assign y5016 = ~1'b0 ;
  assign y5017 = ~n6771 ;
  assign y5018 = ~n6772 ;
  assign y5019 = 1'b0 ;
  assign y5020 = n6773 ;
  assign y5021 = ~1'b0 ;
  assign y5022 = ~n467 ;
  assign y5023 = ~n6775 ;
  assign y5024 = ~1'b0 ;
  assign y5025 = ~1'b0 ;
  assign y5026 = ~1'b0 ;
  assign y5027 = ~n5626 ;
  assign y5028 = ~1'b0 ;
  assign y5029 = n6776 ;
  assign y5030 = ~n6780 ;
  assign y5031 = n6783 ;
  assign y5032 = ~1'b0 ;
  assign y5033 = ~1'b0 ;
  assign y5034 = ~n6784 ;
  assign y5035 = ~1'b0 ;
  assign y5036 = ~1'b0 ;
  assign y5037 = ~1'b0 ;
  assign y5038 = n6785 ;
  assign y5039 = ~n1388 ;
  assign y5040 = ~n6786 ;
  assign y5041 = n5733 ;
  assign y5042 = n6788 ;
  assign y5043 = ~n6789 ;
  assign y5044 = ~1'b0 ;
  assign y5045 = ~n6806 ;
  assign y5046 = ~1'b0 ;
  assign y5047 = ~n294 ;
  assign y5048 = n3589 ;
  assign y5049 = n6808 ;
  assign y5050 = n5794 ;
  assign y5051 = n322 ;
  assign y5052 = ~1'b0 ;
  assign y5053 = ~1'b0 ;
  assign y5054 = ~1'b0 ;
  assign y5055 = ~n6814 ;
  assign y5056 = ~1'b0 ;
  assign y5057 = ~n4883 ;
  assign y5058 = ~n6816 ;
  assign y5059 = ~n2835 ;
  assign y5060 = n6817 ;
  assign y5061 = ~n6823 ;
  assign y5062 = ~1'b0 ;
  assign y5063 = n6826 ;
  assign y5064 = ~1'b0 ;
  assign y5065 = ~1'b0 ;
  assign y5066 = n2435 ;
  assign y5067 = ~n4493 ;
  assign y5068 = 1'b0 ;
  assign y5069 = n6828 ;
  assign y5070 = n6834 ;
  assign y5071 = n6839 ;
  assign y5072 = ~n6843 ;
  assign y5073 = ~n6845 ;
  assign y5074 = ~1'b0 ;
  assign y5075 = 1'b0 ;
  assign y5076 = n6846 ;
  assign y5077 = 1'b0 ;
  assign y5078 = ~n6847 ;
  assign y5079 = ~n6853 ;
  assign y5080 = ~1'b0 ;
  assign y5081 = ~1'b0 ;
  assign y5082 = ~1'b0 ;
  assign y5083 = n6857 ;
  assign y5084 = ~n6860 ;
  assign y5085 = ~1'b0 ;
  assign y5086 = ~n6863 ;
  assign y5087 = ~1'b0 ;
  assign y5088 = ~n6870 ;
  assign y5089 = ~n6871 ;
  assign y5090 = ~n1229 ;
  assign y5091 = ~n6873 ;
  assign y5092 = n6875 ;
  assign y5093 = ~1'b0 ;
  assign y5094 = ~1'b0 ;
  assign y5095 = ~1'b0 ;
  assign y5096 = ~1'b0 ;
  assign y5097 = ~n6881 ;
  assign y5098 = n6884 ;
  assign y5099 = ~n6885 ;
  assign y5100 = ~n6886 ;
  assign y5101 = ~n6890 ;
  assign y5102 = ~1'b0 ;
  assign y5103 = ~1'b0 ;
  assign y5104 = ~1'b0 ;
  assign y5105 = ~n6892 ;
  assign y5106 = n6896 ;
  assign y5107 = ~1'b0 ;
  assign y5108 = ~1'b0 ;
  assign y5109 = ~1'b0 ;
  assign y5110 = ~n628 ;
  assign y5111 = ~1'b0 ;
  assign y5112 = ~1'b0 ;
  assign y5113 = ~1'b0 ;
  assign y5114 = n6899 ;
  assign y5115 = n6900 ;
  assign y5116 = ~n6901 ;
  assign y5117 = ~1'b0 ;
  assign y5118 = ~1'b0 ;
  assign y5119 = ~1'b0 ;
  assign y5120 = n6902 ;
  assign y5121 = n6904 ;
  assign y5122 = ~n1026 ;
  assign y5123 = ~n6911 ;
  assign y5124 = ~1'b0 ;
  assign y5125 = ~1'b0 ;
  assign y5126 = ~n6912 ;
  assign y5127 = ~1'b0 ;
  assign y5128 = ~n6915 ;
  assign y5129 = ~n6919 ;
  assign y5130 = ~1'b0 ;
  assign y5131 = n6920 ;
  assign y5132 = n6921 ;
  assign y5133 = ~1'b0 ;
  assign y5134 = n6922 ;
  assign y5135 = ~1'b0 ;
  assign y5136 = ~1'b0 ;
  assign y5137 = n6923 ;
  assign y5138 = 1'b0 ;
  assign y5139 = n4327 ;
  assign y5140 = ~1'b0 ;
  assign y5141 = ~n6924 ;
  assign y5142 = n6932 ;
  assign y5143 = 1'b0 ;
  assign y5144 = ~1'b0 ;
  assign y5145 = 1'b0 ;
  assign y5146 = ~1'b0 ;
  assign y5147 = n6933 ;
  assign y5148 = ~n6935 ;
  assign y5149 = ~n6937 ;
  assign y5150 = ~1'b0 ;
  assign y5151 = n6938 ;
  assign y5152 = n6939 ;
  assign y5153 = ~1'b0 ;
  assign y5154 = ~n1263 ;
  assign y5155 = ~1'b0 ;
  assign y5156 = ~1'b0 ;
  assign y5157 = ~1'b0 ;
  assign y5158 = ~n6940 ;
  assign y5159 = ~1'b0 ;
  assign y5160 = ~1'b0 ;
  assign y5161 = ~n6942 ;
  assign y5162 = ~n6948 ;
  assign y5163 = ~n6949 ;
  assign y5164 = n6955 ;
  assign y5165 = ~1'b0 ;
  assign y5166 = ~1'b0 ;
  assign y5167 = ~1'b0 ;
  assign y5168 = ~1'b0 ;
  assign y5169 = ~1'b0 ;
  assign y5170 = 1'b0 ;
  assign y5171 = n6957 ;
  assign y5172 = n6958 ;
  assign y5173 = n6965 ;
  assign y5174 = ~1'b0 ;
  assign y5175 = ~1'b0 ;
  assign y5176 = ~1'b0 ;
  assign y5177 = n6970 ;
  assign y5178 = ~n6971 ;
  assign y5179 = ~1'b0 ;
  assign y5180 = ~n6972 ;
  assign y5181 = n6973 ;
  assign y5182 = ~n6979 ;
  assign y5183 = ~1'b0 ;
  assign y5184 = n6983 ;
  assign y5185 = n6986 ;
  assign y5186 = ~n6998 ;
  assign y5187 = n7005 ;
  assign y5188 = ~n7006 ;
  assign y5189 = ~n7008 ;
  assign y5190 = n7013 ;
  assign y5191 = 1'b0 ;
  assign y5192 = n7021 ;
  assign y5193 = n7023 ;
  assign y5194 = ~1'b0 ;
  assign y5195 = ~1'b0 ;
  assign y5196 = ~n7024 ;
  assign y5197 = n7026 ;
  assign y5198 = 1'b0 ;
  assign y5199 = n7032 ;
  assign y5200 = n7033 ;
  assign y5201 = n7040 ;
  assign y5202 = n7041 ;
  assign y5203 = 1'b0 ;
  assign y5204 = n7046 ;
  assign y5205 = 1'b0 ;
  assign y5206 = ~1'b0 ;
  assign y5207 = ~1'b0 ;
  assign y5208 = n7047 ;
  assign y5209 = ~n7049 ;
  assign y5210 = ~n7051 ;
  assign y5211 = n7052 ;
  assign y5212 = n7053 ;
  assign y5213 = n7054 ;
  assign y5214 = n7055 ;
  assign y5215 = ~n7056 ;
  assign y5216 = ~1'b0 ;
  assign y5217 = ~n7057 ;
  assign y5218 = 1'b0 ;
  assign y5219 = ~1'b0 ;
  assign y5220 = ~1'b0 ;
  assign y5221 = ~1'b0 ;
  assign y5222 = ~n6989 ;
  assign y5223 = ~n5551 ;
  assign y5224 = n7063 ;
  assign y5225 = ~n7067 ;
  assign y5226 = ~n3951 ;
  assign y5227 = n5295 ;
  assign y5228 = ~n7070 ;
  assign y5229 = ~n7071 ;
  assign y5230 = ~n86 ;
  assign y5231 = ~1'b0 ;
  assign y5232 = 1'b0 ;
  assign y5233 = 1'b0 ;
  assign y5234 = ~n7072 ;
  assign y5235 = n7075 ;
  assign y5236 = n7077 ;
  assign y5237 = ~1'b0 ;
  assign y5238 = ~1'b0 ;
  assign y5239 = ~n7056 ;
  assign y5240 = ~n2546 ;
  assign y5241 = ~n7079 ;
  assign y5242 = n7080 ;
  assign y5243 = ~n7081 ;
  assign y5244 = ~n7082 ;
  assign y5245 = ~n7083 ;
  assign y5246 = 1'b0 ;
  assign y5247 = ~1'b0 ;
  assign y5248 = n7085 ;
  assign y5249 = ~n60 ;
  assign y5250 = ~n7090 ;
  assign y5251 = ~n7098 ;
  assign y5252 = ~n7100 ;
  assign y5253 = 1'b0 ;
  assign y5254 = ~1'b0 ;
  assign y5255 = n7101 ;
  assign y5256 = n7105 ;
  assign y5257 = ~n6361 ;
  assign y5258 = ~n2148 ;
  assign y5259 = ~n450 ;
  assign y5260 = n7108 ;
  assign y5261 = ~1'b0 ;
  assign y5262 = ~1'b0 ;
  assign y5263 = 1'b0 ;
  assign y5264 = ~1'b0 ;
  assign y5265 = n7109 ;
  assign y5266 = ~n7110 ;
  assign y5267 = 1'b0 ;
  assign y5268 = n7111 ;
  assign y5269 = ~n7113 ;
  assign y5270 = ~1'b0 ;
  assign y5271 = n7114 ;
  assign y5272 = n7115 ;
  assign y5273 = ~n7118 ;
  assign y5274 = ~1'b0 ;
  assign y5275 = ~1'b0 ;
  assign y5276 = ~n7119 ;
  assign y5277 = ~n7121 ;
  assign y5278 = n7122 ;
  assign y5279 = ~1'b0 ;
  assign y5280 = n7123 ;
  assign y5281 = n5726 ;
  assign y5282 = ~1'b0 ;
  assign y5283 = ~1'b0 ;
  assign y5284 = ~n7124 ;
  assign y5285 = n7130 ;
  assign y5286 = n4575 ;
  assign y5287 = ~n7132 ;
  assign y5288 = ~1'b0 ;
  assign y5289 = 1'b0 ;
  assign y5290 = 1'b0 ;
  assign y5291 = ~1'b0 ;
  assign y5292 = n7134 ;
  assign y5293 = ~1'b0 ;
  assign y5294 = ~1'b0 ;
  assign y5295 = ~1'b0 ;
  assign y5296 = ~1'b0 ;
  assign y5297 = ~n7135 ;
  assign y5298 = ~1'b0 ;
  assign y5299 = n7137 ;
  assign y5300 = ~n7139 ;
  assign y5301 = ~n7140 ;
  assign y5302 = n7143 ;
  assign y5303 = n7144 ;
  assign y5304 = n7145 ;
  assign y5305 = ~1'b0 ;
  assign y5306 = ~1'b0 ;
  assign y5307 = ~1'b0 ;
  assign y5308 = ~n7146 ;
  assign y5309 = ~1'b0 ;
  assign y5310 = ~n7147 ;
  assign y5311 = n7148 ;
  assign y5312 = ~1'b0 ;
  assign y5313 = ~1'b0 ;
  assign y5314 = ~1'b0 ;
  assign y5315 = ~n7149 ;
  assign y5316 = ~n7153 ;
  assign y5317 = ~n7154 ;
  assign y5318 = ~n7156 ;
  assign y5319 = n7159 ;
  assign y5320 = n7178 ;
  assign y5321 = ~n7180 ;
  assign y5322 = ~1'b0 ;
  assign y5323 = ~1'b0 ;
  assign y5324 = ~n7181 ;
  assign y5325 = ~1'b0 ;
  assign y5326 = n2692 ;
  assign y5327 = ~n7183 ;
  assign y5328 = ~1'b0 ;
  assign y5329 = ~1'b0 ;
  assign y5330 = ~1'b0 ;
  assign y5331 = ~n7185 ;
  assign y5332 = n4662 ;
  assign y5333 = n7186 ;
  assign y5334 = n4254 ;
  assign y5335 = ~n7191 ;
  assign y5336 = ~n3980 ;
  assign y5337 = ~1'b0 ;
  assign y5338 = ~1'b0 ;
  assign y5339 = ~n7197 ;
  assign y5340 = ~1'b0 ;
  assign y5341 = n7203 ;
  assign y5342 = ~n7214 ;
  assign y5343 = n7222 ;
  assign y5344 = ~n4037 ;
  assign y5345 = ~n7229 ;
  assign y5346 = n6291 ;
  assign y5347 = ~n7233 ;
  assign y5348 = ~1'b0 ;
  assign y5349 = ~n3015 ;
  assign y5350 = n7234 ;
  assign y5351 = ~n7236 ;
  assign y5352 = n7239 ;
  assign y5353 = ~n7240 ;
  assign y5354 = n7247 ;
  assign y5355 = ~1'b0 ;
  assign y5356 = ~n7250 ;
  assign y5357 = ~1'b0 ;
  assign y5358 = ~n7259 ;
  assign y5359 = n419 ;
  assign y5360 = ~1'b0 ;
  assign y5361 = n4763 ;
  assign y5362 = ~1'b0 ;
  assign y5363 = ~1'b0 ;
  assign y5364 = n7260 ;
  assign y5365 = ~1'b0 ;
  assign y5366 = ~n7261 ;
  assign y5367 = ~n7264 ;
  assign y5368 = 1'b0 ;
  assign y5369 = 1'b0 ;
  assign y5370 = ~n7267 ;
  assign y5371 = n7272 ;
  assign y5372 = n7275 ;
  assign y5373 = ~1'b0 ;
  assign y5374 = ~n7278 ;
  assign y5375 = ~1'b0 ;
  assign y5376 = n7279 ;
  assign y5377 = ~1'b0 ;
  assign y5378 = n7281 ;
  assign y5379 = ~1'b0 ;
  assign y5380 = ~1'b0 ;
  assign y5381 = ~1'b0 ;
  assign y5382 = ~1'b0 ;
  assign y5383 = ~1'b0 ;
  assign y5384 = n7282 ;
  assign y5385 = ~n7283 ;
  assign y5386 = ~1'b0 ;
  assign y5387 = ~1'b0 ;
  assign y5388 = ~n764 ;
  assign y5389 = ~1'b0 ;
  assign y5390 = ~n7284 ;
  assign y5391 = ~n7288 ;
  assign y5392 = ~n3539 ;
  assign y5393 = ~1'b0 ;
  assign y5394 = n7296 ;
  assign y5395 = ~n7300 ;
  assign y5396 = ~1'b0 ;
  assign y5397 = n7301 ;
  assign y5398 = ~n7303 ;
  assign y5399 = n7304 ;
  assign y5400 = ~n7305 ;
  assign y5401 = ~1'b0 ;
  assign y5402 = ~1'b0 ;
  assign y5403 = ~n7307 ;
  assign y5404 = n7311 ;
  assign y5405 = ~1'b0 ;
  assign y5406 = ~1'b0 ;
  assign y5407 = ~1'b0 ;
  assign y5408 = ~1'b0 ;
  assign y5409 = ~1'b0 ;
  assign y5410 = ~1'b0 ;
  assign y5411 = n7313 ;
  assign y5412 = ~n7316 ;
  assign y5413 = ~n7322 ;
  assign y5414 = ~n7323 ;
  assign y5415 = ~n7327 ;
  assign y5416 = ~1'b0 ;
  assign y5417 = n7328 ;
  assign y5418 = ~1'b0 ;
  assign y5419 = n7331 ;
  assign y5420 = n7333 ;
  assign y5421 = ~1'b0 ;
  assign y5422 = n5041 ;
  assign y5423 = ~n7336 ;
  assign y5424 = ~1'b0 ;
  assign y5425 = n7341 ;
  assign y5426 = ~1'b0 ;
  assign y5427 = ~n7343 ;
  assign y5428 = ~1'b0 ;
  assign y5429 = n7345 ;
  assign y5430 = ~1'b0 ;
  assign y5431 = n7348 ;
  assign y5432 = 1'b0 ;
  assign y5433 = ~n7353 ;
  assign y5434 = n7355 ;
  assign y5435 = ~1'b0 ;
  assign y5436 = ~n6553 ;
  assign y5437 = ~n7358 ;
  assign y5438 = 1'b0 ;
  assign y5439 = ~1'b0 ;
  assign y5440 = ~n7360 ;
  assign y5441 = ~1'b0 ;
  assign y5442 = ~1'b0 ;
  assign y5443 = 1'b0 ;
  assign y5444 = ~1'b0 ;
  assign y5445 = ~n7363 ;
  assign y5446 = n7364 ;
  assign y5447 = ~1'b0 ;
  assign y5448 = n7368 ;
  assign y5449 = ~1'b0 ;
  assign y5450 = ~1'b0 ;
  assign y5451 = ~n7369 ;
  assign y5452 = ~1'b0 ;
  assign y5453 = ~n7371 ;
  assign y5454 = ~n7374 ;
  assign y5455 = n7375 ;
  assign y5456 = n7376 ;
  assign y5457 = ~1'b0 ;
  assign y5458 = n7377 ;
  assign y5459 = ~1'b0 ;
  assign y5460 = ~1'b0 ;
  assign y5461 = ~n7381 ;
  assign y5462 = ~n7383 ;
  assign y5463 = n7390 ;
  assign y5464 = n7392 ;
  assign y5465 = n7394 ;
  assign y5466 = ~1'b0 ;
  assign y5467 = n7395 ;
  assign y5468 = n7397 ;
  assign y5469 = ~n7400 ;
  assign y5470 = ~1'b0 ;
  assign y5471 = ~n7407 ;
  assign y5472 = ~n7408 ;
  assign y5473 = ~1'b0 ;
  assign y5474 = ~1'b0 ;
  assign y5475 = ~n7410 ;
  assign y5476 = ~n7411 ;
  assign y5477 = ~n7413 ;
  assign y5478 = ~1'b0 ;
  assign y5479 = n7415 ;
  assign y5480 = ~1'b0 ;
  assign y5481 = ~1'b0 ;
  assign y5482 = n7417 ;
  assign y5483 = ~1'b0 ;
  assign y5484 = ~1'b0 ;
  assign y5485 = n2233 ;
  assign y5486 = ~1'b0 ;
  assign y5487 = n7418 ;
  assign y5488 = ~n7427 ;
  assign y5489 = ~n7429 ;
  assign y5490 = ~n7430 ;
  assign y5491 = ~n7431 ;
  assign y5492 = ~n7432 ;
  assign y5493 = ~1'b0 ;
  assign y5494 = ~n7438 ;
  assign y5495 = ~1'b0 ;
  assign y5496 = ~n7439 ;
  assign y5497 = n1118 ;
  assign y5498 = ~n7440 ;
  assign y5499 = ~n7442 ;
  assign y5500 = n7443 ;
  assign y5501 = ~1'b0 ;
  assign y5502 = ~n374 ;
  assign y5503 = ~1'b0 ;
  assign y5504 = ~n7448 ;
  assign y5505 = ~1'b0 ;
  assign y5506 = n7452 ;
  assign y5507 = ~1'b0 ;
  assign y5508 = ~n7454 ;
  assign y5509 = n1186 ;
  assign y5510 = n7456 ;
  assign y5511 = ~1'b0 ;
  assign y5512 = ~1'b0 ;
  assign y5513 = n7459 ;
  assign y5514 = 1'b0 ;
  assign y5515 = n7461 ;
  assign y5516 = ~n7462 ;
  assign y5517 = ~1'b0 ;
  assign y5518 = ~1'b0 ;
  assign y5519 = n7464 ;
  assign y5520 = 1'b0 ;
  assign y5521 = ~n7465 ;
  assign y5522 = ~n7471 ;
  assign y5523 = n7472 ;
  assign y5524 = 1'b0 ;
  assign y5525 = n3767 ;
  assign y5526 = ~n7477 ;
  assign y5527 = ~n7479 ;
  assign y5528 = ~n7483 ;
  assign y5529 = ~n7486 ;
  assign y5530 = ~n1331 ;
  assign y5531 = n2573 ;
  assign y5532 = ~1'b0 ;
  assign y5533 = ~1'b0 ;
  assign y5534 = ~1'b0 ;
  assign y5535 = ~1'b0 ;
  assign y5536 = ~n7487 ;
  assign y5537 = ~n7488 ;
  assign y5538 = n278 ;
  assign y5539 = ~1'b0 ;
  assign y5540 = n7489 ;
  assign y5541 = ~1'b0 ;
  assign y5542 = n6955 ;
  assign y5543 = ~n7491 ;
  assign y5544 = ~1'b0 ;
  assign y5545 = ~1'b0 ;
  assign y5546 = ~1'b0 ;
  assign y5547 = ~n7497 ;
  assign y5548 = n5152 ;
  assign y5549 = ~n7500 ;
  assign y5550 = ~n7501 ;
  assign y5551 = 1'b0 ;
  assign y5552 = ~1'b0 ;
  assign y5553 = ~1'b0 ;
  assign y5554 = ~1'b0 ;
  assign y5555 = ~n2883 ;
  assign y5556 = ~n7502 ;
  assign y5557 = ~1'b0 ;
  assign y5558 = ~1'b0 ;
  assign y5559 = ~1'b0 ;
  assign y5560 = ~n2303 ;
  assign y5561 = ~n68 ;
  assign y5562 = ~1'b0 ;
  assign y5563 = ~1'b0 ;
  assign y5564 = ~n7514 ;
  assign y5565 = 1'b0 ;
  assign y5566 = 1'b0 ;
  assign y5567 = ~1'b0 ;
  assign y5568 = ~n7520 ;
  assign y5569 = n7531 ;
  assign y5570 = ~n7532 ;
  assign y5571 = 1'b0 ;
  assign y5572 = ~n7535 ;
  assign y5573 = ~1'b0 ;
  assign y5574 = 1'b0 ;
  assign y5575 = ~n7542 ;
  assign y5576 = ~1'b0 ;
  assign y5577 = ~n7543 ;
  assign y5578 = ~1'b0 ;
  assign y5579 = n5884 ;
  assign y5580 = 1'b0 ;
  assign y5581 = ~n1917 ;
  assign y5582 = 1'b0 ;
  assign y5583 = n7545 ;
  assign y5584 = ~1'b0 ;
  assign y5585 = ~1'b0 ;
  assign y5586 = ~1'b0 ;
  assign y5587 = ~1'b0 ;
  assign y5588 = n7546 ;
  assign y5589 = ~n7550 ;
  assign y5590 = ~1'b0 ;
  assign y5591 = ~1'b0 ;
  assign y5592 = 1'b0 ;
  assign y5593 = n7552 ;
  assign y5594 = ~n7555 ;
  assign y5595 = ~n1158 ;
  assign y5596 = n7562 ;
  assign y5597 = n7563 ;
  assign y5598 = ~n7564 ;
  assign y5599 = ~1'b0 ;
  assign y5600 = n7566 ;
  assign y5601 = 1'b0 ;
  assign y5602 = n2238 ;
  assign y5603 = ~n7568 ;
  assign y5604 = ~n7570 ;
  assign y5605 = ~1'b0 ;
  assign y5606 = ~1'b0 ;
  assign y5607 = n7576 ;
  assign y5608 = n7578 ;
  assign y5609 = n7579 ;
  assign y5610 = ~1'b0 ;
  assign y5611 = n7580 ;
  assign y5612 = ~n7582 ;
  assign y5613 = ~1'b0 ;
  assign y5614 = ~1'b0 ;
  assign y5615 = ~1'b0 ;
  assign y5616 = ~n7584 ;
  assign y5617 = n7586 ;
  assign y5618 = ~n7588 ;
  assign y5619 = ~n7589 ;
  assign y5620 = ~1'b0 ;
  assign y5621 = ~1'b0 ;
  assign y5622 = ~1'b0 ;
  assign y5623 = ~n3112 ;
  assign y5624 = n7593 ;
  assign y5625 = ~1'b0 ;
  assign y5626 = ~1'b0 ;
  assign y5627 = ~1'b0 ;
  assign y5628 = ~1'b0 ;
  assign y5629 = ~1'b0 ;
  assign y5630 = n7594 ;
  assign y5631 = ~n7601 ;
  assign y5632 = ~n7603 ;
  assign y5633 = n7604 ;
  assign y5634 = ~1'b0 ;
  assign y5635 = ~n7605 ;
  assign y5636 = n7606 ;
  assign y5637 = ~n7607 ;
  assign y5638 = n7609 ;
  assign y5639 = n1856 ;
  assign y5640 = ~n7614 ;
  assign y5641 = ~1'b0 ;
  assign y5642 = n7616 ;
  assign y5643 = n7617 ;
  assign y5644 = n7619 ;
  assign y5645 = ~n7621 ;
  assign y5646 = ~n7622 ;
  assign y5647 = ~n7623 ;
  assign y5648 = ~n7625 ;
  assign y5649 = n7627 ;
  assign y5650 = n7628 ;
  assign y5651 = ~1'b0 ;
  assign y5652 = ~1'b0 ;
  assign y5653 = ~n7630 ;
  assign y5654 = ~n5551 ;
  assign y5655 = ~n7632 ;
  assign y5656 = ~n5252 ;
  assign y5657 = ~n7636 ;
  assign y5658 = ~1'b0 ;
  assign y5659 = ~1'b0 ;
  assign y5660 = ~n7637 ;
  assign y5661 = ~n7639 ;
  assign y5662 = n7641 ;
  assign y5663 = ~n7646 ;
  assign y5664 = ~n7648 ;
  assign y5665 = ~1'b0 ;
  assign y5666 = ~n308 ;
  assign y5667 = ~1'b0 ;
  assign y5668 = ~n7650 ;
  assign y5669 = ~1'b0 ;
  assign y5670 = n3338 ;
  assign y5671 = n7655 ;
  assign y5672 = ~n7657 ;
  assign y5673 = ~1'b0 ;
  assign y5674 = ~1'b0 ;
  assign y5675 = ~1'b0 ;
  assign y5676 = n7658 ;
  assign y5677 = ~n7666 ;
  assign y5678 = ~1'b0 ;
  assign y5679 = ~n7667 ;
  assign y5680 = ~n7668 ;
  assign y5681 = n2261 ;
  assign y5682 = ~1'b0 ;
  assign y5683 = 1'b0 ;
  assign y5684 = ~n5032 ;
  assign y5685 = ~n785 ;
  assign y5686 = ~n339 ;
  assign y5687 = n3533 ;
  assign y5688 = n7669 ;
  assign y5689 = ~n7670 ;
  assign y5690 = ~1'b0 ;
  assign y5691 = ~n7673 ;
  assign y5692 = ~1'b0 ;
  assign y5693 = ~n7674 ;
  assign y5694 = ~n7679 ;
  assign y5695 = ~1'b0 ;
  assign y5696 = n6462 ;
  assign y5697 = ~1'b0 ;
  assign y5698 = n7684 ;
  assign y5699 = ~n7686 ;
  assign y5700 = ~1'b0 ;
  assign y5701 = ~n7688 ;
  assign y5702 = n7689 ;
  assign y5703 = n7691 ;
  assign y5704 = n1704 ;
  assign y5705 = ~n7694 ;
  assign y5706 = n7697 ;
  assign y5707 = ~n7698 ;
  assign y5708 = ~n4923 ;
  assign y5709 = ~n1022 ;
  assign y5710 = ~1'b0 ;
  assign y5711 = n7699 ;
  assign y5712 = n7700 ;
  assign y5713 = ~1'b0 ;
  assign y5714 = ~1'b0 ;
  assign y5715 = ~1'b0 ;
  assign y5716 = 1'b0 ;
  assign y5717 = n7701 ;
  assign y5718 = ~1'b0 ;
  assign y5719 = 1'b0 ;
  assign y5720 = 1'b0 ;
  assign y5721 = ~1'b0 ;
  assign y5722 = n7261 ;
  assign y5723 = n7702 ;
  assign y5724 = ~1'b0 ;
  assign y5725 = 1'b0 ;
  assign y5726 = ~n7707 ;
  assign y5727 = ~1'b0 ;
  assign y5728 = ~n7709 ;
  assign y5729 = n7714 ;
  assign y5730 = 1'b0 ;
  assign y5731 = ~n4559 ;
  assign y5732 = n7715 ;
  assign y5733 = ~n7718 ;
  assign y5734 = n3369 ;
  assign y5735 = ~1'b0 ;
  assign y5736 = ~1'b0 ;
  assign y5737 = ~1'b0 ;
  assign y5738 = ~n7720 ;
  assign y5739 = ~n7722 ;
  assign y5740 = n7724 ;
  assign y5741 = ~n7728 ;
  assign y5742 = n1178 ;
  assign y5743 = n7730 ;
  assign y5744 = ~n7740 ;
  assign y5745 = ~1'b0 ;
  assign y5746 = ~n7744 ;
  assign y5747 = 1'b0 ;
  assign y5748 = ~n7745 ;
  assign y5749 = ~n7764 ;
  assign y5750 = ~1'b0 ;
  assign y5751 = ~n4927 ;
  assign y5752 = ~n7766 ;
  assign y5753 = ~1'b0 ;
  assign y5754 = ~n3938 ;
  assign y5755 = ~1'b0 ;
  assign y5756 = n7769 ;
  assign y5757 = ~1'b0 ;
  assign y5758 = ~1'b0 ;
  assign y5759 = ~n7770 ;
  assign y5760 = ~n7773 ;
  assign y5761 = n7777 ;
  assign y5762 = n7779 ;
  assign y5763 = n7783 ;
  assign y5764 = ~1'b0 ;
  assign y5765 = n7784 ;
  assign y5766 = n7795 ;
  assign y5767 = ~1'b0 ;
  assign y5768 = ~1'b0 ;
  assign y5769 = ~n7798 ;
  assign y5770 = 1'b0 ;
  assign y5771 = n7799 ;
  assign y5772 = n7800 ;
  assign y5773 = ~1'b0 ;
  assign y5774 = ~1'b0 ;
  assign y5775 = n7802 ;
  assign y5776 = ~n7805 ;
  assign y5777 = n7806 ;
  assign y5778 = n7807 ;
  assign y5779 = ~1'b0 ;
  assign y5780 = n7808 ;
  assign y5781 = ~n7810 ;
  assign y5782 = ~n7812 ;
  assign y5783 = ~n7815 ;
  assign y5784 = ~1'b0 ;
  assign y5785 = ~n7819 ;
  assign y5786 = ~n7824 ;
  assign y5787 = ~n7827 ;
  assign y5788 = n7843 ;
  assign y5789 = n7844 ;
  assign y5790 = n7851 ;
  assign y5791 = ~1'b0 ;
  assign y5792 = ~n7855 ;
  assign y5793 = ~n7856 ;
  assign y5794 = ~1'b0 ;
  assign y5795 = n7857 ;
  assign y5796 = ~n7862 ;
  assign y5797 = ~1'b0 ;
  assign y5798 = n7863 ;
  assign y5799 = n4068 ;
  assign y5800 = ~n4085 ;
  assign y5801 = n6944 ;
  assign y5802 = ~1'b0 ;
  assign y5803 = ~1'b0 ;
  assign y5804 = ~1'b0 ;
  assign y5805 = n7864 ;
  assign y5806 = ~1'b0 ;
  assign y5807 = 1'b0 ;
  assign y5808 = 1'b0 ;
  assign y5809 = ~n7867 ;
  assign y5810 = 1'b0 ;
  assign y5811 = n1254 ;
  assign y5812 = n7870 ;
  assign y5813 = n7875 ;
  assign y5814 = ~n7878 ;
  assign y5815 = ~n7880 ;
  assign y5816 = n2732 ;
  assign y5817 = ~n7884 ;
  assign y5818 = n7887 ;
  assign y5819 = ~n7890 ;
  assign y5820 = 1'b0 ;
  assign y5821 = ~1'b0 ;
  assign y5822 = ~n7904 ;
  assign y5823 = n7353 ;
  assign y5824 = n7907 ;
  assign y5825 = ~n7909 ;
  assign y5826 = ~1'b0 ;
  assign y5827 = ~n7910 ;
  assign y5828 = ~1'b0 ;
  assign y5829 = n7914 ;
  assign y5830 = ~1'b0 ;
  assign y5831 = n7915 ;
  assign y5832 = ~1'b0 ;
  assign y5833 = n7918 ;
  assign y5834 = ~1'b0 ;
  assign y5835 = 1'b0 ;
  assign y5836 = n814 ;
  assign y5837 = n7920 ;
  assign y5838 = ~n7921 ;
  assign y5839 = ~n7922 ;
  assign y5840 = n7924 ;
  assign y5841 = n814 ;
  assign y5842 = n942 ;
  assign y5843 = ~1'b0 ;
  assign y5844 = ~1'b0 ;
  assign y5845 = ~1'b0 ;
  assign y5846 = 1'b0 ;
  assign y5847 = ~n7926 ;
  assign y5848 = ~n7928 ;
  assign y5849 = ~n7934 ;
  assign y5850 = ~n7935 ;
  assign y5851 = ~1'b0 ;
  assign y5852 = ~n7940 ;
  assign y5853 = 1'b0 ;
  assign y5854 = ~n7943 ;
  assign y5855 = ~n7947 ;
  assign y5856 = ~1'b0 ;
  assign y5857 = ~1'b0 ;
  assign y5858 = ~1'b0 ;
  assign y5859 = n7948 ;
  assign y5860 = ~1'b0 ;
  assign y5861 = ~n7951 ;
  assign y5862 = n4650 ;
  assign y5863 = 1'b0 ;
  assign y5864 = ~n7952 ;
  assign y5865 = ~1'b0 ;
  assign y5866 = n7954 ;
  assign y5867 = n7958 ;
  assign y5868 = ~1'b0 ;
  assign y5869 = n7959 ;
  assign y5870 = ~1'b0 ;
  assign y5871 = 1'b0 ;
  assign y5872 = ~n7965 ;
  assign y5873 = n7967 ;
  assign y5874 = ~1'b0 ;
  assign y5875 = ~1'b0 ;
  assign y5876 = n7968 ;
  assign y5877 = ~1'b0 ;
  assign y5878 = n7969 ;
  assign y5879 = ~1'b0 ;
  assign y5880 = ~n6571 ;
  assign y5881 = ~1'b0 ;
  assign y5882 = n7970 ;
  assign y5883 = n7973 ;
  assign y5884 = n7975 ;
  assign y5885 = n7978 ;
  assign y5886 = ~1'b0 ;
  assign y5887 = n7980 ;
  assign y5888 = 1'b0 ;
  assign y5889 = ~1'b0 ;
  assign y5890 = n7981 ;
  assign y5891 = n7983 ;
  assign y5892 = ~n7984 ;
  assign y5893 = n7986 ;
  assign y5894 = n6653 ;
  assign y5895 = n7987 ;
  assign y5896 = ~1'b0 ;
  assign y5897 = ~1'b0 ;
  assign y5898 = n7229 ;
  assign y5899 = n2202 ;
  assign y5900 = ~1'b0 ;
  assign y5901 = ~1'b0 ;
  assign y5902 = ~1'b0 ;
  assign y5903 = ~1'b0 ;
  assign y5904 = n1663 ;
  assign y5905 = ~1'b0 ;
  assign y5906 = ~1'b0 ;
  assign y5907 = n7990 ;
  assign y5908 = 1'b0 ;
  assign y5909 = n7991 ;
  assign y5910 = n7992 ;
  assign y5911 = ~1'b0 ;
  assign y5912 = n7995 ;
  assign y5913 = ~n5396 ;
  assign y5914 = ~n7996 ;
  assign y5915 = ~1'b0 ;
  assign y5916 = n7998 ;
  assign y5917 = ~n8000 ;
  assign y5918 = ~1'b0 ;
  assign y5919 = n8001 ;
  assign y5920 = n8002 ;
  assign y5921 = ~n8004 ;
  assign y5922 = ~1'b0 ;
  assign y5923 = ~n8010 ;
  assign y5924 = ~n2027 ;
  assign y5925 = ~n8011 ;
  assign y5926 = ~n8015 ;
  assign y5927 = ~1'b0 ;
  assign y5928 = ~1'b0 ;
  assign y5929 = ~1'b0 ;
  assign y5930 = n8018 ;
  assign y5931 = ~n8019 ;
  assign y5932 = ~n8022 ;
  assign y5933 = n6534 ;
  assign y5934 = ~n1658 ;
  assign y5935 = ~1'b0 ;
  assign y5936 = n8028 ;
  assign y5937 = ~1'b0 ;
  assign y5938 = ~1'b0 ;
  assign y5939 = ~n8030 ;
  assign y5940 = ~1'b0 ;
  assign y5941 = ~n8031 ;
  assign y5942 = n8034 ;
  assign y5943 = n1002 ;
  assign y5944 = ~1'b0 ;
  assign y5945 = ~1'b0 ;
  assign y5946 = ~1'b0 ;
  assign y5947 = n8036 ;
  assign y5948 = n8037 ;
  assign y5949 = n8039 ;
  assign y5950 = n8040 ;
  assign y5951 = ~1'b0 ;
  assign y5952 = ~1'b0 ;
  assign y5953 = ~n8044 ;
  assign y5954 = ~1'b0 ;
  assign y5955 = ~1'b0 ;
  assign y5956 = ~n8047 ;
  assign y5957 = ~1'b0 ;
  assign y5958 = ~1'b0 ;
  assign y5959 = n8050 ;
  assign y5960 = ~1'b0 ;
  assign y5961 = ~n8053 ;
  assign y5962 = n8054 ;
  assign y5963 = ~1'b0 ;
  assign y5964 = n6090 ;
  assign y5965 = ~n8057 ;
  assign y5966 = ~n8059 ;
  assign y5967 = ~1'b0 ;
  assign y5968 = ~1'b0 ;
  assign y5969 = ~1'b0 ;
  assign y5970 = ~1'b0 ;
  assign y5971 = ~n8064 ;
  assign y5972 = ~n8066 ;
  assign y5973 = ~1'b0 ;
  assign y5974 = ~n8067 ;
  assign y5975 = n8068 ;
  assign y5976 = n8069 ;
  assign y5977 = ~n8070 ;
  assign y5978 = ~n8073 ;
  assign y5979 = n8075 ;
  assign y5980 = n8077 ;
  assign y5981 = ~1'b0 ;
  assign y5982 = ~1'b0 ;
  assign y5983 = ~1'b0 ;
  assign y5984 = ~1'b0 ;
  assign y5985 = n8081 ;
  assign y5986 = n8082 ;
  assign y5987 = n8084 ;
  assign y5988 = ~n8086 ;
  assign y5989 = ~1'b0 ;
  assign y5990 = ~1'b0 ;
  assign y5991 = ~n8090 ;
  assign y5992 = n8091 ;
  assign y5993 = n8092 ;
  assign y5994 = ~1'b0 ;
  assign y5995 = ~n6367 ;
  assign y5996 = ~1'b0 ;
  assign y5997 = ~n7221 ;
  assign y5998 = ~n8095 ;
  assign y5999 = ~1'b0 ;
  assign y6000 = ~1'b0 ;
  assign y6001 = ~1'b0 ;
  assign y6002 = n8099 ;
  assign y6003 = ~1'b0 ;
  assign y6004 = ~1'b0 ;
  assign y6005 = ~1'b0 ;
  assign y6006 = ~1'b0 ;
  assign y6007 = n8101 ;
  assign y6008 = ~1'b0 ;
  assign y6009 = n2627 ;
  assign y6010 = 1'b0 ;
  assign y6011 = n8104 ;
  assign y6012 = ~1'b0 ;
  assign y6013 = ~n8105 ;
  assign y6014 = ~n8106 ;
  assign y6015 = ~1'b0 ;
  assign y6016 = ~1'b0 ;
  assign y6017 = ~1'b0 ;
  assign y6018 = ~1'b0 ;
  assign y6019 = ~1'b0 ;
  assign y6020 = n8107 ;
  assign y6021 = ~n8108 ;
  assign y6022 = n8109 ;
  assign y6023 = ~1'b0 ;
  assign y6024 = n8110 ;
  assign y6025 = ~1'b0 ;
  assign y6026 = ~n8114 ;
  assign y6027 = n8115 ;
  assign y6028 = n8116 ;
  assign y6029 = n8117 ;
  assign y6030 = n8119 ;
  assign y6031 = ~n8122 ;
  assign y6032 = n8127 ;
  assign y6033 = ~n84 ;
  assign y6034 = ~1'b0 ;
  assign y6035 = ~n1349 ;
  assign y6036 = ~n8128 ;
  assign y6037 = n8129 ;
  assign y6038 = ~n4320 ;
  assign y6039 = ~1'b0 ;
  assign y6040 = ~1'b0 ;
  assign y6041 = n8134 ;
  assign y6042 = ~n8135 ;
  assign y6043 = ~1'b0 ;
  assign y6044 = ~n8137 ;
  assign y6045 = ~1'b0 ;
  assign y6046 = ~1'b0 ;
  assign y6047 = n8138 ;
  assign y6048 = ~1'b0 ;
  assign y6049 = ~n8140 ;
  assign y6050 = ~1'b0 ;
  assign y6051 = n8143 ;
  assign y6052 = ~1'b0 ;
  assign y6053 = 1'b0 ;
  assign y6054 = ~1'b0 ;
  assign y6055 = ~1'b0 ;
  assign y6056 = ~1'b0 ;
  assign y6057 = ~n8144 ;
  assign y6058 = n8148 ;
  assign y6059 = ~n8151 ;
  assign y6060 = n8155 ;
  assign y6061 = n8156 ;
  assign y6062 = ~1'b0 ;
  assign y6063 = 1'b0 ;
  assign y6064 = n8158 ;
  assign y6065 = n8160 ;
  assign y6066 = ~n8162 ;
  assign y6067 = n8163 ;
  assign y6068 = n8166 ;
  assign y6069 = ~n8169 ;
  assign y6070 = n8171 ;
  assign y6071 = ~1'b0 ;
  assign y6072 = ~1'b0 ;
  assign y6073 = ~n8172 ;
  assign y6074 = ~n8179 ;
  assign y6075 = ~n8184 ;
  assign y6076 = ~n8185 ;
  assign y6077 = ~n8186 ;
  assign y6078 = ~1'b0 ;
  assign y6079 = ~1'b0 ;
  assign y6080 = ~1'b0 ;
  assign y6081 = n8191 ;
  assign y6082 = ~1'b0 ;
  assign y6083 = ~n8192 ;
  assign y6084 = n8195 ;
  assign y6085 = ~1'b0 ;
  assign y6086 = ~n8198 ;
  assign y6087 = ~1'b0 ;
  assign y6088 = n8117 ;
  assign y6089 = n8199 ;
  assign y6090 = ~1'b0 ;
  assign y6091 = n8202 ;
  assign y6092 = ~n8205 ;
  assign y6093 = 1'b0 ;
  assign y6094 = ~1'b0 ;
  assign y6095 = ~n8206 ;
  assign y6096 = n8207 ;
  assign y6097 = n8212 ;
  assign y6098 = ~1'b0 ;
  assign y6099 = 1'b0 ;
  assign y6100 = n8214 ;
  assign y6101 = n8216 ;
  assign y6102 = ~n8217 ;
  assign y6103 = ~1'b0 ;
  assign y6104 = ~n4070 ;
  assign y6105 = 1'b0 ;
  assign y6106 = ~n8218 ;
  assign y6107 = ~1'b0 ;
  assign y6108 = n8219 ;
  assign y6109 = ~n8220 ;
  assign y6110 = ~1'b0 ;
  assign y6111 = n8223 ;
  assign y6112 = n7383 ;
  assign y6113 = n8224 ;
  assign y6114 = ~1'b0 ;
  assign y6115 = ~1'b0 ;
  assign y6116 = n8225 ;
  assign y6117 = n8227 ;
  assign y6118 = ~n8229 ;
  assign y6119 = n2752 ;
  assign y6120 = ~1'b0 ;
  assign y6121 = ~1'b0 ;
  assign y6122 = n3539 ;
  assign y6123 = ~1'b0 ;
  assign y6124 = n8230 ;
  assign y6125 = n8231 ;
  assign y6126 = 1'b0 ;
  assign y6127 = ~1'b0 ;
  assign y6128 = ~1'b0 ;
  assign y6129 = ~1'b0 ;
  assign y6130 = ~n8232 ;
  assign y6131 = ~1'b0 ;
  assign y6132 = ~n8239 ;
  assign y6133 = n8242 ;
  assign y6134 = ~1'b0 ;
  assign y6135 = ~n8244 ;
  assign y6136 = ~n8247 ;
  assign y6137 = ~n8248 ;
  assign y6138 = ~n8249 ;
  assign y6139 = ~1'b0 ;
  assign y6140 = n8253 ;
  assign y6141 = n8256 ;
  assign y6142 = ~n8261 ;
  assign y6143 = n8262 ;
  assign y6144 = ~1'b0 ;
  assign y6145 = n8264 ;
  assign y6146 = ~1'b0 ;
  assign y6147 = ~1'b0 ;
  assign y6148 = ~1'b0 ;
  assign y6149 = n8266 ;
  assign y6150 = n8274 ;
  assign y6151 = n8275 ;
  assign y6152 = ~n8278 ;
  assign y6153 = ~n8280 ;
  assign y6154 = n8281 ;
  assign y6155 = ~1'b0 ;
  assign y6156 = ~1'b0 ;
  assign y6157 = ~1'b0 ;
  assign y6158 = ~1'b0 ;
  assign y6159 = n8282 ;
  assign y6160 = n5860 ;
  assign y6161 = n8285 ;
  assign y6162 = ~1'b0 ;
  assign y6163 = n8288 ;
  assign y6164 = ~1'b0 ;
  assign y6165 = ~n8290 ;
  assign y6166 = n8292 ;
  assign y6167 = ~1'b0 ;
  assign y6168 = ~1'b0 ;
  assign y6169 = ~1'b0 ;
  assign y6170 = ~1'b0 ;
  assign y6171 = n8294 ;
  assign y6172 = ~1'b0 ;
  assign y6173 = n8298 ;
  assign y6174 = 1'b0 ;
  assign y6175 = ~1'b0 ;
  assign y6176 = ~n5663 ;
  assign y6177 = ~1'b0 ;
  assign y6178 = 1'b0 ;
  assign y6179 = ~1'b0 ;
  assign y6180 = n8299 ;
  assign y6181 = ~n8304 ;
  assign y6182 = ~1'b0 ;
  assign y6183 = ~n8305 ;
  assign y6184 = ~n8311 ;
  assign y6185 = ~1'b0 ;
  assign y6186 = ~n7430 ;
  assign y6187 = ~n8314 ;
  assign y6188 = n8316 ;
  assign y6189 = ~n8318 ;
  assign y6190 = n8320 ;
  assign y6191 = ~n8322 ;
  assign y6192 = ~n8323 ;
  assign y6193 = ~1'b0 ;
  assign y6194 = n8324 ;
  assign y6195 = ~n8327 ;
  assign y6196 = ~1'b0 ;
  assign y6197 = ~1'b0 ;
  assign y6198 = n8330 ;
  assign y6199 = n8333 ;
  assign y6200 = ~n8346 ;
  assign y6201 = ~1'b0 ;
  assign y6202 = n2842 ;
  assign y6203 = ~n8347 ;
  assign y6204 = n8350 ;
  assign y6205 = ~n8351 ;
  assign y6206 = ~1'b0 ;
  assign y6207 = n8355 ;
  assign y6208 = ~n8358 ;
  assign y6209 = n8362 ;
  assign y6210 = ~1'b0 ;
  assign y6211 = ~1'b0 ;
  assign y6212 = ~n8368 ;
  assign y6213 = n8370 ;
  assign y6214 = ~x8 ;
  assign y6215 = ~n8372 ;
  assign y6216 = n8373 ;
  assign y6217 = ~1'b0 ;
  assign y6218 = n8377 ;
  assign y6219 = n4778 ;
  assign y6220 = n8381 ;
  assign y6221 = ~1'b0 ;
  assign y6222 = ~1'b0 ;
  assign y6223 = 1'b0 ;
  assign y6224 = n2797 ;
  assign y6225 = ~1'b0 ;
  assign y6226 = ~1'b0 ;
  assign y6227 = ~n8384 ;
  assign y6228 = n1226 ;
  assign y6229 = n8387 ;
  assign y6230 = n8388 ;
  assign y6231 = ~1'b0 ;
  assign y6232 = ~1'b0 ;
  assign y6233 = ~n8391 ;
  assign y6234 = ~n8395 ;
  assign y6235 = ~1'b0 ;
  assign y6236 = n8396 ;
  assign y6237 = ~n8397 ;
  assign y6238 = ~1'b0 ;
  assign y6239 = ~1'b0 ;
  assign y6240 = n8399 ;
  assign y6241 = ~n8402 ;
  assign y6242 = ~n3566 ;
  assign y6243 = ~1'b0 ;
  assign y6244 = ~1'b0 ;
  assign y6245 = ~n1974 ;
  assign y6246 = n8403 ;
  assign y6247 = ~n8406 ;
  assign y6248 = ~n8407 ;
  assign y6249 = n8410 ;
  assign y6250 = ~1'b0 ;
  assign y6251 = ~1'b0 ;
  assign y6252 = 1'b0 ;
  assign y6253 = ~1'b0 ;
  assign y6254 = ~1'b0 ;
  assign y6255 = 1'b0 ;
  assign y6256 = n8414 ;
  assign y6257 = ~1'b0 ;
  assign y6258 = ~1'b0 ;
  assign y6259 = 1'b0 ;
  assign y6260 = n8415 ;
  assign y6261 = ~1'b0 ;
  assign y6262 = n8416 ;
  assign y6263 = ~1'b0 ;
  assign y6264 = ~n8419 ;
  assign y6265 = ~1'b0 ;
  assign y6266 = ~1'b0 ;
  assign y6267 = ~n1117 ;
  assign y6268 = n8421 ;
  assign y6269 = n8422 ;
  assign y6270 = ~n8424 ;
  assign y6271 = n3369 ;
  assign y6272 = ~1'b0 ;
  assign y6273 = ~n8426 ;
  assign y6274 = n8429 ;
  assign y6275 = n8430 ;
  assign y6276 = 1'b0 ;
  assign y6277 = ~1'b0 ;
  assign y6278 = ~1'b0 ;
  assign y6279 = ~n8432 ;
  assign y6280 = ~1'b0 ;
  assign y6281 = ~1'b0 ;
  assign y6282 = 1'b0 ;
  assign y6283 = ~1'b0 ;
  assign y6284 = ~n8437 ;
  assign y6285 = ~1'b0 ;
  assign y6286 = ~1'b0 ;
  assign y6287 = ~n8441 ;
  assign y6288 = n8444 ;
  assign y6289 = ~1'b0 ;
  assign y6290 = ~1'b0 ;
  assign y6291 = ~n8445 ;
  assign y6292 = n4748 ;
  assign y6293 = ~1'b0 ;
  assign y6294 = ~n8448 ;
  assign y6295 = ~1'b0 ;
  assign y6296 = n8451 ;
  assign y6297 = ~1'b0 ;
  assign y6298 = n8452 ;
  assign y6299 = ~1'b0 ;
  assign y6300 = n5046 ;
  assign y6301 = n8457 ;
  assign y6302 = ~1'b0 ;
  assign y6303 = 1'b0 ;
  assign y6304 = n8458 ;
  assign y6305 = n8459 ;
  assign y6306 = ~1'b0 ;
  assign y6307 = ~1'b0 ;
  assign y6308 = ~n4332 ;
  assign y6309 = n8461 ;
  assign y6310 = n5393 ;
  assign y6311 = ~1'b0 ;
  assign y6312 = ~1'b0 ;
  assign y6313 = ~1'b0 ;
  assign y6314 = ~1'b0 ;
  assign y6315 = n8463 ;
  assign y6316 = n8464 ;
  assign y6317 = n8467 ;
  assign y6318 = n8469 ;
  assign y6319 = ~n8470 ;
  assign y6320 = n8472 ;
  assign y6321 = ~1'b0 ;
  assign y6322 = ~1'b0 ;
  assign y6323 = ~1'b0 ;
  assign y6324 = ~1'b0 ;
  assign y6325 = ~1'b0 ;
  assign y6326 = ~1'b0 ;
  assign y6327 = ~n4365 ;
  assign y6328 = ~1'b0 ;
  assign y6329 = n4895 ;
  assign y6330 = ~n8475 ;
  assign y6331 = ~n8477 ;
  assign y6332 = ~n8479 ;
  assign y6333 = 1'b0 ;
  assign y6334 = ~1'b0 ;
  assign y6335 = n8480 ;
  assign y6336 = n2757 ;
  assign y6337 = ~n8482 ;
  assign y6338 = ~n8487 ;
  assign y6339 = ~n8489 ;
  assign y6340 = ~n8490 ;
  assign y6341 = ~1'b0 ;
  assign y6342 = ~1'b0 ;
  assign y6343 = ~1'b0 ;
  assign y6344 = n8491 ;
  assign y6345 = ~n8493 ;
  assign y6346 = ~1'b0 ;
  assign y6347 = n962 ;
  assign y6348 = ~n8494 ;
  assign y6349 = ~n8499 ;
  assign y6350 = ~1'b0 ;
  assign y6351 = ~n8503 ;
  assign y6352 = ~n8510 ;
  assign y6353 = ~1'b0 ;
  assign y6354 = ~n8512 ;
  assign y6355 = n934 ;
  assign y6356 = n7497 ;
  assign y6357 = ~1'b0 ;
  assign y6358 = ~1'b0 ;
  assign y6359 = n8517 ;
  assign y6360 = ~1'b0 ;
  assign y6361 = ~n8521 ;
  assign y6362 = ~1'b0 ;
  assign y6363 = ~1'b0 ;
  assign y6364 = ~1'b0 ;
  assign y6365 = ~1'b0 ;
  assign y6366 = n8524 ;
  assign y6367 = ~n8525 ;
  assign y6368 = ~1'b0 ;
  assign y6369 = ~n8526 ;
  assign y6370 = n501 ;
  assign y6371 = ~1'b0 ;
  assign y6372 = n8529 ;
  assign y6373 = ~n8530 ;
  assign y6374 = ~1'b0 ;
  assign y6375 = ~n1961 ;
  assign y6376 = n8534 ;
  assign y6377 = ~1'b0 ;
  assign y6378 = ~n8540 ;
  assign y6379 = n8541 ;
  assign y6380 = ~n8543 ;
  assign y6381 = n8546 ;
  assign y6382 = ~1'b0 ;
  assign y6383 = ~n8548 ;
  assign y6384 = ~1'b0 ;
  assign y6385 = ~n8549 ;
  assign y6386 = ~1'b0 ;
  assign y6387 = n8550 ;
  assign y6388 = n8551 ;
  assign y6389 = n8553 ;
  assign y6390 = n8555 ;
  assign y6391 = ~n8557 ;
  assign y6392 = n8559 ;
  assign y6393 = ~1'b0 ;
  assign y6394 = ~n8561 ;
  assign y6395 = ~1'b0 ;
  assign y6396 = ~n8562 ;
  assign y6397 = ~1'b0 ;
  assign y6398 = ~n695 ;
  assign y6399 = n8564 ;
  assign y6400 = ~1'b0 ;
  assign y6401 = ~1'b0 ;
  assign y6402 = ~n8567 ;
  assign y6403 = n8014 ;
  assign y6404 = n8571 ;
  assign y6405 = ~1'b0 ;
  assign y6406 = ~n8573 ;
  assign y6407 = ~n8575 ;
  assign y6408 = ~1'b0 ;
  assign y6409 = 1'b0 ;
  assign y6410 = ~n8579 ;
  assign y6411 = n8582 ;
  assign y6412 = ~1'b0 ;
  assign y6413 = ~1'b0 ;
  assign y6414 = n8583 ;
  assign y6415 = n8587 ;
  assign y6416 = n8594 ;
  assign y6417 = ~1'b0 ;
  assign y6418 = n8595 ;
  assign y6419 = 1'b0 ;
  assign y6420 = ~1'b0 ;
  assign y6421 = ~n8596 ;
  assign y6422 = ~1'b0 ;
  assign y6423 = ~1'b0 ;
  assign y6424 = n8599 ;
  assign y6425 = ~n8601 ;
  assign y6426 = ~1'b0 ;
  assign y6427 = n8605 ;
  assign y6428 = ~n8608 ;
  assign y6429 = ~n8609 ;
  assign y6430 = ~n8611 ;
  assign y6431 = 1'b0 ;
  assign y6432 = n8616 ;
  assign y6433 = n8619 ;
  assign y6434 = 1'b0 ;
  assign y6435 = ~1'b0 ;
  assign y6436 = ~1'b0 ;
  assign y6437 = ~n8620 ;
  assign y6438 = n8623 ;
  assign y6439 = ~1'b0 ;
  assign y6440 = ~1'b0 ;
  assign y6441 = ~1'b0 ;
  assign y6442 = n8624 ;
  assign y6443 = ~n8625 ;
  assign y6444 = ~n8626 ;
  assign y6445 = n8627 ;
  assign y6446 = ~n8628 ;
  assign y6447 = n8629 ;
  assign y6448 = ~n8643 ;
  assign y6449 = ~n8644 ;
  assign y6450 = n4954 ;
  assign y6451 = ~1'b0 ;
  assign y6452 = n8648 ;
  assign y6453 = ~1'b0 ;
  assign y6454 = n8652 ;
  assign y6455 = ~n1172 ;
  assign y6456 = ~n8653 ;
  assign y6457 = ~1'b0 ;
  assign y6458 = n8656 ;
  assign y6459 = ~1'b0 ;
  assign y6460 = n8657 ;
  assign y6461 = ~n8659 ;
  assign y6462 = ~1'b0 ;
  assign y6463 = n8664 ;
  assign y6464 = ~n8665 ;
  assign y6465 = 1'b0 ;
  assign y6466 = ~n2321 ;
  assign y6467 = n8667 ;
  assign y6468 = ~1'b0 ;
  assign y6469 = ~n8668 ;
  assign y6470 = ~n8669 ;
  assign y6471 = n8670 ;
  assign y6472 = ~n8672 ;
  assign y6473 = ~n8151 ;
  assign y6474 = n8674 ;
  assign y6475 = ~1'b0 ;
  assign y6476 = ~1'b0 ;
  assign y6477 = n8681 ;
  assign y6478 = n8539 ;
  assign y6479 = ~n7310 ;
  assign y6480 = ~1'b0 ;
  assign y6481 = 1'b0 ;
  assign y6482 = ~n8684 ;
  assign y6483 = 1'b0 ;
  assign y6484 = 1'b0 ;
  assign y6485 = ~n8686 ;
  assign y6486 = ~1'b0 ;
  assign y6487 = ~1'b0 ;
  assign y6488 = n8687 ;
  assign y6489 = ~n8689 ;
  assign y6490 = ~1'b0 ;
  assign y6491 = ~n6249 ;
  assign y6492 = ~1'b0 ;
  assign y6493 = ~n2964 ;
  assign y6494 = ~1'b0 ;
  assign y6495 = ~n8703 ;
  assign y6496 = ~n8704 ;
  assign y6497 = n8707 ;
  assign y6498 = n8708 ;
  assign y6499 = ~n8710 ;
  assign y6500 = ~1'b0 ;
  assign y6501 = ~n8711 ;
  assign y6502 = ~1'b0 ;
  assign y6503 = n8081 ;
  assign y6504 = n8717 ;
  assign y6505 = n8718 ;
  assign y6506 = ~1'b0 ;
  assign y6507 = ~n8719 ;
  assign y6508 = ~n1041 ;
  assign y6509 = ~n8723 ;
  assign y6510 = n8726 ;
  assign y6511 = n8728 ;
  assign y6512 = n1298 ;
  assign y6513 = ~n8729 ;
  assign y6514 = ~1'b0 ;
  assign y6515 = ~n8732 ;
  assign y6516 = ~n8734 ;
  assign y6517 = ~1'b0 ;
  assign y6518 = ~n5256 ;
  assign y6519 = ~1'b0 ;
  assign y6520 = n8739 ;
  assign y6521 = ~1'b0 ;
  assign y6522 = n8745 ;
  assign y6523 = ~1'b0 ;
  assign y6524 = ~n8747 ;
  assign y6525 = ~1'b0 ;
  assign y6526 = n8751 ;
  assign y6527 = ~1'b0 ;
  assign y6528 = ~1'b0 ;
  assign y6529 = ~n3269 ;
  assign y6530 = ~n8756 ;
  assign y6531 = ~1'b0 ;
  assign y6532 = ~n8757 ;
  assign y6533 = ~1'b0 ;
  assign y6534 = ~n8760 ;
  assign y6535 = n8764 ;
  assign y6536 = ~1'b0 ;
  assign y6537 = ~1'b0 ;
  assign y6538 = ~n8765 ;
  assign y6539 = ~n8768 ;
  assign y6540 = ~1'b0 ;
  assign y6541 = ~1'b0 ;
  assign y6542 = n8773 ;
  assign y6543 = n8775 ;
  assign y6544 = n8064 ;
  assign y6545 = ~1'b0 ;
  assign y6546 = ~n4927 ;
  assign y6547 = n8779 ;
  assign y6548 = ~n8780 ;
  assign y6549 = ~n8783 ;
  assign y6550 = ~1'b0 ;
  assign y6551 = n8785 ;
  assign y6552 = ~n8792 ;
  assign y6553 = ~n8793 ;
  assign y6554 = n159 ;
  assign y6555 = ~n4748 ;
  assign y6556 = n8797 ;
  assign y6557 = n532 ;
  assign y6558 = ~n8798 ;
  assign y6559 = n8802 ;
  assign y6560 = ~n8803 ;
  assign y6561 = n8804 ;
  assign y6562 = ~1'b0 ;
  assign y6563 = n8811 ;
  assign y6564 = n8812 ;
  assign y6565 = n8813 ;
  assign y6566 = n5501 ;
  assign y6567 = ~n8814 ;
  assign y6568 = ~n6546 ;
  assign y6569 = ~n8819 ;
  assign y6570 = n2642 ;
  assign y6571 = ~n8820 ;
  assign y6572 = n8823 ;
  assign y6573 = ~1'b0 ;
  assign y6574 = n8824 ;
  assign y6575 = ~n8826 ;
  assign y6576 = n5774 ;
  assign y6577 = n8829 ;
  assign y6578 = n8832 ;
  assign y6579 = 1'b0 ;
  assign y6580 = ~n8838 ;
  assign y6581 = n8841 ;
  assign y6582 = ~1'b0 ;
  assign y6583 = n8843 ;
  assign y6584 = n8845 ;
  assign y6585 = ~n8846 ;
  assign y6586 = 1'b0 ;
  assign y6587 = ~n8847 ;
  assign y6588 = ~1'b0 ;
  assign y6589 = ~n8848 ;
  assign y6590 = ~n8851 ;
  assign y6591 = ~n8853 ;
  assign y6592 = 1'b0 ;
  assign y6593 = n8854 ;
  assign y6594 = ~1'b0 ;
  assign y6595 = ~n8855 ;
  assign y6596 = ~n8857 ;
  assign y6597 = ~1'b0 ;
  assign y6598 = ~n8858 ;
  assign y6599 = ~n8862 ;
  assign y6600 = n8863 ;
  assign y6601 = n8866 ;
  assign y6602 = ~1'b0 ;
  assign y6603 = ~1'b0 ;
  assign y6604 = ~1'b0 ;
  assign y6605 = ~n8869 ;
  assign y6606 = ~1'b0 ;
  assign y6607 = ~n8870 ;
  assign y6608 = ~n8872 ;
  assign y6609 = ~n1110 ;
  assign y6610 = n8877 ;
  assign y6611 = ~1'b0 ;
  assign y6612 = ~1'b0 ;
  assign y6613 = ~n8879 ;
  assign y6614 = ~n8883 ;
  assign y6615 = ~n8884 ;
  assign y6616 = ~1'b0 ;
  assign y6617 = ~n8885 ;
  assign y6618 = ~n8887 ;
  assign y6619 = n8889 ;
  assign y6620 = ~n8893 ;
  assign y6621 = n8896 ;
  assign y6622 = n8897 ;
  assign y6623 = ~1'b0 ;
  assign y6624 = ~n8898 ;
  assign y6625 = ~1'b0 ;
  assign y6626 = ~1'b0 ;
  assign y6627 = ~n8900 ;
  assign y6628 = ~n2414 ;
  assign y6629 = ~1'b0 ;
  assign y6630 = 1'b0 ;
  assign y6631 = n8902 ;
  assign y6632 = ~n8904 ;
  assign y6633 = n8905 ;
  assign y6634 = n8908 ;
  assign y6635 = ~n8910 ;
  assign y6636 = ~1'b0 ;
  assign y6637 = ~n8915 ;
  assign y6638 = ~1'b0 ;
  assign y6639 = n8919 ;
  assign y6640 = ~1'b0 ;
  assign y6641 = ~1'b0 ;
  assign y6642 = ~n8921 ;
  assign y6643 = ~1'b0 ;
  assign y6644 = n8923 ;
  assign y6645 = ~1'b0 ;
  assign y6646 = ~1'b0 ;
  assign y6647 = ~n8925 ;
  assign y6648 = n8928 ;
  assign y6649 = n8932 ;
  assign y6650 = ~1'b0 ;
  assign y6651 = n8933 ;
  assign y6652 = ~n8935 ;
  assign y6653 = n8941 ;
  assign y6654 = ~n8942 ;
  assign y6655 = 1'b0 ;
  assign y6656 = ~1'b0 ;
  assign y6657 = n8944 ;
  assign y6658 = ~n8945 ;
  assign y6659 = ~n3089 ;
  assign y6660 = ~1'b0 ;
  assign y6661 = ~1'b0 ;
  assign y6662 = ~1'b0 ;
  assign y6663 = ~n8946 ;
  assign y6664 = n6009 ;
  assign y6665 = ~n8947 ;
  assign y6666 = ~n8948 ;
  assign y6667 = ~1'b0 ;
  assign y6668 = ~n8951 ;
  assign y6669 = 1'b0 ;
  assign y6670 = n7350 ;
  assign y6671 = ~1'b0 ;
  assign y6672 = ~1'b0 ;
  assign y6673 = n8957 ;
  assign y6674 = ~n8959 ;
  assign y6675 = n8488 ;
  assign y6676 = 1'b0 ;
  assign y6677 = ~n8965 ;
  assign y6678 = ~1'b0 ;
  assign y6679 = ~1'b0 ;
  assign y6680 = ~1'b0 ;
  assign y6681 = ~1'b0 ;
  assign y6682 = n8966 ;
  assign y6683 = ~1'b0 ;
  assign y6684 = n8971 ;
  assign y6685 = 1'b0 ;
  assign y6686 = ~1'b0 ;
  assign y6687 = n8972 ;
  assign y6688 = ~1'b0 ;
  assign y6689 = n8973 ;
  assign y6690 = ~n8976 ;
  assign y6691 = n8977 ;
  assign y6692 = ~n8980 ;
  assign y6693 = ~n8986 ;
  assign y6694 = n8987 ;
  assign y6695 = n4934 ;
  assign y6696 = n8988 ;
  assign y6697 = ~n8989 ;
  assign y6698 = n2680 ;
  assign y6699 = n8990 ;
  assign y6700 = ~1'b0 ;
  assign y6701 = n8991 ;
  assign y6702 = ~1'b0 ;
  assign y6703 = n8992 ;
  assign y6704 = n8993 ;
  assign y6705 = ~n8995 ;
  assign y6706 = ~n8998 ;
  assign y6707 = ~n8999 ;
  assign y6708 = n9000 ;
  assign y6709 = n339 ;
  assign y6710 = ~n9008 ;
  assign y6711 = ~n9009 ;
  assign y6712 = n9010 ;
  assign y6713 = ~n9011 ;
  assign y6714 = ~n5516 ;
  assign y6715 = n9012 ;
  assign y6716 = ~n9015 ;
  assign y6717 = n9017 ;
  assign y6718 = ~n9018 ;
  assign y6719 = ~n9019 ;
  assign y6720 = ~1'b0 ;
  assign y6721 = ~1'b0 ;
  assign y6722 = ~1'b0 ;
  assign y6723 = ~1'b0 ;
  assign y6724 = n9020 ;
  assign y6725 = ~1'b0 ;
  assign y6726 = ~n7597 ;
  assign y6727 = n9024 ;
  assign y6728 = ~n9026 ;
  assign y6729 = ~n9030 ;
  assign y6730 = ~n9036 ;
  assign y6731 = ~n9038 ;
  assign y6732 = ~1'b0 ;
  assign y6733 = ~1'b0 ;
  assign y6734 = ~n9039 ;
  assign y6735 = ~n9041 ;
  assign y6736 = n9043 ;
  assign y6737 = ~n2933 ;
  assign y6738 = ~1'b0 ;
  assign y6739 = n9045 ;
  assign y6740 = n9046 ;
  assign y6741 = ~n9047 ;
  assign y6742 = ~1'b0 ;
  assign y6743 = ~1'b0 ;
  assign y6744 = ~n9048 ;
  assign y6745 = n6876 ;
  assign y6746 = ~n9051 ;
  assign y6747 = n9052 ;
  assign y6748 = n9055 ;
  assign y6749 = ~1'b0 ;
  assign y6750 = ~1'b0 ;
  assign y6751 = ~n9060 ;
  assign y6752 = ~1'b0 ;
  assign y6753 = n6536 ;
  assign y6754 = n9061 ;
  assign y6755 = ~1'b0 ;
  assign y6756 = ~1'b0 ;
  assign y6757 = ~n9062 ;
  assign y6758 = n9064 ;
  assign y6759 = n9066 ;
  assign y6760 = ~1'b0 ;
  assign y6761 = 1'b0 ;
  assign y6762 = ~1'b0 ;
  assign y6763 = ~n9067 ;
  assign y6764 = ~n9070 ;
  assign y6765 = ~1'b0 ;
  assign y6766 = ~1'b0 ;
  assign y6767 = ~n4700 ;
  assign y6768 = ~n2269 ;
  assign y6769 = n9077 ;
  assign y6770 = n9082 ;
  assign y6771 = n9083 ;
  assign y6772 = ~n2311 ;
  assign y6773 = n9084 ;
  assign y6774 = n9085 ;
  assign y6775 = n9086 ;
  assign y6776 = 1'b0 ;
  assign y6777 = ~n9092 ;
  assign y6778 = ~n9099 ;
  assign y6779 = ~1'b0 ;
  assign y6780 = ~1'b0 ;
  assign y6781 = 1'b0 ;
  assign y6782 = ~n9103 ;
  assign y6783 = ~n9104 ;
  assign y6784 = ~n159 ;
  assign y6785 = n9105 ;
  assign y6786 = ~1'b0 ;
  assign y6787 = n9107 ;
  assign y6788 = n9108 ;
  assign y6789 = ~n9109 ;
  assign y6790 = n489 ;
  assign y6791 = ~n7483 ;
  assign y6792 = n9117 ;
  assign y6793 = ~n9119 ;
  assign y6794 = ~n9121 ;
  assign y6795 = n9124 ;
  assign y6796 = ~1'b0 ;
  assign y6797 = ~1'b0 ;
  assign y6798 = n9126 ;
  assign y6799 = n9128 ;
  assign y6800 = n9130 ;
  assign y6801 = n428 ;
  assign y6802 = ~1'b0 ;
  assign y6803 = n3150 ;
  assign y6804 = ~n9132 ;
  assign y6805 = ~1'b0 ;
  assign y6806 = ~n9134 ;
  assign y6807 = n9135 ;
  assign y6808 = ~1'b0 ;
  assign y6809 = ~n9136 ;
  assign y6810 = ~1'b0 ;
  assign y6811 = n670 ;
  assign y6812 = ~1'b0 ;
  assign y6813 = n9140 ;
  assign y6814 = ~1'b0 ;
  assign y6815 = n9141 ;
  assign y6816 = ~1'b0 ;
  assign y6817 = n9149 ;
  assign y6818 = ~n9151 ;
  assign y6819 = ~1'b0 ;
  assign y6820 = ~1'b0 ;
  assign y6821 = ~n6250 ;
  assign y6822 = n9153 ;
  assign y6823 = ~n9155 ;
  assign y6824 = ~1'b0 ;
  assign y6825 = n9157 ;
  assign y6826 = ~1'b0 ;
  assign y6827 = ~1'b0 ;
  assign y6828 = ~1'b0 ;
  assign y6829 = n9159 ;
  assign y6830 = ~n9161 ;
  assign y6831 = ~1'b0 ;
  assign y6832 = ~n9164 ;
  assign y6833 = ~n9169 ;
  assign y6834 = ~1'b0 ;
  assign y6835 = 1'b0 ;
  assign y6836 = ~n9170 ;
  assign y6837 = n9171 ;
  assign y6838 = ~1'b0 ;
  assign y6839 = ~n3095 ;
  assign y6840 = ~1'b0 ;
  assign y6841 = ~n9172 ;
  assign y6842 = n9174 ;
  assign y6843 = ~n9176 ;
  assign y6844 = n6114 ;
  assign y6845 = ~1'b0 ;
  assign y6846 = n9177 ;
  assign y6847 = ~1'b0 ;
  assign y6848 = n9180 ;
  assign y6849 = ~1'b0 ;
  assign y6850 = ~1'b0 ;
  assign y6851 = ~n9182 ;
  assign y6852 = ~1'b0 ;
  assign y6853 = n9186 ;
  assign y6854 = ~1'b0 ;
  assign y6855 = n1233 ;
  assign y6856 = n9188 ;
  assign y6857 = ~1'b0 ;
  assign y6858 = n9191 ;
  assign y6859 = ~n9192 ;
  assign y6860 = ~1'b0 ;
  assign y6861 = ~1'b0 ;
  assign y6862 = 1'b0 ;
  assign y6863 = ~n9193 ;
  assign y6864 = n9194 ;
  assign y6865 = ~1'b0 ;
  assign y6866 = ~n9198 ;
  assign y6867 = ~n9199 ;
  assign y6868 = ~n9204 ;
  assign y6869 = n9208 ;
  assign y6870 = n1834 ;
  assign y6871 = ~1'b0 ;
  assign y6872 = n9210 ;
  assign y6873 = ~1'b0 ;
  assign y6874 = n9212 ;
  assign y6875 = ~n2261 ;
  assign y6876 = n9213 ;
  assign y6877 = ~1'b0 ;
  assign y6878 = n9216 ;
  assign y6879 = n3394 ;
  assign y6880 = ~1'b0 ;
  assign y6881 = ~n9217 ;
  assign y6882 = ~1'b0 ;
  assign y6883 = n9220 ;
  assign y6884 = n9222 ;
  assign y6885 = n9223 ;
  assign y6886 = ~1'b0 ;
  assign y6887 = ~n9225 ;
  assign y6888 = ~n9230 ;
  assign y6889 = ~n9233 ;
  assign y6890 = ~1'b0 ;
  assign y6891 = n9235 ;
  assign y6892 = n9236 ;
  assign y6893 = ~1'b0 ;
  assign y6894 = n9237 ;
  assign y6895 = ~n9240 ;
  assign y6896 = 1'b0 ;
  assign y6897 = n9251 ;
  assign y6898 = ~n9252 ;
  assign y6899 = n9253 ;
  assign y6900 = ~n9261 ;
  assign y6901 = ~n9263 ;
  assign y6902 = n9265 ;
  assign y6903 = ~n9268 ;
  assign y6904 = ~n9270 ;
  assign y6905 = n9276 ;
  assign y6906 = ~n9280 ;
  assign y6907 = ~n9282 ;
  assign y6908 = ~1'b0 ;
  assign y6909 = ~1'b0 ;
  assign y6910 = n9284 ;
  assign y6911 = n9004 ;
  assign y6912 = ~1'b0 ;
  assign y6913 = ~n2967 ;
  assign y6914 = ~n9286 ;
  assign y6915 = ~1'b0 ;
  assign y6916 = n9287 ;
  assign y6917 = ~n9289 ;
  assign y6918 = ~1'b0 ;
  assign y6919 = n9290 ;
  assign y6920 = ~n9294 ;
  assign y6921 = ~n9296 ;
  assign y6922 = n3007 ;
  assign y6923 = ~n9298 ;
  assign y6924 = ~1'b0 ;
  assign y6925 = ~n9299 ;
  assign y6926 = n9302 ;
  assign y6927 = n9304 ;
  assign y6928 = ~n9309 ;
  assign y6929 = ~1'b0 ;
  assign y6930 = n9313 ;
  assign y6931 = ~n9316 ;
  assign y6932 = ~1'b0 ;
  assign y6933 = ~n9322 ;
  assign y6934 = ~n7674 ;
  assign y6935 = n9325 ;
  assign y6936 = n9327 ;
  assign y6937 = ~n9332 ;
  assign y6938 = ~1'b0 ;
  assign y6939 = ~n9334 ;
  assign y6940 = ~n9335 ;
  assign y6941 = ~n9347 ;
  assign y6942 = ~1'b0 ;
  assign y6943 = n9348 ;
  assign y6944 = n9350 ;
  assign y6945 = ~n9355 ;
  assign y6946 = ~n9359 ;
  assign y6947 = ~1'b0 ;
  assign y6948 = n9360 ;
  assign y6949 = n9363 ;
  assign y6950 = ~n9368 ;
  assign y6951 = n3007 ;
  assign y6952 = ~1'b0 ;
  assign y6953 = n9370 ;
  assign y6954 = ~1'b0 ;
  assign y6955 = n9372 ;
  assign y6956 = ~1'b0 ;
  assign y6957 = ~1'b0 ;
  assign y6958 = ~1'b0 ;
  assign y6959 = n9373 ;
  assign y6960 = ~1'b0 ;
  assign y6961 = ~1'b0 ;
  assign y6962 = n9374 ;
  assign y6963 = ~1'b0 ;
  assign y6964 = ~1'b0 ;
  assign y6965 = ~1'b0 ;
  assign y6966 = 1'b0 ;
  assign y6967 = ~1'b0 ;
  assign y6968 = n9379 ;
  assign y6969 = 1'b0 ;
  assign y6970 = n9381 ;
  assign y6971 = n9384 ;
  assign y6972 = ~1'b0 ;
  assign y6973 = ~n2254 ;
  assign y6974 = ~1'b0 ;
  assign y6975 = n9385 ;
  assign y6976 = ~n376 ;
  assign y6977 = ~1'b0 ;
  assign y6978 = ~1'b0 ;
  assign y6979 = ~1'b0 ;
  assign y6980 = ~1'b0 ;
  assign y6981 = ~n9394 ;
  assign y6982 = n9396 ;
  assign y6983 = ~n9397 ;
  assign y6984 = n9402 ;
  assign y6985 = n9406 ;
  assign y6986 = 1'b0 ;
  assign y6987 = ~n9408 ;
  assign y6988 = ~1'b0 ;
  assign y6989 = ~1'b0 ;
  assign y6990 = ~n9409 ;
  assign y6991 = ~1'b0 ;
  assign y6992 = ~n9411 ;
  assign y6993 = ~1'b0 ;
  assign y6994 = ~1'b0 ;
  assign y6995 = ~1'b0 ;
  assign y6996 = ~1'b0 ;
  assign y6997 = ~n9412 ;
  assign y6998 = ~n9413 ;
  assign y6999 = ~1'b0 ;
  assign y7000 = ~1'b0 ;
  assign y7001 = n9414 ;
  assign y7002 = ~n9416 ;
  assign y7003 = ~1'b0 ;
  assign y7004 = ~n9419 ;
  assign y7005 = ~1'b0 ;
  assign y7006 = n9420 ;
  assign y7007 = ~1'b0 ;
  assign y7008 = ~1'b0 ;
  assign y7009 = ~1'b0 ;
  assign y7010 = ~n9424 ;
  assign y7011 = n9425 ;
  assign y7012 = n1947 ;
  assign y7013 = n116 ;
  assign y7014 = 1'b0 ;
  assign y7015 = ~1'b0 ;
  assign y7016 = ~n9432 ;
  assign y7017 = ~1'b0 ;
  assign y7018 = n3845 ;
  assign y7019 = ~1'b0 ;
  assign y7020 = ~n9434 ;
  assign y7021 = ~n9442 ;
  assign y7022 = ~n9444 ;
  assign y7023 = ~n9446 ;
  assign y7024 = 1'b0 ;
  assign y7025 = ~1'b0 ;
  assign y7026 = ~1'b0 ;
  assign y7027 = ~n3569 ;
  assign y7028 = ~1'b0 ;
  assign y7029 = ~1'b0 ;
  assign y7030 = ~1'b0 ;
  assign y7031 = ~n9447 ;
  assign y7032 = n9448 ;
  assign y7033 = ~1'b0 ;
  assign y7034 = ~1'b0 ;
  assign y7035 = ~1'b0 ;
  assign y7036 = 1'b0 ;
  assign y7037 = n9451 ;
  assign y7038 = n9452 ;
  assign y7039 = n9471 ;
  assign y7040 = ~1'b0 ;
  assign y7041 = n9479 ;
  assign y7042 = n9483 ;
  assign y7043 = ~1'b0 ;
  assign y7044 = ~1'b0 ;
  assign y7045 = ~1'b0 ;
  assign y7046 = n9490 ;
  assign y7047 = ~1'b0 ;
  assign y7048 = ~n8107 ;
  assign y7049 = 1'b0 ;
  assign y7050 = ~n9491 ;
  assign y7051 = ~1'b0 ;
  assign y7052 = ~n2681 ;
  assign y7053 = n9495 ;
  assign y7054 = ~n9496 ;
  assign y7055 = ~n4533 ;
  assign y7056 = n9498 ;
  assign y7057 = ~1'b0 ;
  assign y7058 = 1'b0 ;
  assign y7059 = n9502 ;
  assign y7060 = ~1'b0 ;
  assign y7061 = n9506 ;
  assign y7062 = ~n9507 ;
  assign y7063 = n1730 ;
  assign y7064 = ~1'b0 ;
  assign y7065 = n9510 ;
  assign y7066 = ~1'b0 ;
  assign y7067 = 1'b0 ;
  assign y7068 = 1'b0 ;
  assign y7069 = ~n9512 ;
  assign y7070 = ~n9514 ;
  assign y7071 = ~n9516 ;
  assign y7072 = ~n9518 ;
  assign y7073 = ~1'b0 ;
  assign y7074 = ~n9520 ;
  assign y7075 = 1'b0 ;
  assign y7076 = ~1'b0 ;
  assign y7077 = ~n9521 ;
  assign y7078 = ~n9523 ;
  assign y7079 = ~1'b0 ;
  assign y7080 = ~n3822 ;
  assign y7081 = ~n9524 ;
  assign y7082 = ~1'b0 ;
  assign y7083 = ~n9527 ;
  assign y7084 = ~1'b0 ;
  assign y7085 = n9528 ;
  assign y7086 = ~n3946 ;
  assign y7087 = ~n9530 ;
  assign y7088 = ~1'b0 ;
  assign y7089 = ~n9536 ;
  assign y7090 = ~1'b0 ;
  assign y7091 = n9542 ;
  assign y7092 = ~n9545 ;
  assign y7093 = ~1'b0 ;
  assign y7094 = ~n9546 ;
  assign y7095 = n9548 ;
  assign y7096 = ~n9549 ;
  assign y7097 = ~1'b0 ;
  assign y7098 = ~1'b0 ;
  assign y7099 = ~1'b0 ;
  assign y7100 = ~n9550 ;
  assign y7101 = ~1'b0 ;
  assign y7102 = ~n9551 ;
  assign y7103 = ~1'b0 ;
  assign y7104 = 1'b0 ;
  assign y7105 = n9552 ;
  assign y7106 = 1'b0 ;
  assign y7107 = ~n9557 ;
  assign y7108 = n9559 ;
  assign y7109 = ~n9561 ;
  assign y7110 = n9562 ;
  assign y7111 = ~n9564 ;
  assign y7112 = ~n9569 ;
  assign y7113 = n9401 ;
  assign y7114 = ~n9571 ;
  assign y7115 = ~1'b0 ;
  assign y7116 = ~1'b0 ;
  assign y7117 = n9572 ;
  assign y7118 = ~1'b0 ;
  assign y7119 = ~1'b0 ;
  assign y7120 = 1'b0 ;
  assign y7121 = ~1'b0 ;
  assign y7122 = ~n9573 ;
  assign y7123 = ~n216 ;
  assign y7124 = ~n9575 ;
  assign y7125 = 1'b0 ;
  assign y7126 = ~n895 ;
  assign y7127 = n9576 ;
  assign y7128 = ~n9578 ;
  assign y7129 = ~n9580 ;
  assign y7130 = ~n9581 ;
  assign y7131 = 1'b0 ;
  assign y7132 = ~n4449 ;
  assign y7133 = n9583 ;
  assign y7134 = ~1'b0 ;
  assign y7135 = n9586 ;
  assign y7136 = ~n2905 ;
  assign y7137 = ~n9589 ;
  assign y7138 = ~1'b0 ;
  assign y7139 = ~1'b0 ;
  assign y7140 = ~1'b0 ;
  assign y7141 = ~1'b0 ;
  assign y7142 = ~n9590 ;
  assign y7143 = ~n9591 ;
  assign y7144 = ~n3206 ;
  assign y7145 = n9594 ;
  assign y7146 = ~1'b0 ;
  assign y7147 = n9595 ;
  assign y7148 = ~n9596 ;
  assign y7149 = ~n9597 ;
  assign y7150 = n9602 ;
  assign y7151 = n9606 ;
  assign y7152 = n9610 ;
  assign y7153 = ~1'b0 ;
  assign y7154 = n9611 ;
  assign y7155 = ~1'b0 ;
  assign y7156 = ~n9613 ;
  assign y7157 = ~1'b0 ;
  assign y7158 = ~1'b0 ;
  assign y7159 = n9614 ;
  assign y7160 = ~1'b0 ;
  assign y7161 = n5952 ;
  assign y7162 = ~1'b0 ;
  assign y7163 = n9616 ;
  assign y7164 = n9617 ;
  assign y7165 = n9620 ;
  assign y7166 = ~1'b0 ;
  assign y7167 = ~1'b0 ;
  assign y7168 = ~1'b0 ;
  assign y7169 = ~n9623 ;
  assign y7170 = ~1'b0 ;
  assign y7171 = n9625 ;
  assign y7172 = 1'b0 ;
  assign y7173 = ~1'b0 ;
  assign y7174 = ~1'b0 ;
  assign y7175 = 1'b0 ;
  assign y7176 = n9626 ;
  assign y7177 = n163 ;
  assign y7178 = ~1'b0 ;
  assign y7179 = n9634 ;
  assign y7180 = n9638 ;
  assign y7181 = ~n273 ;
  assign y7182 = ~n9643 ;
  assign y7183 = ~1'b0 ;
  assign y7184 = ~1'b0 ;
  assign y7185 = ~1'b0 ;
  assign y7186 = 1'b0 ;
  assign y7187 = n1620 ;
  assign y7188 = n9645 ;
  assign y7189 = n9646 ;
  assign y7190 = ~1'b0 ;
  assign y7191 = ~n9647 ;
  assign y7192 = n9651 ;
  assign y7193 = ~1'b0 ;
  assign y7194 = n3382 ;
  assign y7195 = ~1'b0 ;
  assign y7196 = ~n6944 ;
  assign y7197 = n9652 ;
  assign y7198 = ~1'b0 ;
  assign y7199 = ~1'b0 ;
  assign y7200 = ~n9657 ;
  assign y7201 = n9659 ;
  assign y7202 = n9660 ;
  assign y7203 = ~1'b0 ;
  assign y7204 = n9661 ;
  assign y7205 = ~n9662 ;
  assign y7206 = ~n9663 ;
  assign y7207 = ~1'b0 ;
  assign y7208 = 1'b0 ;
  assign y7209 = ~n9668 ;
  assign y7210 = 1'b0 ;
  assign y7211 = ~1'b0 ;
  assign y7212 = ~n9672 ;
  assign y7213 = n9677 ;
  assign y7214 = ~1'b0 ;
  assign y7215 = n4196 ;
  assign y7216 = 1'b0 ;
  assign y7217 = n9684 ;
  assign y7218 = n9689 ;
  assign y7219 = ~1'b0 ;
  assign y7220 = ~1'b0 ;
  assign y7221 = ~1'b0 ;
  assign y7222 = ~n9691 ;
  assign y7223 = ~1'b0 ;
  assign y7224 = ~n9696 ;
  assign y7225 = ~n9698 ;
  assign y7226 = ~n9702 ;
  assign y7227 = n9703 ;
  assign y7228 = ~1'b0 ;
  assign y7229 = ~n9705 ;
  assign y7230 = n9712 ;
  assign y7231 = ~1'b0 ;
  assign y7232 = ~1'b0 ;
  assign y7233 = ~n9713 ;
  assign y7234 = n3265 ;
  assign y7235 = n9715 ;
  assign y7236 = ~n9717 ;
  assign y7237 = n9718 ;
  assign y7238 = ~1'b0 ;
  assign y7239 = ~n512 ;
  assign y7240 = n9722 ;
  assign y7241 = ~1'b0 ;
  assign y7242 = n470 ;
  assign y7243 = ~1'b0 ;
  assign y7244 = n1246 ;
  assign y7245 = n9723 ;
  assign y7246 = ~1'b0 ;
  assign y7247 = ~n9725 ;
  assign y7248 = 1'b0 ;
  assign y7249 = ~1'b0 ;
  assign y7250 = 1'b0 ;
  assign y7251 = n5388 ;
  assign y7252 = ~1'b0 ;
  assign y7253 = ~n9726 ;
  assign y7254 = ~n9727 ;
  assign y7255 = n5971 ;
  assign y7256 = ~1'b0 ;
  assign y7257 = 1'b0 ;
  assign y7258 = ~n9730 ;
  assign y7259 = n4412 ;
  assign y7260 = n9733 ;
  assign y7261 = n9736 ;
  assign y7262 = 1'b0 ;
  assign y7263 = n9737 ;
  assign y7264 = n4322 ;
  assign y7265 = ~n9741 ;
  assign y7266 = ~1'b0 ;
  assign y7267 = n9743 ;
  assign y7268 = ~n9744 ;
  assign y7269 = 1'b0 ;
  assign y7270 = ~n461 ;
  assign y7271 = n9746 ;
  assign y7272 = ~n9751 ;
  assign y7273 = ~n9754 ;
  assign y7274 = ~n9756 ;
  assign y7275 = ~n9757 ;
  assign y7276 = 1'b0 ;
  assign y7277 = ~n9759 ;
  assign y7278 = n9760 ;
  assign y7279 = ~1'b0 ;
  assign y7280 = ~n9764 ;
  assign y7281 = n9765 ;
  assign y7282 = n9770 ;
  assign y7283 = ~n9771 ;
  assign y7284 = ~n9776 ;
  assign y7285 = ~n9778 ;
  assign y7286 = n9781 ;
  assign y7287 = ~1'b0 ;
  assign y7288 = n9787 ;
  assign y7289 = n9789 ;
  assign y7290 = ~1'b0 ;
  assign y7291 = n4784 ;
  assign y7292 = ~1'b0 ;
  assign y7293 = ~n9791 ;
  assign y7294 = ~n9793 ;
  assign y7295 = n9794 ;
  assign y7296 = ~n5871 ;
  assign y7297 = n9796 ;
  assign y7298 = ~n9799 ;
  assign y7299 = ~1'b0 ;
  assign y7300 = ~1'b0 ;
  assign y7301 = n9801 ;
  assign y7302 = ~1'b0 ;
  assign y7303 = n9802 ;
  assign y7304 = ~n9805 ;
  assign y7305 = ~1'b0 ;
  assign y7306 = n9806 ;
  assign y7307 = ~1'b0 ;
  assign y7308 = ~1'b0 ;
  assign y7309 = ~1'b0 ;
  assign y7310 = ~1'b0 ;
  assign y7311 = ~1'b0 ;
  assign y7312 = ~n9810 ;
  assign y7313 = ~1'b0 ;
  assign y7314 = ~n9814 ;
  assign y7315 = n715 ;
  assign y7316 = n9816 ;
  assign y7317 = ~n9817 ;
  assign y7318 = n9822 ;
  assign y7319 = n9824 ;
  assign y7320 = ~1'b0 ;
  assign y7321 = ~n9827 ;
  assign y7322 = n9828 ;
  assign y7323 = ~n8581 ;
  assign y7324 = ~n9829 ;
  assign y7325 = ~n9835 ;
  assign y7326 = ~n3670 ;
  assign y7327 = n9836 ;
  assign y7328 = ~n6025 ;
  assign y7329 = ~n9838 ;
  assign y7330 = ~1'b0 ;
  assign y7331 = ~1'b0 ;
  assign y7332 = n9841 ;
  assign y7333 = ~1'b0 ;
  assign y7334 = ~1'b0 ;
  assign y7335 = ~1'b0 ;
  assign y7336 = ~1'b0 ;
  assign y7337 = ~1'b0 ;
  assign y7338 = n9843 ;
  assign y7339 = ~1'b0 ;
  assign y7340 = ~n9845 ;
  assign y7341 = ~n9848 ;
  assign y7342 = ~1'b0 ;
  assign y7343 = ~n9850 ;
  assign y7344 = ~n9851 ;
  assign y7345 = ~1'b0 ;
  assign y7346 = ~1'b0 ;
  assign y7347 = ~1'b0 ;
  assign y7348 = n9852 ;
  assign y7349 = ~n9855 ;
  assign y7350 = ~n9857 ;
  assign y7351 = n9858 ;
  assign y7352 = n9859 ;
  assign y7353 = ~1'b0 ;
  assign y7354 = n278 ;
  assign y7355 = n4623 ;
  assign y7356 = ~n7442 ;
  assign y7357 = ~n9862 ;
  assign y7358 = ~n9867 ;
  assign y7359 = n9868 ;
  assign y7360 = n9870 ;
  assign y7361 = n9872 ;
  assign y7362 = ~1'b0 ;
  assign y7363 = ~1'b0 ;
  assign y7364 = ~1'b0 ;
  assign y7365 = ~1'b0 ;
  assign y7366 = ~1'b0 ;
  assign y7367 = ~1'b0 ;
  assign y7368 = ~1'b0 ;
  assign y7369 = n9873 ;
  assign y7370 = ~1'b0 ;
  assign y7371 = ~n9880 ;
  assign y7372 = ~n9882 ;
  assign y7373 = n1690 ;
  assign y7374 = ~n9883 ;
  assign y7375 = n9884 ;
  assign y7376 = n9888 ;
  assign y7377 = n9890 ;
  assign y7378 = n9892 ;
  assign y7379 = ~1'b0 ;
  assign y7380 = ~n9894 ;
  assign y7381 = n9895 ;
  assign y7382 = ~n9899 ;
  assign y7383 = n9900 ;
  assign y7384 = ~1'b0 ;
  assign y7385 = n9901 ;
  assign y7386 = ~n3507 ;
  assign y7387 = n9905 ;
  assign y7388 = n9910 ;
  assign y7389 = ~n9922 ;
  assign y7390 = n9923 ;
  assign y7391 = ~n5972 ;
  assign y7392 = ~1'b0 ;
  assign y7393 = ~n9930 ;
  assign y7394 = n9931 ;
  assign y7395 = n9934 ;
  assign y7396 = ~1'b0 ;
  assign y7397 = ~1'b0 ;
  assign y7398 = n4246 ;
  assign y7399 = ~n9935 ;
  assign y7400 = n9940 ;
  assign y7401 = n9941 ;
  assign y7402 = ~1'b0 ;
  assign y7403 = n9942 ;
  assign y7404 = ~1'b0 ;
  assign y7405 = ~1'b0 ;
  assign y7406 = n3793 ;
  assign y7407 = ~1'b0 ;
  assign y7408 = n30 ;
  assign y7409 = n9951 ;
  assign y7410 = n9955 ;
  assign y7411 = ~n9957 ;
  assign y7412 = ~1'b0 ;
  assign y7413 = n9959 ;
  assign y7414 = ~n9961 ;
  assign y7415 = ~1'b0 ;
  assign y7416 = n9964 ;
  assign y7417 = ~1'b0 ;
  assign y7418 = ~n9965 ;
  assign y7419 = ~1'b0 ;
  assign y7420 = ~n9966 ;
  assign y7421 = n9969 ;
  assign y7422 = ~1'b0 ;
  assign y7423 = ~1'b0 ;
  assign y7424 = n4799 ;
  assign y7425 = ~n9971 ;
  assign y7426 = ~1'b0 ;
  assign y7427 = ~n9979 ;
  assign y7428 = ~1'b0 ;
  assign y7429 = ~1'b0 ;
  assign y7430 = ~1'b0 ;
  assign y7431 = 1'b0 ;
  assign y7432 = ~1'b0 ;
  assign y7433 = n8617 ;
  assign y7434 = ~1'b0 ;
  assign y7435 = n9981 ;
  assign y7436 = n9982 ;
  assign y7437 = ~1'b0 ;
  assign y7438 = n5131 ;
  assign y7439 = ~n9983 ;
  assign y7440 = ~n9985 ;
  assign y7441 = n9987 ;
  assign y7442 = 1'b0 ;
  assign y7443 = ~n9988 ;
  assign y7444 = ~1'b0 ;
  assign y7445 = ~1'b0 ;
  assign y7446 = ~1'b0 ;
  assign y7447 = ~n9989 ;
  assign y7448 = ~n9990 ;
  assign y7449 = n9991 ;
  assign y7450 = n9992 ;
  assign y7451 = n9996 ;
  assign y7452 = n9998 ;
  assign y7453 = ~1'b0 ;
  assign y7454 = ~n9999 ;
  assign y7455 = n10000 ;
  assign y7456 = ~1'b0 ;
  assign y7457 = n10005 ;
  assign y7458 = ~1'b0 ;
  assign y7459 = 1'b0 ;
  assign y7460 = ~n10011 ;
  assign y7461 = n10018 ;
  assign y7462 = n10024 ;
  assign y7463 = ~n10026 ;
  assign y7464 = n10030 ;
  assign y7465 = ~n7488 ;
  assign y7466 = ~1'b0 ;
  assign y7467 = n10031 ;
  assign y7468 = ~1'b0 ;
  assign y7469 = n10032 ;
  assign y7470 = ~n10036 ;
  assign y7471 = ~1'b0 ;
  assign y7472 = ~n10040 ;
  assign y7473 = ~1'b0 ;
  assign y7474 = ~1'b0 ;
  assign y7475 = n10041 ;
  assign y7476 = ~n3718 ;
  assign y7477 = ~n10043 ;
  assign y7478 = ~n10044 ;
  assign y7479 = n10046 ;
  assign y7480 = 1'b0 ;
  assign y7481 = ~n10047 ;
  assign y7482 = n10048 ;
  assign y7483 = ~n10052 ;
  assign y7484 = n8829 ;
  assign y7485 = ~1'b0 ;
  assign y7486 = ~n10053 ;
  assign y7487 = ~1'b0 ;
  assign y7488 = n10055 ;
  assign y7489 = ~1'b0 ;
  assign y7490 = ~n10056 ;
  assign y7491 = n4580 ;
  assign y7492 = ~n10059 ;
  assign y7493 = n10060 ;
  assign y7494 = n10063 ;
  assign y7495 = ~1'b0 ;
  assign y7496 = 1'b0 ;
  assign y7497 = n10064 ;
  assign y7498 = ~1'b0 ;
  assign y7499 = ~n10066 ;
  assign y7500 = ~1'b0 ;
  assign y7501 = ~n10067 ;
  assign y7502 = ~1'b0 ;
  assign y7503 = ~n4551 ;
  assign y7504 = n10069 ;
  assign y7505 = ~n10071 ;
  assign y7506 = n10076 ;
  assign y7507 = n1227 ;
  assign y7508 = ~n10077 ;
  assign y7509 = n10078 ;
  assign y7510 = ~n10080 ;
  assign y7511 = n9221 ;
  assign y7512 = ~1'b0 ;
  assign y7513 = ~1'b0 ;
  assign y7514 = ~n10083 ;
  assign y7515 = ~n10085 ;
  assign y7516 = n10086 ;
  assign y7517 = n2109 ;
  assign y7518 = 1'b0 ;
  assign y7519 = ~n10089 ;
  assign y7520 = n10092 ;
  assign y7521 = n1067 ;
  assign y7522 = ~n10096 ;
  assign y7523 = ~n1555 ;
  assign y7524 = ~1'b0 ;
  assign y7525 = ~n10099 ;
  assign y7526 = ~n4404 ;
  assign y7527 = 1'b0 ;
  assign y7528 = ~1'b0 ;
  assign y7529 = ~n10100 ;
  assign y7530 = ~1'b0 ;
  assign y7531 = ~1'b0 ;
  assign y7532 = ~n10101 ;
  assign y7533 = ~1'b0 ;
  assign y7534 = ~n6001 ;
  assign y7535 = ~1'b0 ;
  assign y7536 = 1'b0 ;
  assign y7537 = n10104 ;
  assign y7538 = ~n10106 ;
  assign y7539 = ~1'b0 ;
  assign y7540 = n10112 ;
  assign y7541 = ~n10113 ;
  assign y7542 = n10115 ;
  assign y7543 = ~n10118 ;
  assign y7544 = n10119 ;
  assign y7545 = ~1'b0 ;
  assign y7546 = n6764 ;
  assign y7547 = 1'b0 ;
  assign y7548 = n10123 ;
  assign y7549 = ~1'b0 ;
  assign y7550 = ~1'b0 ;
  assign y7551 = ~n10126 ;
  assign y7552 = n10128 ;
  assign y7553 = n727 ;
  assign y7554 = ~n1957 ;
  assign y7555 = ~1'b0 ;
  assign y7556 = ~n10131 ;
  assign y7557 = n10133 ;
  assign y7558 = ~n10134 ;
  assign y7559 = n6150 ;
  assign y7560 = n10137 ;
  assign y7561 = ~1'b0 ;
  assign y7562 = n10144 ;
  assign y7563 = ~1'b0 ;
  assign y7564 = ~n10149 ;
  assign y7565 = ~n10151 ;
  assign y7566 = n10155 ;
  assign y7567 = ~n2148 ;
  assign y7568 = 1'b0 ;
  assign y7569 = ~n10156 ;
  assign y7570 = n10157 ;
  assign y7571 = n8031 ;
  assign y7572 = ~1'b0 ;
  assign y7573 = 1'b0 ;
  assign y7574 = n3965 ;
  assign y7575 = ~1'b0 ;
  assign y7576 = ~1'b0 ;
  assign y7577 = ~1'b0 ;
  assign y7578 = ~n10159 ;
  assign y7579 = n10163 ;
  assign y7580 = ~1'b0 ;
  assign y7581 = ~1'b0 ;
  assign y7582 = ~n10165 ;
  assign y7583 = n10167 ;
  assign y7584 = n10168 ;
  assign y7585 = n10171 ;
  assign y7586 = ~n144 ;
  assign y7587 = ~1'b0 ;
  assign y7588 = n10175 ;
  assign y7589 = ~1'b0 ;
  assign y7590 = ~1'b0 ;
  assign y7591 = ~n10177 ;
  assign y7592 = ~n10178 ;
  assign y7593 = ~1'b0 ;
  assign y7594 = ~n389 ;
  assign y7595 = ~n10180 ;
  assign y7596 = ~n10182 ;
  assign y7597 = n10188 ;
  assign y7598 = n10192 ;
  assign y7599 = ~n10193 ;
  assign y7600 = n2686 ;
  assign y7601 = n10195 ;
  assign y7602 = n10200 ;
  assign y7603 = n10201 ;
  assign y7604 = ~n10202 ;
  assign y7605 = ~1'b0 ;
  assign y7606 = ~n10206 ;
  assign y7607 = n10208 ;
  assign y7608 = ~n7639 ;
  assign y7609 = n10210 ;
  assign y7610 = ~1'b0 ;
  assign y7611 = 1'b0 ;
  assign y7612 = n715 ;
  assign y7613 = ~n10212 ;
  assign y7614 = ~1'b0 ;
  assign y7615 = n10216 ;
  assign y7616 = ~1'b0 ;
  assign y7617 = n2919 ;
  assign y7618 = ~1'b0 ;
  assign y7619 = ~n10223 ;
  assign y7620 = n10224 ;
  assign y7621 = n10226 ;
  assign y7622 = ~1'b0 ;
  assign y7623 = n1209 ;
  assign y7624 = ~n10229 ;
  assign y7625 = ~1'b0 ;
  assign y7626 = ~1'b0 ;
  assign y7627 = ~n10233 ;
  assign y7628 = ~n10241 ;
  assign y7629 = ~n10246 ;
  assign y7630 = ~1'b0 ;
  assign y7631 = ~1'b0 ;
  assign y7632 = ~n10247 ;
  assign y7633 = ~n10251 ;
  assign y7634 = n10252 ;
  assign y7635 = n7955 ;
  assign y7636 = ~n10253 ;
  assign y7637 = ~n10260 ;
  assign y7638 = ~n10264 ;
  assign y7639 = ~1'b0 ;
  assign y7640 = ~1'b0 ;
  assign y7641 = ~n6481 ;
  assign y7642 = ~1'b0 ;
  assign y7643 = ~1'b0 ;
  assign y7644 = ~1'b0 ;
  assign y7645 = ~n10266 ;
  assign y7646 = n10267 ;
  assign y7647 = n10268 ;
  assign y7648 = ~n10269 ;
  assign y7649 = n10280 ;
  assign y7650 = ~1'b0 ;
  assign y7651 = n9029 ;
  assign y7652 = ~n10282 ;
  assign y7653 = ~n10284 ;
  assign y7654 = n10285 ;
  assign y7655 = ~n10286 ;
  assign y7656 = ~1'b0 ;
  assign y7657 = n10289 ;
  assign y7658 = n10292 ;
  assign y7659 = n10296 ;
  assign y7660 = n10298 ;
  assign y7661 = ~n10307 ;
  assign y7662 = ~n3670 ;
  assign y7663 = ~1'b0 ;
  assign y7664 = ~n10310 ;
  assign y7665 = ~1'b0 ;
  assign y7666 = n10312 ;
  assign y7667 = 1'b0 ;
  assign y7668 = ~n10313 ;
  assign y7669 = n10318 ;
  assign y7670 = ~1'b0 ;
  assign y7671 = ~n10320 ;
  assign y7672 = ~n10321 ;
  assign y7673 = n3581 ;
  assign y7674 = ~n10322 ;
  assign y7675 = n10323 ;
  assign y7676 = ~n10325 ;
  assign y7677 = ~1'b0 ;
  assign y7678 = ~n10328 ;
  assign y7679 = ~1'b0 ;
  assign y7680 = ~n10329 ;
  assign y7681 = ~1'b0 ;
  assign y7682 = ~1'b0 ;
  assign y7683 = ~n10330 ;
  assign y7684 = ~1'b0 ;
  assign y7685 = ~1'b0 ;
  assign y7686 = ~n10333 ;
  assign y7687 = 1'b0 ;
  assign y7688 = ~n10105 ;
  assign y7689 = ~1'b0 ;
  assign y7690 = ~1'b0 ;
  assign y7691 = ~n10335 ;
  assign y7692 = ~1'b0 ;
  assign y7693 = ~1'b0 ;
  assign y7694 = n3483 ;
  assign y7695 = ~1'b0 ;
  assign y7696 = ~1'b0 ;
  assign y7697 = ~1'b0 ;
  assign y7698 = ~n10338 ;
  assign y7699 = ~1'b0 ;
  assign y7700 = ~1'b0 ;
  assign y7701 = ~n10339 ;
  assign y7702 = 1'b0 ;
  assign y7703 = n10343 ;
  assign y7704 = ~1'b0 ;
  assign y7705 = ~n10345 ;
  assign y7706 = ~n10348 ;
  assign y7707 = ~1'b0 ;
  assign y7708 = ~n10349 ;
  assign y7709 = ~1'b0 ;
  assign y7710 = n10352 ;
  assign y7711 = ~1'b0 ;
  assign y7712 = ~n10355 ;
  assign y7713 = ~n10356 ;
  assign y7714 = n10357 ;
  assign y7715 = ~n10360 ;
  assign y7716 = ~n3708 ;
  assign y7717 = ~n10361 ;
  assign y7718 = n10367 ;
  assign y7719 = ~n10369 ;
  assign y7720 = ~1'b0 ;
  assign y7721 = ~n10370 ;
  assign y7722 = n10372 ;
  assign y7723 = ~n10374 ;
  assign y7724 = ~1'b0 ;
  assign y7725 = ~1'b0 ;
  assign y7726 = n3295 ;
  assign y7727 = ~n10378 ;
  assign y7728 = n10379 ;
  assign y7729 = ~n10382 ;
  assign y7730 = ~n8326 ;
  assign y7731 = ~n1232 ;
  assign y7732 = ~n8322 ;
  assign y7733 = ~1'b0 ;
  assign y7734 = n10384 ;
  assign y7735 = n10387 ;
  assign y7736 = n10390 ;
  assign y7737 = ~n10391 ;
  assign y7738 = n10393 ;
  assign y7739 = ~n10399 ;
  assign y7740 = ~1'b0 ;
  assign y7741 = n10401 ;
  assign y7742 = 1'b0 ;
  assign y7743 = ~1'b0 ;
  assign y7744 = ~n10405 ;
  assign y7745 = ~n10414 ;
  assign y7746 = ~1'b0 ;
  assign y7747 = ~1'b0 ;
  assign y7748 = n10419 ;
  assign y7749 = n10420 ;
  assign y7750 = n10422 ;
  assign y7751 = ~1'b0 ;
  assign y7752 = ~n10423 ;
  assign y7753 = ~1'b0 ;
  assign y7754 = n4855 ;
  assign y7755 = ~1'b0 ;
  assign y7756 = 1'b0 ;
  assign y7757 = n10424 ;
  assign y7758 = ~n4449 ;
  assign y7759 = ~n1165 ;
  assign y7760 = ~n10426 ;
  assign y7761 = n10428 ;
  assign y7762 = n940 ;
  assign y7763 = ~n10430 ;
  assign y7764 = ~n10432 ;
  assign y7765 = ~1'b0 ;
  assign y7766 = ~1'b0 ;
  assign y7767 = ~1'b0 ;
  assign y7768 = n1165 ;
  assign y7769 = n10434 ;
  assign y7770 = ~1'b0 ;
  assign y7771 = n9055 ;
  assign y7772 = n10439 ;
  assign y7773 = n10444 ;
  assign y7774 = n10448 ;
  assign y7775 = n10449 ;
  assign y7776 = n10459 ;
  assign y7777 = ~n10463 ;
  assign y7778 = ~1'b0 ;
  assign y7779 = n10472 ;
  assign y7780 = ~1'b0 ;
  assign y7781 = ~1'b0 ;
  assign y7782 = n9954 ;
  assign y7783 = ~n10479 ;
  assign y7784 = ~n10480 ;
  assign y7785 = 1'b0 ;
  assign y7786 = n10482 ;
  assign y7787 = ~n10487 ;
  assign y7788 = n10489 ;
  assign y7789 = n10490 ;
  assign y7790 = ~1'b0 ;
  assign y7791 = n10492 ;
  assign y7792 = ~1'b0 ;
  assign y7793 = n1370 ;
  assign y7794 = ~1'b0 ;
  assign y7795 = n10493 ;
  assign y7796 = ~1'b0 ;
  assign y7797 = ~1'b0 ;
  assign y7798 = 1'b0 ;
  assign y7799 = n10495 ;
  assign y7800 = ~n10499 ;
  assign y7801 = n10500 ;
  assign y7802 = ~n10502 ;
  assign y7803 = ~1'b0 ;
  assign y7804 = n10507 ;
  assign y7805 = 1'b0 ;
  assign y7806 = n10508 ;
  assign y7807 = ~1'b0 ;
  assign y7808 = ~1'b0 ;
  assign y7809 = ~n10509 ;
  assign y7810 = ~n5559 ;
  assign y7811 = n10512 ;
  assign y7812 = ~n10514 ;
  assign y7813 = n6191 ;
  assign y7814 = ~n10517 ;
  assign y7815 = n10519 ;
  assign y7816 = ~1'b0 ;
  assign y7817 = n10523 ;
  assign y7818 = ~1'b0 ;
  assign y7819 = 1'b0 ;
  assign y7820 = ~1'b0 ;
  assign y7821 = ~n7377 ;
  assign y7822 = ~1'b0 ;
  assign y7823 = n10524 ;
  assign y7824 = 1'b0 ;
  assign y7825 = ~1'b0 ;
  assign y7826 = 1'b0 ;
  assign y7827 = ~1'b0 ;
  assign y7828 = ~1'b0 ;
  assign y7829 = ~1'b0 ;
  assign y7830 = 1'b0 ;
  assign y7831 = ~1'b0 ;
  assign y7832 = ~n10530 ;
  assign y7833 = n10531 ;
  assign y7834 = n10532 ;
  assign y7835 = ~1'b0 ;
  assign y7836 = ~n10533 ;
  assign y7837 = n10534 ;
  assign y7838 = ~n10535 ;
  assign y7839 = ~1'b0 ;
  assign y7840 = ~1'b0 ;
  assign y7841 = 1'b0 ;
  assign y7842 = ~n10536 ;
  assign y7843 = n6709 ;
  assign y7844 = ~n10537 ;
  assign y7845 = n10538 ;
  assign y7846 = n10539 ;
  assign y7847 = n10541 ;
  assign y7848 = ~n1020 ;
  assign y7849 = n10543 ;
  assign y7850 = ~n10546 ;
  assign y7851 = ~n9697 ;
  assign y7852 = ~1'b0 ;
  assign y7853 = ~1'b0 ;
  assign y7854 = ~1'b0 ;
  assign y7855 = ~n8969 ;
  assign y7856 = ~1'b0 ;
  assign y7857 = n10547 ;
  assign y7858 = n3100 ;
  assign y7859 = ~1'b0 ;
  assign y7860 = ~n10553 ;
  assign y7861 = ~n10554 ;
  assign y7862 = ~n10560 ;
  assign y7863 = ~1'b0 ;
  assign y7864 = ~n10273 ;
  assign y7865 = ~n10565 ;
  assign y7866 = ~n4613 ;
  assign y7867 = n10569 ;
  assign y7868 = n10572 ;
  assign y7869 = ~n1637 ;
  assign y7870 = n10575 ;
  assign y7871 = n10576 ;
  assign y7872 = n3187 ;
  assign y7873 = ~1'b0 ;
  assign y7874 = n10579 ;
  assign y7875 = ~1'b0 ;
  assign y7876 = ~1'b0 ;
  assign y7877 = n10580 ;
  assign y7878 = ~1'b0 ;
  assign y7879 = n10583 ;
  assign y7880 = n10584 ;
  assign y7881 = ~n10586 ;
  assign y7882 = ~1'b0 ;
  assign y7883 = ~1'b0 ;
  assign y7884 = ~n10590 ;
  assign y7885 = ~1'b0 ;
  assign y7886 = ~n10591 ;
  assign y7887 = ~n10592 ;
  assign y7888 = ~n3608 ;
  assign y7889 = ~1'b0 ;
  assign y7890 = ~n10593 ;
  assign y7891 = ~n10598 ;
  assign y7892 = n10599 ;
  assign y7893 = ~1'b0 ;
  assign y7894 = ~n10603 ;
  assign y7895 = ~1'b0 ;
  assign y7896 = ~1'b0 ;
  assign y7897 = ~1'b0 ;
  assign y7898 = ~n10604 ;
  assign y7899 = n10605 ;
  assign y7900 = n10607 ;
  assign y7901 = ~1'b0 ;
  assign y7902 = n10608 ;
  assign y7903 = n10610 ;
  assign y7904 = ~n10612 ;
  assign y7905 = ~1'b0 ;
  assign y7906 = n10617 ;
  assign y7907 = ~n10619 ;
  assign y7908 = ~n10624 ;
  assign y7909 = ~1'b0 ;
  assign y7910 = n10630 ;
  assign y7911 = ~n10631 ;
  assign y7912 = ~1'b0 ;
  assign y7913 = n10632 ;
  assign y7914 = n10633 ;
  assign y7915 = 1'b0 ;
  assign y7916 = ~n10634 ;
  assign y7917 = ~1'b0 ;
  assign y7918 = ~n10637 ;
  assign y7919 = ~n10643 ;
  assign y7920 = ~n10644 ;
  assign y7921 = ~1'b0 ;
  assign y7922 = n10645 ;
  assign y7923 = ~n10646 ;
  assign y7924 = ~n10648 ;
  assign y7925 = ~1'b0 ;
  assign y7926 = ~n10653 ;
  assign y7927 = n10656 ;
  assign y7928 = 1'b0 ;
  assign y7929 = n1765 ;
  assign y7930 = 1'b0 ;
  assign y7931 = ~1'b0 ;
  assign y7932 = ~n10657 ;
  assign y7933 = ~n9499 ;
  assign y7934 = ~1'b0 ;
  assign y7935 = ~n1316 ;
  assign y7936 = ~1'b0 ;
  assign y7937 = ~n2943 ;
  assign y7938 = n10659 ;
  assign y7939 = ~1'b0 ;
  assign y7940 = n10661 ;
  assign y7941 = ~1'b0 ;
  assign y7942 = ~1'b0 ;
  assign y7943 = ~1'b0 ;
  assign y7944 = ~n10662 ;
  assign y7945 = ~n4126 ;
  assign y7946 = ~n10668 ;
  assign y7947 = ~1'b0 ;
  assign y7948 = ~n10670 ;
  assign y7949 = n10672 ;
  assign y7950 = ~1'b0 ;
  assign y7951 = n10673 ;
  assign y7952 = ~n10674 ;
  assign y7953 = n10675 ;
  assign y7954 = n10682 ;
  assign y7955 = ~n10686 ;
  assign y7956 = ~1'b0 ;
  assign y7957 = ~1'b0 ;
  assign y7958 = ~1'b0 ;
  assign y7959 = n10689 ;
  assign y7960 = ~1'b0 ;
  assign y7961 = ~n10692 ;
  assign y7962 = 1'b0 ;
  assign y7963 = n2449 ;
  assign y7964 = ~1'b0 ;
  assign y7965 = ~n3645 ;
  assign y7966 = ~n10704 ;
  assign y7967 = ~1'b0 ;
  assign y7968 = ~1'b0 ;
  assign y7969 = ~1'b0 ;
  assign y7970 = ~1'b0 ;
  assign y7971 = n10706 ;
  assign y7972 = ~1'b0 ;
  assign y7973 = n340 ;
  assign y7974 = n6419 ;
  assign y7975 = n10707 ;
  assign y7976 = ~1'b0 ;
  assign y7977 = n10658 ;
  assign y7978 = ~1'b0 ;
  assign y7979 = n6539 ;
  assign y7980 = n10708 ;
  assign y7981 = n10709 ;
  assign y7982 = ~n10717 ;
  assign y7983 = ~1'b0 ;
  assign y7984 = ~n10718 ;
  assign y7985 = ~1'b0 ;
  assign y7986 = ~n10719 ;
  assign y7987 = ~n10723 ;
  assign y7988 = ~1'b0 ;
  assign y7989 = ~1'b0 ;
  assign y7990 = ~1'b0 ;
  assign y7991 = n10727 ;
  assign y7992 = n10728 ;
  assign y7993 = ~1'b0 ;
  assign y7994 = n10729 ;
  assign y7995 = ~1'b0 ;
  assign y7996 = ~1'b0 ;
  assign y7997 = n10736 ;
  assign y7998 = ~n4840 ;
  assign y7999 = ~n10739 ;
  assign y8000 = ~1'b0 ;
  assign y8001 = ~1'b0 ;
  assign y8002 = ~1'b0 ;
  assign y8003 = ~1'b0 ;
  assign y8004 = ~n10740 ;
  assign y8005 = n10741 ;
  assign y8006 = n10743 ;
  assign y8007 = ~n10747 ;
  assign y8008 = n10751 ;
  assign y8009 = n10752 ;
  assign y8010 = ~1'b0 ;
  assign y8011 = n10755 ;
  assign y8012 = ~n10758 ;
  assign y8013 = n10761 ;
  assign y8014 = ~n10762 ;
  assign y8015 = ~1'b0 ;
  assign y8016 = n2220 ;
  assign y8017 = 1'b0 ;
  assign y8018 = ~n10763 ;
  assign y8019 = ~1'b0 ;
  assign y8020 = ~1'b0 ;
  assign y8021 = ~1'b0 ;
  assign y8022 = ~n10765 ;
  assign y8023 = n10766 ;
  assign y8024 = ~n10767 ;
  assign y8025 = ~1'b0 ;
  assign y8026 = n10769 ;
  assign y8027 = ~1'b0 ;
  assign y8028 = ~n273 ;
  assign y8029 = ~1'b0 ;
  assign y8030 = ~n10770 ;
  assign y8031 = ~n10772 ;
  assign y8032 = ~n3632 ;
  assign y8033 = ~n10774 ;
  assign y8034 = ~n10776 ;
  assign y8035 = n10778 ;
  assign y8036 = n10780 ;
  assign y8037 = ~n10781 ;
  assign y8038 = ~1'b0 ;
  assign y8039 = n10782 ;
  assign y8040 = n10785 ;
  assign y8041 = ~1'b0 ;
  assign y8042 = ~1'b0 ;
  assign y8043 = ~1'b0 ;
  assign y8044 = ~n10788 ;
  assign y8045 = ~1'b0 ;
  assign y8046 = n10795 ;
  assign y8047 = ~n10796 ;
  assign y8048 = n10798 ;
  assign y8049 = 1'b0 ;
  assign y8050 = 1'b0 ;
  assign y8051 = ~n10799 ;
  assign y8052 = 1'b0 ;
  assign y8053 = ~1'b0 ;
  assign y8054 = ~1'b0 ;
  assign y8055 = ~n10803 ;
  assign y8056 = n10807 ;
  assign y8057 = ~1'b0 ;
  assign y8058 = ~1'b0 ;
  assign y8059 = n10808 ;
  assign y8060 = ~n10809 ;
  assign y8061 = n10814 ;
  assign y8062 = ~n10818 ;
  assign y8063 = n10822 ;
  assign y8064 = ~n954 ;
  assign y8065 = ~1'b0 ;
  assign y8066 = n10823 ;
  assign y8067 = ~1'b0 ;
  assign y8068 = ~1'b0 ;
  assign y8069 = ~1'b0 ;
  assign y8070 = n10824 ;
  assign y8071 = ~n10825 ;
  assign y8072 = ~n10826 ;
  assign y8073 = ~1'b0 ;
  assign y8074 = 1'b0 ;
  assign y8075 = ~1'b0 ;
  assign y8076 = ~1'b0 ;
  assign y8077 = ~1'b0 ;
  assign y8078 = ~1'b0 ;
  assign y8079 = ~1'b0 ;
  assign y8080 = n10827 ;
  assign y8081 = n10829 ;
  assign y8082 = ~1'b0 ;
  assign y8083 = n10830 ;
  assign y8084 = n724 ;
  assign y8085 = ~1'b0 ;
  assign y8086 = n10833 ;
  assign y8087 = ~n4522 ;
  assign y8088 = ~n10834 ;
  assign y8089 = ~n10836 ;
  assign y8090 = n10837 ;
  assign y8091 = 1'b0 ;
  assign y8092 = n10841 ;
  assign y8093 = ~1'b0 ;
  assign y8094 = ~1'b0 ;
  assign y8095 = ~n10845 ;
  assign y8096 = ~n10849 ;
  assign y8097 = ~n6610 ;
  assign y8098 = ~1'b0 ;
  assign y8099 = ~1'b0 ;
  assign y8100 = ~n10850 ;
  assign y8101 = 1'b0 ;
  assign y8102 = ~n1003 ;
  assign y8103 = n10852 ;
  assign y8104 = ~n10853 ;
  assign y8105 = ~1'b0 ;
  assign y8106 = ~1'b0 ;
  assign y8107 = ~n10856 ;
  assign y8108 = ~n10864 ;
  assign y8109 = n10865 ;
  assign y8110 = ~n10871 ;
  assign y8111 = n10874 ;
  assign y8112 = ~n10877 ;
  assign y8113 = ~1'b0 ;
  assign y8114 = ~1'b0 ;
  assign y8115 = n10880 ;
  assign y8116 = ~1'b0 ;
  assign y8117 = ~n10881 ;
  assign y8118 = ~1'b0 ;
  assign y8119 = 1'b0 ;
  assign y8120 = ~n7646 ;
  assign y8121 = n10882 ;
  assign y8122 = n10884 ;
  assign y8123 = n10885 ;
  assign y8124 = ~1'b0 ;
  assign y8125 = ~1'b0 ;
  assign y8126 = n10886 ;
  assign y8127 = n7090 ;
  assign y8128 = n6102 ;
  assign y8129 = ~1'b0 ;
  assign y8130 = n2371 ;
  assign y8131 = 1'b0 ;
  assign y8132 = n10899 ;
  assign y8133 = ~n10902 ;
  assign y8134 = 1'b0 ;
  assign y8135 = n10903 ;
  assign y8136 = ~n10906 ;
  assign y8137 = ~1'b0 ;
  assign y8138 = n10909 ;
  assign y8139 = ~n10913 ;
  assign y8140 = ~1'b0 ;
  assign y8141 = n10914 ;
  assign y8142 = ~n10916 ;
  assign y8143 = ~1'b0 ;
  assign y8144 = n10919 ;
  assign y8145 = 1'b0 ;
  assign y8146 = ~1'b0 ;
  assign y8147 = ~1'b0 ;
  assign y8148 = ~n10922 ;
  assign y8149 = ~1'b0 ;
  assign y8150 = ~n10923 ;
  assign y8151 = ~1'b0 ;
  assign y8152 = 1'b0 ;
  assign y8153 = ~n10924 ;
  assign y8154 = n10925 ;
  assign y8155 = ~n7483 ;
  assign y8156 = ~n10926 ;
  assign y8157 = ~1'b0 ;
  assign y8158 = ~1'b0 ;
  assign y8159 = ~1'b0 ;
  assign y8160 = ~n10930 ;
  assign y8161 = n3880 ;
  assign y8162 = n10933 ;
  assign y8163 = ~1'b0 ;
  assign y8164 = ~1'b0 ;
  assign y8165 = ~1'b0 ;
  assign y8166 = ~n10934 ;
  assign y8167 = ~1'b0 ;
  assign y8168 = ~1'b0 ;
  assign y8169 = n10938 ;
  assign y8170 = n10940 ;
  assign y8171 = ~n7239 ;
  assign y8172 = ~1'b0 ;
  assign y8173 = ~n10945 ;
  assign y8174 = n10947 ;
  assign y8175 = ~n10950 ;
  assign y8176 = n8707 ;
  assign y8177 = n10951 ;
  assign y8178 = ~n10958 ;
  assign y8179 = ~n10963 ;
  assign y8180 = ~1'b0 ;
  assign y8181 = ~n10964 ;
  assign y8182 = ~n10965 ;
  assign y8183 = n10968 ;
  assign y8184 = ~1'b0 ;
  assign y8185 = ~n10970 ;
  assign y8186 = ~1'b0 ;
  assign y8187 = ~n10975 ;
  assign y8188 = n10977 ;
  assign y8189 = ~n10983 ;
  assign y8190 = ~n10984 ;
  assign y8191 = ~n10985 ;
  assign y8192 = n10991 ;
  assign y8193 = ~n10992 ;
  assign y8194 = n10995 ;
  assign y8195 = n10996 ;
  assign y8196 = ~n10998 ;
  assign y8197 = ~1'b0 ;
  assign y8198 = ~n9966 ;
  assign y8199 = n11000 ;
  assign y8200 = ~n11002 ;
  assign y8201 = ~n11005 ;
  assign y8202 = ~1'b0 ;
  assign y8203 = ~n5566 ;
  assign y8204 = ~n11007 ;
  assign y8205 = ~n11010 ;
  assign y8206 = ~n11012 ;
  assign y8207 = ~1'b0 ;
  assign y8208 = ~1'b0 ;
  assign y8209 = ~1'b0 ;
  assign y8210 = n38 ;
  assign y8211 = ~n11016 ;
  assign y8212 = ~1'b0 ;
  assign y8213 = ~1'b0 ;
  assign y8214 = ~n11020 ;
  assign y8215 = ~1'b0 ;
  assign y8216 = ~1'b0 ;
  assign y8217 = ~n11023 ;
  assign y8218 = ~1'b0 ;
  assign y8219 = ~1'b0 ;
  assign y8220 = n11026 ;
  assign y8221 = n11027 ;
  assign y8222 = ~1'b0 ;
  assign y8223 = n3046 ;
  assign y8224 = n6011 ;
  assign y8225 = ~1'b0 ;
  assign y8226 = ~n11032 ;
  assign y8227 = n11035 ;
  assign y8228 = ~n11037 ;
  assign y8229 = n11040 ;
  assign y8230 = ~1'b0 ;
  assign y8231 = ~1'b0 ;
  assign y8232 = n11042 ;
  assign y8233 = ~1'b0 ;
  assign y8234 = ~n11050 ;
  assign y8235 = ~1'b0 ;
  assign y8236 = ~n11051 ;
  assign y8237 = n11055 ;
  assign y8238 = 1'b0 ;
  assign y8239 = ~1'b0 ;
  assign y8240 = n9667 ;
  assign y8241 = n11056 ;
  assign y8242 = n11065 ;
  assign y8243 = ~1'b0 ;
  assign y8244 = ~n11069 ;
  assign y8245 = ~n11071 ;
  assign y8246 = n6558 ;
  assign y8247 = ~1'b0 ;
  assign y8248 = ~1'b0 ;
  assign y8249 = ~n11076 ;
  assign y8250 = n11077 ;
  assign y8251 = ~1'b0 ;
  assign y8252 = ~n11081 ;
  assign y8253 = ~1'b0 ;
  assign y8254 = ~1'b0 ;
  assign y8255 = ~1'b0 ;
  assign y8256 = n11085 ;
  assign y8257 = n11088 ;
  assign y8258 = 1'b0 ;
  assign y8259 = n105 ;
  assign y8260 = ~n11089 ;
  assign y8261 = ~1'b0 ;
  assign y8262 = ~1'b0 ;
  assign y8263 = ~n11093 ;
  assign y8264 = n11106 ;
  assign y8265 = ~1'b0 ;
  assign y8266 = n11107 ;
  assign y8267 = ~n11108 ;
  assign y8268 = n11115 ;
  assign y8269 = n11116 ;
  assign y8270 = ~1'b0 ;
  assign y8271 = ~1'b0 ;
  assign y8272 = ~1'b0 ;
  assign y8273 = ~1'b0 ;
  assign y8274 = n11120 ;
  assign y8275 = ~1'b0 ;
  assign y8276 = ~n11122 ;
  assign y8277 = ~n11123 ;
  assign y8278 = n11124 ;
  assign y8279 = ~1'b0 ;
  assign y8280 = n11126 ;
  assign y8281 = ~1'b0 ;
  assign y8282 = ~1'b0 ;
  assign y8283 = ~n11127 ;
  assign y8284 = ~1'b0 ;
  assign y8285 = ~1'b0 ;
  assign y8286 = ~n11131 ;
  assign y8287 = ~n11132 ;
  assign y8288 = n11133 ;
  assign y8289 = ~1'b0 ;
  assign y8290 = n9512 ;
  assign y8291 = ~n11136 ;
  assign y8292 = ~1'b0 ;
  assign y8293 = ~1'b0 ;
  assign y8294 = ~n11152 ;
  assign y8295 = n11153 ;
  assign y8296 = n11157 ;
  assign y8297 = n4308 ;
  assign y8298 = ~n2462 ;
  assign y8299 = n11158 ;
  assign y8300 = n11160 ;
  assign y8301 = 1'b0 ;
  assign y8302 = n11175 ;
  assign y8303 = ~1'b0 ;
  assign y8304 = ~n30 ;
  assign y8305 = ~n11177 ;
  assign y8306 = ~n11182 ;
  assign y8307 = ~n11186 ;
  assign y8308 = ~1'b0 ;
  assign y8309 = 1'b0 ;
  assign y8310 = ~1'b0 ;
  assign y8311 = n11188 ;
  assign y8312 = ~1'b0 ;
  assign y8313 = ~1'b0 ;
  assign y8314 = ~1'b0 ;
  assign y8315 = ~1'b0 ;
  assign y8316 = ~1'b0 ;
  assign y8317 = ~1'b0 ;
  assign y8318 = ~n11189 ;
  assign y8319 = ~1'b0 ;
  assign y8320 = ~1'b0 ;
  assign y8321 = 1'b0 ;
  assign y8322 = 1'b0 ;
  assign y8323 = n11193 ;
  assign y8324 = n11203 ;
  assign y8325 = ~1'b0 ;
  assign y8326 = ~1'b0 ;
  assign y8327 = ~n11204 ;
  assign y8328 = n11207 ;
  assign y8329 = ~1'b0 ;
  assign y8330 = ~1'b0 ;
  assign y8331 = ~n671 ;
  assign y8332 = ~n2377 ;
  assign y8333 = ~n11209 ;
  assign y8334 = ~1'b0 ;
  assign y8335 = ~n3931 ;
  assign y8336 = ~n11210 ;
  assign y8337 = ~1'b0 ;
  assign y8338 = ~1'b0 ;
  assign y8339 = ~n11211 ;
  assign y8340 = ~n11216 ;
  assign y8341 = n11222 ;
  assign y8342 = ~1'b0 ;
  assign y8343 = ~n4538 ;
  assign y8344 = ~n11224 ;
  assign y8345 = ~1'b0 ;
  assign y8346 = ~1'b0 ;
  assign y8347 = n11232 ;
  assign y8348 = ~1'b0 ;
  assign y8349 = ~n11237 ;
  assign y8350 = n11037 ;
  assign y8351 = ~n11238 ;
  assign y8352 = ~1'b0 ;
  assign y8353 = ~n11239 ;
  assign y8354 = n333 ;
  assign y8355 = ~n11246 ;
  assign y8356 = ~n11250 ;
  assign y8357 = ~n11253 ;
  assign y8358 = ~n11255 ;
  assign y8359 = ~n541 ;
  assign y8360 = n11256 ;
  assign y8361 = ~1'b0 ;
  assign y8362 = n11261 ;
  assign y8363 = 1'b0 ;
  assign y8364 = n11264 ;
  assign y8365 = ~1'b0 ;
  assign y8366 = ~1'b0 ;
  assign y8367 = ~n11266 ;
  assign y8368 = ~1'b0 ;
  assign y8369 = ~1'b0 ;
  assign y8370 = n11267 ;
  assign y8371 = n11268 ;
  assign y8372 = ~n677 ;
  assign y8373 = ~n11270 ;
  assign y8374 = n11272 ;
  assign y8375 = n7920 ;
  assign y8376 = n11274 ;
  assign y8377 = ~n11275 ;
  assign y8378 = ~1'b0 ;
  assign y8379 = ~n11276 ;
  assign y8380 = ~n11279 ;
  assign y8381 = ~n11281 ;
  assign y8382 = ~1'b0 ;
  assign y8383 = 1'b0 ;
  assign y8384 = ~n11293 ;
  assign y8385 = n11294 ;
  assign y8386 = ~1'b0 ;
  assign y8387 = ~n11295 ;
  assign y8388 = ~1'b0 ;
  assign y8389 = n11296 ;
  assign y8390 = ~1'b0 ;
  assign y8391 = ~1'b0 ;
  assign y8392 = ~1'b0 ;
  assign y8393 = ~n11299 ;
  assign y8394 = ~n11301 ;
  assign y8395 = ~1'b0 ;
  assign y8396 = ~n11302 ;
  assign y8397 = ~1'b0 ;
  assign y8398 = ~n11304 ;
  assign y8399 = ~1'b0 ;
  assign y8400 = ~1'b0 ;
  assign y8401 = ~n11307 ;
  assign y8402 = n11315 ;
  assign y8403 = n11316 ;
  assign y8404 = ~1'b0 ;
  assign y8405 = ~1'b0 ;
  assign y8406 = ~1'b0 ;
  assign y8407 = ~1'b0 ;
  assign y8408 = n11317 ;
  assign y8409 = ~n11321 ;
  assign y8410 = n11323 ;
  assign y8411 = ~n11326 ;
  assign y8412 = ~n1208 ;
  assign y8413 = n11329 ;
  assign y8414 = ~n11330 ;
  assign y8415 = ~n11335 ;
  assign y8416 = ~1'b0 ;
  assign y8417 = ~n11340 ;
  assign y8418 = ~n11342 ;
  assign y8419 = ~n11343 ;
  assign y8420 = 1'b0 ;
  assign y8421 = 1'b0 ;
  assign y8422 = ~n11346 ;
  assign y8423 = n3526 ;
  assign y8424 = n11348 ;
  assign y8425 = n11349 ;
  assign y8426 = ~n11351 ;
  assign y8427 = ~n11353 ;
  assign y8428 = ~1'b0 ;
  assign y8429 = ~1'b0 ;
  assign y8430 = ~n1943 ;
  assign y8431 = ~1'b0 ;
  assign y8432 = ~1'b0 ;
  assign y8433 = 1'b0 ;
  assign y8434 = ~1'b0 ;
  assign y8435 = n443 ;
  assign y8436 = n11355 ;
  assign y8437 = ~n11357 ;
  assign y8438 = ~n6170 ;
  assign y8439 = ~1'b0 ;
  assign y8440 = n2847 ;
  assign y8441 = ~1'b0 ;
  assign y8442 = ~n11358 ;
  assign y8443 = ~n11360 ;
  assign y8444 = ~1'b0 ;
  assign y8445 = ~n7217 ;
  assign y8446 = ~1'b0 ;
  assign y8447 = 1'b0 ;
  assign y8448 = ~1'b0 ;
  assign y8449 = ~1'b0 ;
  assign y8450 = ~1'b0 ;
  assign y8451 = n11361 ;
  assign y8452 = ~1'b0 ;
  assign y8453 = n11363 ;
  assign y8454 = ~n685 ;
  assign y8455 = n11367 ;
  assign y8456 = ~n11368 ;
  assign y8457 = ~n11369 ;
  assign y8458 = ~n11371 ;
  assign y8459 = ~1'b0 ;
  assign y8460 = ~n8330 ;
  assign y8461 = ~n11374 ;
  assign y8462 = n11375 ;
  assign y8463 = ~1'b0 ;
  assign y8464 = n11379 ;
  assign y8465 = ~1'b0 ;
  assign y8466 = 1'b0 ;
  assign y8467 = ~n4070 ;
  assign y8468 = ~1'b0 ;
  assign y8469 = ~1'b0 ;
  assign y8470 = ~1'b0 ;
  assign y8471 = n11385 ;
  assign y8472 = ~n5161 ;
  assign y8473 = ~1'b0 ;
  assign y8474 = ~n11389 ;
  assign y8475 = n11390 ;
  assign y8476 = ~1'b0 ;
  assign y8477 = ~n11391 ;
  assign y8478 = ~n11393 ;
  assign y8479 = 1'b0 ;
  assign y8480 = ~1'b0 ;
  assign y8481 = n9758 ;
  assign y8482 = ~1'b0 ;
  assign y8483 = n11394 ;
  assign y8484 = ~n11397 ;
  assign y8485 = ~1'b0 ;
  assign y8486 = ~1'b0 ;
  assign y8487 = n7077 ;
  assign y8488 = n11400 ;
  assign y8489 = n8081 ;
  assign y8490 = ~1'b0 ;
  assign y8491 = ~1'b0 ;
  assign y8492 = ~n11401 ;
  assign y8493 = 1'b0 ;
  assign y8494 = ~1'b0 ;
  assign y8495 = n11402 ;
  assign y8496 = ~n11404 ;
  assign y8497 = ~n7609 ;
  assign y8498 = ~1'b0 ;
  assign y8499 = n8158 ;
  assign y8500 = ~n11405 ;
  assign y8501 = ~1'b0 ;
  assign y8502 = ~1'b0 ;
  assign y8503 = ~n11406 ;
  assign y8504 = ~1'b0 ;
  assign y8505 = n11409 ;
  assign y8506 = n11410 ;
  assign y8507 = ~1'b0 ;
  assign y8508 = ~n11412 ;
  assign y8509 = ~1'b0 ;
  assign y8510 = ~n11413 ;
  assign y8511 = n11415 ;
  assign y8512 = ~1'b0 ;
  assign y8513 = n11419 ;
  assign y8514 = ~n10525 ;
  assign y8515 = ~n695 ;
  assign y8516 = ~1'b0 ;
  assign y8517 = n11423 ;
  assign y8518 = ~n11425 ;
  assign y8519 = ~n817 ;
  assign y8520 = ~n9567 ;
  assign y8521 = ~1'b0 ;
  assign y8522 = ~n11426 ;
  assign y8523 = n11429 ;
  assign y8524 = ~n11431 ;
  assign y8525 = n11434 ;
  assign y8526 = ~n11435 ;
  assign y8527 = ~n7465 ;
  assign y8528 = ~n11436 ;
  assign y8529 = ~n8639 ;
  assign y8530 = ~n11437 ;
  assign y8531 = ~n11438 ;
  assign y8532 = ~1'b0 ;
  assign y8533 = ~n11439 ;
  assign y8534 = ~1'b0 ;
  assign y8535 = ~1'b0 ;
  assign y8536 = ~1'b0 ;
  assign y8537 = ~n11444 ;
  assign y8538 = ~n5701 ;
  assign y8539 = ~n11447 ;
  assign y8540 = 1'b0 ;
  assign y8541 = ~n11448 ;
  assign y8542 = n227 ;
  assign y8543 = ~1'b0 ;
  assign y8544 = ~1'b0 ;
  assign y8545 = ~1'b0 ;
  assign y8546 = n9149 ;
  assign y8547 = ~n11449 ;
  assign y8548 = n11452 ;
  assign y8549 = ~1'b0 ;
  assign y8550 = ~1'b0 ;
  assign y8551 = ~1'b0 ;
  assign y8552 = ~1'b0 ;
  assign y8553 = ~1'b0 ;
  assign y8554 = ~n11458 ;
  assign y8555 = ~1'b0 ;
  assign y8556 = n11462 ;
  assign y8557 = n11465 ;
  assign y8558 = ~1'b0 ;
  assign y8559 = ~1'b0 ;
  assign y8560 = ~1'b0 ;
  assign y8561 = ~n11471 ;
  assign y8562 = ~n11478 ;
  assign y8563 = ~1'b0 ;
  assign y8564 = ~n11479 ;
  assign y8565 = ~n11481 ;
  assign y8566 = ~n11485 ;
  assign y8567 = ~n11486 ;
  assign y8568 = ~n11491 ;
  assign y8569 = ~1'b0 ;
  assign y8570 = ~1'b0 ;
  assign y8571 = n11492 ;
  assign y8572 = 1'b0 ;
  assign y8573 = ~1'b0 ;
  assign y8574 = n11493 ;
  assign y8575 = 1'b0 ;
  assign y8576 = n11499 ;
  assign y8577 = 1'b0 ;
  assign y8578 = n1004 ;
  assign y8579 = ~n11501 ;
  assign y8580 = n11503 ;
  assign y8581 = ~n11506 ;
  assign y8582 = ~1'b0 ;
  assign y8583 = ~1'b0 ;
  assign y8584 = ~1'b0 ;
  assign y8585 = ~1'b0 ;
  assign y8586 = ~n11510 ;
  assign y8587 = n11513 ;
  assign y8588 = ~1'b0 ;
  assign y8589 = ~1'b0 ;
  assign y8590 = ~n11514 ;
  assign y8591 = ~n11515 ;
  assign y8592 = n1431 ;
  assign y8593 = n11516 ;
  assign y8594 = n11518 ;
  assign y8595 = ~1'b0 ;
  assign y8596 = n11524 ;
  assign y8597 = ~1'b0 ;
  assign y8598 = n11525 ;
  assign y8599 = ~n11528 ;
  assign y8600 = ~n11531 ;
  assign y8601 = n11542 ;
  assign y8602 = ~1'b0 ;
  assign y8603 = ~n11543 ;
  assign y8604 = ~1'b0 ;
  assign y8605 = ~n11545 ;
  assign y8606 = ~1'b0 ;
  assign y8607 = ~1'b0 ;
  assign y8608 = ~n11546 ;
  assign y8609 = ~n11548 ;
  assign y8610 = ~1'b0 ;
  assign y8611 = ~1'b0 ;
  assign y8612 = ~1'b0 ;
  assign y8613 = n11552 ;
  assign y8614 = ~1'b0 ;
  assign y8615 = ~1'b0 ;
  assign y8616 = ~n11555 ;
  assign y8617 = n11561 ;
  assign y8618 = ~n3452 ;
  assign y8619 = n11562 ;
  assign y8620 = ~n11568 ;
  assign y8621 = ~1'b0 ;
  assign y8622 = ~1'b0 ;
  assign y8623 = ~n11570 ;
  assign y8624 = 1'b0 ;
  assign y8625 = ~1'b0 ;
  assign y8626 = ~n11582 ;
  assign y8627 = n7439 ;
  assign y8628 = ~1'b0 ;
  assign y8629 = ~n11583 ;
  assign y8630 = ~1'b0 ;
  assign y8631 = ~1'b0 ;
  assign y8632 = ~1'b0 ;
  assign y8633 = ~1'b0 ;
  assign y8634 = ~n11584 ;
  assign y8635 = n11587 ;
  assign y8636 = ~n11588 ;
  assign y8637 = n11591 ;
  assign y8638 = n11592 ;
  assign y8639 = n11597 ;
  assign y8640 = n11598 ;
  assign y8641 = n11600 ;
  assign y8642 = 1'b0 ;
  assign y8643 = ~n9036 ;
  assign y8644 = ~1'b0 ;
  assign y8645 = n11602 ;
  assign y8646 = n11603 ;
  assign y8647 = ~n11604 ;
  assign y8648 = ~n11612 ;
  assign y8649 = ~1'b0 ;
  assign y8650 = ~1'b0 ;
  assign y8651 = ~1'b0 ;
  assign y8652 = ~1'b0 ;
  assign y8653 = ~1'b0 ;
  assign y8654 = 1'b0 ;
  assign y8655 = ~n11615 ;
  assign y8656 = ~n11618 ;
  assign y8657 = ~n9733 ;
  assign y8658 = ~1'b0 ;
  assign y8659 = ~1'b0 ;
  assign y8660 = ~1'b0 ;
  assign y8661 = ~n11619 ;
  assign y8662 = ~n9412 ;
  assign y8663 = ~n11623 ;
  assign y8664 = ~n11624 ;
  assign y8665 = ~n11626 ;
  assign y8666 = n11627 ;
  assign y8667 = n11629 ;
  assign y8668 = ~n11633 ;
  assign y8669 = ~1'b0 ;
  assign y8670 = ~1'b0 ;
  assign y8671 = n11634 ;
  assign y8672 = n11635 ;
  assign y8673 = ~n11637 ;
  assign y8674 = ~1'b0 ;
  assign y8675 = ~1'b0 ;
  assign y8676 = ~1'b0 ;
  assign y8677 = n11638 ;
  assign y8678 = ~n11644 ;
  assign y8679 = n11646 ;
  assign y8680 = n137 ;
  assign y8681 = ~1'b0 ;
  assign y8682 = ~n11653 ;
  assign y8683 = n11654 ;
  assign y8684 = ~1'b0 ;
  assign y8685 = ~1'b0 ;
  assign y8686 = ~n8396 ;
  assign y8687 = ~n11656 ;
  assign y8688 = n11658 ;
  assign y8689 = ~n11660 ;
  assign y8690 = ~1'b0 ;
  assign y8691 = ~1'b0 ;
  assign y8692 = ~n11662 ;
  assign y8693 = ~n10191 ;
  assign y8694 = n11664 ;
  assign y8695 = ~1'b0 ;
  assign y8696 = ~1'b0 ;
  assign y8697 = ~1'b0 ;
  assign y8698 = ~1'b0 ;
  assign y8699 = ~n11667 ;
  assign y8700 = n11669 ;
  assign y8701 = ~1'b0 ;
  assign y8702 = n4875 ;
  assign y8703 = n11670 ;
  assign y8704 = ~1'b0 ;
  assign y8705 = ~1'b0 ;
  assign y8706 = n11674 ;
  assign y8707 = ~1'b0 ;
  assign y8708 = n11676 ;
  assign y8709 = ~n3501 ;
  assign y8710 = n9228 ;
  assign y8711 = ~n11678 ;
  assign y8712 = n11679 ;
  assign y8713 = 1'b0 ;
  assign y8714 = n11680 ;
  assign y8715 = ~1'b0 ;
  assign y8716 = n11684 ;
  assign y8717 = n11686 ;
  assign y8718 = ~1'b0 ;
  assign y8719 = ~n11687 ;
  assign y8720 = ~1'b0 ;
  assign y8721 = ~1'b0 ;
  assign y8722 = ~1'b0 ;
  assign y8723 = ~1'b0 ;
  assign y8724 = ~1'b0 ;
  assign y8725 = ~n11690 ;
  assign y8726 = 1'b0 ;
  assign y8727 = n11692 ;
  assign y8728 = ~1'b0 ;
  assign y8729 = ~1'b0 ;
  assign y8730 = ~n11693 ;
  assign y8731 = ~1'b0 ;
  assign y8732 = n11694 ;
  assign y8733 = n11696 ;
  assign y8734 = ~n11700 ;
  assign y8735 = n6332 ;
  assign y8736 = 1'b0 ;
  assign y8737 = ~n11711 ;
  assign y8738 = n11712 ;
  assign y8739 = ~n5111 ;
  assign y8740 = ~n11714 ;
  assign y8741 = ~1'b0 ;
  assign y8742 = n11717 ;
  assign y8743 = ~1'b0 ;
  assign y8744 = ~1'b0 ;
  assign y8745 = ~n5409 ;
  assign y8746 = ~n11718 ;
  assign y8747 = ~n11720 ;
  assign y8748 = ~1'b0 ;
  assign y8749 = ~n11721 ;
  assign y8750 = n11723 ;
  assign y8751 = n11726 ;
  assign y8752 = ~1'b0 ;
  assign y8753 = n11729 ;
  assign y8754 = ~1'b0 ;
  assign y8755 = ~1'b0 ;
  assign y8756 = n11732 ;
  assign y8757 = n364 ;
  assign y8758 = ~n11733 ;
  assign y8759 = n11734 ;
  assign y8760 = ~1'b0 ;
  assign y8761 = ~1'b0 ;
  assign y8762 = ~n11737 ;
  assign y8763 = ~n1465 ;
  assign y8764 = n11738 ;
  assign y8765 = ~1'b0 ;
  assign y8766 = ~1'b0 ;
  assign y8767 = n11740 ;
  assign y8768 = n11750 ;
  assign y8769 = n11751 ;
  assign y8770 = ~n11753 ;
  assign y8771 = ~n7381 ;
  assign y8772 = ~n11755 ;
  assign y8773 = ~1'b0 ;
  assign y8774 = n11756 ;
  assign y8775 = ~1'b0 ;
  assign y8776 = ~n11758 ;
  assign y8777 = n11760 ;
  assign y8778 = n11763 ;
  assign y8779 = n11765 ;
  assign y8780 = ~n11770 ;
  assign y8781 = n11771 ;
  assign y8782 = ~n11772 ;
  assign y8783 = n11773 ;
  assign y8784 = ~1'b0 ;
  assign y8785 = 1'b0 ;
  assign y8786 = ~1'b0 ;
  assign y8787 = n11775 ;
  assign y8788 = ~1'b0 ;
  assign y8789 = 1'b0 ;
  assign y8790 = ~1'b0 ;
  assign y8791 = n11776 ;
  assign y8792 = n11778 ;
  assign y8793 = ~1'b0 ;
  assign y8794 = n958 ;
  assign y8795 = n11782 ;
  assign y8796 = ~1'b0 ;
  assign y8797 = ~1'b0 ;
  assign y8798 = n11783 ;
  assign y8799 = ~1'b0 ;
  assign y8800 = 1'b0 ;
  assign y8801 = n11784 ;
  assign y8802 = ~1'b0 ;
  assign y8803 = n11787 ;
  assign y8804 = ~n11794 ;
  assign y8805 = n11796 ;
  assign y8806 = ~n11797 ;
  assign y8807 = n11798 ;
  assign y8808 = ~n4311 ;
  assign y8809 = n1829 ;
  assign y8810 = n11192 ;
  assign y8811 = ~n11800 ;
  assign y8812 = ~1'b0 ;
  assign y8813 = ~1'b0 ;
  assign y8814 = n11804 ;
  assign y8815 = ~n11806 ;
  assign y8816 = n3951 ;
  assign y8817 = n11807 ;
  assign y8818 = ~n2910 ;
  assign y8819 = n11809 ;
  assign y8820 = ~1'b0 ;
  assign y8821 = ~n11818 ;
  assign y8822 = n11821 ;
  assign y8823 = ~1'b0 ;
  assign y8824 = ~n11824 ;
  assign y8825 = ~n11826 ;
  assign y8826 = ~n11827 ;
  assign y8827 = n11829 ;
  assign y8828 = ~1'b0 ;
  assign y8829 = 1'b0 ;
  assign y8830 = ~n6094 ;
  assign y8831 = ~1'b0 ;
  assign y8832 = ~1'b0 ;
  assign y8833 = n11834 ;
  assign y8834 = 1'b0 ;
  assign y8835 = ~n11837 ;
  assign y8836 = ~n11838 ;
  assign y8837 = ~n11844 ;
  assign y8838 = ~n9799 ;
  assign y8839 = ~n11847 ;
  assign y8840 = ~1'b0 ;
  assign y8841 = ~n11848 ;
  assign y8842 = ~n11850 ;
  assign y8843 = n11851 ;
  assign y8844 = ~1'b0 ;
  assign y8845 = ~n11852 ;
  assign y8846 = n11854 ;
  assign y8847 = ~1'b0 ;
  assign y8848 = ~1'b0 ;
  assign y8849 = ~1'b0 ;
  assign y8850 = n11861 ;
  assign y8851 = n11862 ;
  assign y8852 = ~n11864 ;
  assign y8853 = ~n3697 ;
  assign y8854 = ~1'b0 ;
  assign y8855 = ~n11866 ;
  assign y8856 = n11869 ;
  assign y8857 = ~1'b0 ;
  assign y8858 = ~n11874 ;
  assign y8859 = ~n11875 ;
  assign y8860 = 1'b0 ;
  assign y8861 = ~n11885 ;
  assign y8862 = ~1'b0 ;
  assign y8863 = n11886 ;
  assign y8864 = ~1'b0 ;
  assign y8865 = ~1'b0 ;
  assign y8866 = ~n11891 ;
  assign y8867 = n11894 ;
  assign y8868 = ~1'b0 ;
  assign y8869 = ~n11900 ;
  assign y8870 = n11907 ;
  assign y8871 = ~1'b0 ;
  assign y8872 = n11909 ;
  assign y8873 = ~1'b0 ;
  assign y8874 = 1'b0 ;
  assign y8875 = ~n11912 ;
  assign y8876 = ~n11916 ;
  assign y8877 = n11917 ;
  assign y8878 = ~n11926 ;
  assign y8879 = ~n107 ;
  assign y8880 = ~1'b0 ;
  assign y8881 = ~n11927 ;
  assign y8882 = ~n11929 ;
  assign y8883 = ~n11937 ;
  assign y8884 = n11938 ;
  assign y8885 = ~1'b0 ;
  assign y8886 = ~n481 ;
  assign y8887 = ~1'b0 ;
  assign y8888 = n11943 ;
  assign y8889 = ~n11956 ;
  assign y8890 = n2607 ;
  assign y8891 = n11959 ;
  assign y8892 = n11961 ;
  assign y8893 = n11965 ;
  assign y8894 = ~1'b0 ;
  assign y8895 = ~1'b0 ;
  assign y8896 = ~n11967 ;
  assign y8897 = ~n11969 ;
  assign y8898 = ~1'b0 ;
  assign y8899 = ~n3843 ;
  assign y8900 = n11970 ;
  assign y8901 = n11971 ;
  assign y8902 = n11972 ;
  assign y8903 = n11973 ;
  assign y8904 = ~1'b0 ;
  assign y8905 = ~1'b0 ;
  assign y8906 = n11977 ;
  assign y8907 = n11980 ;
  assign y8908 = ~1'b0 ;
  assign y8909 = ~1'b0 ;
  assign y8910 = n11981 ;
  assign y8911 = n3099 ;
  assign y8912 = ~n9535 ;
  assign y8913 = ~1'b0 ;
  assign y8914 = ~n11982 ;
  assign y8915 = n11988 ;
  assign y8916 = n4799 ;
  assign y8917 = n11990 ;
  assign y8918 = ~n11992 ;
  assign y8919 = ~n11994 ;
  assign y8920 = ~1'b0 ;
  assign y8921 = n11998 ;
  assign y8922 = ~n12002 ;
  assign y8923 = n12005 ;
  assign y8924 = ~n12006 ;
  assign y8925 = ~1'b0 ;
  assign y8926 = 1'b0 ;
  assign y8927 = ~1'b0 ;
  assign y8928 = ~1'b0 ;
  assign y8929 = ~n12013 ;
  assign y8930 = n12014 ;
  assign y8931 = ~n12019 ;
  assign y8932 = ~1'b0 ;
  assign y8933 = n12021 ;
  assign y8934 = 1'b0 ;
  assign y8935 = n12022 ;
  assign y8936 = ~n12026 ;
  assign y8937 = ~n12028 ;
  assign y8938 = ~1'b0 ;
  assign y8939 = n12029 ;
  assign y8940 = ~1'b0 ;
  assign y8941 = ~n12033 ;
  assign y8942 = ~n12037 ;
  assign y8943 = ~n12045 ;
  assign y8944 = ~n10057 ;
  assign y8945 = ~n12049 ;
  assign y8946 = n4358 ;
  assign y8947 = n12050 ;
  assign y8948 = ~n12051 ;
  assign y8949 = 1'b0 ;
  assign y8950 = ~n12054 ;
  assign y8951 = ~n5551 ;
  assign y8952 = ~n12056 ;
  assign y8953 = 1'b0 ;
  assign y8954 = n12059 ;
  assign y8955 = n12062 ;
  assign y8956 = ~1'b0 ;
  assign y8957 = n12064 ;
  assign y8958 = ~1'b0 ;
  assign y8959 = ~n12066 ;
  assign y8960 = n12067 ;
  assign y8961 = ~n12072 ;
  assign y8962 = ~n12073 ;
  assign y8963 = ~n12076 ;
  assign y8964 = ~1'b0 ;
  assign y8965 = ~n12080 ;
  assign y8966 = ~n12082 ;
  assign y8967 = ~n12087 ;
  assign y8968 = ~n12092 ;
  assign y8969 = ~1'b0 ;
  assign y8970 = ~1'b0 ;
  assign y8971 = n12099 ;
  assign y8972 = n439 ;
  assign y8973 = n12104 ;
  assign y8974 = ~n12108 ;
  assign y8975 = n12109 ;
  assign y8976 = ~1'b0 ;
  assign y8977 = ~n12111 ;
  assign y8978 = ~n12121 ;
  assign y8979 = ~1'b0 ;
  assign y8980 = n6270 ;
  assign y8981 = ~n12123 ;
  assign y8982 = n12155 ;
  assign y8983 = ~n12159 ;
  assign y8984 = ~n9507 ;
  assign y8985 = n5877 ;
  assign y8986 = ~n12162 ;
  assign y8987 = n12163 ;
  assign y8988 = n12165 ;
  assign y8989 = n12170 ;
  assign y8990 = ~n12171 ;
  assign y8991 = n12172 ;
  assign y8992 = n12173 ;
  assign y8993 = ~1'b0 ;
  assign y8994 = ~1'b0 ;
  assign y8995 = ~1'b0 ;
  assign y8996 = n12178 ;
  assign y8997 = n12180 ;
  assign y8998 = ~n12184 ;
  assign y8999 = ~n2222 ;
  assign y9000 = ~1'b0 ;
  assign y9001 = ~1'b0 ;
  assign y9002 = ~1'b0 ;
  assign y9003 = ~n12185 ;
  assign y9004 = ~n12186 ;
  assign y9005 = ~1'b0 ;
  assign y9006 = n12187 ;
  assign y9007 = ~1'b0 ;
  assign y9008 = ~n6071 ;
  assign y9009 = n12188 ;
  assign y9010 = n12189 ;
  assign y9011 = ~n12192 ;
  assign y9012 = n12195 ;
  assign y9013 = ~1'b0 ;
  assign y9014 = ~1'b0 ;
  assign y9015 = ~1'b0 ;
  assign y9016 = ~n12198 ;
  assign y9017 = ~n12203 ;
  assign y9018 = 1'b0 ;
  assign y9019 = n907 ;
  assign y9020 = ~1'b0 ;
  assign y9021 = n12209 ;
  assign y9022 = ~n12210 ;
  assign y9023 = 1'b0 ;
  assign y9024 = ~1'b0 ;
  assign y9025 = n12212 ;
  assign y9026 = ~n12214 ;
  assign y9027 = n2819 ;
  assign y9028 = ~n12218 ;
  assign y9029 = ~n12224 ;
  assign y9030 = n6249 ;
  assign y9031 = ~1'b0 ;
  assign y9032 = ~n9491 ;
  assign y9033 = n12225 ;
  assign y9034 = ~n12227 ;
  assign y9035 = n12232 ;
  assign y9036 = 1'b0 ;
  assign y9037 = ~n12237 ;
  assign y9038 = n12238 ;
  assign y9039 = n12239 ;
  assign y9040 = ~n12240 ;
  assign y9041 = ~n12241 ;
  assign y9042 = ~n12242 ;
  assign y9043 = ~n12245 ;
  assign y9044 = ~1'b0 ;
  assign y9045 = ~1'b0 ;
  assign y9046 = ~n12248 ;
  assign y9047 = ~n12251 ;
  assign y9048 = ~1'b0 ;
  assign y9049 = 1'b0 ;
  assign y9050 = ~n12253 ;
  assign y9051 = ~1'b0 ;
  assign y9052 = ~n12254 ;
  assign y9053 = n4748 ;
  assign y9054 = ~1'b0 ;
  assign y9055 = ~n594 ;
  assign y9056 = 1'b0 ;
  assign y9057 = ~n12257 ;
  assign y9058 = ~n12259 ;
  assign y9059 = ~n12261 ;
  assign y9060 = ~1'b0 ;
  assign y9061 = ~n12263 ;
  assign y9062 = ~n12264 ;
  assign y9063 = ~1'b0 ;
  assign y9064 = ~1'b0 ;
  assign y9065 = n12265 ;
  assign y9066 = ~n12266 ;
  assign y9067 = n12268 ;
  assign y9068 = n12269 ;
  assign y9069 = n3116 ;
  assign y9070 = n12273 ;
  assign y9071 = n12274 ;
  assign y9072 = ~n12276 ;
  assign y9073 = ~n12278 ;
  assign y9074 = n3897 ;
  assign y9075 = n12280 ;
  assign y9076 = ~n12283 ;
  assign y9077 = ~n12284 ;
  assign y9078 = ~1'b0 ;
  assign y9079 = 1'b0 ;
  assign y9080 = ~1'b0 ;
  assign y9081 = ~n12286 ;
  assign y9082 = n12288 ;
  assign y9083 = n12289 ;
  assign y9084 = ~1'b0 ;
  assign y9085 = ~1'b0 ;
  assign y9086 = n12295 ;
  assign y9087 = n12298 ;
  assign y9088 = ~1'b0 ;
  assign y9089 = ~n12302 ;
  assign y9090 = ~n12303 ;
  assign y9091 = ~n12306 ;
  assign y9092 = ~1'b0 ;
  assign y9093 = n12308 ;
  assign y9094 = ~1'b0 ;
  assign y9095 = ~n12310 ;
  assign y9096 = 1'b0 ;
  assign y9097 = ~n12312 ;
  assign y9098 = n12313 ;
  assign y9099 = n12317 ;
  assign y9100 = ~n12318 ;
  assign y9101 = ~n12327 ;
  assign y9102 = n12328 ;
  assign y9103 = ~1'b0 ;
  assign y9104 = ~1'b0 ;
  assign y9105 = ~1'b0 ;
  assign y9106 = n12333 ;
  assign y9107 = ~1'b0 ;
  assign y9108 = ~1'b0 ;
  assign y9109 = n12345 ;
  assign y9110 = ~1'b0 ;
  assign y9111 = ~1'b0 ;
  assign y9112 = n12347 ;
  assign y9113 = ~n12349 ;
  assign y9114 = n12350 ;
  assign y9115 = ~1'b0 ;
  assign y9116 = ~1'b0 ;
  assign y9117 = ~n12353 ;
  assign y9118 = ~1'b0 ;
  assign y9119 = ~1'b0 ;
  assign y9120 = ~1'b0 ;
  assign y9121 = n12357 ;
  assign y9122 = n12360 ;
  assign y9123 = n12361 ;
  assign y9124 = ~n12362 ;
  assign y9125 = n12363 ;
  assign y9126 = ~n2519 ;
  assign y9127 = ~n10180 ;
  assign y9128 = ~n12364 ;
  assign y9129 = ~n12368 ;
  assign y9130 = ~1'b0 ;
  assign y9131 = ~1'b0 ;
  assign y9132 = n12370 ;
  assign y9133 = ~n12374 ;
  assign y9134 = ~n12376 ;
  assign y9135 = ~n12378 ;
  assign y9136 = n12379 ;
  assign y9137 = ~1'b0 ;
  assign y9138 = ~1'b0 ;
  assign y9139 = ~1'b0 ;
  assign y9140 = n12381 ;
  assign y9141 = ~n12382 ;
  assign y9142 = ~1'b0 ;
  assign y9143 = n12383 ;
  assign y9144 = ~1'b0 ;
  assign y9145 = ~n12385 ;
  assign y9146 = ~n12386 ;
  assign y9147 = n12387 ;
  assign y9148 = ~1'b0 ;
  assign y9149 = 1'b0 ;
  assign y9150 = n12388 ;
  assign y9151 = n12390 ;
  assign y9152 = ~n3423 ;
  assign y9153 = ~n12391 ;
  assign y9154 = ~1'b0 ;
  assign y9155 = ~1'b0 ;
  assign y9156 = ~1'b0 ;
  assign y9157 = n12393 ;
  assign y9158 = n2063 ;
  assign y9159 = ~n12395 ;
  assign y9160 = ~n12396 ;
  assign y9161 = ~n12398 ;
  assign y9162 = 1'b0 ;
  assign y9163 = ~1'b0 ;
  assign y9164 = ~1'b0 ;
  assign y9165 = ~n12399 ;
  assign y9166 = ~n12400 ;
  assign y9167 = n12401 ;
  assign y9168 = ~n2362 ;
  assign y9169 = n12404 ;
  assign y9170 = ~1'b0 ;
  assign y9171 = n12406 ;
  assign y9172 = ~n12411 ;
  assign y9173 = ~n12412 ;
  assign y9174 = ~1'b0 ;
  assign y9175 = ~1'b0 ;
  assign y9176 = ~1'b0 ;
  assign y9177 = ~1'b0 ;
  assign y9178 = ~n12414 ;
  assign y9179 = n12416 ;
  assign y9180 = n12417 ;
  assign y9181 = ~n12419 ;
  assign y9182 = n12420 ;
  assign y9183 = n12421 ;
  assign y9184 = ~1'b0 ;
  assign y9185 = ~n12424 ;
  assign y9186 = ~n12425 ;
  assign y9187 = n12427 ;
  assign y9188 = ~1'b0 ;
  assign y9189 = n12428 ;
  assign y9190 = ~n12429 ;
  assign y9191 = ~1'b0 ;
  assign y9192 = ~1'b0 ;
  assign y9193 = ~1'b0 ;
  assign y9194 = n12433 ;
  assign y9195 = ~n1331 ;
  assign y9196 = ~1'b0 ;
  assign y9197 = n12436 ;
  assign y9198 = ~n12438 ;
  assign y9199 = n12441 ;
  assign y9200 = ~1'b0 ;
  assign y9201 = ~1'b0 ;
  assign y9202 = n12442 ;
  assign y9203 = n12444 ;
  assign y9204 = n12452 ;
  assign y9205 = ~n12458 ;
  assign y9206 = n12462 ;
  assign y9207 = ~n12467 ;
  assign y9208 = ~1'b0 ;
  assign y9209 = ~n12470 ;
  assign y9210 = n12475 ;
  assign y9211 = ~1'b0 ;
  assign y9212 = ~n4842 ;
  assign y9213 = ~n12477 ;
  assign y9214 = n12481 ;
  assign y9215 = 1'b0 ;
  assign y9216 = n12484 ;
  assign y9217 = ~1'b0 ;
  assign y9218 = ~1'b0 ;
  assign y9219 = ~n12487 ;
  assign y9220 = n12488 ;
  assign y9221 = ~n4914 ;
  assign y9222 = n12489 ;
  assign y9223 = ~n12495 ;
  assign y9224 = n10470 ;
  assign y9225 = ~1'b0 ;
  assign y9226 = n12497 ;
  assign y9227 = ~1'b0 ;
  assign y9228 = ~1'b0 ;
  assign y9229 = n12500 ;
  assign y9230 = ~1'b0 ;
  assign y9231 = 1'b0 ;
  assign y9232 = n12502 ;
  assign y9233 = n12503 ;
  assign y9234 = n12505 ;
  assign y9235 = ~1'b0 ;
  assign y9236 = ~1'b0 ;
  assign y9237 = ~n12507 ;
  assign y9238 = n5575 ;
  assign y9239 = 1'b0 ;
  assign y9240 = n7920 ;
  assign y9241 = ~n12512 ;
  assign y9242 = n12513 ;
  assign y9243 = ~n12517 ;
  assign y9244 = ~1'b0 ;
  assign y9245 = ~n52 ;
  assign y9246 = ~n12518 ;
  assign y9247 = ~n12521 ;
  assign y9248 = n12526 ;
  assign y9249 = ~1'b0 ;
  assign y9250 = ~n12527 ;
  assign y9251 = n12530 ;
  assign y9252 = ~n12532 ;
  assign y9253 = ~n12533 ;
  assign y9254 = ~1'b0 ;
  assign y9255 = ~1'b0 ;
  assign y9256 = n12534 ;
  assign y9257 = ~n12537 ;
  assign y9258 = 1'b0 ;
  assign y9259 = ~1'b0 ;
  assign y9260 = ~n12539 ;
  assign y9261 = ~n12541 ;
  assign y9262 = 1'b0 ;
  assign y9263 = ~n12547 ;
  assign y9264 = n8900 ;
  assign y9265 = ~n12553 ;
  assign y9266 = ~1'b0 ;
  assign y9267 = ~1'b0 ;
  assign y9268 = ~n4424 ;
  assign y9269 = n7737 ;
  assign y9270 = ~n12555 ;
  assign y9271 = ~1'b0 ;
  assign y9272 = n12562 ;
  assign y9273 = n12563 ;
  assign y9274 = n12566 ;
  assign y9275 = ~1'b0 ;
  assign y9276 = ~n12626 ;
  assign y9277 = ~1'b0 ;
  assign y9278 = ~n9540 ;
  assign y9279 = n12629 ;
  assign y9280 = ~n5643 ;
  assign y9281 = ~1'b0 ;
  assign y9282 = n12630 ;
  assign y9283 = n12632 ;
  assign y9284 = ~1'b0 ;
  assign y9285 = ~1'b0 ;
  assign y9286 = ~n12637 ;
  assign y9287 = n12639 ;
  assign y9288 = n12641 ;
  assign y9289 = n12642 ;
  assign y9290 = ~1'b0 ;
  assign y9291 = ~1'b0 ;
  assign y9292 = ~n12645 ;
  assign y9293 = ~1'b0 ;
  assign y9294 = ~n3452 ;
  assign y9295 = ~1'b0 ;
  assign y9296 = ~1'b0 ;
  assign y9297 = ~n12651 ;
  assign y9298 = ~n12652 ;
  assign y9299 = n12655 ;
  assign y9300 = ~1'b0 ;
  assign y9301 = ~n4545 ;
  assign y9302 = ~n12656 ;
  assign y9303 = n12657 ;
  assign y9304 = ~n12660 ;
  assign y9305 = ~n12664 ;
  assign y9306 = ~1'b0 ;
  assign y9307 = ~n12665 ;
  assign y9308 = ~n12666 ;
  assign y9309 = n12303 ;
  assign y9310 = ~n12667 ;
  assign y9311 = n12671 ;
  assign y9312 = ~1'b0 ;
  assign y9313 = ~1'b0 ;
  assign y9314 = n12672 ;
  assign y9315 = ~n12678 ;
  assign y9316 = 1'b0 ;
  assign y9317 = ~1'b0 ;
  assign y9318 = ~n3162 ;
  assign y9319 = ~n12680 ;
  assign y9320 = n6889 ;
  assign y9321 = n12681 ;
  assign y9322 = ~n940 ;
  assign y9323 = ~n12683 ;
  assign y9324 = ~1'b0 ;
  assign y9325 = ~1'b0 ;
  assign y9326 = n12687 ;
  assign y9327 = n2856 ;
  assign y9328 = ~n12689 ;
  assign y9329 = ~n12690 ;
  assign y9330 = ~1'b0 ;
  assign y9331 = ~1'b0 ;
  assign y9332 = ~1'b0 ;
  assign y9333 = ~1'b0 ;
  assign y9334 = n12692 ;
  assign y9335 = ~n4131 ;
  assign y9336 = ~1'b0 ;
  assign y9337 = ~1'b0 ;
  assign y9338 = n3946 ;
  assign y9339 = ~1'b0 ;
  assign y9340 = ~n12696 ;
  assign y9341 = ~n12698 ;
  assign y9342 = ~n12699 ;
  assign y9343 = ~n12703 ;
  assign y9344 = ~n12705 ;
  assign y9345 = ~n12710 ;
  assign y9346 = ~n12711 ;
  assign y9347 = ~1'b0 ;
  assign y9348 = n11087 ;
  assign y9349 = ~n12713 ;
  assign y9350 = ~n12714 ;
  assign y9351 = n2903 ;
  assign y9352 = ~1'b0 ;
  assign y9353 = ~1'b0 ;
  assign y9354 = ~n12717 ;
  assign y9355 = n5498 ;
  assign y9356 = ~1'b0 ;
  assign y9357 = ~n12719 ;
  assign y9358 = n12720 ;
  assign y9359 = n12738 ;
  assign y9360 = ~1'b0 ;
  assign y9361 = n12746 ;
  assign y9362 = ~n12749 ;
  assign y9363 = ~1'b0 ;
  assign y9364 = ~n12752 ;
  assign y9365 = ~1'b0 ;
  assign y9366 = n12754 ;
  assign y9367 = n12756 ;
  assign y9368 = n12757 ;
  assign y9369 = ~1'b0 ;
  assign y9370 = 1'b0 ;
  assign y9371 = ~n3434 ;
  assign y9372 = ~1'b0 ;
  assign y9373 = n12758 ;
  assign y9374 = ~n5554 ;
  assign y9375 = ~1'b0 ;
  assign y9376 = n12760 ;
  assign y9377 = ~n12763 ;
  assign y9378 = 1'b0 ;
  assign y9379 = n12770 ;
  assign y9380 = ~n12721 ;
  assign y9381 = 1'b0 ;
  assign y9382 = ~n3855 ;
  assign y9383 = ~1'b0 ;
  assign y9384 = 1'b0 ;
  assign y9385 = n12772 ;
  assign y9386 = n12773 ;
  assign y9387 = n12776 ;
  assign y9388 = n12779 ;
  assign y9389 = n12784 ;
  assign y9390 = ~1'b0 ;
  assign y9391 = ~1'b0 ;
  assign y9392 = ~1'b0 ;
  assign y9393 = 1'b0 ;
  assign y9394 = n12785 ;
  assign y9395 = n12787 ;
  assign y9396 = ~n12791 ;
  assign y9397 = ~1'b0 ;
  assign y9398 = ~n12795 ;
  assign y9399 = ~1'b0 ;
  assign y9400 = ~1'b0 ;
  assign y9401 = ~n3019 ;
  assign y9402 = n12797 ;
  assign y9403 = n12800 ;
  assign y9404 = ~n12803 ;
  assign y9405 = n12807 ;
  assign y9406 = ~1'b0 ;
  assign y9407 = n12808 ;
  assign y9408 = ~1'b0 ;
  assign y9409 = 1'b0 ;
  assign y9410 = ~n12810 ;
  assign y9411 = n12811 ;
  assign y9412 = ~n12852 ;
  assign y9413 = n6015 ;
  assign y9414 = ~1'b0 ;
  assign y9415 = ~1'b0 ;
  assign y9416 = ~n12853 ;
  assign y9417 = ~1'b0 ;
  assign y9418 = ~1'b0 ;
  assign y9419 = ~1'b0 ;
  assign y9420 = 1'b0 ;
  assign y9421 = n11690 ;
  assign y9422 = n940 ;
  assign y9423 = ~1'b0 ;
  assign y9424 = n12854 ;
  assign y9425 = ~n12856 ;
  assign y9426 = ~n484 ;
  assign y9427 = n581 ;
  assign y9428 = ~1'b0 ;
  assign y9429 = ~n12863 ;
  assign y9430 = ~1'b0 ;
  assign y9431 = ~n12865 ;
  assign y9432 = ~1'b0 ;
  assign y9433 = n12868 ;
  assign y9434 = n6418 ;
  assign y9435 = n12873 ;
  assign y9436 = n12879 ;
  assign y9437 = ~1'b0 ;
  assign y9438 = n12880 ;
  assign y9439 = ~1'b0 ;
  assign y9440 = n12881 ;
  assign y9441 = ~1'b0 ;
  assign y9442 = 1'b0 ;
  assign y9443 = ~n12886 ;
  assign y9444 = n12887 ;
  assign y9445 = ~n12892 ;
  assign y9446 = ~n12893 ;
  assign y9447 = 1'b0 ;
  assign y9448 = 1'b0 ;
  assign y9449 = ~n12896 ;
  assign y9450 = ~n12901 ;
  assign y9451 = n12904 ;
  assign y9452 = ~n12906 ;
  assign y9453 = ~n2017 ;
  assign y9454 = ~1'b0 ;
  assign y9455 = ~1'b0 ;
  assign y9456 = 1'b0 ;
  assign y9457 = ~n12907 ;
  assign y9458 = ~n7419 ;
  assign y9459 = ~n832 ;
  assign y9460 = ~n12908 ;
  assign y9461 = ~1'b0 ;
  assign y9462 = ~n12909 ;
  assign y9463 = ~1'b0 ;
  assign y9464 = 1'b0 ;
  assign y9465 = ~1'b0 ;
  assign y9466 = ~n12910 ;
  assign y9467 = ~n12912 ;
  assign y9468 = n3007 ;
  assign y9469 = ~n12916 ;
  assign y9470 = ~n12917 ;
  assign y9471 = ~1'b0 ;
  assign y9472 = ~1'b0 ;
  assign y9473 = ~n12918 ;
  assign y9474 = ~1'b0 ;
  assign y9475 = n12925 ;
  assign y9476 = ~1'b0 ;
  assign y9477 = ~1'b0 ;
  assign y9478 = 1'b0 ;
  assign y9479 = n12926 ;
  assign y9480 = ~1'b0 ;
  assign y9481 = ~n12928 ;
  assign y9482 = n12934 ;
  assign y9483 = ~1'b0 ;
  assign y9484 = ~1'b0 ;
  assign y9485 = n12935 ;
  assign y9486 = n12939 ;
  assign y9487 = n12940 ;
  assign y9488 = ~n12942 ;
  assign y9489 = ~1'b0 ;
  assign y9490 = ~n12946 ;
  assign y9491 = ~n12950 ;
  assign y9492 = n12955 ;
  assign y9493 = ~1'b0 ;
  assign y9494 = ~n12961 ;
  assign y9495 = ~n12963 ;
  assign y9496 = ~n12964 ;
  assign y9497 = ~n12966 ;
  assign y9498 = ~1'b0 ;
  assign y9499 = 1'b0 ;
  assign y9500 = n12967 ;
  assign y9501 = n12969 ;
  assign y9502 = ~n12972 ;
  assign y9503 = n12974 ;
  assign y9504 = ~n12976 ;
  assign y9505 = ~1'b0 ;
  assign y9506 = ~1'b0 ;
  assign y9507 = ~n6942 ;
  assign y9508 = ~n12977 ;
  assign y9509 = ~1'b0 ;
  assign y9510 = ~n9483 ;
  assign y9511 = n12978 ;
  assign y9512 = n12980 ;
  assign y9513 = n12981 ;
  assign y9514 = ~1'b0 ;
  assign y9515 = n12984 ;
  assign y9516 = ~n12985 ;
  assign y9517 = ~1'b0 ;
  assign y9518 = ~n12986 ;
  assign y9519 = ~n3781 ;
  assign y9520 = ~n12987 ;
  assign y9521 = n12989 ;
  assign y9522 = ~n3008 ;
  assign y9523 = ~1'b0 ;
  assign y9524 = ~1'b0 ;
  assign y9525 = ~n12991 ;
  assign y9526 = ~n8995 ;
  assign y9527 = ~1'b0 ;
  assign y9528 = ~1'b0 ;
  assign y9529 = 1'b0 ;
  assign y9530 = ~n12992 ;
  assign y9531 = n12998 ;
  assign y9532 = ~1'b0 ;
  assign y9533 = n9252 ;
  assign y9534 = ~1'b0 ;
  assign y9535 = n12999 ;
  assign y9536 = ~n6818 ;
  assign y9537 = ~n8175 ;
  assign y9538 = n13000 ;
  assign y9539 = 1'b0 ;
  assign y9540 = ~1'b0 ;
  assign y9541 = ~n13005 ;
  assign y9542 = ~1'b0 ;
  assign y9543 = ~1'b0 ;
  assign y9544 = ~1'b0 ;
  assign y9545 = ~n13009 ;
  assign y9546 = n13010 ;
  assign y9547 = ~n5947 ;
  assign y9548 = ~n2856 ;
  assign y9549 = ~n13011 ;
  assign y9550 = ~1'b0 ;
  assign y9551 = ~n13013 ;
  assign y9552 = ~1'b0 ;
  assign y9553 = ~n13016 ;
  assign y9554 = ~1'b0 ;
  assign y9555 = n11299 ;
  assign y9556 = ~1'b0 ;
  assign y9557 = ~1'b0 ;
  assign y9558 = 1'b0 ;
  assign y9559 = ~1'b0 ;
  assign y9560 = ~n13019 ;
  assign y9561 = 1'b0 ;
  assign y9562 = ~n13021 ;
  assign y9563 = n13022 ;
  assign y9564 = ~1'b0 ;
  assign y9565 = 1'b0 ;
  assign y9566 = n13023 ;
  assign y9567 = ~n6046 ;
  assign y9568 = n13025 ;
  assign y9569 = n13027 ;
  assign y9570 = ~1'b0 ;
  assign y9571 = ~1'b0 ;
  assign y9572 = n2482 ;
  assign y9573 = n13028 ;
  assign y9574 = ~1'b0 ;
  assign y9575 = n13029 ;
  assign y9576 = n13032 ;
  assign y9577 = ~1'b0 ;
  assign y9578 = 1'b0 ;
  assign y9579 = n4193 ;
  assign y9580 = n13035 ;
  assign y9581 = ~1'b0 ;
  assign y9582 = ~1'b0 ;
  assign y9583 = n13037 ;
  assign y9584 = n13040 ;
  assign y9585 = ~n13042 ;
  assign y9586 = n13043 ;
  assign y9587 = ~n13048 ;
  assign y9588 = ~1'b0 ;
  assign y9589 = ~n13051 ;
  assign y9590 = ~1'b0 ;
  assign y9591 = n13052 ;
  assign y9592 = ~1'b0 ;
  assign y9593 = ~1'b0 ;
  assign y9594 = ~1'b0 ;
  assign y9595 = n13054 ;
  assign y9596 = ~n13064 ;
  assign y9597 = ~1'b0 ;
  assign y9598 = ~1'b0 ;
  assign y9599 = 1'b0 ;
  assign y9600 = n10837 ;
  assign y9601 = ~n13066 ;
  assign y9602 = ~n13067 ;
  assign y9603 = ~1'b0 ;
  assign y9604 = ~n13071 ;
  assign y9605 = ~n13072 ;
  assign y9606 = n13073 ;
  assign y9607 = ~n13076 ;
  assign y9608 = ~n13079 ;
  assign y9609 = ~1'b0 ;
  assign y9610 = n13080 ;
  assign y9611 = ~1'b0 ;
  assign y9612 = ~1'b0 ;
  assign y9613 = ~n13083 ;
  assign y9614 = ~n13086 ;
  assign y9615 = n13089 ;
  assign y9616 = ~n13091 ;
  assign y9617 = ~n13093 ;
  assign y9618 = ~1'b0 ;
  assign y9619 = ~n6875 ;
  assign y9620 = ~1'b0 ;
  assign y9621 = ~n13095 ;
  assign y9622 = n13104 ;
  assign y9623 = ~1'b0 ;
  assign y9624 = n13106 ;
  assign y9625 = n13109 ;
  assign y9626 = ~n13110 ;
  assign y9627 = ~1'b0 ;
  assign y9628 = n2321 ;
  assign y9629 = ~1'b0 ;
  assign y9630 = ~n227 ;
  assign y9631 = ~1'b0 ;
  assign y9632 = ~1'b0 ;
  assign y9633 = n5075 ;
  assign y9634 = n11671 ;
  assign y9635 = n13111 ;
  assign y9636 = 1'b0 ;
  assign y9637 = n13113 ;
  assign y9638 = 1'b0 ;
  assign y9639 = ~n13116 ;
  assign y9640 = ~n13118 ;
  assign y9641 = n13120 ;
  assign y9642 = n246 ;
  assign y9643 = n13125 ;
  assign y9644 = ~1'b0 ;
  assign y9645 = 1'b0 ;
  assign y9646 = ~n13126 ;
  assign y9647 = ~1'b0 ;
  assign y9648 = n12170 ;
  assign y9649 = ~n13128 ;
  assign y9650 = ~n13130 ;
  assign y9651 = ~n13139 ;
  assign y9652 = n13140 ;
  assign y9653 = ~n13149 ;
  assign y9654 = n13151 ;
  assign y9655 = ~1'b0 ;
  assign y9656 = ~1'b0 ;
  assign y9657 = n13153 ;
  assign y9658 = ~1'b0 ;
  assign y9659 = ~1'b0 ;
  assign y9660 = ~1'b0 ;
  assign y9661 = ~1'b0 ;
  assign y9662 = n13155 ;
  assign y9663 = n13156 ;
  assign y9664 = ~1'b0 ;
  assign y9665 = ~1'b0 ;
  assign y9666 = ~n13162 ;
  assign y9667 = n11965 ;
  assign y9668 = ~1'b0 ;
  assign y9669 = ~n13164 ;
  assign y9670 = n13168 ;
  assign y9671 = n13170 ;
  assign y9672 = ~n13171 ;
  assign y9673 = n13173 ;
  assign y9674 = ~n13174 ;
  assign y9675 = 1'b0 ;
  assign y9676 = ~n13177 ;
  assign y9677 = ~n13179 ;
  assign y9678 = ~n13181 ;
  assign y9679 = ~1'b0 ;
  assign y9680 = ~1'b0 ;
  assign y9681 = ~n13184 ;
  assign y9682 = ~n13188 ;
  assign y9683 = ~n13191 ;
  assign y9684 = ~1'b0 ;
  assign y9685 = n13194 ;
  assign y9686 = ~n13195 ;
  assign y9687 = n10282 ;
  assign y9688 = n13196 ;
  assign y9689 = 1'b0 ;
  assign y9690 = n13201 ;
  assign y9691 = n13204 ;
  assign y9692 = ~1'b0 ;
  assign y9693 = n13209 ;
  assign y9694 = ~n13217 ;
  assign y9695 = ~n13219 ;
  assign y9696 = ~1'b0 ;
  assign y9697 = 1'b0 ;
  assign y9698 = n8823 ;
  assign y9699 = n13223 ;
  assign y9700 = n13241 ;
  assign y9701 = ~n13250 ;
  assign y9702 = ~1'b0 ;
  assign y9703 = n13253 ;
  assign y9704 = n13261 ;
  assign y9705 = ~n13263 ;
  assign y9706 = ~1'b0 ;
  assign y9707 = n13265 ;
  assign y9708 = n13266 ;
  assign y9709 = ~n13268 ;
  assign y9710 = ~n13270 ;
  assign y9711 = ~n13275 ;
  assign y9712 = ~n13279 ;
  assign y9713 = ~1'b0 ;
  assign y9714 = ~n13282 ;
  assign y9715 = ~1'b0 ;
  assign y9716 = n3485 ;
  assign y9717 = ~1'b0 ;
  assign y9718 = ~1'b0 ;
  assign y9719 = ~n9195 ;
  assign y9720 = 1'b0 ;
  assign y9721 = ~1'b0 ;
  assign y9722 = ~1'b0 ;
  assign y9723 = ~n13283 ;
  assign y9724 = ~1'b0 ;
  assign y9725 = ~1'b0 ;
  assign y9726 = n13285 ;
  assign y9727 = n13291 ;
  assign y9728 = 1'b0 ;
  assign y9729 = ~n13292 ;
  assign y9730 = n13295 ;
  assign y9731 = n13298 ;
  assign y9732 = ~1'b0 ;
  assign y9733 = ~n13299 ;
  assign y9734 = ~n13301 ;
  assign y9735 = n13304 ;
  assign y9736 = ~n13306 ;
  assign y9737 = ~1'b0 ;
  assign y9738 = 1'b0 ;
  assign y9739 = ~n13310 ;
  assign y9740 = 1'b0 ;
  assign y9741 = ~1'b0 ;
  assign y9742 = ~n13312 ;
  assign y9743 = ~n13322 ;
  assign y9744 = n2166 ;
  assign y9745 = ~1'b0 ;
  assign y9746 = ~n13332 ;
  assign y9747 = ~n5481 ;
  assign y9748 = ~n13334 ;
  assign y9749 = ~n13336 ;
  assign y9750 = ~n12687 ;
  assign y9751 = ~1'b0 ;
  assign y9752 = n13337 ;
  assign y9753 = ~n13340 ;
  assign y9754 = ~n13341 ;
  assign y9755 = n13344 ;
  assign y9756 = ~1'b0 ;
  assign y9757 = n13346 ;
  assign y9758 = n13348 ;
  assign y9759 = ~n8629 ;
  assign y9760 = n9823 ;
  assign y9761 = ~n13352 ;
  assign y9762 = n13354 ;
  assign y9763 = ~n13356 ;
  assign y9764 = n13358 ;
  assign y9765 = n13359 ;
  assign y9766 = n13362 ;
  assign y9767 = n13363 ;
  assign y9768 = ~n13366 ;
  assign y9769 = n13367 ;
  assign y9770 = n13369 ;
  assign y9771 = ~1'b0 ;
  assign y9772 = ~1'b0 ;
  assign y9773 = ~n1157 ;
  assign y9774 = n13371 ;
  assign y9775 = ~n13372 ;
  assign y9776 = ~n13375 ;
  assign y9777 = ~1'b0 ;
  assign y9778 = ~n13377 ;
  assign y9779 = n13378 ;
  assign y9780 = n13379 ;
  assign y9781 = ~n13380 ;
  assign y9782 = n13382 ;
  assign y9783 = n5915 ;
  assign y9784 = ~n13386 ;
  assign y9785 = ~n13387 ;
  assign y9786 = ~1'b0 ;
  assign y9787 = n13388 ;
  assign y9788 = ~1'b0 ;
  assign y9789 = ~1'b0 ;
  assign y9790 = 1'b0 ;
  assign y9791 = 1'b0 ;
  assign y9792 = ~n6493 ;
  assign y9793 = ~n13389 ;
  assign y9794 = ~n13390 ;
  assign y9795 = n13395 ;
  assign y9796 = ~1'b0 ;
  assign y9797 = ~n13397 ;
  assign y9798 = ~1'b0 ;
  assign y9799 = ~1'b0 ;
  assign y9800 = ~n13398 ;
  assign y9801 = ~n13404 ;
  assign y9802 = n13411 ;
  assign y9803 = n9569 ;
  assign y9804 = ~1'b0 ;
  assign y9805 = ~n13414 ;
  assign y9806 = n13424 ;
  assign y9807 = ~n13427 ;
  assign y9808 = ~1'b0 ;
  assign y9809 = ~1'b0 ;
  assign y9810 = ~1'b0 ;
  assign y9811 = ~n13430 ;
  assign y9812 = ~1'b0 ;
  assign y9813 = n13434 ;
  assign y9814 = n977 ;
  assign y9815 = ~1'b0 ;
  assign y9816 = n13438 ;
  assign y9817 = ~n8764 ;
  assign y9818 = ~n13420 ;
  assign y9819 = ~n13439 ;
  assign y9820 = ~1'b0 ;
  assign y9821 = n13440 ;
  assign y9822 = ~1'b0 ;
  assign y9823 = ~n13443 ;
  assign y9824 = ~n11645 ;
  assign y9825 = ~n13444 ;
  assign y9826 = ~1'b0 ;
  assign y9827 = ~1'b0 ;
  assign y9828 = n13447 ;
  assign y9829 = ~1'b0 ;
  assign y9830 = ~n13449 ;
  assign y9831 = ~n13450 ;
  assign y9832 = ~n13455 ;
  assign y9833 = ~1'b0 ;
  assign y9834 = n13462 ;
  assign y9835 = ~1'b0 ;
  assign y9836 = 1'b0 ;
  assign y9837 = n13467 ;
  assign y9838 = ~1'b0 ;
  assign y9839 = n13473 ;
  assign y9840 = n13474 ;
  assign y9841 = n13476 ;
  assign y9842 = 1'b0 ;
  assign y9843 = ~n13478 ;
  assign y9844 = ~1'b0 ;
  assign y9845 = ~n158 ;
  assign y9846 = ~n13480 ;
  assign y9847 = n6444 ;
  assign y9848 = ~n1631 ;
  assign y9849 = ~n13481 ;
  assign y9850 = ~1'b0 ;
  assign y9851 = ~n13482 ;
  assign y9852 = n13485 ;
  assign y9853 = ~1'b0 ;
  assign y9854 = ~n13488 ;
  assign y9855 = ~n13492 ;
  assign y9856 = n13494 ;
  assign y9857 = ~n13518 ;
  assign y9858 = ~n13521 ;
  assign y9859 = ~n13526 ;
  assign y9860 = ~n13527 ;
  assign y9861 = ~n13528 ;
  assign y9862 = ~1'b0 ;
  assign y9863 = n517 ;
  assign y9864 = ~1'b0 ;
  assign y9865 = ~n10541 ;
  assign y9866 = n13530 ;
  assign y9867 = ~n13531 ;
  assign y9868 = ~n13532 ;
  assign y9869 = ~n13536 ;
  assign y9870 = ~n13540 ;
  assign y9871 = n13544 ;
  assign y9872 = ~1'b0 ;
  assign y9873 = n13547 ;
  assign y9874 = n13551 ;
  assign y9875 = ~1'b0 ;
  assign y9876 = 1'b0 ;
  assign y9877 = n13554 ;
  assign y9878 = ~1'b0 ;
  assign y9879 = n13555 ;
  assign y9880 = ~n13561 ;
  assign y9881 = n13566 ;
  assign y9882 = ~n13569 ;
  assign y9883 = ~n13571 ;
  assign y9884 = ~1'b0 ;
  assign y9885 = n13572 ;
  assign y9886 = n13576 ;
  assign y9887 = ~n13577 ;
  assign y9888 = ~1'b0 ;
  assign y9889 = n13578 ;
  assign y9890 = n7599 ;
  assign y9891 = 1'b0 ;
  assign y9892 = ~n13581 ;
  assign y9893 = ~1'b0 ;
  assign y9894 = ~1'b0 ;
  assign y9895 = ~1'b0 ;
  assign y9896 = n13584 ;
  assign y9897 = ~1'b0 ;
  assign y9898 = n13585 ;
  assign y9899 = ~1'b0 ;
  assign y9900 = ~1'b0 ;
  assign y9901 = ~1'b0 ;
  assign y9902 = n13586 ;
  assign y9903 = 1'b0 ;
  assign y9904 = ~n13590 ;
  assign y9905 = ~n13594 ;
  assign y9906 = ~n13595 ;
  assign y9907 = ~n13596 ;
  assign y9908 = 1'b0 ;
  assign y9909 = ~1'b0 ;
  assign y9910 = ~1'b0 ;
  assign y9911 = ~n1229 ;
  assign y9912 = n13597 ;
  assign y9913 = ~n13599 ;
  assign y9914 = ~1'b0 ;
  assign y9915 = ~1'b0 ;
  assign y9916 = ~n13600 ;
  assign y9917 = ~n13601 ;
  assign y9918 = ~1'b0 ;
  assign y9919 = n13607 ;
  assign y9920 = ~n5056 ;
  assign y9921 = ~n13611 ;
  assign y9922 = n13613 ;
  assign y9923 = ~1'b0 ;
  assign y9924 = ~1'b0 ;
  assign y9925 = ~n5111 ;
  assign y9926 = n12388 ;
  assign y9927 = ~1'b0 ;
  assign y9928 = ~1'b0 ;
  assign y9929 = ~1'b0 ;
  assign y9930 = ~1'b0 ;
  assign y9931 = ~1'b0 ;
  assign y9932 = ~1'b0 ;
  assign y9933 = n13614 ;
  assign y9934 = n13615 ;
  assign y9935 = n13617 ;
  assign y9936 = 1'b0 ;
  assign y9937 = ~1'b0 ;
  assign y9938 = n13618 ;
  assign y9939 = n13619 ;
  assign y9940 = n13043 ;
  assign y9941 = ~1'b0 ;
  assign y9942 = ~n1565 ;
  assign y9943 = n13620 ;
  assign y9944 = n13621 ;
  assign y9945 = n13622 ;
  assign y9946 = ~1'b0 ;
  assign y9947 = n13624 ;
  assign y9948 = ~n13626 ;
  assign y9949 = n13627 ;
  assign y9950 = ~1'b0 ;
  assign y9951 = ~1'b0 ;
  assign y9952 = n13633 ;
  assign y9953 = ~1'b0 ;
  assign y9954 = ~n13634 ;
  assign y9955 = ~n7933 ;
  assign y9956 = ~1'b0 ;
  assign y9957 = ~n1174 ;
  assign y9958 = n13635 ;
  assign y9959 = ~n13637 ;
  assign y9960 = ~1'b0 ;
  assign y9961 = ~1'b0 ;
  assign y9962 = n13639 ;
  assign y9963 = ~1'b0 ;
  assign y9964 = ~1'b0 ;
  assign y9965 = ~n13641 ;
  assign y9966 = n13644 ;
  assign y9967 = ~1'b0 ;
  assign y9968 = ~1'b0 ;
  assign y9969 = ~n13646 ;
  assign y9970 = ~n13648 ;
  assign y9971 = 1'b0 ;
  assign y9972 = 1'b0 ;
  assign y9973 = ~n13650 ;
  assign y9974 = n13654 ;
  assign y9975 = ~n13656 ;
  assign y9976 = ~n13657 ;
  assign y9977 = n13658 ;
  assign y9978 = n13663 ;
  assign y9979 = ~n13665 ;
  assign y9980 = ~n13667 ;
  assign y9981 = ~n9966 ;
  assign y9982 = ~1'b0 ;
  assign y9983 = ~1'b0 ;
  assign y9984 = ~n13670 ;
  assign y9985 = ~1'b0 ;
  assign y9986 = ~n13673 ;
  assign y9987 = ~1'b0 ;
  assign y9988 = ~1'b0 ;
  assign y9989 = ~1'b0 ;
  assign y9990 = ~n13676 ;
  assign y9991 = ~n13681 ;
  assign y9992 = ~n13683 ;
  assign y9993 = ~n13685 ;
  assign y9994 = n13686 ;
  assign y9995 = ~1'b0 ;
  assign y9996 = ~n13687 ;
  assign y9997 = n13688 ;
  assign y9998 = ~1'b0 ;
  assign y9999 = ~1'b0 ;
  assign y10000 = ~n13689 ;
  assign y10001 = n13690 ;
  assign y10002 = n13694 ;
  assign y10003 = ~1'b0 ;
  assign y10004 = n13696 ;
  assign y10005 = ~1'b0 ;
  assign y10006 = ~n882 ;
  assign y10007 = ~n13698 ;
  assign y10008 = ~n11272 ;
  assign y10009 = ~1'b0 ;
  assign y10010 = ~1'b0 ;
  assign y10011 = n13699 ;
  assign y10012 = ~1'b0 ;
  assign y10013 = n5141 ;
  assign y10014 = ~1'b0 ;
  assign y10015 = ~1'b0 ;
  assign y10016 = ~1'b0 ;
  assign y10017 = ~n13702 ;
  assign y10018 = ~n13707 ;
  assign y10019 = ~n13599 ;
  assign y10020 = ~n13708 ;
  assign y10021 = 1'b0 ;
  assign y10022 = ~1'b0 ;
  assign y10023 = ~1'b0 ;
  assign y10024 = n13710 ;
  assign y10025 = n4221 ;
  assign y10026 = ~n13711 ;
  assign y10027 = ~1'b0 ;
  assign y10028 = n13714 ;
  assign y10029 = ~n82 ;
  assign y10030 = ~1'b0 ;
  assign y10031 = n13719 ;
  assign y10032 = ~1'b0 ;
  assign y10033 = ~n13720 ;
  assign y10034 = ~1'b0 ;
  assign y10035 = ~1'b0 ;
  assign y10036 = n13721 ;
  assign y10037 = ~1'b0 ;
  assign y10038 = ~n13726 ;
  assign y10039 = ~n13729 ;
  assign y10040 = ~n13735 ;
  assign y10041 = ~1'b0 ;
  assign y10042 = ~1'b0 ;
  assign y10043 = ~1'b0 ;
  assign y10044 = n13737 ;
  assign y10045 = ~n13738 ;
  assign y10046 = ~n13741 ;
  assign y10047 = ~n13742 ;
  assign y10048 = ~1'b0 ;
  assign y10049 = ~1'b0 ;
  assign y10050 = ~n6764 ;
  assign y10051 = n13745 ;
  assign y10052 = ~1'b0 ;
  assign y10053 = ~n13747 ;
  assign y10054 = n13749 ;
  assign y10055 = n13751 ;
  assign y10056 = ~n8135 ;
  assign y10057 = ~n13753 ;
  assign y10058 = ~n13755 ;
  assign y10059 = ~1'b0 ;
  assign y10060 = ~1'b0 ;
  assign y10061 = n13758 ;
  assign y10062 = ~n3604 ;
  assign y10063 = n13759 ;
  assign y10064 = ~1'b0 ;
  assign y10065 = ~n13760 ;
  assign y10066 = n13761 ;
  assign y10067 = ~1'b0 ;
  assign y10068 = n13762 ;
  assign y10069 = ~n13771 ;
  assign y10070 = ~1'b0 ;
  assign y10071 = ~n13772 ;
  assign y10072 = ~n5823 ;
  assign y10073 = n13773 ;
  assign y10074 = n13776 ;
  assign y10075 = ~1'b0 ;
  assign y10076 = ~n13777 ;
  assign y10077 = ~1'b0 ;
  assign y10078 = n7079 ;
  assign y10079 = n13784 ;
  assign y10080 = n13791 ;
  assign y10081 = ~1'b0 ;
  assign y10082 = n13792 ;
  assign y10083 = ~n13793 ;
  assign y10084 = ~n13799 ;
  assign y10085 = ~n13801 ;
  assign y10086 = 1'b0 ;
  assign y10087 = n13803 ;
  assign y10088 = ~n7512 ;
  assign y10089 = n13805 ;
  assign y10090 = ~n13808 ;
  assign y10091 = ~n13810 ;
  assign y10092 = n13811 ;
  assign y10093 = ~1'b0 ;
  assign y10094 = 1'b0 ;
  assign y10095 = ~1'b0 ;
  assign y10096 = ~n13815 ;
  assign y10097 = n13817 ;
  assign y10098 = ~1'b0 ;
  assign y10099 = ~1'b0 ;
  assign y10100 = ~n13819 ;
  assign y10101 = n13820 ;
  assign y10102 = ~n13821 ;
  assign y10103 = ~1'b0 ;
  assign y10104 = ~1'b0 ;
  assign y10105 = ~1'b0 ;
  assign y10106 = n13824 ;
  assign y10107 = ~n612 ;
  assign y10108 = ~1'b0 ;
  assign y10109 = ~1'b0 ;
  assign y10110 = n13827 ;
  assign y10111 = ~1'b0 ;
  assign y10112 = n13828 ;
  assign y10113 = ~1'b0 ;
  assign y10114 = ~n13829 ;
  assign y10115 = n7904 ;
  assign y10116 = ~n353 ;
  assign y10117 = ~1'b0 ;
  assign y10118 = n13831 ;
  assign y10119 = n13832 ;
  assign y10120 = ~1'b0 ;
  assign y10121 = ~1'b0 ;
  assign y10122 = ~n13836 ;
  assign y10123 = ~1'b0 ;
  assign y10124 = ~1'b0 ;
  assign y10125 = n1008 ;
  assign y10126 = n13838 ;
  assign y10127 = n13841 ;
  assign y10128 = n13842 ;
  assign y10129 = n13843 ;
  assign y10130 = n13844 ;
  assign y10131 = n13845 ;
  assign y10132 = ~1'b0 ;
  assign y10133 = ~n13846 ;
  assign y10134 = ~n13848 ;
  assign y10135 = ~n2923 ;
  assign y10136 = n13851 ;
  assign y10137 = n13852 ;
  assign y10138 = n13853 ;
  assign y10139 = ~1'b0 ;
  assign y10140 = ~n13854 ;
  assign y10141 = ~1'b0 ;
  assign y10142 = n13859 ;
  assign y10143 = ~1'b0 ;
  assign y10144 = ~n13864 ;
  assign y10145 = ~n13865 ;
  assign y10146 = n13867 ;
  assign y10147 = 1'b0 ;
  assign y10148 = ~n13870 ;
  assign y10149 = ~n13875 ;
  assign y10150 = ~n13876 ;
  assign y10151 = ~n3037 ;
  assign y10152 = ~n13878 ;
  assign y10153 = n3946 ;
  assign y10154 = ~n13879 ;
  assign y10155 = ~1'b0 ;
  assign y10156 = n13882 ;
  assign y10157 = ~n13883 ;
  assign y10158 = n10567 ;
  assign y10159 = n13884 ;
  assign y10160 = ~n13885 ;
  assign y10161 = ~n13887 ;
  assign y10162 = ~1'b0 ;
  assign y10163 = ~1'b0 ;
  assign y10164 = ~1'b0 ;
  assign y10165 = n13888 ;
  assign y10166 = n13890 ;
  assign y10167 = ~n13892 ;
  assign y10168 = n13893 ;
  assign y10169 = n13895 ;
  assign y10170 = n13896 ;
  assign y10171 = n13900 ;
  assign y10172 = ~1'b0 ;
  assign y10173 = ~1'b0 ;
  assign y10174 = n13901 ;
  assign y10175 = ~n13903 ;
  assign y10176 = ~1'b0 ;
  assign y10177 = ~1'b0 ;
  assign y10178 = n13904 ;
  assign y10179 = ~1'b0 ;
  assign y10180 = ~1'b0 ;
  assign y10181 = n13906 ;
  assign y10182 = ~1'b0 ;
  assign y10183 = ~n10589 ;
  assign y10184 = n13907 ;
  assign y10185 = ~n13911 ;
  assign y10186 = ~1'b0 ;
  assign y10187 = ~n13913 ;
  assign y10188 = ~1'b0 ;
  assign y10189 = ~n13915 ;
  assign y10190 = ~1'b0 ;
  assign y10191 = n13918 ;
  assign y10192 = 1'b0 ;
  assign y10193 = ~n13921 ;
  assign y10194 = 1'b0 ;
  assign y10195 = ~n8392 ;
  assign y10196 = ~n13923 ;
  assign y10197 = ~n13924 ;
  assign y10198 = n13925 ;
  assign y10199 = ~1'b0 ;
  assign y10200 = n13929 ;
  assign y10201 = ~1'b0 ;
  assign y10202 = ~n13930 ;
  assign y10203 = 1'b0 ;
  assign y10204 = ~1'b0 ;
  assign y10205 = n13931 ;
  assign y10206 = n13937 ;
  assign y10207 = ~n13939 ;
  assign y10208 = ~1'b0 ;
  assign y10209 = ~1'b0 ;
  assign y10210 = ~n13941 ;
  assign y10211 = n13945 ;
  assign y10212 = ~1'b0 ;
  assign y10213 = n13946 ;
  assign y10214 = n13947 ;
  assign y10215 = n13951 ;
  assign y10216 = 1'b0 ;
  assign y10217 = ~1'b0 ;
  assign y10218 = ~1'b0 ;
  assign y10219 = n13952 ;
  assign y10220 = ~1'b0 ;
  assign y10221 = ~1'b0 ;
  assign y10222 = n13953 ;
  assign y10223 = n13954 ;
  assign y10224 = ~1'b0 ;
  assign y10225 = ~1'b0 ;
  assign y10226 = ~1'b0 ;
  assign y10227 = n13957 ;
  assign y10228 = n13962 ;
  assign y10229 = n13963 ;
  assign y10230 = n13964 ;
  assign y10231 = n13970 ;
  assign y10232 = n13971 ;
  assign y10233 = n13973 ;
  assign y10234 = ~n13979 ;
  assign y10235 = ~1'b0 ;
  assign y10236 = 1'b0 ;
  assign y10237 = ~n13984 ;
  assign y10238 = ~1'b0 ;
  assign y10239 = n13986 ;
  assign y10240 = ~n13990 ;
  assign y10241 = ~n13994 ;
  assign y10242 = n13999 ;
  assign y10243 = ~1'b0 ;
  assign y10244 = ~n14003 ;
  assign y10245 = n14005 ;
  assign y10246 = n14007 ;
  assign y10247 = n5011 ;
  assign y10248 = n14035 ;
  assign y10249 = n14036 ;
  assign y10250 = ~n14045 ;
  assign y10251 = ~n14050 ;
  assign y10252 = n14052 ;
  assign y10253 = n14053 ;
  assign y10254 = n14055 ;
  assign y10255 = ~n14056 ;
  assign y10256 = ~1'b0 ;
  assign y10257 = n14057 ;
  assign y10258 = n14062 ;
  assign y10259 = n14063 ;
  assign y10260 = ~1'b0 ;
  assign y10261 = n14064 ;
  assign y10262 = ~1'b0 ;
  assign y10263 = ~n14067 ;
  assign y10264 = ~1'b0 ;
  assign y10265 = n14068 ;
  assign y10266 = ~1'b0 ;
  assign y10267 = ~1'b0 ;
  assign y10268 = n414 ;
  assign y10269 = n14069 ;
  assign y10270 = ~1'b0 ;
  assign y10271 = ~1'b0 ;
  assign y10272 = ~1'b0 ;
  assign y10273 = ~n2291 ;
  assign y10274 = ~n14071 ;
  assign y10275 = ~n14072 ;
  assign y10276 = ~1'b0 ;
  assign y10277 = n14073 ;
  assign y10278 = ~n14074 ;
  assign y10279 = ~1'b0 ;
  assign y10280 = ~1'b0 ;
  assign y10281 = n14078 ;
  assign y10282 = ~n14082 ;
  assign y10283 = ~n14084 ;
  assign y10284 = ~1'b0 ;
  assign y10285 = ~n14088 ;
  assign y10286 = ~n14091 ;
  assign y10287 = n14092 ;
  assign y10288 = ~n14093 ;
  assign y10289 = ~n14095 ;
  assign y10290 = ~1'b0 ;
  assign y10291 = n14096 ;
  assign y10292 = ~1'b0 ;
  assign y10293 = n12293 ;
  assign y10294 = n917 ;
  assign y10295 = ~1'b0 ;
  assign y10296 = ~1'b0 ;
  assign y10297 = n14102 ;
  assign y10298 = ~n14108 ;
  assign y10299 = n14112 ;
  assign y10300 = ~n14115 ;
  assign y10301 = ~n14120 ;
  assign y10302 = n14126 ;
  assign y10303 = ~1'b0 ;
  assign y10304 = ~1'b0 ;
  assign y10305 = ~1'b0 ;
  assign y10306 = n14129 ;
  assign y10307 = n14133 ;
  assign y10308 = ~1'b0 ;
  assign y10309 = n14135 ;
  assign y10310 = ~1'b0 ;
  assign y10311 = n14141 ;
  assign y10312 = n14143 ;
  assign y10313 = ~1'b0 ;
  assign y10314 = n14144 ;
  assign y10315 = n14147 ;
  assign y10316 = ~n14148 ;
  assign y10317 = ~n14149 ;
  assign y10318 = 1'b0 ;
  assign y10319 = ~n8653 ;
  assign y10320 = ~1'b0 ;
  assign y10321 = 1'b0 ;
  assign y10322 = n14152 ;
  assign y10323 = 1'b0 ;
  assign y10324 = n14153 ;
  assign y10325 = ~n14157 ;
  assign y10326 = ~1'b0 ;
  assign y10327 = n14158 ;
  assign y10328 = n14159 ;
  assign y10329 = 1'b0 ;
  assign y10330 = ~1'b0 ;
  assign y10331 = ~1'b0 ;
  assign y10332 = ~1'b0 ;
  assign y10333 = n14160 ;
  assign y10334 = ~1'b0 ;
  assign y10335 = n14162 ;
  assign y10336 = n14165 ;
  assign y10337 = ~1'b0 ;
  assign y10338 = n14166 ;
  assign y10339 = ~n14169 ;
  assign y10340 = 1'b0 ;
  assign y10341 = n14170 ;
  assign y10342 = n14177 ;
  assign y10343 = ~n14182 ;
  assign y10344 = n14184 ;
  assign y10345 = ~1'b0 ;
  assign y10346 = ~n14187 ;
  assign y10347 = ~1'b0 ;
  assign y10348 = ~n14190 ;
  assign y10349 = ~1'b0 ;
  assign y10350 = n14192 ;
  assign y10351 = n14194 ;
  assign y10352 = ~1'b0 ;
  assign y10353 = ~1'b0 ;
  assign y10354 = ~1'b0 ;
  assign y10355 = n14202 ;
  assign y10356 = ~1'b0 ;
  assign y10357 = ~1'b0 ;
  assign y10358 = ~n14204 ;
  assign y10359 = ~1'b0 ;
  assign y10360 = n14207 ;
  assign y10361 = ~1'b0 ;
  assign y10362 = ~1'b0 ;
  assign y10363 = ~1'b0 ;
  assign y10364 = n2607 ;
  assign y10365 = ~n14208 ;
  assign y10366 = n14209 ;
  assign y10367 = n14210 ;
  assign y10368 = ~n1840 ;
  assign y10369 = ~n14215 ;
  assign y10370 = n14217 ;
  assign y10371 = ~1'b0 ;
  assign y10372 = n14218 ;
  assign y10373 = n6775 ;
  assign y10374 = n9747 ;
  assign y10375 = ~1'b0 ;
  assign y10376 = ~1'b0 ;
  assign y10377 = ~n14224 ;
  assign y10378 = ~n14228 ;
  assign y10379 = ~n3791 ;
  assign y10380 = ~1'b0 ;
  assign y10381 = ~n14229 ;
  assign y10382 = ~1'b0 ;
  assign y10383 = ~n14231 ;
  assign y10384 = ~1'b0 ;
  assign y10385 = ~n14233 ;
  assign y10386 = n6633 ;
  assign y10387 = ~n14235 ;
  assign y10388 = n364 ;
  assign y10389 = n374 ;
  assign y10390 = ~1'b0 ;
  assign y10391 = 1'b0 ;
  assign y10392 = 1'b0 ;
  assign y10393 = ~1'b0 ;
  assign y10394 = ~n14240 ;
  assign y10395 = n14241 ;
  assign y10396 = ~n14243 ;
  assign y10397 = ~n14245 ;
  assign y10398 = ~n14246 ;
  assign y10399 = ~n14248 ;
  assign y10400 = n14249 ;
  assign y10401 = n14251 ;
  assign y10402 = ~1'b0 ;
  assign y10403 = n14253 ;
  assign y10404 = 1'b0 ;
  assign y10405 = ~1'b0 ;
  assign y10406 = ~n14255 ;
  assign y10407 = ~n14256 ;
  assign y10408 = ~n14259 ;
  assign y10409 = ~n7008 ;
  assign y10410 = ~n14260 ;
  assign y10411 = n14261 ;
  assign y10412 = ~1'b0 ;
  assign y10413 = ~1'b0 ;
  assign y10414 = ~1'b0 ;
  assign y10415 = n14262 ;
  assign y10416 = 1'b0 ;
  assign y10417 = ~n14264 ;
  assign y10418 = ~1'b0 ;
  assign y10419 = ~n14268 ;
  assign y10420 = ~n14269 ;
  assign y10421 = n14270 ;
  assign y10422 = ~n14274 ;
  assign y10423 = n14275 ;
  assign y10424 = ~n14277 ;
  assign y10425 = ~n14278 ;
  assign y10426 = 1'b0 ;
  assign y10427 = n14279 ;
  assign y10428 = ~1'b0 ;
  assign y10429 = ~n10378 ;
  assign y10430 = ~n14301 ;
  assign y10431 = ~1'b0 ;
  assign y10432 = ~1'b0 ;
  assign y10433 = ~n14304 ;
  assign y10434 = ~n14305 ;
  assign y10435 = ~n12708 ;
  assign y10436 = n14309 ;
  assign y10437 = n14310 ;
  assign y10438 = n14312 ;
  assign y10439 = ~1'b0 ;
  assign y10440 = n14313 ;
  assign y10441 = ~n216 ;
  assign y10442 = ~1'b0 ;
  assign y10443 = ~n14315 ;
  assign y10444 = ~1'b0 ;
  assign y10445 = 1'b0 ;
  assign y10446 = n14323 ;
  assign y10447 = ~1'b0 ;
  assign y10448 = n14325 ;
  assign y10449 = ~1'b0 ;
  assign y10450 = n14329 ;
  assign y10451 = ~n14343 ;
  assign y10452 = n14346 ;
  assign y10453 = ~n14348 ;
  assign y10454 = ~n14349 ;
  assign y10455 = ~n14350 ;
  assign y10456 = n14355 ;
  assign y10457 = ~n7886 ;
  assign y10458 = n14356 ;
  assign y10459 = ~n14358 ;
  assign y10460 = ~n14360 ;
  assign y10461 = n14367 ;
  assign y10462 = ~1'b0 ;
  assign y10463 = 1'b0 ;
  assign y10464 = n14369 ;
  assign y10465 = ~1'b0 ;
  assign y10466 = ~1'b0 ;
  assign y10467 = ~1'b0 ;
  assign y10468 = 1'b0 ;
  assign y10469 = ~n3032 ;
  assign y10470 = ~1'b0 ;
  assign y10471 = ~n14370 ;
  assign y10472 = ~1'b0 ;
  assign y10473 = n14371 ;
  assign y10474 = 1'b0 ;
  assign y10475 = ~n14372 ;
  assign y10476 = n14385 ;
  assign y10477 = ~1'b0 ;
  assign y10478 = ~n14386 ;
  assign y10479 = n14391 ;
  assign y10480 = n14392 ;
  assign y10481 = ~1'b0 ;
  assign y10482 = ~1'b0 ;
  assign y10483 = 1'b0 ;
  assign y10484 = ~1'b0 ;
  assign y10485 = ~1'b0 ;
  assign y10486 = ~1'b0 ;
  assign y10487 = n14393 ;
  assign y10488 = 1'b0 ;
  assign y10489 = ~n1804 ;
  assign y10490 = n14394 ;
  assign y10491 = ~n14395 ;
  assign y10492 = ~1'b0 ;
  assign y10493 = ~n14396 ;
  assign y10494 = ~1'b0 ;
  assign y10495 = ~1'b0 ;
  assign y10496 = ~1'b0 ;
  assign y10497 = ~1'b0 ;
  assign y10498 = n14397 ;
  assign y10499 = ~n14398 ;
  assign y10500 = ~n14400 ;
  assign y10501 = ~n4000 ;
  assign y10502 = n14401 ;
  assign y10503 = n14404 ;
  assign y10504 = ~1'b0 ;
  assign y10505 = ~n14410 ;
  assign y10506 = n14414 ;
  assign y10507 = n14415 ;
  assign y10508 = ~1'b0 ;
  assign y10509 = n14418 ;
  assign y10510 = ~1'b0 ;
  assign y10511 = ~1'b0 ;
  assign y10512 = n14420 ;
  assign y10513 = ~n14423 ;
  assign y10514 = ~n14424 ;
  assign y10515 = ~n6375 ;
  assign y10516 = ~n1175 ;
  assign y10517 = ~1'b0 ;
  assign y10518 = ~n14425 ;
  assign y10519 = ~n14427 ;
  assign y10520 = n14435 ;
  assign y10521 = n14436 ;
  assign y10522 = ~n14443 ;
  assign y10523 = ~1'b0 ;
  assign y10524 = ~n592 ;
  assign y10525 = ~1'b0 ;
  assign y10526 = n14445 ;
  assign y10527 = ~1'b0 ;
  assign y10528 = n7850 ;
  assign y10529 = ~1'b0 ;
  assign y10530 = ~1'b0 ;
  assign y10531 = ~n14448 ;
  assign y10532 = ~n14457 ;
  assign y10533 = n14458 ;
  assign y10534 = 1'b0 ;
  assign y10535 = n1958 ;
  assign y10536 = ~n14463 ;
  assign y10537 = n14469 ;
  assign y10538 = 1'b0 ;
  assign y10539 = ~1'b0 ;
  assign y10540 = n2546 ;
  assign y10541 = n14470 ;
  assign y10542 = 1'b0 ;
  assign y10543 = n14471 ;
  assign y10544 = ~1'b0 ;
  assign y10545 = n14473 ;
  assign y10546 = n14474 ;
  assign y10547 = n14476 ;
  assign y10548 = n14478 ;
  assign y10549 = ~n14483 ;
  assign y10550 = ~1'b0 ;
  assign y10551 = ~n14486 ;
  assign y10552 = ~1'b0 ;
  assign y10553 = n14488 ;
  assign y10554 = n14490 ;
  assign y10555 = n14491 ;
  assign y10556 = ~n14492 ;
  assign y10557 = ~1'b0 ;
  assign y10558 = ~n844 ;
  assign y10559 = ~n13578 ;
  assign y10560 = n11763 ;
  assign y10561 = n14495 ;
  assign y10562 = ~n14496 ;
  assign y10563 = ~1'b0 ;
  assign y10564 = ~n14498 ;
  assign y10565 = n1523 ;
  assign y10566 = ~n7360 ;
  assign y10567 = ~1'b0 ;
  assign y10568 = ~1'b0 ;
  assign y10569 = ~1'b0 ;
  assign y10570 = n14502 ;
  assign y10571 = ~1'b0 ;
  assign y10572 = ~1'b0 ;
  assign y10573 = ~n14512 ;
  assign y10574 = ~1'b0 ;
  assign y10575 = n14513 ;
  assign y10576 = ~n11405 ;
  assign y10577 = ~n14517 ;
  assign y10578 = ~1'b0 ;
  assign y10579 = ~1'b0 ;
  assign y10580 = n14520 ;
  assign y10581 = n14523 ;
  assign y10582 = ~n220 ;
  assign y10583 = ~1'b0 ;
  assign y10584 = ~n14528 ;
  assign y10585 = n14531 ;
  assign y10586 = ~1'b0 ;
  assign y10587 = n14532 ;
  assign y10588 = n14535 ;
  assign y10589 = ~n14536 ;
  assign y10590 = n14539 ;
  assign y10591 = ~n14541 ;
  assign y10592 = n14547 ;
  assign y10593 = ~1'b0 ;
  assign y10594 = n14549 ;
  assign y10595 = ~n14552 ;
  assign y10596 = n11698 ;
  assign y10597 = n14554 ;
  assign y10598 = ~1'b0 ;
  assign y10599 = ~1'b0 ;
  assign y10600 = ~n14556 ;
  assign y10601 = n14557 ;
  assign y10602 = ~n14559 ;
  assign y10603 = ~1'b0 ;
  assign y10604 = ~1'b0 ;
  assign y10605 = ~1'b0 ;
  assign y10606 = ~1'b0 ;
  assign y10607 = n14560 ;
  assign y10608 = ~1'b0 ;
  assign y10609 = ~n14561 ;
  assign y10610 = n14563 ;
  assign y10611 = ~1'b0 ;
  assign y10612 = ~n14564 ;
  assign y10613 = n14568 ;
  assign y10614 = ~1'b0 ;
  assign y10615 = n14570 ;
  assign y10616 = ~1'b0 ;
  assign y10617 = ~1'b0 ;
  assign y10618 = ~n14573 ;
  assign y10619 = n14574 ;
  assign y10620 = ~n3527 ;
  assign y10621 = ~1'b0 ;
  assign y10622 = n1441 ;
  assign y10623 = n14586 ;
  assign y10624 = ~1'b0 ;
  assign y10625 = ~n5779 ;
  assign y10626 = ~1'b0 ;
  assign y10627 = 1'b0 ;
  assign y10628 = n14587 ;
  assign y10629 = n14588 ;
  assign y10630 = ~n14591 ;
  assign y10631 = n14593 ;
  assign y10632 = ~1'b0 ;
  assign y10633 = ~1'b0 ;
  assign y10634 = ~1'b0 ;
  assign y10635 = n14595 ;
  assign y10636 = ~1'b0 ;
  assign y10637 = 1'b0 ;
  assign y10638 = ~1'b0 ;
  assign y10639 = ~1'b0 ;
  assign y10640 = ~1'b0 ;
  assign y10641 = ~1'b0 ;
  assign y10642 = n14600 ;
  assign y10643 = ~1'b0 ;
  assign y10644 = ~1'b0 ;
  assign y10645 = n14602 ;
  assign y10646 = ~n14603 ;
  assign y10647 = ~1'b0 ;
  assign y10648 = n14607 ;
  assign y10649 = n14612 ;
  assign y10650 = n14616 ;
  assign y10651 = n11479 ;
  assign y10652 = n14619 ;
  assign y10653 = n14620 ;
  assign y10654 = ~n14624 ;
  assign y10655 = 1'b0 ;
  assign y10656 = ~1'b0 ;
  assign y10657 = ~1'b0 ;
  assign y10658 = ~n865 ;
  assign y10659 = ~1'b0 ;
  assign y10660 = ~n14625 ;
  assign y10661 = n14639 ;
  assign y10662 = ~n14642 ;
  assign y10663 = n14644 ;
  assign y10664 = n14645 ;
  assign y10665 = n758 ;
  assign y10666 = n4937 ;
  assign y10667 = n14646 ;
  assign y10668 = n14649 ;
  assign y10669 = ~1'b0 ;
  assign y10670 = ~1'b0 ;
  assign y10671 = ~n14650 ;
  assign y10672 = ~1'b0 ;
  assign y10673 = ~n14651 ;
  assign y10674 = ~1'b0 ;
  assign y10675 = ~1'b0 ;
  assign y10676 = ~1'b0 ;
  assign y10677 = ~1'b0 ;
  assign y10678 = ~n14653 ;
  assign y10679 = ~n14654 ;
  assign y10680 = ~1'b0 ;
  assign y10681 = ~n13266 ;
  assign y10682 = n14657 ;
  assign y10683 = n14660 ;
  assign y10684 = n10352 ;
  assign y10685 = ~1'b0 ;
  assign y10686 = n14662 ;
  assign y10687 = n14664 ;
  assign y10688 = ~n14665 ;
  assign y10689 = n14667 ;
  assign y10690 = ~1'b0 ;
  assign y10691 = n14672 ;
  assign y10692 = ~1'b0 ;
  assign y10693 = n308 ;
  assign y10694 = ~n14674 ;
  assign y10695 = n661 ;
  assign y10696 = ~n14675 ;
  assign y10697 = n14676 ;
  assign y10698 = n14677 ;
  assign y10699 = ~1'b0 ;
  assign y10700 = ~n3774 ;
  assign y10701 = n14682 ;
  assign y10702 = n14684 ;
  assign y10703 = ~1'b0 ;
  assign y10704 = ~n14688 ;
  assign y10705 = ~n14692 ;
  assign y10706 = ~1'b0 ;
  assign y10707 = ~n14699 ;
  assign y10708 = ~n1316 ;
  assign y10709 = ~n14702 ;
  assign y10710 = ~1'b0 ;
  assign y10711 = ~1'b0 ;
  assign y10712 = ~1'b0 ;
  assign y10713 = ~n14708 ;
  assign y10714 = ~n14709 ;
  assign y10715 = n14710 ;
  assign y10716 = n13960 ;
  assign y10717 = ~n14715 ;
  assign y10718 = ~1'b0 ;
  assign y10719 = ~1'b0 ;
  assign y10720 = ~n14720 ;
  assign y10721 = n14721 ;
  assign y10722 = n14724 ;
  assign y10723 = n14725 ;
  assign y10724 = ~n14727 ;
  assign y10725 = ~n7227 ;
  assign y10726 = ~1'b0 ;
  assign y10727 = ~n14730 ;
  assign y10728 = ~1'b0 ;
  assign y10729 = ~1'b0 ;
  assign y10730 = n14732 ;
  assign y10731 = ~1'b0 ;
  assign y10732 = 1'b0 ;
  assign y10733 = n14733 ;
  assign y10734 = n14735 ;
  assign y10735 = n14736 ;
  assign y10736 = ~1'b0 ;
  assign y10737 = n14741 ;
  assign y10738 = n14744 ;
  assign y10739 = n7599 ;
  assign y10740 = n14745 ;
  assign y10741 = ~1'b0 ;
  assign y10742 = ~1'b0 ;
  assign y10743 = ~n14748 ;
  assign y10744 = n14757 ;
  assign y10745 = ~1'b0 ;
  assign y10746 = n14764 ;
  assign y10747 = ~1'b0 ;
  assign y10748 = ~1'b0 ;
  assign y10749 = n14765 ;
  assign y10750 = ~1'b0 ;
  assign y10751 = ~n1303 ;
  assign y10752 = ~n14766 ;
  assign y10753 = ~n14767 ;
  assign y10754 = n14768 ;
  assign y10755 = ~n14770 ;
  assign y10756 = ~1'b0 ;
  assign y10757 = n14771 ;
  assign y10758 = 1'b0 ;
  assign y10759 = n14084 ;
  assign y10760 = n14772 ;
  assign y10761 = 1'b0 ;
  assign y10762 = ~n14777 ;
  assign y10763 = ~1'b0 ;
  assign y10764 = ~n14779 ;
  assign y10765 = ~1'b0 ;
  assign y10766 = n10734 ;
  assign y10767 = ~1'b0 ;
  assign y10768 = ~1'b0 ;
  assign y10769 = n14782 ;
  assign y10770 = ~n4469 ;
  assign y10771 = ~n14786 ;
  assign y10772 = n2301 ;
  assign y10773 = ~n14788 ;
  assign y10774 = n14789 ;
  assign y10775 = 1'b0 ;
  assign y10776 = ~1'b0 ;
  assign y10777 = n14793 ;
  assign y10778 = ~n246 ;
  assign y10779 = ~n14798 ;
  assign y10780 = ~1'b0 ;
  assign y10781 = ~1'b0 ;
  assign y10782 = ~n5030 ;
  assign y10783 = ~1'b0 ;
  assign y10784 = n3077 ;
  assign y10785 = ~n14800 ;
  assign y10786 = n14803 ;
  assign y10787 = ~n14804 ;
  assign y10788 = ~1'b0 ;
  assign y10789 = n14811 ;
  assign y10790 = n14812 ;
  assign y10791 = ~n14813 ;
  assign y10792 = n14817 ;
  assign y10793 = ~n14822 ;
  assign y10794 = ~n7369 ;
  assign y10795 = ~n14422 ;
  assign y10796 = ~1'b0 ;
  assign y10797 = n14825 ;
  assign y10798 = ~n14826 ;
  assign y10799 = ~1'b0 ;
  assign y10800 = ~1'b0 ;
  assign y10801 = n14828 ;
  assign y10802 = ~1'b0 ;
  assign y10803 = ~1'b0 ;
  assign y10804 = n14832 ;
  assign y10805 = ~n14834 ;
  assign y10806 = ~1'b0 ;
  assign y10807 = ~n14836 ;
  assign y10808 = ~n3813 ;
  assign y10809 = ~n14839 ;
  assign y10810 = ~1'b0 ;
  assign y10811 = ~1'b0 ;
  assign y10812 = n14840 ;
  assign y10813 = ~1'b0 ;
  assign y10814 = ~1'b0 ;
  assign y10815 = ~n14844 ;
  assign y10816 = n14845 ;
  assign y10817 = ~n9490 ;
  assign y10818 = n14850 ;
  assign y10819 = ~1'b0 ;
  assign y10820 = ~1'b0 ;
  assign y10821 = ~1'b0 ;
  assign y10822 = ~n14852 ;
  assign y10823 = n14860 ;
  assign y10824 = ~n14862 ;
  assign y10825 = ~1'b0 ;
  assign y10826 = ~1'b0 ;
  assign y10827 = ~n14867 ;
  assign y10828 = ~n14876 ;
  assign y10829 = ~n14881 ;
  assign y10830 = ~1'b0 ;
  assign y10831 = n14882 ;
  assign y10832 = ~1'b0 ;
  assign y10833 = n14891 ;
  assign y10834 = ~n1772 ;
  assign y10835 = n14896 ;
  assign y10836 = ~n14897 ;
  assign y10837 = ~1'b0 ;
  assign y10838 = ~1'b0 ;
  assign y10839 = ~1'b0 ;
  assign y10840 = ~n14899 ;
  assign y10841 = ~1'b0 ;
  assign y10842 = ~1'b0 ;
  assign y10843 = n14901 ;
  assign y10844 = ~1'b0 ;
  assign y10845 = n7135 ;
  assign y10846 = ~n14905 ;
  assign y10847 = ~n14906 ;
  assign y10848 = ~1'b0 ;
  assign y10849 = ~n14907 ;
  assign y10850 = 1'b0 ;
  assign y10851 = ~1'b0 ;
  assign y10852 = 1'b0 ;
  assign y10853 = ~n14914 ;
  assign y10854 = n4840 ;
  assign y10855 = ~1'b0 ;
  assign y10856 = ~n14924 ;
  assign y10857 = n14929 ;
  assign y10858 = ~n14930 ;
  assign y10859 = 1'b0 ;
  assign y10860 = ~n14937 ;
  assign y10861 = ~1'b0 ;
  assign y10862 = n14942 ;
  assign y10863 = n6272 ;
  assign y10864 = n14943 ;
  assign y10865 = ~n14944 ;
  assign y10866 = ~n14945 ;
  assign y10867 = ~1'b0 ;
  assign y10868 = ~n10358 ;
  assign y10869 = ~1'b0 ;
  assign y10870 = n14947 ;
  assign y10871 = ~1'b0 ;
  assign y10872 = ~1'b0 ;
  assign y10873 = n14948 ;
  assign y10874 = ~n8705 ;
  assign y10875 = ~1'b0 ;
  assign y10876 = ~n14951 ;
  assign y10877 = n14957 ;
  assign y10878 = ~n14963 ;
  assign y10879 = ~n14966 ;
  assign y10880 = ~n14967 ;
  assign y10881 = ~1'b0 ;
  assign y10882 = ~1'b0 ;
  assign y10883 = ~1'b0 ;
  assign y10884 = ~n14971 ;
  assign y10885 = ~n14976 ;
  assign y10886 = n14978 ;
  assign y10887 = ~1'b0 ;
  assign y10888 = n14980 ;
  assign y10889 = n14982 ;
  assign y10890 = ~1'b0 ;
  assign y10891 = n14983 ;
  assign y10892 = n14986 ;
  assign y10893 = 1'b0 ;
  assign y10894 = ~1'b0 ;
  assign y10895 = ~1'b0 ;
  assign y10896 = n14987 ;
  assign y10897 = ~1'b0 ;
  assign y10898 = ~1'b0 ;
  assign y10899 = ~n14988 ;
  assign y10900 = 1'b0 ;
  assign y10901 = n14990 ;
  assign y10902 = ~1'b0 ;
  assign y10903 = n14992 ;
  assign y10904 = ~n14998 ;
  assign y10905 = ~n15002 ;
  assign y10906 = 1'b0 ;
  assign y10907 = n15004 ;
  assign y10908 = n2939 ;
  assign y10909 = ~n15005 ;
  assign y10910 = n15010 ;
  assign y10911 = n6900 ;
  assign y10912 = ~1'b0 ;
  assign y10913 = n15012 ;
  assign y10914 = ~1'b0 ;
  assign y10915 = 1'b0 ;
  assign y10916 = ~n15013 ;
  assign y10917 = n15014 ;
  assign y10918 = ~n12252 ;
  assign y10919 = ~n15016 ;
  assign y10920 = ~1'b0 ;
  assign y10921 = n15020 ;
  assign y10922 = n15021 ;
  assign y10923 = n15025 ;
  assign y10924 = ~1'b0 ;
  assign y10925 = n15026 ;
  assign y10926 = ~1'b0 ;
  assign y10927 = ~n15029 ;
  assign y10928 = n12421 ;
  assign y10929 = ~1'b0 ;
  assign y10930 = n15032 ;
  assign y10931 = ~1'b0 ;
  assign y10932 = n15033 ;
  assign y10933 = ~n15040 ;
  assign y10934 = ~1'b0 ;
  assign y10935 = ~1'b0 ;
  assign y10936 = 1'b0 ;
  assign y10937 = n15043 ;
  assign y10938 = ~1'b0 ;
  assign y10939 = n15045 ;
  assign y10940 = n7668 ;
  assign y10941 = ~n15048 ;
  assign y10942 = ~n5409 ;
  assign y10943 = ~1'b0 ;
  assign y10944 = ~n542 ;
  assign y10945 = n15056 ;
  assign y10946 = 1'b0 ;
  assign y10947 = n15057 ;
  assign y10948 = n15058 ;
  assign y10949 = ~1'b0 ;
  assign y10950 = ~n5573 ;
  assign y10951 = ~1'b0 ;
  assign y10952 = n15062 ;
  assign y10953 = ~1'b0 ;
  assign y10954 = ~n5205 ;
  assign y10955 = n5905 ;
  assign y10956 = ~n15063 ;
  assign y10957 = ~n15067 ;
  assign y10958 = ~n4022 ;
  assign y10959 = ~n15068 ;
  assign y10960 = ~n15071 ;
  assign y10961 = ~1'b0 ;
  assign y10962 = ~n15075 ;
  assign y10963 = ~1'b0 ;
  assign y10964 = ~n15077 ;
  assign y10965 = ~n678 ;
  assign y10966 = ~n6322 ;
  assign y10967 = 1'b0 ;
  assign y10968 = ~n15078 ;
  assign y10969 = ~n15086 ;
  assign y10970 = 1'b0 ;
  assign y10971 = n15093 ;
  assign y10972 = ~n15095 ;
  assign y10973 = n9544 ;
  assign y10974 = ~1'b0 ;
  assign y10975 = ~1'b0 ;
  assign y10976 = n15096 ;
  assign y10977 = ~n15097 ;
  assign y10978 = n15101 ;
  assign y10979 = ~n15105 ;
  assign y10980 = ~1'b0 ;
  assign y10981 = ~n15108 ;
  assign y10982 = ~n6714 ;
  assign y10983 = ~1'b0 ;
  assign y10984 = ~n15109 ;
  assign y10985 = ~1'b0 ;
  assign y10986 = ~1'b0 ;
  assign y10987 = n1851 ;
  assign y10988 = ~n15114 ;
  assign y10989 = ~1'b0 ;
  assign y10990 = n15115 ;
  assign y10991 = ~1'b0 ;
  assign y10992 = ~1'b0 ;
  assign y10993 = ~n15116 ;
  assign y10994 = n15119 ;
  assign y10995 = ~n15121 ;
  assign y10996 = 1'b0 ;
  assign y10997 = ~1'b0 ;
  assign y10998 = n15122 ;
  assign y10999 = ~1'b0 ;
  assign y11000 = ~1'b0 ;
  assign y11001 = n15126 ;
  assign y11002 = ~1'b0 ;
  assign y11003 = n15128 ;
  assign y11004 = ~n15132 ;
  assign y11005 = 1'b0 ;
  assign y11006 = ~n15134 ;
  assign y11007 = ~n15135 ;
  assign y11008 = n15137 ;
  assign y11009 = ~n15139 ;
  assign y11010 = ~n15144 ;
  assign y11011 = 1'b0 ;
  assign y11012 = ~1'b0 ;
  assign y11013 = n15146 ;
  assign y11014 = ~n15151 ;
  assign y11015 = ~n4075 ;
  assign y11016 = ~n15152 ;
  assign y11017 = n3318 ;
  assign y11018 = n9523 ;
  assign y11019 = 1'b0 ;
  assign y11020 = ~n15154 ;
  assign y11021 = ~n15156 ;
  assign y11022 = ~1'b0 ;
  assign y11023 = ~1'b0 ;
  assign y11024 = ~1'b0 ;
  assign y11025 = 1'b0 ;
  assign y11026 = ~1'b0 ;
  assign y11027 = ~1'b0 ;
  assign y11028 = ~n15157 ;
  assign y11029 = ~n8206 ;
  assign y11030 = ~n15161 ;
  assign y11031 = ~1'b0 ;
  assign y11032 = n11866 ;
  assign y11033 = 1'b0 ;
  assign y11034 = n15162 ;
  assign y11035 = ~n15163 ;
  assign y11036 = ~n15166 ;
  assign y11037 = ~1'b0 ;
  assign y11038 = n15168 ;
  assign y11039 = n15169 ;
  assign y11040 = n15172 ;
  assign y11041 = n2589 ;
  assign y11042 = ~1'b0 ;
  assign y11043 = n15175 ;
  assign y11044 = ~n15177 ;
  assign y11045 = n15181 ;
  assign y11046 = ~1'b0 ;
  assign y11047 = ~n15185 ;
  assign y11048 = ~n15189 ;
  assign y11049 = ~1'b0 ;
  assign y11050 = n246 ;
  assign y11051 = ~1'b0 ;
  assign y11052 = n15191 ;
  assign y11053 = ~n15192 ;
  assign y11054 = ~n11235 ;
  assign y11055 = ~1'b0 ;
  assign y11056 = ~1'b0 ;
  assign y11057 = ~1'b0 ;
  assign y11058 = n15193 ;
  assign y11059 = ~n15194 ;
  assign y11060 = ~1'b0 ;
  assign y11061 = ~1'b0 ;
  assign y11062 = n15196 ;
  assign y11063 = ~1'b0 ;
  assign y11064 = ~1'b0 ;
  assign y11065 = ~1'b0 ;
  assign y11066 = ~1'b0 ;
  assign y11067 = n15199 ;
  assign y11068 = ~1'b0 ;
  assign y11069 = ~n10423 ;
  assign y11070 = n15205 ;
  assign y11071 = ~1'b0 ;
  assign y11072 = ~n15207 ;
  assign y11073 = ~1'b0 ;
  assign y11074 = n15208 ;
  assign y11075 = ~1'b0 ;
  assign y11076 = ~n15212 ;
  assign y11077 = ~1'b0 ;
  assign y11078 = ~1'b0 ;
  assign y11079 = ~n13689 ;
  assign y11080 = ~1'b0 ;
  assign y11081 = ~n15214 ;
  assign y11082 = ~n15218 ;
  assign y11083 = 1'b0 ;
  assign y11084 = ~n7181 ;
  assign y11085 = ~1'b0 ;
  assign y11086 = ~1'b0 ;
  assign y11087 = ~n37 ;
  assign y11088 = 1'b0 ;
  assign y11089 = ~n15222 ;
  assign y11090 = n15223 ;
  assign y11091 = 1'b0 ;
  assign y11092 = 1'b0 ;
  assign y11093 = ~1'b0 ;
  assign y11094 = n15224 ;
  assign y11095 = ~n15229 ;
  assign y11096 = 1'b0 ;
  assign y11097 = ~n1316 ;
  assign y11098 = ~n15231 ;
  assign y11099 = ~n15232 ;
  assign y11100 = ~1'b0 ;
  assign y11101 = ~1'b0 ;
  assign y11102 = ~1'b0 ;
  assign y11103 = n15233 ;
  assign y11104 = ~1'b0 ;
  assign y11105 = ~1'b0 ;
  assign y11106 = ~n15240 ;
  assign y11107 = ~n15241 ;
  assign y11108 = ~1'b0 ;
  assign y11109 = ~1'b0 ;
  assign y11110 = n15244 ;
  assign y11111 = n9143 ;
  assign y11112 = ~n15245 ;
  assign y11113 = ~n15246 ;
  assign y11114 = ~1'b0 ;
  assign y11115 = ~1'b0 ;
  assign y11116 = ~n15249 ;
  assign y11117 = ~1'b0 ;
  assign y11118 = n15252 ;
  assign y11119 = ~n15256 ;
  assign y11120 = ~n15258 ;
  assign y11121 = ~n83 ;
  assign y11122 = n15261 ;
  assign y11123 = ~n15262 ;
  assign y11124 = n15263 ;
  assign y11125 = ~1'b0 ;
  assign y11126 = n15265 ;
  assign y11127 = ~n15266 ;
  assign y11128 = n15271 ;
  assign y11129 = 1'b0 ;
  assign y11130 = ~1'b0 ;
  assign y11131 = n15273 ;
  assign y11132 = n15274 ;
  assign y11133 = n15276 ;
  assign y11134 = ~1'b0 ;
  assign y11135 = ~n15278 ;
  assign y11136 = ~n15281 ;
  assign y11137 = ~n15284 ;
  assign y11138 = ~1'b0 ;
  assign y11139 = n15285 ;
  assign y11140 = 1'b0 ;
  assign y11141 = ~1'b0 ;
  assign y11142 = n15287 ;
  assign y11143 = ~1'b0 ;
  assign y11144 = ~1'b0 ;
  assign y11145 = ~n15289 ;
  assign y11146 = ~n15291 ;
  assign y11147 = n15292 ;
  assign y11148 = ~n15294 ;
  assign y11149 = ~n9447 ;
  assign y11150 = n3687 ;
  assign y11151 = ~1'b0 ;
  assign y11152 = ~n15297 ;
  assign y11153 = 1'b0 ;
  assign y11154 = n15298 ;
  assign y11155 = n15299 ;
  assign y11156 = n15300 ;
  assign y11157 = n15302 ;
  assign y11158 = ~1'b0 ;
  assign y11159 = 1'b0 ;
  assign y11160 = ~n15304 ;
  assign y11161 = 1'b0 ;
  assign y11162 = ~1'b0 ;
  assign y11163 = 1'b0 ;
  assign y11164 = ~n15307 ;
  assign y11165 = n15308 ;
  assign y11166 = ~n15309 ;
  assign y11167 = n15310 ;
  assign y11168 = ~n4526 ;
  assign y11169 = ~1'b0 ;
  assign y11170 = ~n15312 ;
  assign y11171 = ~n15318 ;
  assign y11172 = ~1'b0 ;
  assign y11173 = ~n15319 ;
  assign y11174 = ~n15325 ;
  assign y11175 = ~n15326 ;
  assign y11176 = n15328 ;
  assign y11177 = ~n15329 ;
  assign y11178 = ~1'b0 ;
  assign y11179 = n15330 ;
  assign y11180 = n15332 ;
  assign y11181 = ~n15333 ;
  assign y11182 = ~n15361 ;
  assign y11183 = ~n364 ;
  assign y11184 = n15362 ;
  assign y11185 = n15364 ;
  assign y11186 = 1'b0 ;
  assign y11187 = 1'b0 ;
  assign y11188 = ~n15366 ;
  assign y11189 = ~1'b0 ;
  assign y11190 = n15372 ;
  assign y11191 = 1'b0 ;
  assign y11192 = ~x10 ;
  assign y11193 = ~1'b0 ;
  assign y11194 = ~n15379 ;
  assign y11195 = ~1'b0 ;
  assign y11196 = n15380 ;
  assign y11197 = ~1'b0 ;
  assign y11198 = ~n15381 ;
  assign y11199 = ~1'b0 ;
  assign y11200 = ~n15385 ;
  assign y11201 = ~n15394 ;
  assign y11202 = ~n15398 ;
  assign y11203 = 1'b0 ;
  assign y11204 = n15399 ;
  assign y11205 = ~1'b0 ;
  assign y11206 = n15400 ;
  assign y11207 = n15403 ;
  assign y11208 = ~1'b0 ;
  assign y11209 = ~1'b0 ;
  assign y11210 = ~1'b0 ;
  assign y11211 = ~n15404 ;
  assign y11212 = ~1'b0 ;
  assign y11213 = n15406 ;
  assign y11214 = n13656 ;
  assign y11215 = n15407 ;
  assign y11216 = ~1'b0 ;
  assign y11217 = ~n15409 ;
  assign y11218 = ~n15410 ;
  assign y11219 = ~1'b0 ;
  assign y11220 = ~1'b0 ;
  assign y11221 = n15411 ;
  assign y11222 = 1'b0 ;
  assign y11223 = ~1'b0 ;
  assign y11224 = n15412 ;
  assign y11225 = ~n15414 ;
  assign y11226 = n15415 ;
  assign y11227 = n15418 ;
  assign y11228 = ~1'b0 ;
  assign y11229 = 1'b0 ;
  assign y11230 = n2235 ;
  assign y11231 = n15419 ;
  assign y11232 = n15424 ;
  assign y11233 = ~1'b0 ;
  assign y11234 = n15426 ;
  assign y11235 = ~1'b0 ;
  assign y11236 = ~1'b0 ;
  assign y11237 = ~1'b0 ;
  assign y11238 = ~1'b0 ;
  assign y11239 = ~1'b0 ;
  assign y11240 = ~n4552 ;
  assign y11241 = n15427 ;
  assign y11242 = ~1'b0 ;
  assign y11243 = n15430 ;
  assign y11244 = ~n2324 ;
  assign y11245 = ~n15433 ;
  assign y11246 = n15434 ;
  assign y11247 = n15435 ;
  assign y11248 = n15437 ;
  assign y11249 = 1'b0 ;
  assign y11250 = ~n15441 ;
  assign y11251 = ~1'b0 ;
  assign y11252 = ~n15444 ;
  assign y11253 = ~n15448 ;
  assign y11254 = n15451 ;
  assign y11255 = n15454 ;
  assign y11256 = n15455 ;
  assign y11257 = ~n13682 ;
  assign y11258 = n15456 ;
  assign y11259 = ~1'b0 ;
  assign y11260 = ~1'b0 ;
  assign y11261 = ~n15457 ;
  assign y11262 = n15458 ;
  assign y11263 = ~n15459 ;
  assign y11264 = 1'b0 ;
  assign y11265 = ~1'b0 ;
  assign y11266 = ~n15461 ;
  assign y11267 = n15463 ;
  assign y11268 = n15465 ;
  assign y11269 = ~n15467 ;
  assign y11270 = ~1'b0 ;
  assign y11271 = n15468 ;
  assign y11272 = n3368 ;
  assign y11273 = ~1'b0 ;
  assign y11274 = n13083 ;
  assign y11275 = ~n15469 ;
  assign y11276 = ~1'b0 ;
  assign y11277 = n15476 ;
  assign y11278 = ~n15478 ;
  assign y11279 = n1995 ;
  assign y11280 = ~1'b0 ;
  assign y11281 = ~n15479 ;
  assign y11282 = n15480 ;
  assign y11283 = ~1'b0 ;
  assign y11284 = ~n15481 ;
  assign y11285 = ~1'b0 ;
  assign y11286 = n15483 ;
  assign y11287 = n15484 ;
  assign y11288 = ~1'b0 ;
  assign y11289 = ~1'b0 ;
  assign y11290 = ~n15488 ;
  assign y11291 = ~1'b0 ;
  assign y11292 = ~n15490 ;
  assign y11293 = ~1'b0 ;
  assign y11294 = ~n15493 ;
  assign y11295 = n15495 ;
  assign y11296 = n15497 ;
  assign y11297 = n15499 ;
  assign y11298 = n15507 ;
  assign y11299 = ~1'b0 ;
  assign y11300 = ~n15512 ;
  assign y11301 = n15514 ;
  assign y11302 = ~1'b0 ;
  assign y11303 = ~n15518 ;
  assign y11304 = n15519 ;
  assign y11305 = 1'b0 ;
  assign y11306 = ~n15520 ;
  assign y11307 = n15525 ;
  assign y11308 = ~n15529 ;
  assign y11309 = ~1'b0 ;
  assign y11310 = 1'b0 ;
  assign y11311 = 1'b0 ;
  assign y11312 = ~1'b0 ;
  assign y11313 = ~1'b0 ;
  assign y11314 = ~n15533 ;
  assign y11315 = n15534 ;
  assign y11316 = ~1'b0 ;
  assign y11317 = ~1'b0 ;
  assign y11318 = n15541 ;
  assign y11319 = ~n15542 ;
  assign y11320 = ~1'b0 ;
  assign y11321 = ~1'b0 ;
  assign y11322 = n8763 ;
  assign y11323 = ~1'b0 ;
  assign y11324 = ~n15543 ;
  assign y11325 = ~n15546 ;
  assign y11326 = n15552 ;
  assign y11327 = ~1'b0 ;
  assign y11328 = ~n15555 ;
  assign y11329 = ~n15557 ;
  assign y11330 = 1'b0 ;
  assign y11331 = ~n15559 ;
  assign y11332 = ~1'b0 ;
  assign y11333 = n15560 ;
  assign y11334 = ~1'b0 ;
  assign y11335 = ~n15569 ;
  assign y11336 = n15572 ;
  assign y11337 = n15574 ;
  assign y11338 = n15577 ;
  assign y11339 = n15579 ;
  assign y11340 = ~1'b0 ;
  assign y11341 = n15583 ;
  assign y11342 = ~n15588 ;
  assign y11343 = n15591 ;
  assign y11344 = ~n15595 ;
  assign y11345 = ~n15597 ;
  assign y11346 = ~n15600 ;
  assign y11347 = ~n15605 ;
  assign y11348 = ~x3 ;
  assign y11349 = ~1'b0 ;
  assign y11350 = n15606 ;
  assign y11351 = ~1'b0 ;
  assign y11352 = ~1'b0 ;
  assign y11353 = ~1'b0 ;
  assign y11354 = ~n15611 ;
  assign y11355 = ~n15614 ;
  assign y11356 = n7572 ;
  assign y11357 = n15615 ;
  assign y11358 = ~1'b0 ;
  assign y11359 = n15618 ;
  assign y11360 = ~1'b0 ;
  assign y11361 = ~1'b0 ;
  assign y11362 = ~n15623 ;
  assign y11363 = ~n15624 ;
  assign y11364 = ~1'b0 ;
  assign y11365 = n11535 ;
  assign y11366 = ~1'b0 ;
  assign y11367 = n15625 ;
  assign y11368 = n15626 ;
  assign y11369 = ~n15627 ;
  assign y11370 = ~1'b0 ;
  assign y11371 = n15631 ;
  assign y11372 = ~1'b0 ;
  assign y11373 = ~1'b0 ;
  assign y11374 = ~n15633 ;
  assign y11375 = ~1'b0 ;
  assign y11376 = n639 ;
  assign y11377 = n15635 ;
  assign y11378 = ~n15637 ;
  assign y11379 = ~1'b0 ;
  assign y11380 = ~n5947 ;
  assign y11381 = n15639 ;
  assign y11382 = ~n10223 ;
  assign y11383 = n15642 ;
  assign y11384 = ~n15644 ;
  assign y11385 = ~1'b0 ;
  assign y11386 = n15648 ;
  assign y11387 = n15649 ;
  assign y11388 = n1117 ;
  assign y11389 = ~n15655 ;
  assign y11390 = ~n15137 ;
  assign y11391 = ~n15657 ;
  assign y11392 = ~n15659 ;
  assign y11393 = ~n15664 ;
  assign y11394 = ~n15670 ;
  assign y11395 = ~1'b0 ;
  assign y11396 = ~1'b0 ;
  assign y11397 = n15671 ;
  assign y11398 = ~1'b0 ;
  assign y11399 = ~n8820 ;
  assign y11400 = ~1'b0 ;
  assign y11401 = ~n4189 ;
  assign y11402 = ~1'b0 ;
  assign y11403 = ~1'b0 ;
  assign y11404 = n15672 ;
  assign y11405 = n15675 ;
  assign y11406 = ~1'b0 ;
  assign y11407 = n15676 ;
  assign y11408 = ~1'b0 ;
  assign y11409 = ~1'b0 ;
  assign y11410 = n15057 ;
  assign y11411 = ~1'b0 ;
  assign y11412 = ~n15677 ;
  assign y11413 = n15678 ;
  assign y11414 = n15680 ;
  assign y11415 = n13886 ;
  assign y11416 = ~n15682 ;
  assign y11417 = ~1'b0 ;
  assign y11418 = ~1'b0 ;
  assign y11419 = ~n15683 ;
  assign y11420 = ~n15684 ;
  assign y11421 = n4357 ;
  assign y11422 = n10805 ;
  assign y11423 = n15686 ;
  assign y11424 = ~n15688 ;
  assign y11425 = ~n15689 ;
  assign y11426 = ~1'b0 ;
  assign y11427 = n15690 ;
  assign y11428 = n15691 ;
  assign y11429 = ~n15694 ;
  assign y11430 = ~n15696 ;
  assign y11431 = ~1'b0 ;
  assign y11432 = n10080 ;
  assign y11433 = ~1'b0 ;
  assign y11434 = ~1'b0 ;
  assign y11435 = n15697 ;
  assign y11436 = ~1'b0 ;
  assign y11437 = n15701 ;
  assign y11438 = ~1'b0 ;
  assign y11439 = ~1'b0 ;
  assign y11440 = ~n15705 ;
  assign y11441 = n15706 ;
  assign y11442 = ~n15707 ;
  assign y11443 = 1'b0 ;
  assign y11444 = ~1'b0 ;
  assign y11445 = n15709 ;
  assign y11446 = ~1'b0 ;
  assign y11447 = ~1'b0 ;
  assign y11448 = 1'b0 ;
  assign y11449 = ~n15712 ;
  assign y11450 = ~n15713 ;
  assign y11451 = ~n15714 ;
  assign y11452 = n15715 ;
  assign y11453 = ~n15720 ;
  assign y11454 = n15721 ;
  assign y11455 = ~1'b0 ;
  assign y11456 = ~1'b0 ;
  assign y11457 = ~1'b0 ;
  assign y11458 = ~1'b0 ;
  assign y11459 = ~1'b0 ;
  assign y11460 = ~n15723 ;
  assign y11461 = n15724 ;
  assign y11462 = ~n15747 ;
  assign y11463 = ~1'b0 ;
  assign y11464 = ~1'b0 ;
  assign y11465 = n15749 ;
  assign y11466 = n15750 ;
  assign y11467 = ~1'b0 ;
  assign y11468 = n15760 ;
  assign y11469 = ~1'b0 ;
  assign y11470 = n15761 ;
  assign y11471 = ~1'b0 ;
  assign y11472 = ~n15766 ;
  assign y11473 = ~n15768 ;
  assign y11474 = ~1'b0 ;
  assign y11475 = n15773 ;
  assign y11476 = ~1'b0 ;
  assign y11477 = ~1'b0 ;
  assign y11478 = ~1'b0 ;
  assign y11479 = ~n15781 ;
  assign y11480 = ~1'b0 ;
  assign y11481 = ~1'b0 ;
  assign y11482 = ~n15782 ;
  assign y11483 = 1'b0 ;
  assign y11484 = ~1'b0 ;
  assign y11485 = n6770 ;
  assign y11486 = ~1'b0 ;
  assign y11487 = ~n15784 ;
  assign y11488 = ~1'b0 ;
  assign y11489 = ~n15786 ;
  assign y11490 = ~n15797 ;
  assign y11491 = n741 ;
  assign y11492 = ~1'b0 ;
  assign y11493 = ~1'b0 ;
  assign y11494 = n15799 ;
  assign y11495 = ~n15801 ;
  assign y11496 = ~1'b0 ;
  assign y11497 = n15802 ;
  assign y11498 = ~1'b0 ;
  assign y11499 = ~n15804 ;
  assign y11500 = n15811 ;
  assign y11501 = ~1'b0 ;
  assign y11502 = ~1'b0 ;
  assign y11503 = n15812 ;
  assign y11504 = ~n15816 ;
  assign y11505 = n15818 ;
  assign y11506 = ~n2547 ;
  assign y11507 = ~1'b0 ;
  assign y11508 = ~1'b0 ;
  assign y11509 = 1'b0 ;
  assign y11510 = n9751 ;
  assign y11511 = ~n15822 ;
  assign y11512 = ~1'b0 ;
  assign y11513 = ~n15823 ;
  assign y11514 = ~1'b0 ;
  assign y11515 = ~1'b0 ;
  assign y11516 = ~1'b0 ;
  assign y11517 = ~1'b0 ;
  assign y11518 = ~1'b0 ;
  assign y11519 = ~1'b0 ;
  assign y11520 = ~n15835 ;
  assign y11521 = ~1'b0 ;
  assign y11522 = ~n15838 ;
  assign y11523 = ~1'b0 ;
  assign y11524 = n15840 ;
  assign y11525 = n15842 ;
  assign y11526 = 1'b0 ;
  assign y11527 = ~1'b0 ;
  assign y11528 = ~1'b0 ;
  assign y11529 = n15844 ;
  assign y11530 = ~1'b0 ;
  assign y11531 = n15847 ;
  assign y11532 = ~n10876 ;
  assign y11533 = n15851 ;
  assign y11534 = ~n15857 ;
  assign y11535 = ~n15862 ;
  assign y11536 = ~1'b0 ;
  assign y11537 = n15863 ;
  assign y11538 = ~n15864 ;
  assign y11539 = ~1'b0 ;
  assign y11540 = 1'b0 ;
  assign y11541 = ~n15867 ;
  assign y11542 = ~n15871 ;
  assign y11543 = ~1'b0 ;
  assign y11544 = n15872 ;
  assign y11545 = n15875 ;
  assign y11546 = ~n15878 ;
  assign y11547 = ~n15890 ;
  assign y11548 = ~1'b0 ;
  assign y11549 = ~1'b0 ;
  assign y11550 = n15894 ;
  assign y11551 = n15895 ;
  assign y11552 = n15897 ;
  assign y11553 = ~1'b0 ;
  assign y11554 = ~1'b0 ;
  assign y11555 = n15902 ;
  assign y11556 = n15904 ;
  assign y11557 = ~n7981 ;
  assign y11558 = ~1'b0 ;
  assign y11559 = ~n15905 ;
  assign y11560 = ~1'b0 ;
  assign y11561 = 1'b0 ;
  assign y11562 = ~n15909 ;
  assign y11563 = ~1'b0 ;
  assign y11564 = n15913 ;
  assign y11565 = n15918 ;
  assign y11566 = ~1'b0 ;
  assign y11567 = ~1'b0 ;
  assign y11568 = n12440 ;
  assign y11569 = ~1'b0 ;
  assign y11570 = ~1'b0 ;
  assign y11571 = ~n15920 ;
  assign y11572 = ~1'b0 ;
  assign y11573 = ~n15925 ;
  assign y11574 = ~1'b0 ;
  assign y11575 = ~n15926 ;
  assign y11576 = ~1'b0 ;
  assign y11577 = ~1'b0 ;
  assign y11578 = n15928 ;
  assign y11579 = ~1'b0 ;
  assign y11580 = ~1'b0 ;
  assign y11581 = ~n1687 ;
  assign y11582 = ~n15930 ;
  assign y11583 = ~n15932 ;
  assign y11584 = n12972 ;
  assign y11585 = ~1'b0 ;
  assign y11586 = ~n15933 ;
  assign y11587 = ~n15948 ;
  assign y11588 = n15952 ;
  assign y11589 = ~1'b0 ;
  assign y11590 = ~n15958 ;
  assign y11591 = ~n15959 ;
  assign y11592 = ~n15960 ;
  assign y11593 = ~1'b0 ;
  assign y11594 = ~1'b0 ;
  assign y11595 = ~1'b0 ;
  assign y11596 = ~n15963 ;
  assign y11597 = ~n9745 ;
  assign y11598 = ~1'b0 ;
  assign y11599 = n15965 ;
  assign y11600 = n2842 ;
  assign y11601 = ~1'b0 ;
  assign y11602 = ~1'b0 ;
  assign y11603 = n15966 ;
  assign y11604 = ~n15977 ;
  assign y11605 = ~1'b0 ;
  assign y11606 = ~1'b0 ;
  assign y11607 = n15978 ;
  assign y11608 = ~1'b0 ;
  assign y11609 = ~n15979 ;
  assign y11610 = ~n15985 ;
  assign y11611 = n15991 ;
  assign y11612 = ~1'b0 ;
  assign y11613 = ~n15992 ;
  assign y11614 = ~1'b0 ;
  assign y11615 = ~1'b0 ;
  assign y11616 = n15994 ;
  assign y11617 = n16004 ;
  assign y11618 = n16007 ;
  assign y11619 = ~1'b0 ;
  assign y11620 = 1'b0 ;
  assign y11621 = ~1'b0 ;
  assign y11622 = ~1'b0 ;
  assign y11623 = ~n16009 ;
  assign y11624 = ~1'b0 ;
  assign y11625 = ~n16010 ;
  assign y11626 = n16018 ;
  assign y11627 = n16022 ;
  assign y11628 = ~n16024 ;
  assign y11629 = ~1'b0 ;
  assign y11630 = ~1'b0 ;
  assign y11631 = n14539 ;
  assign y11632 = ~1'b0 ;
  assign y11633 = ~1'b0 ;
  assign y11634 = n2912 ;
  assign y11635 = n11100 ;
  assign y11636 = ~1'b0 ;
  assign y11637 = ~n16027 ;
  assign y11638 = ~n16029 ;
  assign y11639 = ~1'b0 ;
  assign y11640 = n9155 ;
  assign y11641 = n16030 ;
  assign y11642 = n16031 ;
  assign y11643 = n233 ;
  assign y11644 = n16032 ;
  assign y11645 = ~n16035 ;
  assign y11646 = ~n16036 ;
  assign y11647 = ~1'b0 ;
  assign y11648 = ~n16040 ;
  assign y11649 = 1'b0 ;
  assign y11650 = n16042 ;
  assign y11651 = ~n16046 ;
  assign y11652 = ~1'b0 ;
  assign y11653 = ~1'b0 ;
  assign y11654 = ~1'b0 ;
  assign y11655 = ~1'b0 ;
  assign y11656 = 1'b0 ;
  assign y11657 = ~n16047 ;
  assign y11658 = ~n7597 ;
  assign y11659 = n16050 ;
  assign y11660 = ~n12343 ;
  assign y11661 = ~1'b0 ;
  assign y11662 = n16054 ;
  assign y11663 = ~1'b0 ;
  assign y11664 = ~1'b0 ;
  assign y11665 = ~1'b0 ;
  assign y11666 = ~n16055 ;
  assign y11667 = ~n16057 ;
  assign y11668 = ~1'b0 ;
  assign y11669 = ~1'b0 ;
  assign y11670 = 1'b0 ;
  assign y11671 = 1'b0 ;
  assign y11672 = ~1'b0 ;
  assign y11673 = ~1'b0 ;
  assign y11674 = ~n16058 ;
  assign y11675 = ~n16062 ;
  assign y11676 = ~n16064 ;
  assign y11677 = ~1'b0 ;
  assign y11678 = ~n16066 ;
  assign y11679 = n16067 ;
  assign y11680 = ~1'b0 ;
  assign y11681 = ~1'b0 ;
  assign y11682 = ~n16069 ;
  assign y11683 = n16073 ;
  assign y11684 = ~n16074 ;
  assign y11685 = ~1'b0 ;
  assign y11686 = ~1'b0 ;
  assign y11687 = ~1'b0 ;
  assign y11688 = ~n16076 ;
  assign y11689 = ~n16082 ;
  assign y11690 = n16084 ;
  assign y11691 = ~n16090 ;
  assign y11692 = ~n16092 ;
  assign y11693 = ~1'b0 ;
  assign y11694 = ~1'b0 ;
  assign y11695 = n16095 ;
  assign y11696 = n16098 ;
  assign y11697 = ~n16099 ;
  assign y11698 = ~1'b0 ;
  assign y11699 = ~1'b0 ;
  assign y11700 = n7714 ;
  assign y11701 = ~1'b0 ;
  assign y11702 = n16101 ;
  assign y11703 = ~n16102 ;
  assign y11704 = ~1'b0 ;
  assign y11705 = ~1'b0 ;
  assign y11706 = ~1'b0 ;
  assign y11707 = ~1'b0 ;
  assign y11708 = ~1'b0 ;
  assign y11709 = ~1'b0 ;
  assign y11710 = ~1'b0 ;
  assign y11711 = 1'b0 ;
  assign y11712 = ~1'b0 ;
  assign y11713 = ~1'b0 ;
  assign y11714 = n16104 ;
  assign y11715 = ~1'b0 ;
  assign y11716 = n16107 ;
  assign y11717 = ~1'b0 ;
  assign y11718 = ~n16057 ;
  assign y11719 = n16110 ;
  assign y11720 = ~1'b0 ;
  assign y11721 = ~n16117 ;
  assign y11722 = n16118 ;
  assign y11723 = n16119 ;
  assign y11724 = ~n16122 ;
  assign y11725 = ~1'b0 ;
  assign y11726 = ~n16126 ;
  assign y11727 = ~n16127 ;
  assign y11728 = 1'b0 ;
  assign y11729 = n16130 ;
  assign y11730 = ~n16132 ;
  assign y11731 = ~n16133 ;
  assign y11732 = ~n588 ;
  assign y11733 = ~n16135 ;
  assign y11734 = ~n16137 ;
  assign y11735 = n16141 ;
  assign y11736 = ~n16143 ;
  assign y11737 = ~n16145 ;
  assign y11738 = ~n16146 ;
  assign y11739 = ~1'b0 ;
  assign y11740 = n16147 ;
  assign y11741 = ~n16150 ;
  assign y11742 = ~1'b0 ;
  assign y11743 = n395 ;
  assign y11744 = n16151 ;
  assign y11745 = n16155 ;
  assign y11746 = n16156 ;
  assign y11747 = 1'b0 ;
  assign y11748 = n16157 ;
  assign y11749 = n16160 ;
  assign y11750 = ~n16162 ;
  assign y11751 = ~1'b0 ;
  assign y11752 = ~1'b0 ;
  assign y11753 = ~1'b0 ;
  assign y11754 = ~n5465 ;
  assign y11755 = ~n16163 ;
  assign y11756 = ~1'b0 ;
  assign y11757 = ~1'b0 ;
  assign y11758 = n16164 ;
  assign y11759 = ~n16166 ;
  assign y11760 = ~n2326 ;
  assign y11761 = n16167 ;
  assign y11762 = ~1'b0 ;
  assign y11763 = n16168 ;
  assign y11764 = ~n16173 ;
  assign y11765 = ~n16176 ;
  assign y11766 = ~n16180 ;
  assign y11767 = n16182 ;
  assign y11768 = ~n16184 ;
  assign y11769 = ~1'b0 ;
  assign y11770 = ~1'b0 ;
  assign y11771 = ~n16185 ;
  assign y11772 = ~n16188 ;
  assign y11773 = ~n16190 ;
  assign y11774 = ~1'b0 ;
  assign y11775 = n16194 ;
  assign y11776 = n4231 ;
  assign y11777 = n16196 ;
  assign y11778 = ~n16198 ;
  assign y11779 = 1'b0 ;
  assign y11780 = n16202 ;
  assign y11781 = ~1'b0 ;
  assign y11782 = ~n16203 ;
  assign y11783 = ~n16206 ;
  assign y11784 = ~n16207 ;
  assign y11785 = n16211 ;
  assign y11786 = ~n16216 ;
  assign y11787 = ~1'b0 ;
  assign y11788 = 1'b0 ;
  assign y11789 = ~n16218 ;
  assign y11790 = n16219 ;
  assign y11791 = n16221 ;
  assign y11792 = ~n16224 ;
  assign y11793 = ~n16228 ;
  assign y11794 = ~n16231 ;
  assign y11795 = ~1'b0 ;
  assign y11796 = ~1'b0 ;
  assign y11797 = ~n16235 ;
  assign y11798 = 1'b0 ;
  assign y11799 = ~1'b0 ;
  assign y11800 = n16236 ;
  assign y11801 = n16237 ;
  assign y11802 = n16240 ;
  assign y11803 = ~n16242 ;
  assign y11804 = n16243 ;
  assign y11805 = ~n16246 ;
  assign y11806 = ~n16247 ;
  assign y11807 = ~n16249 ;
  assign y11808 = ~1'b0 ;
  assign y11809 = ~n16253 ;
  assign y11810 = ~n2922 ;
  assign y11811 = n16255 ;
  assign y11812 = ~1'b0 ;
  assign y11813 = ~1'b0 ;
  assign y11814 = 1'b0 ;
  assign y11815 = ~n13870 ;
  assign y11816 = n16257 ;
  assign y11817 = n16259 ;
  assign y11818 = n16260 ;
  assign y11819 = n16261 ;
  assign y11820 = n11039 ;
  assign y11821 = n16262 ;
  assign y11822 = n16263 ;
  assign y11823 = ~n16264 ;
  assign y11824 = n16266 ;
  assign y11825 = ~n16269 ;
  assign y11826 = n16272 ;
  assign y11827 = n16273 ;
  assign y11828 = ~1'b0 ;
  assign y11829 = ~1'b0 ;
  assign y11830 = ~1'b0 ;
  assign y11831 = ~1'b0 ;
  assign y11832 = ~n16275 ;
  assign y11833 = ~1'b0 ;
  assign y11834 = ~n16279 ;
  assign y11835 = ~1'b0 ;
  assign y11836 = ~n2914 ;
  assign y11837 = ~1'b0 ;
  assign y11838 = ~n16281 ;
  assign y11839 = n16286 ;
  assign y11840 = ~n4207 ;
  assign y11841 = n16289 ;
  assign y11842 = ~n16292 ;
  assign y11843 = n16294 ;
  assign y11844 = ~1'b0 ;
  assign y11845 = ~1'b0 ;
  assign y11846 = 1'b0 ;
  assign y11847 = ~1'b0 ;
  assign y11848 = n16295 ;
  assign y11849 = ~n16300 ;
  assign y11850 = ~1'b0 ;
  assign y11851 = n16301 ;
  assign y11852 = ~n16308 ;
  assign y11853 = ~n16309 ;
  assign y11854 = n16313 ;
  assign y11855 = ~n16315 ;
  assign y11856 = ~1'b0 ;
  assign y11857 = n16320 ;
  assign y11858 = n16321 ;
  assign y11859 = n16324 ;
  assign y11860 = n16325 ;
  assign y11861 = ~n16328 ;
  assign y11862 = ~n16330 ;
  assign y11863 = ~1'b0 ;
  assign y11864 = ~n16333 ;
  assign y11865 = ~1'b0 ;
  assign y11866 = ~n16334 ;
  assign y11867 = ~1'b0 ;
  assign y11868 = n16335 ;
  assign y11869 = n16336 ;
  assign y11870 = ~n16338 ;
  assign y11871 = ~1'b0 ;
  assign y11872 = n16339 ;
  assign y11873 = ~1'b0 ;
  assign y11874 = ~n16340 ;
  assign y11875 = n16343 ;
  assign y11876 = ~1'b0 ;
  assign y11877 = ~n16346 ;
  assign y11878 = ~n16347 ;
  assign y11879 = ~1'b0 ;
  assign y11880 = n16351 ;
  assign y11881 = n16353 ;
  assign y11882 = ~1'b0 ;
  assign y11883 = n16354 ;
  assign y11884 = ~1'b0 ;
  assign y11885 = n16355 ;
  assign y11886 = ~n15598 ;
  assign y11887 = ~1'b0 ;
  assign y11888 = n16338 ;
  assign y11889 = ~n9739 ;
  assign y11890 = ~n16357 ;
  assign y11891 = n16359 ;
  assign y11892 = ~1'b0 ;
  assign y11893 = n8262 ;
  assign y11894 = ~1'b0 ;
  assign y11895 = n16360 ;
  assign y11896 = ~n16362 ;
  assign y11897 = ~1'b0 ;
  assign y11898 = ~1'b0 ;
  assign y11899 = ~1'b0 ;
  assign y11900 = n9185 ;
  assign y11901 = n2800 ;
  assign y11902 = n16365 ;
  assign y11903 = ~1'b0 ;
  assign y11904 = ~1'b0 ;
  assign y11905 = ~n16368 ;
  assign y11906 = 1'b0 ;
  assign y11907 = ~1'b0 ;
  assign y11908 = ~1'b0 ;
  assign y11909 = ~1'b0 ;
  assign y11910 = ~1'b0 ;
  assign y11911 = ~1'b0 ;
  assign y11912 = ~1'b0 ;
  assign y11913 = ~n16370 ;
  assign y11914 = ~n1572 ;
  assign y11915 = 1'b0 ;
  assign y11916 = ~n16371 ;
  assign y11917 = 1'b0 ;
  assign y11918 = ~n16375 ;
  assign y11919 = ~n16377 ;
  assign y11920 = ~1'b0 ;
  assign y11921 = ~1'b0 ;
  assign y11922 = n16381 ;
  assign y11923 = ~1'b0 ;
  assign y11924 = ~1'b0 ;
  assign y11925 = n16384 ;
  assign y11926 = ~n11309 ;
  assign y11927 = ~1'b0 ;
  assign y11928 = ~n16389 ;
  assign y11929 = ~n16397 ;
  assign y11930 = n16398 ;
  assign y11931 = ~n16400 ;
  assign y11932 = n16403 ;
  assign y11933 = n16404 ;
  assign y11934 = ~1'b0 ;
  assign y11935 = ~1'b0 ;
  assign y11936 = ~n11027 ;
  assign y11937 = ~n16406 ;
  assign y11938 = ~n16409 ;
  assign y11939 = n16411 ;
  assign y11940 = ~n16412 ;
  assign y11941 = ~n16415 ;
  assign y11942 = n16417 ;
  assign y11943 = ~n16420 ;
  assign y11944 = ~1'b0 ;
  assign y11945 = ~n16421 ;
  assign y11946 = n764 ;
  assign y11947 = n16423 ;
  assign y11948 = n16424 ;
  assign y11949 = n16427 ;
  assign y11950 = ~1'b0 ;
  assign y11951 = ~1'b0 ;
  assign y11952 = ~n16428 ;
  assign y11953 = ~1'b0 ;
  assign y11954 = n16429 ;
  assign y11955 = n1070 ;
  assign y11956 = ~n16433 ;
  assign y11957 = ~n16442 ;
  assign y11958 = n16455 ;
  assign y11959 = n10551 ;
  assign y11960 = ~n16458 ;
  assign y11961 = ~1'b0 ;
  assign y11962 = 1'b0 ;
  assign y11963 = ~1'b0 ;
  assign y11964 = ~n16459 ;
  assign y11965 = n16460 ;
  assign y11966 = ~n16461 ;
  assign y11967 = n16462 ;
  assign y11968 = ~n16468 ;
  assign y11969 = ~1'b0 ;
  assign y11970 = ~n5994 ;
  assign y11971 = ~1'b0 ;
  assign y11972 = ~n16469 ;
  assign y11973 = n16470 ;
  assign y11974 = ~n16472 ;
  assign y11975 = ~n16473 ;
  assign y11976 = ~1'b0 ;
  assign y11977 = ~n16475 ;
  assign y11978 = n16478 ;
  assign y11979 = n16482 ;
  assign y11980 = ~n16485 ;
  assign y11981 = ~n16486 ;
  assign y11982 = ~n16487 ;
  assign y11983 = ~n16489 ;
  assign y11984 = ~1'b0 ;
  assign y11985 = ~1'b0 ;
  assign y11986 = n16490 ;
  assign y11987 = n16492 ;
  assign y11988 = n16500 ;
  assign y11989 = ~n16501 ;
  assign y11990 = ~1'b0 ;
  assign y11991 = ~1'b0 ;
  assign y11992 = ~n16502 ;
  assign y11993 = ~1'b0 ;
  assign y11994 = ~n16505 ;
  assign y11995 = ~1'b0 ;
  assign y11996 = ~1'b0 ;
  assign y11997 = ~1'b0 ;
  assign y11998 = ~1'b0 ;
  assign y11999 = n16506 ;
  assign y12000 = ~1'b0 ;
  assign y12001 = ~1'b0 ;
  assign y12002 = ~n16511 ;
  assign y12003 = ~n16512 ;
  assign y12004 = ~n16515 ;
  assign y12005 = n16516 ;
  assign y12006 = ~n6721 ;
  assign y12007 = ~n16518 ;
  assign y12008 = ~1'b0 ;
  assign y12009 = ~1'b0 ;
  assign y12010 = 1'b0 ;
  assign y12011 = ~n16519 ;
  assign y12012 = ~n16525 ;
  assign y12013 = ~n16529 ;
  assign y12014 = ~n16535 ;
  assign y12015 = ~1'b0 ;
  assign y12016 = ~n16539 ;
  assign y12017 = ~n7868 ;
  assign y12018 = ~1'b0 ;
  assign y12019 = ~1'b0 ;
  assign y12020 = ~1'b0 ;
  assign y12021 = ~n16541 ;
  assign y12022 = ~n16543 ;
  assign y12023 = ~n16544 ;
  assign y12024 = ~n16550 ;
  assign y12025 = ~1'b0 ;
  assign y12026 = ~1'b0 ;
  assign y12027 = ~1'b0 ;
  assign y12028 = ~1'b0 ;
  assign y12029 = n16552 ;
  assign y12030 = ~n16554 ;
  assign y12031 = ~n16556 ;
  assign y12032 = 1'b0 ;
  assign y12033 = ~1'b0 ;
  assign y12034 = ~1'b0 ;
  assign y12035 = ~n16558 ;
  assign y12036 = n16561 ;
  assign y12037 = n10965 ;
  assign y12038 = ~n16565 ;
  assign y12039 = n16566 ;
  assign y12040 = ~1'b0 ;
  assign y12041 = n16568 ;
  assign y12042 = ~n1437 ;
  assign y12043 = n16572 ;
  assign y12044 = ~1'b0 ;
  assign y12045 = ~n16575 ;
  assign y12046 = ~n1786 ;
  assign y12047 = ~1'b0 ;
  assign y12048 = ~1'b0 ;
  assign y12049 = n5528 ;
  assign y12050 = ~n16579 ;
  assign y12051 = ~1'b0 ;
  assign y12052 = n16580 ;
  assign y12053 = n16582 ;
  assign y12054 = ~n16584 ;
  assign y12055 = ~1'b0 ;
  assign y12056 = n16585 ;
  assign y12057 = ~1'b0 ;
  assign y12058 = ~n16586 ;
  assign y12059 = n16588 ;
  assign y12060 = ~1'b0 ;
  assign y12061 = n16591 ;
  assign y12062 = ~n16596 ;
  assign y12063 = ~n16606 ;
  assign y12064 = ~n16610 ;
  assign y12065 = ~1'b0 ;
  assign y12066 = n16611 ;
  assign y12067 = n16612 ;
  assign y12068 = ~1'b0 ;
  assign y12069 = ~1'b0 ;
  assign y12070 = ~n5284 ;
  assign y12071 = n16613 ;
  assign y12072 = n16615 ;
  assign y12073 = ~1'b0 ;
  assign y12074 = ~n16617 ;
  assign y12075 = n16621 ;
  assign y12076 = ~1'b0 ;
  assign y12077 = 1'b0 ;
  assign y12078 = ~1'b0 ;
  assign y12079 = ~1'b0 ;
  assign y12080 = ~n16627 ;
  assign y12081 = ~1'b0 ;
  assign y12082 = n16630 ;
  assign y12083 = ~n4000 ;
  assign y12084 = n16631 ;
  assign y12085 = ~1'b0 ;
  assign y12086 = ~1'b0 ;
  assign y12087 = n16632 ;
  assign y12088 = n16633 ;
  assign y12089 = n16634 ;
  assign y12090 = ~n16635 ;
  assign y12091 = ~n16638 ;
  assign y12092 = ~n16639 ;
  assign y12093 = n16640 ;
  assign y12094 = n16641 ;
  assign y12095 = n2456 ;
  assign y12096 = ~1'b0 ;
  assign y12097 = ~1'b0 ;
  assign y12098 = ~n16646 ;
  assign y12099 = ~1'b0 ;
  assign y12100 = ~n16648 ;
  assign y12101 = ~1'b0 ;
  assign y12102 = ~1'b0 ;
  assign y12103 = n16650 ;
  assign y12104 = ~n16655 ;
  assign y12105 = ~1'b0 ;
  assign y12106 = n16659 ;
  assign y12107 = ~n16661 ;
  assign y12108 = ~1'b0 ;
  assign y12109 = ~n16490 ;
  assign y12110 = n16663 ;
  assign y12111 = x9 ;
  assign y12112 = ~1'b0 ;
  assign y12113 = n16666 ;
  assign y12114 = ~n16670 ;
  assign y12115 = ~n16672 ;
  assign y12116 = ~1'b0 ;
  assign y12117 = 1'b0 ;
  assign y12118 = ~1'b0 ;
  assign y12119 = ~1'b0 ;
  assign y12120 = ~1'b0 ;
  assign y12121 = ~1'b0 ;
  assign y12122 = n16674 ;
  assign y12123 = ~1'b0 ;
  assign y12124 = ~1'b0 ;
  assign y12125 = ~n16675 ;
  assign y12126 = ~n16680 ;
  assign y12127 = ~1'b0 ;
  assign y12128 = ~n16682 ;
  assign y12129 = n16684 ;
  assign y12130 = ~1'b0 ;
  assign y12131 = n16687 ;
  assign y12132 = ~n7551 ;
  assign y12133 = ~n8283 ;
  assign y12134 = n16689 ;
  assign y12135 = ~1'b0 ;
  assign y12136 = ~n16695 ;
  assign y12137 = ~1'b0 ;
  assign y12138 = ~n16699 ;
  assign y12139 = ~1'b0 ;
  assign y12140 = ~n7394 ;
  assign y12141 = ~1'b0 ;
  assign y12142 = ~n16700 ;
  assign y12143 = n137 ;
  assign y12144 = n16705 ;
  assign y12145 = ~n1404 ;
  assign y12146 = ~1'b0 ;
  assign y12147 = ~n1212 ;
  assign y12148 = n6477 ;
  assign y12149 = ~n16708 ;
  assign y12150 = n16710 ;
  assign y12151 = ~1'b0 ;
  assign y12152 = ~1'b0 ;
  assign y12153 = n16712 ;
  assign y12154 = ~n11044 ;
  assign y12155 = ~1'b0 ;
  assign y12156 = ~n16713 ;
  assign y12157 = ~1'b0 ;
  assign y12158 = ~1'b0 ;
  assign y12159 = ~1'b0 ;
  assign y12160 = n16716 ;
  assign y12161 = ~1'b0 ;
  assign y12162 = n16721 ;
  assign y12163 = n16726 ;
  assign y12164 = n16729 ;
  assign y12165 = ~n16735 ;
  assign y12166 = n16736 ;
  assign y12167 = n16739 ;
  assign y12168 = n16740 ;
  assign y12169 = ~n16741 ;
  assign y12170 = ~1'b0 ;
  assign y12171 = ~n16744 ;
  assign y12172 = ~n16748 ;
  assign y12173 = ~n16754 ;
  assign y12174 = ~1'b0 ;
  assign y12175 = ~1'b0 ;
  assign y12176 = n8106 ;
  assign y12177 = ~1'b0 ;
  assign y12178 = n16757 ;
  assign y12179 = ~n15021 ;
  assign y12180 = n10759 ;
  assign y12181 = ~n6062 ;
  assign y12182 = n16758 ;
  assign y12183 = ~1'b0 ;
  assign y12184 = ~1'b0 ;
  assign y12185 = ~n16760 ;
  assign y12186 = ~1'b0 ;
  assign y12187 = ~n16765 ;
  assign y12188 = n2667 ;
  assign y12189 = ~n2120 ;
  assign y12190 = n16767 ;
  assign y12191 = ~1'b0 ;
  assign y12192 = ~1'b0 ;
  assign y12193 = n16769 ;
  assign y12194 = ~n16774 ;
  assign y12195 = n16775 ;
  assign y12196 = ~n16780 ;
  assign y12197 = ~n16784 ;
  assign y12198 = n16787 ;
  assign y12199 = ~1'b0 ;
  assign y12200 = ~1'b0 ;
  assign y12201 = ~n16790 ;
  assign y12202 = ~n16791 ;
  assign y12203 = ~n16794 ;
  assign y12204 = ~1'b0 ;
  assign y12205 = n16796 ;
  assign y12206 = n3429 ;
  assign y12207 = ~n16799 ;
  assign y12208 = n16804 ;
  assign y12209 = ~n16812 ;
  assign y12210 = ~1'b0 ;
  assign y12211 = ~n16816 ;
  assign y12212 = n16818 ;
  assign y12213 = ~1'b0 ;
  assign y12214 = ~n16819 ;
  assign y12215 = ~1'b0 ;
  assign y12216 = ~n16821 ;
  assign y12217 = ~n16824 ;
  assign y12218 = ~1'b0 ;
  assign y12219 = ~n16825 ;
  assign y12220 = n16831 ;
  assign y12221 = ~1'b0 ;
  assign y12222 = ~n16832 ;
  assign y12223 = n16833 ;
  assign y12224 = ~1'b0 ;
  assign y12225 = n16837 ;
  assign y12226 = ~n4286 ;
  assign y12227 = ~1'b0 ;
  assign y12228 = n16843 ;
  assign y12229 = ~1'b0 ;
  assign y12230 = ~1'b0 ;
  assign y12231 = ~1'b0 ;
  assign y12232 = ~1'b0 ;
  assign y12233 = ~1'b0 ;
  assign y12234 = ~n16845 ;
  assign y12235 = n2268 ;
  assign y12236 = ~n16847 ;
  assign y12237 = ~n16850 ;
  assign y12238 = ~n16851 ;
  assign y12239 = ~1'b0 ;
  assign y12240 = n16852 ;
  assign y12241 = ~1'b0 ;
  assign y12242 = ~1'b0 ;
  assign y12243 = ~1'b0 ;
  assign y12244 = ~1'b0 ;
  assign y12245 = n16853 ;
  assign y12246 = ~n16858 ;
  assign y12247 = n4120 ;
  assign y12248 = n367 ;
  assign y12249 = ~1'b0 ;
  assign y12250 = ~n12028 ;
  assign y12251 = ~n16881 ;
  assign y12252 = ~n16884 ;
  assign y12253 = ~1'b0 ;
  assign y12254 = ~n16900 ;
  assign y12255 = n16903 ;
  assign y12256 = ~1'b0 ;
  assign y12257 = ~1'b0 ;
  assign y12258 = n16905 ;
  assign y12259 = ~n16908 ;
  assign y12260 = n16909 ;
  assign y12261 = n16913 ;
  assign y12262 = ~1'b0 ;
  assign y12263 = n16914 ;
  assign y12264 = ~1'b0 ;
  assign y12265 = n16916 ;
  assign y12266 = ~n16918 ;
  assign y12267 = ~1'b0 ;
  assign y12268 = n16919 ;
  assign y12269 = ~1'b0 ;
  assign y12270 = n16922 ;
  assign y12271 = n16925 ;
  assign y12272 = ~1'b0 ;
  assign y12273 = ~n16928 ;
  assign y12274 = ~1'b0 ;
  assign y12275 = ~1'b0 ;
  assign y12276 = n16930 ;
  assign y12277 = ~n16932 ;
  assign y12278 = ~n16938 ;
  assign y12279 = ~n16940 ;
  assign y12280 = ~n16942 ;
  assign y12281 = ~n16945 ;
  assign y12282 = ~1'b0 ;
  assign y12283 = ~1'b0 ;
  assign y12284 = n16946 ;
  assign y12285 = ~1'b0 ;
  assign y12286 = ~n16952 ;
  assign y12287 = ~1'b0 ;
  assign y12288 = ~1'b0 ;
  assign y12289 = ~n16960 ;
  assign y12290 = ~n16963 ;
  assign y12291 = ~1'b0 ;
  assign y12292 = ~1'b0 ;
  assign y12293 = ~1'b0 ;
  assign y12294 = ~n2767 ;
  assign y12295 = n16965 ;
  assign y12296 = ~1'b0 ;
  assign y12297 = n16966 ;
  assign y12298 = ~1'b0 ;
  assign y12299 = ~1'b0 ;
  assign y12300 = ~1'b0 ;
  assign y12301 = n16120 ;
  assign y12302 = n16967 ;
  assign y12303 = n16971 ;
  assign y12304 = ~1'b0 ;
  assign y12305 = ~n7520 ;
  assign y12306 = ~n16974 ;
  assign y12307 = ~n16977 ;
  assign y12308 = n16982 ;
  assign y12309 = n16989 ;
  assign y12310 = ~n16993 ;
  assign y12311 = ~n17006 ;
  assign y12312 = ~1'b0 ;
  assign y12313 = ~n17013 ;
  assign y12314 = ~n7197 ;
  assign y12315 = 1'b0 ;
  assign y12316 = n17017 ;
  assign y12317 = n17018 ;
  assign y12318 = ~1'b0 ;
  assign y12319 = n17019 ;
  assign y12320 = ~1'b0 ;
  assign y12321 = ~n17025 ;
  assign y12322 = ~1'b0 ;
  assign y12323 = ~n17026 ;
  assign y12324 = n17033 ;
  assign y12325 = n17037 ;
  assign y12326 = ~1'b0 ;
  assign y12327 = ~1'b0 ;
  assign y12328 = ~n17040 ;
  assign y12329 = n17048 ;
  assign y12330 = ~1'b0 ;
  assign y12331 = 1'b0 ;
  assign y12332 = n17053 ;
  assign y12333 = ~1'b0 ;
  assign y12334 = ~1'b0 ;
  assign y12335 = ~1'b0 ;
  assign y12336 = ~1'b0 ;
  assign y12337 = ~n17055 ;
  assign y12338 = ~n17056 ;
  assign y12339 = n17059 ;
  assign y12340 = ~1'b0 ;
  assign y12341 = ~1'b0 ;
  assign y12342 = n17060 ;
  assign y12343 = n17063 ;
  assign y12344 = ~n17064 ;
  assign y12345 = ~n4422 ;
  assign y12346 = ~n17065 ;
  assign y12347 = ~1'b0 ;
  assign y12348 = ~1'b0 ;
  assign y12349 = ~1'b0 ;
  assign y12350 = n3674 ;
  assign y12351 = n17066 ;
  assign y12352 = ~n13481 ;
  assign y12353 = ~n17068 ;
  assign y12354 = n17069 ;
  assign y12355 = ~n17070 ;
  assign y12356 = ~1'b0 ;
  assign y12357 = ~n17071 ;
  assign y12358 = n17073 ;
  assign y12359 = n17074 ;
  assign y12360 = ~1'b0 ;
  assign y12361 = n17075 ;
  assign y12362 = ~n17085 ;
  assign y12363 = ~1'b0 ;
  assign y12364 = ~1'b0 ;
  assign y12365 = ~n17086 ;
  assign y12366 = n17088 ;
  assign y12367 = ~1'b0 ;
  assign y12368 = 1'b0 ;
  assign y12369 = ~1'b0 ;
  assign y12370 = ~n17089 ;
  assign y12371 = n17092 ;
  assign y12372 = 1'b0 ;
  assign y12373 = ~1'b0 ;
  assign y12374 = ~1'b0 ;
  assign y12375 = n17093 ;
  assign y12376 = ~n17094 ;
  assign y12377 = n17098 ;
  assign y12378 = ~1'b0 ;
  assign y12379 = ~n17101 ;
  assign y12380 = ~n17103 ;
  assign y12381 = 1'b0 ;
  assign y12382 = n17106 ;
  assign y12383 = ~n17108 ;
  assign y12384 = n17110 ;
  assign y12385 = ~n17111 ;
  assign y12386 = n17112 ;
  assign y12387 = ~1'b0 ;
  assign y12388 = ~n17113 ;
  assign y12389 = n17115 ;
  assign y12390 = ~n16459 ;
  assign y12391 = ~1'b0 ;
  assign y12392 = ~1'b0 ;
  assign y12393 = ~1'b0 ;
  assign y12394 = n17119 ;
  assign y12395 = ~n17125 ;
  assign y12396 = ~n17128 ;
  assign y12397 = ~1'b0 ;
  assign y12398 = ~1'b0 ;
  assign y12399 = ~n17130 ;
  assign y12400 = ~n17132 ;
  assign y12401 = ~1'b0 ;
  assign y12402 = ~1'b0 ;
  assign y12403 = ~1'b0 ;
  assign y12404 = ~n17137 ;
  assign y12405 = ~n3679 ;
  assign y12406 = ~n17140 ;
  assign y12407 = ~1'b0 ;
  assign y12408 = ~n17143 ;
  assign y12409 = 1'b0 ;
  assign y12410 = ~n17146 ;
  assign y12411 = ~1'b0 ;
  assign y12412 = ~n17148 ;
  assign y12413 = ~n17150 ;
  assign y12414 = ~1'b0 ;
  assign y12415 = ~1'b0 ;
  assign y12416 = n17151 ;
  assign y12417 = ~1'b0 ;
  assign y12418 = n17153 ;
  assign y12419 = n17157 ;
  assign y12420 = n17159 ;
  assign y12421 = ~1'b0 ;
  assign y12422 = n17161 ;
  assign y12423 = ~1'b0 ;
  assign y12424 = n17163 ;
  assign y12425 = ~n17165 ;
  assign y12426 = ~1'b0 ;
  assign y12427 = ~n17166 ;
  assign y12428 = ~n17167 ;
  assign y12429 = ~n17170 ;
  assign y12430 = n17171 ;
  assign y12431 = ~1'b0 ;
  assign y12432 = ~1'b0 ;
  assign y12433 = n2339 ;
  assign y12434 = ~1'b0 ;
  assign y12435 = ~1'b0 ;
  assign y12436 = ~1'b0 ;
  assign y12437 = ~n17182 ;
  assign y12438 = n17183 ;
  assign y12439 = ~1'b0 ;
  assign y12440 = n16136 ;
  assign y12441 = ~1'b0 ;
  assign y12442 = ~1'b0 ;
  assign y12443 = ~1'b0 ;
  assign y12444 = ~n17185 ;
  assign y12445 = ~n17186 ;
  assign y12446 = ~n17193 ;
  assign y12447 = ~1'b0 ;
  assign y12448 = ~n17196 ;
  assign y12449 = ~1'b0 ;
  assign y12450 = ~n17201 ;
  assign y12451 = n17202 ;
  assign y12452 = ~1'b0 ;
  assign y12453 = n532 ;
  assign y12454 = ~n17205 ;
  assign y12455 = ~n17209 ;
  assign y12456 = n2129 ;
  assign y12457 = ~n17210 ;
  assign y12458 = 1'b0 ;
  assign y12459 = n17216 ;
  assign y12460 = ~1'b0 ;
  assign y12461 = n17218 ;
  assign y12462 = n17220 ;
  assign y12463 = n528 ;
  assign y12464 = ~n17223 ;
  assign y12465 = ~1'b0 ;
  assign y12466 = n17226 ;
  assign y12467 = ~n17227 ;
  assign y12468 = 1'b0 ;
  assign y12469 = ~1'b0 ;
  assign y12470 = ~n17228 ;
  assign y12471 = ~n17230 ;
  assign y12472 = n3848 ;
  assign y12473 = n17233 ;
  assign y12474 = ~1'b0 ;
  assign y12475 = ~1'b0 ;
  assign y12476 = ~n17241 ;
  assign y12477 = ~1'b0 ;
  assign y12478 = ~n8181 ;
  assign y12479 = ~1'b0 ;
  assign y12480 = ~n246 ;
  assign y12481 = ~1'b0 ;
  assign y12482 = ~1'b0 ;
  assign y12483 = ~1'b0 ;
  assign y12484 = ~n17243 ;
  assign y12485 = ~1'b0 ;
  assign y12486 = n17245 ;
  assign y12487 = ~1'b0 ;
  assign y12488 = ~n17247 ;
  assign y12489 = ~1'b0 ;
  assign y12490 = n13429 ;
  assign y12491 = n17249 ;
  assign y12492 = ~1'b0 ;
  assign y12493 = n17256 ;
  assign y12494 = ~1'b0 ;
  assign y12495 = ~n17258 ;
  assign y12496 = ~1'b0 ;
  assign y12497 = n17260 ;
  assign y12498 = ~1'b0 ;
  assign y12499 = ~n17261 ;
  assign y12500 = ~1'b0 ;
  assign y12501 = ~1'b0 ;
  assign y12502 = ~1'b0 ;
  assign y12503 = n17264 ;
  assign y12504 = n17265 ;
  assign y12505 = n14165 ;
  assign y12506 = n2472 ;
  assign y12507 = ~1'b0 ;
  assign y12508 = ~n6149 ;
  assign y12509 = n17266 ;
  assign y12510 = ~n17268 ;
  assign y12511 = ~n17269 ;
  assign y12512 = ~n8990 ;
  assign y12513 = ~n17277 ;
  assign y12514 = n17279 ;
  assign y12515 = n17284 ;
  assign y12516 = ~1'b0 ;
  assign y12517 = n9008 ;
  assign y12518 = ~1'b0 ;
  assign y12519 = n17285 ;
  assign y12520 = ~n11756 ;
  assign y12521 = n17286 ;
  assign y12522 = n17288 ;
  assign y12523 = ~1'b0 ;
  assign y12524 = ~1'b0 ;
  assign y12525 = ~n17290 ;
  assign y12526 = ~1'b0 ;
  assign y12527 = ~n10876 ;
  assign y12528 = ~1'b0 ;
  assign y12529 = ~n17293 ;
  assign y12530 = ~1'b0 ;
  assign y12531 = ~n17295 ;
  assign y12532 = ~n17299 ;
  assign y12533 = n17300 ;
  assign y12534 = ~n17301 ;
  assign y12535 = ~1'b0 ;
  assign y12536 = ~1'b0 ;
  assign y12537 = ~n17302 ;
  assign y12538 = n17305 ;
  assign y12539 = ~1'b0 ;
  assign y12540 = ~1'b0 ;
  assign y12541 = ~n17306 ;
  assign y12542 = ~1'b0 ;
  assign y12543 = ~n17308 ;
  assign y12544 = ~1'b0 ;
  assign y12545 = ~1'b0 ;
  assign y12546 = ~n10037 ;
  assign y12547 = ~n15790 ;
  assign y12548 = n9252 ;
  assign y12549 = ~1'b0 ;
  assign y12550 = n17313 ;
  assign y12551 = ~n17316 ;
  assign y12552 = ~1'b0 ;
  assign y12553 = ~1'b0 ;
  assign y12554 = n1627 ;
  assign y12555 = ~1'b0 ;
  assign y12556 = ~1'b0 ;
  assign y12557 = 1'b0 ;
  assign y12558 = n17317 ;
  assign y12559 = ~1'b0 ;
  assign y12560 = ~n17319 ;
  assign y12561 = n17325 ;
  assign y12562 = ~n17328 ;
  assign y12563 = ~1'b0 ;
  assign y12564 = n17329 ;
  assign y12565 = ~1'b0 ;
  assign y12566 = ~n17334 ;
  assign y12567 = ~1'b0 ;
  assign y12568 = ~1'b0 ;
  assign y12569 = 1'b0 ;
  assign y12570 = 1'b0 ;
  assign y12571 = ~n17346 ;
  assign y12572 = n17348 ;
  assign y12573 = ~n4668 ;
  assign y12574 = n1067 ;
  assign y12575 = ~1'b0 ;
  assign y12576 = ~n17351 ;
  assign y12577 = ~n17353 ;
  assign y12578 = ~n17356 ;
  assign y12579 = n17358 ;
  assign y12580 = ~n17360 ;
  assign y12581 = ~1'b0 ;
  assign y12582 = ~1'b0 ;
  assign y12583 = ~1'b0 ;
  assign y12584 = ~n17363 ;
  assign y12585 = ~1'b0 ;
  assign y12586 = ~n6442 ;
  assign y12587 = ~1'b0 ;
  assign y12588 = ~1'b0 ;
  assign y12589 = ~1'b0 ;
  assign y12590 = n17365 ;
  assign y12591 = n17366 ;
  assign y12592 = ~n17370 ;
  assign y12593 = ~n17371 ;
  assign y12594 = ~1'b0 ;
  assign y12595 = ~1'b0 ;
  assign y12596 = 1'b0 ;
  assign y12597 = ~n17372 ;
  assign y12598 = ~n17381 ;
  assign y12599 = ~n17386 ;
  assign y12600 = ~1'b0 ;
  assign y12601 = ~1'b0 ;
  assign y12602 = ~1'b0 ;
  assign y12603 = n17388 ;
  assign y12604 = ~n17389 ;
  assign y12605 = ~n17392 ;
  assign y12606 = ~n17394 ;
  assign y12607 = n8692 ;
  assign y12608 = n17395 ;
  assign y12609 = ~1'b0 ;
  assign y12610 = ~n17398 ;
  assign y12611 = ~1'b0 ;
  assign y12612 = n17431 ;
  assign y12613 = ~n17432 ;
  assign y12614 = ~n6242 ;
  assign y12615 = n17438 ;
  assign y12616 = ~1'b0 ;
  assign y12617 = ~n17441 ;
  assign y12618 = ~1'b0 ;
  assign y12619 = ~n3606 ;
  assign y12620 = ~n17444 ;
  assign y12621 = ~1'b0 ;
  assign y12622 = ~n1937 ;
  assign y12623 = n17445 ;
  assign y12624 = n17447 ;
  assign y12625 = ~1'b0 ;
  assign y12626 = ~n17449 ;
  assign y12627 = ~n17452 ;
  assign y12628 = ~1'b0 ;
  assign y12629 = ~n17461 ;
  assign y12630 = ~n812 ;
  assign y12631 = ~1'b0 ;
  assign y12632 = ~n17462 ;
  assign y12633 = ~n17464 ;
  assign y12634 = n4328 ;
  assign y12635 = n17465 ;
  assign y12636 = 1'b0 ;
  assign y12637 = n17468 ;
  assign y12638 = n13481 ;
  assign y12639 = ~n17469 ;
  assign y12640 = ~1'b0 ;
  assign y12641 = 1'b0 ;
  assign y12642 = ~1'b0 ;
  assign y12643 = ~1'b0 ;
  assign y12644 = ~n17474 ;
  assign y12645 = n17475 ;
  assign y12646 = ~1'b0 ;
  assign y12647 = n17478 ;
  assign y12648 = ~1'b0 ;
  assign y12649 = ~n17481 ;
  assign y12650 = n17482 ;
  assign y12651 = ~n17484 ;
  assign y12652 = ~1'b0 ;
  assign y12653 = ~n17486 ;
  assign y12654 = ~n17487 ;
  assign y12655 = ~n17488 ;
  assign y12656 = ~n17490 ;
  assign y12657 = ~n17493 ;
  assign y12658 = ~1'b0 ;
  assign y12659 = ~1'b0 ;
  assign y12660 = 1'b0 ;
  assign y12661 = ~n17495 ;
  assign y12662 = ~n17498 ;
  assign y12663 = n17504 ;
  assign y12664 = n17506 ;
  assign y12665 = ~1'b0 ;
  assign y12666 = n17509 ;
  assign y12667 = ~1'b0 ;
  assign y12668 = ~1'b0 ;
  assign y12669 = ~n17514 ;
  assign y12670 = ~n17516 ;
  assign y12671 = ~n6462 ;
  assign y12672 = ~n17517 ;
  assign y12673 = ~1'b0 ;
  assign y12674 = ~1'b0 ;
  assign y12675 = n17524 ;
  assign y12676 = 1'b0 ;
  assign y12677 = n17528 ;
  assign y12678 = ~1'b0 ;
  assign y12679 = n17530 ;
  assign y12680 = ~n17533 ;
  assign y12681 = ~n17534 ;
  assign y12682 = 1'b0 ;
  assign y12683 = 1'b0 ;
  assign y12684 = n17538 ;
  assign y12685 = n3418 ;
  assign y12686 = n17541 ;
  assign y12687 = ~n17547 ;
  assign y12688 = ~1'b0 ;
  assign y12689 = n17548 ;
  assign y12690 = n17549 ;
  assign y12691 = ~n17550 ;
  assign y12692 = ~n17551 ;
  assign y12693 = ~n17553 ;
  assign y12694 = ~1'b0 ;
  assign y12695 = ~1'b0 ;
  assign y12696 = n17557 ;
  assign y12697 = n3873 ;
  assign y12698 = ~n17558 ;
  assign y12699 = ~1'b0 ;
  assign y12700 = n17561 ;
  assign y12701 = n17564 ;
  assign y12702 = ~n17565 ;
  assign y12703 = ~1'b0 ;
  assign y12704 = ~n17567 ;
  assign y12705 = n17568 ;
  assign y12706 = ~n16840 ;
  assign y12707 = n17571 ;
  assign y12708 = ~n17573 ;
  assign y12709 = ~1'b0 ;
  assign y12710 = ~1'b0 ;
  assign y12711 = ~n17574 ;
  assign y12712 = ~n17579 ;
  assign y12713 = ~n7644 ;
  assign y12714 = n17584 ;
  assign y12715 = 1'b0 ;
  assign y12716 = n17586 ;
  assign y12717 = ~n17588 ;
  assign y12718 = ~1'b0 ;
  assign y12719 = n17589 ;
  assign y12720 = n10987 ;
  assign y12721 = n17591 ;
  assign y12722 = n17592 ;
  assign y12723 = ~n17596 ;
  assign y12724 = n17598 ;
  assign y12725 = ~1'b0 ;
  assign y12726 = n17599 ;
  assign y12727 = ~n17600 ;
  assign y12728 = ~1'b0 ;
  assign y12729 = ~1'b0 ;
  assign y12730 = n17601 ;
  assign y12731 = ~n17605 ;
  assign y12732 = n6834 ;
  assign y12733 = ~1'b0 ;
  assign y12734 = ~n17608 ;
  assign y12735 = n17610 ;
  assign y12736 = ~1'b0 ;
  assign y12737 = ~1'b0 ;
  assign y12738 = ~n942 ;
  assign y12739 = ~n17612 ;
  assign y12740 = ~1'b0 ;
  assign y12741 = n17613 ;
  assign y12742 = ~1'b0 ;
  assign y12743 = ~n17615 ;
  assign y12744 = ~n17617 ;
  assign y12745 = ~n17620 ;
  assign y12746 = ~1'b0 ;
  assign y12747 = ~n17621 ;
  assign y12748 = n17624 ;
  assign y12749 = ~1'b0 ;
  assign y12750 = ~1'b0 ;
  assign y12751 = ~1'b0 ;
  assign y12752 = ~1'b0 ;
  assign y12753 = ~n17625 ;
  assign y12754 = ~1'b0 ;
  assign y12755 = ~1'b0 ;
  assign y12756 = ~1'b0 ;
  assign y12757 = ~n17628 ;
  assign y12758 = n17634 ;
  assign y12759 = 1'b0 ;
  assign y12760 = ~1'b0 ;
  assign y12761 = ~n17636 ;
  assign y12762 = ~n1722 ;
  assign y12763 = n17638 ;
  assign y12764 = ~n17639 ;
  assign y12765 = ~n17640 ;
  assign y12766 = ~1'b0 ;
  assign y12767 = n5218 ;
  assign y12768 = n17642 ;
  assign y12769 = ~n17643 ;
  assign y12770 = 1'b0 ;
  assign y12771 = n17650 ;
  assign y12772 = ~1'b0 ;
  assign y12773 = ~n17651 ;
  assign y12774 = ~n17652 ;
  assign y12775 = ~n17653 ;
  assign y12776 = ~1'b0 ;
  assign y12777 = n5254 ;
  assign y12778 = n17655 ;
  assign y12779 = ~1'b0 ;
  assign y12780 = ~1'b0 ;
  assign y12781 = ~1'b0 ;
  assign y12782 = ~n10174 ;
  assign y12783 = ~1'b0 ;
  assign y12784 = 1'b0 ;
  assign y12785 = ~1'b0 ;
  assign y12786 = ~1'b0 ;
  assign y12787 = 1'b0 ;
  assign y12788 = ~n17657 ;
  assign y12789 = n6133 ;
  assign y12790 = ~1'b0 ;
  assign y12791 = ~n17665 ;
  assign y12792 = n17669 ;
  assign y12793 = ~1'b0 ;
  assign y12794 = n17670 ;
  assign y12795 = n2751 ;
  assign y12796 = n17671 ;
  assign y12797 = n17674 ;
  assign y12798 = ~1'b0 ;
  assign y12799 = ~1'b0 ;
  assign y12800 = n17675 ;
  assign y12801 = n17678 ;
  assign y12802 = ~1'b0 ;
  assign y12803 = ~1'b0 ;
  assign y12804 = ~1'b0 ;
  assign y12805 = n17680 ;
  assign y12806 = ~n17682 ;
  assign y12807 = ~1'b0 ;
  assign y12808 = n17687 ;
  assign y12809 = n17049 ;
  assign y12810 = ~n12457 ;
  assign y12811 = ~1'b0 ;
  assign y12812 = ~1'b0 ;
  assign y12813 = ~1'b0 ;
  assign y12814 = ~n17688 ;
  assign y12815 = n17691 ;
  assign y12816 = ~1'b0 ;
  assign y12817 = ~n17692 ;
  assign y12818 = ~n8069 ;
  assign y12819 = n17695 ;
  assign y12820 = ~n17701 ;
  assign y12821 = ~1'b0 ;
  assign y12822 = ~n17702 ;
  assign y12823 = ~1'b0 ;
  assign y12824 = ~n17703 ;
  assign y12825 = n17704 ;
  assign y12826 = ~1'b0 ;
  assign y12827 = n13083 ;
  assign y12828 = n17711 ;
  assign y12829 = 1'b0 ;
  assign y12830 = n17713 ;
  assign y12831 = ~1'b0 ;
  assign y12832 = n17717 ;
  assign y12833 = n17728 ;
  assign y12834 = n17734 ;
  assign y12835 = ~1'b0 ;
  assign y12836 = ~1'b0 ;
  assign y12837 = ~1'b0 ;
  assign y12838 = ~1'b0 ;
  assign y12839 = ~n4544 ;
  assign y12840 = ~1'b0 ;
  assign y12841 = ~1'b0 ;
  assign y12842 = ~1'b0 ;
  assign y12843 = 1'b0 ;
  assign y12844 = n13432 ;
  assign y12845 = ~n17736 ;
  assign y12846 = 1'b0 ;
  assign y12847 = ~n17742 ;
  assign y12848 = n17744 ;
  assign y12849 = n17746 ;
  assign y12850 = ~1'b0 ;
  assign y12851 = ~1'b0 ;
  assign y12852 = ~n17748 ;
  assign y12853 = 1'b0 ;
  assign y12854 = n56 ;
  assign y12855 = 1'b0 ;
  assign y12856 = ~1'b0 ;
  assign y12857 = ~n17754 ;
  assign y12858 = ~n17758 ;
  assign y12859 = n17759 ;
  assign y12860 = ~n1058 ;
  assign y12861 = ~n612 ;
  assign y12862 = ~n852 ;
  assign y12863 = n17760 ;
  assign y12864 = ~1'b0 ;
  assign y12865 = ~n17761 ;
  assign y12866 = n17762 ;
  assign y12867 = 1'b0 ;
  assign y12868 = ~n17764 ;
  assign y12869 = n17765 ;
  assign y12870 = n17766 ;
  assign y12871 = n17771 ;
  assign y12872 = ~1'b0 ;
  assign y12873 = ~1'b0 ;
  assign y12874 = ~n17772 ;
  assign y12875 = ~1'b0 ;
  assign y12876 = n17779 ;
  assign y12877 = ~n2157 ;
  assign y12878 = n12730 ;
  assign y12879 = ~1'b0 ;
  assign y12880 = ~n17780 ;
  assign y12881 = ~1'b0 ;
  assign y12882 = ~n17781 ;
  assign y12883 = ~1'b0 ;
  assign y12884 = ~1'b0 ;
  assign y12885 = ~n17790 ;
  assign y12886 = ~n17794 ;
  assign y12887 = n4799 ;
  assign y12888 = ~n2547 ;
  assign y12889 = ~1'b0 ;
  assign y12890 = ~n17796 ;
  assign y12891 = ~1'b0 ;
  assign y12892 = ~n17800 ;
  assign y12893 = n17802 ;
  assign y12894 = ~n17804 ;
  assign y12895 = ~n324 ;
  assign y12896 = ~n17806 ;
  assign y12897 = ~n17807 ;
  assign y12898 = ~1'b0 ;
  assign y12899 = ~n17809 ;
  assign y12900 = ~n17812 ;
  assign y12901 = ~1'b0 ;
  assign y12902 = ~n17813 ;
  assign y12903 = ~1'b0 ;
  assign y12904 = 1'b0 ;
  assign y12905 = 1'b0 ;
  assign y12906 = ~n17816 ;
  assign y12907 = ~1'b0 ;
  assign y12908 = n17817 ;
  assign y12909 = n7160 ;
  assign y12910 = ~1'b0 ;
  assign y12911 = n17818 ;
  assign y12912 = n17821 ;
  assign y12913 = n17827 ;
  assign y12914 = ~n17833 ;
  assign y12915 = ~1'b0 ;
  assign y12916 = ~n17835 ;
  assign y12917 = ~1'b0 ;
  assign y12918 = ~n17837 ;
  assign y12919 = ~n17838 ;
  assign y12920 = n17839 ;
  assign y12921 = ~1'b0 ;
  assign y12922 = ~1'b0 ;
  assign y12923 = ~1'b0 ;
  assign y12924 = n17841 ;
  assign y12925 = ~1'b0 ;
  assign y12926 = n5530 ;
  assign y12927 = n17844 ;
  assign y12928 = ~n8292 ;
  assign y12929 = ~n1469 ;
  assign y12930 = 1'b0 ;
  assign y12931 = ~1'b0 ;
  assign y12932 = n17846 ;
  assign y12933 = ~1'b0 ;
  assign y12934 = ~n17853 ;
  assign y12935 = ~n8295 ;
  assign y12936 = ~n17854 ;
  assign y12937 = ~n17856 ;
  assign y12938 = n9963 ;
  assign y12939 = ~n4449 ;
  assign y12940 = n12073 ;
  assign y12941 = n17857 ;
  assign y12942 = n17859 ;
  assign y12943 = ~n17864 ;
  assign y12944 = ~1'b0 ;
  assign y12945 = ~n17866 ;
  assign y12946 = ~1'b0 ;
  assign y12947 = n17867 ;
  assign y12948 = ~n17868 ;
  assign y12949 = ~1'b0 ;
  assign y12950 = n17875 ;
  assign y12951 = n17877 ;
  assign y12952 = ~n17881 ;
  assign y12953 = ~n17884 ;
  assign y12954 = ~1'b0 ;
  assign y12955 = n17885 ;
  assign y12956 = n1854 ;
  assign y12957 = n17887 ;
  assign y12958 = ~1'b0 ;
  assign y12959 = ~n17890 ;
  assign y12960 = 1'b0 ;
  assign y12961 = ~n16660 ;
  assign y12962 = n16225 ;
  assign y12963 = ~n17895 ;
  assign y12964 = ~n17896 ;
  assign y12965 = 1'b0 ;
  assign y12966 = ~1'b0 ;
  assign y12967 = ~1'b0 ;
  assign y12968 = ~n17897 ;
  assign y12969 = ~1'b0 ;
  assign y12970 = ~1'b0 ;
  assign y12971 = n17899 ;
  assign y12972 = n17900 ;
  assign y12973 = ~1'b0 ;
  assign y12974 = ~1'b0 ;
  assign y12975 = ~1'b0 ;
  assign y12976 = n15875 ;
  assign y12977 = ~n17901 ;
  assign y12978 = ~1'b0 ;
  assign y12979 = n17907 ;
  assign y12980 = n17911 ;
  assign y12981 = n17912 ;
  assign y12982 = 1'b0 ;
  assign y12983 = n17918 ;
  assign y12984 = n17926 ;
  assign y12985 = ~1'b0 ;
  assign y12986 = ~n17931 ;
  assign y12987 = ~1'b0 ;
  assign y12988 = ~1'b0 ;
  assign y12989 = ~1'b0 ;
  assign y12990 = n17934 ;
  assign y12991 = n17936 ;
  assign y12992 = n17939 ;
  assign y12993 = n17940 ;
  assign y12994 = ~n17942 ;
  assign y12995 = n17943 ;
  assign y12996 = ~n17946 ;
  assign y12997 = ~n17947 ;
  assign y12998 = ~1'b0 ;
  assign y12999 = ~1'b0 ;
  assign y13000 = ~n17951 ;
  assign y13001 = ~1'b0 ;
  assign y13002 = ~1'b0 ;
  assign y13003 = ~1'b0 ;
  assign y13004 = ~n17953 ;
  assign y13005 = ~n17956 ;
  assign y13006 = n11308 ;
  assign y13007 = ~n17957 ;
  assign y13008 = ~n17959 ;
  assign y13009 = n17963 ;
  assign y13010 = ~1'b0 ;
  assign y13011 = ~1'b0 ;
  assign y13012 = ~1'b0 ;
  assign y13013 = n17964 ;
  assign y13014 = n17965 ;
  assign y13015 = ~n17974 ;
  assign y13016 = n17976 ;
  assign y13017 = ~n17986 ;
  assign y13018 = ~1'b0 ;
  assign y13019 = n17987 ;
  assign y13020 = n17989 ;
  assign y13021 = ~1'b0 ;
  assign y13022 = ~1'b0 ;
  assign y13023 = n17992 ;
  assign y13024 = ~n17993 ;
  assign y13025 = n17996 ;
  assign y13026 = ~1'b0 ;
  assign y13027 = ~1'b0 ;
  assign y13028 = ~n17998 ;
  assign y13029 = ~1'b0 ;
  assign y13030 = n18001 ;
  assign y13031 = ~1'b0 ;
  assign y13032 = ~n18003 ;
  assign y13033 = ~1'b0 ;
  assign y13034 = ~n960 ;
  assign y13035 = n18004 ;
  assign y13036 = ~1'b0 ;
  assign y13037 = ~n16713 ;
  assign y13038 = ~n1851 ;
  assign y13039 = ~n18005 ;
  assign y13040 = ~n18010 ;
  assign y13041 = ~1'b0 ;
  assign y13042 = n18013 ;
  assign y13043 = ~n17449 ;
  assign y13044 = ~1'b0 ;
  assign y13045 = ~1'b0 ;
  assign y13046 = n18019 ;
  assign y13047 = ~1'b0 ;
  assign y13048 = ~n7818 ;
  assign y13049 = n3402 ;
  assign y13050 = n18021 ;
  assign y13051 = ~1'b0 ;
  assign y13052 = ~n18024 ;
  assign y13053 = ~1'b0 ;
  assign y13054 = ~n18025 ;
  assign y13055 = ~n104 ;
  assign y13056 = ~n18028 ;
  assign y13057 = ~n16483 ;
  assign y13058 = ~1'b0 ;
  assign y13059 = ~1'b0 ;
  assign y13060 = n8183 ;
  assign y13061 = ~1'b0 ;
  assign y13062 = n18030 ;
  assign y13063 = ~1'b0 ;
  assign y13064 = ~1'b0 ;
  assign y13065 = ~n18031 ;
  assign y13066 = ~n18032 ;
  assign y13067 = ~1'b0 ;
  assign y13068 = ~n18033 ;
  assign y13069 = n18034 ;
  assign y13070 = ~n18039 ;
  assign y13071 = n18043 ;
  assign y13072 = ~n3576 ;
  assign y13073 = ~n18045 ;
  assign y13074 = ~1'b0 ;
  assign y13075 = ~1'b0 ;
  assign y13076 = ~1'b0 ;
  assign y13077 = ~n18047 ;
  assign y13078 = ~n18049 ;
  assign y13079 = ~n18051 ;
  assign y13080 = ~1'b0 ;
  assign y13081 = ~1'b0 ;
  assign y13082 = ~n18055 ;
  assign y13083 = ~n18061 ;
  assign y13084 = n18062 ;
  assign y13085 = ~n18069 ;
  assign y13086 = ~1'b0 ;
  assign y13087 = ~1'b0 ;
  assign y13088 = ~1'b0 ;
  assign y13089 = ~1'b0 ;
  assign y13090 = ~1'b0 ;
  assign y13091 = ~n18072 ;
  assign y13092 = n18073 ;
  assign y13093 = ~1'b0 ;
  assign y13094 = n15319 ;
  assign y13095 = ~1'b0 ;
  assign y13096 = ~1'b0 ;
  assign y13097 = ~1'b0 ;
  assign y13098 = n18074 ;
  assign y13099 = 1'b0 ;
  assign y13100 = ~1'b0 ;
  assign y13101 = ~n18081 ;
  assign y13102 = n14549 ;
  assign y13103 = ~1'b0 ;
  assign y13104 = 1'b0 ;
  assign y13105 = n5612 ;
  assign y13106 = 1'b0 ;
  assign y13107 = ~n18082 ;
  assign y13108 = ~1'b0 ;
  assign y13109 = ~1'b0 ;
  assign y13110 = ~1'b0 ;
  assign y13111 = ~1'b0 ;
  assign y13112 = ~1'b0 ;
  assign y13113 = ~1'b0 ;
  assign y13114 = ~1'b0 ;
  assign y13115 = ~1'b0 ;
  assign y13116 = n18083 ;
  assign y13117 = n18084 ;
  assign y13118 = n18086 ;
  assign y13119 = n18087 ;
  assign y13120 = n9359 ;
  assign y13121 = n18088 ;
  assign y13122 = ~n18090 ;
  assign y13123 = 1'b0 ;
  assign y13124 = n18093 ;
  assign y13125 = n18097 ;
  assign y13126 = ~1'b0 ;
  assign y13127 = n18100 ;
  assign y13128 = n18103 ;
  assign y13129 = n7439 ;
  assign y13130 = n18107 ;
  assign y13131 = n18109 ;
  assign y13132 = ~n18110 ;
  assign y13133 = ~n18112 ;
  assign y13134 = ~n18114 ;
  assign y13135 = ~n18116 ;
  assign y13136 = ~n18118 ;
  assign y13137 = ~n18123 ;
  assign y13138 = 1'b0 ;
  assign y13139 = ~n18127 ;
  assign y13140 = ~1'b0 ;
  assign y13141 = ~n18128 ;
  assign y13142 = ~n18130 ;
  assign y13143 = ~1'b0 ;
  assign y13144 = n18132 ;
  assign y13145 = 1'b0 ;
  assign y13146 = n18136 ;
  assign y13147 = ~1'b0 ;
  assign y13148 = n2910 ;
  assign y13149 = ~1'b0 ;
  assign y13150 = ~1'b0 ;
  assign y13151 = ~1'b0 ;
  assign y13152 = ~n18138 ;
  assign y13153 = n18139 ;
  assign y13154 = ~1'b0 ;
  assign y13155 = ~n18142 ;
  assign y13156 = ~n12113 ;
  assign y13157 = ~n18144 ;
  assign y13158 = n6206 ;
  assign y13159 = n15233 ;
  assign y13160 = n18145 ;
  assign y13161 = ~1'b0 ;
  assign y13162 = ~1'b0 ;
  assign y13163 = ~1'b0 ;
  assign y13164 = n18147 ;
  assign y13165 = n18150 ;
  assign y13166 = n18152 ;
  assign y13167 = ~n18154 ;
  assign y13168 = ~1'b0 ;
  assign y13169 = ~1'b0 ;
  assign y13170 = ~n18156 ;
  assign y13171 = n18159 ;
  assign y13172 = ~n18170 ;
  assign y13173 = n18173 ;
  assign y13174 = n18174 ;
  assign y13175 = ~1'b0 ;
  assign y13176 = n18175 ;
  assign y13177 = n18176 ;
  assign y13178 = ~n18178 ;
  assign y13179 = ~1'b0 ;
  assign y13180 = n18179 ;
  assign y13181 = ~n18181 ;
  assign y13182 = n18185 ;
  assign y13183 = ~1'b0 ;
  assign y13184 = ~n18188 ;
  assign y13185 = n18189 ;
  assign y13186 = ~n18190 ;
  assign y13187 = ~n18192 ;
  assign y13188 = ~n18193 ;
  assign y13189 = n9315 ;
  assign y13190 = ~1'b0 ;
  assign y13191 = ~n18200 ;
  assign y13192 = ~1'b0 ;
  assign y13193 = n18201 ;
  assign y13194 = ~1'b0 ;
  assign y13195 = ~n18203 ;
  assign y13196 = ~1'b0 ;
  assign y13197 = n18205 ;
  assign y13198 = ~1'b0 ;
  assign y13199 = ~n18211 ;
  assign y13200 = ~1'b0 ;
  assign y13201 = ~1'b0 ;
  assign y13202 = n18212 ;
  assign y13203 = ~1'b0 ;
  assign y13204 = ~1'b0 ;
  assign y13205 = n18213 ;
  assign y13206 = n18218 ;
  assign y13207 = ~1'b0 ;
  assign y13208 = ~n18219 ;
  assign y13209 = n18226 ;
  assign y13210 = ~n18227 ;
  assign y13211 = ~n18228 ;
  assign y13212 = ~1'b0 ;
  assign y13213 = n4247 ;
  assign y13214 = n18231 ;
  assign y13215 = n1326 ;
  assign y13216 = n553 ;
  assign y13217 = ~1'b0 ;
  assign y13218 = ~1'b0 ;
  assign y13219 = n18233 ;
  assign y13220 = n18237 ;
  assign y13221 = n18239 ;
  assign y13222 = ~1'b0 ;
  assign y13223 = ~n18241 ;
  assign y13224 = ~1'b0 ;
  assign y13225 = ~n18242 ;
  assign y13226 = ~n18247 ;
  assign y13227 = 1'b0 ;
  assign y13228 = ~n18248 ;
  assign y13229 = n14998 ;
  assign y13230 = ~n18250 ;
  assign y13231 = ~n18255 ;
  assign y13232 = ~1'b0 ;
  assign y13233 = ~n18258 ;
  assign y13234 = ~1'b0 ;
  assign y13235 = ~n18259 ;
  assign y13236 = ~n18261 ;
  assign y13237 = ~1'b0 ;
  assign y13238 = ~n18262 ;
  assign y13239 = ~n18266 ;
  assign y13240 = n18267 ;
  assign y13241 = ~1'b0 ;
  assign y13242 = ~1'b0 ;
  assign y13243 = ~1'b0 ;
  assign y13244 = n18268 ;
  assign y13245 = n11833 ;
  assign y13246 = n18270 ;
  assign y13247 = ~n18271 ;
  assign y13248 = ~n18272 ;
  assign y13249 = ~n18276 ;
  assign y13250 = n18288 ;
  assign y13251 = ~n18289 ;
  assign y13252 = ~n7574 ;
  assign y13253 = ~n18292 ;
  assign y13254 = n18293 ;
  assign y13255 = 1'b0 ;
  assign y13256 = n18294 ;
  assign y13257 = ~n18297 ;
  assign y13258 = ~n18299 ;
  assign y13259 = ~n18300 ;
  assign y13260 = n18302 ;
  assign y13261 = n18303 ;
  assign y13262 = ~n18304 ;
  assign y13263 = ~n18305 ;
  assign y13264 = n18307 ;
  assign y13265 = 1'b0 ;
  assign y13266 = 1'b0 ;
  assign y13267 = ~1'b0 ;
  assign y13268 = ~n18310 ;
  assign y13269 = ~n18311 ;
  assign y13270 = ~n18312 ;
  assign y13271 = ~1'b0 ;
  assign y13272 = n18316 ;
  assign y13273 = ~n18319 ;
  assign y13274 = n11802 ;
  assign y13275 = ~1'b0 ;
  assign y13276 = ~n18320 ;
  assign y13277 = ~n18322 ;
  assign y13278 = n18324 ;
  assign y13279 = ~n18325 ;
  assign y13280 = n18328 ;
  assign y13281 = ~1'b0 ;
  assign y13282 = n18330 ;
  assign y13283 = ~n18332 ;
  assign y13284 = n18334 ;
  assign y13285 = ~1'b0 ;
  assign y13286 = ~1'b0 ;
  assign y13287 = ~1'b0 ;
  assign y13288 = ~1'b0 ;
  assign y13289 = ~n18336 ;
  assign y13290 = ~1'b0 ;
  assign y13291 = ~n18337 ;
  assign y13292 = ~1'b0 ;
  assign y13293 = ~1'b0 ;
  assign y13294 = n18340 ;
  assign y13295 = n18344 ;
  assign y13296 = ~n18346 ;
  assign y13297 = ~1'b0 ;
  assign y13298 = ~n1178 ;
  assign y13299 = 1'b0 ;
  assign y13300 = 1'b0 ;
  assign y13301 = ~n5744 ;
  assign y13302 = ~n18348 ;
  assign y13303 = ~1'b0 ;
  assign y13304 = ~1'b0 ;
  assign y13305 = ~1'b0 ;
  assign y13306 = n1704 ;
  assign y13307 = ~n18350 ;
  assign y13308 = ~1'b0 ;
  assign y13309 = ~n18357 ;
  assign y13310 = ~1'b0 ;
  assign y13311 = n5205 ;
  assign y13312 = n18358 ;
  assign y13313 = ~n18359 ;
  assign y13314 = n18361 ;
  assign y13315 = n18363 ;
  assign y13316 = ~1'b0 ;
  assign y13317 = ~n18366 ;
  assign y13318 = ~n18375 ;
  assign y13319 = ~1'b0 ;
  assign y13320 = ~n4748 ;
  assign y13321 = n18378 ;
  assign y13322 = n8863 ;
  assign y13323 = ~n18380 ;
  assign y13324 = ~n9531 ;
  assign y13325 = n18381 ;
  assign y13326 = ~1'b0 ;
  assign y13327 = ~1'b0 ;
  assign y13328 = ~1'b0 ;
  assign y13329 = n18382 ;
  assign y13330 = ~n18385 ;
  assign y13331 = ~n18388 ;
  assign y13332 = ~n8596 ;
  assign y13333 = ~1'b0 ;
  assign y13334 = ~n18391 ;
  assign y13335 = ~n3217 ;
  assign y13336 = ~n18276 ;
  assign y13337 = n18392 ;
  assign y13338 = ~1'b0 ;
  assign y13339 = ~1'b0 ;
  assign y13340 = ~n18398 ;
  assign y13341 = n1463 ;
  assign y13342 = n10994 ;
  assign y13343 = n18400 ;
  assign y13344 = ~1'b0 ;
  assign y13345 = ~n18402 ;
  assign y13346 = n18407 ;
  assign y13347 = ~n18408 ;
  assign y13348 = ~1'b0 ;
  assign y13349 = ~1'b0 ;
  assign y13350 = ~n18414 ;
  assign y13351 = ~1'b0 ;
  assign y13352 = ~1'b0 ;
  assign y13353 = 1'b0 ;
  assign y13354 = ~1'b0 ;
  assign y13355 = n18415 ;
  assign y13356 = n18422 ;
  assign y13357 = ~1'b0 ;
  assign y13358 = ~1'b0 ;
  assign y13359 = n18423 ;
  assign y13360 = ~n18432 ;
  assign y13361 = n632 ;
  assign y13362 = ~1'b0 ;
  assign y13363 = ~1'b0 ;
  assign y13364 = n18433 ;
  assign y13365 = n8429 ;
  assign y13366 = ~n18445 ;
  assign y13367 = ~1'b0 ;
  assign y13368 = ~1'b0 ;
  assign y13369 = ~n18446 ;
  assign y13370 = 1'b0 ;
  assign y13371 = ~1'b0 ;
  assign y13372 = ~n18448 ;
  assign y13373 = n18451 ;
  assign y13374 = ~n18456 ;
  assign y13375 = ~n18464 ;
  assign y13376 = n18468 ;
  assign y13377 = n18469 ;
  assign y13378 = ~1'b0 ;
  assign y13379 = ~1'b0 ;
  assign y13380 = ~n18472 ;
  assign y13381 = n1961 ;
  assign y13382 = ~1'b0 ;
  assign y13383 = ~1'b0 ;
  assign y13384 = n7419 ;
  assign y13385 = ~n15942 ;
  assign y13386 = n18473 ;
  assign y13387 = n11042 ;
  assign y13388 = n18474 ;
  assign y13389 = n18476 ;
  assign y13390 = ~1'b0 ;
  assign y13391 = ~n18480 ;
  assign y13392 = ~n18483 ;
  assign y13393 = ~1'b0 ;
  assign y13394 = ~1'b0 ;
  assign y13395 = ~n18484 ;
  assign y13396 = ~n18487 ;
  assign y13397 = ~1'b0 ;
  assign y13398 = n18488 ;
  assign y13399 = ~n18492 ;
  assign y13400 = ~n18496 ;
  assign y13401 = ~n18503 ;
  assign y13402 = ~1'b0 ;
  assign y13403 = ~n1090 ;
  assign y13404 = ~1'b0 ;
  assign y13405 = n18505 ;
  assign y13406 = ~1'b0 ;
  assign y13407 = ~1'b0 ;
  assign y13408 = n18506 ;
  assign y13409 = ~n18508 ;
  assign y13410 = n3237 ;
  assign y13411 = n18509 ;
  assign y13412 = ~1'b0 ;
  assign y13413 = ~n18511 ;
  assign y13414 = ~1'b0 ;
  assign y13415 = n18515 ;
  assign y13416 = n18518 ;
  assign y13417 = n18519 ;
  assign y13418 = ~1'b0 ;
  assign y13419 = n18520 ;
  assign y13420 = ~n18521 ;
  assign y13421 = ~n18522 ;
  assign y13422 = n18526 ;
  assign y13423 = ~n18533 ;
  assign y13424 = ~1'b0 ;
  assign y13425 = n3500 ;
  assign y13426 = ~n18536 ;
  assign y13427 = n18537 ;
  assign y13428 = ~1'b0 ;
  assign y13429 = 1'b0 ;
  assign y13430 = ~n18545 ;
  assign y13431 = ~n18548 ;
  assign y13432 = ~n18554 ;
  assign y13433 = n18555 ;
  assign y13434 = ~1'b0 ;
  assign y13435 = ~n18556 ;
  assign y13436 = ~n18560 ;
  assign y13437 = n18562 ;
  assign y13438 = ~1'b0 ;
  assign y13439 = n18563 ;
  assign y13440 = n18564 ;
  assign y13441 = ~1'b0 ;
  assign y13442 = 1'b0 ;
  assign y13443 = ~1'b0 ;
  assign y13444 = ~1'b0 ;
  assign y13445 = ~n18568 ;
  assign y13446 = ~1'b0 ;
  assign y13447 = n18569 ;
  assign y13448 = n18572 ;
  assign y13449 = ~n18574 ;
  assign y13450 = ~1'b0 ;
  assign y13451 = ~1'b0 ;
  assign y13452 = n18575 ;
  assign y13453 = ~n18580 ;
  assign y13454 = n18581 ;
  assign y13455 = ~n18582 ;
  assign y13456 = n12354 ;
  assign y13457 = 1'b0 ;
  assign y13458 = ~n18583 ;
  assign y13459 = ~1'b0 ;
  assign y13460 = n18585 ;
  assign y13461 = ~1'b0 ;
  assign y13462 = ~n17057 ;
  assign y13463 = n18588 ;
  assign y13464 = ~1'b0 ;
  assign y13465 = ~n18589 ;
  assign y13466 = ~n5726 ;
  assign y13467 = ~1'b0 ;
  assign y13468 = ~1'b0 ;
  assign y13469 = 1'b0 ;
  assign y13470 = n18590 ;
  assign y13471 = ~n18593 ;
  assign y13472 = ~n18600 ;
  assign y13473 = n512 ;
  assign y13474 = ~1'b0 ;
  assign y13475 = ~1'b0 ;
  assign y13476 = ~n18601 ;
  assign y13477 = ~n18603 ;
  assign y13478 = n18605 ;
  assign y13479 = ~n18607 ;
  assign y13480 = ~1'b0 ;
  assign y13481 = ~1'b0 ;
  assign y13482 = n4485 ;
  assign y13483 = ~1'b0 ;
  assign y13484 = ~n18608 ;
  assign y13485 = ~1'b0 ;
  assign y13486 = ~1'b0 ;
  assign y13487 = ~n18614 ;
  assign y13488 = ~1'b0 ;
  assign y13489 = ~1'b0 ;
  assign y13490 = ~n18618 ;
  assign y13491 = ~1'b0 ;
  assign y13492 = n18619 ;
  assign y13493 = n18622 ;
  assign y13494 = ~1'b0 ;
  assign y13495 = ~1'b0 ;
  assign y13496 = ~n18623 ;
  assign y13497 = ~1'b0 ;
  assign y13498 = 1'b0 ;
  assign y13499 = ~1'b0 ;
  assign y13500 = ~n18626 ;
  assign y13501 = n18629 ;
  assign y13502 = ~n18632 ;
  assign y13503 = ~n18634 ;
  assign y13504 = ~n18635 ;
  assign y13505 = ~1'b0 ;
  assign y13506 = n18636 ;
  assign y13507 = ~1'b0 ;
  assign y13508 = ~1'b0 ;
  assign y13509 = ~n14422 ;
  assign y13510 = 1'b0 ;
  assign y13511 = 1'b0 ;
  assign y13512 = n18637 ;
  assign y13513 = ~n1368 ;
  assign y13514 = ~1'b0 ;
  assign y13515 = ~1'b0 ;
  assign y13516 = n18638 ;
  assign y13517 = n18641 ;
  assign y13518 = ~1'b0 ;
  assign y13519 = ~n36 ;
  assign y13520 = ~1'b0 ;
  assign y13521 = n1069 ;
  assign y13522 = n18642 ;
  assign y13523 = n18643 ;
  assign y13524 = ~n14683 ;
  assign y13525 = ~n18646 ;
  assign y13526 = ~n18648 ;
  assign y13527 = n18650 ;
  assign y13528 = ~n18651 ;
  assign y13529 = ~1'b0 ;
  assign y13530 = ~n18654 ;
  assign y13531 = ~1'b0 ;
  assign y13532 = n18662 ;
  assign y13533 = n18664 ;
  assign y13534 = n18666 ;
  assign y13535 = ~1'b0 ;
  assign y13536 = n18710 ;
  assign y13537 = ~n18712 ;
  assign y13538 = ~n310 ;
  assign y13539 = n18716 ;
  assign y13540 = ~n18717 ;
  assign y13541 = ~n18719 ;
  assign y13542 = ~n18720 ;
  assign y13543 = ~1'b0 ;
  assign y13544 = ~n18722 ;
  assign y13545 = ~1'b0 ;
  assign y13546 = ~1'b0 ;
  assign y13547 = ~1'b0 ;
  assign y13548 = ~1'b0 ;
  assign y13549 = ~1'b0 ;
  assign y13550 = ~n18727 ;
  assign y13551 = n18733 ;
  assign y13552 = n18738 ;
  assign y13553 = ~1'b0 ;
  assign y13554 = ~1'b0 ;
  assign y13555 = n4492 ;
  assign y13556 = ~1'b0 ;
  assign y13557 = n18739 ;
  assign y13558 = 1'b0 ;
  assign y13559 = ~n18740 ;
  assign y13560 = ~n18741 ;
  assign y13561 = 1'b0 ;
  assign y13562 = ~1'b0 ;
  assign y13563 = ~n12669 ;
  assign y13564 = ~1'b0 ;
  assign y13565 = ~n18749 ;
  assign y13566 = ~n3037 ;
  assign y13567 = 1'b0 ;
  assign y13568 = ~n18751 ;
  assign y13569 = n18753 ;
  assign y13570 = ~1'b0 ;
  assign y13571 = n18755 ;
  assign y13572 = ~1'b0 ;
  assign y13573 = 1'b0 ;
  assign y13574 = ~1'b0 ;
  assign y13575 = ~n18756 ;
  assign y13576 = 1'b0 ;
  assign y13577 = ~n18759 ;
  assign y13578 = n18762 ;
  assign y13579 = ~n18763 ;
  assign y13580 = ~1'b0 ;
  assign y13581 = ~1'b0 ;
  assign y13582 = ~1'b0 ;
  assign y13583 = n18766 ;
  assign y13584 = n18767 ;
  assign y13585 = n18777 ;
  assign y13586 = ~1'b0 ;
  assign y13587 = n18778 ;
  assign y13588 = ~n14804 ;
  assign y13589 = 1'b0 ;
  assign y13590 = n18783 ;
  assign y13591 = ~1'b0 ;
  assign y13592 = ~n263 ;
  assign y13593 = ~n18785 ;
  assign y13594 = ~1'b0 ;
  assign y13595 = n229 ;
  assign y13596 = ~n18786 ;
  assign y13597 = n18789 ;
  assign y13598 = ~1'b0 ;
  assign y13599 = n18790 ;
  assign y13600 = n11684 ;
  assign y13601 = ~n18791 ;
  assign y13602 = ~n18792 ;
  assign y13603 = ~n18793 ;
  assign y13604 = ~1'b0 ;
  assign y13605 = ~1'b0 ;
  assign y13606 = ~n18795 ;
  assign y13607 = ~1'b0 ;
  assign y13608 = n18798 ;
  assign y13609 = n2681 ;
  assign y13610 = ~1'b0 ;
  assign y13611 = ~n18800 ;
  assign y13612 = ~1'b0 ;
  assign y13613 = n18802 ;
  assign y13614 = n18803 ;
  assign y13615 = n18804 ;
  assign y13616 = ~n14224 ;
  assign y13617 = ~n18805 ;
  assign y13618 = ~1'b0 ;
  assign y13619 = ~1'b0 ;
  assign y13620 = ~n18808 ;
  assign y13621 = ~1'b0 ;
  assign y13622 = ~1'b0 ;
  assign y13623 = ~n18809 ;
  assign y13624 = n18814 ;
  assign y13625 = n18818 ;
  assign y13626 = n18822 ;
  assign y13627 = ~n18824 ;
  assign y13628 = n18832 ;
  assign y13629 = ~1'b0 ;
  assign y13630 = n18833 ;
  assign y13631 = ~n18838 ;
  assign y13632 = ~1'b0 ;
  assign y13633 = ~n18841 ;
  assign y13634 = n9461 ;
  assign y13635 = n18842 ;
  assign y13636 = ~1'b0 ;
  assign y13637 = ~n18843 ;
  assign y13638 = ~n18848 ;
  assign y13639 = ~1'b0 ;
  assign y13640 = ~1'b0 ;
  assign y13641 = n6001 ;
  assign y13642 = ~n10965 ;
  assign y13643 = ~n18850 ;
  assign y13644 = n18851 ;
  assign y13645 = ~1'b0 ;
  assign y13646 = n14789 ;
  assign y13647 = n18852 ;
  assign y13648 = ~n18855 ;
  assign y13649 = ~n18859 ;
  assign y13650 = 1'b0 ;
  assign y13651 = ~n18862 ;
  assign y13652 = ~n18863 ;
  assign y13653 = ~1'b0 ;
  assign y13654 = ~n18866 ;
  assign y13655 = ~1'b0 ;
  assign y13656 = ~n8665 ;
  assign y13657 = ~n2842 ;
  assign y13658 = n18867 ;
  assign y13659 = ~1'b0 ;
  assign y13660 = ~1'b0 ;
  assign y13661 = ~1'b0 ;
  assign y13662 = n18868 ;
  assign y13663 = n18871 ;
  assign y13664 = ~n18873 ;
  assign y13665 = n18880 ;
  assign y13666 = ~1'b0 ;
  assign y13667 = ~1'b0 ;
  assign y13668 = ~1'b0 ;
  assign y13669 = 1'b0 ;
  assign y13670 = n18883 ;
  assign y13671 = ~1'b0 ;
  assign y13672 = ~1'b0 ;
  assign y13673 = n18884 ;
  assign y13674 = ~n18885 ;
  assign y13675 = n1399 ;
  assign y13676 = ~n291 ;
  assign y13677 = n6194 ;
  assign y13678 = ~n18888 ;
  assign y13679 = ~n18891 ;
  assign y13680 = ~n18892 ;
  assign y13681 = n18893 ;
  assign y13682 = ~n18894 ;
  assign y13683 = ~1'b0 ;
  assign y13684 = n18899 ;
  assign y13685 = ~1'b0 ;
  assign y13686 = ~n18908 ;
  assign y13687 = ~1'b0 ;
  assign y13688 = ~n18910 ;
  assign y13689 = ~n18915 ;
  assign y13690 = ~n18918 ;
  assign y13691 = ~1'b0 ;
  assign y13692 = ~n7612 ;
  assign y13693 = ~1'b0 ;
  assign y13694 = n18919 ;
  assign y13695 = n18925 ;
  assign y13696 = ~1'b0 ;
  assign y13697 = ~1'b0 ;
  assign y13698 = n18930 ;
  assign y13699 = ~n18935 ;
  assign y13700 = n18936 ;
  assign y13701 = ~1'b0 ;
  assign y13702 = n18937 ;
  assign y13703 = n18939 ;
  assign y13704 = ~n18947 ;
  assign y13705 = ~1'b0 ;
  assign y13706 = ~1'b0 ;
  assign y13707 = ~1'b0 ;
  assign y13708 = ~1'b0 ;
  assign y13709 = ~1'b0 ;
  assign y13710 = ~n18951 ;
  assign y13711 = ~1'b0 ;
  assign y13712 = ~1'b0 ;
  assign y13713 = 1'b0 ;
  assign y13714 = n18958 ;
  assign y13715 = ~1'b0 ;
  assign y13716 = ~1'b0 ;
  assign y13717 = n11044 ;
  assign y13718 = ~n18960 ;
  assign y13719 = ~n18965 ;
  assign y13720 = n236 ;
  assign y13721 = ~n18968 ;
  assign y13722 = ~n18971 ;
  assign y13723 = ~1'b0 ;
  assign y13724 = ~n18973 ;
  assign y13725 = ~1'b0 ;
  assign y13726 = n18976 ;
  assign y13727 = n18977 ;
  assign y13728 = ~1'b0 ;
  assign y13729 = ~1'b0 ;
  assign y13730 = ~1'b0 ;
  assign y13731 = n18979 ;
  assign y13732 = ~1'b0 ;
  assign y13733 = ~n10019 ;
  assign y13734 = ~1'b0 ;
  assign y13735 = ~n18983 ;
  assign y13736 = ~n18990 ;
  assign y13737 = n4533 ;
  assign y13738 = ~1'b0 ;
  assign y13739 = ~n18996 ;
  assign y13740 = n4756 ;
  assign y13741 = n18997 ;
  assign y13742 = n19000 ;
  assign y13743 = n19003 ;
  assign y13744 = ~n19005 ;
  assign y13745 = ~1'b0 ;
  assign y13746 = ~1'b0 ;
  assign y13747 = n6133 ;
  assign y13748 = n14120 ;
  assign y13749 = ~n10718 ;
  assign y13750 = ~n19007 ;
  assign y13751 = n2680 ;
  assign y13752 = n19009 ;
  assign y13753 = ~1'b0 ;
  assign y13754 = ~1'b0 ;
  assign y13755 = n19010 ;
  assign y13756 = ~1'b0 ;
  assign y13757 = n19011 ;
  assign y13758 = ~1'b0 ;
  assign y13759 = n19012 ;
  assign y13760 = ~n19015 ;
  assign y13761 = ~n19016 ;
  assign y13762 = ~n19019 ;
  assign y13763 = ~n2209 ;
  assign y13764 = ~1'b0 ;
  assign y13765 = n19024 ;
  assign y13766 = 1'b0 ;
  assign y13767 = ~1'b0 ;
  assign y13768 = ~1'b0 ;
  assign y13769 = ~n5698 ;
  assign y13770 = ~n19025 ;
  assign y13771 = ~n19026 ;
  assign y13772 = ~n19034 ;
  assign y13773 = ~n19039 ;
  assign y13774 = ~n19040 ;
  assign y13775 = ~n19041 ;
  assign y13776 = ~n10277 ;
  assign y13777 = ~1'b0 ;
  assign y13778 = ~1'b0 ;
  assign y13779 = n19044 ;
  assign y13780 = 1'b0 ;
  assign y13781 = ~1'b0 ;
  assign y13782 = ~n19050 ;
  assign y13783 = ~1'b0 ;
  assign y13784 = ~1'b0 ;
  assign y13785 = ~n19053 ;
  assign y13786 = n19066 ;
  assign y13787 = ~1'b0 ;
  assign y13788 = ~n19069 ;
  assign y13789 = ~1'b0 ;
  assign y13790 = n19075 ;
  assign y13791 = ~1'b0 ;
  assign y13792 = 1'b0 ;
  assign y13793 = n19077 ;
  assign y13794 = ~1'b0 ;
  assign y13795 = ~1'b0 ;
  assign y13796 = 1'b0 ;
  assign y13797 = ~n19080 ;
  assign y13798 = ~1'b0 ;
  assign y13799 = n19081 ;
  assign y13800 = 1'b0 ;
  assign y13801 = n19082 ;
  assign y13802 = n19087 ;
  assign y13803 = ~1'b0 ;
  assign y13804 = ~n3311 ;
  assign y13805 = ~n19090 ;
  assign y13806 = ~1'b0 ;
  assign y13807 = n9351 ;
  assign y13808 = ~n19091 ;
  assign y13809 = ~1'b0 ;
  assign y13810 = ~n19092 ;
  assign y13811 = n1100 ;
  assign y13812 = ~n19095 ;
  assign y13813 = ~1'b0 ;
  assign y13814 = ~n19096 ;
  assign y13815 = ~n19097 ;
  assign y13816 = n19105 ;
  assign y13817 = ~1'b0 ;
  assign y13818 = ~n19109 ;
  assign y13819 = ~n19110 ;
  assign y13820 = ~1'b0 ;
  assign y13821 = ~n19111 ;
  assign y13822 = ~1'b0 ;
  assign y13823 = ~1'b0 ;
  assign y13824 = ~1'b0 ;
  assign y13825 = ~1'b0 ;
  assign y13826 = n19113 ;
  assign y13827 = 1'b0 ;
  assign y13828 = ~1'b0 ;
  assign y13829 = ~n19115 ;
  assign y13830 = n19116 ;
  assign y13831 = ~1'b0 ;
  assign y13832 = ~1'b0 ;
  assign y13833 = ~1'b0 ;
  assign y13834 = ~n18735 ;
  assign y13835 = ~n19120 ;
  assign y13836 = n19121 ;
  assign y13837 = ~n19122 ;
  assign y13838 = n19124 ;
  assign y13839 = ~1'b0 ;
  assign y13840 = n19126 ;
  assign y13841 = n6250 ;
  assign y13842 = ~n19135 ;
  assign y13843 = n19136 ;
  assign y13844 = n19137 ;
  assign y13845 = n19140 ;
  assign y13846 = ~1'b0 ;
  assign y13847 = ~1'b0 ;
  assign y13848 = n19141 ;
  assign y13849 = ~1'b0 ;
  assign y13850 = n19142 ;
  assign y13851 = ~n19143 ;
  assign y13852 = ~1'b0 ;
  assign y13853 = n19146 ;
  assign y13854 = n19149 ;
  assign y13855 = ~1'b0 ;
  assign y13856 = n19150 ;
  assign y13857 = ~1'b0 ;
  assign y13858 = ~1'b0 ;
  assign y13859 = ~n2082 ;
  assign y13860 = ~n19151 ;
  assign y13861 = 1'b0 ;
  assign y13862 = ~1'b0 ;
  assign y13863 = ~n19155 ;
  assign y13864 = n19156 ;
  assign y13865 = 1'b0 ;
  assign y13866 = ~1'b0 ;
  assign y13867 = n19158 ;
  assign y13868 = ~n19160 ;
  assign y13869 = n19161 ;
  assign y13870 = n19165 ;
  assign y13871 = ~n15482 ;
  assign y13872 = ~1'b0 ;
  assign y13873 = ~n19167 ;
  assign y13874 = ~1'b0 ;
  assign y13875 = n19169 ;
  assign y13876 = n19172 ;
  assign y13877 = ~1'b0 ;
  assign y13878 = ~1'b0 ;
  assign y13879 = n19173 ;
  assign y13880 = ~1'b0 ;
  assign y13881 = n12390 ;
  assign y13882 = 1'b0 ;
  assign y13883 = ~n19182 ;
  assign y13884 = ~1'b0 ;
  assign y13885 = n19183 ;
  assign y13886 = ~n19185 ;
  assign y13887 = ~1'b0 ;
  assign y13888 = 1'b0 ;
  assign y13889 = n19186 ;
  assign y13890 = ~n4428 ;
  assign y13891 = ~n19187 ;
  assign y13892 = ~1'b0 ;
  assign y13893 = n19193 ;
  assign y13894 = n19197 ;
  assign y13895 = n19204 ;
  assign y13896 = ~1'b0 ;
  assign y13897 = ~1'b0 ;
  assign y13898 = ~n19205 ;
  assign y13899 = ~1'b0 ;
  assign y13900 = n19207 ;
  assign y13901 = n7117 ;
  assign y13902 = n19213 ;
  assign y13903 = ~n19215 ;
  assign y13904 = ~n19217 ;
  assign y13905 = n19219 ;
  assign y13906 = ~n19223 ;
  assign y13907 = ~1'b0 ;
  assign y13908 = ~n19224 ;
  assign y13909 = 1'b0 ;
  assign y13910 = 1'b0 ;
  assign y13911 = ~1'b0 ;
  assign y13912 = ~1'b0 ;
  assign y13913 = ~n19228 ;
  assign y13914 = ~n12454 ;
  assign y13915 = n19231 ;
  assign y13916 = ~n30 ;
  assign y13917 = ~n19233 ;
  assign y13918 = n19234 ;
  assign y13919 = n19236 ;
  assign y13920 = ~1'b0 ;
  assign y13921 = n19237 ;
  assign y13922 = n19240 ;
  assign y13923 = ~n5180 ;
  assign y13924 = n19243 ;
  assign y13925 = ~1'b0 ;
  assign y13926 = ~1'b0 ;
  assign y13927 = ~1'b0 ;
  assign y13928 = n19245 ;
  assign y13929 = 1'b0 ;
  assign y13930 = ~1'b0 ;
  assign y13931 = ~n19246 ;
  assign y13932 = ~1'b0 ;
  assign y13933 = ~n19249 ;
  assign y13934 = ~1'b0 ;
  assign y13935 = n19255 ;
  assign y13936 = ~n19258 ;
  assign y13937 = 1'b0 ;
  assign y13938 = ~n19260 ;
  assign y13939 = n19261 ;
  assign y13940 = ~1'b0 ;
  assign y13941 = ~1'b0 ;
  assign y13942 = ~n19264 ;
  assign y13943 = ~n19266 ;
  assign y13944 = n19292 ;
  assign y13945 = ~n19293 ;
  assign y13946 = 1'b0 ;
  assign y13947 = ~n10194 ;
  assign y13948 = n19296 ;
  assign y13949 = n19299 ;
  assign y13950 = ~1'b0 ;
  assign y13951 = ~n19307 ;
  assign y13952 = ~n19312 ;
  assign y13953 = ~1'b0 ;
  assign y13954 = ~1'b0 ;
  assign y13955 = n19316 ;
  assign y13956 = 1'b0 ;
  assign y13957 = n19318 ;
  assign y13958 = ~n19319 ;
  assign y13959 = 1'b0 ;
  assign y13960 = ~n19325 ;
  assign y13961 = ~1'b0 ;
  assign y13962 = ~n19328 ;
  assign y13963 = ~1'b0 ;
  assign y13964 = ~1'b0 ;
  assign y13965 = n510 ;
  assign y13966 = ~1'b0 ;
  assign y13967 = ~n19329 ;
  assign y13968 = n19330 ;
  assign y13969 = n2342 ;
  assign y13970 = ~1'b0 ;
  assign y13971 = n18856 ;
  assign y13972 = ~n19332 ;
  assign y13973 = ~1'b0 ;
  assign y13974 = ~1'b0 ;
  assign y13975 = ~1'b0 ;
  assign y13976 = n19345 ;
  assign y13977 = ~n19350 ;
  assign y13978 = n16473 ;
  assign y13979 = ~1'b0 ;
  assign y13980 = ~n19354 ;
  assign y13981 = 1'b0 ;
  assign y13982 = ~n19359 ;
  assign y13983 = n19361 ;
  assign y13984 = n19365 ;
  assign y13985 = ~n297 ;
  assign y13986 = ~n19369 ;
  assign y13987 = n19370 ;
  assign y13988 = n19372 ;
  assign y13989 = ~n17263 ;
  assign y13990 = ~1'b0 ;
  assign y13991 = n15416 ;
  assign y13992 = n19374 ;
  assign y13993 = ~n19378 ;
  assign y13994 = 1'b0 ;
  assign y13995 = ~1'b0 ;
  assign y13996 = n19387 ;
  assign y13997 = ~1'b0 ;
  assign y13998 = n19389 ;
  assign y13999 = n19391 ;
  assign y14000 = 1'b0 ;
  assign y14001 = ~1'b0 ;
  assign y14002 = ~n19392 ;
  assign y14003 = n19394 ;
  assign y14004 = ~1'b0 ;
  assign y14005 = ~1'b0 ;
  assign y14006 = ~1'b0 ;
  assign y14007 = ~1'b0 ;
  assign y14008 = ~n19398 ;
  assign y14009 = n5438 ;
  assign y14010 = n19399 ;
  assign y14011 = ~1'b0 ;
  assign y14012 = ~n19400 ;
  assign y14013 = ~1'b0 ;
  assign y14014 = ~1'b0 ;
  assign y14015 = ~1'b0 ;
  assign y14016 = ~n6658 ;
  assign y14017 = ~1'b0 ;
  assign y14018 = n19401 ;
  assign y14019 = n19402 ;
  assign y14020 = ~1'b0 ;
  assign y14021 = n19403 ;
  assign y14022 = ~n19404 ;
  assign y14023 = n19406 ;
  assign y14024 = n4757 ;
  assign y14025 = n19411 ;
  assign y14026 = n19414 ;
  assign y14027 = ~n5303 ;
  assign y14028 = ~n19415 ;
  assign y14029 = ~1'b0 ;
  assign y14030 = n19416 ;
  assign y14031 = 1'b0 ;
  assign y14032 = ~n19417 ;
  assign y14033 = ~1'b0 ;
  assign y14034 = ~1'b0 ;
  assign y14035 = n19419 ;
  assign y14036 = n19421 ;
  assign y14037 = n19425 ;
  assign y14038 = ~n19427 ;
  assign y14039 = ~n11389 ;
  assign y14040 = ~1'b0 ;
  assign y14041 = ~1'b0 ;
  assign y14042 = n19429 ;
  assign y14043 = ~1'b0 ;
  assign y14044 = n19430 ;
  assign y14045 = ~n13766 ;
  assign y14046 = ~1'b0 ;
  assign y14047 = ~n19431 ;
  assign y14048 = ~1'b0 ;
  assign y14049 = ~1'b0 ;
  assign y14050 = ~1'b0 ;
  assign y14051 = n19437 ;
  assign y14052 = ~1'b0 ;
  assign y14053 = n5897 ;
  assign y14054 = n19438 ;
  assign y14055 = ~n19439 ;
  assign y14056 = ~1'b0 ;
  assign y14057 = ~n19441 ;
  assign y14058 = ~1'b0 ;
  assign y14059 = ~n19443 ;
  assign y14060 = ~1'b0 ;
  assign y14061 = n19444 ;
  assign y14062 = ~1'b0 ;
  assign y14063 = ~1'b0 ;
  assign y14064 = ~1'b0 ;
  assign y14065 = ~1'b0 ;
  assign y14066 = ~n19445 ;
  assign y14067 = ~n19453 ;
  assign y14068 = ~1'b0 ;
  assign y14069 = n19457 ;
  assign y14070 = ~1'b0 ;
  assign y14071 = ~n19463 ;
  assign y14072 = ~n19466 ;
  assign y14073 = ~1'b0 ;
  assign y14074 = ~n19474 ;
  assign y14075 = 1'b0 ;
  assign y14076 = n19475 ;
  assign y14077 = ~1'b0 ;
  assign y14078 = ~n512 ;
  assign y14079 = n19479 ;
  assign y14080 = ~n19480 ;
  assign y14081 = ~1'b0 ;
  assign y14082 = ~1'b0 ;
  assign y14083 = ~n19484 ;
  assign y14084 = ~n19488 ;
  assign y14085 = ~1'b0 ;
  assign y14086 = ~n19492 ;
  assign y14087 = 1'b0 ;
  assign y14088 = n19493 ;
  assign y14089 = n19498 ;
  assign y14090 = ~1'b0 ;
  assign y14091 = ~1'b0 ;
  assign y14092 = ~n19499 ;
  assign y14093 = ~n19502 ;
  assign y14094 = ~n19503 ;
  assign y14095 = ~n19509 ;
  assign y14096 = ~n1879 ;
  assign y14097 = ~1'b0 ;
  assign y14098 = ~1'b0 ;
  assign y14099 = ~n19511 ;
  assign y14100 = ~1'b0 ;
  assign y14101 = ~1'b0 ;
  assign y14102 = ~n19512 ;
  assign y14103 = ~n19514 ;
  assign y14104 = ~1'b0 ;
  assign y14105 = ~1'b0 ;
  assign y14106 = n19516 ;
  assign y14107 = n19518 ;
  assign y14108 = ~1'b0 ;
  assign y14109 = 1'b0 ;
  assign y14110 = n2699 ;
  assign y14111 = ~1'b0 ;
  assign y14112 = ~n9286 ;
  assign y14113 = ~1'b0 ;
  assign y14114 = n19519 ;
  assign y14115 = ~n19521 ;
  assign y14116 = ~1'b0 ;
  assign y14117 = n19522 ;
  assign y14118 = ~n19524 ;
  assign y14119 = n19530 ;
  assign y14120 = ~1'b0 ;
  assign y14121 = ~1'b0 ;
  assign y14122 = n19532 ;
  assign y14123 = n19534 ;
  assign y14124 = ~n19535 ;
  assign y14125 = n6149 ;
  assign y14126 = n1186 ;
  assign y14127 = n19537 ;
  assign y14128 = ~1'b0 ;
  assign y14129 = n19539 ;
  assign y14130 = ~1'b0 ;
  assign y14131 = ~1'b0 ;
  assign y14132 = ~1'b0 ;
  assign y14133 = ~n19540 ;
  assign y14134 = ~n19549 ;
  assign y14135 = ~1'b0 ;
  assign y14136 = ~1'b0 ;
  assign y14137 = ~1'b0 ;
  assign y14138 = ~1'b0 ;
  assign y14139 = n19550 ;
  assign y14140 = n19553 ;
  assign y14141 = ~1'b0 ;
  assign y14142 = ~n19554 ;
  assign y14143 = n19555 ;
  assign y14144 = ~n19557 ;
  assign y14145 = ~1'b0 ;
  assign y14146 = n19560 ;
  assign y14147 = ~1'b0 ;
  assign y14148 = n19561 ;
  assign y14149 = ~1'b0 ;
  assign y14150 = n19563 ;
  assign y14151 = 1'b0 ;
  assign y14152 = n19567 ;
  assign y14153 = ~n19570 ;
  assign y14154 = ~n19573 ;
  assign y14155 = n19574 ;
  assign y14156 = ~1'b0 ;
  assign y14157 = ~1'b0 ;
  assign y14158 = ~1'b0 ;
  assign y14159 = ~1'b0 ;
  assign y14160 = ~1'b0 ;
  assign y14161 = n19575 ;
  assign y14162 = n16275 ;
  assign y14163 = n19576 ;
  assign y14164 = ~n532 ;
  assign y14165 = n19578 ;
  assign y14166 = ~1'b0 ;
  assign y14167 = ~n19579 ;
  assign y14168 = n19581 ;
  assign y14169 = n19585 ;
  assign y14170 = n19586 ;
  assign y14171 = n19592 ;
  assign y14172 = ~1'b0 ;
  assign y14173 = ~n19594 ;
  assign y14174 = n19595 ;
  assign y14175 = ~n19602 ;
  assign y14176 = ~1'b0 ;
  assign y14177 = ~1'b0 ;
  assign y14178 = ~n19608 ;
  assign y14179 = ~1'b0 ;
  assign y14180 = ~1'b0 ;
  assign y14181 = ~n19609 ;
  assign y14182 = 1'b0 ;
  assign y14183 = ~1'b0 ;
  assign y14184 = ~n3692 ;
  assign y14185 = 1'b0 ;
  assign y14186 = n19612 ;
  assign y14187 = ~n19614 ;
  assign y14188 = ~1'b0 ;
  assign y14189 = n113 ;
  assign y14190 = ~1'b0 ;
  assign y14191 = ~1'b0 ;
  assign y14192 = ~n19615 ;
  assign y14193 = n19621 ;
  assign y14194 = n19622 ;
  assign y14195 = n19624 ;
  assign y14196 = n19626 ;
  assign y14197 = ~n19627 ;
  assign y14198 = ~1'b0 ;
  assign y14199 = n19628 ;
  assign y14200 = ~1'b0 ;
  assign y14201 = n19630 ;
  assign y14202 = ~1'b0 ;
  assign y14203 = n19631 ;
  assign y14204 = n19632 ;
  assign y14205 = ~n1704 ;
  assign y14206 = ~n19635 ;
  assign y14207 = ~1'b0 ;
  assign y14208 = ~1'b0 ;
  assign y14209 = n19637 ;
  assign y14210 = n19648 ;
  assign y14211 = ~n19649 ;
  assign y14212 = ~1'b0 ;
  assign y14213 = ~n19650 ;
  assign y14214 = ~1'b0 ;
  assign y14215 = n19651 ;
  assign y14216 = ~n19653 ;
  assign y14217 = ~n19654 ;
  assign y14218 = n19655 ;
  assign y14219 = ~1'b0 ;
  assign y14220 = n19658 ;
  assign y14221 = ~n19659 ;
  assign y14222 = n19663 ;
  assign y14223 = ~1'b0 ;
  assign y14224 = ~1'b0 ;
  assign y14225 = ~n227 ;
  assign y14226 = n19664 ;
  assign y14227 = ~1'b0 ;
  assign y14228 = n19666 ;
  assign y14229 = ~n19667 ;
  assign y14230 = n19668 ;
  assign y14231 = ~1'b0 ;
  assign y14232 = ~n19670 ;
  assign y14233 = ~n19671 ;
  assign y14234 = ~1'b0 ;
  assign y14235 = n19674 ;
  assign y14236 = ~1'b0 ;
  assign y14237 = 1'b0 ;
  assign y14238 = n19675 ;
  assign y14239 = n19680 ;
  assign y14240 = ~1'b0 ;
  assign y14241 = ~n13608 ;
  assign y14242 = ~n19681 ;
  assign y14243 = ~1'b0 ;
  assign y14244 = n2120 ;
  assign y14245 = ~1'b0 ;
  assign y14246 = ~1'b0 ;
  assign y14247 = 1'b0 ;
  assign y14248 = ~n19683 ;
  assign y14249 = ~n19685 ;
  assign y14250 = n19686 ;
  assign y14251 = n19693 ;
  assign y14252 = ~1'b0 ;
  assign y14253 = ~1'b0 ;
  assign y14254 = ~1'b0 ;
  assign y14255 = n19695 ;
  assign y14256 = ~1'b0 ;
  assign y14257 = ~1'b0 ;
  assign y14258 = 1'b0 ;
  assign y14259 = n19696 ;
  assign y14260 = ~n19698 ;
  assign y14261 = ~n15979 ;
  assign y14262 = n19702 ;
  assign y14263 = ~n13248 ;
  assign y14264 = ~n19704 ;
  assign y14265 = ~n19705 ;
  assign y14266 = n19706 ;
  assign y14267 = ~n19709 ;
  assign y14268 = n19711 ;
  assign y14269 = ~n19712 ;
  assign y14270 = n19714 ;
  assign y14271 = ~1'b0 ;
  assign y14272 = n19715 ;
  assign y14273 = n19720 ;
  assign y14274 = n19724 ;
  assign y14275 = ~n19730 ;
  assign y14276 = ~n19732 ;
  assign y14277 = n19733 ;
  assign y14278 = ~1'b0 ;
  assign y14279 = ~1'b0 ;
  assign y14280 = n19734 ;
  assign y14281 = ~1'b0 ;
  assign y14282 = ~1'b0 ;
  assign y14283 = 1'b0 ;
  assign y14284 = ~n5541 ;
  assign y14285 = ~n19739 ;
  assign y14286 = ~1'b0 ;
  assign y14287 = ~1'b0 ;
  assign y14288 = ~1'b0 ;
  assign y14289 = ~n19740 ;
  assign y14290 = n2571 ;
  assign y14291 = ~n19742 ;
  assign y14292 = ~1'b0 ;
  assign y14293 = ~1'b0 ;
  assign y14294 = n19743 ;
  assign y14295 = ~1'b0 ;
  assign y14296 = ~n19748 ;
  assign y14297 = n19749 ;
  assign y14298 = ~1'b0 ;
  assign y14299 = ~n19752 ;
  assign y14300 = n19753 ;
  assign y14301 = ~1'b0 ;
  assign y14302 = n19754 ;
  assign y14303 = ~1'b0 ;
  assign y14304 = 1'b0 ;
  assign y14305 = 1'b0 ;
  assign y14306 = n19755 ;
  assign y14307 = n11834 ;
  assign y14308 = ~1'b0 ;
  assign y14309 = ~1'b0 ;
  assign y14310 = ~1'b0 ;
  assign y14311 = ~n19756 ;
  assign y14312 = ~1'b0 ;
  assign y14313 = ~1'b0 ;
  assign y14314 = ~1'b0 ;
  assign y14315 = n19760 ;
  assign y14316 = ~1'b0 ;
  assign y14317 = n6433 ;
  assign y14318 = ~1'b0 ;
  assign y14319 = ~n19761 ;
  assign y14320 = n709 ;
  assign y14321 = ~1'b0 ;
  assign y14322 = n19763 ;
  assign y14323 = n19765 ;
  assign y14324 = ~n19767 ;
  assign y14325 = ~n19769 ;
  assign y14326 = ~1'b0 ;
  assign y14327 = n2882 ;
  assign y14328 = ~1'b0 ;
  assign y14329 = ~n19771 ;
  assign y14330 = ~1'b0 ;
  assign y14331 = ~1'b0 ;
  assign y14332 = ~1'b0 ;
  assign y14333 = ~n19773 ;
  assign y14334 = ~1'b0 ;
  assign y14335 = ~1'b0 ;
  assign y14336 = ~n19778 ;
  assign y14337 = n19781 ;
  assign y14338 = ~n19783 ;
  assign y14339 = ~1'b0 ;
  assign y14340 = ~1'b0 ;
  assign y14341 = n19784 ;
  assign y14342 = n19786 ;
  assign y14343 = ~1'b0 ;
  assign y14344 = n19788 ;
  assign y14345 = ~1'b0 ;
  assign y14346 = ~n19796 ;
  assign y14347 = ~n9008 ;
  assign y14348 = n19801 ;
  assign y14349 = ~n19804 ;
  assign y14350 = n19806 ;
  assign y14351 = ~1'b0 ;
  assign y14352 = ~1'b0 ;
  assign y14353 = ~n10923 ;
  assign y14354 = n19808 ;
  assign y14355 = n19816 ;
  assign y14356 = ~1'b0 ;
  assign y14357 = ~1'b0 ;
  assign y14358 = ~1'b0 ;
  assign y14359 = ~n19818 ;
  assign y14360 = ~n19819 ;
  assign y14361 = ~1'b0 ;
  assign y14362 = ~n19820 ;
  assign y14363 = ~1'b0 ;
  assign y14364 = ~1'b0 ;
  assign y14365 = ~1'b0 ;
  assign y14366 = ~1'b0 ;
  assign y14367 = 1'b0 ;
  assign y14368 = ~1'b0 ;
  assign y14369 = ~n14266 ;
  assign y14370 = n47 ;
  assign y14371 = n10357 ;
  assign y14372 = ~1'b0 ;
  assign y14373 = n18011 ;
  assign y14374 = ~n2789 ;
  assign y14375 = 1'b0 ;
  assign y14376 = ~n5830 ;
  assign y14377 = 1'b0 ;
  assign y14378 = ~n19827 ;
  assign y14379 = ~n19828 ;
  assign y14380 = ~1'b0 ;
  assign y14381 = ~1'b0 ;
  assign y14382 = 1'b0 ;
  assign y14383 = ~n19829 ;
  assign y14384 = ~n6451 ;
  assign y14385 = ~1'b0 ;
  assign y14386 = ~1'b0 ;
  assign y14387 = ~1'b0 ;
  assign y14388 = n19830 ;
  assign y14389 = ~1'b0 ;
  assign y14390 = n19832 ;
  assign y14391 = ~1'b0 ;
  assign y14392 = n19834 ;
  assign y14393 = n19836 ;
  assign y14394 = ~n52 ;
  assign y14395 = n19837 ;
  assign y14396 = ~n19840 ;
  assign y14397 = ~n19847 ;
  assign y14398 = ~1'b0 ;
  assign y14399 = ~1'b0 ;
  assign y14400 = ~1'b0 ;
  assign y14401 = n19850 ;
  assign y14402 = n19851 ;
  assign y14403 = n19852 ;
  assign y14404 = n19853 ;
  assign y14405 = n19857 ;
  assign y14406 = n19864 ;
  assign y14407 = ~n19865 ;
  assign y14408 = ~1'b0 ;
  assign y14409 = n19868 ;
  assign y14410 = ~n19869 ;
  assign y14411 = ~n19877 ;
  assign y14412 = ~1'b0 ;
  assign y14413 = ~1'b0 ;
  assign y14414 = ~n19879 ;
  assign y14415 = ~n19881 ;
  assign y14416 = ~n5780 ;
  assign y14417 = 1'b0 ;
  assign y14418 = ~1'b0 ;
  assign y14419 = n19882 ;
  assign y14420 = ~n19894 ;
  assign y14421 = n19897 ;
  assign y14422 = ~1'b0 ;
  assign y14423 = n19899 ;
  assign y14424 = ~1'b0 ;
  assign y14425 = ~n19900 ;
  assign y14426 = ~1'b0 ;
  assign y14427 = ~1'b0 ;
  assign y14428 = ~n19902 ;
  assign y14429 = n17974 ;
  assign y14430 = ~n19904 ;
  assign y14431 = ~n19905 ;
  assign y14432 = n5815 ;
  assign y14433 = n19906 ;
  assign y14434 = n19910 ;
  assign y14435 = ~n19911 ;
  assign y14436 = ~1'b0 ;
  assign y14437 = n2322 ;
  assign y14438 = n19913 ;
  assign y14439 = n6440 ;
  assign y14440 = n19914 ;
  assign y14441 = n19915 ;
  assign y14442 = ~1'b0 ;
  assign y14443 = ~1'b0 ;
  assign y14444 = ~n19932 ;
  assign y14445 = n19933 ;
  assign y14446 = ~1'b0 ;
  assign y14447 = n68 ;
  assign y14448 = ~n19937 ;
  assign y14449 = ~1'b0 ;
  assign y14450 = ~1'b0 ;
  assign y14451 = ~n19940 ;
  assign y14452 = n6120 ;
  assign y14453 = n19941 ;
  assign y14454 = n19943 ;
  assign y14455 = ~1'b0 ;
  assign y14456 = n19945 ;
  assign y14457 = n19954 ;
  assign y14458 = ~1'b0 ;
  assign y14459 = ~n19956 ;
  assign y14460 = ~n7472 ;
  assign y14461 = ~1'b0 ;
  assign y14462 = ~1'b0 ;
  assign y14463 = ~1'b0 ;
  assign y14464 = ~1'b0 ;
  assign y14465 = ~1'b0 ;
  assign y14466 = ~1'b0 ;
  assign y14467 = ~1'b0 ;
  assign y14468 = ~n3679 ;
  assign y14469 = ~1'b0 ;
  assign y14470 = 1'b0 ;
  assign y14471 = ~n19966 ;
  assign y14472 = ~n19968 ;
  assign y14473 = ~1'b0 ;
  assign y14474 = ~1'b0 ;
  assign y14475 = ~1'b0 ;
  assign y14476 = ~n19970 ;
  assign y14477 = ~1'b0 ;
  assign y14478 = 1'b0 ;
  assign y14479 = ~1'b0 ;
  assign y14480 = ~n14385 ;
  assign y14481 = ~1'b0 ;
  assign y14482 = ~1'b0 ;
  assign y14483 = ~n19973 ;
  assign y14484 = ~n7767 ;
  assign y14485 = ~n19974 ;
  assign y14486 = ~1'b0 ;
  assign y14487 = n19985 ;
  assign y14488 = ~1'b0 ;
  assign y14489 = ~1'b0 ;
  assign y14490 = ~1'b0 ;
  assign y14491 = n19986 ;
  assign y14492 = ~n19988 ;
  assign y14493 = ~n19990 ;
  assign y14494 = n520 ;
  assign y14495 = ~n55 ;
  assign y14496 = n19996 ;
  assign y14497 = ~n20000 ;
  assign y14498 = ~n20006 ;
  assign y14499 = n20010 ;
  assign y14500 = n20011 ;
  assign y14501 = ~1'b0 ;
  assign y14502 = n20012 ;
  assign y14503 = ~n20013 ;
  assign y14504 = ~n3320 ;
  assign y14505 = 1'b0 ;
  assign y14506 = n20017 ;
  assign y14507 = ~1'b0 ;
  assign y14508 = ~n20019 ;
  assign y14509 = ~1'b0 ;
  assign y14510 = n20022 ;
  assign y14511 = ~1'b0 ;
  assign y14512 = ~n20028 ;
  assign y14513 = ~n20029 ;
  assign y14514 = n20031 ;
  assign y14515 = ~1'b0 ;
  assign y14516 = n20033 ;
  assign y14517 = ~1'b0 ;
  assign y14518 = ~1'b0 ;
  assign y14519 = n20036 ;
  assign y14520 = ~n20037 ;
  assign y14521 = ~1'b0 ;
  assign y14522 = n3124 ;
  assign y14523 = n20039 ;
  assign y14524 = ~1'b0 ;
  assign y14525 = n20040 ;
  assign y14526 = ~1'b0 ;
  assign y14527 = ~n20042 ;
  assign y14528 = ~1'b0 ;
  assign y14529 = n20045 ;
  assign y14530 = ~1'b0 ;
  assign y14531 = n20046 ;
  assign y14532 = ~1'b0 ;
  assign y14533 = ~1'b0 ;
  assign y14534 = n20047 ;
  assign y14535 = n20048 ;
  assign y14536 = ~1'b0 ;
  assign y14537 = ~1'b0 ;
  assign y14538 = n19803 ;
  assign y14539 = ~n20050 ;
  assign y14540 = ~n20053 ;
  assign y14541 = ~n18771 ;
  assign y14542 = ~n20054 ;
  assign y14543 = n20055 ;
  assign y14544 = ~1'b0 ;
  assign y14545 = ~1'b0 ;
  assign y14546 = ~n20059 ;
  assign y14547 = ~1'b0 ;
  assign y14548 = ~n20060 ;
  assign y14549 = ~n20061 ;
  assign y14550 = ~1'b0 ;
  assign y14551 = 1'b0 ;
  assign y14552 = ~n13118 ;
  assign y14553 = ~n20069 ;
  assign y14554 = n20071 ;
  assign y14555 = ~n11222 ;
  assign y14556 = ~n3718 ;
  assign y14557 = n20078 ;
  assign y14558 = ~n20081 ;
  assign y14559 = n2041 ;
  assign y14560 = ~n20082 ;
  assign y14561 = ~1'b0 ;
  assign y14562 = ~1'b0 ;
  assign y14563 = ~1'b0 ;
  assign y14564 = ~n20084 ;
  assign y14565 = n20086 ;
  assign y14566 = ~n20089 ;
  assign y14567 = ~1'b0 ;
  assign y14568 = ~1'b0 ;
  assign y14569 = n20091 ;
  assign y14570 = n20092 ;
  assign y14571 = ~n20096 ;
  assign y14572 = n20098 ;
  assign y14573 = n20099 ;
  assign y14574 = ~n20100 ;
  assign y14575 = n20101 ;
  assign y14576 = n2083 ;
  assign y14577 = ~n20102 ;
  assign y14578 = ~1'b0 ;
  assign y14579 = n20103 ;
  assign y14580 = ~1'b0 ;
  assign y14581 = ~1'b0 ;
  assign y14582 = n20107 ;
  assign y14583 = ~n20112 ;
  assign y14584 = ~1'b0 ;
  assign y14585 = ~n20115 ;
  assign y14586 = n12099 ;
  assign y14587 = ~1'b0 ;
  assign y14588 = ~1'b0 ;
  assign y14589 = ~1'b0 ;
  assign y14590 = n20118 ;
  assign y14591 = n20119 ;
  assign y14592 = ~1'b0 ;
  assign y14593 = n594 ;
  assign y14594 = ~1'b0 ;
  assign y14595 = ~n20122 ;
  assign y14596 = ~1'b0 ;
  assign y14597 = n20126 ;
  assign y14598 = n20129 ;
  assign y14599 = n866 ;
  assign y14600 = ~1'b0 ;
  assign y14601 = ~1'b0 ;
  assign y14602 = n20130 ;
  assign y14603 = ~1'b0 ;
  assign y14604 = n20132 ;
  assign y14605 = ~n20133 ;
  assign y14606 = ~n20134 ;
  assign y14607 = n20135 ;
  assign y14608 = ~1'b0 ;
  assign y14609 = n20136 ;
  assign y14610 = ~n20138 ;
  assign y14611 = n20139 ;
  assign y14612 = 1'b0 ;
  assign y14613 = ~1'b0 ;
  assign y14614 = ~n16518 ;
  assign y14615 = ~1'b0 ;
  assign y14616 = ~n20142 ;
  assign y14617 = n20143 ;
  assign y14618 = ~n20145 ;
  assign y14619 = ~n20148 ;
  assign y14620 = n20184 ;
  assign y14621 = n20187 ;
  assign y14622 = ~n20189 ;
  assign y14623 = ~n20190 ;
  assign y14624 = ~n20191 ;
  assign y14625 = n20192 ;
  assign y14626 = ~1'b0 ;
  assign y14627 = n20194 ;
  assign y14628 = ~1'b0 ;
  assign y14629 = ~n6381 ;
  assign y14630 = ~n20195 ;
  assign y14631 = n20198 ;
  assign y14632 = n20203 ;
  assign y14633 = ~n20204 ;
  assign y14634 = ~n20205 ;
  assign y14635 = ~n20208 ;
  assign y14636 = ~1'b0 ;
  assign y14637 = ~1'b0 ;
  assign y14638 = n20210 ;
  assign y14639 = n20214 ;
  assign y14640 = n20221 ;
  assign y14641 = ~n20222 ;
  assign y14642 = n20225 ;
  assign y14643 = ~1'b0 ;
  assign y14644 = ~1'b0 ;
  assign y14645 = ~n20230 ;
  assign y14646 = ~n20232 ;
  assign y14647 = ~1'b0 ;
  assign y14648 = 1'b0 ;
  assign y14649 = ~n20233 ;
  assign y14650 = ~n20235 ;
  assign y14651 = n20237 ;
  assign y14652 = ~1'b0 ;
  assign y14653 = ~n4906 ;
  assign y14654 = ~1'b0 ;
  assign y14655 = ~1'b0 ;
  assign y14656 = n20238 ;
  assign y14657 = n20242 ;
  assign y14658 = n20243 ;
  assign y14659 = ~n20244 ;
  assign y14660 = 1'b0 ;
  assign y14661 = ~1'b0 ;
  assign y14662 = ~n17383 ;
  assign y14663 = 1'b0 ;
  assign y14664 = ~1'b0 ;
  assign y14665 = ~1'b0 ;
  assign y14666 = n20245 ;
  assign y14667 = ~1'b0 ;
  assign y14668 = ~n20246 ;
  assign y14669 = n20248 ;
  assign y14670 = ~1'b0 ;
  assign y14671 = ~n20249 ;
  assign y14672 = n20252 ;
  assign y14673 = ~n294 ;
  assign y14674 = ~n20253 ;
  assign y14675 = ~n20254 ;
  assign y14676 = n11533 ;
  assign y14677 = n6333 ;
  assign y14678 = ~n20255 ;
  assign y14679 = n20258 ;
  assign y14680 = ~1'b0 ;
  assign y14681 = n7596 ;
  assign y14682 = ~n20263 ;
  assign y14683 = n20266 ;
  assign y14684 = ~1'b0 ;
  assign y14685 = ~n20267 ;
  assign y14686 = ~n20272 ;
  assign y14687 = ~1'b0 ;
  assign y14688 = ~n20275 ;
  assign y14689 = n3533 ;
  assign y14690 = 1'b0 ;
  assign y14691 = n20276 ;
  assign y14692 = n20278 ;
  assign y14693 = n20280 ;
  assign y14694 = 1'b0 ;
  assign y14695 = ~1'b0 ;
  assign y14696 = n20281 ;
  assign y14697 = n20283 ;
  assign y14698 = n20284 ;
  assign y14699 = ~n20286 ;
  assign y14700 = ~1'b0 ;
  assign y14701 = n1922 ;
  assign y14702 = ~1'b0 ;
  assign y14703 = ~1'b0 ;
  assign y14704 = ~1'b0 ;
  assign y14705 = ~n20287 ;
  assign y14706 = n20289 ;
  assign y14707 = n20290 ;
  assign y14708 = n20291 ;
  assign y14709 = ~n20292 ;
  assign y14710 = n2662 ;
  assign y14711 = ~n20296 ;
  assign y14712 = n20301 ;
  assign y14713 = ~n20303 ;
  assign y14714 = n20304 ;
  assign y14715 = n20309 ;
  assign y14716 = ~n20310 ;
  assign y14717 = n20311 ;
  assign y14718 = ~n20312 ;
  assign y14719 = ~1'b0 ;
  assign y14720 = ~n20315 ;
  assign y14721 = ~1'b0 ;
  assign y14722 = n20317 ;
  assign y14723 = ~n20320 ;
  assign y14724 = n20321 ;
  assign y14725 = ~n20324 ;
  assign y14726 = n20325 ;
  assign y14727 = 1'b0 ;
  assign y14728 = ~1'b0 ;
  assign y14729 = n20328 ;
  assign y14730 = n20333 ;
  assign y14731 = ~1'b0 ;
  assign y14732 = ~1'b0 ;
  assign y14733 = n20334 ;
  assign y14734 = ~1'b0 ;
  assign y14735 = ~n20339 ;
  assign y14736 = ~1'b0 ;
  assign y14737 = ~1'b0 ;
  assign y14738 = ~n20342 ;
  assign y14739 = ~1'b0 ;
  assign y14740 = ~1'b0 ;
  assign y14741 = ~1'b0 ;
  assign y14742 = n20347 ;
  assign y14743 = ~n20351 ;
  assign y14744 = n20353 ;
  assign y14745 = ~1'b0 ;
  assign y14746 = ~1'b0 ;
  assign y14747 = ~n20354 ;
  assign y14748 = n19937 ;
  assign y14749 = n20356 ;
  assign y14750 = ~1'b0 ;
  assign y14751 = ~1'b0 ;
  assign y14752 = ~1'b0 ;
  assign y14753 = n20357 ;
  assign y14754 = n8054 ;
  assign y14755 = ~n20359 ;
  assign y14756 = n20360 ;
  assign y14757 = ~n20361 ;
  assign y14758 = n20363 ;
  assign y14759 = n20365 ;
  assign y14760 = ~n20372 ;
  assign y14761 = ~n20374 ;
  assign y14762 = n20379 ;
  assign y14763 = 1'b0 ;
  assign y14764 = ~n20383 ;
  assign y14765 = ~n19896 ;
  assign y14766 = n20386 ;
  assign y14767 = ~1'b0 ;
  assign y14768 = 1'b0 ;
  assign y14769 = ~1'b0 ;
  assign y14770 = ~1'b0 ;
  assign y14771 = n20387 ;
  assign y14772 = ~1'b0 ;
  assign y14773 = ~n20389 ;
  assign y14774 = ~1'b0 ;
  assign y14775 = n7346 ;
  assign y14776 = 1'b0 ;
  assign y14777 = ~1'b0 ;
  assign y14778 = ~n20391 ;
  assign y14779 = ~1'b0 ;
  assign y14780 = ~n20392 ;
  assign y14781 = ~1'b0 ;
  assign y14782 = ~1'b0 ;
  assign y14783 = n9061 ;
  assign y14784 = ~n20394 ;
  assign y14785 = n4730 ;
  assign y14786 = ~n20397 ;
  assign y14787 = ~1'b0 ;
  assign y14788 = ~1'b0 ;
  assign y14789 = n20400 ;
  assign y14790 = n20401 ;
  assign y14791 = ~n20402 ;
  assign y14792 = ~n20411 ;
  assign y14793 = ~1'b0 ;
  assign y14794 = ~1'b0 ;
  assign y14795 = ~1'b0 ;
  assign y14796 = ~n20412 ;
  assign y14797 = ~n20414 ;
  assign y14798 = n20416 ;
  assign y14799 = n20417 ;
  assign y14800 = n20419 ;
  assign y14801 = n20420 ;
  assign y14802 = n20422 ;
  assign y14803 = 1'b0 ;
  assign y14804 = ~1'b0 ;
  assign y14805 = ~n20423 ;
  assign y14806 = n20425 ;
  assign y14807 = n20427 ;
  assign y14808 = ~n20428 ;
  assign y14809 = n20430 ;
  assign y14810 = ~1'b0 ;
  assign y14811 = ~n20432 ;
  assign y14812 = ~1'b0 ;
  assign y14813 = ~n20434 ;
  assign y14814 = ~1'b0 ;
  assign y14815 = ~n20436 ;
  assign y14816 = n7674 ;
  assign y14817 = ~1'b0 ;
  assign y14818 = n20425 ;
  assign y14819 = n20439 ;
  assign y14820 = ~1'b0 ;
  assign y14821 = ~n20441 ;
  assign y14822 = ~n20443 ;
  assign y14823 = 1'b0 ;
  assign y14824 = ~n20447 ;
  assign y14825 = ~1'b0 ;
  assign y14826 = ~n20449 ;
  assign y14827 = 1'b0 ;
  assign y14828 = ~n20451 ;
  assign y14829 = ~n14454 ;
  assign y14830 = n20454 ;
  assign y14831 = ~n20461 ;
  assign y14832 = n20467 ;
  assign y14833 = ~1'b0 ;
  assign y14834 = ~n20468 ;
  assign y14835 = ~1'b0 ;
  assign y14836 = ~n20469 ;
  assign y14837 = ~1'b0 ;
  assign y14838 = n20470 ;
  assign y14839 = ~1'b0 ;
  assign y14840 = ~n20472 ;
  assign y14841 = ~n19934 ;
  assign y14842 = ~1'b0 ;
  assign y14843 = ~1'b0 ;
  assign y14844 = ~n20473 ;
  assign y14845 = 1'b0 ;
  assign y14846 = n20474 ;
  assign y14847 = ~n20476 ;
  assign y14848 = n20478 ;
  assign y14849 = ~n20482 ;
  assign y14850 = n20483 ;
  assign y14851 = ~n20486 ;
  assign y14852 = ~n4740 ;
  assign y14853 = n20488 ;
  assign y14854 = ~n20490 ;
  assign y14855 = ~1'b0 ;
  assign y14856 = 1'b0 ;
  assign y14857 = ~n20493 ;
  assign y14858 = n20496 ;
  assign y14859 = ~1'b0 ;
  assign y14860 = ~1'b0 ;
  assign y14861 = ~1'b0 ;
  assign y14862 = ~1'b0 ;
  assign y14863 = ~n20501 ;
  assign y14864 = ~1'b0 ;
  assign y14865 = n20503 ;
  assign y14866 = n20504 ;
  assign y14867 = 1'b0 ;
  assign y14868 = ~1'b0 ;
  assign y14869 = ~n20510 ;
  assign y14870 = n20511 ;
  assign y14871 = ~n20512 ;
  assign y14872 = n20513 ;
  assign y14873 = 1'b0 ;
  assign y14874 = ~n15028 ;
  assign y14875 = ~1'b0 ;
  assign y14876 = ~n20514 ;
  assign y14877 = ~n20515 ;
  assign y14878 = n20516 ;
  assign y14879 = ~1'b0 ;
  assign y14880 = 1'b0 ;
  assign y14881 = ~1'b0 ;
  assign y14882 = ~n20520 ;
  assign y14883 = n20521 ;
  assign y14884 = ~1'b0 ;
  assign y14885 = ~1'b0 ;
  assign y14886 = n20522 ;
  assign y14887 = n20523 ;
  assign y14888 = ~n20527 ;
  assign y14889 = ~1'b0 ;
  assign y14890 = n20528 ;
  assign y14891 = n16906 ;
  assign y14892 = n20533 ;
  assign y14893 = 1'b0 ;
  assign y14894 = ~n16918 ;
  assign y14895 = ~1'b0 ;
  assign y14896 = ~n20539 ;
  assign y14897 = ~n20541 ;
  assign y14898 = ~n20547 ;
  assign y14899 = n20549 ;
  assign y14900 = ~n20551 ;
  assign y14901 = ~1'b0 ;
  assign y14902 = ~1'b0 ;
  assign y14903 = n20552 ;
  assign y14904 = n20553 ;
  assign y14905 = ~n20558 ;
  assign y14906 = 1'b0 ;
  assign y14907 = ~1'b0 ;
  assign y14908 = n1233 ;
  assign y14909 = n20561 ;
  assign y14910 = n20567 ;
  assign y14911 = ~1'b0 ;
  assign y14912 = ~1'b0 ;
  assign y14913 = n11089 ;
  assign y14914 = ~1'b0 ;
  assign y14915 = n4193 ;
  assign y14916 = n20569 ;
  assign y14917 = ~1'b0 ;
  assign y14918 = ~n20572 ;
  assign y14919 = n20575 ;
  assign y14920 = n20576 ;
  assign y14921 = ~n20581 ;
  assign y14922 = ~1'b0 ;
  assign y14923 = n20582 ;
  assign y14924 = n20585 ;
  assign y14925 = ~1'b0 ;
  assign y14926 = n20586 ;
  assign y14927 = ~n20588 ;
  assign y14928 = ~1'b0 ;
  assign y14929 = n20589 ;
  assign y14930 = ~n20591 ;
  assign y14931 = n2825 ;
  assign y14932 = ~1'b0 ;
  assign y14933 = n20593 ;
  assign y14934 = ~n20594 ;
  assign y14935 = ~n20595 ;
  assign y14936 = n7304 ;
  assign y14937 = ~1'b0 ;
  assign y14938 = ~1'b0 ;
  assign y14939 = ~n20597 ;
  assign y14940 = ~n20604 ;
  assign y14941 = ~n7271 ;
  assign y14942 = ~1'b0 ;
  assign y14943 = ~1'b0 ;
  assign y14944 = ~n374 ;
  assign y14945 = ~1'b0 ;
  assign y14946 = n20605 ;
  assign y14947 = n20607 ;
  assign y14948 = n20611 ;
  assign y14949 = ~n20612 ;
  assign y14950 = n9634 ;
  assign y14951 = ~n20614 ;
  assign y14952 = ~n20618 ;
  assign y14953 = n20620 ;
  assign y14954 = ~1'b0 ;
  assign y14955 = ~n10514 ;
  assign y14956 = ~n20626 ;
  assign y14957 = ~n20628 ;
  assign y14958 = ~1'b0 ;
  assign y14959 = ~1'b0 ;
  assign y14960 = ~n20631 ;
  assign y14961 = ~1'b0 ;
  assign y14962 = ~1'b0 ;
  assign y14963 = ~1'b0 ;
  assign y14964 = 1'b0 ;
  assign y14965 = ~n20637 ;
  assign y14966 = ~n20640 ;
  assign y14967 = ~n20641 ;
  assign y14968 = ~1'b0 ;
  assign y14969 = ~n20644 ;
  assign y14970 = ~n20645 ;
  assign y14971 = ~1'b0 ;
  assign y14972 = ~n20648 ;
  assign y14973 = ~1'b0 ;
  assign y14974 = ~n3137 ;
  assign y14975 = n20649 ;
  assign y14976 = ~n20656 ;
  assign y14977 = ~n20659 ;
  assign y14978 = ~1'b0 ;
  assign y14979 = n20664 ;
  assign y14980 = n20666 ;
  assign y14981 = 1'b0 ;
  assign y14982 = n20669 ;
  assign y14983 = ~1'b0 ;
  assign y14984 = ~1'b0 ;
  assign y14985 = 1'b0 ;
  assign y14986 = ~1'b0 ;
  assign y14987 = ~1'b0 ;
  assign y14988 = ~1'b0 ;
  assign y14989 = n20670 ;
  assign y14990 = ~n20672 ;
  assign y14991 = ~n20674 ;
  assign y14992 = ~n20676 ;
  assign y14993 = ~n20677 ;
  assign y14994 = ~n20681 ;
  assign y14995 = n20684 ;
  assign y14996 = ~n20686 ;
  assign y14997 = ~n20688 ;
  assign y14998 = ~1'b0 ;
  assign y14999 = ~1'b0 ;
  assign y15000 = 1'b0 ;
  assign y15001 = n638 ;
  assign y15002 = n20690 ;
  assign y15003 = ~n20692 ;
  assign y15004 = n16491 ;
  assign y15005 = ~1'b0 ;
  assign y15006 = ~1'b0 ;
  assign y15007 = ~1'b0 ;
  assign y15008 = ~n20693 ;
  assign y15009 = n20700 ;
  assign y15010 = ~n15402 ;
  assign y15011 = ~1'b0 ;
  assign y15012 = n13327 ;
  assign y15013 = ~1'b0 ;
  assign y15014 = n20708 ;
  assign y15015 = n20709 ;
  assign y15016 = ~n20710 ;
  assign y15017 = n20715 ;
  assign y15018 = n20716 ;
  assign y15019 = ~n20718 ;
  assign y15020 = ~n20721 ;
  assign y15021 = ~1'b0 ;
  assign y15022 = ~n20725 ;
  assign y15023 = n20729 ;
  assign y15024 = n20731 ;
  assign y15025 = n20733 ;
  assign y15026 = n20735 ;
  assign y15027 = ~n20742 ;
  assign y15028 = ~n20744 ;
  assign y15029 = n20745 ;
  assign y15030 = ~n20751 ;
  assign y15031 = n20753 ;
  assign y15032 = ~1'b0 ;
  assign y15033 = n20754 ;
  assign y15034 = ~1'b0 ;
  assign y15035 = ~1'b0 ;
  assign y15036 = ~1'b0 ;
  assign y15037 = ~1'b0 ;
  assign y15038 = ~1'b0 ;
  assign y15039 = ~n20755 ;
  assign y15040 = n20760 ;
  assign y15041 = ~1'b0 ;
  assign y15042 = n15912 ;
  assign y15043 = n20763 ;
  assign y15044 = ~n5972 ;
  assign y15045 = ~n20766 ;
  assign y15046 = ~n13585 ;
  assign y15047 = ~1'b0 ;
  assign y15048 = ~n20767 ;
  assign y15049 = ~1'b0 ;
  assign y15050 = 1'b0 ;
  assign y15051 = ~1'b0 ;
  assign y15052 = ~1'b0 ;
  assign y15053 = n20768 ;
  assign y15054 = ~1'b0 ;
  assign y15055 = n20771 ;
  assign y15056 = ~1'b0 ;
  assign y15057 = ~1'b0 ;
  assign y15058 = ~n20772 ;
  assign y15059 = ~n20775 ;
  assign y15060 = ~n20777 ;
  assign y15061 = ~n20778 ;
  assign y15062 = ~1'b0 ;
  assign y15063 = n20779 ;
  assign y15064 = n20780 ;
  assign y15065 = ~1'b0 ;
  assign y15066 = ~1'b0 ;
  assign y15067 = ~n20781 ;
  assign y15068 = n11174 ;
  assign y15069 = ~n20782 ;
  assign y15070 = ~1'b0 ;
  assign y15071 = ~n20783 ;
  assign y15072 = ~n20788 ;
  assign y15073 = ~1'b0 ;
  assign y15074 = ~n17115 ;
  assign y15075 = n4535 ;
  assign y15076 = ~1'b0 ;
  assign y15077 = ~n20789 ;
  assign y15078 = n20790 ;
  assign y15079 = ~1'b0 ;
  assign y15080 = ~n20792 ;
  assign y15081 = 1'b0 ;
  assign y15082 = ~1'b0 ;
  assign y15083 = ~n20807 ;
  assign y15084 = ~n20809 ;
  assign y15085 = n20813 ;
  assign y15086 = ~1'b0 ;
  assign y15087 = n20814 ;
  assign y15088 = ~n10824 ;
  assign y15089 = ~n20818 ;
  assign y15090 = ~1'b0 ;
  assign y15091 = n20819 ;
  assign y15092 = n20820 ;
  assign y15093 = ~1'b0 ;
  assign y15094 = ~1'b0 ;
  assign y15095 = ~n20822 ;
  assign y15096 = ~1'b0 ;
  assign y15097 = ~n20826 ;
  assign y15098 = n20833 ;
  assign y15099 = ~n20841 ;
  assign y15100 = n20846 ;
  assign y15101 = ~1'b0 ;
  assign y15102 = ~n1001 ;
  assign y15103 = ~1'b0 ;
  assign y15104 = ~1'b0 ;
  assign y15105 = ~1'b0 ;
  assign y15106 = ~n20848 ;
  assign y15107 = ~1'b0 ;
  assign y15108 = ~n20849 ;
  assign y15109 = n3061 ;
  assign y15110 = ~n20850 ;
  assign y15111 = n20871 ;
  assign y15112 = ~n13661 ;
  assign y15113 = ~1'b0 ;
  assign y15114 = 1'b0 ;
  assign y15115 = ~1'b0 ;
  assign y15116 = ~n20872 ;
  assign y15117 = ~1'b0 ;
  assign y15118 = ~n20873 ;
  assign y15119 = ~1'b0 ;
  assign y15120 = ~1'b0 ;
  assign y15121 = ~1'b0 ;
  assign y15122 = ~n20875 ;
  assign y15123 = ~n20892 ;
  assign y15124 = ~1'b0 ;
  assign y15125 = ~1'b0 ;
  assign y15126 = ~1'b0 ;
  assign y15127 = n20900 ;
  assign y15128 = ~n20904 ;
  assign y15129 = ~1'b0 ;
  assign y15130 = n764 ;
  assign y15131 = ~n20942 ;
  assign y15132 = n20943 ;
  assign y15133 = n13798 ;
  assign y15134 = ~1'b0 ;
  assign y15135 = n11272 ;
  assign y15136 = ~n20945 ;
  assign y15137 = n20946 ;
  assign y15138 = n20947 ;
  assign y15139 = n20948 ;
  assign y15140 = ~n20951 ;
  assign y15141 = ~n20954 ;
  assign y15142 = n20955 ;
  assign y15143 = ~n20956 ;
  assign y15144 = 1'b0 ;
  assign y15145 = ~1'b0 ;
  assign y15146 = n20957 ;
  assign y15147 = ~n20959 ;
  assign y15148 = n20961 ;
  assign y15149 = n20962 ;
  assign y15150 = n20964 ;
  assign y15151 = n616 ;
  assign y15152 = ~1'b0 ;
  assign y15153 = ~1'b0 ;
  assign y15154 = ~1'b0 ;
  assign y15155 = ~n20968 ;
  assign y15156 = ~1'b0 ;
  assign y15157 = ~n20969 ;
  assign y15158 = ~1'b0 ;
  assign y15159 = ~1'b0 ;
  assign y15160 = ~1'b0 ;
  assign y15161 = n20970 ;
  assign y15162 = n20972 ;
  assign y15163 = ~n14256 ;
  assign y15164 = ~n20974 ;
  assign y15165 = ~1'b0 ;
  assign y15166 = n20976 ;
  assign y15167 = ~n9431 ;
  assign y15168 = ~1'b0 ;
  assign y15169 = ~n20989 ;
  assign y15170 = ~n10551 ;
  assign y15171 = n20990 ;
  assign y15172 = ~n20992 ;
  assign y15173 = ~1'b0 ;
  assign y15174 = n20996 ;
  assign y15175 = ~1'b0 ;
  assign y15176 = ~1'b0 ;
  assign y15177 = n20998 ;
  assign y15178 = ~1'b0 ;
  assign y15179 = ~n20999 ;
  assign y15180 = ~1'b0 ;
  assign y15181 = ~1'b0 ;
  assign y15182 = n21001 ;
  assign y15183 = ~1'b0 ;
  assign y15184 = n21005 ;
  assign y15185 = ~n21008 ;
  assign y15186 = n21011 ;
  assign y15187 = ~n8627 ;
  assign y15188 = n21014 ;
  assign y15189 = 1'b0 ;
  assign y15190 = ~n21015 ;
  assign y15191 = n18415 ;
  assign y15192 = ~1'b0 ;
  assign y15193 = 1'b0 ;
  assign y15194 = n21017 ;
  assign y15195 = ~1'b0 ;
  assign y15196 = 1'b0 ;
  assign y15197 = n21019 ;
  assign y15198 = n21021 ;
  assign y15199 = n21025 ;
  assign y15200 = 1'b0 ;
  assign y15201 = ~1'b0 ;
  assign y15202 = ~1'b0 ;
  assign y15203 = ~1'b0 ;
  assign y15204 = ~n21029 ;
  assign y15205 = n21033 ;
  assign y15206 = n16007 ;
  assign y15207 = n21037 ;
  assign y15208 = n21039 ;
  assign y15209 = ~n21041 ;
  assign y15210 = n21042 ;
  assign y15211 = ~1'b0 ;
  assign y15212 = ~n21043 ;
  assign y15213 = ~1'b0 ;
  assign y15214 = 1'b0 ;
  assign y15215 = ~1'b0 ;
  assign y15216 = n21045 ;
  assign y15217 = n21049 ;
  assign y15218 = ~1'b0 ;
  assign y15219 = n21051 ;
  assign y15220 = ~1'b0 ;
  assign y15221 = ~1'b0 ;
  assign y15222 = ~n21055 ;
  assign y15223 = n21056 ;
  assign y15224 = ~1'b0 ;
  assign y15225 = ~1'b0 ;
  assign y15226 = ~1'b0 ;
  assign y15227 = n21057 ;
  assign y15228 = ~1'b0 ;
  assign y15229 = n501 ;
  assign y15230 = n21061 ;
  assign y15231 = ~1'b0 ;
  assign y15232 = n21062 ;
  assign y15233 = n21063 ;
  assign y15234 = n21068 ;
  assign y15235 = n5632 ;
  assign y15236 = n21069 ;
  assign y15237 = n21075 ;
  assign y15238 = n21076 ;
  assign y15239 = ~1'b0 ;
  assign y15240 = n21081 ;
  assign y15241 = ~1'b0 ;
  assign y15242 = ~1'b0 ;
  assign y15243 = ~1'b0 ;
  assign y15244 = n6944 ;
  assign y15245 = ~n21084 ;
  assign y15246 = 1'b0 ;
  assign y15247 = ~1'b0 ;
  assign y15248 = ~n21086 ;
  assign y15249 = ~n21087 ;
  assign y15250 = ~n21088 ;
  assign y15251 = ~n21090 ;
  assign y15252 = ~n21091 ;
  assign y15253 = ~1'b0 ;
  assign y15254 = ~n21096 ;
  assign y15255 = ~1'b0 ;
  assign y15256 = ~1'b0 ;
  assign y15257 = ~n21098 ;
  assign y15258 = ~n5192 ;
  assign y15259 = n21109 ;
  assign y15260 = ~n21112 ;
  assign y15261 = 1'b0 ;
  assign y15262 = n21113 ;
  assign y15263 = n21114 ;
  assign y15264 = ~1'b0 ;
  assign y15265 = n21116 ;
  assign y15266 = ~1'b0 ;
  assign y15267 = ~1'b0 ;
  assign y15268 = ~n1847 ;
  assign y15269 = ~n21121 ;
  assign y15270 = ~n21123 ;
  assign y15271 = ~n21124 ;
  assign y15272 = ~n21126 ;
  assign y15273 = n21129 ;
  assign y15274 = n21130 ;
  assign y15275 = ~n21132 ;
  assign y15276 = n21138 ;
  assign y15277 = ~1'b0 ;
  assign y15278 = ~1'b0 ;
  assign y15279 = ~n21139 ;
  assign y15280 = ~n21141 ;
  assign y15281 = ~n21143 ;
  assign y15282 = n21144 ;
  assign y15283 = n19347 ;
  assign y15284 = ~1'b0 ;
  assign y15285 = n21145 ;
  assign y15286 = ~1'b0 ;
  assign y15287 = n21146 ;
  assign y15288 = ~1'b0 ;
  assign y15289 = ~1'b0 ;
  assign y15290 = ~1'b0 ;
  assign y15291 = ~1'b0 ;
  assign y15292 = 1'b0 ;
  assign y15293 = ~n21148 ;
  assign y15294 = 1'b0 ;
  assign y15295 = n21149 ;
  assign y15296 = n21153 ;
  assign y15297 = ~n21156 ;
  assign y15298 = ~1'b0 ;
  assign y15299 = ~1'b0 ;
  assign y15300 = ~n21162 ;
  assign y15301 = 1'b0 ;
  assign y15302 = ~1'b0 ;
  assign y15303 = ~n10141 ;
  assign y15304 = ~1'b0 ;
  assign y15305 = n21169 ;
  assign y15306 = ~1'b0 ;
  assign y15307 = ~n21170 ;
  assign y15308 = 1'b0 ;
  assign y15309 = ~n21173 ;
  assign y15310 = ~n21174 ;
  assign y15311 = ~1'b0 ;
  assign y15312 = ~1'b0 ;
  assign y15313 = ~n21175 ;
  assign y15314 = n21189 ;
  assign y15315 = n21195 ;
  assign y15316 = ~1'b0 ;
  assign y15317 = 1'b0 ;
  assign y15318 = n9758 ;
  assign y15319 = ~1'b0 ;
  assign y15320 = ~1'b0 ;
  assign y15321 = ~1'b0 ;
  assign y15322 = n21196 ;
  assign y15323 = ~1'b0 ;
  assign y15324 = n21198 ;
  assign y15325 = ~1'b0 ;
  assign y15326 = ~1'b0 ;
  assign y15327 = ~n21201 ;
  assign y15328 = ~1'b0 ;
  assign y15329 = ~n11849 ;
  assign y15330 = ~n21202 ;
  assign y15331 = ~1'b0 ;
  assign y15332 = ~1'b0 ;
  assign y15333 = ~n2209 ;
  assign y15334 = ~1'b0 ;
  assign y15335 = ~n37 ;
  assign y15336 = ~1'b0 ;
  assign y15337 = ~n21207 ;
  assign y15338 = ~1'b0 ;
  assign y15339 = n4714 ;
  assign y15340 = n5554 ;
  assign y15341 = ~1'b0 ;
  assign y15342 = n21208 ;
  assign y15343 = ~1'b0 ;
  assign y15344 = n21209 ;
  assign y15345 = n21211 ;
  assign y15346 = n21216 ;
  assign y15347 = n21220 ;
  assign y15348 = ~n21222 ;
  assign y15349 = ~n21223 ;
  assign y15350 = ~1'b0 ;
  assign y15351 = n21224 ;
  assign y15352 = ~n21227 ;
  assign y15353 = n21231 ;
  assign y15354 = ~1'b0 ;
  assign y15355 = n21232 ;
  assign y15356 = ~n5643 ;
  assign y15357 = ~n21234 ;
  assign y15358 = ~1'b0 ;
  assign y15359 = n1323 ;
  assign y15360 = n21241 ;
  assign y15361 = ~n21242 ;
  assign y15362 = n21243 ;
  assign y15363 = ~1'b0 ;
  assign y15364 = n21244 ;
  assign y15365 = ~1'b0 ;
  assign y15366 = ~n13800 ;
  assign y15367 = ~n21245 ;
  assign y15368 = n21248 ;
  assign y15369 = n13898 ;
  assign y15370 = ~n21250 ;
  assign y15371 = n21252 ;
  assign y15372 = ~n21254 ;
  assign y15373 = ~1'b0 ;
  assign y15374 = n18365 ;
  assign y15375 = n21255 ;
  assign y15376 = ~n21258 ;
  assign y15377 = n21272 ;
  assign y15378 = n21273 ;
  assign y15379 = n21280 ;
  assign y15380 = ~n4700 ;
  assign y15381 = ~1'b0 ;
  assign y15382 = ~n21281 ;
  assign y15383 = ~n10658 ;
  assign y15384 = n21283 ;
  assign y15385 = ~1'b0 ;
  assign y15386 = ~n21284 ;
  assign y15387 = ~n21286 ;
  assign y15388 = ~n21288 ;
  assign y15389 = ~n21289 ;
  assign y15390 = ~n21290 ;
  assign y15391 = n20492 ;
  assign y15392 = n21292 ;
  assign y15393 = ~1'b0 ;
  assign y15394 = ~n8067 ;
  assign y15395 = n21298 ;
  assign y15396 = ~1'b0 ;
  assign y15397 = 1'b0 ;
  assign y15398 = n21300 ;
  assign y15399 = ~n21320 ;
  assign y15400 = ~n9060 ;
  assign y15401 = ~1'b0 ;
  assign y15402 = ~1'b0 ;
  assign y15403 = n21322 ;
  assign y15404 = 1'b0 ;
  assign y15405 = n21328 ;
  assign y15406 = ~n21329 ;
  assign y15407 = n21331 ;
  assign y15408 = ~1'b0 ;
  assign y15409 = ~1'b0 ;
  assign y15410 = n21335 ;
  assign y15411 = n21342 ;
  assign y15412 = ~n21346 ;
  assign y15413 = ~n21350 ;
  assign y15414 = ~1'b0 ;
  assign y15415 = ~1'b0 ;
  assign y15416 = ~1'b0 ;
  assign y15417 = n21355 ;
  assign y15418 = ~1'b0 ;
  assign y15419 = ~n21358 ;
  assign y15420 = ~1'b0 ;
  assign y15421 = ~1'b0 ;
  assign y15422 = ~1'b0 ;
  assign y15423 = n9898 ;
  assign y15424 = ~1'b0 ;
  assign y15425 = ~1'b0 ;
  assign y15426 = ~n21359 ;
  assign y15427 = ~n21361 ;
  assign y15428 = ~1'b0 ;
  assign y15429 = ~1'b0 ;
  assign y15430 = ~1'b0 ;
  assign y15431 = n21362 ;
  assign y15432 = n21366 ;
  assign y15433 = n21368 ;
  assign y15434 = n21370 ;
  assign y15435 = ~n18355 ;
  assign y15436 = ~n21371 ;
  assign y15437 = ~n21372 ;
  assign y15438 = n9180 ;
  assign y15439 = ~1'b0 ;
  assign y15440 = n21375 ;
  assign y15441 = ~n21378 ;
  assign y15442 = ~n21380 ;
  assign y15443 = ~n21382 ;
  assign y15444 = ~1'b0 ;
  assign y15445 = ~n21384 ;
  assign y15446 = ~n21385 ;
  assign y15447 = n21387 ;
  assign y15448 = ~n21391 ;
  assign y15449 = ~n21397 ;
  assign y15450 = n21401 ;
  assign y15451 = 1'b0 ;
  assign y15452 = n21402 ;
  assign y15453 = ~n21405 ;
  assign y15454 = ~n21409 ;
  assign y15455 = ~n21410 ;
  assign y15456 = ~n21412 ;
  assign y15457 = ~1'b0 ;
  assign y15458 = n21414 ;
  assign y15459 = n11673 ;
  assign y15460 = ~1'b0 ;
  assign y15461 = ~n21416 ;
  assign y15462 = n21418 ;
  assign y15463 = n21424 ;
  assign y15464 = ~1'b0 ;
  assign y15465 = ~1'b0 ;
  assign y15466 = ~1'b0 ;
  assign y15467 = ~n21426 ;
  assign y15468 = ~1'b0 ;
  assign y15469 = n21427 ;
  assign y15470 = ~n21432 ;
  assign y15471 = ~1'b0 ;
  assign y15472 = ~n21435 ;
  assign y15473 = ~1'b0 ;
  assign y15474 = n1480 ;
  assign y15475 = ~1'b0 ;
  assign y15476 = 1'b0 ;
  assign y15477 = ~n21437 ;
  assign y15478 = ~n21446 ;
  assign y15479 = n21447 ;
  assign y15480 = 1'b0 ;
  assign y15481 = ~1'b0 ;
  assign y15482 = ~n21449 ;
  assign y15483 = ~n21450 ;
  assign y15484 = n17914 ;
  assign y15485 = ~1'b0 ;
  assign y15486 = ~1'b0 ;
  assign y15487 = ~n21452 ;
  assign y15488 = ~n21455 ;
  assign y15489 = ~1'b0 ;
  assign y15490 = n21457 ;
  assign y15491 = ~n21460 ;
  assign y15492 = ~n21467 ;
  assign y15493 = ~n21468 ;
  assign y15494 = ~1'b0 ;
  assign y15495 = ~n21477 ;
  assign y15496 = n21479 ;
  assign y15497 = ~1'b0 ;
  assign y15498 = ~1'b0 ;
  assign y15499 = ~1'b0 ;
  assign y15500 = n21480 ;
  assign y15501 = n21482 ;
  assign y15502 = ~1'b0 ;
  assign y15503 = n21484 ;
  assign y15504 = n21485 ;
  assign y15505 = ~n21487 ;
  assign y15506 = n21491 ;
  assign y15507 = ~1'b0 ;
  assign y15508 = n21500 ;
  assign y15509 = ~n21502 ;
  assign y15510 = ~n15441 ;
  assign y15511 = ~n165 ;
  assign y15512 = ~1'b0 ;
  assign y15513 = ~n21504 ;
  assign y15514 = n21505 ;
  assign y15515 = ~n20115 ;
  assign y15516 = 1'b0 ;
  assign y15517 = n21506 ;
  assign y15518 = ~n21507 ;
  assign y15519 = n21508 ;
  assign y15520 = ~1'b0 ;
  assign y15521 = ~1'b0 ;
  assign y15522 = n21511 ;
  assign y15523 = ~1'b0 ;
  assign y15524 = ~1'b0 ;
  assign y15525 = ~n21512 ;
  assign y15526 = 1'b0 ;
  assign y15527 = n21513 ;
  assign y15528 = n21517 ;
  assign y15529 = ~n21519 ;
  assign y15530 = ~n21522 ;
  assign y15531 = ~n21524 ;
  assign y15532 = ~n21525 ;
  assign y15533 = ~n21526 ;
  assign y15534 = ~1'b0 ;
  assign y15535 = n21527 ;
  assign y15536 = ~1'b0 ;
  assign y15537 = n21531 ;
  assign y15538 = ~n21538 ;
  assign y15539 = 1'b0 ;
  assign y15540 = ~n21542 ;
  assign y15541 = ~1'b0 ;
  assign y15542 = ~1'b0 ;
  assign y15543 = ~1'b0 ;
  assign y15544 = 1'b0 ;
  assign y15545 = ~1'b0 ;
  assign y15546 = ~1'b0 ;
  assign y15547 = n4303 ;
  assign y15548 = n21543 ;
  assign y15549 = n8622 ;
  assign y15550 = ~n21544 ;
  assign y15551 = ~1'b0 ;
  assign y15552 = ~1'b0 ;
  assign y15553 = n19402 ;
  assign y15554 = ~n21545 ;
  assign y15555 = n21546 ;
  assign y15556 = n21547 ;
  assign y15557 = ~1'b0 ;
  assign y15558 = ~n688 ;
  assign y15559 = ~1'b0 ;
  assign y15560 = ~1'b0 ;
  assign y15561 = n21554 ;
  assign y15562 = ~1'b0 ;
  assign y15563 = n21556 ;
  assign y15564 = n21557 ;
  assign y15565 = n21560 ;
  assign y15566 = n21561 ;
  assign y15567 = ~n21562 ;
  assign y15568 = ~n21567 ;
  assign y15569 = 1'b0 ;
  assign y15570 = n21568 ;
  assign y15571 = ~n21569 ;
  assign y15572 = ~1'b0 ;
  assign y15573 = ~n21574 ;
  assign y15574 = n21583 ;
  assign y15575 = ~n21589 ;
  assign y15576 = 1'b0 ;
  assign y15577 = ~1'b0 ;
  assign y15578 = ~n21590 ;
  assign y15579 = ~1'b0 ;
  assign y15580 = ~1'b0 ;
  assign y15581 = ~1'b0 ;
  assign y15582 = n21591 ;
  assign y15583 = ~n21594 ;
  assign y15584 = 1'b0 ;
  assign y15585 = ~1'b0 ;
  assign y15586 = ~n21603 ;
  assign y15587 = ~n423 ;
  assign y15588 = ~1'b0 ;
  assign y15589 = ~n21605 ;
  assign y15590 = ~n21607 ;
  assign y15591 = ~n21609 ;
  assign y15592 = ~1'b0 ;
  assign y15593 = 1'b0 ;
  assign y15594 = ~n21610 ;
  assign y15595 = ~n21611 ;
  assign y15596 = ~1'b0 ;
  assign y15597 = ~1'b0 ;
  assign y15598 = ~n21612 ;
  assign y15599 = ~1'b0 ;
  assign y15600 = n21613 ;
  assign y15601 = ~n7609 ;
  assign y15602 = n21619 ;
  assign y15603 = n21622 ;
  assign y15604 = n21625 ;
  assign y15605 = 1'b0 ;
  assign y15606 = n21628 ;
  assign y15607 = ~n21629 ;
  assign y15608 = 1'b0 ;
  assign y15609 = n21631 ;
  assign y15610 = n21632 ;
  assign y15611 = n21635 ;
  assign y15612 = ~n21636 ;
  assign y15613 = ~n9776 ;
  assign y15614 = ~n13461 ;
  assign y15615 = ~n21638 ;
  assign y15616 = n21640 ;
  assign y15617 = ~1'b0 ;
  assign y15618 = n21641 ;
  assign y15619 = 1'b0 ;
  assign y15620 = ~n21642 ;
  assign y15621 = n21644 ;
  assign y15622 = ~n21647 ;
  assign y15623 = ~n21649 ;
  assign y15624 = ~n21650 ;
  assign y15625 = ~n21653 ;
  assign y15626 = n21654 ;
  assign y15627 = ~1'b0 ;
  assign y15628 = n17623 ;
  assign y15629 = ~1'b0 ;
  assign y15630 = ~1'b0 ;
  assign y15631 = ~1'b0 ;
  assign y15632 = ~n21655 ;
  assign y15633 = ~1'b0 ;
  assign y15634 = ~n21656 ;
  assign y15635 = ~n616 ;
  assign y15636 = ~n21657 ;
  assign y15637 = ~n10427 ;
  assign y15638 = ~1'b0 ;
  assign y15639 = ~n21658 ;
  assign y15640 = n1959 ;
  assign y15641 = ~n21660 ;
  assign y15642 = n21667 ;
  assign y15643 = n21669 ;
  assign y15644 = n21672 ;
  assign y15645 = ~n21674 ;
  assign y15646 = n15668 ;
  assign y15647 = n21677 ;
  assign y15648 = ~n21680 ;
  assign y15649 = ~n21681 ;
  assign y15650 = n21683 ;
  assign y15651 = ~1'b0 ;
  assign y15652 = n21684 ;
  assign y15653 = ~n21685 ;
  assign y15654 = n21686 ;
  assign y15655 = ~n21714 ;
  assign y15656 = ~1'b0 ;
  assign y15657 = ~1'b0 ;
  assign y15658 = ~1'b0 ;
  assign y15659 = ~n21718 ;
  assign y15660 = n21719 ;
  assign y15661 = ~1'b0 ;
  assign y15662 = ~n21720 ;
  assign y15663 = ~n21721 ;
  assign y15664 = ~n5334 ;
  assign y15665 = n3803 ;
  assign y15666 = ~1'b0 ;
  assign y15667 = ~n21724 ;
  assign y15668 = n21727 ;
  assign y15669 = ~n21728 ;
  assign y15670 = ~n21729 ;
  assign y15671 = ~1'b0 ;
  assign y15672 = ~1'b0 ;
  assign y15673 = 1'b0 ;
  assign y15674 = n21730 ;
  assign y15675 = ~n21731 ;
  assign y15676 = ~n15324 ;
  assign y15677 = ~1'b0 ;
  assign y15678 = ~1'b0 ;
  assign y15679 = ~1'b0 ;
  assign y15680 = n21733 ;
  assign y15681 = ~1'b0 ;
  assign y15682 = ~1'b0 ;
  assign y15683 = n21734 ;
  assign y15684 = ~1'b0 ;
  assign y15685 = ~n6674 ;
  assign y15686 = ~1'b0 ;
  assign y15687 = n21735 ;
  assign y15688 = ~n21737 ;
  assign y15689 = n21742 ;
  assign y15690 = ~n21743 ;
  assign y15691 = n21746 ;
  assign y15692 = n21751 ;
  assign y15693 = 1'b0 ;
  assign y15694 = ~1'b0 ;
  assign y15695 = ~1'b0 ;
  assign y15696 = ~1'b0 ;
  assign y15697 = ~n21753 ;
  assign y15698 = ~n21754 ;
  assign y15699 = ~1'b0 ;
  assign y15700 = ~n21756 ;
  assign y15701 = n21757 ;
  assign y15702 = n21762 ;
  assign y15703 = ~1'b0 ;
  assign y15704 = n21765 ;
  assign y15705 = ~1'b0 ;
  assign y15706 = ~1'b0 ;
  assign y15707 = ~n21769 ;
  assign y15708 = ~n21778 ;
  assign y15709 = n21781 ;
  assign y15710 = n16120 ;
  assign y15711 = ~n21783 ;
  assign y15712 = 1'b0 ;
  assign y15713 = ~n13966 ;
  assign y15714 = n21785 ;
  assign y15715 = ~1'b0 ;
  assign y15716 = ~n21787 ;
  assign y15717 = ~n21791 ;
  assign y15718 = ~1'b0 ;
  assign y15719 = n21793 ;
  assign y15720 = ~1'b0 ;
  assign y15721 = ~1'b0 ;
  assign y15722 = ~n21798 ;
  assign y15723 = ~1'b0 ;
  assign y15724 = ~1'b0 ;
  assign y15725 = ~1'b0 ;
  assign y15726 = ~1'b0 ;
  assign y15727 = ~1'b0 ;
  assign y15728 = ~1'b0 ;
  assign y15729 = n21799 ;
  assign y15730 = ~n21800 ;
  assign y15731 = ~1'b0 ;
  assign y15732 = ~1'b0 ;
  assign y15733 = ~n21804 ;
  assign y15734 = n21805 ;
  assign y15735 = n21806 ;
  assign y15736 = ~1'b0 ;
  assign y15737 = ~n21807 ;
  assign y15738 = ~1'b0 ;
  assign y15739 = n21808 ;
  assign y15740 = n21809 ;
  assign y15741 = ~1'b0 ;
  assign y15742 = ~1'b0 ;
  assign y15743 = ~n9565 ;
  assign y15744 = 1'b0 ;
  assign y15745 = ~n21812 ;
  assign y15746 = ~n73 ;
  assign y15747 = n8798 ;
  assign y15748 = n21823 ;
  assign y15749 = ~1'b0 ;
  assign y15750 = n3641 ;
  assign y15751 = n21829 ;
  assign y15752 = n21831 ;
  assign y15753 = ~n21833 ;
  assign y15754 = ~1'b0 ;
  assign y15755 = ~1'b0 ;
  assign y15756 = ~1'b0 ;
  assign y15757 = ~n21834 ;
  assign y15758 = ~n21837 ;
  assign y15759 = n21841 ;
  assign y15760 = ~1'b0 ;
  assign y15761 = ~1'b0 ;
  assign y15762 = ~n21844 ;
  assign y15763 = ~n21850 ;
  assign y15764 = ~1'b0 ;
  assign y15765 = 1'b0 ;
  assign y15766 = ~n15400 ;
  assign y15767 = n21858 ;
  assign y15768 = n21859 ;
  assign y15769 = n2150 ;
  assign y15770 = ~n21864 ;
  assign y15771 = ~1'b0 ;
  assign y15772 = ~n21866 ;
  assign y15773 = ~1'b0 ;
  assign y15774 = ~1'b0 ;
  assign y15775 = n6107 ;
  assign y15776 = 1'b0 ;
  assign y15777 = ~n21868 ;
  assign y15778 = ~n21870 ;
  assign y15779 = ~n6286 ;
  assign y15780 = n21872 ;
  assign y15781 = n21874 ;
  assign y15782 = ~n4964 ;
  assign y15783 = ~1'b0 ;
  assign y15784 = ~n21876 ;
  assign y15785 = ~1'b0 ;
  assign y15786 = ~1'b0 ;
  assign y15787 = n444 ;
  assign y15788 = n21877 ;
  assign y15789 = ~n8979 ;
  assign y15790 = ~n8488 ;
  assign y15791 = ~n13861 ;
  assign y15792 = ~1'b0 ;
  assign y15793 = ~n21880 ;
  assign y15794 = ~n21882 ;
  assign y15795 = ~n21886 ;
  assign y15796 = n21888 ;
  assign y15797 = ~n14515 ;
  assign y15798 = ~1'b0 ;
  assign y15799 = ~n21890 ;
  assign y15800 = n21892 ;
  assign y15801 = ~1'b0 ;
  assign y15802 = ~1'b0 ;
  assign y15803 = ~1'b0 ;
  assign y15804 = ~n21936 ;
  assign y15805 = ~1'b0 ;
  assign y15806 = 1'b0 ;
  assign y15807 = n21938 ;
  assign y15808 = ~n21941 ;
  assign y15809 = ~1'b0 ;
  assign y15810 = ~1'b0 ;
  assign y15811 = n21942 ;
  assign y15812 = ~1'b0 ;
  assign y15813 = n21944 ;
  assign y15814 = ~1'b0 ;
  assign y15815 = ~n21945 ;
  assign y15816 = n1650 ;
  assign y15817 = n21947 ;
  assign y15818 = n21950 ;
  assign y15819 = ~n21952 ;
  assign y15820 = ~n21955 ;
  assign y15821 = ~1'b0 ;
  assign y15822 = ~n21956 ;
  assign y15823 = ~1'b0 ;
  assign y15824 = n21958 ;
  assign y15825 = ~1'b0 ;
  assign y15826 = ~1'b0 ;
  assign y15827 = ~1'b0 ;
  assign y15828 = ~n21960 ;
  assign y15829 = n21963 ;
  assign y15830 = ~1'b0 ;
  assign y15831 = n21965 ;
  assign y15832 = ~n21966 ;
  assign y15833 = ~1'b0 ;
  assign y15834 = ~1'b0 ;
  assign y15835 = ~n21969 ;
  assign y15836 = n21973 ;
  assign y15837 = ~n21975 ;
  assign y15838 = ~n13482 ;
  assign y15839 = ~n21976 ;
  assign y15840 = ~n21978 ;
  assign y15841 = ~n2626 ;
  assign y15842 = n17537 ;
  assign y15843 = ~n21979 ;
  assign y15844 = ~1'b0 ;
  assign y15845 = ~n21981 ;
  assign y15846 = ~n21984 ;
  assign y15847 = ~n21986 ;
  assign y15848 = ~n12105 ;
  assign y15849 = ~n21987 ;
  assign y15850 = n21988 ;
  assign y15851 = 1'b0 ;
  assign y15852 = ~n21990 ;
  assign y15853 = ~n21992 ;
  assign y15854 = ~n21996 ;
  assign y15855 = n21997 ;
  assign y15856 = ~n22000 ;
  assign y15857 = ~1'b0 ;
  assign y15858 = ~1'b0 ;
  assign y15859 = ~1'b0 ;
  assign y15860 = ~n22028 ;
  assign y15861 = n22029 ;
  assign y15862 = n22031 ;
  assign y15863 = ~1'b0 ;
  assign y15864 = ~1'b0 ;
  assign y15865 = ~1'b0 ;
  assign y15866 = ~1'b0 ;
  assign y15867 = n22033 ;
  assign y15868 = n14044 ;
  assign y15869 = ~n22034 ;
  assign y15870 = ~n22037 ;
  assign y15871 = ~n22038 ;
  assign y15872 = n22041 ;
  assign y15873 = ~1'b0 ;
  assign y15874 = n22042 ;
  assign y15875 = ~n22044 ;
  assign y15876 = ~n22045 ;
  assign y15877 = ~1'b0 ;
  assign y15878 = ~n22046 ;
  assign y15879 = ~n22047 ;
  assign y15880 = ~n22048 ;
  assign y15881 = ~n22049 ;
  assign y15882 = 1'b0 ;
  assign y15883 = ~n22050 ;
  assign y15884 = ~1'b0 ;
  assign y15885 = n22052 ;
  assign y15886 = n8312 ;
  assign y15887 = ~n15092 ;
  assign y15888 = ~1'b0 ;
  assign y15889 = n22053 ;
  assign y15890 = ~1'b0 ;
  assign y15891 = ~n16853 ;
  assign y15892 = ~n4883 ;
  assign y15893 = n22061 ;
  assign y15894 = ~n7610 ;
  assign y15895 = n3968 ;
  assign y15896 = n22063 ;
  assign y15897 = n13028 ;
  assign y15898 = n19333 ;
  assign y15899 = ~1'b0 ;
  assign y15900 = n22065 ;
  assign y15901 = ~1'b0 ;
  assign y15902 = n22066 ;
  assign y15903 = ~1'b0 ;
  assign y15904 = ~1'b0 ;
  assign y15905 = ~1'b0 ;
  assign y15906 = n22068 ;
  assign y15907 = ~1'b0 ;
  assign y15908 = ~1'b0 ;
  assign y15909 = ~n22074 ;
  assign y15910 = n22078 ;
  assign y15911 = n22079 ;
  assign y15912 = ~1'b0 ;
  assign y15913 = ~1'b0 ;
  assign y15914 = n22080 ;
  assign y15915 = ~1'b0 ;
  assign y15916 = ~n216 ;
  assign y15917 = ~1'b0 ;
  assign y15918 = ~1'b0 ;
  assign y15919 = ~n22081 ;
  assign y15920 = ~n22084 ;
  assign y15921 = 1'b0 ;
  assign y15922 = ~1'b0 ;
  assign y15923 = n22086 ;
  assign y15924 = n22092 ;
  assign y15925 = n22094 ;
  assign y15926 = ~1'b0 ;
  assign y15927 = n22098 ;
  assign y15928 = ~n13431 ;
  assign y15929 = n22101 ;
  assign y15930 = n22103 ;
  assign y15931 = ~n22104 ;
  assign y15932 = n20965 ;
  assign y15933 = n22106 ;
  assign y15934 = ~1'b0 ;
  assign y15935 = n22111 ;
  assign y15936 = n21145 ;
  assign y15937 = n22112 ;
  assign y15938 = ~n8648 ;
  assign y15939 = ~1'b0 ;
  assign y15940 = ~1'b0 ;
  assign y15941 = n3636 ;
  assign y15942 = n22114 ;
  assign y15943 = ~1'b0 ;
  assign y15944 = n22115 ;
  assign y15945 = ~n18845 ;
  assign y15946 = ~n22117 ;
  assign y15947 = ~1'b0 ;
  assign y15948 = ~1'b0 ;
  assign y15949 = ~n22118 ;
  assign y15950 = ~n22122 ;
  assign y15951 = ~n22124 ;
  assign y15952 = ~n22126 ;
  assign y15953 = ~n22129 ;
  assign y15954 = ~1'b0 ;
  assign y15955 = ~n22130 ;
  assign y15956 = ~1'b0 ;
  assign y15957 = n8946 ;
  assign y15958 = ~n22131 ;
  assign y15959 = ~n22133 ;
  assign y15960 = n22140 ;
  assign y15961 = n22141 ;
  assign y15962 = n13579 ;
  assign y15963 = 1'b0 ;
  assign y15964 = ~1'b0 ;
  assign y15965 = n12341 ;
  assign y15966 = ~1'b0 ;
  assign y15967 = n22143 ;
  assign y15968 = ~1'b0 ;
  assign y15969 = ~1'b0 ;
  assign y15970 = ~1'b0 ;
  assign y15971 = ~1'b0 ;
  assign y15972 = ~1'b0 ;
  assign y15973 = n22144 ;
  assign y15974 = n22145 ;
  assign y15975 = 1'b0 ;
  assign y15976 = n22147 ;
  assign y15977 = ~1'b0 ;
  assign y15978 = ~n22150 ;
  assign y15979 = n22156 ;
  assign y15980 = ~1'b0 ;
  assign y15981 = n22159 ;
  assign y15982 = n22160 ;
  assign y15983 = ~n10920 ;
  assign y15984 = ~n22163 ;
  assign y15985 = ~n22164 ;
  assign y15986 = ~n22166 ;
  assign y15987 = n22169 ;
  assign y15988 = 1'b0 ;
  assign y15989 = n22170 ;
  assign y15990 = n22173 ;
  assign y15991 = ~1'b0 ;
  assign y15992 = ~n22177 ;
  assign y15993 = ~1'b0 ;
  assign y15994 = ~n22179 ;
  assign y15995 = ~1'b0 ;
  assign y15996 = ~n11472 ;
  assign y15997 = ~1'b0 ;
  assign y15998 = n22181 ;
  assign y15999 = n22182 ;
  assign y16000 = n22183 ;
  assign y16001 = ~n22187 ;
  assign y16002 = ~1'b0 ;
  assign y16003 = ~1'b0 ;
  assign y16004 = 1'b0 ;
  assign y16005 = ~n22191 ;
  assign y16006 = ~n22192 ;
  assign y16007 = ~1'b0 ;
  assign y16008 = ~1'b0 ;
  assign y16009 = ~1'b0 ;
  assign y16010 = ~1'b0 ;
  assign y16011 = n1155 ;
  assign y16012 = ~1'b0 ;
  assign y16013 = n22193 ;
  assign y16014 = ~n22198 ;
  assign y16015 = n22203 ;
  assign y16016 = ~n9088 ;
  assign y16017 = n22205 ;
  assign y16018 = 1'b0 ;
  assign y16019 = n22206 ;
  assign y16020 = ~n22207 ;
  assign y16021 = ~n22208 ;
  assign y16022 = n22209 ;
  assign y16023 = n2141 ;
  assign y16024 = ~1'b0 ;
  assign y16025 = ~1'b0 ;
  assign y16026 = n22210 ;
  assign y16027 = ~1'b0 ;
  assign y16028 = n8309 ;
  assign y16029 = ~n22211 ;
  assign y16030 = n22216 ;
  assign y16031 = ~1'b0 ;
  assign y16032 = n22217 ;
  assign y16033 = ~1'b0 ;
  assign y16034 = ~n22218 ;
  assign y16035 = ~1'b0 ;
  assign y16036 = n22219 ;
  assign y16037 = ~1'b0 ;
  assign y16038 = ~1'b0 ;
  assign y16039 = ~1'b0 ;
  assign y16040 = n22221 ;
  assign y16041 = n22227 ;
  assign y16042 = ~1'b0 ;
  assign y16043 = n22229 ;
  assign y16044 = 1'b0 ;
  assign y16045 = ~1'b0 ;
  assign y16046 = ~n22236 ;
  assign y16047 = n22237 ;
  assign y16048 = ~n22240 ;
  assign y16049 = 1'b0 ;
  assign y16050 = ~n22242 ;
  assign y16051 = ~1'b0 ;
  assign y16052 = ~1'b0 ;
  assign y16053 = ~n22246 ;
  assign y16054 = n22249 ;
  assign y16055 = ~n22251 ;
  assign y16056 = ~1'b0 ;
  assign y16057 = ~n3672 ;
  assign y16058 = ~n22252 ;
  assign y16059 = ~n22253 ;
  assign y16060 = ~1'b0 ;
  assign y16061 = n22254 ;
  assign y16062 = n22256 ;
  assign y16063 = 1'b0 ;
  assign y16064 = n22257 ;
  assign y16065 = ~n22263 ;
  assign y16066 = ~1'b0 ;
  assign y16067 = n22267 ;
  assign y16068 = n22270 ;
  assign y16069 = ~n22271 ;
  assign y16070 = n22274 ;
  assign y16071 = ~n22278 ;
  assign y16072 = n22279 ;
  assign y16073 = ~n22281 ;
  assign y16074 = ~1'b0 ;
  assign y16075 = ~1'b0 ;
  assign y16076 = ~1'b0 ;
  assign y16077 = n18267 ;
  assign y16078 = n22287 ;
  assign y16079 = n22288 ;
  assign y16080 = ~n22290 ;
  assign y16081 = n22293 ;
  assign y16082 = ~1'b0 ;
  assign y16083 = ~n22294 ;
  assign y16084 = ~n22295 ;
  assign y16085 = ~1'b0 ;
  assign y16086 = ~n22299 ;
  assign y16087 = n22300 ;
  assign y16088 = n22301 ;
  assign y16089 = 1'b0 ;
  assign y16090 = n8401 ;
  assign y16091 = ~1'b0 ;
  assign y16092 = ~1'b0 ;
  assign y16093 = ~1'b0 ;
  assign y16094 = ~n22303 ;
  assign y16095 = ~n22307 ;
  assign y16096 = ~1'b0 ;
  assign y16097 = ~1'b0 ;
  assign y16098 = ~1'b0 ;
  assign y16099 = 1'b0 ;
  assign y16100 = n22308 ;
  assign y16101 = ~1'b0 ;
  assign y16102 = ~1'b0 ;
  assign y16103 = n22309 ;
  assign y16104 = ~1'b0 ;
  assign y16105 = ~n12565 ;
  assign y16106 = ~n22311 ;
  assign y16107 = ~1'b0 ;
  assign y16108 = n22312 ;
  assign y16109 = n22313 ;
  assign y16110 = n22314 ;
  assign y16111 = ~1'b0 ;
  assign y16112 = ~1'b0 ;
  assign y16113 = ~1'b0 ;
  assign y16114 = ~n22316 ;
  assign y16115 = n22317 ;
  assign y16116 = ~n22328 ;
  assign y16117 = ~1'b0 ;
  assign y16118 = ~n22331 ;
  assign y16119 = ~1'b0 ;
  assign y16120 = ~n22334 ;
  assign y16121 = n22337 ;
  assign y16122 = ~1'b0 ;
  assign y16123 = ~1'b0 ;
  assign y16124 = ~n22339 ;
  assign y16125 = n22340 ;
  assign y16126 = ~1'b0 ;
  assign y16127 = n22342 ;
  assign y16128 = ~1'b0 ;
  assign y16129 = ~1'b0 ;
  assign y16130 = n22346 ;
  assign y16131 = n22349 ;
  assign y16132 = ~1'b0 ;
  assign y16133 = n22357 ;
  assign y16134 = ~n22360 ;
  assign y16135 = n22362 ;
  assign y16136 = ~n17256 ;
  assign y16137 = n22365 ;
  assign y16138 = ~1'b0 ;
  assign y16139 = n22367 ;
  assign y16140 = n14254 ;
  assign y16141 = ~1'b0 ;
  assign y16142 = ~1'b0 ;
  assign y16143 = n4361 ;
  assign y16144 = ~1'b0 ;
  assign y16145 = ~n22370 ;
  assign y16146 = ~n460 ;
  assign y16147 = ~n22373 ;
  assign y16148 = ~n4851 ;
  assign y16149 = n22377 ;
  assign y16150 = ~1'b0 ;
  assign y16151 = n22378 ;
  assign y16152 = ~n22379 ;
  assign y16153 = ~1'b0 ;
  assign y16154 = n22383 ;
  assign y16155 = ~1'b0 ;
  assign y16156 = n22384 ;
  assign y16157 = n22385 ;
  assign y16158 = ~1'b0 ;
  assign y16159 = ~1'b0 ;
  assign y16160 = ~1'b0 ;
  assign y16161 = 1'b0 ;
  assign y16162 = ~n22386 ;
  assign y16163 = ~1'b0 ;
  assign y16164 = ~1'b0 ;
  assign y16165 = ~n22387 ;
  assign y16166 = n22390 ;
  assign y16167 = n7767 ;
  assign y16168 = ~1'b0 ;
  assign y16169 = n22391 ;
  assign y16170 = n22392 ;
  assign y16171 = ~1'b0 ;
  assign y16172 = 1'b0 ;
  assign y16173 = ~1'b0 ;
  assign y16174 = n22398 ;
  assign y16175 = ~n22403 ;
  assign y16176 = n22404 ;
  assign y16177 = ~1'b0 ;
  assign y16178 = n22405 ;
  assign y16179 = ~n22411 ;
  assign y16180 = 1'b0 ;
  assign y16181 = ~1'b0 ;
  assign y16182 = n22415 ;
  assign y16183 = ~1'b0 ;
  assign y16184 = n22416 ;
  assign y16185 = ~n22418 ;
  assign y16186 = ~1'b0 ;
  assign y16187 = n16533 ;
  assign y16188 = ~n194 ;
  assign y16189 = ~1'b0 ;
  assign y16190 = 1'b0 ;
  assign y16191 = n22419 ;
  assign y16192 = n22420 ;
  assign y16193 = ~n22422 ;
  assign y16194 = ~1'b0 ;
  assign y16195 = n22425 ;
  assign y16196 = ~1'b0 ;
  assign y16197 = n22427 ;
  assign y16198 = 1'b0 ;
  assign y16199 = n22429 ;
  assign y16200 = 1'b0 ;
  assign y16201 = ~1'b0 ;
  assign y16202 = n22431 ;
  assign y16203 = ~n22433 ;
  assign y16204 = n3586 ;
  assign y16205 = n22434 ;
  assign y16206 = ~1'b0 ;
  assign y16207 = ~1'b0 ;
  assign y16208 = ~1'b0 ;
  assign y16209 = ~n22438 ;
  assign y16210 = ~1'b0 ;
  assign y16211 = ~1'b0 ;
  assign y16212 = ~1'b0 ;
  assign y16213 = n133 ;
  assign y16214 = ~1'b0 ;
  assign y16215 = ~n22439 ;
  assign y16216 = ~n22442 ;
  assign y16217 = ~1'b0 ;
  assign y16218 = ~n22445 ;
  assign y16219 = ~n22451 ;
  assign y16220 = ~1'b0 ;
  assign y16221 = n22452 ;
  assign y16222 = ~n22455 ;
  assign y16223 = ~n22460 ;
  assign y16224 = ~n22463 ;
  assign y16225 = ~n22465 ;
  assign y16226 = ~n9281 ;
  assign y16227 = n22466 ;
  assign y16228 = ~1'b0 ;
  assign y16229 = ~n22470 ;
  assign y16230 = ~n3940 ;
  assign y16231 = ~n22471 ;
  assign y16232 = ~n22474 ;
  assign y16233 = ~1'b0 ;
  assign y16234 = ~n22475 ;
  assign y16235 = ~1'b0 ;
  assign y16236 = ~1'b0 ;
  assign y16237 = n14571 ;
  assign y16238 = n22476 ;
  assign y16239 = n22480 ;
  assign y16240 = n22482 ;
  assign y16241 = ~1'b0 ;
  assign y16242 = ~n22483 ;
  assign y16243 = ~1'b0 ;
  assign y16244 = n22489 ;
  assign y16245 = ~n22491 ;
  assign y16246 = ~n22492 ;
  assign y16247 = ~1'b0 ;
  assign y16248 = ~1'b0 ;
  assign y16249 = n22494 ;
  assign y16250 = n22495 ;
  assign y16251 = ~1'b0 ;
  assign y16252 = n22497 ;
  assign y16253 = ~1'b0 ;
  assign y16254 = n22498 ;
  assign y16255 = 1'b0 ;
  assign y16256 = ~1'b0 ;
  assign y16257 = ~n22502 ;
  assign y16258 = ~1'b0 ;
  assign y16259 = ~1'b0 ;
  assign y16260 = n9158 ;
  assign y16261 = ~n22503 ;
  assign y16262 = ~n22504 ;
  assign y16263 = n22507 ;
  assign y16264 = n22508 ;
  assign y16265 = ~n22509 ;
  assign y16266 = ~1'b0 ;
  assign y16267 = ~1'b0 ;
  assign y16268 = ~n22525 ;
  assign y16269 = ~1'b0 ;
  assign y16270 = ~n108 ;
  assign y16271 = ~1'b0 ;
  assign y16272 = ~n22529 ;
  assign y16273 = n9309 ;
  assign y16274 = ~n22530 ;
  assign y16275 = ~1'b0 ;
  assign y16276 = n22532 ;
  assign y16277 = n22534 ;
  assign y16278 = ~n6631 ;
  assign y16279 = n22538 ;
  assign y16280 = ~1'b0 ;
  assign y16281 = n22539 ;
  assign y16282 = ~1'b0 ;
  assign y16283 = ~1'b0 ;
  assign y16284 = ~1'b0 ;
  assign y16285 = ~n22540 ;
  assign y16286 = ~n22542 ;
  assign y16287 = 1'b0 ;
  assign y16288 = ~n22544 ;
  assign y16289 = ~1'b0 ;
  assign y16290 = n5749 ;
  assign y16291 = n22545 ;
  assign y16292 = n22548 ;
  assign y16293 = ~n22563 ;
  assign y16294 = n22564 ;
  assign y16295 = 1'b0 ;
  assign y16296 = n22565 ;
  assign y16297 = ~1'b0 ;
  assign y16298 = ~1'b0 ;
  assign y16299 = n22566 ;
  assign y16300 = ~1'b0 ;
  assign y16301 = ~1'b0 ;
  assign y16302 = ~n22568 ;
  assign y16303 = n22569 ;
  assign y16304 = n18013 ;
  assign y16305 = n1590 ;
  assign y16306 = ~1'b0 ;
  assign y16307 = ~n22570 ;
  assign y16308 = ~n22573 ;
  assign y16309 = n4211 ;
  assign y16310 = ~n22575 ;
  assign y16311 = ~1'b0 ;
  assign y16312 = ~n22576 ;
  assign y16313 = ~1'b0 ;
  assign y16314 = n22579 ;
  assign y16315 = n22580 ;
  assign y16316 = ~n18462 ;
  assign y16317 = n22584 ;
  assign y16318 = ~n22588 ;
  assign y16319 = ~n18172 ;
  assign y16320 = ~1'b0 ;
  assign y16321 = ~n22590 ;
  assign y16322 = ~1'b0 ;
  assign y16323 = ~1'b0 ;
  assign y16324 = ~1'b0 ;
  assign y16325 = n22591 ;
  assign y16326 = ~n18716 ;
  assign y16327 = n6034 ;
  assign y16328 = ~1'b0 ;
  assign y16329 = ~1'b0 ;
  assign y16330 = ~1'b0 ;
  assign y16331 = n22401 ;
  assign y16332 = 1'b0 ;
  assign y16333 = n22592 ;
  assign y16334 = n22595 ;
  assign y16335 = ~n22600 ;
  assign y16336 = ~1'b0 ;
  assign y16337 = n22604 ;
  assign y16338 = ~n22608 ;
  assign y16339 = ~n5005 ;
  assign y16340 = ~n22612 ;
  assign y16341 = n22613 ;
  assign y16342 = n22614 ;
  assign y16343 = ~n22615 ;
  assign y16344 = n22616 ;
  assign y16345 = ~n22619 ;
  assign y16346 = ~n22622 ;
  assign y16347 = ~n8561 ;
  assign y16348 = n22624 ;
  assign y16349 = ~1'b0 ;
  assign y16350 = ~n8409 ;
  assign y16351 = n13782 ;
  assign y16352 = ~1'b0 ;
  assign y16353 = ~n22625 ;
  assign y16354 = ~n22628 ;
  assign y16355 = ~1'b0 ;
  assign y16356 = n22633 ;
  assign y16357 = n22634 ;
  assign y16358 = n11731 ;
  assign y16359 = ~n22635 ;
  assign y16360 = n22641 ;
  assign y16361 = ~1'b0 ;
  assign y16362 = n22644 ;
  assign y16363 = ~n22646 ;
  assign y16364 = ~n22650 ;
  assign y16365 = ~1'b0 ;
  assign y16366 = n22652 ;
  assign y16367 = n22654 ;
  assign y16368 = n22658 ;
  assign y16369 = ~n22570 ;
  assign y16370 = ~1'b0 ;
  assign y16371 = ~n22659 ;
  assign y16372 = n9306 ;
  assign y16373 = n22661 ;
  assign y16374 = ~1'b0 ;
  assign y16375 = ~1'b0 ;
  assign y16376 = n22668 ;
  assign y16377 = ~n22670 ;
  assign y16378 = n22671 ;
  assign y16379 = n22672 ;
  assign y16380 = ~1'b0 ;
  assign y16381 = n22674 ;
  assign y16382 = ~1'b0 ;
  assign y16383 = ~n22676 ;
  assign y16384 = ~1'b0 ;
  assign y16385 = n22677 ;
  assign y16386 = n22681 ;
  assign y16387 = ~1'b0 ;
  assign y16388 = ~1'b0 ;
  assign y16389 = ~n4009 ;
  assign y16390 = ~1'b0 ;
  assign y16391 = n6408 ;
  assign y16392 = ~n22683 ;
  assign y16393 = ~n5532 ;
  assign y16394 = n22685 ;
  assign y16395 = n22686 ;
  assign y16396 = n22688 ;
  assign y16397 = 1'b0 ;
  assign y16398 = n22689 ;
  assign y16399 = n22691 ;
  assign y16400 = ~1'b0 ;
  assign y16401 = ~n22692 ;
  assign y16402 = ~n16689 ;
  assign y16403 = ~n22696 ;
  assign y16404 = ~n22698 ;
  assign y16405 = ~n22704 ;
  assign y16406 = n22705 ;
  assign y16407 = ~n11915 ;
  assign y16408 = n4077 ;
  assign y16409 = n22706 ;
  assign y16410 = 1'b0 ;
  assign y16411 = n12045 ;
  assign y16412 = ~n22708 ;
  assign y16413 = n22712 ;
  assign y16414 = ~1'b0 ;
  assign y16415 = n22714 ;
  assign y16416 = ~n22717 ;
  assign y16417 = ~n22719 ;
  assign y16418 = n22720 ;
  assign y16419 = n22722 ;
  assign y16420 = ~1'b0 ;
  assign y16421 = ~n22726 ;
  assign y16422 = n22728 ;
  assign y16423 = n22730 ;
  assign y16424 = ~1'b0 ;
  assign y16425 = 1'b0 ;
  assign y16426 = ~n22731 ;
  assign y16427 = n22733 ;
  assign y16428 = ~n2593 ;
  assign y16429 = ~1'b0 ;
  assign y16430 = ~n22735 ;
  assign y16431 = ~1'b0 ;
  assign y16432 = ~1'b0 ;
  assign y16433 = ~n22736 ;
  assign y16434 = ~n22737 ;
  assign y16435 = 1'b0 ;
  assign y16436 = ~1'b0 ;
  assign y16437 = n22740 ;
  assign y16438 = n22746 ;
  assign y16439 = ~1'b0 ;
  assign y16440 = n22748 ;
  assign y16441 = n6929 ;
  assign y16442 = n22749 ;
  assign y16443 = ~n22751 ;
  assign y16444 = n22753 ;
  assign y16445 = ~n22754 ;
  assign y16446 = ~1'b0 ;
  assign y16447 = n22756 ;
  assign y16448 = ~1'b0 ;
  assign y16449 = ~n22759 ;
  assign y16450 = ~n22765 ;
  assign y16451 = ~1'b0 ;
  assign y16452 = n22767 ;
  assign y16453 = ~1'b0 ;
  assign y16454 = ~n22768 ;
  assign y16455 = ~1'b0 ;
  assign y16456 = ~1'b0 ;
  assign y16457 = ~n22770 ;
  assign y16458 = ~1'b0 ;
  assign y16459 = ~1'b0 ;
  assign y16460 = ~1'b0 ;
  assign y16461 = n22772 ;
  assign y16462 = ~1'b0 ;
  assign y16463 = ~1'b0 ;
  assign y16464 = ~n11388 ;
  assign y16465 = n22775 ;
  assign y16466 = ~n22779 ;
  assign y16467 = ~n22780 ;
  assign y16468 = 1'b0 ;
  assign y16469 = ~1'b0 ;
  assign y16470 = n22781 ;
  assign y16471 = n19012 ;
  assign y16472 = ~1'b0 ;
  assign y16473 = ~1'b0 ;
  assign y16474 = ~n11131 ;
  assign y16475 = ~1'b0 ;
  assign y16476 = ~1'b0 ;
  assign y16477 = n22782 ;
  assign y16478 = ~n22785 ;
  assign y16479 = ~n22787 ;
  assign y16480 = ~1'b0 ;
  assign y16481 = ~n16541 ;
  assign y16482 = ~n22789 ;
  assign y16483 = ~1'b0 ;
  assign y16484 = ~n22792 ;
  assign y16485 = ~1'b0 ;
  assign y16486 = ~n22795 ;
  assign y16487 = ~1'b0 ;
  assign y16488 = ~1'b0 ;
  assign y16489 = n22797 ;
  assign y16490 = n22804 ;
  assign y16491 = ~n22806 ;
  assign y16492 = ~n22807 ;
  assign y16493 = 1'b0 ;
  assign y16494 = n22809 ;
  assign y16495 = n22811 ;
  assign y16496 = ~1'b0 ;
  assign y16497 = ~n22817 ;
  assign y16498 = n22823 ;
  assign y16499 = n22828 ;
  assign y16500 = ~n22829 ;
  assign y16501 = ~n22831 ;
  assign y16502 = ~n22832 ;
  assign y16503 = n22835 ;
  assign y16504 = n22836 ;
  assign y16505 = ~n22837 ;
  assign y16506 = ~n22838 ;
  assign y16507 = n22845 ;
  assign y16508 = n2910 ;
  assign y16509 = ~1'b0 ;
  assign y16510 = n22849 ;
  assign y16511 = ~1'b0 ;
  assign y16512 = ~n10060 ;
  assign y16513 = n22850 ;
  assign y16514 = ~n22851 ;
  assign y16515 = ~1'b0 ;
  assign y16516 = ~n22853 ;
  assign y16517 = n4247 ;
  assign y16518 = ~n22855 ;
  assign y16519 = ~n22856 ;
  assign y16520 = 1'b0 ;
  assign y16521 = ~1'b0 ;
  assign y16522 = ~1'b0 ;
  assign y16523 = n22857 ;
  assign y16524 = n22859 ;
  assign y16525 = ~n22861 ;
  assign y16526 = ~1'b0 ;
  assign y16527 = ~1'b0 ;
  assign y16528 = ~1'b0 ;
  assign y16529 = 1'b0 ;
  assign y16530 = ~n22864 ;
  assign y16531 = ~n12697 ;
  assign y16532 = n22865 ;
  assign y16533 = ~1'b0 ;
  assign y16534 = n22870 ;
  assign y16535 = ~n22872 ;
  assign y16536 = ~n22873 ;
  assign y16537 = ~1'b0 ;
  assign y16538 = n22874 ;
  assign y16539 = ~1'b0 ;
  assign y16540 = ~n22878 ;
  assign y16541 = ~n22879 ;
  assign y16542 = ~1'b0 ;
  assign y16543 = ~n22882 ;
  assign y16544 = n22885 ;
  assign y16545 = n22887 ;
  assign y16546 = ~n22888 ;
  assign y16547 = ~n22889 ;
  assign y16548 = ~n22892 ;
  assign y16549 = ~1'b0 ;
  assign y16550 = ~1'b0 ;
  assign y16551 = 1'b0 ;
  assign y16552 = ~n22893 ;
  assign y16553 = ~1'b0 ;
  assign y16554 = n22898 ;
  assign y16555 = n22901 ;
  assign y16556 = ~n22903 ;
  assign y16557 = ~n22909 ;
  assign y16558 = ~1'b0 ;
  assign y16559 = n22911 ;
  assign y16560 = n4258 ;
  assign y16561 = n22912 ;
  assign y16562 = n2482 ;
  assign y16563 = ~1'b0 ;
  assign y16564 = ~1'b0 ;
  assign y16565 = ~1'b0 ;
  assign y16566 = ~1'b0 ;
  assign y16567 = ~n22914 ;
  assign y16568 = ~n22915 ;
  assign y16569 = ~n22916 ;
  assign y16570 = n22919 ;
  assign y16571 = ~n22920 ;
  assign y16572 = ~n22922 ;
  assign y16573 = ~n7851 ;
  assign y16574 = n22926 ;
  assign y16575 = ~1'b0 ;
  assign y16576 = ~n22930 ;
  assign y16577 = ~n22932 ;
  assign y16578 = ~1'b0 ;
  assign y16579 = ~1'b0 ;
  assign y16580 = ~n22937 ;
  assign y16581 = ~1'b0 ;
  assign y16582 = ~n22945 ;
  assign y16583 = n22946 ;
  assign y16584 = ~1'b0 ;
  assign y16585 = n22947 ;
  assign y16586 = ~n22954 ;
  assign y16587 = n22955 ;
  assign y16588 = ~1'b0 ;
  assign y16589 = n21023 ;
  assign y16590 = ~n22956 ;
  assign y16591 = ~n22958 ;
  assign y16592 = ~n22960 ;
  assign y16593 = ~n22961 ;
  assign y16594 = ~1'b0 ;
  assign y16595 = ~n22963 ;
  assign y16596 = ~n22965 ;
  assign y16597 = n22967 ;
  assign y16598 = n22969 ;
  assign y16599 = n7210 ;
  assign y16600 = n6846 ;
  assign y16601 = ~n22972 ;
  assign y16602 = 1'b0 ;
  assign y16603 = ~1'b0 ;
  assign y16604 = ~1'b0 ;
  assign y16605 = ~1'b0 ;
  assign y16606 = ~1'b0 ;
  assign y16607 = n22983 ;
  assign y16608 = n6454 ;
  assign y16609 = ~1'b0 ;
  assign y16610 = ~n22984 ;
  assign y16611 = ~1'b0 ;
  assign y16612 = ~1'b0 ;
  assign y16613 = ~1'b0 ;
  assign y16614 = n22988 ;
  assign y16615 = n22989 ;
  assign y16616 = ~1'b0 ;
  assign y16617 = ~1'b0 ;
  assign y16618 = n675 ;
  assign y16619 = n22995 ;
  assign y16620 = ~1'b0 ;
  assign y16621 = ~1'b0 ;
  assign y16622 = ~n22998 ;
  assign y16623 = n294 ;
  assign y16624 = ~n23000 ;
  assign y16625 = n23001 ;
  assign y16626 = ~n23005 ;
  assign y16627 = ~n23006 ;
  assign y16628 = ~1'b0 ;
  assign y16629 = ~1'b0 ;
  assign y16630 = ~1'b0 ;
  assign y16631 = ~1'b0 ;
  assign y16632 = 1'b0 ;
  assign y16633 = ~1'b0 ;
  assign y16634 = n23007 ;
  assign y16635 = ~n23010 ;
  assign y16636 = ~1'b0 ;
  assign y16637 = n527 ;
  assign y16638 = n23014 ;
  assign y16639 = ~1'b0 ;
  assign y16640 = n36 ;
  assign y16641 = ~n4979 ;
  assign y16642 = n23016 ;
  assign y16643 = n23020 ;
  assign y16644 = n23021 ;
  assign y16645 = ~1'b0 ;
  assign y16646 = ~1'b0 ;
  assign y16647 = n23025 ;
  assign y16648 = n23027 ;
  assign y16649 = ~1'b0 ;
  assign y16650 = n23028 ;
  assign y16651 = ~n23029 ;
  assign y16652 = n23030 ;
  assign y16653 = ~1'b0 ;
  assign y16654 = ~n23034 ;
  assign y16655 = ~1'b0 ;
  assign y16656 = ~1'b0 ;
  assign y16657 = ~1'b0 ;
  assign y16658 = 1'b0 ;
  assign y16659 = ~1'b0 ;
  assign y16660 = n23035 ;
  assign y16661 = n23036 ;
  assign y16662 = n23037 ;
  assign y16663 = ~1'b0 ;
  assign y16664 = ~n23038 ;
  assign y16665 = ~n23041 ;
  assign y16666 = ~n23046 ;
  assign y16667 = n23047 ;
  assign y16668 = ~n23049 ;
  assign y16669 = ~1'b0 ;
  assign y16670 = ~n23052 ;
  assign y16671 = n23055 ;
  assign y16672 = ~1'b0 ;
  assign y16673 = ~1'b0 ;
  assign y16674 = n23058 ;
  assign y16675 = ~n14317 ;
  assign y16676 = ~n23059 ;
  assign y16677 = ~1'b0 ;
  assign y16678 = ~1'b0 ;
  assign y16679 = ~1'b0 ;
  assign y16680 = n23062 ;
  assign y16681 = n23065 ;
  assign y16682 = ~n23066 ;
  assign y16683 = ~1'b0 ;
  assign y16684 = ~1'b0 ;
  assign y16685 = ~1'b0 ;
  assign y16686 = ~n23068 ;
  assign y16687 = ~1'b0 ;
  assign y16688 = ~1'b0 ;
  assign y16689 = ~1'b0 ;
  assign y16690 = n23069 ;
  assign y16691 = ~1'b0 ;
  assign y16692 = ~1'b0 ;
  assign y16693 = 1'b0 ;
  assign y16694 = ~n23071 ;
  assign y16695 = ~n2736 ;
  assign y16696 = n23072 ;
  assign y16697 = 1'b0 ;
  assign y16698 = ~1'b0 ;
  assign y16699 = ~n23074 ;
  assign y16700 = ~1'b0 ;
  assign y16701 = ~n23077 ;
  assign y16702 = 1'b0 ;
  assign y16703 = ~1'b0 ;
  assign y16704 = ~n23080 ;
  assign y16705 = n23081 ;
  assign y16706 = ~1'b0 ;
  assign y16707 = n23086 ;
  assign y16708 = 1'b0 ;
  assign y16709 = n23091 ;
  assign y16710 = ~n23093 ;
  assign y16711 = ~1'b0 ;
  assign y16712 = ~n9811 ;
  assign y16713 = ~1'b0 ;
  assign y16714 = ~n6173 ;
  assign y16715 = n23095 ;
  assign y16716 = ~1'b0 ;
  assign y16717 = ~n23103 ;
  assign y16718 = n23109 ;
  assign y16719 = n23111 ;
  assign y16720 = ~1'b0 ;
  assign y16721 = n9372 ;
  assign y16722 = ~1'b0 ;
  assign y16723 = n18923 ;
  assign y16724 = n23113 ;
  assign y16725 = ~n23116 ;
  assign y16726 = n23117 ;
  assign y16727 = ~1'b0 ;
  assign y16728 = ~n23118 ;
  assign y16729 = ~n23119 ;
  assign y16730 = ~n5336 ;
  assign y16731 = ~1'b0 ;
  assign y16732 = ~n23121 ;
  assign y16733 = ~n23137 ;
  assign y16734 = n23143 ;
  assign y16735 = n23145 ;
  assign y16736 = ~n23146 ;
  assign y16737 = ~1'b0 ;
  assign y16738 = ~n23147 ;
  assign y16739 = ~1'b0 ;
  assign y16740 = n23148 ;
  assign y16741 = ~n23152 ;
  assign y16742 = ~n23156 ;
  assign y16743 = ~n23159 ;
  assign y16744 = ~n17145 ;
  assign y16745 = 1'b0 ;
  assign y16746 = ~n2784 ;
  assign y16747 = ~1'b0 ;
  assign y16748 = ~n11542 ;
  assign y16749 = ~n23160 ;
  assign y16750 = ~n23163 ;
  assign y16751 = ~n23164 ;
  assign y16752 = ~n23174 ;
  assign y16753 = ~1'b0 ;
  assign y16754 = ~1'b0 ;
  assign y16755 = ~1'b0 ;
  assign y16756 = n23175 ;
  assign y16757 = n2569 ;
  assign y16758 = ~n23176 ;
  assign y16759 = ~n23178 ;
  assign y16760 = n21428 ;
  assign y16761 = n23179 ;
  assign y16762 = ~n23181 ;
  assign y16763 = ~n23182 ;
  assign y16764 = ~n23183 ;
  assign y16765 = ~n23188 ;
  assign y16766 = ~1'b0 ;
  assign y16767 = n3848 ;
  assign y16768 = ~1'b0 ;
  assign y16769 = n23190 ;
  assign y16770 = n23191 ;
  assign y16771 = ~1'b0 ;
  assign y16772 = ~1'b0 ;
  assign y16773 = ~n1081 ;
  assign y16774 = ~n23194 ;
  assign y16775 = ~1'b0 ;
  assign y16776 = ~n23195 ;
  assign y16777 = ~1'b0 ;
  assign y16778 = n23197 ;
  assign y16779 = ~1'b0 ;
  assign y16780 = n23200 ;
  assign y16781 = ~n7188 ;
  assign y16782 = n23202 ;
  assign y16783 = ~n23203 ;
  assign y16784 = ~1'b0 ;
  assign y16785 = ~n23205 ;
  assign y16786 = n23206 ;
  assign y16787 = ~1'b0 ;
  assign y16788 = n23210 ;
  assign y16789 = ~1'b0 ;
  assign y16790 = ~n23213 ;
  assign y16791 = ~1'b0 ;
  assign y16792 = n23215 ;
  assign y16793 = ~n23218 ;
  assign y16794 = n23224 ;
  assign y16795 = ~1'b0 ;
  assign y16796 = ~1'b0 ;
  assign y16797 = n23227 ;
  assign y16798 = ~n23230 ;
  assign y16799 = ~1'b0 ;
  assign y16800 = ~1'b0 ;
  assign y16801 = ~n23232 ;
  assign y16802 = ~1'b0 ;
  assign y16803 = ~n23234 ;
  assign y16804 = ~n3219 ;
  assign y16805 = n23236 ;
  assign y16806 = ~1'b0 ;
  assign y16807 = ~1'b0 ;
  assign y16808 = ~1'b0 ;
  assign y16809 = n23244 ;
  assign y16810 = ~1'b0 ;
  assign y16811 = ~n23252 ;
  assign y16812 = ~1'b0 ;
  assign y16813 = ~1'b0 ;
  assign y16814 = 1'b0 ;
  assign y16815 = n18463 ;
  assign y16816 = ~1'b0 ;
  assign y16817 = n23254 ;
  assign y16818 = ~n23259 ;
  assign y16819 = ~1'b0 ;
  assign y16820 = ~n23266 ;
  assign y16821 = ~n23271 ;
  assign y16822 = ~1'b0 ;
  assign y16823 = n12368 ;
  assign y16824 = ~n23273 ;
  assign y16825 = ~1'b0 ;
  assign y16826 = ~1'b0 ;
  assign y16827 = ~n23277 ;
  assign y16828 = ~1'b0 ;
  assign y16829 = n23278 ;
  assign y16830 = n23280 ;
  assign y16831 = ~1'b0 ;
  assign y16832 = n23283 ;
  assign y16833 = ~n23293 ;
  assign y16834 = ~n23296 ;
  assign y16835 = ~1'b0 ;
  assign y16836 = ~n23297 ;
  assign y16837 = 1'b0 ;
  assign y16838 = ~1'b0 ;
  assign y16839 = n23309 ;
  assign y16840 = ~1'b0 ;
  assign y16841 = ~n23310 ;
  assign y16842 = ~1'b0 ;
  assign y16843 = ~n23313 ;
  assign y16844 = n23314 ;
  assign y16845 = ~1'b0 ;
  assign y16846 = n8116 ;
  assign y16847 = ~1'b0 ;
  assign y16848 = ~1'b0 ;
  assign y16849 = n23317 ;
  assign y16850 = ~1'b0 ;
  assign y16851 = n23325 ;
  assign y16852 = ~n8922 ;
  assign y16853 = n2721 ;
  assign y16854 = ~1'b0 ;
  assign y16855 = n23327 ;
  assign y16856 = n23332 ;
  assign y16857 = n16422 ;
  assign y16858 = ~1'b0 ;
  assign y16859 = 1'b0 ;
  assign y16860 = ~n23338 ;
  assign y16861 = ~n23341 ;
  assign y16862 = ~1'b0 ;
  assign y16863 = ~n23342 ;
  assign y16864 = ~1'b0 ;
  assign y16865 = ~n23343 ;
  assign y16866 = ~1'b0 ;
  assign y16867 = ~1'b0 ;
  assign y16868 = n23345 ;
  assign y16869 = ~n3378 ;
  assign y16870 = ~n23346 ;
  assign y16871 = n20342 ;
  assign y16872 = ~n23350 ;
  assign y16873 = ~1'b0 ;
  assign y16874 = n23351 ;
  assign y16875 = ~n21168 ;
  assign y16876 = ~1'b0 ;
  assign y16877 = ~n23352 ;
  assign y16878 = n23353 ;
  assign y16879 = ~n23354 ;
  assign y16880 = ~1'b0 ;
  assign y16881 = n23355 ;
  assign y16882 = ~n23356 ;
  assign y16883 = ~n23358 ;
  assign y16884 = ~n23371 ;
  assign y16885 = n23373 ;
  assign y16886 = ~n23375 ;
  assign y16887 = ~1'b0 ;
  assign y16888 = ~1'b0 ;
  assign y16889 = ~n23377 ;
  assign y16890 = n23380 ;
  assign y16891 = ~1'b0 ;
  assign y16892 = ~n23385 ;
  assign y16893 = ~n16156 ;
  assign y16894 = ~1'b0 ;
  assign y16895 = ~1'b0 ;
  assign y16896 = n23386 ;
  assign y16897 = ~n23388 ;
  assign y16898 = ~n23392 ;
  assign y16899 = 1'b0 ;
  assign y16900 = n23399 ;
  assign y16901 = ~n23400 ;
  assign y16902 = ~1'b0 ;
  assign y16903 = ~1'b0 ;
  assign y16904 = ~n5032 ;
  assign y16905 = ~1'b0 ;
  assign y16906 = ~n23402 ;
  assign y16907 = ~n23408 ;
  assign y16908 = n13839 ;
  assign y16909 = ~n23410 ;
  assign y16910 = n23416 ;
  assign y16911 = ~1'b0 ;
  assign y16912 = ~1'b0 ;
  assign y16913 = ~1'b0 ;
  assign y16914 = ~1'b0 ;
  assign y16915 = ~n23418 ;
  assign y16916 = ~n23419 ;
  assign y16917 = n23421 ;
  assign y16918 = ~1'b0 ;
  assign y16919 = ~n23437 ;
  assign y16920 = n23444 ;
  assign y16921 = ~1'b0 ;
  assign y16922 = n20380 ;
  assign y16923 = ~n9004 ;
  assign y16924 = ~1'b0 ;
  assign y16925 = ~1'b0 ;
  assign y16926 = n23446 ;
  assign y16927 = ~1'b0 ;
  assign y16928 = n23447 ;
  assign y16929 = ~1'b0 ;
  assign y16930 = ~1'b0 ;
  assign y16931 = ~n21854 ;
  assign y16932 = ~1'b0 ;
  assign y16933 = ~n23450 ;
  assign y16934 = ~n23454 ;
  assign y16935 = n23455 ;
  assign y16936 = n23459 ;
  assign y16937 = ~n23461 ;
  assign y16938 = n23463 ;
  assign y16939 = ~n23464 ;
  assign y16940 = 1'b0 ;
  assign y16941 = ~1'b0 ;
  assign y16942 = ~n23466 ;
  assign y16943 = ~1'b0 ;
  assign y16944 = n23468 ;
  assign y16945 = ~1'b0 ;
  assign y16946 = ~1'b0 ;
  assign y16947 = ~n23472 ;
  assign y16948 = ~1'b0 ;
  assign y16949 = ~n23475 ;
  assign y16950 = ~n23477 ;
  assign y16951 = ~n23478 ;
  assign y16952 = ~1'b0 ;
  assign y16953 = n23480 ;
  assign y16954 = ~n23482 ;
  assign y16955 = n23488 ;
  assign y16956 = ~n23490 ;
  assign y16957 = n8019 ;
  assign y16958 = ~1'b0 ;
  assign y16959 = n12948 ;
  assign y16960 = n23491 ;
  assign y16961 = n23493 ;
  assign y16962 = n23498 ;
  assign y16963 = ~1'b0 ;
  assign y16964 = ~1'b0 ;
  assign y16965 = n612 ;
  assign y16966 = n23502 ;
  assign y16967 = n23510 ;
  assign y16968 = ~n23512 ;
  assign y16969 = ~1'b0 ;
  assign y16970 = n23514 ;
  assign y16971 = n23515 ;
  assign y16972 = ~n23516 ;
  assign y16973 = n23517 ;
  assign y16974 = 1'b0 ;
  assign y16975 = ~n23519 ;
  assign y16976 = n23521 ;
  assign y16977 = 1'b0 ;
  assign y16978 = n23522 ;
  assign y16979 = ~n23525 ;
  assign y16980 = ~1'b0 ;
  assign y16981 = ~n7227 ;
  assign y16982 = ~1'b0 ;
  assign y16983 = ~n3816 ;
  assign y16984 = ~1'b0 ;
  assign y16985 = ~1'b0 ;
  assign y16986 = ~1'b0 ;
  assign y16987 = n23528 ;
  assign y16988 = ~n23530 ;
  assign y16989 = ~1'b0 ;
  assign y16990 = ~n18286 ;
  assign y16991 = n23533 ;
  assign y16992 = ~1'b0 ;
  assign y16993 = ~n23536 ;
  assign y16994 = ~n1961 ;
  assign y16995 = ~n23539 ;
  assign y16996 = ~1'b0 ;
  assign y16997 = n23540 ;
  assign y16998 = ~1'b0 ;
  assign y16999 = ~n23542 ;
  assign y17000 = ~n23543 ;
  assign y17001 = ~1'b0 ;
  assign y17002 = n10587 ;
  assign y17003 = ~1'b0 ;
  assign y17004 = n19175 ;
  assign y17005 = ~1'b0 ;
  assign y17006 = ~1'b0 ;
  assign y17007 = ~1'b0 ;
  assign y17008 = ~1'b0 ;
  assign y17009 = ~1'b0 ;
  assign y17010 = n23548 ;
  assign y17011 = ~1'b0 ;
  assign y17012 = n23551 ;
  assign y17013 = 1'b0 ;
  assign y17014 = ~n23553 ;
  assign y17015 = ~n14809 ;
  assign y17016 = ~n23555 ;
  assign y17017 = ~1'b0 ;
  assign y17018 = n23558 ;
  assign y17019 = ~n23560 ;
  assign y17020 = n23566 ;
  assign y17021 = ~1'b0 ;
  assign y17022 = n23567 ;
  assign y17023 = ~1'b0 ;
  assign y17024 = n23568 ;
  assign y17025 = ~1'b0 ;
  assign y17026 = ~1'b0 ;
  assign y17027 = n23571 ;
  assign y17028 = n23577 ;
  assign y17029 = n23579 ;
  assign y17030 = n9619 ;
  assign y17031 = ~n23591 ;
  assign y17032 = 1'b0 ;
  assign y17033 = 1'b0 ;
  assign y17034 = ~n23597 ;
  assign y17035 = ~1'b0 ;
  assign y17036 = n23600 ;
  assign y17037 = n23604 ;
  assign y17038 = ~1'b0 ;
  assign y17039 = n23607 ;
  assign y17040 = ~1'b0 ;
  assign y17041 = n23614 ;
  assign y17042 = ~1'b0 ;
  assign y17043 = n23617 ;
  assign y17044 = ~1'b0 ;
  assign y17045 = ~1'b0 ;
  assign y17046 = ~n7388 ;
  assign y17047 = ~n23618 ;
  assign y17048 = ~n6218 ;
  assign y17049 = n23622 ;
  assign y17050 = ~1'b0 ;
  assign y17051 = ~n23628 ;
  assign y17052 = n23629 ;
  assign y17053 = ~1'b0 ;
  assign y17054 = ~1'b0 ;
  assign y17055 = ~n9548 ;
  assign y17056 = ~n23631 ;
  assign y17057 = n23635 ;
  assign y17058 = n23637 ;
  assign y17059 = ~1'b0 ;
  assign y17060 = n23639 ;
  assign y17061 = ~n23645 ;
  assign y17062 = n23647 ;
  assign y17063 = ~1'b0 ;
  assign y17064 = ~1'b0 ;
  assign y17065 = ~1'b0 ;
  assign y17066 = ~n23649 ;
  assign y17067 = ~1'b0 ;
  assign y17068 = ~1'b0 ;
  assign y17069 = n23650 ;
  assign y17070 = ~n23653 ;
  assign y17071 = ~1'b0 ;
  assign y17072 = ~1'b0 ;
  assign y17073 = n23655 ;
  assign y17074 = ~n5206 ;
  assign y17075 = ~n23674 ;
  assign y17076 = ~n23676 ;
  assign y17077 = ~n23679 ;
  assign y17078 = ~1'b0 ;
  assign y17079 = ~n23683 ;
  assign y17080 = ~n23686 ;
  assign y17081 = n23687 ;
  assign y17082 = n23691 ;
  assign y17083 = ~1'b0 ;
  assign y17084 = n23692 ;
  assign y17085 = n23694 ;
  assign y17086 = ~n6698 ;
  assign y17087 = ~n21587 ;
  assign y17088 = ~n23695 ;
  assign y17089 = n23696 ;
  assign y17090 = n23699 ;
  assign y17091 = n9703 ;
  assign y17092 = ~1'b0 ;
  assign y17093 = ~n23700 ;
  assign y17094 = n23702 ;
  assign y17095 = 1'b0 ;
  assign y17096 = n23707 ;
  assign y17097 = n8377 ;
  assign y17098 = ~n23710 ;
  assign y17099 = n23724 ;
  assign y17100 = n4750 ;
  assign y17101 = n843 ;
  assign y17102 = ~n23726 ;
  assign y17103 = n23728 ;
  assign y17104 = ~n23729 ;
  assign y17105 = ~n6955 ;
  assign y17106 = ~1'b0 ;
  assign y17107 = ~1'b0 ;
  assign y17108 = ~n23730 ;
  assign y17109 = n23736 ;
  assign y17110 = n23740 ;
  assign y17111 = n23741 ;
  assign y17112 = n23742 ;
  assign y17113 = ~1'b0 ;
  assign y17114 = ~n23745 ;
  assign y17115 = ~1'b0 ;
  assign y17116 = ~n23749 ;
  assign y17117 = ~1'b0 ;
  assign y17118 = n23751 ;
  assign y17119 = ~n23752 ;
  assign y17120 = n23754 ;
  assign y17121 = n23755 ;
  assign y17122 = n23757 ;
  assign y17123 = n23758 ;
  assign y17124 = ~1'b0 ;
  assign y17125 = ~1'b0 ;
  assign y17126 = n375 ;
  assign y17127 = ~n23761 ;
  assign y17128 = ~1'b0 ;
  assign y17129 = n23765 ;
  assign y17130 = ~n23768 ;
  assign y17131 = ~n23769 ;
  assign y17132 = n5833 ;
  assign y17133 = ~n13748 ;
  assign y17134 = 1'b0 ;
  assign y17135 = ~1'b0 ;
  assign y17136 = ~n23774 ;
  assign y17137 = ~1'b0 ;
  assign y17138 = ~n23778 ;
  assign y17139 = ~1'b0 ;
  assign y17140 = n23781 ;
  assign y17141 = n23785 ;
  assign y17142 = ~1'b0 ;
  assign y17143 = ~n23786 ;
  assign y17144 = n23788 ;
  assign y17145 = n23790 ;
  assign y17146 = ~1'b0 ;
  assign y17147 = ~n23792 ;
  assign y17148 = 1'b0 ;
  assign y17149 = ~n23797 ;
  assign y17150 = ~1'b0 ;
  assign y17151 = ~1'b0 ;
  assign y17152 = n23804 ;
  assign y17153 = n21961 ;
  assign y17154 = ~1'b0 ;
  assign y17155 = ~1'b0 ;
  assign y17156 = ~1'b0 ;
  assign y17157 = ~1'b0 ;
  assign y17158 = ~n23807 ;
  assign y17159 = ~n23813 ;
  assign y17160 = ~1'b0 ;
  assign y17161 = ~n23814 ;
  assign y17162 = n23815 ;
  assign y17163 = ~n11245 ;
  assign y17164 = ~1'b0 ;
  assign y17165 = n23817 ;
  assign y17166 = ~n23726 ;
  assign y17167 = ~1'b0 ;
  assign y17168 = ~1'b0 ;
  assign y17169 = ~n23822 ;
  assign y17170 = ~n5892 ;
  assign y17171 = n23826 ;
  assign y17172 = ~1'b0 ;
  assign y17173 = ~1'b0 ;
  assign y17174 = ~1'b0 ;
  assign y17175 = 1'b0 ;
  assign y17176 = n23828 ;
  assign y17177 = ~n23831 ;
  assign y17178 = ~1'b0 ;
  assign y17179 = n23833 ;
  assign y17180 = ~n23835 ;
  assign y17181 = n23838 ;
  assign y17182 = ~n23839 ;
  assign y17183 = ~1'b0 ;
  assign y17184 = ~1'b0 ;
  assign y17185 = n23841 ;
  assign y17186 = 1'b0 ;
  assign y17187 = ~1'b0 ;
  assign y17188 = ~1'b0 ;
  assign y17189 = ~n23842 ;
  assign y17190 = ~1'b0 ;
  assign y17191 = ~n23846 ;
  assign y17192 = 1'b0 ;
  assign y17193 = ~1'b0 ;
  assign y17194 = 1'b0 ;
  assign y17195 = n23847 ;
  assign y17196 = ~n23849 ;
  assign y17197 = ~1'b0 ;
  assign y17198 = ~1'b0 ;
  assign y17199 = ~1'b0 ;
  assign y17200 = n23851 ;
  assign y17201 = ~1'b0 ;
  assign y17202 = n23852 ;
  assign y17203 = 1'b0 ;
  assign y17204 = ~1'b0 ;
  assign y17205 = ~1'b0 ;
  assign y17206 = ~1'b0 ;
  assign y17207 = 1'b0 ;
  assign y17208 = ~n23854 ;
  assign y17209 = ~n23857 ;
  assign y17210 = ~1'b0 ;
  assign y17211 = ~n23859 ;
  assign y17212 = ~1'b0 ;
  assign y17213 = n23860 ;
  assign y17214 = n23861 ;
  assign y17215 = ~n23863 ;
  assign y17216 = ~1'b0 ;
  assign y17217 = ~n11973 ;
  assign y17218 = n23864 ;
  assign y17219 = ~n23867 ;
  assign y17220 = n23868 ;
  assign y17221 = ~n23869 ;
  assign y17222 = 1'b0 ;
  assign y17223 = ~n23870 ;
  assign y17224 = n23871 ;
  assign y17225 = n23876 ;
  assign y17226 = ~1'b0 ;
  assign y17227 = ~1'b0 ;
  assign y17228 = ~1'b0 ;
  assign y17229 = ~1'b0 ;
  assign y17230 = ~n23878 ;
  assign y17231 = ~n14429 ;
  assign y17232 = ~1'b0 ;
  assign y17233 = ~n23884 ;
  assign y17234 = ~n23886 ;
  assign y17235 = n879 ;
  assign y17236 = ~n23888 ;
  assign y17237 = ~1'b0 ;
  assign y17238 = ~1'b0 ;
  assign y17239 = ~1'b0 ;
  assign y17240 = ~1'b0 ;
  assign y17241 = ~1'b0 ;
  assign y17242 = ~n23890 ;
  assign y17243 = ~1'b0 ;
  assign y17244 = ~n23891 ;
  assign y17245 = ~1'b0 ;
  assign y17246 = n23892 ;
  assign y17247 = n23898 ;
  assign y17248 = ~1'b0 ;
  assign y17249 = n23901 ;
  assign y17250 = ~n23904 ;
  assign y17251 = ~1'b0 ;
  assign y17252 = n23905 ;
  assign y17253 = n23907 ;
  assign y17254 = ~1'b0 ;
  assign y17255 = ~1'b0 ;
  assign y17256 = n13977 ;
  assign y17257 = ~n23915 ;
  assign y17258 = ~1'b0 ;
  assign y17259 = ~n10548 ;
  assign y17260 = n23919 ;
  assign y17261 = n23924 ;
  assign y17262 = ~n23927 ;
  assign y17263 = n23929 ;
  assign y17264 = ~1'b0 ;
  assign y17265 = ~n23930 ;
  assign y17266 = ~1'b0 ;
  assign y17267 = ~1'b0 ;
  assign y17268 = ~n23931 ;
  assign y17269 = ~1'b0 ;
  assign y17270 = n3947 ;
  assign y17271 = ~1'b0 ;
  assign y17272 = ~n23935 ;
  assign y17273 = ~1'b0 ;
  assign y17274 = n23939 ;
  assign y17275 = ~n23941 ;
  assign y17276 = ~n23942 ;
  assign y17277 = 1'b0 ;
  assign y17278 = ~1'b0 ;
  assign y17279 = 1'b0 ;
  assign y17280 = n23944 ;
  assign y17281 = ~1'b0 ;
  assign y17282 = ~n23946 ;
  assign y17283 = ~n23947 ;
  assign y17284 = ~n23950 ;
  assign y17285 = ~n942 ;
  assign y17286 = ~1'b0 ;
  assign y17287 = ~1'b0 ;
  assign y17288 = ~1'b0 ;
  assign y17289 = ~n18289 ;
  assign y17290 = n23952 ;
  assign y17291 = ~n23954 ;
  assign y17292 = ~n23955 ;
  assign y17293 = n23956 ;
  assign y17294 = n23957 ;
  assign y17295 = ~1'b0 ;
  assign y17296 = n23964 ;
  assign y17297 = ~n23967 ;
  assign y17298 = n23968 ;
  assign y17299 = ~n23970 ;
  assign y17300 = ~n23973 ;
  assign y17301 = 1'b0 ;
  assign y17302 = ~n23978 ;
  assign y17303 = ~n23980 ;
  assign y17304 = ~n23985 ;
  assign y17305 = ~1'b0 ;
  assign y17306 = n23990 ;
  assign y17307 = ~n23993 ;
  assign y17308 = n23994 ;
  assign y17309 = ~n9191 ;
  assign y17310 = ~1'b0 ;
  assign y17311 = n22984 ;
  assign y17312 = n23996 ;
  assign y17313 = n23998 ;
  assign y17314 = ~n23999 ;
  assign y17315 = n24003 ;
  assign y17316 = ~n24007 ;
  assign y17317 = ~n24008 ;
  assign y17318 = ~n3384 ;
  assign y17319 = n24009 ;
  assign y17320 = ~n24010 ;
  assign y17321 = ~1'b0 ;
  assign y17322 = n24011 ;
  assign y17323 = n24015 ;
  assign y17324 = ~1'b0 ;
  assign y17325 = n24018 ;
  assign y17326 = ~n17592 ;
  assign y17327 = ~n16779 ;
  assign y17328 = ~n24019 ;
  assign y17329 = ~1'b0 ;
  assign y17330 = ~n24020 ;
  assign y17331 = ~n24022 ;
  assign y17332 = n24023 ;
  assign y17333 = ~1'b0 ;
  assign y17334 = n24024 ;
  assign y17335 = n24026 ;
  assign y17336 = n21109 ;
  assign y17337 = ~n24027 ;
  assign y17338 = ~1'b0 ;
  assign y17339 = n24029 ;
  assign y17340 = ~n24033 ;
  assign y17341 = ~n24035 ;
  assign y17342 = n10191 ;
  assign y17343 = ~1'b0 ;
  assign y17344 = ~n18408 ;
  assign y17345 = ~1'b0 ;
  assign y17346 = n24038 ;
  assign y17347 = ~1'b0 ;
  assign y17348 = n24044 ;
  assign y17349 = ~n24049 ;
  assign y17350 = ~n5269 ;
  assign y17351 = ~n24051 ;
  assign y17352 = n24052 ;
  assign y17353 = ~1'b0 ;
  assign y17354 = ~n24055 ;
  assign y17355 = ~1'b0 ;
  assign y17356 = ~n24057 ;
  assign y17357 = ~n24058 ;
  assign y17358 = ~1'b0 ;
  assign y17359 = ~n17119 ;
  assign y17360 = n24059 ;
  assign y17361 = n24061 ;
  assign y17362 = n24063 ;
  assign y17363 = ~1'b0 ;
  assign y17364 = ~1'b0 ;
  assign y17365 = n24066 ;
  assign y17366 = 1'b0 ;
  assign y17367 = n24067 ;
  assign y17368 = ~n24073 ;
  assign y17369 = ~1'b0 ;
  assign y17370 = n24074 ;
  assign y17371 = ~1'b0 ;
  assign y17372 = n3007 ;
  assign y17373 = n24076 ;
  assign y17374 = ~1'b0 ;
  assign y17375 = ~n1989 ;
  assign y17376 = ~1'b0 ;
  assign y17377 = n24077 ;
  assign y17378 = n13334 ;
  assign y17379 = n24084 ;
  assign y17380 = n24086 ;
  assign y17381 = ~1'b0 ;
  assign y17382 = n4419 ;
  assign y17383 = n24090 ;
  assign y17384 = ~1'b0 ;
  assign y17385 = ~n24091 ;
  assign y17386 = n24092 ;
  assign y17387 = n24094 ;
  assign y17388 = ~1'b0 ;
  assign y17389 = ~1'b0 ;
  assign y17390 = ~n24099 ;
  assign y17391 = 1'b0 ;
  assign y17392 = n24101 ;
  assign y17393 = 1'b0 ;
  assign y17394 = n24103 ;
  assign y17395 = ~n24104 ;
  assign y17396 = ~1'b0 ;
  assign y17397 = ~n24108 ;
  assign y17398 = ~1'b0 ;
  assign y17399 = n24109 ;
  assign y17400 = ~1'b0 ;
  assign y17401 = n24110 ;
  assign y17402 = ~n24118 ;
  assign y17403 = ~n24119 ;
  assign y17404 = 1'b0 ;
  assign y17405 = ~1'b0 ;
  assign y17406 = n24123 ;
  assign y17407 = ~n24124 ;
  assign y17408 = ~1'b0 ;
  assign y17409 = ~1'b0 ;
  assign y17410 = n24125 ;
  assign y17411 = ~1'b0 ;
  assign y17412 = ~n24128 ;
  assign y17413 = ~1'b0 ;
  assign y17414 = 1'b0 ;
  assign y17415 = n23794 ;
  assign y17416 = ~1'b0 ;
  assign y17417 = ~n22898 ;
  assign y17418 = 1'b0 ;
  assign y17419 = ~1'b0 ;
  assign y17420 = n24132 ;
  assign y17421 = n24133 ;
  assign y17422 = ~1'b0 ;
  assign y17423 = ~1'b0 ;
  assign y17424 = ~n24135 ;
  assign y17425 = ~1'b0 ;
  assign y17426 = ~n4095 ;
  assign y17427 = n24137 ;
  assign y17428 = ~1'b0 ;
  assign y17429 = ~1'b0 ;
  assign y17430 = ~1'b0 ;
  assign y17431 = ~n24138 ;
  assign y17432 = n11723 ;
  assign y17433 = ~1'b0 ;
  assign y17434 = ~n24139 ;
  assign y17435 = ~n8917 ;
  assign y17436 = ~1'b0 ;
  assign y17437 = n24141 ;
  assign y17438 = ~n24142 ;
  assign y17439 = n24145 ;
  assign y17440 = n24151 ;
  assign y17441 = n24152 ;
  assign y17442 = ~1'b0 ;
  assign y17443 = ~n24158 ;
  assign y17444 = n632 ;
  assign y17445 = ~n24161 ;
  assign y17446 = ~n24162 ;
  assign y17447 = ~n4700 ;
  assign y17448 = n24167 ;
  assign y17449 = ~1'b0 ;
  assign y17450 = n24169 ;
  assign y17451 = ~n24171 ;
  assign y17452 = ~n24175 ;
  assign y17453 = n24177 ;
  assign y17454 = n24181 ;
  assign y17455 = ~n24183 ;
  assign y17456 = ~1'b0 ;
  assign y17457 = ~1'b0 ;
  assign y17458 = n18832 ;
  assign y17459 = ~1'b0 ;
  assign y17460 = 1'b0 ;
  assign y17461 = ~1'b0 ;
  assign y17462 = ~1'b0 ;
  assign y17463 = n24185 ;
  assign y17464 = ~1'b0 ;
  assign y17465 = n24186 ;
  assign y17466 = ~n24195 ;
  assign y17467 = ~n24198 ;
  assign y17468 = ~n24202 ;
  assign y17469 = ~1'b0 ;
  assign y17470 = n24206 ;
  assign y17471 = n12325 ;
  assign y17472 = ~1'b0 ;
  assign y17473 = ~1'b0 ;
  assign y17474 = ~1'b0 ;
  assign y17475 = ~1'b0 ;
  assign y17476 = n24207 ;
  assign y17477 = ~n24209 ;
  assign y17478 = ~n24211 ;
  assign y17479 = ~1'b0 ;
  assign y17480 = n24212 ;
  assign y17481 = ~n6889 ;
  assign y17482 = 1'b0 ;
  assign y17483 = ~n24213 ;
  assign y17484 = n24217 ;
  assign y17485 = ~n24218 ;
  assign y17486 = ~n24220 ;
  assign y17487 = ~n24222 ;
  assign y17488 = ~n24223 ;
  assign y17489 = n24225 ;
  assign y17490 = ~n24227 ;
  assign y17491 = ~1'b0 ;
  assign y17492 = n24229 ;
  assign y17493 = ~1'b0 ;
  assign y17494 = ~n24231 ;
  assign y17495 = ~n24232 ;
  assign y17496 = ~n24233 ;
  assign y17497 = 1'b0 ;
  assign y17498 = ~1'b0 ;
  assign y17499 = ~1'b0 ;
  assign y17500 = n24235 ;
  assign y17501 = ~n24238 ;
  assign y17502 = ~1'b0 ;
  assign y17503 = ~n24240 ;
  assign y17504 = n2932 ;
  assign y17505 = ~1'b0 ;
  assign y17506 = ~n24242 ;
  assign y17507 = n24251 ;
  assign y17508 = ~1'b0 ;
  assign y17509 = ~1'b0 ;
  assign y17510 = ~1'b0 ;
  assign y17511 = ~n24252 ;
  assign y17512 = ~n24254 ;
  assign y17513 = ~n24255 ;
  assign y17514 = ~1'b0 ;
  assign y17515 = 1'b0 ;
  assign y17516 = 1'b0 ;
  assign y17517 = ~1'b0 ;
  assign y17518 = n24259 ;
  assign y17519 = n24265 ;
  assign y17520 = n24270 ;
  assign y17521 = ~1'b0 ;
  assign y17522 = 1'b0 ;
  assign y17523 = n24275 ;
  assign y17524 = n24277 ;
  assign y17525 = n24279 ;
  assign y17526 = ~1'b0 ;
  assign y17527 = ~n24288 ;
  assign y17528 = n24291 ;
  assign y17529 = ~1'b0 ;
  assign y17530 = n24293 ;
  assign y17531 = n7787 ;
  assign y17532 = ~1'b0 ;
  assign y17533 = ~n16573 ;
  assign y17534 = ~1'b0 ;
  assign y17535 = n24297 ;
  assign y17536 = n24299 ;
  assign y17537 = n24300 ;
  assign y17538 = ~n24302 ;
  assign y17539 = n24305 ;
  assign y17540 = 1'b0 ;
  assign y17541 = ~n24307 ;
  assign y17542 = n24312 ;
  assign y17543 = ~1'b0 ;
  assign y17544 = ~1'b0 ;
  assign y17545 = ~1'b0 ;
  assign y17546 = ~n24315 ;
  assign y17547 = ~1'b0 ;
  assign y17548 = ~1'b0 ;
  assign y17549 = 1'b0 ;
  assign y17550 = n24318 ;
  assign y17551 = ~1'b0 ;
  assign y17552 = ~1'b0 ;
  assign y17553 = ~1'b0 ;
  assign y17554 = n24320 ;
  assign y17555 = n24324 ;
  assign y17556 = ~n24325 ;
  assign y17557 = 1'b0 ;
  assign y17558 = ~1'b0 ;
  assign y17559 = ~1'b0 ;
  assign y17560 = ~n24328 ;
  assign y17561 = ~n24329 ;
  assign y17562 = n170 ;
  assign y17563 = n24332 ;
  assign y17564 = ~n24333 ;
  assign y17565 = n23493 ;
  assign y17566 = ~1'b0 ;
  assign y17567 = ~1'b0 ;
  assign y17568 = ~n24335 ;
  assign y17569 = n24339 ;
  assign y17570 = ~1'b0 ;
  assign y17571 = ~1'b0 ;
  assign y17572 = ~n24340 ;
  assign y17573 = n24341 ;
  assign y17574 = n24346 ;
  assign y17575 = ~1'b0 ;
  assign y17576 = ~n24347 ;
  assign y17577 = n24351 ;
  assign y17578 = ~1'b0 ;
  assign y17579 = ~1'b0 ;
  assign y17580 = n24352 ;
  assign y17581 = ~n24355 ;
  assign y17582 = n24360 ;
  assign y17583 = n24361 ;
  assign y17584 = ~1'b0 ;
  assign y17585 = ~1'b0 ;
  assign y17586 = ~1'b0 ;
  assign y17587 = ~n24365 ;
  assign y17588 = ~n24367 ;
  assign y17589 = n2157 ;
  assign y17590 = n24368 ;
  assign y17591 = ~1'b0 ;
  assign y17592 = n24370 ;
  assign y17593 = n24371 ;
  assign y17594 = ~1'b0 ;
  assign y17595 = ~1'b0 ;
  assign y17596 = ~1'b0 ;
  assign y17597 = ~1'b0 ;
  assign y17598 = ~n24372 ;
  assign y17599 = ~1'b0 ;
  assign y17600 = n12999 ;
  assign y17601 = ~n24373 ;
  assign y17602 = 1'b0 ;
  assign y17603 = ~1'b0 ;
  assign y17604 = ~1'b0 ;
  assign y17605 = ~n24378 ;
  assign y17606 = ~n24382 ;
  assign y17607 = ~n8973 ;
  assign y17608 = n24384 ;
  assign y17609 = ~n24386 ;
  assign y17610 = n24390 ;
  assign y17611 = n2242 ;
  assign y17612 = n24391 ;
  assign y17613 = ~1'b0 ;
  assign y17614 = n13847 ;
  assign y17615 = ~1'b0 ;
  assign y17616 = n24393 ;
  assign y17617 = ~n24396 ;
  assign y17618 = ~n24397 ;
  assign y17619 = n24398 ;
  assign y17620 = n24399 ;
  assign y17621 = ~n24401 ;
  assign y17622 = 1'b0 ;
  assign y17623 = n497 ;
  assign y17624 = ~1'b0 ;
  assign y17625 = n24405 ;
  assign y17626 = ~n24407 ;
  assign y17627 = ~1'b0 ;
  assign y17628 = ~n24408 ;
  assign y17629 = ~1'b0 ;
  assign y17630 = ~n24410 ;
  assign y17631 = ~1'b0 ;
  assign y17632 = n24413 ;
  assign y17633 = ~n24415 ;
  assign y17634 = ~n24424 ;
  assign y17635 = 1'b0 ;
  assign y17636 = n24427 ;
  assign y17637 = n24431 ;
  assign y17638 = ~n15879 ;
  assign y17639 = n24437 ;
  assign y17640 = ~n15100 ;
  assign y17641 = ~n24441 ;
  assign y17642 = n24445 ;
  assign y17643 = ~1'b0 ;
  assign y17644 = ~n24448 ;
  assign y17645 = ~n24449 ;
  assign y17646 = n24452 ;
  assign y17647 = ~1'b0 ;
  assign y17648 = n24455 ;
  assign y17649 = ~1'b0 ;
  assign y17650 = n24458 ;
  assign y17651 = ~n24460 ;
  assign y17652 = ~1'b0 ;
  assign y17653 = ~1'b0 ;
  assign y17654 = ~1'b0 ;
  assign y17655 = ~n24465 ;
  assign y17656 = ~n321 ;
  assign y17657 = 1'b0 ;
  assign y17658 = ~n24475 ;
  assign y17659 = ~1'b0 ;
  assign y17660 = ~n24477 ;
  assign y17661 = ~1'b0 ;
  assign y17662 = ~1'b0 ;
  assign y17663 = n7237 ;
  assign y17664 = 1'b0 ;
  assign y17665 = n24478 ;
  assign y17666 = ~1'b0 ;
  assign y17667 = ~1'b0 ;
  assign y17668 = ~n4735 ;
  assign y17669 = 1'b0 ;
  assign y17670 = 1'b0 ;
  assign y17671 = 1'b0 ;
  assign y17672 = ~1'b0 ;
  assign y17673 = ~n24479 ;
  assign y17674 = ~n24482 ;
  assign y17675 = n24483 ;
  assign y17676 = n24488 ;
  assign y17677 = n24491 ;
  assign y17678 = ~1'b0 ;
  assign y17679 = n24492 ;
  assign y17680 = n24494 ;
  assign y17681 = ~n24496 ;
  assign y17682 = ~n4897 ;
  assign y17683 = ~n24498 ;
  assign y17684 = ~n24501 ;
  assign y17685 = ~1'b0 ;
  assign y17686 = ~1'b0 ;
  assign y17687 = ~1'b0 ;
  assign y17688 = n24502 ;
  assign y17689 = n24503 ;
  assign y17690 = ~n24506 ;
  assign y17691 = n24507 ;
  assign y17692 = ~n24511 ;
  assign y17693 = ~n8282 ;
  assign y17694 = ~n24515 ;
  assign y17695 = n24516 ;
  assign y17696 = ~n24520 ;
  assign y17697 = ~n16219 ;
  assign y17698 = ~1'b0 ;
  assign y17699 = ~1'b0 ;
  assign y17700 = ~1'b0 ;
  assign y17701 = ~1'b0 ;
  assign y17702 = n24522 ;
  assign y17703 = ~1'b0 ;
  assign y17704 = ~n24524 ;
  assign y17705 = ~1'b0 ;
  assign y17706 = ~1'b0 ;
  assign y17707 = ~n24528 ;
  assign y17708 = n24530 ;
  assign y17709 = n24532 ;
  assign y17710 = ~1'b0 ;
  assign y17711 = n24533 ;
  assign y17712 = n24534 ;
  assign y17713 = ~1'b0 ;
  assign y17714 = ~n24535 ;
  assign y17715 = n5308 ;
  assign y17716 = 1'b0 ;
  assign y17717 = ~1'b0 ;
  assign y17718 = ~n24536 ;
  assign y17719 = ~n24538 ;
  assign y17720 = ~n24539 ;
  assign y17721 = ~n24541 ;
  assign y17722 = ~n24546 ;
  assign y17723 = ~n2687 ;
  assign y17724 = ~n24548 ;
  assign y17725 = 1'b0 ;
  assign y17726 = ~1'b0 ;
  assign y17727 = ~1'b0 ;
  assign y17728 = n24550 ;
  assign y17729 = n7023 ;
  assign y17730 = n24551 ;
  assign y17731 = ~n24555 ;
  assign y17732 = n24559 ;
  assign y17733 = n24560 ;
  assign y17734 = ~n24561 ;
  assign y17735 = n24562 ;
  assign y17736 = ~1'b0 ;
  assign y17737 = n24566 ;
  assign y17738 = n24567 ;
  assign y17739 = n24568 ;
  assign y17740 = ~1'b0 ;
  assign y17741 = n24570 ;
  assign y17742 = n24571 ;
  assign y17743 = ~1'b0 ;
  assign y17744 = ~1'b0 ;
  assign y17745 = n24576 ;
  assign y17746 = ~1'b0 ;
  assign y17747 = ~1'b0 ;
  assign y17748 = n24579 ;
  assign y17749 = n13857 ;
  assign y17750 = ~1'b0 ;
  assign y17751 = ~1'b0 ;
  assign y17752 = n9023 ;
  assign y17753 = ~1'b0 ;
  assign y17754 = n24582 ;
  assign y17755 = 1'b0 ;
  assign y17756 = ~n24584 ;
  assign y17757 = n24586 ;
  assign y17758 = ~n24587 ;
  assign y17759 = n8330 ;
  assign y17760 = ~1'b0 ;
  assign y17761 = n24589 ;
  assign y17762 = ~1'b0 ;
  assign y17763 = n3074 ;
  assign y17764 = ~n24593 ;
  assign y17765 = ~n24596 ;
  assign y17766 = ~1'b0 ;
  assign y17767 = n24599 ;
  assign y17768 = ~1'b0 ;
  assign y17769 = n24600 ;
  assign y17770 = ~n24602 ;
  assign y17771 = ~1'b0 ;
  assign y17772 = n10751 ;
  assign y17773 = ~n8547 ;
  assign y17774 = n24608 ;
  assign y17775 = n21799 ;
  assign y17776 = 1'b0 ;
  assign y17777 = ~n21962 ;
  assign y17778 = ~1'b0 ;
  assign y17779 = ~1'b0 ;
  assign y17780 = ~1'b0 ;
  assign y17781 = ~1'b0 ;
  assign y17782 = ~n24612 ;
  assign y17783 = 1'b0 ;
  assign y17784 = 1'b0 ;
  assign y17785 = ~1'b0 ;
  assign y17786 = ~1'b0 ;
  assign y17787 = n24613 ;
  assign y17788 = n20312 ;
  assign y17789 = 1'b0 ;
  assign y17790 = ~1'b0 ;
  assign y17791 = ~n24618 ;
  assign y17792 = ~1'b0 ;
  assign y17793 = n3800 ;
  assign y17794 = ~n24619 ;
  assign y17795 = n24620 ;
  assign y17796 = n24624 ;
  assign y17797 = 1'b0 ;
  assign y17798 = 1'b0 ;
  assign y17799 = ~n24626 ;
  assign y17800 = n24627 ;
  assign y17801 = n24629 ;
  assign y17802 = ~1'b0 ;
  assign y17803 = ~n24631 ;
  assign y17804 = ~n24641 ;
  assign y17805 = ~n400 ;
  assign y17806 = ~n24642 ;
  assign y17807 = ~1'b0 ;
  assign y17808 = ~n24643 ;
  assign y17809 = ~1'b0 ;
  assign y17810 = n24645 ;
  assign y17811 = 1'b0 ;
  assign y17812 = ~1'b0 ;
  assign y17813 = ~1'b0 ;
  assign y17814 = ~1'b0 ;
  assign y17815 = n24647 ;
  assign y17816 = ~n14692 ;
  assign y17817 = ~n24654 ;
  assign y17818 = ~1'b0 ;
  assign y17819 = ~n24656 ;
  assign y17820 = n24657 ;
  assign y17821 = n24659 ;
  assign y17822 = ~n24660 ;
  assign y17823 = ~1'b0 ;
  assign y17824 = n24662 ;
  assign y17825 = n713 ;
  assign y17826 = ~1'b0 ;
  assign y17827 = n24664 ;
  assign y17828 = ~1'b0 ;
  assign y17829 = 1'b0 ;
  assign y17830 = ~1'b0 ;
  assign y17831 = ~1'b0 ;
  assign y17832 = n13845 ;
  assign y17833 = ~n24665 ;
  assign y17834 = ~n24674 ;
  assign y17835 = ~1'b0 ;
  assign y17836 = ~n4186 ;
  assign y17837 = n24678 ;
  assign y17838 = n24679 ;
  assign y17839 = ~n24680 ;
  assign y17840 = ~n24682 ;
  assign y17841 = ~n24685 ;
  assign y17842 = n24690 ;
  assign y17843 = n24692 ;
  assign y17844 = ~1'b0 ;
  assign y17845 = ~n24694 ;
  assign y17846 = ~n24697 ;
  assign y17847 = ~n4061 ;
  assign y17848 = ~n5918 ;
  assign y17849 = ~1'b0 ;
  assign y17850 = ~1'b0 ;
  assign y17851 = ~1'b0 ;
  assign y17852 = ~1'b0 ;
  assign y17853 = 1'b0 ;
  assign y17854 = ~n24701 ;
  assign y17855 = ~1'b0 ;
  assign y17856 = n24702 ;
  assign y17857 = n24704 ;
  assign y17858 = n24705 ;
  assign y17859 = n10257 ;
  assign y17860 = 1'b0 ;
  assign y17861 = ~1'b0 ;
  assign y17862 = 1'b0 ;
  assign y17863 = ~1'b0 ;
  assign y17864 = ~1'b0 ;
  assign y17865 = ~n24707 ;
  assign y17866 = ~n24710 ;
  assign y17867 = ~1'b0 ;
  assign y17868 = n24711 ;
  assign y17869 = ~1'b0 ;
  assign y17870 = ~n24715 ;
  assign y17871 = ~n24717 ;
  assign y17872 = ~1'b0 ;
  assign y17873 = ~1'b0 ;
  assign y17874 = ~1'b0 ;
  assign y17875 = n24719 ;
  assign y17876 = ~1'b0 ;
  assign y17877 = n24721 ;
  assign y17878 = n24727 ;
  assign y17879 = ~1'b0 ;
  assign y17880 = ~n24729 ;
  assign y17881 = n415 ;
  assign y17882 = ~1'b0 ;
  assign y17883 = ~n22852 ;
  assign y17884 = 1'b0 ;
  assign y17885 = ~1'b0 ;
  assign y17886 = ~1'b0 ;
  assign y17887 = n11309 ;
  assign y17888 = n24732 ;
  assign y17889 = n24733 ;
  assign y17890 = ~1'b0 ;
  assign y17891 = ~1'b0 ;
  assign y17892 = n24755 ;
  assign y17893 = ~1'b0 ;
  assign y17894 = n24757 ;
  assign y17895 = ~n24760 ;
  assign y17896 = ~n24764 ;
  assign y17897 = ~1'b0 ;
  assign y17898 = ~1'b0 ;
  assign y17899 = n24765 ;
  assign y17900 = ~n24768 ;
  assign y17901 = n24770 ;
  assign y17902 = ~n24775 ;
  assign y17903 = ~1'b0 ;
  assign y17904 = ~1'b0 ;
  assign y17905 = n24777 ;
  assign y17906 = ~n24780 ;
  assign y17907 = ~1'b0 ;
  assign y17908 = ~n24781 ;
  assign y17909 = ~n2567 ;
  assign y17910 = n24783 ;
  assign y17911 = ~1'b0 ;
  assign y17912 = ~1'b0 ;
  assign y17913 = ~n24815 ;
  assign y17914 = ~1'b0 ;
  assign y17915 = n24827 ;
  assign y17916 = ~n24830 ;
  assign y17917 = 1'b0 ;
  assign y17918 = 1'b0 ;
  assign y17919 = ~1'b0 ;
  assign y17920 = ~n1243 ;
  assign y17921 = ~n24831 ;
  assign y17922 = 1'b0 ;
  assign y17923 = ~1'b0 ;
  assign y17924 = ~n24833 ;
  assign y17925 = ~1'b0 ;
  assign y17926 = n24835 ;
  assign y17927 = n24839 ;
  assign y17928 = ~1'b0 ;
  assign y17929 = ~n15525 ;
  assign y17930 = ~1'b0 ;
  assign y17931 = 1'b0 ;
  assign y17932 = ~n14916 ;
  assign y17933 = ~n24845 ;
  assign y17934 = ~n24850 ;
  assign y17935 = n24852 ;
  assign y17936 = n24853 ;
  assign y17937 = n24856 ;
  assign y17938 = ~n24860 ;
  assign y17939 = n24862 ;
  assign y17940 = n24864 ;
  assign y17941 = ~1'b0 ;
  assign y17942 = ~1'b0 ;
  assign y17943 = ~1'b0 ;
  assign y17944 = n24865 ;
  assign y17945 = ~1'b0 ;
  assign y17946 = ~n7720 ;
  assign y17947 = ~1'b0 ;
  assign y17948 = n24867 ;
  assign y17949 = ~n24869 ;
  assign y17950 = n24873 ;
  assign y17951 = ~n24874 ;
  assign y17952 = ~n24878 ;
  assign y17953 = n24880 ;
  assign y17954 = n6847 ;
  assign y17955 = 1'b0 ;
  assign y17956 = ~1'b0 ;
  assign y17957 = ~n24882 ;
  assign y17958 = n24885 ;
  assign y17959 = ~n24886 ;
  assign y17960 = 1'b0 ;
  assign y17961 = 1'b0 ;
  assign y17962 = n24889 ;
  assign y17963 = ~1'b0 ;
  assign y17964 = ~n24891 ;
  assign y17965 = ~n24895 ;
  assign y17966 = n24897 ;
  assign y17967 = n24900 ;
  assign y17968 = n24902 ;
  assign y17969 = n13698 ;
  assign y17970 = ~n24903 ;
  assign y17971 = ~1'b0 ;
  assign y17972 = ~n24908 ;
  assign y17973 = ~n5684 ;
  assign y17974 = ~n8793 ;
  assign y17975 = ~1'b0 ;
  assign y17976 = ~1'b0 ;
  assign y17977 = ~n24911 ;
  assign y17978 = ~n24914 ;
  assign y17979 = ~1'b0 ;
  assign y17980 = ~1'b0 ;
  assign y17981 = 1'b0 ;
  assign y17982 = ~1'b0 ;
  assign y17983 = 1'b0 ;
  assign y17984 = ~1'b0 ;
  assign y17985 = ~n24917 ;
  assign y17986 = n24920 ;
  assign y17987 = ~1'b0 ;
  assign y17988 = ~1'b0 ;
  assign y17989 = n24927 ;
  assign y17990 = ~1'b0 ;
  assign y17991 = 1'b0 ;
  assign y17992 = n24931 ;
  assign y17993 = n24932 ;
  assign y17994 = ~1'b0 ;
  assign y17995 = n24933 ;
  assign y17996 = ~n24935 ;
  assign y17997 = ~1'b0 ;
  assign y17998 = ~1'b0 ;
  assign y17999 = n24938 ;
  assign y18000 = n24939 ;
  assign y18001 = ~n24952 ;
  assign y18002 = ~1'b0 ;
  assign y18003 = ~1'b0 ;
  assign y18004 = n15092 ;
  assign y18005 = ~n24953 ;
  assign y18006 = ~n24954 ;
  assign y18007 = ~n24956 ;
  assign y18008 = ~1'b0 ;
  assign y18009 = n24957 ;
  assign y18010 = ~1'b0 ;
  assign y18011 = ~n24958 ;
  assign y18012 = 1'b0 ;
  assign y18013 = n24959 ;
  assign y18014 = ~n24961 ;
  assign y18015 = n24962 ;
  assign y18016 = ~n24963 ;
  assign y18017 = ~n24965 ;
  assign y18018 = ~1'b0 ;
  assign y18019 = ~1'b0 ;
  assign y18020 = ~n24967 ;
  assign y18021 = ~1'b0 ;
  assign y18022 = ~1'b0 ;
  assign y18023 = ~n24969 ;
  assign y18024 = ~1'b0 ;
  assign y18025 = ~1'b0 ;
  assign y18026 = ~1'b0 ;
  assign y18027 = ~1'b0 ;
  assign y18028 = ~n24972 ;
  assign y18029 = ~1'b0 ;
  assign y18030 = n24975 ;
  assign y18031 = ~1'b0 ;
  assign y18032 = n24981 ;
  assign y18033 = ~n9201 ;
  assign y18034 = ~n24982 ;
  assign y18035 = ~n18201 ;
  assign y18036 = ~n24987 ;
  assign y18037 = n185 ;
  assign y18038 = ~1'b0 ;
  assign y18039 = n24988 ;
  assign y18040 = n24989 ;
  assign y18041 = n24994 ;
  assign y18042 = ~1'b0 ;
  assign y18043 = ~n24997 ;
  assign y18044 = ~n24998 ;
  assign y18045 = n25000 ;
  assign y18046 = ~1'b0 ;
  assign y18047 = n25001 ;
  assign y18048 = n25003 ;
  assign y18049 = n25004 ;
  assign y18050 = n25005 ;
  assign y18051 = n25009 ;
  assign y18052 = n25012 ;
  assign y18053 = ~1'b0 ;
  assign y18054 = ~1'b0 ;
  assign y18055 = 1'b0 ;
  assign y18056 = ~n25013 ;
  assign y18057 = ~1'b0 ;
  assign y18058 = ~1'b0 ;
  assign y18059 = ~1'b0 ;
  assign y18060 = ~1'b0 ;
  assign y18061 = ~n1169 ;
  assign y18062 = ~1'b0 ;
  assign y18063 = n19400 ;
  assign y18064 = 1'b0 ;
  assign y18065 = ~n25015 ;
  assign y18066 = n25017 ;
  assign y18067 = ~1'b0 ;
  assign y18068 = n25018 ;
  assign y18069 = ~1'b0 ;
  assign y18070 = n25020 ;
  assign y18071 = ~1'b0 ;
  assign y18072 = ~1'b0 ;
  assign y18073 = ~1'b0 ;
  assign y18074 = ~n25023 ;
  assign y18075 = 1'b0 ;
  assign y18076 = ~1'b0 ;
  assign y18077 = ~1'b0 ;
  assign y18078 = ~1'b0 ;
  assign y18079 = n25026 ;
  assign y18080 = ~1'b0 ;
  assign y18081 = ~1'b0 ;
  assign y18082 = ~1'b0 ;
  assign y18083 = ~1'b0 ;
  assign y18084 = n25028 ;
  assign y18085 = n25033 ;
  assign y18086 = ~n5273 ;
  assign y18087 = ~n25036 ;
  assign y18088 = ~1'b0 ;
  assign y18089 = n153 ;
  assign y18090 = ~1'b0 ;
  assign y18091 = ~n25037 ;
  assign y18092 = n25038 ;
  assign y18093 = ~1'b0 ;
  assign y18094 = ~n25039 ;
  assign y18095 = ~n25041 ;
  assign y18096 = ~n25045 ;
  assign y18097 = ~1'b0 ;
  assign y18098 = ~n25047 ;
  assign y18099 = n25048 ;
  assign y18100 = ~n25051 ;
  assign y18101 = ~n25053 ;
  assign y18102 = ~n25055 ;
  assign y18103 = ~1'b0 ;
  assign y18104 = ~1'b0 ;
  assign y18105 = ~1'b0 ;
  assign y18106 = n25058 ;
  assign y18107 = ~n25059 ;
  assign y18108 = ~n25060 ;
  assign y18109 = ~n25061 ;
  assign y18110 = ~1'b0 ;
  assign y18111 = ~1'b0 ;
  assign y18112 = ~1'b0 ;
  assign y18113 = ~1'b0 ;
  assign y18114 = ~n25063 ;
  assign y18115 = ~n25065 ;
  assign y18116 = ~n25066 ;
  assign y18117 = ~1'b0 ;
  assign y18118 = ~1'b0 ;
  assign y18119 = ~n25068 ;
  assign y18120 = ~n1772 ;
  assign y18121 = ~1'b0 ;
  assign y18122 = ~1'b0 ;
  assign y18123 = n25072 ;
  assign y18124 = n25073 ;
  assign y18125 = 1'b0 ;
  assign y18126 = n25075 ;
  assign y18127 = 1'b0 ;
  assign y18128 = n25076 ;
  assign y18129 = ~1'b0 ;
  assign y18130 = n25079 ;
  assign y18131 = ~1'b0 ;
  assign y18132 = ~1'b0 ;
  assign y18133 = n9240 ;
  assign y18134 = ~n25081 ;
  assign y18135 = ~n25083 ;
  assign y18136 = ~n11319 ;
  assign y18137 = n25085 ;
  assign y18138 = n25088 ;
  assign y18139 = ~n25089 ;
  assign y18140 = ~n25092 ;
  assign y18141 = n25099 ;
  assign y18142 = ~n25100 ;
  assign y18143 = ~1'b0 ;
  assign y18144 = ~1'b0 ;
  assign y18145 = ~n7718 ;
  assign y18146 = n25105 ;
  assign y18147 = ~n25106 ;
  assign y18148 = n25111 ;
  assign y18149 = n25113 ;
  assign y18150 = ~n25116 ;
  assign y18151 = ~1'b0 ;
  assign y18152 = n25120 ;
  assign y18153 = ~n25127 ;
  assign y18154 = ~n25130 ;
  assign y18155 = ~n25131 ;
  assign y18156 = n25134 ;
  assign y18157 = ~n8656 ;
  assign y18158 = ~n25138 ;
  assign y18159 = ~1'b0 ;
  assign y18160 = ~1'b0 ;
  assign y18161 = ~n25139 ;
  assign y18162 = ~1'b0 ;
  assign y18163 = ~1'b0 ;
  assign y18164 = n25144 ;
  assign y18165 = ~1'b0 ;
  assign y18166 = ~n25146 ;
  assign y18167 = n25147 ;
  assign y18168 = n25148 ;
  assign y18169 = n25151 ;
  assign y18170 = ~n25154 ;
  assign y18171 = ~1'b0 ;
  assign y18172 = n10635 ;
  assign y18173 = ~1'b0 ;
  assign y18174 = n3333 ;
  assign y18175 = n25155 ;
  assign y18176 = 1'b0 ;
  assign y18177 = ~1'b0 ;
  assign y18178 = ~n25157 ;
  assign y18179 = ~1'b0 ;
  assign y18180 = ~1'b0 ;
  assign y18181 = ~n25161 ;
  assign y18182 = n25163 ;
  assign y18183 = ~1'b0 ;
  assign y18184 = n25164 ;
  assign y18185 = ~1'b0 ;
  assign y18186 = n25170 ;
  assign y18187 = ~1'b0 ;
  assign y18188 = ~1'b0 ;
  assign y18189 = ~1'b0 ;
  assign y18190 = ~n4070 ;
  assign y18191 = n25172 ;
  assign y18192 = ~n25177 ;
  assign y18193 = n25180 ;
  assign y18194 = ~n25181 ;
  assign y18195 = ~1'b0 ;
  assign y18196 = ~n25188 ;
  assign y18197 = ~n25190 ;
  assign y18198 = ~1'b0 ;
  assign y18199 = ~1'b0 ;
  assign y18200 = 1'b0 ;
  assign y18201 = n25195 ;
  assign y18202 = ~n25196 ;
  assign y18203 = n25199 ;
  assign y18204 = ~1'b0 ;
  assign y18205 = ~1'b0 ;
  assign y18206 = ~1'b0 ;
  assign y18207 = ~n25207 ;
  assign y18208 = n25209 ;
  assign y18209 = ~n25215 ;
  assign y18210 = ~1'b0 ;
  assign y18211 = ~1'b0 ;
  assign y18212 = n25216 ;
  assign y18213 = n25217 ;
  assign y18214 = ~1'b0 ;
  assign y18215 = ~1'b0 ;
  assign y18216 = ~n25220 ;
  assign y18217 = ~1'b0 ;
  assign y18218 = n21752 ;
  assign y18219 = ~1'b0 ;
  assign y18220 = ~1'b0 ;
  assign y18221 = ~1'b0 ;
  assign y18222 = ~n25222 ;
  assign y18223 = ~1'b0 ;
  assign y18224 = ~1'b0 ;
  assign y18225 = 1'b0 ;
  assign y18226 = ~n25225 ;
  assign y18227 = ~n25229 ;
  assign y18228 = n25233 ;
  assign y18229 = ~1'b0 ;
  assign y18230 = ~n25234 ;
  assign y18231 = ~1'b0 ;
  assign y18232 = n25131 ;
  assign y18233 = ~n25235 ;
  assign y18234 = ~1'b0 ;
  assign y18235 = ~n13618 ;
  assign y18236 = ~n25236 ;
  assign y18237 = n25237 ;
  assign y18238 = n11442 ;
  assign y18239 = ~1'b0 ;
  assign y18240 = n25239 ;
  assign y18241 = ~1'b0 ;
  assign y18242 = n23692 ;
  assign y18243 = n25241 ;
  assign y18244 = ~1'b0 ;
  assign y18245 = ~1'b0 ;
  assign y18246 = 1'b0 ;
  assign y18247 = n25242 ;
  assign y18248 = ~1'b0 ;
  assign y18249 = ~1'b0 ;
  assign y18250 = n1029 ;
  assign y18251 = ~n25244 ;
  assign y18252 = ~1'b0 ;
  assign y18253 = ~n25247 ;
  assign y18254 = ~1'b0 ;
  assign y18255 = ~n25249 ;
  assign y18256 = ~n5628 ;
  assign y18257 = ~n25252 ;
  assign y18258 = n6194 ;
  assign y18259 = ~1'b0 ;
  assign y18260 = n25256 ;
  assign y18261 = ~1'b0 ;
  assign y18262 = ~1'b0 ;
  assign y18263 = ~n25263 ;
  assign y18264 = ~n643 ;
  assign y18265 = ~1'b0 ;
  assign y18266 = n25267 ;
  assign y18267 = n13523 ;
  assign y18268 = n25269 ;
  assign y18269 = ~1'b0 ;
  assign y18270 = 1'b0 ;
  assign y18271 = ~1'b0 ;
  assign y18272 = ~1'b0 ;
  assign y18273 = ~1'b0 ;
  assign y18274 = ~1'b0 ;
  assign y18275 = ~n25271 ;
  assign y18276 = n25272 ;
  assign y18277 = ~n2476 ;
  assign y18278 = n8897 ;
  assign y18279 = ~n25277 ;
  assign y18280 = ~1'b0 ;
  assign y18281 = ~1'b0 ;
  assign y18282 = ~n25280 ;
  assign y18283 = ~n25283 ;
  assign y18284 = n25285 ;
  assign y18285 = ~n25287 ;
  assign y18286 = ~n25288 ;
  assign y18287 = ~1'b0 ;
  assign y18288 = ~1'b0 ;
  assign y18289 = ~n25289 ;
  assign y18290 = n23975 ;
  assign y18291 = n25290 ;
  assign y18292 = n16835 ;
  assign y18293 = n25293 ;
  assign y18294 = ~1'b0 ;
  assign y18295 = n25297 ;
  assign y18296 = n25298 ;
  assign y18297 = ~n25300 ;
  assign y18298 = 1'b0 ;
  assign y18299 = 1'b0 ;
  assign y18300 = ~n25302 ;
  assign y18301 = ~n25303 ;
  assign y18302 = n25304 ;
  assign y18303 = ~n25310 ;
  assign y18304 = ~n25314 ;
  assign y18305 = 1'b0 ;
  assign y18306 = n25315 ;
  assign y18307 = ~n25316 ;
  assign y18308 = ~1'b0 ;
  assign y18309 = ~1'b0 ;
  assign y18310 = ~n6454 ;
  assign y18311 = ~1'b0 ;
  assign y18312 = ~n2978 ;
  assign y18313 = 1'b0 ;
  assign y18314 = ~1'b0 ;
  assign y18315 = n25318 ;
  assign y18316 = n25320 ;
  assign y18317 = ~n25321 ;
  assign y18318 = ~n25325 ;
  assign y18319 = n25327 ;
  assign y18320 = ~1'b0 ;
  assign y18321 = ~n25329 ;
  assign y18322 = n25330 ;
  assign y18323 = ~1'b0 ;
  assign y18324 = ~n25333 ;
  assign y18325 = ~1'b0 ;
  assign y18326 = ~1'b0 ;
  assign y18327 = ~1'b0 ;
  assign y18328 = ~n25336 ;
  assign y18329 = n25338 ;
  assign y18330 = ~n25340 ;
  assign y18331 = ~1'b0 ;
  assign y18332 = ~1'b0 ;
  assign y18333 = ~n25341 ;
  assign y18334 = n1034 ;
  assign y18335 = ~1'b0 ;
  assign y18336 = ~1'b0 ;
  assign y18337 = ~n25343 ;
  assign y18338 = ~1'b0 ;
  assign y18339 = ~1'b0 ;
  assign y18340 = ~1'b0 ;
  assign y18341 = ~1'b0 ;
  assign y18342 = ~n25344 ;
  assign y18343 = n25346 ;
  assign y18344 = ~1'b0 ;
  assign y18345 = n25349 ;
  assign y18346 = n25350 ;
  assign y18347 = ~n25352 ;
  assign y18348 = n25354 ;
  assign y18349 = n25360 ;
  assign y18350 = ~1'b0 ;
  assign y18351 = ~1'b0 ;
  assign y18352 = ~1'b0 ;
  assign y18353 = n25364 ;
  assign y18354 = ~1'b0 ;
  assign y18355 = ~1'b0 ;
  assign y18356 = ~1'b0 ;
  assign y18357 = n25368 ;
  assign y18358 = ~1'b0 ;
  assign y18359 = ~1'b0 ;
  assign y18360 = ~n25373 ;
  assign y18361 = 1'b0 ;
  assign y18362 = 1'b0 ;
  assign y18363 = ~1'b0 ;
  assign y18364 = ~n10438 ;
  assign y18365 = n25376 ;
  assign y18366 = n7679 ;
  assign y18367 = n25377 ;
  assign y18368 = ~n25378 ;
  assign y18369 = n25379 ;
  assign y18370 = n25380 ;
  assign y18371 = ~1'b0 ;
  assign y18372 = ~n25390 ;
  assign y18373 = ~n25398 ;
  assign y18374 = 1'b0 ;
  assign y18375 = ~n25399 ;
  assign y18376 = ~1'b0 ;
  assign y18377 = ~1'b0 ;
  assign y18378 = n25403 ;
  assign y18379 = n25404 ;
  assign y18380 = n25409 ;
  assign y18381 = ~1'b0 ;
  assign y18382 = ~n25413 ;
  assign y18383 = n25414 ;
  assign y18384 = ~1'b0 ;
  assign y18385 = n25415 ;
  assign y18386 = ~1'b0 ;
  assign y18387 = ~1'b0 ;
  assign y18388 = n25419 ;
  assign y18389 = n25421 ;
  assign y18390 = ~1'b0 ;
  assign y18391 = ~1'b0 ;
  assign y18392 = 1'b0 ;
  assign y18393 = 1'b0 ;
  assign y18394 = 1'b0 ;
  assign y18395 = ~n25424 ;
  assign y18396 = 1'b0 ;
  assign y18397 = ~n1370 ;
  assign y18398 = ~1'b0 ;
  assign y18399 = ~n25426 ;
  assign y18400 = ~1'b0 ;
  assign y18401 = ~n25427 ;
  assign y18402 = ~1'b0 ;
  assign y18403 = n18594 ;
  assign y18404 = n25429 ;
  assign y18405 = ~1'b0 ;
  assign y18406 = n25431 ;
  assign y18407 = ~1'b0 ;
  assign y18408 = n13839 ;
  assign y18409 = ~1'b0 ;
  assign y18410 = ~n25432 ;
  assign y18411 = ~1'b0 ;
  assign y18412 = ~1'b0 ;
  assign y18413 = ~1'b0 ;
  assign y18414 = ~n25434 ;
  assign y18415 = n25436 ;
  assign y18416 = ~n25438 ;
  assign y18417 = ~1'b0 ;
  assign y18418 = ~1'b0 ;
  assign y18419 = ~1'b0 ;
  assign y18420 = ~n25441 ;
  assign y18421 = n25447 ;
  assign y18422 = ~n25448 ;
  assign y18423 = n25450 ;
  assign y18424 = ~n25452 ;
  assign y18425 = ~n25453 ;
  assign y18426 = n501 ;
  assign y18427 = ~1'b0 ;
  assign y18428 = ~1'b0 ;
  assign y18429 = n5140 ;
  assign y18430 = ~n25454 ;
  assign y18431 = ~n25455 ;
  assign y18432 = ~n25458 ;
  assign y18433 = ~1'b0 ;
  assign y18434 = n25462 ;
  assign y18435 = n25465 ;
  assign y18436 = ~n25469 ;
  assign y18437 = ~1'b0 ;
  assign y18438 = ~1'b0 ;
  assign y18439 = n25470 ;
  assign y18440 = n25471 ;
  assign y18441 = ~1'b0 ;
  assign y18442 = n20283 ;
  assign y18443 = ~1'b0 ;
  assign y18444 = n21943 ;
  assign y18445 = ~n25478 ;
  assign y18446 = n21985 ;
  assign y18447 = n25480 ;
  assign y18448 = n25483 ;
  assign y18449 = n25484 ;
  assign y18450 = ~1'b0 ;
  assign y18451 = ~1'b0 ;
  assign y18452 = ~1'b0 ;
  assign y18453 = ~1'b0 ;
  assign y18454 = ~n2723 ;
  assign y18455 = ~1'b0 ;
  assign y18456 = ~n25486 ;
  assign y18457 = n25488 ;
  assign y18458 = ~1'b0 ;
  assign y18459 = ~n25489 ;
  assign y18460 = n14429 ;
  assign y18461 = ~1'b0 ;
  assign y18462 = n25490 ;
  assign y18463 = ~1'b0 ;
  assign y18464 = ~n25493 ;
  assign y18465 = ~n25494 ;
  assign y18466 = ~1'b0 ;
  assign y18467 = ~n25497 ;
  assign y18468 = ~1'b0 ;
  assign y18469 = ~n25499 ;
  assign y18470 = ~1'b0 ;
  assign y18471 = ~n284 ;
  assign y18472 = ~n25502 ;
  assign y18473 = ~1'b0 ;
  assign y18474 = n25503 ;
  assign y18475 = ~1'b0 ;
  assign y18476 = n11308 ;
  assign y18477 = ~1'b0 ;
  assign y18478 = n25507 ;
  assign y18479 = ~1'b0 ;
  assign y18480 = ~n25509 ;
  assign y18481 = ~n25511 ;
  assign y18482 = ~n25514 ;
  assign y18483 = ~1'b0 ;
  assign y18484 = ~n25517 ;
  assign y18485 = ~n25519 ;
  assign y18486 = n11842 ;
  assign y18487 = n25521 ;
  assign y18488 = n25523 ;
  assign y18489 = ~n25539 ;
  assign y18490 = n25540 ;
  assign y18491 = ~n25541 ;
  assign y18492 = ~1'b0 ;
  assign y18493 = ~1'b0 ;
  assign y18494 = ~1'b0 ;
  assign y18495 = ~n25542 ;
  assign y18496 = n21509 ;
  assign y18497 = ~1'b0 ;
  assign y18498 = ~1'b0 ;
  assign y18499 = ~1'b0 ;
  assign y18500 = n13492 ;
  assign y18501 = ~n25543 ;
  assign y18502 = ~1'b0 ;
  assign y18503 = n25545 ;
  assign y18504 = n25548 ;
  assign y18505 = ~1'b0 ;
  assign y18506 = n25549 ;
  assign y18507 = n25552 ;
  assign y18508 = 1'b0 ;
  assign y18509 = ~1'b0 ;
  assign y18510 = n25555 ;
  assign y18511 = n25557 ;
  assign y18512 = ~1'b0 ;
  assign y18513 = n25558 ;
  assign y18514 = n25562 ;
  assign y18515 = 1'b0 ;
  assign y18516 = n25563 ;
  assign y18517 = ~1'b0 ;
  assign y18518 = n25568 ;
  assign y18519 = ~n25570 ;
  assign y18520 = n25572 ;
  assign y18521 = ~1'b0 ;
  assign y18522 = ~1'b0 ;
  assign y18523 = ~1'b0 ;
  assign y18524 = n25575 ;
  assign y18525 = ~n25577 ;
  assign y18526 = n25579 ;
  assign y18527 = n11931 ;
  assign y18528 = ~n25580 ;
  assign y18529 = ~n25581 ;
  assign y18530 = ~1'b0 ;
  assign y18531 = n25585 ;
  assign y18532 = ~1'b0 ;
  assign y18533 = n25587 ;
  assign y18534 = ~n25589 ;
  assign y18535 = n25592 ;
  assign y18536 = ~n25593 ;
  assign y18537 = ~n25594 ;
  assign y18538 = n25597 ;
  assign y18539 = ~1'b0 ;
  assign y18540 = ~1'b0 ;
  assign y18541 = n25598 ;
  assign y18542 = n25600 ;
  assign y18543 = ~1'b0 ;
  assign y18544 = ~n25602 ;
  assign y18545 = ~n25605 ;
  assign y18546 = ~n25606 ;
  assign y18547 = ~1'b0 ;
  assign y18548 = ~1'b0 ;
  assign y18549 = ~n25607 ;
  assign y18550 = n25612 ;
  assign y18551 = ~n25616 ;
  assign y18552 = n25617 ;
  assign y18553 = ~1'b0 ;
  assign y18554 = n6234 ;
  assign y18555 = n25619 ;
  assign y18556 = ~1'b0 ;
  assign y18557 = ~1'b0 ;
  assign y18558 = n25620 ;
  assign y18559 = ~n25624 ;
  assign y18560 = n25625 ;
  assign y18561 = n25626 ;
  assign y18562 = ~1'b0 ;
  assign y18563 = ~1'b0 ;
  assign y18564 = 1'b0 ;
  assign y18565 = n15167 ;
  assign y18566 = ~n10126 ;
  assign y18567 = ~1'b0 ;
  assign y18568 = ~1'b0 ;
  assign y18569 = ~n25628 ;
  assign y18570 = 1'b0 ;
  assign y18571 = ~n25632 ;
  assign y18572 = n25635 ;
  assign y18573 = 1'b0 ;
  assign y18574 = ~n25636 ;
  assign y18575 = ~n25638 ;
  assign y18576 = n25640 ;
  assign y18577 = n25642 ;
  assign y18578 = n25644 ;
  assign y18579 = ~n25645 ;
  assign y18580 = n25647 ;
  assign y18581 = ~1'b0 ;
  assign y18582 = n25651 ;
  assign y18583 = n25656 ;
  assign y18584 = ~n25657 ;
  assign y18585 = 1'b0 ;
  assign y18586 = ~n7440 ;
  assign y18587 = ~n25658 ;
  assign y18588 = n25661 ;
  assign y18589 = n128 ;
  assign y18590 = ~1'b0 ;
  assign y18591 = n25665 ;
  assign y18592 = n25666 ;
  assign y18593 = n25668 ;
  assign y18594 = ~1'b0 ;
  assign y18595 = n25671 ;
  assign y18596 = ~n25673 ;
  assign y18597 = ~n25676 ;
  assign y18598 = ~n25678 ;
  assign y18599 = n25679 ;
  assign y18600 = ~1'b0 ;
  assign y18601 = 1'b0 ;
  assign y18602 = n7395 ;
  assign y18603 = ~n25680 ;
  assign y18604 = n12280 ;
  assign y18605 = ~1'b0 ;
  assign y18606 = ~n25682 ;
  assign y18607 = n25683 ;
  assign y18608 = 1'b0 ;
  assign y18609 = ~1'b0 ;
  assign y18610 = n25685 ;
  assign y18611 = ~n25686 ;
  assign y18612 = n25690 ;
  assign y18613 = ~1'b0 ;
  assign y18614 = ~n25691 ;
  assign y18615 = ~n25695 ;
  assign y18616 = ~n25698 ;
  assign y18617 = ~n1188 ;
  assign y18618 = n25699 ;
  assign y18619 = ~1'b0 ;
  assign y18620 = ~1'b0 ;
  assign y18621 = ~n25703 ;
  assign y18622 = ~1'b0 ;
  assign y18623 = ~n25707 ;
  assign y18624 = ~1'b0 ;
  assign y18625 = n25708 ;
  assign y18626 = ~1'b0 ;
  assign y18627 = n25709 ;
  assign y18628 = ~1'b0 ;
  assign y18629 = ~1'b0 ;
  assign y18630 = ~1'b0 ;
  assign y18631 = ~n25711 ;
  assign y18632 = ~n25715 ;
  assign y18633 = ~1'b0 ;
  assign y18634 = ~1'b0 ;
  assign y18635 = n25717 ;
  assign y18636 = ~n25718 ;
  assign y18637 = ~n25719 ;
  assign y18638 = ~n25721 ;
  assign y18639 = n25724 ;
  assign y18640 = n25725 ;
  assign y18641 = ~n25729 ;
  assign y18642 = n25730 ;
  assign y18643 = n4742 ;
  assign y18644 = ~1'b0 ;
  assign y18645 = ~n25731 ;
  assign y18646 = n25740 ;
  assign y18647 = n25742 ;
  assign y18648 = ~1'b0 ;
  assign y18649 = ~1'b0 ;
  assign y18650 = ~1'b0 ;
  assign y18651 = n25744 ;
  assign y18652 = ~n25745 ;
  assign y18653 = n25747 ;
  assign y18654 = ~1'b0 ;
  assign y18655 = ~1'b0 ;
  assign y18656 = ~n25750 ;
  assign y18657 = ~n25753 ;
  assign y18658 = ~1'b0 ;
  assign y18659 = ~1'b0 ;
  assign y18660 = n25754 ;
  assign y18661 = ~n25755 ;
  assign y18662 = ~1'b0 ;
  assign y18663 = ~1'b0 ;
  assign y18664 = n25757 ;
  assign y18665 = ~1'b0 ;
  assign y18666 = ~n25758 ;
  assign y18667 = ~n172 ;
  assign y18668 = ~1'b0 ;
  assign y18669 = ~1'b0 ;
  assign y18670 = ~1'b0 ;
  assign y18671 = ~1'b0 ;
  assign y18672 = n25759 ;
  assign y18673 = ~n25760 ;
  assign y18674 = ~1'b0 ;
  assign y18675 = ~1'b0 ;
  assign y18676 = n25761 ;
  assign y18677 = ~1'b0 ;
  assign y18678 = ~n25768 ;
  assign y18679 = ~1'b0 ;
  assign y18680 = ~n25769 ;
  assign y18681 = n25771 ;
  assign y18682 = ~1'b0 ;
  assign y18683 = ~n25777 ;
  assign y18684 = ~1'b0 ;
  assign y18685 = ~n25784 ;
  assign y18686 = n3567 ;
  assign y18687 = ~1'b0 ;
  assign y18688 = ~n25785 ;
  assign y18689 = ~n25786 ;
  assign y18690 = n25787 ;
  assign y18691 = ~1'b0 ;
  assign y18692 = n25792 ;
  assign y18693 = ~1'b0 ;
  assign y18694 = n25794 ;
  assign y18695 = ~1'b0 ;
  assign y18696 = 1'b0 ;
  assign y18697 = ~1'b0 ;
  assign y18698 = n25795 ;
  assign y18699 = ~n1306 ;
  assign y18700 = ~1'b0 ;
  assign y18701 = ~1'b0 ;
  assign y18702 = n25798 ;
  assign y18703 = ~1'b0 ;
  assign y18704 = ~n25799 ;
  assign y18705 = ~1'b0 ;
  assign y18706 = ~1'b0 ;
  assign y18707 = ~n25801 ;
  assign y18708 = ~n9778 ;
  assign y18709 = n25805 ;
  assign y18710 = ~n25806 ;
  assign y18711 = ~n5428 ;
  assign y18712 = ~n25809 ;
  assign y18713 = n25810 ;
  assign y18714 = ~1'b0 ;
  assign y18715 = ~n25814 ;
  assign y18716 = 1'b0 ;
  assign y18717 = n25815 ;
  assign y18718 = 1'b0 ;
  assign y18719 = ~n25816 ;
  assign y18720 = ~n25818 ;
  assign y18721 = ~1'b0 ;
  assign y18722 = ~n25819 ;
  assign y18723 = ~1'b0 ;
  assign y18724 = ~n25822 ;
  assign y18725 = n25825 ;
  assign y18726 = ~n25826 ;
  assign y18727 = ~n1430 ;
  assign y18728 = ~n25830 ;
  assign y18729 = n25832 ;
  assign y18730 = ~1'b0 ;
  assign y18731 = ~1'b0 ;
  assign y18732 = ~1'b0 ;
  assign y18733 = ~n25834 ;
  assign y18734 = ~1'b0 ;
  assign y18735 = ~n25836 ;
  assign y18736 = ~n596 ;
  assign y18737 = ~n25837 ;
  assign y18738 = ~n25841 ;
  assign y18739 = ~1'b0 ;
  assign y18740 = n1950 ;
  assign y18741 = n25843 ;
  assign y18742 = ~1'b0 ;
  assign y18743 = 1'b0 ;
  assign y18744 = n25849 ;
  assign y18745 = n2196 ;
  assign y18746 = n25855 ;
  assign y18747 = n25856 ;
  assign y18748 = ~n25859 ;
  assign y18749 = ~n25861 ;
  assign y18750 = ~1'b0 ;
  assign y18751 = ~n25863 ;
  assign y18752 = ~n25864 ;
  assign y18753 = ~1'b0 ;
  assign y18754 = n25865 ;
  assign y18755 = ~1'b0 ;
  assign y18756 = ~1'b0 ;
  assign y18757 = n25867 ;
  assign y18758 = ~1'b0 ;
  assign y18759 = ~1'b0 ;
  assign y18760 = n25872 ;
  assign y18761 = ~1'b0 ;
  assign y18762 = ~n25873 ;
  assign y18763 = n25875 ;
  assign y18764 = ~n25876 ;
  assign y18765 = ~1'b0 ;
  assign y18766 = ~n25882 ;
  assign y18767 = ~n25890 ;
  assign y18768 = ~1'b0 ;
  assign y18769 = ~n25894 ;
  assign y18770 = ~n2460 ;
  assign y18771 = ~1'b0 ;
  assign y18772 = ~n25896 ;
  assign y18773 = n13414 ;
  assign y18774 = ~n25898 ;
  assign y18775 = ~1'b0 ;
  assign y18776 = n25899 ;
  assign y18777 = n25900 ;
  assign y18778 = ~n25901 ;
  assign y18779 = n25903 ;
  assign y18780 = ~1'b0 ;
  assign y18781 = ~n25905 ;
  assign y18782 = ~1'b0 ;
  assign y18783 = ~n25908 ;
  assign y18784 = n10414 ;
  assign y18785 = ~n25910 ;
  assign y18786 = ~n25913 ;
  assign y18787 = ~1'b0 ;
  assign y18788 = ~1'b0 ;
  assign y18789 = n25919 ;
  assign y18790 = ~1'b0 ;
  assign y18791 = n25921 ;
  assign y18792 = n25922 ;
  assign y18793 = n25923 ;
  assign y18794 = ~1'b0 ;
  assign y18795 = ~1'b0 ;
  assign y18796 = n25924 ;
  assign y18797 = n15984 ;
  assign y18798 = n10551 ;
  assign y18799 = ~n25927 ;
  assign y18800 = ~n25933 ;
  assign y18801 = ~n25935 ;
  assign y18802 = ~1'b0 ;
  assign y18803 = ~n25938 ;
  assign y18804 = n25939 ;
  assign y18805 = 1'b0 ;
  assign y18806 = 1'b0 ;
  assign y18807 = 1'b0 ;
  assign y18808 = ~n25942 ;
  assign y18809 = ~1'b0 ;
  assign y18810 = ~1'b0 ;
  assign y18811 = ~n25944 ;
  assign y18812 = n25946 ;
  assign y18813 = ~n25947 ;
  assign y18814 = ~1'b0 ;
  assign y18815 = ~1'b0 ;
  assign y18816 = n4742 ;
  assign y18817 = n25948 ;
  assign y18818 = n25949 ;
  assign y18819 = ~n25956 ;
  assign y18820 = n25957 ;
  assign y18821 = n25958 ;
  assign y18822 = n25959 ;
  assign y18823 = ~1'b0 ;
  assign y18824 = ~1'b0 ;
  assign y18825 = ~n25960 ;
  assign y18826 = ~n25961 ;
  assign y18827 = n25962 ;
  assign y18828 = ~1'b0 ;
  assign y18829 = ~1'b0 ;
  assign y18830 = ~n25963 ;
  assign y18831 = n25967 ;
  assign y18832 = n25968 ;
  assign y18833 = ~1'b0 ;
  assign y18834 = ~n23118 ;
  assign y18835 = ~1'b0 ;
  assign y18836 = n25969 ;
  assign y18837 = ~n5580 ;
  assign y18838 = n25970 ;
  assign y18839 = n25971 ;
  assign y18840 = ~1'b0 ;
  assign y18841 = n25972 ;
  assign y18842 = ~n7179 ;
  assign y18843 = ~n15655 ;
  assign y18844 = ~n25975 ;
  assign y18845 = ~n25976 ;
  assign y18846 = ~n25982 ;
  assign y18847 = ~n25983 ;
  assign y18848 = ~n25984 ;
  assign y18849 = ~n25985 ;
  assign y18850 = n25986 ;
  assign y18851 = 1'b0 ;
  assign y18852 = n25988 ;
  assign y18853 = ~1'b0 ;
  assign y18854 = n25989 ;
  assign y18855 = ~n7511 ;
  assign y18856 = ~1'b0 ;
  assign y18857 = ~1'b0 ;
  assign y18858 = ~n25992 ;
  assign y18859 = ~1'b0 ;
  assign y18860 = ~n25993 ;
  assign y18861 = ~n25996 ;
  assign y18862 = ~n26000 ;
  assign y18863 = ~n26005 ;
  assign y18864 = ~1'b0 ;
  assign y18865 = n26006 ;
  assign y18866 = n26011 ;
  assign y18867 = n26013 ;
  assign y18868 = n26014 ;
  assign y18869 = ~1'b0 ;
  assign y18870 = n26015 ;
  assign y18871 = ~1'b0 ;
  assign y18872 = ~1'b0 ;
  assign y18873 = ~n9090 ;
  assign y18874 = 1'b0 ;
  assign y18875 = ~n26016 ;
  assign y18876 = ~n26022 ;
  assign y18877 = ~n26023 ;
  assign y18878 = ~n15162 ;
  assign y18879 = ~1'b0 ;
  assign y18880 = ~n10273 ;
  assign y18881 = ~1'b0 ;
  assign y18882 = ~1'b0 ;
  assign y18883 = ~1'b0 ;
  assign y18884 = ~1'b0 ;
  assign y18885 = ~n26025 ;
  assign y18886 = ~1'b0 ;
  assign y18887 = ~1'b0 ;
  assign y18888 = n26027 ;
  assign y18889 = n26028 ;
  assign y18890 = ~n26030 ;
  assign y18891 = ~n26032 ;
  assign y18892 = n26034 ;
  assign y18893 = ~n26035 ;
  assign y18894 = n26036 ;
  assign y18895 = ~1'b0 ;
  assign y18896 = ~1'b0 ;
  assign y18897 = ~n26037 ;
  assign y18898 = ~1'b0 ;
  assign y18899 = 1'b0 ;
  assign y18900 = 1'b0 ;
  assign y18901 = 1'b0 ;
  assign y18902 = ~1'b0 ;
  assign y18903 = n3738 ;
  assign y18904 = n26039 ;
  assign y18905 = n976 ;
  assign y18906 = ~1'b0 ;
  assign y18907 = ~1'b0 ;
  assign y18908 = ~n26043 ;
  assign y18909 = ~1'b0 ;
  assign y18910 = ~1'b0 ;
  assign y18911 = n26046 ;
  assign y18912 = n26049 ;
  assign y18913 = ~n26050 ;
  assign y18914 = ~n26052 ;
  assign y18915 = n26054 ;
  assign y18916 = ~1'b0 ;
  assign y18917 = ~n26056 ;
  assign y18918 = n26058 ;
  assign y18919 = ~1'b0 ;
  assign y18920 = ~1'b0 ;
  assign y18921 = ~n19175 ;
  assign y18922 = n26062 ;
  assign y18923 = ~1'b0 ;
  assign y18924 = ~1'b0 ;
  assign y18925 = n26063 ;
  assign y18926 = ~1'b0 ;
  assign y18927 = ~1'b0 ;
  assign y18928 = ~n26065 ;
  assign y18929 = n26067 ;
  assign y18930 = ~n26074 ;
  assign y18931 = ~1'b0 ;
  assign y18932 = ~1'b0 ;
  assign y18933 = ~n13990 ;
  assign y18934 = ~n26075 ;
  assign y18935 = n26076 ;
  assign y18936 = n17969 ;
  assign y18937 = n26079 ;
  assign y18938 = ~1'b0 ;
  assign y18939 = ~1'b0 ;
  assign y18940 = ~1'b0 ;
  assign y18941 = ~1'b0 ;
  assign y18942 = n26083 ;
  assign y18943 = ~n26084 ;
  assign y18944 = ~1'b0 ;
  assign y18945 = ~n26086 ;
  assign y18946 = 1'b0 ;
  assign y18947 = n26087 ;
  assign y18948 = n21366 ;
  assign y18949 = 1'b0 ;
  assign y18950 = n26096 ;
  assign y18951 = ~n15287 ;
  assign y18952 = ~1'b0 ;
  assign y18953 = ~1'b0 ;
  assign y18954 = ~1'b0 ;
  assign y18955 = ~n2822 ;
  assign y18956 = ~1'b0 ;
  assign y18957 = n26099 ;
  assign y18958 = ~n26103 ;
  assign y18959 = ~n26107 ;
  assign y18960 = ~1'b0 ;
  assign y18961 = ~n26108 ;
  assign y18962 = ~1'b0 ;
  assign y18963 = n26109 ;
  assign y18964 = ~n799 ;
  assign y18965 = 1'b0 ;
  assign y18966 = ~1'b0 ;
  assign y18967 = ~n26116 ;
  assign y18968 = n26118 ;
  assign y18969 = ~n6272 ;
  assign y18970 = ~1'b0 ;
  assign y18971 = ~n5468 ;
  assign y18972 = n26122 ;
  assign y18973 = 1'b0 ;
  assign y18974 = ~1'b0 ;
  assign y18975 = ~n26124 ;
  assign y18976 = ~n26126 ;
  assign y18977 = ~n26127 ;
  assign y18978 = n26130 ;
  assign y18979 = ~n26131 ;
  assign y18980 = ~n26132 ;
  assign y18981 = ~1'b0 ;
  assign y18982 = ~n26141 ;
  assign y18983 = 1'b0 ;
  assign y18984 = ~n26142 ;
  assign y18985 = n26143 ;
  assign y18986 = ~n26144 ;
  assign y18987 = n26147 ;
  assign y18988 = ~n26148 ;
  assign y18989 = n26153 ;
  assign y18990 = n26159 ;
  assign y18991 = n26168 ;
  assign y18992 = n26169 ;
  assign y18993 = ~n26171 ;
  assign y18994 = ~n26179 ;
  assign y18995 = ~1'b0 ;
  assign y18996 = ~n26180 ;
  assign y18997 = ~1'b0 ;
  assign y18998 = n26183 ;
  assign y18999 = ~n26184 ;
  assign y19000 = n26185 ;
  assign y19001 = 1'b0 ;
  assign y19002 = ~1'b0 ;
  assign y19003 = ~1'b0 ;
  assign y19004 = ~1'b0 ;
  assign y19005 = ~1'b0 ;
  assign y19006 = ~n26186 ;
  assign y19007 = n26187 ;
  assign y19008 = ~n26188 ;
  assign y19009 = ~n26189 ;
  assign y19010 = ~1'b0 ;
  assign y19011 = n26190 ;
  assign y19012 = n26194 ;
  assign y19013 = n26195 ;
  assign y19014 = ~n26196 ;
  assign y19015 = ~1'b0 ;
  assign y19016 = ~n26197 ;
  assign y19017 = ~1'b0 ;
  assign y19018 = ~n26200 ;
  assign y19019 = ~n26201 ;
  assign y19020 = ~1'b0 ;
  assign y19021 = ~n17921 ;
  assign y19022 = ~1'b0 ;
  assign y19023 = n26206 ;
  assign y19024 = ~n5934 ;
  assign y19025 = ~n26209 ;
  assign y19026 = ~x7 ;
  assign y19027 = n26210 ;
  assign y19028 = n14398 ;
  assign y19029 = ~1'b0 ;
  assign y19030 = ~1'b0 ;
  assign y19031 = n26211 ;
  assign y19032 = ~1'b0 ;
  assign y19033 = ~n26214 ;
  assign y19034 = n26215 ;
  assign y19035 = 1'b0 ;
  assign y19036 = ~n6385 ;
  assign y19037 = ~1'b0 ;
  assign y19038 = n26225 ;
  assign y19039 = ~1'b0 ;
  assign y19040 = ~1'b0 ;
  assign y19041 = n26227 ;
  assign y19042 = n26228 ;
  assign y19043 = ~n26231 ;
  assign y19044 = n26233 ;
  assign y19045 = ~n26234 ;
  assign y19046 = ~n26237 ;
  assign y19047 = ~n26239 ;
  assign y19048 = n26242 ;
  assign y19049 = ~1'b0 ;
  assign y19050 = n26247 ;
  assign y19051 = ~n26251 ;
  assign y19052 = 1'b0 ;
  assign y19053 = ~1'b0 ;
  assign y19054 = ~n26255 ;
  assign y19055 = n26256 ;
  assign y19056 = n26257 ;
  assign y19057 = ~n3154 ;
  assign y19058 = ~1'b0 ;
  assign y19059 = n26259 ;
  assign y19060 = ~n3025 ;
  assign y19061 = n26262 ;
  assign y19062 = ~n26265 ;
  assign y19063 = ~1'b0 ;
  assign y19064 = ~n26277 ;
  assign y19065 = n26278 ;
  assign y19066 = ~1'b0 ;
  assign y19067 = ~1'b0 ;
  assign y19068 = ~1'b0 ;
  assign y19069 = ~1'b0 ;
  assign y19070 = ~1'b0 ;
  assign y19071 = ~n26281 ;
  assign y19072 = ~1'b0 ;
  assign y19073 = ~1'b0 ;
  assign y19074 = n26284 ;
  assign y19075 = n26290 ;
  assign y19076 = ~n26291 ;
  assign y19077 = n26293 ;
  assign y19078 = ~n11690 ;
  assign y19079 = ~n26296 ;
  assign y19080 = ~1'b0 ;
  assign y19081 = 1'b0 ;
  assign y19082 = ~1'b0 ;
  assign y19083 = ~1'b0 ;
  assign y19084 = ~n26299 ;
  assign y19085 = n20762 ;
  assign y19086 = ~n26301 ;
  assign y19087 = ~1'b0 ;
  assign y19088 = ~1'b0 ;
  assign y19089 = n26309 ;
  assign y19090 = n26310 ;
  assign y19091 = n26314 ;
  assign y19092 = ~n26315 ;
  assign y19093 = n26316 ;
  assign y19094 = ~n26318 ;
  assign y19095 = 1'b0 ;
  assign y19096 = n26320 ;
  assign y19097 = ~1'b0 ;
  assign y19098 = ~1'b0 ;
  assign y19099 = ~n26322 ;
  assign y19100 = ~n26323 ;
  assign y19101 = ~n26324 ;
  assign y19102 = ~1'b0 ;
  assign y19103 = ~1'b0 ;
  assign y19104 = ~1'b0 ;
  assign y19105 = n7497 ;
  assign y19106 = ~1'b0 ;
  assign y19107 = ~1'b0 ;
  assign y19108 = 1'b0 ;
  assign y19109 = ~1'b0 ;
  assign y19110 = ~1'b0 ;
  assign y19111 = ~n26326 ;
  assign y19112 = n26327 ;
  assign y19113 = n26329 ;
  assign y19114 = n26330 ;
  assign y19115 = ~1'b0 ;
  assign y19116 = ~1'b0 ;
  assign y19117 = ~1'b0 ;
  assign y19118 = ~n26333 ;
  assign y19119 = n26335 ;
  assign y19120 = ~n26337 ;
  assign y19121 = ~1'b0 ;
  assign y19122 = n22107 ;
  assign y19123 = ~n26339 ;
  assign y19124 = n607 ;
  assign y19125 = ~n26342 ;
  assign y19126 = ~n23788 ;
  assign y19127 = n26345 ;
  assign y19128 = n9670 ;
  assign y19129 = ~1'b0 ;
  assign y19130 = ~n26347 ;
  assign y19131 = n25324 ;
  assign y19132 = n26349 ;
  assign y19133 = n26350 ;
  assign y19134 = ~1'b0 ;
  assign y19135 = ~1'b0 ;
  assign y19136 = ~1'b0 ;
  assign y19137 = ~1'b0 ;
  assign y19138 = 1'b0 ;
  assign y19139 = ~n26356 ;
  assign y19140 = ~1'b0 ;
  assign y19141 = ~1'b0 ;
  assign y19142 = ~n26360 ;
  assign y19143 = n26365 ;
  assign y19144 = ~n26367 ;
  assign y19145 = ~1'b0 ;
  assign y19146 = ~1'b0 ;
  assign y19147 = ~1'b0 ;
  assign y19148 = ~n14403 ;
  assign y19149 = ~1'b0 ;
  assign y19150 = n25106 ;
  assign y19151 = ~n26370 ;
  assign y19152 = ~n26372 ;
  assign y19153 = ~1'b0 ;
  assign y19154 = ~1'b0 ;
  assign y19155 = ~1'b0 ;
  assign y19156 = ~1'b0 ;
  assign y19157 = ~1'b0 ;
  assign y19158 = n26375 ;
  assign y19159 = ~1'b0 ;
  assign y19160 = ~n16300 ;
  assign y19161 = ~1'b0 ;
  assign y19162 = n12657 ;
  assign y19163 = n26376 ;
  assign y19164 = ~1'b0 ;
  assign y19165 = n26377 ;
  assign y19166 = ~1'b0 ;
  assign y19167 = n26379 ;
  assign y19168 = ~n26380 ;
  assign y19169 = ~n26381 ;
  assign y19170 = n13953 ;
  assign y19171 = n20109 ;
  assign y19172 = ~1'b0 ;
  assign y19173 = ~n26387 ;
  assign y19174 = n24577 ;
  assign y19175 = ~1'b0 ;
  assign y19176 = ~1'b0 ;
  assign y19177 = n26390 ;
  assign y19178 = ~n26391 ;
  assign y19179 = n6037 ;
  assign y19180 = ~n26392 ;
  assign y19181 = ~1'b0 ;
  assign y19182 = ~n26394 ;
  assign y19183 = ~1'b0 ;
  assign y19184 = n26395 ;
  assign y19185 = n4299 ;
  assign y19186 = ~n10215 ;
  assign y19187 = ~1'b0 ;
  assign y19188 = n26399 ;
  assign y19189 = 1'b0 ;
  assign y19190 = ~n26402 ;
  assign y19191 = n11425 ;
  assign y19192 = ~1'b0 ;
  assign y19193 = ~n26407 ;
  assign y19194 = ~1'b0 ;
  assign y19195 = ~1'b0 ;
  assign y19196 = ~n26413 ;
  assign y19197 = 1'b0 ;
  assign y19198 = ~n26420 ;
  assign y19199 = ~n26421 ;
  assign y19200 = n19068 ;
  assign y19201 = ~n26423 ;
  assign y19202 = ~1'b0 ;
  assign y19203 = n26426 ;
  assign y19204 = ~n7736 ;
  assign y19205 = n26428 ;
  assign y19206 = n26434 ;
  assign y19207 = n26446 ;
  assign y19208 = 1'b0 ;
  assign y19209 = ~1'b0 ;
  assign y19210 = n26447 ;
  assign y19211 = ~1'b0 ;
  assign y19212 = 1'b0 ;
  assign y19213 = ~n26448 ;
  assign y19214 = ~1'b0 ;
  assign y19215 = ~1'b0 ;
  assign y19216 = ~1'b0 ;
  assign y19217 = ~n26450 ;
  assign y19218 = ~1'b0 ;
  assign y19219 = n26452 ;
  assign y19220 = ~n26462 ;
  assign y19221 = ~1'b0 ;
  assign y19222 = n26464 ;
  assign y19223 = ~1'b0 ;
  assign y19224 = n216 ;
  assign y19225 = n26466 ;
  assign y19226 = ~n495 ;
  assign y19227 = ~1'b0 ;
  assign y19228 = n26467 ;
  assign y19229 = ~n26468 ;
  assign y19230 = n26469 ;
  assign y19231 = ~n26471 ;
  assign y19232 = ~1'b0 ;
  assign y19233 = n26473 ;
  assign y19234 = ~n26474 ;
  assign y19235 = 1'b0 ;
  assign y19236 = ~n26475 ;
  assign y19237 = ~n26478 ;
  assign y19238 = ~n26479 ;
  assign y19239 = ~n26483 ;
  assign y19240 = ~n26486 ;
  assign y19241 = ~n26488 ;
  assign y19242 = n26489 ;
  assign y19243 = n26493 ;
  assign y19244 = ~1'b0 ;
  assign y19245 = n26497 ;
  assign y19246 = ~n15591 ;
  assign y19247 = ~n26500 ;
  assign y19248 = n26502 ;
  assign y19249 = ~n26505 ;
  assign y19250 = n26507 ;
  assign y19251 = ~1'b0 ;
  assign y19252 = ~1'b0 ;
  assign y19253 = ~1'b0 ;
  assign y19254 = n26510 ;
  assign y19255 = ~n26512 ;
  assign y19256 = n26513 ;
  assign y19257 = ~n1266 ;
  assign y19258 = ~1'b0 ;
  assign y19259 = ~1'b0 ;
  assign y19260 = ~1'b0 ;
  assign y19261 = ~n26516 ;
  assign y19262 = n26518 ;
  assign y19263 = ~n16834 ;
  assign y19264 = n26519 ;
  assign y19265 = ~1'b0 ;
  assign y19266 = n26520 ;
  assign y19267 = n1815 ;
  assign y19268 = ~1'b0 ;
  assign y19269 = ~1'b0 ;
  assign y19270 = n26523 ;
  assign y19271 = ~n26525 ;
  assign y19272 = 1'b0 ;
  assign y19273 = n26526 ;
  assign y19274 = n26528 ;
  assign y19275 = n26529 ;
  assign y19276 = ~n26530 ;
  assign y19277 = n26531 ;
  assign y19278 = 1'b0 ;
  assign y19279 = ~1'b0 ;
  assign y19280 = ~1'b0 ;
  assign y19281 = 1'b0 ;
  assign y19282 = n26532 ;
  assign y19283 = ~1'b0 ;
  assign y19284 = n26534 ;
  assign y19285 = ~1'b0 ;
  assign y19286 = ~1'b0 ;
  assign y19287 = ~1'b0 ;
  assign y19288 = n26538 ;
  assign y19289 = ~n26549 ;
  assign y19290 = ~n26550 ;
  assign y19291 = 1'b0 ;
  assign y19292 = 1'b0 ;
  assign y19293 = n7180 ;
  assign y19294 = ~1'b0 ;
  assign y19295 = ~n26551 ;
  assign y19296 = ~n26554 ;
  assign y19297 = ~1'b0 ;
  assign y19298 = ~1'b0 ;
  assign y19299 = ~n26555 ;
  assign y19300 = ~n26564 ;
  assign y19301 = ~1'b0 ;
  assign y19302 = ~n26565 ;
  assign y19303 = n11561 ;
  assign y19304 = n26567 ;
  assign y19305 = 1'b0 ;
  assign y19306 = n24370 ;
  assign y19307 = ~n26568 ;
  assign y19308 = ~1'b0 ;
  assign y19309 = ~n26571 ;
  assign y19310 = ~n26572 ;
  assign y19311 = ~n26573 ;
  assign y19312 = ~n26574 ;
  assign y19313 = ~n26583 ;
  assign y19314 = n3219 ;
  assign y19315 = ~1'b0 ;
  assign y19316 = ~1'b0 ;
  assign y19317 = ~n26589 ;
  assign y19318 = n26594 ;
  assign y19319 = ~n17564 ;
  assign y19320 = n26596 ;
  assign y19321 = ~n26597 ;
  assign y19322 = ~1'b0 ;
  assign y19323 = ~n26602 ;
  assign y19324 = n26609 ;
  assign y19325 = ~n26612 ;
  assign y19326 = ~1'b0 ;
  assign y19327 = n15481 ;
  assign y19328 = ~n26131 ;
  assign y19329 = ~1'b0 ;
  assign y19330 = ~1'b0 ;
  assign y19331 = n26614 ;
  assign y19332 = ~n26615 ;
  assign y19333 = ~n26616 ;
  assign y19334 = ~n16672 ;
  assign y19335 = ~1'b0 ;
  assign y19336 = ~n6525 ;
  assign y19337 = ~1'b0 ;
  assign y19338 = n26618 ;
  assign y19339 = ~1'b0 ;
  assign y19340 = n26621 ;
  assign y19341 = ~1'b0 ;
  assign y19342 = ~n26624 ;
  assign y19343 = ~n26625 ;
  assign y19344 = ~1'b0 ;
  assign y19345 = ~n26626 ;
  assign y19346 = ~n26628 ;
  assign y19347 = n980 ;
  assign y19348 = 1'b0 ;
  assign y19349 = n26632 ;
  assign y19350 = ~1'b0 ;
  assign y19351 = ~1'b0 ;
  assign y19352 = n26636 ;
  assign y19353 = ~n26637 ;
  assign y19354 = ~1'b0 ;
  assign y19355 = n26638 ;
  assign y19356 = ~n26639 ;
  assign y19357 = n26640 ;
  assign y19358 = ~n26642 ;
  assign y19359 = ~1'b0 ;
  assign y19360 = ~n26643 ;
  assign y19361 = n26645 ;
  assign y19362 = n26648 ;
  assign y19363 = ~n26650 ;
  assign y19364 = n26652 ;
  assign y19365 = ~1'b0 ;
  assign y19366 = n26659 ;
  assign y19367 = ~n26663 ;
  assign y19368 = n26666 ;
  assign y19369 = ~1'b0 ;
  assign y19370 = n8984 ;
  assign y19371 = ~1'b0 ;
  assign y19372 = ~n26668 ;
  assign y19373 = ~1'b0 ;
  assign y19374 = ~n26670 ;
  assign y19375 = ~n4720 ;
  assign y19376 = n26672 ;
  assign y19377 = ~1'b0 ;
  assign y19378 = ~1'b0 ;
  assign y19379 = n38 ;
  assign y19380 = ~n26673 ;
  assign y19381 = ~n26675 ;
  assign y19382 = n26678 ;
  assign y19383 = n26681 ;
  assign y19384 = ~1'b0 ;
  assign y19385 = ~1'b0 ;
  assign y19386 = n26683 ;
  assign y19387 = ~n10635 ;
  assign y19388 = 1'b0 ;
  assign y19389 = ~n19306 ;
  assign y19390 = ~n26685 ;
  assign y19391 = ~n26706 ;
  assign y19392 = ~1'b0 ;
  assign y19393 = ~n26707 ;
  assign y19394 = ~1'b0 ;
  assign y19395 = ~n26710 ;
  assign y19396 = n26712 ;
  assign y19397 = ~n26714 ;
  assign y19398 = ~n26718 ;
  assign y19399 = ~n26720 ;
  assign y19400 = ~1'b0 ;
  assign y19401 = ~n26725 ;
  assign y19402 = ~1'b0 ;
  assign y19403 = ~n26726 ;
  assign y19404 = ~1'b0 ;
  assign y19405 = ~1'b0 ;
  assign y19406 = ~n26729 ;
  assign y19407 = ~n26731 ;
  assign y19408 = ~1'b0 ;
  assign y19409 = ~n26732 ;
  assign y19410 = n26733 ;
  assign y19411 = ~1'b0 ;
  assign y19412 = n2078 ;
  assign y19413 = ~1'b0 ;
  assign y19414 = ~1'b0 ;
  assign y19415 = ~1'b0 ;
  assign y19416 = ~1'b0 ;
  assign y19417 = ~1'b0 ;
  assign y19418 = ~n13451 ;
  assign y19419 = n26738 ;
  assign y19420 = ~n26739 ;
  assign y19421 = ~n26740 ;
  assign y19422 = ~1'b0 ;
  assign y19423 = n12494 ;
  assign y19424 = ~1'b0 ;
  assign y19425 = ~n26741 ;
  assign y19426 = n26742 ;
  assign y19427 = ~n23910 ;
  assign y19428 = ~1'b0 ;
  assign y19429 = ~n26745 ;
  assign y19430 = ~n26747 ;
  assign y19431 = ~1'b0 ;
  assign y19432 = n26750 ;
  assign y19433 = n26754 ;
  assign y19434 = ~n5551 ;
  assign y19435 = ~n5397 ;
  assign y19436 = n26758 ;
  assign y19437 = ~n26765 ;
  assign y19438 = ~n26767 ;
  assign y19439 = n26770 ;
  assign y19440 = ~n26775 ;
  assign y19441 = n26776 ;
  assign y19442 = ~n8186 ;
  assign y19443 = n16745 ;
  assign y19444 = ~1'b0 ;
  assign y19445 = n26778 ;
  assign y19446 = ~1'b0 ;
  assign y19447 = n26782 ;
  assign y19448 = n26786 ;
  assign y19449 = n26787 ;
  assign y19450 = ~n26790 ;
  assign y19451 = 1'b0 ;
  assign y19452 = n26791 ;
  assign y19453 = n26792 ;
  assign y19454 = n26795 ;
  assign y19455 = n26803 ;
  assign y19456 = ~n26804 ;
  assign y19457 = n26825 ;
  assign y19458 = ~n310 ;
  assign y19459 = ~n8648 ;
  assign y19460 = 1'b0 ;
  assign y19461 = ~1'b0 ;
  assign y19462 = n26826 ;
  assign y19463 = n26827 ;
  assign y19464 = ~n26829 ;
  assign y19465 = n26830 ;
  assign y19466 = ~1'b0 ;
  assign y19467 = ~1'b0 ;
  assign y19468 = ~1'b0 ;
  assign y19469 = ~n26833 ;
  assign y19470 = ~1'b0 ;
  assign y19471 = ~n26835 ;
  assign y19472 = n26836 ;
  assign y19473 = ~1'b0 ;
  assign y19474 = ~1'b0 ;
  assign y19475 = n26837 ;
  assign y19476 = ~n26838 ;
  assign y19477 = n26842 ;
  assign y19478 = n26845 ;
  assign y19479 = ~1'b0 ;
  assign y19480 = ~n26847 ;
  assign y19481 = ~n332 ;
  assign y19482 = ~n26849 ;
  assign y19483 = ~n26851 ;
  assign y19484 = n23477 ;
  assign y19485 = n26852 ;
  assign y19486 = ~1'b0 ;
  assign y19487 = ~1'b0 ;
  assign y19488 = ~n26853 ;
  assign y19489 = ~n26856 ;
  assign y19490 = n26857 ;
  assign y19491 = ~1'b0 ;
  assign y19492 = n26858 ;
  assign y19493 = ~n5182 ;
  assign y19494 = ~1'b0 ;
  assign y19495 = ~n175 ;
  assign y19496 = ~1'b0 ;
  assign y19497 = n26859 ;
  assign y19498 = ~1'b0 ;
  assign y19499 = ~n26862 ;
  assign y19500 = ~n23894 ;
  assign y19501 = n26863 ;
  assign y19502 = n26876 ;
  assign y19503 = n26877 ;
  assign y19504 = n26879 ;
  assign y19505 = ~n26881 ;
  assign y19506 = n26882 ;
  assign y19507 = n26883 ;
  assign y19508 = ~1'b0 ;
  assign y19509 = ~1'b0 ;
  assign y19510 = ~1'b0 ;
  assign y19511 = ~n26885 ;
  assign y19512 = ~1'b0 ;
  assign y19513 = ~n6689 ;
  assign y19514 = ~n20621 ;
  assign y19515 = n869 ;
  assign y19516 = ~1'b0 ;
  assign y19517 = n9372 ;
  assign y19518 = ~1'b0 ;
  assign y19519 = 1'b0 ;
  assign y19520 = ~n26886 ;
  assign y19521 = ~n6009 ;
  assign y19522 = 1'b0 ;
  assign y19523 = ~1'b0 ;
  assign y19524 = ~n26889 ;
  assign y19525 = 1'b0 ;
  assign y19526 = ~1'b0 ;
  assign y19527 = 1'b0 ;
  assign y19528 = ~1'b0 ;
  assign y19529 = ~1'b0 ;
  assign y19530 = 1'b0 ;
  assign y19531 = ~1'b0 ;
  assign y19532 = ~1'b0 ;
  assign y19533 = 1'b0 ;
  assign y19534 = ~n13917 ;
  assign y19535 = n26895 ;
  assign y19536 = ~n26897 ;
  assign y19537 = n1017 ;
  assign y19538 = ~1'b0 ;
  assign y19539 = ~n26899 ;
  assign y19540 = ~1'b0 ;
  assign y19541 = n11656 ;
  assign y19542 = n26900 ;
  assign y19543 = ~n26901 ;
  assign y19544 = ~n23355 ;
  assign y19545 = ~1'b0 ;
  assign y19546 = ~n2784 ;
  assign y19547 = n26902 ;
  assign y19548 = ~n14694 ;
  assign y19549 = ~n26904 ;
  assign y19550 = ~n26905 ;
  assign y19551 = n26907 ;
  assign y19552 = n26912 ;
  assign y19553 = ~1'b0 ;
  assign y19554 = n26915 ;
  assign y19555 = ~n26920 ;
  assign y19556 = ~1'b0 ;
  assign y19557 = ~1'b0 ;
  assign y19558 = ~1'b0 ;
  assign y19559 = n26926 ;
  assign y19560 = ~n26932 ;
  assign y19561 = ~n26936 ;
  assign y19562 = n26942 ;
  assign y19563 = n26944 ;
  assign y19564 = ~n26945 ;
  assign y19565 = ~1'b0 ;
  assign y19566 = n26946 ;
  assign y19567 = n26948 ;
  assign y19568 = ~1'b0 ;
  assign y19569 = 1'b0 ;
  assign y19570 = ~n17008 ;
  assign y19571 = ~n26950 ;
  assign y19572 = ~n26953 ;
  assign y19573 = n26957 ;
  assign y19574 = ~1'b0 ;
  assign y19575 = ~n26958 ;
  assign y19576 = n26959 ;
  assign y19577 = ~n26961 ;
  assign y19578 = ~1'b0 ;
  assign y19579 = ~n26963 ;
  assign y19580 = ~n26970 ;
  assign y19581 = n26975 ;
  assign y19582 = n19171 ;
  assign y19583 = ~n26976 ;
  assign y19584 = n26979 ;
  assign y19585 = n6882 ;
  assign y19586 = ~n26980 ;
  assign y19587 = ~1'b0 ;
  assign y19588 = ~1'b0 ;
  assign y19589 = ~1'b0 ;
  assign y19590 = ~n26982 ;
  assign y19591 = n14393 ;
  assign y19592 = n26983 ;
  assign y19593 = n26984 ;
  assign y19594 = ~n26988 ;
  assign y19595 = ~1'b0 ;
  assign y19596 = n26989 ;
  assign y19597 = ~1'b0 ;
  assign y19598 = ~n26990 ;
  assign y19599 = ~1'b0 ;
  assign y19600 = ~n11018 ;
  assign y19601 = ~1'b0 ;
  assign y19602 = n26991 ;
  assign y19603 = ~1'b0 ;
  assign y19604 = ~1'b0 ;
  assign y19605 = ~1'b0 ;
  assign y19606 = ~n26999 ;
  assign y19607 = ~n27005 ;
  assign y19608 = n27006 ;
  assign y19609 = n27007 ;
  assign y19610 = ~n27009 ;
  assign y19611 = n27010 ;
  assign y19612 = n27013 ;
  assign y19613 = ~1'b0 ;
  assign y19614 = 1'b0 ;
  assign y19615 = ~n27015 ;
  assign y19616 = n27016 ;
  assign y19617 = 1'b0 ;
  assign y19618 = n27018 ;
  assign y19619 = n27022 ;
  assign y19620 = ~n27025 ;
  assign y19621 = ~n12777 ;
  assign y19622 = ~n27031 ;
  assign y19623 = n27034 ;
  assign y19624 = n15983 ;
  assign y19625 = n27037 ;
  assign y19626 = ~1'b0 ;
  assign y19627 = ~n27059 ;
  assign y19628 = ~1'b0 ;
  assign y19629 = n27061 ;
  assign y19630 = ~1'b0 ;
  assign y19631 = ~n27065 ;
  assign y19632 = n8231 ;
  assign y19633 = n27071 ;
  assign y19634 = n27075 ;
  assign y19635 = n27076 ;
  assign y19636 = ~1'b0 ;
  assign y19637 = ~1'b0 ;
  assign y19638 = ~1'b0 ;
  assign y19639 = ~1'b0 ;
  assign y19640 = ~1'b0 ;
  assign y19641 = ~1'b0 ;
  assign y19642 = n27077 ;
  assign y19643 = ~1'b0 ;
  assign y19644 = ~n27078 ;
  assign y19645 = ~1'b0 ;
  assign y19646 = ~n27081 ;
  assign y19647 = ~n27082 ;
  assign y19648 = ~1'b0 ;
  assign y19649 = ~1'b0 ;
  assign y19650 = ~1'b0 ;
  assign y19651 = ~1'b0 ;
  assign y19652 = ~1'b0 ;
  assign y19653 = n27083 ;
  assign y19654 = ~1'b0 ;
  assign y19655 = n7231 ;
  assign y19656 = n27086 ;
  assign y19657 = n27088 ;
  assign y19658 = ~n27089 ;
  assign y19659 = ~1'b0 ;
  assign y19660 = ~n27091 ;
  assign y19661 = n27092 ;
  assign y19662 = ~1'b0 ;
  assign y19663 = ~n23735 ;
  assign y19664 = ~1'b0 ;
  assign y19665 = ~1'b0 ;
  assign y19666 = n27093 ;
  assign y19667 = n27094 ;
  assign y19668 = ~1'b0 ;
  assign y19669 = n27095 ;
  assign y19670 = ~n27102 ;
  assign y19671 = ~n27103 ;
  assign y19672 = ~1'b0 ;
  assign y19673 = ~1'b0 ;
  assign y19674 = ~1'b0 ;
  assign y19675 = ~n8446 ;
  assign y19676 = ~1'b0 ;
  assign y19677 = n27105 ;
  assign y19678 = n27106 ;
  assign y19679 = n27108 ;
  assign y19680 = ~n27109 ;
  assign y19681 = n27110 ;
  assign y19682 = ~1'b0 ;
  assign y19683 = ~n27114 ;
  assign y19684 = ~n27117 ;
  assign y19685 = ~1'b0 ;
  assign y19686 = ~n27120 ;
  assign y19687 = ~n27123 ;
  assign y19688 = n27126 ;
  assign y19689 = ~1'b0 ;
  assign y19690 = ~1'b0 ;
  assign y19691 = ~n27128 ;
  assign y19692 = ~1'b0 ;
  assign y19693 = ~1'b0 ;
  assign y19694 = ~n27129 ;
  assign y19695 = ~n27135 ;
  assign y19696 = ~n27136 ;
  assign y19697 = ~1'b0 ;
  assign y19698 = n27138 ;
  assign y19699 = ~1'b0 ;
  assign y19700 = ~1'b0 ;
  assign y19701 = n27139 ;
  assign y19702 = ~1'b0 ;
  assign y19703 = ~n27140 ;
  assign y19704 = ~1'b0 ;
  assign y19705 = ~n27144 ;
  assign y19706 = n27145 ;
  assign y19707 = ~1'b0 ;
  assign y19708 = ~n27146 ;
  assign y19709 = ~n27153 ;
  assign y19710 = ~1'b0 ;
  assign y19711 = n27156 ;
  assign y19712 = ~1'b0 ;
  assign y19713 = ~n27164 ;
  assign y19714 = ~1'b0 ;
  assign y19715 = n27167 ;
  assign y19716 = n27168 ;
  assign y19717 = ~1'b0 ;
  assign y19718 = ~1'b0 ;
  assign y19719 = ~1'b0 ;
  assign y19720 = ~1'b0 ;
  assign y19721 = ~n27170 ;
  assign y19722 = n27171 ;
  assign y19723 = n27172 ;
  assign y19724 = ~1'b0 ;
  assign y19725 = n27173 ;
  assign y19726 = ~n14411 ;
  assign y19727 = ~n27175 ;
  assign y19728 = ~1'b0 ;
  assign y19729 = n27177 ;
  assign y19730 = ~1'b0 ;
  assign y19731 = ~1'b0 ;
  assign y19732 = ~n2611 ;
  assign y19733 = n24684 ;
  assign y19734 = ~1'b0 ;
  assign y19735 = n27178 ;
  assign y19736 = ~n27186 ;
  assign y19737 = ~n27187 ;
  assign y19738 = n27188 ;
  assign y19739 = ~1'b0 ;
  assign y19740 = n27192 ;
  assign y19741 = ~1'b0 ;
  assign y19742 = ~n27193 ;
  assign y19743 = ~n24106 ;
  assign y19744 = ~n27200 ;
  assign y19745 = ~n27203 ;
  assign y19746 = ~n27207 ;
  assign y19747 = n27209 ;
  assign y19748 = n27212 ;
  assign y19749 = n27213 ;
  assign y19750 = ~1'b0 ;
  assign y19751 = n27217 ;
  assign y19752 = ~1'b0 ;
  assign y19753 = ~n27224 ;
  assign y19754 = ~1'b0 ;
  assign y19755 = 1'b0 ;
  assign y19756 = n27226 ;
  assign y19757 = ~n27230 ;
  assign y19758 = ~n27235 ;
  assign y19759 = ~1'b0 ;
  assign y19760 = ~1'b0 ;
  assign y19761 = 1'b0 ;
  assign y19762 = ~n5206 ;
  assign y19763 = ~n27236 ;
  assign y19764 = ~n27240 ;
  assign y19765 = ~n27242 ;
  assign y19766 = ~1'b0 ;
  assign y19767 = ~1'b0 ;
  assign y19768 = ~n27244 ;
  assign y19769 = ~1'b0 ;
  assign y19770 = ~n20736 ;
  assign y19771 = n27249 ;
  assign y19772 = 1'b0 ;
  assign y19773 = ~1'b0 ;
  assign y19774 = ~1'b0 ;
  assign y19775 = n27251 ;
  assign y19776 = ~1'b0 ;
  assign y19777 = n9942 ;
  assign y19778 = ~n27255 ;
  assign y19779 = ~1'b0 ;
  assign y19780 = ~1'b0 ;
  assign y19781 = n27256 ;
  assign y19782 = ~1'b0 ;
  assign y19783 = ~n27257 ;
  assign y19784 = n27259 ;
  assign y19785 = ~1'b0 ;
  assign y19786 = ~1'b0 ;
  assign y19787 = n60 ;
  assign y19788 = ~1'b0 ;
  assign y19789 = n27260 ;
  assign y19790 = ~1'b0 ;
  assign y19791 = 1'b0 ;
  assign y19792 = n27266 ;
  assign y19793 = n27270 ;
  assign y19794 = ~n27271 ;
  assign y19795 = n2194 ;
  assign y19796 = ~n27272 ;
  assign y19797 = ~n27277 ;
  assign y19798 = 1'b0 ;
  assign y19799 = ~1'b0 ;
  assign y19800 = ~1'b0 ;
  assign y19801 = n27278 ;
  assign y19802 = 1'b0 ;
  assign y19803 = ~n27279 ;
  assign y19804 = ~1'b0 ;
  assign y19805 = ~1'b0 ;
  assign y19806 = n17989 ;
  assign y19807 = n27281 ;
  assign y19808 = n27287 ;
  assign y19809 = ~n27288 ;
  assign y19810 = n17285 ;
  assign y19811 = ~n27296 ;
  assign y19812 = ~1'b0 ;
  assign y19813 = n27297 ;
  assign y19814 = ~1'b0 ;
  assign y19815 = ~1'b0 ;
  assign y19816 = ~n3307 ;
  assign y19817 = n10743 ;
  assign y19818 = ~n18156 ;
  assign y19819 = ~1'b0 ;
  assign y19820 = ~1'b0 ;
  assign y19821 = ~1'b0 ;
  assign y19822 = ~1'b0 ;
  assign y19823 = ~1'b0 ;
  assign y19824 = n27298 ;
  assign y19825 = ~n27300 ;
  assign y19826 = ~1'b0 ;
  assign y19827 = n1396 ;
  assign y19828 = ~1'b0 ;
  assign y19829 = ~n27301 ;
  assign y19830 = ~n7029 ;
  assign y19831 = ~1'b0 ;
  assign y19832 = n27302 ;
  assign y19833 = ~1'b0 ;
  assign y19834 = ~1'b0 ;
  assign y19835 = ~n27306 ;
  assign y19836 = ~1'b0 ;
  assign y19837 = ~1'b0 ;
  assign y19838 = ~n27310 ;
  assign y19839 = ~n27311 ;
  assign y19840 = ~n27313 ;
  assign y19841 = n27314 ;
  assign y19842 = ~1'b0 ;
  assign y19843 = ~n27315 ;
  assign y19844 = 1'b0 ;
  assign y19845 = n27316 ;
  assign y19846 = ~1'b0 ;
  assign y19847 = ~n20700 ;
  assign y19848 = ~n27318 ;
  assign y19849 = ~n18403 ;
  assign y19850 = ~1'b0 ;
  assign y19851 = ~n27320 ;
  assign y19852 = ~1'b0 ;
  assign y19853 = n27323 ;
  assign y19854 = n20076 ;
  assign y19855 = n23237 ;
  assign y19856 = n27325 ;
  assign y19857 = ~1'b0 ;
  assign y19858 = n27326 ;
  assign y19859 = n27327 ;
  assign y19860 = 1'b0 ;
  assign y19861 = ~n27328 ;
  assign y19862 = ~1'b0 ;
  assign y19863 = ~n27329 ;
  assign y19864 = ~1'b0 ;
  assign y19865 = ~n27330 ;
  assign y19866 = n330 ;
  assign y19867 = ~1'b0 ;
  assign y19868 = n27333 ;
  assign y19869 = n27334 ;
  assign y19870 = n27339 ;
  assign y19871 = ~1'b0 ;
  assign y19872 = ~n27340 ;
  assign y19873 = ~n27342 ;
  assign y19874 = ~1'b0 ;
  assign y19875 = ~1'b0 ;
  assign y19876 = ~n27344 ;
  assign y19877 = n27347 ;
  assign y19878 = ~n27350 ;
  assign y19879 = ~1'b0 ;
  assign y19880 = ~1'b0 ;
  assign y19881 = ~n27352 ;
  assign y19882 = 1'b0 ;
  assign y19883 = ~1'b0 ;
  assign y19884 = 1'b0 ;
  assign y19885 = ~1'b0 ;
  assign y19886 = n27353 ;
  assign y19887 = n27354 ;
  assign y19888 = ~1'b0 ;
  assign y19889 = n6185 ;
  assign y19890 = ~1'b0 ;
  assign y19891 = n27355 ;
  assign y19892 = n27356 ;
  assign y19893 = 1'b0 ;
  assign y19894 = ~1'b0 ;
  assign y19895 = ~n27357 ;
  assign y19896 = ~n27359 ;
  assign y19897 = n27361 ;
  assign y19898 = ~n27003 ;
  assign y19899 = ~1'b0 ;
  assign y19900 = ~n27366 ;
  assign y19901 = n27368 ;
  assign y19902 = ~n27370 ;
  assign y19903 = ~1'b0 ;
  assign y19904 = ~1'b0 ;
  assign y19905 = ~n27372 ;
  assign y19906 = ~1'b0 ;
  assign y19907 = n19870 ;
  assign y19908 = n27374 ;
  assign y19909 = ~n27375 ;
  assign y19910 = ~1'b0 ;
  assign y19911 = n27382 ;
  assign y19912 = n27385 ;
  assign y19913 = n27386 ;
  assign y19914 = ~1'b0 ;
  assign y19915 = ~1'b0 ;
  assign y19916 = n1995 ;
  assign y19917 = ~1'b0 ;
  assign y19918 = n27388 ;
  assign y19919 = ~n11067 ;
  assign y19920 = ~1'b0 ;
  assign y19921 = ~n6295 ;
  assign y19922 = ~n27389 ;
  assign y19923 = ~1'b0 ;
  assign y19924 = ~n27393 ;
  assign y19925 = ~1'b0 ;
  assign y19926 = ~1'b0 ;
  assign y19927 = ~n27395 ;
  assign y19928 = ~1'b0 ;
  assign y19929 = n27399 ;
  assign y19930 = ~1'b0 ;
  assign y19931 = ~n512 ;
  assign y19932 = 1'b0 ;
  assign y19933 = ~1'b0 ;
  assign y19934 = ~1'b0 ;
  assign y19935 = 1'b0 ;
  assign y19936 = n27403 ;
  assign y19937 = n27405 ;
  assign y19938 = ~n27406 ;
  assign y19939 = ~1'b0 ;
  assign y19940 = 1'b0 ;
  assign y19941 = ~1'b0 ;
  assign y19942 = ~1'b0 ;
  assign y19943 = 1'b0 ;
  assign y19944 = ~1'b0 ;
  assign y19945 = n27407 ;
  assign y19946 = ~n27410 ;
  assign y19947 = ~1'b0 ;
  assign y19948 = ~1'b0 ;
  assign y19949 = ~n27411 ;
  assign y19950 = ~1'b0 ;
  assign y19951 = ~n3735 ;
  assign y19952 = ~1'b0 ;
  assign y19953 = n27412 ;
  assign y19954 = ~1'b0 ;
  assign y19955 = n27413 ;
  assign y19956 = ~1'b0 ;
  assign y19957 = n27416 ;
  assign y19958 = n5393 ;
  assign y19959 = ~1'b0 ;
  assign y19960 = ~n27419 ;
  assign y19961 = n27422 ;
  assign y19962 = ~1'b0 ;
  assign y19963 = ~1'b0 ;
  assign y19964 = n27425 ;
  assign y19965 = ~1'b0 ;
  assign y19966 = n27426 ;
  assign y19967 = ~n27429 ;
  assign y19968 = 1'b0 ;
  assign y19969 = ~1'b0 ;
  assign y19970 = ~1'b0 ;
  assign y19971 = ~n18776 ;
  assign y19972 = ~1'b0 ;
  assign y19973 = ~1'b0 ;
  assign y19974 = ~1'b0 ;
  assign y19975 = ~n27440 ;
  assign y19976 = n27443 ;
  assign y19977 = ~n25397 ;
  assign y19978 = n27449 ;
  assign y19979 = ~n8198 ;
  assign y19980 = n27451 ;
  assign y19981 = ~n27452 ;
  assign y19982 = n27456 ;
  assign y19983 = ~n18460 ;
  assign y19984 = ~1'b0 ;
  assign y19985 = ~n27463 ;
  assign y19986 = ~1'b0 ;
  assign y19987 = ~n27466 ;
  assign y19988 = n8019 ;
  assign y19989 = 1'b0 ;
  assign y19990 = ~n27468 ;
  assign y19991 = n27469 ;
  assign y19992 = ~1'b0 ;
  assign y19993 = ~n27472 ;
  assign y19994 = ~1'b0 ;
  assign y19995 = ~1'b0 ;
  assign y19996 = n27478 ;
  assign y19997 = ~1'b0 ;
  assign y19998 = n19710 ;
  assign y19999 = n27479 ;
  assign y20000 = ~n27481 ;
  assign y20001 = n27484 ;
  assign y20002 = n27488 ;
  assign y20003 = ~n27489 ;
  assign y20004 = ~1'b0 ;
  assign y20005 = ~1'b0 ;
  assign y20006 = ~n27494 ;
  assign y20007 = ~n27497 ;
  assign y20008 = ~1'b0 ;
  assign y20009 = n27499 ;
  assign y20010 = ~n27501 ;
  assign y20011 = ~n27503 ;
  assign y20012 = n27504 ;
  assign y20013 = ~1'b0 ;
  assign y20014 = ~n14904 ;
  assign y20015 = n27505 ;
  assign y20016 = ~n27507 ;
  assign y20017 = n27508 ;
  assign y20018 = ~1'b0 ;
  assign y20019 = ~1'b0 ;
  assign y20020 = n27517 ;
  assign y20021 = n27518 ;
  assign y20022 = ~1'b0 ;
  assign y20023 = ~1'b0 ;
  assign y20024 = ~n27523 ;
  assign y20025 = ~n27524 ;
  assign y20026 = ~n21468 ;
  assign y20027 = ~1'b0 ;
  assign y20028 = n27527 ;
  assign y20029 = ~1'b0 ;
  assign y20030 = n27528 ;
  assign y20031 = n27530 ;
  assign y20032 = ~1'b0 ;
  assign y20033 = ~1'b0 ;
  assign y20034 = ~1'b0 ;
  assign y20035 = n27532 ;
  assign y20036 = ~n27534 ;
  assign y20037 = ~n27539 ;
  assign y20038 = ~n27541 ;
  assign y20039 = ~1'b0 ;
  assign y20040 = n27542 ;
  assign y20041 = ~n14435 ;
  assign y20042 = ~1'b0 ;
  assign y20043 = n27544 ;
  assign y20044 = 1'b0 ;
  assign y20045 = n27546 ;
  assign y20046 = 1'b0 ;
  assign y20047 = ~n27548 ;
  assign y20048 = ~n27549 ;
  assign y20049 = n3287 ;
  assign y20050 = n1802 ;
  assign y20051 = n27554 ;
  assign y20052 = n17049 ;
  assign y20053 = n23783 ;
  assign y20054 = n27555 ;
  assign y20055 = ~1'b0 ;
  assign y20056 = ~1'b0 ;
  assign y20057 = ~n27556 ;
  assign y20058 = n14590 ;
  assign y20059 = ~1'b0 ;
  assign y20060 = n27557 ;
  assign y20061 = ~1'b0 ;
  assign y20062 = n27561 ;
  assign y20063 = n27562 ;
  assign y20064 = n27567 ;
  assign y20065 = ~1'b0 ;
  assign y20066 = n27573 ;
  assign y20067 = ~n27575 ;
  assign y20068 = ~n27577 ;
  assign y20069 = n23894 ;
  assign y20070 = n27578 ;
  assign y20071 = n6176 ;
  assign y20072 = ~n27579 ;
  assign y20073 = ~1'b0 ;
  assign y20074 = ~1'b0 ;
  assign y20075 = ~n27581 ;
  assign y20076 = ~n27583 ;
  assign y20077 = n27586 ;
  assign y20078 = ~1'b0 ;
  assign y20079 = ~1'b0 ;
  assign y20080 = n27592 ;
  assign y20081 = ~n27594 ;
  assign y20082 = ~1'b0 ;
  assign y20083 = ~1'b0 ;
  assign y20084 = ~n27596 ;
  assign y20085 = ~1'b0 ;
  assign y20086 = ~1'b0 ;
  assign y20087 = ~1'b0 ;
  assign y20088 = ~n27597 ;
  assign y20089 = ~1'b0 ;
  assign y20090 = ~n27599 ;
  assign y20091 = ~n27600 ;
  assign y20092 = ~n27603 ;
  assign y20093 = ~n27608 ;
  assign y20094 = ~n27609 ;
  assign y20095 = ~n27612 ;
  assign y20096 = ~n27614 ;
  assign y20097 = ~n27617 ;
  assign y20098 = ~1'b0 ;
  assign y20099 = ~n27618 ;
  assign y20100 = ~n27626 ;
  assign y20101 = ~n6464 ;
  assign y20102 = 1'b0 ;
  assign y20103 = n7606 ;
  assign y20104 = n27628 ;
  assign y20105 = ~n27633 ;
  assign y20106 = n27637 ;
  assign y20107 = n27638 ;
  assign y20108 = n22835 ;
  assign y20109 = 1'b0 ;
  assign y20110 = n27642 ;
  assign y20111 = n27643 ;
  assign y20112 = ~1'b0 ;
  assign y20113 = ~1'b0 ;
  assign y20114 = ~1'b0 ;
  assign y20115 = n27644 ;
  assign y20116 = ~n27646 ;
  assign y20117 = ~1'b0 ;
  assign y20118 = ~n27651 ;
  assign y20119 = n2278 ;
  assign y20120 = ~1'b0 ;
  assign y20121 = ~n27652 ;
  assign y20122 = ~1'b0 ;
  assign y20123 = ~n27653 ;
  assign y20124 = ~n27654 ;
  assign y20125 = ~n27656 ;
  assign y20126 = n8198 ;
  assign y20127 = n27657 ;
  assign y20128 = n144 ;
  assign y20129 = ~n27659 ;
  assign y20130 = ~1'b0 ;
  assign y20131 = ~n27661 ;
  assign y20132 = n27669 ;
  assign y20133 = n257 ;
  assign y20134 = ~n9134 ;
  assign y20135 = ~n7108 ;
  assign y20136 = ~n27673 ;
  assign y20137 = ~n27675 ;
  assign y20138 = ~n17950 ;
  assign y20139 = ~1'b0 ;
  assign y20140 = n27678 ;
  assign y20141 = ~n27683 ;
  assign y20142 = 1'b0 ;
  assign y20143 = ~n27684 ;
  assign y20144 = n19333 ;
  assign y20145 = ~n27685 ;
  assign y20146 = n27686 ;
  assign y20147 = n27689 ;
  assign y20148 = n27690 ;
  assign y20149 = ~n27691 ;
  assign y20150 = ~1'b0 ;
  assign y20151 = ~1'b0 ;
  assign y20152 = ~1'b0 ;
  assign y20153 = n27693 ;
  assign y20154 = n27694 ;
  assign y20155 = ~1'b0 ;
  assign y20156 = n27696 ;
  assign y20157 = ~1'b0 ;
  assign y20158 = ~1'b0 ;
  assign y20159 = n27698 ;
  assign y20160 = ~n27699 ;
  assign y20161 = ~n27700 ;
  assign y20162 = n17935 ;
  assign y20163 = n27703 ;
  assign y20164 = ~n27706 ;
  assign y20165 = n27708 ;
  assign y20166 = ~1'b0 ;
  assign y20167 = ~1'b0 ;
  assign y20168 = ~1'b0 ;
  assign y20169 = n27716 ;
  assign y20170 = ~n27718 ;
  assign y20171 = ~1'b0 ;
  assign y20172 = ~1'b0 ;
  assign y20173 = ~n27720 ;
  assign y20174 = ~n27723 ;
  assign y20175 = 1'b0 ;
  assign y20176 = ~1'b0 ;
  assign y20177 = 1'b0 ;
  assign y20178 = ~1'b0 ;
  assign y20179 = n27725 ;
  assign y20180 = n27732 ;
  assign y20181 = ~n27734 ;
  assign y20182 = ~1'b0 ;
  assign y20183 = ~1'b0 ;
  assign y20184 = n27735 ;
  assign y20185 = n27739 ;
  assign y20186 = ~1'b0 ;
  assign y20187 = ~1'b0 ;
  assign y20188 = ~n27741 ;
  assign y20189 = ~n27743 ;
  assign y20190 = n27745 ;
  assign y20191 = n27749 ;
  assign y20192 = ~1'b0 ;
  assign y20193 = ~1'b0 ;
  assign y20194 = ~n27752 ;
  assign y20195 = ~1'b0 ;
  assign y20196 = ~n24678 ;
  assign y20197 = n27753 ;
  assign y20198 = ~n27756 ;
  assign y20199 = ~1'b0 ;
  assign y20200 = ~1'b0 ;
  assign y20201 = ~1'b0 ;
  assign y20202 = ~n10617 ;
  assign y20203 = ~1'b0 ;
  assign y20204 = 1'b0 ;
  assign y20205 = n27761 ;
  assign y20206 = ~n27762 ;
  assign y20207 = ~n27764 ;
  assign y20208 = ~1'b0 ;
  assign y20209 = ~1'b0 ;
  assign y20210 = n27767 ;
  assign y20211 = ~1'b0 ;
  assign y20212 = n27769 ;
  assign y20213 = ~1'b0 ;
  assign y20214 = ~n27771 ;
  assign y20215 = ~n27772 ;
  assign y20216 = ~1'b0 ;
  assign y20217 = n27773 ;
  assign y20218 = n1243 ;
  assign y20219 = ~1'b0 ;
  assign y20220 = ~1'b0 ;
  assign y20221 = n27774 ;
  assign y20222 = n5465 ;
  assign y20223 = ~n20264 ;
  assign y20224 = ~n16613 ;
  assign y20225 = ~1'b0 ;
  assign y20226 = n27776 ;
  assign y20227 = n27777 ;
  assign y20228 = ~1'b0 ;
  assign y20229 = ~n27780 ;
  assign y20230 = n27782 ;
  assign y20231 = ~n27783 ;
  assign y20232 = ~n27785 ;
  assign y20233 = ~1'b0 ;
  assign y20234 = n27788 ;
  assign y20235 = ~n27791 ;
  assign y20236 = n27792 ;
  assign y20237 = ~n27793 ;
  assign y20238 = n15259 ;
  assign y20239 = ~n27795 ;
  assign y20240 = ~n27796 ;
  assign y20241 = ~1'b0 ;
  assign y20242 = ~n2176 ;
  assign y20243 = ~1'b0 ;
  assign y20244 = 1'b0 ;
  assign y20245 = n24840 ;
  assign y20246 = ~1'b0 ;
  assign y20247 = n27799 ;
  assign y20248 = ~n27800 ;
  assign y20249 = ~1'b0 ;
  assign y20250 = n27805 ;
  assign y20251 = ~n27809 ;
  assign y20252 = ~1'b0 ;
  assign y20253 = ~n27810 ;
  assign y20254 = ~n22418 ;
  assign y20255 = n18932 ;
  assign y20256 = ~1'b0 ;
  assign y20257 = ~1'b0 ;
  assign y20258 = ~1'b0 ;
  assign y20259 = ~1'b0 ;
  assign y20260 = n27812 ;
  assign y20261 = n27813 ;
  assign y20262 = ~n27814 ;
  assign y20263 = ~1'b0 ;
  assign y20264 = ~n27815 ;
  assign y20265 = ~1'b0 ;
  assign y20266 = n27817 ;
  assign y20267 = ~n27818 ;
  assign y20268 = n27820 ;
  assign y20269 = ~1'b0 ;
  assign y20270 = ~1'b0 ;
  assign y20271 = ~1'b0 ;
  assign y20272 = 1'b0 ;
  assign y20273 = n27824 ;
  assign y20274 = ~1'b0 ;
  assign y20275 = n27826 ;
  assign y20276 = ~n27828 ;
  assign y20277 = ~1'b0 ;
  assign y20278 = ~n2578 ;
  assign y20279 = n27829 ;
  assign y20280 = n7713 ;
  assign y20281 = n27830 ;
  assign y20282 = ~n27833 ;
  assign y20283 = ~1'b0 ;
  assign y20284 = n27839 ;
  assign y20285 = ~1'b0 ;
  assign y20286 = n27840 ;
  assign y20287 = ~n27842 ;
  assign y20288 = n27845 ;
  assign y20289 = ~n27846 ;
  assign y20290 = n27848 ;
  assign y20291 = n27849 ;
  assign y20292 = ~n27850 ;
  assign y20293 = ~n27852 ;
  assign y20294 = n27853 ;
  assign y20295 = ~1'b0 ;
  assign y20296 = 1'b0 ;
  assign y20297 = n27855 ;
  assign y20298 = ~1'b0 ;
  assign y20299 = n2342 ;
  assign y20300 = ~1'b0 ;
  assign y20301 = n27856 ;
  assign y20302 = ~1'b0 ;
  assign y20303 = n27857 ;
  assign y20304 = ~n27859 ;
  assign y20305 = ~n27860 ;
  assign y20306 = ~1'b0 ;
  assign y20307 = ~1'b0 ;
  assign y20308 = ~n27862 ;
  assign y20309 = ~n27866 ;
  assign y20310 = ~1'b0 ;
  assign y20311 = ~1'b0 ;
  assign y20312 = ~1'b0 ;
  assign y20313 = n27871 ;
  assign y20314 = ~n27874 ;
  assign y20315 = n4797 ;
  assign y20316 = ~1'b0 ;
  assign y20317 = ~1'b0 ;
  assign y20318 = ~n27875 ;
  assign y20319 = ~1'b0 ;
  assign y20320 = ~1'b0 ;
  assign y20321 = n27877 ;
  assign y20322 = ~n27878 ;
  assign y20323 = ~n27880 ;
  assign y20324 = ~n7945 ;
  assign y20325 = ~n27881 ;
  assign y20326 = ~1'b0 ;
  assign y20327 = ~n27883 ;
  assign y20328 = ~1'b0 ;
  assign y20329 = ~1'b0 ;
  assign y20330 = n27884 ;
  assign y20331 = 1'b0 ;
  assign y20332 = n27890 ;
  assign y20333 = ~1'b0 ;
  assign y20334 = ~1'b0 ;
  assign y20335 = ~n27891 ;
  assign y20336 = n27893 ;
  assign y20337 = ~n27894 ;
  assign y20338 = n27895 ;
  assign y20339 = ~1'b0 ;
  assign y20340 = ~1'b0 ;
  assign y20341 = n27897 ;
  assign y20342 = ~1'b0 ;
  assign y20343 = ~1'b0 ;
  assign y20344 = ~1'b0 ;
  assign y20345 = n27898 ;
  assign y20346 = ~n27904 ;
  assign y20347 = n27906 ;
  assign y20348 = ~n1833 ;
  assign y20349 = ~1'b0 ;
  assign y20350 = ~n15262 ;
  assign y20351 = n27907 ;
  assign y20352 = n27910 ;
  assign y20353 = ~n27911 ;
  assign y20354 = ~n27913 ;
  assign y20355 = n27915 ;
  assign y20356 = ~1'b0 ;
  assign y20357 = 1'b0 ;
  assign y20358 = n27916 ;
  assign y20359 = ~n27919 ;
  assign y20360 = n27920 ;
  assign y20361 = ~n27924 ;
  assign y20362 = ~n27926 ;
  assign y20363 = ~n12764 ;
  assign y20364 = ~n27930 ;
  assign y20365 = n1193 ;
  assign y20366 = ~1'b0 ;
  assign y20367 = ~n27932 ;
  assign y20368 = ~1'b0 ;
  assign y20369 = ~n27936 ;
  assign y20370 = ~1'b0 ;
  assign y20371 = ~n27937 ;
  assign y20372 = ~n27938 ;
  assign y20373 = ~n27939 ;
  assign y20374 = n27940 ;
  assign y20375 = n27941 ;
  assign y20376 = n27942 ;
  assign y20377 = ~1'b0 ;
  assign y20378 = n27945 ;
  assign y20379 = ~1'b0 ;
  assign y20380 = ~1'b0 ;
  assign y20381 = ~n27949 ;
  assign y20382 = ~1'b0 ;
  assign y20383 = ~n27950 ;
  assign y20384 = ~n27952 ;
  assign y20385 = ~1'b0 ;
  assign y20386 = ~1'b0 ;
  assign y20387 = n14232 ;
  assign y20388 = n27954 ;
  assign y20389 = n27955 ;
  assign y20390 = n27956 ;
  assign y20391 = ~1'b0 ;
  assign y20392 = n27958 ;
  assign y20393 = n1915 ;
  assign y20394 = ~n27959 ;
  assign y20395 = ~n27962 ;
  assign y20396 = n27965 ;
  assign y20397 = ~1'b0 ;
  assign y20398 = n14272 ;
  assign y20399 = ~1'b0 ;
  assign y20400 = ~1'b0 ;
  assign y20401 = ~1'b0 ;
  assign y20402 = ~1'b0 ;
  assign y20403 = ~1'b0 ;
  assign y20404 = ~n27971 ;
  assign y20405 = ~1'b0 ;
  assign y20406 = ~n27974 ;
  assign y20407 = n24146 ;
  assign y20408 = 1'b0 ;
  assign y20409 = ~n27976 ;
  assign y20410 = ~n27978 ;
  assign y20411 = ~n27981 ;
  assign y20412 = ~1'b0 ;
  assign y20413 = n25118 ;
  assign y20414 = n27985 ;
  assign y20415 = n27986 ;
  assign y20416 = ~1'b0 ;
  assign y20417 = ~1'b0 ;
  assign y20418 = n27988 ;
  assign y20419 = ~n27990 ;
  assign y20420 = n27991 ;
  assign y20421 = ~1'b0 ;
  assign y20422 = ~1'b0 ;
  assign y20423 = 1'b0 ;
  assign y20424 = ~1'b0 ;
  assign y20425 = ~n27992 ;
  assign y20426 = ~n22204 ;
  assign y20427 = 1'b0 ;
  assign y20428 = ~1'b0 ;
  assign y20429 = ~n2725 ;
  assign y20430 = n27997 ;
  assign y20431 = ~n28000 ;
  assign y20432 = ~n9213 ;
  assign y20433 = ~n28001 ;
  assign y20434 = ~1'b0 ;
  assign y20435 = ~1'b0 ;
  assign y20436 = 1'b0 ;
  assign y20437 = n28002 ;
  assign y20438 = ~1'b0 ;
  assign y20439 = ~n635 ;
  assign y20440 = n28004 ;
  assign y20441 = ~n28008 ;
  assign y20442 = ~1'b0 ;
  assign y20443 = n28009 ;
  assign y20444 = n28011 ;
  assign y20445 = ~n28013 ;
  assign y20446 = ~1'b0 ;
  assign y20447 = n24313 ;
  assign y20448 = ~1'b0 ;
  assign y20449 = ~1'b0 ;
  assign y20450 = ~1'b0 ;
  assign y20451 = n28015 ;
  assign y20452 = ~1'b0 ;
  assign y20453 = ~n28016 ;
  assign y20454 = ~1'b0 ;
  assign y20455 = ~1'b0 ;
  assign y20456 = ~n28025 ;
  assign y20457 = ~1'b0 ;
  assign y20458 = n28029 ;
  assign y20459 = n28032 ;
  assign y20460 = n28034 ;
  assign y20461 = ~n28035 ;
  assign y20462 = n28040 ;
  assign y20463 = ~1'b0 ;
  assign y20464 = n28043 ;
  assign y20465 = ~n28044 ;
  assign y20466 = ~1'b0 ;
  assign y20467 = ~1'b0 ;
  assign y20468 = 1'b0 ;
  assign y20469 = n28045 ;
  assign y20470 = ~n28046 ;
  assign y20471 = n5603 ;
  assign y20472 = ~1'b0 ;
  assign y20473 = ~1'b0 ;
  assign y20474 = n28048 ;
  assign y20475 = ~n28049 ;
  assign y20476 = n28052 ;
  assign y20477 = ~n28053 ;
  assign y20478 = ~1'b0 ;
  assign y20479 = n28057 ;
  assign y20480 = ~n28058 ;
  assign y20481 = ~1'b0 ;
  assign y20482 = 1'b0 ;
  assign y20483 = n28059 ;
  assign y20484 = n28061 ;
  assign y20485 = ~1'b0 ;
  assign y20486 = n28064 ;
  assign y20487 = ~1'b0 ;
  assign y20488 = 1'b0 ;
  assign y20489 = ~1'b0 ;
  assign y20490 = ~1'b0 ;
  assign y20491 = ~n28065 ;
  assign y20492 = ~1'b0 ;
  assign y20493 = ~n28067 ;
  assign y20494 = ~n28068 ;
  assign y20495 = n28069 ;
  assign y20496 = ~1'b0 ;
  assign y20497 = ~n28070 ;
  assign y20498 = ~1'b0 ;
  assign y20499 = n3138 ;
  assign y20500 = ~1'b0 ;
  assign y20501 = ~n28072 ;
  assign y20502 = ~1'b0 ;
  assign y20503 = ~1'b0 ;
  assign y20504 = n28077 ;
  assign y20505 = ~n28078 ;
  assign y20506 = 1'b0 ;
  assign y20507 = ~n28081 ;
  assign y20508 = n28082 ;
  assign y20509 = ~n28084 ;
  assign y20510 = ~1'b0 ;
  assign y20511 = ~n3718 ;
  assign y20512 = ~n11946 ;
  assign y20513 = ~1'b0 ;
  assign y20514 = ~n28085 ;
  assign y20515 = ~n28086 ;
  assign y20516 = ~n28087 ;
  assign y20517 = ~n28092 ;
  assign y20518 = n28093 ;
  assign y20519 = 1'b0 ;
  assign y20520 = ~1'b0 ;
  assign y20521 = ~1'b0 ;
  assign y20522 = ~n3833 ;
  assign y20523 = ~n28095 ;
  assign y20524 = ~1'b0 ;
  assign y20525 = ~n28097 ;
  assign y20526 = n28099 ;
  assign y20527 = 1'b0 ;
  assign y20528 = ~n28101 ;
  assign y20529 = n28102 ;
  assign y20530 = ~n9692 ;
  assign y20531 = 1'b0 ;
  assign y20532 = ~1'b0 ;
  assign y20533 = n28103 ;
  assign y20534 = ~1'b0 ;
  assign y20535 = ~1'b0 ;
  assign y20536 = n823 ;
  assign y20537 = n13408 ;
  assign y20538 = n28105 ;
  assign y20539 = ~1'b0 ;
  assign y20540 = n28106 ;
  assign y20541 = n28107 ;
  assign y20542 = n28110 ;
  assign y20543 = ~1'b0 ;
  assign y20544 = n28111 ;
  assign y20545 = n28124 ;
  assign y20546 = ~1'b0 ;
  assign y20547 = n2430 ;
  assign y20548 = ~1'b0 ;
  assign y20549 = ~n28126 ;
  assign y20550 = n28128 ;
  assign y20551 = ~1'b0 ;
  assign y20552 = ~n28134 ;
  assign y20553 = ~n28138 ;
  assign y20554 = ~n28141 ;
  assign y20555 = ~n28144 ;
  assign y20556 = ~1'b0 ;
  assign y20557 = ~n28145 ;
  assign y20558 = 1'b0 ;
  assign y20559 = ~1'b0 ;
  assign y20560 = ~n28148 ;
  assign y20561 = ~n3946 ;
  assign y20562 = ~n12053 ;
  assign y20563 = n11582 ;
  assign y20564 = n28149 ;
  assign y20565 = ~n28151 ;
  assign y20566 = n28152 ;
  assign y20567 = ~n28155 ;
  assign y20568 = ~1'b0 ;
  assign y20569 = ~n28157 ;
  assign y20570 = ~n28159 ;
  assign y20571 = n28163 ;
  assign y20572 = ~1'b0 ;
  assign y20573 = ~1'b0 ;
  assign y20574 = ~n28166 ;
  assign y20575 = ~1'b0 ;
  assign y20576 = ~1'b0 ;
  assign y20577 = ~n28168 ;
  assign y20578 = ~n28169 ;
  assign y20579 = ~1'b0 ;
  assign y20580 = n18144 ;
  assign y20581 = n28171 ;
  assign y20582 = ~1'b0 ;
  assign y20583 = ~n12177 ;
  assign y20584 = ~n28172 ;
  assign y20585 = ~1'b0 ;
  assign y20586 = ~1'b0 ;
  assign y20587 = ~1'b0 ;
  assign y20588 = n16199 ;
  assign y20589 = ~1'b0 ;
  assign y20590 = ~n28173 ;
  assign y20591 = ~n28176 ;
  assign y20592 = n28177 ;
  assign y20593 = ~1'b0 ;
  assign y20594 = n28178 ;
  assign y20595 = n22387 ;
  assign y20596 = ~1'b0 ;
  assign y20597 = ~n6992 ;
  assign y20598 = ~n28179 ;
  assign y20599 = ~1'b0 ;
  assign y20600 = ~1'b0 ;
  assign y20601 = ~n28182 ;
  assign y20602 = 1'b0 ;
  assign y20603 = ~n28183 ;
  assign y20604 = n28184 ;
  assign y20605 = n28186 ;
  assign y20606 = ~1'b0 ;
  assign y20607 = ~n28188 ;
  assign y20608 = ~n28190 ;
  assign y20609 = ~1'b0 ;
  assign y20610 = n28192 ;
  assign y20611 = ~1'b0 ;
  assign y20612 = ~n28197 ;
  assign y20613 = ~n28198 ;
  assign y20614 = ~1'b0 ;
  assign y20615 = ~1'b0 ;
  assign y20616 = ~n28203 ;
  assign y20617 = n28205 ;
  assign y20618 = ~1'b0 ;
  assign y20619 = ~1'b0 ;
  assign y20620 = ~n28208 ;
  assign y20621 = n28211 ;
  assign y20622 = ~n28217 ;
  assign y20623 = ~1'b0 ;
  assign y20624 = ~n28220 ;
  assign y20625 = ~1'b0 ;
  assign y20626 = ~n28221 ;
  assign y20627 = ~1'b0 ;
  assign y20628 = ~1'b0 ;
  assign y20629 = ~n28222 ;
  assign y20630 = ~n710 ;
  assign y20631 = ~1'b0 ;
  assign y20632 = ~1'b0 ;
  assign y20633 = ~n14813 ;
  assign y20634 = n28224 ;
  assign y20635 = ~n28225 ;
  assign y20636 = n3131 ;
  assign y20637 = ~n28226 ;
  assign y20638 = ~1'b0 ;
  assign y20639 = ~1'b0 ;
  assign y20640 = 1'b0 ;
  assign y20641 = n28227 ;
  assign y20642 = ~n28228 ;
  assign y20643 = ~1'b0 ;
  assign y20644 = ~n28230 ;
  assign y20645 = ~n3803 ;
  assign y20646 = n28231 ;
  assign y20647 = ~1'b0 ;
  assign y20648 = 1'b0 ;
  assign y20649 = n28234 ;
  assign y20650 = n28237 ;
  assign y20651 = ~1'b0 ;
  assign y20652 = n28240 ;
  assign y20653 = ~1'b0 ;
  assign y20654 = ~1'b0 ;
  assign y20655 = ~1'b0 ;
  assign y20656 = ~n28241 ;
  assign y20657 = ~n28242 ;
  assign y20658 = n28243 ;
  assign y20659 = ~1'b0 ;
  assign y20660 = ~n28247 ;
  assign y20661 = n1471 ;
  assign y20662 = ~1'b0 ;
  assign y20663 = n7523 ;
  assign y20664 = ~1'b0 ;
  assign y20665 = ~n28250 ;
  assign y20666 = ~n28253 ;
  assign y20667 = n28255 ;
  assign y20668 = n28256 ;
  assign y20669 = n25874 ;
  assign y20670 = ~n28257 ;
  assign y20671 = ~n4700 ;
  assign y20672 = ~n28258 ;
  assign y20673 = n28262 ;
  assign y20674 = ~1'b0 ;
  assign y20675 = ~1'b0 ;
  assign y20676 = n28264 ;
  assign y20677 = n28267 ;
  assign y20678 = ~n28269 ;
  assign y20679 = n1194 ;
  assign y20680 = ~n28270 ;
  assign y20681 = ~1'b0 ;
  assign y20682 = ~1'b0 ;
  assign y20683 = ~n28271 ;
  assign y20684 = n28272 ;
  assign y20685 = n28274 ;
  assign y20686 = ~1'b0 ;
  assign y20687 = 1'b0 ;
  assign y20688 = 1'b0 ;
  assign y20689 = n28275 ;
  assign y20690 = ~n28278 ;
  assign y20691 = ~n28280 ;
  assign y20692 = ~n9885 ;
  assign y20693 = ~1'b0 ;
  assign y20694 = n9561 ;
  assign y20695 = n28284 ;
  assign y20696 = ~1'b0 ;
  assign y20697 = n28285 ;
  assign y20698 = n28288 ;
  assign y20699 = ~n28289 ;
  assign y20700 = ~n28291 ;
  assign y20701 = n28293 ;
  assign y20702 = ~1'b0 ;
  assign y20703 = ~n28297 ;
  assign y20704 = ~1'b0 ;
  assign y20705 = ~1'b0 ;
  assign y20706 = n28302 ;
  assign y20707 = ~1'b0 ;
  assign y20708 = ~1'b0 ;
  assign y20709 = ~1'b0 ;
  assign y20710 = n28304 ;
  assign y20711 = ~1'b0 ;
  assign y20712 = ~1'b0 ;
  assign y20713 = ~1'b0 ;
  assign y20714 = n28306 ;
  assign y20715 = ~n28310 ;
  assign y20716 = ~n28311 ;
  assign y20717 = ~1'b0 ;
  assign y20718 = n28312 ;
  assign y20719 = ~1'b0 ;
  assign y20720 = ~n28314 ;
  assign y20721 = ~n28318 ;
  assign y20722 = ~1'b0 ;
  assign y20723 = ~n11167 ;
  assign y20724 = ~1'b0 ;
  assign y20725 = ~1'b0 ;
  assign y20726 = ~n8397 ;
  assign y20727 = ~1'b0 ;
  assign y20728 = ~n28320 ;
  assign y20729 = ~1'b0 ;
  assign y20730 = ~n28321 ;
  assign y20731 = ~n13776 ;
  assign y20732 = n28325 ;
  assign y20733 = ~1'b0 ;
  assign y20734 = n4668 ;
  assign y20735 = n28329 ;
  assign y20736 = ~1'b0 ;
  assign y20737 = ~n12028 ;
  assign y20738 = n28332 ;
  assign y20739 = ~1'b0 ;
  assign y20740 = ~1'b0 ;
  assign y20741 = ~n28335 ;
  assign y20742 = ~n28337 ;
  assign y20743 = ~1'b0 ;
  assign y20744 = n28339 ;
  assign y20745 = ~1'b0 ;
  assign y20746 = n13065 ;
  assign y20747 = ~n28347 ;
  assign y20748 = ~1'b0 ;
  assign y20749 = ~1'b0 ;
  assign y20750 = ~1'b0 ;
  assign y20751 = ~1'b0 ;
  assign y20752 = ~1'b0 ;
  assign y20753 = ~n28358 ;
  assign y20754 = ~n28359 ;
  assign y20755 = n28361 ;
  assign y20756 = n133 ;
  assign y20757 = n28362 ;
  assign y20758 = ~1'b0 ;
  assign y20759 = ~n28364 ;
  assign y20760 = ~n28367 ;
  assign y20761 = ~1'b0 ;
  assign y20762 = ~1'b0 ;
  assign y20763 = ~n28368 ;
  assign y20764 = n28369 ;
  assign y20765 = ~1'b0 ;
  assign y20766 = 1'b0 ;
  assign y20767 = ~1'b0 ;
  assign y20768 = n28373 ;
  assign y20769 = ~n28374 ;
  assign y20770 = ~1'b0 ;
  assign y20771 = ~1'b0 ;
  assign y20772 = 1'b0 ;
  assign y20773 = n28377 ;
  assign y20774 = ~n28378 ;
  assign y20775 = ~1'b0 ;
  assign y20776 = ~1'b0 ;
  assign y20777 = n28380 ;
  assign y20778 = n28382 ;
  assign y20779 = ~n28383 ;
  assign y20780 = ~n28385 ;
  assign y20781 = ~n28387 ;
  assign y20782 = n28388 ;
  assign y20783 = ~1'b0 ;
  assign y20784 = n28393 ;
  assign y20785 = ~1'b0 ;
  assign y20786 = ~n2601 ;
  assign y20787 = ~n28395 ;
  assign y20788 = ~1'b0 ;
  assign y20789 = ~n28396 ;
  assign y20790 = 1'b0 ;
  assign y20791 = ~n8792 ;
  assign y20792 = n28397 ;
  assign y20793 = ~1'b0 ;
  assign y20794 = n28398 ;
  assign y20795 = ~1'b0 ;
  assign y20796 = ~n28404 ;
  assign y20797 = ~n28405 ;
  assign y20798 = ~1'b0 ;
  assign y20799 = n28407 ;
  assign y20800 = n28409 ;
  assign y20801 = ~n28413 ;
  assign y20802 = ~1'b0 ;
  assign y20803 = ~1'b0 ;
  assign y20804 = n28415 ;
  assign y20805 = ~1'b0 ;
  assign y20806 = ~n28416 ;
  assign y20807 = ~n11462 ;
  assign y20808 = n28419 ;
  assign y20809 = 1'b0 ;
  assign y20810 = ~n28420 ;
  assign y20811 = n28421 ;
  assign y20812 = ~n28422 ;
  assign y20813 = ~n28423 ;
  assign y20814 = n28424 ;
  assign y20815 = ~n7667 ;
  assign y20816 = ~1'b0 ;
  assign y20817 = ~1'b0 ;
  assign y20818 = n28428 ;
  assign y20819 = ~1'b0 ;
  assign y20820 = ~n28429 ;
  assign y20821 = ~1'b0 ;
  assign y20822 = ~1'b0 ;
  assign y20823 = ~n13527 ;
  assign y20824 = 1'b0 ;
  assign y20825 = ~n23326 ;
  assign y20826 = ~n28433 ;
  assign y20827 = ~n28441 ;
  assign y20828 = n28443 ;
  assign y20829 = n6254 ;
  assign y20830 = ~n28444 ;
  assign y20831 = ~1'b0 ;
  assign y20832 = ~n28445 ;
  assign y20833 = ~1'b0 ;
  assign y20834 = n28486 ;
  assign y20835 = 1'b0 ;
  assign y20836 = n28489 ;
  assign y20837 = ~1'b0 ;
  assign y20838 = ~n28492 ;
  assign y20839 = ~1'b0 ;
  assign y20840 = ~n28493 ;
  assign y20841 = ~1'b0 ;
  assign y20842 = ~1'b0 ;
  assign y20843 = n28495 ;
  assign y20844 = ~1'b0 ;
  assign y20845 = ~n28496 ;
  assign y20846 = n15688 ;
  assign y20847 = ~1'b0 ;
  assign y20848 = n28498 ;
  assign y20849 = ~1'b0 ;
  assign y20850 = 1'b0 ;
  assign y20851 = ~1'b0 ;
  assign y20852 = ~1'b0 ;
  assign y20853 = ~n28499 ;
  assign y20854 = n2949 ;
  assign y20855 = n28501 ;
  assign y20856 = ~n28507 ;
  assign y20857 = ~1'b0 ;
  assign y20858 = n9327 ;
  assign y20859 = ~1'b0 ;
  assign y20860 = n28509 ;
  assign y20861 = ~1'b0 ;
  assign y20862 = ~1'b0 ;
  assign y20863 = ~1'b0 ;
  assign y20864 = ~1'b0 ;
  assign y20865 = n28513 ;
  assign y20866 = ~n17635 ;
  assign y20867 = ~n28521 ;
  assign y20868 = ~1'b0 ;
  assign y20869 = ~1'b0 ;
  assign y20870 = ~n28522 ;
  assign y20871 = ~n28524 ;
  assign y20872 = ~n1602 ;
  assign y20873 = ~1'b0 ;
  assign y20874 = ~1'b0 ;
  assign y20875 = ~n28529 ;
  assign y20876 = ~1'b0 ;
  assign y20877 = n28531 ;
  assign y20878 = ~1'b0 ;
  assign y20879 = n28535 ;
  assign y20880 = ~n28536 ;
  assign y20881 = ~n28540 ;
  assign y20882 = n28541 ;
  assign y20883 = ~1'b0 ;
  assign y20884 = ~n28542 ;
  assign y20885 = ~n28546 ;
  assign y20886 = ~n28548 ;
  assign y20887 = n28549 ;
  assign y20888 = ~1'b0 ;
  assign y20889 = ~1'b0 ;
  assign y20890 = ~n28552 ;
  assign y20891 = ~1'b0 ;
  assign y20892 = ~n28555 ;
  assign y20893 = ~n16289 ;
  assign y20894 = ~n28559 ;
  assign y20895 = ~n28561 ;
  assign y20896 = ~n28562 ;
  assign y20897 = ~n28563 ;
  assign y20898 = ~1'b0 ;
  assign y20899 = ~1'b0 ;
  assign y20900 = ~n28564 ;
  assign y20901 = n28565 ;
  assign y20902 = ~1'b0 ;
  assign y20903 = 1'b0 ;
  assign y20904 = n27783 ;
  assign y20905 = n28583 ;
  assign y20906 = ~1'b0 ;
  assign y20907 = ~n28586 ;
  assign y20908 = ~n28587 ;
  assign y20909 = n28598 ;
  assign y20910 = ~1'b0 ;
  assign y20911 = ~1'b0 ;
  assign y20912 = ~1'b0 ;
  assign y20913 = ~1'b0 ;
  assign y20914 = ~n27572 ;
  assign y20915 = ~n28602 ;
  assign y20916 = ~n28605 ;
  assign y20917 = n28253 ;
  assign y20918 = ~n28609 ;
  assign y20919 = ~n28611 ;
  assign y20920 = ~1'b0 ;
  assign y20921 = ~n28614 ;
  assign y20922 = ~n28616 ;
  assign y20923 = ~1'b0 ;
  assign y20924 = ~1'b0 ;
  assign y20925 = ~n5542 ;
  assign y20926 = n28617 ;
  assign y20927 = n28619 ;
  assign y20928 = 1'b0 ;
  assign y20929 = ~1'b0 ;
  assign y20930 = ~n28621 ;
  assign y20931 = n28624 ;
  assign y20932 = n14537 ;
  assign y20933 = ~1'b0 ;
  assign y20934 = ~1'b0 ;
  assign y20935 = ~1'b0 ;
  assign y20936 = n28625 ;
  assign y20937 = n28626 ;
  assign y20938 = ~n28628 ;
  assign y20939 = ~1'b0 ;
  assign y20940 = 1'b0 ;
  assign y20941 = n26153 ;
  assign y20942 = ~1'b0 ;
  assign y20943 = ~n28630 ;
  assign y20944 = ~1'b0 ;
  assign y20945 = n28633 ;
  assign y20946 = ~n28634 ;
  assign y20947 = ~1'b0 ;
  assign y20948 = ~n28635 ;
  assign y20949 = n28637 ;
  assign y20950 = ~1'b0 ;
  assign y20951 = ~1'b0 ;
  assign y20952 = ~1'b0 ;
  assign y20953 = ~n28640 ;
  assign y20954 = ~n28641 ;
  assign y20955 = ~n28642 ;
  assign y20956 = n28645 ;
  assign y20957 = ~1'b0 ;
  assign y20958 = ~1'b0 ;
  assign y20959 = ~n28646 ;
  assign y20960 = n28647 ;
  assign y20961 = n28648 ;
  assign y20962 = 1'b0 ;
  assign y20963 = 1'b0 ;
  assign y20964 = ~n20197 ;
  assign y20965 = ~1'b0 ;
  assign y20966 = ~1'b0 ;
  assign y20967 = n28649 ;
  assign y20968 = ~n28651 ;
  assign y20969 = ~1'b0 ;
  assign y20970 = ~n28654 ;
  assign y20971 = ~1'b0 ;
  assign y20972 = ~1'b0 ;
  assign y20973 = n28656 ;
  assign y20974 = ~1'b0 ;
  assign y20975 = n28658 ;
  assign y20976 = n28660 ;
  assign y20977 = ~n28661 ;
  assign y20978 = ~n1990 ;
  assign y20979 = n104 ;
  assign y20980 = ~1'b0 ;
  assign y20981 = ~n28668 ;
  assign y20982 = ~n28669 ;
  assign y20983 = 1'b0 ;
  assign y20984 = ~1'b0 ;
  assign y20985 = ~1'b0 ;
  assign y20986 = ~1'b0 ;
  assign y20987 = n28670 ;
  assign y20988 = ~1'b0 ;
  assign y20989 = n14834 ;
  assign y20990 = n28671 ;
  assign y20991 = n28672 ;
  assign y20992 = ~1'b0 ;
  assign y20993 = ~n28678 ;
  assign y20994 = n9111 ;
  assign y20995 = ~n28680 ;
  assign y20996 = n28682 ;
  assign y20997 = ~1'b0 ;
  assign y20998 = n28684 ;
  assign y20999 = ~1'b0 ;
  assign y21000 = n28685 ;
  assign y21001 = ~1'b0 ;
  assign y21002 = ~n28687 ;
  assign y21003 = n28689 ;
  assign y21004 = n28694 ;
  assign y21005 = ~1'b0 ;
  assign y21006 = n28695 ;
  assign y21007 = ~n28698 ;
  assign y21008 = n28717 ;
  assign y21009 = ~n28718 ;
  assign y21010 = ~n28719 ;
  assign y21011 = ~n28720 ;
  assign y21012 = n28721 ;
  assign y21013 = ~n28722 ;
  assign y21014 = n28725 ;
  assign y21015 = ~1'b0 ;
  assign y21016 = ~n28727 ;
  assign y21017 = ~1'b0 ;
  assign y21018 = n28728 ;
  assign y21019 = ~n28731 ;
  assign y21020 = ~n28735 ;
  assign y21021 = ~n28737 ;
  assign y21022 = ~1'b0 ;
  assign y21023 = n28739 ;
  assign y21024 = ~1'b0 ;
  assign y21025 = ~n28740 ;
  assign y21026 = ~n25671 ;
  assign y21027 = n28741 ;
  assign y21028 = ~n28749 ;
  assign y21029 = ~n28751 ;
  assign y21030 = ~1'b0 ;
  assign y21031 = n28752 ;
  assign y21032 = ~1'b0 ;
  assign y21033 = ~1'b0 ;
  assign y21034 = ~1'b0 ;
  assign y21035 = ~n28753 ;
  assign y21036 = ~1'b0 ;
  assign y21037 = ~1'b0 ;
  assign y21038 = ~1'b0 ;
  assign y21039 = ~n28754 ;
  assign y21040 = n28755 ;
  assign y21041 = n28759 ;
  assign y21042 = ~n28765 ;
  assign y21043 = ~n24909 ;
  assign y21044 = ~n28769 ;
  assign y21045 = n28771 ;
  assign y21046 = ~n1950 ;
  assign y21047 = ~n28773 ;
  assign y21048 = ~n28777 ;
  assign y21049 = ~1'b0 ;
  assign y21050 = ~1'b0 ;
  assign y21051 = ~1'b0 ;
  assign y21052 = ~1'b0 ;
  assign y21053 = ~1'b0 ;
  assign y21054 = ~1'b0 ;
  assign y21055 = ~1'b0 ;
  assign y21056 = n20342 ;
  assign y21057 = n23611 ;
  assign y21058 = n28780 ;
  assign y21059 = ~n15549 ;
  assign y21060 = ~1'b0 ;
  assign y21061 = ~1'b0 ;
  assign y21062 = n28783 ;
  assign y21063 = ~1'b0 ;
  assign y21064 = ~n28785 ;
  assign y21065 = n28802 ;
  assign y21066 = ~1'b0 ;
  assign y21067 = ~1'b0 ;
  assign y21068 = ~1'b0 ;
  assign y21069 = ~1'b0 ;
  assign y21070 = ~1'b0 ;
  assign y21071 = ~1'b0 ;
  assign y21072 = ~n7181 ;
  assign y21073 = ~n28806 ;
  assign y21074 = ~1'b0 ;
  assign y21075 = ~n28808 ;
  assign y21076 = ~n28810 ;
  assign y21077 = ~1'b0 ;
  assign y21078 = ~n28811 ;
  assign y21079 = ~1'b0 ;
  assign y21080 = n28813 ;
  assign y21081 = ~1'b0 ;
  assign y21082 = ~n28814 ;
  assign y21083 = ~1'b0 ;
  assign y21084 = ~n28817 ;
  assign y21085 = ~n28821 ;
  assign y21086 = n28824 ;
  assign y21087 = n28828 ;
  assign y21088 = ~1'b0 ;
  assign y21089 = ~1'b0 ;
  assign y21090 = 1'b0 ;
  assign y21091 = ~1'b0 ;
  assign y21092 = ~n23566 ;
  assign y21093 = ~n28832 ;
  assign y21094 = ~1'b0 ;
  assign y21095 = ~1'b0 ;
  assign y21096 = n28835 ;
  assign y21097 = ~1'b0 ;
  assign y21098 = ~n28838 ;
  assign y21099 = ~n28839 ;
  assign y21100 = ~1'b0 ;
  assign y21101 = 1'b0 ;
  assign y21102 = ~1'b0 ;
  assign y21103 = ~n28842 ;
  assign y21104 = ~1'b0 ;
  assign y21105 = n28843 ;
  assign y21106 = ~n28844 ;
  assign y21107 = ~1'b0 ;
  assign y21108 = ~n13034 ;
  assign y21109 = n28846 ;
  assign y21110 = n5424 ;
  assign y21111 = ~n28849 ;
  assign y21112 = n28852 ;
  assign y21113 = ~1'b0 ;
  assign y21114 = ~1'b0 ;
  assign y21115 = n28856 ;
  assign y21116 = n28858 ;
  assign y21117 = ~1'b0 ;
  assign y21118 = n28860 ;
  assign y21119 = ~1'b0 ;
  assign y21120 = ~1'b0 ;
  assign y21121 = ~1'b0 ;
  assign y21122 = ~1'b0 ;
  assign y21123 = ~1'b0 ;
  assign y21124 = n4840 ;
  assign y21125 = ~1'b0 ;
  assign y21126 = n1766 ;
  assign y21127 = ~1'b0 ;
  assign y21128 = ~1'b0 ;
  assign y21129 = ~n18873 ;
  assign y21130 = ~n28863 ;
  assign y21131 = ~n28865 ;
  assign y21132 = n28869 ;
  assign y21133 = ~n28870 ;
  assign y21134 = ~1'b0 ;
  assign y21135 = ~n12922 ;
  assign y21136 = ~1'b0 ;
  assign y21137 = ~1'b0 ;
  assign y21138 = n28872 ;
  assign y21139 = ~n28874 ;
  assign y21140 = n28875 ;
  assign y21141 = n28877 ;
  assign y21142 = n28878 ;
  assign y21143 = ~n28885 ;
  assign y21144 = ~n28887 ;
  assign y21145 = n28890 ;
  assign y21146 = ~1'b0 ;
  assign y21147 = ~n14805 ;
  assign y21148 = ~1'b0 ;
  assign y21149 = ~1'b0 ;
  assign y21150 = ~1'b0 ;
  assign y21151 = n28891 ;
  assign y21152 = n14670 ;
  assign y21153 = ~n28896 ;
  assign y21154 = n28897 ;
  assign y21155 = ~1'b0 ;
  assign y21156 = n28899 ;
  assign y21157 = ~n28900 ;
  assign y21158 = ~1'b0 ;
  assign y21159 = ~1'b0 ;
  assign y21160 = ~1'b0 ;
  assign y21161 = ~1'b0 ;
  assign y21162 = n28901 ;
  assign y21163 = ~1'b0 ;
  assign y21164 = ~n28902 ;
  assign y21165 = n28904 ;
  assign y21166 = ~n28905 ;
  assign y21167 = ~n28908 ;
  assign y21168 = ~n28909 ;
  assign y21169 = ~1'b0 ;
  assign y21170 = ~1'b0 ;
  assign y21171 = ~1'b0 ;
  assign y21172 = ~n5493 ;
  assign y21173 = ~n28911 ;
  assign y21174 = ~1'b0 ;
  assign y21175 = ~1'b0 ;
  assign y21176 = ~1'b0 ;
  assign y21177 = ~n28912 ;
  assign y21178 = ~n15707 ;
  assign y21179 = ~n28913 ;
  assign y21180 = ~1'b0 ;
  assign y21181 = n28914 ;
  assign y21182 = ~1'b0 ;
  assign y21183 = ~n28921 ;
  assign y21184 = ~n28924 ;
  assign y21185 = ~n28926 ;
  assign y21186 = ~1'b0 ;
  assign y21187 = n28928 ;
  assign y21188 = ~1'b0 ;
  assign y21189 = n28929 ;
  assign y21190 = ~n28930 ;
  assign y21191 = n28934 ;
  assign y21192 = ~n28938 ;
  assign y21193 = ~n25493 ;
  assign y21194 = ~n28939 ;
  assign y21195 = ~1'b0 ;
  assign y21196 = ~n2223 ;
  assign y21197 = ~n28940 ;
  assign y21198 = ~1'b0 ;
  assign y21199 = ~n28942 ;
  assign y21200 = ~n28945 ;
  assign y21201 = n3947 ;
  assign y21202 = n20486 ;
  assign y21203 = ~1'b0 ;
  assign y21204 = ~1'b0 ;
  assign y21205 = ~1'b0 ;
  assign y21206 = ~n28947 ;
  assign y21207 = n13564 ;
  assign y21208 = n28950 ;
  assign y21209 = ~1'b0 ;
  assign y21210 = n28951 ;
  assign y21211 = ~1'b0 ;
  assign y21212 = ~n28952 ;
  assign y21213 = n28955 ;
  assign y21214 = n28958 ;
  assign y21215 = n28959 ;
  assign y21216 = n28960 ;
  assign y21217 = ~1'b0 ;
  assign y21218 = ~1'b0 ;
  assign y21219 = ~n28961 ;
  assign y21220 = ~n28962 ;
  assign y21221 = ~1'b0 ;
  assign y21222 = ~n28967 ;
  assign y21223 = ~n28969 ;
  assign y21224 = ~1'b0 ;
  assign y21225 = n28971 ;
  assign y21226 = n28974 ;
  assign y21227 = ~n28976 ;
  assign y21228 = ~n28978 ;
  assign y21229 = n28981 ;
  assign y21230 = ~1'b0 ;
  assign y21231 = n28984 ;
  assign y21232 = 1'b0 ;
  assign y21233 = ~n18538 ;
  assign y21234 = ~1'b0 ;
  assign y21235 = n28986 ;
  assign y21236 = ~n1810 ;
  assign y21237 = ~n28990 ;
  assign y21238 = 1'b0 ;
  assign y21239 = n28993 ;
  assign y21240 = n28997 ;
  assign y21241 = ~1'b0 ;
  assign y21242 = n28999 ;
  assign y21243 = ~1'b0 ;
  assign y21244 = n29002 ;
  assign y21245 = ~n11844 ;
  assign y21246 = ~n29003 ;
  assign y21247 = ~n646 ;
  assign y21248 = ~n29005 ;
  assign y21249 = ~1'b0 ;
  assign y21250 = ~n11061 ;
  assign y21251 = ~n29009 ;
  assign y21252 = n29010 ;
  assign y21253 = n29011 ;
  assign y21254 = ~1'b0 ;
  assign y21255 = ~n11673 ;
  assign y21256 = n29013 ;
  assign y21257 = ~n29014 ;
  assign y21258 = n29015 ;
  assign y21259 = ~1'b0 ;
  assign y21260 = n2934 ;
  assign y21261 = ~1'b0 ;
  assign y21262 = n29024 ;
  assign y21263 = ~1'b0 ;
  assign y21264 = ~n29026 ;
  assign y21265 = n29031 ;
  assign y21266 = ~n29032 ;
  assign y21267 = ~n29036 ;
  assign y21268 = ~1'b0 ;
  assign y21269 = ~n29037 ;
  assign y21270 = n29041 ;
  assign y21271 = n29043 ;
  assign y21272 = 1'b0 ;
  assign y21273 = ~1'b0 ;
  assign y21274 = ~n29045 ;
  assign y21275 = n29048 ;
  assign y21276 = ~1'b0 ;
  assign y21277 = ~1'b0 ;
  assign y21278 = ~1'b0 ;
  assign y21279 = n29049 ;
  assign y21280 = ~1'b0 ;
  assign y21281 = n29052 ;
  assign y21282 = ~1'b0 ;
  assign y21283 = ~n6142 ;
  assign y21284 = ~n29053 ;
  assign y21285 = ~n29054 ;
  assign y21286 = ~1'b0 ;
  assign y21287 = ~n29055 ;
  assign y21288 = n29063 ;
  assign y21289 = ~n29064 ;
  assign y21290 = n29067 ;
  assign y21291 = ~1'b0 ;
  assign y21292 = ~1'b0 ;
  assign y21293 = 1'b0 ;
  assign y21294 = n29070 ;
  assign y21295 = n21711 ;
  assign y21296 = ~n29075 ;
  assign y21297 = ~n29079 ;
  assign y21298 = ~1'b0 ;
  assign y21299 = ~1'b0 ;
  assign y21300 = 1'b0 ;
  assign y21301 = ~n18433 ;
  assign y21302 = n29081 ;
  assign y21303 = ~1'b0 ;
  assign y21304 = ~1'b0 ;
  assign y21305 = ~n29083 ;
  assign y21306 = n29084 ;
  assign y21307 = ~n29085 ;
  assign y21308 = ~n29086 ;
  assign y21309 = ~n29087 ;
  assign y21310 = ~1'b0 ;
  assign y21311 = ~1'b0 ;
  assign y21312 = 1'b0 ;
  assign y21313 = ~n29089 ;
  assign y21314 = ~1'b0 ;
  assign y21315 = ~n29094 ;
  assign y21316 = n29095 ;
  assign y21317 = n29099 ;
  assign y21318 = ~1'b0 ;
  assign y21319 = n29100 ;
  assign y21320 = ~1'b0 ;
  assign y21321 = ~1'b0 ;
  assign y21322 = ~n29101 ;
  assign y21323 = ~1'b0 ;
  assign y21324 = ~1'b0 ;
  assign y21325 = ~n24512 ;
  assign y21326 = n29102 ;
  assign y21327 = 1'b0 ;
  assign y21328 = n29105 ;
  assign y21329 = ~n29109 ;
  assign y21330 = n29110 ;
  assign y21331 = ~n29113 ;
  assign y21332 = n29115 ;
  assign y21333 = n29116 ;
  assign y21334 = n29119 ;
  assign y21335 = ~1'b0 ;
  assign y21336 = ~1'b0 ;
  assign y21337 = n29120 ;
  assign y21338 = ~n29122 ;
  assign y21339 = 1'b0 ;
  assign y21340 = ~1'b0 ;
  assign y21341 = 1'b0 ;
  assign y21342 = ~1'b0 ;
  assign y21343 = n18595 ;
  assign y21344 = ~1'b0 ;
  assign y21345 = ~1'b0 ;
  assign y21346 = n29123 ;
  assign y21347 = n18455 ;
  assign y21348 = ~1'b0 ;
  assign y21349 = ~n29124 ;
  assign y21350 = n2124 ;
  assign y21351 = ~1'b0 ;
  assign y21352 = n29126 ;
  assign y21353 = ~1'b0 ;
  assign y21354 = n29130 ;
  assign y21355 = ~n3304 ;
  assign y21356 = n29133 ;
  assign y21357 = ~1'b0 ;
  assign y21358 = ~n29136 ;
  assign y21359 = ~1'b0 ;
  assign y21360 = n29139 ;
  assign y21361 = ~n29140 ;
  assign y21362 = ~1'b0 ;
  assign y21363 = ~n29142 ;
  assign y21364 = ~n29143 ;
  assign y21365 = ~n18355 ;
  assign y21366 = 1'b0 ;
  assign y21367 = ~1'b0 ;
  assign y21368 = ~n29146 ;
  assign y21369 = n29149 ;
  assign y21370 = n29150 ;
  assign y21371 = ~n29151 ;
  assign y21372 = ~n29152 ;
  assign y21373 = n715 ;
  assign y21374 = ~n29154 ;
  assign y21375 = ~n29157 ;
  assign y21376 = ~1'b0 ;
  assign y21377 = n29158 ;
  assign y21378 = ~n29164 ;
  assign y21379 = ~n29165 ;
  assign y21380 = n29169 ;
  assign y21381 = n29171 ;
  assign y21382 = n29173 ;
  assign y21383 = n813 ;
  assign y21384 = ~1'b0 ;
  assign y21385 = ~n29175 ;
  assign y21386 = ~n29176 ;
  assign y21387 = ~n29179 ;
  assign y21388 = n29182 ;
  assign y21389 = ~1'b0 ;
  assign y21390 = ~1'b0 ;
  assign y21391 = 1'b0 ;
  assign y21392 = ~1'b0 ;
  assign y21393 = ~n29187 ;
  assign y21394 = n29192 ;
  assign y21395 = ~n29198 ;
  assign y21396 = n29199 ;
  assign y21397 = n29203 ;
  assign y21398 = n29204 ;
  assign y21399 = ~1'b0 ;
  assign y21400 = n29208 ;
  assign y21401 = 1'b0 ;
  assign y21402 = 1'b0 ;
  assign y21403 = ~n10877 ;
  assign y21404 = n29209 ;
  assign y21405 = n29210 ;
  assign y21406 = ~1'b0 ;
  assign y21407 = n29212 ;
  assign y21408 = ~n29219 ;
  assign y21409 = ~1'b0 ;
  assign y21410 = n29221 ;
  assign y21411 = ~1'b0 ;
  assign y21412 = ~1'b0 ;
  assign y21413 = ~1'b0 ;
  assign y21414 = ~1'b0 ;
  assign y21415 = n29222 ;
  assign y21416 = ~n29224 ;
  assign y21417 = n29228 ;
  assign y21418 = n29229 ;
  assign y21419 = n29232 ;
  assign y21420 = n29233 ;
  assign y21421 = n29234 ;
  assign y21422 = ~n29236 ;
  assign y21423 = ~n29237 ;
  assign y21424 = ~1'b0 ;
  assign y21425 = ~n29240 ;
  assign y21426 = n29245 ;
  assign y21427 = ~n29246 ;
  assign y21428 = n29249 ;
  assign y21429 = n29250 ;
  assign y21430 = n26522 ;
  assign y21431 = ~n29251 ;
  assign y21432 = ~n29256 ;
  assign y21433 = 1'b0 ;
  assign y21434 = ~1'b0 ;
  assign y21435 = ~n29257 ;
  assign y21436 = n29259 ;
  assign y21437 = n29261 ;
  assign y21438 = ~n29264 ;
  assign y21439 = ~1'b0 ;
  assign y21440 = 1'b0 ;
  assign y21441 = ~n29265 ;
  assign y21442 = n29267 ;
  assign y21443 = n29268 ;
  assign y21444 = ~n29271 ;
  assign y21445 = n29277 ;
  assign y21446 = ~n29278 ;
  assign y21447 = n29281 ;
  assign y21448 = ~n29284 ;
  assign y21449 = ~n7646 ;
  assign y21450 = ~n29286 ;
  assign y21451 = ~n29287 ;
  assign y21452 = ~1'b0 ;
  assign y21453 = ~n29288 ;
  assign y21454 = ~n29289 ;
  assign y21455 = n29290 ;
  assign y21456 = n29291 ;
  assign y21457 = ~1'b0 ;
  assign y21458 = n5399 ;
  assign y21459 = ~n29299 ;
  assign y21460 = ~n29300 ;
  assign y21461 = ~1'b0 ;
  assign y21462 = ~n16477 ;
  assign y21463 = ~n29303 ;
  assign y21464 = ~1'b0 ;
  assign y21465 = ~1'b0 ;
  assign y21466 = ~n29313 ;
  assign y21467 = ~1'b0 ;
  assign y21468 = ~1'b0 ;
  assign y21469 = ~n29317 ;
  assign y21470 = n29319 ;
  assign y21471 = ~1'b0 ;
  assign y21472 = ~n29321 ;
  assign y21473 = n3710 ;
  assign y21474 = ~1'b0 ;
  assign y21475 = ~n29323 ;
  assign y21476 = ~n29337 ;
  assign y21477 = n27708 ;
  assign y21478 = ~1'b0 ;
  assign y21479 = n29340 ;
  assign y21480 = ~n29341 ;
  assign y21481 = n29347 ;
  assign y21482 = ~n29348 ;
  assign y21483 = ~n29349 ;
  assign y21484 = n29352 ;
  assign y21485 = 1'b0 ;
  assign y21486 = ~1'b0 ;
  assign y21487 = n29354 ;
  assign y21488 = n29356 ;
  assign y21489 = ~1'b0 ;
  assign y21490 = ~n29362 ;
  assign y21491 = ~1'b0 ;
  assign y21492 = ~n29365 ;
  assign y21493 = n29368 ;
  assign y21494 = ~1'b0 ;
  assign y21495 = n29374 ;
  assign y21496 = n29375 ;
  assign y21497 = n29376 ;
  assign y21498 = n13911 ;
  assign y21499 = ~n29377 ;
  assign y21500 = ~n29380 ;
  assign y21501 = n29381 ;
  assign y21502 = n29384 ;
  assign y21503 = ~n29386 ;
  assign y21504 = n29390 ;
  assign y21505 = n29392 ;
  assign y21506 = n29394 ;
  assign y21507 = ~1'b0 ;
  assign y21508 = ~1'b0 ;
  assign y21509 = ~n16454 ;
  assign y21510 = ~n29416 ;
  assign y21511 = ~1'b0 ;
  assign y21512 = n29420 ;
  assign y21513 = n8800 ;
  assign y21514 = ~1'b0 ;
  assign y21515 = ~1'b0 ;
  assign y21516 = ~n29421 ;
  assign y21517 = ~n29425 ;
  assign y21518 = ~1'b0 ;
  assign y21519 = ~n29426 ;
  assign y21520 = n4167 ;
  assign y21521 = ~1'b0 ;
  assign y21522 = ~1'b0 ;
  assign y21523 = 1'b0 ;
  assign y21524 = ~1'b0 ;
  assign y21525 = ~1'b0 ;
  assign y21526 = ~1'b0 ;
  assign y21527 = n29428 ;
  assign y21528 = ~n29429 ;
  assign y21529 = ~1'b0 ;
  assign y21530 = ~1'b0 ;
  assign y21531 = n29436 ;
  assign y21532 = ~1'b0 ;
  assign y21533 = 1'b0 ;
  assign y21534 = n29437 ;
  assign y21535 = ~1'b0 ;
  assign y21536 = n29438 ;
  assign y21537 = ~n29440 ;
  assign y21538 = ~n29441 ;
  assign y21539 = ~1'b0 ;
  assign y21540 = n12180 ;
  assign y21541 = 1'b0 ;
  assign y21542 = ~n29444 ;
  assign y21543 = ~1'b0 ;
  assign y21544 = n29445 ;
  assign y21545 = ~n10470 ;
  assign y21546 = n29447 ;
  assign y21547 = n29450 ;
  assign y21548 = ~n29451 ;
  assign y21549 = n29452 ;
  assign y21550 = ~1'b0 ;
  assign y21551 = n29453 ;
  assign y21552 = ~1'b0 ;
  assign y21553 = ~1'b0 ;
  assign y21554 = ~1'b0 ;
  assign y21555 = ~1'b0 ;
  assign y21556 = n29454 ;
  assign y21557 = ~1'b0 ;
  assign y21558 = n29456 ;
  assign y21559 = ~1'b0 ;
  assign y21560 = ~n29459 ;
  assign y21561 = ~n11763 ;
  assign y21562 = ~1'b0 ;
  assign y21563 = n29460 ;
  assign y21564 = ~1'b0 ;
  assign y21565 = ~1'b0 ;
  assign y21566 = ~n2927 ;
  assign y21567 = n29463 ;
  assign y21568 = n29469 ;
  assign y21569 = ~1'b0 ;
  assign y21570 = 1'b0 ;
  assign y21571 = ~n29470 ;
  assign y21572 = ~n26761 ;
  assign y21573 = 1'b0 ;
  assign y21574 = n29471 ;
  assign y21575 = ~n29472 ;
  assign y21576 = 1'b0 ;
  assign y21577 = ~n36 ;
  assign y21578 = n29474 ;
  assign y21579 = ~n29478 ;
  assign y21580 = ~1'b0 ;
  assign y21581 = ~1'b0 ;
  assign y21582 = 1'b0 ;
  assign y21583 = n29481 ;
  assign y21584 = ~n29483 ;
  assign y21585 = n29484 ;
  assign y21586 = ~1'b0 ;
  assign y21587 = ~n29488 ;
  assign y21588 = ~n29491 ;
  assign y21589 = ~n29495 ;
  assign y21590 = n29497 ;
  assign y21591 = n17523 ;
  assign y21592 = n3414 ;
  assign y21593 = n22597 ;
  assign y21594 = ~n14725 ;
  assign y21595 = ~1'b0 ;
  assign y21596 = ~1'b0 ;
  assign y21597 = n29501 ;
  assign y21598 = ~1'b0 ;
  assign y21599 = ~1'b0 ;
  assign y21600 = ~1'b0 ;
  assign y21601 = ~n29503 ;
  assign y21602 = n29506 ;
  assign y21603 = 1'b0 ;
  assign y21604 = ~1'b0 ;
  assign y21605 = n29507 ;
  assign y21606 = ~1'b0 ;
  assign y21607 = n29510 ;
  assign y21608 = ~1'b0 ;
  assign y21609 = ~n29512 ;
  assign y21610 = ~1'b0 ;
  assign y21611 = n29513 ;
  assign y21612 = ~1'b0 ;
  assign y21613 = ~n29514 ;
  assign y21614 = n29517 ;
  assign y21615 = ~1'b0 ;
  assign y21616 = n29518 ;
  assign y21617 = ~1'b0 ;
  assign y21618 = ~n29520 ;
  assign y21619 = ~1'b0 ;
  assign y21620 = n29522 ;
  assign y21621 = ~1'b0 ;
  assign y21622 = ~n29524 ;
  assign y21623 = ~1'b0 ;
  assign y21624 = ~1'b0 ;
  assign y21625 = ~n29525 ;
  assign y21626 = 1'b0 ;
  assign y21627 = ~1'b0 ;
  assign y21628 = ~n29526 ;
  assign y21629 = ~1'b0 ;
  assign y21630 = n12542 ;
  assign y21631 = 1'b0 ;
  assign y21632 = ~n29528 ;
  assign y21633 = ~1'b0 ;
  assign y21634 = n29530 ;
  assign y21635 = ~1'b0 ;
  assign y21636 = ~1'b0 ;
  assign y21637 = 1'b0 ;
  assign y21638 = ~1'b0 ;
  assign y21639 = n29532 ;
  assign y21640 = ~n29533 ;
  assign y21641 = ~n29535 ;
  assign y21642 = ~n29536 ;
  assign y21643 = n29537 ;
  assign y21644 = ~n29539 ;
  assign y21645 = 1'b0 ;
  assign y21646 = n29543 ;
  assign y21647 = ~n29544 ;
  assign y21648 = ~1'b0 ;
  assign y21649 = n29545 ;
  assign y21650 = 1'b0 ;
  assign y21651 = ~1'b0 ;
  assign y21652 = n1000 ;
  assign y21653 = ~1'b0 ;
  assign y21654 = n29546 ;
  assign y21655 = ~1'b0 ;
  assign y21656 = n1879 ;
  assign y21657 = ~1'b0 ;
  assign y21658 = ~1'b0 ;
  assign y21659 = ~1'b0 ;
  assign y21660 = ~1'b0 ;
  assign y21661 = ~1'b0 ;
  assign y21662 = ~1'b0 ;
  assign y21663 = n29552 ;
  assign y21664 = ~n7231 ;
  assign y21665 = ~n29554 ;
  assign y21666 = ~1'b0 ;
  assign y21667 = n29558 ;
  assign y21668 = ~1'b0 ;
  assign y21669 = ~1'b0 ;
  assign y21670 = n29560 ;
  assign y21671 = ~n29567 ;
  assign y21672 = ~n29572 ;
  assign y21673 = ~n29575 ;
  assign y21674 = ~n29576 ;
  assign y21675 = n29578 ;
  assign y21676 = ~1'b0 ;
  assign y21677 = ~1'b0 ;
  assign y21678 = ~1'b0 ;
  assign y21679 = ~n29579 ;
  assign y21680 = ~n9321 ;
  assign y21681 = ~1'b0 ;
  assign y21682 = ~1'b0 ;
  assign y21683 = ~1'b0 ;
  assign y21684 = n29589 ;
  assign y21685 = ~n29590 ;
  assign y21686 = ~1'b0 ;
  assign y21687 = ~1'b0 ;
  assign y21688 = ~n29591 ;
  assign y21689 = 1'b0 ;
  assign y21690 = ~1'b0 ;
  assign y21691 = n29593 ;
  assign y21692 = ~n29595 ;
  assign y21693 = n29597 ;
  assign y21694 = n29599 ;
  assign y21695 = ~1'b0 ;
  assign y21696 = ~1'b0 ;
  assign y21697 = ~n29600 ;
  assign y21698 = ~n2578 ;
  assign y21699 = ~1'b0 ;
  assign y21700 = ~n29200 ;
  assign y21701 = n29602 ;
  assign y21702 = ~1'b0 ;
  assign y21703 = n29603 ;
  assign y21704 = ~1'b0 ;
  assign y21705 = n29607 ;
  assign y21706 = ~n4303 ;
  assign y21707 = ~1'b0 ;
  assign y21708 = ~1'b0 ;
  assign y21709 = ~n29608 ;
  assign y21710 = ~n29609 ;
  assign y21711 = 1'b0 ;
  assign y21712 = ~n1926 ;
  assign y21713 = ~n29611 ;
  assign y21714 = ~1'b0 ;
  assign y21715 = ~1'b0 ;
  assign y21716 = ~n29612 ;
  assign y21717 = n29613 ;
  assign y21718 = n29617 ;
  assign y21719 = 1'b0 ;
  assign y21720 = n29620 ;
  assign y21721 = ~1'b0 ;
  assign y21722 = n29621 ;
  assign y21723 = ~n29622 ;
  assign y21724 = ~1'b0 ;
  assign y21725 = ~1'b0 ;
  assign y21726 = ~n29624 ;
  assign y21727 = ~n29626 ;
  assign y21728 = n29629 ;
  assign y21729 = n29631 ;
  assign y21730 = ~1'b0 ;
  assign y21731 = ~n29632 ;
  assign y21732 = ~n1250 ;
  assign y21733 = ~n29633 ;
  assign y21734 = ~1'b0 ;
  assign y21735 = ~1'b0 ;
  assign y21736 = n29635 ;
  assign y21737 = n29642 ;
  assign y21738 = n29643 ;
  assign y21739 = ~1'b0 ;
  assign y21740 = ~1'b0 ;
  assign y21741 = ~n29645 ;
  assign y21742 = ~1'b0 ;
  assign y21743 = ~n29649 ;
  assign y21744 = ~n29650 ;
  assign y21745 = ~n29655 ;
  assign y21746 = ~n29657 ;
  assign y21747 = ~n29662 ;
  assign y21748 = n29663 ;
  assign y21749 = ~n29664 ;
  assign y21750 = ~1'b0 ;
  assign y21751 = n29665 ;
  assign y21752 = n29667 ;
  assign y21753 = n10973 ;
  assign y21754 = ~n29668 ;
  assign y21755 = n29670 ;
  assign y21756 = n29671 ;
  assign y21757 = n29672 ;
  assign y21758 = ~n29673 ;
  assign y21759 = ~1'b0 ;
  assign y21760 = n29674 ;
  assign y21761 = ~1'b0 ;
  assign y21762 = n17010 ;
  assign y21763 = ~1'b0 ;
  assign y21764 = ~n9116 ;
  assign y21765 = n29678 ;
  assign y21766 = ~n29679 ;
  assign y21767 = ~n29681 ;
  assign y21768 = ~1'b0 ;
  assign y21769 = n8466 ;
  assign y21770 = n29688 ;
  assign y21771 = n29689 ;
  assign y21772 = ~1'b0 ;
  assign y21773 = n29690 ;
  assign y21774 = n29692 ;
  assign y21775 = n29693 ;
  assign y21776 = n29698 ;
  assign y21777 = ~1'b0 ;
  assign y21778 = ~1'b0 ;
  assign y21779 = n29699 ;
  assign y21780 = n29700 ;
  assign y21781 = ~n29702 ;
  assign y21782 = n29705 ;
  assign y21783 = ~n29707 ;
  assign y21784 = ~1'b0 ;
  assign y21785 = n29710 ;
  assign y21786 = ~n29712 ;
  assign y21787 = n19484 ;
  assign y21788 = ~n29714 ;
  assign y21789 = n29715 ;
  assign y21790 = ~1'b0 ;
  assign y21791 = n29721 ;
  assign y21792 = 1'b0 ;
  assign y21793 = 1'b0 ;
  assign y21794 = ~1'b0 ;
  assign y21795 = ~n538 ;
  assign y21796 = ~1'b0 ;
  assign y21797 = n29723 ;
  assign y21798 = n29724 ;
  assign y21799 = ~n29731 ;
  assign y21800 = 1'b0 ;
  assign y21801 = n14262 ;
  assign y21802 = n29739 ;
  assign y21803 = n29741 ;
  assign y21804 = n29744 ;
  assign y21805 = ~n29747 ;
  assign y21806 = ~1'b0 ;
  assign y21807 = ~n29748 ;
  assign y21808 = ~n29751 ;
  assign y21809 = ~1'b0 ;
  assign y21810 = ~n29753 ;
  assign y21811 = ~n29756 ;
  assign y21812 = ~1'b0 ;
  assign y21813 = n29759 ;
  assign y21814 = ~1'b0 ;
  assign y21815 = ~1'b0 ;
  assign y21816 = n29760 ;
  assign y21817 = ~1'b0 ;
  assign y21818 = ~n29763 ;
  assign y21819 = n29764 ;
  assign y21820 = ~n29768 ;
  assign y21821 = ~n29772 ;
  assign y21822 = ~n29776 ;
  assign y21823 = ~1'b0 ;
  assign y21824 = ~1'b0 ;
  assign y21825 = ~n29777 ;
  assign y21826 = ~n29778 ;
  assign y21827 = ~1'b0 ;
  assign y21828 = n29782 ;
  assign y21829 = ~1'b0 ;
  assign y21830 = n29783 ;
  assign y21831 = n29786 ;
  assign y21832 = n7908 ;
  assign y21833 = ~n29788 ;
  assign y21834 = ~1'b0 ;
  assign y21835 = n24553 ;
  assign y21836 = n29790 ;
  assign y21837 = n29791 ;
  assign y21838 = ~n29795 ;
  assign y21839 = ~1'b0 ;
  assign y21840 = ~1'b0 ;
  assign y21841 = ~n29796 ;
  assign y21842 = ~n29802 ;
  assign y21843 = ~n29804 ;
  assign y21844 = n29805 ;
  assign y21845 = ~1'b0 ;
  assign y21846 = n29806 ;
  assign y21847 = 1'b0 ;
  assign y21848 = ~n29808 ;
  assign y21849 = ~1'b0 ;
  assign y21850 = ~1'b0 ;
  assign y21851 = n29810 ;
  assign y21852 = ~n6462 ;
  assign y21853 = ~1'b0 ;
  assign y21854 = ~1'b0 ;
  assign y21855 = n29818 ;
  assign y21856 = ~n29819 ;
  assign y21857 = ~n29820 ;
  assign y21858 = ~n29821 ;
  assign y21859 = ~1'b0 ;
  assign y21860 = ~n1151 ;
  assign y21861 = ~n29827 ;
  assign y21862 = ~n29828 ;
  assign y21863 = ~n29829 ;
  assign y21864 = n12702 ;
  assign y21865 = n29830 ;
  assign y21866 = ~n29831 ;
  assign y21867 = ~n29832 ;
  assign y21868 = n29833 ;
  assign y21869 = ~n29838 ;
  assign y21870 = ~1'b0 ;
  assign y21871 = ~n7090 ;
  assign y21872 = n29840 ;
  assign y21873 = n29841 ;
  assign y21874 = 1'b0 ;
  assign y21875 = ~n22540 ;
  assign y21876 = n29844 ;
  assign y21877 = ~1'b0 ;
  assign y21878 = ~n29845 ;
  assign y21879 = ~1'b0 ;
  assign y21880 = ~1'b0 ;
  assign y21881 = n28810 ;
  assign y21882 = ~1'b0 ;
  assign y21883 = ~1'b0 ;
  assign y21884 = ~1'b0 ;
  assign y21885 = ~1'b0 ;
  assign y21886 = ~n29846 ;
  assign y21887 = ~n29847 ;
  assign y21888 = ~1'b0 ;
  assign y21889 = ~1'b0 ;
  assign y21890 = ~n29848 ;
  assign y21891 = ~1'b0 ;
  assign y21892 = n29850 ;
  assign y21893 = ~n29853 ;
  assign y21894 = 1'b0 ;
  assign y21895 = n29858 ;
  assign y21896 = n11465 ;
  assign y21897 = ~1'b0 ;
  assign y21898 = n29868 ;
  assign y21899 = n29873 ;
  assign y21900 = ~n29875 ;
  assign y21901 = n29345 ;
  assign y21902 = n29877 ;
  assign y21903 = ~n29880 ;
  assign y21904 = ~1'b0 ;
  assign y21905 = ~n29883 ;
  assign y21906 = ~n29885 ;
  assign y21907 = ~1'b0 ;
  assign y21908 = n29887 ;
  assign y21909 = ~1'b0 ;
  assign y21910 = ~1'b0 ;
  assign y21911 = n29888 ;
  assign y21912 = 1'b0 ;
  assign y21913 = ~1'b0 ;
  assign y21914 = ~n29898 ;
  assign y21915 = ~1'b0 ;
  assign y21916 = n13715 ;
  assign y21917 = ~1'b0 ;
  assign y21918 = ~n29901 ;
  assign y21919 = n29902 ;
  assign y21920 = ~1'b0 ;
  assign y21921 = n10734 ;
  assign y21922 = ~1'b0 ;
  assign y21923 = ~n29903 ;
  assign y21924 = ~n29907 ;
  assign y21925 = ~1'b0 ;
  assign y21926 = ~n29909 ;
  assign y21927 = ~1'b0 ;
  assign y21928 = n29911 ;
  assign y21929 = ~n29913 ;
  assign y21930 = ~n29914 ;
  assign y21931 = ~1'b0 ;
  assign y21932 = n29916 ;
  assign y21933 = n29918 ;
  assign y21934 = ~1'b0 ;
  assign y21935 = n29919 ;
  assign y21936 = ~1'b0 ;
  assign y21937 = n29921 ;
  assign y21938 = ~1'b0 ;
  assign y21939 = n3799 ;
  assign y21940 = ~1'b0 ;
  assign y21941 = n29923 ;
  assign y21942 = ~n29925 ;
  assign y21943 = ~n29927 ;
  assign y21944 = ~n29928 ;
  assign y21945 = n29929 ;
  assign y21946 = n29930 ;
  assign y21947 = ~1'b0 ;
  assign y21948 = ~n29932 ;
  assign y21949 = ~1'b0 ;
  assign y21950 = ~1'b0 ;
  assign y21951 = ~n29933 ;
  assign y21952 = ~1'b0 ;
  assign y21953 = n29935 ;
  assign y21954 = n24652 ;
  assign y21955 = n29937 ;
  assign y21956 = n29939 ;
  assign y21957 = ~1'b0 ;
  assign y21958 = ~n29942 ;
  assign y21959 = ~1'b0 ;
  assign y21960 = n10816 ;
  assign y21961 = n15552 ;
  assign y21962 = n1565 ;
  assign y21963 = ~1'b0 ;
  assign y21964 = ~1'b0 ;
  assign y21965 = ~n29948 ;
  assign y21966 = ~n29949 ;
  assign y21967 = ~n12303 ;
  assign y21968 = n29951 ;
  assign y21969 = ~n29955 ;
  assign y21970 = ~n29956 ;
  assign y21971 = ~1'b0 ;
  assign y21972 = 1'b0 ;
  assign y21973 = ~1'b0 ;
  assign y21974 = ~n29957 ;
  assign y21975 = ~n29959 ;
  assign y21976 = ~n29961 ;
  assign y21977 = n29965 ;
  assign y21978 = ~n29967 ;
  assign y21979 = ~n29971 ;
  assign y21980 = ~1'b0 ;
  assign y21981 = n10778 ;
  assign y21982 = n29975 ;
  assign y21983 = n29976 ;
  assign y21984 = 1'b0 ;
  assign y21985 = n29977 ;
  assign y21986 = ~1'b0 ;
  assign y21987 = ~n2539 ;
  assign y21988 = ~n29979 ;
  assign y21989 = ~1'b0 ;
  assign y21990 = ~1'b0 ;
  assign y21991 = n29980 ;
  assign y21992 = ~1'b0 ;
  assign y21993 = ~n29981 ;
  assign y21994 = ~1'b0 ;
  assign y21995 = n13962 ;
  assign y21996 = ~1'b0 ;
  assign y21997 = 1'b0 ;
  assign y21998 = ~1'b0 ;
  assign y21999 = ~1'b0 ;
  assign y22000 = ~n29982 ;
  assign y22001 = ~1'b0 ;
  assign y22002 = n29983 ;
  assign y22003 = ~1'b0 ;
  assign y22004 = ~1'b0 ;
  assign y22005 = n29986 ;
  assign y22006 = ~1'b0 ;
  assign y22007 = ~n29989 ;
  assign y22008 = ~1'b0 ;
  assign y22009 = ~1'b0 ;
  assign y22010 = ~n29991 ;
  assign y22011 = n29995 ;
  assign y22012 = ~1'b0 ;
  assign y22013 = ~1'b0 ;
  assign y22014 = n29997 ;
  assign y22015 = ~1'b0 ;
  assign y22016 = n29999 ;
  assign y22017 = n30000 ;
  assign y22018 = ~1'b0 ;
  assign y22019 = ~1'b0 ;
  assign y22020 = n30001 ;
  assign y22021 = n30004 ;
  assign y22022 = ~n30007 ;
  assign y22023 = n30009 ;
  assign y22024 = n30013 ;
  assign y22025 = ~1'b0 ;
  assign y22026 = ~1'b0 ;
  assign y22027 = ~1'b0 ;
  assign y22028 = n30014 ;
  assign y22029 = 1'b0 ;
  assign y22030 = ~1'b0 ;
  assign y22031 = ~1'b0 ;
  assign y22032 = ~1'b0 ;
  assign y22033 = n30018 ;
  assign y22034 = ~n30020 ;
  assign y22035 = ~1'b0 ;
  assign y22036 = ~n30022 ;
  assign y22037 = n9536 ;
  assign y22038 = n4092 ;
  assign y22039 = n30023 ;
  assign y22040 = n30027 ;
  assign y22041 = ~n25453 ;
  assign y22042 = ~n30041 ;
  assign y22043 = ~n30042 ;
  assign y22044 = n30043 ;
  assign y22045 = ~n30045 ;
  assign y22046 = ~n30049 ;
  assign y22047 = ~n22676 ;
  assign y22048 = n30051 ;
  assign y22049 = ~1'b0 ;
  assign y22050 = ~1'b0 ;
  assign y22051 = 1'b0 ;
  assign y22052 = n30052 ;
  assign y22053 = n30054 ;
  assign y22054 = n30055 ;
  assign y22055 = ~1'b0 ;
  assign y22056 = ~n12280 ;
  assign y22057 = n30057 ;
  assign y22058 = ~1'b0 ;
  assign y22059 = ~1'b0 ;
  assign y22060 = ~1'b0 ;
  assign y22061 = ~1'b0 ;
  assign y22062 = n30063 ;
  assign y22063 = n30065 ;
  assign y22064 = n30066 ;
  assign y22065 = ~1'b0 ;
  assign y22066 = ~1'b0 ;
  assign y22067 = ~1'b0 ;
  assign y22068 = ~1'b0 ;
  assign y22069 = n30067 ;
  assign y22070 = n30071 ;
  assign y22071 = ~1'b0 ;
  assign y22072 = ~n30073 ;
  assign y22073 = 1'b0 ;
  assign y22074 = ~1'b0 ;
  assign y22075 = n30074 ;
  assign y22076 = ~n30075 ;
  assign y22077 = ~1'b0 ;
  assign y22078 = ~1'b0 ;
  assign y22079 = n30076 ;
  assign y22080 = ~n30086 ;
  assign y22081 = 1'b0 ;
  assign y22082 = ~n30089 ;
  assign y22083 = ~n30090 ;
  assign y22084 = ~1'b0 ;
  assign y22085 = n30092 ;
  assign y22086 = ~n30095 ;
  assign y22087 = n30099 ;
  assign y22088 = ~1'b0 ;
  assign y22089 = n30102 ;
  assign y22090 = ~n30107 ;
  assign y22091 = ~n30108 ;
  assign y22092 = n11604 ;
  assign y22093 = ~1'b0 ;
  assign y22094 = n30110 ;
  assign y22095 = ~n30113 ;
  assign y22096 = ~n30117 ;
  assign y22097 = n30118 ;
  assign y22098 = ~n30119 ;
  assign y22099 = ~1'b0 ;
  assign y22100 = ~n29777 ;
  assign y22101 = ~1'b0 ;
  assign y22102 = ~n30121 ;
  assign y22103 = n30125 ;
  assign y22104 = ~n30127 ;
  assign y22105 = ~n30129 ;
  assign y22106 = n30130 ;
  assign y22107 = ~1'b0 ;
  assign y22108 = ~1'b0 ;
  assign y22109 = ~n15864 ;
  assign y22110 = ~n12002 ;
  assign y22111 = ~n30131 ;
  assign y22112 = ~n30134 ;
  assign y22113 = ~1'b0 ;
  assign y22114 = n30135 ;
  assign y22115 = n30139 ;
  assign y22116 = n159 ;
  assign y22117 = n30140 ;
  assign y22118 = ~n30142 ;
  assign y22119 = ~1'b0 ;
  assign y22120 = ~1'b0 ;
  assign y22121 = 1'b0 ;
  assign y22122 = ~1'b0 ;
  assign y22123 = ~n30144 ;
  assign y22124 = ~n30150 ;
  assign y22125 = n27240 ;
  assign y22126 = n30152 ;
  assign y22127 = ~1'b0 ;
  assign y22128 = ~n30154 ;
  assign y22129 = ~n30158 ;
  assign y22130 = ~n23975 ;
  assign y22131 = ~n30159 ;
  assign y22132 = ~n30162 ;
  assign y22133 = ~1'b0 ;
  assign y22134 = 1'b0 ;
  assign y22135 = ~1'b0 ;
  assign y22136 = n30165 ;
  assign y22137 = ~n1834 ;
  assign y22138 = n30189 ;
  assign y22139 = 1'b0 ;
  assign y22140 = ~1'b0 ;
  assign y22141 = n566 ;
  assign y22142 = n30190 ;
  assign y22143 = ~1'b0 ;
  assign y22144 = n30192 ;
  assign y22145 = ~n30194 ;
  assign y22146 = ~1'b0 ;
  assign y22147 = n30197 ;
  assign y22148 = ~1'b0 ;
  assign y22149 = ~n30198 ;
  assign y22150 = ~1'b0 ;
  assign y22151 = 1'b0 ;
  assign y22152 = ~n30199 ;
  assign y22153 = ~n30202 ;
  assign y22154 = n30204 ;
  assign y22155 = ~1'b0 ;
  assign y22156 = ~1'b0 ;
  assign y22157 = ~1'b0 ;
  assign y22158 = n30205 ;
  assign y22159 = n30208 ;
  assign y22160 = ~n30209 ;
  assign y22161 = ~1'b0 ;
  assign y22162 = ~1'b0 ;
  assign y22163 = n30212 ;
  assign y22164 = n30214 ;
  assign y22165 = ~1'b0 ;
  assign y22166 = ~1'b0 ;
  assign y22167 = n30218 ;
  assign y22168 = n30219 ;
  assign y22169 = ~1'b0 ;
  assign y22170 = n30220 ;
  assign y22171 = ~1'b0 ;
  assign y22172 = n30222 ;
  assign y22173 = n30226 ;
  assign y22174 = ~1'b0 ;
  assign y22175 = n30227 ;
  assign y22176 = n30229 ;
  assign y22177 = n30231 ;
  assign y22178 = n30232 ;
  assign y22179 = ~1'b0 ;
  assign y22180 = n30233 ;
  assign y22181 = n30237 ;
  assign y22182 = ~1'b0 ;
  assign y22183 = n30239 ;
  assign y22184 = ~n395 ;
  assign y22185 = ~1'b0 ;
  assign y22186 = ~1'b0 ;
  assign y22187 = ~n30243 ;
  assign y22188 = ~n19591 ;
  assign y22189 = ~1'b0 ;
  assign y22190 = n30246 ;
  assign y22191 = ~n27199 ;
  assign y22192 = ~1'b0 ;
  assign y22193 = ~n30250 ;
  assign y22194 = ~n3196 ;
  assign y22195 = 1'b0 ;
  assign y22196 = ~n30256 ;
  assign y22197 = ~n30257 ;
  assign y22198 = ~1'b0 ;
  assign y22199 = ~1'b0 ;
  assign y22200 = n30258 ;
  assign y22201 = ~1'b0 ;
  assign y22202 = ~1'b0 ;
  assign y22203 = ~1'b0 ;
  assign y22204 = ~1'b0 ;
  assign y22205 = n10061 ;
  assign y22206 = ~1'b0 ;
  assign y22207 = ~1'b0 ;
  assign y22208 = ~n30259 ;
  assign y22209 = n12697 ;
  assign y22210 = ~n2198 ;
  assign y22211 = ~1'b0 ;
  assign y22212 = ~1'b0 ;
  assign y22213 = ~1'b0 ;
  assign y22214 = n30260 ;
  assign y22215 = ~1'b0 ;
  assign y22216 = ~n30261 ;
  assign y22217 = 1'b0 ;
  assign y22218 = ~n4805 ;
  assign y22219 = ~n30262 ;
  assign y22220 = n27548 ;
  assign y22221 = ~1'b0 ;
  assign y22222 = n30264 ;
  assign y22223 = ~1'b0 ;
  assign y22224 = ~n13555 ;
  assign y22225 = ~n5049 ;
  assign y22226 = ~1'b0 ;
  assign y22227 = ~1'b0 ;
  assign y22228 = ~n17891 ;
  assign y22229 = ~1'b0 ;
  assign y22230 = n3221 ;
  assign y22231 = ~n30267 ;
  assign y22232 = ~n30269 ;
  assign y22233 = ~1'b0 ;
  assign y22234 = ~1'b0 ;
  assign y22235 = ~n30270 ;
  assign y22236 = ~n30275 ;
  assign y22237 = ~n30276 ;
  assign y22238 = ~1'b0 ;
  assign y22239 = ~1'b0 ;
  assign y22240 = ~n30278 ;
  assign y22241 = 1'b0 ;
  assign y22242 = n30283 ;
  assign y22243 = ~1'b0 ;
  assign y22244 = ~1'b0 ;
  assign y22245 = 1'b0 ;
  assign y22246 = ~n30284 ;
  assign y22247 = n30287 ;
  assign y22248 = ~n30291 ;
  assign y22249 = n30292 ;
  assign y22250 = ~n30293 ;
  assign y22251 = ~n30296 ;
  assign y22252 = n2911 ;
  assign y22253 = ~1'b0 ;
  assign y22254 = ~n30300 ;
  assign y22255 = ~1'b0 ;
  assign y22256 = ~1'b0 ;
  assign y22257 = ~n30301 ;
  assign y22258 = ~1'b0 ;
  assign y22259 = ~1'b0 ;
  assign y22260 = ~1'b0 ;
  assign y22261 = ~1'b0 ;
  assign y22262 = n30303 ;
  assign y22263 = ~1'b0 ;
  assign y22264 = ~n30304 ;
  assign y22265 = ~1'b0 ;
  assign y22266 = ~n30309 ;
  assign y22267 = ~1'b0 ;
  assign y22268 = ~1'b0 ;
  assign y22269 = n30311 ;
  assign y22270 = ~1'b0 ;
  assign y22271 = ~n30316 ;
  assign y22272 = ~1'b0 ;
  assign y22273 = ~n30320 ;
  assign y22274 = ~n30321 ;
  assign y22275 = n30322 ;
  assign y22276 = ~n30330 ;
  assign y22277 = ~1'b0 ;
  assign y22278 = ~n30333 ;
  assign y22279 = ~n9359 ;
  assign y22280 = n30334 ;
  assign y22281 = n30335 ;
  assign y22282 = ~1'b0 ;
  assign y22283 = ~n7439 ;
  assign y22284 = n30409 ;
  assign y22285 = ~n30411 ;
  assign y22286 = n30412 ;
  assign y22287 = ~1'b0 ;
  assign y22288 = ~1'b0 ;
  assign y22289 = ~n30414 ;
  assign y22290 = ~n30416 ;
  assign y22291 = 1'b0 ;
  assign y22292 = n3682 ;
  assign y22293 = ~1'b0 ;
  assign y22294 = n30419 ;
  assign y22295 = ~n30423 ;
  assign y22296 = n30424 ;
  assign y22297 = ~1'b0 ;
  assign y22298 = ~n30430 ;
  assign y22299 = ~1'b0 ;
  assign y22300 = ~1'b0 ;
  assign y22301 = 1'b0 ;
  assign y22302 = n30431 ;
  assign y22303 = n30432 ;
  assign y22304 = ~n30435 ;
  assign y22305 = n30436 ;
  assign y22306 = ~n27531 ;
  assign y22307 = ~1'b0 ;
  assign y22308 = n7395 ;
  assign y22309 = ~n5277 ;
  assign y22310 = n980 ;
  assign y22311 = ~1'b0 ;
  assign y22312 = ~1'b0 ;
  assign y22313 = n12973 ;
  assign y22314 = ~1'b0 ;
  assign y22315 = ~n30438 ;
  assign y22316 = ~1'b0 ;
  assign y22317 = ~1'b0 ;
  assign y22318 = ~1'b0 ;
  assign y22319 = ~1'b0 ;
  assign y22320 = ~1'b0 ;
  assign y22321 = ~1'b0 ;
  assign y22322 = ~n30446 ;
  assign y22323 = ~n30448 ;
  assign y22324 = n15030 ;
  assign y22325 = ~n30449 ;
  assign y22326 = ~1'b0 ;
  assign y22327 = ~n30450 ;
  assign y22328 = n30455 ;
  assign y22329 = ~n30460 ;
  assign y22330 = ~1'b0 ;
  assign y22331 = ~n30464 ;
  assign y22332 = ~n30466 ;
  assign y22333 = ~1'b0 ;
  assign y22334 = n6622 ;
  assign y22335 = n7754 ;
  assign y22336 = n30468 ;
  assign y22337 = ~1'b0 ;
  assign y22338 = ~n30469 ;
  assign y22339 = 1'b0 ;
  assign y22340 = ~1'b0 ;
  assign y22341 = ~n8275 ;
  assign y22342 = ~n30471 ;
  assign y22343 = ~1'b0 ;
  assign y22344 = ~n30472 ;
  assign y22345 = ~n500 ;
  assign y22346 = n30473 ;
  assign y22347 = 1'b0 ;
  assign y22348 = n30475 ;
  assign y22349 = n30481 ;
  assign y22350 = n5280 ;
  assign y22351 = n30483 ;
  assign y22352 = 1'b0 ;
  assign y22353 = 1'b0 ;
  assign y22354 = ~n30485 ;
  assign y22355 = ~1'b0 ;
  assign y22356 = n30488 ;
  assign y22357 = ~1'b0 ;
  assign y22358 = ~n30490 ;
  assign y22359 = n30491 ;
  assign y22360 = n30493 ;
  assign y22361 = ~n30496 ;
  assign y22362 = n30498 ;
  assign y22363 = ~1'b0 ;
  assign y22364 = ~n10858 ;
  assign y22365 = ~n30499 ;
  assign y22366 = n25419 ;
  assign y22367 = n30507 ;
  assign y22368 = ~n21764 ;
  assign y22369 = ~1'b0 ;
  assign y22370 = 1'b0 ;
  assign y22371 = ~n30508 ;
  assign y22372 = n30514 ;
  assign y22373 = n30516 ;
  assign y22374 = ~1'b0 ;
  assign y22375 = ~1'b0 ;
  assign y22376 = ~n30517 ;
  assign y22377 = ~n30522 ;
  assign y22378 = n30526 ;
  assign y22379 = ~1'b0 ;
  assign y22380 = ~1'b0 ;
  assign y22381 = ~n30530 ;
  assign y22382 = ~1'b0 ;
  assign y22383 = n30535 ;
  assign y22384 = ~n30536 ;
  assign y22385 = ~1'b0 ;
  assign y22386 = ~n26899 ;
  assign y22387 = n30538 ;
  assign y22388 = ~1'b0 ;
  assign y22389 = ~1'b0 ;
  assign y22390 = ~n30539 ;
  assign y22391 = n30540 ;
  assign y22392 = ~n970 ;
  assign y22393 = ~n30542 ;
  assign y22394 = ~1'b0 ;
  assign y22395 = ~1'b0 ;
  assign y22396 = ~1'b0 ;
  assign y22397 = n30543 ;
  assign y22398 = 1'b0 ;
  assign y22399 = ~1'b0 ;
  assign y22400 = ~1'b0 ;
  assign y22401 = ~1'b0 ;
  assign y22402 = ~1'b0 ;
  assign y22403 = n30544 ;
  assign y22404 = n30545 ;
  assign y22405 = ~n30547 ;
  assign y22406 = n997 ;
  assign y22407 = n27535 ;
  assign y22408 = ~n30554 ;
  assign y22409 = ~1'b0 ;
  assign y22410 = n13961 ;
  assign y22411 = ~1'b0 ;
  assign y22412 = ~1'b0 ;
  assign y22413 = n30557 ;
  assign y22414 = n30559 ;
  assign y22415 = ~n7951 ;
  assign y22416 = ~1'b0 ;
  assign y22417 = ~1'b0 ;
  assign y22418 = n30560 ;
  assign y22419 = ~1'b0 ;
  assign y22420 = n30564 ;
  assign y22421 = ~1'b0 ;
  assign y22422 = ~n30567 ;
  assign y22423 = ~n30568 ;
  assign y22424 = n30590 ;
  assign y22425 = ~n30592 ;
  assign y22426 = ~1'b0 ;
  assign y22427 = ~n30595 ;
  assign y22428 = ~n30596 ;
  assign y22429 = n30598 ;
  assign y22430 = ~n30602 ;
  assign y22431 = ~1'b0 ;
  assign y22432 = ~1'b0 ;
  assign y22433 = n30604 ;
  assign y22434 = n30607 ;
  assign y22435 = n30610 ;
  assign y22436 = ~1'b0 ;
  assign y22437 = n30612 ;
  assign y22438 = ~1'b0 ;
  assign y22439 = ~1'b0 ;
  assign y22440 = n30615 ;
  assign y22441 = ~n30617 ;
  assign y22442 = n30619 ;
  assign y22443 = ~1'b0 ;
  assign y22444 = ~1'b0 ;
  assign y22445 = ~n30620 ;
  assign y22446 = ~n30623 ;
  assign y22447 = n30624 ;
  assign y22448 = n30625 ;
  assign y22449 = n30628 ;
  assign y22450 = ~n30631 ;
  assign y22451 = n30633 ;
  assign y22452 = n227 ;
  assign y22453 = ~n30635 ;
  assign y22454 = ~n30637 ;
  assign y22455 = ~n30641 ;
  assign y22456 = x11 ;
  assign y22457 = ~n30642 ;
  assign y22458 = n30643 ;
  assign y22459 = n30646 ;
  assign y22460 = ~1'b0 ;
  assign y22461 = n30649 ;
  assign y22462 = ~n30650 ;
  assign y22463 = n30652 ;
  assign y22464 = n30653 ;
  assign y22465 = n30656 ;
  assign y22466 = ~n3158 ;
  assign y22467 = ~n27272 ;
  assign y22468 = ~n30659 ;
  assign y22469 = 1'b0 ;
  assign y22470 = n30663 ;
  assign y22471 = n30665 ;
  assign y22472 = ~1'b0 ;
  assign y22473 = ~1'b0 ;
  assign y22474 = n21613 ;
  assign y22475 = n30672 ;
  assign y22476 = ~1'b0 ;
  assign y22477 = ~1'b0 ;
  assign y22478 = n30673 ;
  assign y22479 = ~1'b0 ;
  assign y22480 = ~1'b0 ;
  assign y22481 = 1'b0 ;
  assign y22482 = 1'b0 ;
  assign y22483 = ~1'b0 ;
  assign y22484 = ~n30675 ;
  assign y22485 = n30679 ;
  assign y22486 = ~n30680 ;
  assign y22487 = n9370 ;
  assign y22488 = n30682 ;
  assign y22489 = ~1'b0 ;
  assign y22490 = n25711 ;
  assign y22491 = ~n30684 ;
  assign y22492 = ~n30689 ;
  assign y22493 = ~1'b0 ;
  assign y22494 = ~n30691 ;
  assign y22495 = ~n30694 ;
  assign y22496 = n30698 ;
  assign y22497 = ~1'b0 ;
  assign y22498 = n30699 ;
  assign y22499 = ~n30705 ;
  assign y22500 = n30710 ;
  assign y22501 = n30713 ;
  assign y22502 = ~1'b0 ;
  assign y22503 = ~1'b0 ;
  assign y22504 = n17008 ;
  assign y22505 = ~n30714 ;
  assign y22506 = ~1'b0 ;
  assign y22507 = ~1'b0 ;
  assign y22508 = ~n30715 ;
  assign y22509 = 1'b0 ;
  assign y22510 = ~n30716 ;
  assign y22511 = ~n30717 ;
  assign y22512 = ~1'b0 ;
  assign y22513 = n29144 ;
  assign y22514 = 1'b0 ;
  assign y22515 = ~n30718 ;
  assign y22516 = ~1'b0 ;
  assign y22517 = ~1'b0 ;
  assign y22518 = ~1'b0 ;
  assign y22519 = ~n30720 ;
  assign y22520 = ~1'b0 ;
  assign y22521 = n30722 ;
  assign y22522 = ~n30723 ;
  assign y22523 = ~1'b0 ;
  assign y22524 = n30724 ;
  assign y22525 = ~n30725 ;
  assign y22526 = n30734 ;
  assign y22527 = ~n30736 ;
  assign y22528 = n30738 ;
  assign y22529 = n30739 ;
  assign y22530 = ~1'b0 ;
  assign y22531 = ~n30740 ;
  assign y22532 = ~1'b0 ;
  assign y22533 = ~1'b0 ;
  assign y22534 = n5634 ;
  assign y22535 = n12985 ;
  assign y22536 = ~1'b0 ;
  assign y22537 = ~n30741 ;
  assign y22538 = ~n5347 ;
  assign y22539 = ~n30743 ;
  assign y22540 = ~1'b0 ;
  assign y22541 = ~1'b0 ;
  assign y22542 = ~1'b0 ;
  assign y22543 = ~n30744 ;
  assign y22544 = n30745 ;
  assign y22545 = n30746 ;
  assign y22546 = ~1'b0 ;
  assign y22547 = ~1'b0 ;
  assign y22548 = ~1'b0 ;
  assign y22549 = n30748 ;
  assign y22550 = n30749 ;
  assign y22551 = n1277 ;
  assign y22552 = n21767 ;
  assign y22553 = ~1'b0 ;
  assign y22554 = ~1'b0 ;
  assign y22555 = ~1'b0 ;
  assign y22556 = ~n30752 ;
  assign y22557 = ~1'b0 ;
  assign y22558 = ~1'b0 ;
  assign y22559 = n30755 ;
  assign y22560 = ~1'b0 ;
  assign y22561 = ~1'b0 ;
  assign y22562 = ~n30756 ;
  assign y22563 = ~1'b0 ;
  assign y22564 = n30757 ;
  assign y22565 = n30758 ;
  assign y22566 = n30759 ;
  assign y22567 = ~1'b0 ;
  assign y22568 = n30760 ;
  assign y22569 = ~n30763 ;
  assign y22570 = n30765 ;
  assign y22571 = ~1'b0 ;
  assign y22572 = ~n30767 ;
  assign y22573 = ~n30768 ;
  assign y22574 = n30771 ;
  assign y22575 = ~n30773 ;
  assign y22576 = ~1'b0 ;
  assign y22577 = ~n30775 ;
  assign y22578 = n30776 ;
  assign y22579 = ~1'b0 ;
  assign y22580 = ~1'b0 ;
  assign y22581 = ~1'b0 ;
  assign y22582 = ~1'b0 ;
  assign y22583 = ~1'b0 ;
  assign y22584 = ~n30777 ;
  assign y22585 = ~n30778 ;
  assign y22586 = ~n17923 ;
  assign y22587 = n30781 ;
  assign y22588 = n30782 ;
  assign y22589 = ~1'b0 ;
  assign y22590 = ~1'b0 ;
  assign y22591 = ~1'b0 ;
  assign y22592 = ~n30786 ;
  assign y22593 = ~1'b0 ;
  assign y22594 = ~n30787 ;
  assign y22595 = ~n30788 ;
  assign y22596 = ~n30789 ;
  assign y22597 = n8047 ;
  assign y22598 = n30790 ;
  assign y22599 = ~n30791 ;
  assign y22600 = ~1'b0 ;
  assign y22601 = ~n30792 ;
  assign y22602 = n30793 ;
  assign y22603 = ~1'b0 ;
  assign y22604 = ~1'b0 ;
  assign y22605 = n30799 ;
  assign y22606 = n30800 ;
  assign y22607 = n30801 ;
  assign y22608 = ~1'b0 ;
  assign y22609 = n30802 ;
  assign y22610 = ~1'b0 ;
  assign y22611 = ~n30804 ;
  assign y22612 = ~1'b0 ;
  assign y22613 = n30806 ;
  assign y22614 = ~1'b0 ;
  assign y22615 = 1'b0 ;
  assign y22616 = ~1'b0 ;
  assign y22617 = n30807 ;
  assign y22618 = n906 ;
  assign y22619 = ~n30808 ;
  assign y22620 = ~1'b0 ;
  assign y22621 = ~n30810 ;
  assign y22622 = ~1'b0 ;
  assign y22623 = ~n27748 ;
  assign y22624 = ~n14790 ;
  assign y22625 = n19315 ;
  assign y22626 = n30812 ;
  assign y22627 = ~1'b0 ;
  assign y22628 = ~n2790 ;
  assign y22629 = n30814 ;
  assign y22630 = n6436 ;
  assign y22631 = ~1'b0 ;
  assign y22632 = ~1'b0 ;
  assign y22633 = ~n13606 ;
  assign y22634 = ~n23869 ;
  assign y22635 = ~1'b0 ;
  assign y22636 = ~n30816 ;
  assign y22637 = ~1'b0 ;
  assign y22638 = ~1'b0 ;
  assign y22639 = n30819 ;
  assign y22640 = ~1'b0 ;
  assign y22641 = ~n30820 ;
  assign y22642 = 1'b0 ;
  assign y22643 = ~n203 ;
  assign y22644 = ~1'b0 ;
  assign y22645 = 1'b0 ;
  assign y22646 = ~n30822 ;
  assign y22647 = ~n30823 ;
  assign y22648 = ~n30824 ;
  assign y22649 = n30826 ;
  assign y22650 = n30827 ;
  assign y22651 = n30829 ;
  assign y22652 = n30831 ;
  assign y22653 = n30834 ;
  assign y22654 = ~1'b0 ;
  assign y22655 = ~1'b0 ;
  assign y22656 = ~1'b0 ;
  assign y22657 = n30838 ;
  assign y22658 = ~n30840 ;
  assign y22659 = ~n30841 ;
  assign y22660 = ~1'b0 ;
  assign y22661 = ~n30844 ;
  assign y22662 = n30847 ;
  assign y22663 = n30848 ;
  assign y22664 = ~1'b0 ;
  assign y22665 = ~1'b0 ;
  assign y22666 = ~1'b0 ;
  assign y22667 = ~n28390 ;
  assign y22668 = n30852 ;
  assign y22669 = n30858 ;
  assign y22670 = 1'b0 ;
  assign y22671 = ~1'b0 ;
  assign y22672 = n30859 ;
  assign y22673 = 1'b0 ;
  assign y22674 = ~n30860 ;
  assign y22675 = ~1'b0 ;
  assign y22676 = ~n157 ;
  assign y22677 = 1'b0 ;
  assign y22678 = n6281 ;
  assign y22679 = n30866 ;
  assign y22680 = ~n30867 ;
  assign y22681 = ~n30868 ;
  assign y22682 = ~n30869 ;
  assign y22683 = n30870 ;
  assign y22684 = ~1'b0 ;
  assign y22685 = ~1'b0 ;
  assign y22686 = ~n30871 ;
  assign y22687 = ~1'b0 ;
  assign y22688 = ~1'b0 ;
  assign y22689 = ~n30872 ;
  assign y22690 = ~n30873 ;
  assign y22691 = n30877 ;
  assign y22692 = ~1'b0 ;
  assign y22693 = n30885 ;
  assign y22694 = n30889 ;
  assign y22695 = ~1'b0 ;
  assign y22696 = n30892 ;
  assign y22697 = n25662 ;
  assign y22698 = n30893 ;
  assign y22699 = n30895 ;
  assign y22700 = n30897 ;
  assign y22701 = n22070 ;
  assign y22702 = n30901 ;
  assign y22703 = n30903 ;
  assign y22704 = ~n30907 ;
  assign y22705 = ~1'b0 ;
  assign y22706 = ~1'b0 ;
  assign y22707 = ~n30908 ;
  assign y22708 = ~1'b0 ;
  assign y22709 = ~1'b0 ;
  assign y22710 = ~1'b0 ;
  assign y22711 = n30910 ;
  assign y22712 = ~n30912 ;
  assign y22713 = ~1'b0 ;
  assign y22714 = ~1'b0 ;
  assign y22715 = ~1'b0 ;
  assign y22716 = n30920 ;
  assign y22717 = ~1'b0 ;
  assign y22718 = n30927 ;
  assign y22719 = ~n30930 ;
  assign y22720 = ~1'b0 ;
  assign y22721 = ~1'b0 ;
  assign y22722 = n30932 ;
  assign y22723 = n121 ;
  assign y22724 = ~1'b0 ;
  assign y22725 = ~n30935 ;
  assign y22726 = ~1'b0 ;
  assign y22727 = n30938 ;
  assign y22728 = ~1'b0 ;
  assign y22729 = n30939 ;
  assign y22730 = ~1'b0 ;
  assign y22731 = n26401 ;
  assign y22732 = ~n30942 ;
  assign y22733 = ~1'b0 ;
  assign y22734 = ~n30943 ;
  assign y22735 = ~n30946 ;
  assign y22736 = ~1'b0 ;
  assign y22737 = ~n30948 ;
  assign y22738 = ~1'b0 ;
  assign y22739 = n6644 ;
  assign y22740 = ~n30949 ;
  assign y22741 = ~1'b0 ;
  assign y22742 = n11590 ;
  assign y22743 = n8994 ;
  assign y22744 = ~1'b0 ;
  assign y22745 = ~n30951 ;
  assign y22746 = ~1'b0 ;
  assign y22747 = ~n30954 ;
  assign y22748 = n7449 ;
  assign y22749 = ~1'b0 ;
  assign y22750 = ~1'b0 ;
  assign y22751 = ~n30958 ;
  assign y22752 = ~1'b0 ;
  assign y22753 = n16024 ;
  assign y22754 = ~n30959 ;
  assign y22755 = ~n30960 ;
  assign y22756 = n30961 ;
  assign y22757 = ~1'b0 ;
  assign y22758 = n30965 ;
  assign y22759 = ~1'b0 ;
  assign y22760 = ~n30966 ;
  assign y22761 = ~1'b0 ;
  assign y22762 = n30970 ;
  assign y22763 = ~1'b0 ;
  assign y22764 = ~n30971 ;
  assign y22765 = ~n30972 ;
  assign y22766 = ~n6658 ;
  assign y22767 = ~1'b0 ;
  assign y22768 = ~1'b0 ;
  assign y22769 = 1'b0 ;
  assign y22770 = n30973 ;
  assign y22771 = ~n30975 ;
  assign y22772 = ~1'b0 ;
  assign y22773 = ~n13861 ;
  assign y22774 = ~1'b0 ;
  assign y22775 = n30976 ;
  assign y22776 = n30977 ;
  assign y22777 = ~n10521 ;
  assign y22778 = ~1'b0 ;
  assign y22779 = ~1'b0 ;
  assign y22780 = n30979 ;
  assign y22781 = ~1'b0 ;
  assign y22782 = n30980 ;
  assign y22783 = 1'b0 ;
  assign y22784 = ~n30983 ;
  assign y22785 = ~1'b0 ;
  assign y22786 = n30990 ;
  assign y22787 = n30993 ;
  assign y22788 = n30995 ;
  assign y22789 = ~1'b0 ;
  assign y22790 = ~n30996 ;
  assign y22791 = ~n30998 ;
  assign y22792 = n17537 ;
  assign y22793 = n5564 ;
  assign y22794 = ~1'b0 ;
  assign y22795 = ~1'b0 ;
  assign y22796 = ~1'b0 ;
  assign y22797 = ~n31005 ;
  assign y22798 = n31006 ;
  assign y22799 = ~1'b0 ;
  assign y22800 = ~1'b0 ;
  assign y22801 = n31010 ;
  assign y22802 = ~1'b0 ;
  assign y22803 = ~n6679 ;
  assign y22804 = ~n31012 ;
  assign y22805 = n378 ;
  assign y22806 = ~n31016 ;
  assign y22807 = ~1'b0 ;
  assign y22808 = n31017 ;
  assign y22809 = n31018 ;
  assign y22810 = ~1'b0 ;
  assign y22811 = ~n31021 ;
  assign y22812 = n31022 ;
  assign y22813 = ~n31025 ;
  assign y22814 = n31026 ;
  assign y22815 = ~1'b0 ;
  assign y22816 = n31027 ;
  assign y22817 = n31029 ;
  assign y22818 = ~1'b0 ;
  assign y22819 = n31030 ;
  assign y22820 = ~n31032 ;
  assign y22821 = ~1'b0 ;
  assign y22822 = ~1'b0 ;
  assign y22823 = ~n1518 ;
  assign y22824 = 1'b0 ;
  assign y22825 = ~1'b0 ;
  assign y22826 = ~n31034 ;
  assign y22827 = n10973 ;
  assign y22828 = ~n31035 ;
  assign y22829 = n31039 ;
  assign y22830 = ~n31042 ;
  assign y22831 = ~1'b0 ;
  assign y22832 = n31043 ;
  assign y22833 = ~n10777 ;
  assign y22834 = n8917 ;
  assign y22835 = ~n31044 ;
  assign y22836 = ~n13777 ;
  assign y22837 = ~1'b0 ;
  assign y22838 = ~1'b0 ;
  assign y22839 = ~n31046 ;
  assign y22840 = 1'b0 ;
  assign y22841 = ~n6695 ;
  assign y22842 = ~n31048 ;
  assign y22843 = ~n31049 ;
  assign y22844 = ~1'b0 ;
  assign y22845 = 1'b0 ;
  assign y22846 = n31053 ;
  assign y22847 = ~1'b0 ;
  assign y22848 = ~n1086 ;
  assign y22849 = n31055 ;
  assign y22850 = n31058 ;
  assign y22851 = n31063 ;
  assign y22852 = n94 ;
  assign y22853 = ~n31064 ;
  assign y22854 = ~1'b0 ;
  assign y22855 = ~n31065 ;
  assign y22856 = ~1'b0 ;
  assign y22857 = ~n31066 ;
  assign y22858 = ~1'b0 ;
  assign y22859 = ~n31067 ;
  assign y22860 = n31071 ;
  assign y22861 = ~n31072 ;
  assign y22862 = ~1'b0 ;
  assign y22863 = ~1'b0 ;
  assign y22864 = ~1'b0 ;
  assign y22865 = n31073 ;
  assign y22866 = n31074 ;
  assign y22867 = ~n8320 ;
  assign y22868 = n22233 ;
  assign y22869 = ~1'b0 ;
  assign y22870 = n31075 ;
  assign y22871 = 1'b0 ;
  assign y22872 = ~n31076 ;
  assign y22873 = n31077 ;
  assign y22874 = ~n31083 ;
  assign y22875 = ~1'b0 ;
  assign y22876 = n4300 ;
  assign y22877 = ~n2202 ;
  assign y22878 = ~1'b0 ;
  assign y22879 = ~n31086 ;
  assign y22880 = ~n3037 ;
  assign y22881 = ~n31088 ;
  assign y22882 = ~1'b0 ;
  assign y22883 = n31090 ;
  assign y22884 = ~n4578 ;
  assign y22885 = ~1'b0 ;
  assign y22886 = ~n31091 ;
  assign y22887 = ~1'b0 ;
  assign y22888 = ~n31092 ;
  assign y22889 = n31093 ;
  assign y22890 = ~1'b0 ;
  assign y22891 = ~1'b0 ;
  assign y22892 = ~n7417 ;
  assign y22893 = n462 ;
  assign y22894 = n31094 ;
  assign y22895 = ~n31095 ;
  assign y22896 = ~n31096 ;
  assign y22897 = ~1'b0 ;
  assign y22898 = n31098 ;
  assign y22899 = ~1'b0 ;
  assign y22900 = ~1'b0 ;
  assign y22901 = ~n31100 ;
  assign y22902 = ~1'b0 ;
  assign y22903 = ~1'b0 ;
  assign y22904 = ~n31103 ;
  assign y22905 = ~n31104 ;
  assign y22906 = ~n31105 ;
  assign y22907 = ~1'b0 ;
  assign y22908 = ~1'b0 ;
  assign y22909 = n31109 ;
  assign y22910 = ~1'b0 ;
  assign y22911 = ~1'b0 ;
  assign y22912 = ~n4625 ;
  assign y22913 = n31113 ;
  assign y22914 = ~1'b0 ;
  assign y22915 = ~n31116 ;
  assign y22916 = ~n31117 ;
  assign y22917 = ~1'b0 ;
  assign y22918 = n26940 ;
  assign y22919 = ~1'b0 ;
  assign y22920 = n31120 ;
  assign y22921 = ~1'b0 ;
  assign y22922 = ~n31123 ;
  assign y22923 = ~n31124 ;
  assign y22924 = ~n31126 ;
  assign y22925 = n31127 ;
  assign y22926 = ~1'b0 ;
  assign y22927 = n31131 ;
  assign y22928 = ~n31134 ;
  assign y22929 = ~1'b0 ;
  assign y22930 = 1'b0 ;
  assign y22931 = ~1'b0 ;
  assign y22932 = n31135 ;
  assign y22933 = n31138 ;
  assign y22934 = ~n31143 ;
  assign y22935 = n11308 ;
  assign y22936 = ~1'b0 ;
  assign y22937 = ~1'b0 ;
  assign y22938 = ~1'b0 ;
  assign y22939 = ~1'b0 ;
  assign y22940 = ~n31144 ;
  assign y22941 = ~1'b0 ;
  assign y22942 = n31149 ;
  assign y22943 = ~1'b0 ;
  assign y22944 = ~1'b0 ;
  assign y22945 = n18882 ;
  assign y22946 = ~1'b0 ;
  assign y22947 = n31150 ;
  assign y22948 = n7273 ;
  assign y22949 = n31151 ;
  assign y22950 = ~1'b0 ;
  assign y22951 = ~1'b0 ;
  assign y22952 = ~1'b0 ;
  assign y22953 = ~n31155 ;
  assign y22954 = ~n31157 ;
  assign y22955 = n31158 ;
  assign y22956 = ~n31161 ;
  assign y22957 = n31164 ;
  assign y22958 = 1'b0 ;
  assign y22959 = ~n385 ;
  assign y22960 = ~n14418 ;
  assign y22961 = ~n31165 ;
  assign y22962 = ~1'b0 ;
  assign y22963 = ~n31169 ;
  assign y22964 = ~n31175 ;
  assign y22965 = n31176 ;
  assign y22966 = ~1'b0 ;
  assign y22967 = n31177 ;
  assign y22968 = n31179 ;
  assign y22969 = n31180 ;
  assign y22970 = n31182 ;
  assign y22971 = ~n31183 ;
  assign y22972 = n31185 ;
  assign y22973 = ~1'b0 ;
  assign y22974 = ~n31186 ;
  assign y22975 = ~1'b0 ;
  assign y22976 = n25996 ;
  assign y22977 = ~n31188 ;
  assign y22978 = ~n31190 ;
  assign y22979 = ~1'b0 ;
  assign y22980 = n3237 ;
  assign y22981 = ~n31191 ;
  assign y22982 = n31193 ;
  assign y22983 = n31195 ;
  assign y22984 = n31198 ;
  assign y22985 = n3394 ;
  assign y22986 = n31200 ;
  assign y22987 = n31202 ;
  assign y22988 = ~n31203 ;
  assign y22989 = n31205 ;
  assign y22990 = n31207 ;
  assign y22991 = n11588 ;
  assign y22992 = ~n31208 ;
  assign y22993 = ~1'b0 ;
  assign y22994 = ~n31210 ;
  assign y22995 = ~n31216 ;
  assign y22996 = ~1'b0 ;
  assign y22997 = ~n25783 ;
  assign y22998 = n31217 ;
  assign y22999 = n31220 ;
  assign y23000 = n31223 ;
  assign y23001 = ~n31224 ;
  assign y23002 = 1'b0 ;
  assign y23003 = ~1'b0 ;
  assign y23004 = ~1'b0 ;
  assign y23005 = n31226 ;
  assign y23006 = ~n31227 ;
  assign y23007 = n31231 ;
  assign y23008 = ~n31232 ;
  assign y23009 = n31238 ;
  assign y23010 = ~n31240 ;
  assign y23011 = n31245 ;
  assign y23012 = ~n31246 ;
  assign y23013 = n31247 ;
  assign y23014 = n31248 ;
  assign y23015 = ~n31255 ;
  assign y23016 = ~n31257 ;
  assign y23017 = ~n31258 ;
  assign y23018 = n31259 ;
  assign y23019 = ~n31262 ;
  assign y23020 = n22924 ;
  assign y23021 = ~1'b0 ;
  assign y23022 = ~1'b0 ;
  assign y23023 = n31266 ;
  assign y23024 = ~1'b0 ;
  assign y23025 = n31267 ;
  assign y23026 = n31268 ;
  assign y23027 = ~n10421 ;
  assign y23028 = ~1'b0 ;
  assign y23029 = ~n31270 ;
  assign y23030 = ~n31277 ;
  assign y23031 = ~1'b0 ;
  assign y23032 = ~1'b0 ;
  assign y23033 = n31279 ;
  assign y23034 = 1'b0 ;
  assign y23035 = ~1'b0 ;
  assign y23036 = ~n31281 ;
  assign y23037 = ~1'b0 ;
  assign y23038 = ~1'b0 ;
  assign y23039 = ~n2896 ;
  assign y23040 = ~n31282 ;
  assign y23041 = ~n31283 ;
  assign y23042 = ~1'b0 ;
  assign y23043 = ~1'b0 ;
  assign y23044 = ~1'b0 ;
  assign y23045 = n31284 ;
  assign y23046 = n31286 ;
  assign y23047 = ~1'b0 ;
  assign y23048 = ~1'b0 ;
  assign y23049 = 1'b0 ;
  assign y23050 = ~1'b0 ;
  assign y23051 = n31289 ;
  assign y23052 = n31291 ;
  assign y23053 = n31295 ;
  assign y23054 = ~1'b0 ;
  assign y23055 = ~n31297 ;
  assign y23056 = ~1'b0 ;
  assign y23057 = n31298 ;
  assign y23058 = ~n31299 ;
  assign y23059 = ~n5271 ;
  assign y23060 = ~1'b0 ;
  assign y23061 = n31304 ;
  assign y23062 = n6360 ;
  assign y23063 = ~1'b0 ;
  assign y23064 = n31306 ;
  assign y23065 = n31309 ;
  assign y23066 = ~1'b0 ;
  assign y23067 = ~1'b0 ;
  assign y23068 = ~1'b0 ;
  assign y23069 = ~n24611 ;
  assign y23070 = ~n2759 ;
  assign y23071 = ~n24598 ;
  assign y23072 = ~n31313 ;
  assign y23073 = ~n31315 ;
  assign y23074 = ~1'b0 ;
  assign y23075 = ~1'b0 ;
  assign y23076 = n15787 ;
  assign y23077 = ~1'b0 ;
  assign y23078 = ~1'b0 ;
  assign y23079 = ~1'b0 ;
  assign y23080 = ~1'b0 ;
  assign y23081 = n31316 ;
  assign y23082 = ~n31322 ;
  assign y23083 = ~n31324 ;
  assign y23084 = n31325 ;
  assign y23085 = ~1'b0 ;
  assign y23086 = n12468 ;
  assign y23087 = ~n31326 ;
  assign y23088 = ~1'b0 ;
  assign y23089 = ~1'b0 ;
  assign y23090 = ~1'b0 ;
  assign y23091 = ~n31329 ;
  assign y23092 = n31330 ;
  assign y23093 = n31332 ;
  assign y23094 = ~1'b0 ;
  assign y23095 = ~1'b0 ;
  assign y23096 = ~n31334 ;
  assign y23097 = ~n27408 ;
  assign y23098 = ~n31336 ;
  assign y23099 = n1416 ;
  assign y23100 = ~n31339 ;
  assign y23101 = n31343 ;
  assign y23102 = n31344 ;
  assign y23103 = ~n31345 ;
  assign y23104 = ~1'b0 ;
  assign y23105 = ~n31346 ;
  assign y23106 = ~1'b0 ;
  assign y23107 = ~n31348 ;
  assign y23108 = n31349 ;
  assign y23109 = n7459 ;
  assign y23110 = n31350 ;
  assign y23111 = n31351 ;
  assign y23112 = ~1'b0 ;
  assign y23113 = ~1'b0 ;
  assign y23114 = n31352 ;
  assign y23115 = ~1'b0 ;
  assign y23116 = n31353 ;
  assign y23117 = ~n31354 ;
  assign y23118 = n31359 ;
  assign y23119 = n31364 ;
  assign y23120 = n31366 ;
  assign y23121 = ~1'b0 ;
  assign y23122 = n31368 ;
  assign y23123 = ~n31369 ;
  assign y23124 = ~n31371 ;
  assign y23125 = n31372 ;
  assign y23126 = n31373 ;
  assign y23127 = ~n7949 ;
  assign y23128 = ~1'b0 ;
  assign y23129 = ~1'b0 ;
  assign y23130 = n31378 ;
  assign y23131 = 1'b0 ;
  assign y23132 = ~n2817 ;
  assign y23133 = ~n31379 ;
  assign y23134 = ~1'b0 ;
  assign y23135 = 1'b0 ;
  assign y23136 = n9439 ;
  assign y23137 = ~1'b0 ;
  assign y23138 = ~n31381 ;
  assign y23139 = n18288 ;
  assign y23140 = ~1'b0 ;
  assign y23141 = ~1'b0 ;
  assign y23142 = n31382 ;
  assign y23143 = ~n241 ;
  assign y23144 = ~1'b0 ;
  assign y23145 = ~n31384 ;
  assign y23146 = 1'b0 ;
  assign y23147 = ~n31386 ;
  assign y23148 = ~1'b0 ;
  assign y23149 = ~1'b0 ;
  assign y23150 = n16827 ;
  assign y23151 = 1'b0 ;
  assign y23152 = ~1'b0 ;
  assign y23153 = n31388 ;
  assign y23154 = n31389 ;
  assign y23155 = ~1'b0 ;
  assign y23156 = ~1'b0 ;
  assign y23157 = ~n31402 ;
  assign y23158 = ~n31404 ;
  assign y23159 = ~n31405 ;
  assign y23160 = ~1'b0 ;
  assign y23161 = n31406 ;
  assign y23162 = n31410 ;
  assign y23163 = n31414 ;
  assign y23164 = n31415 ;
  assign y23165 = ~n31417 ;
  assign y23166 = ~1'b0 ;
  assign y23167 = ~n31419 ;
  assign y23168 = n31420 ;
  assign y23169 = ~1'b0 ;
  assign y23170 = n31424 ;
  assign y23171 = ~1'b0 ;
  assign y23172 = ~1'b0 ;
  assign y23173 = ~n31427 ;
  assign y23174 = n8040 ;
  assign y23175 = n31429 ;
  assign y23176 = n7450 ;
  assign y23177 = ~n31430 ;
  assign y23178 = n31431 ;
  assign y23179 = n31436 ;
  assign y23180 = ~n31438 ;
  assign y23181 = ~1'b0 ;
  assign y23182 = ~n1790 ;
  assign y23183 = n31441 ;
  assign y23184 = n31443 ;
  assign y23185 = ~1'b0 ;
  assign y23186 = ~n31448 ;
  assign y23187 = n31449 ;
  assign y23188 = n31451 ;
  assign y23189 = ~1'b0 ;
  assign y23190 = ~1'b0 ;
  assign y23191 = n31452 ;
  assign y23192 = n31453 ;
  assign y23193 = ~n31455 ;
  assign y23194 = ~1'b0 ;
  assign y23195 = ~n31456 ;
  assign y23196 = 1'b0 ;
  assign y23197 = n31460 ;
  assign y23198 = n31461 ;
  assign y23199 = n31463 ;
  assign y23200 = ~1'b0 ;
  assign y23201 = n31464 ;
  assign y23202 = ~1'b0 ;
  assign y23203 = ~n31467 ;
  assign y23204 = n19371 ;
  assign y23205 = n7606 ;
  assign y23206 = ~1'b0 ;
  assign y23207 = n31468 ;
  assign y23208 = n31469 ;
  assign y23209 = ~n31473 ;
  assign y23210 = n31477 ;
  assign y23211 = ~n31479 ;
  assign y23212 = ~n31481 ;
  assign y23213 = ~1'b0 ;
  assign y23214 = ~1'b0 ;
  assign y23215 = n2842 ;
  assign y23216 = ~n31482 ;
  assign y23217 = ~n31483 ;
  assign y23218 = n31486 ;
  assign y23219 = ~1'b0 ;
  assign y23220 = ~n31491 ;
  assign y23221 = ~1'b0 ;
  assign y23222 = n31495 ;
  assign y23223 = n31496 ;
  assign y23224 = ~1'b0 ;
  assign y23225 = n24520 ;
  assign y23226 = n19735 ;
  assign y23227 = n31497 ;
  assign y23228 = n31498 ;
  assign y23229 = ~n31499 ;
  assign y23230 = ~1'b0 ;
  assign y23231 = n31502 ;
  assign y23232 = ~1'b0 ;
  assign y23233 = ~n31505 ;
  assign y23234 = n11178 ;
  assign y23235 = n31508 ;
  assign y23236 = ~n31509 ;
  assign y23237 = ~n31510 ;
  assign y23238 = n31511 ;
  assign y23239 = ~n31512 ;
  assign y23240 = ~1'b0 ;
  assign y23241 = 1'b0 ;
  assign y23242 = ~1'b0 ;
  assign y23243 = ~n31517 ;
  assign y23244 = n31518 ;
  assign y23245 = ~1'b0 ;
  assign y23246 = n31519 ;
  assign y23247 = n14622 ;
  assign y23248 = ~n31522 ;
  assign y23249 = ~n9702 ;
  assign y23250 = n29486 ;
  assign y23251 = ~1'b0 ;
  assign y23252 = n31523 ;
  assign y23253 = 1'b0 ;
  assign y23254 = ~n24816 ;
  assign y23255 = ~n31526 ;
  assign y23256 = n14674 ;
  assign y23257 = ~n31528 ;
  assign y23258 = ~n31529 ;
  assign y23259 = ~1'b0 ;
  assign y23260 = ~1'b0 ;
  assign y23261 = n31532 ;
  assign y23262 = n13775 ;
  assign y23263 = ~1'b0 ;
  assign y23264 = ~1'b0 ;
  assign y23265 = n18317 ;
  assign y23266 = n17021 ;
  assign y23267 = ~1'b0 ;
  assign y23268 = ~1'b0 ;
  assign y23269 = ~n31539 ;
  assign y23270 = ~n31540 ;
  assign y23271 = n10992 ;
  assign y23272 = ~n9245 ;
  assign y23273 = ~n31542 ;
  assign y23274 = n31543 ;
  assign y23275 = 1'b0 ;
  assign y23276 = ~1'b0 ;
  assign y23277 = ~n31545 ;
  assign y23278 = ~1'b0 ;
  assign y23279 = ~1'b0 ;
  assign y23280 = n31550 ;
  assign y23281 = ~1'b0 ;
  assign y23282 = n31551 ;
  assign y23283 = ~n31555 ;
  assign y23284 = ~n31557 ;
  assign y23285 = ~n31558 ;
  assign y23286 = ~1'b0 ;
  assign y23287 = ~1'b0 ;
  assign y23288 = n2075 ;
  assign y23289 = ~1'b0 ;
  assign y23290 = 1'b0 ;
  assign y23291 = ~1'b0 ;
  assign y23292 = ~n31560 ;
  assign y23293 = ~1'b0 ;
  assign y23294 = ~n31562 ;
  assign y23295 = n31567 ;
  assign y23296 = n31568 ;
  assign y23297 = ~n31573 ;
  assign y23298 = ~n31576 ;
  assign y23299 = n31577 ;
  assign y23300 = ~n31579 ;
  assign y23301 = ~n31603 ;
  assign y23302 = 1'b0 ;
  assign y23303 = ~n31604 ;
  assign y23304 = ~n31607 ;
  assign y23305 = ~n6486 ;
  assign y23306 = n29468 ;
  assign y23307 = ~n6084 ;
  assign y23308 = n31609 ;
  assign y23309 = ~n31612 ;
  assign y23310 = ~1'b0 ;
  assign y23311 = ~1'b0 ;
  assign y23312 = n31614 ;
  assign y23313 = ~1'b0 ;
  assign y23314 = n31616 ;
  assign y23315 = ~1'b0 ;
  assign y23316 = ~n1300 ;
  assign y23317 = ~n31619 ;
  assign y23318 = ~n31623 ;
  assign y23319 = ~n31626 ;
  assign y23320 = ~n31627 ;
  assign y23321 = ~n31628 ;
  assign y23322 = n1328 ;
  assign y23323 = ~1'b0 ;
  assign y23324 = n31632 ;
  assign y23325 = ~1'b0 ;
  assign y23326 = ~1'b0 ;
  assign y23327 = ~n31633 ;
  assign y23328 = n31638 ;
  assign y23329 = n31639 ;
  assign y23330 = ~1'b0 ;
  assign y23331 = ~1'b0 ;
  assign y23332 = ~1'b0 ;
  assign y23333 = ~n31640 ;
  assign y23334 = n31641 ;
  assign y23335 = n31644 ;
  assign y23336 = ~n31648 ;
  assign y23337 = ~1'b0 ;
  assign y23338 = ~1'b0 ;
  assign y23339 = ~n31651 ;
  assign y23340 = n31652 ;
  assign y23341 = n31653 ;
  assign y23342 = n31659 ;
  assign y23343 = ~n31662 ;
  assign y23344 = ~1'b0 ;
  assign y23345 = ~n31663 ;
  assign y23346 = ~1'b0 ;
  assign y23347 = ~n13901 ;
  assign y23348 = ~1'b0 ;
  assign y23349 = ~1'b0 ;
  assign y23350 = n31669 ;
  assign y23351 = n31671 ;
  assign y23352 = ~n31673 ;
  assign y23353 = ~1'b0 ;
  assign y23354 = ~n31674 ;
  assign y23355 = ~n31676 ;
  assign y23356 = ~1'b0 ;
  assign y23357 = ~1'b0 ;
  assign y23358 = n31677 ;
  assign y23359 = ~1'b0 ;
  assign y23360 = ~1'b0 ;
  assign y23361 = n18836 ;
  assign y23362 = ~1'b0 ;
  assign y23363 = ~n31680 ;
  assign y23364 = ~1'b0 ;
  assign y23365 = ~1'b0 ;
  assign y23366 = ~1'b0 ;
  assign y23367 = ~n31682 ;
  assign y23368 = ~n31683 ;
  assign y23369 = n31687 ;
  assign y23370 = 1'b0 ;
  assign y23371 = 1'b0 ;
  assign y23372 = n31691 ;
  assign y23373 = ~n31692 ;
  assign y23374 = ~1'b0 ;
  assign y23375 = ~1'b0 ;
  assign y23376 = n31696 ;
  assign y23377 = ~n31700 ;
  assign y23378 = ~n31702 ;
  assign y23379 = n4327 ;
  assign y23380 = ~1'b0 ;
  assign y23381 = ~1'b0 ;
  assign y23382 = n31703 ;
  assign y23383 = n31704 ;
  assign y23384 = ~1'b0 ;
  assign y23385 = ~1'b0 ;
  assign y23386 = n31705 ;
  assign y23387 = 1'b0 ;
  assign y23388 = ~1'b0 ;
  assign y23389 = n31708 ;
  assign y23390 = n26707 ;
  assign y23391 = ~1'b0 ;
  assign y23392 = n31709 ;
  assign y23393 = n31711 ;
  assign y23394 = n31712 ;
  assign y23395 = ~n31713 ;
  assign y23396 = ~1'b0 ;
  assign y23397 = ~n31716 ;
  assign y23398 = ~1'b0 ;
  assign y23399 = ~n31717 ;
  assign y23400 = ~n31718 ;
  assign y23401 = ~1'b0 ;
  assign y23402 = n31723 ;
  assign y23403 = ~n31726 ;
  assign y23404 = ~n31730 ;
  assign y23405 = ~n31732 ;
  assign y23406 = n31734 ;
  assign y23407 = ~1'b0 ;
  assign y23408 = ~1'b0 ;
  assign y23409 = n31737 ;
  assign y23410 = ~1'b0 ;
  assign y23411 = ~1'b0 ;
  assign y23412 = ~n31739 ;
  assign y23413 = n31740 ;
  assign y23414 = ~n31742 ;
  assign y23415 = ~1'b0 ;
  assign y23416 = ~1'b0 ;
  assign y23417 = ~n31745 ;
  assign y23418 = ~1'b0 ;
  assign y23419 = ~1'b0 ;
  assign y23420 = ~1'b0 ;
  assign y23421 = ~n31746 ;
  assign y23422 = ~n31747 ;
  assign y23423 = ~n6279 ;
  assign y23424 = ~n31748 ;
  assign y23425 = 1'b0 ;
  assign y23426 = ~n31749 ;
  assign y23427 = ~1'b0 ;
  assign y23428 = n31753 ;
  assign y23429 = n31755 ;
  assign y23430 = n31759 ;
  assign y23431 = n31760 ;
  assign y23432 = n31761 ;
  assign y23433 = n31764 ;
  assign y23434 = ~1'b0 ;
  assign y23435 = n31768 ;
  assign y23436 = n31770 ;
  assign y23437 = n31772 ;
  assign y23438 = ~n31773 ;
  assign y23439 = ~1'b0 ;
  assign y23440 = n21399 ;
  assign y23441 = n31774 ;
  assign y23442 = ~n1394 ;
  assign y23443 = ~1'b0 ;
  assign y23444 = 1'b0 ;
  assign y23445 = ~1'b0 ;
  assign y23446 = ~1'b0 ;
  assign y23447 = n31782 ;
  assign y23448 = ~1'b0 ;
  assign y23449 = ~1'b0 ;
  assign y23450 = ~n31785 ;
  assign y23451 = ~n31788 ;
  assign y23452 = ~n31789 ;
  assign y23453 = ~n31792 ;
  assign y23454 = n9451 ;
  assign y23455 = ~1'b0 ;
  assign y23456 = ~1'b0 ;
  assign y23457 = ~1'b0 ;
  assign y23458 = n31796 ;
  assign y23459 = n31797 ;
  assign y23460 = ~n31798 ;
  assign y23461 = ~1'b0 ;
  assign y23462 = ~n31804 ;
  assign y23463 = n818 ;
  assign y23464 = n31805 ;
  assign y23465 = ~1'b0 ;
  assign y23466 = n31806 ;
  assign y23467 = ~n31807 ;
  assign y23468 = ~1'b0 ;
  assign y23469 = ~n31808 ;
  assign y23470 = n15038 ;
  assign y23471 = n30248 ;
  assign y23472 = 1'b0 ;
  assign y23473 = ~n31813 ;
  assign y23474 = ~1'b0 ;
  assign y23475 = ~1'b0 ;
  assign y23476 = ~1'b0 ;
  assign y23477 = ~1'b0 ;
  assign y23478 = ~1'b0 ;
  assign y23479 = n31818 ;
  assign y23480 = n31821 ;
  assign y23481 = n31822 ;
  assign y23482 = ~1'b0 ;
  assign y23483 = ~1'b0 ;
  assign y23484 = n31828 ;
  assign y23485 = ~n25051 ;
  assign y23486 = n31829 ;
  assign y23487 = n31830 ;
  assign y23488 = ~1'b0 ;
  assign y23489 = n31832 ;
  assign y23490 = ~1'b0 ;
  assign y23491 = ~1'b0 ;
  assign y23492 = ~1'b0 ;
  assign y23493 = n31834 ;
  assign y23494 = n31836 ;
  assign y23495 = n5002 ;
  assign y23496 = ~1'b0 ;
  assign y23497 = ~n31838 ;
  assign y23498 = n31839 ;
  assign y23499 = ~1'b0 ;
  assign y23500 = n31840 ;
  assign y23501 = 1'b0 ;
  assign y23502 = ~n31842 ;
  assign y23503 = ~1'b0 ;
  assign y23504 = ~n31844 ;
  assign y23505 = ~1'b0 ;
  assign y23506 = n31846 ;
  assign y23507 = ~1'b0 ;
  assign y23508 = ~1'b0 ;
  assign y23509 = ~1'b0 ;
  assign y23510 = n31848 ;
  assign y23511 = ~n4337 ;
  assign y23512 = n4924 ;
  assign y23513 = ~1'b0 ;
  assign y23514 = n31850 ;
  assign y23515 = n27807 ;
  assign y23516 = n31852 ;
  assign y23517 = 1'b0 ;
  assign y23518 = n31853 ;
  assign y23519 = ~1'b0 ;
  assign y23520 = n31855 ;
  assign y23521 = n31859 ;
  assign y23522 = ~1'b0 ;
  assign y23523 = ~1'b0 ;
  assign y23524 = ~n31860 ;
  assign y23525 = n31863 ;
  assign y23526 = ~n31877 ;
  assign y23527 = ~1'b0 ;
  assign y23528 = ~1'b0 ;
  assign y23529 = n31878 ;
  assign y23530 = ~n1015 ;
  assign y23531 = 1'b0 ;
  assign y23532 = n31879 ;
  assign y23533 = ~1'b0 ;
  assign y23534 = ~1'b0 ;
  assign y23535 = n31885 ;
  assign y23536 = ~n31887 ;
  assign y23537 = ~n31888 ;
  assign y23538 = ~1'b0 ;
  assign y23539 = ~n31891 ;
  assign y23540 = n31893 ;
  assign y23541 = ~1'b0 ;
  assign y23542 = ~n31896 ;
  assign y23543 = n31898 ;
  assign y23544 = 1'b0 ;
  assign y23545 = ~1'b0 ;
  assign y23546 = ~n31900 ;
  assign y23547 = ~1'b0 ;
  assign y23548 = ~1'b0 ;
  assign y23549 = ~n31903 ;
  assign y23550 = n31905 ;
  assign y23551 = ~n31907 ;
  assign y23552 = n31908 ;
  assign y23553 = ~1'b0 ;
  assign y23554 = ~n31910 ;
  assign y23555 = ~1'b0 ;
  assign y23556 = ~n31913 ;
  assign y23557 = ~n31914 ;
  assign y23558 = ~1'b0 ;
  assign y23559 = n31917 ;
  assign y23560 = ~n31919 ;
  assign y23561 = ~1'b0 ;
  assign y23562 = ~n31920 ;
  assign y23563 = ~n31921 ;
  assign y23564 = ~n31925 ;
  assign y23565 = ~n31927 ;
  assign y23566 = ~n31930 ;
  assign y23567 = ~1'b0 ;
  assign y23568 = ~1'b0 ;
  assign y23569 = ~1'b0 ;
  assign y23570 = ~1'b0 ;
  assign y23571 = n31934 ;
  assign y23572 = ~1'b0 ;
  assign y23573 = n31936 ;
  assign y23574 = n31938 ;
  assign y23575 = n31939 ;
  assign y23576 = ~1'b0 ;
  assign y23577 = ~n31941 ;
  assign y23578 = ~1'b0 ;
  assign y23579 = ~n31942 ;
  assign y23580 = ~n31943 ;
  assign y23581 = ~n31950 ;
  assign y23582 = n31952 ;
  assign y23583 = ~1'b0 ;
  assign y23584 = ~n31953 ;
  assign y23585 = n20027 ;
  assign y23586 = ~n1034 ;
  assign y23587 = n31955 ;
  assign y23588 = ~1'b0 ;
  assign y23589 = ~1'b0 ;
  assign y23590 = 1'b0 ;
  assign y23591 = ~1'b0 ;
  assign y23592 = ~n13277 ;
  assign y23593 = ~1'b0 ;
  assign y23594 = n31958 ;
  assign y23595 = n31961 ;
  assign y23596 = ~1'b0 ;
  assign y23597 = ~1'b0 ;
  assign y23598 = n31962 ;
  assign y23599 = ~1'b0 ;
  assign y23600 = n31966 ;
  assign y23601 = ~n31968 ;
  assign y23602 = ~n935 ;
  assign y23603 = ~1'b0 ;
  assign y23604 = ~n31969 ;
  assign y23605 = ~1'b0 ;
  assign y23606 = n31975 ;
  assign y23607 = n31978 ;
  assign y23608 = ~n21456 ;
  assign y23609 = ~1'b0 ;
  assign y23610 = n20508 ;
  assign y23611 = ~n31980 ;
  assign y23612 = n31981 ;
  assign y23613 = ~n21173 ;
  assign y23614 = n10719 ;
  assign y23615 = ~1'b0 ;
  assign y23616 = ~n31982 ;
  assign y23617 = ~n5205 ;
  assign y23618 = n13990 ;
  assign y23619 = ~1'b0 ;
  assign y23620 = n31984 ;
  assign y23621 = n31985 ;
  assign y23622 = ~n31986 ;
  assign y23623 = n31991 ;
  assign y23624 = ~1'b0 ;
  assign y23625 = ~n31996 ;
  assign y23626 = ~n32000 ;
  assign y23627 = ~1'b0 ;
  assign y23628 = ~1'b0 ;
  assign y23629 = ~n9843 ;
  assign y23630 = ~n32001 ;
  assign y23631 = ~1'b0 ;
  assign y23632 = ~n167 ;
  assign y23633 = n32002 ;
  assign y23634 = n32003 ;
  assign y23635 = ~n158 ;
  assign y23636 = ~1'b0 ;
  assign y23637 = ~n32005 ;
  assign y23638 = ~n32008 ;
  assign y23639 = ~1'b0 ;
  assign y23640 = ~1'b0 ;
  assign y23641 = n32009 ;
  assign y23642 = ~1'b0 ;
  assign y23643 = n32012 ;
  assign y23644 = n32014 ;
  assign y23645 = 1'b0 ;
  assign y23646 = n32015 ;
  assign y23647 = ~n32022 ;
  assign y23648 = ~1'b0 ;
  assign y23649 = n32024 ;
  assign y23650 = ~1'b0 ;
  assign y23651 = ~n32025 ;
  assign y23652 = ~1'b0 ;
  assign y23653 = ~1'b0 ;
  assign y23654 = ~n2083 ;
  assign y23655 = ~1'b0 ;
  assign y23656 = ~1'b0 ;
  assign y23657 = ~1'b0 ;
  assign y23658 = n32028 ;
  assign y23659 = n32037 ;
  assign y23660 = ~1'b0 ;
  assign y23661 = ~1'b0 ;
  assign y23662 = n32042 ;
  assign y23663 = ~1'b0 ;
  assign y23664 = ~n19175 ;
  assign y23665 = n32043 ;
  assign y23666 = ~1'b0 ;
  assign y23667 = ~n32046 ;
  assign y23668 = ~1'b0 ;
  assign y23669 = n32047 ;
  assign y23670 = n32048 ;
  assign y23671 = ~1'b0 ;
  assign y23672 = ~1'b0 ;
  assign y23673 = ~n32050 ;
  assign y23674 = ~1'b0 ;
  assign y23675 = n32054 ;
  assign y23676 = ~1'b0 ;
  assign y23677 = ~1'b0 ;
  assign y23678 = ~n8016 ;
  assign y23679 = n32055 ;
  assign y23680 = ~n32056 ;
  assign y23681 = ~1'b0 ;
  assign y23682 = n32057 ;
  assign y23683 = n32058 ;
  assign y23684 = ~n7811 ;
  assign y23685 = n32059 ;
  assign y23686 = 1'b0 ;
  assign y23687 = ~1'b0 ;
  assign y23688 = n32062 ;
  assign y23689 = ~1'b0 ;
  assign y23690 = ~n32063 ;
  assign y23691 = ~n32064 ;
  assign y23692 = ~n32065 ;
  assign y23693 = ~1'b0 ;
  assign y23694 = ~n32067 ;
  assign y23695 = ~n15430 ;
  assign y23696 = ~n32069 ;
  assign y23697 = ~n32072 ;
  assign y23698 = ~1'b0 ;
  assign y23699 = ~1'b0 ;
  assign y23700 = ~1'b0 ;
  assign y23701 = ~1'b0 ;
  assign y23702 = 1'b0 ;
  assign y23703 = ~1'b0 ;
  assign y23704 = ~n32075 ;
  assign y23705 = ~n32077 ;
  assign y23706 = 1'b0 ;
  assign y23707 = ~n32080 ;
  assign y23708 = ~n5857 ;
  assign y23709 = 1'b0 ;
  assign y23710 = ~n22777 ;
  assign y23711 = ~n32083 ;
  assign y23712 = n32084 ;
  assign y23713 = 1'b0 ;
  assign y23714 = ~1'b0 ;
  assign y23715 = ~1'b0 ;
  assign y23716 = n32088 ;
  assign y23717 = ~1'b0 ;
  assign y23718 = 1'b0 ;
  assign y23719 = ~1'b0 ;
  assign y23720 = n32095 ;
  assign y23721 = ~n30080 ;
  assign y23722 = n3820 ;
  assign y23723 = n32098 ;
  assign y23724 = n32099 ;
  assign y23725 = ~n32102 ;
  assign y23726 = ~n15183 ;
  assign y23727 = n32104 ;
  assign y23728 = ~1'b0 ;
  assign y23729 = ~1'b0 ;
  assign y23730 = ~1'b0 ;
  assign y23731 = n32105 ;
  assign y23732 = 1'b0 ;
  assign y23733 = n24602 ;
  assign y23734 = n32106 ;
  assign y23735 = ~n1740 ;
  assign y23736 = ~n32108 ;
  assign y23737 = ~1'b0 ;
  assign y23738 = ~1'b0 ;
  assign y23739 = n32109 ;
  assign y23740 = ~1'b0 ;
  assign y23741 = n2644 ;
  assign y23742 = ~1'b0 ;
  assign y23743 = ~1'b0 ;
  assign y23744 = ~1'b0 ;
  assign y23745 = ~1'b0 ;
  assign y23746 = ~1'b0 ;
  assign y23747 = ~n4597 ;
  assign y23748 = ~n32110 ;
  assign y23749 = n32111 ;
  assign y23750 = ~n32116 ;
  assign y23751 = ~1'b0 ;
  assign y23752 = n32120 ;
  assign y23753 = ~1'b0 ;
  assign y23754 = ~n32122 ;
  assign y23755 = n32125 ;
  assign y23756 = ~n32128 ;
  assign y23757 = n32129 ;
  assign y23758 = ~n32131 ;
  assign y23759 = ~n32132 ;
  assign y23760 = ~1'b0 ;
  assign y23761 = n32136 ;
  assign y23762 = ~1'b0 ;
  assign y23763 = n32137 ;
  assign y23764 = ~1'b0 ;
  assign y23765 = n32140 ;
  assign y23766 = ~n32142 ;
  assign y23767 = n32146 ;
  assign y23768 = n6875 ;
  assign y23769 = ~1'b0 ;
  assign y23770 = ~1'b0 ;
  assign y23771 = ~1'b0 ;
  assign y23772 = n32147 ;
  assign y23773 = ~n10578 ;
  assign y23774 = n10853 ;
  assign y23775 = ~1'b0 ;
  assign y23776 = ~1'b0 ;
  assign y23777 = ~n32149 ;
  assign y23778 = ~1'b0 ;
  assign y23779 = n32156 ;
  assign y23780 = ~n32158 ;
  assign y23781 = ~1'b0 ;
  assign y23782 = n12229 ;
  assign y23783 = ~1'b0 ;
  assign y23784 = n32159 ;
  assign y23785 = ~n32160 ;
  assign y23786 = ~n11438 ;
  assign y23787 = n32162 ;
  assign y23788 = ~1'b0 ;
  assign y23789 = ~n32163 ;
  assign y23790 = ~n22273 ;
  assign y23791 = ~n32169 ;
  assign y23792 = ~n17617 ;
  assign y23793 = n12494 ;
  assign y23794 = n32174 ;
  assign y23795 = ~1'b0 ;
  assign y23796 = ~1'b0 ;
  assign y23797 = ~n32177 ;
  assign y23798 = ~n32178 ;
  assign y23799 = ~1'b0 ;
  assign y23800 = ~n32181 ;
  assign y23801 = ~n32183 ;
  assign y23802 = ~1'b0 ;
  assign y23803 = ~1'b0 ;
  assign y23804 = n32184 ;
  assign y23805 = ~n32185 ;
  assign y23806 = ~1'b0 ;
  assign y23807 = ~n32186 ;
  assign y23808 = n32187 ;
  assign y23809 = n32188 ;
  assign y23810 = n32190 ;
  assign y23811 = n32192 ;
  assign y23812 = ~n32196 ;
  assign y23813 = n32204 ;
  assign y23814 = n32206 ;
  assign y23815 = ~n32210 ;
  assign y23816 = n32212 ;
  assign y23817 = ~1'b0 ;
  assign y23818 = n32213 ;
  assign y23819 = n32214 ;
  assign y23820 = ~n32216 ;
  assign y23821 = n32217 ;
  assign y23822 = ~n32221 ;
  assign y23823 = ~n32233 ;
  assign y23824 = ~1'b0 ;
  assign y23825 = ~n32238 ;
  assign y23826 = ~n32243 ;
  assign y23827 = ~n18845 ;
  assign y23828 = n32245 ;
  assign y23829 = ~n32248 ;
  assign y23830 = ~1'b0 ;
  assign y23831 = ~1'b0 ;
  assign y23832 = n12020 ;
  assign y23833 = ~n32249 ;
  assign y23834 = ~1'b0 ;
  assign y23835 = ~n32251 ;
  assign y23836 = n32252 ;
  assign y23837 = n32256 ;
  assign y23838 = ~n32257 ;
  assign y23839 = n32039 ;
  assign y23840 = ~n32258 ;
  assign y23841 = ~1'b0 ;
  assign y23842 = 1'b0 ;
  assign y23843 = ~1'b0 ;
  assign y23844 = n32259 ;
  assign y23845 = ~1'b0 ;
  assign y23846 = ~1'b0 ;
  assign y23847 = ~n10157 ;
  assign y23848 = n17861 ;
  assign y23849 = ~1'b0 ;
  assign y23850 = ~n32260 ;
  assign y23851 = ~1'b0 ;
  assign y23852 = n32261 ;
  assign y23853 = ~1'b0 ;
  assign y23854 = ~1'b0 ;
  assign y23855 = ~1'b0 ;
  assign y23856 = n32263 ;
  assign y23857 = ~n32264 ;
  assign y23858 = ~1'b0 ;
  assign y23859 = n32274 ;
  assign y23860 = ~n4970 ;
  assign y23861 = ~1'b0 ;
  assign y23862 = n32277 ;
  assign y23863 = ~1'b0 ;
  assign y23864 = ~n32285 ;
  assign y23865 = ~1'b0 ;
  assign y23866 = n32286 ;
  assign y23867 = ~n32289 ;
  assign y23868 = ~n32291 ;
  assign y23869 = ~n31065 ;
  assign y23870 = ~1'b0 ;
  assign y23871 = n32293 ;
  assign y23872 = n32294 ;
  assign y23873 = n32296 ;
  assign y23874 = ~1'b0 ;
  assign y23875 = ~n32301 ;
  assign y23876 = ~1'b0 ;
  assign y23877 = ~n32303 ;
  assign y23878 = ~1'b0 ;
  assign y23879 = ~1'b0 ;
  assign y23880 = n27441 ;
  assign y23881 = ~1'b0 ;
  assign y23882 = n32308 ;
  assign y23883 = ~1'b0 ;
  assign y23884 = ~n32315 ;
  assign y23885 = ~1'b0 ;
  assign y23886 = ~n128 ;
  assign y23887 = n32316 ;
  assign y23888 = n32320 ;
  assign y23889 = ~1'b0 ;
  assign y23890 = ~n32322 ;
  assign y23891 = ~1'b0 ;
  assign y23892 = ~n32325 ;
  assign y23893 = ~1'b0 ;
  assign y23894 = n32326 ;
  assign y23895 = ~n31161 ;
  assign y23896 = ~n26955 ;
  assign y23897 = ~n32327 ;
  assign y23898 = ~1'b0 ;
  assign y23899 = ~n32329 ;
  assign y23900 = ~n32330 ;
  assign y23901 = ~n2835 ;
  assign y23902 = n32331 ;
  assign y23903 = ~n32332 ;
  assign y23904 = ~1'b0 ;
  assign y23905 = ~1'b0 ;
  assign y23906 = ~1'b0 ;
  assign y23907 = ~1'b0 ;
  assign y23908 = ~n32333 ;
  assign y23909 = ~n32334 ;
  assign y23910 = n32337 ;
  assign y23911 = ~1'b0 ;
  assign y23912 = n1344 ;
  assign y23913 = ~1'b0 ;
  assign y23914 = ~n32340 ;
  assign y23915 = ~1'b0 ;
  assign y23916 = ~n32342 ;
  assign y23917 = ~n32343 ;
  assign y23918 = ~1'b0 ;
  assign y23919 = ~1'b0 ;
  assign y23920 = ~n32344 ;
  assign y23921 = ~1'b0 ;
  assign y23922 = ~1'b0 ;
  assign y23923 = ~n32345 ;
  assign y23924 = ~1'b0 ;
  assign y23925 = ~n32348 ;
  assign y23926 = n32351 ;
  assign y23927 = ~n32353 ;
  assign y23928 = ~n32354 ;
  assign y23929 = n32355 ;
  assign y23930 = ~1'b0 ;
  assign y23931 = ~1'b0 ;
  assign y23932 = n8539 ;
  assign y23933 = n32356 ;
  assign y23934 = ~1'b0 ;
  assign y23935 = ~n32363 ;
  assign y23936 = ~n32365 ;
  assign y23937 = ~1'b0 ;
  assign y23938 = ~n32367 ;
  assign y23939 = ~n608 ;
  assign y23940 = n32369 ;
  assign y23941 = n32371 ;
  assign y23942 = 1'b0 ;
  assign y23943 = n13397 ;
  assign y23944 = ~1'b0 ;
  assign y23945 = ~n32372 ;
  assign y23946 = ~n32374 ;
  assign y23947 = n32376 ;
  assign y23948 = ~1'b0 ;
  assign y23949 = ~1'b0 ;
  assign y23950 = ~n32381 ;
  assign y23951 = ~n32382 ;
  assign y23952 = ~1'b0 ;
  assign y23953 = ~1'b0 ;
  assign y23954 = ~1'b0 ;
  assign y23955 = n32383 ;
  assign y23956 = ~n32384 ;
  assign y23957 = ~1'b0 ;
  assign y23958 = ~1'b0 ;
  assign y23959 = ~1'b0 ;
  assign y23960 = ~n1284 ;
  assign y23961 = ~1'b0 ;
  assign y23962 = ~n32385 ;
  assign y23963 = ~n536 ;
  assign y23964 = ~n32387 ;
  assign y23965 = ~1'b0 ;
  assign y23966 = n32391 ;
  assign y23967 = ~1'b0 ;
  assign y23968 = ~1'b0 ;
  assign y23969 = ~1'b0 ;
  assign y23970 = ~1'b0 ;
  assign y23971 = ~1'b0 ;
  assign y23972 = n32393 ;
  assign y23973 = ~n32396 ;
  assign y23974 = ~n32401 ;
  assign y23975 = 1'b0 ;
  assign y23976 = 1'b0 ;
  assign y23977 = n32402 ;
  assign y23978 = ~1'b0 ;
  assign y23979 = ~n32403 ;
  assign y23980 = ~1'b0 ;
  assign y23981 = ~n32407 ;
  assign y23982 = ~n17668 ;
  assign y23983 = ~1'b0 ;
  assign y23984 = ~1'b0 ;
  assign y23985 = n32413 ;
  assign y23986 = 1'b0 ;
  assign y23987 = n32414 ;
  assign y23988 = ~1'b0 ;
  assign y23989 = ~1'b0 ;
  assign y23990 = ~n32418 ;
  assign y23991 = n32419 ;
  assign y23992 = ~n15549 ;
  assign y23993 = ~1'b0 ;
  assign y23994 = ~1'b0 ;
  assign y23995 = ~1'b0 ;
  assign y23996 = n32422 ;
  assign y23997 = ~n32423 ;
  assign y23998 = 1'b0 ;
  assign y23999 = ~1'b0 ;
  assign y24000 = 1'b0 ;
  assign y24001 = ~1'b0 ;
  assign y24002 = n32425 ;
  assign y24003 = n32428 ;
  assign y24004 = ~1'b0 ;
  assign y24005 = ~n32431 ;
  assign y24006 = n32432 ;
  assign y24007 = ~n32433 ;
  assign y24008 = ~1'b0 ;
  assign y24009 = n32437 ;
  assign y24010 = ~n32439 ;
  assign y24011 = ~n128 ;
  assign y24012 = ~n32441 ;
  assign y24013 = n32444 ;
  assign y24014 = ~1'b0 ;
  assign y24015 = n32445 ;
  assign y24016 = n32448 ;
  assign y24017 = n32449 ;
  assign y24018 = n32453 ;
  assign y24019 = n32455 ;
  assign y24020 = ~1'b0 ;
  assign y24021 = n32136 ;
  assign y24022 = ~n32459 ;
  assign y24023 = n32461 ;
  assign y24024 = n32466 ;
  assign y24025 = ~1'b0 ;
  assign y24026 = 1'b0 ;
  assign y24027 = n32468 ;
  assign y24028 = ~n32469 ;
  assign y24029 = ~n32473 ;
  assign y24030 = ~n25962 ;
  assign y24031 = n32474 ;
  assign y24032 = ~1'b0 ;
  assign y24033 = ~1'b0 ;
  assign y24034 = n32476 ;
  assign y24035 = ~1'b0 ;
  assign y24036 = n32479 ;
  assign y24037 = ~n32480 ;
  assign y24038 = ~1'b0 ;
  assign y24039 = ~n22877 ;
  assign y24040 = ~1'b0 ;
  assign y24041 = ~n32484 ;
  assign y24042 = n23764 ;
  assign y24043 = n32485 ;
  assign y24044 = n32488 ;
  assign y24045 = ~n32489 ;
  assign y24046 = ~n32495 ;
  assign y24047 = n26398 ;
  assign y24048 = ~1'b0 ;
  assign y24049 = ~n4422 ;
  assign y24050 = ~1'b0 ;
  assign y24051 = ~n32500 ;
  assign y24052 = ~1'b0 ;
  assign y24053 = n32503 ;
  assign y24054 = ~n32506 ;
  assign y24055 = ~1'b0 ;
  assign y24056 = ~1'b0 ;
  assign y24057 = ~n32507 ;
  assign y24058 = ~1'b0 ;
  assign y24059 = ~n32508 ;
  assign y24060 = n32510 ;
  assign y24061 = ~1'b0 ;
  assign y24062 = n32511 ;
  assign y24063 = ~1'b0 ;
  assign y24064 = ~n32516 ;
  assign y24065 = ~n32517 ;
  assign y24066 = n13051 ;
  assign y24067 = ~n32519 ;
  assign y24068 = ~1'b0 ;
  assign y24069 = n32522 ;
  assign y24070 = 1'b0 ;
  assign y24071 = ~n24013 ;
  assign y24072 = n32523 ;
  assign y24073 = n32525 ;
  assign y24074 = ~1'b0 ;
  assign y24075 = n32527 ;
  assign y24076 = n32528 ;
  assign y24077 = 1'b0 ;
  assign y24078 = n32529 ;
  assign y24079 = ~1'b0 ;
  assign y24080 = ~1'b0 ;
  assign y24081 = n32530 ;
  assign y24082 = ~n32534 ;
  assign y24083 = n32536 ;
  assign y24084 = ~1'b0 ;
  assign y24085 = ~n32537 ;
  assign y24086 = ~n32538 ;
  assign y24087 = ~1'b0 ;
  assign y24088 = n32542 ;
  assign y24089 = ~n32546 ;
  assign y24090 = n32548 ;
  assign y24091 = ~n32550 ;
  assign y24092 = ~n32553 ;
  assign y24093 = ~1'b0 ;
  assign y24094 = ~n32555 ;
  assign y24095 = ~1'b0 ;
  assign y24096 = ~1'b0 ;
  assign y24097 = ~n32557 ;
  assign y24098 = n32559 ;
  assign y24099 = ~1'b0 ;
  assign y24100 = ~1'b0 ;
  assign y24101 = n32562 ;
  assign y24102 = ~n32564 ;
  assign y24103 = ~1'b0 ;
  assign y24104 = n32566 ;
  assign y24105 = n32568 ;
  assign y24106 = 1'b0 ;
  assign y24107 = ~n32570 ;
  assign y24108 = ~n32573 ;
  assign y24109 = ~n32575 ;
  assign y24110 = ~n32577 ;
  assign y24111 = ~1'b0 ;
  assign y24112 = 1'b0 ;
  assign y24113 = ~n32580 ;
  assign y24114 = ~n32581 ;
  assign y24115 = ~n32582 ;
  assign y24116 = ~1'b0 ;
  assign y24117 = n18156 ;
  assign y24118 = n32583 ;
  assign y24119 = n32584 ;
  assign y24120 = ~1'b0 ;
  assign y24121 = ~n32585 ;
  assign y24122 = ~1'b0 ;
  assign y24123 = ~1'b0 ;
  assign y24124 = ~n32590 ;
  assign y24125 = ~n32591 ;
  assign y24126 = ~n32592 ;
  assign y24127 = ~1'b0 ;
  assign y24128 = ~n32594 ;
  assign y24129 = 1'b0 ;
  assign y24130 = ~1'b0 ;
  assign y24131 = ~n32595 ;
  assign y24132 = n32597 ;
  assign y24133 = n18352 ;
  assign y24134 = ~1'b0 ;
  assign y24135 = ~n32598 ;
  assign y24136 = n32599 ;
  assign y24137 = n32604 ;
  assign y24138 = n32606 ;
  assign y24139 = ~n21822 ;
  assign y24140 = n32608 ;
  assign y24141 = ~1'b0 ;
  assign y24142 = n32609 ;
  assign y24143 = ~1'b0 ;
  assign y24144 = ~n32610 ;
  assign y24145 = ~1'b0 ;
  assign y24146 = ~1'b0 ;
  assign y24147 = n32612 ;
  assign y24148 = ~1'b0 ;
  assign y24149 = n32613 ;
  assign y24150 = ~1'b0 ;
  assign y24151 = ~n32615 ;
  assign y24152 = ~1'b0 ;
  assign y24153 = ~1'b0 ;
  assign y24154 = n32618 ;
  assign y24155 = ~1'b0 ;
  assign y24156 = ~1'b0 ;
  assign y24157 = ~1'b0 ;
  assign y24158 = ~1'b0 ;
  assign y24159 = n4862 ;
  assign y24160 = n32619 ;
  assign y24161 = ~n899 ;
  assign y24162 = n32621 ;
  assign y24163 = n32624 ;
  assign y24164 = n8161 ;
  assign y24165 = ~1'b0 ;
  assign y24166 = ~n32634 ;
  assign y24167 = n32637 ;
  assign y24168 = n32639 ;
  assign y24169 = ~n32640 ;
  assign y24170 = ~n32641 ;
  assign y24171 = ~1'b0 ;
  assign y24172 = ~n32642 ;
  assign y24173 = n32643 ;
  assign y24174 = ~1'b0 ;
  assign y24175 = ~n7794 ;
  assign y24176 = ~n32646 ;
  assign y24177 = n32648 ;
  assign y24178 = n32651 ;
  assign y24179 = 1'b0 ;
  assign y24180 = ~1'b0 ;
  assign y24181 = ~1'b0 ;
  assign y24182 = ~n32653 ;
  assign y24183 = 1'b0 ;
  assign y24184 = ~1'b0 ;
  assign y24185 = ~n32660 ;
  assign y24186 = ~1'b0 ;
  assign y24187 = ~n32662 ;
  assign y24188 = n6476 ;
  assign y24189 = ~n32663 ;
  assign y24190 = ~1'b0 ;
  assign y24191 = n24909 ;
  assign y24192 = n3394 ;
  assign y24193 = n32665 ;
  assign y24194 = ~1'b0 ;
  assign y24195 = n32669 ;
  assign y24196 = ~n32673 ;
  assign y24197 = ~1'b0 ;
  assign y24198 = ~1'b0 ;
  assign y24199 = ~1'b0 ;
  assign y24200 = n32676 ;
  assign y24201 = n25407 ;
  assign y24202 = n32678 ;
  assign y24203 = ~n32679 ;
  assign y24204 = ~n32682 ;
  assign y24205 = ~1'b0 ;
  assign y24206 = ~1'b0 ;
  assign y24207 = n13278 ;
  assign y24208 = n17572 ;
  assign y24209 = ~n32683 ;
  assign y24210 = ~n32684 ;
  assign y24211 = ~n32685 ;
  assign y24212 = n32687 ;
  assign y24213 = ~n32688 ;
  assign y24214 = ~n32689 ;
  assign y24215 = ~n32690 ;
  assign y24216 = ~1'b0 ;
  assign y24217 = n32692 ;
  assign y24218 = ~n32694 ;
  assign y24219 = n32695 ;
  assign y24220 = n32697 ;
  assign y24221 = ~1'b0 ;
  assign y24222 = ~n32699 ;
  assign y24223 = 1'b0 ;
  assign y24224 = ~n32703 ;
  assign y24225 = ~1'b0 ;
  assign y24226 = n32704 ;
  assign y24227 = ~n32707 ;
  assign y24228 = ~n32708 ;
  assign y24229 = 1'b0 ;
  assign y24230 = ~1'b0 ;
  assign y24231 = ~1'b0 ;
  assign y24232 = n32711 ;
  assign y24233 = ~n32713 ;
  assign y24234 = ~n5046 ;
  assign y24235 = ~1'b0 ;
  assign y24236 = ~1'b0 ;
  assign y24237 = n32714 ;
  assign y24238 = n32715 ;
  assign y24239 = n32716 ;
  assign y24240 = 1'b0 ;
  assign y24241 = ~1'b0 ;
  assign y24242 = ~n11258 ;
  assign y24243 = ~n758 ;
  assign y24244 = ~1'b0 ;
  assign y24245 = n32717 ;
  assign y24246 = ~n32720 ;
  assign y24247 = ~n32723 ;
  assign y24248 = ~n32724 ;
  assign y24249 = ~n32725 ;
  assign y24250 = ~1'b0 ;
  assign y24251 = n25625 ;
  assign y24252 = n32726 ;
  assign y24253 = ~1'b0 ;
  assign y24254 = ~n32728 ;
  assign y24255 = ~n32731 ;
  assign y24256 = ~n32733 ;
  assign y24257 = ~n32736 ;
  assign y24258 = n32758 ;
  assign y24259 = n32759 ;
  assign y24260 = ~1'b0 ;
  assign y24261 = ~n32761 ;
  assign y24262 = ~1'b0 ;
  assign y24263 = n32763 ;
  assign y24264 = ~1'b0 ;
  assign y24265 = n16423 ;
  assign y24266 = n32767 ;
  assign y24267 = ~n32768 ;
  assign y24268 = ~1'b0 ;
  assign y24269 = n32769 ;
  assign y24270 = ~n32772 ;
  assign y24271 = 1'b0 ;
  assign y24272 = n32774 ;
  assign y24273 = ~n32776 ;
  assign y24274 = n32780 ;
  assign y24275 = n32782 ;
  assign y24276 = ~1'b0 ;
  assign y24277 = 1'b0 ;
  assign y24278 = n32783 ;
  assign y24279 = ~n6714 ;
  assign y24280 = ~n32784 ;
  assign y24281 = ~1'b0 ;
  assign y24282 = n21424 ;
  assign y24283 = ~n32786 ;
  assign y24284 = n32787 ;
  assign y24285 = ~n9480 ;
  assign y24286 = ~n32790 ;
  assign y24287 = ~n32792 ;
  assign y24288 = ~n32795 ;
  assign y24289 = ~n32799 ;
  assign y24290 = ~1'b0 ;
  assign y24291 = ~n32800 ;
  assign y24292 = ~n32801 ;
  assign y24293 = ~1'b0 ;
  assign y24294 = ~n32804 ;
  assign y24295 = n32806 ;
  assign y24296 = ~1'b0 ;
  assign y24297 = n32808 ;
  assign y24298 = ~1'b0 ;
  assign y24299 = n32813 ;
  assign y24300 = n32815 ;
  assign y24301 = ~1'b0 ;
  assign y24302 = ~1'b0 ;
  assign y24303 = n32819 ;
  assign y24304 = ~n32821 ;
  assign y24305 = ~n32822 ;
  assign y24306 = n9012 ;
  assign y24307 = ~n32823 ;
  assign y24308 = n32824 ;
  assign y24309 = ~n32825 ;
  assign y24310 = ~n32827 ;
  assign y24311 = ~1'b0 ;
  assign y24312 = ~1'b0 ;
  assign y24313 = ~1'b0 ;
  assign y24314 = ~n32828 ;
  assign y24315 = n32830 ;
  assign y24316 = ~n32831 ;
  assign y24317 = ~1'b0 ;
  assign y24318 = n32833 ;
  assign y24319 = ~n32839 ;
  assign y24320 = ~n32840 ;
  assign y24321 = ~1'b0 ;
  assign y24322 = n257 ;
  assign y24323 = n32841 ;
  assign y24324 = ~n32843 ;
  assign y24325 = n30520 ;
  assign y24326 = ~n32846 ;
  assign y24327 = ~1'b0 ;
  assign y24328 = ~1'b0 ;
  assign y24329 = n2107 ;
  assign y24330 = n23589 ;
  assign y24331 = ~1'b0 ;
  assign y24332 = ~1'b0 ;
  assign y24333 = ~n32849 ;
  assign y24334 = n32850 ;
  assign y24335 = ~n32853 ;
  assign y24336 = n32854 ;
  assign y24337 = n12473 ;
  assign y24338 = ~1'b0 ;
  assign y24339 = n1072 ;
  assign y24340 = ~1'b0 ;
  assign y24341 = n32855 ;
  assign y24342 = ~n32857 ;
  assign y24343 = ~1'b0 ;
  assign y24344 = n32859 ;
  assign y24345 = ~n32860 ;
  assign y24346 = ~n32861 ;
  assign y24347 = n32864 ;
  assign y24348 = ~1'b0 ;
  assign y24349 = ~1'b0 ;
  assign y24350 = ~1'b0 ;
  assign y24351 = ~1'b0 ;
  assign y24352 = ~1'b0 ;
  assign y24353 = n32867 ;
  assign y24354 = ~n32868 ;
  assign y24355 = n32870 ;
  assign y24356 = ~1'b0 ;
  assign y24357 = ~n32872 ;
  assign y24358 = ~n32874 ;
  assign y24359 = ~1'b0 ;
  assign y24360 = n32876 ;
  assign y24361 = ~1'b0 ;
  assign y24362 = n32877 ;
  assign y24363 = ~n32878 ;
  assign y24364 = ~1'b0 ;
  assign y24365 = ~1'b0 ;
  assign y24366 = ~1'b0 ;
  assign y24367 = ~n32879 ;
  assign y24368 = ~1'b0 ;
  assign y24369 = ~n32883 ;
  assign y24370 = ~n32885 ;
  assign y24371 = n32886 ;
  assign y24372 = n32887 ;
  assign y24373 = ~n32889 ;
  assign y24374 = n32890 ;
  assign y24375 = ~1'b0 ;
  assign y24376 = n32892 ;
  assign y24377 = ~1'b0 ;
  assign y24378 = ~n32893 ;
  assign y24379 = ~n32895 ;
  assign y24380 = ~n32899 ;
  assign y24381 = ~1'b0 ;
  assign y24382 = n32900 ;
  assign y24383 = ~n32903 ;
  assign y24384 = ~1'b0 ;
  assign y24385 = n32905 ;
  assign y24386 = n32906 ;
  assign y24387 = n32908 ;
  assign y24388 = ~n7688 ;
  assign y24389 = n32909 ;
  assign y24390 = ~n32910 ;
  assign y24391 = ~n32918 ;
  assign y24392 = 1'b0 ;
  assign y24393 = n32920 ;
  assign y24394 = ~1'b0 ;
  assign y24395 = ~n32921 ;
  assign y24396 = ~1'b0 ;
  assign y24397 = n32923 ;
  assign y24398 = ~n32925 ;
  assign y24399 = ~n32929 ;
  assign y24400 = n28015 ;
  assign y24401 = n32930 ;
  assign y24402 = ~1'b0 ;
  assign y24403 = ~n32933 ;
  assign y24404 = n12487 ;
  assign y24405 = ~1'b0 ;
  assign y24406 = ~n32934 ;
  assign y24407 = ~1'b0 ;
  assign y24408 = ~1'b0 ;
  assign y24409 = n32936 ;
  assign y24410 = ~n3299 ;
  assign y24411 = ~1'b0 ;
  assign y24412 = ~1'b0 ;
  assign y24413 = ~1'b0 ;
  assign y24414 = ~n859 ;
  assign y24415 = ~1'b0 ;
  assign y24416 = ~1'b0 ;
  assign y24417 = ~1'b0 ;
  assign y24418 = ~n32938 ;
  assign y24419 = n32939 ;
  assign y24420 = ~n2526 ;
  assign y24421 = n14326 ;
  assign y24422 = ~n8192 ;
  assign y24423 = ~1'b0 ;
  assign y24424 = n32941 ;
  assign y24425 = n32942 ;
  assign y24426 = ~1'b0 ;
  assign y24427 = n26905 ;
  assign y24428 = n32944 ;
  assign y24429 = n1169 ;
  assign y24430 = ~1'b0 ;
  assign y24431 = n32947 ;
  assign y24432 = n32951 ;
  assign y24433 = ~1'b0 ;
  assign y24434 = n32952 ;
  assign y24435 = ~1'b0 ;
  assign y24436 = ~1'b0 ;
  assign y24437 = ~1'b0 ;
  assign y24438 = ~1'b0 ;
  assign y24439 = ~n16440 ;
  assign y24440 = n10641 ;
  assign y24441 = ~n32953 ;
  assign y24442 = ~1'b0 ;
  assign y24443 = ~1'b0 ;
  assign y24444 = ~n2212 ;
  assign y24445 = n32955 ;
  assign y24446 = ~1'b0 ;
  assign y24447 = n32956 ;
  assign y24448 = ~1'b0 ;
  assign y24449 = n32958 ;
  assign y24450 = ~n25878 ;
  assign y24451 = ~1'b0 ;
  assign y24452 = n32616 ;
  assign y24453 = ~n32960 ;
  assign y24454 = ~n19158 ;
  assign y24455 = n32961 ;
  assign y24456 = n32962 ;
  assign y24457 = 1'b0 ;
  assign y24458 = ~n32963 ;
  assign y24459 = ~1'b0 ;
  assign y24460 = n852 ;
  assign y24461 = ~n32967 ;
  assign y24462 = ~1'b0 ;
  assign y24463 = ~1'b0 ;
  assign y24464 = ~n32968 ;
  assign y24465 = n32969 ;
  assign y24466 = ~n32971 ;
  assign y24467 = ~1'b0 ;
  assign y24468 = ~n32972 ;
  assign y24469 = ~n116 ;
  assign y24470 = ~n32973 ;
  assign y24471 = ~1'b0 ;
  assign y24472 = ~n32974 ;
  assign y24473 = n32975 ;
  assign y24474 = n32978 ;
  assign y24475 = ~1'b0 ;
  assign y24476 = n32979 ;
  assign y24477 = ~1'b0 ;
  assign y24478 = ~n32982 ;
  assign y24479 = n32984 ;
  assign y24480 = ~n32985 ;
  assign y24481 = ~1'b0 ;
  assign y24482 = n31943 ;
  assign y24483 = ~1'b0 ;
  assign y24484 = n32988 ;
  assign y24485 = n32991 ;
  assign y24486 = 1'b0 ;
  assign y24487 = n32997 ;
  assign y24488 = ~n32998 ;
  assign y24489 = ~1'b0 ;
  assign y24490 = ~n32999 ;
  assign y24491 = ~n8071 ;
  assign y24492 = n33001 ;
  assign y24493 = ~1'b0 ;
  assign y24494 = n6040 ;
  assign y24495 = n33002 ;
  assign y24496 = ~n33004 ;
  assign y24497 = 1'b0 ;
  assign y24498 = 1'b0 ;
  assign y24499 = ~1'b0 ;
  assign y24500 = ~1'b0 ;
  assign y24501 = n33006 ;
  assign y24502 = n33007 ;
  assign y24503 = n33008 ;
  assign y24504 = n33010 ;
  assign y24505 = n33011 ;
  assign y24506 = ~1'b0 ;
  assign y24507 = ~1'b0 ;
  assign y24508 = ~1'b0 ;
  assign y24509 = ~1'b0 ;
  assign y24510 = n33012 ;
  assign y24511 = ~n33016 ;
  assign y24512 = ~1'b0 ;
  assign y24513 = ~1'b0 ;
  assign y24514 = ~1'b0 ;
  assign y24515 = ~n33017 ;
  assign y24516 = n33020 ;
  assign y24517 = ~n33022 ;
  assign y24518 = n33023 ;
  assign y24519 = ~1'b0 ;
  assign y24520 = n2014 ;
  assign y24521 = ~1'b0 ;
  assign y24522 = ~1'b0 ;
  assign y24523 = ~1'b0 ;
  assign y24524 = ~n33025 ;
  assign y24525 = ~n33026 ;
  assign y24526 = ~1'b0 ;
  assign y24527 = n33027 ;
  assign y24528 = n33032 ;
  assign y24529 = ~n33033 ;
  assign y24530 = n29530 ;
  assign y24531 = ~1'b0 ;
  assign y24532 = ~n33036 ;
  assign y24533 = n33038 ;
  assign y24534 = ~1'b0 ;
  assign y24535 = n13594 ;
  assign y24536 = ~n33039 ;
  assign y24537 = n2817 ;
  assign y24538 = ~1'b0 ;
  assign y24539 = ~n18200 ;
  assign y24540 = n9524 ;
  assign y24541 = ~1'b0 ;
  assign y24542 = 1'b0 ;
  assign y24543 = n33040 ;
  assign y24544 = ~n33041 ;
  assign y24545 = n33042 ;
  assign y24546 = ~1'b0 ;
  assign y24547 = n33045 ;
  assign y24548 = ~1'b0 ;
  assign y24549 = ~1'b0 ;
  assign y24550 = ~n33046 ;
  assign y24551 = 1'b0 ;
  assign y24552 = n33047 ;
  assign y24553 = n28490 ;
  assign y24554 = ~n33050 ;
  assign y24555 = n33052 ;
  assign y24556 = ~1'b0 ;
  assign y24557 = ~1'b0 ;
  assign y24558 = ~n33055 ;
  assign y24559 = ~n33058 ;
  assign y24560 = ~1'b0 ;
  assign y24561 = n33063 ;
  assign y24562 = 1'b0 ;
  assign y24563 = ~n33066 ;
  assign y24564 = ~1'b0 ;
  assign y24565 = ~n33067 ;
  assign y24566 = n33070 ;
  assign y24567 = ~1'b0 ;
  assign y24568 = ~1'b0 ;
  assign y24569 = ~n33071 ;
  assign y24570 = ~1'b0 ;
  assign y24571 = ~1'b0 ;
  assign y24572 = ~n33072 ;
  assign y24573 = n17891 ;
  assign y24574 = n33073 ;
  assign y24575 = ~n33074 ;
  assign y24576 = ~1'b0 ;
  assign y24577 = ~1'b0 ;
  assign y24578 = ~1'b0 ;
  assign y24579 = ~n33075 ;
  assign y24580 = n33080 ;
  assign y24581 = ~1'b0 ;
  assign y24582 = n33090 ;
  assign y24583 = n33092 ;
  assign y24584 = ~n33096 ;
  assign y24585 = ~1'b0 ;
  assign y24586 = ~n33100 ;
  assign y24587 = ~1'b0 ;
  assign y24588 = ~1'b0 ;
  assign y24589 = ~n33101 ;
  assign y24590 = n33103 ;
  assign y24591 = ~n33105 ;
  assign y24592 = ~1'b0 ;
  assign y24593 = n33107 ;
  assign y24594 = ~n33108 ;
  assign y24595 = ~n33109 ;
  assign y24596 = ~n33110 ;
  assign y24597 = ~n33113 ;
  assign y24598 = n7110 ;
  assign y24599 = ~1'b0 ;
  assign y24600 = 1'b0 ;
  assign y24601 = ~1'b0 ;
  assign y24602 = 1'b0 ;
  assign y24603 = ~n820 ;
  assign y24604 = ~n33114 ;
  assign y24605 = ~1'b0 ;
  assign y24606 = ~1'b0 ;
  assign y24607 = ~n2370 ;
  assign y24608 = ~1'b0 ;
  assign y24609 = ~1'b0 ;
  assign y24610 = ~1'b0 ;
  assign y24611 = n33117 ;
  assign y24612 = ~1'b0 ;
  assign y24613 = n33120 ;
  assign y24614 = ~1'b0 ;
  assign y24615 = ~n33132 ;
  assign y24616 = ~n33136 ;
  assign y24617 = n33138 ;
  assign y24618 = ~n33139 ;
  assign y24619 = ~n33144 ;
  assign y24620 = 1'b0 ;
  assign y24621 = n11931 ;
  assign y24622 = n33145 ;
  assign y24623 = n13903 ;
  assign y24624 = ~1'b0 ;
  assign y24625 = n33146 ;
  assign y24626 = ~1'b0 ;
  assign y24627 = n33151 ;
  assign y24628 = ~1'b0 ;
  assign y24629 = n33153 ;
  assign y24630 = ~1'b0 ;
  assign y24631 = ~n33156 ;
  assign y24632 = n1139 ;
  assign y24633 = ~1'b0 ;
  assign y24634 = ~1'b0 ;
  assign y24635 = ~n33157 ;
  assign y24636 = ~1'b0 ;
  assign y24637 = ~1'b0 ;
  assign y24638 = ~1'b0 ;
  assign y24639 = ~n33159 ;
  assign y24640 = n33160 ;
  assign y24641 = ~1'b0 ;
  assign y24642 = 1'b0 ;
  assign y24643 = ~n33163 ;
  assign y24644 = ~n33166 ;
  assign y24645 = ~n33177 ;
  assign y24646 = ~1'b0 ;
  assign y24647 = n33178 ;
  assign y24648 = ~1'b0 ;
  assign y24649 = ~n11758 ;
  assign y24650 = ~1'b0 ;
  assign y24651 = ~1'b0 ;
  assign y24652 = ~1'b0 ;
  assign y24653 = 1'b0 ;
  assign y24654 = 1'b0 ;
  assign y24655 = n33180 ;
  assign y24656 = ~1'b0 ;
  assign y24657 = ~n33181 ;
  assign y24658 = ~1'b0 ;
  assign y24659 = ~1'b0 ;
  assign y24660 = ~n33183 ;
  assign y24661 = ~n33187 ;
  assign y24662 = ~n33191 ;
  assign y24663 = ~n33192 ;
  assign y24664 = 1'b0 ;
  assign y24665 = n31537 ;
  assign y24666 = ~1'b0 ;
  assign y24667 = ~1'b0 ;
  assign y24668 = n33194 ;
  assign y24669 = ~1'b0 ;
  assign y24670 = ~1'b0 ;
  assign y24671 = ~n33196 ;
  assign y24672 = ~1'b0 ;
  assign y24673 = ~1'b0 ;
  assign y24674 = ~n33199 ;
  assign y24675 = ~1'b0 ;
  assign y24676 = ~1'b0 ;
  assign y24677 = n33204 ;
  assign y24678 = ~n33208 ;
  assign y24679 = 1'b0 ;
  assign y24680 = n33212 ;
  assign y24681 = ~1'b0 ;
  assign y24682 = ~n33216 ;
  assign y24683 = ~n33219 ;
  assign y24684 = ~n33221 ;
  assign y24685 = ~n33222 ;
  assign y24686 = ~n33223 ;
  assign y24687 = n33225 ;
  assign y24688 = ~n33226 ;
  assign y24689 = ~n170 ;
  assign y24690 = 1'b0 ;
  assign y24691 = ~1'b0 ;
  assign y24692 = ~1'b0 ;
  assign y24693 = ~n33227 ;
  assign y24694 = ~n33229 ;
  assign y24695 = n24241 ;
  assign y24696 = ~1'b0 ;
  assign y24697 = ~1'b0 ;
  assign y24698 = ~n5360 ;
  assign y24699 = ~1'b0 ;
  assign y24700 = ~n33231 ;
  assign y24701 = n1622 ;
  assign y24702 = ~n33232 ;
  assign y24703 = ~1'b0 ;
  assign y24704 = n33235 ;
  assign y24705 = n33236 ;
  assign y24706 = n23764 ;
  assign y24707 = n33237 ;
  assign y24708 = ~1'b0 ;
  assign y24709 = ~n21330 ;
  assign y24710 = ~1'b0 ;
  assign y24711 = ~n33240 ;
  assign y24712 = ~n33241 ;
  assign y24713 = ~1'b0 ;
  assign y24714 = ~1'b0 ;
  assign y24715 = ~n33244 ;
  assign y24716 = ~1'b0 ;
  assign y24717 = n33248 ;
  assign y24718 = ~1'b0 ;
  assign y24719 = ~1'b0 ;
  assign y24720 = n33251 ;
  assign y24721 = ~1'b0 ;
  assign y24722 = 1'b0 ;
  assign y24723 = n33252 ;
  assign y24724 = n33258 ;
  assign y24725 = n33263 ;
  assign y24726 = ~n33265 ;
  assign y24727 = ~1'b0 ;
  assign y24728 = ~n33267 ;
  assign y24729 = ~1'b0 ;
  assign y24730 = n33271 ;
  assign y24731 = ~n1152 ;
  assign y24732 = n33272 ;
  assign y24733 = n33275 ;
  assign y24734 = 1'b0 ;
  assign y24735 = ~1'b0 ;
  assign y24736 = ~1'b0 ;
  assign y24737 = ~n33281 ;
  assign y24738 = ~n33282 ;
  assign y24739 = ~1'b0 ;
  assign y24740 = ~n33285 ;
  assign y24741 = ~1'b0 ;
  assign y24742 = n33289 ;
  assign y24743 = ~1'b0 ;
  assign y24744 = ~n33291 ;
  assign y24745 = ~n33292 ;
  assign y24746 = ~1'b0 ;
  assign y24747 = n33293 ;
  assign y24748 = ~n33297 ;
  assign y24749 = n33300 ;
  assign y24750 = ~1'b0 ;
  assign y24751 = ~1'b0 ;
  assign y24752 = ~1'b0 ;
  assign y24753 = ~1'b0 ;
  assign y24754 = ~n33301 ;
  assign y24755 = ~1'b0 ;
  assign y24756 = ~n33303 ;
  assign y24757 = n33304 ;
  assign y24758 = ~1'b0 ;
  assign y24759 = n33305 ;
  assign y24760 = ~1'b0 ;
  assign y24761 = n12736 ;
  assign y24762 = ~n33309 ;
  assign y24763 = n3907 ;
  assign y24764 = ~n33311 ;
  assign y24765 = ~1'b0 ;
  assign y24766 = ~n33315 ;
  assign y24767 = ~n2754 ;
  assign y24768 = ~1'b0 ;
  assign y24769 = n3188 ;
  assign y24770 = ~n33316 ;
  assign y24771 = ~1'b0 ;
  assign y24772 = ~1'b0 ;
  assign y24773 = n33317 ;
  assign y24774 = ~n33318 ;
  assign y24775 = ~n33319 ;
  assign y24776 = 1'b0 ;
  assign y24777 = ~n33325 ;
  assign y24778 = ~1'b0 ;
  assign y24779 = ~n33326 ;
  assign y24780 = ~1'b0 ;
  assign y24781 = ~1'b0 ;
  assign y24782 = n33332 ;
  assign y24783 = ~n33334 ;
  assign y24784 = ~n33336 ;
  assign y24785 = ~n33337 ;
  assign y24786 = ~1'b0 ;
  assign y24787 = n33340 ;
  assign y24788 = ~n33345 ;
  assign y24789 = ~1'b0 ;
  assign y24790 = ~1'b0 ;
  assign y24791 = ~1'b0 ;
  assign y24792 = ~n33349 ;
  assign y24793 = ~n33350 ;
  assign y24794 = ~1'b0 ;
  assign y24795 = n33351 ;
  assign y24796 = ~n33353 ;
  assign y24797 = ~n17104 ;
  assign y24798 = n33355 ;
  assign y24799 = n33356 ;
  assign y24800 = ~1'b0 ;
  assign y24801 = ~1'b0 ;
  assign y24802 = ~n33357 ;
  assign y24803 = n33360 ;
  assign y24804 = n33361 ;
  assign y24805 = n33362 ;
  assign y24806 = n16313 ;
  assign y24807 = n33364 ;
  assign y24808 = ~1'b0 ;
  assign y24809 = n33366 ;
  assign y24810 = n33368 ;
  assign y24811 = n33369 ;
  assign y24812 = ~n33376 ;
  assign y24813 = ~n19770 ;
  assign y24814 = ~1'b0 ;
  assign y24815 = ~n33377 ;
  assign y24816 = ~n33379 ;
  assign y24817 = ~n18921 ;
  assign y24818 = 1'b0 ;
  assign y24819 = n33380 ;
  assign y24820 = ~n33382 ;
  assign y24821 = n33383 ;
  assign y24822 = n33384 ;
  assign y24823 = ~1'b0 ;
  assign y24824 = ~n33388 ;
  assign y24825 = ~n813 ;
  assign y24826 = ~n33390 ;
  assign y24827 = ~1'b0 ;
  assign y24828 = n3078 ;
  assign y24829 = ~1'b0 ;
  assign y24830 = n33391 ;
  assign y24831 = n33392 ;
  assign y24832 = ~n1790 ;
  assign y24833 = n33393 ;
  assign y24834 = 1'b0 ;
  assign y24835 = ~1'b0 ;
  assign y24836 = ~1'b0 ;
  assign y24837 = 1'b0 ;
  assign y24838 = n33395 ;
  assign y24839 = 1'b0 ;
  assign y24840 = ~1'b0 ;
  assign y24841 = n33398 ;
  assign y24842 = n29843 ;
  assign y24843 = ~n33401 ;
  assign y24844 = ~n33402 ;
  assign y24845 = n33404 ;
  assign y24846 = n33407 ;
  assign y24847 = n33411 ;
  assign y24848 = n33412 ;
  assign y24849 = n33414 ;
  assign y24850 = ~n33417 ;
  assign y24851 = ~n33419 ;
  assign y24852 = n33420 ;
  assign y24853 = ~1'b0 ;
  assign y24854 = ~n33421 ;
  assign y24855 = ~1'b0 ;
  assign y24856 = ~1'b0 ;
  assign y24857 = n33425 ;
  assign y24858 = ~n33426 ;
  assign y24859 = ~1'b0 ;
  assign y24860 = n33427 ;
  assign y24861 = ~n25074 ;
  assign y24862 = n33428 ;
  assign y24863 = ~1'b0 ;
  assign y24864 = 1'b0 ;
  assign y24865 = ~1'b0 ;
  assign y24866 = n1086 ;
  assign y24867 = n33430 ;
  assign y24868 = n33431 ;
  assign y24869 = ~n33433 ;
  assign y24870 = ~n33434 ;
  assign y24871 = n33435 ;
  assign y24872 = n4921 ;
  assign y24873 = ~1'b0 ;
  assign y24874 = n33436 ;
  assign y24875 = n33443 ;
  assign y24876 = ~n33447 ;
  assign y24877 = ~n33449 ;
  assign y24878 = ~n33452 ;
  assign y24879 = ~n33454 ;
  assign y24880 = ~n33455 ;
  assign y24881 = n33456 ;
  assign y24882 = ~n33457 ;
  assign y24883 = ~1'b0 ;
  assign y24884 = ~1'b0 ;
  assign y24885 = n33458 ;
  assign y24886 = ~1'b0 ;
  assign y24887 = n33460 ;
  assign y24888 = ~n33463 ;
  assign y24889 = ~n33468 ;
  assign y24890 = n25633 ;
  assign y24891 = ~1'b0 ;
  assign y24892 = ~1'b0 ;
  assign y24893 = ~n33469 ;
  assign y24894 = ~n20727 ;
  assign y24895 = n33470 ;
  assign y24896 = n33472 ;
  assign y24897 = ~n33473 ;
  assign y24898 = ~n33474 ;
  assign y24899 = n33476 ;
  assign y24900 = ~1'b0 ;
  assign y24901 = ~1'b0 ;
  assign y24902 = n33482 ;
  assign y24903 = ~1'b0 ;
  assign y24904 = ~1'b0 ;
  assign y24905 = ~1'b0 ;
  assign y24906 = ~n33485 ;
  assign y24907 = ~1'b0 ;
  assign y24908 = ~1'b0 ;
  assign y24909 = n33488 ;
  assign y24910 = ~1'b0 ;
  assign y24911 = ~n33490 ;
  assign y24912 = ~n24284 ;
  assign y24913 = n33492 ;
  assign y24914 = ~n14624 ;
  assign y24915 = ~n33493 ;
  assign y24916 = ~n33495 ;
  assign y24917 = ~n33501 ;
  assign y24918 = n33504 ;
  assign y24919 = ~1'b0 ;
  assign y24920 = ~1'b0 ;
  assign y24921 = ~1'b0 ;
  assign y24922 = ~1'b0 ;
  assign y24923 = n33505 ;
  assign y24924 = ~n33506 ;
  assign y24925 = ~n33509 ;
  assign y24926 = n33513 ;
  assign y24927 = n33514 ;
  assign y24928 = ~1'b0 ;
  assign y24929 = n33515 ;
  assign y24930 = ~1'b0 ;
  assign y24931 = ~1'b0 ;
  assign y24932 = n33517 ;
  assign y24933 = n33520 ;
  assign y24934 = ~n5726 ;
  assign y24935 = ~1'b0 ;
  assign y24936 = ~1'b0 ;
  assign y24937 = n33522 ;
  assign y24938 = n33523 ;
  assign y24939 = ~1'b0 ;
  assign y24940 = n30262 ;
  assign y24941 = ~n15923 ;
  assign y24942 = n33524 ;
  assign y24943 = ~n33526 ;
  assign y24944 = ~n9746 ;
  assign y24945 = ~n33529 ;
  assign y24946 = n33531 ;
  assign y24947 = ~1'b0 ;
  assign y24948 = n33534 ;
  assign y24949 = ~1'b0 ;
  assign y24950 = ~n33536 ;
  assign y24951 = n33538 ;
  assign y24952 = ~n33542 ;
  assign y24953 = ~n2233 ;
  assign y24954 = ~1'b0 ;
  assign y24955 = ~1'b0 ;
  assign y24956 = n33546 ;
  assign y24957 = ~n33547 ;
  assign y24958 = n11666 ;
  assign y24959 = ~n33549 ;
  assign y24960 = ~1'b0 ;
  assign y24961 = n33554 ;
  assign y24962 = ~n33557 ;
  assign y24963 = ~n33559 ;
  assign y24964 = n33561 ;
  assign y24965 = ~n33562 ;
  assign y24966 = ~n33565 ;
  assign y24967 = ~1'b0 ;
  assign y24968 = ~n33566 ;
  assign y24969 = ~1'b0 ;
  assign y24970 = ~n33569 ;
  assign y24971 = ~1'b0 ;
  assign y24972 = ~1'b0 ;
  assign y24973 = n33571 ;
  assign y24974 = ~n15904 ;
  assign y24975 = n33574 ;
  assign y24976 = ~n1054 ;
  assign y24977 = ~n33577 ;
  assign y24978 = ~1'b0 ;
  assign y24979 = ~1'b0 ;
  assign y24980 = n33578 ;
  assign y24981 = n33581 ;
  assign y24982 = ~n4482 ;
  assign y24983 = n33583 ;
  assign y24984 = n33586 ;
  assign y24985 = n510 ;
  assign y24986 = ~n33589 ;
  assign y24987 = ~1'b0 ;
  assign y24988 = ~n33590 ;
  assign y24989 = n33592 ;
  assign y24990 = ~n33593 ;
  assign y24991 = ~1'b0 ;
  assign y24992 = ~n33594 ;
  assign y24993 = n33595 ;
  assign y24994 = ~n33597 ;
  assign y24995 = n33602 ;
  assign y24996 = n33604 ;
  assign y24997 = ~1'b0 ;
  assign y24998 = ~1'b0 ;
  assign y24999 = ~n33605 ;
  assign y25000 = ~1'b0 ;
  assign y25001 = ~n33608 ;
  assign y25002 = ~1'b0 ;
  assign y25003 = n33611 ;
  assign y25004 = ~n33612 ;
  assign y25005 = ~n33619 ;
  assign y25006 = ~1'b0 ;
  assign y25007 = ~1'b0 ;
  assign y25008 = n33620 ;
  assign y25009 = n33623 ;
  assign y25010 = n33627 ;
  assign y25011 = ~n33631 ;
  assign y25012 = ~1'b0 ;
  assign y25013 = ~1'b0 ;
  assign y25014 = ~1'b0 ;
  assign y25015 = ~1'b0 ;
  assign y25016 = ~n33633 ;
  assign y25017 = n33634 ;
  assign y25018 = ~1'b0 ;
  assign y25019 = ~n33637 ;
  assign y25020 = ~n33639 ;
  assign y25021 = n24838 ;
  assign y25022 = ~n33642 ;
  assign y25023 = ~n26595 ;
  assign y25024 = ~1'b0 ;
  assign y25025 = ~1'b0 ;
  assign y25026 = n33644 ;
  assign y25027 = n33648 ;
  assign y25028 = ~1'b0 ;
  assign y25029 = ~1'b0 ;
  assign y25030 = ~n6579 ;
  assign y25031 = ~1'b0 ;
  assign y25032 = ~n323 ;
  assign y25033 = ~n33650 ;
  assign y25034 = n33651 ;
  assign y25035 = ~n33652 ;
  assign y25036 = ~n33653 ;
  assign y25037 = ~1'b0 ;
  assign y25038 = n33658 ;
  assign y25039 = n33660 ;
  assign y25040 = 1'b0 ;
  assign y25041 = n33662 ;
  assign y25042 = ~n33666 ;
  assign y25043 = ~1'b0 ;
  assign y25044 = ~n1960 ;
  assign y25045 = ~1'b0 ;
  assign y25046 = n9717 ;
  assign y25047 = ~n1705 ;
  assign y25048 = n33668 ;
  assign y25049 = ~n33674 ;
  assign y25050 = ~n33676 ;
  assign y25051 = n33677 ;
  assign y25052 = ~1'b0 ;
  assign y25053 = ~1'b0 ;
  assign y25054 = ~n33680 ;
  assign y25055 = ~1'b0 ;
  assign y25056 = 1'b0 ;
  assign y25057 = ~1'b0 ;
  assign y25058 = ~1'b0 ;
  assign y25059 = ~n33682 ;
  assign y25060 = ~1'b0 ;
  assign y25061 = ~1'b0 ;
  assign y25062 = n33697 ;
  assign y25063 = n33698 ;
  assign y25064 = ~1'b0 ;
  assign y25065 = 1'b0 ;
  assign y25066 = ~n6958 ;
  assign y25067 = ~1'b0 ;
  assign y25068 = 1'b0 ;
  assign y25069 = n12980 ;
  assign y25070 = n33702 ;
  assign y25071 = n33703 ;
  assign y25072 = ~1'b0 ;
  assign y25073 = ~n33706 ;
  assign y25074 = ~n33709 ;
  assign y25075 = n158 ;
  assign y25076 = n33711 ;
  assign y25077 = n33713 ;
  assign y25078 = ~1'b0 ;
  assign y25079 = ~1'b0 ;
  assign y25080 = ~1'b0 ;
  assign y25081 = ~n33718 ;
  assign y25082 = ~1'b0 ;
  assign y25083 = ~1'b0 ;
  assign y25084 = ~n33722 ;
  assign y25085 = ~n33723 ;
  assign y25086 = ~n33724 ;
  assign y25087 = ~1'b0 ;
  assign y25088 = ~n33725 ;
  assign y25089 = n24041 ;
  assign y25090 = ~1'b0 ;
  assign y25091 = n33729 ;
  assign y25092 = n33731 ;
  assign y25093 = ~n25230 ;
  assign y25094 = ~n33732 ;
  assign y25095 = ~1'b0 ;
  assign y25096 = ~n2141 ;
  assign y25097 = ~1'b0 ;
  assign y25098 = ~1'b0 ;
  assign y25099 = ~n33736 ;
  assign y25100 = n9910 ;
  assign y25101 = ~1'b0 ;
  assign y25102 = ~n33738 ;
  assign y25103 = ~n33739 ;
  assign y25104 = ~1'b0 ;
  assign y25105 = n33742 ;
  assign y25106 = ~1'b0 ;
  assign y25107 = n33745 ;
  assign y25108 = ~n33747 ;
  assign y25109 = ~n33748 ;
  assign y25110 = n33750 ;
  assign y25111 = ~1'b0 ;
  assign y25112 = ~n33751 ;
  assign y25113 = ~1'b0 ;
  assign y25114 = n33753 ;
  assign y25115 = ~n33759 ;
  assign y25116 = ~1'b0 ;
  assign y25117 = n33760 ;
  assign y25118 = ~n33773 ;
  assign y25119 = n33778 ;
  assign y25120 = 1'b0 ;
  assign y25121 = ~1'b0 ;
  assign y25122 = ~n33779 ;
  assign y25123 = n33780 ;
  assign y25124 = ~1'b0 ;
  assign y25125 = n33781 ;
  assign y25126 = n33783 ;
  assign y25127 = ~n33784 ;
  assign y25128 = ~n33786 ;
  assign y25129 = ~1'b0 ;
  assign y25130 = ~1'b0 ;
  assign y25131 = ~1'b0 ;
  assign y25132 = ~n33789 ;
  assign y25133 = n33793 ;
  assign y25134 = ~n7112 ;
  assign y25135 = n33794 ;
  assign y25136 = ~1'b0 ;
  assign y25137 = ~1'b0 ;
  assign y25138 = ~n33797 ;
  assign y25139 = ~n33802 ;
  assign y25140 = ~1'b0 ;
  assign y25141 = ~1'b0 ;
  assign y25142 = ~n33803 ;
  assign y25143 = n33807 ;
  assign y25144 = ~1'b0 ;
  assign y25145 = ~n31281 ;
  assign y25146 = ~1'b0 ;
  assign y25147 = ~1'b0 ;
  assign y25148 = ~n33809 ;
  assign y25149 = n33810 ;
  assign y25150 = ~1'b0 ;
  assign y25151 = n33811 ;
  assign y25152 = n1060 ;
  assign y25153 = n33812 ;
  assign y25154 = n33816 ;
  assign y25155 = n33818 ;
  assign y25156 = ~n33820 ;
  assign y25157 = ~n33821 ;
  assign y25158 = ~n33822 ;
  assign y25159 = n33830 ;
  assign y25160 = ~1'b0 ;
  assign y25161 = 1'b0 ;
  assign y25162 = n33834 ;
  assign y25163 = ~1'b0 ;
  assign y25164 = ~n257 ;
  assign y25165 = n33837 ;
  assign y25166 = ~n33839 ;
  assign y25167 = ~1'b0 ;
  assign y25168 = ~1'b0 ;
  assign y25169 = n5727 ;
  assign y25170 = ~1'b0 ;
  assign y25171 = n33840 ;
  assign y25172 = ~1'b0 ;
  assign y25173 = n2894 ;
  assign y25174 = ~n33841 ;
  assign y25175 = ~n33847 ;
  assign y25176 = 1'b0 ;
  assign y25177 = 1'b0 ;
  assign y25178 = 1'b0 ;
  assign y25179 = n33848 ;
  assign y25180 = n33849 ;
  assign y25181 = n33853 ;
  assign y25182 = n33854 ;
  assign y25183 = n33856 ;
  assign y25184 = ~1'b0 ;
  assign y25185 = ~n19628 ;
  assign y25186 = ~1'b0 ;
  assign y25187 = ~n33859 ;
  assign y25188 = ~n33860 ;
  assign y25189 = 1'b0 ;
  assign y25190 = n33861 ;
  assign y25191 = ~1'b0 ;
  assign y25192 = ~n8446 ;
  assign y25193 = ~1'b0 ;
  assign y25194 = ~n33863 ;
  assign y25195 = n33865 ;
  assign y25196 = ~n33868 ;
  assign y25197 = n33870 ;
  assign y25198 = 1'b0 ;
  assign y25199 = ~n33871 ;
  assign y25200 = n33872 ;
  assign y25201 = ~1'b0 ;
  assign y25202 = ~n33875 ;
  assign y25203 = 1'b0 ;
  assign y25204 = n33876 ;
  assign y25205 = ~n33877 ;
  assign y25206 = n33878 ;
  assign y25207 = ~1'b0 ;
  assign y25208 = n33882 ;
  assign y25209 = ~n33886 ;
  assign y25210 = ~n33889 ;
  assign y25211 = ~n28666 ;
  assign y25212 = ~n33892 ;
  assign y25213 = ~n33893 ;
  assign y25214 = ~n33895 ;
  assign y25215 = n33896 ;
  assign y25216 = ~1'b0 ;
  assign y25217 = ~n33902 ;
  assign y25218 = ~1'b0 ;
  assign y25219 = ~1'b0 ;
  assign y25220 = ~n33903 ;
  assign y25221 = n33904 ;
  assign y25222 = n33905 ;
  assign y25223 = n33906 ;
  assign y25224 = ~1'b0 ;
  assign y25225 = ~1'b0 ;
  assign y25226 = n33909 ;
  assign y25227 = n33913 ;
  assign y25228 = n33917 ;
  assign y25229 = n33918 ;
  assign y25230 = n33921 ;
  assign y25231 = n33926 ;
  assign y25232 = ~n33927 ;
  assign y25233 = ~1'b0 ;
  assign y25234 = ~1'b0 ;
  assign y25235 = n2109 ;
  assign y25236 = n33932 ;
  assign y25237 = ~n33933 ;
  assign y25238 = n33934 ;
  assign y25239 = ~n33936 ;
  assign y25240 = ~n33941 ;
  assign y25241 = ~1'b0 ;
  assign y25242 = n33942 ;
  assign y25243 = n33944 ;
  assign y25244 = ~n33945 ;
  assign y25245 = ~1'b0 ;
  assign y25246 = ~n33949 ;
  assign y25247 = ~1'b0 ;
  assign y25248 = ~n33953 ;
  assign y25249 = ~1'b0 ;
  assign y25250 = ~1'b0 ;
  assign y25251 = n33954 ;
  assign y25252 = ~1'b0 ;
  assign y25253 = ~1'b0 ;
  assign y25254 = n33956 ;
  assign y25255 = n33957 ;
  assign y25256 = ~1'b0 ;
  assign y25257 = ~n32070 ;
  assign y25258 = n33962 ;
  assign y25259 = ~1'b0 ;
  assign y25260 = ~n33964 ;
  assign y25261 = ~n33967 ;
  assign y25262 = ~1'b0 ;
  assign y25263 = ~n33971 ;
  assign y25264 = ~1'b0 ;
  assign y25265 = ~1'b0 ;
  assign y25266 = n33976 ;
  assign y25267 = n5551 ;
  assign y25268 = n3497 ;
  assign y25269 = n33977 ;
  assign y25270 = ~1'b0 ;
  assign y25271 = ~1'b0 ;
  assign y25272 = n33978 ;
  assign y25273 = 1'b0 ;
  assign y25274 = ~1'b0 ;
  assign y25275 = n33979 ;
  assign y25276 = ~n33980 ;
  assign y25277 = n33981 ;
  assign y25278 = ~n2896 ;
  assign y25279 = ~1'b0 ;
  assign y25280 = ~1'b0 ;
  assign y25281 = ~1'b0 ;
  assign y25282 = ~n33983 ;
  assign y25283 = n2092 ;
  assign y25284 = ~1'b0 ;
  assign y25285 = ~n33985 ;
  assign y25286 = ~n33991 ;
  assign y25287 = 1'b0 ;
  assign y25288 = n33993 ;
  assign y25289 = n13813 ;
  assign y25290 = ~n33995 ;
  assign y25291 = n33997 ;
  assign y25292 = n34002 ;
  assign y25293 = n34003 ;
  assign y25294 = ~n34009 ;
  assign y25295 = ~n34013 ;
  assign y25296 = ~n4361 ;
  assign y25297 = ~1'b0 ;
  assign y25298 = ~n34016 ;
  assign y25299 = ~n34017 ;
  assign y25300 = ~1'b0 ;
  assign y25301 = ~1'b0 ;
  assign y25302 = n34020 ;
  assign y25303 = ~1'b0 ;
  assign y25304 = ~1'b0 ;
  assign y25305 = ~n34022 ;
  assign y25306 = ~n34026 ;
  assign y25307 = ~1'b0 ;
  assign y25308 = 1'b0 ;
  assign y25309 = 1'b0 ;
  assign y25310 = n9443 ;
  assign y25311 = n34029 ;
  assign y25312 = n34032 ;
  assign y25313 = n34033 ;
  assign y25314 = ~1'b0 ;
  assign y25315 = n34035 ;
  assign y25316 = 1'b0 ;
  assign y25317 = n34036 ;
  assign y25318 = 1'b0 ;
  assign y25319 = ~1'b0 ;
  assign y25320 = ~1'b0 ;
  assign y25321 = n34040 ;
  assign y25322 = ~1'b0 ;
  assign y25323 = n34042 ;
  assign y25324 = ~n22365 ;
  assign y25325 = 1'b0 ;
  assign y25326 = ~n34046 ;
  assign y25327 = ~n34047 ;
  assign y25328 = ~n34048 ;
  assign y25329 = ~1'b0 ;
  assign y25330 = n34050 ;
  assign y25331 = ~1'b0 ;
  assign y25332 = ~1'b0 ;
  assign y25333 = ~n34053 ;
  assign y25334 = ~n34056 ;
  assign y25335 = ~1'b0 ;
  assign y25336 = n34057 ;
  assign y25337 = ~1'b0 ;
  assign y25338 = n34058 ;
  assign y25339 = n34059 ;
  assign y25340 = n34060 ;
  assign y25341 = n34061 ;
  assign y25342 = ~n34063 ;
  assign y25343 = n34065 ;
  assign y25344 = n34071 ;
  assign y25345 = ~1'b0 ;
  assign y25346 = ~n34072 ;
  assign y25347 = n34073 ;
  assign y25348 = n34075 ;
  assign y25349 = n34077 ;
  assign y25350 = n34078 ;
  assign y25351 = n34083 ;
  assign y25352 = n34084 ;
  assign y25353 = ~n34086 ;
  assign y25354 = ~n34092 ;
  assign y25355 = n34095 ;
  assign y25356 = ~1'b0 ;
  assign y25357 = n8092 ;
  assign y25358 = n34096 ;
  assign y25359 = n34103 ;
  assign y25360 = ~n34105 ;
  assign y25361 = ~n34107 ;
  assign y25362 = n34114 ;
  assign y25363 = ~n9998 ;
  assign y25364 = n34116 ;
  assign y25365 = ~1'b0 ;
  assign y25366 = ~n34118 ;
  assign y25367 = 1'b0 ;
  assign y25368 = ~n33098 ;
  assign y25369 = n34120 ;
  assign y25370 = n34127 ;
  assign y25371 = ~n34129 ;
  assign y25372 = n34132 ;
  assign y25373 = ~1'b0 ;
  assign y25374 = n34134 ;
  assign y25375 = n34135 ;
  assign y25376 = n34139 ;
  assign y25377 = ~n31467 ;
  assign y25378 = ~n34141 ;
  assign y25379 = n34142 ;
  assign y25380 = ~1'b0 ;
  assign y25381 = ~1'b0 ;
  assign y25382 = ~1'b0 ;
  assign y25383 = ~1'b0 ;
  assign y25384 = ~1'b0 ;
  assign y25385 = ~1'b0 ;
  assign y25386 = n34143 ;
  assign y25387 = ~n34144 ;
  assign y25388 = ~n34149 ;
  assign y25389 = ~1'b0 ;
  assign y25390 = n1950 ;
  assign y25391 = ~n34151 ;
  assign y25392 = ~1'b0 ;
  assign y25393 = 1'b0 ;
  assign y25394 = ~n34153 ;
  assign y25395 = ~1'b0 ;
  assign y25396 = n34154 ;
  assign y25397 = ~1'b0 ;
  assign y25398 = n34156 ;
  assign y25399 = ~n34160 ;
  assign y25400 = ~1'b0 ;
  assign y25401 = ~1'b0 ;
  assign y25402 = 1'b0 ;
  assign y25403 = ~n34161 ;
  assign y25404 = n34162 ;
  assign y25405 = n2642 ;
  assign y25406 = ~1'b0 ;
  assign y25407 = ~1'b0 ;
  assign y25408 = ~1'b0 ;
  assign y25409 = n34163 ;
  assign y25410 = ~1'b0 ;
  assign y25411 = ~n34164 ;
  assign y25412 = ~1'b0 ;
  assign y25413 = ~1'b0 ;
  assign y25414 = ~1'b0 ;
  assign y25415 = ~1'b0 ;
  assign y25416 = ~n290 ;
  assign y25417 = n34167 ;
  assign y25418 = n9222 ;
  assign y25419 = 1'b0 ;
  assign y25420 = ~1'b0 ;
  assign y25421 = ~n34171 ;
  assign y25422 = n75 ;
  assign y25423 = n6168 ;
  assign y25424 = ~1'b0 ;
  assign y25425 = ~1'b0 ;
  assign y25426 = ~n34174 ;
  assign y25427 = ~n34175 ;
  assign y25428 = n34177 ;
  assign y25429 = ~n27235 ;
  assign y25430 = ~n34179 ;
  assign y25431 = ~n34183 ;
  assign y25432 = n34185 ;
  assign y25433 = n6955 ;
  assign y25434 = ~1'b0 ;
  assign y25435 = ~1'b0 ;
  assign y25436 = ~n34186 ;
  assign y25437 = ~1'b0 ;
  assign y25438 = 1'b0 ;
  assign y25439 = ~1'b0 ;
  assign y25440 = n18538 ;
  assign y25441 = ~1'b0 ;
  assign y25442 = ~1'b0 ;
  assign y25443 = ~n34188 ;
  assign y25444 = n34189 ;
  assign y25445 = n34191 ;
  assign y25446 = ~1'b0 ;
  assign y25447 = n34195 ;
  assign y25448 = ~1'b0 ;
  assign y25449 = ~1'b0 ;
  assign y25450 = ~n34196 ;
  assign y25451 = ~n12126 ;
  assign y25452 = ~n1202 ;
  assign y25453 = ~n34197 ;
  assign y25454 = n34198 ;
  assign y25455 = n34200 ;
  assign y25456 = ~n34201 ;
  assign y25457 = n34202 ;
  assign y25458 = ~n34203 ;
  assign y25459 = ~1'b0 ;
  assign y25460 = n34204 ;
  assign y25461 = n34206 ;
  assign y25462 = ~1'b0 ;
  assign y25463 = 1'b0 ;
  assign y25464 = ~1'b0 ;
  assign y25465 = n34207 ;
  assign y25466 = n34212 ;
  assign y25467 = n34216 ;
  assign y25468 = ~1'b0 ;
  assign y25469 = ~n20425 ;
  assign y25470 = ~n34218 ;
  assign y25471 = ~1'b0 ;
  assign y25472 = n34219 ;
  assign y25473 = ~1'b0 ;
  assign y25474 = ~n34221 ;
  assign y25475 = ~1'b0 ;
  assign y25476 = ~n34222 ;
  assign y25477 = n34226 ;
  assign y25478 = n34231 ;
  assign y25479 = ~n21059 ;
  assign y25480 = ~1'b0 ;
  assign y25481 = n34235 ;
  assign y25482 = ~1'b0 ;
  assign y25483 = 1'b0 ;
  assign y25484 = n13091 ;
  assign y25485 = ~1'b0 ;
  assign y25486 = ~n34239 ;
  assign y25487 = ~n34241 ;
  assign y25488 = n34242 ;
  assign y25489 = n34243 ;
  assign y25490 = ~n34244 ;
  assign y25491 = n12053 ;
  assign y25492 = ~n34246 ;
  assign y25493 = n34247 ;
  assign y25494 = ~n34249 ;
  assign y25495 = n34254 ;
  assign y25496 = ~1'b0 ;
  assign y25497 = ~n5259 ;
  assign y25498 = ~1'b0 ;
  assign y25499 = ~n34255 ;
  assign y25500 = ~1'b0 ;
  assign y25501 = 1'b0 ;
  assign y25502 = ~1'b0 ;
  assign y25503 = ~1'b0 ;
  assign y25504 = ~1'b0 ;
  assign y25505 = n34257 ;
  assign y25506 = n2452 ;
  assign y25507 = ~n5508 ;
  assign y25508 = ~1'b0 ;
  assign y25509 = n34262 ;
  assign y25510 = n34266 ;
  assign y25511 = ~1'b0 ;
  assign y25512 = ~1'b0 ;
  assign y25513 = ~1'b0 ;
  assign y25514 = ~1'b0 ;
  assign y25515 = n5030 ;
  assign y25516 = n34267 ;
  assign y25517 = 1'b0 ;
  assign y25518 = n34269 ;
  assign y25519 = ~1'b0 ;
  assign y25520 = n34270 ;
  assign y25521 = n34272 ;
  assign y25522 = ~1'b0 ;
  assign y25523 = ~n34273 ;
  assign y25524 = n34274 ;
  assign y25525 = ~n34276 ;
  assign y25526 = ~1'b0 ;
  assign y25527 = n34277 ;
  assign y25528 = ~n34278 ;
  assign y25529 = 1'b0 ;
  assign y25530 = ~n34280 ;
  assign y25531 = ~1'b0 ;
  assign y25532 = ~n34281 ;
  assign y25533 = n34282 ;
  assign y25534 = ~n34286 ;
  assign y25535 = ~1'b0 ;
  assign y25536 = ~n23596 ;
  assign y25537 = ~n34291 ;
  assign y25538 = ~n34293 ;
  assign y25539 = ~1'b0 ;
  assign y25540 = ~1'b0 ;
  assign y25541 = ~1'b0 ;
  assign y25542 = ~1'b0 ;
  assign y25543 = n34294 ;
  assign y25544 = ~1'b0 ;
  assign y25545 = n34295 ;
  assign y25546 = ~n14771 ;
  assign y25547 = ~n34298 ;
  assign y25548 = ~1'b0 ;
  assign y25549 = ~1'b0 ;
  assign y25550 = ~n24439 ;
  assign y25551 = ~1'b0 ;
  assign y25552 = ~n34301 ;
  assign y25553 = n34305 ;
  assign y25554 = ~n1472 ;
  assign y25555 = n34310 ;
  assign y25556 = ~n34315 ;
  assign y25557 = ~1'b0 ;
  assign y25558 = ~n34318 ;
  assign y25559 = n10245 ;
  assign y25560 = n34320 ;
  assign y25561 = ~n34338 ;
  assign y25562 = ~n34348 ;
  assign y25563 = 1'b0 ;
  assign y25564 = ~1'b0 ;
  assign y25565 = ~1'b0 ;
  assign y25566 = n34349 ;
  assign y25567 = ~1'b0 ;
  assign y25568 = ~n34351 ;
  assign y25569 = ~1'b0 ;
  assign y25570 = n34352 ;
  assign y25571 = ~n34353 ;
  assign y25572 = ~1'b0 ;
  assign y25573 = ~1'b0 ;
  assign y25574 = n857 ;
  assign y25575 = ~1'b0 ;
  assign y25576 = ~n34355 ;
  assign y25577 = ~n34359 ;
  assign y25578 = ~1'b0 ;
  assign y25579 = n6904 ;
  assign y25580 = n34361 ;
  assign y25581 = n1297 ;
  assign y25582 = n34362 ;
  assign y25583 = ~n34363 ;
  assign y25584 = n10899 ;
  assign y25585 = n34365 ;
  assign y25586 = ~n19981 ;
  assign y25587 = 1'b0 ;
  assign y25588 = ~n34366 ;
  assign y25589 = n34367 ;
  assign y25590 = ~1'b0 ;
  assign y25591 = ~n34369 ;
  assign y25592 = n34373 ;
  assign y25593 = ~n34374 ;
  assign y25594 = ~n34375 ;
  assign y25595 = ~1'b0 ;
  assign y25596 = ~n34377 ;
  assign y25597 = ~n34381 ;
  assign y25598 = n34382 ;
  assign y25599 = ~1'b0 ;
  assign y25600 = n34383 ;
  assign y25601 = ~n34385 ;
  assign y25602 = ~n19433 ;
  assign y25603 = ~1'b0 ;
  assign y25604 = n32136 ;
  assign y25605 = ~n34386 ;
  assign y25606 = ~1'b0 ;
  assign y25607 = n34388 ;
  assign y25608 = ~n34394 ;
  assign y25609 = ~n34395 ;
  assign y25610 = n34397 ;
  assign y25611 = 1'b0 ;
  assign y25612 = ~n34403 ;
  assign y25613 = ~1'b0 ;
  assign y25614 = ~n34405 ;
  assign y25615 = ~1'b0 ;
  assign y25616 = ~n34410 ;
  assign y25617 = ~n34413 ;
  assign y25618 = ~1'b0 ;
  assign y25619 = ~n34417 ;
  assign y25620 = n34418 ;
  assign y25621 = n27337 ;
  assign y25622 = 1'b0 ;
  assign y25623 = ~1'b0 ;
  assign y25624 = 1'b0 ;
  assign y25625 = n34420 ;
  assign y25626 = ~1'b0 ;
  assign y25627 = ~n34422 ;
  assign y25628 = n1756 ;
  assign y25629 = ~1'b0 ;
  assign y25630 = n34423 ;
  assign y25631 = ~1'b0 ;
  assign y25632 = ~1'b0 ;
  assign y25633 = ~n34426 ;
  assign y25634 = ~1'b0 ;
  assign y25635 = ~1'b0 ;
  assign y25636 = ~1'b0 ;
  assign y25637 = ~n34431 ;
  assign y25638 = n34433 ;
  assign y25639 = n34435 ;
  assign y25640 = ~n11624 ;
  assign y25641 = n34437 ;
  assign y25642 = ~1'b0 ;
  assign y25643 = ~n34441 ;
  assign y25644 = ~n34443 ;
  assign y25645 = ~n20954 ;
  assign y25646 = n12304 ;
  assign y25647 = ~n34446 ;
  assign y25648 = n34447 ;
  assign y25649 = ~1'b0 ;
  assign y25650 = ~1'b0 ;
  assign y25651 = ~1'b0 ;
  assign y25652 = n34449 ;
  assign y25653 = n5915 ;
  assign y25654 = ~1'b0 ;
  assign y25655 = n34452 ;
  assign y25656 = n34453 ;
  assign y25657 = n34454 ;
  assign y25658 = ~n34455 ;
  assign y25659 = n34460 ;
  assign y25660 = ~1'b0 ;
  assign y25661 = n34462 ;
  assign y25662 = n34463 ;
  assign y25663 = ~n34465 ;
  assign y25664 = ~n34467 ;
  assign y25665 = ~1'b0 ;
  assign y25666 = n34468 ;
  assign y25667 = n34469 ;
  assign y25668 = ~1'b0 ;
  assign y25669 = n34474 ;
  assign y25670 = n34476 ;
  assign y25671 = 1'b0 ;
  assign y25672 = ~1'b0 ;
  assign y25673 = n34480 ;
  assign y25674 = ~1'b0 ;
  assign y25675 = ~1'b0 ;
  assign y25676 = n34481 ;
  assign y25677 = 1'b0 ;
  assign y25678 = ~1'b0 ;
  assign y25679 = n11835 ;
  assign y25680 = ~1'b0 ;
  assign y25681 = ~n34483 ;
  assign y25682 = 1'b0 ;
  assign y25683 = ~1'b0 ;
  assign y25684 = ~n34485 ;
  assign y25685 = n34488 ;
  assign y25686 = ~1'b0 ;
  assign y25687 = ~1'b0 ;
  assign y25688 = ~n34491 ;
  assign y25689 = n34492 ;
  assign y25690 = ~1'b0 ;
  assign y25691 = ~1'b0 ;
  assign y25692 = ~n34494 ;
  assign y25693 = n34497 ;
  assign y25694 = ~1'b0 ;
  assign y25695 = ~1'b0 ;
  assign y25696 = n34499 ;
  assign y25697 = 1'b0 ;
  assign y25698 = ~1'b0 ;
  assign y25699 = ~n34501 ;
  assign y25700 = ~n34504 ;
  assign y25701 = ~1'b0 ;
  assign y25702 = ~n34505 ;
  assign y25703 = ~n34506 ;
  assign y25704 = ~1'b0 ;
  assign y25705 = ~1'b0 ;
  assign y25706 = n34509 ;
  assign y25707 = ~1'b0 ;
  assign y25708 = ~1'b0 ;
  assign y25709 = ~1'b0 ;
  assign y25710 = n34510 ;
  assign y25711 = ~n34512 ;
  assign y25712 = ~n34518 ;
  assign y25713 = ~1'b0 ;
  assign y25714 = n34523 ;
  assign y25715 = ~1'b0 ;
  assign y25716 = n15093 ;
  assign y25717 = ~n23727 ;
  assign y25718 = ~n34525 ;
  assign y25719 = ~n34526 ;
  assign y25720 = ~n34527 ;
  assign y25721 = ~1'b0 ;
  assign y25722 = ~n34530 ;
  assign y25723 = ~1'b0 ;
  assign y25724 = ~1'b0 ;
  assign y25725 = n34531 ;
  assign y25726 = n34533 ;
  assign y25727 = n34535 ;
  assign y25728 = ~1'b0 ;
  assign y25729 = ~n34537 ;
  assign y25730 = n34541 ;
  assign y25731 = ~1'b0 ;
  assign y25732 = ~1'b0 ;
  assign y25733 = n34542 ;
  assign y25734 = ~n34545 ;
  assign y25735 = n34547 ;
  assign y25736 = ~n34549 ;
  assign y25737 = ~1'b0 ;
  assign y25738 = ~1'b0 ;
  assign y25739 = ~n34551 ;
  assign y25740 = ~1'b0 ;
  assign y25741 = ~n34553 ;
  assign y25742 = ~1'b0 ;
  assign y25743 = ~n34554 ;
  assign y25744 = ~1'b0 ;
  assign y25745 = ~1'b0 ;
  assign y25746 = ~1'b0 ;
  assign y25747 = ~1'b0 ;
  assign y25748 = ~n34555 ;
  assign y25749 = ~n34557 ;
  assign y25750 = n34560 ;
  assign y25751 = n34564 ;
  assign y25752 = ~n34569 ;
  assign y25753 = ~1'b0 ;
  assign y25754 = ~1'b0 ;
  assign y25755 = n34570 ;
  assign y25756 = ~1'b0 ;
  assign y25757 = ~n34571 ;
  assign y25758 = ~n34572 ;
  assign y25759 = ~1'b0 ;
  assign y25760 = ~1'b0 ;
  assign y25761 = ~n34573 ;
  assign y25762 = n34575 ;
  assign y25763 = ~n37 ;
  assign y25764 = ~1'b0 ;
  assign y25765 = n34576 ;
  assign y25766 = ~n34578 ;
  assign y25767 = ~n11463 ;
  assign y25768 = ~n34582 ;
  assign y25769 = ~n34583 ;
  assign y25770 = n34607 ;
  assign y25771 = ~n34608 ;
  assign y25772 = n34612 ;
  assign y25773 = n6422 ;
  assign y25774 = ~1'b0 ;
  assign y25775 = ~1'b0 ;
  assign y25776 = n34613 ;
  assign y25777 = n34614 ;
  assign y25778 = ~n34615 ;
  assign y25779 = x4 ;
  assign y25780 = ~n34618 ;
  assign y25781 = n34627 ;
  assign y25782 = n34636 ;
  assign y25783 = ~1'b0 ;
  assign y25784 = ~n9218 ;
  assign y25785 = ~n34638 ;
  assign y25786 = 1'b0 ;
  assign y25787 = n34641 ;
  assign y25788 = n21338 ;
  assign y25789 = n34644 ;
  assign y25790 = n34646 ;
  assign y25791 = ~1'b0 ;
  assign y25792 = ~n34648 ;
  assign y25793 = n34655 ;
  assign y25794 = n34657 ;
  assign y25795 = ~1'b0 ;
  assign y25796 = ~1'b0 ;
  assign y25797 = n34658 ;
  assign y25798 = n34659 ;
  assign y25799 = n34660 ;
  assign y25800 = ~1'b0 ;
  assign y25801 = n34661 ;
  assign y25802 = ~n34662 ;
  assign y25803 = n34664 ;
  assign y25804 = n34667 ;
  assign y25805 = ~n811 ;
  assign y25806 = ~1'b0 ;
  assign y25807 = 1'b0 ;
  assign y25808 = ~n34670 ;
  assign y25809 = ~1'b0 ;
  assign y25810 = ~1'b0 ;
  assign y25811 = ~n34675 ;
  assign y25812 = n34680 ;
  assign y25813 = n34684 ;
  assign y25814 = ~1'b0 ;
  assign y25815 = ~1'b0 ;
  assign y25816 = ~1'b0 ;
  assign y25817 = ~1'b0 ;
  assign y25818 = ~1'b0 ;
  assign y25819 = 1'b0 ;
  assign y25820 = ~n34687 ;
  assign y25821 = ~1'b0 ;
  assign y25822 = ~1'b0 ;
  assign y25823 = ~1'b0 ;
  assign y25824 = ~n34688 ;
  assign y25825 = ~n34690 ;
  assign y25826 = n34703 ;
  assign y25827 = ~1'b0 ;
  assign y25828 = ~n34705 ;
  assign y25829 = ~n34706 ;
  assign y25830 = ~1'b0 ;
  assign y25831 = ~1'b0 ;
  assign y25832 = ~1'b0 ;
  assign y25833 = n34707 ;
  assign y25834 = 1'b0 ;
  assign y25835 = ~n2316 ;
  assign y25836 = ~1'b0 ;
  assign y25837 = ~n34710 ;
  assign y25838 = n6295 ;
  assign y25839 = ~n34716 ;
  assign y25840 = n34718 ;
  assign y25841 = ~n34727 ;
  assign y25842 = ~n6433 ;
  assign y25843 = n34732 ;
  assign y25844 = n34734 ;
  assign y25845 = ~1'b0 ;
  assign y25846 = ~1'b0 ;
  assign y25847 = ~1'b0 ;
  assign y25848 = ~n34735 ;
  assign y25849 = ~n28103 ;
  assign y25850 = ~1'b0 ;
  assign y25851 = ~n34736 ;
  assign y25852 = n34740 ;
  assign y25853 = ~n34744 ;
  assign y25854 = n769 ;
  assign y25855 = ~n34746 ;
  assign y25856 = n34747 ;
  assign y25857 = n22048 ;
  assign y25858 = ~1'b0 ;
  assign y25859 = ~1'b0 ;
  assign y25860 = ~1'b0 ;
  assign y25861 = ~1'b0 ;
  assign y25862 = ~1'b0 ;
  assign y25863 = ~1'b0 ;
  assign y25864 = ~n34750 ;
  assign y25865 = ~n17675 ;
  assign y25866 = 1'b0 ;
  assign y25867 = ~1'b0 ;
  assign y25868 = n34752 ;
  assign y25869 = n34753 ;
  assign y25870 = n34762 ;
  assign y25871 = n34763 ;
  assign y25872 = n34764 ;
  assign y25873 = ~1'b0 ;
  assign y25874 = n34766 ;
  assign y25875 = ~n34767 ;
  assign y25876 = ~1'b0 ;
  assign y25877 = n34770 ;
  assign y25878 = ~1'b0 ;
  assign y25879 = ~1'b0 ;
  assign y25880 = ~n34772 ;
  assign y25881 = ~n34774 ;
  assign y25882 = ~n5000 ;
  assign y25883 = n34777 ;
  assign y25884 = ~n34779 ;
  assign y25885 = ~1'b0 ;
  assign y25886 = n34780 ;
  assign y25887 = ~n25411 ;
  assign y25888 = ~1'b0 ;
  assign y25889 = ~n34782 ;
  assign y25890 = ~1'b0 ;
  assign y25891 = ~1'b0 ;
  assign y25892 = n34787 ;
  assign y25893 = n34788 ;
  assign y25894 = ~n34789 ;
  assign y25895 = ~n34791 ;
  assign y25896 = ~n34794 ;
  assign y25897 = n34795 ;
  assign y25898 = ~n34797 ;
  assign y25899 = ~1'b0 ;
  assign y25900 = n34800 ;
  assign y25901 = ~n34802 ;
  assign y25902 = n2233 ;
  assign y25903 = n34808 ;
  assign y25904 = ~1'b0 ;
  assign y25905 = 1'b0 ;
  assign y25906 = ~1'b0 ;
  assign y25907 = ~1'b0 ;
  assign y25908 = ~n34809 ;
  assign y25909 = n3131 ;
  assign y25910 = ~1'b0 ;
  assign y25911 = ~n34810 ;
  assign y25912 = n34811 ;
  assign y25913 = ~n34813 ;
  assign y25914 = ~n34816 ;
  assign y25915 = n34820 ;
  assign y25916 = ~1'b0 ;
  assign y25917 = n34821 ;
  assign y25918 = n34822 ;
  assign y25919 = ~n16153 ;
  assign y25920 = n34826 ;
  assign y25921 = n34828 ;
  assign y25922 = ~1'b0 ;
  assign y25923 = 1'b0 ;
  assign y25924 = ~n34829 ;
  assign y25925 = n34836 ;
  assign y25926 = ~1'b0 ;
  assign y25927 = ~n34838 ;
  assign y25928 = ~1'b0 ;
  assign y25929 = ~1'b0 ;
  assign y25930 = ~n34839 ;
  assign y25931 = ~1'b0 ;
  assign y25932 = ~n34842 ;
  assign y25933 = 1'b0 ;
  assign y25934 = n34844 ;
  assign y25935 = ~1'b0 ;
  assign y25936 = ~n34846 ;
  assign y25937 = ~n34848 ;
  assign y25938 = n34849 ;
  assign y25939 = ~1'b0 ;
  assign y25940 = n33239 ;
  assign y25941 = n17161 ;
  assign y25942 = n34852 ;
  assign y25943 = ~n34854 ;
  assign y25944 = ~1'b0 ;
  assign y25945 = ~1'b0 ;
  assign y25946 = 1'b0 ;
  assign y25947 = n34856 ;
  assign y25948 = ~n34858 ;
  assign y25949 = ~1'b0 ;
  assign y25950 = ~n34859 ;
  assign y25951 = n34860 ;
  assign y25952 = ~1'b0 ;
  assign y25953 = ~1'b0 ;
  assign y25954 = 1'b0 ;
  assign y25955 = n34861 ;
  assign y25956 = ~n34865 ;
  assign y25957 = ~n19439 ;
  assign y25958 = ~1'b0 ;
  assign y25959 = ~1'b0 ;
  assign y25960 = ~1'b0 ;
  assign y25961 = ~n34866 ;
  assign y25962 = n34868 ;
  assign y25963 = ~n34869 ;
  assign y25964 = 1'b0 ;
  assign y25965 = n34871 ;
  assign y25966 = ~n1233 ;
  assign y25967 = n34873 ;
  assign y25968 = ~1'b0 ;
  assign y25969 = n532 ;
  assign y25970 = ~n34874 ;
  assign y25971 = ~1'b0 ;
  assign y25972 = ~1'b0 ;
  assign y25973 = n21683 ;
  assign y25974 = ~1'b0 ;
  assign y25975 = n2155 ;
  assign y25976 = n34875 ;
  assign y25977 = 1'b0 ;
  assign y25978 = n34876 ;
  assign y25979 = n34881 ;
  assign y25980 = ~n34884 ;
  assign y25981 = ~n34885 ;
  assign y25982 = n34889 ;
  assign y25983 = 1'b0 ;
  assign y25984 = ~n34890 ;
  assign y25985 = ~n34892 ;
  assign y25986 = ~n34894 ;
  assign y25987 = n6770 ;
  assign y25988 = 1'b0 ;
  assign y25989 = n33060 ;
  assign y25990 = ~1'b0 ;
  assign y25991 = ~1'b0 ;
  assign y25992 = n34901 ;
  assign y25993 = ~1'b0 ;
  assign y25994 = 1'b0 ;
  assign y25995 = ~n14226 ;
  assign y25996 = n34902 ;
  assign y25997 = ~1'b0 ;
  assign y25998 = ~n34903 ;
  assign y25999 = n19117 ;
  assign y26000 = n34904 ;
  assign y26001 = ~n34905 ;
  assign y26002 = n34906 ;
  assign y26003 = ~n34907 ;
  assign y26004 = n34910 ;
  assign y26005 = ~1'b0 ;
  assign y26006 = ~1'b0 ;
  assign y26007 = ~n34912 ;
  assign y26008 = ~n14975 ;
  assign y26009 = n5162 ;
  assign y26010 = 1'b0 ;
  assign y26011 = ~n1777 ;
  assign y26012 = ~1'b0 ;
  assign y26013 = ~1'b0 ;
  assign y26014 = ~n34913 ;
  assign y26015 = n34936 ;
  assign y26016 = ~1'b0 ;
  assign y26017 = n34938 ;
  assign y26018 = n34939 ;
  assign y26019 = n534 ;
  assign y26020 = n34943 ;
  assign y26021 = ~n34945 ;
  assign y26022 = ~1'b0 ;
  assign y26023 = ~n34946 ;
  assign y26024 = n34950 ;
  assign y26025 = ~1'b0 ;
  assign y26026 = ~1'b0 ;
  assign y26027 = ~1'b0 ;
  assign y26028 = ~1'b0 ;
  assign y26029 = ~n34952 ;
  assign y26030 = 1'b0 ;
  assign y26031 = n34954 ;
  assign y26032 = n34956 ;
  assign y26033 = n3730 ;
  assign y26034 = ~1'b0 ;
  assign y26035 = 1'b0 ;
  assign y26036 = ~n34957 ;
  assign y26037 = 1'b0 ;
  assign y26038 = n34960 ;
  assign y26039 = ~n34961 ;
  assign y26040 = n34964 ;
  assign y26041 = ~1'b0 ;
  assign y26042 = n21847 ;
  assign y26043 = n34965 ;
  assign y26044 = ~n34079 ;
  assign y26045 = ~1'b0 ;
  assign y26046 = ~1'b0 ;
  assign y26047 = n34967 ;
  assign y26048 = ~1'b0 ;
  assign y26049 = ~n34970 ;
  assign y26050 = ~1'b0 ;
  assign y26051 = ~1'b0 ;
  assign y26052 = ~n34972 ;
  assign y26053 = n33806 ;
  assign y26054 = n34973 ;
  assign y26055 = ~1'b0 ;
  assign y26056 = n518 ;
  assign y26057 = ~1'b0 ;
  assign y26058 = n34974 ;
  assign y26059 = 1'b0 ;
  assign y26060 = ~1'b0 ;
  assign y26061 = n34978 ;
  assign y26062 = ~n34983 ;
  assign y26063 = ~n2526 ;
  assign y26064 = ~n34986 ;
  assign y26065 = ~n34994 ;
  assign y26066 = ~n35000 ;
  assign y26067 = ~n35007 ;
  assign y26068 = n24371 ;
  assign y26069 = ~1'b0 ;
  assign y26070 = n35008 ;
  assign y26071 = ~1'b0 ;
  assign y26072 = ~1'b0 ;
  assign y26073 = n35009 ;
  assign y26074 = n35012 ;
  assign y26075 = n615 ;
  assign y26076 = ~1'b0 ;
  assign y26077 = ~n35014 ;
  assign y26078 = ~1'b0 ;
  assign y26079 = ~n35015 ;
  assign y26080 = ~n35017 ;
  assign y26081 = ~1'b0 ;
  assign y26082 = n35018 ;
  assign y26083 = ~1'b0 ;
  assign y26084 = ~1'b0 ;
  assign y26085 = ~n35019 ;
  assign y26086 = ~n3371 ;
  assign y26087 = ~1'b0 ;
  assign y26088 = ~1'b0 ;
  assign y26089 = ~1'b0 ;
  assign y26090 = ~1'b0 ;
  assign y26091 = ~1'b0 ;
  assign y26092 = ~n35022 ;
  assign y26093 = ~n35023 ;
  assign y26094 = n35025 ;
  assign y26095 = n33977 ;
  assign y26096 = ~n35026 ;
  assign y26097 = n35027 ;
  assign y26098 = ~n35029 ;
  assign y26099 = n35030 ;
  assign y26100 = ~n35032 ;
  assign y26101 = ~1'b0 ;
  assign y26102 = ~1'b0 ;
  assign y26103 = ~n35034 ;
  assign y26104 = ~1'b0 ;
  assign y26105 = ~n35035 ;
  assign y26106 = ~1'b0 ;
  assign y26107 = ~1'b0 ;
  assign y26108 = ~1'b0 ;
  assign y26109 = ~1'b0 ;
  assign y26110 = n35038 ;
  assign y26111 = ~n35039 ;
  assign y26112 = 1'b0 ;
  assign y26113 = n35041 ;
  assign y26114 = ~1'b0 ;
  assign y26115 = n35043 ;
  assign y26116 = ~n5952 ;
  assign y26117 = ~1'b0 ;
  assign y26118 = ~1'b0 ;
  assign y26119 = ~1'b0 ;
  assign y26120 = ~1'b0 ;
  assign y26121 = n9980 ;
  assign y26122 = n35045 ;
  assign y26123 = 1'b0 ;
  assign y26124 = ~1'b0 ;
  assign y26125 = n35046 ;
  assign y26126 = ~n35048 ;
  assign y26127 = ~n35049 ;
  assign y26128 = ~1'b0 ;
  assign y26129 = ~1'b0 ;
  assign y26130 = n35054 ;
  assign y26131 = 1'b0 ;
  assign y26132 = ~1'b0 ;
  assign y26133 = n35056 ;
  assign y26134 = n35057 ;
  assign y26135 = n35058 ;
  assign y26136 = ~n35063 ;
  assign y26137 = n35065 ;
  assign y26138 = ~n35066 ;
  assign y26139 = n35067 ;
  assign y26140 = n35069 ;
  assign y26141 = ~n35070 ;
  assign y26142 = ~n35072 ;
  assign y26143 = n35074 ;
  assign y26144 = n3722 ;
  assign y26145 = n35075 ;
  assign y26146 = ~n35076 ;
  assign y26147 = ~n35078 ;
  assign y26148 = ~n35080 ;
  assign y26149 = n35082 ;
  assign y26150 = ~n35087 ;
  assign y26151 = ~n35088 ;
  assign y26152 = ~1'b0 ;
  assign y26153 = ~n35089 ;
  assign y26154 = ~1'b0 ;
  assign y26155 = ~1'b0 ;
  assign y26156 = n35091 ;
  assign y26157 = n8099 ;
  assign y26158 = ~n1214 ;
  assign y26159 = ~1'b0 ;
  assign y26160 = ~n4927 ;
  assign y26161 = n35092 ;
  assign y26162 = ~n35094 ;
  assign y26163 = n35098 ;
  assign y26164 = ~1'b0 ;
  assign y26165 = ~n35099 ;
  assign y26166 = n35100 ;
  assign y26167 = 1'b0 ;
  assign y26168 = 1'b0 ;
  assign y26169 = n35102 ;
  assign y26170 = ~1'b0 ;
  assign y26171 = n35103 ;
  assign y26172 = n31709 ;
  assign y26173 = ~n35105 ;
  assign y26174 = ~1'b0 ;
  assign y26175 = ~n35107 ;
  assign y26176 = n7812 ;
  assign y26177 = ~n35109 ;
  assign y26178 = n35111 ;
  assign y26179 = ~n35113 ;
  assign y26180 = n35114 ;
  assign y26181 = 1'b0 ;
  assign y26182 = ~n1426 ;
  assign y26183 = n35115 ;
  assign y26184 = n35116 ;
  assign y26185 = 1'b0 ;
  assign y26186 = n35118 ;
  assign y26187 = ~1'b0 ;
  assign y26188 = ~n19099 ;
  assign y26189 = ~n35122 ;
  assign y26190 = n7352 ;
  assign y26191 = ~n35123 ;
  assign y26192 = 1'b0 ;
  assign y26193 = ~n35125 ;
  assign y26194 = ~1'b0 ;
  assign y26195 = n35127 ;
  assign y26196 = ~n35134 ;
  assign y26197 = ~1'b0 ;
  assign y26198 = ~1'b0 ;
  assign y26199 = n35137 ;
  assign y26200 = n35140 ;
  assign y26201 = ~1'b0 ;
  assign y26202 = ~n35141 ;
  assign y26203 = ~n35142 ;
  assign y26204 = ~n35150 ;
  assign y26205 = n35151 ;
  assign y26206 = ~1'b0 ;
  assign y26207 = ~1'b0 ;
  assign y26208 = ~n9463 ;
  assign y26209 = ~n35153 ;
  assign y26210 = n35154 ;
  assign y26211 = ~n15713 ;
  assign y26212 = ~1'b0 ;
  assign y26213 = ~1'b0 ;
  assign y26214 = 1'b0 ;
  assign y26215 = ~n35160 ;
  assign y26216 = ~1'b0 ;
  assign y26217 = 1'b0 ;
  assign y26218 = ~n35161 ;
  assign y26219 = ~1'b0 ;
  assign y26220 = ~n17737 ;
  assign y26221 = 1'b0 ;
  assign y26222 = ~n16777 ;
  assign y26223 = ~1'b0 ;
  assign y26224 = ~1'b0 ;
  assign y26225 = ~1'b0 ;
  assign y26226 = ~n5905 ;
  assign y26227 = ~1'b0 ;
  assign y26228 = ~n35162 ;
  assign y26229 = 1'b0 ;
  assign y26230 = ~n7156 ;
  assign y26231 = ~1'b0 ;
  assign y26232 = n35164 ;
  assign y26233 = n35165 ;
  assign y26234 = ~1'b0 ;
  assign y26235 = ~1'b0 ;
  assign y26236 = ~n35168 ;
  assign y26237 = n35170 ;
  assign y26238 = ~1'b0 ;
  assign y26239 = ~1'b0 ;
  assign y26240 = ~1'b0 ;
  assign y26241 = ~n35171 ;
  assign y26242 = n35173 ;
  assign y26243 = ~n35174 ;
  assign y26244 = 1'b0 ;
  assign y26245 = n35175 ;
  assign y26246 = ~1'b0 ;
  assign y26247 = ~n35176 ;
  assign y26248 = ~n20787 ;
  assign y26249 = n35177 ;
  assign y26250 = ~n1486 ;
  assign y26251 = ~1'b0 ;
  assign y26252 = n35179 ;
  assign y26253 = 1'b0 ;
  assign y26254 = ~n35180 ;
  assign y26255 = ~1'b0 ;
  assign y26256 = n35186 ;
  assign y26257 = ~n35189 ;
  assign y26258 = ~1'b0 ;
  assign y26259 = ~1'b0 ;
  assign y26260 = n35190 ;
  assign y26261 = ~1'b0 ;
  assign y26262 = n10909 ;
  assign y26263 = n31520 ;
  assign y26264 = ~1'b0 ;
  assign y26265 = ~n10798 ;
  assign y26266 = n35192 ;
  assign y26267 = ~1'b0 ;
  assign y26268 = ~1'b0 ;
  assign y26269 = n35193 ;
  assign y26270 = 1'b0 ;
  assign y26271 = n35194 ;
  assign y26272 = ~1'b0 ;
  assign y26273 = ~1'b0 ;
  assign y26274 = ~n35201 ;
  assign y26275 = ~n35202 ;
  assign y26276 = ~n28323 ;
  assign y26277 = n35204 ;
  assign y26278 = n35205 ;
  assign y26279 = n35206 ;
  assign y26280 = ~1'b0 ;
  assign y26281 = ~n35208 ;
  assign y26282 = ~n35211 ;
  assign y26283 = ~1'b0 ;
  assign y26284 = n35215 ;
  assign y26285 = ~1'b0 ;
  assign y26286 = n7657 ;
  assign y26287 = ~n35217 ;
  assign y26288 = n35219 ;
  assign y26289 = 1'b0 ;
  assign y26290 = ~1'b0 ;
  assign y26291 = n35221 ;
  assign y26292 = n35224 ;
  assign y26293 = n35226 ;
  assign y26294 = n35227 ;
  assign y26295 = ~1'b0 ;
  assign y26296 = ~n35229 ;
  assign y26297 = n35231 ;
  assign y26298 = 1'b0 ;
  assign y26299 = n35237 ;
  assign y26300 = n35238 ;
  assign y26301 = n35242 ;
  assign y26302 = ~n35243 ;
  assign y26303 = ~1'b0 ;
  assign y26304 = ~1'b0 ;
  assign y26305 = n3414 ;
  assign y26306 = ~1'b0 ;
  assign y26307 = 1'b0 ;
  assign y26308 = ~1'b0 ;
  assign y26309 = n35244 ;
  assign y26310 = ~1'b0 ;
  assign y26311 = ~1'b0 ;
  assign y26312 = n35247 ;
  assign y26313 = n23650 ;
  assign y26314 = n35250 ;
  assign y26315 = ~1'b0 ;
  assign y26316 = ~1'b0 ;
  assign y26317 = n35252 ;
  assign y26318 = 1'b0 ;
  assign y26319 = n35253 ;
  assign y26320 = ~n35255 ;
  assign y26321 = ~n35258 ;
  assign y26322 = ~1'b0 ;
  assign y26323 = ~1'b0 ;
  assign y26324 = n35259 ;
  assign y26325 = ~1'b0 ;
  assign y26326 = n35263 ;
  assign y26327 = n8930 ;
  assign y26328 = n35264 ;
  assign y26329 = ~1'b0 ;
  assign y26330 = ~1'b0 ;
  assign y26331 = ~1'b0 ;
  assign y26332 = n35266 ;
  assign y26333 = ~n35267 ;
  assign y26334 = ~n35268 ;
  assign y26335 = ~n35269 ;
  assign y26336 = n35272 ;
  assign y26337 = ~1'b0 ;
  assign y26338 = ~1'b0 ;
  assign y26339 = ~n35273 ;
  assign y26340 = n9186 ;
  assign y26341 = ~n35276 ;
  assign y26342 = ~n35278 ;
  assign y26343 = ~n18821 ;
  assign y26344 = ~1'b0 ;
  assign y26345 = ~1'b0 ;
  assign y26346 = ~1'b0 ;
  assign y26347 = ~1'b0 ;
  assign y26348 = ~1'b0 ;
  assign y26349 = n35279 ;
  assign y26350 = 1'b0 ;
  assign y26351 = n35281 ;
  assign y26352 = ~1'b0 ;
  assign y26353 = n35283 ;
  assign y26354 = ~1'b0 ;
  assign y26355 = ~n11837 ;
  assign y26356 = ~n35284 ;
  assign y26357 = ~n35286 ;
  assign y26358 = n35288 ;
  assign y26359 = n35291 ;
  assign y26360 = ~n35293 ;
  assign y26361 = ~1'b0 ;
  assign y26362 = 1'b0 ;
  assign y26363 = n35295 ;
  assign y26364 = n10131 ;
  assign y26365 = ~n35296 ;
  assign y26366 = ~n35298 ;
  assign y26367 = ~1'b0 ;
  assign y26368 = n35301 ;
  assign y26369 = ~n35304 ;
  assign y26370 = ~n35305 ;
  assign y26371 = n35308 ;
  assign y26372 = ~1'b0 ;
  assign y26373 = 1'b0 ;
  assign y26374 = ~1'b0 ;
  assign y26375 = ~n35310 ;
  assign y26376 = ~n5186 ;
  assign y26377 = n1067 ;
  assign y26378 = ~n35320 ;
  assign y26379 = ~n35322 ;
  assign y26380 = ~1'b0 ;
  assign y26381 = n35324 ;
  assign y26382 = ~1'b0 ;
  assign y26383 = n35327 ;
  assign y26384 = ~n35328 ;
  assign y26385 = ~1'b0 ;
  assign y26386 = ~1'b0 ;
  assign y26387 = n7029 ;
  assign y26388 = ~1'b0 ;
  assign y26389 = n35330 ;
  assign y26390 = ~1'b0 ;
  assign y26391 = ~1'b0 ;
  assign y26392 = ~1'b0 ;
  assign y26393 = n35332 ;
  assign y26394 = ~1'b0 ;
  assign y26395 = ~n35333 ;
  assign y26396 = ~n35335 ;
  assign y26397 = ~n35338 ;
  assign y26398 = ~n35344 ;
  assign y26399 = n35347 ;
  assign y26400 = 1'b0 ;
  assign y26401 = ~n35350 ;
  assign y26402 = n35351 ;
  assign y26403 = n35352 ;
  assign y26404 = n35353 ;
  assign y26405 = n35355 ;
  assign y26406 = n35357 ;
  assign y26407 = ~n35360 ;
  assign y26408 = ~1'b0 ;
  assign y26409 = n35363 ;
  assign y26410 = ~1'b0 ;
  assign y26411 = ~1'b0 ;
  assign y26412 = ~n35364 ;
  assign y26413 = n35365 ;
  assign y26414 = n35366 ;
  assign y26415 = ~1'b0 ;
  assign y26416 = ~1'b0 ;
  assign y26417 = ~n35368 ;
  assign y26418 = ~n35372 ;
  assign y26419 = 1'b0 ;
  assign y26420 = n35375 ;
  assign y26421 = ~n35376 ;
  assign y26422 = ~1'b0 ;
  assign y26423 = n9907 ;
  assign y26424 = ~1'b0 ;
  assign y26425 = ~1'b0 ;
  assign y26426 = n35377 ;
  assign y26427 = ~1'b0 ;
  assign y26428 = 1'b0 ;
  assign y26429 = ~n35380 ;
  assign y26430 = n35381 ;
  assign y26431 = n35382 ;
  assign y26432 = n35385 ;
  assign y26433 = n7344 ;
  assign y26434 = ~n35387 ;
  assign y26435 = ~1'b0 ;
  assign y26436 = n35389 ;
  assign y26437 = ~n35393 ;
  assign y26438 = n35395 ;
  assign y26439 = ~1'b0 ;
  assign y26440 = ~n35396 ;
  assign y26441 = 1'b0 ;
  assign y26442 = n35398 ;
  assign y26443 = ~n35401 ;
  assign y26444 = ~n35402 ;
  assign y26445 = ~n35403 ;
  assign y26446 = n35405 ;
  assign y26447 = ~n35407 ;
  assign y26448 = ~1'b0 ;
  assign y26449 = ~1'b0 ;
  assign y26450 = ~1'b0 ;
  assign y26451 = n35409 ;
  assign y26452 = ~n35417 ;
  assign y26453 = n35420 ;
  assign y26454 = ~1'b0 ;
  assign y26455 = ~n24655 ;
  assign y26456 = ~n35421 ;
  assign y26457 = ~n35424 ;
  assign y26458 = n35426 ;
  assign y26459 = ~n35432 ;
  assign y26460 = n35433 ;
  assign y26461 = ~1'b0 ;
  assign y26462 = ~n35434 ;
  assign y26463 = ~1'b0 ;
  assign y26464 = ~n35439 ;
  assign y26465 = ~1'b0 ;
  assign y26466 = ~1'b0 ;
  assign y26467 = ~1'b0 ;
  assign y26468 = ~1'b0 ;
  assign y26469 = n35441 ;
  assign y26470 = 1'b0 ;
  assign y26471 = n35446 ;
  assign y26472 = n35447 ;
  assign y26473 = n35449 ;
  assign y26474 = ~1'b0 ;
  assign y26475 = n35450 ;
  assign y26476 = ~n35451 ;
  assign y26477 = n35454 ;
  assign y26478 = ~1'b0 ;
  assign y26479 = ~n13766 ;
  assign y26480 = ~1'b0 ;
  assign y26481 = ~1'b0 ;
  assign y26482 = n35455 ;
  assign y26483 = ~1'b0 ;
  assign y26484 = ~n159 ;
  assign y26485 = n35458 ;
  assign y26486 = ~n35460 ;
  assign y26487 = ~n35465 ;
  assign y26488 = ~n35466 ;
  assign y26489 = n35469 ;
  assign y26490 = ~1'b0 ;
  assign y26491 = n35470 ;
  assign y26492 = n22135 ;
  assign y26493 = ~n3613 ;
  assign y26494 = n35472 ;
  assign y26495 = ~1'b0 ;
  assign y26496 = ~1'b0 ;
  assign y26497 = ~n35473 ;
  assign y26498 = ~1'b0 ;
  assign y26499 = ~n35474 ;
  assign y26500 = ~n35475 ;
  assign y26501 = ~1'b0 ;
  assign y26502 = ~1'b0 ;
  assign y26503 = n9072 ;
  assign y26504 = ~1'b0 ;
  assign y26505 = ~1'b0 ;
  assign y26506 = ~n35478 ;
  assign y26507 = ~n35479 ;
  assign y26508 = n35480 ;
  assign y26509 = n35485 ;
  assign y26510 = ~n35489 ;
  assign y26511 = ~1'b0 ;
  assign y26512 = ~1'b0 ;
  assign y26513 = n35493 ;
  assign y26514 = ~n35494 ;
  assign y26515 = ~n35498 ;
  assign y26516 = ~1'b0 ;
  assign y26517 = ~n35500 ;
  assign y26518 = n35501 ;
  assign y26519 = ~n35502 ;
  assign y26520 = ~1'b0 ;
  assign y26521 = ~n35505 ;
  assign y26522 = ~1'b0 ;
  assign y26523 = ~n35509 ;
  assign y26524 = ~1'b0 ;
  assign y26525 = ~n35511 ;
  assign y26526 = 1'b0 ;
  assign y26527 = n35514 ;
  assign y26528 = ~n35517 ;
  assign y26529 = ~n35518 ;
  assign y26530 = ~1'b0 ;
  assign y26531 = ~n35521 ;
  assign y26532 = ~1'b0 ;
  assign y26533 = ~1'b0 ;
  assign y26534 = ~n35524 ;
  assign y26535 = ~n35525 ;
  assign y26536 = ~1'b0 ;
  assign y26537 = ~1'b0 ;
  assign y26538 = ~n35529 ;
  assign y26539 = ~1'b0 ;
  assign y26540 = n35530 ;
  assign y26541 = ~n35537 ;
  assign y26542 = ~n35543 ;
  assign y26543 = ~n35544 ;
  assign y26544 = ~1'b0 ;
  assign y26545 = ~n469 ;
  assign y26546 = ~n35549 ;
  assign y26547 = ~n33138 ;
  assign y26548 = ~n2377 ;
  assign y26549 = ~1'b0 ;
  assign y26550 = ~1'b0 ;
  assign y26551 = ~n35550 ;
  assign y26552 = n4522 ;
  assign y26553 = n35551 ;
  assign y26554 = n35552 ;
  assign y26555 = 1'b0 ;
  assign y26556 = ~1'b0 ;
  assign y26557 = n35553 ;
  assign y26558 = ~1'b0 ;
  assign y26559 = n35554 ;
  assign y26560 = n35555 ;
  assign y26561 = ~n35556 ;
  assign y26562 = ~n35562 ;
  assign y26563 = ~n35563 ;
  assign y26564 = ~1'b0 ;
  assign y26565 = ~n35566 ;
  assign y26566 = ~n4469 ;
  assign y26567 = n35568 ;
  assign y26568 = ~1'b0 ;
  assign y26569 = n35569 ;
  assign y26570 = ~1'b0 ;
  assign y26571 = n35570 ;
  assign y26572 = ~n35573 ;
  assign y26573 = ~1'b0 ;
  assign y26574 = ~1'b0 ;
  assign y26575 = ~n35575 ;
  assign y26576 = ~1'b0 ;
  assign y26577 = ~1'b0 ;
  assign y26578 = ~1'b0 ;
  assign y26579 = ~n35576 ;
  assign y26580 = n35577 ;
  assign y26581 = ~n35578 ;
  assign y26582 = ~1'b0 ;
  assign y26583 = ~n35579 ;
  assign y26584 = ~1'b0 ;
  assign y26585 = n35580 ;
  assign y26586 = ~1'b0 ;
  assign y26587 = n35583 ;
  assign y26588 = ~1'b0 ;
  assign y26589 = ~1'b0 ;
  assign y26590 = n35586 ;
  assign y26591 = ~n35588 ;
  assign y26592 = ~n35590 ;
  assign y26593 = ~1'b0 ;
  assign y26594 = ~n35592 ;
  assign y26595 = ~n35596 ;
  assign y26596 = ~n35597 ;
  assign y26597 = ~1'b0 ;
  assign y26598 = ~1'b0 ;
  assign y26599 = ~n35600 ;
  assign y26600 = ~n35601 ;
  assign y26601 = 1'b0 ;
  assign y26602 = n35604 ;
  assign y26603 = ~n35610 ;
  assign y26604 = ~1'b0 ;
  assign y26605 = ~n35617 ;
  assign y26606 = ~n35621 ;
  assign y26607 = n21369 ;
  assign y26608 = ~1'b0 ;
  assign y26609 = ~1'b0 ;
  assign y26610 = n35625 ;
  assign y26611 = ~1'b0 ;
  assign y26612 = ~1'b0 ;
  assign y26613 = ~n35629 ;
  assign y26614 = ~1'b0 ;
  assign y26615 = ~n19565 ;
  assign y26616 = n35632 ;
  assign y26617 = n35634 ;
  assign y26618 = ~n35638 ;
  assign y26619 = ~1'b0 ;
  assign y26620 = ~1'b0 ;
  assign y26621 = n35639 ;
  assign y26622 = ~1'b0 ;
  assign y26623 = ~n5130 ;
  assign y26624 = ~n35640 ;
  assign y26625 = 1'b0 ;
  assign y26626 = ~1'b0 ;
  assign y26627 = n35643 ;
  assign y26628 = n35647 ;
  assign y26629 = n35649 ;
  assign y26630 = n14051 ;
  assign y26631 = ~1'b0 ;
  assign y26632 = ~1'b0 ;
  assign y26633 = ~n35651 ;
  assign y26634 = ~1'b0 ;
  assign y26635 = ~1'b0 ;
  assign y26636 = ~1'b0 ;
  assign y26637 = n35654 ;
  assign y26638 = n35656 ;
  assign y26639 = n35659 ;
  assign y26640 = n35660 ;
  assign y26641 = ~1'b0 ;
  assign y26642 = n24025 ;
  assign y26643 = n4115 ;
  assign y26644 = n2047 ;
  assign y26645 = ~1'b0 ;
  assign y26646 = 1'b0 ;
  assign y26647 = 1'b0 ;
  assign y26648 = n35661 ;
  assign y26649 = n35664 ;
  assign y26650 = n35665 ;
  assign y26651 = ~n35666 ;
  assign y26652 = ~n35667 ;
  assign y26653 = n35668 ;
  assign y26654 = ~1'b0 ;
  assign y26655 = ~n28684 ;
  assign y26656 = ~n35670 ;
  assign y26657 = n35671 ;
  assign y26658 = ~1'b0 ;
  assign y26659 = n35675 ;
  assign y26660 = ~1'b0 ;
  assign y26661 = n35678 ;
  assign y26662 = ~1'b0 ;
  assign y26663 = ~n35680 ;
  assign y26664 = ~1'b0 ;
  assign y26665 = ~1'b0 ;
  assign y26666 = ~1'b0 ;
  assign y26667 = n35682 ;
  assign y26668 = n35685 ;
  assign y26669 = ~n35686 ;
  assign y26670 = ~n35687 ;
  assign y26671 = ~1'b0 ;
  assign y26672 = ~n35688 ;
  assign y26673 = ~1'b0 ;
  assign y26674 = n35691 ;
  assign y26675 = n35692 ;
  assign y26676 = ~1'b0 ;
  assign y26677 = n35696 ;
  assign y26678 = ~n35699 ;
  assign y26679 = ~n35704 ;
  assign y26680 = ~1'b0 ;
  assign y26681 = ~n6764 ;
  assign y26682 = ~1'b0 ;
  assign y26683 = ~n35705 ;
  assign y26684 = ~n35708 ;
  assign y26685 = ~n35709 ;
  assign y26686 = n10414 ;
  assign y26687 = ~1'b0 ;
  assign y26688 = n35711 ;
  assign y26689 = ~1'b0 ;
  assign y26690 = ~1'b0 ;
  assign y26691 = ~n35712 ;
  assign y26692 = ~1'b0 ;
  assign y26693 = n35714 ;
  assign y26694 = ~1'b0 ;
  assign y26695 = ~1'b0 ;
  assign y26696 = n35715 ;
  assign y26697 = n35716 ;
  assign y26698 = n8876 ;
  assign y26699 = ~n35717 ;
  assign y26700 = ~1'b0 ;
  assign y26701 = ~n15205 ;
  assign y26702 = n35719 ;
  assign y26703 = ~n1151 ;
  assign y26704 = ~1'b0 ;
  assign y26705 = ~n35722 ;
  assign y26706 = n35724 ;
  assign y26707 = ~1'b0 ;
  assign y26708 = ~1'b0 ;
  assign y26709 = n35728 ;
  assign y26710 = ~1'b0 ;
  assign y26711 = n35733 ;
  assign y26712 = ~n8227 ;
  assign y26713 = ~n13597 ;
  assign y26714 = n35737 ;
  assign y26715 = n35740 ;
  assign y26716 = ~n35741 ;
  assign y26717 = n68 ;
  assign y26718 = n35742 ;
  assign y26719 = n35743 ;
  assign y26720 = ~n35744 ;
  assign y26721 = ~n5832 ;
  assign y26722 = n35745 ;
  assign y26723 = n35747 ;
  assign y26724 = ~1'b0 ;
  assign y26725 = 1'b0 ;
  assign y26726 = 1'b0 ;
  assign y26727 = ~n35748 ;
  assign y26728 = n35751 ;
  assign y26729 = ~1'b0 ;
  assign y26730 = n35753 ;
  assign y26731 = n35758 ;
  assign y26732 = 1'b0 ;
  assign y26733 = ~n24825 ;
  assign y26734 = n35760 ;
  assign y26735 = ~n16490 ;
  assign y26736 = n35765 ;
  assign y26737 = ~1'b0 ;
  assign y26738 = ~n35766 ;
  assign y26739 = ~n35770 ;
  assign y26740 = n35771 ;
  assign y26741 = n35772 ;
  assign y26742 = n35773 ;
  assign y26743 = ~1'b0 ;
  assign y26744 = ~1'b0 ;
  assign y26745 = n35774 ;
  assign y26746 = n13679 ;
  assign y26747 = ~n35658 ;
  assign y26748 = n35776 ;
  assign y26749 = n35778 ;
  assign y26750 = ~1'b0 ;
  assign y26751 = n35779 ;
  assign y26752 = ~n35780 ;
  assign y26753 = ~1'b0 ;
  assign y26754 = n35783 ;
  assign y26755 = ~1'b0 ;
  assign y26756 = ~1'b0 ;
  assign y26757 = ~1'b0 ;
  assign y26758 = n35785 ;
  assign y26759 = n12694 ;
  assign y26760 = ~n539 ;
  assign y26761 = n35786 ;
  assign y26762 = ~1'b0 ;
  assign y26763 = ~n35788 ;
  assign y26764 = n29618 ;
  assign y26765 = ~n35789 ;
  assign y26766 = 1'b0 ;
  assign y26767 = ~1'b0 ;
  assign y26768 = ~1'b0 ;
  assign y26769 = ~1'b0 ;
  assign y26770 = ~1'b0 ;
  assign y26771 = n5836 ;
  assign y26772 = ~1'b0 ;
  assign y26773 = n35797 ;
  assign y26774 = ~1'b0 ;
  assign y26775 = n35798 ;
  assign y26776 = 1'b0 ;
  assign y26777 = ~n799 ;
  assign y26778 = n35800 ;
  assign y26779 = n2566 ;
  assign y26780 = ~1'b0 ;
  assign y26781 = n35802 ;
  assign y26782 = n26388 ;
  assign y26783 = ~1'b0 ;
  assign y26784 = n35804 ;
  assign y26785 = n35806 ;
  assign y26786 = ~n10580 ;
  assign y26787 = ~n35813 ;
  assign y26788 = ~n35814 ;
  assign y26789 = ~n35815 ;
  assign y26790 = ~1'b0 ;
  assign y26791 = ~1'b0 ;
  assign y26792 = n35817 ;
  assign y26793 = ~n35821 ;
  assign y26794 = n35822 ;
  assign y26795 = n35825 ;
  assign y26796 = ~1'b0 ;
  assign y26797 = ~1'b0 ;
  assign y26798 = ~n35826 ;
  assign y26799 = ~n35829 ;
  assign y26800 = ~n28775 ;
  assign y26801 = ~1'b0 ;
  assign y26802 = 1'b0 ;
  assign y26803 = n35830 ;
  assign y26804 = ~1'b0 ;
  assign y26805 = ~1'b0 ;
  assign y26806 = ~1'b0 ;
  assign y26807 = ~n35832 ;
  assign y26808 = ~1'b0 ;
  assign y26809 = n35834 ;
  assign y26810 = ~1'b0 ;
  assign y26811 = n290 ;
  assign y26812 = ~1'b0 ;
  assign y26813 = ~1'b0 ;
  assign y26814 = n35835 ;
  assign y26815 = ~n5258 ;
  assign y26816 = n35836 ;
  assign y26817 = ~1'b0 ;
  assign y26818 = ~n35841 ;
  assign y26819 = n35843 ;
  assign y26820 = n35844 ;
  assign y26821 = ~n35845 ;
  assign y26822 = n35849 ;
  assign y26823 = ~n35850 ;
  assign y26824 = ~n35852 ;
  assign y26825 = ~1'b0 ;
  assign y26826 = ~n27139 ;
  assign y26827 = ~n35853 ;
  assign y26828 = ~1'b0 ;
  assign y26829 = ~n263 ;
  assign y26830 = n35854 ;
  assign y26831 = 1'b0 ;
  assign y26832 = ~1'b0 ;
  assign y26833 = ~n35855 ;
  assign y26834 = n35857 ;
  assign y26835 = ~n35858 ;
  assign y26836 = ~n35154 ;
  assign y26837 = n35859 ;
  assign y26838 = ~n35863 ;
  assign y26839 = n35864 ;
  assign y26840 = ~n35865 ;
  assign y26841 = ~1'b0 ;
  assign y26842 = ~n35866 ;
  assign y26843 = ~1'b0 ;
  assign y26844 = 1'b0 ;
  assign y26845 = ~n13261 ;
  assign y26846 = n35867 ;
  assign y26847 = n35869 ;
  assign y26848 = ~1'b0 ;
  assign y26849 = ~1'b0 ;
  assign y26850 = n35871 ;
  assign y26851 = ~1'b0 ;
  assign y26852 = ~n35873 ;
  assign y26853 = ~n35877 ;
  assign y26854 = n1054 ;
  assign y26855 = ~n35878 ;
  assign y26856 = ~n35881 ;
  assign y26857 = 1'b0 ;
  assign y26858 = ~n35884 ;
  assign y26859 = ~n35886 ;
  assign y26860 = n35888 ;
  assign y26861 = ~1'b0 ;
  assign y26862 = ~1'b0 ;
  assign y26863 = ~1'b0 ;
  assign y26864 = ~1'b0 ;
  assign y26865 = n35890 ;
  assign y26866 = ~n35894 ;
  assign y26867 = ~1'b0 ;
  assign y26868 = ~1'b0 ;
  assign y26869 = ~1'b0 ;
  assign y26870 = n35895 ;
  assign y26871 = n16182 ;
  assign y26872 = n35897 ;
  assign y26873 = ~1'b0 ;
  assign y26874 = ~1'b0 ;
  assign y26875 = n35898 ;
  assign y26876 = n35900 ;
  assign y26877 = ~n35901 ;
  assign y26878 = 1'b0 ;
  assign y26879 = n35906 ;
  assign y26880 = ~1'b0 ;
  assign y26881 = ~n35907 ;
  assign y26882 = n35909 ;
  assign y26883 = ~n35913 ;
  assign y26884 = ~1'b0 ;
  assign y26885 = n35914 ;
  assign y26886 = ~n35916 ;
  assign y26887 = n35922 ;
  assign y26888 = ~1'b0 ;
  assign y26889 = ~n35923 ;
  assign y26890 = ~1'b0 ;
  assign y26891 = ~1'b0 ;
  assign y26892 = 1'b0 ;
  assign y26893 = 1'b0 ;
  assign y26894 = ~n35925 ;
  assign y26895 = n35926 ;
  assign y26896 = ~n35928 ;
  assign y26897 = ~n1992 ;
  assign y26898 = ~1'b0 ;
  assign y26899 = ~1'b0 ;
  assign y26900 = ~n35932 ;
  assign y26901 = n35936 ;
  assign y26902 = ~1'b0 ;
  assign y26903 = ~n35939 ;
  assign y26904 = ~1'b0 ;
  assign y26905 = ~1'b0 ;
  assign y26906 = ~1'b0 ;
  assign y26907 = n35940 ;
  assign y26908 = ~1'b0 ;
  assign y26909 = ~1'b0 ;
  assign y26910 = n35943 ;
  assign y26911 = ~1'b0 ;
  assign y26912 = ~1'b0 ;
  assign y26913 = ~1'b0 ;
  assign y26914 = n35945 ;
  assign y26915 = ~1'b0 ;
  assign y26916 = n35947 ;
  assign y26917 = n35948 ;
  assign y26918 = n35949 ;
  assign y26919 = ~n35951 ;
  assign y26920 = n374 ;
  assign y26921 = n35952 ;
  assign y26922 = ~1'b0 ;
  assign y26923 = ~1'b0 ;
  assign y26924 = ~n35954 ;
  assign y26925 = ~1'b0 ;
  assign y26926 = n738 ;
  assign y26927 = 1'b0 ;
  assign y26928 = n35972 ;
  assign y26929 = n35974 ;
  assign y26930 = 1'b0 ;
  assign y26931 = ~n30547 ;
  assign y26932 = ~n35976 ;
  assign y26933 = ~1'b0 ;
  assign y26934 = 1'b0 ;
  assign y26935 = ~1'b0 ;
  assign y26936 = ~1'b0 ;
  assign y26937 = ~1'b0 ;
  assign y26938 = ~1'b0 ;
  assign y26939 = ~n35977 ;
  assign y26940 = n35981 ;
  assign y26941 = ~n35982 ;
  assign y26942 = ~n35983 ;
  assign y26943 = ~1'b0 ;
  assign y26944 = ~1'b0 ;
  assign y26945 = ~1'b0 ;
  assign y26946 = n35986 ;
  assign y26947 = n35988 ;
  assign y26948 = n35991 ;
  assign y26949 = ~n35993 ;
  assign y26950 = ~1'b0 ;
  assign y26951 = n35997 ;
  assign y26952 = ~n35999 ;
  assign y26953 = ~1'b0 ;
  assign y26954 = n36001 ;
  assign y26955 = n36012 ;
  assign y26956 = n36015 ;
  assign y26957 = ~n36017 ;
  assign y26958 = n36019 ;
  assign y26959 = ~n36021 ;
  assign y26960 = ~1'b0 ;
  assign y26961 = n36027 ;
  assign y26962 = ~n36030 ;
  assign y26963 = ~1'b0 ;
  assign y26964 = ~n36031 ;
  assign y26965 = ~n36032 ;
  assign y26966 = ~1'b0 ;
  assign y26967 = ~n36035 ;
  assign y26968 = ~n36036 ;
  assign y26969 = ~1'b0 ;
  assign y26970 = 1'b0 ;
  assign y26971 = n23638 ;
  assign y26972 = ~n36038 ;
  assign y26973 = n36039 ;
  assign y26974 = ~n36040 ;
  assign y26975 = ~n36041 ;
  assign y26976 = ~1'b0 ;
  assign y26977 = ~1'b0 ;
  assign y26978 = 1'b0 ;
  assign y26979 = 1'b0 ;
  assign y26980 = ~n36045 ;
  assign y26981 = n36047 ;
  assign y26982 = ~n14181 ;
  assign y26983 = n36048 ;
  assign y26984 = n36051 ;
  assign y26985 = n181 ;
  assign y26986 = ~1'b0 ;
  assign y26987 = ~n36056 ;
  assign y26988 = 1'b0 ;
  assign y26989 = ~1'b0 ;
  assign y26990 = n36057 ;
  assign y26991 = ~n36059 ;
  assign y26992 = ~1'b0 ;
  assign y26993 = n36060 ;
  assign y26994 = ~n36062 ;
  assign y26995 = ~1'b0 ;
  assign y26996 = ~n25194 ;
  assign y26997 = ~1'b0 ;
  assign y26998 = n36064 ;
  assign y26999 = ~n36065 ;
  assign y27000 = ~1'b0 ;
  assign y27001 = n36069 ;
  assign y27002 = ~1'b0 ;
  assign y27003 = n36071 ;
  assign y27004 = ~1'b0 ;
  assign y27005 = ~1'b0 ;
  assign y27006 = ~1'b0 ;
  assign y27007 = ~1'b0 ;
  assign y27008 = n36072 ;
  assign y27009 = ~1'b0 ;
  assign y27010 = ~1'b0 ;
  assign y27011 = n36074 ;
  assign y27012 = ~n36077 ;
  assign y27013 = n36079 ;
  assign y27014 = ~n15875 ;
  assign y27015 = n36084 ;
  assign y27016 = n36087 ;
  assign y27017 = ~1'b0 ;
  assign y27018 = ~n36088 ;
  assign y27019 = n36094 ;
  assign y27020 = ~1'b0 ;
  assign y27021 = n89 ;
  assign y27022 = ~n36096 ;
  assign y27023 = n1048 ;
  assign y27024 = ~n4228 ;
  assign y27025 = n36097 ;
  assign y27026 = ~n2554 ;
  assign y27027 = ~n28992 ;
  assign y27028 = ~n26295 ;
  assign y27029 = ~n36099 ;
  assign y27030 = 1'b0 ;
  assign y27031 = ~n36101 ;
  assign y27032 = ~n36102 ;
  assign y27033 = ~n36103 ;
  assign y27034 = ~n36104 ;
  assign y27035 = n36109 ;
  assign y27036 = ~1'b0 ;
  assign y27037 = n36112 ;
  assign y27038 = n36114 ;
  assign y27039 = ~1'b0 ;
  assign y27040 = ~n36115 ;
  assign y27041 = n36127 ;
  assign y27042 = ~1'b0 ;
  assign y27043 = n36133 ;
  assign y27044 = ~1'b0 ;
  assign y27045 = n36135 ;
  assign y27046 = n36136 ;
  assign y27047 = n36137 ;
  assign y27048 = ~1'b0 ;
  assign y27049 = n36141 ;
  assign y27050 = n1693 ;
  assign y27051 = ~n36144 ;
  assign y27052 = 1'b0 ;
  assign y27053 = n36146 ;
  assign y27054 = ~n36147 ;
  assign y27055 = n36149 ;
  assign y27056 = ~1'b0 ;
  assign y27057 = n19884 ;
  assign y27058 = ~n36151 ;
  assign y27059 = n13386 ;
  assign y27060 = ~1'b0 ;
  assign y27061 = ~1'b0 ;
  assign y27062 = n6847 ;
  assign y27063 = n10059 ;
  assign y27064 = ~n36155 ;
  assign y27065 = n36183 ;
  assign y27066 = ~1'b0 ;
  assign y27067 = ~1'b0 ;
  assign y27068 = n36184 ;
  assign y27069 = ~n36185 ;
  assign y27070 = n36190 ;
  assign y27071 = ~n36193 ;
  assign y27072 = ~1'b0 ;
  assign y27073 = n36195 ;
  assign y27074 = ~1'b0 ;
  assign y27075 = n36196 ;
  assign y27076 = n8248 ;
  assign y27077 = n36198 ;
  assign y27078 = ~n36199 ;
  assign y27079 = ~n36200 ;
  assign y27080 = ~n36204 ;
  assign y27081 = ~1'b0 ;
  assign y27082 = n36205 ;
  assign y27083 = ~1'b0 ;
  assign y27084 = n36206 ;
  assign y27085 = ~1'b0 ;
  assign y27086 = ~n36208 ;
  assign y27087 = ~1'b0 ;
  assign y27088 = ~n36209 ;
  assign y27089 = n36210 ;
  assign y27090 = ~n36212 ;
  assign y27091 = n36213 ;
  assign y27092 = n36215 ;
  assign y27093 = ~1'b0 ;
  assign y27094 = ~1'b0 ;
  assign y27095 = ~1'b0 ;
  assign y27096 = n36219 ;
  assign y27097 = ~n36223 ;
  assign y27098 = ~n36225 ;
  assign y27099 = ~1'b0 ;
  assign y27100 = ~n23854 ;
  assign y27101 = ~n36227 ;
  assign y27102 = ~1'b0 ;
  assign y27103 = n36234 ;
  assign y27104 = n17632 ;
  assign y27105 = ~1'b0 ;
  assign y27106 = n36236 ;
  assign y27107 = ~n36240 ;
  assign y27108 = n36241 ;
  assign y27109 = ~n36243 ;
  assign y27110 = ~1'b0 ;
  assign y27111 = ~1'b0 ;
  assign y27112 = n36244 ;
  assign y27113 = n36245 ;
  assign y27114 = n36247 ;
  assign y27115 = ~1'b0 ;
  assign y27116 = n36252 ;
  assign y27117 = ~n36253 ;
  assign y27118 = ~n4163 ;
  assign y27119 = ~1'b0 ;
  assign y27120 = ~1'b0 ;
  assign y27121 = ~n36254 ;
  assign y27122 = n36255 ;
  assign y27123 = ~n36257 ;
  assign y27124 = ~1'b0 ;
  assign y27125 = 1'b0 ;
  assign y27126 = 1'b0 ;
  assign y27127 = n36258 ;
  assign y27128 = n36261 ;
  assign y27129 = ~n36263 ;
  assign y27130 = ~n36264 ;
  assign y27131 = n36266 ;
  assign y27132 = n36269 ;
  assign y27133 = ~1'b0 ;
  assign y27134 = ~n36270 ;
  assign y27135 = ~n36273 ;
  assign y27136 = n36274 ;
  assign y27137 = ~n36276 ;
  assign y27138 = ~n36281 ;
  assign y27139 = ~1'b0 ;
  assign y27140 = 1'b0 ;
  assign y27141 = n36284 ;
  assign y27142 = ~n36287 ;
  assign y27143 = ~1'b0 ;
  assign y27144 = ~n36288 ;
  assign y27145 = ~1'b0 ;
  assign y27146 = ~1'b0 ;
  assign y27147 = n36292 ;
  assign y27148 = ~1'b0 ;
  assign y27149 = ~1'b0 ;
  assign y27150 = n10395 ;
  assign y27151 = n36293 ;
  assign y27152 = n457 ;
  assign y27153 = ~n2604 ;
  assign y27154 = n36295 ;
  assign y27155 = ~n16482 ;
  assign y27156 = 1'b0 ;
  assign y27157 = ~1'b0 ;
  assign y27158 = ~1'b0 ;
  assign y27159 = ~1'b0 ;
  assign y27160 = n17598 ;
  assign y27161 = ~n36300 ;
  assign y27162 = n24640 ;
  assign y27163 = ~1'b0 ;
  assign y27164 = ~n36303 ;
  assign y27165 = ~1'b0 ;
  assign y27166 = n36305 ;
  assign y27167 = ~1'b0 ;
  assign y27168 = n36306 ;
  assign y27169 = ~n36308 ;
  assign y27170 = ~n36309 ;
  assign y27171 = ~n36310 ;
  assign y27172 = 1'b0 ;
  assign y27173 = ~n1811 ;
  assign y27174 = ~1'b0 ;
  assign y27175 = n36311 ;
  assign y27176 = n36312 ;
  assign y27177 = n36313 ;
  assign y27178 = ~n36315 ;
  assign y27179 = 1'b0 ;
  assign y27180 = n36316 ;
  assign y27181 = ~n8080 ;
  assign y27182 = ~1'b0 ;
  assign y27183 = ~n36318 ;
  assign y27184 = ~1'b0 ;
  assign y27185 = n36320 ;
  assign y27186 = ~n36323 ;
  assign y27187 = ~1'b0 ;
  assign y27188 = ~1'b0 ;
  assign y27189 = n36326 ;
  assign y27190 = ~1'b0 ;
  assign y27191 = 1'b0 ;
  assign y27192 = ~n36328 ;
  assign y27193 = ~n36330 ;
  assign y27194 = ~1'b0 ;
  assign y27195 = 1'b0 ;
  assign y27196 = ~n36333 ;
  assign y27197 = n36335 ;
  assign y27198 = ~1'b0 ;
  assign y27199 = ~n36336 ;
  assign y27200 = n12768 ;
  assign y27201 = ~n36337 ;
  assign y27202 = n36338 ;
  assign y27203 = n36339 ;
  assign y27204 = ~1'b0 ;
  assign y27205 = n36341 ;
  assign y27206 = ~1'b0 ;
  assign y27207 = ~n36342 ;
  assign y27208 = ~n4446 ;
  assign y27209 = ~n36343 ;
  assign y27210 = ~n36345 ;
  assign y27211 = ~1'b0 ;
  assign y27212 = ~n36347 ;
  assign y27213 = ~1'b0 ;
  assign y27214 = ~1'b0 ;
  assign y27215 = ~1'b0 ;
  assign y27216 = n36350 ;
  assign y27217 = ~n25674 ;
  assign y27218 = ~n36352 ;
  assign y27219 = ~n3411 ;
  assign y27220 = ~n20100 ;
  assign y27221 = ~n36353 ;
  assign y27222 = ~n36356 ;
  assign y27223 = n16979 ;
  assign y27224 = ~1'b0 ;
  assign y27225 = ~1'b0 ;
  assign y27226 = ~n36357 ;
  assign y27227 = ~n36358 ;
  assign y27228 = ~n8320 ;
  assign y27229 = n19938 ;
  assign y27230 = ~1'b0 ;
  assign y27231 = ~1'b0 ;
  assign y27232 = ~n36359 ;
  assign y27233 = ~n36363 ;
  assign y27234 = ~1'b0 ;
  assign y27235 = ~1'b0 ;
  assign y27236 = n36364 ;
  assign y27237 = ~n36366 ;
  assign y27238 = n36368 ;
  assign y27239 = ~1'b0 ;
  assign y27240 = 1'b0 ;
  assign y27241 = n36373 ;
  assign y27242 = 1'b0 ;
  assign y27243 = ~n36374 ;
  assign y27244 = 1'b0 ;
  assign y27245 = n36375 ;
  assign y27246 = ~n36376 ;
  assign y27247 = ~n36378 ;
  assign y27248 = ~1'b0 ;
  assign y27249 = ~1'b0 ;
  assign y27250 = ~n36379 ;
  assign y27251 = n36380 ;
  assign y27252 = ~n7701 ;
  assign y27253 = ~n36382 ;
  assign y27254 = ~n2244 ;
  assign y27255 = n36383 ;
  assign y27256 = ~1'b0 ;
  assign y27257 = n4927 ;
  assign y27258 = n28513 ;
  assign y27259 = ~1'b0 ;
  assign y27260 = ~1'b0 ;
  assign y27261 = ~1'b0 ;
  assign y27262 = n36385 ;
  assign y27263 = ~1'b0 ;
  assign y27264 = n33461 ;
  assign y27265 = ~1'b0 ;
  assign y27266 = 1'b0 ;
  assign y27267 = ~1'b0 ;
  assign y27268 = ~n36386 ;
  assign y27269 = n36389 ;
  assign y27270 = n36391 ;
  assign y27271 = ~n36392 ;
  assign y27272 = ~n36396 ;
  assign y27273 = n36397 ;
  assign y27274 = ~n36406 ;
  assign y27275 = n36408 ;
  assign y27276 = ~1'b0 ;
  assign y27277 = ~n36409 ;
  assign y27278 = ~n36410 ;
  assign y27279 = n36415 ;
  assign y27280 = ~1'b0 ;
  assign y27281 = ~n36418 ;
  assign y27282 = ~1'b0 ;
  assign y27283 = n36419 ;
  assign y27284 = ~n36421 ;
  assign y27285 = ~1'b0 ;
  assign y27286 = n4501 ;
  assign y27287 = ~n36422 ;
  assign y27288 = ~1'b0 ;
  assign y27289 = n36423 ;
  assign y27290 = ~n36425 ;
  assign y27291 = ~1'b0 ;
  assign y27292 = ~n36428 ;
  assign y27293 = ~n36430 ;
  assign y27294 = ~1'b0 ;
  assign y27295 = ~n2366 ;
  assign y27296 = ~1'b0 ;
  assign y27297 = ~n36432 ;
  assign y27298 = ~1'b0 ;
  assign y27299 = ~n36433 ;
  assign y27300 = ~n36435 ;
  assign y27301 = n36440 ;
  assign y27302 = ~n36441 ;
  assign y27303 = 1'b0 ;
  assign y27304 = n36444 ;
  assign y27305 = ~n36447 ;
  assign y27306 = ~1'b0 ;
  assign y27307 = ~n36450 ;
  assign y27308 = ~n36451 ;
  assign y27309 = ~1'b0 ;
  assign y27310 = n36453 ;
  assign y27311 = ~1'b0 ;
  assign y27312 = ~1'b0 ;
  assign y27313 = ~1'b0 ;
  assign y27314 = n36456 ;
  assign y27315 = ~1'b0 ;
  assign y27316 = n36457 ;
  assign y27317 = ~1'b0 ;
  assign y27318 = ~1'b0 ;
  assign y27319 = 1'b0 ;
  assign y27320 = ~n36458 ;
  assign y27321 = 1'b0 ;
  assign y27322 = n36459 ;
  assign y27323 = ~1'b0 ;
  assign y27324 = n36460 ;
  assign y27325 = ~n36462 ;
  assign y27326 = ~1'b0 ;
  assign y27327 = n36465 ;
  assign y27328 = ~1'b0 ;
  assign y27329 = n36466 ;
  assign y27330 = ~1'b0 ;
  assign y27331 = ~1'b0 ;
  assign y27332 = n36467 ;
  assign y27333 = ~n36474 ;
  assign y27334 = 1'b0 ;
  assign y27335 = n36475 ;
  assign y27336 = ~n36476 ;
  assign y27337 = ~1'b0 ;
  assign y27338 = ~1'b0 ;
  assign y27339 = ~n36478 ;
  assign y27340 = ~n36481 ;
  assign y27341 = ~1'b0 ;
  assign y27342 = ~1'b0 ;
  assign y27343 = ~1'b0 ;
  assign y27344 = ~1'b0 ;
  assign y27345 = ~n36483 ;
  assign y27346 = n36484 ;
  assign y27347 = n36488 ;
  assign y27348 = ~1'b0 ;
  assign y27349 = n36493 ;
  assign y27350 = ~1'b0 ;
  assign y27351 = n1241 ;
  assign y27352 = ~n36494 ;
  assign y27353 = 1'b0 ;
  assign y27354 = n36496 ;
  assign y27355 = n36497 ;
  assign y27356 = ~1'b0 ;
  assign y27357 = ~1'b0 ;
  assign y27358 = ~n36498 ;
  assign y27359 = 1'b0 ;
  assign y27360 = ~n36501 ;
  assign y27361 = ~n8156 ;
  assign y27362 = ~1'b0 ;
  assign y27363 = ~1'b0 ;
  assign y27364 = ~n36505 ;
  assign y27365 = ~1'b0 ;
  assign y27366 = ~n36506 ;
  assign y27367 = n36511 ;
  assign y27368 = ~1'b0 ;
  assign y27369 = n36515 ;
  assign y27370 = ~n36517 ;
  assign y27371 = ~n36519 ;
  assign y27372 = ~1'b0 ;
  assign y27373 = ~1'b0 ;
  assign y27374 = n36522 ;
  assign y27375 = n36523 ;
  assign y27376 = n36524 ;
  assign y27377 = n36526 ;
  assign y27378 = ~n36531 ;
  assign y27379 = ~n36533 ;
  assign y27380 = ~1'b0 ;
  assign y27381 = 1'b0 ;
  assign y27382 = ~1'b0 ;
  assign y27383 = ~1'b0 ;
  assign y27384 = n5338 ;
  assign y27385 = n36534 ;
  assign y27386 = ~1'b0 ;
  assign y27387 = ~1'b0 ;
  assign y27388 = n36536 ;
  assign y27389 = ~1'b0 ;
  assign y27390 = ~1'b0 ;
  assign y27391 = n21963 ;
  assign y27392 = ~n36537 ;
  assign y27393 = ~1'b0 ;
  assign y27394 = ~1'b0 ;
  assign y27395 = ~1'b0 ;
  assign y27396 = n16186 ;
  assign y27397 = n36539 ;
  assign y27398 = ~1'b0 ;
  assign y27399 = ~n36542 ;
  assign y27400 = n36547 ;
  assign y27401 = n36551 ;
  assign y27402 = ~n36554 ;
  assign y27403 = ~1'b0 ;
  assign y27404 = n8767 ;
  assign y27405 = ~1'b0 ;
  assign y27406 = ~n36555 ;
  assign y27407 = ~n36556 ;
  assign y27408 = ~n36557 ;
  assign y27409 = n36559 ;
  assign y27410 = ~n36562 ;
  assign y27411 = ~n21123 ;
  assign y27412 = ~1'b0 ;
  assign y27413 = n36566 ;
  assign y27414 = ~n6185 ;
  assign y27415 = ~1'b0 ;
  assign y27416 = ~n36567 ;
  assign y27417 = n36568 ;
  assign y27418 = ~1'b0 ;
  assign y27419 = ~n33253 ;
  assign y27420 = ~n36569 ;
  assign y27421 = ~n36571 ;
  assign y27422 = ~1'b0 ;
  assign y27423 = ~n36574 ;
  assign y27424 = ~1'b0 ;
  assign y27425 = ~n36575 ;
  assign y27426 = ~n15166 ;
  assign y27427 = ~1'b0 ;
  assign y27428 = ~n36577 ;
  assign y27429 = n36579 ;
  assign y27430 = ~1'b0 ;
  assign y27431 = ~1'b0 ;
  assign y27432 = ~1'b0 ;
  assign y27433 = ~n36581 ;
  assign y27434 = ~n36583 ;
  assign y27435 = ~n36585 ;
  assign y27436 = ~1'b0 ;
  assign y27437 = ~1'b0 ;
  assign y27438 = n36588 ;
  assign y27439 = ~1'b0 ;
  assign y27440 = ~1'b0 ;
  assign y27441 = n36590 ;
  assign y27442 = ~1'b0 ;
  assign y27443 = ~n36592 ;
  assign y27444 = ~n36599 ;
  assign y27445 = ~1'b0 ;
  assign y27446 = n36600 ;
  assign y27447 = ~1'b0 ;
  assign y27448 = ~1'b0 ;
  assign y27449 = ~n36602 ;
  assign y27450 = ~1'b0 ;
  assign y27451 = n36605 ;
  assign y27452 = ~1'b0 ;
  assign y27453 = ~n36606 ;
  assign y27454 = ~1'b0 ;
  assign y27455 = ~n36607 ;
  assign y27456 = ~1'b0 ;
  assign y27457 = ~1'b0 ;
  assign y27458 = 1'b0 ;
  assign y27459 = n36612 ;
  assign y27460 = ~1'b0 ;
  assign y27461 = n36617 ;
  assign y27462 = ~1'b0 ;
  assign y27463 = n36619 ;
  assign y27464 = ~1'b0 ;
  assign y27465 = ~1'b0 ;
  assign y27466 = ~n5701 ;
  assign y27467 = ~n36621 ;
  assign y27468 = ~n36623 ;
  assign y27469 = n36625 ;
  assign y27470 = ~n36628 ;
  assign y27471 = ~n36630 ;
  assign y27472 = ~n36632 ;
  assign y27473 = ~1'b0 ;
  assign y27474 = ~1'b0 ;
  assign y27475 = ~1'b0 ;
  assign y27476 = ~1'b0 ;
  assign y27477 = ~1'b0 ;
  assign y27478 = n36634 ;
  assign y27479 = ~n36635 ;
  assign y27480 = ~1'b0 ;
  assign y27481 = n36637 ;
  assign y27482 = ~1'b0 ;
  assign y27483 = ~1'b0 ;
  assign y27484 = ~1'b0 ;
  assign y27485 = ~1'b0 ;
  assign y27486 = ~1'b0 ;
  assign y27487 = ~n36640 ;
  assign y27488 = ~n36645 ;
  assign y27489 = ~n36647 ;
  assign y27490 = ~1'b0 ;
  assign y27491 = ~n4024 ;
  assign y27492 = ~n36649 ;
  assign y27493 = ~1'b0 ;
  assign y27494 = ~1'b0 ;
  assign y27495 = ~1'b0 ;
  assign y27496 = n36651 ;
  assign y27497 = n36652 ;
  assign y27498 = ~1'b0 ;
  assign y27499 = n36659 ;
  assign y27500 = ~1'b0 ;
  assign y27501 = n36660 ;
  assign y27502 = ~1'b0 ;
  assign y27503 = n36661 ;
  assign y27504 = n36665 ;
  assign y27505 = n36667 ;
  assign y27506 = n36672 ;
  assign y27507 = ~n36674 ;
  assign y27508 = n24366 ;
  assign y27509 = n36677 ;
  assign y27510 = ~n36680 ;
  assign y27511 = ~n36683 ;
  assign y27512 = ~1'b0 ;
  assign y27513 = ~n36684 ;
  assign y27514 = ~n23119 ;
  assign y27515 = n36686 ;
  assign y27516 = n36688 ;
  assign y27517 = ~n36689 ;
  assign y27518 = ~1'b0 ;
  assign y27519 = ~n36693 ;
  assign y27520 = ~1'b0 ;
  assign y27521 = 1'b0 ;
  assign y27522 = ~1'b0 ;
  assign y27523 = n36696 ;
  assign y27524 = ~n36701 ;
  assign y27525 = ~1'b0 ;
  assign y27526 = 1'b0 ;
  assign y27527 = n36703 ;
  assign y27528 = ~n36707 ;
  assign y27529 = ~n36708 ;
  assign y27530 = ~1'b0 ;
  assign y27531 = n36710 ;
  assign y27532 = ~1'b0 ;
  assign y27533 = n36713 ;
  assign y27534 = ~n36719 ;
  assign y27535 = ~1'b0 ;
  assign y27536 = ~1'b0 ;
  assign y27537 = ~1'b0 ;
  assign y27538 = n36721 ;
  assign y27539 = n36724 ;
  assign y27540 = ~1'b0 ;
  assign y27541 = ~n4560 ;
  assign y27542 = ~1'b0 ;
  assign y27543 = n36727 ;
  assign y27544 = ~n36731 ;
  assign y27545 = ~1'b0 ;
  assign y27546 = ~1'b0 ;
  assign y27547 = ~n36735 ;
  assign y27548 = ~n36736 ;
  assign y27549 = ~n36739 ;
  assign y27550 = n36740 ;
  assign y27551 = n36741 ;
  assign y27552 = n36746 ;
  assign y27553 = n36747 ;
  assign y27554 = n36751 ;
  assign y27555 = ~1'b0 ;
  assign y27556 = ~n36541 ;
  assign y27557 = n159 ;
  assign y27558 = ~n36752 ;
  assign y27559 = ~n36753 ;
  assign y27560 = ~1'b0 ;
  assign y27561 = ~1'b0 ;
  assign y27562 = n88 ;
  assign y27563 = n36754 ;
  assign y27564 = ~1'b0 ;
  assign y27565 = ~1'b0 ;
  assign y27566 = n36755 ;
  assign y27567 = ~1'b0 ;
  assign y27568 = ~n36757 ;
  assign y27569 = ~1'b0 ;
  assign y27570 = n2418 ;
  assign y27571 = n36760 ;
  assign y27572 = ~1'b0 ;
  assign y27573 = ~1'b0 ;
  assign y27574 = ~n36762 ;
  assign y27575 = ~1'b0 ;
  assign y27576 = n36764 ;
  assign y27577 = ~n36767 ;
  assign y27578 = ~n16368 ;
  assign y27579 = ~1'b0 ;
  assign y27580 = n29661 ;
  assign y27581 = ~1'b0 ;
  assign y27582 = n36771 ;
  assign y27583 = ~1'b0 ;
  assign y27584 = ~n36775 ;
  assign y27585 = ~n36778 ;
  assign y27586 = ~n36780 ;
  assign y27587 = n8446 ;
  assign y27588 = ~1'b0 ;
  assign y27589 = n36781 ;
  assign y27590 = ~1'b0 ;
  assign y27591 = n36782 ;
  assign y27592 = ~1'b0 ;
  assign y27593 = ~1'b0 ;
  assign y27594 = ~1'b0 ;
  assign y27595 = ~n36784 ;
  assign y27596 = 1'b0 ;
  assign y27597 = n36788 ;
  assign y27598 = ~1'b0 ;
  assign y27599 = n36791 ;
  assign y27600 = ~n36794 ;
  assign y27601 = ~1'b0 ;
  assign y27602 = ~1'b0 ;
  assign y27603 = ~n36796 ;
  assign y27604 = n2280 ;
  assign y27605 = ~1'b0 ;
  assign y27606 = ~n4790 ;
  assign y27607 = ~1'b0 ;
  assign y27608 = n36798 ;
  assign y27609 = n36803 ;
  assign y27610 = n13701 ;
  assign y27611 = ~n36805 ;
  assign y27612 = ~n33823 ;
  assign y27613 = n36806 ;
  assign y27614 = ~1'b0 ;
  assign y27615 = ~1'b0 ;
  assign y27616 = ~1'b0 ;
  assign y27617 = 1'b0 ;
  assign y27618 = ~1'b0 ;
  assign y27619 = ~1'b0 ;
  assign y27620 = n36807 ;
  assign y27621 = ~1'b0 ;
  assign y27622 = ~1'b0 ;
  assign y27623 = ~n36811 ;
  assign y27624 = ~1'b0 ;
  assign y27625 = n36812 ;
  assign y27626 = ~n36814 ;
  assign y27627 = n17092 ;
  assign y27628 = ~1'b0 ;
  assign y27629 = ~n36818 ;
  assign y27630 = ~n36820 ;
  assign y27631 = n1441 ;
  assign y27632 = n36821 ;
  assign y27633 = ~n36823 ;
  assign y27634 = ~1'b0 ;
  assign y27635 = n36825 ;
  assign y27636 = ~n5853 ;
  assign y27637 = ~1'b0 ;
  assign y27638 = ~1'b0 ;
  assign y27639 = ~1'b0 ;
  assign y27640 = ~1'b0 ;
  assign y27641 = ~n36826 ;
  assign y27642 = ~n6907 ;
  assign y27643 = n36827 ;
  assign y27644 = ~n36828 ;
  assign y27645 = ~1'b0 ;
  assign y27646 = ~1'b0 ;
  assign y27647 = ~n36829 ;
  assign y27648 = 1'b0 ;
  assign y27649 = ~1'b0 ;
  assign y27650 = n36830 ;
  assign y27651 = ~1'b0 ;
  assign y27652 = n36832 ;
  assign y27653 = n36835 ;
  assign y27654 = ~n36838 ;
  assign y27655 = n9483 ;
  assign y27656 = ~n36842 ;
  assign y27657 = ~n36843 ;
  assign y27658 = ~n36845 ;
  assign y27659 = ~n19910 ;
  assign y27660 = n708 ;
  assign y27661 = ~n36846 ;
  assign y27662 = n36849 ;
  assign y27663 = n36850 ;
  assign y27664 = ~1'b0 ;
  assign y27665 = ~1'b0 ;
  assign y27666 = ~1'b0 ;
  assign y27667 = ~n36851 ;
  assign y27668 = n36853 ;
  assign y27669 = n36854 ;
  assign y27670 = ~n5281 ;
  assign y27671 = n36857 ;
  assign y27672 = ~n36858 ;
  assign y27673 = ~1'b0 ;
  assign y27674 = ~1'b0 ;
  assign y27675 = n36859 ;
  assign y27676 = ~1'b0 ;
  assign y27677 = ~1'b0 ;
  assign y27678 = n5610 ;
  assign y27679 = ~n36860 ;
  assign y27680 = ~1'b0 ;
  assign y27681 = n36862 ;
  assign y27682 = n33933 ;
  assign y27683 = n36863 ;
  assign y27684 = n36864 ;
  assign y27685 = n36865 ;
  assign y27686 = ~n36866 ;
  assign y27687 = ~n36868 ;
  assign y27688 = ~n36870 ;
  assign y27689 = ~n36871 ;
  assign y27690 = ~1'b0 ;
  assign y27691 = n36874 ;
  assign y27692 = ~1'b0 ;
  assign y27693 = n36875 ;
  assign y27694 = ~1'b0 ;
  assign y27695 = ~1'b0 ;
  assign y27696 = ~1'b0 ;
  assign y27697 = ~n36876 ;
  assign y27698 = ~n36878 ;
  assign y27699 = n14450 ;
  assign y27700 = ~1'b0 ;
  assign y27701 = ~1'b0 ;
  assign y27702 = ~1'b0 ;
  assign y27703 = ~n36884 ;
  assign y27704 = ~n36885 ;
  assign y27705 = ~1'b0 ;
  assign y27706 = n36890 ;
  assign y27707 = n36892 ;
  assign y27708 = n36894 ;
  assign y27709 = 1'b0 ;
  assign y27710 = n18453 ;
  assign y27711 = ~n36898 ;
  assign y27712 = 1'b0 ;
  assign y27713 = ~1'b0 ;
  assign y27714 = n24228 ;
  assign y27715 = n36901 ;
  assign y27716 = ~n36903 ;
  assign y27717 = 1'b0 ;
  assign y27718 = ~1'b0 ;
  assign y27719 = n36905 ;
  assign y27720 = ~1'b0 ;
  assign y27721 = n36906 ;
  assign y27722 = ~n36907 ;
  assign y27723 = ~1'b0 ;
  assign y27724 = ~n36909 ;
  assign y27725 = ~n36925 ;
  assign y27726 = ~1'b0 ;
  assign y27727 = n36927 ;
  assign y27728 = n36935 ;
  assign y27729 = n36938 ;
  assign y27730 = n36940 ;
  assign y27731 = ~n32051 ;
  assign y27732 = n18717 ;
  assign y27733 = ~1'b0 ;
  assign y27734 = ~n36943 ;
  assign y27735 = ~1'b0 ;
  assign y27736 = n36945 ;
  assign y27737 = ~1'b0 ;
  assign y27738 = ~n36947 ;
  assign y27739 = n36948 ;
  assign y27740 = n36950 ;
  assign y27741 = ~1'b0 ;
  assign y27742 = n8341 ;
  assign y27743 = 1'b0 ;
  assign y27744 = n36952 ;
  assign y27745 = ~1'b0 ;
  assign y27746 = ~1'b0 ;
  assign y27747 = ~1'b0 ;
  assign y27748 = 1'b0 ;
  assign y27749 = n36953 ;
  assign y27750 = 1'b0 ;
  assign y27751 = ~n36954 ;
  assign y27752 = ~1'b0 ;
  assign y27753 = 1'b0 ;
  assign y27754 = ~1'b0 ;
  assign y27755 = n16288 ;
  assign y27756 = 1'b0 ;
  assign y27757 = n36955 ;
  assign y27758 = ~n36957 ;
  assign y27759 = ~n36958 ;
  assign y27760 = 1'b0 ;
  assign y27761 = n16938 ;
  assign y27762 = ~1'b0 ;
  assign y27763 = n36959 ;
  assign y27764 = n36963 ;
  assign y27765 = ~1'b0 ;
  assign y27766 = ~1'b0 ;
  assign y27767 = n36966 ;
  assign y27768 = ~n36968 ;
  assign y27769 = ~n36973 ;
  assign y27770 = ~n36974 ;
  assign y27771 = ~1'b0 ;
  assign y27772 = ~n36977 ;
  assign y27773 = ~n6929 ;
  assign y27774 = ~1'b0 ;
  assign y27775 = ~1'b0 ;
  assign y27776 = n36983 ;
  assign y27777 = ~1'b0 ;
  assign y27778 = ~n36986 ;
  assign y27779 = n36988 ;
  assign y27780 = n36989 ;
  assign y27781 = ~n36994 ;
  assign y27782 = n36999 ;
  assign y27783 = ~1'b0 ;
  assign y27784 = ~1'b0 ;
  assign y27785 = n37000 ;
  assign y27786 = ~1'b0 ;
  assign y27787 = ~1'b0 ;
  assign y27788 = 1'b0 ;
  assign y27789 = n37001 ;
  assign y27790 = n37007 ;
  assign y27791 = ~n37008 ;
  assign y27792 = ~n37011 ;
  assign y27793 = ~1'b0 ;
  assign y27794 = n37013 ;
  assign y27795 = ~1'b0 ;
  assign y27796 = ~n37016 ;
  assign y27797 = n14381 ;
  assign y27798 = ~n37023 ;
  assign y27799 = n37026 ;
  assign y27800 = ~n37028 ;
  assign y27801 = ~n37029 ;
  assign y27802 = n37031 ;
  assign y27803 = n37032 ;
  assign y27804 = n37033 ;
  assign y27805 = n37035 ;
  assign y27806 = ~n37037 ;
  assign y27807 = ~1'b0 ;
  assign y27808 = n37041 ;
  assign y27809 = n37043 ;
  assign y27810 = ~1'b0 ;
  assign y27811 = ~n37044 ;
  assign y27812 = ~n37046 ;
  assign y27813 = n1401 ;
  assign y27814 = ~1'b0 ;
  assign y27815 = ~1'b0 ;
  assign y27816 = ~n37050 ;
  assign y27817 = ~n30686 ;
  assign y27818 = ~n37056 ;
  assign y27819 = ~n1070 ;
  assign y27820 = 1'b0 ;
  assign y27821 = ~1'b0 ;
  assign y27822 = n37058 ;
  assign y27823 = ~1'b0 ;
  assign y27824 = ~1'b0 ;
  assign y27825 = ~1'b0 ;
  assign y27826 = ~n37061 ;
  assign y27827 = ~n37062 ;
  assign y27828 = ~1'b0 ;
  assign y27829 = n37064 ;
  assign y27830 = ~n37065 ;
  assign y27831 = ~n37074 ;
  assign y27832 = 1'b0 ;
  assign y27833 = ~1'b0 ;
  assign y27834 = ~1'b0 ;
  assign y27835 = 1'b0 ;
  assign y27836 = ~1'b0 ;
  assign y27837 = ~n37075 ;
  assign y27838 = ~n37078 ;
  assign y27839 = n37080 ;
  assign y27840 = n37081 ;
  assign y27841 = ~n6955 ;
  assign y27842 = n37082 ;
  assign y27843 = n37083 ;
  assign y27844 = n599 ;
  assign y27845 = ~1'b0 ;
  assign y27846 = n8706 ;
  assign y27847 = ~n31167 ;
  assign y27848 = ~1'b0 ;
  assign y27849 = ~n37084 ;
  assign y27850 = n37085 ;
  assign y27851 = ~1'b0 ;
  assign y27852 = ~1'b0 ;
  assign y27853 = ~1'b0 ;
  assign y27854 = ~1'b0 ;
  assign y27855 = ~1'b0 ;
  assign y27856 = n37086 ;
  assign y27857 = ~n37088 ;
  assign y27858 = ~1'b0 ;
  assign y27859 = n37089 ;
  assign y27860 = ~n37092 ;
  assign y27861 = ~n23718 ;
  assign y27862 = ~n1883 ;
  assign y27863 = ~n37095 ;
  assign y27864 = ~1'b0 ;
  assign y27865 = n37098 ;
  assign y27866 = ~n37099 ;
  assign y27867 = n37107 ;
  assign y27868 = ~1'b0 ;
  assign y27869 = ~n2136 ;
  assign y27870 = ~n37111 ;
  assign y27871 = ~1'b0 ;
  assign y27872 = ~n37119 ;
  assign y27873 = n37120 ;
  assign y27874 = ~1'b0 ;
  assign y27875 = n37123 ;
  assign y27876 = ~n37124 ;
  assign y27877 = n37126 ;
  assign y27878 = ~n1447 ;
  assign y27879 = ~1'b0 ;
  assign y27880 = ~n37128 ;
  assign y27881 = ~1'b0 ;
  assign y27882 = ~1'b0 ;
  assign y27883 = n37129 ;
  assign y27884 = ~n37132 ;
  assign y27885 = ~1'b0 ;
  assign y27886 = ~1'b0 ;
  assign y27887 = ~1'b0 ;
  assign y27888 = ~1'b0 ;
  assign y27889 = n37137 ;
  assign y27890 = ~1'b0 ;
  assign y27891 = n27582 ;
  assign y27892 = ~1'b0 ;
  assign y27893 = ~1'b0 ;
  assign y27894 = 1'b0 ;
  assign y27895 = ~n37141 ;
  assign y27896 = n37143 ;
  assign y27897 = n36529 ;
  assign y27898 = ~1'b0 ;
  assign y27899 = ~1'b0 ;
  assign y27900 = n37149 ;
  assign y27901 = n37150 ;
  assign y27902 = n2269 ;
  assign y27903 = ~n37151 ;
  assign y27904 = ~n26003 ;
  assign y27905 = ~1'b0 ;
  assign y27906 = n37153 ;
  assign y27907 = ~1'b0 ;
  assign y27908 = n37154 ;
  assign y27909 = ~1'b0 ;
  assign y27910 = n37155 ;
  assign y27911 = n37158 ;
  assign y27912 = ~1'b0 ;
  assign y27913 = ~n37161 ;
  assign y27914 = 1'b0 ;
  assign y27915 = ~n37163 ;
  assign y27916 = ~n37165 ;
  assign y27917 = ~1'b0 ;
  assign y27918 = ~1'b0 ;
  assign y27919 = ~1'b0 ;
  assign y27920 = n37170 ;
  assign y27921 = ~n37171 ;
  assign y27922 = ~1'b0 ;
  assign y27923 = ~n37172 ;
  assign y27924 = ~1'b0 ;
  assign y27925 = ~n133 ;
  assign y27926 = ~1'b0 ;
  assign y27927 = ~n37173 ;
  assign y27928 = n37175 ;
  assign y27929 = ~1'b0 ;
  assign y27930 = n10638 ;
  assign y27931 = n37176 ;
  assign y27932 = ~1'b0 ;
  assign y27933 = n37177 ;
  assign y27934 = n37180 ;
  assign y27935 = ~1'b0 ;
  assign y27936 = ~1'b0 ;
  assign y27937 = 1'b0 ;
  assign y27938 = ~1'b0 ;
  assign y27939 = ~1'b0 ;
  assign y27940 = n37181 ;
  assign y27941 = ~n37183 ;
  assign y27942 = ~1'b0 ;
  assign y27943 = 1'b0 ;
  assign y27944 = ~n37189 ;
  assign y27945 = ~1'b0 ;
  assign y27946 = n37190 ;
  assign y27947 = ~n37192 ;
  assign y27948 = ~n37195 ;
  assign y27949 = n5660 ;
  assign y27950 = n20101 ;
  assign y27951 = ~1'b0 ;
  assign y27952 = n37200 ;
  assign y27953 = n37201 ;
  assign y27954 = ~1'b0 ;
  assign y27955 = n37202 ;
  assign y27956 = ~1'b0 ;
  assign y27957 = ~1'b0 ;
  assign y27958 = n37203 ;
  assign y27959 = ~1'b0 ;
  assign y27960 = ~n37204 ;
  assign y27961 = ~n4952 ;
  assign y27962 = ~n37207 ;
  assign y27963 = ~n37208 ;
  assign y27964 = ~1'b0 ;
  assign y27965 = ~n37212 ;
  assign y27966 = n37214 ;
  assign y27967 = ~1'b0 ;
  assign y27968 = n37216 ;
  assign y27969 = ~1'b0 ;
  assign y27970 = ~1'b0 ;
  assign y27971 = n37219 ;
  assign y27972 = 1'b0 ;
  assign y27973 = ~1'b0 ;
  assign y27974 = ~n37222 ;
  assign y27975 = ~n37223 ;
  assign y27976 = ~n37226 ;
  assign y27977 = ~1'b0 ;
  assign y27978 = ~1'b0 ;
  assign y27979 = ~n30687 ;
  assign y27980 = ~n37227 ;
  assign y27981 = n37233 ;
  assign y27982 = ~n37234 ;
  assign y27983 = ~1'b0 ;
  assign y27984 = ~1'b0 ;
  assign y27985 = ~n37236 ;
  assign y27986 = ~n37237 ;
  assign y27987 = 1'b0 ;
  assign y27988 = ~1'b0 ;
  assign y27989 = ~1'b0 ;
  assign y27990 = n37239 ;
  assign y27991 = ~1'b0 ;
  assign y27992 = ~n37240 ;
  assign y27993 = ~n27302 ;
  assign y27994 = n37243 ;
  assign y27995 = ~n37246 ;
  assign y27996 = ~n18417 ;
  assign y27997 = ~1'b0 ;
  assign y27998 = ~1'b0 ;
  assign y27999 = 1'b0 ;
  assign y28000 = ~1'b0 ;
  assign y28001 = n37248 ;
  assign y28002 = n37249 ;
  assign y28003 = ~1'b0 ;
  assign y28004 = ~1'b0 ;
  assign y28005 = ~n37251 ;
  assign y28006 = ~1'b0 ;
  assign y28007 = ~n37255 ;
  assign y28008 = ~n37259 ;
  assign y28009 = ~1'b0 ;
  assign y28010 = ~1'b0 ;
  assign y28011 = ~1'b0 ;
  assign y28012 = ~n37263 ;
  assign y28013 = n37268 ;
  assign y28014 = ~n37269 ;
  assign y28015 = ~n35297 ;
  assign y28016 = n6254 ;
  assign y28017 = ~1'b0 ;
  assign y28018 = ~1'b0 ;
  assign y28019 = n37272 ;
  assign y28020 = ~1'b0 ;
  assign y28021 = n37273 ;
  assign y28022 = ~1'b0 ;
  assign y28023 = ~n37274 ;
  assign y28024 = ~n37276 ;
  assign y28025 = ~1'b0 ;
  assign y28026 = 1'b0 ;
  assign y28027 = n37277 ;
  assign y28028 = ~1'b0 ;
  assign y28029 = ~1'b0 ;
  assign y28030 = ~1'b0 ;
  assign y28031 = n37280 ;
  assign y28032 = n37283 ;
  assign y28033 = ~1'b0 ;
  assign y28034 = n37284 ;
  assign y28035 = n37288 ;
  assign y28036 = ~1'b0 ;
  assign y28037 = ~n37289 ;
  assign y28038 = ~1'b0 ;
  assign y28039 = ~1'b0 ;
  assign y28040 = ~1'b0 ;
  assign y28041 = ~1'b0 ;
  assign y28042 = ~n37296 ;
  assign y28043 = n37297 ;
  assign y28044 = n37299 ;
  assign y28045 = ~n37302 ;
  assign y28046 = ~1'b0 ;
  assign y28047 = ~n37306 ;
  assign y28048 = ~1'b0 ;
  assign y28049 = ~1'b0 ;
  assign y28050 = ~1'b0 ;
  assign y28051 = ~1'b0 ;
  assign y28052 = ~n37309 ;
  assign y28053 = ~n37311 ;
  assign y28054 = ~n37313 ;
  assign y28055 = ~1'b0 ;
  assign y28056 = ~1'b0 ;
  assign y28057 = ~n37314 ;
  assign y28058 = ~n37318 ;
  assign y28059 = ~1'b0 ;
  assign y28060 = ~n37322 ;
  assign y28061 = ~1'b0 ;
  assign y28062 = n37323 ;
  assign y28063 = ~1'b0 ;
  assign y28064 = ~n37326 ;
  assign y28065 = ~n37327 ;
  assign y28066 = ~1'b0 ;
  assign y28067 = ~n37328 ;
  assign y28068 = ~n37334 ;
  assign y28069 = ~n37336 ;
  assign y28070 = ~1'b0 ;
  assign y28071 = n37338 ;
  assign y28072 = ~n37339 ;
  assign y28073 = ~1'b0 ;
  assign y28074 = ~1'b0 ;
  assign y28075 = ~n37341 ;
  assign y28076 = ~1'b0 ;
  assign y28077 = 1'b0 ;
  assign y28078 = ~1'b0 ;
  assign y28079 = ~1'b0 ;
  assign y28080 = ~n37343 ;
  assign y28081 = ~n37349 ;
  assign y28082 = ~1'b0 ;
  assign y28083 = ~n37350 ;
  assign y28084 = ~1'b0 ;
  assign y28085 = 1'b0 ;
  assign y28086 = ~1'b0 ;
  assign y28087 = ~n37351 ;
  assign y28088 = ~1'b0 ;
  assign y28089 = ~n37353 ;
  assign y28090 = ~n37354 ;
  assign y28091 = n37356 ;
  assign y28092 = n28938 ;
  assign y28093 = ~n37358 ;
  assign y28094 = n37361 ;
  assign y28095 = 1'b0 ;
  assign y28096 = ~1'b0 ;
  assign y28097 = ~1'b0 ;
  assign y28098 = n37362 ;
  assign y28099 = ~1'b0 ;
  assign y28100 = n37364 ;
  assign y28101 = 1'b0 ;
  assign y28102 = ~n37365 ;
  assign y28103 = n37367 ;
  assign y28104 = ~n3193 ;
  assign y28105 = ~1'b0 ;
  assign y28106 = ~1'b0 ;
  assign y28107 = ~1'b0 ;
  assign y28108 = n37370 ;
  assign y28109 = n37374 ;
  assign y28110 = ~n37376 ;
  assign y28111 = ~1'b0 ;
  assign y28112 = ~1'b0 ;
  assign y28113 = ~n382 ;
  assign y28114 = ~n37378 ;
  assign y28115 = ~n17176 ;
  assign y28116 = n37382 ;
  assign y28117 = ~1'b0 ;
  assign y28118 = n37384 ;
  assign y28119 = n37387 ;
  assign y28120 = n37388 ;
  assign y28121 = ~1'b0 ;
  assign y28122 = ~n37391 ;
  assign y28123 = ~n37396 ;
  assign y28124 = n37397 ;
  assign y28125 = ~1'b0 ;
  assign y28126 = ~1'b0 ;
  assign y28127 = ~n37398 ;
  assign y28128 = ~n24451 ;
  assign y28129 = 1'b0 ;
  assign y28130 = n3361 ;
  assign y28131 = ~1'b0 ;
  assign y28132 = n37400 ;
  assign y28133 = ~1'b0 ;
  assign y28134 = ~1'b0 ;
  assign y28135 = n37402 ;
  assign y28136 = ~1'b0 ;
  assign y28137 = ~1'b0 ;
  assign y28138 = n37405 ;
  assign y28139 = ~1'b0 ;
  assign y28140 = n37408 ;
  assign y28141 = n37414 ;
  assign y28142 = ~n37416 ;
  assign y28143 = ~1'b0 ;
  assign y28144 = n37422 ;
  assign y28145 = ~1'b0 ;
  assign y28146 = ~1'b0 ;
  assign y28147 = ~1'b0 ;
  assign y28148 = n37428 ;
  assign y28149 = ~n37434 ;
  assign y28150 = 1'b0 ;
  assign y28151 = n37435 ;
  assign y28152 = ~1'b0 ;
  assign y28153 = 1'b0 ;
  assign y28154 = ~n37436 ;
  assign y28155 = n37438 ;
  assign y28156 = ~n164 ;
  assign y28157 = ~1'b0 ;
  assign y28158 = ~n37440 ;
  assign y28159 = n37444 ;
  assign y28160 = n37446 ;
  assign y28161 = ~1'b0 ;
  assign y28162 = ~n37448 ;
  assign y28163 = ~n37449 ;
  assign y28164 = ~1'b0 ;
  assign y28165 = n37451 ;
  assign y28166 = ~n37452 ;
  assign y28167 = n37455 ;
  assign y28168 = ~1'b0 ;
  assign y28169 = ~1'b0 ;
  assign y28170 = ~n37456 ;
  assign y28171 = n37457 ;
  assign y28172 = ~1'b0 ;
  assign y28173 = n37458 ;
  assign y28174 = ~n37463 ;
  assign y28175 = n37464 ;
  assign y28176 = n37466 ;
  assign y28177 = ~n37467 ;
  assign y28178 = ~1'b0 ;
  assign y28179 = n37469 ;
  assign y28180 = n37470 ;
  assign y28181 = ~n37476 ;
  assign y28182 = ~1'b0 ;
  assign y28183 = ~n37483 ;
  assign y28184 = n5632 ;
  assign y28185 = n37485 ;
  assign y28186 = ~1'b0 ;
  assign y28187 = ~n37486 ;
  assign y28188 = ~n19327 ;
  assign y28189 = ~1'b0 ;
  assign y28190 = ~n3670 ;
  assign y28191 = n37489 ;
  assign y28192 = ~1'b0 ;
  assign y28193 = ~n24049 ;
  assign y28194 = 1'b0 ;
  assign y28195 = n37493 ;
  assign y28196 = 1'b0 ;
  assign y28197 = ~n37494 ;
  assign y28198 = ~1'b0 ;
  assign y28199 = ~1'b0 ;
  assign y28200 = ~1'b0 ;
  assign y28201 = ~1'b0 ;
  assign y28202 = ~1'b0 ;
  assign y28203 = ~n37495 ;
  assign y28204 = ~n18403 ;
  assign y28205 = 1'b0 ;
  assign y28206 = n37501 ;
  assign y28207 = n37508 ;
  assign y28208 = n37512 ;
  assign y28209 = n37514 ;
  assign y28210 = n37516 ;
  assign y28211 = ~n37519 ;
  assign y28212 = ~n37525 ;
  assign y28213 = n37527 ;
  assign y28214 = ~1'b0 ;
  assign y28215 = ~1'b0 ;
  assign y28216 = n37528 ;
  assign y28217 = n11915 ;
  assign y28218 = ~1'b0 ;
  assign y28219 = ~1'b0 ;
  assign y28220 = ~1'b0 ;
  assign y28221 = n37530 ;
  assign y28222 = ~1'b0 ;
  assign y28223 = ~n37533 ;
  assign y28224 = ~1'b0 ;
  assign y28225 = ~1'b0 ;
  assign y28226 = n685 ;
  assign y28227 = n37534 ;
  assign y28228 = n37535 ;
  assign y28229 = ~1'b0 ;
  assign y28230 = ~n37538 ;
  assign y28231 = n5537 ;
  assign y28232 = ~1'b0 ;
  assign y28233 = ~1'b0 ;
  assign y28234 = ~1'b0 ;
  assign y28235 = ~1'b0 ;
  assign y28236 = ~1'b0 ;
  assign y28237 = ~n37541 ;
  assign y28238 = ~1'b0 ;
  assign y28239 = ~1'b0 ;
  assign y28240 = ~1'b0 ;
  assign y28241 = ~n37542 ;
  assign y28242 = ~1'b0 ;
  assign y28243 = ~n37544 ;
  assign y28244 = n37546 ;
  assign y28245 = n37547 ;
  assign y28246 = ~1'b0 ;
  assign y28247 = ~1'b0 ;
  assign y28248 = ~n37549 ;
  assign y28249 = ~n5251 ;
  assign y28250 = 1'b0 ;
  assign y28251 = ~n37550 ;
  assign y28252 = ~n37554 ;
  assign y28253 = ~n11246 ;
  assign y28254 = 1'b0 ;
  assign y28255 = ~n37555 ;
  assign y28256 = ~n37559 ;
  assign y28257 = ~1'b0 ;
  assign y28258 = ~n37560 ;
  assign y28259 = n37565 ;
  assign y28260 = ~n37567 ;
  assign y28261 = ~n16972 ;
  assign y28262 = n37568 ;
  assign y28263 = ~n37570 ;
  assign y28264 = ~n37571 ;
  assign y28265 = ~n37572 ;
  assign y28266 = n37573 ;
  assign y28267 = ~1'b0 ;
  assign y28268 = ~1'b0 ;
  assign y28269 = ~1'b0 ;
  assign y28270 = ~1'b0 ;
  assign y28271 = n37576 ;
  assign y28272 = n37580 ;
  assign y28273 = ~1'b0 ;
  assign y28274 = ~1'b0 ;
  assign y28275 = n37583 ;
  assign y28276 = 1'b0 ;
  assign y28277 = ~1'b0 ;
  assign y28278 = n13327 ;
  assign y28279 = ~1'b0 ;
  assign y28280 = n37585 ;
  assign y28281 = ~1'b0 ;
  assign y28282 = ~n37587 ;
  assign y28283 = ~n37589 ;
  assign y28284 = n37592 ;
  assign y28285 = n37595 ;
  assign y28286 = ~1'b0 ;
  assign y28287 = ~1'b0 ;
  assign y28288 = ~1'b0 ;
  assign y28289 = ~1'b0 ;
  assign y28290 = n37598 ;
  assign y28291 = n37600 ;
  assign y28292 = n15912 ;
  assign y28293 = n37602 ;
  assign y28294 = 1'b0 ;
  assign y28295 = n37603 ;
  assign y28296 = ~n37605 ;
  assign y28297 = ~n37606 ;
  assign y28298 = n37607 ;
  assign y28299 = ~1'b0 ;
  assign y28300 = ~n37608 ;
  assign y28301 = ~n23376 ;
  assign y28302 = n2497 ;
  assign y28303 = ~n37610 ;
  assign y28304 = n37612 ;
  assign y28305 = ~1'b0 ;
  assign y28306 = ~1'b0 ;
  assign y28307 = ~n7460 ;
  assign y28308 = ~1'b0 ;
  assign y28309 = ~n37613 ;
  assign y28310 = 1'b0 ;
  assign y28311 = n37614 ;
  assign y28312 = ~1'b0 ;
  assign y28313 = n37616 ;
  assign y28314 = ~n37620 ;
  assign y28315 = ~1'b0 ;
  assign y28316 = n2830 ;
  assign y28317 = ~n37621 ;
  assign y28318 = n37627 ;
  assign y28319 = ~1'b0 ;
  assign y28320 = n37631 ;
  assign y28321 = n37632 ;
  assign y28322 = ~1'b0 ;
  assign y28323 = n37636 ;
  assign y28324 = ~n37638 ;
  assign y28325 = ~n37640 ;
  assign y28326 = n37641 ;
  assign y28327 = n24412 ;
  assign y28328 = 1'b0 ;
  assign y28329 = ~n37642 ;
  assign y28330 = ~n37645 ;
  assign y28331 = ~1'b0 ;
  assign y28332 = ~n37646 ;
  assign y28333 = ~1'b0 ;
  assign y28334 = n1531 ;
  assign y28335 = ~n37647 ;
  assign y28336 = ~n31196 ;
  assign y28337 = ~1'b0 ;
  assign y28338 = ~n37649 ;
  assign y28339 = ~1'b0 ;
  assign y28340 = ~1'b0 ;
  assign y28341 = ~n20330 ;
  assign y28342 = ~n37655 ;
  assign y28343 = ~1'b0 ;
  assign y28344 = n37657 ;
  assign y28345 = ~n37658 ;
  assign y28346 = n37659 ;
  assign y28347 = n37661 ;
  assign y28348 = ~n37665 ;
  assign y28349 = ~1'b0 ;
  assign y28350 = n37667 ;
  assign y28351 = n37668 ;
  assign y28352 = ~n37669 ;
  assign y28353 = ~1'b0 ;
  assign y28354 = ~n37670 ;
  assign y28355 = n31948 ;
  assign y28356 = ~1'b0 ;
  assign y28357 = ~n37675 ;
  assign y28358 = n37676 ;
  assign y28359 = ~n24260 ;
  assign y28360 = n37680 ;
  assign y28361 = n14647 ;
  assign y28362 = ~1'b0 ;
  assign y28363 = ~1'b0 ;
  assign y28364 = 1'b0 ;
  assign y28365 = ~1'b0 ;
  assign y28366 = ~n6194 ;
  assign y28367 = n37683 ;
  assign y28368 = n37684 ;
  assign y28369 = n37685 ;
  assign y28370 = ~1'b0 ;
  assign y28371 = n37690 ;
  assign y28372 = ~n37692 ;
  assign y28373 = ~1'b0 ;
  assign y28374 = ~1'b0 ;
  assign y28375 = ~1'b0 ;
  assign y28376 = n615 ;
  assign y28377 = ~1'b0 ;
  assign y28378 = ~1'b0 ;
  assign y28379 = n37693 ;
  assign y28380 = n37696 ;
  assign y28381 = 1'b0 ;
  assign y28382 = ~n10066 ;
  assign y28383 = n37697 ;
  assign y28384 = ~1'b0 ;
  assign y28385 = ~n37698 ;
  assign y28386 = ~1'b0 ;
  assign y28387 = ~1'b0 ;
  assign y28388 = ~1'b0 ;
  assign y28389 = n35500 ;
  assign y28390 = n37700 ;
  assign y28391 = n34018 ;
  assign y28392 = n37701 ;
  assign y28393 = 1'b0 ;
  assign y28394 = n2256 ;
  assign y28395 = ~1'b0 ;
  assign y28396 = ~n37706 ;
  assign y28397 = ~1'b0 ;
  assign y28398 = n37707 ;
  assign y28399 = ~n2431 ;
  assign y28400 = ~n37712 ;
  assign y28401 = n7416 ;
  assign y28402 = ~1'b0 ;
  assign y28403 = ~1'b0 ;
  assign y28404 = ~n37715 ;
  assign y28405 = 1'b0 ;
  assign y28406 = ~n37716 ;
  assign y28407 = ~n37717 ;
  assign y28408 = n37719 ;
  assign y28409 = ~n37720 ;
  assign y28410 = ~n10596 ;
  assign y28411 = ~n37723 ;
  assign y28412 = ~n19109 ;
  assign y28413 = n6374 ;
  assign y28414 = ~n37725 ;
  assign y28415 = ~1'b0 ;
  assign y28416 = ~1'b0 ;
  assign y28417 = n37726 ;
  assign y28418 = n27434 ;
  assign y28419 = ~1'b0 ;
  assign y28420 = ~n37727 ;
  assign y28421 = n20954 ;
  assign y28422 = ~1'b0 ;
  assign y28423 = ~1'b0 ;
  assign y28424 = n2929 ;
  assign y28425 = ~n37728 ;
  assign y28426 = ~n37729 ;
  assign y28427 = ~n37730 ;
  assign y28428 = n37731 ;
  assign y28429 = 1'b0 ;
  assign y28430 = ~1'b0 ;
  assign y28431 = ~n37738 ;
  assign y28432 = n37740 ;
  assign y28433 = 1'b0 ;
  assign y28434 = n37741 ;
  assign y28435 = ~1'b0 ;
  assign y28436 = 1'b0 ;
  assign y28437 = n37743 ;
  assign y28438 = n37744 ;
  assign y28439 = 1'b0 ;
  assign y28440 = ~n37746 ;
  assign y28441 = ~n37751 ;
  assign y28442 = ~1'b0 ;
  assign y28443 = ~1'b0 ;
  assign y28444 = n16656 ;
  assign y28445 = ~1'b0 ;
  assign y28446 = ~n37763 ;
  assign y28447 = ~n12721 ;
  assign y28448 = ~1'b0 ;
  assign y28449 = ~1'b0 ;
  assign y28450 = ~1'b0 ;
  assign y28451 = ~n37765 ;
  assign y28452 = n37766 ;
  assign y28453 = ~1'b0 ;
  assign y28454 = n37770 ;
  assign y28455 = ~n37771 ;
  assign y28456 = ~n37774 ;
  assign y28457 = n37775 ;
  assign y28458 = ~n29159 ;
  assign y28459 = 1'b0 ;
  assign y28460 = ~n37779 ;
  assign y28461 = ~1'b0 ;
  assign y28462 = n37780 ;
  assign y28463 = ~1'b0 ;
  assign y28464 = ~n37781 ;
  assign y28465 = ~n37784 ;
  assign y28466 = ~1'b0 ;
  assign y28467 = ~1'b0 ;
  assign y28468 = ~n37789 ;
  assign y28469 = ~n29524 ;
  assign y28470 = ~1'b0 ;
  assign y28471 = ~1'b0 ;
  assign y28472 = n37792 ;
  assign y28473 = ~1'b0 ;
  assign y28474 = n37793 ;
  assign y28475 = n37794 ;
  assign y28476 = ~n37797 ;
  assign y28477 = ~1'b0 ;
  assign y28478 = ~1'b0 ;
  assign y28479 = ~n37799 ;
  assign y28480 = n37800 ;
  assign y28481 = n7355 ;
  assign y28482 = ~1'b0 ;
  assign y28483 = ~n37802 ;
  assign y28484 = ~n37803 ;
  assign y28485 = ~1'b0 ;
  assign y28486 = ~n37807 ;
  assign y28487 = ~n37809 ;
  assign y28488 = ~n37811 ;
  assign y28489 = ~1'b0 ;
  assign y28490 = ~n37813 ;
  assign y28491 = n3743 ;
  assign y28492 = ~1'b0 ;
  assign y28493 = ~1'b0 ;
  assign y28494 = ~n37816 ;
  assign y28495 = ~1'b0 ;
  assign y28496 = ~1'b0 ;
  assign y28497 = n37817 ;
  assign y28498 = n37823 ;
  assign y28499 = n15329 ;
  assign y28500 = n5180 ;
  assign y28501 = 1'b0 ;
  assign y28502 = ~1'b0 ;
  assign y28503 = ~n12298 ;
  assign y28504 = n37824 ;
  assign y28505 = ~1'b0 ;
  assign y28506 = ~n37825 ;
  assign y28507 = ~1'b0 ;
  assign y28508 = ~1'b0 ;
  assign y28509 = ~1'b0 ;
  assign y28510 = ~1'b0 ;
  assign y28511 = ~1'b0 ;
  assign y28512 = ~1'b0 ;
  assign y28513 = ~n37827 ;
  assign y28514 = ~n29340 ;
  assign y28515 = n37830 ;
  assign y28516 = ~1'b0 ;
  assign y28517 = ~n2680 ;
  assign y28518 = ~n37835 ;
  assign y28519 = ~1'b0 ;
  assign y28520 = ~1'b0 ;
  assign y28521 = n37838 ;
  assign y28522 = 1'b0 ;
  assign y28523 = ~n37840 ;
  assign y28524 = n37841 ;
  assign y28525 = 1'b0 ;
  assign y28526 = n37842 ;
  assign y28527 = ~n37843 ;
  assign y28528 = ~n29397 ;
  assign y28529 = ~1'b0 ;
  assign y28530 = ~1'b0 ;
  assign y28531 = ~1'b0 ;
  assign y28532 = n37844 ;
  assign y28533 = ~n37845 ;
  assign y28534 = n16792 ;
  assign y28535 = n37846 ;
  assign y28536 = 1'b0 ;
  assign y28537 = ~n37848 ;
  assign y28538 = ~1'b0 ;
  assign y28539 = ~n37852 ;
  assign y28540 = n5005 ;
  assign y28541 = n37854 ;
  assign y28542 = ~1'b0 ;
  assign y28543 = n4112 ;
  assign y28544 = ~1'b0 ;
  assign y28545 = ~n37857 ;
  assign y28546 = ~n37860 ;
  assign y28547 = n17673 ;
  assign y28548 = ~n36495 ;
  assign y28549 = ~1'b0 ;
  assign y28550 = ~n37861 ;
  assign y28551 = ~n37864 ;
  assign y28552 = ~n37866 ;
  assign y28553 = ~n29860 ;
  assign y28554 = ~1'b0 ;
  assign y28555 = ~1'b0 ;
  assign y28556 = 1'b0 ;
  assign y28557 = ~1'b0 ;
  assign y28558 = ~1'b0 ;
  assign y28559 = n37868 ;
  assign y28560 = ~n37869 ;
  assign y28561 = ~1'b0 ;
  assign y28562 = ~1'b0 ;
  assign y28563 = ~n37870 ;
  assign y28564 = ~1'b0 ;
  assign y28565 = ~n37873 ;
  assign y28566 = ~1'b0 ;
  assign y28567 = ~n37877 ;
  assign y28568 = ~n37878 ;
  assign y28569 = ~1'b0 ;
  assign y28570 = ~1'b0 ;
  assign y28571 = ~1'b0 ;
  assign y28572 = ~1'b0 ;
  assign y28573 = ~n2813 ;
  assign y28574 = n12045 ;
  assign y28575 = ~1'b0 ;
  assign y28576 = ~1'b0 ;
  assign y28577 = n37881 ;
  assign y28578 = ~1'b0 ;
  assign y28579 = ~1'b0 ;
  assign y28580 = ~1'b0 ;
  assign y28581 = ~n37883 ;
  assign y28582 = ~1'b0 ;
  assign y28583 = n37887 ;
  assign y28584 = ~1'b0 ;
  assign y28585 = ~n622 ;
  assign y28586 = ~n37891 ;
  assign y28587 = ~n37892 ;
  assign y28588 = ~n37893 ;
  assign y28589 = ~n37894 ;
  assign y28590 = ~n32911 ;
  assign y28591 = n19633 ;
  assign y28592 = n37897 ;
  assign y28593 = ~n37898 ;
  assign y28594 = ~n37900 ;
  assign y28595 = ~n6753 ;
  assign y28596 = ~n7855 ;
  assign y28597 = ~1'b0 ;
  assign y28598 = ~n37906 ;
  assign y28599 = ~1'b0 ;
  assign y28600 = n30066 ;
  assign y28601 = ~1'b0 ;
  assign y28602 = ~n37907 ;
  assign y28603 = ~n12058 ;
  assign y28604 = n37908 ;
  assign y28605 = ~1'b0 ;
  assign y28606 = n37909 ;
  assign y28607 = ~1'b0 ;
  assign y28608 = n37911 ;
  assign y28609 = n37912 ;
  assign y28610 = ~1'b0 ;
  assign y28611 = n37913 ;
  assign y28612 = n37915 ;
  assign y28613 = n37917 ;
  assign y28614 = ~n37919 ;
  assign y28615 = ~n1954 ;
  assign y28616 = ~n37923 ;
  assign y28617 = n37926 ;
  assign y28618 = ~1'b0 ;
  assign y28619 = n37928 ;
  assign y28620 = n37929 ;
  assign y28621 = ~n37930 ;
  assign y28622 = ~n37934 ;
  assign y28623 = ~n37940 ;
  assign y28624 = ~n6585 ;
  assign y28625 = n37943 ;
  assign y28626 = n37945 ;
  assign y28627 = 1'b0 ;
  assign y28628 = ~n37946 ;
  assign y28629 = ~1'b0 ;
  assign y28630 = ~n37948 ;
  assign y28631 = ~1'b0 ;
  assign y28632 = ~n37949 ;
  assign y28633 = ~1'b0 ;
  assign y28634 = n37955 ;
  assign y28635 = ~n37958 ;
  assign y28636 = n37959 ;
  assign y28637 = ~1'b0 ;
  assign y28638 = 1'b0 ;
  assign y28639 = ~1'b0 ;
  assign y28640 = ~1'b0 ;
  assign y28641 = n37960 ;
  assign y28642 = ~1'b0 ;
  assign y28643 = n37965 ;
  assign y28644 = n37968 ;
  assign y28645 = ~n37971 ;
  assign y28646 = n37972 ;
  assign y28647 = 1'b0 ;
  assign y28648 = ~n37974 ;
  assign y28649 = ~n13928 ;
  assign y28650 = ~n14189 ;
  assign y28651 = ~1'b0 ;
  assign y28652 = ~1'b0 ;
  assign y28653 = n37976 ;
  assign y28654 = ~1'b0 ;
  assign y28655 = n37977 ;
  assign y28656 = n37995 ;
  assign y28657 = n37996 ;
  assign y28658 = n37999 ;
  assign y28659 = n38000 ;
  assign y28660 = ~1'b0 ;
  assign y28661 = ~1'b0 ;
  assign y28662 = ~n38004 ;
  assign y28663 = ~1'b0 ;
  assign y28664 = ~n38005 ;
  assign y28665 = ~1'b0 ;
  assign y28666 = ~1'b0 ;
  assign y28667 = ~n38010 ;
  assign y28668 = ~1'b0 ;
  assign y28669 = ~n38015 ;
  assign y28670 = 1'b0 ;
  assign y28671 = n38017 ;
  assign y28672 = n2348 ;
  assign y28673 = ~1'b0 ;
  assign y28674 = ~1'b0 ;
  assign y28675 = ~n38019 ;
  assign y28676 = ~1'b0 ;
  assign y28677 = ~n38022 ;
  assign y28678 = n38023 ;
  assign y28679 = n38025 ;
  assign y28680 = n38027 ;
  assign y28681 = ~n38028 ;
  assign y28682 = n38036 ;
  assign y28683 = n38038 ;
  assign y28684 = ~n38039 ;
  assign y28685 = n31275 ;
  assign y28686 = n9409 ;
  assign y28687 = ~1'b0 ;
  assign y28688 = ~1'b0 ;
  assign y28689 = ~1'b0 ;
  assign y28690 = n38040 ;
  assign y28691 = ~1'b0 ;
  assign y28692 = ~1'b0 ;
  assign y28693 = ~n38041 ;
  assign y28694 = n38044 ;
  assign y28695 = ~n38055 ;
  assign y28696 = n14748 ;
  assign y28697 = ~n11164 ;
  assign y28698 = ~1'b0 ;
  assign y28699 = n20644 ;
  assign y28700 = n29918 ;
  assign y28701 = ~n38056 ;
  assign y28702 = ~n38058 ;
  assign y28703 = n38063 ;
  assign y28704 = ~1'b0 ;
  assign y28705 = ~1'b0 ;
  assign y28706 = n38065 ;
  assign y28707 = ~n38066 ;
  assign y28708 = n507 ;
  assign y28709 = ~1'b0 ;
  assign y28710 = n38067 ;
  assign y28711 = ~1'b0 ;
  assign y28712 = n38069 ;
  assign y28713 = ~n1106 ;
  assign y28714 = ~1'b0 ;
  assign y28715 = ~n38073 ;
  assign y28716 = ~n38075 ;
  assign y28717 = ~n38076 ;
  assign y28718 = 1'b0 ;
  assign y28719 = ~n38078 ;
  assign y28720 = ~1'b0 ;
  assign y28721 = n38079 ;
  assign y28722 = ~1'b0 ;
  assign y28723 = ~n38080 ;
  assign y28724 = ~n38089 ;
  assign y28725 = ~1'b0 ;
  assign y28726 = ~1'b0 ;
  assign y28727 = ~1'b0 ;
  assign y28728 = n38090 ;
  assign y28729 = ~n38093 ;
  assign y28730 = ~1'b0 ;
  assign y28731 = ~n38096 ;
  assign y28732 = n38098 ;
  assign y28733 = n38101 ;
  assign y28734 = ~n20808 ;
  assign y28735 = ~n38104 ;
  assign y28736 = n789 ;
  assign y28737 = n38106 ;
  assign y28738 = ~1'b0 ;
  assign y28739 = n38108 ;
  assign y28740 = n38111 ;
  assign y28741 = ~1'b0 ;
  assign y28742 = ~1'b0 ;
  assign y28743 = ~n38112 ;
  assign y28744 = ~1'b0 ;
  assign y28745 = n26656 ;
  assign y28746 = n38116 ;
  assign y28747 = n22362 ;
  assign y28748 = ~1'b0 ;
  assign y28749 = ~n4748 ;
  assign y28750 = n38117 ;
  assign y28751 = ~1'b0 ;
  assign y28752 = ~1'b0 ;
  assign y28753 = ~1'b0 ;
  assign y28754 = n14306 ;
  assign y28755 = ~1'b0 ;
  assign y28756 = n38119 ;
  assign y28757 = n38120 ;
  assign y28758 = ~n38121 ;
  assign y28759 = ~n38122 ;
  assign y28760 = ~n38126 ;
  assign y28761 = ~n38129 ;
  assign y28762 = ~1'b0 ;
  assign y28763 = ~1'b0 ;
  assign y28764 = n38130 ;
  assign y28765 = n7506 ;
  assign y28766 = ~n18296 ;
  assign y28767 = ~1'b0 ;
  assign y28768 = n38131 ;
  assign y28769 = 1'b0 ;
  assign y28770 = n38132 ;
  assign y28771 = ~n38133 ;
  assign y28772 = ~1'b0 ;
  assign y28773 = n38136 ;
  assign y28774 = n38138 ;
  assign y28775 = n38139 ;
  assign y28776 = ~n19632 ;
  assign y28777 = ~1'b0 ;
  assign y28778 = ~n38140 ;
  assign y28779 = ~n38141 ;
  assign y28780 = ~n38144 ;
  assign y28781 = ~n38146 ;
  assign y28782 = ~1'b0 ;
  assign y28783 = n38149 ;
  assign y28784 = ~1'b0 ;
  assign y28785 = ~1'b0 ;
  assign y28786 = ~n38150 ;
  assign y28787 = ~1'b0 ;
  assign y28788 = ~1'b0 ;
  assign y28789 = ~1'b0 ;
  assign y28790 = ~1'b0 ;
  assign y28791 = n38151 ;
  assign y28792 = 1'b0 ;
  assign y28793 = n38155 ;
  assign y28794 = ~1'b0 ;
  assign y28795 = n38160 ;
  assign y28796 = n38162 ;
  assign y28797 = ~1'b0 ;
  assign y28798 = ~1'b0 ;
  assign y28799 = n38163 ;
  assign y28800 = ~1'b0 ;
  assign y28801 = n38164 ;
  assign y28802 = ~n38167 ;
  assign y28803 = ~n38168 ;
  assign y28804 = ~1'b0 ;
  assign y28805 = 1'b0 ;
  assign y28806 = ~1'b0 ;
  assign y28807 = n38169 ;
  assign y28808 = ~1'b0 ;
  assign y28809 = ~n38170 ;
  assign y28810 = 1'b0 ;
  assign y28811 = ~1'b0 ;
  assign y28812 = n38171 ;
  assign y28813 = n997 ;
  assign y28814 = n38179 ;
  assign y28815 = ~1'b0 ;
  assign y28816 = ~1'b0 ;
  assign y28817 = ~n38180 ;
  assign y28818 = n38181 ;
  assign y28819 = ~n38185 ;
  assign y28820 = n38187 ;
  assign y28821 = ~n38189 ;
  assign y28822 = ~1'b0 ;
  assign y28823 = ~1'b0 ;
  assign y28824 = n38191 ;
  assign y28825 = ~n38193 ;
  assign y28826 = ~1'b0 ;
  assign y28827 = ~n38194 ;
  assign y28828 = ~n38197 ;
  assign y28829 = n38198 ;
  assign y28830 = ~1'b0 ;
  assign y28831 = n16438 ;
  assign y28832 = n38201 ;
  assign y28833 = 1'b0 ;
  assign y28834 = 1'b0 ;
  assign y28835 = n38202 ;
  assign y28836 = ~n38204 ;
  assign y28837 = ~1'b0 ;
  assign y28838 = ~1'b0 ;
  assign y28839 = ~1'b0 ;
  assign y28840 = n38206 ;
  assign y28841 = n38209 ;
  assign y28842 = ~1'b0 ;
  assign y28843 = ~1'b0 ;
  assign y28844 = n38210 ;
  assign y28845 = n1152 ;
  assign y28846 = n38211 ;
  assign y28847 = ~n38215 ;
  assign y28848 = ~n38218 ;
  assign y28849 = ~n38223 ;
  assign y28850 = 1'b0 ;
  assign y28851 = ~n4297 ;
  assign y28852 = ~n38228 ;
  assign y28853 = ~1'b0 ;
  assign y28854 = ~n38230 ;
  assign y28855 = ~n38232 ;
  assign y28856 = n38233 ;
  assign y28857 = ~n4633 ;
  assign y28858 = ~n38234 ;
  assign y28859 = n38238 ;
  assign y28860 = ~1'b0 ;
  assign y28861 = ~1'b0 ;
  assign y28862 = ~n14100 ;
  assign y28863 = ~n21767 ;
  assign y28864 = n38240 ;
  assign y28865 = ~1'b0 ;
  assign y28866 = n38242 ;
  assign y28867 = ~1'b0 ;
  assign y28868 = ~n38247 ;
  assign y28869 = n38248 ;
  assign y28870 = ~1'b0 ;
  assign y28871 = ~1'b0 ;
  assign y28872 = ~1'b0 ;
  assign y28873 = ~1'b0 ;
  assign y28874 = ~1'b0 ;
  assign y28875 = 1'b0 ;
  assign y28876 = ~n38258 ;
  assign y28877 = n16491 ;
  assign y28878 = ~1'b0 ;
  assign y28879 = n38261 ;
  assign y28880 = ~1'b0 ;
  assign y28881 = n38262 ;
  assign y28882 = ~n38265 ;
  assign y28883 = n38274 ;
  assign y28884 = ~n38275 ;
  assign y28885 = n38279 ;
  assign y28886 = ~1'b0 ;
  assign y28887 = ~1'b0 ;
  assign y28888 = ~n38280 ;
  assign y28889 = ~n38286 ;
  assign y28890 = ~n22165 ;
  assign y28891 = ~n38287 ;
  assign y28892 = ~1'b0 ;
  assign y28893 = ~1'b0 ;
  assign y28894 = ~n38291 ;
  assign y28895 = ~1'b0 ;
  assign y28896 = n38292 ;
  assign y28897 = ~1'b0 ;
  assign y28898 = ~n38294 ;
  assign y28899 = ~n38297 ;
  assign y28900 = ~n38299 ;
  assign y28901 = n38300 ;
  assign y28902 = ~n38303 ;
  assign y28903 = ~1'b0 ;
  assign y28904 = n5180 ;
  assign y28905 = ~n20010 ;
  assign y28906 = ~1'b0 ;
  assign y28907 = ~1'b0 ;
  assign y28908 = ~n38304 ;
  assign y28909 = ~n38305 ;
  assign y28910 = ~n38306 ;
  assign y28911 = n38308 ;
  assign y28912 = ~1'b0 ;
  assign y28913 = ~1'b0 ;
  assign y28914 = ~n38310 ;
  assign y28915 = ~1'b0 ;
  assign y28916 = ~1'b0 ;
  assign y28917 = ~1'b0 ;
  assign y28918 = n9335 ;
  assign y28919 = ~1'b0 ;
  assign y28920 = n38313 ;
  assign y28921 = n12507 ;
  assign y28922 = ~1'b0 ;
  assign y28923 = n38318 ;
  assign y28924 = ~1'b0 ;
  assign y28925 = ~1'b0 ;
  assign y28926 = n38321 ;
  assign y28927 = n9448 ;
  assign y28928 = 1'b0 ;
  assign y28929 = ~1'b0 ;
  assign y28930 = n38322 ;
  assign y28931 = n38325 ;
  assign y28932 = ~n38328 ;
  assign y28933 = ~n38329 ;
  assign y28934 = ~1'b0 ;
  assign y28935 = n38331 ;
  assign y28936 = ~n37538 ;
  assign y28937 = 1'b0 ;
  assign y28938 = n38332 ;
  assign y28939 = ~n38334 ;
  assign y28940 = ~n11827 ;
  assign y28941 = ~1'b0 ;
  assign y28942 = n38336 ;
  assign y28943 = ~n38339 ;
  assign y28944 = ~n38341 ;
  assign y28945 = ~n38342 ;
  assign y28946 = ~1'b0 ;
  assign y28947 = ~n158 ;
  assign y28948 = ~n38343 ;
  assign y28949 = ~n38345 ;
  assign y28950 = ~1'b0 ;
  assign y28951 = ~1'b0 ;
  assign y28952 = ~n12343 ;
  assign y28953 = ~n38352 ;
  assign y28954 = ~n38354 ;
  assign y28955 = n38356 ;
  assign y28956 = 1'b0 ;
  assign y28957 = ~1'b0 ;
  assign y28958 = n3424 ;
  assign y28959 = ~n38358 ;
  assign y28960 = ~1'b0 ;
  assign y28961 = ~1'b0 ;
  assign y28962 = n38359 ;
  assign y28963 = n38360 ;
  assign y28964 = n27537 ;
  assign y28965 = n38364 ;
  assign y28966 = n38367 ;
  assign y28967 = ~1'b0 ;
  assign y28968 = ~1'b0 ;
  assign y28969 = n38375 ;
  assign y28970 = n14785 ;
  assign y28971 = ~n38377 ;
  assign y28972 = ~1'b0 ;
  assign y28973 = n38378 ;
  assign y28974 = ~1'b0 ;
  assign y28975 = ~1'b0 ;
  assign y28976 = ~n38379 ;
  assign y28977 = n38380 ;
  assign y28978 = ~n38381 ;
  assign y28979 = ~n38383 ;
  assign y28980 = ~1'b0 ;
  assign y28981 = ~n38384 ;
  assign y28982 = ~n38385 ;
  assign y28983 = ~n38388 ;
  assign y28984 = ~1'b0 ;
  assign y28985 = ~n38390 ;
  assign y28986 = n38391 ;
  assign y28987 = ~1'b0 ;
  assign y28988 = ~n38393 ;
  assign y28989 = n75 ;
  assign y28990 = ~1'b0 ;
  assign y28991 = 1'b0 ;
  assign y28992 = ~n38397 ;
  assign y28993 = n38398 ;
  assign y28994 = ~n38400 ;
  assign y28995 = ~1'b0 ;
  assign y28996 = ~1'b0 ;
  assign y28997 = 1'b0 ;
  assign y28998 = n38403 ;
  assign y28999 = ~n3585 ;
  assign y29000 = n13815 ;
  assign y29001 = ~n38404 ;
  assign y29002 = n38405 ;
  assign y29003 = ~1'b0 ;
  assign y29004 = ~1'b0 ;
  assign y29005 = ~1'b0 ;
  assign y29006 = n38406 ;
  assign y29007 = ~1'b0 ;
  assign y29008 = ~1'b0 ;
  assign y29009 = n38407 ;
  assign y29010 = n38408 ;
  assign y29011 = ~n38409 ;
  assign y29012 = n38411 ;
  assign y29013 = ~1'b0 ;
  assign y29014 = ~n6025 ;
  assign y29015 = n38414 ;
  assign y29016 = ~1'b0 ;
  assign y29017 = ~1'b0 ;
  assign y29018 = ~n2462 ;
  assign y29019 = n38416 ;
  assign y29020 = ~1'b0 ;
  assign y29021 = ~1'b0 ;
  assign y29022 = ~n2136 ;
  assign y29023 = n3273 ;
  assign y29024 = n38418 ;
  assign y29025 = ~n38421 ;
  assign y29026 = ~1'b0 ;
  assign y29027 = ~n38422 ;
  assign y29028 = ~1'b0 ;
  assign y29029 = 1'b0 ;
  assign y29030 = ~n38423 ;
  assign y29031 = ~n38424 ;
  assign y29032 = ~1'b0 ;
  assign y29033 = ~1'b0 ;
  assign y29034 = 1'b0 ;
  assign y29035 = n38426 ;
  assign y29036 = n3743 ;
  assign y29037 = ~1'b0 ;
  assign y29038 = 1'b0 ;
  assign y29039 = ~1'b0 ;
  assign y29040 = ~1'b0 ;
  assign y29041 = ~1'b0 ;
  assign y29042 = ~n38427 ;
  assign y29043 = n33350 ;
  assign y29044 = ~1'b0 ;
  assign y29045 = ~1'b0 ;
  assign y29046 = ~1'b0 ;
  assign y29047 = n37644 ;
  assign y29048 = ~1'b0 ;
  assign y29049 = ~1'b0 ;
  assign y29050 = ~1'b0 ;
  assign y29051 = ~n4898 ;
  assign y29052 = 1'b0 ;
  assign y29053 = ~n38428 ;
  assign y29054 = ~1'b0 ;
  assign y29055 = ~1'b0 ;
  assign y29056 = ~1'b0 ;
  assign y29057 = n38429 ;
  assign y29058 = ~1'b0 ;
  assign y29059 = n38430 ;
  assign y29060 = n10787 ;
  assign y29061 = ~1'b0 ;
  assign y29062 = n11055 ;
  assign y29063 = ~1'b0 ;
  assign y29064 = ~1'b0 ;
  assign y29065 = ~1'b0 ;
  assign y29066 = n38431 ;
  assign y29067 = n38436 ;
  assign y29068 = ~n38438 ;
  assign y29069 = ~1'b0 ;
  assign y29070 = n22429 ;
  assign y29071 = n38440 ;
  assign y29072 = ~1'b0 ;
  assign y29073 = ~n38441 ;
  assign y29074 = ~1'b0 ;
  assign y29075 = ~1'b0 ;
  assign y29076 = 1'b0 ;
  assign y29077 = ~n38442 ;
  assign y29078 = ~1'b0 ;
  assign y29079 = n38447 ;
  assign y29080 = ~n33048 ;
  assign y29081 = 1'b0 ;
  assign y29082 = n38448 ;
  assign y29083 = ~1'b0 ;
  assign y29084 = n38450 ;
  assign y29085 = ~1'b0 ;
  assign y29086 = n38455 ;
  assign y29087 = ~1'b0 ;
  assign y29088 = ~n38460 ;
  assign y29089 = n38463 ;
  assign y29090 = ~1'b0 ;
  assign y29091 = ~1'b0 ;
  assign y29092 = ~n26827 ;
  assign y29093 = ~1'b0 ;
  assign y29094 = ~n38465 ;
  assign y29095 = ~1'b0 ;
  assign y29096 = 1'b0 ;
  assign y29097 = 1'b0 ;
  assign y29098 = ~1'b0 ;
  assign y29099 = ~1'b0 ;
  assign y29100 = ~n38467 ;
  assign y29101 = ~1'b0 ;
  assign y29102 = ~1'b0 ;
  assign y29103 = ~n38469 ;
  assign y29104 = ~n38473 ;
  assign y29105 = ~n38474 ;
  assign y29106 = ~1'b0 ;
  assign y29107 = ~n38477 ;
  assign y29108 = ~1'b0 ;
  assign y29109 = ~n38478 ;
  assign y29110 = n29221 ;
  assign y29111 = ~n38483 ;
  assign y29112 = ~1'b0 ;
  assign y29113 = ~1'b0 ;
  assign y29114 = 1'b0 ;
  assign y29115 = n38486 ;
  assign y29116 = ~1'b0 ;
  assign y29117 = n294 ;
  assign y29118 = ~n38487 ;
  assign y29119 = n38493 ;
  assign y29120 = ~1'b0 ;
  assign y29121 = ~n38498 ;
  assign y29122 = ~1'b0 ;
  assign y29123 = ~1'b0 ;
  assign y29124 = n2927 ;
  assign y29125 = ~1'b0 ;
  assign y29126 = ~n38500 ;
  assign y29127 = n38504 ;
  assign y29128 = 1'b0 ;
  assign y29129 = ~n38506 ;
  assign y29130 = n38508 ;
  assign y29131 = n3268 ;
  assign y29132 = ~n38509 ;
  assign y29133 = ~n38512 ;
  assign y29134 = n38519 ;
  assign y29135 = n38520 ;
  assign y29136 = ~1'b0 ;
  assign y29137 = ~n38522 ;
  assign y29138 = ~1'b0 ;
  assign y29139 = ~1'b0 ;
  assign y29140 = ~1'b0 ;
  assign y29141 = ~1'b0 ;
  assign y29142 = ~1'b0 ;
  assign y29143 = ~1'b0 ;
  assign y29144 = n38523 ;
  assign y29145 = ~1'b0 ;
  assign y29146 = n37126 ;
  assign y29147 = ~1'b0 ;
  assign y29148 = n38525 ;
  assign y29149 = n16791 ;
  assign y29150 = ~n38526 ;
  assign y29151 = ~n40 ;
  assign y29152 = ~n38531 ;
  assign y29153 = n38532 ;
  assign y29154 = ~1'b0 ;
  assign y29155 = n38538 ;
  assign y29156 = ~1'b0 ;
  assign y29157 = ~n29049 ;
  assign y29158 = ~n38540 ;
  assign y29159 = 1'b0 ;
  assign y29160 = ~1'b0 ;
  assign y29161 = ~n38542 ;
  assign y29162 = ~n38545 ;
  assign y29163 = n38546 ;
  assign y29164 = ~n38548 ;
  assign y29165 = ~n38552 ;
  assign y29166 = ~n3674 ;
  assign y29167 = ~n38554 ;
  assign y29168 = ~1'b0 ;
  assign y29169 = ~n9484 ;
  assign y29170 = ~n38557 ;
  assign y29171 = ~n38561 ;
  assign y29172 = n38563 ;
  assign y29173 = n38569 ;
  assign y29174 = n38570 ;
  assign y29175 = n38571 ;
  assign y29176 = n3718 ;
  assign y29177 = ~1'b0 ;
  assign y29178 = ~1'b0 ;
  assign y29179 = ~1'b0 ;
  assign y29180 = n38572 ;
  assign y29181 = ~1'b0 ;
  assign y29182 = ~1'b0 ;
  assign y29183 = n38573 ;
  assign y29184 = ~n38576 ;
  assign y29185 = ~n38577 ;
  assign y29186 = ~1'b0 ;
  assign y29187 = ~1'b0 ;
  assign y29188 = ~n38579 ;
  assign y29189 = 1'b0 ;
  assign y29190 = ~n38581 ;
  assign y29191 = ~n38584 ;
  assign y29192 = n38586 ;
  assign y29193 = ~n38588 ;
  assign y29194 = n38589 ;
  assign y29195 = ~1'b0 ;
  assign y29196 = n38591 ;
  assign y29197 = n38595 ;
  assign y29198 = ~n20517 ;
  assign y29199 = ~1'b0 ;
  assign y29200 = ~n38597 ;
  assign y29201 = ~n33386 ;
  assign y29202 = ~n38599 ;
  assign y29203 = ~1'b0 ;
  assign y29204 = n38600 ;
  assign y29205 = 1'b0 ;
  assign y29206 = n38601 ;
  assign y29207 = ~1'b0 ;
  assign y29208 = n38602 ;
  assign y29209 = ~1'b0 ;
  assign y29210 = 1'b0 ;
  assign y29211 = n38604 ;
  assign y29212 = ~n1435 ;
  assign y29213 = ~1'b0 ;
  assign y29214 = n38608 ;
  assign y29215 = n38614 ;
  assign y29216 = ~1'b0 ;
  assign y29217 = ~1'b0 ;
  assign y29218 = ~1'b0 ;
  assign y29219 = ~1'b0 ;
  assign y29220 = ~n38616 ;
  assign y29221 = ~n38618 ;
  assign y29222 = ~1'b0 ;
  assign y29223 = n38619 ;
  assign y29224 = n38623 ;
  assign y29225 = 1'b0 ;
  assign y29226 = n38625 ;
  assign y29227 = ~1'b0 ;
  assign y29228 = n38626 ;
  assign y29229 = ~1'b0 ;
  assign y29230 = n38627 ;
  assign y29231 = ~1'b0 ;
  assign y29232 = ~n38629 ;
  assign y29233 = ~1'b0 ;
  assign y29234 = ~n38635 ;
  assign y29235 = ~n38638 ;
  assign y29236 = ~1'b0 ;
  assign y29237 = ~1'b0 ;
  assign y29238 = ~1'b0 ;
  assign y29239 = n38641 ;
  assign y29240 = ~n22832 ;
  assign y29241 = n11931 ;
  assign y29242 = n38644 ;
  assign y29243 = ~n38646 ;
  assign y29244 = ~n38652 ;
  assign y29245 = n38653 ;
  assign y29246 = ~1'b0 ;
  assign y29247 = n38654 ;
  assign y29248 = ~1'b0 ;
  assign y29249 = n38655 ;
  assign y29250 = ~1'b0 ;
  assign y29251 = ~n1065 ;
  assign y29252 = ~1'b0 ;
  assign y29253 = ~n38658 ;
  assign y29254 = n38659 ;
  assign y29255 = n38662 ;
  assign y29256 = ~n38665 ;
  assign y29257 = ~n38667 ;
  assign y29258 = ~n38668 ;
  assign y29259 = n38669 ;
  assign y29260 = ~n38676 ;
  assign y29261 = n38677 ;
  assign y29262 = ~1'b0 ;
  assign y29263 = ~n7815 ;
  assign y29264 = ~1'b0 ;
  assign y29265 = ~n7754 ;
  assign y29266 = ~n38678 ;
  assign y29267 = ~n9233 ;
  assign y29268 = ~n38679 ;
  assign y29269 = n9675 ;
  assign y29270 = n38683 ;
  assign y29271 = ~n38684 ;
  assign y29272 = ~n38685 ;
  assign y29273 = n38687 ;
  assign y29274 = n38711 ;
  assign y29275 = n38714 ;
  assign y29276 = n35046 ;
  assign y29277 = ~n37812 ;
  assign y29278 = n38716 ;
  assign y29279 = ~1'b0 ;
  assign y29280 = ~n38717 ;
  assign y29281 = n38719 ;
  assign y29282 = ~1'b0 ;
  assign y29283 = ~1'b0 ;
  assign y29284 = ~n8453 ;
  assign y29285 = n38722 ;
  assign y29286 = ~n38724 ;
  assign y29287 = ~1'b0 ;
  assign y29288 = ~1'b0 ;
  assign y29289 = ~n38727 ;
  assign y29290 = ~n38728 ;
  assign y29291 = ~1'b0 ;
  assign y29292 = n38731 ;
  assign y29293 = ~n19944 ;
  assign y29294 = ~1'b0 ;
  assign y29295 = ~n38732 ;
  assign y29296 = ~n38734 ;
  assign y29297 = ~1'b0 ;
  assign y29298 = ~n38735 ;
  assign y29299 = ~n38736 ;
  assign y29300 = ~n1337 ;
  assign y29301 = ~n38737 ;
  assign y29302 = ~1'b0 ;
  assign y29303 = ~n38766 ;
  assign y29304 = ~1'b0 ;
  assign y29305 = ~n38767 ;
  assign y29306 = n5189 ;
  assign y29307 = ~n38769 ;
  assign y29308 = n38774 ;
  assign y29309 = n27037 ;
  assign y29310 = ~n38775 ;
  assign y29311 = ~n38777 ;
  assign y29312 = n38778 ;
  assign y29313 = ~n38780 ;
  assign y29314 = ~1'b0 ;
  assign y29315 = ~1'b0 ;
  assign y29316 = 1'b0 ;
  assign y29317 = n38781 ;
  assign y29318 = n38782 ;
  assign y29319 = n38783 ;
  assign y29320 = n38785 ;
  assign y29321 = ~1'b0 ;
  assign y29322 = n38786 ;
  assign y29323 = 1'b0 ;
  assign y29324 = ~1'b0 ;
  assign y29325 = n38787 ;
  assign y29326 = ~n9416 ;
  assign y29327 = ~1'b0 ;
  assign y29328 = ~1'b0 ;
  assign y29329 = 1'b0 ;
  assign y29330 = n38788 ;
  assign y29331 = ~1'b0 ;
  assign y29332 = n6159 ;
  assign y29333 = ~1'b0 ;
  assign y29334 = ~n38789 ;
  assign y29335 = ~n38790 ;
  assign y29336 = n16156 ;
  assign y29337 = ~1'b0 ;
  assign y29338 = n20240 ;
  assign y29339 = ~1'b0 ;
  assign y29340 = ~n38796 ;
  assign y29341 = ~n38797 ;
  assign y29342 = ~1'b0 ;
  assign y29343 = ~n38799 ;
  assign y29344 = n38803 ;
  assign y29345 = n8319 ;
  assign y29346 = ~1'b0 ;
  assign y29347 = ~1'b0 ;
  assign y29348 = ~1'b0 ;
  assign y29349 = n38804 ;
  assign y29350 = ~n38805 ;
  assign y29351 = n38808 ;
  assign y29352 = ~n38822 ;
  assign y29353 = ~n38824 ;
  assign y29354 = ~1'b0 ;
  assign y29355 = n38829 ;
  assign y29356 = ~1'b0 ;
  assign y29357 = ~1'b0 ;
  assign y29358 = ~1'b0 ;
  assign y29359 = ~n726 ;
  assign y29360 = 1'b0 ;
  assign y29361 = n33287 ;
  assign y29362 = n38830 ;
  assign y29363 = n28364 ;
  assign y29364 = ~n38840 ;
  assign y29365 = ~1'b0 ;
  assign y29366 = ~n38845 ;
  assign y29367 = ~n23341 ;
  assign y29368 = ~1'b0 ;
  assign y29369 = ~1'b0 ;
  assign y29370 = n38847 ;
  assign y29371 = ~n33218 ;
  assign y29372 = ~1'b0 ;
  assign y29373 = ~n38850 ;
  assign y29374 = ~1'b0 ;
  assign y29375 = n38851 ;
  assign y29376 = n38853 ;
  assign y29377 = ~n38857 ;
  assign y29378 = n2922 ;
  assign y29379 = n38863 ;
  assign y29380 = ~1'b0 ;
  assign y29381 = n38865 ;
  assign y29382 = ~1'b0 ;
  assign y29383 = ~n26331 ;
  assign y29384 = ~n38867 ;
  assign y29385 = ~n13125 ;
  assign y29386 = ~n7958 ;
  assign y29387 = ~n4823 ;
  assign y29388 = n38888 ;
  assign y29389 = ~1'b0 ;
  assign y29390 = ~1'b0 ;
  assign y29391 = ~n38889 ;
  assign y29392 = n2235 ;
  assign y29393 = 1'b0 ;
  assign y29394 = 1'b0 ;
  assign y29395 = ~1'b0 ;
  assign y29396 = ~1'b0 ;
  assign y29397 = ~n38891 ;
  assign y29398 = ~n38892 ;
  assign y29399 = ~n29740 ;
  assign y29400 = n38896 ;
  assign y29401 = ~n38897 ;
  assign y29402 = ~n38899 ;
  assign y29403 = ~n38902 ;
  assign y29404 = ~1'b0 ;
  assign y29405 = n38903 ;
  assign y29406 = ~n38905 ;
  assign y29407 = ~n38908 ;
  assign y29408 = ~1'b0 ;
  assign y29409 = ~n38910 ;
  assign y29410 = ~1'b0 ;
  assign y29411 = ~n38912 ;
  assign y29412 = n38915 ;
  assign y29413 = ~1'b0 ;
  assign y29414 = ~1'b0 ;
  assign y29415 = ~n15276 ;
  assign y29416 = ~1'b0 ;
  assign y29417 = ~1'b0 ;
  assign y29418 = ~1'b0 ;
  assign y29419 = ~n128 ;
  assign y29420 = n38916 ;
  assign y29421 = n38918 ;
  assign y29422 = n38919 ;
  assign y29423 = ~1'b0 ;
  assign y29424 = n38924 ;
  assign y29425 = n38926 ;
  assign y29426 = ~1'b0 ;
  assign y29427 = ~n38929 ;
  assign y29428 = ~1'b0 ;
  assign y29429 = ~1'b0 ;
  assign y29430 = ~1'b0 ;
  assign y29431 = n38931 ;
  assign y29432 = ~n38934 ;
  assign y29433 = ~1'b0 ;
  assign y29434 = ~n38935 ;
  assign y29435 = ~n38945 ;
  assign y29436 = n38948 ;
  assign y29437 = n38949 ;
  assign y29438 = ~1'b0 ;
  assign y29439 = n38954 ;
  assign y29440 = ~n38956 ;
  assign y29441 = ~1'b0 ;
  assign y29442 = ~n38961 ;
  assign y29443 = n38962 ;
  assign y29444 = ~1'b0 ;
  assign y29445 = ~1'b0 ;
  assign y29446 = ~1'b0 ;
  assign y29447 = n9252 ;
  assign y29448 = n38963 ;
  assign y29449 = ~1'b0 ;
  assign y29450 = ~1'b0 ;
  assign y29451 = ~n38964 ;
  assign y29452 = n14213 ;
  assign y29453 = ~n36593 ;
  assign y29454 = n38965 ;
  assign y29455 = ~1'b0 ;
  assign y29456 = 1'b0 ;
  assign y29457 = n38967 ;
  assign y29458 = ~1'b0 ;
  assign y29459 = n38969 ;
  assign y29460 = ~n38972 ;
  assign y29461 = ~n38979 ;
  assign y29462 = ~n38982 ;
  assign y29463 = ~1'b0 ;
  assign y29464 = ~n38983 ;
  assign y29465 = ~1'b0 ;
  assign y29466 = n21560 ;
  assign y29467 = ~1'b0 ;
  assign y29468 = n38986 ;
  assign y29469 = ~1'b0 ;
  assign y29470 = n38989 ;
  assign y29471 = ~1'b0 ;
  assign y29472 = ~n38992 ;
  assign y29473 = ~1'b0 ;
  assign y29474 = n38998 ;
  assign y29475 = n39000 ;
  assign y29476 = ~1'b0 ;
  assign y29477 = n39004 ;
  assign y29478 = ~n39006 ;
  assign y29479 = ~n39011 ;
  assign y29480 = 1'b0 ;
  assign y29481 = ~n17500 ;
  assign y29482 = ~n39012 ;
  assign y29483 = ~1'b0 ;
  assign y29484 = n5174 ;
  assign y29485 = 1'b0 ;
  assign y29486 = ~1'b0 ;
  assign y29487 = ~1'b0 ;
  assign y29488 = n39013 ;
  assign y29489 = n39015 ;
  assign y29490 = n39018 ;
  assign y29491 = ~n39019 ;
  assign y29492 = ~1'b0 ;
  assign y29493 = ~n39023 ;
  assign y29494 = ~1'b0 ;
  assign y29495 = n3418 ;
  assign y29496 = ~1'b0 ;
  assign y29497 = n39025 ;
  assign y29498 = ~n39026 ;
  assign y29499 = ~n39030 ;
  assign y29500 = ~1'b0 ;
  assign y29501 = ~n39031 ;
  assign y29502 = 1'b0 ;
  assign y29503 = ~n39035 ;
  assign y29504 = ~n39040 ;
  assign y29505 = ~n39046 ;
  assign y29506 = n21615 ;
  assign y29507 = 1'b0 ;
  assign y29508 = ~n39051 ;
  assign y29509 = n14418 ;
  assign y29510 = n39052 ;
  assign y29511 = n39053 ;
  assign y29512 = ~1'b0 ;
  assign y29513 = ~n39055 ;
  assign y29514 = n39057 ;
  assign y29515 = n39058 ;
  assign y29516 = ~1'b0 ;
  assign y29517 = ~1'b0 ;
  assign y29518 = ~1'b0 ;
  assign y29519 = n39059 ;
  assign y29520 = ~1'b0 ;
  assign y29521 = n39061 ;
  assign y29522 = n39063 ;
  assign y29523 = ~1'b0 ;
  assign y29524 = ~1'b0 ;
  assign y29525 = ~n39065 ;
  assign y29526 = n39066 ;
  assign y29527 = n16190 ;
  assign y29528 = n39068 ;
  assign y29529 = ~n743 ;
  assign y29530 = ~1'b0 ;
  assign y29531 = n39069 ;
  assign y29532 = ~n39070 ;
  assign y29533 = n39075 ;
  assign y29534 = ~1'b0 ;
  assign y29535 = n27837 ;
  assign y29536 = ~1'b0 ;
  assign y29537 = n39076 ;
  assign y29538 = ~1'b0 ;
  assign y29539 = ~1'b0 ;
  assign y29540 = 1'b0 ;
  assign y29541 = n39078 ;
  assign y29542 = ~1'b0 ;
  assign y29543 = ~1'b0 ;
  assign y29544 = ~n27840 ;
  assign y29545 = ~n39080 ;
  assign y29546 = ~n39082 ;
  assign y29547 = n39083 ;
  assign y29548 = ~1'b0 ;
  assign y29549 = n39084 ;
  assign y29550 = n39085 ;
  assign y29551 = ~1'b0 ;
  assign y29552 = n15765 ;
  assign y29553 = n39087 ;
  assign y29554 = ~1'b0 ;
  assign y29555 = ~1'b0 ;
  assign y29556 = ~n39089 ;
  assign y29557 = ~1'b0 ;
  assign y29558 = ~1'b0 ;
  assign y29559 = ~1'b0 ;
  assign y29560 = ~n39091 ;
  assign y29561 = n21636 ;
  assign y29562 = ~n39093 ;
  assign y29563 = n7289 ;
  assign y29564 = n39097 ;
  assign y29565 = n39099 ;
  assign y29566 = n39100 ;
  assign y29567 = n39102 ;
  assign y29568 = ~1'b0 ;
  assign y29569 = ~1'b0 ;
  assign y29570 = ~n39107 ;
  assign y29571 = n39110 ;
  assign y29572 = ~1'b0 ;
  assign y29573 = ~1'b0 ;
  assign y29574 = ~1'b0 ;
  assign y29575 = ~1'b0 ;
  assign y29576 = ~n39113 ;
  assign y29577 = n2065 ;
  assign y29578 = n39116 ;
  assign y29579 = ~1'b0 ;
  assign y29580 = ~n39117 ;
  assign y29581 = ~1'b0 ;
  assign y29582 = n39121 ;
  assign y29583 = ~n39132 ;
  assign y29584 = 1'b0 ;
  assign y29585 = ~1'b0 ;
  assign y29586 = ~1'b0 ;
  assign y29587 = n39136 ;
  assign y29588 = ~n39137 ;
  assign y29589 = ~n13760 ;
  assign y29590 = ~n39140 ;
  assign y29591 = n39142 ;
  assign y29592 = ~n39145 ;
  assign y29593 = ~1'b0 ;
  assign y29594 = ~1'b0 ;
  assign y29595 = n39146 ;
  assign y29596 = ~n39149 ;
  assign y29597 = ~n39150 ;
  assign y29598 = ~1'b0 ;
  assign y29599 = ~n39151 ;
  assign y29600 = ~1'b0 ;
  assign y29601 = ~n39152 ;
  assign y29602 = ~1'b0 ;
  assign y29603 = ~n4865 ;
  assign y29604 = ~1'b0 ;
  assign y29605 = n39159 ;
  assign y29606 = n39160 ;
  assign y29607 = n39161 ;
  assign y29608 = n39163 ;
  assign y29609 = ~1'b0 ;
  assign y29610 = ~n1350 ;
  assign y29611 = ~1'b0 ;
  assign y29612 = ~1'b0 ;
  assign y29613 = n39166 ;
  assign y29614 = n39168 ;
  assign y29615 = n39171 ;
  assign y29616 = ~1'b0 ;
  assign y29617 = ~n39175 ;
  assign y29618 = n39177 ;
  assign y29619 = 1'b0 ;
  assign y29620 = ~1'b0 ;
  assign y29621 = ~n39180 ;
  assign y29622 = ~1'b0 ;
  assign y29623 = n39181 ;
  assign y29624 = ~1'b0 ;
  assign y29625 = n39186 ;
  assign y29626 = n7083 ;
  assign y29627 = n14887 ;
  assign y29628 = n39188 ;
  assign y29629 = n39190 ;
  assign y29630 = ~1'b0 ;
  assign y29631 = 1'b0 ;
  assign y29632 = ~n39191 ;
  assign y29633 = ~n39192 ;
  assign y29634 = ~n39195 ;
  assign y29635 = ~1'b0 ;
  assign y29636 = ~1'b0 ;
  assign y29637 = ~1'b0 ;
  assign y29638 = ~1'b0 ;
  assign y29639 = n39196 ;
  assign y29640 = ~n39198 ;
  assign y29641 = 1'b0 ;
  assign y29642 = ~n39199 ;
  assign y29643 = n39200 ;
  assign y29644 = ~n39201 ;
  assign y29645 = n39204 ;
  assign y29646 = ~1'b0 ;
  assign y29647 = ~n39205 ;
  assign y29648 = n39206 ;
  assign y29649 = n39207 ;
  assign y29650 = ~n27313 ;
  assign y29651 = n39209 ;
  assign y29652 = ~n1620 ;
  assign y29653 = ~n39212 ;
  assign y29654 = ~1'b0 ;
  assign y29655 = ~1'b0 ;
  assign y29656 = n17973 ;
  assign y29657 = n39213 ;
  assign y29658 = ~n310 ;
  assign y29659 = ~1'b0 ;
  assign y29660 = ~n39218 ;
  assign y29661 = ~n39220 ;
  assign y29662 = ~1'b0 ;
  assign y29663 = ~n7590 ;
  assign y29664 = ~n39221 ;
  assign y29665 = ~1'b0 ;
  assign y29666 = ~1'b0 ;
  assign y29667 = ~1'b0 ;
  assign y29668 = n39223 ;
  assign y29669 = ~1'b0 ;
  assign y29670 = n39224 ;
  assign y29671 = ~1'b0 ;
  assign y29672 = ~1'b0 ;
  assign y29673 = n39225 ;
  assign y29674 = n39226 ;
  assign y29675 = n39231 ;
  assign y29676 = n39235 ;
  assign y29677 = 1'b0 ;
  assign y29678 = ~1'b0 ;
  assign y29679 = ~n39236 ;
  assign y29680 = ~1'b0 ;
  assign y29681 = ~n39237 ;
  assign y29682 = n4883 ;
  assign y29683 = n39238 ;
  assign y29684 = n3446 ;
  assign y29685 = ~n39241 ;
  assign y29686 = n39245 ;
  assign y29687 = ~1'b0 ;
  assign y29688 = ~1'b0 ;
  assign y29689 = n37300 ;
  assign y29690 = ~n16270 ;
  assign y29691 = ~n39246 ;
  assign y29692 = ~1'b0 ;
  assign y29693 = ~n39248 ;
  assign y29694 = ~1'b0 ;
  assign y29695 = n39251 ;
  assign y29696 = ~1'b0 ;
  assign y29697 = ~n5933 ;
  assign y29698 = ~1'b0 ;
  assign y29699 = n39253 ;
  assign y29700 = ~n39254 ;
  assign y29701 = ~1'b0 ;
  assign y29702 = ~1'b0 ;
  assign y29703 = ~n39259 ;
  assign y29704 = ~n39260 ;
  assign y29705 = n39261 ;
  assign y29706 = n39263 ;
  assign y29707 = ~n5534 ;
  assign y29708 = n39268 ;
  assign y29709 = n39269 ;
  assign y29710 = ~n39273 ;
  assign y29711 = ~1'b0 ;
  assign y29712 = ~1'b0 ;
  assign y29713 = n39274 ;
  assign y29714 = n39277 ;
  assign y29715 = ~n39278 ;
  assign y29716 = n14647 ;
  assign y29717 = ~n39280 ;
  assign y29718 = ~n39281 ;
  assign y29719 = ~1'b0 ;
  assign y29720 = ~n39285 ;
  assign y29721 = ~n39288 ;
  assign y29722 = ~1'b0 ;
  assign y29723 = n39289 ;
  assign y29724 = n39290 ;
  assign y29725 = ~n39296 ;
  assign y29726 = ~1'b0 ;
  assign y29727 = n39297 ;
  assign y29728 = ~1'b0 ;
  assign y29729 = n39298 ;
  assign y29730 = n39300 ;
  assign y29731 = n39303 ;
  assign y29732 = n39305 ;
  assign y29733 = n39307 ;
  assign y29734 = ~1'b0 ;
  assign y29735 = n39308 ;
  assign y29736 = 1'b0 ;
  assign y29737 = ~1'b0 ;
  assign y29738 = ~1'b0 ;
  assign y29739 = n20030 ;
  assign y29740 = n39309 ;
  assign y29741 = ~n39310 ;
  assign y29742 = n39313 ;
  assign y29743 = n39314 ;
  assign y29744 = ~1'b0 ;
  assign y29745 = n16619 ;
  assign y29746 = ~n39317 ;
  assign y29747 = ~n3593 ;
  assign y29748 = ~1'b0 ;
  assign y29749 = 1'b0 ;
  assign y29750 = n2889 ;
  assign y29751 = ~1'b0 ;
  assign y29752 = ~n39318 ;
  assign y29753 = n14460 ;
  assign y29754 = n39319 ;
  assign y29755 = ~n7948 ;
  assign y29756 = ~1'b0 ;
  assign y29757 = n39321 ;
  assign y29758 = 1'b0 ;
  assign y29759 = ~1'b0 ;
  assign y29760 = ~n39322 ;
  assign y29761 = ~1'b0 ;
  assign y29762 = ~1'b0 ;
  assign y29763 = ~1'b0 ;
  assign y29764 = 1'b0 ;
  assign y29765 = ~1'b0 ;
  assign y29766 = ~n39323 ;
  assign y29767 = ~1'b0 ;
  assign y29768 = ~1'b0 ;
  assign y29769 = ~n39327 ;
  assign y29770 = n39332 ;
  assign y29771 = ~1'b0 ;
  assign y29772 = ~1'b0 ;
  assign y29773 = ~1'b0 ;
  assign y29774 = ~n39336 ;
  assign y29775 = n39337 ;
  assign y29776 = ~n39338 ;
  assign y29777 = ~n39342 ;
  assign y29778 = ~1'b0 ;
  assign y29779 = n8011 ;
  assign y29780 = ~n22185 ;
  assign y29781 = ~1'b0 ;
  assign y29782 = 1'b0 ;
  assign y29783 = ~n39345 ;
  assign y29784 = n39347 ;
  assign y29785 = ~1'b0 ;
  assign y29786 = ~1'b0 ;
  assign y29787 = ~1'b0 ;
  assign y29788 = ~n39350 ;
  assign y29789 = 1'b0 ;
  assign y29790 = ~1'b0 ;
  assign y29791 = n25094 ;
  assign y29792 = ~n39353 ;
  assign y29793 = ~n39354 ;
  assign y29794 = ~n39355 ;
  assign y29795 = 1'b0 ;
  assign y29796 = ~1'b0 ;
  assign y29797 = ~1'b0 ;
  assign y29798 = n39357 ;
  assign y29799 = ~n22218 ;
  assign y29800 = ~1'b0 ;
  assign y29801 = ~1'b0 ;
  assign y29802 = n39358 ;
  assign y29803 = ~1'b0 ;
  assign y29804 = n19724 ;
  assign y29805 = ~n39359 ;
  assign y29806 = ~1'b0 ;
  assign y29807 = n39360 ;
  assign y29808 = ~1'b0 ;
  assign y29809 = ~1'b0 ;
  assign y29810 = n23318 ;
  assign y29811 = n39362 ;
  assign y29812 = ~1'b0 ;
  assign y29813 = ~n36446 ;
  assign y29814 = n22353 ;
  assign y29815 = n39364 ;
  assign y29816 = ~n39368 ;
  assign y29817 = ~1'b0 ;
  assign y29818 = n39370 ;
  assign y29819 = ~1'b0 ;
  assign y29820 = n39372 ;
  assign y29821 = ~n39378 ;
  assign y29822 = n39380 ;
  assign y29823 = n39384 ;
  assign y29824 = ~1'b0 ;
  assign y29825 = n39386 ;
  assign y29826 = ~n39391 ;
  assign y29827 = ~1'b0 ;
  assign y29828 = n28198 ;
  assign y29829 = ~n39392 ;
  assign y29830 = ~n39394 ;
  assign y29831 = ~n39397 ;
  assign y29832 = ~1'b0 ;
  assign y29833 = ~n39399 ;
  assign y29834 = ~1'b0 ;
  assign y29835 = ~1'b0 ;
  assign y29836 = n39404 ;
  assign y29837 = ~1'b0 ;
  assign y29838 = ~n39410 ;
  assign y29839 = n39411 ;
  assign y29840 = ~1'b0 ;
  assign y29841 = n39413 ;
  assign y29842 = ~n39416 ;
  assign y29843 = n39418 ;
  assign y29844 = 1'b0 ;
  assign y29845 = ~1'b0 ;
  assign y29846 = ~n39420 ;
  assign y29847 = ~n6096 ;
  assign y29848 = ~1'b0 ;
  assign y29849 = n39421 ;
  assign y29850 = ~1'b0 ;
  assign y29851 = ~1'b0 ;
  assign y29852 = ~1'b0 ;
  assign y29853 = n39424 ;
  assign y29854 = ~1'b0 ;
  assign y29855 = n39425 ;
  assign y29856 = ~1'b0 ;
  assign y29857 = 1'b0 ;
  assign y29858 = n39430 ;
  assign y29859 = n39431 ;
  assign y29860 = ~1'b0 ;
  assign y29861 = ~n39432 ;
  assign y29862 = ~1'b0 ;
  assign y29863 = ~1'b0 ;
  assign y29864 = ~1'b0 ;
  assign y29865 = ~1'b0 ;
  assign y29866 = n16151 ;
  assign y29867 = n39433 ;
  assign y29868 = n26142 ;
  assign y29869 = ~n39435 ;
  assign y29870 = ~1'b0 ;
  assign y29871 = n39439 ;
  assign y29872 = ~n39440 ;
  assign y29873 = n39445 ;
  assign y29874 = ~1'b0 ;
  assign y29875 = ~1'b0 ;
  assign y29876 = n17755 ;
  assign y29877 = n39446 ;
  assign y29878 = n39447 ;
  assign y29879 = ~1'b0 ;
  assign y29880 = ~1'b0 ;
  assign y29881 = n39448 ;
  assign y29882 = n39451 ;
  assign y29883 = ~1'b0 ;
  assign y29884 = ~1'b0 ;
  assign y29885 = ~1'b0 ;
  assign y29886 = ~n24036 ;
  assign y29887 = ~1'b0 ;
  assign y29888 = ~n39455 ;
  assign y29889 = n39457 ;
  assign y29890 = n39462 ;
  assign y29891 = ~n39463 ;
  assign y29892 = ~1'b0 ;
  assign y29893 = ~1'b0 ;
  assign y29894 = n39464 ;
  assign y29895 = n39466 ;
  assign y29896 = ~1'b0 ;
  assign y29897 = ~1'b0 ;
  assign y29898 = ~n39468 ;
  assign y29899 = n39470 ;
  assign y29900 = n39473 ;
  assign y29901 = ~1'b0 ;
  assign y29902 = ~1'b0 ;
  assign y29903 = ~1'b0 ;
  assign y29904 = n39475 ;
  assign y29905 = ~1'b0 ;
  assign y29906 = n33906 ;
  assign y29907 = ~n39476 ;
  assign y29908 = 1'b0 ;
  assign y29909 = ~n39478 ;
  assign y29910 = ~n39479 ;
  assign y29911 = ~n39482 ;
  assign y29912 = n31695 ;
  assign y29913 = ~1'b0 ;
  assign y29914 = ~n39486 ;
  assign y29915 = ~1'b0 ;
  assign y29916 = ~1'b0 ;
  assign y29917 = ~1'b0 ;
  assign y29918 = n39487 ;
  assign y29919 = n39489 ;
  assign y29920 = n39490 ;
  assign y29921 = ~1'b0 ;
  assign y29922 = ~1'b0 ;
  assign y29923 = ~n39491 ;
  assign y29924 = ~n39492 ;
  assign y29925 = n39495 ;
  assign y29926 = n39496 ;
  assign y29927 = n39499 ;
  assign y29928 = ~n39502 ;
  assign y29929 = 1'b0 ;
  assign y29930 = n39503 ;
  assign y29931 = ~n39505 ;
  assign y29932 = ~n19041 ;
  assign y29933 = n39507 ;
  assign y29934 = ~1'b0 ;
  assign y29935 = ~1'b0 ;
  assign y29936 = n39508 ;
  assign y29937 = ~1'b0 ;
  assign y29938 = 1'b0 ;
  assign y29939 = ~1'b0 ;
  assign y29940 = ~1'b0 ;
  assign y29941 = n39511 ;
  assign y29942 = n30480 ;
  assign y29943 = n39512 ;
  assign y29944 = ~n39516 ;
  assign y29945 = n19733 ;
  assign y29946 = ~n39518 ;
  assign y29947 = n39519 ;
  assign y29948 = n39520 ;
  assign y29949 = ~n39523 ;
  assign y29950 = ~1'b0 ;
  assign y29951 = ~1'b0 ;
  assign y29952 = ~n39526 ;
  assign y29953 = ~n39530 ;
  assign y29954 = n39532 ;
  assign y29955 = ~1'b0 ;
  assign y29956 = ~n39535 ;
  assign y29957 = ~1'b0 ;
  assign y29958 = ~1'b0 ;
  assign y29959 = n39536 ;
  assign y29960 = ~n39540 ;
  assign y29961 = ~1'b0 ;
  assign y29962 = ~1'b0 ;
  assign y29963 = ~n39541 ;
  assign y29964 = ~n39544 ;
  assign y29965 = ~n39549 ;
  assign y29966 = ~n39550 ;
  assign y29967 = ~1'b0 ;
  assign y29968 = ~1'b0 ;
  assign y29969 = ~n595 ;
  assign y29970 = n39551 ;
  assign y29971 = n39555 ;
  assign y29972 = ~1'b0 ;
  assign y29973 = ~n39558 ;
  assign y29974 = n39560 ;
  assign y29975 = ~n39564 ;
  assign y29976 = n39565 ;
  assign y29977 = ~1'b0 ;
  assign y29978 = ~1'b0 ;
  assign y29979 = ~1'b0 ;
  assign y29980 = n39574 ;
  assign y29981 = ~n11735 ;
  assign y29982 = 1'b0 ;
  assign y29983 = ~n10228 ;
  assign y29984 = n39578 ;
  assign y29985 = ~1'b0 ;
  assign y29986 = ~1'b0 ;
  assign y29987 = ~1'b0 ;
  assign y29988 = ~1'b0 ;
  assign y29989 = ~1'b0 ;
  assign y29990 = ~1'b0 ;
  assign y29991 = ~n39581 ;
  assign y29992 = ~n39583 ;
  assign y29993 = n39584 ;
  assign y29994 = ~1'b0 ;
  assign y29995 = ~n8452 ;
  assign y29996 = n39585 ;
  assign y29997 = ~1'b0 ;
  assign y29998 = ~n29694 ;
  assign y29999 = n39587 ;
  assign y30000 = 1'b0 ;
  assign y30001 = n34432 ;
  assign y30002 = ~n39592 ;
  assign y30003 = n39594 ;
  assign y30004 = ~n39596 ;
  assign y30005 = ~1'b0 ;
  assign y30006 = ~n2185 ;
  assign y30007 = ~n39597 ;
  assign y30008 = ~1'b0 ;
  assign y30009 = n17259 ;
  assign y30010 = ~1'b0 ;
  assign y30011 = ~1'b0 ;
  assign y30012 = ~1'b0 ;
  assign y30013 = ~n39598 ;
  assign y30014 = ~n39606 ;
  assign y30015 = n39608 ;
  assign y30016 = ~1'b0 ;
  assign y30017 = ~n39609 ;
  assign y30018 = n39610 ;
  assign y30019 = n39616 ;
  assign y30020 = ~n39618 ;
  assign y30021 = ~1'b0 ;
  assign y30022 = n39619 ;
  assign y30023 = ~n39620 ;
  assign y30024 = ~1'b0 ;
  assign y30025 = ~n39626 ;
  assign y30026 = n31730 ;
  assign y30027 = ~1'b0 ;
  assign y30028 = n39627 ;
  assign y30029 = ~n39628 ;
  assign y30030 = 1'b0 ;
  assign y30031 = ~1'b0 ;
  assign y30032 = n39631 ;
  assign y30033 = ~n39632 ;
  assign y30034 = ~n32622 ;
  assign y30035 = ~1'b0 ;
  assign y30036 = n39633 ;
  assign y30037 = n2148 ;
  assign y30038 = n28804 ;
  assign y30039 = ~n39634 ;
  assign y30040 = ~1'b0 ;
  assign y30041 = n39635 ;
  assign y30042 = n39636 ;
  assign y30043 = ~1'b0 ;
  assign y30044 = n39637 ;
  assign y30045 = ~1'b0 ;
  assign y30046 = n39641 ;
  assign y30047 = n11127 ;
  assign y30048 = ~1'b0 ;
  assign y30049 = ~1'b0 ;
  assign y30050 = ~n39642 ;
  assign y30051 = ~n39643 ;
  assign y30052 = ~1'b0 ;
  assign y30053 = ~1'b0 ;
  assign y30054 = n39644 ;
  assign y30055 = ~n39645 ;
  assign y30056 = ~n10822 ;
  assign y30057 = ~1'b0 ;
  assign y30058 = ~1'b0 ;
  assign y30059 = n39647 ;
  assign y30060 = ~n39651 ;
  assign y30061 = ~n39653 ;
  assign y30062 = n39655 ;
  assign y30063 = ~1'b0 ;
  assign y30064 = ~n39658 ;
  assign y30065 = ~n9024 ;
  assign y30066 = ~1'b0 ;
  assign y30067 = n39659 ;
  assign y30068 = ~n39660 ;
  assign y30069 = ~1'b0 ;
  assign y30070 = n39662 ;
  assign y30071 = n39672 ;
  assign y30072 = n39673 ;
  assign y30073 = ~1'b0 ;
  assign y30074 = ~1'b0 ;
  assign y30075 = ~n39675 ;
  assign y30076 = ~1'b0 ;
  assign y30077 = n609 ;
  assign y30078 = ~n5826 ;
  assign y30079 = ~n39676 ;
  assign y30080 = ~n9083 ;
  assign y30081 = ~n39677 ;
  assign y30082 = ~n39678 ;
  assign y30083 = ~1'b0 ;
  assign y30084 = ~n39680 ;
  assign y30085 = ~1'b0 ;
  assign y30086 = ~1'b0 ;
  assign y30087 = n10271 ;
  assign y30088 = ~1'b0 ;
  assign y30089 = n39681 ;
  assign y30090 = n39682 ;
  assign y30091 = n39683 ;
  assign y30092 = ~n39685 ;
  assign y30093 = n39687 ;
  assign y30094 = n39688 ;
  assign y30095 = ~1'b0 ;
  assign y30096 = n19138 ;
  assign y30097 = ~n39690 ;
  assign y30098 = n39692 ;
  assign y30099 = ~n39693 ;
  assign y30100 = ~1'b0 ;
  assign y30101 = ~1'b0 ;
  assign y30102 = ~n39694 ;
  assign y30103 = ~1'b0 ;
  assign y30104 = ~n39695 ;
  assign y30105 = n39698 ;
  assign y30106 = ~n5541 ;
  assign y30107 = n39699 ;
  assign y30108 = ~1'b0 ;
  assign y30109 = ~n39700 ;
  assign y30110 = n39704 ;
  assign y30111 = ~1'b0 ;
  assign y30112 = ~n39707 ;
  assign y30113 = n2245 ;
  assign y30114 = ~n39708 ;
  assign y30115 = n39709 ;
  assign y30116 = ~1'b0 ;
  assign y30117 = n39710 ;
  assign y30118 = ~1'b0 ;
  assign y30119 = ~n39711 ;
  assign y30120 = n39716 ;
  assign y30121 = n39717 ;
  assign y30122 = 1'b0 ;
  assign y30123 = ~1'b0 ;
  assign y30124 = ~n28732 ;
  assign y30125 = ~1'b0 ;
  assign y30126 = n39720 ;
  assign y30127 = n39724 ;
  assign y30128 = n39726 ;
  assign y30129 = ~1'b0 ;
  assign y30130 = ~1'b0 ;
  assign y30131 = ~n39730 ;
  assign y30132 = n39732 ;
  assign y30133 = ~1'b0 ;
  assign y30134 = n39734 ;
  assign y30135 = ~n10177 ;
  assign y30136 = n36714 ;
  assign y30137 = ~n39735 ;
  assign y30138 = ~1'b0 ;
  assign y30139 = ~1'b0 ;
  assign y30140 = n39737 ;
  assign y30141 = n39744 ;
  assign y30142 = n39745 ;
  assign y30143 = ~1'b0 ;
  assign y30144 = ~n39747 ;
  assign y30145 = n31999 ;
  assign y30146 = n31617 ;
  assign y30147 = ~1'b0 ;
  assign y30148 = ~1'b0 ;
  assign y30149 = n39751 ;
  assign y30150 = ~n39753 ;
  assign y30151 = ~n39756 ;
  assign y30152 = ~n39758 ;
  assign y30153 = ~n29973 ;
  assign y30154 = ~1'b0 ;
  assign y30155 = ~n39765 ;
  assign y30156 = n39768 ;
  assign y30157 = ~n39773 ;
  assign y30158 = ~1'b0 ;
  assign y30159 = n11047 ;
  assign y30160 = ~n39774 ;
  assign y30161 = ~1'b0 ;
  assign y30162 = ~1'b0 ;
  assign y30163 = ~1'b0 ;
  assign y30164 = ~1'b0 ;
  assign y30165 = ~n39777 ;
  assign y30166 = n39778 ;
  assign y30167 = n39781 ;
  assign y30168 = n39783 ;
  assign y30169 = ~n31748 ;
  assign y30170 = ~n14417 ;
  assign y30171 = n39784 ;
  assign y30172 = n7109 ;
  assign y30173 = n39787 ;
  assign y30174 = ~1'b0 ;
  assign y30175 = ~n39788 ;
  assign y30176 = n39789 ;
  assign y30177 = ~n39790 ;
  assign y30178 = n39792 ;
  assign y30179 = ~1'b0 ;
  assign y30180 = ~n39794 ;
  assign y30181 = ~n39798 ;
  assign y30182 = ~1'b0 ;
  assign y30183 = n39800 ;
  assign y30184 = n39801 ;
  assign y30185 = ~n39802 ;
  assign y30186 = ~n39803 ;
  assign y30187 = ~n39805 ;
  assign y30188 = 1'b0 ;
  assign y30189 = n39807 ;
  assign y30190 = n39809 ;
  assign y30191 = n17266 ;
  assign y30192 = 1'b0 ;
  assign y30193 = ~n39812 ;
  assign y30194 = ~n39814 ;
  assign y30195 = ~1'b0 ;
  assign y30196 = ~1'b0 ;
  assign y30197 = ~1'b0 ;
  assign y30198 = ~1'b0 ;
  assign y30199 = ~n39816 ;
  assign y30200 = ~n39817 ;
  assign y30201 = ~1'b0 ;
  assign y30202 = ~1'b0 ;
  assign y30203 = ~n39819 ;
  assign y30204 = ~n39820 ;
  assign y30205 = ~1'b0 ;
  assign y30206 = ~1'b0 ;
  assign y30207 = n39822 ;
  assign y30208 = ~n39823 ;
  assign y30209 = ~n39825 ;
  assign y30210 = ~n15672 ;
  assign y30211 = ~n39827 ;
  assign y30212 = n39832 ;
  assign y30213 = ~n39835 ;
  assign y30214 = ~1'b0 ;
  assign y30215 = ~1'b0 ;
  assign y30216 = ~1'b0 ;
  assign y30217 = ~1'b0 ;
  assign y30218 = ~1'b0 ;
  assign y30219 = n39839 ;
  assign y30220 = n10680 ;
  assign y30221 = 1'b0 ;
  assign y30222 = ~n3452 ;
  assign y30223 = ~1'b0 ;
  assign y30224 = ~n39840 ;
  assign y30225 = n12974 ;
  assign y30226 = ~1'b0 ;
  assign y30227 = n39841 ;
  assign y30228 = ~n977 ;
  assign y30229 = n39842 ;
  assign y30230 = ~1'b0 ;
  assign y30231 = n39844 ;
  assign y30232 = ~n39848 ;
  assign y30233 = ~n31779 ;
  assign y30234 = n39849 ;
  assign y30235 = ~1'b0 ;
  assign y30236 = ~1'b0 ;
  assign y30237 = n39850 ;
  assign y30238 = ~1'b0 ;
  assign y30239 = ~n39852 ;
  assign y30240 = ~1'b0 ;
  assign y30241 = n8358 ;
  assign y30242 = ~1'b0 ;
  assign y30243 = ~n39853 ;
  assign y30244 = ~n39856 ;
  assign y30245 = n39857 ;
  assign y30246 = ~1'b0 ;
  assign y30247 = ~n39858 ;
  assign y30248 = n39862 ;
  assign y30249 = 1'b0 ;
  assign y30250 = n39866 ;
  assign y30251 = ~n39540 ;
  assign y30252 = ~n39867 ;
  assign y30253 = ~1'b0 ;
  assign y30254 = ~1'b0 ;
  assign y30255 = ~1'b0 ;
  assign y30256 = ~1'b0 ;
  assign y30257 = n39869 ;
  assign y30258 = n39870 ;
  assign y30259 = ~n39883 ;
  assign y30260 = ~n39885 ;
  assign y30261 = ~n39887 ;
  assign y30262 = ~n39889 ;
  assign y30263 = ~n39893 ;
  assign y30264 = ~1'b0 ;
  assign y30265 = ~n39895 ;
  assign y30266 = ~1'b0 ;
  assign y30267 = ~n39898 ;
  assign y30268 = n39900 ;
  assign y30269 = n37484 ;
  assign y30270 = n21648 ;
  assign y30271 = n39902 ;
  assign y30272 = n39903 ;
  assign y30273 = ~n39905 ;
  assign y30274 = n39907 ;
  assign y30275 = ~n39916 ;
  assign y30276 = ~1'b0 ;
  assign y30277 = ~1'b0 ;
  assign y30278 = ~1'b0 ;
  assign y30279 = ~1'b0 ;
  assign y30280 = ~1'b0 ;
  assign y30281 = 1'b0 ;
  assign y30282 = ~n39917 ;
  assign y30283 = 1'b0 ;
  assign y30284 = ~1'b0 ;
  assign y30285 = 1'b0 ;
  assign y30286 = n39922 ;
  assign y30287 = ~n39923 ;
  assign y30288 = ~1'b0 ;
  assign y30289 = ~1'b0 ;
  assign y30290 = ~1'b0 ;
  assign y30291 = n286 ;
  assign y30292 = ~1'b0 ;
  assign y30293 = ~n39925 ;
  assign y30294 = ~n39927 ;
  assign y30295 = n39928 ;
  assign y30296 = n39929 ;
  assign y30297 = n39930 ;
  assign y30298 = ~n39931 ;
  assign y30299 = n39934 ;
  assign y30300 = ~n39938 ;
  assign y30301 = n39939 ;
  assign y30302 = ~n39943 ;
  assign y30303 = n39945 ;
  assign y30304 = ~1'b0 ;
  assign y30305 = n4757 ;
  assign y30306 = ~n39946 ;
  assign y30307 = 1'b0 ;
  assign y30308 = ~n39948 ;
  assign y30309 = 1'b0 ;
  assign y30310 = n39951 ;
  assign y30311 = ~1'b0 ;
  assign y30312 = ~n39952 ;
  assign y30313 = ~1'b0 ;
  assign y30314 = ~n39954 ;
  assign y30315 = ~1'b0 ;
  assign y30316 = ~n39956 ;
  assign y30317 = ~n39957 ;
  assign y30318 = ~n39959 ;
  assign y30319 = ~1'b0 ;
  assign y30320 = n39964 ;
  assign y30321 = ~n39967 ;
  assign y30322 = ~1'b0 ;
  assign y30323 = ~n39973 ;
  assign y30324 = ~1'b0 ;
  assign y30325 = 1'b0 ;
  assign y30326 = n39974 ;
  assign y30327 = ~n39975 ;
  assign y30328 = ~n39976 ;
  assign y30329 = n39979 ;
  assign y30330 = ~1'b0 ;
  assign y30331 = n39981 ;
  assign y30332 = n39984 ;
  assign y30333 = n39987 ;
  assign y30334 = n39989 ;
  assign y30335 = n39991 ;
  assign y30336 = ~1'b0 ;
  assign y30337 = 1'b0 ;
  assign y30338 = 1'b0 ;
  assign y30339 = n2023 ;
  assign y30340 = n10887 ;
  assign y30341 = ~1'b0 ;
  assign y30342 = ~n39995 ;
  assign y30343 = ~n39998 ;
  assign y30344 = n40000 ;
  assign y30345 = n40004 ;
  assign y30346 = ~n40009 ;
  assign y30347 = n29901 ;
  assign y30348 = n40010 ;
  assign y30349 = ~n5948 ;
  assign y30350 = ~n1314 ;
  assign y30351 = ~n40011 ;
  assign y30352 = n9335 ;
  assign y30353 = n40015 ;
  assign y30354 = ~n40017 ;
  assign y30355 = ~1'b0 ;
  assign y30356 = ~n15302 ;
  assign y30357 = ~n40018 ;
  assign y30358 = n40020 ;
  assign y30359 = ~1'b0 ;
  assign y30360 = ~1'b0 ;
  assign y30361 = n40024 ;
  assign y30362 = n40027 ;
  assign y30363 = n17695 ;
  assign y30364 = ~1'b0 ;
  assign y30365 = n25310 ;
  assign y30366 = 1'b0 ;
  assign y30367 = ~n40029 ;
  assign y30368 = ~n40030 ;
  assign y30369 = ~n40033 ;
  assign y30370 = ~1'b0 ;
  assign y30371 = n40034 ;
  assign y30372 = ~1'b0 ;
  assign y30373 = ~1'b0 ;
  assign y30374 = ~n40035 ;
  assign y30375 = ~1'b0 ;
  assign y30376 = ~n33103 ;
  assign y30377 = n40036 ;
  assign y30378 = ~n40037 ;
  assign y30379 = n2148 ;
  assign y30380 = n40040 ;
  assign y30381 = ~n40042 ;
  assign y30382 = n40043 ;
  assign y30383 = n40047 ;
  assign y30384 = ~1'b0 ;
  assign y30385 = ~n20277 ;
  assign y30386 = ~n40048 ;
  assign y30387 = ~n40050 ;
  assign y30388 = ~1'b0 ;
  assign y30389 = n40053 ;
  assign y30390 = ~1'b0 ;
  assign y30391 = ~n40055 ;
  assign y30392 = ~1'b0 ;
  assign y30393 = ~n40057 ;
  assign y30394 = n40058 ;
  assign y30395 = ~1'b0 ;
  assign y30396 = ~1'b0 ;
  assign y30397 = ~1'b0 ;
  assign y30398 = 1'b0 ;
  assign y30399 = n40059 ;
  assign y30400 = n1838 ;
  assign y30401 = ~1'b0 ;
  assign y30402 = n40061 ;
  assign y30403 = ~n7455 ;
  assign y30404 = ~1'b0 ;
  assign y30405 = n40062 ;
  assign y30406 = n1143 ;
  assign y30407 = n11802 ;
  assign y30408 = n15901 ;
  assign y30409 = n40064 ;
  assign y30410 = n40067 ;
  assign y30411 = 1'b0 ;
  assign y30412 = ~n40069 ;
  assign y30413 = n40070 ;
  assign y30414 = ~n40071 ;
  assign y30415 = ~1'b0 ;
  assign y30416 = ~n40074 ;
  assign y30417 = ~1'b0 ;
  assign y30418 = n40075 ;
  assign y30419 = ~1'b0 ;
  assign y30420 = ~n40076 ;
  assign y30421 = ~n40077 ;
  assign y30422 = n2615 ;
  assign y30423 = ~1'b0 ;
  assign y30424 = ~n40078 ;
  assign y30425 = ~n12207 ;
  assign y30426 = n40081 ;
  assign y30427 = n40084 ;
  assign y30428 = ~n20450 ;
  assign y30429 = ~1'b0 ;
  assign y30430 = n40086 ;
  assign y30431 = ~n40090 ;
  assign y30432 = n40093 ;
  assign y30433 = n40095 ;
  assign y30434 = ~n40096 ;
  assign y30435 = n40099 ;
  assign y30436 = n40100 ;
  assign y30437 = 1'b0 ;
  assign y30438 = n40103 ;
  assign y30439 = ~1'b0 ;
  assign y30440 = ~1'b0 ;
  assign y30441 = n40105 ;
  assign y30442 = ~n40106 ;
  assign y30443 = n40109 ;
  assign y30444 = ~n40110 ;
  assign y30445 = n40112 ;
  assign y30446 = ~n40114 ;
  assign y30447 = n40115 ;
  assign y30448 = 1'b0 ;
  assign y30449 = n40116 ;
  assign y30450 = ~1'b0 ;
  assign y30451 = ~1'b0 ;
  assign y30452 = ~n40119 ;
  assign y30453 = ~1'b0 ;
  assign y30454 = ~1'b0 ;
  assign y30455 = ~1'b0 ;
  assign y30456 = ~n40121 ;
  assign y30457 = n40123 ;
  assign y30458 = ~n40124 ;
  assign y30459 = ~1'b0 ;
  assign y30460 = n40125 ;
  assign y30461 = n19181 ;
  assign y30462 = ~n40126 ;
  assign y30463 = ~n40127 ;
  assign y30464 = n39146 ;
  assign y30465 = ~n39994 ;
  assign y30466 = ~n40129 ;
  assign y30467 = ~1'b0 ;
  assign y30468 = ~n9002 ;
  assign y30469 = ~n40131 ;
  assign y30470 = ~n40132 ;
  assign y30471 = n6373 ;
  assign y30472 = ~1'b0 ;
  assign y30473 = n40133 ;
  assign y30474 = n40137 ;
  assign y30475 = ~n40138 ;
  assign y30476 = ~1'b0 ;
  assign y30477 = ~1'b0 ;
  assign y30478 = n40139 ;
  assign y30479 = ~n40142 ;
  assign y30480 = n40143 ;
  assign y30481 = ~n40146 ;
  assign y30482 = ~1'b0 ;
  assign y30483 = ~1'b0 ;
  assign y30484 = n40147 ;
  assign y30485 = ~1'b0 ;
  assign y30486 = ~1'b0 ;
  assign y30487 = n40152 ;
  assign y30488 = ~1'b0 ;
  assign y30489 = n40155 ;
  assign y30490 = ~n40157 ;
  assign y30491 = ~1'b0 ;
  assign y30492 = ~n40160 ;
  assign y30493 = ~1'b0 ;
  assign y30494 = ~1'b0 ;
  assign y30495 = ~n40161 ;
  assign y30496 = n40163 ;
  assign y30497 = ~1'b0 ;
  assign y30498 = ~1'b0 ;
  assign y30499 = ~n40164 ;
  assign y30500 = 1'b0 ;
  assign y30501 = ~n40166 ;
  assign y30502 = ~1'b0 ;
  assign y30503 = n40167 ;
  assign y30504 = ~1'b0 ;
  assign y30505 = n40170 ;
  assign y30506 = n40171 ;
  assign y30507 = 1'b0 ;
  assign y30508 = ~n40174 ;
  assign y30509 = n7375 ;
  assign y30510 = ~1'b0 ;
  assign y30511 = ~1'b0 ;
  assign y30512 = n22627 ;
  assign y30513 = 1'b0 ;
  assign y30514 = n40175 ;
  assign y30515 = ~n40179 ;
  assign y30516 = n5202 ;
  assign y30517 = 1'b0 ;
  assign y30518 = ~1'b0 ;
  assign y30519 = ~n40182 ;
  assign y30520 = ~1'b0 ;
  assign y30521 = n40183 ;
  assign y30522 = ~1'b0 ;
  assign y30523 = ~1'b0 ;
  assign y30524 = 1'b0 ;
  assign y30525 = n40191 ;
  assign y30526 = ~1'b0 ;
  assign y30527 = ~1'b0 ;
  assign y30528 = ~n40192 ;
  assign y30529 = ~n40194 ;
  assign y30530 = n40195 ;
  assign y30531 = ~1'b0 ;
  assign y30532 = ~1'b0 ;
  assign y30533 = ~n40197 ;
  assign y30534 = ~n40198 ;
  assign y30535 = ~n40200 ;
  assign y30536 = n40201 ;
  assign y30537 = n40203 ;
  assign y30538 = ~n40206 ;
  assign y30539 = ~n40212 ;
  assign y30540 = n40213 ;
  assign y30541 = ~1'b0 ;
  assign y30542 = n40214 ;
  assign y30543 = ~1'b0 ;
  assign y30544 = ~n40215 ;
  assign y30545 = ~n40217 ;
  assign y30546 = ~1'b0 ;
  assign y30547 = ~1'b0 ;
  assign y30548 = ~1'b0 ;
  assign y30549 = n40218 ;
  assign y30550 = ~1'b0 ;
  assign y30551 = ~1'b0 ;
  assign y30552 = ~1'b0 ;
  assign y30553 = n40220 ;
  assign y30554 = ~1'b0 ;
  assign y30555 = ~n40222 ;
  assign y30556 = ~1'b0 ;
  assign y30557 = ~1'b0 ;
  assign y30558 = ~n40224 ;
  assign y30559 = ~n40225 ;
  assign y30560 = ~n40226 ;
  assign y30561 = ~n17068 ;
  assign y30562 = ~n40232 ;
  assign y30563 = ~n40234 ;
  assign y30564 = ~n40237 ;
  assign y30565 = ~n9531 ;
  assign y30566 = ~1'b0 ;
  assign y30567 = ~1'b0 ;
  assign y30568 = ~1'b0 ;
  assign y30569 = ~n40239 ;
  assign y30570 = n40240 ;
  assign y30571 = n40243 ;
  assign y30572 = ~1'b0 ;
  assign y30573 = n40245 ;
  assign y30574 = ~1'b0 ;
  assign y30575 = ~n40246 ;
  assign y30576 = n40247 ;
  assign y30577 = ~1'b0 ;
  assign y30578 = ~n40248 ;
  assign y30579 = ~1'b0 ;
  assign y30580 = n40250 ;
  assign y30581 = n40252 ;
  assign y30582 = n15166 ;
  assign y30583 = ~n40256 ;
  assign y30584 = n40257 ;
  assign y30585 = ~n40258 ;
  assign y30586 = ~1'b0 ;
  assign y30587 = ~1'b0 ;
  assign y30588 = ~1'b0 ;
  assign y30589 = ~1'b0 ;
  assign y30590 = ~1'b0 ;
  assign y30591 = ~n40262 ;
  assign y30592 = n40264 ;
  assign y30593 = ~n40267 ;
  assign y30594 = n40269 ;
  assign y30595 = ~n40270 ;
  assign y30596 = ~n40272 ;
  assign y30597 = ~n40275 ;
  assign y30598 = ~1'b0 ;
  assign y30599 = ~n21651 ;
  assign y30600 = 1'b0 ;
  assign y30601 = ~n40277 ;
  assign y30602 = ~n40280 ;
  assign y30603 = n17895 ;
  assign y30604 = n7394 ;
  assign y30605 = ~n40282 ;
  assign y30606 = ~n40283 ;
  assign y30607 = ~n40284 ;
  assign y30608 = ~1'b0 ;
  assign y30609 = ~n40285 ;
  assign y30610 = ~1'b0 ;
  assign y30611 = n40286 ;
  assign y30612 = ~n40287 ;
  assign y30613 = ~n40288 ;
  assign y30614 = n40289 ;
  assign y30615 = ~n1631 ;
  assign y30616 = ~1'b0 ;
  assign y30617 = ~1'b0 ;
  assign y30618 = n40291 ;
  assign y30619 = ~n40293 ;
  assign y30620 = ~n90 ;
  assign y30621 = ~1'b0 ;
  assign y30622 = n40295 ;
  assign y30623 = ~n40298 ;
  assign y30624 = 1'b0 ;
  assign y30625 = ~n40300 ;
  assign y30626 = ~1'b0 ;
  assign y30627 = ~1'b0 ;
  assign y30628 = ~n40301 ;
  assign y30629 = 1'b0 ;
  assign y30630 = n40303 ;
  assign y30631 = ~1'b0 ;
  assign y30632 = ~n40306 ;
  assign y30633 = n40310 ;
  assign y30634 = ~n31019 ;
  assign y30635 = x3 ;
  assign y30636 = ~1'b0 ;
  assign y30637 = ~1'b0 ;
  assign y30638 = ~1'b0 ;
  assign y30639 = ~1'b0 ;
  assign y30640 = ~1'b0 ;
  assign y30641 = ~1'b0 ;
  assign y30642 = n40312 ;
  assign y30643 = 1'b0 ;
  assign y30644 = n40313 ;
  assign y30645 = ~1'b0 ;
  assign y30646 = n40314 ;
  assign y30647 = ~1'b0 ;
  assign y30648 = ~1'b0 ;
  assign y30649 = ~1'b0 ;
  assign y30650 = ~n40315 ;
  assign y30651 = ~1'b0 ;
  assign y30652 = ~n40318 ;
  assign y30653 = n40319 ;
  assign y30654 = n15439 ;
  assign y30655 = ~1'b0 ;
  assign y30656 = ~1'b0 ;
  assign y30657 = n40322 ;
  assign y30658 = ~n40324 ;
  assign y30659 = ~1'b0 ;
  assign y30660 = ~n40325 ;
  assign y30661 = ~1'b0 ;
  assign y30662 = ~1'b0 ;
  assign y30663 = 1'b0 ;
  assign y30664 = ~n40331 ;
  assign y30665 = ~1'b0 ;
  assign y30666 = ~n2311 ;
  assign y30667 = ~1'b0 ;
  assign y30668 = ~n3022 ;
  assign y30669 = ~1'b0 ;
  assign y30670 = n40332 ;
  assign y30671 = n40334 ;
  assign y30672 = n21479 ;
  assign y30673 = n40336 ;
  assign y30674 = n40337 ;
  assign y30675 = n40338 ;
  assign y30676 = 1'b0 ;
  assign y30677 = ~1'b0 ;
  assign y30678 = ~1'b0 ;
  assign y30679 = n40341 ;
  assign y30680 = ~1'b0 ;
  assign y30681 = ~1'b0 ;
  assign y30682 = ~n40342 ;
  assign y30683 = ~1'b0 ;
  assign y30684 = n40343 ;
  assign y30685 = ~n40344 ;
  assign y30686 = n40346 ;
  assign y30687 = ~1'b0 ;
  assign y30688 = ~1'b0 ;
  assign y30689 = ~1'b0 ;
  assign y30690 = n40348 ;
  assign y30691 = n40349 ;
  assign y30692 = n24667 ;
  assign y30693 = ~1'b0 ;
  assign y30694 = ~n40351 ;
  assign y30695 = n21498 ;
  assign y30696 = n507 ;
  assign y30697 = ~n40352 ;
  assign y30698 = ~n40354 ;
  assign y30699 = ~1'b0 ;
  assign y30700 = ~n40355 ;
  assign y30701 = ~n15536 ;
  assign y30702 = ~1'b0 ;
  assign y30703 = ~n40358 ;
  assign y30704 = n1875 ;
  assign y30705 = ~1'b0 ;
  assign y30706 = ~1'b0 ;
  assign y30707 = ~n19879 ;
  assign y30708 = ~n40360 ;
  assign y30709 = ~n40364 ;
  assign y30710 = ~1'b0 ;
  assign y30711 = ~n40369 ;
  assign y30712 = n38574 ;
  assign y30713 = ~1'b0 ;
  assign y30714 = ~1'b0 ;
  assign y30715 = n40372 ;
  assign y30716 = n40375 ;
  assign y30717 = ~1'b0 ;
  assign y30718 = ~n40376 ;
  assign y30719 = n1856 ;
  assign y30720 = ~1'b0 ;
  assign y30721 = n39253 ;
  assign y30722 = ~1'b0 ;
  assign y30723 = ~n37976 ;
  assign y30724 = n40378 ;
  assign y30725 = ~n40380 ;
  assign y30726 = n40381 ;
  assign y30727 = ~1'b0 ;
  assign y30728 = n40382 ;
  assign y30729 = ~n40383 ;
  assign y30730 = ~1'b0 ;
  assign y30731 = ~1'b0 ;
  assign y30732 = ~1'b0 ;
  assign y30733 = ~1'b0 ;
  assign y30734 = n40385 ;
  assign y30735 = n40388 ;
  assign y30736 = n40392 ;
  assign y30737 = ~n40396 ;
  assign y30738 = ~1'b0 ;
  assign y30739 = ~1'b0 ;
  assign y30740 = ~n40401 ;
  assign y30741 = ~1'b0 ;
  assign y30742 = n40405 ;
  assign y30743 = n29515 ;
  assign y30744 = ~n39150 ;
  assign y30745 = ~n40411 ;
  assign y30746 = ~n40412 ;
  assign y30747 = ~1'b0 ;
  assign y30748 = n40413 ;
  assign y30749 = ~1'b0 ;
  assign y30750 = 1'b0 ;
  assign y30751 = n40416 ;
  assign y30752 = ~n40419 ;
  assign y30753 = ~n40420 ;
  assign y30754 = ~n40422 ;
  assign y30755 = 1'b0 ;
  assign y30756 = ~1'b0 ;
  assign y30757 = ~1'b0 ;
  assign y30758 = ~n40424 ;
  assign y30759 = 1'b0 ;
  assign y30760 = ~1'b0 ;
  assign y30761 = 1'b0 ;
  assign y30762 = ~1'b0 ;
  assign y30763 = n40425 ;
  assign y30764 = ~1'b0 ;
  assign y30765 = ~1'b0 ;
  assign y30766 = ~1'b0 ;
  assign y30767 = ~n1056 ;
  assign y30768 = ~1'b0 ;
  assign y30769 = ~n40426 ;
  assign y30770 = ~1'b0 ;
  assign y30771 = 1'b0 ;
  assign y30772 = ~1'b0 ;
  assign y30773 = ~1'b0 ;
  assign y30774 = ~n40428 ;
  assign y30775 = ~1'b0 ;
  assign y30776 = n40431 ;
  assign y30777 = ~1'b0 ;
  assign y30778 = n40432 ;
  assign y30779 = n40433 ;
  assign y30780 = ~n40436 ;
  assign y30781 = ~1'b0 ;
  assign y30782 = ~n40439 ;
  assign y30783 = ~n40442 ;
  assign y30784 = ~1'b0 ;
  assign y30785 = ~1'b0 ;
  assign y30786 = ~n40444 ;
  assign y30787 = n40447 ;
  assign y30788 = ~1'b0 ;
  assign y30789 = ~n40448 ;
  assign y30790 = n40452 ;
  assign y30791 = ~n17354 ;
  assign y30792 = ~n40455 ;
  assign y30793 = n40457 ;
  assign y30794 = n40460 ;
  assign y30795 = ~n40467 ;
  assign y30796 = ~1'b0 ;
  assign y30797 = ~n40468 ;
  assign y30798 = ~n40471 ;
  assign y30799 = ~n40473 ;
  assign y30800 = ~1'b0 ;
  assign y30801 = 1'b0 ;
  assign y30802 = ~n40479 ;
  assign y30803 = n40483 ;
  assign y30804 = ~n40485 ;
  assign y30805 = ~n40486 ;
  assign y30806 = n40487 ;
  assign y30807 = ~1'b0 ;
  assign y30808 = n40488 ;
  assign y30809 = ~n40489 ;
  assign y30810 = ~1'b0 ;
  assign y30811 = ~1'b0 ;
  assign y30812 = ~n18532 ;
  assign y30813 = n40496 ;
  assign y30814 = ~1'b0 ;
  assign y30815 = ~n40497 ;
  assign y30816 = ~n40498 ;
  assign y30817 = ~1'b0 ;
  assign y30818 = n40501 ;
  assign y30819 = n40504 ;
  assign y30820 = ~1'b0 ;
  assign y30821 = ~n40505 ;
  assign y30822 = n40507 ;
  assign y30823 = 1'b0 ;
  assign y30824 = n20897 ;
  assign y30825 = n40508 ;
  assign y30826 = ~n40511 ;
  assign y30827 = ~n40512 ;
  assign y30828 = ~n40514 ;
  assign y30829 = n40516 ;
  assign y30830 = ~n40522 ;
  assign y30831 = ~1'b0 ;
  assign y30832 = ~1'b0 ;
  assign y30833 = ~1'b0 ;
  assign y30834 = n40526 ;
  assign y30835 = n40527 ;
  assign y30836 = ~1'b0 ;
  assign y30837 = ~n40532 ;
  assign y30838 = n40536 ;
  assign y30839 = 1'b0 ;
  assign y30840 = ~n40538 ;
  assign y30841 = ~1'b0 ;
  assign y30842 = ~n40540 ;
  assign y30843 = 1'b0 ;
  assign y30844 = ~1'b0 ;
  assign y30845 = n40547 ;
  assign y30846 = n40548 ;
  assign y30847 = ~n40552 ;
  assign y30848 = ~1'b0 ;
  assign y30849 = ~1'b0 ;
  assign y30850 = ~1'b0 ;
  assign y30851 = n40553 ;
  assign y30852 = ~n40554 ;
  assign y30853 = n40556 ;
  assign y30854 = ~1'b0 ;
  assign y30855 = ~n40557 ;
  assign y30856 = ~n40558 ;
  assign y30857 = ~1'b0 ;
  assign y30858 = ~n40559 ;
  assign y30859 = n27497 ;
  assign y30860 = ~n40560 ;
  assign y30861 = 1'b0 ;
  assign y30862 = ~1'b0 ;
  assign y30863 = ~n40562 ;
  assign y30864 = ~n40564 ;
  assign y30865 = ~n29296 ;
  assign y30866 = ~1'b0 ;
  assign y30867 = ~n40570 ;
  assign y30868 = n40572 ;
  assign y30869 = ~n40574 ;
  assign y30870 = n26020 ;
  assign y30871 = n40575 ;
  assign y30872 = 1'b0 ;
  assign y30873 = n40576 ;
  assign y30874 = ~n40577 ;
  assign y30875 = n8459 ;
  assign y30876 = n40578 ;
  assign y30877 = ~1'b0 ;
  assign y30878 = ~n40581 ;
  assign y30879 = 1'b0 ;
  assign y30880 = ~n40583 ;
  assign y30881 = ~n840 ;
  assign y30882 = n40585 ;
  assign y30883 = ~1'b0 ;
  assign y30884 = ~n40586 ;
  assign y30885 = ~1'b0 ;
  assign y30886 = n40587 ;
  assign y30887 = 1'b0 ;
  assign y30888 = ~1'b0 ;
  assign y30889 = 1'b0 ;
  assign y30890 = ~n40588 ;
  assign y30891 = ~1'b0 ;
  assign y30892 = ~1'b0 ;
  assign y30893 = ~1'b0 ;
  assign y30894 = ~n40590 ;
  assign y30895 = ~1'b0 ;
  assign y30896 = ~1'b0 ;
  assign y30897 = ~1'b0 ;
  assign y30898 = ~1'b0 ;
  assign y30899 = n40591 ;
  assign y30900 = ~1'b0 ;
  assign y30901 = ~1'b0 ;
  assign y30902 = ~n40592 ;
  assign y30903 = ~n40594 ;
  assign y30904 = ~1'b0 ;
  assign y30905 = ~1'b0 ;
  assign y30906 = ~1'b0 ;
  assign y30907 = ~1'b0 ;
  assign y30908 = ~n1932 ;
  assign y30909 = ~n6892 ;
  assign y30910 = ~n40595 ;
  assign y30911 = ~n40596 ;
  assign y30912 = ~n40597 ;
  assign y30913 = ~1'b0 ;
  assign y30914 = ~n40599 ;
  assign y30915 = ~1'b0 ;
  assign y30916 = ~1'b0 ;
  assign y30917 = ~1'b0 ;
  assign y30918 = n7970 ;
  assign y30919 = ~1'b0 ;
  assign y30920 = n40601 ;
  assign y30921 = ~n40603 ;
  assign y30922 = ~1'b0 ;
  assign y30923 = n40605 ;
  assign y30924 = ~n40607 ;
  assign y30925 = ~n40609 ;
  assign y30926 = n40610 ;
  assign y30927 = ~n40617 ;
  assign y30928 = n40618 ;
  assign y30929 = ~1'b0 ;
  assign y30930 = n40619 ;
  assign y30931 = n40620 ;
  assign y30932 = n40623 ;
  assign y30933 = ~n40624 ;
  assign y30934 = n40625 ;
  assign y30935 = ~1'b0 ;
  assign y30936 = ~1'b0 ;
  assign y30937 = ~1'b0 ;
  assign y30938 = ~n40626 ;
  assign y30939 = 1'b0 ;
  assign y30940 = ~n40627 ;
  assign y30941 = ~n40628 ;
  assign y30942 = ~1'b0 ;
  assign y30943 = n40629 ;
  assign y30944 = n9306 ;
  assign y30945 = ~n4389 ;
  assign y30946 = ~1'b0 ;
  assign y30947 = ~1'b0 ;
  assign y30948 = ~1'b0 ;
  assign y30949 = n40631 ;
  assign y30950 = 1'b0 ;
  assign y30951 = n40633 ;
  assign y30952 = n40634 ;
  assign y30953 = n40636 ;
  assign y30954 = ~n40638 ;
  assign y30955 = ~n1693 ;
  assign y30956 = n40639 ;
  assign y30957 = ~1'b0 ;
  assign y30958 = 1'b0 ;
  assign y30959 = ~n40640 ;
  assign y30960 = n18375 ;
  assign y30961 = ~1'b0 ;
  assign y30962 = n40641 ;
  assign y30963 = n11000 ;
  assign y30964 = ~1'b0 ;
  assign y30965 = ~1'b0 ;
  assign y30966 = ~1'b0 ;
  assign y30967 = n40642 ;
  assign y30968 = ~n40645 ;
  assign y30969 = ~n40647 ;
  assign y30970 = ~1'b0 ;
  assign y30971 = ~n40648 ;
  assign y30972 = ~n40650 ;
  assign y30973 = n40652 ;
  assign y30974 = ~n40655 ;
  assign y30975 = n40658 ;
  assign y30976 = ~n40659 ;
  assign y30977 = ~n40660 ;
  assign y30978 = n592 ;
  assign y30979 = ~n19138 ;
  assign y30980 = ~n40661 ;
  assign y30981 = ~n40662 ;
  assign y30982 = ~1'b0 ;
  assign y30983 = ~1'b0 ;
  assign y30984 = n40663 ;
  assign y30985 = n40664 ;
  assign y30986 = n40667 ;
  assign y30987 = n23066 ;
  assign y30988 = ~1'b0 ;
  assign y30989 = ~n40671 ;
  assign y30990 = ~1'b0 ;
  assign y30991 = n40674 ;
  assign y30992 = n40675 ;
  assign y30993 = ~1'b0 ;
  assign y30994 = n40676 ;
  assign y30995 = ~1'b0 ;
  assign y30996 = ~1'b0 ;
  assign y30997 = n40677 ;
  assign y30998 = n40678 ;
  assign y30999 = ~1'b0 ;
  assign y31000 = n40679 ;
  assign y31001 = ~n40681 ;
  assign y31002 = 1'b0 ;
  assign y31003 = n1043 ;
  assign y31004 = ~n40682 ;
  assign y31005 = ~n1873 ;
  assign y31006 = n40683 ;
  assign y31007 = ~n40685 ;
  assign y31008 = ~1'b0 ;
  assign y31009 = ~1'b0 ;
  assign y31010 = ~1'b0 ;
  assign y31011 = n30938 ;
  assign y31012 = ~1'b0 ;
  assign y31013 = n40688 ;
  assign y31014 = ~1'b0 ;
  assign y31015 = ~1'b0 ;
  assign y31016 = ~1'b0 ;
  assign y31017 = n40689 ;
  assign y31018 = ~1'b0 ;
  assign y31019 = 1'b0 ;
  assign y31020 = ~n12906 ;
  assign y31021 = ~1'b0 ;
  assign y31022 = n6091 ;
  assign y31023 = ~n40692 ;
  assign y31024 = ~n40693 ;
  assign y31025 = n12789 ;
  assign y31026 = ~1'b0 ;
  assign y31027 = ~1'b0 ;
  assign y31028 = ~n40695 ;
  assign y31029 = ~1'b0 ;
  assign y31030 = n22707 ;
  assign y31031 = n40696 ;
  assign y31032 = n40697 ;
  assign y31033 = n40698 ;
  assign y31034 = n40699 ;
  assign y31035 = n40700 ;
  assign y31036 = n6383 ;
  assign y31037 = ~1'b0 ;
  assign y31038 = n40704 ;
  assign y31039 = ~n30999 ;
  assign y31040 = n40707 ;
  assign y31041 = ~1'b0 ;
  assign y31042 = n40710 ;
  assign y31043 = n40712 ;
  assign y31044 = ~n40714 ;
  assign y31045 = n40715 ;
  assign y31046 = n40716 ;
  assign y31047 = ~1'b0 ;
  assign y31048 = ~n40720 ;
  assign y31049 = ~1'b0 ;
  assign y31050 = n40723 ;
  assign y31051 = ~1'b0 ;
  assign y31052 = 1'b0 ;
  assign y31053 = ~n40724 ;
  assign y31054 = ~1'b0 ;
  assign y31055 = n5813 ;
  assign y31056 = 1'b0 ;
  assign y31057 = n40725 ;
  assign y31058 = ~n40726 ;
  assign y31059 = n40729 ;
  assign y31060 = ~n40730 ;
  assign y31061 = ~n40733 ;
  assign y31062 = ~1'b0 ;
  assign y31063 = n12912 ;
  assign y31064 = n40734 ;
  assign y31065 = ~1'b0 ;
  assign y31066 = ~1'b0 ;
  assign y31067 = ~1'b0 ;
  assign y31068 = ~n40735 ;
  assign y31069 = ~n40739 ;
  assign y31070 = n15783 ;
  assign y31071 = n19062 ;
  assign y31072 = ~1'b0 ;
  assign y31073 = ~n40740 ;
  assign y31074 = ~1'b0 ;
  assign y31075 = n40741 ;
  assign y31076 = 1'b0 ;
  assign y31077 = ~1'b0 ;
  assign y31078 = ~n40743 ;
  assign y31079 = n40744 ;
  assign y31080 = ~n40746 ;
  assign y31081 = n6371 ;
  assign y31082 = ~1'b0 ;
  assign y31083 = n40748 ;
  assign y31084 = ~1'b0 ;
  assign y31085 = n40749 ;
  assign y31086 = ~1'b0 ;
  assign y31087 = ~1'b0 ;
  assign y31088 = ~n40753 ;
  assign y31089 = ~n40754 ;
  assign y31090 = n40757 ;
  assign y31091 = ~1'b0 ;
  assign y31092 = ~1'b0 ;
  assign y31093 = ~1'b0 ;
  assign y31094 = 1'b0 ;
  assign y31095 = n40759 ;
  assign y31096 = n40761 ;
  assign y31097 = ~n40763 ;
  assign y31098 = ~1'b0 ;
  assign y31099 = n40765 ;
  assign y31100 = n40766 ;
  assign y31101 = ~1'b0 ;
  assign y31102 = n40768 ;
  assign y31103 = ~1'b0 ;
  assign y31104 = ~1'b0 ;
  assign y31105 = ~1'b0 ;
  assign y31106 = ~1'b0 ;
  assign y31107 = ~1'b0 ;
  assign y31108 = ~1'b0 ;
  assign y31109 = n6695 ;
  assign y31110 = ~1'b0 ;
  assign y31111 = ~n2491 ;
  assign y31112 = ~1'b0 ;
  assign y31113 = ~1'b0 ;
  assign y31114 = n6014 ;
  assign y31115 = ~1'b0 ;
  assign y31116 = ~n8692 ;
  assign y31117 = ~n40770 ;
  assign y31118 = ~n40771 ;
  assign y31119 = n40776 ;
  assign y31120 = ~n40782 ;
  assign y31121 = ~1'b0 ;
  assign y31122 = n40783 ;
  assign y31123 = ~1'b0 ;
  assign y31124 = n40785 ;
  assign y31125 = 1'b0 ;
  assign y31126 = 1'b0 ;
  assign y31127 = ~n40786 ;
  assign y31128 = 1'b0 ;
  assign y31129 = ~n40788 ;
  assign y31130 = 1'b0 ;
  assign y31131 = ~n40789 ;
  assign y31132 = 1'b0 ;
  assign y31133 = n24598 ;
  assign y31134 = ~1'b0 ;
  assign y31135 = n40791 ;
  assign y31136 = ~1'b0 ;
  assign y31137 = ~n40792 ;
  assign y31138 = ~1'b0 ;
  assign y31139 = ~n30469 ;
  assign y31140 = 1'b0 ;
  assign y31141 = ~1'b0 ;
  assign y31142 = ~1'b0 ;
  assign y31143 = ~1'b0 ;
  assign y31144 = ~n40793 ;
  assign y31145 = n40795 ;
  assign y31146 = n40796 ;
  assign y31147 = ~1'b0 ;
  assign y31148 = ~n40799 ;
  assign y31149 = n9270 ;
  assign y31150 = ~1'b0 ;
  assign y31151 = ~n40800 ;
  assign y31152 = ~n40802 ;
  assign y31153 = ~1'b0 ;
  assign y31154 = n40805 ;
  assign y31155 = n2734 ;
  assign y31156 = ~1'b0 ;
  assign y31157 = ~1'b0 ;
  assign y31158 = ~1'b0 ;
  assign y31159 = ~n40808 ;
  assign y31160 = n40810 ;
  assign y31161 = n40814 ;
  assign y31162 = ~1'b0 ;
  assign y31163 = 1'b0 ;
  assign y31164 = n40818 ;
  assign y31165 = n40819 ;
  assign y31166 = ~1'b0 ;
  assign y31167 = ~n40820 ;
  assign y31168 = ~n13183 ;
  assign y31169 = ~n40822 ;
  assign y31170 = ~n40823 ;
  assign y31171 = 1'b0 ;
  assign y31172 = ~n40824 ;
  assign y31173 = 1'b0 ;
  assign y31174 = n20676 ;
  assign y31175 = ~1'b0 ;
  assign y31176 = ~n40825 ;
  assign y31177 = ~n40826 ;
  assign y31178 = ~1'b0 ;
  assign y31179 = ~1'b0 ;
  assign y31180 = ~1'b0 ;
  assign y31181 = ~n40830 ;
  assign y31182 = ~1'b0 ;
  assign y31183 = ~n40831 ;
  assign y31184 = n27061 ;
  assign y31185 = ~1'b0 ;
  assign y31186 = ~1'b0 ;
  assign y31187 = n19841 ;
  assign y31188 = ~1'b0 ;
  assign y31189 = ~n40832 ;
  assign y31190 = ~1'b0 ;
  assign y31191 = ~n40834 ;
  assign y31192 = ~n40837 ;
  assign y31193 = n40838 ;
  assign y31194 = n6077 ;
  assign y31195 = ~1'b0 ;
  assign y31196 = ~n40842 ;
  assign y31197 = ~1'b0 ;
  assign y31198 = n40844 ;
  assign y31199 = n40845 ;
  assign y31200 = ~n4270 ;
  assign y31201 = 1'b0 ;
  assign y31202 = ~1'b0 ;
  assign y31203 = ~n40847 ;
  assign y31204 = ~n40850 ;
  assign y31205 = ~n40855 ;
  assign y31206 = 1'b0 ;
  assign y31207 = n40856 ;
  assign y31208 = ~n40857 ;
  assign y31209 = ~n40858 ;
  assign y31210 = ~1'b0 ;
  assign y31211 = n40860 ;
  assign y31212 = ~n40862 ;
  assign y31213 = n13382 ;
  assign y31214 = n40865 ;
  assign y31215 = ~1'b0 ;
  assign y31216 = ~n40868 ;
  assign y31217 = n40869 ;
  assign y31218 = ~1'b0 ;
  assign y31219 = ~n40870 ;
  assign y31220 = ~1'b0 ;
  assign y31221 = ~n23814 ;
  assign y31222 = ~n40874 ;
  assign y31223 = ~1'b0 ;
  assign y31224 = ~n40876 ;
  assign y31225 = ~1'b0 ;
  assign y31226 = ~1'b0 ;
  assign y31227 = ~n40737 ;
  assign y31228 = n40879 ;
  assign y31229 = n23501 ;
  assign y31230 = n40881 ;
  assign y31231 = ~n40882 ;
  assign y31232 = n40884 ;
  assign y31233 = ~n40886 ;
  assign y31234 = ~1'b0 ;
  assign y31235 = ~n40887 ;
  assign y31236 = n14877 ;
  assign y31237 = n40889 ;
  assign y31238 = ~1'b0 ;
  assign y31239 = n40892 ;
  assign y31240 = ~n40894 ;
  assign y31241 = ~1'b0 ;
  assign y31242 = n40895 ;
  assign y31243 = ~n40896 ;
  assign y31244 = ~n40897 ;
  assign y31245 = ~n6458 ;
  assign y31246 = ~1'b0 ;
  assign y31247 = ~1'b0 ;
  assign y31248 = ~n40900 ;
  assign y31249 = n40901 ;
  assign y31250 = ~n29080 ;
  assign y31251 = n40902 ;
  assign y31252 = ~1'b0 ;
  assign y31253 = ~n9422 ;
  assign y31254 = n40903 ;
  assign y31255 = ~1'b0 ;
  assign y31256 = n40904 ;
  assign y31257 = n40906 ;
  assign y31258 = 1'b0 ;
  assign y31259 = n40907 ;
  assign y31260 = n40909 ;
  assign y31261 = n40912 ;
  assign y31262 = ~1'b0 ;
  assign y31263 = n23690 ;
  assign y31264 = ~n40913 ;
  assign y31265 = ~1'b0 ;
  assign y31266 = ~n40916 ;
  assign y31267 = ~1'b0 ;
  assign y31268 = 1'b0 ;
  assign y31269 = ~n40920 ;
  assign y31270 = ~n440 ;
  assign y31271 = n40922 ;
  assign y31272 = ~n13841 ;
  assign y31273 = ~n40926 ;
  assign y31274 = ~n40930 ;
  assign y31275 = ~n25192 ;
  assign y31276 = 1'b0 ;
  assign y31277 = ~1'b0 ;
  assign y31278 = ~1'b0 ;
  assign y31279 = ~n40932 ;
  assign y31280 = n40933 ;
  assign y31281 = ~1'b0 ;
  assign y31282 = n40949 ;
  assign y31283 = ~n40950 ;
  assign y31284 = ~1'b0 ;
  assign y31285 = ~1'b0 ;
  assign y31286 = n40952 ;
  assign y31287 = ~n40955 ;
  assign y31288 = ~1'b0 ;
  assign y31289 = ~n1283 ;
  assign y31290 = 1'b0 ;
  assign y31291 = ~n40957 ;
  assign y31292 = n40958 ;
  assign y31293 = n40961 ;
  assign y31294 = n40963 ;
  assign y31295 = ~1'b0 ;
  assign y31296 = ~n12883 ;
  assign y31297 = ~n40964 ;
  assign y31298 = ~1'b0 ;
  assign y31299 = ~1'b0 ;
  assign y31300 = ~1'b0 ;
  assign y31301 = 1'b0 ;
  assign y31302 = ~1'b0 ;
  assign y31303 = ~n15196 ;
  assign y31304 = ~1'b0 ;
  assign y31305 = n40967 ;
  assign y31306 = ~n28011 ;
  assign y31307 = ~n40971 ;
  assign y31308 = ~1'b0 ;
  assign y31309 = ~n7668 ;
  assign y31310 = ~1'b0 ;
  assign y31311 = n40973 ;
  assign y31312 = n40975 ;
  assign y31313 = ~1'b0 ;
  assign y31314 = n40979 ;
  assign y31315 = ~1'b0 ;
  assign y31316 = ~1'b0 ;
  assign y31317 = 1'b0 ;
  assign y31318 = n40980 ;
  assign y31319 = n29066 ;
  assign y31320 = ~1'b0 ;
  assign y31321 = ~1'b0 ;
  assign y31322 = ~n40985 ;
  assign y31323 = ~1'b0 ;
  assign y31324 = ~n40986 ;
  assign y31325 = ~1'b0 ;
  assign y31326 = ~1'b0 ;
  assign y31327 = n40996 ;
  assign y31328 = n40998 ;
  assign y31329 = ~n40999 ;
  assign y31330 = n41001 ;
  assign y31331 = ~n41002 ;
  assign y31332 = ~n41005 ;
  assign y31333 = n41007 ;
  assign y31334 = ~1'b0 ;
  assign y31335 = ~1'b0 ;
  assign y31336 = ~1'b0 ;
  assign y31337 = n3791 ;
  assign y31338 = ~1'b0 ;
  assign y31339 = n41008 ;
  assign y31340 = ~n5284 ;
  assign y31341 = ~1'b0 ;
  assign y31342 = ~1'b0 ;
  assign y31343 = n18227 ;
  assign y31344 = ~1'b0 ;
  assign y31345 = ~1'b0 ;
  assign y31346 = n33697 ;
  assign y31347 = n41009 ;
  assign y31348 = ~1'b0 ;
  assign y31349 = 1'b0 ;
  assign y31350 = ~n41011 ;
  assign y31351 = ~n41014 ;
  assign y31352 = n41016 ;
  assign y31353 = ~1'b0 ;
  assign y31354 = ~1'b0 ;
  assign y31355 = ~n31709 ;
  assign y31356 = ~n41019 ;
  assign y31357 = ~1'b0 ;
  assign y31358 = ~1'b0 ;
  assign y31359 = n20590 ;
  assign y31360 = ~n41024 ;
  assign y31361 = n9578 ;
  assign y31362 = ~n41025 ;
  assign y31363 = n41026 ;
  assign y31364 = ~1'b0 ;
  assign y31365 = ~1'b0 ;
  assign y31366 = ~n41028 ;
  assign y31367 = n41031 ;
  assign y31368 = ~1'b0 ;
  assign y31369 = ~n41032 ;
  assign y31370 = ~1'b0 ;
  assign y31371 = n41036 ;
  assign y31372 = n5046 ;
  assign y31373 = ~n30107 ;
  assign y31374 = ~n41038 ;
  assign y31375 = n41041 ;
  assign y31376 = n41044 ;
  assign y31377 = ~1'b0 ;
  assign y31378 = ~n31498 ;
  assign y31379 = 1'b0 ;
  assign y31380 = ~n41045 ;
  assign y31381 = ~n41050 ;
  assign y31382 = n41053 ;
  assign y31383 = ~1'b0 ;
  assign y31384 = ~n41054 ;
  assign y31385 = 1'b0 ;
  assign y31386 = n41055 ;
  assign y31387 = ~n41056 ;
  assign y31388 = ~1'b0 ;
  assign y31389 = ~1'b0 ;
  assign y31390 = ~1'b0 ;
  assign y31391 = ~1'b0 ;
  assign y31392 = n41058 ;
  assign y31393 = ~1'b0 ;
  assign y31394 = ~n23253 ;
  assign y31395 = n41060 ;
  assign y31396 = ~1'b0 ;
  assign y31397 = ~1'b0 ;
  assign y31398 = n41065 ;
  assign y31399 = ~n41066 ;
  assign y31400 = n10851 ;
  assign y31401 = ~n41067 ;
  assign y31402 = ~1'b0 ;
  assign y31403 = n41069 ;
  assign y31404 = ~1'b0 ;
  assign y31405 = n41071 ;
  assign y31406 = n41072 ;
  assign y31407 = ~n15873 ;
  assign y31408 = n41075 ;
  assign y31409 = ~n41082 ;
  assign y31410 = n41084 ;
  assign y31411 = n41086 ;
  assign y31412 = ~1'b0 ;
  assign y31413 = ~1'b0 ;
  assign y31414 = ~1'b0 ;
  assign y31415 = n41087 ;
  assign y31416 = ~1'b0 ;
  assign y31417 = ~n41088 ;
  assign y31418 = ~n41089 ;
  assign y31419 = ~1'b0 ;
  assign y31420 = ~1'b0 ;
  assign y31421 = ~n41093 ;
  assign y31422 = ~1'b0 ;
  assign y31423 = n41095 ;
  assign y31424 = ~n41097 ;
  assign y31425 = ~1'b0 ;
  assign y31426 = n41099 ;
  assign y31427 = 1'b0 ;
  assign y31428 = ~n34487 ;
  assign y31429 = ~n41100 ;
  assign y31430 = ~1'b0 ;
  assign y31431 = ~n41102 ;
  assign y31432 = n41106 ;
  assign y31433 = ~1'b0 ;
  assign y31434 = ~n41110 ;
  assign y31435 = ~n41111 ;
  assign y31436 = ~1'b0 ;
  assign y31437 = ~1'b0 ;
  assign y31438 = n10729 ;
  assign y31439 = n41116 ;
  assign y31440 = n41117 ;
  assign y31441 = ~1'b0 ;
  assign y31442 = ~1'b0 ;
  assign y31443 = ~1'b0 ;
  assign y31444 = 1'b0 ;
  assign y31445 = n41119 ;
  assign y31446 = ~n39698 ;
  assign y31447 = n41120 ;
  assign y31448 = ~1'b0 ;
  assign y31449 = n11766 ;
  assign y31450 = n41121 ;
  assign y31451 = ~1'b0 ;
  assign y31452 = ~n22924 ;
  assign y31453 = ~1'b0 ;
  assign y31454 = n41124 ;
  assign y31455 = ~1'b0 ;
  assign y31456 = ~1'b0 ;
  assign y31457 = ~1'b0 ;
  assign y31458 = ~1'b0 ;
  assign y31459 = n41126 ;
  assign y31460 = ~n41128 ;
  assign y31461 = ~n41129 ;
  assign y31462 = n41134 ;
  assign y31463 = ~n41139 ;
  assign y31464 = n41140 ;
  assign y31465 = n41141 ;
  assign y31466 = ~1'b0 ;
  assign y31467 = ~1'b0 ;
  assign y31468 = ~n41144 ;
  assign y31469 = ~1'b0 ;
  assign y31470 = ~n41154 ;
  assign y31471 = n41155 ;
  assign y31472 = ~n33057 ;
  assign y31473 = ~n41158 ;
  assign y31474 = ~1'b0 ;
  assign y31475 = ~1'b0 ;
  assign y31476 = ~n41160 ;
  assign y31477 = n41161 ;
  assign y31478 = ~n41163 ;
  assign y31479 = ~n28253 ;
  assign y31480 = ~1'b0 ;
  assign y31481 = ~1'b0 ;
  assign y31482 = ~1'b0 ;
  assign y31483 = ~n41165 ;
  assign y31484 = ~1'b0 ;
  assign y31485 = ~1'b0 ;
  assign y31486 = ~n616 ;
  assign y31487 = ~n41167 ;
  assign y31488 = n41168 ;
  assign y31489 = ~1'b0 ;
  assign y31490 = ~n41169 ;
  assign y31491 = ~1'b0 ;
  assign y31492 = ~n4436 ;
  assign y31493 = ~n41170 ;
  assign y31494 = n41171 ;
  assign y31495 = ~1'b0 ;
  assign y31496 = ~1'b0 ;
  assign y31497 = ~n41173 ;
  assign y31498 = n41174 ;
  assign y31499 = ~n41176 ;
  assign y31500 = ~1'b0 ;
  assign y31501 = ~1'b0 ;
  assign y31502 = n41178 ;
  assign y31503 = 1'b0 ;
  assign y31504 = ~n41179 ;
  assign y31505 = ~n41181 ;
  assign y31506 = n41189 ;
  assign y31507 = ~1'b0 ;
  assign y31508 = ~1'b0 ;
  assign y31509 = ~n41191 ;
  assign y31510 = 1'b0 ;
  assign y31511 = ~1'b0 ;
  assign y31512 = n41194 ;
  assign y31513 = n41196 ;
  assign y31514 = ~1'b0 ;
  assign y31515 = 1'b0 ;
  assign y31516 = n41197 ;
  assign y31517 = ~n41199 ;
  assign y31518 = ~1'b0 ;
  assign y31519 = n41203 ;
  assign y31520 = n3326 ;
  assign y31521 = ~1'b0 ;
  assign y31522 = n41206 ;
  assign y31523 = ~1'b0 ;
  assign y31524 = ~1'b0 ;
  assign y31525 = ~n41210 ;
  assign y31526 = n1316 ;
  assign y31527 = ~n41212 ;
  assign y31528 = ~1'b0 ;
  assign y31529 = ~1'b0 ;
  assign y31530 = ~1'b0 ;
  assign y31531 = ~1'b0 ;
  assign y31532 = ~1'b0 ;
  assign y31533 = ~1'b0 ;
  assign y31534 = n41213 ;
  assign y31535 = ~1'b0 ;
  assign y31536 = ~n41218 ;
  assign y31537 = 1'b0 ;
  assign y31538 = ~n8750 ;
  assign y31539 = ~1'b0 ;
  assign y31540 = ~n41219 ;
  assign y31541 = ~1'b0 ;
  assign y31542 = ~1'b0 ;
  assign y31543 = ~n41221 ;
  assign y31544 = ~n41222 ;
  assign y31545 = n41223 ;
  assign y31546 = ~n34642 ;
  assign y31547 = ~1'b0 ;
  assign y31548 = n41224 ;
  assign y31549 = ~n41226 ;
  assign y31550 = ~n41227 ;
  assign y31551 = ~1'b0 ;
  assign y31552 = ~1'b0 ;
  assign y31553 = n41232 ;
  assign y31554 = ~1'b0 ;
  assign y31555 = n41238 ;
  assign y31556 = ~n41240 ;
  assign y31557 = n41241 ;
  assign y31558 = ~1'b0 ;
  assign y31559 = ~n18923 ;
  assign y31560 = n41242 ;
  assign y31561 = ~n41244 ;
  assign y31562 = n33517 ;
  assign y31563 = n41245 ;
  assign y31564 = n41249 ;
  assign y31565 = n41252 ;
  assign y31566 = ~1'b0 ;
  assign y31567 = ~n41253 ;
  assign y31568 = ~n8084 ;
  assign y31569 = ~n41254 ;
  assign y31570 = ~1'b0 ;
  assign y31571 = n41255 ;
  assign y31572 = ~n41256 ;
  assign y31573 = ~n41260 ;
  assign y31574 = ~1'b0 ;
  assign y31575 = ~1'b0 ;
  assign y31576 = n41261 ;
  assign y31577 = n41262 ;
  assign y31578 = n41263 ;
  assign y31579 = ~n41265 ;
  assign y31580 = ~n41266 ;
  assign y31581 = ~1'b0 ;
  assign y31582 = n41271 ;
  assign y31583 = ~1'b0 ;
  assign y31584 = ~1'b0 ;
  assign y31585 = n41273 ;
  assign y31586 = ~1'b0 ;
  assign y31587 = n28764 ;
  assign y31588 = ~n41274 ;
  assign y31589 = ~n41276 ;
  assign y31590 = 1'b0 ;
  assign y31591 = ~1'b0 ;
  assign y31592 = n41277 ;
  assign y31593 = n41279 ;
  assign y31594 = n41284 ;
  assign y31595 = ~n10664 ;
  assign y31596 = ~1'b0 ;
  assign y31597 = ~n41288 ;
  assign y31598 = ~1'b0 ;
  assign y31599 = ~1'b0 ;
  assign y31600 = n41289 ;
  assign y31601 = ~1'b0 ;
  assign y31602 = ~1'b0 ;
  assign y31603 = ~1'b0 ;
  assign y31604 = n41291 ;
  assign y31605 = n24313 ;
  assign y31606 = n41292 ;
  assign y31607 = ~1'b0 ;
  assign y31608 = ~n41293 ;
  assign y31609 = ~1'b0 ;
  assign y31610 = ~1'b0 ;
  assign y31611 = n1140 ;
  assign y31612 = n41295 ;
  assign y31613 = ~1'b0 ;
  assign y31614 = n30 ;
  assign y31615 = 1'b0 ;
  assign y31616 = ~n13478 ;
  assign y31617 = ~1'b0 ;
  assign y31618 = ~1'b0 ;
  assign y31619 = ~n41297 ;
  assign y31620 = ~n41301 ;
  assign y31621 = n41305 ;
  assign y31622 = n41306 ;
  assign y31623 = ~1'b0 ;
  assign y31624 = n41308 ;
  assign y31625 = ~n41298 ;
  assign y31626 = n41309 ;
  assign y31627 = ~n41311 ;
  assign y31628 = ~n41315 ;
  assign y31629 = ~1'b0 ;
  assign y31630 = ~1'b0 ;
  assign y31631 = ~n41320 ;
  assign y31632 = n2882 ;
  assign y31633 = n41322 ;
  assign y31634 = n13715 ;
  assign y31635 = ~1'b0 ;
  assign y31636 = n41323 ;
  assign y31637 = ~1'b0 ;
  assign y31638 = ~1'b0 ;
  assign y31639 = ~n41324 ;
  assign y31640 = ~n41326 ;
  assign y31641 = ~1'b0 ;
  assign y31642 = ~1'b0 ;
  assign y31643 = 1'b0 ;
  assign y31644 = n41327 ;
  assign y31645 = ~n41331 ;
  assign y31646 = ~n41333 ;
  assign y31647 = ~n41335 ;
  assign y31648 = ~n41336 ;
  assign y31649 = ~1'b0 ;
  assign y31650 = ~n41338 ;
  assign y31651 = ~n41344 ;
  assign y31652 = ~n41345 ;
  assign y31653 = ~1'b0 ;
  assign y31654 = 1'b0 ;
  assign y31655 = ~n41347 ;
  assign y31656 = ~1'b0 ;
  assign y31657 = ~n41349 ;
  assign y31658 = ~n41351 ;
  assign y31659 = ~1'b0 ;
  assign y31660 = ~1'b0 ;
  assign y31661 = ~1'b0 ;
  assign y31662 = ~1'b0 ;
  assign y31663 = ~1'b0 ;
  assign y31664 = n31800 ;
  assign y31665 = n41353 ;
  assign y31666 = n41354 ;
  assign y31667 = n41358 ;
  assign y31668 = ~n41360 ;
  assign y31669 = ~n41366 ;
  assign y31670 = ~1'b0 ;
  assign y31671 = ~1'b0 ;
  assign y31672 = ~1'b0 ;
  assign y31673 = 1'b0 ;
  assign y31674 = ~n34939 ;
  assign y31675 = n41368 ;
  assign y31676 = ~n10403 ;
  assign y31677 = n41369 ;
  assign y31678 = ~n41372 ;
  assign y31679 = n41373 ;
  assign y31680 = ~n41377 ;
  assign y31681 = ~n18505 ;
  assign y31682 = ~1'b0 ;
  assign y31683 = ~1'b0 ;
  assign y31684 = ~1'b0 ;
  assign y31685 = n41378 ;
  assign y31686 = ~1'b0 ;
  assign y31687 = n41381 ;
  assign y31688 = ~n41383 ;
  assign y31689 = ~n41385 ;
  assign y31690 = ~n8208 ;
  assign y31691 = ~1'b0 ;
  assign y31692 = ~n41388 ;
  assign y31693 = ~n41390 ;
  assign y31694 = ~1'b0 ;
  assign y31695 = 1'b0 ;
  assign y31696 = n41391 ;
  assign y31697 = ~n41394 ;
  assign y31698 = ~1'b0 ;
  assign y31699 = ~n41397 ;
  assign y31700 = n41398 ;
  assign y31701 = 1'b0 ;
  assign y31702 = ~n41407 ;
  assign y31703 = ~n7395 ;
  assign y31704 = ~1'b0 ;
  assign y31705 = ~n41408 ;
  assign y31706 = ~n41410 ;
  assign y31707 = ~n41414 ;
  assign y31708 = n3382 ;
  assign y31709 = ~n5101 ;
  assign y31710 = ~1'b0 ;
  assign y31711 = ~1'b0 ;
  assign y31712 = ~n41416 ;
  assign y31713 = ~n11827 ;
  assign y31714 = ~n41417 ;
  assign y31715 = n1048 ;
  assign y31716 = ~1'b0 ;
  assign y31717 = ~1'b0 ;
  assign y31718 = ~1'b0 ;
  assign y31719 = ~n2876 ;
  assign y31720 = ~n41420 ;
  assign y31721 = n41421 ;
  assign y31722 = ~1'b0 ;
  assign y31723 = n41427 ;
  assign y31724 = ~n41429 ;
  assign y31725 = n41430 ;
  assign y31726 = ~1'b0 ;
  assign y31727 = ~1'b0 ;
  assign y31728 = ~1'b0 ;
  assign y31729 = n41432 ;
  assign y31730 = ~n41433 ;
  assign y31731 = ~1'b0 ;
  assign y31732 = n41434 ;
  assign y31733 = ~n41437 ;
  assign y31734 = n41438 ;
  assign y31735 = n41441 ;
  assign y31736 = n41442 ;
  assign y31737 = 1'b0 ;
  assign y31738 = ~1'b0 ;
  assign y31739 = ~n41450 ;
  assign y31740 = ~1'b0 ;
  assign y31741 = ~1'b0 ;
  assign y31742 = ~1'b0 ;
  assign y31743 = ~1'b0 ;
  assign y31744 = ~1'b0 ;
  assign y31745 = ~n41452 ;
  assign y31746 = ~n29790 ;
  assign y31747 = ~1'b0 ;
  assign y31748 = n41453 ;
  assign y31749 = ~n41459 ;
  assign y31750 = ~n41462 ;
  assign y31751 = ~n41465 ;
  assign y31752 = n41466 ;
  assign y31753 = ~n41468 ;
  assign y31754 = ~1'b0 ;
  assign y31755 = n41471 ;
  assign y31756 = ~n41475 ;
  assign y31757 = ~n3483 ;
  assign y31758 = n41478 ;
  assign y31759 = ~n41480 ;
  assign y31760 = n41482 ;
  assign y31761 = n41486 ;
  assign y31762 = n41487 ;
  assign y31763 = ~n41490 ;
  assign y31764 = n41492 ;
  assign y31765 = 1'b0 ;
  assign y31766 = ~n41493 ;
  assign y31767 = n41494 ;
  assign y31768 = ~n23402 ;
  assign y31769 = 1'b0 ;
  assign y31770 = n41495 ;
  assign y31771 = ~n41496 ;
  assign y31772 = n7955 ;
  assign y31773 = ~n41499 ;
  assign y31774 = ~1'b0 ;
  assign y31775 = ~1'b0 ;
  assign y31776 = ~n41508 ;
  assign y31777 = n41509 ;
  assign y31778 = ~1'b0 ;
  assign y31779 = ~n8046 ;
  assign y31780 = ~1'b0 ;
  assign y31781 = ~n41512 ;
  assign y31782 = ~1'b0 ;
  assign y31783 = n41513 ;
  assign y31784 = ~1'b0 ;
  assign y31785 = n41514 ;
  assign y31786 = ~1'b0 ;
  assign y31787 = ~1'b0 ;
  assign y31788 = n41515 ;
  assign y31789 = ~1'b0 ;
  assign y31790 = ~1'b0 ;
  assign y31791 = 1'b0 ;
  assign y31792 = ~n41516 ;
  assign y31793 = ~n41517 ;
  assign y31794 = ~1'b0 ;
  assign y31795 = n41518 ;
  assign y31796 = ~n41520 ;
  assign y31797 = n20975 ;
  assign y31798 = ~1'b0 ;
  assign y31799 = ~n41521 ;
  assign y31800 = ~1'b0 ;
  assign y31801 = n41522 ;
  assign y31802 = ~n906 ;
  assign y31803 = ~1'b0 ;
  assign y31804 = ~1'b0 ;
  assign y31805 = ~n41524 ;
  assign y31806 = ~n17391 ;
  assign y31807 = n41525 ;
  assign y31808 = ~n41527 ;
  assign y31809 = ~1'b0 ;
  assign y31810 = n41529 ;
  assign y31811 = ~n36387 ;
  assign y31812 = ~n41534 ;
  assign y31813 = ~1'b0 ;
  assign y31814 = ~1'b0 ;
  assign y31815 = n39975 ;
  assign y31816 = ~1'b0 ;
  assign y31817 = ~n13865 ;
  assign y31818 = n41535 ;
  assign y31819 = ~1'b0 ;
  assign y31820 = n41536 ;
  assign y31821 = n41539 ;
  assign y31822 = n41541 ;
  assign y31823 = 1'b0 ;
  assign y31824 = ~1'b0 ;
  assign y31825 = ~1'b0 ;
  assign y31826 = n41544 ;
  assign y31827 = n41545 ;
  assign y31828 = n41546 ;
  assign y31829 = ~1'b0 ;
  assign y31830 = n41548 ;
  assign y31831 = 1'b0 ;
  assign y31832 = ~n41549 ;
  assign y31833 = n41550 ;
  assign y31834 = ~1'b0 ;
  assign y31835 = n7056 ;
  assign y31836 = ~1'b0 ;
  assign y31837 = ~1'b0 ;
  assign y31838 = ~1'b0 ;
  assign y31839 = ~n41551 ;
  assign y31840 = ~1'b0 ;
  assign y31841 = ~n31679 ;
  assign y31842 = ~n41553 ;
  assign y31843 = ~n41554 ;
  assign y31844 = ~1'b0 ;
  assign y31845 = ~n41556 ;
  assign y31846 = n41557 ;
  assign y31847 = ~n41558 ;
  assign y31848 = ~n19112 ;
  assign y31849 = ~1'b0 ;
  assign y31850 = ~1'b0 ;
  assign y31851 = 1'b0 ;
  assign y31852 = n10548 ;
  assign y31853 = ~n41560 ;
  assign y31854 = n41561 ;
  assign y31855 = ~1'b0 ;
  assign y31856 = ~1'b0 ;
  assign y31857 = ~n8561 ;
  assign y31858 = n41563 ;
  assign y31859 = ~n41566 ;
  assign y31860 = ~1'b0 ;
  assign y31861 = ~1'b0 ;
  assign y31862 = ~n41567 ;
  assign y31863 = ~1'b0 ;
  assign y31864 = ~1'b0 ;
  assign y31865 = n16629 ;
  assign y31866 = ~1'b0 ;
  assign y31867 = ~1'b0 ;
  assign y31868 = ~n41574 ;
  assign y31869 = ~n41576 ;
  assign y31870 = ~n41580 ;
  assign y31871 = ~n41582 ;
  assign y31872 = n41583 ;
  assign y31873 = n41584 ;
  assign y31874 = ~1'b0 ;
  assign y31875 = ~n41585 ;
  assign y31876 = ~n29144 ;
  assign y31877 = n41586 ;
  assign y31878 = ~n41588 ;
  assign y31879 = ~n10784 ;
  assign y31880 = ~1'b0 ;
  assign y31881 = n41590 ;
  assign y31882 = ~1'b0 ;
  assign y31883 = n41593 ;
  assign y31884 = n41594 ;
  assign y31885 = ~1'b0 ;
  assign y31886 = ~1'b0 ;
  assign y31887 = n41597 ;
  assign y31888 = ~1'b0 ;
  assign y31889 = ~n41598 ;
  assign y31890 = n41599 ;
  assign y31891 = ~n41601 ;
  assign y31892 = ~1'b0 ;
  assign y31893 = ~1'b0 ;
  assign y31894 = ~n41603 ;
  assign y31895 = ~1'b0 ;
  assign y31896 = ~1'b0 ;
  assign y31897 = 1'b0 ;
  assign y31898 = n567 ;
  assign y31899 = ~n41604 ;
  assign y31900 = n41606 ;
  assign y31901 = ~n41608 ;
  assign y31902 = n41611 ;
  assign y31903 = ~n41612 ;
  assign y31904 = 1'b0 ;
  assign y31905 = ~n41615 ;
  assign y31906 = ~1'b0 ;
  assign y31907 = 1'b0 ;
  assign y31908 = ~n41617 ;
  assign y31909 = ~n41618 ;
  assign y31910 = n41620 ;
  assign y31911 = n41622 ;
  assign y31912 = n41623 ;
  assign y31913 = 1'b0 ;
  assign y31914 = ~1'b0 ;
  assign y31915 = ~n41624 ;
  assign y31916 = n41626 ;
  assign y31917 = ~n41627 ;
  assign y31918 = n41629 ;
  assign y31919 = ~n41631 ;
  assign y31920 = ~n41635 ;
  assign y31921 = ~1'b0 ;
  assign y31922 = n41636 ;
  assign y31923 = n41639 ;
  assign y31924 = ~1'b0 ;
  assign y31925 = ~n39267 ;
  assign y31926 = ~n41641 ;
  assign y31927 = n41644 ;
  assign y31928 = n41645 ;
  assign y31929 = ~1'b0 ;
  assign y31930 = ~1'b0 ;
  assign y31931 = 1'b0 ;
  assign y31932 = 1'b0 ;
  assign y31933 = ~1'b0 ;
  assign y31934 = ~n41646 ;
  assign y31935 = ~n40225 ;
  assign y31936 = n41647 ;
  assign y31937 = ~1'b0 ;
  assign y31938 = ~n41648 ;
  assign y31939 = n41651 ;
  assign y31940 = n41653 ;
  assign y31941 = n41654 ;
  assign y31942 = ~n41657 ;
  assign y31943 = ~1'b0 ;
  assign y31944 = n19595 ;
  assign y31945 = 1'b0 ;
  assign y31946 = ~n41659 ;
  assign y31947 = ~1'b0 ;
  assign y31948 = n41660 ;
  assign y31949 = n11735 ;
  assign y31950 = 1'b0 ;
  assign y31951 = ~1'b0 ;
  assign y31952 = ~1'b0 ;
  assign y31953 = ~n41662 ;
  assign y31954 = ~1'b0 ;
  assign y31955 = ~1'b0 ;
  assign y31956 = ~n41664 ;
  assign y31957 = n41665 ;
  assign y31958 = 1'b0 ;
  assign y31959 = ~1'b0 ;
  assign y31960 = ~n41666 ;
  assign y31961 = n31329 ;
  assign y31962 = n41671 ;
  assign y31963 = 1'b0 ;
  assign y31964 = n41673 ;
  assign y31965 = ~1'b0 ;
  assign y31966 = ~1'b0 ;
  assign y31967 = ~n41675 ;
  assign y31968 = ~n41677 ;
  assign y31969 = ~n12196 ;
  assign y31970 = ~1'b0 ;
  assign y31971 = 1'b0 ;
  assign y31972 = 1'b0 ;
  assign y31973 = n41679 ;
  assign y31974 = ~n41680 ;
  assign y31975 = ~n41681 ;
  assign y31976 = ~n41682 ;
  assign y31977 = n41691 ;
  assign y31978 = ~n41693 ;
  assign y31979 = ~1'b0 ;
  assign y31980 = ~1'b0 ;
  assign y31981 = ~n41694 ;
  assign y31982 = ~1'b0 ;
  assign y31983 = ~n41697 ;
  assign y31984 = n41699 ;
  assign y31985 = n3399 ;
  assign y31986 = n6610 ;
  assign y31987 = ~1'b0 ;
  assign y31988 = ~1'b0 ;
  assign y31989 = ~1'b0 ;
  assign y31990 = 1'b0 ;
  assign y31991 = ~n34190 ;
  assign y31992 = n41701 ;
  assign y31993 = ~n41703 ;
  assign y31994 = ~1'b0 ;
  assign y31995 = ~1'b0 ;
  assign y31996 = n41705 ;
  assign y31997 = ~n41706 ;
  assign y31998 = n41707 ;
  assign y31999 = n41709 ;
  assign y32000 = ~1'b0 ;
  assign y32001 = ~1'b0 ;
  assign y32002 = n41710 ;
  assign y32003 = 1'b0 ;
  assign y32004 = ~1'b0 ;
  assign y32005 = ~1'b0 ;
  assign y32006 = 1'b0 ;
  assign y32007 = n41713 ;
  assign y32008 = ~n41715 ;
  assign y32009 = n41717 ;
  assign y32010 = ~1'b0 ;
  assign y32011 = ~n40228 ;
  assign y32012 = ~1'b0 ;
  assign y32013 = 1'b0 ;
  assign y32014 = ~1'b0 ;
  assign y32015 = ~n41718 ;
  assign y32016 = 1'b0 ;
  assign y32017 = ~1'b0 ;
  assign y32018 = n41720 ;
  assign y32019 = ~n41722 ;
  assign y32020 = ~n41724 ;
  assign y32021 = 1'b0 ;
  assign y32022 = ~1'b0 ;
  assign y32023 = ~1'b0 ;
  assign y32024 = n41726 ;
  assign y32025 = ~1'b0 ;
  assign y32026 = ~n41732 ;
  assign y32027 = ~n41735 ;
  assign y32028 = 1'b0 ;
  assign y32029 = n5412 ;
  assign y32030 = ~n41741 ;
  assign y32031 = ~n41743 ;
  assign y32032 = ~1'b0 ;
  assign y32033 = ~1'b0 ;
  assign y32034 = 1'b0 ;
endmodule
